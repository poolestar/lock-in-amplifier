`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
R/f6FeJ0QLro/ha58bTY8NKxDKKO+q15gtVmuO+X1HoPKFvrmCJfIKY2+7Y4Wuzatwd/djCDDzbj
Lz/cs4hVvg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lvJVFxu1g3pXdpkq1DD/m9B6mZRZl1z25RnVPa2Pqa1r9owDEtgzfIY4YDwmNQWPtDZsGSa+gEVc
uqLBz0NWoe/TiDsviZj2qMM4pCFiMScHidDdqY7hiOFolMJLOulI7mQ0fiA5T+heXQGYdREM/Qxj
GFB/xJTL+k8zIvuECHc=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
a5PKA7Wq+G9niejwJOtSNs4IYuZHc8JqbN6w2EefAaPj+yqsVOpcNJaAPUuj6cFCMp7VN9w85Z05
FkFSxCcUs7RmQu3uWLGNQezUuGW/d6OS7GYPf4MRX9mK7q0fMkS51Hl+4n0QkyxOcB8Z84+JB4dc
KwKO49DHwZGhr+GGEZQ=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Jcb8JNchDQSiulaqmbTXpOUYbMkdd6d293bW8sxozNV2U0p6APpmuBEA/7+1IWt2cownZDUiOKbh
vpwDhXEdV3JarZHTGsXiIAWpt1Vb8QcOd4sKL7UeP47aQzH/7PSfm+5VaJ53FRa9Re0Yyiy+xiDq
5WVXsB9CYYUn/nWLUbEWGdBizGZnmhwxGfWdJHz5tlSnRgJn1ZXc9UpXaugB8C9Yfndn1hGYi2LE
tSAxdQ3IeR2usZtM/poSve0h0ybGzEZxjlKK0JJwlaNPwKJMIqwSNyeYlhN7d22YGRW4es59Wp2f
gGsqis3PqJ7NiPAfwd+Yjbzi7svUdzwMx+pfWA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JtZntbd26RdNOdSV6FB7P8Axt3WOPCRpCpwgQKzPy2bHyy1xOosVNfEGfOCxVQ1nZWYD5L94l8eL
17GOiNRzQ89J9xdECYcyMVwbwDQV1nQpWX+6FTvcVdecK+hQyFs+2Yn5HH/kbbObpoIJz9gCxUmF
BH71W4+J+zEZKiu9xnknefZOhniAzDyKNKc9y3UI0pUoJmpv4HVR3XBXMkvPo+wnxzA3wtzrZnpl
ABbEwNwHOUX4HT6JHiiyy8C6BQBDHp/2srtR9XQdv04gJ1JjPTHdrdHy/7xZ4ufKW1UJ666d1b2L
SBegWiCzIFgbSKTujiY2Ob2b6lsDW+W+JjzIzQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
U7NH9yg0f8tUSSiMzO2ZV0vdPTPVgwBRvvyiarSitGa0/REvP3ado3WY4HYt7rtUt6whHqYlgSz4
hK41g8yCOnMvqeHIQnhbMDDd1y7QyRgOUBuZB71vrBBw871SocSq9FNklLclETG0J7Khywsw8So0
HUBpgiZ9bVTO8LU+2SabnPD3ChIt7NLLDHs9/z7JnEqXPf7KiCTdIFM8Szq2mSAw2Q6DTv+cYfYJ
HRazXb4a76QvTIBZbtKXyaOLgRURM4WFVAPBZp/T6h91uV2D4iz5NecaV46d2ZFMpc/6K5y/I4l1
GU+vKtfSH1upfbz5itvG/2sn98hh9hrtmMHXNQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 67920)
`protect data_block
9tJTcCtZHraGI/8rPIzcvmKMbEp4F+jGZJSBm3QWbTQ5vrn4RDbw/8Jq5i6aq5ocst7TsGm0Kls1
DlFr2r1Knh1F680aNjq/ohknlxqFDDizmXniQV7obs2+W4BBDY8tCOaE3D4ULW9kk6XrHBsN8h0X
cgtOuKF2LWOkFobMrWe/O98xzbdg70+W77iTyx/+z5uoIofjnaXXrtSY6kZpdUvrsBk0zsnsCscf
Doo9LeVp4vKEtYjoyaBYu77+wE+OJrTCJ/OHpzYsbuhmtMUrKLDAkoKcUPWLPQBZFAmdA/sdnhP2
wM2wAPTKqVYwko/Azxmg0Lt7UMTey8MXxKaLays3QM25sbju1CkYiQl6PiICFcncHWNLOsiS9/2s
MGtursRzYhvi82lzYn1UaLbMuqO17Yr0xdacy6EtjdHqIICX/y4mR8nxKdk3Fv05/r3q20Qi6ENZ
TSbCq1pUmz2fxIb86b3xPOEhyH3HWMX0ayW3eTAmQFgYlwHgNKR9onqge6GjaL07T1FkSS8xKsUn
G2k6qo81jFTChQ//1r5cecyoeIehzB1iyhdez6zWTpDLJD4bBNiB8enikTBH08X2tGWOEvC3+mTv
oRNN3vu5XJY2kfWdLIDu77DP31xuxb66pL+WcjuiC0KtIpcpe39gOW+LdWMMkAo8BW+cCraW1q4Z
5vLZRahSHXSHo9koSPwwj5WP58ffsRqfna/DV+N+LUaodXPrnOj55zx4J698rONLVCMR8t3QXtzR
/b80pUVwp9HCZ6bZT9AE09lP4QCy27RVx/UbHQ0wywm9xGulpq1UC7Tum2KGlMNe3UBgh7JRz/2h
0idOJPiWlrBpAYLlui5iANE59D/ljnEQMnUCQTx47X4gesjI2zmozrNMWLNt+ePYHQGI8DCMDTn/
B5TF5TC0TOlke2wuMcEk7jUTnxjYe1/QHcucQKSwpRYQ3RXvEKXd8yxeP15zzMwjeCuaMTJeCOhQ
YQcJd/ceYOdSKdohkUtrMC4QxkBRE6ayNt6xpU+ld3n1nZ7FaMvYmKVLNyuPz+qMO3yr84DeEkv3
fhZdyKOUGp24ASSFl90Ib+rTv8ot7ksC4x8g36u9Sd6rEKxUD7n8p8uZAzrj/YEwqbWQxKJ1cTPL
Iny9BszuctZ4tgq+7MFVe52IRy9XQDanNe1XrMDcGvNr0Zf4YWYHAVv4qsUqtN4APSqCwIQE/ktk
dhfZ8WAkLR3W+2hN27JWa44E5TYR8JtxYS1DIp4XuFmx79jZaQp3/zE72Kiy6m/Mc+nWCaHgFpDf
QDKrdPDb7qWVHtZtCki+GUXhECujdWKeOPU10IuPhj8aNBo1s6D0QC0ChmWJcPCotZQLutNLMwQJ
MUytl0cifd+D+tpJa/h04ygH2orrvvVx+kS3zM5HckoBE+5nR2bpwdbXRzg+dUYu0J7nffR3tH7w
2lwxmGCpgTQ1ej6g9uFKNQhyswvj9gWsOTTgKetaowJl1licIvL5wPzaKs1z3laZKddeZ74xCLc2
F7e5aOocWoFxJYvKqtVCp5xrbJPZabnaptlzBngSlZS7gBKHu22/dk54KzGZnPYL7Po0BQac+oDz
izxdj9f489cp1dEZ8YWI4qYyV6d3WNeSCnha+89R3MbAKlDM7OyvXexB25xqyRq/RtOGejaO84m/
EYPNPBrt9u4FVVQCblEpX2vOnjmTBCQ+XWMx4AFNEeWn/wUINCvRjTsUmx5OKBfEkxd8DDdANTJg
FQWFskiYhpddSbW1OfxnuiKOFpOAtH7e6eMpgPQj8Ui90B+r+Od2UaeoStscZ9bioDcPv1GiOjA+
8caPra+lVVP8CdaN9YKQyfzNXfQiKBO1g/rpEWEcJ1Wosq2AW/ykBBvIMZ1tAsGluyJ70nySQNV+
joE+Yeqc1lkSq+vecLhGc5I1J/gVcSPFKPR4S5yu38a3wwHx8FOuB/KDtHIsGQAORt2ZgblljRz3
gdyElRihFR0g3aaan1TUW7lFNO7SOGS38skBzw3BJXmGJpDwg6V77Fga2Iq4/0ZNXJhLis9nAkBd
3Pw/yEnszyTk4qb0Z95BGqoD3PJAsx8UN0cV1YsvBBw9pvFhq4ANSVcMY0cifsIX2NKY8qzL6JFD
g14P+bJax57SdikFhV7+4VbJazniMig3x6K4IZ4g3suJg7AG/szKt6NqIhPvgSVNeK9msqyjEwzI
JPUlfw42hdg94TkvO7O9zyG1K6tGBS8c76HN7E/tQy3WGewP+jKCec5fY3FgNfkJMhmMsW1xA2HX
BLxTEqZVBbz+8lTWZFIyv8gZJ3P6ZXweE8atLoV87e1PKWYRrc6w/J3ApmdFjwdZOIjhZwjPIMBL
9ycISJyc0fcGEu9LGnHkgiJEEjSDnpwN/FIdkubDbiCW4unCSpF69UbHVpv685DNveeD7Lw7jCQM
crnDyyM04Kf39VuwZTO7dYIkL6s/NvVFRp4IT6ru8+ZLXGTeltm1euXWNCQSzs2oTLxNjwaxtfrF
0sXjFkT7Y+T8tGBGxAV0Rf40R3w2FgBpYkDB+1ZeS45ZG7RkRzKUtWj+zZFpBtfE1AzWU98QgVzT
7uIAQZG8cxdUDdAwJ2aA/TofG5ARg2cHDjYwDF81CgFMoym4TNFkDnntsDHUyE6f7FCPt/VJ8bf8
toSqEkzU1FWidDuAndU45mWXGbZFaaiPvM3IgnUIgOY585hIUWUfEzIcr3OHw0nhs3KwE9OCIXbC
AhD3se/to5GxZI9YraKQmmcXLapqJABSvWzG7mdpVJ2M//uyNf151fowyx8tf5ZIyx3OP46qNc9L
k/bTEmjLQTpd8x1ukjwnUVcwUiejt5ar5v9yEonfZDgr6iKouCxAkmkKLN2KGlPmz94TIAlRe+uU
J6Cq7w9UMf4ADUEgxv6+x1jKQ93bZ78FyoaYkiARZPMLUBL6TbFwp/HgRs6GGfUPKXUFO1qc8DVw
weRx0mL17+Uk0fw7YrsoW1WlRrQgORg17NCQ6MkqPnvWiiLkOUh6c9gQweYGyDlycZMmXT3cdKda
wFemXn429hrPqbqTpyanvDDI8oCLDWyrcAQehxLh5HC1D1ObnJW5Hz6rjw3swpYWW1jUEFrtCt5H
T6mZqmmO4yZrC3b/YQltyQRjcTfSEveGhN5OiaXYiGKYhVriHNoDbM7JNvo0oZOikcTM7EMm1XZk
lOegz1w1OXEueNpCCUXW3LtDvaJd5fWoqREQq9+ahAISJYcmE8c+pFHoDIbzwuMahxiC4t0dHAfO
Aw6K/zV1e6fIfCuCzZ/3tTffCIPeC2esqwlgOxxTEIDGDc52a4vVZaWVlecxVzpl6C8fTtyRVwih
t8zc7bKYZZp+5yjA/7M7nynN0NnINEF81N2b33+WE3Vc0KZW59DD+4UI09K2hYxobO9GN733dbfZ
SX23i2b7AuDLJPRBouF2kiIQo2WqaTQaWeVhGecJncmMONJGNxfjplaI9w9hz8imjJjZmnm+CLZb
sOVoYh/AGJUcMGyPERFNxkZ14ssRRriDqwGaUc7eqX79KgPjM+Yhjz6qj3gds+k5VS3bMdIDrBHV
lqArY7jhBYovvKWDDUZs/DBbgq7g+z7r1Ht9xXCkpoWsvI5DIpE5xl7hBHCC/j7OCjgNN2EzCuAd
iuuqkl9+T96E8i+Av/6cH7yvgAXrtMlMGCdJxwmC0ZxAGSua863pUikyOb+oQ+bVH+FYmIX8yGMH
hyHQ4mXqa2l0p/d1QLWn7QG5Po/Zatc3XXA3Lkj0cTJKWefw2+jcbcj5AbEUh1XK7Hy6h+bV8Rzs
OyPJxqfTzX6sTwqrTNKNu6FNixyVQ2JzcxJ1Sq9gdrbIGHHNgDUqj4iiQQdRujdTqYUhsq4i5kzI
8zIW7+pri/Nw9CGzI+0Tnr9cJbfktTs8R2oSS/Wps+E/HdvzucwMF7t+yPxUEVmAuqrXzaJ3eQME
jcneIU8jfvmnozFzdoxk2fLxqeZcYXWa5d2mxETIZz5x3F0yuf+cNs9vTwnncfFqy8N2Hw19NnPy
/MrEn3G8aTT0/jTdug4gOB+xfLk6vil25BT0xb0NaDztPtE6aMmZKkSk4oVqyeevA6WQfqJWHtoO
8VaTjrB0D42lxeT1rfae0ablWflbZFOksXTxCVrwxSa4VrdXEaFXZx2ae2bX3OzmZZyM7+5iq3CH
6zDiH3seSKUM80ieXnJ8/xlPdmzq6AN1uQzlUFIW4ywkcBDvWuzmIE3uyTwGPaiACsN1TumXrbS4
F0f7rHPD3RSudH7uy82RSMq7DEBJZl0KHRpQ9rPFuj0PyAHHUN4Uclq1v+ANoUKVfMVh0U8O03uC
U4AgF6YMjY1DAKQLhjmBeWHF3OdUu5mJPP9/nToQe/K77lMoi3VLTTvHlvudRzGCD/4906kpl/vj
UrJrErG35TiECK2HfqqmXEAP/jTDYetrUpl3D+3omQYMTo+pX66IkGoFMrYmCjGD1m9ll6bB8JuO
zeqbsb5E5eTjGcZTzu+Po0ps8FUAR4eBEy5mXuaybWBSWR2su/zOMra/EXkzAkYSH17sdS0lhvPa
huOpaBVm21RHi+dYsyFnqrq8TTDeXRcsJTax/uCYL46N5/HQaNeqkYJs28Hz2Kx1+gfoJWTtMBiA
Fb0jt4yFyozcL4HAclt0duIty2bYdevfG8K933Oaf9pilHuEMteuHhjTV602VrCNXJAKjUQQUMuL
pho3XsuD12T99ZHaiklwpjIb5ncuP96vB0jJhnO0jxRmcGezDDI/qxEvN1Otf2scQX7u7fr57QWO
tu3t6ta3S89o3Z0N4dyVzzIo4lEjuQkfp/KaSsj37orMtHIEfNVEEFFr2hreRe2MTlio9ZLtkYX6
yIhjAyKIognV5XGYyvyFR1WWtoWnBkYxGhzNtr5oU1Je7xPVkKo5wXHJo+fuZGULtNSzlQsbLY6c
4koYd0+GGfVOqFNqjDDu/mX2Yt+DQqTXv3WDCJ975Z/DpCQSZsKg7m3cC0kGa5Aqxixw1ZnAGleN
KewgJjC3HmKujOjq//HVoM0JLZwPLA6WjZtw0+fdPkM3kfEzU54WDllZ9qF6hTMYpStDgAX6tZ7g
3XrtZo1ESz+Rvgs4dndH6IAQ6lvmMZPEwRJ1ZNoyd8CQ63op+a8cOon9J4NEwg0h3puA3vnzwP0i
qweZRgq8yOQy8YSUotTb6aHY6tgafyo3PumVxBYzk7mS2m8p4rhZZ7ADeZREHWHAd9ARqERAgyI2
L2Qcgxgor59m6Ts4mstwmaq1T6tfldkK2bwPyIUkgn7kCq2kYNQtCKyJQREkLkcNn1keHVx/6Kt/
LPoTwD59z66xJRk9GFP04JvoLuoVIb3NADd79Q9u0Qvf6HehIf8ChaAbmzHmU2O1+0/PtoFAGpX4
JxTc7n5gQ/rY465FeWX+d1875DQffD1uBZKq9LKbe9xoV+NGAyJZk+ywulTGvmS3lL0GkrrjbAiz
lGOKATaBYLawIQ4U8fOtZvYyvR4BnMhJIhaUZUqjV8lsytrbYJOBQw5C/C/rpZd9Tr46TgGkBkcX
rwA/TmuYgRaztEcxxVGEGSlR4ZsnNBAM4k/1VLg/HJUtNqM1ZFo52laorp1Lz7MnEgcF8iexPqsn
57L0XzyBUAS1vT0FaO4hrx21ekQaGG1fBileTX+T3Z5OLYlbQijVcMqiwbQlbaJjJXtNhHJhfDrf
otvVbBzM11YRW1UGgp45jWOoG6/IkD51gAyYU5P2670kVxOgg0Qs1VVt6G0n2EczpxU3TtT2ndp5
ywn7K6Od+96mrvTcc9H1vqfbAZDtzv9vkCY87Q52ur5oTCLuLbHHDJNofVN6F5nMX8/VDbW4vBiJ
0INkKfhuKYZ9Abxt5k022N0GF5AXhBPDGQmhzOmw8ZLXAomgznS285NZL10mAyRhLd6m5kKvF8j+
Ku5GWQSctWSnONlj0cOus54c6Oec5mVXDS9w0TmglvjMbLJN34GwLMr7UugAhITklYS/+paIK/eD
8RZLZ3GIPlyexg0SokU1RUOx2mEb4rx63UvVVeYR9gGj9xVHMpD9q7Ap/nldhQrM8gBTaC/eWtQZ
b4roQl6e7ki2hf3gOkMUaE+F5bXwKB8yiOmO8MhKm2KIOgPF3+ksKJpcN5CROuVJ5G7Pzs7lM6o+
r+QNgomQ5sjwYXYBhG4Ix4hXKGAbuffyu6m0rQ3+cRxoGjHYLKdKE9OS+HAiu02FZt6ZKnxqnUfb
sZq/NQVyDGI02lq9k6L1Mib1Rnu8qSavAQ/IDLU++dDjQm3UzcXrceOwzBZ9QmOqDJkBcYqxw5CY
bIUzc6Hluij9xRjXHYQckE0yJx3xMMt5EeAQ4iRS2fzGMwmQDfgYD7s3naFvK6smR3K9Zkpl7OS9
ulGkYMiGq016OzNWryoB5wg3eai6ae9IiF5v1Ryiz2S0/kb3Beuq3mfJfN25q/4hj1egG1iSoLRA
afrnQoJ8gDsb0YjsMSLEk29YtLl9MqKf121VbRxeLOAUQdoJnFet/PpTB3sh4H+SB9e0md+STicQ
W8iB9RDXQOQk8x/7543Qgg0LfPE0Y0lH3uSJrYQZK5KFtnO81QFy0rTdPtSDcA/0hTEsmJcOKfZ9
IyRZz3hR62nXn+N73bjZxysa9581JfH89Ucyk8mkmC3fJU5fg2X7XUXunFEGooRli/cY+NluDcne
YMYGunp/+PcEYqZXS29ZZdRmYnsgefhlLditbS4bZKqolt+LN9TLCzxDQsqIiuSP8at4UDLKRt0h
EjnXaYPoUgX1GxE8qIO/mHm+y6L5HN5/JlJyBccmseZG28TR0r6Yl/YUGDh8yQ3vi/E1XD2gyoU7
xXNSaVVn+VNLAN0eB3RzVYAy5MfCPayCl5+F4P3N9Nii1s2XLpr9FVeL9Nuzh1rs59r6umOo8vPd
O5iP8lRQ5DCbZcXuBt6NkqTin2X+wymQBQC0bnAVHZWrGR1ER0qF5iB//c5AyDN/bKVBHwgpKwNS
PVGJqdvwrM8UWDt3zYYbrs3meR8E71WFrHZaGTYmbzfQSZ0FnlP2wIAQpm5I8u6jlf5McHVow9Iq
mX2r/29tc8ZS/y4WxumVDiqpkLGnKaBgRvfw1j2AWCzrM6O0VUPNPPJlGWHTWclPZL9d356uK0Sg
I48JcjuCetsfIKmly33jm2vWIHwF6Z9a552sG8i1qgq6pYJl5JJY5yHtmVt5Qw8vAj70Qo1td3ug
E/uO4c+9mWPljyou/7tF5/w19avlv17Pqpp9kK4QJMXS1wVyBKQHoXJTVtMMsW0rvE0TVfTNpltB
fIa39wqDi5Ar/FJBzNxJO/q9gOEXM0u+lIyIaSfMXn/tWxS7r9gaDfP/vGkmQFeQu867SKt5pvfM
JwJW5+V5CI/p4Y8RX7AqsEjb2PnIHVRMCYeWqxciRVwJA2umy15LWGwHnJFzHj/CQ8a89uacSc40
sU/+dPk2EHZCugCb2mxh5eJe8kpr4Xsn4X4xjACBgytcbt/sSUmUuDfmVMGNyMy1lmbjFROmLEBT
9p6m7Xvbf3pCHIfusNlaKdlsAdfg+EnE6kcwziAzLYb6b1rWZBluNYWBc9+yOnf7omCfsknXCwcJ
/kzBIrklW328oKD5ZQ925xQbf/SK0d1hZG2/HeGttRcrNmwiTjGiNlDorjcz1JkVweA4DAejfPdk
k3yygzIMuPha2nQymQualTNRN1rm1hfkrhw/AN9VdFrRcv5UJtsYYiFmk1qFSe8NO/wQB8WGrDPR
MskGf3ANylVT4Zw6F6JTaqtv1ujW1HWpjAETTgIc7ON2wrW+g8NPWtGCtSH3uSrWCaoq600ToXeR
y28zwmMFpBqTEZf9KDm3afwH+0QSSRH9+xpWG/4jxpeNvr3nJHTKKlH7hSTOh8Iwh8Id3QVRPNTD
4UUtY/tiTF+5ZukBBrcEulQek+sbtPbjtjp70z8vwXJlJ5juw6Cn0FIHyFsEB3gZl0IKep9ygDgr
ktkbue3tUhgEujt/uGdosTJWJkKMZX7gl4JdF7Gvxp4woFLkB5TYnnz2ll494Sbjbiyd3t/uzFjj
zz9sN9oXp+VUvZci8vYi5dzhA3BKiq84c5xbow+Qb+uTrpNRRVFuV1hszq/xu7hGUXGb/L6xidUF
jus8WPRvrBeLj4LyRY7D5MzdO2U72nYPgdSX0spp+qqOri8rZ5yqVOIsuihfT+KwROJSFIOhVU4G
ZqbwcQz2yuz0hqY9YwmMYMwaRpIO+IifBOtEsFSsuLbZW0+fTzD9NfknHKb6E+88E631U0y/JxsB
Zx2mpTUJq38TXVVLX7G4aKdWda+g5GJrs9FRJu51RNdvlumNHEpgD3UoHmdAGEa4uUPNbVx1A7Jd
LBXvhdqnLAmVPwrwUgAUuuFg3VKo0BNz4P/b44JPNEDcX2fLqY5L0GBf2c+z8mmP65r4s6XJqvYV
wbOPjmj11UdxcXMTalUwnePGUSwIK9FxR50hE0X0brOLrM0SnceaA9nb9CCH+shura4kC04OETX3
HHPX490LRg/flYYkh+dOpzMreKIgFezgsSn7V1XTNIIw8Xv75QVn4Vuz93HgbJDqBmkj08rLkbLu
5pmFyrlj5A3oLqecInKVWPiZjEVVJOKx00TjhgY84eSiJFTF945awuUX59+oLa0Gl6w2vf1hlVGt
AQx5VTfPtTX8GU+tmFC0eY2x0MzCKkvsM3da04qWpB/o/FsAcUR6szSQ9EYZ+WMiOfBYR9HMeomQ
GsFWI9YM6zGOCrfetDaRAUJmgXnDK/4OkOumGopZM2k9lXorzI6zZLPqbGFxrQXgjtKK37DlOyeh
HoIre6r+7aYidQM1I5TiPN36vFp4/CbUsLG54f6BVypd1i0J2iGpwYi9IzXLUAQEivRFu/tcA1yG
FNzK0+sIhMkewGgbcjti/BJW1IaUdwkexeEOk4jnr2HiZQy+vb2vlB70Sm7RL70lUtgUJ8EglB90
2RUjlLubPBQvT5Ui2Is/+MHbtC1ljt/7I7i2Nw9YFqAOZ/MhrL3PEUZQ/fBMmYr/6rbAFe8IIycy
NAdkBfLU+L4YboIGCQ6vhyF64+3oo+5GKJ4u/I0SA7RF1KP1ikH00FFB5J4wDExbtokiaC3PytdS
5MO+ixlAwppM3A1ZuvPoURCquf4i2NA+o3uxNOwrgGLsW6tzFxCEOXP3rxxyU+AUbcQM4eJAdt/n
6GCjNHo+UZAz4DpuvIRX2Jg/PeyknR2nvqOOQRfZzBbXvED0DCp1cP6pGs0frmFx8V/lnenvZX7F
3MO6ZXOvFkzn2vdFe/e7oPCYbxsFYZ9rza9UHe/rQgS2VASpBWUvffW/qXo59gQSoKEjCzR6Yl1g
LjYip0l/dbz8c7j7OuIgzQ1VsKL5sZUbQZ8z3jG51lgUiUY5QwAY6D82VVpExpevYJsU6UST+9fk
5+OD6AzDBqTmDHWXbJxxOn04Wa8UShFwpWSKUjCsD8q8VpVR+vTEvNthEwVIvncAcMzC/qUOxfJ+
Tmuy4u2hiCOF9lbZQgYQIddcP5/R8PvYST2XTIGG9TWDv8y+w3DS2LcaARtANaF9/JgTymM/wWpm
UBSo5MI7dpR2iKg0Bc38ezhPQvfR9DGdO+uZI9ORMFxtTU29laYIKUJa19lIZtFOq6IhV3A1Ipfb
wFrcGeip7ZQIVE/j4HpSkexiB1h2Xid1vhcx+ZEsyYSOTOCKUbFMyUlFLVMe0Pu+IxIAP3070gUV
5C0LGm1S4iFkIA+cSRurZXQwVGGGYzpI8i4xkYv78gXrsc/KfQEfdTeQ3+eJoNBZ5X2wxk5gDFf/
SAsMEYU/Nf7U8ah8p+nEiyaQhBeF22f3AZu5AtwUJXPrqmIC5O7Msf3nfxPJr3ea0cgJIxMo4Tva
MmSfi4g/l7TjBU+t0HYhl3cloFM4k7GSSt7tNQlALwYvMcCn+EdiHu+OFmOKB0L1C+Q2Kn2YcHB4
3tJmnoJfLxCfS5uLt4npNstacewYfDIwq3uFjFthnefVkRMRjwigRrHCddPe+vPWQkd9vFbtxjTg
+BehEOipSMy87r3bjsSyESV1ksjt8JEtaVGgIBw2F678jmXTZ/ISBFU98C8jET6t3ftW2yfistmY
WK6OvhuNhFK/o7PdS4uteN91p2sy93HW7hiVTXEFFwHEbYGHqHMDh8mn531ysOeoJUbNlKUxai9X
BZR5gBlQbFTNPDj3LL5sWp0vinHsdCLPW1lHw8osZufz3w9eB22RFXCmOzODETXJZbyAD0u0ujga
CJ0a+qL5Ra0d3LLNScAmkPqmQvNCCcgxccdeaOO9sRa/TFhRehZZXe76xiv9HaRCL2Z/L8ry06A6
R1i++Pxh2Q6cLrm71JMFInVp4LwBxed//DRPaZv45BvsemR9bE3XCvfVEoqZ3vSen0Ut+ZpZnNI8
OTMFdq3XZ4eioUSILEGGBopveIQ6iy1pL2k0BPjsECJr6BNl8bNP7UsiyySls4ZA8X8Q0tZM9XXI
bSJiI9RCJE1xpQf0ARTlUm2sC99apg7jobAec1DCsDJLUOMD2b7An+HgnP32zCit8F/bK3eC/yuW
rbq2fr+L+ZC692G/XgaIW3E2JwWkbTcVQRnbO/eUcvlXwG96cuSQiywIX6NZKyQ9VaaMUwK/90Hp
cOwv6cCt2mkEVaKuN+y5n7XevM1qtIg1y74kr+U6DvhwkZ/FWSi92NpOM/Qvik4Ct6wsLv24avz/
M9ca82eli5pnl/yNJjI+YakE+oxuu7fcS5/ydPH4+bu+YkceWsbOvgXGZypsJx7Rl3yiu9GFDRXd
gUYjlFF/p9dKwBR89+QDrjUUGmV5ESoSsE3l0xYMhQNLGj4H3jlRv2zdySnGfyyAI3dcJ5vbDubE
vA9Fxn+Tr8LrxYImv0gfCRL4EhZR8F4Aajpp1Om31Isz0m3iGtnBYfE04JpgG/LCn1EenRS2mCMk
8OnVXnfDtYPDDhFF+8XvlbsQZRe4g/sgnqBC+3s3Axjm48ez34tZN3bqdKgmPhW4wxp04b1j/tz8
BCPOJk/NY2VlUZzu7mQ/RKychp+OTTxQt85tSFwrhquC5dzJM2bl+j+unznKSxBvDkXFZ9pysUzm
lyYdmhfCtclUUTyeELu4dal46xsaYKJhNpSNFZm5k5sQhxVMbfm1TVxr7t/jfmT/Vin/uhHqCCku
5T3Dx7CPoszmMb7Ebt3jYWpCpwu9g5atr0OUMNM+4hW2i1ut9dRgZBijI9WyvidKrqatb8AhH5H3
mCCrkg9rV8EkBVFG483WL/q3X+4vDXKSysS7BLfGWmzhe+GgST22wZUKjDMDF5Y/qgs+HMw1++0b
k906Sud2RQRTtW9se+ibro/NgI6jtY6EKxoioCNPPeDngNlJMw9OSD93EmS+dQgnw+S42AkeLmom
f4icFFF7zHMX8/WEnVWGA9eO3R2iZO2kOINmU+vNxN9guYdzXh0T77+nvJ1ZJGVukRQw312ArfDb
9AZ6VYi1pB6ViXTfcl0FdQQMQ0+NB7gdXKd2wjwSe+fHxQn73l7r7xjKP1UwTFfRSLKTnBQDnDjU
4P0XAgC/QvC3dOP0ecY+nxYUKUTWg4xGDLMz95Y7omKdjEkPf6Vmnq0UtIq/jfZAoR/2rId9270h
6/ujibfsaP/ITeONdvTpT0fuu7+LS8IR78x9yL6GihC+GTJKFlR06HGWvHhI9zlgzbFysgIlqsx3
fNPud2xZflqrDGQ2rilf3kg+33IrMw4AqCQYCV7ArIhkoxlaIe/C9pz/3yBxcBh3XQ4zEyoBgVhu
R97KJOXLxyDoJp3OmL5QRLxNO7oUY7LvqZq5lbpk2SsEyxpU6rNEVJman3li0/fKS83QMPNDmFoJ
YHUr2xubRNbyNuhWRE482hPfzVJhb2yXTaLpje2L434XbKqqIum4FenM4QrCy3zdSqYWdzQAwAN0
7eZg25/2FsuGcoiBXqkqoOlZACFKDIRst0G2xC9+Ccvh3XoPn0RZf3ByuyW6/S5qpobKvXa/O7Sr
/8N4lV7Ega3u6Zg3wy2Nsm7IYlZwYhT4scG0EAQFBBwJKbjq8apPpAkJHZUHA8cImw5ckgFMu3kd
9W+RmyiyHwH32RYapg0mK6x4R+9BLi7DjMSNphIJLe1e5LjjI1ZvGan9iN213h5d9Fkzj+zcSF8t
pva/I2qqB0U3VVfH0um/4er3p6FccwCVqm415ivj8kcWjAWu0EN7HtVZRq1ms5kYWA6Lnjuf3Ehj
DxBIO697A1ehNxQ4NPE94RMPPszcTYAjc+7b5Z+dF6go1u6olt3v294yR2tmFNvwuJIReHzAswY0
kV6cmTI/MqRNEsfZv1CMNvYFEts1mb5OUVbDpJGFK+n8M7huQg7+6G88ism2p2cLyzUkqolDA11h
2u1Ks+A043XdmjzmuJgbzGEerNw9WjU6qQCdNtiuKQlQlb+oChGDi1y19oSnArRkslCO8S0vyo/i
qjybufct/uJoVFnXTFxSO3W4kOvHUGkMbIauhG2V9tzQxQP+YWZjyvXS7X0VE1j0On09/w/wYS7u
hHXr5iL36NO/ozZgaKoarJ12YfZ5nLb8NJbVGtMxZaxumod32jd1KE1CpMUmGwMQ2UuGiqUQajse
TypOR7t+dNYvjb0Vr0gCoCNyEQ8EJRyAVHG1vlabZnOmBHvwhE/bSkDVaMX7E4YysjYOdMz4Ipkd
VF+/XNpsOg1kXXWUVJcLfoUr/eKU80B4j+23dlR1vzamgQYeRMWU8kmXxLjE+QOvwhsfCLTizlMw
V0mCo3IJW0zAM3wM8Gh+NFXpE5S1mXhA8Y9dnPOBuj9LE6RSADAA882RPviOsG/2ot1hIVbfV5OK
jT8iRupgsm6xJzSYfpjGsmsGBFCQKbZ+af4ROO6fkVsIMJHPqrFcvRRAlXqYZoMJsb0mJA2qtV62
hLNd4F2aprrfecTZzGr54wwrUUHUlelUFFC/37vKDHB3SkuNUY/ogxzLgeJCEg4Q6esY78AuCjRE
Vb+WS0uqA0P7+pGpkzJfdd//7/vEWM3f017oziiaSraUREV64kauIEyD//1caaV0rOfbq0ZupTRw
u5GBuGiQKASSmvKScTGVU1r4b7h8QD3Zlh7u/AJPvhvsmocP1xEomyhINtUQ6uPdwq9fZiBlDfd1
01eLeNkYsP5LHJ1F/JraJ2Dc8r9vBEXYnD/wBaUiwwUWvvjjjTOpfkDHZ3umy2dztr3Vo48xOT0x
NEIj/LJe8g0Pgg1yU0aNslsmhHx6ZHqSoLAVex4Ho1F8hLnpCckFtaH0cv9fg10XvRrW5Z9pauXo
oTFOQT4M+CRWm9c0HblsL9Bsj/M6//RpF8RpVWq/otZgw55GRHc/YnfzLZcXQz8fy8tOvy1SU37z
xa6vmRI2CMfbX27lBk0rb+E86dG2Qkje8HEWzLmHsUrAdoqquu6vFJ9Ph40A1VQWpxIPrvTOQE3s
UUs63z1xeiq4Ivy6/zmyCrG6RTTq6IMwE2gEo093Qc9plXV6++xSkDtUXA7JEKaehIdDcEcC6HQg
oi+x2w5+yVzsRXoQHrnyTHgd2ariUK6OR87CB6DaPbfu5YgKr+4WJIP23POWd0if6TNHAZm0H6Z1
/AMKHHxMDi72uXGREnjNnq0P3XYKp3oNr2bbpffsoAsSLEWscaudw+FKTZ+OsI/iXnSIAPXRCD1U
Ea64pTY6yhRkXde7dOZpSY48PIZ2LRqkeUEVZZgMtVN2cIS+oLIsvARQo9cdOe/Nm+xdRFz1osdV
gkMHp1d3d4ARvFXLNEeGk8MhdaMif4QlwLdR5UO83WqykZ3I7jeElV1erceuKz/HNK24Q3GfAift
+0tUgAatgv0zBZHxzMoAUSxh4yIRFIZ2s1JKmI74+r81lzHJPVKiuszbjLSgliL5XQGy5gsKJMz0
/boqAVDgusl0+pEB6mzl2yoYr53EyeiccJxzPFM5ygWxpRAhGj6xalk/zbkOTIZIL8WHGdIwx7hE
pdNoLXRj7CBaFuu/hUNvDVik05drEiCCE8eVcff0kpjM2HI1lGlWW+Vov67Ox5P1De8HxsnPZuA9
UlUU0j9ak98NPHkVba6X9SZxDeaq/sgReF5wAeDDj/drcfPufTUKNTOXEdBpZXRu1OhS51DyOWXY
go5QUSbMK7n9EcVGLZhfyt273DE83bQaB86GEmKtc3jW+JlGWjL9OmW+WqBS5xtIhFl7v5oO1elC
qmeEzg+kCwbFWs/xXVeVd9IjxvqQpGLuR2TQk93JsyeU0G2ISoeBEOzBXt7hw2vmvrXj+o8YnSeM
bkvGUxOuia060g1EhHK68DmaP+6O+vnf7VpV9mWPtluELh9cUNND3vPBx3nIFhI/wdi+Hzm9emZk
77WkCBGFrfYOpp0tY5wv1NkzBg4HD7wWnw9yfc087z6TY0qllKxLmWFIzCtOaCgObhwYDAPlKnlQ
dWL+zyAqoKAzqFBp67RzvqLq6NW6V0ohTbUgp6167I+yvjmPjRu9+WPFqtA8Y7U92m5vNq75ylQk
l1oy4BCCUWlUWmTenBlZ+EQVOvlo4fX37JOwUxu3BUc8rOjgRQ6VYrDOaeqdXcBRSlbvfWMfzkwJ
zgEBO6pttcmOr1L9Hvby6O6yh68H1oaXCGX6dh32+UpWyd6AUg9ggbNAzs6JU6tulK2crqQiu0je
j/vGMDjCeEXKXjtSo9ktb3p0ZMxHYN4bk0PRdgAq+TSgAfEd2niwXi2v3LQpXZ/oPjvzNyB+5QmW
T7DoBTvcY2m7LBHJj5ueZ+dI+0c0C8k4x4CNufunW+Xrpp2UixgjOjd9k6WpVIYn+i/Chf8C65ec
ULgVqctE1W6CcoCb981lPvbtT8vWXOnxW2ef37oyYgMvRNl8POPrABhoujBhnpUqVgXqPc/hWE66
k8yxjCQy/nn64HSNuv1M+r7X0M3FPgGLQ7PNYI3jLAutDbV5NHOF9jFCkB+J50dMttDamhDYgRco
rGPacmIg1KETMs757iLA837e0x79Po1Z4hJN/9QnISaTTJpx2/Iq76l21BIFc/UjXBRNm6GsyWOn
KHVwr1zmZq2nrisTfaZ9IpIx9RLzsRutiOQhrPC7jmK5k/IZZCr2N/7H+IpKVs2/RzOvhI2OHmqX
FeGVkUoOXaWiuq/1tmf5LjAEgIP/K89W9ciQpTO7KhytfgNZuUtHbGXz1Qd6K5uDiHPHIAnDQNU/
IE6h8EA9c7ReCW0C3h524FphZNMHNID3X2a9gU0XOiEJopKEXsgjMldN9ors8+Kk9sXJGfwTbFSR
q0XbqWBQAxm2rzxhacEN/gDvmAZU80UzwsCZIY5hNxAtiFMbt221UXVBMNYn8RoHbt5zy/DLS4L9
ViOOacDhco1H94tsyYsLIUGFsz6A/PBPHdfwObhNL0+0dQkiRZoiKOjDN86f0u+Yh2mYk0d+/T0F
pdrQ1bz3YoTcbBdJh3o+ocOxp9wpk0zMq5YW9X8qb0WG8oxED9b2nhKBwXSEdAgDqCCIVCaxXnBq
JivlUeekVRsMxHLVChD4jNj4ATZFGpgC4vWPWZbH+exIMYFwJD9dVg/4Zf77f/sOxplK25D7Vi/l
6Ew44/DPCF6cZARKU/3ZGXShY++wirVUw3r1fKsySgY2+FQRxth/ywQw7mPBwQnjfQXLn/xNjiQo
xPrdTpbLmOCB9XEeK1vwQp4qEZNp4YX0C8ot4JWcJViQ/wpmTdeLWZzP/UOKhkLeZ+FZxL8Kw3iZ
nHVVsRME1vZWN+jpRPhj6diutWQP3AiQMo78cx7utqyw1F6Pm9EMFY/w+rnbzUy8At9+M09FxnVJ
lJRAeiBalKnxV2iV+H4RF4fZv3mNN37+1MA2PnGGlq4sb/XoKHCkm3RiXV6J5B7L6VuylidW/xvN
R+rJL97P0Sv4DblSZpuBsZ2B/z5ZSmUKenakwTmMA9Gi+ua9n+ACX4PmrradTT7/WqMpvnT5zwP8
qnonr0pMzY5VBz9Eg7M4m1cNZa5Q/SDn3giGfeteLS0bsa8qnOi3Qlc4pcZk3UkQC9bnZaMSU7mU
W2cIoHZARgagoH5Pdy+/0wY65AgmIkxAQnORrxKzw/k/kmxb7LBC2pVC10oJaq0nNHvwg9y+M1Fs
8j8rus5BCkkCqYHrICgJq0a+wfE7+Oyaj9op0i+1Z1IUplyn8byO65/K6nod6mSWb0axvDG6XV7N
t+11MPxKnPHtDvJ8DFBPw05ky4mOf4Llga1876IA38SJX3YVDiwoAMlvoL6auy8r7c5KeF/Y2Gjs
1iGwecLufBglv5lNxVm1mdHSmNhEj0Wn41FuaintM0UJjyGII+AI+9qZw6DbuC9DYfzE8tbrtNgO
/JeIewMtItaDui8SX+8cZJO5l4Ydqv0+JTSxuXKMjOGCHY6SD0kkFcbMADpl5JrheMWq68fkGTby
imff7/vDO4XXbiZNLsdoE3Bw3xxip0CE6Tw+BLsysRbGJHBTu0REt2jX29FDKaG/eVEvUmhxu5yQ
QnbAG7hk9mElZiqWK+6nUiZOQZD3h30c4R82TlQ+Bgva0AxCacroMF4HeRSu5zJilaweOlcljDLW
bQRbmX45uB7+J5XzBvpG1JPlw9DzrSgLp+I/aPKuP46NFBHZJ0YkWaQCO0kVE/MMDYjJrUEQ2+Xc
LDB9nDOMUrgL3cFx8IUVwQdT82xO7yg/lQtn2BEt1Od4cxZyK7Nf1ut923Fllupel7WxfOUuhMog
AeW2fVl69bQPwpW50aj/sXR/xf7sT/2m8UOYLBBu8W+7OuoWTgolWFlFMAGaW0i2rMvi4YMsHfOf
uR58qA5YQ7rat4eJjGCL7fCS/MCQ45ZjLe8gIM24hFeEePNhDSZ1op8DTy2X9xeIfafhMG1vNUHK
Cexxw972Tuwj4mhGkp/P0JrtSD4QhZHhFihphLeFg9i4Ne4dhNzvIX7wxHVOjBI6pt/xZ3YaLQoB
pkF1Xc0UutBQfSTBRT35eDle8nWdASOYXpEguZgiFZsQN01Tr4etiQTWm4jZ9i/GO6MbOQ52oG6N
/76Agu4iJOV9j3YI/Id7lFw49KJwc5fDEHXhz5Ba0f5VyRVgp0M+A4LCSB3QOCllWbHN7NxyLMeM
GDCAlb99QHC3DxGGqpf7oK5UoNHg5vxRYELBBdqbihfzl6jzC/U7qoDwuGOHDojFv+2iETTEnrEb
u05iEdaMmi/VcwZNchBMosYRdUvV053jJGmZBMv7mmGBwtklRiELjoneppFKQFZ/YAKOmT3zFIjD
sGMDNtl+jDVmYJLutJxrE6U+cZnMnKoxSfz5quxaJ3skdP9Weg4182bNiZeFcWKHHlAWIaCP/tKr
XL3/cLEhsHKSwnWVd2NUqoCQFwGERAHqznWvlK64949llZzoADFxU6liO8XbfUA9GpuqJDDINCwm
6BSNo3FEttPykeugTxPlV0XQLMYkW/BTnGwf2BmMd59dECYMuNXXRkDcwL11fifumfUZOTN/08dE
QQ7/HyvfL/YnBV0vdlMLtzMBJWVLwpdXOkLOrADv8cB95sMnmMHunkaz3/L/EjYkF/1qizer+l4S
nxzzaFj+gZcdEPzhYbgxKbvPmI9HtRE+egfiW6FnTntR0fgweVmEyAM8KeJkFVFzf8+Jv5qLQKyJ
XpH82ySzcmxQHWP5grpbarLjV0dbIse6nbammU5Br5KrmZqeY5My4ZSP+JHx3A7799CmUuhQrv88
giHmg57uapiDEB6+TFurxViRBrTHTI41n1kHtUMR0pxfZ5Ys6OPZSDcfwCx9Wm5mC+59p6NHiM23
vupoWamlI5p72f0fBWmFfijYSCPlruqGGJKkHtPVkLTY6q24F3tZIhqJxgMt9XKiLrfE2c77epnx
63FLCJ3vzUH+mIYDWDqTNa7XFBU/JpQrdLhtUdxh5WfLkuirl/dtSGqml2nbAyLeXDiJbyIiy/V9
IIVdw62002ZGFRZrP8+aw6V27uL16jgoUH7bfbfg4/hr60Y6W+1qz2LDGbv99klj7gEv3wml/e8j
FAAM8Q+OuTw4kgC9L6lfhNSWhN+T+xjfcvkEoSxf4re9qX4gdWz2dWAZugiZoAzOStiSaJw4kvwJ
9XxPXaxguEqDWWCe6qYz+S6XGMrzsnDf5XxCrENCpUIzbdfuesHzkGmcrrQ14Fd45CKNHpILjDUs
+6SDik01/3yez+PaRXSlnuEjiJXjwEPijPHTfYVdiukWv8hxIPimhxD3N+x+roZTrFQDiovvuapg
UWuJVzhnqONcUzZ3OxzteDYpmVQpFbmsSnmJGHYjEv4ZY8Fq2+N575cy2tzUYZ1MuUzMk31lymNR
EZ4HA5UEVzzdiDGOLhrLU1ATwSb9M81929zE2R2HBWt95Zgv82n3u3Bma9x/4iv8yYZFlZDMvH2L
ru4bJp2cmmHfggPlk0QjsTZhYh/XEIyoq9uEvKunq6ii0qEhAO/ovd0uJWdpZN/YL1//wRglGKAp
n0ZmDOsu8ZliF9+0NoVRID4y3H/pAFecAYvOBo/NDCAQPSn/K0z7n+xt2+aD4bdjgVVALFNDwYN0
4dJhPTcHcQyuHtZ4JQxyuWAsA5Mw4eyeOrqNH7YSUBwK/B81FHUEHDDSUBOHVxFZAUhJhCMJ8uU3
+BjmpO5O0hpvScN0oD6KgWU9Kobth34GxauB6u99PuvIzpCwDMyjCXNl7mOyneHGHihEGXPFayA/
cztL42xJAONv44Cn5bAz5DWZ90KLTARGl/quiQxpyr7znJIfxyFLOJJDRH54RLD7UBNrESccR4Lf
Bq08QJauu1mtfNnerUb2JNZXyCg7iONkVf0zTO8pUirfUla93lz67t/U4qFnJfhiK43O87YSqqNf
gxnadNmDU/u9SFygBI3Pual14MGuL6VdJoWzUDcLW7/vnbLo9/3RGJtkweM9RwUsPUD40jjyh34E
QGJXLDeJRzVC0Qkqxi0KXesAWx77dtk7KTzmzYhv2HZrZ4E2c+9AmtUS1eSlzWr+COq+ryMob5CO
9zHoZ9iSjrtc9xBeozVEYjDVBieeRAY82myOU+1I64f8YnGcV/BU94rgpONz3/t1yjIrZZfCRGDP
gdCoH+qblqdsjMQ76bM+jCvWbS+cnls3zAAuERrlXjgnpb3XwFdotr2LkiOOD4YdMUyllMR9feK6
LlMS+iWWBa3rWM2v9mIizMkTJoPxVOD4sWyMca2IlasQSxU/KWQXVlX30vqhqS9InYZxI/7T1WP/
NWEBH6MDS8oGKBBNgzV0bDyuaVwDFq4n3R5m1mym95DT4S3jfQkmelGDcl009SMSMLpXJ3ZBSRdo
lwn5YEZvmu/qlHTBKZvMWbagfGicBV7wmCvzNmsDUa6y5TDhMPusrAoh+NCmTeK8gTdeF2vCMbeT
g8nuzqLSlrMO3uyCFMaPhgwYhyRSyI7X6aF7edbnFTIYLNde1cZHCbLYdOGGPXMM1ThfGGiDylM7
wwJhPbroHtn7ApYKVf3DGeF6zMtIO5IR0ogpg2zUC2xc5e+m7WHTx86bBksxZqjbrHhw6NDR7OPj
SvxYn44qN0UnvFoNzpWxhkrfKp+lyvqOgzxNc7XnMPSsguJSqJnP2TK6oWbmvTEUrSf3rBHutFSH
moE2SyizMCu8+BrzxPvD9jdbkbWaGkfJaMK+ZjmuZxHsgtR0a2BGDXsz/yLK0I9ZazMo6cx7UM5C
6lNfNEVPVA6c6iwYycA2+8KSQ0kps0V3PsS0QQZUQC7DIb4+GYxq1sSBuKHqSEsL6zve3y/xL90N
JeuxgPwgrF+8RtfWE4Cj0ZGlUXNug9IgH3nFtYw4NZF0Epx0ts4tSQtWAxMwf1kPE4QPipsnzjRH
xsnujXX6B8wupa88Vxek4H/JerHRESnmIsvohQDvW2g346zxHHMTDVt9EcgS9fgCWF6mlnsp05Ji
Gm5ut2iRiI9X0eQAZx5dLAKQftkCJgdgjhhBuxPHGEUqBRzDyIC7GcDma9k2bdClp60K3SUEjQVh
6o7tlhfXafz8Pm5IbXnwaML54c6ZHvxc8AuUF4156uocYsOnaXvtGPX//fmYqjexx7RheyOU5s77
PRb/HCtzvghwxDm5KhxCVCXzXIvw0cUkVfM8S97c9L26K2d/mH5NXmZb5PBK0Y+afTAMVNMlPkn/
8+y5Zv339NqWzwVu+GN9eP1V8TW4OUv3+rzGgAGZiBcKoP9GecdNywLl8aVi8YN70F4KKOhF9nYK
1ucr2f80bQdfKblsiQSoserLp02Yr40lZLnAyIAkIjlwSu2jUZo3jo2h/uTSfZD90rmPXg75SBkx
cUCXyK18h6Xyep3FKmkZywnd9dESf7oTtG2Ui2umDLr3QAdO4ApE7Qn73KfPmmV3+g6lO44EhPlF
oWWmbEgsQpOvsudIt149Fcr+07IkW73isebIXztzq6hNiCfXpLEsoIYdKtMBkhF5E32qOK/8N7i7
F+NyOkvZVAVCnAPq9/AL+tPKOGtQRwksOy9580svwSsq86mJWmzZSwRde4OKWrixoTYmNntyMgb4
gIyrfdHcdq+KMtev4J0Rx7gIDtapEBS1TCZf4U1iKnfBKwgMocKEV1pHlJZ0vH6kJycvmiaMwMeO
sQ10jHGLvdrdOPz1V4KkxBzOWyhQjLSBu1laHAheuvunLdONUYQu4MJpK9OxzPrMY5/eU4dzelst
7QyV7Ic4Aojp5T0cy4ZbYbdMqLkTfw+12VhIHtvG9GJPE34/w4lzxj3vuUBXq7Gl/ybOBwKAK3lU
XVy9hA8xEvdZvub59khcuBXQXCyY2DsOv9DFlUNr9sXzy4snMNQmXDTqhAthPz9KtUwc8wLHRfki
by1e1das2Ls+TPPc127lpsWPy6VnbIcsDE7eRxxaEPGP0jO0Flf3rAptQCaHQ18aBFXzvlmUZSdY
sL47+4Tza/vKlHeR8ExSfI5Si01uSyIT8rM8ZRDCOrpxf6j62MjEhnKqCrZgrj4tadAjpNyh8PcO
XEQH5haNjbVeZoD5grat/sFBqCWGbaYm/RJNJ7nTRB5/r7f5zjLTzNZwKlcUgu7sII9k5bl+LvRs
wsX8lVP36GJSUZvQFWC8k70XLatyxW7bd8uAUNRUH92bMKh8ACyUUWoECFLfst4bqJXsmYo/4fzl
IPTUl7e00K46oNcLuBaaIjG9nht4FZBjGxI2BpSYiGHEywjOfZ+xs0caDbbAMt4QF6ZUd4+02sEB
tC3dgCgmLgY+0fDEzRY9o/+ftsRf297VsLeKr6vKnxw5dLEA/DtcEV/16xX+BUvGGnjq+8yK2Yto
N/lAZo2/jCzy24JckNXsoOxbDfROAuj16iFim3p+ooUNM21jTNO3nJ+zf52i5Z0OVE11MIjGJvew
E4DRsJOMPe4p/RcMSC6SrKpHMAn6eeQhC262LgqBpL51xZh8zkkjrQi8zXTrrIQVGFXHvIpBAVuU
tBn+3cn+yQXAPrlvrYVxiZDTfJs8ZHz/aQRKv2SJreTTCv/uHQZsTOXOhGWdmWpizzzE0XhbvQfr
3Ba7IdNyN36zwLbwKaobqNkDuSTApuBXHG52c4pRfn58QIzn+D123d956dNJDZAk2tzUdS2SYMp9
WIf4BSG9kB12vqXnu0CS02xsTGzS/SzO45FXXh11+txbF1D9uM/+ZtOhZK944FjZPHnHbEr+3W7y
qsUxLXqRkLQvRITKSF7t6IhyWyJrrfLjrxqooN0Ucnm+lWy2DO1GlYvqRT57cApLUaKWYcKUzU6C
CB5yXw/MbgNoyeSDlSqiOt3KweDt1WJSJxxIrglIJE4TowpFUQkt4HRrJLqXBYfFqPMzbVWvv80w
Ef1nbdA+NbzysBCtv6Nh5yZMtEOM3T+lqV6Sw8fWP8loSmWMcvXE+QLa8ZzNiUWREYlwfhlz98Gr
iFEH+yIKN5d2BvcIR5zYM1D/vavGhZxC9CqQ9TSvxDxjjE2Eg4+gFsfn9UAJqTTRSLzsGD0utQM3
yqBjfzkOz8XmCKr5ibhbwr6FuAXfti1kEhTWTYzsC4bGFD9vPbsIcN6aDTIaCWR0AQISCY6nrdWY
G/u9QwmKSwwcySV3H3Qr/dnsHm8jatCQCWFmqjSYKpL8/xW92HBZ592NK1Y3oLBsiRMKEUE5NMgg
wPoVK8ZqeU5qQidFWBAy6wxJZ7LTjftYjgZ0yfU9RjgubaUveHiam0dFbuSK0Oz29zs//ZCriGPS
gleJJKDPIoVkKUQWClHkL9p3n1Ie1pW6VrioxAU+qUIpjBlErhE4PJ1j3eRmu5OzyddAD0bTvePE
JjC2xhJiprRgWp8LZLCOnemvppqp/o3nJKOaC8m8ydU3RnamP784SuZbCOBFlYaBatw/4ocHP90w
HeH95RjEvU9dKQHplrLx78OphjLNGq73jRAZ0yCsYLrCrmtUUvLft158TkEvRr1iyCD3XnrQlCZ2
SJ1u207I8B26KOrwLigmCchaFUr1s0JRLXdPL2rNu+/oqfLy3lG4QRIBu4b1zCWvYLqloQxB7z5R
gSbMXfYg33svS+0hzYFjMfMPdHTaHMUaKl/38hwklZXyHFJ9UeZS0jb4DbfbyteHyyGep/XXWuxE
POeUFjyo4/RrQlA/k/qcI8J+vmUc1tan2kssE95pMc1Mghzqad9mYkj+8T5Oje3ZHbPKF93NLut/
yHozxM9QcNncEPLDKkyIQcxBn1dF9kZN7/YDOPY36BTzn76EWbN9HbElvsV7xe17UDZTQ6ejzpdU
ycFBu1SQWO6atHUBFvx1CaPEJNHHdQSOrni32OYE8+SmJ6nSSrCNJAwbwBdVfiHJ+N4hTM/fSJRz
dxe+vZyIzaYA6mhBUANAUZ3RjHUw7RWqoRStxlnJXnQVxHm1nsRxk39m0xYhyzsCO+noezyqa1oI
OGIHFBUqBgSfEPMgW6eWOau2LgojcPSB6Xuq4xXYGwjLKIcPFwgZkE2m5yAnmTYv3qwSTkagE0e5
NCMpNJ/tuWy2VhEQDjYVOeiiemGsHBaMVj/RNgRK7LKl9WF2IifBJmpe5hFLV8/pQaS0sxU796yI
ytD9rWzigUHngQUIHDQYVhRE8pR+xSvsBTqXukRGaWge2ZxeIbAbinM3xAWMJ6UHPdapDLUwvBHg
cGxsKGbK8jTqulUdKBdCiN3ajRswO+29OAGJQ7Z2mHOP9W3yPbB+VJUJMpdk3p693eLVpFTudqlb
byauSH1zXx24XHCdZz3T9nWxw8XLRMCh3MsG3UERLBGpyT3q7T7MS+ddn35xhr4XWFbCKUVboLRZ
WHLZkt05z+J/WYtaitB8M32fe+0I9nI99c8cJgDluLDwiP8AQLFjdhlGm9A/mwjKcqmwV4xrfshl
j95zNKM0cUK9LgT4cRLuOJtzQPnIZ+C3CaE6Q3pz/odQkDEwbubDdM3lz06BcmI3QJgJJqhqeZcM
f14OY6tn7gdfWb9xKXlafiBVu3u+irIQSqJVqJ+kle3qcWZV8YOd41xVcF0TZ52D+1+Gy3y4+f6y
UgrBTxcGAlqVcnQbgm7aI4B6ZWYTMlTu8PbWaIIPbRKgTnisR63N+65mQZXcr4/mdi/d++mknBBI
PQCLaDkERXIbkmac/LCtjRzuQkJeYzqlWVqJIhtMayv5nSCU0fhJpFZAWocuHMla8hr7xWQuCiXW
qd2/g40AA3zMjDRjQuTQo7lBmMhI2kqtxsS3xaslgkbuJAvBN75K5udr4uWjwaWO3Xh+N8v4WTKc
SKo/w9jkzc7Q/848Ic2IYZivaxdJnd/H9+yJXsUoMp5K3+j6bRjtDdja0g9EuiXOGrDw8ZGG8PNo
1tCyJfpzsOwlTpOHCloVxR3yCVsuxkFC82/kIInhPSOFDaAIUIeXX6heuffO6aIokHsfVdYUCr5E
BQsbxC279dEY9g77glqegWGQM4ww/TgEFyxTi+ZW/V9wOY3t2gLSzZlwDqA/8zCLco6/g9dkYHjj
0uSrJ5DiFwQT0oJ0qLVjf81rHmT8/IRMoQto3qoeW7gDNnAqEqRgHZ+HCJDMjan9JBMNYR1/nNvR
Jzsfn2j8F5lXwHMtXPIcFLu40Hf44h9WdA18aiIKmXdfcLriLalabHHxq2XZTqdgX3MVC/ftImcq
MssKyBDfOAHE26IA86eFHRw/C8Dz4AGcPlSZZtfzCtAWdXkc6DayorJZ91rYhyW4JNp4U3QNC6lw
RwVUEEU/wQ1X86WYi6MNVfiAB6OR5edxWGbcoftuWTKJrHsk+XnqnMVWh0dpsVvoILYUGtz1S97l
9qDxaKOee93/M3nk25gXShz6AsbrNk/+hHaVDEZ82qW2EV5k0eTQzHSwKqYYBFdq8hrOFVZb2rYy
nm3yoGVQutWnrsgSuFbfgYZUymzyibN6ZMZrFdW8+w14IN0vLYQ8DVnp+A8ujjjVRBUm5AeE6K8f
u3OqY7SJyevWJOZawdEZpIxDVibtTDoowpyWe9oRHPd/y/pO2Hee7YSl8EyQZzq6hGPoqwmqu8Yo
KQ8wdivjY/CioItHrKI76Sy9u918U+QOrSpcXaITkTvY4s3yQzrC7HNjpc9cWrAyEqIrz43HSR5H
JxSPJpfYykdYKSHfCUiLBLQBFIdrbKXqPfgau4WivxHS6ifFA1HGZ/ltDL71WkS51TinaOm2pdAM
LAahE9dlXjPResn2jHlWVZZWNoJQ0ToG6lM742/SV5Y5sETCRZcb4E0SRsp7ajeOy+6+OJEG5ZIw
YOeJrRrMhuyT+bY0hrvWAvrprxY+KK3Tk7qO+I+Vy3aG+3JPC+1lu0FQKXIGEfxzxX8SX7eIoqDs
33oCepXLhDf4iBwzdvj1Y9PkNs19usc2UelZrVmLijzmmuUQeTju+vqWJMo0rqJoh5CHmrpAGY2m
jfbQ4ERy8n9OLZmmeoWPaPzhZHc1p8yDGg1SKi/5pcnkRrxJxHxAvOnVPfvTn3eRsS1LybTyJvwH
5g9Sf+m7hNeIcXiYgM9klcBHUlud7ZKAQ5Yv0Fqabxu53troToqZGqcAIWLw30kSghxWBykHY4bL
A79KkRuh30u2DUa9EmnrEHc9weN5uZEBYbH1S0wuT7MOyuwrHLuPvO0uLkdoxLCxj1Gts+7kGV0n
KVfha6An2XHrfqO5Gyw9wFcmA0rPIYdhMi7APycJe3osVo//QKTUkaD3c0lKQZcLzzOXrKKYn8XF
+sXre5/jszgvncb8KwMNeudtOfbMbqMQcpPhcPlrpFKEs2fq3zdf/Njs7cWtU8B5kvLsTExe6TFA
kQfHchL6LK7bchXF2hzOP1FutuhYdXHZ20CmqkNiqh33iBcSHQfCnwOkt8UiwXnjs1cexKd6wph0
jC0Zr9Fv+b1CV/ye+FBK1XvNiKRU2gc6qqz0egGQsC4I7i0IZ+8+4/U3OauZsxV3VJKTba2BNpVp
rEQPpk4tBOHAtqNCFe1q3bqd4MprM5IpgWiEDg+uvD6O9WP4lgOaJ33wFmz2kyLZZLYqTPSDGrrY
QuEKv000dEQYTLAEunGod5b6JFzGJHT8RdUEEbnYtEbTtlB854m1xVqXCZg7QxOXe+ELmNwJ2OMn
Yq1vt6G8e0wBx7Lr49jOg+aOKmvs6gaj0gEl+wc3oSdYZMCF0rRzq3BpelNg1yyRw3RFv3omoSOb
xpR1rsqNDXZ8nn3WP/iWBr1O1vMBF50gXSiXkWlKMUdYhldHqM7z8FVtk522S8fNJNd7WxgG5MSz
0IeHOtt43y+RAUJXPBA3J05p2WvUHkXpdlPaeg389xm+OTsgmYrAmHy7bXASbuNQ4Kv+F6Nppd8s
bsiLySjAkUiddQVPBYIrfuSuPqNItn4z4401UUwaB+eZ74nxNcnwKhZRI/iJevLmt/ZFOya5duNd
YUINAOQ1bAWwfVw1kKSJsxRklSJljYVZ/f1q1sKbhT4ms3Q8gnOCuWRf3W3tM7pG71VspQ/u8mv5
VEE1En5Abn8YBj0hcitZjoW6eb+MW4UU/ii94DI8jH88nGgIglNDA2ov6p+mZRnIdrpLuGDkiKbr
XsihED9k7P9ZXX9BQKhKP/L1LPKWDkimG2/cXXF1yocfFlSIOVNXXaohi0LDteAlzHpNs8qUhUwk
+NWZT34q0IpFiqj49xFuJygMtEDjhCHdONh22VuLwQ1Vk8A9KuxhiNcF/lYdbKdcxoG7tXT8fB9e
qeijQZx1TJ9c1c178g9FXd/oBuvMPIwaHR0S3Bk8AsOiLytwfwOQVl8X9olQ9IXmz/S5wm0WVXc3
BH7QES5q2GvXJcSNNUrLxc2ENeb0RlrJjTP8gSP4JZrwUTdD5qmBQmHsJgiVyzKgLve4yjDzBtHq
0QyOlZ9B4nsn9JQi1zWByFXs6eOg1/KBZuSWJQagKpVxqdLvMufAOMvoFSgf6VDthe0MdG9kJsmL
Nwy0c2ZVrKkm6yuijA5mAHf/mOuri3+pv8pgPWPI8qlh8X+gAHp7e9xM0GZEmCZGBZjQYT+Eyw97
GLFBt1IoAU3tI1KokXWSH9SkHrOz+vLKBxonYSMSJmwp370TCJRR17bXkVOxC2NwsYnJbJ8TOlZF
GU8eMRGWtgeqlCgcvWN7iSICdOcvJb5sMfD5/EUlnv/wv9EQkTI/FFM0hMkGnsPhudRVPeY02J0I
N+qcRmL/G/MHE/5tl/9lbs5a5cTxha4d5fz5Wj0cyQ9yGDJv13vrJNdx6r5t1vMibKvNC+PaVIE+
yOT3egconrEa32DIJAwN54ySOXxgKLiZ5Rn+5uFhK1qgCII1UuIUTYY11oOlABr54dE9BNO9+85B
VXE/8tGXlyTsq8Jdc3da2acRH4zDLXFovG/TZNeimNbDeijhwnotQ9U9X1Z3Aws95I223EThTYf9
VEiEL9val5dhfNRY+ZplBLb1XiQOO1I33B29MT7cKNZR7acqcKLRDYmIf4xT0PXIM3c5CjnbXSsl
FiRr9YZNN27AAGmgB7FZBQRpjP7i/5IhqavFvevXEjqQ0Bj8GguQ4pE+JRvVV2s5KgSZ+WFP33T5
/Etg0qJikhQ/6ZRN0WfMlKuttlwjYB9/4vFqr9b1A/qfmBkLEFN3cXYEUuy2VHAgOPd/hnGFVf6C
kPtUcbifYP3NNBd70HFsS0OCPW+5Nejuen3zMZCOFbQOR/BvKIS/RFjgG4na67QpivhfXvpLbcWS
hQss0wuj0akV88bj7xgaQ1l4MjE6TGvN/Owln6beTk1Kw2IyvCAfpDSVr+xFw3QTHVi7egvjJL5g
4T4zwLeX1wpGn3A5kIrfvMwPF2nZpB7vKnMA61GtWT6DN3mCJkpyRL2Jj3PFGQDYjwgX6vfv1m30
r9fb8e9Gt9IkXoBryhk00mVRkvlDJRuYA/YGB+SqWmvPJqWM9jGBwd4nIdz9gbPJ1St/MOG3Pa3z
oDDBeDO1LFF/Mh3zCsMiXAIaoix6ospmVzYUTjok+zU1nsV3D2zoVGEULjxYFNGuAK3reB5NAGQf
jkY+0msF8U/ORQv6XQDrp+YceScgyOfAiJxHfgAbUXMGRn1lmm3kKORyDigEczl+07ka5mdFH+li
OscRNAmKRaFo6Pchm0hkaYEffte5TfZBHKo7gPFCquLbH9xGg1l4OPPWLfA1B5RQfqUfywt7fFpm
VBeFE2BnRTpq8FlRXvWrhEATjxr/lF4BmQ+QeKBPU2kczh27kySUNi8u3x2CDmhZqH48OfmMAtNz
KJbOz8KMy3tO5ERZa9Tj1V5Ky8sVdPCyaQfdvkzFzemwdbDfFrAqKxgCPAgvY2mOF9A/dF8ioNzE
REPVeJTyzOhbkvFK4XZ5d2R3YfMTX9PMEdb5dt+NTuqqn68+fT4tGGLEGk9v5d4lfVuqOZrBnN4L
7qd4JSAwsIdmStkWLFPq1aNrf36QkfHnrLTnKsRhJIJdiA4m3RrG86w/27Ivc/dxTV+ZrBPkwa08
4jqu4J8uEUZ440pAhIRYeNyJQtk1MSd5W3HfJRGib9K6kkazEz5SsD11nnVO5e2HvzZMbbfirMdv
pAajbw4+yYqhoMV1yFMjYik41dcPPUix/Zh/jYl3dpIVy2L8NmlwhxuP7v3S/iCfyxY0KNkSZRu7
y2oX6zv9RSCQQyateSNYA2C2itSxK0/is7hJLP0M1ZbhvO5ajZIrGU703/+D9cU3rwf+lOffwj8h
HKbW8OUoyJ0vI+6KskFYIPuTnexFZnHZR01P02Td3h4FjXISPusiRozawKnIsnfWYJHf+yXfCL/3
KsZQQ+NGnRh0XdGsn0+J+wvKmH7crWtPa2Tkzhoz5MfmoRLaEKVZq9EYMT41VZw1XNbqZG8mtHku
H2PhMtVTpw13OOYnL6lNeg79gmaMoiNGud9c6NLpc2W5Vc+sCjAIZqyxi46v+dtTMwOcStrEs1zp
MmyagbAgtnYkAfxDODpiW1Ca0BZsM5duUTiS5ITv+C0T6WAGvyg/yt+LQrsQb6TE0JLhejd8TaLi
z8s/ir0X93Qh6oIASjeab18M0pPbW74hISQsuBfe615Gqh/82JWavqGuuAI+fiUNTkWlyUi9xKNt
jbMfBO2ag76dgcam7JtSZz2aLNvR6NbsvoGuhCL42stzpTFSbmU5eiuurDm0zsREgYaJzH11TgG7
9nFf0Fmy/MGNErb7tP2W7SznMT3FedFxcgHsee6Gg4/X28GZDZI+ntpXUXUJALbE8OLIx18ineSx
Yj3xFwoEKoeiSEuS/bSx+/zn4kKBilTFUC/rYNoGGxQ2/CiLxwiU3z5W9u57ydy6G4nxouUPGInG
eed1Dk7+32bsoWyLcPwDPK7dPexXMTiRGN9ojhgflGYv7AHUqy6B3Wo2ON0OjTFasDLLVNSCafj0
tt0SeZPXyrMaplw3HorMlQ/ey+wIpdVpTk6i2e/Gc8iI7n1Y82uZDJZ1xXD0lDKuFCXt/y+HAK/Y
rsbW9869u4p2j8KzR/saVWcNZyV9KDvCAobrrpfZ07mEm0qERmS5u0djKi9VsKwmOMTjkr+oSDkB
bbOWSvfNEfnj+buo0X3lcjF+zGXYulR5HdZ7NFzSYvumrGV+96FooQiK2FGhlMsjwIEUXEWcfEEp
rfVnuYKOmz8INVaE0SeRStoH60SF6Uuw+you1go6Rg2UiYjQbTDMGZyquH3pcVUfw3+FyDcMcFXd
uWn+sSCCh910STPWFprxvnpG8s8vMMdZ59LCfCGbm8aU7cgrt7YYAI+mxj3uwh10/KdmQVQR7mU2
yI0pPkhjuPx/RZFhkJiPh2jW7IsBYsC2zWbgChY8D/4coqZyprZqnArCgI3CYJZ+P+eoL7lEEn+e
TPyHL8kifPbqLKs14TGPEtg4Az+kpV3ZHbBzcPMHDZ1pYiMC+q99Mu2mFIhIBHm6gIW2oIlfY6lC
XzFEMoByejJXoGEK+Jo+sju7+PLlPWR4d5jKp7sIEsy0vZepJzuXDXsgCeDMSNM+3LZFUFJ4UZ9W
aH/tPKs0QSrr9c1jIT4Tqu3lnMUuzQPhN7Rl8bbGCIzRBW90eKSmkgw6V9QBpOkXygub255/Pk1d
GJ/9yiR++KheqthbdWXxukvMhr0SRuAkPW9sD8+5HcdjjfERX4Or6q0R5nPS1/DU+sEfwNI0h83s
bpYkj3DGuukPjE8pEXjgFm5/Zg1xb9c5TMQ2xEVHfymk1muAbQF5GtgokwzCkzokqBAVcaNbPb7t
LkiHQ6cCPwigJcF9UNZMy/2N8HjXFzW1OQjvYHFsEk5BJjqSxQBxHFBqHUFxMhWtLmNqsxvZh9Lg
Q7kG9qZOtYcQilwE6R8vWMv84sSIb2MEWKIRi1oKCgaVB+HAaVJte9r0J4A+GDegGGdtzEeMxwyj
DozkfwZ+uoNnVkWqffypqIooFyaKtQt5deeOpAF+9B4QUgB9kqZItLAYByyp5jsygRggahMugjQr
VYuc0QJHZ0H7vvR0rZN6gTAZvr6ijcMBoxYhPYgUfM6YRoWcMYXLT19IjbQpXSY1jU7oAx2cluWA
lMVtK4ykJhyrkCHEu4PVH55u1TmjglyD2LiT1cUV0YsGADrQ3lzo9Ouob5MHmUUeT/tk0b8URM6J
YBZr2vnYrm3cs8qDmhZYqxiwAyQysSc5IBkObM9ZAl+dKW6sXfa1lKOLBU/5LfwQan0DXy6Lv8hj
sNnTTwYCIch0GuQLxyqoChYRinyMCgSSC2CvvTeHjq1mpqiOysp1oetxMrTid+SVirFGpChc+TgP
yH2rTET34AvDOSh0//x8o14CXSjN7UQJsjERaVvw5j3T0myg7SkKy2spf0lvEI+2n9Tg0KUPUobB
CfXsUktBAG0ggLaohUeqp+E58dhgeXhBX9RfmFAfkNyT5S1csrL9l5at6Zhqf3HMhWeN2m+66dXS
52G4izZeCObhMZgkLvk9xSltygllwziwehXuyHQDcJR6k10eX/5iNdgh2puEIx1ofGTrwHExHKSU
jcBmD+DUzB7+sIeizBQ7KzMT02BOgXSj0QE9D3fnt7eCP+Pfr9V1+nEnHfcnj+JmU2HuZYajTMMp
u4QnD5sPFYHg0URUIFULJrCmlPjv0/tiL5eUsOk/2LibNm+Z4EZnxlMX8o+ZH4ye1dn+HSex8JVu
4zDQc581rEK/4WC677y3qtSCHhFhqBEPeiLQJx0VnkylfTctxjMx3oLzj6B3MptRhiek9OQfEaNp
7w/cauQVQJKERsx7gYUgK9U3iVuueX3++lVRps4Nel4v9/Y3C6bWT0/gSBxk7NxjT7t0BAzTmSg6
qfV+zgKTdx7bDwaxyte+/t0FLqxMpztrgfLd2NZze57pyF2n6fZ5RnlQOmO7u/cUQRWn7t9MvXKs
JXjXcxbV8TZPXbLrZW5A/X/Q6qZs7MGsFxPosrUA4OZz3NvhyB+UdMzM6N3EuvJmdnujOSD6DT3u
fjU0ztX+fBQV48L3yRrCMrT9iZ9qPS4Z58dm4asP0Wl/wywiz6YglFj7oZ+QyXOPS9T+EREcVQ3J
/ONjxp8c2zCIsFoVnXhlQC2laV2DDJU5fVHWLTECZKPIAglI4HOCWOUXnKmscceUJ8KIpk2Tw8gL
jGRZzPwXv9UeatFaGO0Px0bCYZPePmRJLAzRaP0d+cT9BQLSBw1B6vfKwpL09HvLZ/EcmK5q39VQ
fnRtd6eZIh6j9MWdj/yeOnX3d/Vn/zkSZW7D/VKocI+FLuaAidM+YX85KDdVps43V2O+egJH3M/W
/WRdDQIjQ/DiYxWvgx0p2dXTnH6ox+0966fPh+U38BJU5+TSIE8yxweJ9TBmVVq7rX4CVxSiTAKa
aY5pULT8kX6EoLwezBOoVISAK+bDOxPXgo2OzXxcF7jDcncM2ejuTfJp+ivyxJPyFpV5IqRhMDsT
fL/vF7sYxfquk0gatY48FRWK1Y1DhqPamipQr0XbmF9pkC5ZU0qNgwoC6cZSWttHw3eEfCA2+WlK
iZIRG4crKjw7Smmn4Ndcn1T/wcptb4xuhFeApZa/A/4S63W2u8xqcSY/6ZjxwRSaMwE0etCK34HO
xp++dhiY2BodcwELSOH450uH093Nayp9oRNkrQgp3jXulW202KjsZtf07iOinriH4xdK0Fz4ehAP
SmqbjGrj2jbVMb8hDWGjmwArV4j0Qat9UEXKKy/scymphec7QTR8I1cpfGLTBlAOXkSA4a6jAaJb
BVLEt0MKAS6VtRMaooDAemBpeBegGTYPpp7AGz9CYLnI8K1Lij/b7oksQkmRCoTOVww2cmrmEdBR
cmnkcq12LL2JkDJFvYdOvJvqf17USNz4708w/urplDl9sG37IfawQ3UVoglEZh9SYys+m7dnbW8C
VN5Bzv9XkjIwU5Py7xOoOXmYUezIsjZBtD5LC2bIvfsDRFn3hrmrfJYMRBlVtga0jAXOpmALHxFe
G+BK09vfWVMXzECZ/ksbM3VNM+DLJ0zpYEadbQrHnRtWfDG9XNbE8D5I2L4zinRSHkyxSIgxByo0
r5NjgPqJwvAkWKOP/mYO85FW92hQTF1fmpL2fRKOHG40lqj6dvq7j+pdWhhryQfROjZr39Dp/mLK
ACxRVqMWx5g6D225UUbGsrjIu6KtXrq7pW6B6j+VnOLrA5CfuUdfHX3SGpxEAvuHgYXKn0EroaKy
thyB3VLJJisP8AwJHNS5HtBFg0VuuOSa97Xaci8yMrbYWtXijQxd2WadRaLAIPU66Wr2Ymys5W/1
dHyd4fq6RBpCYRKtRn08FIMAtuPESO9OwE7uhTthgU/S7WR61Qcf3O+0lZ6j6blctX4LadSY794y
dxmByWo1K/q1j6CelWzY/lxP7WzPutHjExbM7SpLrAx7TDLzzHfOHnJ+ILDIKh2bQlA3NxcRWo3x
AVFdxW65Oz5pN3irU8ZrGJnfdM5MattGRp6IoiMwqfHS4v4aWsjgAmagjyyWjmhERpJCK7luagoN
vpMZCk/aNG8TR8Iah6QyyZh8wZtK2op1c4LuzzaPJGn8Ssxb7OGj5CT/PTNhfizuZeD/TdYSHRPP
BnO8PFo8bSlGjFnausro4/COQ+rC1grJLSQClgNs9psLIcNk+YzesuVcVawwv9dr0SkZpS/zwSPT
nXRdOoV1bsCAls/k6VxdfK9hZdr+GZguwsc9RbngQR2PNxZYi1eHvhO5yRnxeLZPB1hTeo8HUmUq
DFr9BHg55pPbJxvLnPC0gQVwGilKPzGrU45hgtem1jfXsnT2Bw/aeTXZV/Z9JBpM8nUUCcJc3Wu2
UiVs13/PNxZ7R/U/6tdg2wKAKsfuVD1e8prunJv5QLot9Ifg/flt62Xa5wbawqFMLafSvvn78OCh
kv3YnxPY1qFuTNMFjfp2IAzqPTF5ycZcAJYxkZsrEyxhmxOv6qFUAL00o/ZxgZCwdk755DU0vFlD
jzyzGK5nUTqj3jYqb0G95MjTgYL9rnBdJCIrznY4bUxB35wPiaZDmFeMjiF38m7+ypOmP7y6wik/
Hhz14MjE/tBu+cH46BR3GSZ2hX/xnaJa7+mGJdk0q8BJw4HJqgY0qUdPfbY8N7uyAt/6suleOD7Y
GPYXw/QuC0RyOxenM3fBDkYBe5qNYM8DRVjkceqzA9T/UY0heeAqXj/p1cRFmbxHUD/IPAq6KFa5
wxexX5iF1dnBH5+Hy0w3FKfAAo1suW0W64fXVlKYhLMXt0VJtwsbfeWSjQKkNLddcl5pYYxxVDNz
/BRtNEyQZt7OFV9QJlMtFqI/Oj7XuRiielSi3O6I9yRHQZMIRFGotjTv6UPHSRAcfOI2GrtKLBD0
ujJZbubkUcgjYosjuyHgUsK+b9scvv8UfE9ObcKG21U42WFO6DGrnhN8G0AnJBKOX90yikk5Zh3R
EaLBoEvc/g6Ll3HWGmlsjA6lqQogULdGRCxWfSQNTEjYWhMU1wB+nmHWpaXk1cTRGynv5lDn3LdO
fpNcRduWMB7PYONFQOTNKgyeYpqmkpSpowEFoS1eHRzY5PIJlK5YqUIYtOlprdatwPpsmFwD0Y8a
4odkgLSo4q6cQtMO10Ay1NNU48MwQw7shyHzUvKW23exsjjm04hLkaBF6/aRbWrha7A8NJcBwAda
3zTn/drvG39AXfP4fdbbmjVJCajMit9lyXnLl2rkRrKs4Re3pei0TUCAZb9k35SC3U3diQpbXBED
SXtXuakstt1anKTn+z6llH7t0cmaO9/fbITjOuvq4dG6gK+xhcUyFtI9V+TZaKPPKqnOSnvKlPy4
aBwNnhAJqjqc3wGaAqjEhI/S9OvXNhpix75Je1KV5guNFdQUjwgewO3pdPCjzn6GpinBMuT+KEYg
Kbfkn6SZ7Nxg55fewWwJg+B4DVSHbNcDc/KGgru397aawAP2zVxAte1UePTGFx+9e9uf9AkXIDSP
/NXge1W59vwAvGS+4/38iIPTanhaq6UMCO5/JIwHPEskazug8IVVeggkqTE6vsyuoKQPNUlP0ICs
t1w/7p8kSO4eJRWYe8sgVObIo8jLqCIodEqD9k1oFvVRKsNXNnX3Mp8q8EkqwuXuWspWGxeRXqmd
/aP8eefDWEBKsZpnqXuL0PRRFrqRB8HlA0clO9QCOlMm8oMoUNY+P/KmwdTzJM+Ar69k3S9FJGBp
wc/8bpstcGI8H1bIj8SXNXZQExdrIY9ZggzZ7zeh8bHwn6dL0nv4NgZ7hPSEmSKQBBJR8iccqBev
KLG3e2q1DolMSaN48qbY68HEYB2+SRJDAXBmWcLQKpHECG37oCvVzYh2DT45BlMjk3ZCTBwykxts
eOKdTmvYPwAUykuCXw0LDX2Xgsl6YeC1XXIt/wYO/jCNJvuEyjlMNalq1iTQSfoAS0u91mLgd44C
4eVs/SykXITJjsYSJKNI8ogMYnYJ4AtcGtv1VpTEnLac6XRE0EjsoonSEz46EICfpkYYDcWO5V/x
OnbH/rcbRHQe++iIBkif59irUpRlk4xhC3ZTX/FT2rkH+L5a35RZyYcYFZgL/2PYXtrw837s3imu
Zi82fBIkzv7H54aX8qsncV2RLC5TzcDPZRA7s6g0pjLKrISkuTjy7F6+5oVlSLW1IrixcIKJm8YF
SNRVEy1EQg/c1ehDXB/Kl2q+nQ599PfOYeGkFwEodRAljI+ch/jIeuyoKeHcsy7h7zOW2/sO9aQy
sRWiVj64WedInoupbWFnAptwZS3s7rw39QR7zEpXuNRr16hLoK43X3Qj2hDUdxuHBJNZ28SFs+iD
nDRhqzDhWo2916nmln7ZvJ8iW9wAM6SuRp2lwHiFhyjE6ZCA/koyKrMcbfWZAKZY0/1MQdA1cWWQ
9CRf1QpSBuOUiitnzfuJv5J7ZdPtQ61PAFPgYcaD8jTGoL5L3QfWoQ3SoEF/quYVCWlQHq7FhokH
iFuDs4CGlUXb98iDJJzgaS0pIdrKzlQX+0Q5Oq/bhigTaNLCgAvlQInzSYdcpnykSFzxxdnciI85
As+o1blgzGde1uJID9wyqyZ5BDdB1qDeV8f9RR77CwBoCyuQ5h5iRZunvZeruVjtt6qe7B0n2AkX
IkzxTFfaKWt+K7uG3uLfWKOBptBQ0AJNbmQOBDAP9ZsMrbxlSApjJlRkc8KoDOKzBcNl2HQ6ary1
pdj08duveqyr0cdmOQh56Xfz9uFsUHy4+h/ENpzw7kYQQVAe6gfndF94bHWi6XHleSiDgfszVjoh
zZuTYg5NU9ETKxifsLpM5qF2gu81WLE52JjyfF7iBiWYZ6EIXp+X26FmZdshOZJkZlIjvZqmaoEm
RzUzv2OMLFzkSGMiL5AR3WfLAm62u/6bM9R1o4Nqia7dBfePdgZtAUrBPZQHuJCoKqxNfrSnTt/1
mfm//sH1EKPDo5DyUv3fTh7WdQ0/F7mFeY7qd2pIIEmlSRBgorLK2p2OLnSfN2xdJhSqFu9L8X/i
lU7aZaC22yV9f5BIhNSfmGRPBw3/iVbVV281u3Q60DXZFTmH8CzyJ+cHYu849VhVcpSUymiELGyH
1UAvIVUZV3Osvxch+/FRsgW/Haeee1YDUubJ1mxQXZjardjYmBzMOfCk/nJlEmMMkBn/JY/Mu/+Q
b8JBio8YyaYlFVwqbeF8fT9gQHWUNFbkSteELt3cbxOME1ZA5Obnq4iCoLsKF48J/zaGI146BlwQ
IkPRfXyYDOiW22lb2q6DwO/wF2d3qmPbrhS79XReHqT/h8Gi4v6aAm54XMVh8lczJJKt5ZSCW9rT
5fK2yKs1dy+34Z95gaoa/00v5O0CFWJqGj8TPar7mJcgqSSk+ak3ohRoG15cEUqwiDl2U5ny5ilM
yQYq39HmUWkCOjTFbt9NfxKz3LywUIDSr0SUG6llLRFEUvjf68EfRh+zk19u7fiYw1x87R9qrQhg
62rMzRaFgBNj9AO2wK7E5wL9s/jRhScMaB5OaCRdtB+IqpeS/J45YhK9d4fenGn5ym/JS8AYFAka
c0dQb2hfOagSVcxRW+tl5LS2euJu5dWwANbs8EaNtHE+jEPBr36iFt6eb98/0R8igrpMDlj7kbOG
8SaEMQk+5D8Urxup1yxi+AtMHBMweKbmTC0FYBBCWqDriqzujPLF5t0uz2YFJkGv/iSumVazEGCz
puQQJxe18uUEINGO9AuzGo4xPUEzWqvEZ0Qbe2l4TwydYwCtmLG7i2bZMT3HUA+xhZqVuxPd2BV5
OBN/2xOzR7LkOSDVlIroqTXxuhZod0eH/ejkZsv+ol5yYLlP3WWcJiddetBg8tqT/Tsbmv90tL6Q
Bbym2HX9+meMV3zE55L+hSEpZo7RRZ0bFHql6L6XAM9k37SOxevp5EbeZDHRvH+07CcvkYInNEsx
tT9SheRZ768491F4a5Aupzcvg0BNSZmQarZ1Lb1h282h0+Q7zA4EfSRM6zT4xc5A3XDdpAX5w9JA
VKsrSvEQW4LCO51MxWCCRceiosJLXjYrTH95GhnfnykAw9BKDyc3GgJz2KYf7tZMNiBTZvNz32vn
qFtkZu8Fc7gv25RgjB3Xc+H2vcRkQUBy73c/co5XD7YNg7EAONnUZtItfuMZv4WfLlXk9i8tMA6+
xtfLNfEtptcCUBJ/0vBCff4nJ628O3cHmr/zMPBHz2waaAPB7jWvzw78SwyeQEecM/zZ/a79iBLQ
PV4TjxkUh/+TpeK582nrORv76bxzDyrtsw0JyZUdPgZginsfW/0Yq974shfGNGMy4RaTvyYh1Rhg
pZgY0sY9LZrYD9K1MYieMdCoWYAKXQz3KBHRU3N4OVOIswAiz23L/tJuWP6YZNmXI9d61Tiuwrzb
vBxXeJSqccPGao8uMgO7kcfaOZzhjmWeI434e/mnTC5O3N8ZLg5ir74H4nisEziVLxIhgAyJ9MyA
Byp7m9S/m9ljTpW1ePDn/J4tY5t+z8BhPg5dM2JsCav5JSaydro1tHtt/t6qh7XybdMQB2hTIj/+
NRjWCtwIkxZoEvjSdzd0oF2Dnx1zgBj228eeB8yiojsmYIgybIcrAjtrkbV0swxs0MkfuoEHbJ3f
K0rv+3qM8AdE4nhvp0TxV826bgKIoIYW8/Wou7aA6bXGBWPkMWO+1KxBSOOugdH8xBxaSQdWXORH
3dmgJ1C5hj5F0YGr1jwUa8cCvqaaJS+rxsXtgNcetwO4sKTeSztIWDWmfkk9SjQ6HjXe7z8CRuWL
mlPmP5PAm7gJN7nhxCrvp2BCkNitQAuA9wfjfxcgKc31SegEqIuJcZ4na0Ee+9BjAE6hgCqUN+9j
mc2sQAYzqyF8Z2xfC5OQE7bj5TSO9Qf2q7Bnx/cNaUJv2HM4HZe42Ay8sfXtteA44+wZze86bL+N
Nejs0JTl0C6tX0KslWQkKCfzN5vFbSILoskj7I9Xp3vXjIrHqtYDL3irX+p8j+Cn01TtAWdS0I66
49AJ4IPLuN9zgHf3ORD5Rk5+SGgV7uLfBoNsldZIe16drzRaOBuRjsund5SXZrU+rsdU9o3g5TVW
uNh+M4wpcF8pTgP0wkYtTzjhzbWmuIoXoNLgkUc09BD988KWNA6OH7vLb29qv+WkYqbcx8f7bsbG
hmAJQ6zYAdGyIi8gCofqHq609fnq6PrfsoLoHUq9496+EjZ7KUcG7uCCxvPaTVsaf0kLPdqge+y6
+IUZypWRxC+KX2Xip6nCVka4pguy+14KA0mwBQzzqLM6houkGFhDSZ3RJLzcejcke6iKzez90Vwf
GSowE9jiidmNhsNFqO241une7fxcbOmjxeKj1K765owGcI7RK+7JeGWJzNC6Ynoqqmui4ikypM3F
cNViyTX1fRIHyyD2XwNuwyZzKgkk2NHY+nAE5GY76cW91/ojpzfcfc2sibCtheetle72kPj6jQcw
05T4E9QB8ghzWg/0jFQxZk1mtvIFm2d9X4M44t2Y+/iHo9HCj7m6IWKv6NdqIqp1uWyEXQeZS7NG
TXI+iDsCwpgLXhgL8TmgD3ZC30L5i7RPEBfOTtLKsERBLzYjgajzfOhso476v+/JLcWauSTkscgP
RXwwgS0XneIZ1D0RT6xvWsnUaI/N6/Ptg1CLL+XYVI5pkuODcu0Q/C4Nuonvu7kxjzXubZvzL91Y
+1Y4r8wsAkl4lSXAR9uop0aAFr5g80oq/C7Md7z13I1zQg4scy6hdVEjKAcPkbPGvzbx5iHrQxl+
cvs+OcxBJkHGqm7i2eTmGSJkpPLZk/uj3jn2qjdHt7PPr0hqzibkpGmILd1XYqnDadMC+5fyUpm7
n+MJBFuWK2x67BoMPA3uyB5YR7wZKSOMI1ABZ8TTXiOq6T6LawgQvEXXoZGkHgxJoYO62lGxMaha
p2Gd8+QvdK8meKp42fawhMWgIVKaOFkAz34ObsxXWl4LNju0j4C7VaUngOuCVtJUSAYDVdOUt9vx
vEu+iBpisQXNHbuagQ7A9CzSfmfaEH4VLBA4RQ1c3dpmrl8g4HLvaM4h7AJX1usceYsFj1WZ7n8N
wqd/c2YF962PVpkeLYv34HanQcbU0NySClz61IECiCGQfs/6Pzauffqq5Psif7saLabRebzJhxNo
kSddsyokG3tOMHqORv++RqkMtTS0pLYGHFJ+XGGXQQbZnarnC07pPsTpGCgy+kbVOSh1yfv3GWvv
R4CAckYomJisWqKs3Fu8nJWmaSVUj75s2r13yRyWEkuZNkh9AZrMx6/GHFP7LnlJ6sJf7prFsab7
U2Em2E6Q0xh/xtq3qXFS5QHarkK8u2qJ85kexYi5lvGMq/PZbM0M4csG3AMKk25DW8+X8iUAMGj1
KsskRISEZF1CBbMh5OWdIuOJTbkkRZfltwm4AnI8xP7Y1jJ94wA8nIcg/rItpY2zucj2GqbuNxkK
yLn301mN9+UC4XlC1hxsoxSBA8+L9Ud5SiJ/AX+cOI+y56lbflkdw9Q6cjCvp2kkVwBSK54Q2u9b
d4FCWVmb8R/kxEvLTG0vVSErrv0uvx5QGhj55Pyx1wK5gV5s7hS19PmZVRKienkTZEB/p/H6KR6E
H00c0cerpiwxB4o0IyQzHj31zESdIyRU0gghGFIn/Ezt1Ahz9AHBEPHTPZhtKHn+2RpKdgqJbu7n
cZrpQR820589PwmvvPbSZJoxfgP0jjgBIHmqH4iWuVVg9drSQeHGkT0EwWAka4CdiqIvvoJ/JEpT
g3ldQRw4F26D0WgcsJOvdj7VRtd9iKLPkKUKQ6FR2L6AhrNi+N1dydFRh+iSR6LtJ8iILhP4N3No
pgXtI8g/8WRGiXo9fV3d8lh40a3zhsfBvBN3nDVmD/etVCsmTa4ffdsN8Al6Ar0quP6f9fm/pIgQ
Rim4VlYSzAQ7z1qBzXV4u+dnyOfjEBGbnUpx/GYG+D6p96qAU2T2QFfYssJo/vO7+/5mKjnIWeOt
N2WbmROxjUY85VXjLIEONQAWet4oq2fPiUN0grBA2QTk8/SGRqbu+eWxIWglUvOSfsO/WaAWc1a3
z9+PRV/TGJn4FA23pJvn6JO528+HEzes9zuxmWVuwLDUU+sDNvHm0NpiuevngdHuqRloAy4qPrx0
ihtxnsgKxAFqi4rHJ+BU/aWVlwqtWW+wnJgZXwvFCWHg+jRZZ+/nmUFPeWbfSxiiogMK7sMuGW4X
/7ku94oxJqgCyQgNvCHiPwBW4U9LE7qTIhp4J89ulWXYK3Jm//6jBSPND653504laTXQq2kMhMe6
z0ub4Ue6RRQ9dLurtLHrzUvlsOzjiC0v5G8wzfcRKUyHMu55GRfjhPbHPG8wORhQlIUtewaZQGhr
PwQO+uDAZXAjrojdYv+ID+xNU+e0qw8v4iKTNk5seWoExtoeUaM8jIhxqWbbFCAludwfzn2ipvjf
NoZUXIq4NXs5nqB9RwUaG4YmQbbj8yMMQLj3Faaq5aUU+uzo3Q32t9E0s1pJftwMhwIRFaj2m4c1
XeD6ni4m+90984qvTmHPij8PgdMVH5fwin0go3rma5kRjIRQoaG8C4ou68GCRMt3IHnTyMNaA8So
uLMLTfi56SbAMHaIvhTLg1/ve7NdPNqv9H/j6J5NmlUDxF6xehJgldxxaXNqR7OMe9pynqAYB+U6
BYI/IMhgscXQuJA8HNCxyilIU6ZKIm4MyE4WPxHiF8syl+lAz+wJEKTpEjW3PvDOhhVV/xZGAg61
NDoQC2EoKmaNPP1mRBwLZaV223sl6VwFBkElUNCoF3Jyigrppgh82TPFb+2O7Gr5F+lxYHWbJ/Eo
5iH9cbisE0ai8jU1sqqROAsVF/SkliTn8+0c4f71ZJrDtAz04KMQqemGp/D2uxmrBkJQ2bQEe8SC
7aDsdqtZp58k2791TFt6t0kjdJCL1jVi8OYozLkZ+AUAeQ+XeNW86z36aXeUJ/JXDXKRC3J3eduH
JNor1qKhgdRsLMJcrQ+KOhl8RTTxDWFQXFELdlPtz3rtZT4/P9m6qJEzL1I4AOHQmlvmXoWIB+ME
Cl2u5PS54kli5TAqtPb896zN/bKDSXwkR1kf57mz50z0WlyXXU32bF0LwM2ZVQ6twkK2OYsGIjZI
769MYNofDrb7D8xBeBOS6ei4Fsk5/GYBSFJa8iaC5e6jP2C4Hig08D4spe7yQxZuvmrVAbAJp8qQ
3/VzNOTOH+FXLr60TV55e1MtI8VYamiIGuPq3WvX2J6Y9tQGb0/RzRPOEzo6kdbTYt88sZVNq/01
qmHW29YiUiW5sio8Zgcrqs4SX9S/rL6HWlc7M0Ndo5UI5n+S4kKEfMZwGbGB+wmqzzC3jGWxDLdF
DoGDehQKCOWAyKmpcCRW5ZgaPDBd7B49ay3kyS498+eBwd4Nsy9tM/okfsSqEUO7peXDobPW4hK6
qHoYVPnEktG1SzF/if0aEnqBgEZZlOUqms7W+N3AxS60rqC7gKAQt12wuJLEstgcziQBma0SFzlx
X/Al4Je+oBBkx52kRQ7sErJrgt0sEXskd9SJ35KhaiOOmENFoK56CcJWbJmDn5b4DMsT2C1XRF1j
F/WuRi2+5hh3+/a/4hkSobw+qEeM+87wgjE2Pce4JNq/xmAJvZ9aLjN5KQ9oa9fwGDHvx+WAngwy
uEX5WFZXKIpFv/iwy2yjfkLPklzspHCQW4487MyT/DnWzw4TTRyfMUgzh7jUsNkJpl/DGlNWCmwt
6Ut4MHqAUoPglfG7ImD2q5bDXOUNKwlGJNPXqEg3j6O/BZw728ddyKacbYbBjcvZjSIK4cVn/NF5
W3WanLGAvYNhknXDZ9H75kTS3dkFsrIsnHu7e4nDbge3BoBAgNzOtoM6R2WLljbKfqHPfG6F+7bK
IlYtZA937CFE3mqTAiSUT861Yui3K0CoEIbLxr4diLf0OSo5WnMDmeN2MqlL2WTjUyooHmQ0q+ju
d/OA0yMUDdCY3yVKixYw0J2JqWaNDjzkv5wf7PP9h91mGuVnTBTEa6ArqeWfBZ1gl/pFLlAqW/JY
ngKBADZfYp6FqHmzUZckjyoA8nJoPvdhLlFpKvrpnjq5thYo/UVZR02PJIm3Ndl6pTyMvcQiYEDd
YFWS1mv2jMJOMfwIdJjMibXsQXLlGjyOOCqmN0VEzq1hrD6d5OoItAuWuCC1QLYWRfypb8fVA6/P
rcSGdkNo2knX+s41Bn9ygdMohHm1FmqRu1/tsqalE75OPOsSbrzO9cQA5QpC/61tLafW5fWM0TBk
6lYLqU57n5zks/+BSuD2QT6Hc4fMFuI0QzTt9vQQF799tY3UIHfxacieD/WC3OZxPzAYZKMD6QFm
ZurEg/vEW8i0nugm10xTGpOTVbeQ2MzCUIiCkLebsjCMRydUATNBTyX6P97gHQV7+6BwfD/pAECN
BRYlSjLBeLVCURncnSvp5cyjEnpY+r1lEv7QnECJ7HIb2RNARiESipaT8SoFE2Z4fPbV+ZyVKK+Q
YNZjaNcufRvHx63p3ndqZgXlf/9k4idxaBI1TbIoL2FAU6Zm1gyw8jmJvipQDyo1zU5/Yrq3TFkm
W4jr7aAoTiui43WfIeVmHnW0c18MQ4zsPLpkmi3teqln+JJ3jOkBQDnG//qYM4aki5yO7H/1AmKl
JWA+AXJXWwjMdiSi9iVGtUOvS1oP+0kyhlTbvjsU13qtXmShnwfZoBuzqyKz78cOV8nclUdSwljL
yf/XBXcntBYEcGxHGdNXDvdWagSK+GB+VTiw9kqtprhOPhS8/fEbQMZ0HbpeC9g5EP+nt5ZXkrCQ
fPDmpNWkyNop8iGNmtGUoVnFNPB94hkry8mi7xbKubCWQGa4Esal1mx6Oa13AtDn+v9uFhR/VUsF
+Pkopo9Bz76gh/WjRMJTvthtkxUttJwSswH8fDeqekUaMcVwdGTq7KacRcrKxkgW3Cy2R65zYA+Y
GrAEfB/qNWJjDbyQybpbSkiX/mrojWFI+3NoMqS4c5it3WA4ZzSsvw67hsZqACWk8okrgEB1eqZ0
LrV55f/3VCH5t/F4kWU1vrH7sttgN96LoGdZgs9X79ikISLV+M/7rCxCO7IilA3UJEVbP9czBxgN
eJLwcUESJEm3vG//xvULXDrjHJXm6mVCP4Kd5xsxVp6kdyj+Ujkrn26qKt/ywTP5H4mkUYcwnUWq
V0YJUUsgawPtp3ANjqQq00Qw5kK4gs43AbwCTAVIHXKKelY20dVhBBjRJWlMb6WdJomovBNu/k7w
2d7RqXjkOOfEyW/qIVSck8V2NELrEo3kzDZsVhzSSIofoCAF3ubx3ljvZYb41i/heNXZ5IFBOVac
w8oPEBzq4g9AIEpVC7wUiKK1tTcFE4BmSEeFk5BxjgV0IlqWDijtaxKxWCYNdr8m9i9TagQuTzuC
JbECTO/bO5mPBjkoBLYBVGBuecO202bP6JUji0urxw/iv6lhhUpuf/jUv+mSwRnfB8vGXkIILPzo
Vnplikc/fubSH8jlaeuIqt5czsWxgYRws3OQYVnd362G+Mva9+nqxMMhyEgSVczQJ9QCWvl4whH8
04eseiun5Ww0f4bOT6m4wwG40lg5ZySD0eH8bTBTctKBAsJW04RJohtVA175pUtttUdR0I1iKjFz
ejBD3GwhlxvOjhyKp0Zlg1Ao/09RAQ8wLRRH8twVMgjnxiwxHXRC+5uUD9z0QKTzFhFYaypwqR5o
YOV4cUMOShFBZqZvjsct4/pFA/CsIJqm7AU5GbIgUA/lvgY77NEmCTib5KyFnc0/uRSOD/9LedUO
mnt/DX/Sq5PovBMRPn/E0ePyqwn2wDBkjPQAB6WV6UItjWQikir/t1pi4SaKBVbV+NBeQ1E8KH7d
AfTiMP5HeM9hhBzaTzS3UbVts6JqHYm7shjpSP5oUTqmtB+eT4V47vzJiCsO/GDPXQ9P0QRDW83N
kcMuxGCWsTVNjDxALlQH0s+N/P7FBTPIjnX8oz3r1+qQ/rZ+4gOHl4ktt04QVqIXV5AL9qyQ61Py
MeXCrNeWdLmcqf4ycXneMTG7Afsb+CgjRrDRSdf5MVGWpfOGBCh+FObwNfuZCotbOEbTOJheEd6v
PDJkKd3wkFgoJOf3pUdjarDLpvA84C+AsIcqYiYO3ys+4qMJm8zGp1w1Pw7/ef6xMDr4fndLJkQV
UYmeF9d1El2DH0rDtMPKCz7V73SLQZzC1SdL61DjudMVaViKeqXIr5jDK/PqLLqrEK9WNCsvCmMQ
uzk13P7hg9JEwdB9KL2DY3U9AuRSuobbUr67DFcIuoTXMZ8vbZYFQ5D/lVM5LnTIkwhyH7TEKpGR
rF1kzZ13VmGsB7RHBxcYV0LV2W8uuOeJC+0iaOiNR98mGulv+G/WLJ7yqAE21GUHk0SZhcxNuEnH
ElPfBW4pMeZfOmHI09/8SL2JeRRnCt6dQUOPHTyaazu+E7pp0mi+Q5hfrnlupgzkXGN1pV0vw+2R
QO6ArG3Tjw3FE5DOm6NqwJBUAc7v1WlnSKcb2mR9ON9B6EoaW9k6VXgY7epAUm8jG8r1rGX1NLy4
eEyC3z7VI7ah53FuPL6eLZy4hrJmbQ26A6nHcbnx+BjVYJGt3Vd30ziL/B8O8oNZjYpqoWGtjurm
St5jF1I8puxjICUbZUT8K9Fp0FxZskUsrJsdFejbBbooAPDjY0u2J5Gqu/IshY/8UiKlsLlXsq6a
7KBr+1g9K95pQepZgcbk+eAtBPk/k5S/3M1iGongi0O2F9Aosq/hfCBs+mrcXvlgguR8aAY8RoxO
bFgGqoHIYQt1abxpym9MALKIlrLgoJpbja0gcSBY6UdtGRQzQ/IO1bcufhRvCMW/0KfWTe6ykkHW
1hZoEEqXNLL2qIScUOroHXhtt+KLIO6h0wP4MCpPJKpqbJY992XewULjVIG3vOwGULsepiA00M28
O+C3ItMWPihUkCY4XpBMIO8r5T4GrlgwPAkJDURGKYYBFXtwPFdcSExOXhmYNrFexEvO4xMJvRb6
x94VDjG36NE+V0W71RDl6L2HCi9VwDH5tcwsqzzF9Y5YKNhPzE3CdJ2cXFb9K5nfw4cuGFZYHB8i
pDFjBS2g0jl7EOS3Yy0K791DjBdFssjPhkZGPgAcBDxj+QB5qZkDKv7ya6QCIar3ibAmOPJqAb1a
mZD9MXS5F13hErEdfPwV72N84emn7zuvbscBzMWt8AtU023782ekpp+geVabuVR9DCL7hSe/pPsY
c7WgTm1YeWP4kPhvapJu6mZ2NdGGM6TjFa91dqN+KUw59oFMZhvIwvZqg4pyujNFXBIOFbScL3AY
P6TrywXp5RXt0NLcKl1rFDLH52k+wdr/gQxNRTNvGOCFL8ait3jo/PBxIMsl8huwCEOSJRivV5Wl
l5fyxkXSe/VhuVNni8FsGOMeiP121Kerbb4c82QDDsQgJcmMmi16tZ+3PTr7f5vLGb4pRAmkR3Qd
mt7f8XKRqxetQ5aK98/FVagouTz4RR36ZFiiYaOZpEc7wyZC1JRbHyXzoN2UKRAPuNKfBi5kORwm
rypAiDRxmN2+qBm3GoHcNhg0HGmNJ1OfLkAi5ha5tfgOYHUdfhNeMNvcOBLYobWJ4ti5SstTY8tt
UE7G2MNYcHjDjQkGYcmHRJZonWKzwiebx5tNWz6oo23kVOAs+JxmvlQkpBshzVgD2S6P+JeDK858
wQFwsRc05HfM9ukmZ2s8iyF2459vPRVzo0UYy4S2QOSgf6WWgyMMFUNbermkRSQSDoMLLi5NlMZh
3gYYDnOTs0zaa8MkSovdw3XnCdnydD2qulSS6nhf2/iOQAhaWXjbv0r5rDrhocO/9b3wvB5ZwN0i
I4E9nNUuHjU50Y5H1lGYCpNTnMuQSBvc6olFntVER2HIKiWpVdalzqKsGsj9FXf9/UTwN4FHhWdJ
xRA8xWOoH2jXbRz2bXlgkcfx2K4e7kVPMzwvnE+GGKE84H+0YYUfR9cpB6sKutQBtHFWIxrZAUo1
SbGJBmZG4MuzpSpoopQpffihwQ2T944ynFi6B2PCdYZB68/NTFgnLwy20x6LTM3y24Qleo+l3CNn
LYLUdpMs6LTLnVWpD57cEaJMMx2GZYQxibEU4lm62uClpkrGPN28XovsWuzmvsAqND65rVKcDNsc
eKiFHoI7m50DfBdHfWJBlGMtcEiLGDUu8ticLD6URjQmYQ21eR6aTK1UWjobaiIGOwnmdNKFzmLF
cl+LSjb59VkwJroKUJ9Y4Uz5TXmV8x/ZIWlJSRPPo7Vih1WlUO1ZdXj9BTQXaeALNgpYL2Sc7/sE
jgSvETKh8CZClGbmuY/st9yb+iuqmlM0PRrBZ3jrEjt9aDei3GFUnaXwaBMs8nZw+y48udJ/99wj
yM1PcUuwwrdMLLh/IcTi0eZWJmu9W49ETDLehWeLsnXhVqafM0Aduq8QsHfv3sduGOqFOtNsppXU
dWta0rcwtOxJq8vg7fK3ZFITP3Ngdrwyo6KkzTn7DuyFpb1vQfdg0qFFJX/Z0/cjiS/5RDFaI6qu
haY2v/2P7ocLGsaCnO5CTHCDINrGIFrLlPgGWAsBZ8nwqEmnu/P4Il6t7qfl5aibJp2Ut/8w9lmC
ACFA/+XSTXQrBGOiRKD7XTI/N1By0Dvnc5uuKX5rqfE/8ME1nuxwx4TcPNipPK7wNglZo3IyZOGi
ntyyrjwO8pE+XhpYBxxQ3ObmypoVHHYw2MJgIjCwORr2t5FaTnCn9MF/m3ka1/75mwRmzNM7ZJTj
hq50Ub+UZyIUyOrPYIXE/T1VyFGarEr1rHGuThY6A/xrL3I2uPZ2Ik3m3kDnXeWNEEi1bsfQSMI7
gAWHnRfQ+VjtxXohhBud0Tqv1AVTKOPrr3oPEL1xwcsCP3ulCSQnGs7F7HyNeNHX4BbMZPEfSjwB
OyL+lzGLCpcxiWeKWqnoP3BIeRXn0/ro5HkJVELBNE2vJi1oLYzloWBhRfh5VMm42iq+nOxvbLt8
HWITam97FohVL7MjbcTZOCLJfwB9qU80DKk+/P3NfS5+lg0YefejvipWuydFliwZUhqp2IFnM2QG
AUJzoXpykIsdjCVpVEf4fkBrVda3Jz9PYGtkT40b7t3VW1hEdpWiGLzH6xBGn6Acerc3jc7lrKfv
UBMgtTxQvUegI/ii10csHdm+4bzgKldM9VoOgvsUh2aEnuFd1P2YY8/UzM8OU9oEkl89N5I3ztIP
vOfy7/lQlnE6RdGz/zwOPIK6KM5zqPc7mkVTWNdMk6HZti+70SEVdxLLimIo5SAdYIyKlgkR9lLq
Blcx+0NztMtSQJ4jmv9KY4d0fB3QENeB8ehi7PVxQGwUJQIaWd9+T74e6zW5uCvKpbSP2HGFu56g
VCd5fb5GF91SUVpM0PdhrdnSM8Z61V09O32U1ryNKP68M7jVPyAyst0uSKaUB3XecjVnwob4GmW8
jpW/HK0G0TbF3fC49VNphCpvJLUDxGwtb7MCshcXIYWZyQmtyGr37ClvE1aKCzPNVGulDHXAq+EQ
XV72osx2orTXxINtMqJZYOiLEmuiZcuyfmhLBgyrNbz+zuvXct5GUbuRLlDcoYWd+/rBWP/MgF8P
ZE+6AtW7QFOrSxy1nYbTzYKtLvLNG1zSCGz9eaIHoxqDd37dUPuqHjdSjN+Y1+ULsyixbiHPY0zc
NIazNQOy/HsOK9KexClOUFR4UgMzhrkfUEbLLDHHGnCvNpNND4QmvV8sHRbrrnBdZnHr0M6FrjPB
vSXU+P+tUpdncvmNo7OTrfB850UlYSvmQGSayfUTereuKDv3U+eyTOvR+Bx4DYqYaFavUkyycHff
+zEgk042AlRXpA0X8zb2pduvZHdbmGNRQRlpAWSRc4MPz2gyY7Qh1/uegIWay7OTjO/+VOcnSWCU
1gzD4eUfaDeuVzFEQtHvCx7oesJi/YzNppVATRBsET4KDYcV+5pyt29y8sY6z9Za8SFB0+ZzxFRh
mFXXS5Hh4XzwQ43x1IQKA5W0o2tuWW0eRnOtpqqq55rxyhWvB1fNNuB6yrBMjdzL9Ny8U8gQmsQ9
swO4ZFksA0gTh7idGP9vuTGvQfmq5nDqwgjg6B9Wetus/W9ZVvJUCtTyq59o7lsXW7WPfnxsjzvh
KEoM44pE/lHinXeigxH+mFIYlgI4zupc9A6fB3qIbetaJZV8w6LHVvCM3ypuj+mmt7m3/N6LyGAf
faJmXBTv9keP2ISXeC3NgFHWjR/B9VTuEJhxdo2rUjRHBvnrf+KrTncdbQARzzuRSHVdtdufwew9
3UPWTjURzeBmqljELgdq9GSdZjb9wJZZbjVFMXMNCar5xlnqGpPfTRmnBvsiutmCUcjG8eK4H8Rr
84UEST+3U7IklcTHPOsTQnUBTNjSB5QclRTwyT/H7R6y/2QEX7iBKUS5eSeLltFXJnZWN4man9eN
nSZKgyo4UtJyq1Oi0SN9qqYnYix1g0CzcmLgoniMurQzWCXKWxCaVa0xIJNxcCsnZKagzviVICFF
Vj30gZHEoRTBtG5clXvGkS+7nG2a/z8rc72D2g/KXDR47453L/iKMcj2EcfVZszebPN4oYt6WrWp
ErQgSWj3+4AH4B2K1tB3EW4nsZaDeG1PPMuLDh58Kjxv0gOurl0IGEAnoDS/BWo2RZ51ZbZfPAU5
vpN8EHjUKwzhp2ETkTpY+oRU0ceBUx+qT10G1lsXg4/6imv4cjwzqpoMlOLSLPaO//0tNrNLnk8R
Mf/RRNJKPxv0ieDMgdadbK0i7J4jP9Ll1fT8EuoV0RYYInm6XjYqX4pz2PpkB88/LmN2b3xmZEld
1XdCbqOkOa9k7i/Mm/b+b9mzVlq9eaYtQ1GPjyRl8sAWtVvoGiCn1VmjSjFpISRz1D/POv5bzoEw
gH++V4JOV9pZt6/tutSkTq0VN+wn5A9EtIE8bWEsSZaKN9h1R8sHX0u2n0vzBJSSA/ENWqRix82u
QQT5gVh4V2Bhqau4QXYP/bhQcc6Fj3KVyXajL9jjSSNhVikZZjv/NhANWbmqJWNiORYeXiBtdjTd
uK8J8sQTUbLbc6D02IfoO0hq/cMq2LVwKbZPeGcG+1+9c0uQyr5w7Zloy7mtX/VYhLUnIlbjImt8
jXOOuX2VqmxnTrPxFmnG9jqrokoRZhPgcVq1JSAFyTdUFVvEq2uyB13Fg+c+mm5seQT1ijWpKolx
nNmXKhgRGc5XsjU7Dv/AEQ3q/gsj+9SYQnxUQddOaDNm7ZbA4oCYmasyxzckm4m10AncZ736IUdU
ki+SJ4VkgE7pOEEbYtcAtHIZZBYQBVO+9Tc2SjtjbfvduTfKcCYdBnKEkOdcOBt2FFwYnbkGxHiT
oILcRA9UsJWi/JdM5oVnTOiWykznmUv8T5Fw0dNmq7fvFYPRG86Xm0UNzFAq0ZU5VWuXiPKP27P/
qgSiKdacRm/4agTVWMzwp0yCi97b6E3r6frcaHh/31yZqvQYQoesaDVL6CHknPu9uqhASk11J6uK
U5qxE6bw59UnyakafwhfhRZNxyShHBybNIQsmE5M3YUKah/iMy9zsCvQZFGLDa29fiq2KvQeyhKU
4Lwkxo8AqAzYB0hGJWNfhQ7ENPW/mxTIllufH8ScwbCEd4flytM+mCxRh1T8tPB2MOOLQ3OX9Cei
7CpcbKYpigLrQhcyvbJPkNzM+yATFNhwsrDIAoaP6olQSmRk7Xz07QUHqbex/6gn81jk1z5NtGd3
y3ofxjIBTZffl1rU29Chk9zNzMgwe7he/nFtv9tl3Sdg+knj0ccOLLDy4qFkQtuRMBDdCxiwvwke
FKCZ46bbeYG10IYqBf/RRkQW1B3vSq+iph1ND7l9koh+2bPLh2XwxcmvKBTVIbMszkgd9Y/j9JON
Vgh5h9hdRi+gOsZVuJ9j+IBjMrnDLag6uj82BA4h1sEt2gVkS8wn4bkt1EVhnn+bGw8CALk9BfBo
pNyX1DuY1ab45wtKVVlHfrjuqTFDhuNT12rFWNVtrWFTsJTccnkcvYiJ0BvkFm1iZpPCYe23qncG
10k/HyXUKvieKJSp5XgvrPix2CBcRmK6378RK2g5hMMVdWKsE3xE3BDIfhel62geGYOAQJEcdRWe
zX9Hr1qPz+G1bkNlnCqBX86EmjBUDrejaIanfriDe6YKU1NAkKu6NSLpzEonq0sEyAJwn+zSjw9t
/PzQhmZvvbHagfRJDd54BwJ5DZZI7gfhp0wQiArmvG6xfb4zh+yFyVIO0iUMpvsGYImTOOUuXM33
NNufVQo3LMWE3YvFUwRJxNxEONJvujoFUJiblDpReac8wmuzRFKPS3xjNcTvFjFsMOzC6HixW5ey
uT04X6sJ3ojnCosE4xDd5IzrXJDAb64ehHvczfexW2Y1jbXP82C22YVVAnZNSH5ze0wEX5XrXrzH
A+g48EgVzIZqJ169je0fBfoboU2fds8hveq7wAL/QYYpdOWdgEInfmT5NEfMG5u8y0pLJQDsh26F
ayQDqCS7VRcLjXyzA9/Z+eIw6IZUZpD1emMmh14CZU5xvnb2lfiK41W8RtUl4EK4ALA+H0up93yh
PCwdmMkTlnobmofhNTMv512flOVPUHMxxkoq2BxHaAcCvH3s1p7nmOocvDopptB8ICw1YTT/H0BO
I8U5X2DOn4GHtt5Bn/cYIszHwlZyigfEGHlh4GhFJTJdjbuRu+cUGDCSvWqSY7RPLskG4ey2XKfc
bXpcImz49hNBuOdMCGb/5m3KXbae09KNyS+vsZWKF8/ljQKwVuf41FdzTvhohFdeVqQXlvE/U3nk
OwGcP1su6+o8ounbYR3EmZFkMOsH4MgCvxCa4Hy3eOXjNn8IwRrU8g12DL6R3nIgpwmcWWw1nrfV
4AzIxDwNKiXTEjalH/Z0fm1OUXZmXn0JHopaaiiIDLZo1FhsD47M2Ymv9IhDzObfbbCcnLWDpb0S
9wF+8WJgEqOwBgkl6jG/pGGzIkZmmOBDhhZd7jEK4Ob71cPDMaDNlJdIwzEVybGot+XIiP+Yp3rk
WL7N9PIG/tY0YAyTUukNhvCXtSnDjQsoPLKbt+DfMB6Fiduv46Zp/w2Z1/FFZS4dYcDcOpjv++9s
BxDwXS1LUdPNX7mGPJPGdh/Hp5QfFxN+4nMmprb0cD/cgQf3xkXifl5+yBApzfk2aR6jDZoIUVkv
hWlWjPXS5NwE2rtisOtQbfu0n5EQWbMwC20UnH5bZkHq/ZEVYr3xI6cF36WKiGNrpKEyrs/VLoTN
Vht+6M9X3tiuBHWRXXZ9YLxMqTTDlr9UJEZxh0yxelOcScfJFxzAh/yaBZBzqC6kN2VSqItkzt6G
22/0Aa58MQnngs5oJ5kNs66aZBjWLdbI+QJs5lwacGdszUcVQ49qcQgNTzn0OnQVemrFAiV1qKtv
7BaIYkcxA3PV+KdiDYlmVt7566MxVUkDdwqlG77YzD4jafCymIQRzOJWVm/FkuXC/auTR3JDUi0S
Vlsj9jAqXZQm3f40kwDg40ylwC6zAUS8xWKaRKYQSqDVKpKM0YmrAfit0T5hENYdLM6+8kNZAz89
gVk1Fc11bpN4T/MYxqkK25F/qqudhXIe1aV2GQDaIK01OprnK4aUxO9huF/L6GKbW/yR2vAcIKhA
fNCJNqpSn1I4i+kd5YqajpcVSW0OO/9E46vxPuMicFh5qtL4U+9CpEdBbXThiI9P3JJ4SU8gWN0M
4x0cO6HifBz/Tqz6h7dSUFV7SsqlrkWek4M3s8ig9RA1boViAlFWUUF4EDZLBvlm6zQ4Lw8F21S8
rNuuIg7VCNXjgH6Emr42yUTYl80+9z3GclzVKRVXmB7S+KUoIZgqdC19G4gMBO88ppObpeqliPFg
bhHcB3bjO9rlrhTGT8NZ9GccoZ44DVA7FX3TrnoHe9EBlfY3WWgM/sVEJPxcAnWsp9Y5bixxaHMZ
vMzxY3e56R6iCm83adgFlTYn1mIid6MAyo8dyzDTQwjOm9XfSkz+kyUdap2d+ASYKlHJUimONr4p
8Q8OGTXtDzmeB7EgzWq/YMn/OhiqjZmECXQmUVzEMtL6NWTUkHM2q2hV3lOuL7x19RJ99boRbQXJ
p2JgCa6N6RhvmbK1npuhPWU3vvK7KQ+g3Lwb4r/LHLukYrfO8cYsSuGdez0cAXhC/48oAKDI3TP6
m0JSLpcDG0DBS2syFw7a6GgtS3E1RLEEkJUAr/Kvp4Cp5FcZgwNzVtBHBK14MXyeofyNB7ev8wkN
9QRSsF/L8HsvqRIljXfzWvv2BxsaZ3OwW2kstSfykdfjjKPhqk8oa4n8L2jYzxofr5PBO87n5JBv
6SHKhKlIAvFOFW8jbva2BUnqKi3zTAVh3z9G/G5QtJ9u21KHXLIvKowy5EvuPgaxqd3SN9cfvxWx
mGBykVsramSEoJx3Lp/2ezyy/T2B5cp5ogkdwQ5PtmfRU+2dZLg/NBM2ml+xXKFOfrCSRiWlSVFB
LAJqpsMxLWumwLIMd89Zi/wIwnM7zDNx1/cne/A054kCclm9X0q0Y7gWpzGeUAzGcXomZ3T3FfYM
gOzurHM7eu/p2NvvGOWFJ7Ms2/AJeSwnkuOmPJA5DYQ8t0zcw1yCrnPZa/TdGRnm10z3fVkZ2A0R
QF56xIEsVso2dYuBbniBFXKLOHoXxNY1Ii3oWcf9H1qXWM6aeScj+lJZAW8HkSmaWkeEsiXB/FQh
Nr8VUkh+m7HZk2M5edRGa22HxTh8FZuD+c9BaUKH87HZGQv/Y1+MqJH3mXhLbK3CAm4fmOfwjgl4
puGtatPkouA1hoGl1+TjijazD05KKHkkEFJhZPLe4J4kWHO3KY/zgVaTnN0CzwyH6r/UDwuHs86m
DoALCeiNzn/a367+Nv86TnHEfY2z+TjdcJIBUMizRoJIUgcNup+kUGqBspQl+FMljdXJ5xTJHmzf
s1Y391MI/HUZYSq8AdJlJJSLDmOrGzvngwKlm9+KqZJerz3dusLtEm0SmW9KGVglZxCGfJNNkJUY
DrEcnXEnLPfsqu9m1ygnr7ADFDVwllHMc85UaXo1ECooiKp9Cuye5tAheiEqe4YCIAK3UIE1kwuw
KLZc78K32XSzZqszxWev+JgOZkbLTl0UZcdAwEnbwqntupvImoXbEQGRPvPujgFZrpGhCCGksg0T
7cKKLcUBIFj6kXDHv9ErGZtv3G6D/KYtXV2zlJg1kQwLR7vP25DULFLm8dDtixLA2LT/NoenS5V8
h0oXw0uQbE8AbwZxK+TXbKdEoWNVkBQPhtiTEQIA1RpljheDSXSy7cJ5GLbwsHw9BoOethqcrq+1
keoY1eqbX0gT/9S1UuW3xliglfT7g+CoW6DkFWV+cKkNbKk7pQBktIxSg4JqbPqGU8Pqhi+oyND7
UcTet9rxrvLoxCsMiQsWRyj0xETbSZJVDFGiJb27FaLQPFhsmZr9USwhAF8CD8enFc9UyOQWnNcp
2HvLaL8Snjx2RFsVKbqWQyNXgsKKYTJojPpcP13OFzyVD58DMYlVKrosDDBN+lG50ccz5pu/2DbE
qjoAZK+q68th/cIt/YH+ELxP2V9KjBuIL1iw1Oj/o2yCOrZfQ4cfNTLEoX2VwUYG0aGJEcJAWGqV
VZ9fNZI/fKDgu1OdOYaLZBp+Dv6eF0/zftf6KtyqS+WCEfHYrGIWRY6Vd8c0RVkcQBKP38HyYevM
FvEtF0yDaSu/yiIc1B4/RwnHIN04k/Mcp9lYm4oNVkrgpysDFHjmLcSMAjH6Qz/zEijioEaSTPbx
N4O6uG6r5yLyZafUZy2A5iaKrG5hdMkoIHNcDOtX8t9R3sz6x4ed5ksYHwlkcb56jlE5wPW/9Gi0
N/1E677EcaFbimobnEz6KM9eIoY37gFWy7Qp6T9SoMlyXMFuTJd1CtifkaxYCG9DswqlrBB+l42O
lUj+gVV4bkPr+hmBoNRR8Mg8b6Fp+8JnUUOCr7SxAYkREHP8ByUhtGKMIKz5LQwtriJof33Lk+Ie
+E83jw4HvYdiAHxzRoLHCF4RjhQGjwt+RG8lXpNPGYSGpArIFBFZ+bsboP9AnZiW1ooZfgLbG1V+
HfGKrxkeg6u7OgvEUAabArdaWXwtdrl43vUlqOyOC0tcvmBxA/i93OVaHkp6iDSQeO6zxomJuZp1
hflnX1BxYsCSuaT3RTyDNBoXn5uL8Q0xfXI2FbQTPPkOjaTmjl+hUhfl4Snwx5x/Ouqv3srRWlGB
Jwf/vocw8qAvxYYuA2A1CgFaKdJSYV41VeqeNgigboQgPB3WDJxvcsd87yX3xT9Kws7mH3KyKOk1
kkFHZICRXKcgVc+p3BN0u1vENITCwFkj64o71KY2sfHJMjYrtcKnN/jrxvr9egXeX5Kb/n+5lfcb
WfcmRG4kWh/02G3zxyfGVtxN88lJTl7XDiB+QS12kt2BggkCmwtLJPJzxtXBK78hQcAdmv3mFUeZ
GgCabRHoWyUjhnW+9m1Ob6hkq0nwVCY2tC8RUNvQdmK5wn0THPfCrBFX1i7NwPqCPykzRIMDN2qx
lULlW5EQMcGNEfjFTq7Co66IkMREfUUZNWeTU0L7wbJ/y5hMxN+mnY+9+7krFTPy0Ck4NHPfQ7OL
DXDrv5GyCYD4a8NWh0+f4jYW8t2wviSIdMzrG4R3afDmmEmNnI4lEcsHjcY6LYv/fszo1kKnQrnb
UzCXJJHgodwu0KODQfVb3YJOjtqKtkhOssY028iIisTqjrCurqDhOiDpw3WgRXBEteRoSWlHdZdP
ZAtNIF1Saq7LM73yg7OA8ofk5EI4sYOvFFAlRwKGSb9LYRc9b3rXBRYPBoPSAQl3/8bllewoLD9X
0aSnXkx7PkRZChCleJhOxQHReuZaNSMEyd4lCMOY1bhy8B4gTmIel5YLGTn5lx4hnvPSKs588Bpg
BaRTT1fdFsLwbrXIYaYhZIYOjVRKHom/tWo1rBsu9W7YYna4Il/snQAuzxwL6EG7W3Xkf3VRSKVT
Tm15pdbFvnfo9lEmn3npT+P8lkUbEqvrEffRDbEd1gZ2mSfhP91KXKmV/rrop+Vc4HVuNBovdoxl
3NgloxRDvmoSHgSaHmwwiPOES8JiWyX+10SR+xCC1x3PDpmwax8gfhOg/6CRKWHsZC6jk6j++lF+
ABNKKrTi5NJrB13oIombgKSj7XKOuOB8zIDv2O25Q44w38Lz4qDLpDqsUn/x7zU+P9fWMc4Gp1mY
p+YSddXbxVxVyrYpauydQ8UWTi6Sl62cZ63KuvK9ZRQBiTSloKI4coR6GsMfRoway3NXScmPpswO
5RSc8tb2t1t/KclEHuOQDbKZ9vOa0oCwQ7aBNm5A9L3guACp/AyZLPbXK+sLU7xscVJt3Dy3A0Kk
uc1nSN+yrWd4Ic2XmgaTRls6eZ58KZOLjrvNINqbiZF3UAWx1fnc/jJ4uZWbJTs+iq1xtfoiwDzW
+lBaOsXjXxwRdxZm3Lalg7siLJ41a2i7tqVb301HegLx1qHo6yuzQol4XFHTdFOc962CLWi0X0q9
sHArrm8710wzVWAaXZmwfgYpIuhNIfizzOY7wWw6IyMj/pIJ1Q93QVH/xSTsiFmrEu631WRcHTbH
wTWJV7WUB9xuiS9VL45UZ/BM8nR+Jvj+jkwA18BCoj89kAArtbA8Iqp6V+HJKIPFcv3kLJc+0gwg
nsR2LQF2OGGQm8TAJee9EYDo7r6KGtsT7AeFWZSLv/RexlM0BCogDaS47inBueW6I3HEjSH5qejw
WGEP/68yqXFsSZ+ajtQQYf3pa38e+gA6ejvwpbxI/FZp3UgRN9oWRyoeI7VkCgjuQAVedcuYn29T
7tffyYp1G5X1nHPD/WHIRBi2zJZvULRRBtdRWj8/r0HZYQfdY/XB+EMkPBUKgpwHvuBK2iU0/Pi0
rHU5HGKyBQjEj3tE+AdhQVvOuTfUC+5i7s5XUwHEXdhnosc3YVu4E5vajSmHjvoAPphMjggZwNoR
EdQb/FmCGLyWpEjelCnabu8lK0qbYCvnZUk6JB85QPs1a1dQup3z6J1RsOKHLpYBrJ/E5ZKYuvl2
ZGFrUX4NkOO8wI4lFzTo6D0XGUKnj+242xQgOkYFxiUl6LTLr4F/prWRupOAHqUbJqzWy+rBd3qg
QhKEUjyZByvun5xo6MJK5RJ0vgn04ZtfdTQEZLZsKTgQqi7TwsEbMOQzljqHcN1uGihEoHI9eit8
KlQ79L884rW0ucqofq3DouMwawav6E6txXoPRBrgPxJv2AxQyJD8JsGeIzsrfhI8uBC3f7sy2mAz
pE3Qr9rJ/4kKcTZFWCY5kuq4+jg6eMnbF2YtcWFplSaAJ/rRl1V1NDG7UUxGYADYHZP8p2M+FDCx
u/STtaBzxGdQsgCAWVy1Yp6qiVIeKnlnfyLKX/RY8KipZGAV9uyv635AeyykUBUsV70m2t0NAHFl
avefiJUaFvB5oRTsUmkk6rmqSX8OtfaXdE50p5biIPOgCqF13kgwU4L0mYd/azMbZCMyeco76Gr3
iFuseBc1ebduPEvwZ6eAddpk4+kFv0HuAesdwXeVUwF3vWzUP5Q6CAEwosxpNRe4cqPjAlltB5+n
Ltm2T2YKF+v9Q0QcNFyTYpm/2VjtmP0WKnlvhfzqb+kRokieJHi3HSfV0bSKTvv7e2IN28845Qo/
Uwp37vGspE44l11BkfYoXpfbC3B2Jcr3OyFwf/On7GgEMusDAAasRP8SaDUCui9mYnsMw9HRL+KJ
eKWCrrgUDJ/ULX5WJwOdiDLErqp6u/z0rKpHtjAx3xb+owfSQi+JBkzOFgFbLoSpt2P3GFS0iJjK
8lkX/TBsFUN6JeFIrCm3G14SBA7zOyk03VgKfmhbDReiImVfyO0rBLkzyXTBrMFTdeu9CS0oBk+Q
8tINhU3hF+HYZjvW2xETTvKvqK4xR+3iLzX4toLiLUxkSG49n9mgeDbpor27rGyBnHTJyr2/qyNI
x9ltldnSCeKoDLQ3DRQznIxdwmC0hzlPb++F6uRCKdw6bQfwSkqgMg208TgkSHUERWI8aCEtTwJC
e382RJZkc0dkY8kRx1kh0GByWEyp8wnpAoFwm1uz6vyaOQVN/iublm8J/80YYY/3qBduMvxuHJep
f6a9Avf63+Y7w2N9D/B6IT+KcREeVvRz54M2IJRKPCguSK7F9K3cfzYEWgqiZZTkMp7ljdVsqbpQ
mTZMwwEIMDqx8FeIwfnO2n3XJ1167orDWTG1A+xHpxtRzjEmx+I7P9bTzco2e2KSpqxZfF1fYNVq
dMMNsH60U4J9igwPGkrDZBtCq8xnwDkdEn2QeaNu/FirM0DXohRTpN0sJE1wTOtyALdXPJdfMNGB
fFFrlEGxx4IIoFRZw75RPDaikL2IO+AhJlgJSj/zl5yiwUkMiqq/jU4XJzVifUQ/fe+S127X5ej7
OZkU82HrCsuc9dRq9VHOU2QU6XxtoQLLJi4i8z6S6w8koWdvS/7ofYrdt4wsMfwgsHZ9VfUZzMve
c4nnWnA52qLwZIMuuVdarwH8g+kLiq3UwujXo+3vNNVKOu8DL9CJsq8NmtNmpxLt4Ld8ilsHZxr/
1gzL6G9paH+khse7Zhn8c4NCm2zEAyFpODtXadoglAFLC/1cyzP46cLQGUXUyA4DuMTouVw1bN5Q
Qa8xWWTwPg75Qss6tUymlHrpsTzebKBuv5e54o9G7qdIcqStGT3/waR8bCzHlm3sGQHSD1QWDANU
2hdwAhqcM2bJK8OZRbyzkrziFJPW3YEQU2jzjnqoMFudNUw7/GHu7s0pLJXD1U1SXqRMrwSQTEjF
q8OxxhnlxgW5vj3TletfUJCA29ssRzOU4RJdLGaGy0nnNJ9Uzsw1yJhi1AeBvh5j0U/3mW+ACsdx
DLyGMJwIjSlveKoKYQ7KBRSDKNL6eVnDQdNXq81YGz7xN3+YbmWgRYMBX+D72OPdVSoy9nC5HTZi
ZUC1FzCZK0T3QPUjTU9QZywVyanOu2SEmqzqwEa3cqwO20BdD02IFZLZwaaYyEPlHnJQClgu7PJY
kGhzfWHlm2RFwZc9gzxDGZGpalTHJ9CH9AREqg5OkPCo5OJQjVwPDbyvcsDkINgynoD9PI9+DiGV
TCsia05pKMkIZqr/RB0oIzJ28Fd1IMPvjUrYdshwc3HdDe52e2EwDpHi5WM+/hW99ICkCiNvrtHR
/1BNl1rXe61pFWThnOqiFz8iy6l7JM22TvhN6M9Dnkg0MjPUyzA3Y0iPFwB+IiQwB5yRC1fFbCqg
NrPGOc7ldT3fMEK95Wy7NRr3II/p0Kk/jhOWbf+aCiNwlD341DsvRmjtAoePO7GIwrZHShmHNHld
ieFKINl9QaXJlU4I2XoKkZXV+aDmltDB7In7BkXK0thSorCINdZobhPOb8V1+bLqIueZFU5IcSrU
BWO0s+ZxddCZ1731KVUaBjc+xd+gxZ9Tc0/zDCfAJ3S0sosLt3Q6b5w4zgjI0imex2rE4aZY0BTD
mDxnnemfmhsbgpl1+h8A1TD6DarafPMPIE1tFgC7rNuX4aICuEcjwJmEJwkK4twUqDXaqexuILzb
5fnublikh4gAaq1axlsvJiY7UQ2+6rvm/z+AUFT2J+CqqRavQM+Itr6O8pqVQjEuntmuiHpHl3o0
GKknwdJfhQddK86rA6Nw/4fFgkazifxIixl7by1dmaGig1dU8Qx+YEVqg9hdAU3wbXVrqvRa1jaL
mF93y64LAT5J3LprBw8CSbn3sLhDsEwnG8dvOQAD1GGVuiBchJXmmW6MciGuBu6Isqqnm99ERgOj
hLwMyEJJS7NdMPgrA9WHOUWtE45xAx/C5v31//JubSk17J2KsRkYvMzE5Z5iNHNSHWi22U8tCVp1
3oFas9NTCMI+Al1jkX68VNEQ2KPundYMusG22KivQk9cxYA8fA7XIueq2Dx1gYOULnx6Yeb9QINm
GuYgWbR2K168mymd1JF+c3CvJhmaN6LTGLXZa2muJqk6mbi64sGll+omKj/D9CyiaDDin3ajJcdU
mCRKWOc77c8tdUC1gKUk5abYGY5QTqBn7wPj5WxPXnNaYsHmNR4wr/xqDjQyroyxZGRweKoeg5XY
PfQds7gIymXt6WT3mKv90woP/+Si2Sp+2z+abet/SPgDl5vd8XWtxG1A1gC3A1WQQP/TOKD8zGPR
gXbvqv+OLjIya9bdxXoNfjt+fg51/7aBIqS3S6drh9SWyS/GG3ctzakescaLmrhNrnodk7vKVp2s
GgYyIu2ZsTu4EARiVC87WP1vPtnQ64dUsuFERLpfw6V+NDb5y/i5Iol7XGtjgwV+iu8rpUNbsj4B
HTEQa0eKzLVzWmjXUaDXj79+BdMNqMEv3aImyTJVAtVxBZy42XlRy2Xi/z5cnZ9Z1eOPxddggtwz
0ZF25+5ocA4pAV1ASigsv71zMhrocOxxYtmhxQKA5Fs+0yhlAIzxdd1GjVWIEvvKtGZJmp7isD/c
EYndlXI3EcwZjXWm6l5eP2un/fjoUNq9/S6nF9xajI2Wck7BXaK4B9nzeMIltfjKSd3xxLTuyCxV
RoA64M3elNFvSnR5gcz+UzgEW8A6ucun7ZsOT8t2yHhLf/vkiD5Z2Vf8KUkf4Eby7eecHZgpQ003
YODw32N4QShs08SGJxbqhASWAJSb6t02MQySd65XWvEblEWVXNaiqoIs1N5objSfvXYxqnLT70D4
X8IYuJakG+7+DpDQzm+YKwHuvoZ4uv0Z9Z8Qvuaiv9JZxATPOdHwtwy3IvNuSvsHf1x47CfrnPsx
ayelr7a+rKtN2RL2J6ryHkgjADwTELRXDZLQ2iOUlFRXmcE2CMcNgW5YZFBGyF/V2TwhUPwm1ptx
4olxaOwT3VnxXpkRiJsVaYOa02K44oAjcWf7PnYLGwwaKFppvCuifzslj19bNSP9vtMQNlDRhSHX
cVtwJxRqRh3BopP89IAoOgd7ce8Q8FFZS7seCn4Pf8Wjexw01QenVOziq6Ev/mGyV2yvFBRRc/GD
Y2cMVA5YM9NV7pwMChAO0FhqHl+VYYwCOMIHCKNrruFhZuY0lopdk8nUBAov2tOYnwTEqJAzkp1C
nAXdEHrhnN5DNVqmy3rMHRB8JjeqPeSiefugbm9NvQfc+WJIY5sPce9Uh/F4V4utLGHaukl411ni
QoBV9Nv6AmHUfn/RrCWghl4LOVkm44ZRrkSZQSEHhtDImOpHzoB19e5oc5vXp7i7d8DU3M06UTJN
+YgP+jwOiyWPl/HktL89lYE2HJSP7OlZ0ni1hS7U2jAv5Y5K2gcSWq8R8bDJ0ytz5Thshsmki8FD
UasvT6GyH5ZJuXzxXP+MCHONEvZGVdiiv9LH3y4bhcgrmkTEl/rDy36kpLGqWfRWVaLkFHJNkt+C
RbtQLcpiYnxc1T7IjDdR0qnMY+hJnEVNXLeH49/mw3Hoq1S8LKw+0Z9hkfJJpRWTH+9AO2B5b7+8
hlQE1Z2z2yLhEjJlTEtCGBWybOQvCcoAM0wEc4a/cSIQFDkKQ6oW24TxZozmREbWOtZsu9iN0Lz3
PRRZnKrUGvbxaMuFXde9biqKTqcPF72gg6JjjQGWiSHw0vvijxN0v7xqYVo7yEuTYR/S3vdW9Ec2
g/5KRxHGIFO8P6OhoPC7hNQTAOtFXVvb32kHSkgX9QohDSxxUYCXZOslvL33kSxnMXQH6r9F/PXe
JTaiPijSIfDeW1QMjI9e3AF7guUyqjTdAweZu+zXtepp6M5mBinvzKEwnfykbO0O43JaC5sfIejP
ybHkFY6MbHNeJi+HopUmbqDPNXZFtPmldQGRK2uGPYJ5zOJd2eFLIlqVbd2GNy5sTR3B/7NDc2wu
oTnTWPt1QQosk3jTCzBM27O/LwQ/LNiL6E4nRQG/lsuHL3g50JKS+gPUe33d2ffkUQ+ir/VXkn6h
gMb4uu5jEJxVqVDjID2y/3+GwxBBo1K61Cruoca3kgoArGdlNZ8XwkaXpNvJvfeEZ3VdmvugPW6N
2uChFZ4jZ7vhceI85EkcrW1cR2AORcfpBJj/RfkdI6m6N/YLROI6am/wdSNfIjfaogvMDlteI1x0
4lYl6hYFGdNgPiuq0xXx2AIHZN54hO7JIIfHJLhFXF6MVjLzYOHV7FHET1MVoWwbjZaPusA0OwMD
6yDL/R5TCZbyHA5mMYx/TKtRJc3D5T4JIi+xjT15J1Dvc8I0yu1RqVr5RydT+NsdiZ1Q1ovVzsKY
EYzDfbBW0HnX8CAUJPTJsqBBSCOgg0VEVDksu5cm0m5HRoxtTGO4aD/8ILXbyXxr5zBniRuOQdNo
P6+C1fEbQRymVuRQ6XQK6RnTaoj8piX6z5frhh3ogepwmYoe7uT9BwImsqdXZj8VSvlDxaLR6j7Q
VlmIlGIXPvHSWoTmviqFnqXtwKT/02/LrJT0KkpLfN2T5LysY98w5KKkf+WGxOPmQ/73if1SJbHH
JYYtCy05BVNoRNNkqrsXhWW1QoVeYyYBoBfWFZK2uQ48RsiZ8wNWs4uCsr/sSgeTGsj4TjgFx9qa
qHtKgOjJkmTXmcovPlXK83zAn6/0Q2irGKJIMRLoz5z4Ln1/RHHRD67gp0G1VhVAB9QSw6+9w0GA
4mc8qXSxJOlzt+IiuvuHXyYSjObKRylOpyUyY+mN80WhY56uok6QsbjNv9rHZBkcAcDkYzfgqHI6
3H63gtYlSUDmlcQ+Oyv+vcDFXA+jtf3pmsgyD7QAt+UFus25mnIeKshm/qo3JMTFdZ3vdeIK/+zf
lyqYTDw41pvun5qUaf8zf2s6Sn+kkp2ThkEOSCeYwIYIidtfNeg9mnO32XK9wUwT/ociRFGBHo8L
o5F6uzKsJR+blFfsJuivoncpRNvC2QG4uutMsYuAV0QO9b3sRpHtZPwJHentbLISfpg4EFHhRo4z
CpV6J1ku4wg5tHKKNH7OYERxy1oywW8LZMBhqEvKKqPKeaTqyvwPBVSI7mm4gPZDj2LsnglfzNqJ
Ip5jSURFk/GwliyDUEVoSSEH5ipi7h12Xf9DpM6CwUML97peCnbq6J4JdTH5tIqqXKeygVymEt+v
pKgsw+EN9xW51BUN7Sqn6zZq48TenOdnzzjspIfl55lmiTHQ3DnMTSilaiRXjxCZOzN5ncw9hXqj
DLZvOV5VgXNk7rsOqNpwSe8P6aJgOmpK1PhT5sJUYb6fwuKsPCrUoyMiOEXNCF3vCTfpqfXSXkq/
baSG6v5GpbuUASq5fZFo2qfb7R15igwUL0r+onB4fasgkvxfem4286x9bU5j5w4Px4X9KGlkcDAd
hmWd0IQkABKvgdHcD02s2rtrx3KfM+PxO/pKXsE7pfyUlUb+9KIYtVnoabHmdS+U3N3PiB78In6S
m1nm266b2nOFYHHHRwkHFzdDebIvgywRz4smBsMPbtFEjzZ98K/mj0L5KUsZNSxKpNFRmD2fLC9g
YCyZn3cZBitc3f3nYi2LEdCmeMc3PQdlgYHfwYRYDDbZ3xK9rLnDbX6aqQY6OLNN1S69o1rgyHjG
A8YT+DegHV8ByHfeECgq4qtvwXy35K4MaHnlIMAt5YFTYaMbhLq6mUNES0DWScRtvH/9+WDf5LVv
23YClQLoGlu3GTEGRfU4VWnmUMSWHFgx+LCtoUcfdPbUassCytRULvJkBr681kTnDP9/HReB8WdI
cM4yAhW+8WCgSu+rbI+Sv0RQLG6RYj8goJirdKhkgscbvITQNLZIRVgGVBm4EbV7a5bGsl4G6aqb
qgSDNZuf0cKsxErZZrAAQC2V1umbnMP5lrIVZmV4CGpbJuhSS+lvFPO4NRvlhKaHMYq2rb5Fjgec
fIasplfD9CIyifGKgna198xPivv3k9m+PQaZYD5r36JC6AMFlW+g/uUB157jhmyznuDByZ4izVcU
wM3sGf8rFSy5ltfUreWj0Db0tryI9gQEFLx1upBUgnXPYCGnA/gg7cBm/cBhJ3H1rEk6JxG4bqTq
0oxgtxMhDgzfuuPskVBc6shSiH+dNEK+QvIoDAAfynTgnjHZexXWTqz5c1gM1HTbrtXFn8vZaf14
q+GfZmVXowLMFGeLJcCGS8khg2GfRGZJx1SclA5IU/fwjrrMOPSIocpamyMrdlac/MOOj3DUcEql
gIJW2wlcNwj+VFJMGTXijzhI0wwjUdjkoJeUTIImk1IojKcW9vIFn0NGIWN+V9CDpB4+/hYrm4Uc
Q/uDvXHIo3Xsx7YL5zVpTnW93DVKFiN51qbDfMO3Gdf3Og6skzzQpfNNtAqWsQPRp9Q1Q0D4ywp5
ZpnIEyUq1YsgA2/m1PnPOP5yWnF7wLNFquX0gOaNZiFvuXdepAZzsGuVoRzXY++uujihjVcXwLAY
bdMz475H23X8cazA+WYydhSVJNAdOmOPQFZTyTf4MLL3UDd7dafje3PNoDx1U1t8UBLVJrKzSuFB
DmuU7nVRydBRaSqCD6SZELrPwE/01MTCPKSa4tkG9CTWONstLAeao5jG4kltEvNWm1xnv6gwtFQD
kSMvgi1HHHhmP4cQK+MD3XE8gzrMSkKwG3km+5885zIitBUGBg9gGxu4jpe+T4BTg0IqXlGrXdkU
z+L6w/58uT6Tww6B8bN5qfd7NWIDgpM4OdIR3XLmMxzAAyLF27jqXat31YFZrJQHvOu9Ifz0M+iU
nHaKo9cIXoNCOaF7drw8bkiy+Z9C5bYcI9TLFvAgoAVmBN403+EgqM1890hKucbh4PuTYgENg1fJ
in3i8JKMau041dpXqQKMvXLH/nTFRKjw8O/TJTHmLgPCEcKmsOCckzlWLgA7dgZ+gxMJnTB5Ncew
PY6S+Rmn2Iin7K2BI1tGmhNSdSlbxvhP91p+KP49jZJiDzTQ/CquCo/k3Vzd+e/nrDCfwsxJMAfM
TpiBfXDXttTx85TVlUQb08VSSBeCpEU/s7XQsxDeC8TkmJe7NmJlE7cEk8gMVbH1tzlFw40XOQfj
UW1fskyEzfe/Fw2EHvs2iD2t3QQ4EMMG2nOxEg1G8KlCbnX6SyJk2Gn1DlwvWfTseubbGkYkXXBi
sRcJMFPEvZCF073XLOt/00/b38jJYqNZST3afimj4Zf0BUYMRMPu1laAhqVkm7VSGqBJrJmsC9Jg
g/KpJtNdClzwC0H5qCteJswV9oIptiZB4GSvSzpvBQLtmSAbWHIGx6RdAQwBOsPZYq1j3Lz5PITw
lDBKKiTjot7hQVO+gJKGJmjPa1ZKHoaeb2kYs+Tn4cjb8DiZSOMo0cauVZgMGHnb5Bhnc/E18+ip
CEgN1jfZ7A49ol43krMA/jgfGfBu6RfHv0fzR2MIT2YjnXyvuu1Vlb/fmNaqvyVhqhbXNXGNJgZY
Z7Yzmv9VQYfFNL/+JYiuvzVl71mJGqwk8BmQpP/C8LaUY861xU+kDPsO8J0fLc8FkhgrcumgidjD
VQcrTL0BCpwo4cWb82+XNnRVmGEWOJGHygvhZR0KVMpTM92bx5JbmvRwednzewFgume4BDBiOPYb
yxpl0g0k31GzbFtmgNE4TgaHCI2T5Fq9gNg7R+ISHkRZjlNN5R5XB8eK7s7L5Tz8KuCFy1ly+q7x
hs50uWYPflL12Z28VYBvy5Jy5WMK8O1tXNUu3biMgZtP32iZa7cbIMKZsKmx2xq5DAHbGEUlxNXa
NxyelcxLawpPeakee+7z8WVFHLuj7U+05Kr1qFqHP+7sNB0633EN5cgdFcQlrVWWg1vSOSKAT9Gx
fhhnUhUI2nxMhpOXtsflYTrJvdgyJX6XnvVx7++tJvw8Zpb6RgFV+rNMeKpK3QB9WNMOluDzyKHT
pbAkgwbXIyi6X//otyuBu2Jlu6C0fsQAeY52F/0UvSc2zuWr3s80bbruULuY+AFAtYMVoTSrQKoA
Y6e3Puh7OeDtbjSuH0XiguBOBNq1lkXdkeLtdD1bZ2HixAwNHTQFY0zTNDa41L28dwaVAXUcOwyx
zPBzHfl69/gqaVwT45qTt0CKAACvUtASVAmS1N3uZM1Cf34BIhF3vLR46tEoxVbsMCQeQSL+jYu5
bGvJ3H383Gnufbl2mFs82AtNpZzdLgkCtC8eYzrr9R8eMDB/R3u6R7czJ47cWZnzyV8FV2NjXdd9
i2wStIIpHxZlOW+QZ+b2Mi0APA1h+p02yBPL0wzBM002rGetKlB7sQ8O4cyJRWHFFb9izHvyF5mX
RTGZmImaPwN0XekMsVTczMEx9R+v8l91XHCkZrXkPJY9KZ1CI3Tfaqkj1knKAAH5OfEUF1EQq2fc
Bhlx4U4EHd2G6tvFW4zVmSqgwc5EN2aTC4EssBbOGZHjdQsAAPw2ACz/efzpCYNL2a7V+KqcSNFt
xF0YJoXNUlpqYz3N6E2VCQD48dTw/JnWBy04UgpB6ziDjoAWqA+yrmH5rnAUyEUrF3kXLmfKNx60
cijWUO5pEgsXZiXyEEcIsTiwMhtG6bUjCtTOxbMoWynMylSSaEBRfUp6Frt664qLhNEYH9dta3yH
Me/Ufd72EdindIuEEOOQNJ9qFSgNjrDao3vVIdLovcj/SMtnGyWCOdX0FakkqOQkQyODd0W5vXSQ
gvFJ21cwL5+CgXIM6ePBgv+lh27k+edvLEPm1xVCrx2ZY/ReVAbsEi7nylfE2Bn+ehYwwOPhL0oJ
OlbHmVWQ0czdl/k/zHvLbxi2iL1zNDufZ3L1dq4kj5oihPjkSGERFa1skjIDQL1jVwvKyeIlQeSe
iOtWpXSENcRgx2SNwpXYT3kErrgJ2iYizBDG2el11QIB32OjQIk+oBiLafZtmRAzTZN6zrnJPSKj
qYJoUPH2sYrpffhqgQMhhlfLaLBgD8DAf8F3Qrhmt03Tuz96xuRg47GGbvvwxYGNgPwHv9UcY5th
uzHL0xGB+nfqO3YHSVSmZADuhykbkwK5Majh8QFotP5x177VFUkSphtqp3oVut2VzQFfUQF8qcur
kzx9hqWpsxcj/CEhXtIe2bIAFfgj1Mq4++RCaOswAL8yN3f9U1s+19n8NlpMocmATbgfp1CtWaB+
yuXc2iffNGsxwO7n7jjjwfYSMEC9bJHCbVTlG19bLgLwN8wDRnTHLFaOgDndHkNlApAZl1/8NMIx
+h4JR6RDVrQqJDmKBkSigcLquaEQVmqtcYxcR012ZvfCeUl116pCSEQCvxCOpVOagdN0iPP2Ksas
p6qiRF8LS49KHz/IK1QHF5AlV+UyFifoczAlUjPN300gdNHMO7XkRV5bJ8oEc+LLXPLIRJRomkhi
x/+VWq30V25BVbkxMEbAmAdseaGXsyNYmuDUY6ih3xDgKrw0ekdn1qA76WxzAVXwklmhWf08ZkC9
9Wag+MGadXiwL/zIZj11mVM4rxPQU6N0Zpn6gV9GQXs7d82Y9L6kZ9QeVSMZOd/YgY6/DJ6+i7WV
fftb9a5NK13Zv8aSonwMiw1MIK4OT7dqd7ISoyvH1Kf9S/HXWZ+6iSeQ5kGWBRioulgybUeOR4+u
n1Feli+QPd3nWOITnmV6lCOwnDu6Rp2PUaFJua32LnFsrv4dc3WHP5FpIY4eM+RcvKa6Q8Q3geLC
9yMph/Ggc1AZNuDmD6EhcdNck4v16oSx9cK0BUTYhJXz1q0/9k8zX2bBXJkb4uI5sAbqrGlTrsNK
Z71hq3J8JXnag1ePBPotyccInhAsxGIuyhulGTvn2Z7ENPgg0nFjmUhIIQrRRmUvyfftFosCcuWG
T+TBmfr7H119POwDHSlJeIdIwYsyd8pgfNYc0frZWqBCZkjlRyIBy2ksEswoqxyarJ1tDQihHue0
7tqCuAZTotEcqLlReGIZ2BpnzRSQx5K7c14TXpekwwvLfTRb/417XY7K3KrEz3iS9MGO6sc5gE1v
b502RMSMNId4BXcd3PhE7pNy6PPh6QjzZpy1npLFWgq6exmHBTV0QikRoLkPm/pVermkd28UorXy
wCSD2q+DIkhM3WKHDJtrQ/TYVe6yRWw8jFKYkZ311QpJICjeN+CT5r3eH29djbXf9IBr2MzB2T1M
cz+7lhgoNr4a3xL8juXdmuCpkWj1EqTTydkCvFK6JvzPMZskNZHJZP4w4VM09/4/Zx6Ocxhn3OJQ
+TIRHsQ4G30zxfk/KwEdXa94O6XOoK5WWyKpHRkxwZ79/P4YB66BNYu4LtfiTWwkTbb15TwGH393
6BgtrVDv2GMFEwbA9b2deAW+MxR07foFemVEFBtASbO6piK+Y1R7YIN2VHTnJuP2gjZKuH+4VwTm
swfMjyxTBJsn9jyt7SQO7D0pY9KUn4iHI2iZxlTq++YYHW87tCSRQUtFdgf34d5P0DWgWoHWkIJ1
RKvlLlCGsWDyPcFu3SGYdNo758rF0yBjlUGf3arjjqh/SqA9xw8jRhK37FtJCk+pdg9EgYg8l+eZ
BwfUTeKZiECXm/DSdIjrDXnzX9okblELb21XJOffUKGkSYFkGGONrapQgcV0XS7xR6MpTE4hkb3K
KLy8aNyNQ3DR31pyS+dZbutzOlrJcRYwEiv9dt95MWaQsWYHFXv6jEPlv1uemA2RFJlkna+CYP2J
lPBW0MeO9SZ2t8Bws9WMHU0NTrmwJW1OZngz2HLlfUjSafK6LiSGQRF9NULxI8989JCZ9lBsq31x
nDIIH+S62ka4JWkEqIldHz7ial3LhFKJpxyqAopD8iSdMB7QjhKARIOnrbk3aFRJ0Gh+U3Wctxgj
jfkciGlBO3lq8GQpOTP3IKXhzXXGsfcNLLTdfT8rgRBhqh6E7/i+Pz3mAkRb8FNLJaYSaqQQHIeq
v36pHoqfZBG3OVqagMB0Ia/S9WJ6BNIMh0XrYNwMb8iQfyBaDsU0L3p4WzF2MXZehkuxQW3AaShu
IPDkTV9jSU+n/JxOP+3TWb3M0y2wg3ZJkhqZBO2jGr+ccmyeIvxVpD5cjyEbqzRjwO+LiTcevbac
7/gGGlMrwsdriBUyTc9rN/zPCNbzGhXVtkMxH2cmgSx3aKzXFO6U0/yYEXO5rhiM40ulqAp/BDrq
FCH03TVdZ4wUEvcvS1Bu/PxRHQdMHE1hdGW95OwnZJKJxEFKPYHXMAuHcQ5Qd2PVflKKBr1iYSZk
o47HJon/PPi8C+2dtZg2U7ohsnY7PFC2Bxp58tnLbtd5e78+el/5XPZuyZs2tNUonuIKfWtuJDn5
XJ3PR8PY/ta8/PoeHvt23qgEG44Cdrcb5SftE0infvz4LGzVvQXKFhG6M4qKnO+S6b9o1bsVBGWi
tHPxlq0rv39bYPuBCKdEDGWmGp7zZpyVabkEia1YnHPalOHV9Jx3+0wXuUDncwTB72xkIlNTKaqH
DZKY+KYELSBxD5AzeHWc9IA2AVg2vFcG1TYj4QVXvfZh1KIf9tkbzadW5a7jifgoWOVxnMSvo0R6
rhwipYvfb97BN5SeS+inilvUD2V1w/mfpTqwblnzDqCY2G1tBvm6uZsOY00ulW3tt3PKXGzLmAFs
Bto7Vy6qTy+fO0nZMp5lH398h/6hcNmLrQxl4QRtKQePF9Etd40vS9PcYyAbX1XuxC6ZPiinQUuU
vT65irUtNO1i3gHVJegALpVXdRLtWzsTnl03U8eBTPSDFN8zGMQ+Vfd/M1HnegM2JJgq/m+667Hs
q2ZRhp2jEHITqbT1a9EPej64HshkGtjClP7ObKRLZ0NJ4k+N2gJL91zzc7oNwPXk9gfm7qhKf+5d
exAW8oQ6zR1iI68rScGNYOzziyS0ZTKNDeGyv6UeZnv+CX2m6ptCv2Yc+3kmERSAPsvF0JFYTtEn
k3E7QzNfFrW4QLeqmna4UlLYMkjucsElvFALsfcUbjhr1OqSPceSrHBtH1Yg8OqQ1u2gk6BWAwKG
GwHAnHWxViNQcJvJdtKMBYad/0kMsWl4hZNBV4CAkaosBi3DxDx1IVx+Wn1exVRzW8Tc9ByBwn08
BTA+z4wiyl+7DTLU7xQihHleRiSbYW3Zyfp37sKtChhICoMAKmfbYkNNmLip8Um8mZXzAl303bSE
TD4saVChew+EE9X0nruP+aPOR3Yc88OnZsbBNRnLtruuUecEAnf0/+7ojfVVHxputPwHS15enwQ/
mvfAtS1iet0SqLrwqESAPj8yNUEAp4iKEmxOZPu9dQAQG4Ubd1l5p0CsOiOWqQ+3RauAN3DuBSmt
zXQakF1LANRy9ZHVmzJ5y9FcHx1sdbSg62mSMNkcsU7F6peOGUMvlyO1cDzHfajQn00YbvdWc8YT
rQs7GU4k9XLkDS6L21e+Jdu7RDdV5DFDR2cbIpMMIW+qcGEyI6fIYYhbKsmLrgUQJWKEXNvaLdW2
k1KKAdL1hXwsO+lxmiGpZvVmPsdRTJWXAdHA+XIzf40+lOZ7AGlNfm28bwhPdbuv6aHabaNypSHB
Q0a0QDCnD/bHompD6Zq84F46NvpZuoNiUO4zDsniU4ORfzd0wTN/lAUe7JHXcBOUNnHH6ppsZ5ta
96TfxRef2g7NPFQegq2gwjUcKvY8IzzCx5m2onSuRfgSC+0RpTqW/8F8rlj1d37H8gxNehyf4ck1
eVr2rzu5w9EkOd27BeC5oW3Di1+H2Er7367g1q7AnFPGHz0Da6LLI/kwj/7f7qHpM15vTuQiXh4y
6H7C6alJqrI4eZNw04d1WOVMTDzeDkYkOCci7FgTMfIdrgIwToWCaGl6Zhz5lMNlHPn9objgvSKw
dUMjqzTEFB+2lo0gaF3xuLZlPwi9IiWQJrRK/iti+EmJhZAtViNLZv98PMlHC1xTQLUXB2739JoQ
M21qh6SxxU9biQQymCbXyT2Pln8Zl7c8RVojXvfdlw2XFg1cB+QA/cIOmp+hpqKb19LCz4OEbFIx
GvTGnd9HDNBeJhTfNpcesbjx+xsikyN2202U6bMiSEdBKnO28lmL8LTKLc+ySAN+tenx7Cga1+iK
1tY24FNeUqr1iNvt2HHXJrPfSJ/Jg5xDZkK5KIQPoptrlOkjX8zs0Dmfi0tB+cXIbfWbRm7Nfafn
WiCWpbzMfSp739wNzF8OVLyrjbjqX0gtEzs8P4yi6KVTNQ2WDLfKPSfiRNEEjCv7/MS2DnnIK/sD
8vbBxuD3nkBrE+7tQkJL/2kEUr48kYsaQHTMwVwA+yShDlspvspfbUDOQDrpI+GESCvWatP91ZWF
XJ2Bc6SL3Rmx+5adhrlARg9yeuBMJxGAoEqi9nLtKN4cf7EFuIGa3X5KXLdhLSgIhfanOO5PFFsV
6EJGGSrglc/vopjU272zmfrMUh0p1cn0QQl+JecoQppn86j9GGoc+1Q0G5M4ZuOc0bk21dKyr4Yp
IAP7sIGVzz6+zP9eSxaJdMP+GxIvetMKoU1cx/4zGBzGT4zCSybBZo1zRUrmUKojznfUfCPTyTEJ
mdNGselEIkrz3WzRshpbthgqfrbHkPXgyQX8wjikMPW7A5oJwOLzg//vHITwwECAarv+uMcQF1rK
L/s+1anRFLYDtpD6sDq8tV0MKspLCerPRR61V5DLdeJysaB+xzhBntLD9ju6pTiwBZVT1toLaf6x
DjKmlu84G+99smPrqWqS91Ri0h+VUSSCZYGMoiAjnlS1Z3uepDUYFGD5O0k1FXrco9x3JBIWW6O3
cAVYAcUk/DzdgpFOwl1zKHw06BJFtncxGlWLGlo46LnvZYy60f+O4ladAwHiqfOVnx8qt9uRQ7/n
rkUvVPTwvj55k2+PFcnuJTDYp+s+UT/PTEYj92xpylFbCLE0jIE0CdhaLmcKMr4Pk0ot5nEaiHZL
vpmlT2IcMG3gJ4LGFJEmtKBcTvU2535AIQL52iGLZoFD9UoNHEYPlfv+3kalq+n6YDkQC+FmxaIV
WvrCTqsD1JLkxkjiEM0FoGhyuxjIZMz8rwDBDeJS6SmZ79kXgiMtO4Tkjxy+6weQbknB8RGNf0QC
yImB4gVq8RFeMBgtBBrclzcNqVtURodkr8pLVKDeYrC78opoKIuCgQhsEBVQ0/hL8/I6BxS+z3uy
e8rq55i55f+xxhYRPvS0PSED95W5mnhWqIl8ps4sjGdy0M5plhi1Mw8T1ge7y5LenBaafKTeB0tP
RQlAwmmfr7GGnpGmDZ+dhNiyscRc5bkcfe/VzcUbjxCwYbUtJ3WL/aXqL/Peqp1UGXvwS0MuZmEB
goTG1BxGhmIqCIhQdC//T4iv/d8asFY7tZuhtac9AQdxEP2is6mieKMKjzNpQJcSEPm3d35DKbEb
hhI3cu2IF6fSUmLWDZYlg+FDrms/p/YBy834qx0mKYpmX+7hEMJi+4Li1TSwLm5BuIGdhhSLULxD
+QuOtoSLetGg4GyGuVkQg+28qMgkGQUEstFcN23t/OdCWETVe9YhswWZFVgaOOEbPoOWQlPItGo4
GdLinyI14dgFIqTf+K4gsVElAxkIokYamY2aLAWK+xwms/bNnSKtrH3iH7x2kLzojBVQrK73RhXi
2ChbaS5T8rl26pSr27Teb69MZ8ptd0IErDBf8TAmQ+QK9bvhNlflMsBeAWWLDA3/oSrM+iNldtLI
ntb7p6XbN7SxRVwy2l2sSGeniuJAvWyOLA+A05/T6OqnkftadyH6ngdqZeEUgnVH6lrcRJW07eq6
plF4BnVef7T+Hrj0F7win1TRvdYSLEHCeOLHIT3LG4v4LbvgGxQAYfV0N4gFTJ7/iCXRzY40jAZi
IJhK2Rjvjk+9HYQSn7EPWLAeJ6vN3Jut3aVw4uWBmGUwcBj+hFUGHIG3wJOIHjX8qyWH9KoJyN1a
Gc97I4ASbymgfVkjgh8tikjADF/k5PKPeN9Tyt5YVtdytyIz1MGdV5MYb3izG4ANYa95VeGrsYjr
kPFs05oxv41f/DwMF2S1tI/hC5eZ0Vto6NMidnIrg/yvvd8Ns4tAYD1U2myXX88vy6yLxC8MwA3g
YuQ3Ek61qfRi7DOBr+YZJi5qNTouFoCtCnf6CV2Gmwpl41+leZLSGZAyay0SqDP3YE4Ec7iajY+f
1rsEWDE4q/f8mUJe92nNSCpSEitdXHP788mVIZXxfqv8RQKgExMYiuSVqkUZN49gJYRRPDpclgdV
BIgSDCxU+NSDmBPaBR0U2/Ksz40sQh+bcAz4AfJO0BCn0tTO/HxTN5ChyzMYF92+03ho2gByv+OG
bazppOu9z/bS3sdg/5eQqPaf1mlOX7mq5t9pe8Z1+V8aiwaQtdWd9zPCn4cgvO2zU65aaSvBccNR
bONF2Mx9DyIst4aVl/iEhaUDte2uo7AdXsMHF1A6+Y68kmDXvfjAZwjy3VfgIwRnvkywCSaZWpNv
eklA/0pgPKlT1QhQnGO7xR1KgC3OR/UEjRoemBEaWoLki1XNBEI9YXyHeMRtxRLrUUcof1qTWit7
1PAi5H8zHIO1uR6AWaxC1YOo0Gsb+Zv0Pt1RvmEINagAVMPbMx0bw17LSZ72dSr6HGP5qSjF+Lhi
8ivUkBLlwFSK0n/OKHoBcZQiHW3vJ0+IoTGdgoUVfciRuO2gjBz3gCT2KvzSkOwNPtQy1AypnweD
s8drL8fW+RFvKxq+R/RxfkuyVkPJCaTZsIJvOlt4hfJGJ+MwD7dV2wNnfCNxoKRPPwUugr/qe0nY
LYBHdD7von0V6KzlDDjN9HECdAS+QnBj1pZv/VaFJJkhdaOvz1Wo25In8IaFSpg0wD4SiM59YMnF
TCoJJKZR+Qt8xkKYhELQrtnSjYuSEecKJxsmqjUxV/MQMmD4ZatHzXTXkRVJXfORYeL9mFudKXgA
eYGygpkZRk0tI0WYloxFDc/HVdPKsHiuPTk4Rvix1fb8yDxYoeenulcbvmlPDpHycb2C431a/qYk
/whSTynu9l9qrTELj+S9ocSho2WW1L08DIw3t3XsrByec/YALnoaskftoKR7Gwrmb/N6PNi2ZwYe
cdG74i8a3gCxuJ3PBlRQYkcqh6TI4AxF9lZukqwk5Fbtz/KPnhwG59DbDvBiGWYELf/XapONYBwA
eqZJliYZqMdH33ESUuSQAQRPYb7nQVisAgh9vemjY1D9XSe5ncY5u7KOw1iFMyNkZ0iO18tg0XXR
cSybcDflz05nHNuvJTMaHHuKfEWP9ceS/uz4O8ROc+zFxaCiakTOAdp5zMkn030f5m9DRzl2L2pq
QCewuiK2BufTqeO+gD7ZXv23XOK47VXD5Qz6H8D8DllMzmwyGYs0nQSMClgYyAGgk9sP4Tm1f5mZ
9SPX3BZXuA2K/9YhqGHM2DO8Je9YHW4RQ4qrKuSixCGhP+1ByFpg3pcHtzNZNEHCE51GtxQ1UBFX
64PMK7VlntpXoKF5uJULZe5ytY7f5axzOsoyVvw2uTqsdn3POc56VJ2r1lpN7iD82F8l0ts9jd5E
kI5boureNXn31TzWQ3YeFlSNAwKMFOOEDeR+rkWLbtUVukfjMwnXiNwYBFaYpYmwn5BnRLQt7lgE
hUrzjdHqgJKyJjrXSgNXbUcJJ8Bt9L9QSJYJMpPsD0AuofvGHUjZ6yOugjSZ+BBymW4KjuZT0K/K
XrvoU0oucu12YDdw60lPD423PM+riN5NdvlIr5NYr21RWPKJVySJSx9yAlP6r32US6UNrzEtyMPg
3Jvdj6xZ37QJncV7hrAoUbjHr7cZe1D/O7PLzaRii1OycfzHIR88nqtu9aQRjQVagGjLlIIeOwTw
/OaRkNaeGS8qR7wHRHqapK9gI6L0dmjCci5LV1OUerTyQEAcldWRQO3sQoovmGUEV/GIPDQf2Ayx
zq+rl/arjh7lE8IJwhIgWwjiE/fJoGfbQ2Dru7gxZH7jpd2NJBAL+482ORmgUWdHk5JRzepClRkg
CCIsaBxIu+gPef5fJkJuX4bs0CbWnKaCL3m66CBuqdVs3oF+9lshkTo/ZspVlpENjYoIbMvIMZxt
2EwXq/87XaJIwAKXNkVYJF6sD1xC1+GMkUnHnHIJUv7NAhvFYufXJHhnAua4t4x5AexPKqOFuATj
rkLrOjdjJbev6oOXfPJZQBsG6kbcdkYOFw1rHnTSvmhM55dR3g/VfYMPLV0mn2fnXjch+xUXqhGV
8RRhkOoUwHtd1dpvJfgHoLGxXwKZ2sNkKl3dp1ROX1G/8MhkGp+QHhDqTQ7yntODTG7owKJUCLFZ
iiMsXlzSr2odP8d4oWjQmXeumvRXmYNCe3+i99e1ULbkRFzZm0E0GyJw6wk7BSDWEXSLtDDn+s7U
W16jCIVYmpGsd+zuBcGmf+TAbHKylqVCOV6rEg+JawfZUSIiMTagNqm6QNWE9XHW/EZLv+j+YLcS
kP4O4Gjy7Zq1+FRfYLvmaB3sm0MENnznBfR9Xn08bfAWkDHIl8iF9AZE9ICUIrJ0OWiwMBhSGt8b
eJ8oyh5FSrBsEPc3BcdeuCYwRyCUtmSf7hDj6F71s03nMaeoM+ZBpVSfwH32qgm2J7425PskD6Rr
soeqCrAVsWn7mp4Xh01W6yeiZL0twFSyods1DdPexrtD2pd11fYHKItpi0MPHebChSwWRnyptEti
e3Ma+Xp/KcOXocYVJnix9mIfYkLC8OFkSZ3UXHnqiZJ8EujXICIH7wRIKj3H7RvsQtsu+h7fHqRx
+eiynt8gGO5jb0PIjGz4Fawy+D7BjKmlOpny70VNXzXc1qBJoI6BAjW+Cr49+KKBiE+YXLichNI/
2DS+TlNkM9We2SLqIXpgtBX+H0MM9NiMu13xH/TPJ8uQGdivtIYi16eEbJesvKdwsnw34f9FQl3Q
juHh5CLT+iI+MjBZrDLdn+J6AYuZQscrnSaa4DwuAdnn+5Nz1Umu0sbd7qIjMOS6yWWzmWGmcdUF
qzubxJuA9JBpQe8baz+x442pI0EU3HPreYdwJ+9QpXOmDkPRwy+QO2pRRrnckHmqTV1CU51Mynxx
zngHImFpefBresKgpLXhWFXiTxB5FEXjDnL2uM3C7qYOfYXHz/AvpfeOYjZvnIulOIG46B8Ch71L
rVa4mPQEncTKKayC6jez70QskyB82o94DIicOPIFVJzgqq/oPoOo7EcyyPM/Rcb1diJtysL1ZRXR
EI5Fv7Cn5OCwH2laEp4wHZgoVCO1bV1T/ohACLVKPXKYAtDD85Tru4xwaXS71nKTAnHPktgWO/K+
udG/K+lGfsx/tH6+FFhXNqpA87HzoPPaeOJ/MZnIMWkSqWtILHiJsQVAbXXRh5PgeTDttqH5jcXj
T7ca1ebPKKndnaBsOr1jDHYJzRzaMPrWz51v2mI8eFHtE4j9jkFy2o1mt1vbTP3Cs1f69bCGrcfk
GzACXOeHNhHHkfP2OtEVsb6hlpo6QfbTlgnP7qUFZE69lhEx54HP40qXryIYrYbPbiEakLj24bYc
jsI0Q288wmALSnrp2hYjw8RTajZdkyb1JoEvij0jP/rgOouCM87wxBF4IAGSzDbY0S9Pk6OgHA60
W4tDkTRSg1LXNm9MvGB1CUlbkzq5Ysc8LlZZBOR6fPr4Ya8ka5BwshTiWulDEgVGl2raUCw1MH2p
nkqdrWYeSx7yX8dkDUvmFhU+hGNUvEWXp9bkHa3eCGEhmE1Y0TQnY+ioOW4gyz0neQid8y0UCDkt
YnvjPGqxmcKJse9L8XyDZvvRbpr4LcpOvZanCbeDPNg9+a0gu9gyJeaXoipsyO0maN9tZsecYbyC
irc1yqMHltFqRGu16Z2typdA389sqCSPy2MDz2FFCgXKaTicjJoQid4ST9SA8YR/DZe4iPcdPu+U
0mQ1TJMBPA5SvHLTW2bKPVshNz+k9r3GacB8tc4tdCidCeMqIZzjfrgu48ZhOKnwbZES41y7A93o
5//GYtWut0jb+EgdZhXUd1PolVZcQkNYwDEBohonHxy4omilTbig5JxpNtPtDJ+++sohH211cwy9
zq0kWwdesQOR2uKJLdhXShM8w2vU/aIrfsuOuY3Izx+AxCjgZFmqpOPPqiKE1FhzhBB8nmd8pPwf
pzmXm2EPKc/XnfhC99c9pSL8XFX4+6+s0BI2FCUTOgEr3BiTiFSEAylWTC3Hprd8pTyr08bAih4x
UJEGAZ7mySS6h6e5Q/gX1lI57qMzcJsEshotPJ5D6ASmJV4ox167tqmv3t+o53zks0Bm4Z6TMH2Y
HT5BDdqao/u6Iy0N8/ADtrcKd+Insw/5RougViB32MM8Y1Cxpa6L93nTrr+8li0emNP3uRfJX/kS
owNW/yG1lPduS3RGbR1QqUv8pkMscgcBnsKUKvivMv09wDqelaix8hQlsNxRZWulggT+VmOsiqfW
djIg3ArF93/q/fcpJkA+vJg3zH02WcLFdylup4JT5IwWeOtLzT1dfxia00JWXpFAR40V7N7DmDMZ
XbAfv0XIICk3C/2gbJbtO44vvDwG+SFf4ZTZ+ahbMJzhkbJVtY5GhJ+qfXzI4sdfFcSOphfbkB5G
m+O55LK/SSjq9wroPTOtb3iNCN2DsN4WdFmplkJL7jtCiyjz+gphCVftUWSpf5UfTtAXfFm1sl+X
oo0+psbF7DaBnRUqrGDUfFRfKpswodQd5Re7NVG6G1d5LV/RzoQ/MtPvvN9Bp+yN1G+sAVNG0vYN
oHz4LeWlxw6yLnbJ2jFIsXTb3btH8mHFBLaOXP0yWz4UryplixhXdmZKGHqltCusSJPImN9Razq0
UPyi9E8Uy/XcO0k37NnyHfHtG96n8++2HaXfP4NvE5lWsTMXmw3gA3dD8VZqTE9QFXsdaRf28igh
I1AdoNITJwPCcua4NeQS5EXQbvYjETu5BunEhgWFgPn3bnjAib7AEDbllSYEL1YL9UYQO+V7uxM3
iPTcRlxFe/kZI2mYdR0LN8DlQQlGS5XS/Mgx7F8CcoQ+CGBDJWIta1nFSA67dfj/CURlqNf3vNAK
etFXp84tfZep67Yhql872+hoPQMa/sYcuTxG4Ljaat+ZJQjuEm9cTyNaHSrQ5gUuM80RxLxc5ivr
IFHCY/W1QkQW1hZKV5ZlxUHTEW7MI2hE9dG0YcS5//zf0zad+suaGgTvgPtF8Ifvk3Ut/lWC2zPK
LhgyUKSu3iXx/TS45qSyKdJYfBE4fms+jFcYqdC6KW1Dg6Jpc0HsiFanjV1WlVBIX/OdOblym5Ep
X1Ar5iws/L1QO9BY4cAdFOxB3One/rT0E+p5d85tvtvteFySmESdDRM2FHMkyLxmJWJy+kHk8Xtj
2BkB2391py7OYNmNKQkLHPwnPRrWRWsZNDsgjcCGqpOgc8Afkr3G3oeoHg7gX0qQSK4tOglAdMxu
9bpSHeQ65TUKc54oleAOJhI0K3LAGzZ0kT38nOJTK7fjc0DQkHsAAkZDueU4iQ+ZHBjh5AB5p6Bu
qvHoCEZumD3tqrBhnFMB4BOcPIHdXeI9WYE06yQ0/+ZQncxqcZl27WAPmghy46BIGbR2nM5JHV/3
CVONk18Yvzo4tTiD2TzDGeYG2sqT7Y/GwSXhyRu/DvTGXL3Uhx0wkJesGszcZBeNnA8Dv3BqP5Kg
GPes9oxNOZ3oq2a/3hgGpbDeOtbpUpo5FD69F4GBAUZlfCejhR9sxaRme/UHoC6wDDHGhogShO9N
ENO3Fs7EinAvFdG7cPJoVPK+6K66UP+aEOKBO6rL8zp9pbkToVa6OImEcGxKuYDpV9ZrQSpk4SeC
JqAXfwn5ZKGS/Rdca0Y4Xv4SDHtlIx4ohhgGHqzTo70rw8oorOl8RKiSAKcI01ASXImtZvhDBMoL
1+ntPjhWk21E61EwITdk9MDN3V1rCeCKZSyWhFv75Qce3lwysfxo3SzcAU0xzcpUBZtdiD2lUrW6
id3eD/XV5s0O8ODz+Fdkf3HQM/9VMVGoIetutMkwYFSBx3zLsdkqEMJtJ+God+hDifZ9Ynlij0zq
mKU0e1wml9exOXRM4dYYm+iG5HPMaaFs8xXBJJoIUc6WQlfQde4nUSNkCF8tdSi3J5JErJCPzdFJ
6iyQIeL03ifVDAkpydGQRNA9yRUpDH62nGF2F1SuMZzJOEYW2orW4NsfCa22yFjLUnSD8qqH/rhG
08WymbRA4NZhkQGPTzlUxIyQYLFWf8156YEmvn0ieMnwWJMUidKaBD4ad2fxUlPPTmZ2K5SSWZEg
sdi2Koe2fwxyAASweGZ4KlzENgknQYELBC4XgoV5AWq++NzJdr5Pnshg2Vp+3E+XlltSg97ydNI0
R5YM/IyAdppd3IDzpkSbe7Ia3o23r+rHhyoYSNJEad5WsueBOxMJEjuCU5yiLc/vT75VwXDRk8sb
//FwndP/yFSBPCr9ATMa+rQrACuQUmjTZsm6HI4Yudkiapj3NhKOVreczCWZByXdGWDjtp8kT0Uq
152uj8FM+RR+NXpi1dh5yQt5h4Q25yWKnWYm22VH10EjywOOiQxH8EwnlJ7tIvv0TB+PDGuz51rZ
ejc4MIwBTaKeBRiUmMyEszPYvpk4tdAwHf23jXGx1hpNK0ysiakxiRfAq8Rj+g/TEdMU47MdfMYA
Bb/2ZbyXweBcMIMHqYT6ud20n5ICP3VABUmwCki5M2Dh+npqyDLHrB9KV1vKIRz8Ao/rNC5cguap
Y2y73srgOFpiFeXehC+bWUP6IuAydQzcEd4rCyCLejt8IxDg0k0UsYhY4wD8EC3TO7PpBO+eKxn0
SRjGvXFgC5DJcR6UB4Tnu/prTbRD7PPSxqZBTlyEX3zpW1pFleTrkTE8oCpB+jv6qRrwn2+BLxU6
pyZUIXEX8HBPzG9tWw5nIIxCqlkCaa+pwkp4b03aJZrsyeJDI2hOVQNSsdzTl8DUWcHM7UQcneXU
JMxz6Mmp/0lYx+Cmr/JnrgNAU5WaLm3pxFHpXYL42qT4bWa3u87d49+0UofCip+1arxENITwQDPr
KgA2prfEJpCfTzQu5Az7jLxqNjw/WxyP2okZ8kgsQsSSFJkRipWNfO3ochuSMeWw1wkC1oWJrxVt
J2oO7L4pcDAhlHZPUXTNUjQt7uE3gLLqtKeNkLSEF2JqFGHMPpcqbpWekrZnJWfSgJ7TkkFbD0My
LTauajWUIzHYJxsg4UGgUjGPuZvNuFmqW/g7/ZNfk+xVZJ19uqqqKWKyU7OvVu6O3jYp10nZllSz
lZnRNrfBDAdt3ssHg+4Chh0MlqDOK/KsItfiBrvrAe4wuVV+3add0vIuoWvx3ASzzfO29KxpmCKI
amCczAAtZ/tjoB8hx+BAh1tut3C8rWSb3xbDwtNs/Q5Ds4bbxVT/SdzATVfS56UPISpIeik/7pHJ
3sL1qIZ8qPTz4+oE5Sn+IkPnEDHYTBIrvYtpiWEJD/IbL5Q7/3wtf4x+xgaBqRDvblwQMXMY3FQc
w9ogNCgoEWTAGRBYekwi7bZMMDoH8PKUsskWREj8db4dfSFFZnM0KRGX9lkGjV+1IePb6K5w/30d
fPo+eOJazwGSj/WQR6Gc/cwM0/B/I2ws8RJ0oj0SL1/AyhQtGocYHYyE93FzQz324wctaegpDjTk
Yc5mpK0+7H0Vg97KscktHfBYqcmPtIUNYZa/v6bdBhWtug8+pkudgFoGmFJCIi8puzx/0KNtyww3
DYOtR34Osmw6UYaaHlWlUNJrUeDfaGhK/QdDrB1CDRHbOGAfYtuj1YId1lE0FKMMRL+L8gLAMFQF
Lej5zV47b2b8LGV0AZr2khXzok2nn1nZB6A/w5XPSDfApLypm+ft9EvtXe5uczSwPkCFbi3YnOsO
Cvew0yf7vU68adZJdeD+Ov8Ty/xYcfRRFC+3yt9jzuTREzysfrDI86gvvXVJVJNBZcoFamYk6Quh
4BhakWxWZeIZjs0U6OTkZ8q+nzwcYDX2OFBz1ahbXmogCgXLfVYw/TzwgtrnIsvLOfYat0rt52cj
ykwcB7+ZJ24bfU3HjMCBdMTzjjhIja8kaBWHoU+HmGc+2qoBHMyDoNU8U9ndf7xtU4qd23rVMDFD
CbZ4sT/mRdhdX8lbQeSKxV5KmFS0sGNeNIcq0wTX4Tfv63mvMOfro0nQj2LKR50PM+IrYgwjWb49
JYLrQVZxtYbsoyIiRo8IxD7oS9vgGz9cKz1ZK1A+IhZXExeQ/UUB0JG2W8CeoqQzaeml7e+dRI6E
7hD+dmt0ZkGRypV1VE7ppVPk6wG/tUUGcoR6EkNYc1ItIvjvvP55qnwe7NEFrC2Wv7OqkRP9xACU
4/tMRSf8JXL7Z2F3oVrKAVrxfdDb945/wUB7LDymidM4EPfikPkY1aXavrATGSXMSAHEfG3OhvjH
JeabmRfuixKTTtLu+zbqLxEgeQcpXSB7WmCcpxZ+ZMNzQ1oWQkWdgkmoXOkhfJET1a+a4QT/x+Sc
G6H+zpq9pYAkM60DvfJtgGhY5YGbDO25ZSL26bd6sFSy/O8AwojlBnORGnfPezTYIsQ8or3Ko0VG
YvDRKyK/RijU+kvbogz5F1/0SpsOfsC7hQ5boiCYlI5ZOTgwd4PglIFO149zwzYRoSMpIRZh+bMg
c+gshf+1VjJMeHQs0dWbk697tmU9Q35iW4kxE6iuNvwRUgeBo2By4xqtRqOfe55EpODM7DeL4pkN
mnfy64VbGrQO+Ih86Azau4cg/nBz+NTf9STauKx3EoUuLX9Oe62V1tSdgqTUwnizk4fDxb2XY54Q
wHkpLDifo/XiEMj2eMb3IprbHgbgIlzPK3UvZIVL9TyguwJSNL2gkJfuOqEnOhWONa/JK8RqxsoA
RQ8EatbgeFPKFzved8tNlOJBmBKO7ly/AbTyzNMZS+Ham1UrIS/lDd9x/lC9Bzg+mdy7H5fPAvoi
48vf1MUC1j5xMo8OhILvMbNoNlkR62Xvk2/ZkTIczMXe8WWJYSVnME8Ba46vvQH1KXoE5ctJBW/H
S0iUUOrCSaSCKyWHbdkRCXo6QBly6QNCRthAlx1jY2rnn08GaqEICiNcp/BIS/BxnhBL20G8DGM+
7b4SzFYCOsFdxxea3BQ3AgsYypDxhMnFx0nCFcO9GsK1vIfMko1DEzLXH+v+2h+7OxyItgg5fYmd
hWYxIvKGmBnJR9jZTNpYtNHMPE2WylBFyzY7bre5ISQXBKj0L9i9gwyB2ycPUbxWuMFZLNWzMgif
C5/HnkRTvxiOdFk38tMcCzT3nSS0W60uPFhImEamGNldtcKhEx6INwvKYWkf+l9YTeYrGwfh8zH6
gHUPCtmHW54dfRKojNRl1WkGGjekREqCKFJf94Y1YT/oxeNpm2iK0gOKqrtA+86noBXWwpwFVImn
qxlAsFLcfOrB36NQ4M+nfDYnEwOwuLhwfE1/s5xiq18gm/3gKWb6Z+edybojwaqxKL/UAOccdlZN
AtruHbk1+vFpl1fFVAUwJOOh/LGUz1SfiFOTTXveiUm/DDDLEITshbv6c9RMwOxeldMiIIsoksUY
TSLhI1eSq8RVbCGkJYEl6y5oGzkBvA6u8Wkv6mL6dp3NRUZuZ9uSq0rA0l+4aAc20UsIVkIm3IDS
lVc1CaBwfTTKAI4kjyXzYx4uWgXVcGF6wXb4FrjJsL5oeiBqF/qefySj1HJdzFfwOd4bN7Z0Qx0p
5vjM9E+eUF3NjlhmtwKiC4Vyt45jGJoLATZ4VXx1SfBYpBZp+ppxuowFxceYe4igg3IS330v79Sa
TPGR0lTbYecT9p0+Coil1RuugL+aluqNp4mhXNfeYwhl9kWJqSRbD/obtLup4EO3HMJU7CZLwzm6
zrqU+MW5ExzCOQQCR0iLv4OEHuXzG0F/Tfq8MrnaVAZ49PKloxnp1Jzck1xlLBz32pJo7gbPyKcu
8aK+RcnhFQWpGnAf1au/EnhJBUIp5jGbd9hr4e/tHLfeSIz9Fq7V+ZJy3/9AzORUsESDV8zzpalL
zbT8Z19ea/73R59Hrhhim1AHPt8zjmx59PvaQXRzdOn0eRaGrxijxIhJN4Gu2HpEFcF77217UQxy
qAWLxPS0ccRfNC+rL2J6PypBK4EB9g2H3rQb9c0/wVdWC4ZaqqzOPjz8WMVRy9s6L41bUFfOowhQ
73EnfKNzDpplohVio7CWNEb3IZhtMS+afzrYF9xbUvcHvRlIQPkWfux9tXhT4mQKbpllbu+/oMaB
bC54zSoMggteRn+VLKeiZXI40UaWjrP+x1kkdMkoSMTyVAUIl7kszMlEifNeo/7VZIeab6iANfhu
h3CHsThh5kAHg/iy+fJ+azaBou19jES5Z8JCUmOKbFbpuTccpC927utg6XgCTqLOplqhS6dVkupM
5FhM0dWILNsZtigqhXYo2UibhOpREyevINhVGUSSaY35g4rcWvlCRNX5FHam5REHzWPQEuwYpVAh
/pMaX3D09mOxGAZUBpbVyzLMrHlsYm/5ZtRrlZievyKLbTrX23UFQ3dJizos6wg1e1wlkSOaqyCK
j7njeJT1+bS0FBfteEv5iCfrRPUyG3A26wgm17p/Ak//zIT1SYdhL0bhgU4Wt8X2qVdDwLpT4WyS
/aAMaF4I0+7QvP9BlfdN0dJ4zuniZlsehRHG9aoasmUtxLcpX4x45W3gMzz+g5t2IEVkP81PV/Kv
Ym35VwgbUYpOWm5G6EARsKAF/uux6OmZ9MeZrVd6HQLDF43um1vBU3nQEa8d+SbN+8jk2Gn0l9o+
Q1oksitTfuFM+TaBrAq2hPDCP6QgpS5ImUJseMtunQ2emRXgyi7sZUpT8fcVzhJAxbsND6+0tBr9
2a9lKNGnivm6+O4ffQsSJl0jpUT9ucy8gghudhvMDwucGurZx6/wp7m3b3YHWi7aDlE89PYNgFJx
NcNR5pSxWiTeyLAQTHRnhtbVVlrpMoMUORhp/DNuSm26Ml1uRBmWfcsK/qYwGc8XB8+APS0hW86I
a35ruFaAOuZJDMQ+MFdVQkGiBfQzV5wX3wffCxvZ/mpU/UG3I8QbW6NwMi29VCGobi4WbGWPFftz
x7+8iaxMcQ3KnRK7Uw3C8BP8gJusOhmsjonw1aqjncfvUS3Gi8J9DjkUP7FNa0LvPq1jdGbzPg5r
8Hm4TyL7E0ONFXQlVqXhPKx00HgEyGEbgfo+3nON8vTsfVSwfsuA0UK5QcuCQrLeIvgHLf5ZYFoA
kSFdeqIN9ltnWzXbNyW06B1MdiX++OClq0FfpGtSq896ubjfQi+RBKBTn489hEU3dMU+C9FBRPPH
FZzN/fl3ELlspJ6vR1xhuNyDZV4YBtzluS9RVQHrIGgaoSG4QCFOd0SyFsyhLLD43MFgdvtbN5NQ
ShJ9Dy/TX7EFpqxkGxj688jV3kw2YV4fcDAepCEboZSqXJ35T8R3DqE2P3zcKxh12WLq2Ev6zzZi
+qPII3ZHKzVJ0ScLt47YXqVlDz6tXS0K3EhdD2BoBiJECL4aFHJyn2Ggx4ABQ6oU3xMqQFaq8lel
Ubz5OlVmNXpc3s7uNF5N2cMR2kuiW8QHSt6GV+JlqHcdhkMKp7toZu6T4k6CqDFkGzHvoK/FOguG
ro6aeCzytvy6V9GNflIX15VrP4SoWSRt3K84J47wohpHrdXFu+9vjG+PO9sKU2PlxY17yswdvvhm
Uyb/YP7Cte/zygxrE+dMRRzy4X3dFAVodKZRqQYBhEJfhdZwpesV6L8jew4ltHpeYWfgq7hjpzgn
XbKMb4MDjYCP+lXOQC49Q1FBjkS20tDg1j/GL05PVFVKP9pocUwitGXJPlk55TmmpIkO24jNGb5g
EXMKSuWZpGSSR+Kca7+OJnT3qAX+OMyTDF6AxjvnpjMOblEGR8rRDjSOsJWf52n/mojgjldTyJYW
x+AIPcPIJ8dkEIsE2DYsn+W5Yn1uJvPpq9xmm+30Rl6PkzHqv15IgipSaaYxaYsYg9QqyK0d8avl
lk7QgdNOkm94lZ7K3nAbKawaA8Z8tng5L5fPPTWz5hZD2QfVgBHjkfPqALylvBnSQ3VAg2HBHfsp
G0hZvA0gQiht6DimD2dOLD+NKm1BDHR71c2APCk90yMGMFPrYUUP3oshRV7yVAXNB1g6kSlAXUw0
nUzq1cfHfvts3DXt9949qgODgXOtmuHLZX4Yf+kyAACP2rVL8Gh0l8Aven3eZG+33WBeXcu3R+SP
UT0/NaVhRYotOGnvaunG1VG9dRtxNkVbSbWr4fpe3glqEzDjOyJTMRkTWOk3cTR5yWQSSE3YJp+N
q0bgdr+oFpke0cfwW7DJCJgNj5vY95SLLBur2luRm93LLEzjvHuWwhbJxECfohnPxpRtryy02RGA
ip3p+8du2Z57eJBHK2EQGjpOCopM1175r4tE5zUaoSZnwpRaZlffjgHlTdFsZfbPhsDCcuThjD+w
tgV6M48TwM+Qtp5gfrmbkayAyWWMYK5l5wt1BTiNUpPXQAlo+xuyiBVqOIowobUbiUjZXLgZtnRB
uDf61QQhf6yPB1brI4SGL62dg3frENrFPBeYf2BgRe9V7/P3V4goODMucW0fF55SQHAFVLGkB5or
8WUe8H4DsfVc3SMiubQ6w6FbR2YG+gjv6lDNc9W5KimcdyQQvZS294UXzHgsb2zhUgxThfyBcjd3
SUMnXFg5cEAVz84pPtSas6dplKtq+MNGg51HsPXZ1azbA9zZzG/RKyfUSPkkCfUJkUc3sbcjRe+Q
fuH1xx9HQMxQzLLDQvU4HNJQqQp6CFr+nRBj9VYGmA0w5jSzOkA8S61evxc4v45fR9X/UyAalGXN
O7RayKBy8h5/JW6wgguZN7rwl6fSHoJ8Nqn+pCQtovEntLfKW1lD+pXt4DMjquuPD0TKm/kTVGiS
b/387oY7NL81wXtIykBwMO2nLhe1xj/Zh6qh10lINeuO8hS5QK3U8MomgS5vwspiem5PY5Y9HqHA
7YMbs+/ZCmbyq9VCviHCFuSGsi2umtWcKth/Y76mrbzoKKUuJP9nlZBqyIMv8j5F/f59Jo6Zg5+0
vYa0QY17vaxhOF4H21o0//gyQC3NR5+fjqed3dI2QcLJl4iLFkxrmx8VlOABiFMu8llur0j/x6oy
m61bkbvFIdi0r7PuLL/BAISDmBGEBDuRaF0yxTS7mvdHvU0GJg+mByOM9g+ZhR04t5mWpUftG8XH
06RUurqC20mLzy42ESWiLmfR473O52JScl6i2KU27gtzqKGzDoebERWRonrOpJiJvwRHofJ2qYgv
TKDeRRtSqfrWTjOSwuwPldWyvVWuiyp4uCWTZNx+gMtlw/CZ9MqplN9ipd9nFWqE5RocQaLbsJgQ
CqUykudaCSOCMvejIVnRpCGBLAJCfnuppDQhdDxQboNQVc5ZT6/RV22kypyNEewXnUs66CDx3Khs
E/XFB9HSihukkz/l5XKqyV53h+kJxSqQtXlu3rU5CBROc6O3lAiDLmDQXOtJ/rWAriZKBofc2kNO
MxDLON989VqF+9Pkw9qB3DLMQGiUrdKwXyRWf8d6TF74Er1GvBIRRtdmNNZtY+chqT4dwI1Avpnx
90QHPsmmi2RYQEv+DYZtXPltW+07hVeqspO4hQQCpUCr4iJbKSs1nMcu4xVqCO/aMwuRQqe865TG
vfFTcs1/9245mACXw80qZEB2B2TdySy29vwAhQpbF+8gPssjoGZpv260mnUuja+nw0XQnqRK28LS
XeVgKevgvg6lR9U1C38lW/wzG09HIP6L6o7UquUZtpDBrKPi2Vli2AP7lXI3ppWzl5IcpTBRgGlF
zHX1kSfYtcfFyUkwOAtv47UCsB/Au9bu9FsF2qruCTA8pbKYxAV614k5aXD/RS0qKoJP7uajkDQZ
UdW/yuJmOwqeLrEb7Y74KcOM8a6Czwvp29MJNIop7Tpiv/KxVbzW+xclWKtQgajYUPf7xQl4vu24
3zxJ4n61+CxQeIYewGM1zILEg1Zlf7qCSM4FLpU/oNu2nxrxi/zbpfLwL3YCRatnh3/lhggmje6w
bfevVQXdyRFt+cksxllhpP615bG7/Ax6zgKImhAW5MU9jtw1a8bvOvZgmybeuGYczIl9mHcWCEKf
Ub37EwUAXqL+WMuDXQ43iKIHH2SOYJggmZA0YmiPATgfJwRlJ/9m11U6TdwJwgiABc1HHQ2xe2mR
ZQv3JS5YAPBhxBdWjAjuFfN/emBFGjoQj28KQmfdy8Y80hsgaQ8kra4ecp34R3CaB979zR3JfwN3
aALN/TMNspiQAAZUd8f23VSpKi66EEf0yNkQCO/l3AdkE1coe4FLZyEtMBdcHnI49LMFfWkvN/E5
gPKEXm53JJHoWsWiRLhYbA3a6oX1U4GxVFhIbQZfWo7WEFjmOYl0sVlyQbQLtHbTqiEu3/0FHeMe
LV4aExLj4CWVP/tJHJHiNee2jnB0mimH1CQGGIleMoIhTjwpm99N8GbJJKc0F19Fu2i1oTFyDgkY
GEPFVlQDuMbocOPmOUReuWn1uc/KcEgkgsMAeBM521J7m8rbKKsTUHpToTs54vUKfuBk+50IgILw
aveabx8defWGPuOgjhviMeAclVcV7i3GxTuRuX43/fnNxSBJesb3EqKLbsGgeUzrVgmlPybnHa7Z
1uNy+Q6Qmnf+bfEyn4YLP4FD47mMzUoOB8ii9rgpjh2VA3Ay3gcg/YKEJ3N5nNh/2eHPgXX2Sb1F
NrGAJIZOXB6qSVVh2XJZH5IsLSD4uLVg7hjisg0lsRON1O9f7EmKyK08AtCTESuJAYaQDLrnatmy
+6So82pkIqS5QhpLgVNwDqL91gMfO5GEeG6WPq2u6eCUrOqCHBtdjNRMd7c/IBJHNrBqS9ry/cEH
MdjjSQBOETFkxh0WNO43PS/orJs/G5LV0GbKdFOYn4EENRx+CBGWYcTUbHwZCR+g3db2N7oXCmEp
BmwKu/PMn/vOJY8EknzGttFtFvcTfwX7zmW9Y92xVn+axkFAGTSUehme40qcOqC4CfECawypZ+Cq
cRO0DE1I6KeD6BE9G15vJertAC8ZaKoCO2HREBH4OPT0wbpfUiq5JcVCFrl5UiywbbcZcxf0NJzU
gWZuZoKkAdeQ9wC4Hgai0g1+o10IdScdBJeup4/jR0xIkhhXItTUPO0QkA7Ss4aYwJY1G6spmScW
cLeRn1ZWLBhDGjlKwUwSdPB3+auiKMbnqa53DEyNiVnadUT5lP0o2CqnEv1AzuFM5dSRQ9r9Tz6F
GBqxGrqZ5WDC0OO1YMs6LVuqkhu4keUwypN+6yfUoXnBVlEmtnax1S4RdJX3r1oJQ84hVy4dumYF
zUbkjFw21/H83CR8eZhENz26hypMG+3qbuZFEmJzznbHKzqcrUUD1jHZ1A7WTdSHYenijsIStqAD
1yaxyjMyv+J1m/BW8Cz9hljfR7W69gNSGNJCGOvmW9OBDaR0L20kNlnJt3JOG5eNp6URB89OK+gQ
VuBjMkpOs/lLNW7jel3vvbq20vR9QxypMqjMtaOs7OODNyG/i4a6vRK0Cv37MqK/ZIc94IxY4P4c
VHj6LtxuREI2Cm3RjRm/43vebKq3jQR0BZCw7I4M3TIVk/sv0IcV4iroZvNpRdpPvuZaXvTBnS66
NzImOVN07Uj9GrhUd+ThuTLtCX/7j5Ky9Hpqg6Fe8vGS4PRQILp/tc/0gbHcuhgfm3mc0/cl3fof
JUkUy6RwsS15K5xCRk0wlxUCQmLueTQu9DaM2yI0J99xjfyABGW18mDEhSrusB2sS6/cABNeB0mZ
HAnnUsnc1GCBSu7ceQ6Dh9WPx1jv8HE42cxvk/KBUX4rac8DGGvNKqhp9Be5Ajy88lIiQfSYKrz9
4mzozIWsCoMCNGR2z0KH8z+dmXKq9WF4SPewkSkiBOfLED5D+Bm0BQiiUCGO5ffZTEFhRkdpCsa+
xAk/pWeE6J/TXj30C2ZztrkCg5lDLsaWGEsL67OBLPLR0rcfqLKBzWvafg4l2VTggtt5/BIoveNC
0E62ioJvEU033eIC939+PRpYGUHmyWDwfXXUF8lWuSGdvoxWH4oqZrJZ0C5hcSebwAkQXEZmqGaa
Lgzlv1ToCSj2VXGVnPjv3D8ikjHpgrUyPSPqzYnVShpN7G6m1BQ+WziU+9MkfB4K7WpmnLdFi7wP
sirhjmz8PwyyTaB74RjgbzcfnEo5AadRQgCNI3YlKV5gH2IysDeIB+BmwRh5x3yUSA6dw5jj3SYM
ozWs9oDZ6ndbxe99yoGoL4MJzfRxZLd6+mK2547EBxHdUM36jSsXHej3Xv+5ZEBh7BdEPjNk3ffT
CEao1kPpwmhhrgnyitDonwoV9ZfkLVU4p/LyWvIWWoTf3bNusz8Pxrhtwned4P2vgjlTu0Pb/ymh
tLX96rzm+shVDt5Lqpe1Mso3v+EKIRevq+mrURanWeStVIdDE14hyHzoWseO4B5YsJyMkUl76SsB
Y34UOAZFsJwaSKbL4OY8zCvH1MvSR2s6oZ7SjklRZTStBkKa4oit23qq2zOLtfAV/tQ+4WMax0yS
l1wqKeyjlGu3SIbapbsSHVAY0w+MZFt80WLlZ6Xoxt8j/fqJH6anvWauuiZ9nbvFZLgaQIUBRtZa
hj8aNEelAPXkNgUvC1pfjTTILB/ReBI0SQCyzM/e2zZtO75tPHU0sVzoLmjKKF3OeCB42FlnficK
+no1nFe60PFil0PudyBeckBDy2vA+DAoZ6NR/Aj+GNmrrtnRHpCBe73r6wwWTWYmSDR8/U6YybuY
Ad0sm38DRw8UBglf5QhD5WeWSMO8/37HMnylQLHkSs7kL3QBGCQGDnerTSMqyLPLI/1w23x0Nqn7
qZa5I3tC/AKXfk2bEcvot0CH/z5ckh4VLX9qpYovE2/sELRjMfaPpZJ7vWv9CauQ+gNF1XORa29U
uwskrnmYI4HIwky4A470cBA6mVvLN7tqoOeCH2mKZFMm1OtoAgKZHhKZXb76cxmUhsVDKUp0XEkh
MxX0UNpFjRkuqPLhkzlixCNlv9Ks+/lcO5KCZNzebk45FhQEP6UXegaPjFDkIM2olrHm1bgfL423
kVYADiU4WFdzAba+sGhQyp4fYX/RvB/8ceDHXEp/7kH6yYBpTZGOKYqda3M3G03taUz+4cDDxZ56
Hnp6AKQdPnhchWfM3MWUTKs286fTOCW2YMcC4oe6hLEh6KurWDW2F3t53nVCQt1vQqmQtUqFcsj8
5hpJmokulPG2nJOxgQWHLrwtSMkMZg2GkDRc+U74dwY9ZMMLoaRzKgNe82ymmz3sNb/ot/LFMwEA
umweNCYzURkYj4AofukVq4lgLJ0Rom5Vn/3OzTwJPr5lrFusw4StnTE/rcrE9pxfMj2kC9FPUU/9
zwQKWg8MbC7GBY+/kEqJb9LlKxC0wRSlBPTYNkYwMt4vOfAiQDa/l12YGYAPWud4BQ54EAZ+CUkS
eWyZgriL8eUjqvEMfAFyegu9rtwgG9oz01yxTBPShYg2mzDhXhffss6XeyWojvIz7xdhIzosB5J1
G6OnAccQYJP+q9I8++KtMcdR2MatMOOgxbQikB4ci4zICitq/Lx9+Mz65U+Pmn9lm2Zf69iGG2Sh
AL3ku+AspAhiVtW5MQtgJYYfy0vnCt/FyDpunUCMDsVOYOOVTDJ1lollBX9eCkkDLA5EFGehr4qy
vOUZ1l98DBKn0dacRmHxbmM315jWBiVd3QzCgvdChHOj8ZFjY0wlMy6IK4u2Cy9d7fUvlEaaX9Se
AdZjhe7oZiFztuKiohcpoPI2/RwrhS0E8nzX7uj3H5OzJ4p51uIYhA+mstEg/WWedrjz8io6ZibR
KhFsLuoYMkR+T01ZZacpXw0PHoF6YwywYTLfTGv7USJ03qzp7CJIU4p/PpRQuM3CIgfjz4SYQU39
zKsO9y5wxJq/OoaBHAA2kIes32PeOBfiNaC4A2HaaUAiWhfVB2FwaZvJlx2pQG/REkXIhpG6jRdU
9sFxzExV3/6ZqU2cMMpTk8XwMGjLrKi/NePNL8/DHklt06Ek3SRy7bBWehu05R5+VlXEZcBgPTfw
pL/BSH0ohLnp97QO6C5EgLVQ9C+9fnstE7ETx6bF9ODzLCiaFEwhLhs9H9b9aHjabz23QGPEkRzf
kxK+KczRDPUrNbmhMk7gXQwSg4i5O+0o2JWiJbLLiz4IXzemM71TZv2JuBUq5bgrNOvCojtDVemb
0p4clFIN/a9AX3N1Ppjojl3ViG06WJXamOGHTtuxyg7JetkC2hlA5l533n0MwEpYshYReDCZZmxN
0hWHBNTrs1M260LtFOSkYp/DJTosQDN5LWu5EtJBd6hSlPiBlMss/N1iqZdS8kueSp/O0LySjvwu
RlmA7S+CGcv9dif6RHASk+ESEPMz0nscoSUE8/xVZXrtUVLMzH7REPUsHKEt8Yk3lG0EmpTe5KcU
qFBBfDBX1vqcFvu3Jmu2TVTZSp9Bg/Kj4HyoP//2uTGgIQv49v7GEsXjp3gFyAqKb52v4r7pWicH
TYty4fKGlNsOIbjQSiqRfMlbQ22QnMDNQpR57lckLvBpbvQLsAHYX2f1RkneQpGyj6qAGlLbS9GF
Yf4/v2B9Pf88FEMDgEtMTn4FTvUr0vl2ycxc7gIlSL+kZdFGlRNSOweC5CvKN2xOFP1ZFVIY1b2K
LPfl/sJKAHS09iA8nG15KHjkcYm0e0ABAkz6bQSVHTCKMhG/MJrOHdyRejR9e3rr1Nzk3DWA2YU3
ojMTDdsGGCwY78xJf0zThqRN0dILHlmoqDTMC7zba90gaSFHQVinQ3FFn2WhRz8vU2+dequNABGd
1gxksnGWr9Gra6g8+J/sUjC++dvEHJnG9um+I074Xkg632qxM2Kwdw22C7EY0XB2g3sf1SBrBl9d
4R0t9fbvZk6vEXPbKMSQhYpwH47Cn6E2WOcGP1guIaCVY2tUWgMASQOyzVqmuTbgDtDh0LPMDzRa
fi7WhftFMdDvsX7850nz4NaFnOkOxssYqNO8CRmdch0kQJr5OBmRpjJ5D+1Rl9HG3f2S75YtErlD
03UXuqhqvsjkqPmdQJfgYi99yGrREkOd41LI/rgnEjnkSojTduS58zQT3dpKsHW1O89ibWn3MlbU
yQY8GEd6VvcungoVazlmnHrt+SBDMcGXZr/rmWyRPYYr+vkKOCyIsUItyBCpI5e3phzHRtnqEJpx
r7qBYznpEeiRFebuLrhfaP/rl4kOpdMnvt4vMKup8nJ2HGg8QO4jyD1swXI1FQ/d0pXRQmRX6QpS
6RitDcjZMs+q0eimuFJ2JgYj1+Us4v9bEvEIY1KuC6qjhs23ejgGtwg1gqXE9bFP7RFvTppSU5da
gqTEUTxKnyZdpyHyZRzLMYvXe9IJBHNU1FuhFHK57US6pAi0fPzUVzWOSZVUETjnW6DVdOtPwMzF
dEBK2DVdIg0cThC6J14D38WFJ2rpYZpiPGnYf3M3g6IVEzPGTOrl5gyFz/6j0HMI1PDlo2Taxm+L
7BIReOHcvIVoMYDEjaxTHIBSm222M0Nwo9Pxaps4ZCTj
`protect end_protected
