`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
U71FUQf0qAsGxfI811Hw7L7fy3nJYTd83JjuLrHeStKqJTUSdPESLymcfn/cVpzfBW2bF3BmYXSP
e5wyjUbgzQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
pWFieWO8oo9hfHkPbS1OEKBGvkAlQMLueuSIE7bWZbT6M/kqq/dye0/px/MdG8aHt5pikgi/t4lz
LuwJbIiNPyrhEa+tgcCOd+vb3cYReHlWv6qj2tNDsdeIKt71eaX1vjVYrragxGzIIBpV0lV9r6kP
KVvXjylDR6lRRoIz//M=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NL/pTlSg2Og5yC3YWVrNMxiSfHO/GibZQp2PQUi2R2a4HnjEylonymvH2vL9j8JouAuk0EFB8tc0
FPakv3CX4TojFCd8gaptzO4C8j2m1/36bqI9Uf+rv6QJs4sPJKomGGlgn1W0EQ98otaSuLPzoswO
7QVhIzc0r7KyYZieWEU=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iV99aGfQcwtekMk3L28+vYpw9Op8htG6fuBIg0zCTnTsG9RIAlgGEYAJA1TMbtP7znscQ9vJtEfT
T2W9slLueLoFJZrjCE/mxALz1CAlD25Ec+I45Zew3XrwE7ALGx0DdVLFvX6rrGYjjDSv4DlIm2VC
6VPRrT0nE7FzO45hOJpJqvRO6QHlNl9OA4qb1iEgAVoqUDz7Q3O1w5yurrFPSx5RObMnWO4Qir4o
LgFRirYZygtHGrCnsFsYiJLWkp+GPNATT9pDv2lpM9NKbSvhFFiGIbQHHydyE66fjDOgmN7gsXCA
UeWavj8i30EH4Fxe6GGfWT0D/Qx7pcscNmPo2Q==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GLCbDl+3CBTQ9mXi3N7iILMMdha19N1H4Xq77fJaHrjhhEYWFsrbEcAlCnAn2Kh520BkwISUGiHX
qhiC60l5dQBrHwPyukWPv6JPp600q2D4tTB4YMXGX59JzIzkFA/QrfOga9Qw0wCvItdYTofCqKo7
eKX3lnG98TeQJ8s8Na7clQL5NcFlbPxzsDOkoCF27W2dAEoIvbTv31NrWkRzh6kEnyUtVfJH1NWV
FG/ORKXULCX73nJx5iFYlTmU7C0VjbqKgPj1iuNvkn0R5JLIQMAtS6mdCRMQoKwPKsaF2wBBoBYk
2rIlVV4P3Xm15ZXC0wxW6lucSgd9Cn7JMSmKHA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wqk2o9IWswI8gqaghcvLi5Mb1OEEF1yuuxRzIAnMyN65arFFPQqZge265OnuRXAV+/iPV0UMsEv6
4dwyuTpRDf8wwbS873M0Q40Lco2/Dam5vuo5sBSb7YIBHHVlW8FOxDEzR9E70T4b82HLX09gCGbS
VHCF3MaIuKHgKOwPoM7xio+IRTmw/QcyxV+ZWxI4gbBzAdJw/7w30WQHXTjlOna/N9/0AC/gf+Ze
AGeCmAx2NVq7WHrX30TUb5uYeV0v1qhZcimC/tGQVg88BfXc/+4efXGKlwNimhMDrAakp9u1bwsa
V8i2/qUMV18HAwJfOTbqZhmb1ioPKYJivmvsDQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 103440)
`protect data_block
tzM02eXxYoxNIN8ZckVIvZNbVYmwmssHdTDeP21oeH1KDHSm1rwtojeIbe4QfTzx2yJ1h+X0rTDC
gfLtAnF7Yxn/MxqzjguJR1CpqX9txfBCCPvs/yHgtQfXgnO8HAVTnMLXrbDSC8QfRjRWUAZ1WiLZ
XS++LHoBmB3+NO+fMnN0N9o2NtLxkaXHbsLFdWkEzo7DtepqUrF51Bkqb3gMMMWsnENsc2GfMUKn
zY/uuuGDUzB4HpIU6SJ2ulkt/AvuW018uRol1iw0CUsyNfkM5wkANCK9PZ9CR/uA7RARrmwl90pR
CRBQMakjGNoj1iVpLlREGDNX2SfFBEun+nQ/e7wumH5rlTNlX0uxJdha/7kd5jOF8Ic/+jHNk1Jt
6Rqhm8i0pn6qsvYl65jF6x/VXI9eBHR90OrtMNpSAtNsf8auBIDFKBytusYQljZyGx5J7F2kGpo8
FqoczuSdBpw5Lgt0wu1xozsLonbcH7PIlbdRSFNRSTJZ3j2MU+1A+KgMv9yIHBz+jTVrT5ApXCLs
vsFHs6EbZgjKbgfT35NcKtk7sFefuY3HT3fm4ZTAJBYCVuh7VL9p6/fof1id/8ISNAuIX0OoCwSh
GZxW0colgLX0rZ6LWeZr0BCDjw+LFrC19R6P93gFaqdKu4BPkdCrkdKT5432ckYbDgIbRZ6mIn5P
FB4jv9wRpw+uBjmhaom7Gebbwj2AjWIVhak03I8WyIgcVGeAYF3kQ+n+AI7OAddE9ViLx17jXgc1
yYpHOpYjHsk2P6Mp5h9B/AJNxc+2TSLRjGNsf+WW9vGyXhXmB/lDcQUMq2Nl9TMtSSjEsZIJvaW5
7bqr6Iyk+8zBFpzyLK52/n0npBqalw/JymAZy6KOKMXPtAXV70v38RVNqvoIwmdwLDvFGXytTViv
Mq85U1xxQjuUFdIgvOPph56aLF/5ZxEpHKaslBpLEr4myUMXeALqijUaxq5GkBV8QxFBXXsk4Zog
L0jg5Tr7gyoArkLX/CNngu5S5IgZecleZM7If/ijG4DKRB+B4tQas2i/2+J7wTceeLJFA+Ey2+HF
ds6lqIAR9JUpB90o2GlzQByPZx3zFZJlhbNMOoub1/KA/Giz6ZsiD3yOMiUuqBS4N3TepP0MQ2qO
0ds1NmjiVmDJYd7N2nktavRMAGmaRlWglJY/3VpXnBcx2vVdJEhLsGw6xUf6F6ThTM/zFArOg1NM
OrtBWeG0bY3F7Tau/2Eb5Ihh7IC2IJXSL1GrlA07mMy5wDIsEnzhxfGOIyhMpa5v7iyHgWF2/1Uw
yBUHd6Vy6Wr9yHc7DqnejlQllw5mD6uDFTzlSpIZFcfg+EvpPwTCcWLwExtZMEdaVu/YACxeyuNj
+UGwdvHvyGoTrhMvj9fEMxJf2uBKMMVofW+nWVKUUY14VD2+6CO7W8fLr6o2DlqDc6cuhaMQWBLJ
/F9i9n55hdK6qborbdPZDj/zZcmyc5J0yFLD28gzbuzw5pzXjirm6vaJwHSjrDqmOwX0z5bx5OFa
oZGnzw/Ga/+BOV2+kyFGreP9mo9n/Npeo3iUmRsnJO0Jo5n9D3r6jZKdpkj4OtWbZ2rO41xFwtw6
/B8JzQA7Tibn7cdu8ebfwXHo/4aL7O7eLjnYdtayFXHFeQPDV3bBwbhX0iYDcZpCQQaUXd8enE59
a87PE1ikIOV1gsUZ31TfI6Jusf6PoSjE5SaqFqGXBJX7StDUPgYUpbBhE32ar+CqE2b3xkhHzTQp
olq1uGfx9lq1BUlUIK94gnefA+2DebtiMJ9qMKIcJFQ4khAfW8WngqZo2kx9tOok4coqppkOpibQ
onea5LArqNwZeGSaKm8VePD8fYLz2SAw9HVHtA8DyUv5CzsC2FZ/nefzXz6KI76MfplMXsYRBC18
iKSFuBitgi+6uldy81W9n7phLveP7EX2eFAgId0LFkfvV/RywFvsdLSE7z20YE2wNMhDNl5RtU4E
R3+jtQZqjSgCpGg10ugbJhur/DZBEOYxVB4D2qC6czvQF6NIaYVc/7Y+Jw+z4ZSb36qMaULq249P
9gpbja2e3m5b04RFE83kJf2UPWRjhUyerBjiCFtJeovEiAV4a6y9NAh2EPEyG4ulYKn6RTK78cYV
QTVzpKmpg2dv0ZzwyrzOnrC1iIVv7c1PRjw/+Qr5RYNhHHOTYnCtmND0oCuPHUYVab2Lw48csFJS
qg8W0ilRUcHR2EODUoEwthveZxok1iqo4EqByZnCqovyl2NHqotDiVe6qvgnEyE0f72mTCoYdzCZ
d5VEx7MYhfCvt9saNV3NlS1skf3pB4dtipu5GjBqRLcKgVvgllj78BbXsjDFyeZC/n0pAdb67CPU
+lr/PdAg3Dj/DGt/w9ajBxsd01Sl32xTYJ9OECwZad8yICtbQTUtaOSVli89inQ7v4TIbuM1LNHY
+W7CjZ3pOLRY4OUtbdUEOBrl48BKydJaiwmsJ9GgQ7leyN0E6IK3yf6n2b6Y1yBWG57Z362Ur7dR
ExUuN5bUX0oXEY1bEaNQ3OV20g6D77orHHe8a+tkT9HlbfLl+W0NfpE2xh1ZVZINbND7wqeU4P7l
mZuvN4IAE/4A2oEe8aUjC3V/FPqAC3IziTPsesjkC0NRkl58BYQyeEtw2//fyFexEBoP8QGnKiO9
bRs+K4e5An59kjxtu/y73NHkooS0Ruvgc+Fwrn1GWhAeetYf0CR1YHNrK1quQjJAuPoGLVV8v65Z
F2nd0kdnZ79ZmgDyeSwByV1KfdAq0mB+HtJvwcqTM8czFZKVvAdEraxJdbQQoo09LItIb0AxbMzP
KwI5j4m9X1BeotgZYkOmqRxcLg/xbUx0XeD0PDToHOLaNtfKr5fTsu3X2wjyAYVvw7VGkbCku8Iq
7Qe7KQ+4NXGOJJSpEfkr1rVlxYGgEcTUeED9kT/dfYuGFAsTApFsL9Z99O0X8Q0Up+6y1i41SbRH
nYEnWzTWHFhJ++7vXi32ads3eGhxoNT3QSHy4BBVEYxMitF6xgFCq40bn/6sEA/dX1ZK4uLAfx/p
YAxB4zpY8KELUh5zWunDAXsjbOpmA8FEjlczW0pVbuF8vG9UusNY4vtUxxbedsKzPMle63sLl3l7
Dqw8fLQK2U/5OeVc/M7dfRGWR8zYXqt4KICeDBgkbeAecBKkA9oiddbzn8ejQgOn3/7SQ772rOSi
rw6Bg1lOOwJ0bEBftAHyySjJ4chEnT4tNWm2Mcsb6SxGivxMtRioFgYYlzr2aiMtFeGUwqCIaEmu
+JrW/ysXko7QP3jUC/kvFyNsEQ3ICJYwyBMIzWEDhsrqXUwyvmLwml8jN1C/QvuRZjSx1/FdsEva
TL0QXWT8DZOpMhYokIbfz7AOuyHxnDUlpEQcmc/KNVmeodoW+77sRGDGTBYplXc+whobxrcvew1L
dqgSI0lP7Syo4L+hxap2G6LZlKuf87NaKIPmIhgMF2n5SiD6jHI5uHwuZploPqR9ZJsRxtE9lvLw
Dsbd6bF1aIRIH0DUw8sRvdMMddZrndV9xQfzZ+5LtNZTYEaHXZMsyVVaEIOK/uVBxzFIQIye8MBa
tQ/Wqe9+udYcVgVDz8LCsen4ItHooPfu4bULuJppubuzyEHNPsiMeShXsWSjHT6iEMQkB6h/+zYM
SsL23rhGpL4uBTTh8S/VIWtj5iJ7tXrfc3U9r1WUqDDYX1uBZD3jxtUacvxT5WZ/3a6sn3Bnio7b
V0j6pu7b89HpJW9MDew7ZHl88mH/gnZ2ThgFHLzznvINQD6uY7xJ8r7pP9wcDMH+S3rVKT6r6A/y
yQvCR4C1QhEx2td99XR2KCWVC/yrDY8F7xzb80yFmGxBlzJLNJzAUWdRKPl3Ogv9mGXnlgmUZFrh
1QGUyM40bmB9NSVAowHzSSieCB9yUe37y+7u+UYafocX1CuJIkDd58fM5broZ6RtfX+PbpgmC6+7
X1fjs2eG1UpXj9dpN4EA2ubI3Cxx+SVhW5qU/0Izve24kUFeBfCI2b5+y7a4fHgkEa4N0MZ8QOBO
YdKUduQNyx5axVQLpWd2GtIpE2KbTtXk8FlgjY31rkVU5kwUTWx+bzcEYYILgH+yqEw0+Gco63fc
Q3l6p/nQYM6RrFF4Y6SKPTP30+2ICOL/rRayX3mQYO3gLTDvTgyklyxq5smCrjOmxTCDtjfVgjQK
VQTiS7tSyjCROYRMpy+G2AW625xMFgpp+GoYCmyIBSnAKT/HdPSmXTreXNCULQMq8a0KRr/7Fvur
egRwFJfYxk071jdfyyu3AwGi+V6g1kZfycryCebp4XIXMac44AysnUvK84H64nMaQdEDL7yYqwx9
zihdC/em3y/JcN3RKLhWKbOevVZu6mF/oikiNuIN71+KwVUDDVI0+SE7Em3HSkNp+W2TH3UTtcjS
508XhzBWw7JiJASkmVlm1jUV2VgcLHjz4Yd82Sm9dOOJ/88LMysdUgCE8S0ETZb5d6VrW9Qu9BaM
yzSjkRQD/5Jp+MxpGiDrFnJ/uQtGUWb6m3VU+FMnxTlvQMhcAOz2oOGZUQntoYYyNBDIQfPHwifw
/2cAO8WWHhg//P8ur6Kqap1ofONlFJ0texDQKL6HCW91OavQhFTXx6rqPUEkvqx5mlBuk37qqXEt
Gx7pLO9e827wyhFp3yuqghQVhkvUBpw4hW2XTJTWw/jfmd1fef3Zir+7ngpzajMk3c25qhNISvFR
VPXn5bpropQo86NRnCx9+AElSv4AG5n53Gbg8deHfKsu4j6nGDOPuQ9xW0XLsnPlkZ/KHj6Smy+3
2QDvNQlePfbTUgl+9h/Ry+wQChMvY3abIGxa3+6++llj/03qggP3A+d1Prg9ZDSFdhc6hYxs5rtV
mLuErgvBG/FC5Ada71gCxCXq1zLIXbdw9Mxk0GiKb37sskc/jcW8sw23VlVoe9o/3OF5/dj4nr2m
C1o07fb7AzZkverHO9WaOdWNaBMR0FKkJXJGB58KIkFNWRbuOh7wUOnweRVWo6tTkYBLSA0DiXJI
q2aAjE/jMoFi2mA1EU2oMaG581NSh24KWMTHWthOpTk/x/R/rVmrnQx7m8wnWsvPlr5vq2cISup0
fsJzvKe/tLAFaDoPzZyDHNzpmovjr9CI6ZYKuqmb6tmH/Cbg5PkqIJbIHMiQEgr29AcP+h54EkHv
PZoYgIuici2Cdg5Hp1Taj+0QUig925e2u23cqQ/FjCg7vGPWj/KtVjUXC8XvQw4/U/tnugejt5CM
8tmK/R4KZa9ycQaSBA48ms6XJxUcvT5dPHL4D0pdmTHoTUINYKHhz0vwzN3JFgNWr/TeVg+/ddq+
yO4awIp4X4Wgh1vTB/yOhG+UETMnznfssS2DJ8BPuz71gjTrbJJNMm+C9hDHPtYsxP92l4nnwkmu
5L6k+7u3UXTvUE+1tb0AQiNqlQXBoaCh+A9RDJSjvhIK1a0itvZdaTRBDtCe54MiC/ObQM6biXA7
uHfUAMXlFGfEUFA8vdHZ7RzzMcwAEo1Bcol4LyL6CboEpuU+W2I3yOdANPSfCZxRLBNgiu1Dp83y
fPjckQbDtBx+ouny0HIX771K86rwsXoR7G/qwFzUJrmxmUWA6pDp3ByTiSL1eZeIP2tlYz01RHPV
QsgFWaHzLFcmdpzDRL7t8bBMPUHtaFbqfEFdRab9ONnNaEZ9MZSKT2miRqFqP79ptphaz/pDTe3L
9VXrijPHmxJVlzLIGjrcNUa6mo+JNcvbplwMYzF42V4kODLnJjanB7/Wh7LxaZdW9vGihE+5IvOh
QNrgYGlfmKKSkCF5soHw9tHVT5qSCgqwf9sHZ1GPaPXwzrp+Gh8OLHkhQkkVpLDxXktVt6uKAmnP
k1tC62W0OknepOXjsctzA7KYgxs5N+ct5P1y6yPu5hjBfngtZGubk7g1TWUr3X5zYJ5bHXVp+1oU
TbablqpyregWoM8jqEbjDYtTpZO0yz1txl+Cjnek8wUpG0ZGt61IdAolQXFIouljeNqGRUDN42m3
7DX9keVNhD1I3W6dl4PGzJnPDYBwDEniyR1F9btchQlrOU+d1Fi2iwjzH7H9jvIDgzXjc+MfnM+s
DE2ZaDF4GFudSD+wofBRkZhu588vKdu0KBf/ktKofzGKlQvA00sJ8P7sxQXefLhAIw0pphYYdiM5
05Wv/KczUa8p8F844gh37+uJa2/VWoxF94MRSxe9DlN0sX9Tgomz0Y51tHDV1sHknHmT5MmpWiQV
5Dy3vQqlKkJfSvub88zP7MAPx4kNwNHYi188VPX31MhMNnT0djQk7uwAuT4yR2LEAH+3jQKFYuFf
iC0pPfyF7UwWN9cUTEA2G1i5nRGCVJOc+UID8dGyOq0k9bL9UaORvyr14xt7RojvNPqpBbFSB0BZ
X93GVILazKF9b6NhwyWLtdlcs2vPXy4pjZzngPB0+L5ClVH2oVRSzhuu+Zw+sQkr4VpNXGW0nkq6
LmZQzd8OY+CDsd+UkjfRKQhn8JHfPon/Lxcy4W3j6fswhHLe7N3cMqF738qSDXo9xnzn/3ksspoq
VTtQWOlJw/VBJmOY1BPCs9Ow4bwpyxIh6Y1aIItROim0knddMpYG4+lZg4C6vTE/XePemwAuf9XX
SKRIbIai3Xroyp2OCRBaIGBL4NmEsrPGfNI4e+T2uzQGC/pf2oqThDggtVZ/ui+sA/+to2EUBOJZ
0vmwL3TjyPXNqYOzGz2DvrRWB5Lx6FX90HnXOT1R1jItxAkjq3MoIAv41IXUSgb/rs88qd7CEExU
8r4HfVj9/hNcpCUTKgAS+YSzpRu7xO9adNn5FfzirZCZ0KOw4bZMNN79TwWwRCdLAN5YWNDrenn+
7uE8pB1rqCwIIU+BOrbXiJAqftdY6EPzgqoN7VGvYKYlCHb9gTm6MNHLUWPUhQzFdMqvk4lTy39F
FK+3tCyFPus2yRMnIYdGzMmCtzZ+jocmn6Z1yY7JHgYX5uB4PgFDwOIFa+Y4aEb1fdrdY6kNV4Y4
dcrhnXzktUEG+7NY/Wi/6KByN5ZzTDJva1pW/Ow2fo5fFq7gBf8PfpZp149tluGZNWDJM3OFjHAL
N8Pc8zTz2r3G/Ry1xlR3yOiQ7JuYVC4izV4BNz4RrvryHx6q1k/edO7aJsIJLiwFyuBso6iV5oFm
z+vUDhHqgwNwlJL/QdfJrCYIeu2JTRG6a3KDywHpv+11QS1B1YNPcOy4DMvVbcGHaxH/sSl024fL
5ZfJGlYPA1N2lyegK3gbGQTMl1tnwehW3gvLeSHkov+HNAdkuWShJDaJpmlCDBDDUip55H59Gph8
IPoSxdPlSBsiOXuODsuZ90z31lQVMEVtIBC96IAln4N0KxwSFBVMynKgmSIF/ksi4t3nu/vxdP4G
eYFbEtvziP4PraagPKGEabmT3UNs3VwtR44ugMJDNTsOCVLPxQTz/fEekParkb362fQmUWaBXVl/
LHwNuQuprR/W91BTY8boZV47xqLQJJwQ6JxqpRAW0+l6uMO9/s3DaYHGEOu8HU2HJ9VQ+ZdYtPdm
r8+drnlfwg/a3Rmvfa689rv+2gVBcTd/ECT3fP/zdXPFE4QBJrX+xUODOKxa/VyU/cSJOeumhp4G
KCmiw/AN+RGjn4HTZxjA3EiBoDh2IEVcEse99sMatGZxRd5l5XFj+h2VIKTbU15j9zSKlSqqcXpd
tR82C0xBidd7iAsxbvtOrbCZ7t+Nns7XTxacI9BKYmFmj64pd2I7CYzgye5BwN8JVkAVRjcPP8DA
YyRGzjw2Hq7KCIWbB0GSZYJa2uRyE4wexGRFH6HN45W/P7J7BWj3Fx/qvOEW+aCrdgUI8v4benz1
SczDI+uG1tK9U683wzZ21WJ+HRQFRJB12Wf9tmeqqKogAn5gIB8WP8VpN+artHYmc3urYKPm2Q0s
wXD3xdyr3yw5Nj6lhe99lWjADs40CbCwOvXpOqGJWrZy8jivkfOSpBonlgZb64bRyEsYMLg98NGo
A4q5Rabss9d9GZbMkMe4tih5TJrS4BxDYpg7a2b/EuAy2jrRezEiz6vO50GpP6av5HUcyBCgZq9Z
LL1p0Pfwazcb9oCcuCYZPedXcqCgKMG87Dom5aifsQCF3njlK7fRLAbrZcObFPWdd6uTJQcKWL5v
RaR52aZectZXyt6uoMiayOoM2zluc/ol+YJ1jGCya//lMJ8Rp691+T+SVvMnM+ehN4urZpyBu9oD
Mpf0qGahHMi4iafsFSfrj9vKNDVhucBOVAQU1C9QY24sX/yulPIot3eOnfGgj+p4otB0SxGFtL+I
tDZcCzH5lyhvygUYiIWy1xvN3lDPcoCmBnDIJVT/yQwz6yarFXUlNAMZDiOYQGwBYzpUD8s/aB4Z
maXomojgSUGVURs766l3ENt4WK5wONRpi/XsfnXZfazqZMowDirIQ4G4SlD5XlTL3YV71aVbHsR9
sHaKXruzwZjKHg2tG0VqwzbyBMAwcys17fsVsgwWtPm19yOcLmw+qsUj9BpXR3O/q4jIMHh6mLzi
UmfzD54taxa21xgH2dhVvd35abFeGzSzv3GZTwPYnZo327ws1uK8xCQpdHCR8fY7l9s6A7OdNUTC
wR+qsu81ef6BCGoZTOP6XBnnNG31nJlrtqSENvnc3ERgZ1gXUs3egBTpq/1Zl+IKSuAglTz7SVMX
UcgZdUvvNgA7fCveevx2daxkuBWqrXYynU5yc1r7yCKIfF5aJ3O78Iqy4wkCWTn9zFnb5gXID1Z+
Qxlie1NvZOPWNXjVrWNtEKHC+quEaFt9U1sV+3d+pqxagsLKRm8MDQd82Rha9o7Qi05Mzt6fWabe
+0y6uwKjVsgEbsliV9IeFPb7CJ79/QWI2hJ3mFIAUj1/kGFnsFzbXWJdlnk+ibynprlNl1NkXQrn
o3490HIaFwPeyPeRi7NVFW6Lic4rKa/rS3Noshe7OTbVpVhimiV87bjffzhR6FOJJJZwTw4k+YiX
0yE7ID/7YmIMms4IWHCxhJhrQTBse83MvcYeeIfHHAD3szWGNSKxcBVcC8tiUpSAoP23vq0ppRz4
alAZRhWI2zNO/42TvsHBHsQGKq7Q4rvAhsANCzdAPpEkfQlAVJS9d3y/K1gZk720P31FCMu1rWHy
dsEJFYfFWpe7rCc8B3+7NnC02qXeYHxKiHquw/DL0yTk9Nfr4uHYz1eSwHIubRoEn8HSAfxYZAG1
i2q464sIIzna6Fr97hcwd/74iQpcDinRrnBpo503Ijt5SC6n/0W8HgV8lWWmz5Hhh6zhL3HQqF2k
9RWA8il1yU6Y1nG9E9HiflVy6/Nop4thUJnRZf3RNYFRVmFvYgrgQaK6wEtgjCPbUb0aHel8Qqu8
c2vHsY+LWZdHXMLnpVoiDcVabMa2I3kkDQ0RWhoSP9WMPFxb1U7+QqqOtz5NcWf4aCnqMVagMMCf
k9XqeYaXDESm7f7QrofjBjUUy0BllDzj8+2v9WdDZ0+c+h5UJ4MYhSQWQovMNg6rx/wIzf503qAv
fUseonihVS8gB8MXIWwmCfZQAVLgyDaIlDJDNgDYvpYYzD5Je6A26/q1K2/tjQoNkKI8e+qKa7vC
ewtvj3gZdYdkWGvyeIH7YkFmSiI3FhfhtH9i+3n8vqR3NkBZdEFReGIjbTryRTWHOtK612jKuNpn
7dBx9eVAxuDw2vrJ9hNyz4jAT1ABiK1JXTv4vfOfhWkIZ6aCJnUF0hdZrT5kibUmG23eXj4adbXh
WXFVVYGU6IZoezdiCoYjv/jFG0fjQ64GcOVm2PnE6xyW1o+1z65oY0/t0Ocvhc+r8PmWf6NTZD/v
VFBn+1WY262OLiKnKrLTMe3kNscNkt0MQzijbq3vz/X8rAnivlYoZaOXhnJP9I+j8XZZkrdefdzz
Zg8+DlCRV12U9jOQx3fr99dGRuem+0ERc1CS9vzLP+sh3i7kdIk4os+ZXxn36npPcwYxjOvt19r6
iNlBoafcJXV+zC9tmJBRN+iIt52DPEO1jqgIOHkztmQPdluZqeQkg1y0b2UOvdifpuHmS1cqCvCq
WjE3icabB5RnPCipEAilBWJyVrdiDbrVcqLPoHLL9EHOrmuwui+USRIBLBP0pIqN/j//mzAqSNDk
IPaCoaq3Frqvy1SFsDyIRhDj7m+a27E21I5EO8gXlHk53Cw3jqTr8i4PTRxTHn/HpYTXAg8b6IoC
pq+zkqxZ+DOhDZsFNWkv0RtQYVmVrkqkMfhnsFAIbslIyZW8FxNFA8Vw7xEc5d3df7xffwoZ2Rt/
ng9E2Zg+bOavSdAEvEmgOcRPE9ezVJtEMwgmiGVYEyHJ67TZTNg+2uotFreORND2JGkMVGi5AMiz
wXs3JAaQitfUPa6HYgg/0x4QqB+JYlnkPH/7Y2ZZbYkwi1j2IPhc5RviJBXQDE574ERpIFBFIoiI
p9Lzc6GBKfobbjKzVLQe/libvntnvLUcAZ8TskEBbyfXkqRS3TVtQ/k21bbjsMk4CjD4ChY7ulYj
Ctc1+rb1grG9cvjE/tOp2etYvvPm00sk9Rb+45/8MJmyv015Oei30n6dPmslbV+v7CTKDTTYXPTS
ryDRYIre6/uxQfaGNQ+P7gPUeZ7iU8cRwhloEm8Bm3ltgh3JdHzQs5GHt6NjTcYREA/aJYUx+q56
6UJPB6m3MUfZu9xK1CIfK1oNKAvNBeEf0JtWQYiZdNJNetslegtaZUmVwMlkoM5t05XwK1E/eP1v
2FW5ya53/UokkXjh1wAlhXCkf7oCs3xh7CBbxrmg+TqUxNdcwayzbxlLScpkOfSpMe06ElFdBMSC
VaIb2DtwFT/LjkWsPPrrFVwxnsBL/5MNTp5lpi5v7r26O4JDz36F2gqdDEqPRUGEihRJrJUegDdB
nYMGZIJycDckmGRiyaU3wKpJVJdEf2iU1zoZj1Gz+tRWtOmlyB2/Cb/a1GcxmwI7aH2fzkOf36yO
NgJr8mlzh4iicgV69O2tYYYYgrfNs00wEQ2k08W9klN97iAgtDB0a2ERkad12fuqjRkNrYQUO2ca
FHOuaJIVBCDhjSTWgy9F87MssaTU9wqnDxmx5fcpJWnojP23nf+lBUqbPByO0HwWnD9MRxTLUhpn
0YNLLv6NeJq7GB91g9uwUKU1xVoMF57hJcuzBa6H/Dk+6phzyD+BHUwuCFjj8y88QcE4YvipO3+/
kBm9irxsUTRLpTsjo/ds073yxd3W6QcPqBtDsAwrnQwgTs4VhR0wOXATDAsyKX6g3BUjsb3lsrVL
bycF6CdyBkuDkmJJLjMHeGvb4rj/9TqOY8xSerR2446bCZOgsJGksGAKW1SdMoymbnCWCYjgFavu
GI0p1+AkN/lOt2UxDdZwWvNJpaPi7y5cXHeZQW6cY9u4divrF4wgj6F0qQsmZ8F7whhRoetIJb41
RnsLZyZXyWPu9b0JEvnjSq9szDeuBliFDGNMM1dXO7mWE15hqGVShPq7wRKfgrGeohqyD4aKA3ZD
8GK7cmjWacr/s35IJEJcKnZcrSq193o4b7DqizYRa7FjUHajWB1LEG42tlku+DHr4DFhm21AD7Zv
XC+YCGbncRbXRTBN+lkOd/dC1slPZB8qkpD5RO9OFMSVEJx/MKOKnKdY6dFy44Rjm6EDCrqoIicE
JXhoWNJygJ7AHxcRlQm93Z4HYAEAYv5nGh1NXNrPiWna46fEyZ94pRJJj9UWunL6wJgfjNxNpW+S
NAzWMwwyBPb0E4pzmT1TFCcBfTeY9kCMgCap46siR2+3CpCUDbkiRWafhdho54nlJ656x0XfAgSZ
uK2HRGmkh2Tt8IQU9e22j+9IedDPzOLQGDEOv2qahTiL9PUwXkUBSZPDabRE8isrNgCZAPw76elO
cHF7XwMNK/8DIJjEGOE39UKfItkYhrqaTwrr+jl/HUQUcAOsl3lMJVPBpKC/dRxfjt5f812JK80H
cPdvo8G99uLq6wZ2JD4Hf19rCprK5UQXxbVIDVEX/PtEfwRlslCia+2OtTKY+a/80O1skwLg/SMy
7Ab7MLpr5YMXrMMg/4fujn++5swG08B9lTC+FVVTyomCKV7iI13pjJDUGqg4oeHuz+4BN87oB0W5
neo+IuKJc5sLPzJ4qfCUFFWhcC53+uAmMh+1S9KDLcvHwlvbEZmMG/NIAJFanQuGA9txznk7PIFD
c2etDYdJ0AM+/twaTSzDKACFPiZryVwZXBpPldekAKkZvZ3WDGY+DhuatmAQi+453pBFL9pMIRYx
60Ydap3+GIxsjwbJJ/NYSVUTLIrUHL5CeOsSQUdyLn2wBgzw7trx8hAuE3+xeCs6EiExWr33z8rp
jf46iu479KuILQt4EPWzBOxe4GjB+dQuhMzZmPJd20MLT+p4DuTrl9eMub8c5OqshpwrZRYLaudB
/1Fp1YUA/fPxStjGyO3aOnmpf9dXtES0QMj88hDYssFtcoetDVwdbwK5DYfLL0Cz7wuSY6ty8le5
vjHzbLHt4jtDjnNGBZzpZeylUTyiMj5SQ2KU5SkMi3Cy2Q1h9zyguHyVm1qhr81LP3PQ5ht4mHXs
Y/EDocVln5ABsbxN8GT3AbPyBoQv99yMCkQuWLDlOMrx5iNi7jIfk6Y29kjY/qTUt1zkDLNVvBew
oqotNY6OHxapKWowLA8yC2qu8JvIbYb4Qx0KEWuAzEP2n22WvpJR6nB961C3Abv7xRrdVdPoPAlu
xQensZO4hxwlefOLho/8zECSJsvoQ9rKyb7JGVg3Y7bvE2bHYesZyBEiR76atzy5+EVhw9Wsa7HH
HyrkAO+1h1UWEoJeoO2qmizOG6GJW2qOjburyA+4TjKrsGptm19noj4jUgvdbWZxiUbjVK9txF7O
Nso8TnIHsiefLi4Fr6s6vvzR0CsGddR42txhShMz3C7GTiVnFpQpBjEFf0EuI1J+6PanSwMOIYVc
7jANTiZd8lT8i1SUAaMwbvZE78inOq0nA5eZoTIlS3tFKh/3L4yvchsQ73NXOMFXazGW6BBHJh+E
qgoIoTBETJo7PoSnminT4cHPq1fyogy47aGS9kaPKDUeWhbn+7/lqUbpVcoAT/ZOLjJJq3bnVsqK
+rLpexpNUlzgL3gwwgJ+OkuNoe8J+Fa+L0OzG/PSFbiFQMvujtN7+5IODU4/mrKl/j5WYn+coPJq
Vwq6B+Ea3gJwrJz8VtiwgOM7bwzrbFo3T+jsECi/9Gg4zF90IjApHaudbCoGDbFb+JkBiBvZFrg+
UflkvcKXlIth2cLBYC2jDfjUnvUcEcaP/lvxooiLsucK8Ft60bVzz+4Ci4+oBZQK/KukwhOJ9ZlF
OQVN6gAFtnBSVmy+mEkNiJPRrnr0tDWy93zr1hBnu1x/LsEJbCRzzUtEeRoXIJaPh0QeVHXoVQIA
T4hi5j+NqXJd4/zsUG/odptJh7m1Nfx+bC/5I8CFWWispnMl501jZ7JOtUJTozQcYnr4APnzpki3
wLdD53n/obPZPeurjN0+tAyFD32wEcJqs1QlpZhDcrq6Pvfu6uJsYc3eDaAZ+qY4m8XO9NvlMAjB
W487V8ZWjSRmjAvfMHylGvl6s3mjkcWnzOmKwLdfUe+V3chmx3c0ezft3F7qOxFrOqOIcKLaZ8IP
wSGAl+7U91CKAMFMKJU2OJBMassq3EKwAxo+Mcwddrk2v4Jb6YeNDFMVwWZ7kaiHWpIuPw0qg1lw
2TjBHvyP40pVh4bOw6609U6rKBspVQX3tS0eFJfskkd7j0NilOkwdLjkzlG7EfHk+6paMXKY33wz
G6XIfmTgVWpd4l1TH82mhChrlbKRol6B+V0SdnHQKIiSsqZ5yL3vcpQs45Q0ll9Hep2NkvesFmL6
bks8pCMgobd5sOVgpfjsW1dcbOTOfOCHzDZDZMbbhi8Iw+aafse5yIZ7rJTV5e0fbxrwozjByyPX
COeqwFx9y446kofrFVoQFACWruphcJl2Udqw1aD+SEffVuvu7WnY2mna/FvvH7tqdsQEkkNgIlkv
qtXxKeWnJLg7SXdlB8uaEuBDqjQCryf2GrJ58PsIajRKnGPO3geetpUIDRUOvbKtAWfDUL39NLq8
0VqU14+OzCMIPffaa+y8/9MbPRiisjJXDX3myLANIjNaxWGyHXi+7DESxNJ4O1LaTeX8Y5qJdDnb
kpjge6vkcPl31pSzEP8q1Ds3jNlvrfQI0zGjr+GcNau9hEbWO0EQi6S/oC3qWZpKfD60aJG+NOU2
P6iipex+kADXsZbob/wnsuZFBZndjfYHk0KaU0U97y1USTs8ZhI8NLgVUrAC4G4ice1WCQM8Th2y
DwIA0IhCH6Am9R9F2YWykYP3vGgVQWYHffVjsy05SWqyB+nzUk9Kj4zTQ7nh4EGw1IZlgvr8mDJE
u/mI2+0yO0+XpEeiwMWYKSsbKhf4QfV3i1bqQkf0kjjztXWaeKJ3JroRi6Ov1OQAvPgFoe0woXZ2
DCG82y+wsoowyiFXMUio+byRFGhtNTQ1mhL7HAXYPvEQpg4r3/WOQL/huSRydctJBDQCpdUYA6G7
hqhO7zJe/+Fwz4Aj7EkCVBRXmR+9eIpx9eC2XgwVm76n05s/mJ07oEfR4JlkHus6V2Ub2ZzEmj7l
c1WPgfK1taM9Ts3JRUmxDb2wv9xDFjWEjh94yyj5YmrdyMSAaw0TVKDKHFH6LXRfWf42fLgSqkhO
jG8ZP8Vf+GzCevX/CGCSrJfcmxJAl3izk76uX4GOMbCzK7od/HKqTMaFDEN7qY/sOS9CjXLeLe1L
qaHH3bsN2j4ON7ujTTAxaXz9TxXccPY5Pd8O4Ap6oqq3m1Gw6W4mBKtBuAOGHrleh9znVpEgt6NB
YRWxQ49DmLn5XrWtUrWvRC4Xe/PG1jsOCiJ6X0QQ0Z6c9LT/b56KohSNNI9ViYSNO4+vrxjTN9+B
Qra3PsIBDyCDY9CONQtirtvjj3tNMcrc7OW+Mp/N0jSU113Zfo0qSGcV4eUGdltZONSwCN1rRLtg
9R5kyaqufid2+UDXpRhfYd9pTdsKVqM51pGx+GJe21kwKw1V7HCgCWOTeN8bdcOoiblndF7IAbwo
QSgawpKKVILFrO8KWhXyktDXw7gDr+dEYJjJ/tsszR/jCW3F7/MvUHTlyds5aF4RsWNCYmNE1hgk
zmTjhyXv1XQL63Bf6b3UEYOBNYuvhydizyHt4Ds09ybrO2CZIjV9CFY7cV5aOkqWwstDktatEUsC
/6ckaKQDSeziRtVcCqSbXW3HcEhTmYU9+qSY3UpxSqanmq4BywyOMwSN3nVJyqzH7r8++5tZVMP6
vWCZcOzYYFLeCCryFKnWFPxq0YY2cPOQIXFuRglPLWmgUtc9jJuI3k4+1SZhitD82TUcvTlxI5ez
HGUQju7xzmv91nkgefa0sSi581OTsuH/tuSOor6E15NXQdYrh6iEPp/Wl9wB2AsebYjHeqc67//U
gckpU/Vv99qHhcJilFkE2n5g97Wq/797ME9Df+kPNHC9vn9YVRQN3tMjzU7rC0jeORojOilh/kNc
ywqdoHubB3avRkf3mID2mY+80gIKBSRPczaeVOmkAqvfLUoIrOj8rKp0yew1bb/RR7iqUD1FA8uz
7iaZeuHtHGmgOBVVurAHrE4kazyY0k2looR3LmVK5CCSV4qPOFB/CjfF5k5FpNe35Yjs58The56t
7yrcWUEjwrVP1S1locNOmqAmLNp0DuC+rPyj3s1Kun/EA2GjVtdCGTMdstEo4jxQi4NbMM+1dX1X
iIE+a6c7lq0D/CEbU4PxroHjpCPqp2l9yAWwPVe6d1sPPSJgqwVqoPDpVrbD3ccdfqpyZiwUQAxb
EYIEHSq6CFmxaXI9RO5I2oi8FkAyd0x/G6pZLvGwa7Tro54E51oCY9uYQ61wJn95UbnZ5PUBM0nJ
Z59asm7BTeXrViD3wXnLh/gfvZ3p0Z18uL3RJpzymMub98oBDpEGmr51gQfrLZCttCDVXtFFhz07
R/YzPFgiyMNGRsR4Q4LN+mI2cASspvcoStYxeqtkgAwQiWGZR9Rx+2jqIjy1nPNJnet3UThsRRLB
RHdhXVd0eA+ViZFm21TO3/+z0LYkOP5AYQ6B0Vz6yn8fZ9fYqwTTGfFpZlBxLBquoOewawlJz533
0gufCmW9JkPBZj5KtvpAmsdXdIoFhTltP4t8Mhn9TsHL5BHp0rsEpo9eihGQKnDSq7j2yVfXPhYc
Jfkst/NIcaLssdamZ/N0KJv6xJqVk3mrdPOdtgOgQug02MpG/OET6m+vg8HFhZDrlRIW2xNPEfUx
sZ/FHZxSs1Rr3C5e/4KPz1NUTXZN366ORrujq/kRCV4Fq2nAg7KHEY5ENt3+6q6B7abiM3uz1gqG
B6ebOUA6F3guEfztHg8HvjMz1xj/ifZ1l/Fyrw68EeN594cEsxucugkAMegjjILZ8zJ2yGfXJ3yL
cPoNV3a1LVZHFETlu7oejAQzzAtCIrjebx8SGNjjpduxaPHTIQ+GK4+ncSqhsb4uE4ZtBF3pcoGW
Gbcf1wMtR4vEXmDrU3XHMFEvoE2aOXSd1WGnRVJpreUyrF2l12tbWthl7HbxBtFBL87kRStdVCYr
NA7C51Lds62ejbGbRLbalYaV15HyEQQT7rzUm/3V2Vx1AypeoBxHJRH3k6utGSb9/O2sX4THaBq+
pulsStchT82JECNHO3CLRKFHcDMlUwZV5+jg2oya4ZKiH/O1U4p44L+BihmyGylXLNBF2fbn9oZA
6pnjlF2cVHhrogDnd92j7XDRr2iykNm65Q+OVriPnA7F5gYQPyh1pThxm/uGTKwGPo4rN1vQ1zXV
E2wsRDGDN16lqiayTKZpPjiuAlo9bjzdfWmAeJAbYMsip5reJz2cXSUmHUWuMeKYeBUpY1RLK0uE
JZqPrPBkKOftVmGnscS8B7oC8VLTmVU5Dcv3YyqGEWYfJyP2NSHUGaGAWfV66V5OpVmReSNfV5h/
X5shl5LICaCw5nsdbKJj5nkH0eH2IlOhOPB8AkSLmsua0bauKRayF9pWCDU4gdJz788gKAU7Zruh
psgTuMhGOPs9xE7Uzr61oqS+oj0Suq4aRiqEKMDyuHynn/VpTF52WmWUJcSlmk2sxtSXpy1tlK5R
D0XKZWY27/Hf0q4+CVnRYF1nzDExZg9asv51JPrJeK4fyhxXWYLXEYZ4C2w7KEkKRMf554vUAtTM
mZ9pn9y/Oe4of/hlbyWWSFKtjmdBGDAjikT/jJiVd93U+u56MBIgci2Ag7b66vSlkbqPvuBiV6VE
z31yD8SWDpFawdfDVpeazgKISOhmDIFhpOZYRUsylzwC/mi/+LQw204coBdDarasEv/vfgqciYH2
FjkVylP8Iu9x3syfTvej9TWLrQTSHqzir0IJQ2spXwrHUlWfTcpoyavv8tLzB6QJuGvruaAn++7N
+90yLjQVulmeFcds8vAw9d0e6j9EdJ3C348aqYmABhts1j5wCf5jr6X7uHKxcHah7ptcNE0aocyw
F56qmB2eq0Ylncb7PHQXoXwtiVJ09TbEd9S0vXTFyjjV0P2xI4J3D8beuSAm+Az8oMrd0EwnVpQr
YyhovwJTUvsqiXYiRvYmSjpc4U8+1xg8bwfcQ052CpCxL9aamGa6D7xZm9ygAq9RKm26J2SBhBj0
whg5Kf+/0TkroIcbmN3um2QsxzCdQje9tFHX4kT3IlICqVKvbmwhJrBoXIvxxOVCsXrE67/vtqHj
1ikIUgKAZHTPP5MoNMZQh2bSi1CXBV0czizeXMMbnqWD/foucsMyJ4DRChLlFD8d9tqC35qeESLq
JTI9Z5SPqTFa43fmOBnWdoDS5agrEW3GdbOZvPpg20x5iHJUmaYC3M7ZU8FAVTJEmGCyK4vyzXNf
YXGuwscu2inWfdtS1txhrDTuZxZTU+r/l/qk+TTeKYWYqqfk7h7vNVuBhKZMh+kMbf/kSIZ02HNQ
BJKoo9fH5P+zUhajE1oL3ChDq1AEjaLFpSot1wyxugX8XmC87fsXtVvahMblKxP1FglpID5ef4rM
005UEQxgcMGsX6eFfUIe2qXzd9Ni2MkLKLkGhhhx+OwXrcKCKvg+6YxBNbgZkO55S4WSmmaZxhOv
IURwcIqHL2n0bSB8xnhKd01Tu3OwcOze1gly+WeCKJHz2FwhkAt/R41gSesMVnVkb3tPDjnwGOWj
PgPLAJ+qHkTVG/qyA+mzbeBsmapyq4MGTPh9AKHyRLhtO0Ut0cB1wk8mOHFYcYmy1PEv4zdS2MAK
+wjZAaspBUlbxau2Hjfkhyple7p4L3cvh0QlQNZ3AgcqfZtIAb+ZqapcfUK9pGMAqSYuP+mJd9KI
O2vVoadvzjwlJx9tYBz9bgng0sSyG0HOa8Kevb8z2c4XoHYFsuVfHK1JWgpTyKs6hjsckSfr7qMB
R8qNQRV3TwXs7QWB4P+BE1f2iVzJGJhxsA7J+Qyd5t044sqv2tE6hkHvRNAprM4TAN/SlF8Qgr7q
XyY1pCdCYOmaVfXbsEwkY51Z4GpstbmbQB3b/nr+2yX/R4VPnTPBtsoL0NjRNVjW/eGFTQBN/FWy
ks/LfG21kRZF9NfDiFHq2ZlMibSHXIFd/A4yp5e3sOIcDRYsNxiMJhInRDZ501lwXVxdqJ5uCGAa
D9G+YdcTSvTF4tj/cxrnFjLaCFdMFENw98kDRxs48DFJLcj2uWIDhIp9MAbD09Kz0CJ55WHTAvnt
gr9nr4RvyFPSgheajN2UGYcTN5q0RkNyIVNjKviU8qFiFwfMui6FDUYRjSbVTb5fBztUMb7HujZL
i3lMHmUzD7wuTuNnlyTtdIYMeJzAxLKzBURFH9Kx1RjH9kNaovG76NfKPIZ2fBdw37GRTVy7cz9U
5DOr/uyjZ9GkoZbd3Yw2C0hXgv7Mr3obXRW3WcvIIfesPa2wMnaUF7jSpOj27cYsJw2cmROBfaRe
OoNcXZn/NkFejEYya/Dj5tUweY/1ofl49ZuwMjQd9Eok/b4bT7osNAzdI5KnW2XIvjtknW8Y6Hak
JQT1JrqdARGajiFwTViUUovcCDotnYCmWnOOCY4TjpetodJ86mMT3oATMUFViHPPL2arcikxzhnP
N2JHSxpMlzmha4J4NaQTyahqQ1RyNqIXLIjUnC12UTf2I52agGWVgeMp2+vGSGYbFGmD1XURHuf7
T5dnlxv328lUtSIwB9t1bx9E/LHlqdr80p4S50nJVj15qR8zO9M6haC9/6OGhgsF0c8vEXKMsPOk
kwn+55qRSjcDsP8RT+xHg+HUwLVFnHgnxuLGGL1sQ/MwD43aL2vszrMbbS776PJtwQvMj3pykyFN
npJ2bEFOdVQEqk5AaOh9c58MrMAhGy2ALbW34EfIZOMXx9SxWsBIMsZn7b0QaKFuNL2jOw/Ho2qW
5zFIaLZtB4xa2xp/uGtXBiTCBwb9k3Hk/O5mQaJ5/nt5tUrbmQrI7u40tKzqCQ5X2m1Zx2AuXUnK
8OIXloK/da4wK3HYgh1aMGIqC06KHmnppXSTFEuteNZUmqhs17ZOJFKKc8jTWA4bJoKcl916do8F
44S7p4h4epHNbegucPdkbvC6jzja9ctrSy1ID1tKjgdrxi3rwdGpdvbWLxx1G2b3WfW2aToeKnSW
ovLyr2qs1uOoLVURJ6ED0FgLu9UPva3+w80KutKQcVJcf/TeOakA/W2P5jmsfHhxzSsbe5ZhctWN
sd+cc0KP3RvW3jgfUcjagOQgqgQpk/320oBKRxq1bBQMlkues8BDnA8CACftHHkYs0fJm/qoe0Nj
t0+nKMeWNIAE2znQI06jKG0xieCABFwgLyEFy4sRUf68ud/wHKXJ3xJSORIAUt/fOcNPoVkwxJ76
nF/p0WdfyqHs5T1MyE4DxGS1/g236nydzSkk5oD0TOj/0K6GUW3DBVl6WCcq+km/7Ge88Pcwam/S
PFBrSinQbQ5APzAlffismPG1Cp+8FCrdy6Xo8QsPPoFz4ZqnQK5C26fC4y+rbp0Jj1SW3fR9zpZy
5ZF6C16IqxguUvulryd8PipMdgWrTslwb2SN5wFZZSolpIgMxpI6tYCX+l2mAMoj0UQ6pXwTmHHN
O5XEE0k27tyW5WiYNZGolxJun1xKYZwuqtEoAxOaxCdH+dxZ70/cAvHGl+I63wfuNqujIqDI8kho
mBql3plquQi9cdBdFo8Pa67pN7/ra0KMEEViwPWLbKbhuBcCs1uohWq6mQH3TV5OfG3ZjHsQXqQD
yYaETQyuZeZwdRd/G+uooghXv52XOFqBFALD5MQik2Kshwk05GIUKtgm9yK5XpMVO9OzhxBmOrWR
P+vBmCbytZLzLfUVReIsGS33WFeIx8nb0XF9HHjH/PqI1jmWZ07Zah22tUNZ7oe/2ntnlpGSOCGX
OJ2r6NdPTe7YQseJYKPt6Kd1YSiXwWdoTDHvyzbigHoZZGGA+WIUuQ2zcQt1FQIYIIHunUaJUbVl
VvPiM0xm1EWbk/U+w6y5bo/YgXB+Mpcf0Kw9tCiKJnj+briCppyjBtAt7qUf+TYwqwEDDavC/wnB
uOO00PXDKiNmSeIbSWOIKnw9abdXcETKWH4/4nAOjU7+KYNVGDOzQy0qUcAMxbjBjlzVqyvRoJYD
TlrJP8Z6oppGTCx6p1nI0FZX44jl36jwZz0boGT26ic6kpgNP/sUcIreOHpTqcP3qvHw5zpH8mlW
s6sQ8cizKUU1Ore2sUF6by7+yqgAfh8gkohddZoNUGk49RhqauSh+r/UDRvqsOFeQ2/qytiPXAaH
ZOga8Wu5wT9b8M5phnt3cwr9bF6YDvF9hQyUaGXDaWno+vKO52/jaibNcBVrjtcrO8qSnjrFiz7O
uFTCJYKmkVBdEriBSfEnBunAH/i27kHYffc3Iw8hVHyA3oK2yqbqmikrhQFf0QXqoEwzOxPE9CPK
GyALBVYu5N3o073ipqmLj1kdA3RWIwV7bIe2KES1C/FQyCU85fLNsQ2bRbwstfP9J4mRfp9yWMJf
sTf0QmNy4EuG9X83GpEID3YgzS5L4mQP2lkJjKtFsGJ7e2JjIYKJ+0E/6trVRiEfWURsyvFyUZTG
EcdE6pxbTB1RbSbjfKeCcy6oK8l+URZ43t/m8aLsnrrbLVOr/I9SElL1Z546qY7H5geeVU+vK2P7
GEqUxtRsIvd1iyP6BtvOSuD/BeMI5DJnIc0X+g/DjbW8fXFjHv5FitsIMZkLEtFMXsP7EtznuIko
XlnWb/uvMmMxhf1wzwCHSwijBbyMftHx7Z8ntrDX5pt/DtgLE+27oCfQZo5TXcj2CGpnUxKQB31l
ZqRIgyL9jToKDq+42jIlcrM3hvil1t1SxBXvPW8mStd9/FR2uifqNeC6xF9ADcfIsU1YlDQ1ToIj
nEedqH1KPkan6q+gnXZHgkH8NFnpxo1PO99uOb43SLawHnc1MJ3DNMcV044R2+1GzsBBsddzIF6U
kP2WvX15PmTner6H9UwVDN7XNcGirqNgTk/zWE6OrNYk+ODQyGt1XOEIgaf9R7nuQ3uK/kD+JhmN
CermjX1NFivqT2CYdKiAyBN9BmEkzRav0m6fQfL88fEzn47XAAogmuqnD/xjBSxykYu6+mPON0yd
1ire1m34jQH280NI2MJ43066z9BDvwZb1wLDDUuxYmkF/fAssHLPU+N/JPramqCJEajpYh+Uxs77
ThMm81LDCYr8COxZIHMJELYoedIwH5V2Nb/Z1KQfX9TWM1ngoLbIUCGVh5yYGd0PyvnsylhbnsDq
tXzLQGDXXRV7so0uldJ83ogMWASW8FR45129+PwvH9FYuJll9O9wHzkGRnBPURCtdlN5sbLlO0ME
tJ3tsv3bxe0TFPGBfMzLXarFKz+CB929c6agWeXI4X+5eLXJzXLZmXgwNwxPoEcgEg6v6tYZriMR
a8nRbvXt+gaq8kt/pAhBb1wf7n8eCX5UWZ6bKMBda3nm/+0/H5xk67TP5kszs0/TMVM8KYpa3VBx
J3n0w+yNmaa6j9RXmQCXJndoa7o/QSGnErpkpBdoc5BDdNu5+wGit3IHifjzfVnpyh2EPyOp5hME
X2hbDTyKT4pMAas/IGsBsJrT79gBJLeSp06mn7reHp8YWoeRene8m9KQnGB8Z4rPZT+lCETwTzrt
GTdIF30NtnHPUSrx+DBbCXlLOFEkFUv3a5QpwD+zdnwXfFz50PO64d+5AjR6x68S83B2WGfrBd4M
LFHndw2FhwM0rMRMjcxENNyVpVt6m8lKQMiOzTuwK9Ar1XpokfwHwUUQA5ijtNTqseKyy9qQPGwZ
pPCWeNfa3dSdHJqhtX2XqeMbFKZLTmoYIxjRLte4cE+JN9Rm0qFfSbS3FWTIyngcAw1k/njDudWk
9K3WgqzeolTQvYx87j3FCZZEIb8exn+hCPLes/MCHYRYysgcep72lPAWFIHd2x7a25jvs0H657BL
8Ke2qemCFUzIZoUvgkX5v2Fd+GHCD6OyISkdxG4sha8HXIwHz5tb8WafqY3NAaLQ3aN39BSdh35b
n5JlRmJq5R1htyHbP60DG9FXNpavKBsfq1JZ4Ql2cDZGulXyCs8CcIUjCGwE6ZYe1NBVZ2evmc+t
kYavGtf5cuOKgVVbkkY4stSKB41zD29v+rLhUy9z6x5uMk/rkicOZfXcJTsvic0vecIZDK6tE0gb
ORPKDQDBk8msBGtyaeQGwySK6zfPUCmEESAsyuE4iOlluopXRFKUgrp0gA1CUcdgBFAMM8AUHX7o
9xwBoSnmjRWWekmJzIEeFqwqLbybdru4DvWbHoUBPfToG/NWs7NboOBVQq+X7svJ4RydMmmkn+z1
IIKNu8ru5NNDH/fb890176ZuJJa4AXVsn7rfOJ0QcYFiOCYIqoAgCqJeBYp6CXJti0X9PoeKyxDo
iYItyHvRc1cRL+u3B5L1no2THNdL9vmo6hR4Z+n2dXq+OwCGkwMms0V5nXqe06FRB3IAgoOjIKJB
KweI8QciuJBUDNgL9jxvvDs3mRUItf2rxUCyd5eL3N9BY8aoVevZKIWEk1ZkqBVOHJz6CixK/9e4
7jioSUCYZxI0Yd8UoxXAV66NZTIkLZjjqoLb6/ZHIKQ9hSo5wvwUCPpprSbCIAZgyOIUGrLxY+Oi
PTvkE/R+ntTYygCjR02DWzN/8FKPzJZ/T/bqsm/4RTJ1yYcuOD7DPCK1xDpN3ScFMcgj3IPAtLCZ
3Zn31i29EXMX8yVrttDwv2oIVhRmnP3y2KrdzSWOtaUiukBiIWw5OMxNBPZ+tl3OLgPox7a6p4vd
UVmMdzPb/CvEHuYg+svcoPDmWQBoUXflfeENwTwhfYbmJ1cFtGy4HOEYwDUneMyr7WCLbF0xk8m8
dUCu1q+mhxW5fstqg3m64wpw7CKYI8DuFNeKptJkBOytc6x/RQZEIsALh0iywKfPlHGSaK5RbkJ8
AnygFnBme/gHb0wlrv8oeSRwL/WrfPX5zzlJ0lyQEfS3nuTvhkE4Bz8aVDsJF/o15ClOWWIwx00T
D0LoR8KlNffnfvkKf/4CO+tLQEZFeVWc/0Fmov/YBdpzeHMc1LkLTl/jIcAm3DEe3vNEsO4Rv08t
HiEl3N5apQkVIkawIyF4QleklVpWUumZOBnWqgBWUXGXnkMIkMX/ZxqCUUjK9I37heo4eJVjGB7r
ldhFOotyKs4HP2O4g6OJbkk/MXrIPTwYoscGho36UfyKrDK7L2nnpS7hitYrrkOzbdKSrEG8Dg0j
77LpSMmoxs8wIEXhRhWgoN9s/gttANoRqCkgf6vvNK1bsSSJD24WIRgNJXV5nzWoYSb/lKbfGeAE
GLONu32NvI2OpPR38z7HI73C0mXuhhDAGkLQjqBLkbf/8wXjfWEnO72CmQgTemRm0bXXlq51vjBU
teBqu+ZpZaXnPrD0v3DLKzPkwzfBZ7SKVQ30nm7lKDoKhpADdoKYYK358OR46XljZIt8gzTQfgPC
+heBiUgYJzmTRz6czkYetY9zKLCCZqdM/HcoqXPUl7v6zfqfJT4aUGaxNfTiWJHV+rNxYdGtu+5L
kTu8AxDFueJ2pPCLeYHTXqDHbpP9NosfcDMVrg/ruCJ63+7whrdplJkm6XrqdJK8wMMBsSDNHWzo
g5J35pB0uKrjPCZtqf83+Y0wcv1zMeleUI3MLKty5/kLkIyXn0/HiYEOmI93cn2Xl058qaGY49r0
aTnX7jukHV6kSZvTPFku+rjAtx8NeU7nbRrAwbjBGxkBcmX6zO6dUs382zYs9DqJ2LpPr9spRw8Z
AbosSnDcGGPq8w0OLSp5wjsKWlrJ3Qmgkuie5Kx0gXnhzMP1U1zT+L9GabNEPdXu9VoBxL1a40Ap
NOi99sG+7xyS8ZWcrk2JDq4C657ni3watt/Pl6qBdkCJ/sieCeu5baemAn0r6Y1gCpxA7/oQ2PPg
3l8IFfvvEIXfcrq0K2PJ897E0+bRuZ1fBiCUu1/fqi40WvYytIo6Rt1Av3Yc789Ls38NzPRHHmyy
04nbcvDsZvMi/DrIujZlSv+WbN61a6fTU3Kb+tD4oandbjOn24zOvXX/h5UCCZm3fL1BQYH5Koh9
lvROCbz6FtdgVltiqLr6a4i+cxs+Ae1ErmDjfox1smWJeerBm1DkpwTB+KpFXwjkyOXyRcvdxClp
Vj0aFbD4NF+jc5RJxGEJrxijuIDG9VgeMVcVV1lzCtZGi7mZ4o7fZmH44ZE3Cht2zVF4rnO6Y4tW
spNTpSBUtAle9fc6j6f0qYZan6Zmhax/qZvx+3MTiDQqVBTsUUK91jPzO4e8LNx11kxpx4BNoJ/d
Vc+PRJSaAHzjajnIk3BUKwGHGDafYJ75DfgEej/vomJeSQ3lGFMkNHTX4auScb1XsHd5UvDU5HXO
HB1sYf6KVp9wNJHxjf0mf4maWeRUhHUR5bvsCRlZqyaJKDKptxagRYLF61PdUWQS71Dl7i35ygbh
ek+KvHGMuYZuQ3xC/RXPsZwBIPZXX4U1FIK+9cvY154IEjBNp4nfAsUo8hLNA47vcY6lxVCDdgCb
26m8oOP16J3yau0IuqRsvwBAGnbEAzEX65u1h6mgl+ku/5ORXq2x/uXjnRnEsGtxrtTnpj3RD/j8
Mse+75Q3gdLShBXxr38FUOvj3r6ZObkHEA+6jbD1Yp3xlIvRjvFaD1pWrwAkki0uJl668HZ69hcR
kJ5J5kpIiuhFfr4PVnEB5paTuiJd57lXPsr4Ng3H4yzU+ALueKIXp1Ah51lUBSPN1WVxjdQAXS5a
NKkeFhMq2RhxbIbJqwmN0+C6WzqdPP3b2DSrdTmH5R818gRI6NGkdgpUyYFCtZdYymHitj9J5Mwa
Ppz/jjiPt31cK5itM492yqy00pO5E781x0yI6V1K/hc4DgvzuVvLdDoBM0l/jwz5WmZPvAnqBjRt
rcQGtdNru7mn8pSrgHZImIafYIu9G/owpMwXTrUskdeC2ydAN+SNjq1sni8KfqETLqe8V5XaHYeh
vA5k18H2rlks3z3/GZeIGaCoF0pN/fdtzzGd3AF8iP52TXe2kF3VjZO3Cz/3vgslpRoLGo+HkT4S
a3EGYVAj8E+y/kb9BWxdYfYa/e0Pv4Jz/2SlfqM9Q2iaLyd7mGt0Zqn5oanIDf5ftuncVRx84Vsj
5ZxoxTQzAMeHRXRqAI75UFeNkJsu3LgUbqo34K9x7YqDXR6GszBQEHh72l9WcxAoC1DQfXTZrSWq
x9aQS0AVuJ57PjoNNP/S1iRl79kKRPnZlv3ycnYKcVqlhDIn8YHdYZja4IkZmKlE7T/tEGsej5oV
7lxh3FiSAFd0N8XwFm59/VKmrtK4LWDdMFHFP+jVlxJ6VSWQ1QZpz3C1FJUSCojfVL6mNRCco1+n
FGooqFgqPSTJ/bdZ3Mfe4k9bmTmLxna6gRHEtet0P/QPY4ehtmMoDxQ7g5YaZKv0CW9KsIzJmkUs
BPKWpTUGb/cYkEdf1Wy6xIgSf2nmoE5Z4ajwr6AS0LmGyPWxbtAQ0l/MFGzJO3/UBCQ42syRzgiU
96lXGMjdI/dVUJ+YrBZPUbuioSpYlV7ucaaBkIvhtialOvFU+plnFJgOUpJYjU9Hxnkkle/NusJK
wezm/HjPz5IkQN+OlEdgW9vnfceK2bZJxOIi857fHqXAbi++dS288cGFwH2myy3HA6r7jHqjkK/N
qTQrw+npmKpWULntDUEQytl56WUk/KlvoThbx8ivPdNjV3m5SuBqTNYPmQE/jRoUh5hxAAJ0YG86
RZhCUSrgcl7j5+9u8DRNoG1unUC2lGNdZklQNDdkosGt7FWS76uKqCeFCpnEZ1W3OtP2ashXjoki
HgKZxFZToyjasRKkGDMzTyRZSH09wMtXlhKKy4by/qveF3YEg06LsmV/pEBiid18z7llJJSp6Exf
S1jfWBSq2SE+LlFNEUJKWZ8jhOn6gD7HDbm481FbU4MINBtwc+r43R3UeORusFiuQMfx6v6WdNNN
9VEa3hsGynnDkM4jAMN1/+PpmN3bB/JsWhgMeemLaI6yxHm9nuZqcThWTYoDvfLnf0S6mWRWvoPS
YTTZkKpztTqGJpI3o0bZ7EtyCX2jvlEh3iwC6KLEf6LPwPWmwMMMZWI10tqzRv2DFatvmzyqGcyu
UnwR8m2COFAys/GhWn8I6EMsj0A0mMPDKp2593j2ue8FJLysYMgYarYgc6MqPtvqpfkqhiqK0+Px
nveHfrygxvznThgnn25P4Gs6Xm2/Y6pYueRw3g4WlO0s4jZWO/fZ1VGL5RTsoxqpmj6JDxZlGPAn
1coAGz2ixohvRQAdDHaN52DZNpSdtopipkFYNtsUc76bUpR1huBcLV60wxhuDm84KiTpeFQqSh/T
b1vYqkRVf2NJqwjqETVfDCHJPEd4tjEbxcGYBrAQJH8qhS/0gmBc5kqhoyDlmcLlSAscTQ+alrxb
vKhvbKoCt9GPH4heOQojSRIHUsW2K1k7VXNNec2J7A/m2ot7xHfdjo7hR9BcO8hgwXt8pqtX95Gt
Vp4DP97eqCMPdgk3nsVq2GoOL+gri9GvrarXCDJAmP44K/vYvBavEUJEA1Q+WVfB6GqIlgDP+0Qd
PMC1V7NERShv2Vjs52tpbHCLBQI7AyUsSg8SXhJCw2Yz4d+TG/EOqyVnXmljJdhAN34BjePaJzbm
4VvzzzR7MKPM9alPyjCiRAL7NqFkRsMLitsWOQfdGWqGRrW7QbQanHHw4Jrk4yYoUuhui7cw4Ifm
RINfZRo3gJS0//gjJ20nzxdxeOOqqNZEl0EKe0vAzaR17bpJF4XFk5CQxWYDE1+UTmwx+fJmgX6k
FFgrjM8n1SynOjRfYnClZiZjsO8hc+DC2QGtIRwe8XG9xzcPKov3aNhu8EX5qYLQfml2/HgzViwb
p2ZhdXiSMlinAdaT3sY4xhNHXVTvnxY+ae75wgnUyeUTHMFYkwGLar08Fxv0RH2tOXqrzfcJ49GT
uD+Mqe5lySDsQ1Pk9264T/SoM/SfhCTisogHhoRzxfGx4W09SyMET3q7mRdE72FvxHR/9Cbdp4Xc
fMH4rh64AxUdPQIygohOO4NW9GeFYRES7XzXuaG2nYhuv40SJ3pP3ROjVcYtSbNXhOoeqmRSAfsj
KNuRgkeQbwveCFeeIK4jAPTi4kfFG+z4yWJVoqc/48W2D23190W66UdSIjstqs5353jHYQwse02Z
1C08RfyPW7NAGfY4TuY7qiMhMQuviEuKntQtbQ087mXkqlwQKrtICz5gwyBJVtOivtqXuyYHceFc
YB2SzwMpZf61l2cfRdxKkqtwcftob2lUE7y1DhDLPdsOszXb0EtTFEX58lRW6A1s5leWIi25bV3o
U51qmqIyKzPg6WnUo+BfgSYpUeuHsgoo/1CQv17s3/imE0zv/u57IcA9JpfkDiNxRlzLDhzoz1s5
nBwsjCuBZ84TsWuPZczZGyYjIPo0SV5PDxYBOFusDKpjF5oBhKNu6BFL1O+GPDsbmx8JSssp1k56
tP8kbTDY8jNz1hZXsghqZJbEuA2TIoYUacM0DrhCbRdHhTOC7Pty387vN+3Rp4E8NFBqtfOwaQ3x
QQq5roWewg4MEKkQhCLG2AjyQgFebHawauvT2j7xWiiBoGIks7kVyNLpAg8+Zy6xByrrbB9t5jtw
k9NoL7cFqoVofuy+llOBDFRSCkUz03qPAlyS4IWAFU9LSgxxhJt2cQ0PBNIMu564cGR4a2PPK6hm
2ke0fA1A4C7poEU2DnaZiRIZCHeyg6bAYPKjOYGGOv1wGn5tXRX32hAkNic6F/GSSBJqGsbyNpdw
pcQwXPtldmi95FXrelybbpwaPjXmVUAQEK7aPFUz799ptUxuEBqEm4dhp/lwIeIWS+7w/Gx1oPqu
Z6EqupD60taBAIr/FJAe7Tr+GFEyL/EWoJIeKWbKEExXv/yWbcZzVN5LU4WSub/85sJl8uXKcm/h
e4DxpA6S5Yju/yWe+TKfxj4xVi8Yu5t/o177Xhx1jIpyZy1jIVKNvWxhvfHeb3AvLhJQTOg51QZy
wmzC9upiIfAx5HcYD0imFYkKleIRv6zPGbr2mTu/KvrsmcBWTqzQQOT4trMuj/QW+cbdWmSK41A0
l+XR6//hp7i3Lu8+9sQQ4B39JwIvrj3myXX1OQZapXzGThdW8mW1twnnV7JgO59gCkfnQBhDtdcg
f9zdCo60MI+yfpWpXluRsez6RQ4VzzoYhGabcNTbKe5W2VbQuBw44qNMU+4sPKwaEOgNOaMkhx8u
uYvpoKd46eaK+mxYN9slkFTNW0mm/X1IW+jVNPRAh1scdvdZ2j0704VNEggsaGbut1rxPUSU5fSy
K47Uj4bU2Sk3rmLG0uCE6+u/0WEgIB4Pc37o2EW9bUC3bG2f3tX7WKAPj2MrUstF9FJVaAfoEs/v
N+LzkzOx9VnAIv3rIsyQtvqDAqRPWuJz3zXSiZLNsNaI78AxSiMksdLEy7NlUJsf9NgjBD3ZpMOW
Jy6lfRbTempQ/dQC5guQfZXWgOTgGuLC3q7D8mrid9Vk+dT/crRXKUkBxdfeOuVpQMqHO6Y0Qaao
52s1LfgjeN6N22hA/FztiXGI5sTMWrc9QNdpuTlzGEjT0m/Lek/w+PEO7ol8UegS1UqPiopzkyT1
MazSHMVmKrHQILXfdOu8aNVl+l80Sd/mmYQa9aSfQffD1xI3XyhQtgYWEJ7KQvwl5GZi13gxOKrl
ngOTK7l0UuJmBGn7nioJF0KPUI0rIytXRfllomQN+/7esaM2IvXahKNMZHg715lnhJWZFapQ3xbE
eFqrbo+m+2yZLp+z085u7QEVXyNnqLRclXgF8VfvMFsKGy8vHwoh4i+wWEO7fQCQ20bsC4elTtuV
4Loy2divJ2VzTtaf4cBNt0txlIPhdRlgMCNAPGwqqzQsyN1vl8s9RtuBkb0fFIYAx0drjyPdfOut
grUy7Muee9ab4ccp0Tuwd6jjN5uEKkObCzsG/h2RRklgXMmjI4ubQtnsSFdeS7F/OePdreTf3/u9
LHvcOnrEDPUIK0BcDDhaKGlp+mmGtZLxXWm5jiH2ElVAFl+Vdrq7EBsDw2iZKkDlYe7JEHkse12G
cdv2W6lMGlmGhHgErJAT5ns9wyBSWGwXi4YZzgqL2zBBpAWywAsnQ1K0p4r7PW2yepJu4hsG4aMa
krhpR3EzfP6qjvnDiQDXPqQaq+FNkfEvJ937iJAHfMhpjJcWWoN41NAtgjepkJQ7rxG1njjBKZ7X
WyBQPDSn5Av3qzE63tVw0MuNYzszJTtrjhuPyUzhHhvTa+EBMkmPNf43Ee0ntGWN4USRDCB1A792
QC04EJ13CeUiyGPDepfF6BZt2MyKE9vfa9ETnGgD9akyxsdZymqZatER9lllHbp6TLReEQoSkkul
UkTGKVGF7Ti8WtgGjQuwvl/FEiMbH9vIQTBnCjX7SoJg0HSrpzIwyV9+euambYCLfnXV3tDkKaQ8
Uc1PNQnPaS2ztsKnvw5B1lNlBJy2JOwIOr2lqr2YHtKab6LnKT8TuJvLTe/IPbTNwZKkYBZIIIJS
47SEXRhXGJpjQ8LZZCiv4hFfVJpJewqMWbuQQREnej1XenGmkCrdaRsX+KnQobCvgBjsfgFZRd9m
B1mkJbE59UfX7WG9WkDOulRO/k4m2YwDU0emfjZiy0DkqV2/UPZ2TivWXJLQHbpe6e+ywZtVnic6
Eylg5qqDaVSYXH/iWlf1QChl3NZ21Qpkq/Z29+tBKXjwm7+MSK36TaWE7MMpvyhujCyfrGC6qyvx
voDeTJxc3Ezn2tQ2s8kV6+4012lH0xslVHDPlvxfld5fEk5j/MoGG1nMQM+iJ0qRW53WsfCV/7x5
3bdx9BsGkupQHJA1DP/1WXRvXUshVxHNWe0dPDq/RvojoJ17dHFU8fu9VjreaL4wUYOfOLzwyZ2X
7irpLzdr/FCsCu6eqRXmYEeEFY0cW1ihW3LMK3Jj6GcAZin+JXbzNnhlYLVJ+hNgVD9DHOKrWNIY
z1ndAczE/4Me+1zX652zvEy6chrGJ4+oQEbnk745U+HoO62ipRXr/vssnu8tOmO49bXlHI0F8kCE
h+wupyP9jbCr+9X9PYPrfP+r+DBC9Wh3DuEtPJ4wikc/p2rteRbS5pj1dTLDKiSXBy17chgObcph
zMlG+8Gt4GTsF2VYstQlrxqS36rzjtvWhGEehmI+sn5KXyoI6S9H8lDUHXo+cUwvkXTlxgYo3J9K
G9HgIjujB2LWf4YERmepdduAVsSx7QdCLB196+bMen3U7tmgK2XpOuEecqCKdfH1NingZ7S+f8RQ
nSMOKv4aR0amd3Fk1FPjt7V3FxM6ZY7DJdwUmcApkUrfNnG1ajDWkXGsAH/g5d8Vb7mDaMqTqKnd
gUCcUUJ6u0+EyjMBm7rxnte5lDPZpuS9/ScTZen1UmokkPL1ussjiPD3/dhOJ6mZcAbwlATZcXqX
6C8H85cDdzBUOAafo5ad/RhDFmlFSGxeymF6jvpC1N/qXj93b9mLKOFOUB86TCKk2n2ZhEwJscGn
Tuu1/MO0BuSHyUJG3Bh/k53vcjfppQo/Knh0gw2JbjKPaOC62SiwrDeA/P0yZZURROsgpyu3I/AM
ZF96XBYFw+LQnx60izwAqyx1qAo0xbV1OWnWolS6wf69HJEug7pMU5Rg7Af0W0okuUIUB3ZGeydN
L9M4Rt+ijFO50cLwEwvGtVKvqJN9RQmNnWyAvsWOvHMIcg8Tf6v6H+GGE5nlRNqOtoA4F+Dc3yEY
Abat8uskMfEey9cKkxXiFz0cBA5FO1kPOAVY2P4hp2Vf24+kezZg2BYD894sSxtqCjMa+awnL4oD
X+ovQ8ZuCQw/lMtZsLHvXZA1yHHdro+V92FDUNMUHgbFodZ0BPCeA9Ju+GxnNOpMOY95LgL7rubK
8FpzwK/smonNU3b23wtA2P/ZQmOKDuyc2lWGBTq8yzyKnpAGzHWQkEGapTNEIpz8g96mrc13URV2
CeLaAw4h1TgBlaTF3+Mi0v7e6tCPHHA4du1Fku3szBv4y44gPfmiHDz8t3FtfkYTimAd132sPBRp
ZYdUke2aDqc7OxGppENyPQaSvj/aBQGHwaFeQY4UiuIuoaUYSZ1moMPGs7i7iepfY5MtIY+CLEjS
/0h/O3RzIAN3BSQ7pSThudAumphZUjPvTU1qZ1ALTvDNtV4L3QiVbaemo2se3uSLOd87n1wJxAtz
Pay0yZrGnHbPjxa1fvn04z6o6iqkpJCUdFu9fm9mLeDZk3BYtYSZvizETqU5Cby+xfs5ziNLaXih
osb7E70f0XFBIKc3zHZmZNS/Xsxnls8eCjiXqebI8zbs/HaOKG+t/pYUKyvoaB9LxOdAWQIHFm8k
eVbqc7MAUNm3kVOlajA67TdvIXcPBHXtQ3IuwoqvumCO03tS64o5pXyk87aIhWJ81a9RRtnlM4ZE
ShLzmXY6STlhlPWCkm35BNRaQw6UEyneVvc290O0QeXnPZcoQb7SilJinS9/vApfXv5OXodNB4n1
31yIKXazODn9hSL7jVx89xwRoyiULN8UBbPEaIp6/pruR8ao9N/10iXMF/NjK7RUCkYzQFewXs14
aOlrujpz+PL2hkr+JVGIoP+7LZTpEv3SyR1s6NvlcVUltTSZ6jkHU/uRH4SDz3r1jWxA8o+1xfQB
ko2C1uaFIIizGzIWwoetj23RTsnS59FhJbsHZXoAGsz+opomgbhtwe5Rl9UdelTQqZdfQXMzu3N0
UpN3NXaLzla7jvo18zkYvzUs5nESsEZVIdcYFYg51GG45GKoD/wQFAnYj+E/o0y/7UTt1mHf+rie
Vjw0nTSxlUkRFFyNOvZQZ9u5kaRiaetwKhq4zDOZnUR6IzW2TwBTHGHjU5Fswem3CTRjBplmxM/x
zcNMlhmbCGTUv/fC1QUVuL16o7GY9W0TW4Q4//b7RyUYX/qkQ1dTwNP7W3JMnGzjTm21YzfZdzku
F9kN7PaIiblBHfrcoSL/33EdtdsSvwJma+YsFwHKAhF42Ng2mM1+Oa1EPFGwF9PN0yr1hjTrdn9b
A6mWpKJdn+di+8wWllDNmOc5nMFwT/qP7b+mwj+VEF9bsS7aIbok9KxfHikpSkrCVDXUkl3blplx
LTKyWuqeYRyjp3qQOD4liP09kVmN93uJ66FUaL4dpZ4h2JcLIzxa6EZOeKyDqpKXgIe4v1kU/kR3
bV3zdNxc7UalddYSZKxQmtLooSd7riCI10IP1dFpuyP/9Hq4FncVwAy6aCAd9uGFTevK7LcXVGB9
OcHrPPEPyjRvZ4sRZG/oMs2iFL8tdbmlHT6ixGGZLFEwYgQbIXPCJMUFEgpRO8inpwrhHTyagTnh
07MEsB/WFtkBxiII1NPVbkbfFK5M1mn6aNa1DaK7p39Tbgaxjj7Y/Gyxwd4d3yH9kXJhfPhTi+BR
65CKEEGxmOAsi+FHTAhFrVDIFlDK+hLvbwHuDq/pt/gapvrqyRsB0Cluif03tiKiK1sIsJu1mZtI
TBtYAwcFZMDRptmUWcL13WhcOe9CLXHMGVtg0yH0H5Z92Ab2pflNM/RlQZJAQs8qgfiRfF075SPR
0dYKf5sFOudf/1dgcnpvlRaD/vkcEZ0soxGrCPiW+njIJ4qDMxZkVaGRKqS//XStwQawmz4w7HjH
D1l+sZhIJ0cEoc8rpUxZhn4upW9MM1GgwOz6JTEAJscJnBTUUJ1Impq1Ab3YQEEug6fzxLrDtgPw
pvK2Q6nO1sXZ31SSFwcyUKztKqGeJUsNgM9MxCh0lrTaOpVxuHmk40O/Xr+JCj0ZrxP4IwJGsfUI
TlZr6PGH2yxMH6H9wm7SBEQa1VfrmtjfP6uSxB2lX6PyXwcZtTgkzCtmKDnACa0F8keC8ruLoQ0m
op2oLSOkp9ddJpOT+KYB1sHEb4fDq5VEZbz5yI/Rqz8Esq2qG6u1/zG1oFvPafK5U6jHhhDPQXAH
wAcsze6YZejnFTZWLcgAmFvpktBCBbbIMwiCbXdVZTuiCPyC3ZIGwWFHcdUJBqBdiD+xeBpP0bBQ
TNNnqMxEWdODP8LDNHjPO7NKba0jou4SNe/HSgqk/qiEsaaZzXkLcTqOxTELOUUgZJu91YYL/2qt
sBmvfLW2mvax/tVsT9mfB02bk/4Xm3n2FcXDbXIf8StiJ3pjX8B+rnFsWoWsgvT8YnoMkl5ss8qs
oAF+KBGWOw5fq21g01rnATqyB3DiwnS84xZWAaf9c7Bgu5tvdHdXOOqTDTUcuyfh7r0e1Khq9YXV
3hb2aSQmyIFaTiesvGgtGcGU5vKKvHWcK7GgkIynmrcOwxmIGig48BhVPaE9ZOM9kk49Tk7W9WSc
c+ii/4eSmhSiDCwOJeknsr5/9MDTXXBiE/r/6wXZy0qJUN/tw29rDnHnCYaVYHDojrj0rD+h5SLb
e859zudY+OFtnDgdgj95OCz97hi3uOxC8uSPvmwAzTBKZAhSdudL95nJgoFZwgvLCRuciPl7ABA0
KWrejVgajQ4hp7WbYR60ZV0EEAHKxfirZjPc5z8l+HfcF3WZ8YKcqa0WQ2IuZVppFnlqTbybRSvh
1UUKQcg3bGBj3j5N3V91/fec9tWwR8f3/HjlRbELMdEKLBxgGot8GUQEIthVsE35Qiy8F0GZlY1d
DWpMU/P1rrp/6dDXHnjkNFhUYdb6CCZ/DNmiKMsXKS0WG32XEqKieDxUw3ymopEh/sEB3LnPGGmR
pbThT5Ve7g13CuHMSmzZuXTROtbZr7M6MUJ93+1bsRMlPssTjDAV+U/Zdsb3O5tLpeWMaEfTMBMw
98dKdMlB7Ak92SnLoeVWcysqZj7ZPOz1j/ipb641LgkwzjRYW6JQBod9BnvU7dWpY6SIb3dEOYND
A/qB28CpyfraXWQN068BUIuEj1ll6ISn/6yJ3xDE5WPO+ffZl65WtZRdEdbsyEnwrWFGm5YOj9nP
a/JvbwUEc9zxjmfsCRBfKKLw/r6mqg2FtRn764IOnv4oFz+LWKViLiSagvRwCd7YlnASJRBose6P
WCrDy4Dna2jAcmWRblha+3CHJbBfBvsauhrGmCgBKbiv4RHtWkfdrwwabAXlJstfocj3twDIWsMW
9lhsTSUxG1k/ZKXlxL6jQJAuNz9zGZUWSOiioqvHZDjLJfnAy+eTvkxH+tkGokF2J1XU2a2TIZyp
OoG0pD24pJmRg26ch1R7VFTZJo0NHVc9qZghS0VWcz4NG+kmpkd0lUjohC1Snqogt+Gnwza5y3bs
V1NOAEqafISUv2yHFcH+xLkc/9zz55BigZ8PslF7eHSQ2yUev/MiiENzu7NdL7TbNbWJu0bniqk/
IyX30MoEkweTiNSD/m09ieTGRbvUe+4am/dRnEmosBZozEzwehaUymjcEiMeihmQ77WONgTF7w9+
xl/5pZHTQ58f1fYso9BrC8YHGDnpGhgoEJrGRX3p517xPdcfUHZZNi81SWKSqMa7tyR1LE6W4fBy
OeemTR8rnAmyCpnp/YuZ6z8aZ3qEqDOzGuHBZRqkljW80ENxIwJZT9GZFeuNX36lXJxXhpe6MZiP
lI26SgPRl92TlxDG6vp3yoQBOfpk3bObuzN+eJeC5jmeZOUKNguIhxhHXNJrimoYlAoz7IeKFarJ
HKX0PBTbzv1lscBO9uvo5XYB4zV2xpgjw3/p4d9Va6pGLqRM03Q1Yiknhdo1e+aHo5giQtdiyBEk
gXD5yIdUCkEzkoJWa2Ydm/LV2s2U0LEFc1g64cQdngj5tHG8dGzgg1b5tD7VRgMr6MGVIud9P6CX
PtEx6zMo/4SxqLXCoXgU2njk5KBNLBR8cY380oLBhdwDhY6QjSvwQ7+ooVR9H8ncFngAfBA4jH18
E1kVaaC0MGcxWsg2Y1DV5oqa9R3Y3b3pIc1c0ATM2ZZRLLxmyTQG2qwTHhQ2b8aUZaRdZ9oF9K96
XjJKfnBuIDqm2t5G2az6Q1T7RGcr0pTBJsCgIeC+cdjv2Bu34l6YZjp255tVYo8odNEu0hrFJYL6
rkzvesiYFdrL4sdzoOpklj5ShizClEzZuh6uKhKsqOyCVxsW13m5k6evlZFp45hlRCqsaTRfD7I7
RuL/JAcCfrzbweSmjeqcwudUUH96JPQPfiwPCfNYB8usaK2tvrDbQhlEYPcywZvfxPDdxKguBhDW
mQqOvIzKgugNAp8JgCbUvv4dyD+JfBIWBsNbwHNNCcRUwyk5Eh8/qEW7MQmhBiiCZ/vMEUSCub5z
0wcZxl5gs1fBn6fQRTAq6onh8Gs8YJJL6OT5GwqT/8Ax5n5jyMmj/G94lNs8u/EtKqufLij2B4A3
BjTc77uDRLXwgpRtBedfl6xlnLskDHrfuecjgoxrURKGVtHxSfT6GuR59A1qqILvkVngjs/rV9gA
D1GIl8FwLF3Q9L9YoUWi13i9MK7u5KL3DkstS67Qj6rA21jhPAQwEntOKFWjwezqKpIfwq+/v9N1
N4qKRRmjSBNaKb6j3SNsPbjBvq6uTHvzsA0WZp5W7CsdwYAbwaWYOEBqBGzf8ucbTe/P4X0Dp6g4
nSLEauj2J4gXAZD4jAL4815v7nV3+cOOqge4+EjgLvU6M0CGVe9dOm0LUVwWxpn1FXTTZufIwLdZ
O+yKaiEppa6Mb1vNXnRr1NUjIQsHsD7ePNlWQRmdf++07E+MCfBZBWNTSKt+0t+NUNN6tEagmSdU
xIHPZKyhINp+WgcJr1hHuLKv+KELIi5NsT52HKBSIrLP6NIDgyxvmprsHiFVvEke/3VHqjxBzWwO
G78saw3vwYdzJ/Cdxix8UM7lOR+9V83ey0c5MY5wfYeQ9S9YOgMwNM21mPWj6VUd0IBM1WIAo5Qk
WkrCYGr5BSjUcAb6vLB2lScSZRwvqLil/MHiCtw8x7bk0Shx+oAVIUxm5HkUbsYrHcB5a/FzUkVb
GRda4tLpzdOLP6rbASxr/OJx5vhSKkR6+tW1GDglBO72S8aT/ftXD59zjZ4qfLKxs6rSufKRtkGh
i8f6FaDp+DJIW9wTbuU0Mgppw2U1gcx3/yuE+X0cg4eF/6ctePa4vbL1/nOl1jAIlIFSPZraY1ko
mZDckQKfjkAN0JdKYNMv2ChNE0+C8uVSF53/gRlGxq18/VkRzmwZlB8ZkMGg6rrXq4VNWV5wejsI
9vzifXyxqQEBs98K4bRuXwD+ubkunsItOxtonLpD15bZ6CevhVOBD0yIxvmor8ENVZ/uQwq/Tbjf
2IiplNJ+e97BfsWnxAQz1UILiTPGHmPEr6wzT0ftSG0PLwtt28s0AzYe7ku6ew7VKV1aUH/3qBRL
xodbakCHckgTRN3RzsT+lEBnLiQ1uEgXA/Vb+hRh3kD9dp9Kk00XrxYPEZ+Dt9KuTK9FiQoYXPFa
tKUZ25bFHlyxCZKKIQHNCAWYiPrqOVAe2xYAbMh+ohhMZeSA9AbDpVBORvFasETUzUeQLiMTzBVT
xPR2VSBU2JOdfv97cxcxsExOb2QioL/iBai/Amo9jTEgqpjyXp6UCG4w5O9FrucQlwmh6IBDBZrE
F9dPfrgWK79CWAAtQcuyEKmu9sFlIxtQyGzmcDt3P9i82OaPqw3LKgMnOqHUIbSi1+BocRFxJfXw
rMNoRCAf3ypzyDuZ0HLpImkIdbX4vwZ2qUpyBKAXWLQ/JsQG1zQwA9+yommOEcPoHe0c40mTT3+K
tPZU3vONvmlbfCGoq4XqqVvEtil5W4LM7HoFM9vRFxwx/wtUQHSMxlh3QYBANeBFqb/Cf9SHxzSi
jI5qSY7tzBWIr7cE0ZSki1wzbfsh375Zft9Th+l2eKtutcunyTXdBUg1md0dPkPWJf+ZdNxFtbYb
DKKgKjTMJCG5jqmsmouVOdVxWt36CgkFij+KRyS/v5ea6kHeUev9LVbKlFnIBHog2zUIIFoGn11t
3EUWxfVn6x4uVXSXwVDSzEZ4ix7svq/VH+NEaY7A+KAz28cgFlyDF8Z+ROVeRddf6xsF2GvIjkyK
G0EMfkIhnXF/VpqPEIrGSMYuGkv3tDHD1dGzUFqxAPA6C+YCrwHhfZfA85biLfVu9rjOOqWzdxMO
GNxu64kovlHmau39cWdcUPzePs+Y8acPkHtbpDhkYwj6AbgqfLHgXYZZAaRCK9vCnKCqonslMOgi
V61MPUsH7bHrn9WfBjCTFUvHKf8wYiUPq+bTy4e1CXGO/LctBkjKM9UR+RCWEz1bXvK1YLFEG+Gl
CCG1iuGhPsKXqJOIOI9rF5Wz40cjzx0fM7woep8W0hIs2/aR3M48vSBPQzpR4gMG5PSESkJj+VI5
hnyl2C8G3rontrGu5PUSeSHq8FIHpdTFSKGNtZtU1anJFDKkGzaqpUZ5Htd4kdWwAM4uKMRhMxtu
+Xxxun5+oP0yYfU3LJcp/CLr3rr4p8MAm3KlPWydY4PdEpQvgFJWaO1hDE0GfgOR/pEJEXTOEL5A
7XV1RqGzY6uPZndIXKw7n0qRuMWV8RNlnna6BfFwMKXHT52KWqb2/pqiSRnU3a6DuCq5VLlPxzfk
Cf1K87M7mSwShaOSkvgKD4VQpluBVrME5jrxW6v3m5lUwvMXeAt3f8g+3RjBzI5q2bJD+i1m0jiq
zSfZPmF7mhHgfU6NG5ltfX67XLFZby28ACFKaarwpIVJgYJ1B9jh15eo+G5cHRTec3AKoSlR6Zhl
5pGOQAbzyKkOUQMN60GX2H/w1aqB7BkPcqkZ/4KSf2fBWZwA0F3l1lHeVEpfHcURU5SQAAGE9ZnY
fVMTAFcdFnB28DGsBGGQBDQh3VvZxR5j/lUMnKuBPZuIUj5YL0H0OuhjqkiUL6l7FjElIb4DCVsb
M0XZIxNeBX84LMK6dcgk4OKIeF1NiYqgZl6llcF1teHTvDTC9eruNpIbAYhovtpsIbrSQBm2LEqf
1DhkPafyo0EefjCoTYi2bDfRWdEBDKdJusfDm4N7qSFRsli9og9+3OJdSS4gMJtTmhaa7+K99pix
rBI/1V2+rJBHmkYzCNH1ew5DNMKxKEVE34Nm63rrRPw18HJpSa/uMaJLDcxUGH8ldy61WCDBpmbQ
hU9vGq92UVb7EhffYdhc9b9iJquhFJqcfg6HvyJbLa2HGKTEa5oa91/8mm4dIMYW7zRaqcslUbMl
/MwRVz4YhG4L3p+X5ZN65Jj8GKy0u6IM5fEiYfbtPn2CreB6gYU65AvxU45RFnog9/txJl0UeYYz
7+PN+uzX1k0wtb1e8MRsHG9eBPCSUCEE5Be65qJHkUHxzdOYst21kQOWwR53r7uKekikdHjQxi42
0XD/PK4DXaKr/IiNw8huJe54BNR0GdgmIjVzaERt/zxKjJ8kOlrt5/v5luahGkWyEnMxkAetZH/N
ymncW2RfYi2giVXkO5O8t6Evc6YCavKGrarFt0RgYSQ0sQWGRAN5Zr0LSLN8LR1v4tPxsrks1AgV
xvKIRW5EiUiGLsqyUlOCePTrTIigKx0/84fmgjSPH5t9Aox6dmUPI52AUi3HtSSot8VrwQAf916a
WSNvmt66pkqYaWTbsIb89+BOg0hcidzc+0zKjg+dLVeiS255ar5TPMCvOvN0BDwYhxcbo0sAC2pZ
k8xgHf71HEeUtSMCelHTSAlsBuM+jwGgZgD1h2XW+8znoEV2oM8tA5B0g39wMrh7618zFM/YTjHm
cxNz8zPJef7bqH9Ai/115S25ulN48I/egx1NoKG05T49RrMDZYFQacQQRq0Rdep4qtW9l9tlswmB
oV3894q3pFOZ+dHz7i7odjQVkoQ3qOCCu1fdjwismy+u66pqERWeVv/Um8rMmCjrFSVrrp+2vl73
X9D2NgfxHIDG9cr0SvR3umoEk4VesyC/oSc9mgvL1SADDY2hYkEKO3Sd0cKmnCYlDJvNMYPPdcrF
MRPtQo6d+ylJX6t6dIaJwhiVNgHlOzMdGOxM306MWUfYpY6nFgyA8FFt4xRohsEUhr+jsBy5SAUq
8twnRdlkvCEK3Chjd8kHShhbY5gPXXL2VyqtejE3KczYhx6hMlNYk1xBhCWOBh+sYvnLBO6zlqjK
HAvjNbGJXGUzTtaFMV7itlqtx6LObs7rCQ0W7cmZhonN8YhWFJsKWn7IO0SOvWYrEwfTXzfICilp
G+OpOuvqYdAurE63vEKDkrhILpjqAafYsMvGKlGJvv4G9vMgChG680yohECiCTpPMfJWaTpHUWJG
nDciZ8YD3OX3XXnOafd5se8AjQdAJvTw2aExfxQeKJSNcqpCZtqckoL5klh9ljoPQ8ofHNp2kSjj
IBA6sOWc73TT62ZoGGPKDjckOmaYAWBTm/USAuVLlXxSWwJK68dEFbwr9+KaKIngQq3CckULcnif
ex8AhFDi/AtN8j2gg+UAhnb22WIHE8K11o2DY7GUrsGLI04Yr45s7WTd920fCdYwjyNGZG0sRS0w
NWSZSNQOuY+d1RbjxK/GVF1NVZE+pek/lEJcxFaE8L6/TMWERDZ+ueKDluY5CqEQX4Z8I8iCox1L
0yRynP4+dyT0gGVGgCaX1nRB7jQLtlT4TI2vF2rB2eqiO9xP+D2QOPYwy0obBnyfdc/RTKAUg66A
T/lIaTG+oEB8knb+nZkWl+NfmpgKCfY0lGzBTiOGTQfNucSk8bf5ngfF/zRJov8XnwjeU0cDy25+
fSrPVj++ZmTJ9pWh4jyQPf/heRtmYbXHGEF/dLREwriutmjwXwQe7UdvLYki0aCdd/gvmPm02xUY
Nvuikj2o3v8zetdvTKb4zivNR0slJ1IFNK5dJFEQtvArFBQp/oEh1HOuYjl5KvgRrFzMMVQinYVu
sle3P5BS2ilcS1oSP0WM5gqf4ku9udG3lDkjUQtSrC731IBO+E2OIlmF5+YhbT4iyOXEOsI0DdmD
J3f9mAVd6jJe69GvM7EbnWUR0T7i58CV/MEyKMgSE2TjXRIyDpSEytLWIYujqX37JfUGyIsPlAh2
Mfv5UIKrwTm5sLjfyMBnI5rxZ44vtQvEX2X/B1vnG1C0j/YiGjpkOZp1fyRFXKEuw3qRMYu53prO
/ThuiZBIepcKQMdZYPpTZTHCMLxde+iusEhNyWMXZbz/4f3zdPINLJXADirgjwqXNrISVF8lhk/K
EbLfYDnFs4vgItfGbiK5lePDvnfbPCDuI7Ufux3rGknECtILslyq9/EJLl/ewNOCRNggbc/sAqig
hhdrZHqX1KegZnFDyJnvzItxjdWCI3lzClrBVB3wQwnJVxzngOHmlkh5Hlj/qgjf01TIKUoriebt
cNJQ+uKAtkEtJDsDROKRWIGATBtuWzwYcst/FaPXlK5idfaUW/ICTdTx3dLbWzKpNF7rlLJSPhPg
RLaDrokgXjDyGt+bAp2Ok/gXNHSzNgNV9SpqgedC+AdNYLZ0aNU36F62Gg8gCD7LwjV8GxMKIQRc
eflkF5DI4htp4SDiUcixVjVHW5SgMNOrPURKYWY+pVBn1wtVOebroZEYyCH9NCoNZHW9pMSigf+D
M0/tdNPjyMxBXooFx4o3q71eTS4vXxZxFEz5nmPIIcSj+k+KlaNNbabRQXxxK/i/XS/JPuSHum83
4W9U9FhfT4gxOkILIOqAsbJ9cenb0NNWmli0IHL10EFqNnsHph1Hi+1r8RuMaAs7uOMOdyv4iWy8
wGfYn09U5Eecyrc9EZkxzEPZ9ocwJ7lrCh7e2lZtCP6rfvyxSjpIf9/S+9hllpYGAkKdoUlADJVb
nZ4KZcFwtIqnRU6Iy0TqV/M1Qr7P35G9khwmwHTlwe4sq7xip/n8aVcLjIJ3RLl/x/DAQhII51/Y
wTNCYY9bNbqRbZlUbvBN8YSXzGks1qv9Porg6xrD0L8uhY9XoSZgA+5HJtq/8ZYGzPPW1HNsW1n/
QQ9MnNNKiCR0Bb6eC0LgCbQE65xbhINpAKLhRCk0tkVD139Gzn6EGwcdfe0nSw0Yfr+jalPKd+p0
OaFUW0rRhjPDP2yrNcXMc8nVTnkJ5okjgHFLs7XaQ5x8emqD7OwZKipLFsZwVcf83KtH23nLXJSe
8LnGTrYu3qk2CgfQc/Vz3dz5dawN74bNfpITwLBO+sgqh/t2FuqpunLkoje7c+v17KLDlzESxqfZ
nU2sKDEPSUkqJzPzhEdUaanPbvxfJkp5yg2T7luX909pb6ruO/hTI2NeoNgvQMz2oaE2W6aCFyef
xFbV89bRECvAqItbXJ465e5vJLeF4/9b+vduYvkx6euYSiumhlgtbPNtkJZjeOZwUNiEjiSMALVv
aZ4mPVkh+SfayLiibPIAVapfHfTjr3mnLjG+JR/KSV4PI/OLreLwFt457ViprVQgfB62ybWxNVdw
w5gpkBR3V6v8tVshldpgB8ljgNF492mm+zVEAeRwThFc5kqEQV14Z/QDjC+Uu8AT4ru1CVFipWS5
1LTzFT4Rta+rzNYsS+iAbdo63uBsaGC2Ag/y+nDSO2JN63h+AefITpk3vW9ZtZRouOD4m7M4tBeK
bn5ABhzihSR/CUSuVKkk50Y1U+grVKJALaNKg3U0ekuODEulvnDXcAUhDoCCGc77TjFW0ZNviChp
ik8tZ6Cfr/FxrqIJAff5RTNBDBv3Nvt/pII4u3gNRIF5lBqEPiSYrUxabYxZOJLueypx7GTWEjEs
mmC4VHS81vgEiybjnFKYTJg1bOBhfNhZET2mGasxJT/ZtIl8QIs8wkV8XROJKv6eo5HnfShmB3QX
AfSwwxjIVOKxJ/2M0qZs5qMzvQMb52465R37/9xvGMRn/GEXQ0sOxMT0O3eRFAAwCIQVBF8gBItx
DNyN8RPxNeZIm3GsGjOX7/e83hywf1ip4HFIGlI+Ivo3/h1AzeKUbLe0TcY4RhBlD6es82uVcq66
o0fm4Ya1MJ6JS2QEr+7rXni4fFkjCMTQRQvRvend+1tRL6+4vULuVhRV0n/lp4vJ+kL3vUemXtps
nBI5NiJ2j9ZMNwP3XR4wqXyukdApWGDq87bbe/RK0YXf46gp9Jsu83TAh7yHIVdiuqRy9ZJkbg0f
0KYHGcKerAiQI2Tg+tHCsYutzonzRiUQfLuZWqIgtzi/JrLBkZYi8NRpueTLBf23vdmwRAAJbf+F
JM3km9Gp6CcyUurP3CyY3pjHYzNocl1zIF5UHojIj2Er5ZK3NIgwGIUAYATRArJG8M/1Qh+iy/v+
nwse2QUVpQOqznYBY1ejkszTxSTPmbiBh+g0yjNvYc6lipYp9KqB+9LKY1lTYex3md0SEcKpzMXL
gYE1992JooNtbOwbHzekFa/QrJ9zwQeY1mjsiswZMa7mtuKeFMzDwn+cl3yZzLkNhLZ8eDjTM237
o+zDo7q6gNttjM5Ocw50fsMGLCZ0Ykv3ahB2w2ZuSrY7FSrMWwgTDBDN4/drqop1YOECig3JU9j3
JwCXbqgDHxHZkHGPU2kLQAI+L7QlQfWbqRvnsUuc67bBi7k26jXJKVRC7vLSPboEIhs1kpzZRTXd
BlVCcrRNvCPPwwNgJD8y33ZHtHInmGy+k9ZbzhXZfUdqrM9HU/CzvNNGHPHAMgqjkndMV4ZaipDX
49Dp/62CkNNhUcp4PlWLVCMkiX20HNjdbDYnwNkadWOR6dT6DGluuZFya6ZyqTGZxe2Kj9P+Zz9o
aI/IKAT6JFZtYWUw7FNFuQ90HdA+ceGb7RcCRapPRoHKZX3bJiEh7bWQBqQ3qMdIB4p0EzVWjkxT
qdxxiFibNINRMV2M4ti4Vbj2lAQiar3PaeduYYRBfDpWxMxRbw/RwdZikDQ1D9pvvfrgTd0drucJ
8lZyEwg/NTjquYXWF5JMfYmTPfgM06r3qbK9wELuDZQPmJNLBR+tuSssuNgrsXX0+5FO3WEoeoxD
aJWUA/IwTxKnUQVcGRSClaS/KM8Le8jm52XUCsy7uGkaSPVVxb1ntKfNx6s81kx6y/jS++IV7iY6
7djzOa6536eSE+N6QX70TVzZw/bYZmiJEQ0LhWoPDRcYjqy5iHwG1Zo9MDuGAGnrdtVJ8/WpjDqx
gZBaOUc5Y9KEIqdVErzc2YrfYnfx83b9ywL/TUMYPh3TO8OnM72+RZ4K1L11KlTanKukA7RzClwU
TzRpnRmzouj79HQBaHJTjuM2GdDPiz0zVEtpfBJOXOieN0CcMVg2ETmOiXOEyYE02j6ekwoHs4qz
W6YpQtRpARyopFkonDNXlfgzWBgQexmpPXQXbuCmtqq9N5Ewj+w1rcWkudLNwQTA5Eao0yH3mJZU
TcucfzuUwBBhFJVLzik9Ln1aRJox1rnT8PUrdGKYx6/zmJVpQyxNxV+35ceBRTUeS52hbONsfBni
llNPBr2ZhmTWqXuTb4b7FnILPSyq8dR0ZWdTAmVzqysIbhkvJhUpIaY3vVroKgbO0yQ6c1oZhfNx
RK8fkSfdABx7B8/BywLCAUk9KfaPA6DRPyWLiuwOC1WYn1nDkIeRVCB7R+bBP4V4UldVjCdKhadn
BTUnbUIzu6iuYap7b1Jwc0fCqmglsqrlln7jIQtGWKqSN1k3cdQR2uOiQqj0YZRYl2egSRGjG+FE
+qnHt+8IponV/Vm51O6n3p5zWgOMsl0GwmCydXKIQlF3QFRS4oQN08hkoYk4UVkZ7M925dqrSEBv
blPRHAdM0RTOdKMXTq0qBsde8T/YumY8LVJsau6Oc55RQo+xaOJVYiwhZ2HkJT5NUYlpZnq5rA77
N+Gu10NZxpN6pA9PSsCc+Lv3YIJNFOGY2Cahb0jWcZ95lZttyy97fD4kM27X5Y/wASlKbN3PDbVT
V0FbIhAsK2xg3+2BVfShohxwKJpqOwOTASkICmxkBazyR8ocXrOgaqzQaox+19enafuYPAo0kkkG
tE8MXK5f4uDqTQix+1ikLljoGUKdghI/3TkvOLREa1WUTkV5c7UE8dOYDC/HkSmpNQnGSrFxIbWs
IVP92iPkTmAIwQjj2tiDoCXkCLrLpaGajtOmeW3ygyCnzRltpR0x8RqGB7QILtE58EdfStxIcY5K
Pvy/q+mum5+oUpP2D8Wq70pqnKFPRsIlxNgtBWJMaYe0gdhdLeLrysM1+6WVaDbEIeak3QbKeVOq
2WyN0JHp7KJDetw8KhGsnA1pMPyCjMcTiNR+BrMEy0XCdX8fiYz2rk2htH83BDZ7YPXZCzt3vlbv
95SwXOwVLx6j8ZmkD+KPYiNQLuzLESKr7qu7t9RXwphYIT10LTBOAYDJPRTsOGWTowniifTA7VJB
A0sfc0CdDAJiCWQKevv25HB4upFAumEU0gXrtIbPGv4mEvbiToLWVBMQj+wJvG0lvyo6YOH0eUA/
WzlOfGa8mkofVR7ljxY4yte9rH8hnt9uoAdaaXWbTgr9sCdE6wceap434nB3zGZmagQL1RUF1XZz
5djnnxqpMCGqmxts4p1kHpK6bz4aZuoHFo+SVFbEU788QEZ4/lHz+IEnBeCZ0Uz5AiG+hDOH9uJ7
8F0jhkfQIcYCkjCFqbGeLT+AF/grp13Iz9Hs94gNe1AaHsJao4g1BUlEVjXgKr6W1Y8e4OTCW+c/
sIuYKvGZekLzofVEGeEUJuDjpYO91tYu2z/nZN688eVULmm7H3KMohMX4je3ELkwb9tM7iy5smdn
TDRk6yoS+m1HkHXOlAVSmZv++nXMn50tiSE6uI6hM/Y6FQsILKFMAtuTBImZ8SA3j1G211/ZrTmf
JCdR3f3Xqr/LRoQO1ZS5qy4rxGjKVkDir4aCH9fPTn16HRWWHFKwgZWvET1rh/WD6FzKUNc7lA4P
POONDPgvXaBHRjuAXve8ZYMIuS5KYT768xIvKHy9K8zlqpaOp/Vog/9jKEkvZbqz3mKvLTm63j9V
/7j6+nrWKCzqviwMdB9X5ow8aA9KawYN+rgHO/7DDN4Bpfpzy0PgJG/GBAYAKBOyMRgH+qgUjI7E
INFIGfdTfeQRQovDO//2ZKLeXOlyg52JSdYCcm+dV2Pj20EltBfVxm/Bt3L+QEZ2iUMgQBBQEI2m
C1tnWhq/0clSKkk0Dqg20zhmuqxctvICxQ2DRfi6VK1gQbjP/ki2L7T8d6dtQEFGNm4/OZ1xV3jZ
1QzBnckqM/agdf3fSZu+s7XfGx3QWJ8vEekHxcUhvOMCB5UScIKDOP9tycX7Nb5dJimwfecCcaS+
fnOlDdNx4048DX5wTVkfnOe0ySPHwKnOU7TH6rLNhT3QA1hRAhSOtfPYzIyzNUsFOJpYe5SP76EV
aL4oDKSQJZcZ0WBa7IW+yiJPFY28jM9BKKfJ3uUU07PVI95gY4ydOrGnNKxDWzLHRV4bGio5XPn8
+7FtRDHWowvo33uTb/jusCMmwLLXJG72d8uWAZCuiv2hMlw6akgZAMtMDFf5b8QMQIpJ0ATdx7h6
lkjmfbNTv4pKQzBSio63bTcOhtrGP4/G55pqk16EY+M04QOq7Aq5OXLbmtpNPHWftII1Kr7CLZdq
Y4VYddvTCb5L/nY0D6h2wJWwdjoE0GN47XzkbMi/u70DCUhsxkLKGEaVaofBAM6DXtj6PUPUtoTI
xkBDqg7YyQQbleIrepxM2bcy85O8JWfE6ZoIE5hhz95nW+itcEEyH7gSUtsPULh1jDpbZ+Y/gSho
4sgebNaQ8z1Lbtx6WP8mixnzV3+wYfoa+Yw/z6ux9xZg3dEExjh+0P7Ew152/e6+809fY+O7BNg2
NKpl50rQT0kOj5tOfa0RUugqtJ1ebemcFclJRtxTMA9TxbBBN66aI4k+AloI49qAcp761Th1CtJw
Q1eZwFsYU0WWctWXYXC6I5lcckXi1h7t2QpianN87dZXHBa6SYJmA9RT0cbdoNRe9vgwc+yqTxyz
528DR68FsOPWwf04qOJq/yqKmE9pwu+d9JrAfh3A++IwgOzfqt68xx0PH8CLo2D5htMwcpBc+3eV
qUe8mO1qpmOyHwdARgU+E/AdWskdiHw5nimHJvjP04QiaFHdM8N3CHaMIi4XM3L+uDvupLM8bpCN
t8s7c4IFF7O4+dvsFJ/PPip12vGui09Zs/ZiYLlRR1G08hdF3hkC5dZWw1loRl222CZDqZYcpXG4
XGDWRYc46TLa86rDohRHv54ZDZEhvMSW3SQGodElxANWOgOprA5eA1IcxfaOxgex0P+Zz7YgSmc+
Kk0fi//ni2y8lWN24PYwgdO3GKEQO3ZevEfJIEwFTJ8PEwEwedrmWY9Cr2aQGxjLRa3DZ3PesfKr
R+Aaxqtk6hJH4RcR7Ui/8cHuNxI1Pd+yweW26CMAIyOF/Fxrz2+rwNSKSOC/0pUYID4waS7NDK8Y
JKP99XwobtLgINodq6DUTlv5VPtK0lFi4sL3gCVy5PvUT/azyeoYw0505MejebILbarFV8xohd5u
1yEiBIllOLRoyCdjxXeay46/Pun4CdC1HT9b9lSlvCU0OtEgL84rAM1CZMSHoC69IQmDEFs/au8O
qXA8FrZg5PlfyeISuZ+2OIevddxL8wwl8fEWEBTWQeSQUMBw2CPUZ1vGDyvKvAvej2PypVh8Yew2
KlFaltVjNF6ZI8qWwGl5nDsD276flKUeeGW6cehi6iD+W4+RqAL5QLASLTpMOJjTTzfDC+ndAdJ2
UXxfrcS5ANNobCetI/3DCVnDO7yrxuXggoQ9s4UILtO4i8qXOEf585rgt0TUQq+4ZPuM61XezjVA
TJ5Y5vyvwm0MhZfdy7nT7MVFTuJmcFHIb6oJimCOrEiM1/Lp5XYhuHPRd10oyG9iiyAEnYHapjFH
vGOfM/5XjCZ6USeQD0toauKQ2mp+zxx+RTt/7vsPsq68QeEiiDVMOiPGAxeiVNLjHfMihtX1aFev
N2x/LVToq41BT6s/EhsO4gHytatvD0EOO2UN4IDScmGYrHz0rpi9ceKaJzSTciFN8VCZX1SnrSGL
vEhSiz66VucGSHwfzcjdC3jhtjGhtGNQ2MZts9HEE/ppKhdvD2L2l2epIWvuXmfIYvdfZ+jZrUxa
5xUuMCUTjA8Vx69Te3EdEVog/hRYmrmoq5QSE8eOyhgEa/g3utYuEOicNKC4q3ryyhbEB6Nydsxe
2uat9bADofvBilLoBE9AGK2jRMwJVF+SfyS/PjuCk/NHUe4q/CcrV1Wj1aEvGbce5lOXrjm08LLA
tYRYH9JokNbcszBgaHtf3JDC+QEIpL3AG7ODuwuuxLdd9oVWMIOznNtk1Mmgjww5lodUk8+XE71A
Xsc7mWhcN+EEa+UFxsTst9epQ0h/rDIDg2uZhKMBzS1GKwNDQML7Iivd+DOUmMfSm+Rmsumnr0XA
eI89XV7hZD1/6qdv/lFgYw5zkGfQkpVabhknl9DZ7GdKI6huogFaDQ/wjgXOf3Xjc2eym+EJGvVX
bGF0jhc48x6AgnGKVUCEmSSGvwblTkHzwivB1PK4h5byxgXWk/x9VYywfQwK8M0te+LHCjYhFwLD
IW8yDIAXTicJuEb1i2+TiL464766e2nxjpLiXKXuwb6cyDtPjT3cVilS2Aa2ZbfDPhqaJSaWSxbL
cJqBnwsu80kkdLcLm/R8vEi0HBRbXftjJWXGyWdNkmbmFV9KVYYtFFtGPxQrNSpCJavnYddveq6M
Duy3TXqN+pk2M20Xv9eZIt5Ov8iLvQEvX6etb2igC7C6cI9aRnl39Px3gSsTB4DGTtvDKd2wryhr
Nsprw0/OrlXdCO4kM/Nbw4Zomf020lx8BLK36ax0k+F8VJejrvCt8rzGE/GH8YrjDaJUM2r00O+R
sw3tb4TtPJivUwcupGZvIcxVCWPLtTwtcnP07xq9Zhf+bs4pgMp+yH8OuoIseHH8vb8m9Km/+1r4
qlYCwktkwDDtLskI0E7otwuby005mIJp0VV6DhRtTj4soTQTLmYuA/+D8T17679+r1QwsQg54Qhs
46XzPV59txp/ppd0MjROh5zsiIq5ee+NFn853F/j1qaowbgipqxw/wRxp0V7uS3XBRcfaETKn0Xq
mMmUvvbLsnL8AEzGyD3ezTTlorJ2Ho5EgoKszYmUmS0jK/K+BaR0ApgAPpw2VN4i4fhDRFC6h++n
bSZR2Bkn5VXgClKwpjQQ9sxULCGg/rHkJrzd39Jr3OyiURb8VmQUgrXmCFDWiF2RwoszZElhRSLX
ASYTFQnYw5vK81eGFeVGjLX8gFYwwJ6pzBBi+i4ZRr/OxoXoWPFCigK0S6i6iGuRoHIVVmzbm8HK
xDz54gjVhbS8bSWGbh5f6C7lpeOyQKKFL/YJ3pX4YDc3uejAtirmsK2KQlnXSA/Ql2St4C4TNsB5
Tplzj1SRpzuAO2UXQnsnVAm51ewmgLeUkIlNBz9wW0i6+Ex+Y5ojn6JC5mrqowGdnFpCB3S9+3i2
qwKJrqOVeXSPkSUOvuFNiP3WdChFlUTpPrd6+SPB2MjnWusk/mGc0Exk+PfoJDrfjv6Zbzw7R8Dj
Z2rXusBeUgA9++Z4HuijcHDD4KjDlGdhLrC5WGTsuNHc9CtpfclH68QiZXCW1oCxnxrAgRQ9vHcp
2bj64JiGojYO+SdWchW7F3pxyl5pHrl+jhMv33MGCBtj3q2kdV/sY0NNxQJPT8QdSphmgXmUcK3j
n9EXMw66jUfI3sJFUWE1TKExVGMhZIccFi4vP5ACBjqeZcF47AbRwJlI08/Q3WpIOb9qlNKpdQmd
hlUWD6a8D2cVatUnmBun+33nRJrugJjIsuNbaYpg+EHR7EIAN2pflzDEN9VvP+ts4evSkUBox+8y
imlQZVC4aA8DBsyFifY2D4y1ZNqKQ+m9s8z7SmxipM2kp3WoKx1UrK+Po3bG3R+/eSL+ydN0F0ZQ
4jDoS0tNdS36fp5NXwHSotomYFftFYc9QQmJLObcoAlz+ugjyz5fNYkOKV3QNwj1/KIFoMP1CWVn
TWB+/bigo2NxIFFnJ3m5d+e3PuLSHDgIPt5gZkg3wNZ2Y/YFRJReShLB4dNumZ9hDQtGq8YJ6fy/
7SmVhWWfU+Yo7DlLqTdckhCMpegjiLlBmt4y2StDPks3JtM6s9pSUBE0oPEV7sBHXDgBCO3vJNPh
1yE7gUovZ/oA5JX0//VIgb0yphEtMZDfyQa9LCeayzFX063EQB8c3k78pHP2ohzflg/QhSV13rk8
pwM3IV+zPaXJmnJCxq4I0C1otQHs4GsDsfrxUopp7Qvj7b/XQWvIGbP01Y2pEoeyFkgrx8mSTnqh
BBEQDGQuzJVsHY+XMry50THtmwqHBuW7YmbnJByM+xbZCcUx8TTgObYOXu9L75M0OV4U+hoREC6u
BaZu/5SZ/XQqnS1Exd3qDhinCpLxU5+q3mWUGmh7Q9spa8+s6MeYus+SnU5P85flQqwtn5DoE6k6
ThBCDp0v8bmXkzR3yrJEboJhhAGBaaMpk7UNgig+7LOvV4qv3wiGolWHKfB4Y7o9BH+eb74QQajP
ZLWZJc8HAuBvi8gMmXQv6Ze5ZsSN1PCOrBrcCuHIMNI3f511nClokn7HuvBJH1UrewHRph1Oby18
HBARoXst/nqzDbzn8InUFkvSPVsU9gnIwYxieQs+i5GIsDTPpX6cZEdI4wNjJcM2jpEpAibJPQJC
Exc8qdi0ugG9meD8SFjsrlzsJN9ybqdImlGeoMVvi9086v8qZf+z6l/2nX6BgCO236mqYXW+EPCb
/MbRQBQhA+Df5UxjgDgq33Cm3/akj9PV+/ixPiDMeLgvdnE1GwS6st5BkEAeEEAbjoJv5AE7hP5L
DrgBOo3i/APsXgT1tHjD24CHfFLRileHkoUJNUc4YYlN2AB2YiXIQTQ62n/V7Egvmr367Nq5+b+c
IMQhKr3qk1CnEaekwT765LbfsOwUKL5G5U9w1fx1fQBzT9MmPOUaECZlDnieZRHZAc2zT2uPE85d
KwXciYtncjJepL1VDFd7ByXv7WotrpBt1lC9SgEtDKSkhqBxi69GZuhRc40hYsDX0/1AHCBNk1T0
RjjgWM8hATGg/QzX5jNtSm81vr1ROdzV300qSOwj9b2I0TguqGMzXQi5RxfY04Bn7c+K7RhgZt7r
dTRcqyymeMk4kZ7hj3ynXVlFs+vI6kC3I/qxOmSXo/tz+I/nTEy8eksh+lqrxLauQpO8B/Jwa6B+
y+PEK2KfAzIhQKI8O6xZRK/KALhx8tQo9uHXDAGdYDllXa35TpQz40Ls4IH5boZaHFEYx2e/XaIH
wQDFvWYtEb0fOwuGk0sWzSf3xS21ibj0SiQQNjQzfW+sNJkyXBshhPShav/lhmLzlmg413bAyRO2
hgTi9dVn1KsPbzB5HPpci0HDxcTpbqQDWpQ/bStw00J6y37sqLUYkE0B1YQz7NKf4VZZRkcqeGRx
mU6Opq/bF4ASJVCsPVDoxl2Rcaz7dbIhK1Xb54ClEjOxssN25Bn1rbNi4y2X5v46cAXWbj0t96AD
67grUcslssObwz90SZR9u1JGpAKrn9VjmCQ5k60HBPrbZEewnzntOFoPmwYt2oEFujN5GbHEzYLj
1UeguZ/5JrVDekLoX8em8YaBynIz7TXlhmTRc0UgWEzQ8VKN/Ps8mXfdgoG+p4jop2SaocjJ7Osh
3m7ertu7ZnKUnabbwDQaloRL1PvNAf3Po39ADQuF/HQ5sBuQ8FjENOtB+BlPeh+AY5fGeoWVjNar
PGINHg46bSv1q2Gstl2bq5VGRWMaAhIdVR+Yv1pYrISaHNKsLGelW4Ef2H+sWRDijQGo6xv3xKhV
/3/5ORJWlqumSs+JR1/vIWTmuvVzNN2iOClfAVH7lmn894xk4GWh5LsXLZzucPSXQWvJ7at4vswY
g+tjzGIpq6CHXgqClzI1T/jjeXXzx7kMSlIgODwchIaxBQUA9oCJUoGDr2LkYuPM8FevuFHWevoO
f92ZI1Vllx9tda90MkIFDvwfK7NsrGVXEyfRHe/BKRSm9fIUCYIP6K+9oPpGO6hGv1JNyDYYktrw
UJ7o11cOiUyLVO1hcrO1V3IVhzmTYAc13zWbtmU+g9WCX0VWAXTCMRIX4ubtJBKfljRZYtlImWd2
ZFLL7RovOZunmAFK2a2yU42g3kd/7bp7aCTEdP2GAATrPeyAB4LRdYNH6tRNkFqc5h8AHChxVXjt
Vl2Fe1sIlZwwwb1kmFrbXrWLxnbBo9Wxx30zQ8oojVkQnQVBv7rx5DB243XfBILQxZlkFRbnp3Ir
fHXHNiSCxIykTkvaG/jtN1Js0GgHFAO89zocc/Ed7JabX0Nm2crvrc0kwU3lNwhiEdMC6RAf2zZ4
duAMMRE2iucwranr2nfo0wu2803PJogHWh1jnaJruLzMj1pIM0uDQO/8x+m07MTW8qS15Ij8n1Hl
XdgwmbQdBSFoivxHYjtSR5EfI4ivaOs+ZhWdpe363VsM+GQnwy0H5rBG3jAn7sVrdh4xKBQPMcr4
hL6PwUY/GUuOwcbPgxEqUY/BlVQX08hkP9TY5ByQ0hupRkO1cEqxrxRE39adCvc3pI8+n2/c7cev
O+vMKVSMyDFv7y5UWGe5cOSfphzRCUujffqFKmq7TDTb89r6CHdFpGWz/S2d4gV9aK+rUWkciTMf
I7DtMtzsjXj+dPU7069TUX5PO6nSyh37wtbKG+HLxFnRsaUL6F4ZwQOKEoQ0DBNocef41iMPEeG5
g62UutyzoERI+GN2+KbOl4Evoq2P8wYoMz3qtW1Lu/4FjkwngdS9uqN4gHb8+fRaUQXRK91VOHQM
4PF4537+NHPM/GaHo7Hgd9QTDrPHVd7brssIjx6gb7KeGkwdzc28QMVSghs2eGCxTKuC2Nu+mFQl
c1ylUwKzYwzxS0dJC/MFTG3qaTlfaWKkdU9RY7yxFgoo3za0uANoH+u7atTDHxKFtMWogHjfC0FZ
ppjrmz3ZCXfvw5jrfoQnUhT+ng8a2JQusZHBkJR5sB3R78Tz4CKcdhaBEU3uoIFTFOr2Lm7Z0jsI
k+sCny0UhBOdgYV4O8ileHU6WNVngMhVxKsYtHaDYsOnnu9BiXhPRtYZ5Laf4b3StEgUsEB9z1kL
c320G+w0TIwoddgz6mrXkz18VxDnaPnjL+C4N9HBzG3JcKf1w16TsbbnL3CnxwSPLU10XDcTX/Mx
RTcMxxRgLV/O5r9lIgORaGnbH6Xygom78qqdcCDYQ2Uywwxv5OK/17UAS/UkuUxhkvk69jWb7BoX
1YBW8cq3mzgk+3LBlQEhnqH6D9iKmBnangp+y028OAZwld+noKAIDDzE8D+VaGHABFZbHmmN5sLT
NpHfP968X4lBHurwE9chMRD/11ca7KZomftDR2Jq5A/1s9Vgokp3YuXagviZFpQK01qJSqRO4jd4
RRXnWyZkApvxFmlBJweCReELgtcsycdz363ZbBcoOf6WcfpqC2+qsoyhUKGQQBW7dMF31Sfopse0
d3xAvm7ubFVbmEYH+pXVdoWv9Txks+fGOoL6WZsl0y4ItPVJNzYDZu8g3RjWVLGDhL0wfUUaObpO
/p7Aqox9F3fwdUvLijPedRfx3Bnh/kixWc0K8QRmM9ytRwtv1ITLK/cPT0K4SK7DpulgSDlxDhYA
LtIUpwI1/cKNheroohZIJdoh/kHnS8s0SHHxZDZNpOLRAsNhSKtgkaW8HNM68UJ4McSnKStKuSBV
FTvPhYInh+gSHMg4SW9hleORGC8kSTjiloHf2D0mAL0oFkx2EFQi3qYF8P/PE+nTYK3O2fmb7Xc2
5Cet4h7TF/deymeaWJKhk3IOsYvQ53YsUyjL4HJLXxBGI7dEifcuAtLpkPp2t1Ff7ttceJbnLdzX
3vUDdm9bbCEHToFjtbgagJ/L75dfRRTVB2u4hLo/g31xzDdK4Bhwd0ZmwJRvg9aKBL+/QQOWYmvH
DmRXTeIQvcQOzpoAks/arPI+BflOYlRHa3PuhGp0PZbvKpkIrkvDjl0h2Yzd+f0MDtT4+G3lo6gT
9Cqp5g9/DGBrSrtkvuiBl8Qx0ewYciN40rUAlSBpu4oXQSLXnW4fS7JllBqqQwIFkG3TV1k5Fxtw
IH44UWeq200Y6yehLkYlb0lwB6PNX1Jd2w36LCwHvyK62D5Nj7Er2tVrykVJ8BE2ZRe5kxPzbQrg
rrrE0ZLAZvIlYrOo13K2P2tK1fPXrELPQLWufD9A4zyhFBNMinzT61gw97ElVvgOOLnhi22fCrpJ
+GYLrnVcvdKiCxpR8yNNgeNLScDNVp4isPwKxTSrEKMa9V2ZVQ8BS8wUrQOi1MRdezk8ewoJXfuV
+ektkbjKToOjuC5IxeCicziB35M1gCGlcUqnsizFAidgSyz39k55HeqLjv2bicbxCHU8f4d8GNyI
nTI4hN3rE4Axt2Yw82rErRUumPUO1cGSF05u4FMQzIPCJ74B1gh9WtHaOvjHbAgWlJqMX0EFahlS
2UJ9N81UipasY8ExxIweXgfm47TkXnlYznxuZjSc+9+fD3m9exQF+gk94VtqlQWPMpc+qhRcsNJU
WLAtG8uAjD2EShTWnyBkAtjMdX2OO+X32olCYQ1pHOoXDVsEf0c5LPd7BhGvGLp6huhDKLJVjtYe
h+k/04wXlm5+g56HGfQ/8L4tRPXMQjWVpr7pPDaMNJCz1ABTf2gFl1e2Hu9xG874P7FknZYoUfDA
/gW0gwKcyOu9zy30Rza0r9tV4mjGbvKtrAhgGYAEwKVvuwlKfbW1my8nuQSikHyJh+yCIDigd5AC
O92AP93FEJV+rp+12GGnWrk+i5ae0IUnFQNLIl30RysqrU9o3dj9t4Z2zaT1SY4H16PX1hO0Hb2i
sLm8U6x8aW/tfOf5BqCpydJK6s5Q9JR8v6sgS41JKZfBVpRWsWzzYzJpAm1/W5yHFWv+TOhrPgo1
6GvR6pAr8AZwJW3d++LHZgp4F6pEi5SnfZjOQgStYfiIO1Dp60XBeeATde9IlVRF0bZl8b9AsAb7
jJb/BmDuFtDPl1jxQqVT31Q5eizkEJJw0ss2Y6RlEgKnr7WIXQCgV5bk7CQvzA9xpRP30BKcBraR
Ft+PnHtqMf+iss846OuL4I6vHmsFbHQ8RSzGNjWMo6gBgxEKjFZtSjPLVB9ffhlQ9utb4BwiG7L9
b84gYd3GimpvuqkCO/gJh5h/T552BMfdBnxLeU+8B0XEsiYEdWlRDBSxsgbVm+jvVf8r9MIQKEQx
OTvXHJoDbSpGM6CFnrZ+U6W/KGTCc/pnZhd1W8/1+XUmyDDLEZSp0XFEfzv3S76dvhY29KNqo7J6
JR5d2ef9L9IhS1RGx6VJdgvsuFv6VIF32pEVxBM3gODxu2o2eAK4LwgHsCKVisg0B/LKCIhMJWP4
+wATms4NsC2tk/IVlmaJ5h/p1dsBvfxAbBB/1cemBvQ486att58sumbAmcv2pRTWBKfHWIi+ufgt
zTNOzF0WMSxK+YFcEpssxcMFXiNnNkb6Aqatn240+3UstJVXmYilg87tgo8UsvcWJXkWEypEyHqp
puYBjvG4NNt1PodqOZaOE6bhrKc4TSN2vJ8wkQwGr0xsHWpbGmMBc9kCSdkw9kQkB/pIMhp1Z4ho
M5Qlm3okGubaudF1g/D02knRuHaZaZKk34bGWF5nVdvuMB1IVblopxSPcTVVV8NDNbbgY3mNqU1P
YUDS9s1Hk0Slm4/HndWbEKr6k3DN/MJ3lrF64DV+ewGOcs/q8yNUemPv6jxNud9FmKKOhbO8tN66
o96pPuC5q1Q7IXlPUkPV7mBHBbUmyyn355sQNBQNgzIrvHmr+0w+tzIfmFGyXWzfRCbf08lQEQFJ
QUhiyDquo1tr6MKyBzmYccaZ+8Ymg84thB9VKQRVAQg4p67/drzd4aoBX0T38NY90pm14Wp4TfeE
Ew5VQljfDW8CfHJMl3LbRrzNTdewoRaKZhyjMbnhEdB5frjAnEMeYeL4RK0NpCYY2h1PiGT/1FJD
tVjNxP3qChE30/b0eZbL291Sf9Y0zk6cGzoMxC5Zrkgny4sqn8AJYMILyatLKCEUbMaGsU8xYnJ6
ZkSTwYO+Wd15nCMj12L46yFsUoA2euTX2c4OPikaUWFjmIAvzHloFVqV7lZf0syANOPZYXJKZU8/
0+4A4t7sjZHj+5h/F2qEzVqzVSLmmA+YPKWHV6nvOyrGlwOBrXOZVw2UcOvYfNJ+1agFFfkM8+PC
LPN9w2dvMzpfF/xLMEPj1EMnjd3arD9Udz7mWnYEALlcxfuTRFl8ISLxVSnDXx29XUs0jc3lWdUt
c1xCOI2t7ZEIVJrPSryePYV6r0W+ZeogB0Jw2XZ39ctwP+PJxxs5Sgrp9nLvoJfyQlr8Y0QZYUos
FttFYKMxQei84FaGrwtNamHGRTK9Rkpag075jUzrLYWAb/tJZebuDG4OI7b2Uyqj6+GSLYF6ReJD
6G/68BeqKYWlSU731VQ34XnwDmQnzU/hhqMV+AMW/9O79EjEwz3Kz4/B7S3VLpkpjgjyuD3QYQKm
Sta/Soj3Ey/Cmjlf0rKvUSCznBXIG+CntyicTRK+wbwIwx2i8k1yIcqkkT1Xwxhp4b9yKDHcPP1N
TuL7TFW/P/Q4SKvmn1cXa7grLIXPdYMjV+Fsn+lU7yYGAQ3Yao/am1RNBNB8/IX1XXFutxhOs6/V
ErBGJ1zWw4Kw2TApomVH4UvZZl+IDdv2BNs1fAjhM5XMKcFr7mOjGhl2TwxTK7YYhhka9l17kIfi
VQX+o3nAgmpwhgukpL2N7kCCsD+5C3u+yMFejgQDeS9jrGNjBcD8PRMccsQ1gHdCVIyBQsoOwRNG
1WVFSd70HHQjS7aPH8Isfy1VskrwPry6Wt75AUMPywk00TMtjR/26e/ix1CDTEfMdxvs8e3TW+sU
MZkyR6mqhqOyWZ+NnT1dNKMAOrmDaHwhPihu05PfOgX1ljOFAF47HTQ8vkGmSCjoR3Dw2+lXnJd5
vrwPo6AoPKJFg/HBto7m1QffZB7O9os7tcODeD7Kuq2GauKx5QA/fPugqdbf+MWABs3YvKWIkScO
A8SNqYv1TWS1Z/LOYYvwd2eQ8Zbdoxak7qJ7aegqx1rjZ74y6p0VtzN6dxKbvs4Hu+jY4WGK120r
uFUY7VqO8T9laCSWRU2eyD/DzUnYFuMo7FIwjBbs8qE3OHxR9//ElV7xc16wotYjtlBn6+qNdO9s
sdglnj3mB8eUSIOz4PxgaycAWhtDD76OMc73ZS70Op4Xtmuo/e0LejN/houxisVUtz4kVgGDz2eW
n/WR5taypdYihCvgE+unvtJ2MQbKRruhTkYcgOsxSL2J77WKiby3moaWze+nRNP2cfDMhdXIkgEL
T0tkgGIpGqKFSKqDL9rpJNvKxYqUA1J12fDT3Mir5st+NJi6BSRytLd97+DPQxK//8BJi+9p4neO
TL8Gl4AR7oz/3EXnzwPlr4OvV8RkjjnjTDk/RVRxdo9gB3Ve6MaZ8ibsU14EhoPqjCQsjxX4XXET
2G7m0goFnsp7g7yvRcnSCLLPidd2vg7DZmHW1mGHsqdV4CTANVzuM9Ed9CB09bkN+JgVwT+mdPOu
KqtYliY8GldHFhkO4ORevPu8C4It2SF3Iap51ur591cI2k7TY5hPWLBF5cDiIkUVbH5BzrMEwefW
aLvt9An86moCLT8t+FBr5agt0rdcB9hssvXBBffXTvjOB6LGtVtMpTvayPJ/xfK9495TXUnSfzus
rTWhckylt1nt+/mZMTKdT+piI9qy2QpGSKmzZiEoqZYZqnr/Ji9+QHDe0VRuJ3Bld2bisUpIJgYF
sLR4Oz6bSkNBcXBrqItWAV7A70AjBueQO26dcgQi8GYJF9zrcgdg4sPr3WBqpdVnWvk5aGQJgeqa
HsAxrXE/7p66xq5PwCR4Le8SlldWs/Gd64mRndy7u5j6YkN4yqiG3kIat+sAztACabRTUpvy/KQl
322yAlQPAAJMEVW6dBO7P3HmFzE97dOGC3Z05lx0/lHW/uTUowA4zJTU9xL1ebZhbzEoiiCemyjj
KpGqFPEg3n0VQ62ccX33N62nk9pz/RtjrNk8zPrGg9k1zTcA/sA+GHiCBYq1aX4Egq+h8Buj9wfV
PlX+XFbmQvTMpQG0lLxVj59rOmAse4qHI9mjJoeECU8KRRzXYcXR4Eyt6vePQyEy9aGTuwy8VQ/i
6c2jD6TBH911h/fmC9sKHnNQWw1MEYm42dRbu2sGVtmtqTkP+cSRVHQOlh/DSkZOm16Uf2EE2bwr
FF3GNv89wm5snQWeqzdnxKk0zXVekFKLP+5lEzEq876ELi0V/QWHZgEmNyxWUKizFfe5v4RxJ4Mp
YbSD/rC73+dSFJreXiPseOqJIeAsFd9OZlEdWw447C0JBZj+2rUPmlpda+vnWWGecFt6InUutjnk
cAjrxMczf6MK44hNAUxoyT0PATwzMSEZ1VmIQ4ywmztsMUbHHlg4E4aXXzkXui9JB9t9x886mfhp
uIK2gldhCP/qolH5yPr6Uv1PzzgKwehXxCkcZqPNkVnZLzBbxFfpVBTjUy4c6t/GXsaharYKqus5
7zfbN20hjyiRJa92Qnfi8PBnqcrH36RdnHh5ULVQyp10mNEdyySDNAWgy/x3CZctdqfRz1+r8Jw5
FId1TtSwawIHAhpGjpgTuK/eUT6Enw7q7mnW6w4y+0IoAtAn9K7fHMocb8PGxR0XTGj26dN7xMrk
4UiuCu1cjaOdfTEFvA1MnxI7RNQppWHHDUw6sux/Xs+llvAjvR/xKpsEcpGvEFjP1w2Wgxjj2QFJ
PLfEW6ze+Xuga0eekanSD7Dwz7Z2TD201RE7SCWFVphPNbA0QyyRKJwamz2w72SUt+J5gg7lklik
CZd3eU+J/HJu6lgFr2gDkTgApMUXgUO7G+JSZAgSeN/VGDo1Uy/UGD/i/OAMtVR18onAXKgeMxc7
P47p6rO3QyhOCzpF2y+FnAwYXb7FMQ9/9I/13Ozuug/+Ez2ma4w9kdMP5omnDSsqP4WbRuQ8Z81p
pC46u2Oa/HWmgiNnMK13iDgZ+32ikgokCVq4+lsx0HeDnnyAikxEyrh7LazRu68SqKsiS7Oc5D5G
+Ho8OczpmecfWdq7HRDPciHpckkndTV1pCaX1v5bXx1WG1A9Su4eCcaK7RbHS0GMGry3D+FLPnLA
Y1sprKe5cvBqHfhkhSYpilpH3ENIa0zg9+0S378e+/X323eEgNni87KWR8CMcWgkQOL6k1BUXip4
qXPBgpRd61J8jabsQd2SVC/M3+HBM+rlecynYP9u14kH6XRAamzQfjsp+3bGKF1z0ALyJ/G4DmMK
ZETFTw2na73eXvbq+GEHpp1YX0uwxu3ctxkeaOs+tH1673l8JtUQM7fJJGVN4lAY2NlSQZN0hz2T
PIAAyAjIfvkkd4WV6bMmYxO6n5w34HRsj8DcMXN/iL1RaCFITwN8ddLW2Cj81rE7INCxiikFZSLO
2fUUal5PUmKSQd00e26Nflt4LG5e0KE3clxmhMDLL4ilL+hJgxngwKxXviiSpCtRdeffIyuxgbwy
otfMQBDPGXNDYHa4UYpBEqWCOzcwhNnTQzHTQiN2jmjnye1aqHJWO/SZ1reL83hfw2ZCmnTT/E0l
fl7pLh8n15CD/NN72CfITWilvf++1NtCIZ4FkZUphINoiILRIJNrh/yE7CuZzS6P9dizCxgpC0L7
AQ4CFmeSX2UsxM6uKsJHu92IDIGB00s3K9Efv+zaCd7DqsdWZY76k8Ake6ii7srwAIcjNtqtEbVQ
IyO9mbILKHB+v+EqWIhR7ybQXgwp9SR7gv6p7nbMbR6NQm+jXczMRRD9oGnKTcKjHMKYAWY6lovR
J+e1njRVCcegaODyxaSaVLMX23ZmG4tKshEHuDUFKO8HLmw2JqghZMfPAkWTC+5YOmC7hnNX7Myb
m5ufxa9OLgTaDO1r3jmm4ILZPWh4E5XIIo4EDZWrIGDOr8OZiMhlXDQtgEbzAsZwb0TTuq1pgRGK
s2ImLMzvmwUp9a4JO6F7yM465gGlE4sMEFJvIQxCS8QHKpUJ2v9ly26e+3fMzY/1KCDCaG5YzoBQ
IU6DXVSUUlp63tKgPH6GMk43rU6Dl8rq5S0Dd7RxTZ3WfB3CfiSAU+Ndo2dj66HlKa5/ie15YqPu
wL//EJeW/yS2WTua3umDMppLCM393JpxHngRnkdZMDKuO3fLqHOGze+FRkf+NLgVcr2tyKCGGbXq
UV/LuhdgA24PLMN1G+2BNIweK2gOmMh2vzfjuiCAqCVEEKcvsYsW8vs9P+vao1zY+HCOjPUE4i59
5emHFZv52AHKzIisvSLDGX+/VFoCKFyuZMLdIr83Ie6up5DpYwQ/B9tJz6ew0RTLBtvRRB0RhWYt
XfGxdVjj8kXxyR3HHoOTj0ZR7zIMpuGthz8iGiMKUW9F80CHsI5RfUIssSC6y074gUOT+qai7HOu
UA21VC757j0McVST2XVmSMGn302oAmfpRqJNzBFyeBGqfMoOZrb/KY/rWrf55HiMUt7dDG0ZU7b5
hOUF2Z+QeA/9ttip8ffyDVsxelQdkoEu8tiDWDTmmiV0URicP96cZyD/O13Z+mCXfReWHx5Pntyk
eAI8+A7NiKQTIjtDhkvEh+JlweHEmP6J1ODIxaeJhchJ2uWk80/RxUGVugQCQbB4c40Q196cmgp5
tIvp95znF5EJY7X1YMaP9dFcMY5iiqKqZ5HFDhUGMz36jzml7rJdSP2hhb3YmOhK8l1x5gdGfkbY
GlxiGlT9U+eVpXZdRB/+6o7BUjBiw3Dc1GpBDeEw1bp0ei127RuLWd7wqA/zJg/W3BrvkBydGI5X
MyIIX+UEEWfDPur4XmCe4zBEyNggjGApZGhSRB6wD0asrG9xM4eDmWszK8hM2zKQMSQ2z+7DkgiN
8oG1BjTqeoI6uy4r7H/7rooyD618KR5oYOUz4OUVK+NmVcFWNrRPbrrE6qzmsQRE12CNiNKUglW9
j4p7s4kttAeRDJH9Wao6Nh/mRkXd6vfFgivvLJ8X+ZWCD+8kE03oHknQRQD5il7dw6zz3AfPmKhT
SSq/NuXbr1qqb3bETMApk3UyqZy1Du1Lo5oX1knWdlwpubbWa3WOrdh/EawENRxhY4bXRy5P7SEQ
U51AhQFgwMIXv5LeenQbYqULbU9fjKbXtKo/V+WXJzNnhk2o3dSw3UY/X4Z6MqvCD4eLqgNochyQ
XjM27rLpP4Ivoj/Z1Dvy2e2sDZQfWjuUm3zqacX0lak4HjQhlAE8Jx5Lk4tH68o8ttn7WasOGJvt
ejDci7BF7Vk49hQxPBfzQ649Y+OnnsyGIn3D2WllyWzABijzMwIw34ABmmMxNdcitKYWy9YRa7i+
6HUQDrwCGn6A5Uy22XuPpkSq0McBioJ2j9VaoLAAnP90ANHXoFtFL3Euz9gZTT+/FwE1eQhOycFa
3IFoqytA2VHGWz2g1OCYD1hJOxVs5px6gVBHmRsnYVa9AT4JWnqqM0KSv2IRmXs53pD9CdK114Oy
H+e6DrB3BP7Taq5LCqIW7KuYl+YHeZjaL5V6CrDARz7Ui2L/saR1t/ehUYTHi3xmWHY3tY7tTr6G
kwK8BTrhgUjyN0w3/J8+Wm1rvyv4RDUueronm7WJprbnp8JabR4fSo65feBmOWfTEvhApCyw8LH2
vmmRvzRKGd7q9uA5YNRr5PxcuIgeJ1i32gfrL2Fcp+ClTMKuikxMcnTmUZfUXe2dGoDXAhVgZMH0
b/JEKs4nklC6Iu22wLxbnqVgHWYTCxPykgx2FGH667Xw0SFhAIVKRyl22CAGa7nT6smf58dpSlOq
wyIwjn8+cuiwsCdllmFG17FAjond5kAsciBzuaIgLl/VvuqrcyHDQy2eAcBlzGqwB+BzszVOCzOY
Tgi2mFPfFtJaeEJ2H1nXqGm3jHWgW5fw0ZMYlLHtees/0WttRlqWidev06XIionqIUewSEuyMWBp
RR+Yc7A3QateNzPFk4DLEyQNsMZlVlto0Hd6YTFTiigpS5/MG1wXYfSYWmdxfMW5HlaCiDL2ae/v
Jc168QOBzfwIdoSuCmvuIMhRN3k2iepRJUOwn5lxARWc6HW8y9lTFAJ96tKbqd4s68oajMLZJJfN
v8MCer8gcS5VTRR1zFWwCRvftLmIg64TlAqtU0XzdKTnK6BbMcRNJgjZiPBRblHiXYXwrQorwDdC
RI1ER7SvCX5oSblBgayPaxcd976gUum7nwpXNKFrTSP/Y18m+fi1LIGsgQ258v2gKwLkaf2Ax6W1
O68JcoY39ZRJJlbuUXDExFFu0G4FbX7wZ9J2w2bPURG8B0/MWAGkI5JjbpWMjkFfEfbVjqSr2D/X
og052fB3023Tys+3rOymvu2BRHYbrPol/Ra6y/0Dl1Hcv9gQBEwNy4nSJ41mcILKI9gNsI7Uiuop
9u+1/eKHUjUWv4xIZ1hw7Y53vFYyGZMKXkOWxgTgQCSwIr3AExnZ+TuIdEZBmcMWMKqHKxQIQGuq
+YAbhsSl7LC5zb0GkzmTZmhdg9XoBrhHFOJb36rgyzlGVNvqEgLePi/b9vRDZw1v7DmLb6vrWIE/
T2d/WZIsLbu69kHbSUGCCJaloS17cxKBQh/4L7a3JGmyLA+YmzUM5KsF0LqV4VhSAFNfbehI8pTP
a4jgBAhCOQcsDG4QuOUahT2SvxE/m7NuBzHVj2BsM95hH+U4Xj5zn9n/+sljcuV4Zt8M9spSLi4E
GC3vBAW8/7wOk5WGrGpOnrwSRya89JD5eUO+BnNKf5aw0HdE9TACAJtH4pMh0a1Kv2sza89eguCJ
8MBijB+MpdgHrhjvMmOHcy16JgO2oZryygunbR0Ezh6E/BcH0JeaULfMSYUOQzo2LSlWIfGgBV5x
KrYekzQkOS19SgpbVOE1o+Y70Lz8FLtjsMyyu6z4Ar23lTi8JXF2BIfYTav9xBtlZOiqvc36Qa9l
USgiyIfpoyJsPHfGmDZZDyhZeCGfuGAlohEOyjxAZerchoDwdVm4++n8VS6i4+oAl87i/RIJSNYh
txxXt0ionciLL3Yeg7Pm+FWRzQLEfxyVPaWWjy0oUgzRQBnuHRzi5LvseVrAjqmuwYAli3m1VNxD
HjFvy2QWB5sAS3FBnZllG1jh4Mb1/KLEuBSv9m711luuNyvkLCsQqgTxJNndIzugDZ16jxdBp57E
mGSrxADNvhTpyTM3bbcvsdlUjlBHdJ7EQ/WU6//YJni9bXtj0wzHVPKUdQiMUXsK2aAKR70vQMEW
YJ0ECKfvVj/NzXbHCEyl4uORn8bARziBV+u3Qw87i3iq3gDG9B4ZdwHjWC4fFHPLhpCQDGSiGKpG
rhpwGCu8rAwK5gv7+RZuJuNFMtG+jbhTZ2Jo2ffdVrDxz4ksN24uItTKONzPecvDD512nzJPuxT2
bIOu6R4fGy5psA9d3EaHcZzehJ5jvzJ2zTOzicmo6HdBfEs1ucnaBKMbEc990gtkXBmX07Al8lpA
/AO3lru3THVD+H5/dwbGN6r/RJBCnPTRSBZJJFlfND0SnT+Q6QbFDQpA2ak4uznK26bIxCja6dBf
sUS2fi0X9duypYglw3BiDhTlcSg+STtG1K4R1oPauYa+B8rdXvYN7MoXDPVwIR8Wb2EWdTSS7FQ3
QQXL43/17yRh99D7KmveO9VMw+Ryt9qvuMRw/grKXVcecIfBz79rGcpZ8enJhxmmPtht1a+xcN0/
xPI4xsyTaKPgzN3GoPkkro2hFq2Rv0Bj1Twv1b2J5JKkXy5/uOaZUwjvJll963nKxT8gfSH4EzW7
ntoXetA9tJ6X5at93IIpZiZAfj9t0NXELifFNX6rnCYOFGhkYYXXJvvNSUfwvsdkXAGE6XIU9pSC
CZrQEw9ksi92/ruH+pANiF+wFZbotWwouKLVqA9SDT8v5KEmnk79m9YgSYXCm8qfaWG/PHtUc0c+
/XVpnt5g8UrQz+F1VAd75V87X7RuzCoPPnGxhnL28fQKsSV/fnU6/RwcMCtAoWePjBDHqk5ENFbH
G+TvHb3Ld1AA7cnCrb/nFoR9T1ND89jYQb42rQ3UpigfUWRBkOzkkP3R0qbBEDWkfQiY7p9ylYJB
PDDcucfEyl4grBtoDcvEkmSi5NKrmQuIMLCBsorRbIvmse49e19xNl+eHTXSP/UPaPyTMWNPnkNY
JYS9nRJnabjnEuPLOUqnH5Mbk1WUeR4oPSv2QzgyQ29zb+v5ELpPpRi0S0B/vH3lVoPobsyWMXxs
gfcYadPoUePFw17TPNfsn5bT2l084QEy6qLuadTbeyNqZb7+KB5ffh7AxiHMXrfwpVmoLR/BNjB2
fauKw+97kqs+Klo28x8AfCWcLlM+pQyV9LVC8cD3fNWpXR1OlqrhySfZsHhJVTL5bR/a/l7tOXRo
q4wQMPDXLVSVqb17Q8/vG3LIKIU4cqIjIezDyWCzrJDifKOTK1ZU45iMgF3G5bO34y6Ihmn+YFkY
QLzr8lW3cl0MZ8kp9JncReOkowGeERiYc7Z1Y78scR/rQyBLvdZ+qCbXExvC9VD9gVo9CyGy4ABh
exxHVMLkkXHkkpwyPlxNtQxt3BOVKsTxgKX3x2881hiun1VQE/oMHZ2ioSikQqzjEqc8JytnS1QD
qWuuaFufWJbTcPXqryy/MmhqEvDd4x8nPfaOyg2AqqfDG0Simph/DlWn2j7TzoskB0jDRL7dKHIn
wmmPEe8ou1Ku7hn0aqcSf+yb7sMDcKwJE7FZA6k1hDgO16FstX44qG+rJYayE5nxX4IFXu+7bLeE
enKmT/nbBCmYBwXlgJtxevnHUqJEnfGzWOD8xWpJnvZifmFv01hLMxxpDUk7kkw1GqWr8N9mYOu8
SPSHFhtuR4lVcIy15ImP9F3kKE/DAapqKHa3Y/RIOpD6mId81p6IkZotfzGzwv748gqluzk3piU4
VRTMycMhe9UeV/XrVt4ongz+y2U+Act/h+oIIjUzgPI3eVsVuYssVPGQuiFiILmrs1lzOs8MDq0L
5hzYswMPvzdZs64LW7H+DCZawIQa4F95GoBCf6eOUrOo/A6xZlzO2SbXsA25kRa+YkJ5tiVlizzw
7f+3tJaP3oI2KTjlGZtt0yf+O/lmOlDM7MEJe1+IqFNO64K98BVmjO2ADxh6yE50rh3yOhcLX11o
br1dih0rWUyZozf+K9ZoHFbrOnDUyZCjtgtI6SzqX/3kufz9SohyD2HTy7wQpkHWS/tcIVADk83T
JXWsjNC8T+R39xlepDTP94khFfkhBotu4CdVTFHLydfnhvjTY+ePt+/U0IckrEhKRCf0l0mYyjsm
qIkhs+8koLZ38brNfAFnIru4bAxz0KTg/57OLa3Gymx6/KpTp1P+w1jrTZx7kp4LKkItC2lG9ws8
dRhIyKeLEpGcIGBkhXSOdqdjncD6HrCdazoK3Y7RDBh6km2RA99wQ9DDlh8IcX2uFgVOZqyEiA5b
G0YzD0f5EWVMtc8lct5r4J9IgNYYffT9UrzIwO6Qj1+cT5zOd0jBEU9fXxyNf4J0Ime0eC0mlOyy
jSD8eeuSRm2dXTtueWmXz6rUbVJaHc7j4/QxnigvbGc29OLZqhxzH+GN3QxixMtgJLcH6jOIpXD7
4BOSLeryTuGjhV456RWaEH+aFxbmZvgzXxe/1b6ixkEc1eIOzKRLH/XxyU5tWJZ6wlaAJtVTHIsE
JKnVE6mwb934vSZHibBWYhylaX9v8eP45ZLZLku/UCR8zn1d9lANE2uX6A6fMacPG6PHxps0NqnX
NcagBfhgZhshR5/zhFHVAr4g2G71j3w+6eWrvmRjvIPaZ1UUK349GGFek/S7d6NYV5OzUWqp9CSq
BmIFQ+AoXv5ro8zkgxt0T1vh5fxHSgKvKgDOIDpC4E6IrvpUAA8cRPWqkqYpzV3tyHM5sQaH54/F
PcIq9m5Y6PyacVBDJYyJJgoBkx9BzD/b79Z62PMPAObPkuI+YS3Lmh/SrbaB2qZpso+70L6s4Iz4
D2cN3+6xQbJt1HBafeCeQm/fG0BBB84rTTJ0jcirgovv0BggdcnKL5P4izmyDWVn5VB01Z34SOjG
nNrLLQ9eTe5eXkb4zSuctJuRTkkv8xGZaun8rUFkI+5CQ/wk99Ro6egOvCik2PLLTB4GRw/hRcvx
sDvgGkI3UlWN/76PhCC2OAMKTGFg9hR4LmZv40CbDuzFUUPt/Hchd50FMh+LqDLVde2Zk7hmU6gE
hBXMUo4EEKNG41aD2SNkoV0aasLkXReqI9U69Uh+TUCeuoBz/wmlzAKMGYYNegG/3xhNwhkLQkgt
SyrfNYPe8QUBlqZWKjMB6aYIsJfHz/MwjJ5UfJGN5AZYA9I5G0YOirBde5FRjf7GKm235wT4wtg9
LyZJVkfRM153RzDQViryw1aGjQhIF8Ifcwo9WvBxXjooXCs7VPM/5v1fI1m4mj/husBrcBSgwoEW
aTjAZGdhPJOs+G/4Nvi9cJZKuUImwjvWzMtD6Da+Zujr8n4qqy7HdBYS2rvXAuAzRQA0XWZHYJ8C
LXOlcahNueyrHvUeucQjl7mz22G8r+UDSPV98CWnsRIroDibUqczhTdB1TORXYo+rcoPjtgDUG8W
Tqj7jN+vfABFB76Lt7Aqn7KUnBLvV9l8x3WKe5nap840Udc6j19bxy9LGppBxQlHyeYCtcTqL/ir
H/Md479I1Pr7Xbd/HKBGtGuF6jRIAvPilNbZWpl5siL1za24B40cxHX0aQt5IswnyjeotSFMN5Ls
lZA/4wNt90+cV8ABuCgzauM3hX94wr7f4nNWRkhOI1lKU4i/pH5Urt8dLJZxO0XJaVBgxO65iml1
JbYtomCutUMnxSAQau1tPD/+a0JXeaDt8M7As6TU8qWPlugcZ5ig1RuWPdoUTnT43EY67j1OAnDt
ZOuIgWlz5yhb1gHTtoIH+W/lev7bg0RE1tEZONWYGqGpD/WeIMxsX9HFi8/lDx3s0Y8J8stJdJmc
7vT+VIuwuRRh8sNz3XrM622cdfLuG5I+47XC7GMb4qU3j3jOQc9Jf7kaWE+gQ8IJAXJWHQ8yN1Ww
nUEhPTCruKj53uBRqmk+FBxKi+UU042bgabXdJasnJHqHGts/ZfzXyI8Otl/qaX0IPeUoOWiIhlA
WSNHp+z0rW32fw06XDT+2TNXll1SceiGUjG78j9aBn0VzFCdGT5wOU5bfdNFfG7sBLLOsR+xFIeg
OeNqLNhILalhfrFbpmDn+dILR+NhULP9xhr6x3I6/FKzD6FqZwegyEJBbM/4+oHDrxBY4GxDtOJ5
0aJ+kMAHi5xmNKwAWR82zKwsn2crdThdxa8J+reBFcrNZWM4CWOm9t8A9RRLeIjCuTdQ9PuSj61e
GhrjC4iS0l+v8lh6eYt9zHizARj/pADkPcZD7cCZLiiZFfcjYQ4C7cP3KPdzn405onHV0Rx3hkE8
3mlWpYwfCDG9RlaL77I4AMlWG0xccDEPsEqXeIUbc0RFc2tnVr5XZXZ6OEHq+7T/Ohk49bWbGpAM
7UrFTRrcH40M3UyMO4hKE/K8USCj1/ql3+UkWi0VUy5vFiygKM4E6VlZ5xT31matXstXJqBsrtvb
OliQXGG/f/qgzNcim3oAJK3BANkfRBHvivATs24TewYVUEoqzwAZythhLJHc3xfaLnc2Fj/4Dhun
Iz61PzJpp9jtwQEpZdeHfJjbHle6a5hqBKsYT7YXrRnR9cFEWYFj7g5OupqfkNGvJccOsFBvXnzV
nmfYyO7ZbslEtYnnRkZ8S92TzJEgNmPQ5siYyMP0ptoF8nxXijilSmZZQBzXPyTD2K2CrNXyFtsW
80ZGNwDI4j8DuiKoRoNIFynS6Kxc2Ega34XgHkUbx8uS8nYqpFJipxBcGuTcQXyQm6XjWr9QwpJl
cEbqLqy/2+vqdyn+ovo894DEgZZFW8n0+M1lNEpTZzGNDXm8oWCjp6K36lQa94+qUW+yCEwC//yJ
XgoVnd1Q5uLnAzqr2Zohc2x3m7a+oKmER+irRnxpXviCmz4wWjyIcSPTI/95K50ph3RNp5bxz4RX
PRLp6nbcglcfCLoQHqvlHCEVE13bZ3pB2xDKmgKXgifQn0uhQeLvfuNM2Br5SGttucahHaRXaD8p
vpMKcCpzajHnPpUl5V8Iagis+xFQXKwPIzxDRNzrEW1bPG3OaFO3jWcIOFQyqUTmizVWwGq8Ump5
fmC0LYEBFAQ5XFLSnjhTovuwMb0ILoh72WW1WzpgXTiyVpEhBKVBlg6hY6soP1gD+oDTsgXaI8uO
RiSsw4rrdVWXaySlw6rhlMFGXr9VhLUhxvJGHQvsC+JXULx51087DFwREEY8uoqkQ5AQpyMwvevg
zr7rqiZh0DaurbTVsXlshFPpJJm5IztrPUzdevhlI144rUu9ZBnadwzJloc0fOlFEJNLonxHNyJm
AhKzv8rHRk2HCjJt+GPiHwRrmSmJryeRW3K1rFq455Zcg0Aat0jfM8M6p3N1tiZVw6yF+/mLziUS
O35eNVFrVSHuupdr05F2craQ/MunCG4dI+OlIWnq7W7bAHIwQjUFxt6QQgzL6MiCnv2QVQ7Grnkc
+kJqcY7Zbw4YavliQU0chmSF99Cw+MSiiiEVGK21ze7gm6/15PKalg7DLAdx63idvD5NuLPqe5iD
rJAdP545rG1EgvUgzxKOkymBDiVyU/smSN35Q6mxZPRkp/LriLb62e+Wk+Vgk9D1GXrd0t1EwOlg
xM6vw5Uf3fKIi+T+qhpGAAt5RC3u5yIkHJwrihCPcryAqQWlpg/AnPEGsEa7LXofLwRkp3VLhPjy
8g0zkoHEZo1YFcoxlpVOcp0qJi9dY/ab3E+aU0dyZOz6GcdC+gtbXE7hdxpagVQCuZZ6CvycCuWe
WM8+tbGP/YP++mwdBjUx/76BiR4XLlNHD+dpWZ2emnqjiYhUZXhlabdUh7q5pzX5XkWJXWT4dY9N
yjVNuPkNUOBsD9R+goSK41l47+MAqdkasppuqFU0g/l0ICzTOz0lTSdws8uig37qVe+V6IkegjGI
3aG1Qth7Hk2QjQwnwlTaE/yH8R6YG+VzPCeQ5Vf1Wxu0cacj/FsLTTNXDmr5s2hQr2BUhpXCf5dF
a+r1ISgHGNoGYK9D3Wev4b1ZMBur/Y70xZdSHtOeOnyj4NnjAd6aBZ05AXOhELc4xRAcISoAiFqW
xx/Qmr+Mlts6s5jjT0CTFZBA4aJChHrEKoT45Yfeyoa75Lhb3bfeGwVbEyfiiMaCsM8Qg0LWVwnq
UkPfwurj+QYYI2uT++PAG/4t7tvnfya9bNQz4/K9UxIoYrU+4tK8jZhukSVfUszc7q7BeqJTXJzP
CJx1lH4WsK/X43v753ghUdoDvjX+BaF0PRI6Ag8r+lNJwGst0u3plAbffZQQjStJkZTTvjPyqCUq
GlZ8lxWgGdT2b9awpgXWHOAWUUAXWTepWsG1RaUU3+VNWKlSo8AHGV8Bbd3gkSDP6VvosKD4OsMo
tvZKbi8BF1YinB3NBS6v7YtiHJ9U1HLnYA76VOtOK5ZpFqD8HsyAMRYAvi7RGfjGdRoTNYeM0xKy
4nVVjrHeX4TFon3dq3A1wlXYbz/Hr5xQc0Gx7rqgXuFJjwi9x8tNeiee8inks9R7GkMHJNNUZz/x
fX5QgPLt6boDDL0tq8cjRf1eNP50p2BPe3ziIcEUyUT4EYGIR78XbN2HVd41U2wLCUFxXHjlWR8+
+jfHc3AkyEFUUx6izQSz5V/4umMcQr2wdvhz//ZM15D6L/TvjFU0e/U5EWdaQmd6nL8gvffuRjXl
tjdgCUCZd9kwi66zXh9kdtcZnRdW9ggRVHVGuRf78ee3iAyDat+ZKuEkg81S6sCpp61scLGVzrix
zh48ww5q2QUySp9/gA/yGDrkvHWgRKWcdRdNyISjToGLvy7MjtPSqBx/ReEcELWHeNKKYQBrsMQY
HQWqalRV5exuqF9o1p44RmnVCLN2RKfMJggFM0fkSJ1nTY25izmYN6qZqLXbgrQeVIm0tEsU+Aga
ZdZNuTfut1jFmQq8ErA2kxr/tOU8nCVWfxOleHqWisD+AsCcyPLt+A11OyPwDn2RvXwZeUU/XQ8E
zRS9i5edhNZnM2MGzgrVVvCVEHSM1LsrnviYAI+P7yXaHTIXVPKJmbeA2KF2m/zlIBQ0kSECUTtu
Fqh+FKR4GpbwkWjdsuAp8XGTJELFdV95rJv/V3MhYy/sqOw8SlKGhN0ErkhyiNCLf/B9xc686Ox+
h2pVgyHhSCaF7hseWPTyqvCv795P15TnaWRtc0i3ATjXBBbCBZ4E11kUdnbcvFW9HTmhKLZkyybw
eb8StSgFEiY2Et4Sr6hpCJD3FMULfK13gbMHDqZeOZOMzRy5UljSS3DUuZVEnbpf/fXNu1J+T3CX
3gV4KKJmg2DIQIzumqXuO6bbjgRTJvRzF4pm3bbRYKFd8WUt+HUcoWRrMWyNM8w7nWpw4+4eNNrK
qDavr7sID1P9ros6YyQXtWKaRlr6SdAX7UGzcXd24pZ88FYzKXINN232rTM3PscZbr2ggCE5glgZ
p/S3IZ4ijP8Ud1p8GBqH6T7CAFXySZwCH3DhZITib/a+IQ6EMk5sV1qQpmOyadbbwVJ7EntlzrdN
j9H8sj0ae23cB+DK0R9d+di5tPYiuIxaepYyZm8ag+rF5ljQzwCG2KwQXGusYjaE7FIJdc3JaZoD
bUXRQwyynWxUomE/VS6qQAze2/Tl59DUi/Waah/mak6KpHQD3h0Nfs8W33o33Pp4Z+UmStrSAjy9
BkXDgfAB/u0SNPlthrt9vK08EdrrVfbJbVEh0KqhUzoLoJYgoAcw+S2MX6p+qRH/GuQFKPk1h5Qb
KPv6vD2fg68zGmIHcP9Y9Aq1cZvwn1/D1wBustPD9QETNLZNfA2PUAZkMs+f/25E6nw8emTniZEK
nwBZSlIWFKmMWSiw8TBG09k1+inINUZwY9ggbzCIWZHYDr/GuaX1zqzHDYtTs3tualIFDYeAczBi
v2VG5ngqQLZQ+gvq7yXmvSm6U6QuXWYODPT9oDRVVfMO1a0EjDMRyL4ICD3oqtdFKSOZmuQQoUgX
J7g4PRQl8ojw/QauPkEkwcaUT+uzumjHb2RPG8udOx+baUPSeC4+VVPzuX2CQoTOPLz0i6sxZ+ip
PK8lblA3NI+n1sJtdeYRmAEZqu+e8dEmNF+bYwhS1hRrZt3XAjYnIbYclQZMz4Bn0RcqaoSxn5mX
1K1QjLFiPZwTbWemrQDOM6IRQMVyG7RPbMIzt7DNmWbWexgCtlPpxr5F8DwbkiDVCP4vYAS34TcA
e310gnPRLypW/brO7TURmEsFTvY3SnZIvXucAR2BxbIxJNY+Odq4LKB3qX6MKGjg2lhWMXudk6Lc
XIRUvtN1AwLYK1+togctd9Lua2COpmHwwrnWkEIbTFGbHW51V8KhkATMrD+ok9cXSplHddWn2Hor
Wbv/CNirR+yCeWIjXEL2cz2kLmxbipbqIyljQlRcz+cfqCjftD8rdoE3x3Rc2M+b5KqvioQ7q6qe
GX5fPj9y1qRrpXH4i/+cHz8gsGiL9E3vhPEy3JJHLsVdCg8FHyZJLvgUQkc64saL9QG8ntJecvnA
KVYEV+tBWfRl5zzXAMDUX4KKs6/PgafHWldMXCL7t4Qg1v1IcUMehOMlkWsKnpr7oA2vhNpuM9J6
CsWwRcCg/KXSEKop97fKW/cO8+45zs7jZZErSXTeRshufMHtfDYKQDvz3WCdnqvyDaMs8xzxZ7lE
gGY6GYMP/H2UOY1wdTHiOYw841Jb+TvYp1GgNTHzLQFmdoDM6FIuaCXsPgpXfUMW04vAJ5CJsCEY
FlpfxS2vRwuvcUkSB14FZtFC6Cbq/kRy/ErZE+dilo9AgYG5zl/DX7ZemsSdf5yCX4eX1sOZ01cm
RoMW6kTurG8r77H99pswCJt0XIdAIvC54vKu741OXhhWL2N7bcxxb7cqBVg7ss9Fu/mnba7vxOKf
Y1FLseDx6kSfQrdF1eoI9xsozA5+dXYhW0LOhq9V++9cbN3DJDfY+F6JLAZ56+pyDnZu2xoSH3gu
ynOyZkxWm9WJPMyy3O/tW7FnAdZcNdhY6FMaCnFtba6fsRBH2PTmLQr7kz5jwl9204+jwCmlA5Mw
4kOMF/Le3fRJaqusEgryGSEl5gdqjI4Y79sLtwJyecwv4i7Mulz6tzhVk28AfdK4rHLf81rRNOnM
6CAeffz3BfNRlwxJvMv+3r9bJ6OMYlGDKTLJVBX/SPCr3UMcJmIj0jM10NGsTk3n8wT67MgMq0eL
9MZPvfYBYwHrbUqL7/O1zkMoiP2tMKXDpDutjs2n7YZyIUbtdTGrYEF8XJud6XzJBkdjh1cxgO5K
GNfV/lne//79VxE2loQb/iPoUUyRl5rXSuvWbBSh/jmf+2EAj5hdRSQzX8nETDADIToJ/MHPHGI5
5+Jm8XosfB/dYtOxy0Tsrlehm29zvzqaRSf2EbZrjYSkaXXx2R4fgjBzup2/+/NOZvKwZfqM491a
YLQD8RfTbGwLvRZx7p3JKtOAdNO75uVsV7RGZX5yi3fD5cVsbZFYDH/Dd/YpCPG5QEbATPtk9ctZ
SuDEfOwxznpTXnJ4pCk0qy+eJq41EoWunQpqebVLfLzT5kupAl5/uGpgT27uVtQcPIDlNRQNHQHL
cxga5VWuPsjin10GIPxgRq05241285hjLwLLtD+lJt7gQ3HPAArtmPcrA2mzrk8ystGegi90QR3d
5tOi46Ma9xurjqy9TQQpdMqTgMfNXhjJHRiYTH5t6wnL72QBCiDWRI2XArDlhMMcWqItHQymyiuE
g5B4VScWIVH8YKVrOMEL5wBKfQHz7pa1no1T5/v5IGLcFPX5MgU3PupbSMRbDNE6H2c9RddlgZfP
xwcnm/VNt9s3rF6MPTenvEfyjsm8GmeUHIawdlQJgQNKtGJ7VoldVcZYFJreozLk0DsCLMY0t5am
p3KYmfj70CTEoX/RIS/khCiaUETLByiA2Sf6VwclLrOni0MU6inn8oJ4KeaBh3n6wMV8ri2ZQ6Bv
PwW8dHFpW/QmVyIZGm5TZD/gLKvhyEmX3XWcl4nSf2wwuA/6JIz9UDr7doHqk4rRG/2/Uco17oit
e4LQPv3tauPaUQY/dp3+yfHquR6OuU/xtdI2KfBycclcB97msqTlW3FnVBHhYrczKudzg1fc0OwJ
UJgrMBO0YphHkPmVqo57YCJolDzTnRtNMQakWi9M9GwqT+Mhj7XEPD00j6HAwgMc7XO5s4HJMG4z
+kUjnXD29L6y4yTk/Kz0iVgz5agYH1qZo/Mtl9UFxgyv5CxFSUpoFlZwc+LwQCCNXIyFXpMukQov
TkoXqybz3Qnu1Tv/eC7nKT2A59hogu5p712Xq6LsZuw2WTx/W+FCeo0MYCRgO15rUQeftoq+8v9O
15vtc+7kazoXK7VGEGqKxgQ5g0z5PR0whMPMEG1CSsJ+lPuSRZv6YStNQZ9xLGq3QA+5BrPKPigH
VXduEle9Yc5O2YDNsYksiNAGIdIV1ApB5Jd9N1KxC0ZL4C+Pg8dJk2+Era7PM2BT4Ia3xuuC0R8c
wjlOCd/PSyIk2kTeSOlo12KktcggKkaQGEXlQKd7BpcrXac3b0MCR6mBrFfaFgQp0djOFaK+5HY+
ddQmHtB1qald6RntnhoJvu1gfQgft30hSXyrOceJUYkUUqcfFFLsQiFiJsg6sj+M1e5fzk2WCNvU
4lmUJh2aDOM1hB8snnlxMB8qn2wdrT6ld+8j2SKIKFikAAisRY4Hx4B49txbPwKUQJ1J3aXLacxa
ppsxmUrxm9a7KoWvk4QxIjy6iTciSCxh9pHD5InyeEePWy8M21y6vVaAs1IgU4WuqaCZRORLYwO5
CWa6thbxYN4IfDHgHWIceHrh3v9Wln/4WxVlUz55KlOOgs+86jasyDE+uVRA1nwdfG1BJB9CrcGu
JSmzCGZ7MplGc+hxxPfZlCG8Q/J2rHnmkaqDehGIO13tyt9BaVm7YcpMx+hz4c85RpdY53/WPPbp
7WytgnW4o4s/dfYYlEiKSMUdHocsskCSzRaCzjyYd0frAuLgAFUaA+I71fXXkFuh+XDu6237cWsu
AJ5oF4iZR/C8LD+GgFwmJ8vWuUTNcTESt5dMQQZ21SmEGb9sYnDMIce8Rl/kaT8ELor4vQyQ/zJ7
1mxyVGLyy78ZNTr+MHFok7+IjnqP2oVe8ycvIf0GU66f/1yxkqbSzjtEXysq1z0JT3GVq9ilpO6Z
vVjbZsf1fLjxI0U9JnLVRBdzsAp+GP+8VxVGoYcVK3pL/q0iH5P1XUpcIqW+KjdeSVEJ+8rlLPYN
Hru7K88MoMa7IPMl0UtW8xA6c8Crg0jXfumI6huzUDBHwBj1Jfz7lsc2fx7PTf6CE7A+lxavEt7t
c5FKSoh3JfYU31vLAYSClPJ+esEN21Ryr13kRRXtZOf//k+50B/tG7lYEgunnpgPQQ0NPufpIvAA
e2xCYfxAEkGpIcOByBVMNm/a4M+Bh5+Oxy4BMgwUhWNVicemNJrfixF5L1EuxSNW5fUE/AuWAO9Q
I8MC58uTVN9Ah+BMqjTB1PxmnpLdnOaXk4bbyOxBaN62/RP12qQoyV49GrTiJ30jdq3yC8t5VjnH
IqyKlxskSFOK0446jg/3YUfnkmyOb/TueFLSdIFIyDcqJTPEYzUPRPEEBv4ArAoEfAhrimgcEXBi
N1f9QvQPtmNuWWxr0e2JE7Ou310moh4sO/AvpDVEAkLfiAuMfVtOKpfdoFJkC1IWT2zAlc7tV02f
OvLgr4fVYr6IeOhdksYpup4hfbH5BE12Oe2jumaPR+PCHePS4jimw/MzEfjvgsOZ+lxnQ6lAj5rh
iv2Eli44GRTOGvH7HE3p5baFr2HhqiMt91zubUfHPghwk2PWNs3oX0qOG9EJjPS8Kt3aTOlTcLhA
SmNjYRKshVMN0dUAZqUxyqclVdibSSe53tGPN68vMXaebkDT+mu4Oak0pZNlLU+SE8SmJvdbabjv
HuStJKApXyoqvQS/uXjSVjTHUE+A2HPLIhPA+wfm/C9FvZ58GLWbBIowVwuWaTGdMeiwfomCIQ6D
ftRXXj6ftCIoYjAbbkWgWN1au0Nct4/6FV2eozDGzhpT+Xffb/KAFO9+CvXtupMg8p2qmFD9dkLN
2RTbr+k/pxSlUb6erUl3Onv55ggJE8UhPbfhaILCcRQq5mscAZevS+8KyPBBFNuwux8Tq6h9RJ3I
MmmPcmClLUC7ZZmxRJMLHINK6AhQZinO2ijfNsW+RbOKzaz5oUorTiNrYwjNdfUGTRUHB42uA/4W
8ZYkvdqiXLY11l6Q1fBf1cpMuS1DH/vnwjOpFamHMM+KVS433rxyhASuUyl0g06aFSfl9xG2yUeX
8gBSShUGSF5ddhWJFB8Cx8xtZbI+d2Qj16NUw3KE1raIvfWk+Uhi2AlVbjK8SX+uKCMyrfK/Ynwl
yjuGLp4OxhbpuwVwcEODm2KtxyUhrc0W5tJDVPuRWck7L5GYsyO+ZX04g2bu1EkOxpDTfXmWCrJx
cLFhGaaPqgVsgPJfrWWnmEyGcxZy4lgr6Kq7I4M1jj2SMGC7kdOt0TRZIxS5XINtz7Qq8gRapQxv
U5Ch6Y1yIy+KkeL3AahdCfnYr2DYfa6J+Ar2/S4uIQ0lt67a2RVyrWQQjIY/g7k9V5ILcDHnKN3c
IIjnSR6CStTV9r4R1XAW5oYd0VpJFzaRjPeP9kpZsGlAc0G874ZCQokcyuuzjP6XHCe3/wyCtTDV
aZkFYheYbZFBpVhSu6AeLKy8/rzKcJZB1nwIss7eV0fD28DcxOCM3Ho1aXUuqVktP7lD9sNq/Xq4
woFBlbXD6sZF+jI+pvbFF4gzw2+wZM3td8ea8QMBBhFRlsl5C2bZHIIaKkDrwTatMBK4lIiXHfao
uAlVuFU11y7kGBQQnFAxnZwtdnu9H7zw5Bww32wShijrPhKmEk0glGBbN4YqEvq2deoKcgPqEqUq
ce+61/fef8biY2UhhPeezJzK5UQlw8qTBF9V9gk4LaCZqc9gV5q1J1HdleO/c/KhTGBIDKYgKKoc
v7rDw81ZaapEmYRDoS44PXwMrPokJdd8+xNB1UB7mRY//9iD7yyU1FJ1rxvRzPsOYxZ0QQQxpm0G
8d2bpYaFRXfJDegOI2XvFa5MCCdIHAJSTIam3KWxgY0z2BIxtNIW9p7SPQ0GlLRgCQ+POaqfvSr7
sSUj0em9lhC7QweqTHUIXyGokTCfignXz1CVpW2PwYXVQUjkPBNO3yrXGrs+uKeUl9R9hWP/92Vh
YBb7C0hUwKcByILrB/TVZLmAw4nmXxjOHYPAz0jpOFTFCRukfNcSPB1jQ5FTaf9KFOVikfMnsFeY
xu6HzSO4QCbOBgMbDBwy5FHxosNRvPS+O8SBXVIZvaUm1FHAt55l0u/vdAEULCDlkZwkA9cbbdNH
c7r1kJP46fgfRm7rR9yfBBpVhVqIZIvjESXzZa6AoOuZq3LnevBdXsTXOI2DlFJcNs6ZOjshjcJ6
WXBRCQKUiGiLAiRENUHYXiy6w1LkV84Be2H1y06RO9wxEZldQi0EU+kRBIYv4bYiD4zR48gpx4qu
TABSwwfQGuzMuOP1gdaGIVGyEMm/XQQINBiu2OjFei42YWmNgmvDOoQfmdJzZlVc/Em/KufkPEQq
mE2XJ0lBb3udpeQgE8x1YyxPmnM03P9zlms9ps/NBbT4+wCJopaZ3rCHBpBN+zF2pMRwNPuvTPL2
0VAs+gK9m37oLv1oav7BYqZgoJSeDhadVwA5imoWdUL+ZnPUmAi7S4o0ecOlh4p1+D+/dV5Eapzh
XRiGuQna+Eim/F444pbv4Y3j8gClyU79M98uwIZB7st5DuZ3mpilIKCJJRShmvjyvjNwll3Kq7Pf
A3fEt9NwzhM2kZjbbhlMN0awDEaT0EHAL3P5XfPfXeIn368r+6g4ytX0hXmKXvVBk5LQfSA5xsFP
UyE4v6UZMBaHbIhDfQnKBNVvYEKs2OZ+gMHd6U3bKdJGLiplC2cA+i/PZFq4lzrx9bpEJ5dM+6wy
DnJyqjboT1sPL++NZ0arIF/hHUzM6D2SPdSHyTDQ6pVvNu7U3whDA81bxnfho8A3Jsn0Wz9914I/
t67bILhrRBtPqcmbENt0ZoId+7qrtwqVFaVeIcFj8euJ7DEhkifrlTmezCzDbLirf5wZUihDcFFI
pvZbmFf/3Lf3wrWOrNKxrGXsFt3aXJJ8RZkv4WOOtVqRrdtuHsUgL8EMO69BQux1bV69WkdwkUde
wmvWfU6KE9R4o9vzmdVZP109dhm/iLGtzyY8yR+nV35JGi4u46EwIbEwTj3UoPkFx3gQVaFlIc+W
nug6fAu3M6VBuqOHw74Dt0BWgZ1XhrSa9BGx9+sOj9Gv+RX9T1cB+VclHL9L6PWXeRrsRNIuyRDV
N8TjErOXbYuuytnc+E61ZEQbxZ0jIko8RAZkv3i2qUGQmx+0ucEVVTDaSS63Kjd2wGWh/lSDmI5g
smJRmsdb5wJTOoXZndxqKtBn/OBHRY88B/rHdu752lviCXZm9OoTeekkSwh74xVmFD6VJoOsig7C
+P3Xi+1HSN+Zm07kCrjMuyo06D61CwFXCa4bu+qtaB3kLCJq/MrVneQJvqXrVs/WJPoz7mtqf1Ps
Z0Z60quWu+38Omcctpn7ExrH+CQaGmhU+rHLsP88jNkDpNJjGcVyJ3bhGXov58VJAkbLukGsgG5/
KUc/ghxdowV8aAeIxmaF5xzoZboNMDppzvfyvAi4L9NKkZxTUVQeF1yKV0Rm+QmwDAVv6t7yXxVm
spJ/BmPwrhofi3rsKngPHhKHTuoMpu87I3+prtPc5c7VztTX0hP0LVGMkR82WuEpULLC9DC0MbIX
BE27yd14vziN1UaN2/qKFZX6j3Py23XyyAsd4oj+CVCMglTFnGhI/O6iwdKFsIYZBEdVkL8gxa3s
mGZx9SHle1vQJ7u8g4PSKoziLuJOdSrFFxU2/aNtNAHJsQ+rL5Jyl/3C3OkVZ5uyc+tWvAwIdPFd
4FuF7KooeJGpEofA1joYDC97meFIP3mGC3fkyIXbqqQsCgfaEsyReMJ1MWpJYDTmMzRUiw9j0v8B
SSkmlniLsHwxzLvo1O6AIDZs7BV9I8yHr8syz0z1H5FIRNFGyMNYmnx6Lc62PNNNp9PorpjvrpIY
ojwQOPYyye7X1Wuny1JuLgKlkNQ68Ax7CPYgn2t/TUxRtqEPKf6nS2Lcb9vFzkdDrDLROQIckmpT
X4egse8CE209Wl6WnIf9ILAsIdvv7i1C32+nWp9n+v+1TxbG2+MC0CZNLJdkgNWkD6A20/vi/IWH
j6CfJPunBzUi82RfRBBUlMbFjRiCRgkmK6+uPdSCyNUk2jvCy421tCg2JUG2LF33SQXSkcyPUARv
35hJuyThlqDVNPgAvjfg3LYKa4ytL+GVN4Mnk5/imo8I4d0JSpj8V7ZDui5IdL1QfUurmq0UPs6k
q2CM+s/USomtDbU8Yy5aJQHE5BcxhwaEnYQiaVhW1nVkKlqYzhMr0p1ZpjNTv0BoPABJeUK5YHqd
iLuq24qekdu4omcNWcdwzZAfvsQVyc28VR1sz0MpU/AHR/pMdmO8gtJ6xnYgS4YGH7WmoQvyFJvo
ekcPiH5GOazq4z8tJGd4qpGAUs+usvxVE3LhZk/BAmviChWzEYbvRlUNhcw1NLqPWLS9cv8XTeHv
IgSPHdacj3FUn5nm5oLvPartlFAQA/kqz3PKGVBCsJOae2o8xqqL78QOPHf7/TVenk5w0k0lL0qB
2wqws9tpmmzMQg0M8aylfn9Hv6m3aCpdG3+GQoE3vvC4pAe1DnS3DriKy91yxBZYU6cHkeByMylY
wpDkNnyIcUZbrjSWjpqKoaCnBPgsc/NL6HmqEpOJaNu9N90wGfzLTXCxGt8sjhrtjIFnansl7FP8
uDcB8Dx8zKpU+H9yr2f5SpYGqud9gUS44qQvo6xaFc669kn02iCmnIM5VRMyiWN+bbbxMvBeoIlN
sAHT91k3qyXU3yB7aAqRlF/xMquEq95CtGfTMLbzdFAVOMrw1+A8Ew4dCKZ+yio856iru8gVJcvD
3jcpOuJro+JWoCVDGzlwVakEK3gQRHPFPQjGWgrEa2E7bdzmWHErAYip5rOrPhBP99dR7pbX+8uZ
6AUJwUfwQLF5sz8A0uc56jRXHxFPUPHhyyV/WTqGu2vJtnVPvbXGN2DBxYqVoOwcQFsKhkgnjkf5
EKKizt5RmQtjpglMGt6eMD3TBNbYHTS7QOECd4FN96dsZ7G2KB+McewhD2KZ6SQK9T+yzGTgkfGR
pJ95PttkOcy5iHNx9ByU59aiohICmPgq6SMGOQsYt1J2xtjzig/RS/q4AZZjaHglHVi0/6qdT/cC
hJmVEDVL2qa/PxAkyVX5lIm9ej6tC6uzxBtq762FBNkpywOICEG8Iflughlva0oeQLndb2mcN6sD
veWBOMSFtWeRIIrObr6acuM5m0l9cDec7tZEv8ASfktuqj/8o6OfgDo8vQ4EbjVET2vDg29P9r2+
qB7BnAtXSCKcSlZYCTEwkmmT9k3aJ5+EGbcnAInqgZ5SdIFuLUu5qqmLH66ql5Rz3FBazn23lwBb
q6hBV0AW6ksNEYlf5/3Koo0XaxvQhUSWkyWavQOELa0yaIlYujikl0zqL/wtjb1bPtR4OncjzXKt
ZFg++uwrBdjFGzYq6AiE7jE8rR5qu6qBrOFCQHuETwjR4x5uenYqXucVuM5soqPLX1MiWX4hKd05
iRhc2oq/5kQ0jq5woIT4Xxmkd9N2Jt7RMtwO34hWVAABfV2YqhmvxLQNazBaFzR1XkSZLfEGNoi+
TcnjpsZhn94lUVapZI1HRPFXu72Zk84TEQ1aC5AMH2kTs99cdrQcbXtrKY/C+2j9agbt4W50gCYZ
/Ze+F+AWtPT+spOdhpGxfJGZ8nTsWG08ktd8SxKdxcFF+WXxbatdp1FlRJ5mnbCmWtgTLqxhMvqh
D+0Umja9gD9bcJrl4gJepGeHw//2NjCZCnhpGKySC85U6bp87/P8C1v1X+jopNsETc72do7dmgoX
maghkA5QQTPUQkVKJhy087bOvObQuOn2abREYmoGP6KSIvXTCMNHSNOJja/1oOYJpSD8Fjb0v6DD
7jjZ3wMdn2K9vG1u3shk3ZzQ9gcoAj0ieqlg1gHxH2aJxOf85JosdL9HLhCvzS4dybV9VGLRbeMV
12vnVRwylMimncmQR1faKpHio8Ao0deqXSdf5WruKcNlqiZEb+o4GH8rm5Fd50Uxnpy8KvGAjh9u
j7aU0puh9Z4GtuQ3YsOs7ZEZZ1VeCeoCyb9jLT/xiUxuSxTJVH+srLBZ3seeDmViNr6MiIt3L2GM
zHrJkzUmk13jkL4H4wGlN5PlGhuiHlBz3uedzBETtJZuuBrtAsq04KZByl/NrnMUPbMrcNBz2t1k
boTqSZh5zoQlYF9VajwOF8pKKyr8W16hZxdESqkFvzgP4z1weo4MfTh5LSgYhQBOy1hxVhHZtoop
mKu/fBZFlqHNjCxVzDxpqo3j4orVGcfniQGgREOeVr29PU0CWEwAjMwL+YYGxR05pP26aqo10b8R
WbDmEnQ/aTeZdvQUX7nKLKU5o11KHBiXXsavN+56UeIagEkXofoH9kt9nBAFaRTSliVzrctgR0e8
7SuwLEshsHf6YmRfaEH6fqWUYKThjPpCGFi5zsEZbqMRC7F525UJcbGNiAsze0ZjJpBIV7fxvxKV
3BxD7jhQCyv8x871lpKgxc99DIf9/Yj9PEXRBxO2+6n5SzD1nskW2rf2RDMeR457CAKEUeGwQVor
TME7zVlH3T+xcmUeFRN1rXPQEdzb+eajaQsbGqtmrMWZhXuPPgpEtT9gNTOjClotUsodzjgF4A3m
aCby5TgtAGkG6N+bLFylqFNVpi0R+QkmclOEjugF+tN7DBNf0hVU0GAh1DaeJ8z2FyuniceaFN2q
MTO6s8JYU58ghNgmewW2YzkvMbyKPAbXcv3WAnDC03gULc22s57WVtB6aZH3cJ9CCTzaEZzv0DRH
1ocTpHim23Bvvgn5soXQifJwz8OsbcUuSKormYRRTG7/zRswaa6rEGZRh4sIiih9wDLntqJeJlD9
VKIgQy1Bpy2RNiBnzxxcp9XOfybLAimkl7eptIPuIIT1PXr8kmrfzwaA28NpoOkDwW6FBBmmDEto
vHN1oy88XZHtcQR+/B5B8jTuZ2qRJljgFUr4+kjXfQ6pNsFTSMnfU1ttQkSnXLRpuF5XoDQd16Pp
R+E7K9S2cATa7fnuJ4R+jkqUeu40xY7mSYM5KDOnEmRDdBRBcihL9hqmfE8VMgxCD7rewsHakMSW
hJFmD+C3T+nNJOzwC+KH43e/Uxej3BBOtZNaSll1xit9Zc8T4q4lvReUzAW9hPpu9EGjcxjic9/Y
kAVWZ/YQ/2YaFrLKYmyBiJoNAKNl0ZCiCmbB6hsu7yxyFcuYSu+6pFQccUh1SdlH8cm4Zo3lgGK7
f7Tar3OW1K6PcqJ/8DDuXKCZTcZY+amdVKjHRWS4HTDjSA26nOsUB6YypQx4fVD85+KuUy42pP+R
zeCEAxoaYBl4oxDG/UCR8zWBa2U/hK059PwAeIbQwy0algfujw8tM9qWBst1MdIwuhXuOsS+WyB6
PKlO4Y9YgIwJXYmT11lSgB4/WcEGmUKrPTbIlbfcs39mhZvJ+1xueK0+dOAvSjZU0lDwuIEfjeJo
H/nTPWHSjiOGbdLABRZ/Im7Bg/r/Gf8SEM9RCS1VsuvLEETfR1pwxeLHzylKupegxAvvzewdNmTr
ueaiKotAOzSjXUhDCETcthLErOz9kr6awTHuPVhT9bN/r2aO+PqPgfP7un/drzuD8wYnfqPbsuiH
NjKcP7qQurUF+kQL95tfpkx1upqOC0Tbr5lrl15aZaH/JTLuU7+xAyb/JXYk89QxQMQ9kwoRSH8r
nFHS0K7rpWkBNzViBQFquLLfk3rDE2XLULI4invWv2yn639FIZOgHGM/HSTVk/cK1CFRYFPIzGxs
s7ABhhJuuL2WXVtCGXisoz5ObZ1CkiTnSh73KYz8g2RsXU9MEA8dt9WTHGQ310ZPl4x2QmR/U8OD
E4Ni0blVA8Lot6CPy/EM/QHT9G7sUCxsJdVsmLoCSk6rbOLnSqkf5wetxWLpTlzOGkNsX2OvZBeq
YG7XEA30eqvKy0617c6Re1voDFH+G1+kHf3Tia8ax8V6pz8rvgOTWbzSv7KJzq6S3EH0E6FrLUyP
EaP9RMTseCoKnZZqh5MwXD2QQM0DpaVSnXTcn6fGJvwO1OZLWjr7pb7+riwmbs2px1MXUxr4l7ir
a9QYzw4it8N3Cve6oSn5lTBDhG93PvtdAm7v+FoqFsbRlQhgIKIWCPS8zZqPBOpKCAcPq3F5rRPn
S/kTTopoYTO+Budu4DPpStE394WqqbZZBw6W+Shjpyj249nVuFkJZu4YJwRzIx7os6HtFwt1o0J3
YdEJD7oZhFpRSfFkXwVT840SsSIKttuewcrKzf/UiQCZBdK2F4ocgkVY5zPTjd6U7YQeyrJ5dZbb
3aNnu6O7I9C0g9mbDd0fheZlzxB/mpXQeTrg1QwRfZjdYxNvT6wAHkc0pPOtqPPDtj7l1BDUNAEN
V3P2/TGVL0NYkpND1YrrikDODc/pLow+mIfWlt9ZAA/yUzwukmDqGz2+5zDgzYCdd8fn9pLPZqi4
E8yj2CA3SVAU4ERSnaOdvRXLHA08/EaQQh7B4XpH48JqygMxLUBRDLcg9uOrIgslW9+tUQ+hQaDc
SKb9tKJI3YGyN5NtNcW46gdsKN6uKw74jxD9+B8f8aSe5BOhJZSzsUazQZBSPBATHRh4ibOizh/m
T98m5HKk7VbExgnmKZ+WEuA23iNnoj0yehwaBku8zKHk5hPsc1t6gvDfTEF5d93pQ4KAknLcUxoC
yBbBtg15/7taMZeH5glhhKy/YXs/5cV4d7FY+0vGO3IKHv24/SNxuAuLsqRM3CHQyeEANiv4t/Gu
oaNC8KmsxeYG1eTifsIYuBMbt+C8xP7ErSN/NcfC6YGkQ8Cv0CtVGu7SPE3HYh7Yx31cekJbe622
5IXIzlYAYxbhugRLwNwrbLEds2yhl1prMv1iKKRrt4Kn7pakuoa594/HnGIgHB0u/Wlo33Qnr/SI
ycnj+Wwy+bj2TYUvR7SCvFIpzHvCToj9MJ/f6iTXJZALxWvzSl6O3xdt1le0HR2jdHb2W+eoR3Rg
t8Zem98vufabgnd0Bs2enpYqnTO3lEoGcdHNvmAUmgMvPTs/o0NtsMNuwTCluuSHm9GzxOvcAalZ
4IqZF21pVpGCjHG29U1rR3ntxXPgeRawuMsvXdXFYuxe5ofJ8MEGPmsUDIW0JGmAjGtp6iVDr1+T
Hw0X7SLNSiwmQtlR0Ggq9jBxT3/yEo5fmB3SbkKlTybm9D8BCeUNdj+WoE2EfGxG5aYE0PIwU+ax
R+R4NYhjV+AiN3+9Jo7IFomSmzkoQ23HXJka9ggyKsqkZ9XF4Kc0HTvaeSijkyRx7qGIVRl+xNS8
2cHZydALjC7vYhmhKwbkDziN71v/jodr/+XifB3adkycdeStJnuhWSsxO5mwEWq2RrGsaO9GqAHS
UzbPQatlEGFDIgYzwNNu+kJ7g17tXfifQ3hL6ERoXBArmYyLO3daMN7Jb1jrmwa/tgVSL31uICJa
VCuuRPR8RTrelqmgRs67nIemrc5jhTeRGsF9QV/0YPwCzzt6eSVIPc0dsEwAXij15kDSW917pssd
FD3Cezf8UELk32/r3ZI9hJAh6eCajEU9OhTFWr5/HYKPkNxUriojE0k7Ptc1pBRQm0krWWDLH+V+
PvX+s8MjAq5ftrYNcHLuiDURnD0+8k4/kcPwsxP9LHj0RDpmRVGfEUQ04U1MhQy33HGTEod+Rf05
kpaRvBs+x1qP1U3FK6ADSnaN5YpQjwAkNhRzp6zqkAwQrTC2mr4yVnd3ekxxmzE0AgEIq6RPVEj8
yAOcHtryD31tVcrlOfJCP4IL0PsV7T1uSHnN0gw6H0hNrRC88MK5l1gMW3Jf7SwfB+MoEtRdLQLk
0JKUAFhqDnEk5mDbsIxU2NO6CQC71TG//qmiDwFomkE3ex2aYFuAdpRB1ICQmr6xstftKCvz71d3
0+3lwO6FOQppl8RD7HnK63Wf+x8u8RpzC9i3cJPC5Q9XxA6uQAGco95tKKL/dUlhogaRWMK4vSKJ
v1fLh88iFMP2qKE7oN9XCBuU5xxHQdb80h0NFL64ALztv/DBWhzw1poCHosKQpUJGW7He0ABfOVO
O8sDb7zuR/Ug8l1AfeuvlFyRnRBRZeo1uj8nRTBvBpaXw6cLzOVsEHJzeGWu/TtFYnjNjhpxjvyX
PcZPGigLgBZx/A851eCcgy9CCQbmyn+GzHC12pPPAzWCrjFRW5/eA5ZIGz9VKGXGkHjmIRz8H0W1
Yhdo55JCSAngYQ80RuEEgnPSj9DV8qSFqdLn6AfsQOePi8QjVv0UuQJAYPy9rSPIRpcZNGfa0mKa
H7QVRp4GxR6ZSCVsMzWT5P4MehzA9W+xMMMhbcFRWNva4/IZTs5KuZBqGB8HkEND/uqasg+/yTrk
s84Re+Pvbb103Z7QlgjhipdOl/hdmIt6YNe+YEq9EDM+K305TZAqepSzYgkcVYGVO1YRRxaFv1Ww
2gK4gtgtTyfXe7VD5aCyYrhmgahEsjj4pL53EL5/F+K5JAPN/wcVHL+Z738ZlTfSlDEEChSHsxCL
5Snbh5hEHZmZFXUmph51euqPDn9WKLMD67EUK9gkbY0L15CZ7FkQd7VBF4kgq6uqXGmlgE3WhOJC
PfCzge6bGqBhfeBuUz234BQrpLiPlsI1MvfTSiPDhPTacrowqYECuZsYDU3d0nyWObyix3ZFf/S8
D7YWiQQVs3nzsi0ghndyOFqBV/rU/fLTZeJkoWIzrPDT2A4q0W7AePnp+GkR5u6gctKFYD1TrzY0
3z6ILi0zwX35vlxz0k24ZR/Z+d6OL/oPmAwcfYAN1DPW8Eh3n4emhn9m+pYoc6TU2bRUWTe+R863
125b3pHEfrjjsgKqYEtDd3GhWPozShOQbqVfU4QwUOU6AbuKkx3rWTJW695oUwFXGUo4mSSZ4GSY
sLq6qzUgoYvrDbf0ARdhxGLPN02nK6dees2Wmsa1jRlPq2U1NSs1vMoOiFec4X81ZlqH5fxpzsoZ
ctYyTKbRLejm3SeLr43s8o3ywveJ7HqpKoGqUo07f7OdSgod9fKY1UaimBt3l/M6f4BS+ab05U/X
TcBHd79fgPEe9y8yglUDU9Gyq5N1uAx6vdU85tpSsptJuvVNUcZp2lWZWW3NIqf9SpPHTKsjVyBf
zI/eIzdA4GPGayZKkNwiCakwvv9YaYn2FA7jgNJmxYnIToqFMvDrJKABb68M4qvwL3j0NDd0CKD5
a8hxJqmcLqdgnAUr4fnTMZkw7dEB/9ZVE4oZWWuROqar/heeWllCFxuCjdW47uduRoZAfD5xxmbh
pm6GOf9M4MQDJ0sEpXij7U5fYzC8ukOG0gej2pGvCnZxCAXgUdVAYDh8UNtuLtCNSihHi3l2LH/9
fyhf6qtPyJjb1e8zxVyIHPIb9HIc1deVL/o9myvcnalpMMsXT8V4dg2ypqWEPJBLplb/L1nARQdK
ZtVle9eyJ8CPGghA96qwZoyr3Xlqp+TH8b+eWm4R/bXEr2GBKYebbQT/6ngzLJrio3mC7ccNj8++
Ic4JcML67ZdF9wrgmhf5Ne6wI0TUxI5TCXQYQTTWFbe4wvaooA4fhpRjA7HgMXDjuNK5QXz1RDod
hkTEqodImOCwYElvWQsQZBq5KAHe4q4QAWBzhNyBMa111nvCmJxauUaFRGPGn/l7TeK+pfd6q4X0
Rezimok8qiIhf0jF/GoR/Dlgp0FYwhABtbK3KLEYBGrco77xrVUoQrp4P51VAelEZTNdrItez2Ax
E3ep6GuMe5pZCfcPbh2GBOHpI5dZmd2egC91Q9kI37EZ/+IXPHwpNMW+d53b5snq6+ePSYsdbgMv
Kf8D5w7nQ97BF/l9XY2U9eWr+iO48V4jSA4bthR9p2gQzR2Tdif7Xr0GBRH5D8kf3p1CJrAhykU6
Uhfwf6g8XhfRlb3Qe7dLJ0V1elp5IPBgGC+c7DMKkNPMl+aVIxLy0eFiFOXlAz8dNydLcNJdbsxX
u1OV9+vuxfQLUkRknI2LrLQaDeANnijNTFMoMSTUZycCCJieX4mHWJQ3b3mnCLkdp/2IHqnVcxE1
bjyX1fIZES3bq4sy/8HeNwwpMLoE/0qnofU7qLPGMSfEOD4JRCksehRT0AWj8m43LLc5XxQAQ56c
3yWQpKdW8kxNPYrWzfcRFwDIhruaHDWmBRrVWor54WT0aHwwDUynzBJK9dAnbSFHVQMH3P00eDpK
vHhmKDqpdhFNqlsbqOFnXDzAn6o5Upf+VjOzzmErqTirjZuus67+EZWIiapM9QVz9FgGcSalulOu
44n1PbY4f0Sf48PdGSWZmz+2MXp5R4RlalY9Y2htWZ6xsa4oeFyMi7PsZ6In71pSKV0ABwFZzd91
0zOG15HmOSulv7yFxg5FP/sMFZc4DCI/bhSuVTEauZgP/HbhYYZHA1fWlCgm8Q0JPYu9OmhbhbHg
e6rSRfuWIaqhN7fHMtQNRgXPb/FgI/znedIJmUj7NVp0wJjK59YSVJB7702ur+pSI71bKRJLFL/T
7EcOdsUztj7pX/RmXaeRV8MczHqZoxO/jIWs7RRc6zIoANGLZ9L95n8CTIY90yNhyA0J4F8y2KhH
gnNNMRkGs03h4EehlkVWiG0iOAEOuDTk3efaVxACLJWIAn3qFxM/ms5uDyyjtA9Wvk5B6ePcKehs
LTYYEKFN8iiwXVJM/mYNSr4DnAwQHZGijWSUGXJPKuRlu1vsRtRNL2JyNTkVKvMgHwHylUPt3eRF
boE68EgGtxHgDe0ZYS6aRlgw5m5tnJB0+zTBrn/L+4hDPpTGUXywEklBiHiTkISLLGkLbCoyawK4
hsv6oqYNauvXpDm2pqvVxRXVQkd76rwNhQp0C/ZUl9SVPrEd3agF0zvnYT2JYy1C0tCKd8220ORZ
mBwd0BpORdMcmXRIezPHt+fioqCY+Iyruw+ZNSUkYrTS+9sCS7crOYHodN/64wYOIbhd+MOYkENG
QkakhTogMMwiGQ4f0/wCw6A/X3FMP2GbFnjlTig49jlvia+vq70kmoUicV+L7+xxRTmtkQFYA0D9
POeQlbNvqPdwupUIgduUWa5w3g2Ncjp6zuANi6NFMSdT08EhqAaNTTw7XeYoK0zdRqigfhzm/LaY
9uaU81Yu3Qp5usH83oHLHkac67W1x7Mg9xgifB447RCJxcMF5pqAqp7XKQN5d6SdUNU+luhu6OIF
D41si5mTeDzvnlUia6Qvs5Yiu7fpTPQW/bGg6s3WpWPaaGWRk8ekE7ELWBLHJWhy0EKTbnjS54bH
ANaLqE2kdi9dk7odebtOBcHFHsuR2eMH7jQpvxrN76+1l4M/KIK/f8yDTE7plw9ijbi1XoUuMfC/
9HL7z0F23IszluXA5ascS2k504bnrTc/ZdCnsqiB8CRM2uwvDFcJ4soD5zOW4ktM2BDgERIU5uGv
vNrKa3u+zntTdW2T0eZr28FufHzu6WhIdy6GTKmY2ACLYYEmFrfdjTI/om+x7hwkKPybWcm2XFt7
UuHtEYLBeHBTCuy/UsYvSwrsnhfT5ic06fzHQsOtEq8y0/l0gO9+1n3iMIDhmENw2XL3PL+PpSyz
R57Ct4n3grdaafFRuXUm74FEv0PSwddI5cNhvs7Q/YdPbK8YGWJWhGv0MC4eOifqbG9MA9rZnhic
aNC0j3fVUq0XSFdsiHS4XZE9n8aSpuPV5fLPpSkf3g+qO+72yeqJ4UIqICY9hYsGTjfEr2miei0L
nxle7QBOpqdf9zrtS6wDjmRtAcotc8LIiHTg1eBDXj29jQQHtdKJubqZZKX+k8ltkmvvpb8kPLPL
3K3GUR3jko/9PVcqIFCOcOPyfW/m+ft4UMWG5+j3jfKEBixp9ayMUzmgVzHdNq42JL/ILQS/QD/Y
tXZFNdPit/hLVxxdTE7TtFl6LtovtR67GmOSl76GhNxJqYxhF2HluP/N78vUpCL7vdM5YbWYiksG
6FOilUc1jWSf2u1HD7Cb3/h17mnQpAGdesRlEhp3PwtnDCHe09vw05ieuGzu8bN73abgwxOu6o07
ii8pXpg0TjUU3YnGvjftEud45XfSOud7A3uYRGZYIBkWCGuP3yZHJZ+Cz6kiZNMNeLN9AuDEie89
fMPZYousvYf6LpunVEpvZ77rTpISDK8f1XKpSpYlutESRGz2goDqluMc+ca5UvBtQoj4rEDJIiOy
atZSIFZZupdhjq0a4A/BJb1whWnPWXIdEhbHJRtUpl4dVPLOAfwu6sP1n/lYGFdF4eVeeiwvv4+X
4XOMJL18SOnyCsJ7KQj+LHiKXgYLXbGeXZU6eQzzR77YbN3+WUdz5OKOTF0rwWItufbIxRvkC9+1
CeEyJAZco+NbnIHoZKy5NJP6BXVg9M8LsT5O0LzxuBe1Dd0bOOd5kCoDlrVr6Rt8qbH8fqMhSlf1
Oaar99F9gXWG6dkHgtOdIL20UfEekciQZQHDFVq2IhmhdhudW4YZqLKU4fZEeM4YYz1hP65yt0GS
6p2A+PI+IVj5bbBEbmMTfGISkltmdKO6sagb3x+H7GqjPvWjDZuukq5h5NawiAuOQjKNqtgLGmeu
NbH9IGjVWl8p00bSLB/3gf907PuqObCvQFMiN9lQsc4kwvazqgyYU6FhQvQY2as1PZ967fKjgNR1
4yBKjOX5mgRXO+IpLjC1UK27lNjy11Ic8zMnyy5sTLU2LVay0iOAskBcODav1pNKYfluCMKDh74f
kU47TJDEbhzswk3oPl5oxVtX+3j+5REBEnTdusnhKk2R9of0q+XrmpxEynr9Ehuc77F7DsnxdD2K
Z4d4sTEVv430sJ/6VSBPiqrdXU/6GPViD9KDp15zA5tEUBpEiKte6oo3PxG9QuA0df65BgLXWjer
3ZBf50kfA1X9Cu0Em4zgVf2vmJfpDD89vuJlwXfgN3M1dkDKqkKdPqdxXqx5dewHLi61JyR/ydJp
lj8/1ptIaqYnxmg48QLZ6QOtTFd7t5C96fKIALn1twsa1WE0E7LqHw3bcIk/mLWQq6UEYM+XROYm
63/pH3ZiozLjqNTkvm0aakjdveK+D1GCO8PCb8GqXzsxGrKLyYVQSmtyfeBqYVDWQEQAMwN6Fdsl
z3wgj/6aMgwG7k5sjx6gpTUAM3QQEFLxt1tRZtuIROOV/p5N5ORk7HVvStdB/iCAjB8T0bO5eCt9
2IRJNhoVaFq4fTr/mS1zs3IEg4YBYY23IypFS9o0MRNBM5EAX/hJsniCNTXxK1usIeSuqsa6fes1
pfJpuizsFmgT3cIls2qrbZEPfniI9HAfNssANkI0lx+BVo+2j0GxddcfvcCRyarZfxs9hNAJSUZk
sE32d6nzh69W09Rk6e9Hr696+KnDpVcnu7SkBHCvN+wSF68cC9LH+MqpbggGsoDbyskWZYNooevC
BuzZem+pvyYLEuaQtMWeUMQqU0MEwb6oHyaN0Qd9ayno7UtYe9sD5vU/rA6PkRZJ9wQ7w2IpvI80
2mB/MhxqEBlx3mP2J/hYTMrsK/JPFpat43aBxtbUZgaeUIAA3WDUhZAFB/L9985VTh7dDesgNFqR
exz0SE8QQhvmiMRWxwkhRYOfvTbGbIIink23b7dsXoNaD3cVAyupaOaMZa5cDyDxNLpzQnXYRLtc
Q/znfOWPdDHFp85ku8Ypfc/0KQbyeazM+XUofY8DKLX57tFZb8amIhJLittXRUbqi3+sESi31LBL
tM+LL7SVZDaWiBvmn0ks4XDT7EeKgnoaQ64xfJgodfxTWnrX0tjOjuiar/YViARyRA7xCQ8CZkNj
Axa8M8Inxtl740fklnt1cO99vLg1A1EBHL2xkLiSSGsJ0/MLThiw8tESocJyALghxorIlJwZDTvF
InaP4rmqVh6UwnoTyyZiGzWPwIxeMaCrlN2oZpWZ+JDFFoD/urY6dL8MKqs+Wi6dgsr+whvp0ys/
/LX5435IihJb8Y27l+ZqA4lw8YLQNQEe0SiqNpvefiTrEmepN3Q/Xcs3TjO3Umkid6OY5n+FXVxV
K02ZXv+ZK6a5TVHRmTVYykhPqMZ3lrDKBIdC4iDPsxVJnLFmsEQbiZ9u5KX0VbGM/aZPabt+YlHw
7T+T+uusZy4KEjIAszQiHvmDNBjNasti/w3QDp+u2h9MKum6mF6NEoCtG1YlFNaJzq3tXKV3SWYd
zFoBknPSN5TNDOyppy+X+1FLEHINTjhJKX1IcuDsEUqNNiHwdUgNRrigBdG6SEaKJuMuQvvsVmMM
tivxrIS7wKj2Qc0pvoff3Z7vX6OE8JSvkJC0PQ7aVBw1yrJHphDNOj0fjPQgSj/07jCowaZSXXDg
aDbEjxXLkn5Qi5vWJ9o382NBsHHcEi4ybh+x8Zw2epqIPKItNocIOfc39vcwc1U9o8PPhuDKQEwN
ouNFLSXIxGLW/ONO74Ai7ChjYxv9J5TqSOn0RymZ/Vo7el0XWrfgMIrcxLgCJf+NwXybp6uctUbP
LY5iJMIChrCOn2n+SeUb35tt4uO8GVnbTTWCo5edfYIpzzTkuXzKbSWCJXVKpngFPrQNVhYLs/Tt
IN9ctv1brSJd5Ru6pEHzsKTxLKMj9aXgQu1WoQLRizfvFNV73aCGRTmK3WN8JwEzr5DDta2TS2mO
7K3WPWdfkVsZPXiyMwbWvNaF3g5KqFKePOVD6m5f+Zt2lF5QcGB50Yo1YFN1yRIsJmuwq8/bGgTE
M5eGNJXvzkMJx3yLxFF4jdnJnPtIk/Dj0rTDKgUiVDiU7B0llRY0R8Mxgp4FbyScFIinasODnQaY
UUlh+2oaZmSIaHY12aRRG9oemrV+8pDi7uTy+PS9A6/auy2oPwy8aPxPYb5p7QfEQ/YlAi/a9fTT
xaWy/PxOSkB6PFrZeWFba1DzpZHmBcP8Qx6VPkAYD8EECqdoMDF6n7dpTk7AFlTd/9Rk5VCOI+Hm
6FYApWb6Vdfn6o6L4h6SixOKe6vOx+9vCF25W2WiQY1LlcuTSQhDQ/Q3cdk4MxRGo8XcLG5D/JeT
G64jjIpLTZLzQ5qEl7AaNaLMoKhLUJKHqNW6gVAdc5/wnkdvq9lZjocdpMXf9iCo5FJP34bfYia1
gZm/2fCKlYRQ9c6Vvek5pUw3lqxLahfiT+ZQRbDrE2mEvkttX9X9KXXKv7dHWpA0z5vsVEr672cu
T9D1mTJzBdB9My1qLnfg/KdSYoAOCLr7gEaZ5JZd9GA8OMFVomnXv+NdAaTgZyNWNEbZ+mJnNSCF
ZRHCjMIlkN3wIuzF6IewsA22uZXiGPQm/Aq0aspYvz6w9aYuAgMjGN2TxONXOdMY2rKQB+5rBfi5
W5caa4clpsQeRGkHWiMSjmtUPYq75g0VgmhfEelmeErTIZXUUmpi6S7uZd1nZjQL0PqNfJneuLPJ
OZMDwXxOcqFhQ50PGallF4MsWS3x2Lsds+kwreB1ojXIB2dlFKBlhqOjhzYGnKpLggGxI3fnWZzh
BnhfUDKLBKA4FqeYbsDwe5WRVI6tENFch4kYjVyDSPUHB622xh1h7lokRIByPlNPD6VaDHAFjbTN
HEccjMhf8laAOBvX1lGRHSlxEBgzxXUogdNzidUgeNnIuW/hqEmdSesQxdleeXFcbWcTPOVgcvZw
IrgY7lwpauRn5ZVisKI+/XYnqYt/TR/91c5Y08Y2pV0YwBqYLxKX9Sc2HXQi/hF0SD7W8jMIZ7QZ
MvKxrPxwyUOQ4fcotLImAWqiCdspu9IM6T2Z5F5StZJypVwF+YWtTluciXnnQVlZbHYo4ezhieuW
lx8V+OkFOM8tUWy2ZMClM48/ntM7ChG3kmqXJIiIHaoyYb7XirkA2Qd+tkpPbW/bqPZ/1gGwSnwy
Nfsu2ADRGPyFe/3AMp0IaXXDX/KhLjY42kOr73wWv5GUInHpu8JMeQSsXdVs8bhUYU4xq8IwaQo+
K4whmOL7a2MkE/uW7lX53HGh/M6ZAblmCntvMP1QeOi9g2deN3Vm9UWD30aRZj/2bn6zTMMuH00w
2d6a2MLvTHtdnM3fJXXBCm9i0g+6aS+0VN3X3yT8F3wbyaUYmNqbEKfwKdYEy+6Qm93q4BgbHzu/
K+ZzEB+zcBPwfGQLhdE1VYeXNhvVjUW5EoXQsLgkKgkFXfxxJJtCPJ8+rFaWVJ6kGV7wm+m3cRFy
87XUSYo6kYn8CelZHADumndtJcbcra2iCXJDfIrCZ0zzyjcQki18W4oivTCtjmlaFRnBDq/yotRb
nxHzpetDyFMzaHRubtWlJi/pPdB2Ppia2Aqc0VteW8EAsDfLRHYSvb9A8A+MSt/McuyDsU3FnsL5
4rE50eiHUcwK1mlExZyKhkawsFrbOPyeA0x+ARHdNZf2WPfYlD+rlAna6uA5x6NADh+ZWqMgy+l1
9j9UKYW2SwWYgX4qTI7uOO6pMLqNva2FdbArEvn2PnXAKn/lDxLbO9nzaafvrLaXzMJn0TzaukSq
BnoE5Hg5dxyHszdi4qmQhtsMGFzBgacFpxCWMNTSiXfvbd4owblTser5ydhcmZKvRxi+N5KtvofG
z4jz6njtiXov+0wZEaQZGE01a+1HnN8cezJh7OeOBVCo6+DDWxAWLU8K+/1ro51EvShVjD7bVnFi
RNwHuE8I7NSBlIMsF6ELn2AqgQYQeQis57MnT0dovYxSmWy6FrynVUpB5rZ23D4EURIsPQtVRhA9
vNgFgtPMtYZhxvPld4zqX8Ir5IRkI3YDgiiWdH3oM/JrcHA+1VQOfZnnbPQIGK8ipHw4QhQjbYTE
HdfV3sWofDOAjmherFzfKkxkRderY1S6CHNyPsSuG8ema2uiUzdt3lp1LTux6y2LuNkGAiNNTWbq
LEXC6IOW654dp55RKF7LJkgMrUvRvGOGLE1s9N0pe4gvJIRbp2Abw4MbFCPng9PU1KUGCrUctRaf
iHh5X3MZDbTkZuCQBezce75W8ypPoV2kvkb28cz/tzg91FJt/cXafCkYVG6mRbsRXc/BIjZcXc7V
IVDDPqapoDk0stBU/bI4hwzssFHUUaJaFLW+ny42pdskgPyRPBsZc651zhnfE8GjeJU7JzmZ40V1
0DMes+dABL1niHh2JUNkdFj8CTLaOPFtd8qeBdrNo9lxxpvzveJ0LJUdfD1n7ZYkRHTFfkbctMy6
yDfE6A5XHkQE3VhEthTa6TvYJ5TIMBiodYx6epYtYrkaF+WDTRmnAQ3613qMpAz36ArjA7B8+ib+
BoPYwNiIay/QUEocOvhK2TAdWHCbsqOj+QhyYcdf4a1NmQ2qGrbI5eCaziov4SjyOYBuRtukk0qb
38F7t5jAuugS0iaEjg9bG5N/vfqGOgCAjnuzqCZBakUyKyijQGFr1SJNw7ggTaUzIBELVue7U+eK
6kpWOgWKys8t0twZUgEEUxKomlJrKIths0N+dIUwOb7k+9Fbx7P+pvf7aETT0SvNBKDTIdDIS6Tt
aiUFLWnYcKcs2stbm7cnR0MIcJdWslz1Y45nt4WVXcOesxEaxdltOKtmkMQ5q0LlMz7FjHPjoddH
sca4nOPgwXinFFfuOCXsenkRTcfg6ndOhBHkqv3OzrnRDi3P0WtssGM58uY9Jy8qei7pgoiDLFWV
J3ew/Q2/ikDhNATlh93XSYw4shIXySaiyWXtkvNfUPAZ8Y080zszxbOu4Rcd9K0PtoJ6BuX/LFK3
g3roQvFStDLQyjZgPrWu1EYXzw/2yhmaB7n57OFtz3mkEW6JD96X2rDYD/zoME4YSecmkpLqaZET
+GewPint9Dll6GLCvM7OgwDaX0nwZ1dtIm65eouW2dpsaH19wyA2ZOjcU0J0tnpV15aI6iDiZcP8
MgSybgF6rwaeNFG19K4IcWO8h1pYyXBFp64X1rHoShZtL9i9LN0tw7UwBx7+yUIBpSsxr5IBfXri
v49Y7a6lPymSThoJgCm+EjZ+rU3JDRrLsuwSaP81yhTpUEdrwKZqqJkLA2JdxvJv+3vqS8R0Wf0I
nEfkmYCTOItWdNBJrU8kKY4hPmt4f/hRJxysLSDyWfzzA7/uTIjEaAmtjp8e8sKu/LnVH2ZZBPDp
RwqbkuOuR3z6qjfHRdGXSa08srJ1/5nivq+J5b2H/061WAtWm7PoG21CTV6FvvRzdPqedHobXGC7
LZhfb3Fl3HgrEi/+EXyQtlqagOD8XR6TESmAqbyOh5193OP2zoDQ9WwR/EBg6tseeX5YB3vRdi6W
dEkiKqIJh7PCFqT78znLeyHdeI5GT+lxiX7Yuyb4o60MBEkUvtXWfJjeOHX7bBLh3EY5yI5nackI
53Ipjg309bkroIr12HfYAf4rgh7XqFjyM2m/5OL0LeNCrmrAKmzNuM3rivWawN/FbQo+0B0YoyGX
WELJhoPGtmeLU9ezyqYcY1h0MFVbE47ANzMKLgR1FfQnCHItC9wCvy1JHGUEPbuiUddy/8wykkW2
Lc8eVB8zUNjf+skOag/Rl+kZaJAUznAftjXAwyichGzb81oz7NoLbgCDB6N2SLdYT5YohK500HRH
fM5M3Mvyzph4s3dAiZhYWV5CmhTf0rKpuK9eVfXg40uGvfFM1ujxLRaQPNZZCY+1Zg0KxfkQm8sy
C9zRxscmAxQWzssYrPDh8bfnqm1YOwsfSJz2RySybw1qV5V4XhyY4a1vFp5WoqagC5UHJDjr7wrc
ZJkh71GBL0HZ0gHXuctErX2SB2pYJUZKsz1Wp37MPAirBoUzaHVbSJ4hql+CnejES8ngFbFC1877
e6GMLf62aMg/o8lev0AMny3mBBkDRyu3NLk7ytwxxxl+RADk5OYe/C3pQVrZerT7e7CyWEtI4Cfc
BzlQura/NQ49d8GGjm6JaSvpR4VWHUidbpoUk6JFnzbCQhp6uf4E0fqqTvsejAe8ukxNU+kdUewP
nKgf9F4Fw9Chfoe9lXFd7pOoydjMALMECCy3+IiPyVd9Zv4NkVSA0owCbviTkuSHwHYAhPHWtD/0
kUpwqHWBH47FXB7Naf4SGQ0jb9lg1n5+LRso6kaW0hNUzyT7ARYFGjYADbT/ZteTiJUoHbEGhS20
hR6jdLtJO8gG3U+T8wrxYOxDWvnkA8olV7Io1Nnzx/FyKQr6gCsf2ChRCDNmqvqRvN11cYh5mYS8
Q4aqGLEC282D+YVgHLtR1ImNKEHl/pffRwSPwGAX3XDDN9xr9oAR9LdFrLs/uuHYC4Ae8P7jgNLp
9Vpm0IvuLOjRqrQDCnF7aLW4KFBe/cmm6Ug4MnljkIeqJf6StQctG0A6Ym8EposD+KpPibfajy9F
G0TdLjL1d2cYQMaCdXZA0fV6kSBv/G2ClxMDG+1q3PoQUrybDc5DneVxEZNOrLYFS2urg30MFO8z
o0LF5m7DcGIdga55DWDk5oBeWTs7gTNM4NBiQbDZypYVaAT9hq/pPrsoSYzBgRBi2bFLYkroksQ2
iFCxg997oUxsax1rHdqRcwKIurVjxE0WmznBCjGJd4Xcq7WB5/GklzTPWjLH5mzE8lpQa2/evX4S
7sDBA5ezLEIbfnmLD2HbBkLf5nqcjFX+3lH3u11bwcpLxZDjshAby/7bf3w/Z8r9RIVDaCdBuWJ/
RzChDJOYUIGGQcJCAkJuap1lUXCeWNfKZMTSe4EIn5ktwJCi6niJr7RbNcMgjNt6PP6BPcYV9wV1
35iy3WyJd3HV6Xj+C1HZTdkh34TWGTpYKqiL+55ppXPQyTnLJWxBYRQvsqK+cUqr7oGE3PdN+bUW
w/oO/fCx4J+uF/tCAHOQQR6f2qEUPMs2Oc97zMOmHuupwbMNMxN7u+jJafc/vObSatzDC6sA1FgX
4O+q9epF/BhuSJbB2zl7MEc038RdOWiqv79l+zSETn4pAY7DijSl3YhcUy5tMBI75b5pisOR+0Tg
+t5EjDT0oPnxrG80Ac8MC2FwesxRE/OXSAYOIYCaYb659qg8TbdLa3P4yYDF95OU/5dsMo49/NVv
i+yl90ICbd5KKOVT87vS1ksFYNmaWF0PY7XQouiW0ZerWKmAxDFZsx01MSiH53znFVVbv++stAcl
K1lRpq3AzDbAgqepsWLL2vy7d5qUwhyWPP9HOYDG/lBBiconzrqs3U35eoUbs6DLc/FYiWOBi8kV
oiCnnB1ce9G1xIg7HuXIDRXo28WWM+zjwp0JfGdvY1iAc0Ws8YZtmeWhtJSMtUR1B5Lzhxtsa8OT
GAt5S61KkmqZzWc1mliY+VBsUJzZOgn4bLm0RLNW5IZJLJZP/45Clqk0GbInb7p0MawAnC5s7c74
rBZPpduf8XZgGBol08N1Z968V0pS0Ey3cyxH08jHAUl2jXfc4OY5Yurf2jk9NVzpN+SwKfy+Ae2z
U7kozd65GuOhM/f6LnxnGrB1Y7uHWWHkWDyICEk4/tkkffKR/Iq0ZTRPk29kMN0I2mGIITvN3/n3
cJqdyOsy5oZXxDacQSiW++/q3GZN771T1LQaMuakwCGfQeZL5XqHTVdmUiVR4uIY1yQvKe+vCmPp
yv/KrthzD7zn0U8ak1WxpWKIQMNqfG2JUrZwTIbfhGrX4Y6KV1zeGcw/flH8zh4tdvpS3klEKHme
7VKiWLxkNWesqUWmimoEcj4fgre/XzOGVXUgb3LkmeZrFMEu3Y+dpRVTYJ7PnGs2JJHH//SwZVUn
oNipGoBwWuQ7Hs5Mg7NZFGsNZCH7bV5lkkytB8dmyrcEonUty3h6SkwXagBRtUN3VAl2WP1N2ggX
UVYtnUzgNNEwlXWaYB8X2BSCVM3fkRKuXRH/tCQEckwdgWNZYrpbaJdmPunxfJh8EETwuPSsPHgb
EzDWFnRMxo+Cd/xRmc1xJzv2BdYDV+spFtBMASL8yJQE4hfOtja6D2KENtWe5VE42Ccxfwtg5ehJ
lo3i3WE1WnuejslDjYn7aw2VmnvMZ+qFVw1X02dPuW6Oqe5J7NNwSFNTuo2JH3oQB6tn+9CnLPro
MMgAb3QwdZ0f5Z1nEVRaNG6IBHfHp1xlE2A67s82MM/zevNCPjuSEfqnpZU2oNWLsBEZ3OlSdxRb
qppGpLM5PQf/Gx3vNLs34CLc1J1e4o98HJ9hHrcdpQCxL2KtX42XliggK42JncpyIYh8r+ihPj6p
ntZQ6d1wDjyZslxmfoWi6bmFj/DxS6uhSweWfylgp80/SXmhIcJsAsbdwL5TxnKQMAL0aFm5VKu1
6AecrPzFZWAKypMJMkeO0M954khky5Qlf6MvzfdrALRwS+/nGjrd/dbYqQy+RqmVn2AWS+sdb17J
8t7RAQqtwhC7Tpm5ybs6FCg1oBaY+QEhkfnG/w8QovalQ4c8kIplPBOGhihug3BpMucJXHtb8x3r
lgh5WhEObJ9WQqK64RBJdiWF/TN+7GPy+VNIdc+AmhLmQJybYXR+GuP5a5mlELxI4yYfNBsQ76Vv
epCpjOZ9Kj0YvZPVUqM+aEw8IL6E1ZJjnns4PZsTR7SJ0hIIyzewH5JJf0FJFDR+XXgQQei7I2IQ
2/q0HwNIr8LzTpNPo95Jfio8JWJgLg3hAJ0lqYSMkELLaCouE28z/fQJX73ggDmO0JV6QE2QEk+0
AnprBeVRC70N7lptYoVsqCIgdgRLNlH4OIX3uiYQMz5aWAwiyu6EmaU87I05blYZk/LJci5LEGbt
R2HXlrDMfFGB3BKZisHHqsl8/bCluodWN2IDuSF9TCR/S9HpM9FZ9SIGVPtVUfQb89razBKhgYw+
rdTO+VgodoNpQ7Rv3YNLvrkvhN6EZPuOKAS0mIZ3ZbySJbIiuOBx+PgnvfP/yCxVT3UvWpSAFkoa
qLIAZwSU663CX3husnWc/ElV8Lv0/nqtcOPEuTGnXO59IVLJ+XyrFtQFybM5zxiHH7AsapLDITf8
s9oY3QowfYVSuhJjtjljE+1dNmOLMSW2aSh9Q3rDVrwZ3bv2Z2oUcanqnI1DIHIIgqoOehVQJgR+
7m6MIcjfuCOrOW81ySi6d9H1pwGP08vCp2+ge862e8Df7KEaxu3LnexOiVffUEkCsHsGVDGy/57M
dEQXnr3lVSG7HP3/ABXl9N8YbGEu2XEZww6euiMapYkjFRb3ntnhuwh+FT3EamdBriJgRKC/u76P
sEUzTunx1T5jWTWtXMpXGCQDP8JhSB+t+6/QZdEn3U1gOtjy2nS9powvGVJBVZ4wV+zYsNA3Xq+P
BCW+Z5IziqTFGUv4K/2kqi+xXvCnKrifMs00WCsg/fZtseHQRkD9Wh4V4JO5BpwWBKdDrGiZqwxI
76iLAu5spkdWecd5ExgZepwijwFb00arzOUzaKxnHfQKscqNFj6kd4Rl6tY+7wl3oz0K166XgDEv
6XfjK9Zn23siODV5JSPEGhLQyq4M+zsBjfIRc3RXlfrMWQzjZ/Hu3wq9wdMQ3ZarYpvMaY0HAxH0
FgkuN3c8CLpLrd6hCD77p7fntbdjK4Xx6pbqqzP2Nfy9rQL1g2iyXed2PqY8l2x8Ac01mkncMaNY
chTYBo2ZBNdbYWMp94AN7z11qVOhwPlv4pLqYxRRp0ykAxoeVHmiI0rytbaU+KaofU07YUoB7Q9j
/yOzCHeQiPNMvyOL+rvT42fOSnDJDEiOTdQvQ+DeWS/WeEmsBv1xhSg42GDTm6b50ST0WxYeJKAe
CJT/Hl2Au//sol2fO6EaMyKrvdWi0coJWN+hTSVg1Ux5CMxGaTP4Jh6cvIw2HFrdVI8EtXg0LWqd
3FBQGUrAIDGmV4EAW+cgloHQgzS8hjH7jBYv09NJKVyV0E/vf5+a9YEsi3Lpds5zNSIuHUl3EpDp
zUEfmlyAqgLnFGMvWDS87vwFF2XZJaWrI2mlqz/g2RFRbwvEGgFHx0/nnaXHTqoxJXDnunyqMGKG
7EHOrpdtQJxBHg5HnNt1yEEA1hjpaFC+TILlMATu+jLyGEwHni899jkKP4PCqLWRPFoEDMumU8/1
8ZvP/S4qJNZCPAzg0wHL44t45bsO7qhGq3n5mMl1zBD5BLWpiy+wev6bLUzzcR0oqHsMx3JzDhqf
GJM3ijS8DK6V2rNXCyxyVLVMwCKlKaXtTncQCBC2wY8NJ8+migy0IYDmthSS3VE+nwUW0g5gsOCl
CSQpBUnQgL+QlZYw5WBU4meSZkoueIPzhg8U/NUmkUzD4kE/OIz9beqLf0P175T6inZefEh4y12i
Un0Z0v+uxBmrC3IRuURTzF/1e5c5Zks282eBGt1+/FoTWVIlcf0+f+fyNpvraBVyxFIfAClloVYH
VADE3hGGHEELaqQIjUpdCKRzsH9af1wmrYlEhz8AMyapFnDMM46qpaKRl8i/BUawwR+8uE97i/rv
B/f00U8ky2QWoJf+cgp978rUfqP4lhqh+o12FpOW/6OS/wCHVLBJc5Lm5qJ6qu0AVyhKl5zzupyn
f4lQ3+BxAOBuIdXwYs4PA8uc5H+z9Fvuy4d6o/+VdsOlc7p4Pwlua5KFCE/o+4rJ7Xsur/iWhBHe
6cbqH0/9TcVYT8tV/tndFFdhKxDa+TyuAv/cBv9BYemrJn3BTo3gg6JtbJQvOvaSNdlh19JnfHTf
7RjRJlslmoKlkSXnD2nuoUavgFm0WbE+bfciWjAYFuPsl5ExRjBj9TGFhzNM0ZYnsquSVRxyDnhz
hTPrK3ksSE4gTF+VldNHZQIjSrK/HeQGMeXjmMMdHUEy6bgQQq8Vb91lPi4NAeIrx5YRHkPwYFYQ
S3NTm0zjlELpzcy0RRR4WnoJnkgEs3bzNXSet++swKG0t+/zfzl1E4vqekWAXWW0j6/RNg0NQ5eS
g0IQeD/L3r7YUwD19uNESTeYRqGLwRFDdOMPMWhSTAE8fGKFG6O80F/eZkDrfrOLrdNwcCav7fvV
QtG4SjfcJkavEnZCaQkSuoSFFY/GfiXQrmb2bBDMn4eDv7kw5EI1dTmch2dtUNMPIxMqJDkhzUdP
naTdHE70tnTnXpL1mFTr+epTWH/zsL9mRswgxDsIstBkRdQCS1SiEYPjcxIWxkVRjWhMsc5wyDby
Ys4rLnNvtDWuQ1Y3RPIH0X/uVP4rbGgwTH/7w0ANDMtBu2toPu+xeiWsOw57JRUIi48hy/WRJIv/
VHp75fwhw/gzWKgMxdb9Xz9f7yeyBgwZmnDuiQypnCYRqPGFe/W2F3sCyCuIaJ0/nzaJZQufvBo4
VdwS1ho+nGcqlWtjMKVtEIIUIPkyc7Z/0KDb/61BiRuD/anBab/pO0/m4g9ntrxeQLZWSMC0cBXX
DvPTMFU1DPliWvhQQXet9YjNY6GVZx+0mmHRIkaByaKRsPfl+fsfOzcc5XmPYRMx9IR+ALnGUizQ
w/WioJWDK37l/OQ8Ges+Vuun5jyJq7hKbswRV8ch6JLp/rp9L3fQpnlgzc2VdMcdsrlvXNYfh1Ew
eu8e4+/oWibbOvvvYPsh+vAgl0BMJaktYmVlRoyLvWV0rCjU1aiPD1VacEXTSHo01Z9gxYiRsOmS
zPtaNmJ8P811InNOHL4IMQuFZDoAVMp3dpYu/KABjueBlWtrTLqj1vMXwI4crlyYHzrhgn3RrHN1
abKig8GmIWz0xPTAAvlJhgXd6eV6+si2yYbDlIjwyG1rKPM5S8RGv1eBHTkzULEB1C4cma/imbOY
+qHrCIMsAaHnmFOk4R80nHZnn+QtjX36YvR/tk/9QE1UTuokz3OkhRMyOsOcP+zY31/di0kQpShq
Q4ogUa9233lTHVyJi0UMSSoyLED5UutbV+PNp3SFVoCtJhZrHDrmKnXW/Nv3x2pu9OQB04w4h1hW
CJhDIbB1pgN+B2EH70PsyjF24b12W7lv9ZwTSC7s22YPsdQT8Wymje67d2OBHCLVsC5igl53EYfB
dovwhxmeyltDrz68p2alSwXyanS3+ct+80bE/qp9sxxALugJo8Bs/J2LuakPBdB/DOwicDmzoSbr
7C9cbpCqHyEKphseJdMK5vXX+VYUq94o357I3VFvBnO5CwduLl+f5kNT0/PU97hEjJlbaTnt7Gd7
jImiinI/2ueD6IEoyO2jIA3Y/+BM95lfA6QDYFHtiI+Wii6tarqbc3xYpwmbMRvtfOrsxx94QXG3
eLChwj5uchkenYYm7oMEb8BzXOYwkOnTsfag+6J1iSxh408VJFO6L6Ahgx5amIOZ4LkhSTRwPv5d
0NEUAOjmodVruczYj6v2bStIBy88C4m0WytyA5mK5EnJrPqrDvI/6nYH+4QLJrIqbLp/AVlzXoPC
vGgKyJNsaJ9LSXRJsiHlPVtgKPUzpl/8FaT63zBaFLRL2kh/fv9Y377ALS7TKGREHoutMI1p7kNz
+8PY6pMiEBIFAeAAfMR03IRe/f6HKpwn1A9nqHOnYc6R6jEWpHIf/lp87CWCoiM30hPjnMRvrSSF
+ARdXZgW7KCZ9iDs8aXURhnrL8poS1TqlJD6Mf/7HKniuT806mYAey1cCfLc0oLEG5kHBnpwsp48
z7rpP1hOftw5UJnu/CnV0uacba7eRkbWRrZaK1dETtkPnZ3tjWgh/34wMcJSyTRUwlPcwpSRKRo8
ZXuK7MAfmWMDTBADbjXbEpgxNiLnONBuhhJ8HVld6+ico7rrViA+Sd4BRi4hPwfAw0v0HQ9qUoX2
Ak9uVwzmbP0tXbJcWw5NSvU65rtbiCSKKScBbDHqcGPUFkkjMmp2QY20ycvOoZurOHsvEhC1ZMlg
tTK0CLV3gwIaOqQcEJdJoBCd27lyX01ihxnIAvzzQ22+3arkyEorVAWHlO22k0ISijEefDjrE7l1
4uxeoTBK4gLXRnGdu2MQKfq56IaeeVMbUWJodfT7RBWVO4B6RPaMMTBXTK6p1Pm3MLQddydrlsk2
BTOLoQrhq60pp5OkUDWd5IZtu5ugjFdHzPkkfLsj0PaB9FoJcKUOrT6u3upohxf/GYQQh5HM9+W4
2Ewg1NA/mUWEwAsS6h6OFIzuvMqHuvkOEICNdbbS6fp52YDqFOhWNX1k/PqeH+HpdVA705kQvky9
z9YOoRsjMpxUee2Mqi6ClZKM0inwNZhKJPO2HHmPN00QRcEuLdnYlA5e8RJpWb+5GhIyehgqqOpK
f+zfXhgDINnTM6DoTiZs1d4F7Eh7MqUTzrnpia6cyWkUeRZIkHVZKoybrh4W070EA+mHHQR39e3X
wHwmWv9nMtF3gVzeGELhUg5qr55nWjWOA86j8QLiHB9H72U7Q07wHB5usaE1QG57KDEBxtaiZ2ow
aa6vagcF8L2yiNJht0otY6yqwpFF01AnpKbgShTrNEAog6Fi/4JhJS1VYBymb2EV8ikHEfOBYN9A
MycfQytL1Q4dwOVszWGDHuzUIUP1xLzNsHE0ADwfhkjVw4+HKizupDMzW7c0K/rCDaSZ3qN9HBQa
fz0mjGX0zLB8RA+TqHf+dJLISPBW8hOicMsCf1/0MSaBUSoiRKsn9oWPMEX5lTUz3F/U7SO7qNJo
6KSjMlwelTovymkdtfXJYcrlSDqnW/EGPFDnsFUgTuuf5owPmWwpueSWCmVXDyQl3l/bIhMt+YBD
buuug6/5Ny/O2+Z7UC3AUy/U/eWkucbzEdMfk3zLcAVnLaNIqTEBjQnBsUz6HAiVy4KrjdNU+saH
ItyAZ6X/GZ0hCRWLyBO9fNw5XmoN2erJuYmOPuvf+14FKX7iFDHE96fjkkoIaBhP0M8lM/ZIEgKt
fvRSdS+IW5SdOlxZsQyhvDUUn/5DAZubvvJEDAkbUo1UlOiXg9YyHYUlmbD41lqUvXxWDPyfkY+R
il1xXFPYhbB5MCOJ/1bDY+zeCNA2zKMbLYKago603mhefLzPooYOipOt2pY5tfRd/IANl1So45BS
P2Xu77BQ9ujkSz83Bctgz8Fe89NhtmFOoHtzRfnLBN73SGPb6RahfQkGNbxaOqXrQF7h6+AP8Wj+
ww2Iqpvw75Fk89khjhjfDAnj1+7tDFppvsP6gSMVk8DkLF/upiZLGOQlV99V9N9Tr24i5sucimIg
H1PFswNagis6jXxVzBi+tjaWfn9nJFXM+/VUibMV0CvzmPRTtQyS7CtGyTSZLJvk7419HgQc+gLo
oI+jPDcJiDSZ42nLbcbjLinrdAsYecUCcFTmpwPXVfnHo/5kGfl4sIrl7n+pZJIuWTrFIn3lE+L4
6tXSBzLFHdQpihTkqaV79/RUQB97Z4E47XTf4A0Zw3PhqK9dWMQ/ko7sPQ12iz7usssj18cpovYo
Ovtc2PtPURoIscB37Tsjy/3GecIp7Am5prEB3TVYNVWKbEd70Zxp8rAAePBGU4P4MVJAywpzUZLf
yEyTu8aZ1nZZxFoHO1AYl60iFPCHr5p+nbWvIpx2uj8t1nJtTCkHqoXNRyqA2uz9+xgCqKO3p18j
+XJ9iT7qPezexLyW86n3cvQIZ/z0gEvnzQHmguDhYT3MAcPsLlQroUISpaLdpk5FGd+Eww8kiXo6
CpUahSok43LKeAdZnd+whRWfG5eRuieh0flcbmG5R5yi2Y+vsj9zBy94SwHmDC+eHGawHlM92VyP
OA/V4n29E2dFArt1O4SPtvn+WC2qbcKgm1Iqzkiln5Xwq8pPgDSEJTGiY1WG5pN1YUvNNqbvEWwe
cUoKVC8ROCj+cU1Fadkn/nxvPIG2hNsgOvZ5OpryomZwbaTV5x6ggK19or4HSsXLpMhWKzKnk7Cd
bkk0rZJyy6jlqdmYGLsUb5t5PMz82o/Un5g+yrGXf7GlVHpVraYhPHmAsB5sInFUAxNNUFzxw7AC
bf00o5eOio86gS9uXagOx3oi04slTPkUDudPeJIbAxJqAuAwHk8h1T5iMTcuSMxWnfd/j6IerJY/
hCgKDnhbWyhjsnaAGAlsyXfLOFy2+ddWByAaZw2dCDq+vbbqSieXNP4BoWFJJ2YuAkEp57lHzH0N
uC0xoAcByTiJvIiTqC006aqTev3efO/11O6mBkJNYIqTCXBanYKH8MWObtu+jZ7xa4bWHYqhSqWE
O9WfYv7vKzYEceHD8fAMjWnXrkHdzHcw8CjFNjZYe9v4Gy1VhGRVgBcbAbsF41ZnpLWoPgRI0Pwr
b9/5pCI/OdNWx4HWPs3nK5Pi7cUbKgaeG2RurxjSYQyKK+Ng+Qfsph9MQM62YklRxOJwsN1oCnOL
YtzhQlEttAdPYmZD1HsQ6lckBaQPR789G7Rw3QdoOuMjaUaje2+9lYtnTwElkosQbkeKTRe69VnP
gtwybG9IzfImBIP3WThWFfLXBqvyhF9HqDxFYegbmSKX7+4vwKHdxRLVKbU7ip4jsXlSWyeYcn/p
x0JyBvH7Ie5ZSGpVQ4x08XptXPs4D15XUnUWH/IMa0eo9GPDB0+UqDqiNBwlszPffx7NcXAgf3lN
pEgYvpyegxt7J8oKe9fDhP53Dt0AEMK/T+gWKi3hUW3+OE/coAgMNF9kyR5UZIEagKqL5YFw3xfX
TmJVbKCfR5yCjIKqw7Y3yqVc3sX+hqVQW28F09winZNbV5ZcgooajyqFa5tBa4wB/OJZGosXNhTA
a//aT8MxJoM7jaZR2G9w6etv/r/McGyA4tKmrIv3II9mqTiahnCzhc8+Uv5U6ZJklkPVhe5cHzP1
M773szAAHgxWQwHj4mPRUMi4MDpaBaGlS1RSl0CJJ4Jf8FLlqw2td/dlXjL+8t7sVtDeVY8AdaM5
0TfBRMq+oH71Y8hxLQV+IbKefJ1MGrtWI8LP3F/g5ZU+M8e+RzNi1aSmmx2JidYmlkSwp1wcuYXg
FyAcoeZSSIyZ9zOaRmyvLMvJji6XpbuK0EJXOGW4ocZ3BqaDiDSR6mCIRauBBobniLbXlXE0xQlt
KmUMe13YNKIFST+m0DI20oZmZ74H5BHL3VJzvXdtTFCjzqx+zYr4Wxkw2HOP5pBEvdbcFS2Ck2fJ
vdNSiHWp1uJybYjhLfKd2q3DxabHNsPAlnPmqBfoKWMHyn3NL6fE3/qjN4n8VYvU8D5kMAXvGSs0
Or4ptplnwlshQzQQrMULWD1zTZDNIHEDpWzQfZJ2u9vMLtYPzn2milqN4AscybTe2aDPXZqZFnU2
0PZKImRFqusn19JNXB1EO0+LnXhEOK4cnSn7ww9Jk1xvJ9GTS9ZhlNIbFNJyiZAL+vFkFwXy/bti
28DxTXwRYbL5PgOjfHX4EMWv79btHkKYt8olwtkJCPIcCo65HWNvNY6468sH6BdlfPnKGBKBfw07
dKbWWSUKGiunTy0BKDWepUCdfQmxlCWuClxjR8OhVqi1dEA8Gj9QsOTkjbe5Bsbpz6ylLim/dCDC
yQ/V7i8zTgdZRV7BxxuZ895fi8jWpjlKd2lTT9mnoS/PD6ETU11eQ1+YLLe8lrAH/lUQHB/fdIFu
SS9L6auP+0G7oyosDC7nFrmszGmYozSQNcj3ltzBZGTvwDe6Oia9eak1gZ/3tutK+hycEFZsA6Eu
+Nmx0ZGrMG8YhvlWglth+Nm9H//M2sc40eVtrlxu1otvzub/hLOikXCwqz8z1sc/FYJkF0jMmUEZ
zI/5VBgBNM39fYyUB6YoXeRmTShVY4MYY6pQtJZz3TcRy/Gr3EmVNvpX7wCbV4JYf1B5N+Xo3tvB
xL6WED7xx2s3xAL9d9nl/e3HxvRmRVaWIVj71IYAqOcYV+DSaH/RzNbUeJcASmWBtuMvbIlYpAjU
K9VWnNpdTWCKkDzDW27qVRycKZkv826qq5eCVUFdzX/t2bGYqCvmyupzkREtElMCVqoq9ZmOLBTy
B/1ilGBXT/zf8KeY8+Wdb5AHbU8DGEof3Bar48d5E+hxEJ8EOpL8qyUqT1WZQrjP+RtY1FXtwEW9
zwmVJu8fKO+PEPElfjvI6UqsjcGkXLgm8P62o0foUUkKGTocvz6oXR/3YzEbu9t5Bj0jZechQpI5
n8GLNKnEmLpK5l0fFll2m1i1iFXmgS22vFkIeuD3KvDOT6VcjfbkV0mnwkzP1WWmKkqqHFT8IO4E
R4D5Vh4kd6To4F1fvekYxc1g5IYbObdKLA1rDN6FQIsxcNKeIo1Dt2X1R0FV1/bevDFuIW2nfB+4
QtvyYXQLZU9jUXDtjFuVvCzHDxGLdD64DSXKmfoFZEX2qt70MnS9I3JJvZTzV7EWvfIzem87aJVg
cprMQZLbZkfVWHRLYX8sXVnoE9CqUtzOHSg3jKcOt5ugAp0gaHXzk4hsqkHuU8H+aF0h9c5Xz8c6
Vy+BBrjwhJPBBZZa4dr2B7vV0iQr4SQs2RtsiuZnNIwDr4+FhOO8i+d4qXfZadgDNNLVOwrlfRFH
miSEdRVYRAsFlWRDVkydDyKnAcuK6cZWJZ41zvy363dMdbQc/2U3Hd162ypbG7OcFNatYPHZD+49
IQHTXnca45WHTpH2aRYQZPdgeLzeoCWoOphtCXFe0K+BghdRzOzeyjQaTXXlJ6zgfQzaRtrIdwOZ
/v059XQRFnKAH/Hfe/ad8gDSMjE570qHhyWoNQTi2bcWgKIJ7heCBacPk1z9vc/4Kn0S2/UOTC1v
/paMjtZfvAvS7DDZZpjngD4jYM55YfBXHs9O6z7KYX7CoX/WzMBAIoonebeoZ86/z/HDuz6Tk1S3
guMQSCFoX85QJbANTEgqnWAmYIzrEIYS3rve2H3F5Pa8f8TO2YG547nI/MGBUnN0qAXHs7Foz24z
2rLXSmK3PFxnTWHCl0Y0By67vbjjlZEDqBpvaQyz9bFKPHOneC5n3uxorOrkbtEPd6A2EDKd1Ngn
KiIVeAlkBkIt32sa97TivTdXwtrN1luUHEyPfuABdGjsLFPWPaEyVSBs+ak9mQzhMnwPFPEhsKmn
ob9ZtSd0pz27A2alFll8+7OhFv4Yw50p8uXYjnXHaDFfBT2Kf8Pz+kv95kxx4T/F2fbZXxOPyty7
wR8+bb6FOpayILYDmoKBr/0wX2S5Q+CYLhyW0WeooTeTeVLrtCy940vmnk0glULuJ1DdBEycu4Rz
SblsMnFzYZOKXsym502+QLxdqhvjzgSnbBkrwq/lFHvx/75nHpr6HnAOzFx7k7mBZcT6RDVs69JH
f78Idyd4Xh0M/Vs/vXd87ILJdfPiKBqqRHq4bxSFIQeCnRjMWWFZplbm0PeDcwFT2iTx4BKwPkJI
klIeuGYkfOMWvP4jwLepE0HyRfxi0vNeI401zK9TYZ/pSOiH6YnDGR7o3SGWq8jM75TG3MMiLiFL
e3YxDhb+K7NcDhotiZvIMqRZRb4LrF/cL1JWQ05TyhSqMcGkoVUIOiaNgcuyBLeXeSb47Mi5ymd0
jP2xp3XDNwPcrojHkvW/53b5YYtb/WEQ9Ea2jvjqRy9o4stNCmb6oN6EgeyeiGtGN5f7AQhlqYRq
OaiT3kkCM8/Hr7cv8D25xdbCXslKY0qT3JUtXCY4PEWK1G5rCxMc4yklypyUKAKuEsVQzNXcmnCe
OlW/zpsDU/uVeNTbrcqf7xIkdrDSASbAXLRa5TLtg8bPdto7YoFnszgWXueE4L/hiAgeKWXuH8Ij
DWvB7+8sWjrmyjSzmpFcG69ck2l5gjDy6SvTEjRnMyYR0e54ns/9KAyyAYS9KJBkJQQjZy+O303w
xKLDgdErNT5AH2cwudvX3kDkkOPKiRxIuUjYo3Zhb+oG1BLcaWf0FbjMmeCNszI0U6aXzhULeoXq
EUm4TUhcqPWWu9l7SgUzBtZHUNlHkP6ONu+kFE/I+iaCPD1vyHomXXLUEOyvakeS43nOvKpv5Nrm
/IXvgC6AZPYzmjH6gNDAruh2IBt6fPsEoMPgI6+pFESPbilGc7qIpepFsS1Vd0Yo8ItZEwNR4XJp
JwW9hc0AbCmBX+wfRrC6gH3o4mkGa0j2If2IhFkyrdBw47mdwKQnja2OeZ9jstfsCk8Zf/P5zggv
gHHg7E2lkxqrwbLiH8LcKvOAqNolsOCo+NJp/g1UiKyj4xH3XslXnW+LrS1YTYq2yDPSazOQuh9N
KnBSVPjDAZuYpmHfEG8mNLHqC5+xlndZatMO6BK1ga64rW9tMSkQ2gBajVH83HfZUz0d9EbndmJy
GyAtyHf2OCxFSkA8wvf/M6Z3aSR7vDDdqfjPmOPujneUqOEiVQxxOYnVg3ORHx3+OpDuYC0w6UGg
4OUSOXaqRp46LdZM+8gZzg82lHx42H3Ra1xrRiL/Bu5+nyhKnYJjRHuqbR1ei5xFvkXGTCfN5aV8
b7xTM7LfBWTw0oLa6ovyNk+BJIKlawxZb6NsQtZ/y0sWYY21Ano+74UvffUcqv4lWD0defnOefLD
z7uGrjPQk7d06wJTIKHPS+cN1kea6tj/jSNpgdYYFcq5k9q3u+5p7iFY5m6OfsbosnsihXbL2ImW
34tZVlnBoXOg4z7wX/d7J8KWywOqc0s41RkZl/aSo3/LUL/FVMpcS7pyMIlnf6Kfc2/jN6uB0gg2
tCMLLW2vkfk8RkSaWMWMF33nUG0NwM5wib2JEVYtkFO4OxdibTD1mEmCWj2NMlHTZ6YcI0oVFMf5
zq7pdwQeBjCbeHudt/cdlBh2FqbArCfyGvkzFtzLRg1mfTHDwI1RV16DwwhYB7Xr+GhiAo9+SNEK
1Vc/4AUZSZ3pG0dp4WshirbIgdPzE6YLAT2wVZaxsAg33uR81CzQEWX1Bw12h8O2aDN1dU6TKezD
DR7p6aid7RtXWXRX1d0YnGvEuWkzFtRN2RJKn+PbiL2bhyIrb5w7D1Wb36y0lXVXp9nhQBgoFNNj
i7fM//HRUpHheP/bGKhy6u8Y9sgcOtog+fxx3/PFRTvfCNBAqHyWClIhTGiZOMOkExs6UsO8053s
nLk6LL8v+HoyseCQuO3ft07zQzhviHUcKD9SVsI+Mf3R3kA03dsWdIwZezPYmEo2oYceoGiT+2u0
EAaiCvZ5DDxvm4OPJiCMSgmwz5v6tmTcc7ymEfQ/QLBJw9Jdpszyd6vcaGEY3rt/76M6uL3lNMJh
CR6UTcIwR8VrWC9v+a6l/f31waPOdrs7shNDQ8TQTCZoOnbwTKBuGVXUOFJGf2o0eugMAcs0aICa
d6+Vrtn5DFK16K745wQQp3ghdlscNZNhZ3+FaKL9pUCgVY4JyeKx/0CvOBzGvDfyGOe3v7xnGE5n
nWAdqgB/qlG9BK7FJiy8mv9Pf0svEbI7vVRrWodMCzrjymuGrunX6Riz1gSyqhu2UE9acX3SZkXA
36aeW60MUFLE7Wgmrfff/5CLl/eCL3jnUBEw1DUtDOWidNbRwYwHl4UBB+x7e/msmdcjIsPoLuZd
NqBJo4bSZ+sHSyFlnLPqJ+7COLa6zIMbXytnihpv/ia0lm8VlvOAQTpYlKuQyoEPMVPJowsN2+LO
0lOwcHHyZOt8R5ufhrMBS5j2mq0w4n8TxBtUuIDDiGFuqglCg3pWrs3sgonDL/w75iYdufSC7myP
im7YGBxQJTW2iNsiW90Na364JJLlG3ABcJ11+hz5ITb8HQeXIcTSL7OMEn2dnPFUQ/4lXUO7GHIC
rdJUwfKR9TJNitvSXld3wQYFfF6cJ+D18xy7jHHXFeTdEYB45/YHNQuyqmFN2fxmPiZwYvEajdv+
61DvuZyrU135b8MtXHfPRIwnz8efjewBRwDixw8tf1CtYysowhheEC6mMEMi4G2qb6Le7A8OVrnv
HM++IYCa03FXtT6OQyjzT1omNFmtxF6UaeQ9BUiK60c6gtKG510P479LDlH7vufDcyIUvDCc4xJT
Wp/xaOulj36/ahT13h9cHjHeH36/Y5mp/rsNv+qUr1WEjAZ40uSv4in27acC5by00d9+SdfjcrvW
O34MhtY2BdURW+MNhQGwAw0oMotDZl8XtOGZkQeczMHELZLF2y3zrWqrEcoi+bERkUsb3gYpt3Eh
dzGPqTpSvAAwcxncGFuxcnKNzIWQwxuo9pWXXLw38ORs6bxSVSXelCVdUDHYmW9oHVRX7a/kaogx
lVGbem6IMKzhQV/QWVs9pJF5kkEMSLpykJQPmKU4N2fFm9vN9UWeB8c+fUOKMDyT55sRBIoQ7muT
90yxNe+DfAXdATRNDv0T+ClYhx5biEYSWB6B/Cx4xxXT8NJ4er/p9KyB2g4ru1AsdqWJWQrQuCI0
h7TkpcIV6pb9MmPzB8GrNhZHne9CYDJL6UiFSpHtFB97ULdgo7AIudsR0huixvM5WRK9a9aEQAvg
TpiZVxUDABmC85d8gz3W2F8Fs8PXU4c7PbreiAI/HEcL1wmKCIVfrKd8dtystFxID+a8+Sxjt0hW
6LUqN1+lHJdsV4B3NhGRmMaCGwi5FFIzdK4xcK9UuW9I7Pq+2sA/DVnSBTt4o5tHs2PMFZ+pvYJq
Y0s6ZRThamHNGk14efie5P/lctzOM4zu2ONk4Kh9lMHaW6nlcAF7WKlmWDIZdPcPnmdFH9zs9r4e
2cxo9KgpIdqXIv5HjOVog5OgN6k+2ahQguCID++fLXxPSnyAfbntREqwLlry8He5UNoZKw6s0FPr
5m3rzXJmqZYfHWu4qachqR9ZqbAjzW3aoGkhuyls6mfTctf4GppbekLCbMx4FRWjfcbkoJQKHtAv
oQCAd8IroAACJHCblL78qZ15QKCJbft0VefFAg8U2gDnewqAk/4NMmDysPis36hgLvnyNmrWHjuu
mJnSP0gbK1Wjr1xNb00qrGuJyr9KBuf03l6RoVtBF9J8DRFb8+R4j/QmCVl/uuF4jdAmR49mw9fo
GWg7bPXYPuSLF5tFFIDqUhde1so+MjoUxlGHOad+9sGs3117DJ4lBaDOFnm04IkC+Z2pYZNTv6RV
6sZ/RKy6r2hldmj53ZCBbtqXA4SZjwvew8f3aktkPqw46Xm5sWs/RtJfBOUPgrBo8zC22KNkEaYA
XBKOOYIfw5YDa17uEDLwrVTaN9i8Ar37G1Y01OpL56onUQFnbPgmBwyNU/owLrX+SxDhfk3JqnaP
pXO+FNlzqBnQbrKpR1+4gN6LjtguGRDtZbnR1Y0iVdQhVwJcVDoAWt7es0EIhUk263OsTqIgCaV+
qeip9AwLYyCbcFC9wXSVlOnysn67IfoV6BdK+ZTLVCBK4YSERKRyGE8GUiLyqha5oJwZcbIHfcZ/
OMNHVysewS1E9d1zcV1h+iUQl3fNXFNA7hFWtLKxJACM/v/c9256stRGvedWMgWdtaPGDN5ufI9T
/GNSawi4dvgBT18IrXgwvCwyS9N33x1JUNu94faLDui33IdWBYwgvly3CrIHCaw0FyBs258PMVSr
gmdI1f02kw5IN6Eue5X1Q+XDiVSFIGQnxwht5tcGHzreJRWfrDLvyy5/ziZsLiW8wA4rAwPouhNt
bpacDWBrbi6SysPMEcSSoqkSnO1rWvBKd+RtS1ikYEz9zF/J8gzy0XgQ9Qylu6A9aw9dk1LUb3EZ
QRnHJnusBtALAkVF2kB9nQP284Q2SNCUyXupi5klNHcCKNlleebTLhjZO0046FmVXCfoY0mfOi08
22cewIbzET6/bIDAUbs6pcdVSnPOufqiJR/iBLGukklfJ0o6d7EO2kfvRlUAmKWwU2u2pN/mBjEB
bLynuGlPoRPfQqTT84Ze+XOWlmv1vA7xdMy2wrDrYAVQkby/73uNEdhUnweqNdocglS856NxsJD1
s3ybCiLmegCq6Iexdic/OAlGib8zg5dzHTSDUzWcZQU+Fv0EAbKTsUdgVWHxxzuyK3qbJAmfnCDu
OokP6C7g8SZV6YIrX1fe7wH2gE8xTx6CEnLQVwjekKVIAi2w9YKXLKPUoLB9wtUmB39H3xwORnmQ
xhiasuXt386+/+IBkPmE8+gDIrx1Psvkaor+/RZe878uGCkET+etuNS9bPuTVJRBpex5yNov45Gl
iGl7LEgFXMwjk4wfV4mztKcbh7p1ypDu0deI4Luxlw0spmLj86YZstKKXSN1rtngjnotnXJBbkBe
hRB1PP7JavqjeTrSqDAMYn+qsBBX6VSi0FFHdCZF8N/rJcC+xy7/WvQd8OiaKoleK3VFffeIlC4V
74D/UeUH4nkwL+eaetfnVf3y4Ye+Zn3pY8EpfbrO9OT3F/NlSXmODhdd+MAevbrMv1SRMqYIlIPM
RurzgeW881nWMLPwG1VBqLz/kOg5/hCr5cstgEDXjAQyHkAWAtw7pCjgv/+NXHvNfiELFT93k8WX
FwC39uBb2X8wPMJX6W03JitylTVIuubs9gZDYynrpAMkP3e9EekNsaRW7kKXMz00ADgBQIRCApJG
/TVAdNFlplmAvG43hTRhSb1rG4ReyjD/VpmeITQsrUUxvzR+C/4yvpJdefKZ/HMJWLauNcXMFJY2
MR1n2mTB1aUMn+bqLlipuCxiWv0oufEwUQ2xbYu8Z8QzyvZfp4XQxucAKVOWG+OnWLUsF3Y30V0b
cLbowX8ZG2gy7zL3sNF40M1KQAv4LGa3/yz+M/woF98EP5Nds24hAR74YSlwEJ4U7FlzHizx/AXC
RnDJ1hUVVEQkUiGKreVeO8cO6wnyfg2Oxvi7yMQCn7cUgBBGnt+62I2VX2oOJCzlmu+FjO9DsvT0
CYrRU/bu16Rqu0ji40MdNbqUYvqeFC+m6tfsaP7Muf00gdEsztvhep91TkM5vpP2oxzux5mJ5F1f
8q7jM8FFKYVFCeh5i7I5U+LsnE1t+PgDVaiWIgVtZOxJcpqed1odnzhBhqFlnjxDzspVzVPhuoP8
fhGweB2j1uZYYNslO0Rl/XalOvR4DOiE7AI5vLeuW+7bgIhDg7TiiDFj9zuHreLwpLh/r/gFK2Nl
lxKR7AUakfT936P9zrvbRVq0D0Mlen+RdNrefSs07OfRqVsALBEdj3JmzKeCBkpvwoREkAquxO3u
TBf8FofZxROYTGixu+LxU9+LhxrdXBdVPBKSw0zwUisJQL8K3qdNw0DGOem0FFMRbwlFNWDI91EO
T2flNDcGCmpBBIh02b7WepSC4vLNcz2qJfb5MbH+MOIf7uCGQ/4fkN04kJrvTKMwF5aoKVY8mygn
MO/MGX1GsLlqujZuERvN/J9cZtRVEmfjvqulyEQXcJl0GB4Eo9vI98Puwn11xVYzg+tWKW4T2p6h
tC/0Y5b0fOcmrLRwoqNk4vuiMCmtJk6vrjPBqXrp7xZkPiIX1xC0VRRSZRbIjTyy19gxmD+y5/vh
P976RuyYPQvFE/hMi0LCUC1p3jHhx2Npu+Ov+OY1UCtWqH7PRpaSztc4c8QBHRMLLo7lJfUKBGHS
sS6z3Tg2wFgDdYSGSa8Y9jJDYOts6+gi/eGqzWIRm/Z+a93bc5vVDkdgtZ4XXJEuknSJi2qOSHAl
GAtUH/jRFKuRZQ+knatBnbHdnex+WAz4c2yn01r8ipT2ycqLU4ZhrIeAWItbpvVcrFuAy3Nj1XZA
A8xETRMFaafgJdMNwmBohxocsgdD53qMujp+5SsFGOw6rPagY1b4pyf/51iUbWfJW14Y87ublQpa
RxbUszXv43pxjhpdTEkTMnhMkJhFT6+xPYvYxC4//ZtHjJWSNEOAlqxw7bpSUPkiS9Tf6e/L/HDr
Sft6AuUKno8FS5YxAxAaIq39PfYdvBbIuY/Wre267L1nKNfZjB4W/yCajn7k3zmtMGnebsBciFWO
EIkiLk45w+pKGOtJXCyZC2uBx6jhVw374P7ukvYxbEr3+JVE4K2XtusorjYSYd/JTlA/bQX84HHT
5n/oF9VKuSVIJ21SxgUFhlLfJ2N0+9A4YZIU1kC/UfnLHUt8btf3SzfS4541ZXy8MxINk+8ejXJj
fX8/R+3TaGrgXmskmFxtD1tPhPuRsp7XlE4xB6PRV353wruSwnhVJIigA6VT4MFUA0Ec3JawmF+h
OvElUnCb0oyF++WSaUCI9653c5okw8Zc8QD82G3FSJbCqHzmacbsPrRlI6gy+d13N3+OfXPsbaa/
9up1cX8coEFo2X4A8ms8LK8KEeBQrgYn19KhYNZcZ/zKApMBWI58RX90+p2i3QbXlSLyzjFv4zxd
Pv+X/feCJzNpUM6pCvw52WwpDynQkQ2T2QfxTtZYMSdxtNMz1p4CSIioQC7t6p4GKFkwn8QNPRC/
UUl7JfNqjIlkRNs7wDaeOwdsUFTYc7RvBg2cdg1BKncSafTns2bhUcnfPU0fK14frt3Jbuphm+Yo
MGXDBX7P7K7B45RogdtdvUtHXILVinSGaC+iZPiUTsKYUxGLp5tpZrrd0g56+z4awBr2ubg57FTE
sX9zO9bvmYXbKoM2dRhqE/0alxpxZ80CY8fGjbZ9t/q4579VNDGEsmg46Hwy/ahwOkofkpJqRNwG
pkBcfSuVqRu0bjSBTUgv8BkwOiB9xUXQ3zqvwerh3Yzf7Qfu0b0QMrl2qIqMOUphCou++PhuG6Sc
/McH8HLP4FBhMYGseR3hBd6nFUiM2AzUI6b+9/0IgQM1YWxH389kDgg/SPJB3TnarV4dfTshGEmd
rsv4DtvESr2ztTjnhbY4FCNeIH0b4/0STjeHd4n4i5wwPzqZqOG8Al7FX21kCEVGNIMPtC4uC7gX
+zbjAlrF/DRY7GZYWL6szGtOZ+LjS0svC3eMFEcVchm56Lo+J3VQ7thf7JLya7PJFNtRZNfLOL74
wSdNLdNnNmtHhfsd/5z81XWzJrTt9o1iaz/s2jcbRw4aMyMuZEDwt9dNFFyG1f39Z/X787wVjNrt
uMISaSR830uQaXUXpR9lZQS/VLIpB5rY+J8WJXZfVYpMIZDF7L2Jj0drQwg2o3BvnRAc6LAp9XgI
jgwvXuNlVsU9TppZjFlQvZZ3LyVUw86a4oc3fHS9ijUykP71QRya+2mHz4INwNk+iB6heLVmsGM3
Ej3UO+2IeVNGyuwCBxkon6JzIK6lGlVgmNsdslCeToChG/IYOrLKBUiy5uBUIeSorQATt4NGTLdZ
BCg4goKKBCd2UVGGyv3rxP8rt2AcSl70LrL18ZVZihW+W2yHm7DzickCl2+noLBtA7TKu0dOffsi
8+Ygx3KQoo6+y+bpBGEyRjyV4e2LAVmhRpGhPl4upQIaXumSycCFThvy0NdRkCRghplzcasuFbmG
qtLSw5LrWz7KX4kbzn6Rvl4YddkGsUs1z6PvLd9DIsXUMUiaX78nvkiARvQ9qXQu3Y27KVtojioA
uPQfETpT8llCe5gy9DpAH9D7U820/IXA4Hx7Vb2Ub/cT40k0tFcH5u17cnTZGZ0+vQS7fglYOups
oX8WAMndy/zD9+UVU5jTSM8s3nTO0qj8C60vepFwhpbhCgXWEqUKgVjMsTU/hglkOFWvGyJJOEMr
4vDBWgJ6xrNXQvlD/anty56jgm0+efivROXTyfLvsNZKv9smf3qcFR/chUJxiAlugwwaGl2ktdG6
PvFJGDrBjmo0JRPsEPtXPBwUAY3Xr695hlvQwf3S9ZCWtAUH8yLf8j2f3KbuNmm8XDZ3wpa4Qu8M
3XsNjJv2PxIhO+sOYFV/OmtCzzN5Mm35evLH3pcCjkOepXp+seKhXPDGhd11Pxt1xqRK3Be9/KB0
Ue/uaEaZDOlKXe9xhy9FE8WdI4RQ+eHKSt+b8E6bubz5RuzcTRqUd4HmmIB3K5i3Ay75y0p4Szey
ZwCo80EAZB5NmBwND01TQRfU1ZPUfkuWB5I2M53yWJoQbOpH2XnqhPtz6D9/IFBPX6trHkhWfqf2
8ScUml+hEa9zEa6bBasq5IAshtc4liTy5wHu3Er7VQkJB4Fx0L8bYYtP8SA489dPWYnOAyeUHohH
qYzjK3a5bjYgMoKtKQ+grxEz6HwKTDo5IC8Agjdx/N+38n3LwzrEOFGwgEI4x/QTg8ReUbWSFaSv
hQBePM5h3Lalej3C/1Zqo7toRRg7KL3WlZkqGoXcRzz140dKuS2YbUtoIwsxukdw5dOotapt7CNL
CtMN4bbKBIPqb21DxVG9QXc8qvpWMX/eHTulaCDGi64MAzDBX8TQWCppPUsRDPBDZbVbooOHzKLw
PSpyj/S8RtSYUyg3caxv94aeS4WqZ/EDtu2TNUw9eUyQsMaSpoETOMeX4AXtp1Tnlbnfk4lycrZf
+a7STx+CftLrQN3m9lSkD4BGXOVPG8EwOQIrMD23oNMVyrAM5aToe3qSs0q3GWK3bNI3RRS7nHV9
u7rFaGng8z0+8viikV6X+8KvJ5NeG/kiXkf40m1JIKFwdQed3v+CbGNOG/+bej3OM1uiTIZwKXUF
638E6OLAfDDotJAqz2AiaKmzvoJEgxzLwRouTgAqIHH3kyQctKWaXBnaXM/h1V92OcZ2M/1Yi5jr
N+ANV2Hv9FgECtctuLXjlvLVeq5AKJ6FmYDOlT0cxG/BlE7anKa8TE6CMMm4IuHYLZneoYMqFAr2
zFZ+yfnszuGrSo5uEouGXk0gFY1NyBGDwNqDY4r6mSqWG2E14rh27Khwkybjsnd5SPkrWeCe+Ch+
Zd5mQ4TAr9/suBlYWwMvIIVKePVCHex+jaf9BHRIg7kuEiXfU2JqLnZWBECK/ZsxoL9/6GqqspfD
2B4A9ubL/vOkwLCmtNK+pMNZeT7wYDPlFMkAvFvrz9P2uzwxS1vZ1koHI57/UhdTKNt0M/wYZQJg
+LZ7lgZrpecLT9u2SeCTKvnNIKiiKv95B5zrhy1XsAuqDfaXMX0XN1KCi040Ncpg5BwUq9KWUNJ3
UTEMpL4gL2aep7WsBhQsv2HjnMJxLJgE3Dsmb7k8W0BdXPsNZqt9wZwH+IjZ1O2i3P+G313l/X+Z
RqJ8xVKLIbjjlHo8xJKI/h9aJYMYFwoxHf//KNJ6ec4EeC0aEs4kjMAl6YLjsu8tytiV/YHuW/zv
rwJ51Bb+GjbOvM7TTaM+slz9n18gmX7rrvGFiQs+zjdEvHMOB5g60kXNnsS5wNmBDloYCn1jLsBH
+1xbjnbLUKpCc2TAnUdT/LvWzB3q3xzSNtibgl5VjqCmTf1/y/i/V+iPVzJRdh3uN1jI6+ZIgLO6
Agj+/wkE/UN8EZdVqf5NzEFAJXujY3YbNx5UCIWHj+yftsNFvaoQW06DcUtu89FcgSVf2DVRURW4
arrhaJ3assRSVBrx+Qb+ZZuOh//pYPVLP+UBLEt/xh3ZWZOUy7vCEnvz+U+PgFxB66KjTud+q+A/
xyNCD+IhmIz8TK3HAJ2v8vLOKp9lGCOIfCesNr7bphgcgcDxOY586Vm5j6Za89XXb9WpVaaP1XH+
UvpVvQY0TGx6Pw1G00s6iXQ2ayDV6AaXOn33VnLHoby6J/FtwJFf02Vh4YAvmemHolsQhEgnq8Pn
U4w6OKMgbhG37w1mg43H6QpiooFAnE4qFxYmIbpsO3NUGPF7h/PlGPQ0CtdBeUotJT/GLwV/mp6d
IcEgcvn/D04pdThuHBZiBfQpB4ADxdQmdUNYGSga30ErAvP4oreJTXxp4Pge/n7xrZQvPSlkAyru
jQuPLAfgRTxwBnfGAb7FphWmq2juu6FmaRLt7xE4l/XIFW3KevnP9YZ1ye+rVOpkb6kI999EwsmI
q8uXUrh4fm+siRIwmusW5zd/fCy1l8x1wkUtqzperOxzix926C2IgpJTwtVOqMNZFVCeVK2RSiHh
9YVZRZ0YFBIPTIQPL3Xfx1kdXCjXwoHEguGnw3q6cu0X833YaaXFL9mF84Ndg48uCtHE/A6G/MDM
JxJwevnuhcfnBrs4LP5/3cLhIFVeOgMTRrYpXmhZq/YX4Y5hlSiOItpofJwKkqooE/rQVV7erJ3n
fSJHNUKWFaC/3XZ9fYck7x4Iyt/JJqkMasoeDCisAsN4kQB62I0TZdXncZAXpyB5zZgbjgo+DnFo
rgbySSUSCrLnJIcveZNXDCMcWpOvjEDmgyvnJ+XMZrVNfOpf+jloI3OC4ndzjgiLt7gRAyqwU6vN
RGEYrrIEyJ7eXfZDCDztmENPHSrmVMfW+X7qzZc5pGM/rv8CXHVGMSG/7AidpkNz9MaTyojP674A
emqvZeR/cNczhvchfyQCuqKl1lyhxxKV9BtSL9FYS3Va4A1mRmlmpBF8bynpNo+te0iN2acOzWuR
HuAm9ZLG/GZ5PcOepfCHxFxjktRHJ+Rx7iQN3pE5l3pik8tIzTd4BNVRvu824O3NZUiCfKLk/UOI
V5RXIJZAEMJHJgc9YFPzkkXBz4nEz2G1xorOXyWLYbU7n7gXR78OzCfx9jOuvUgI4nndK8m/v0+s
gXrAB9TvhsCXCtQWmxpqRCWoHxjnXtMBAkhsikJiLZV7JIRcFiBLOkNt4fI6XxvAEEN3Uf5KOLoA
RgchxIBagw/WwiW0D/JDqbD3I2KgxGAb7zoNyBu6NZI1FDAgytN2x4HYeexGU3rEIJJIghE5b+yA
mfgcwND7MShmZEP5FcQVkkeX88inKQCsSRp3zFPbP1626DBCnRpfOZowMNy8CwCYidHTToXJodl5
bc08EQv2VHSs03z/ffpMx1M77r48Qnd4SpORVVRTSHemuYnhKIyx3atXliflpw3hKvxBFP1s4PqV
wcO+v0RXGOr+FsW0Ot1xCyiV+NZi8NP03YRJEZN0Gi4IWsVCzySqgkLy8KSK1yj8div2/SyZwU+T
3TdKCwBBkmQ39PsDxI8RrhJOjdU0jhNGweqkNsmOcYqX0Uha8fK+h/rnZYXp1dpEKMHcKIWt8ki/
kYaZVCm0KuOy10/kfOhW5i/ppGGuc5Q8ht0LBKovUkys1nr7MCJfkO3wQKpgJbkwov+aD8a27S9t
0RGwbtQxvXax/8GGDmDOgmwPCI4MOcIIScSGWlr0mjd8KHieDViRLNAZScVkgvRUPC2LczaPPzCc
UCkSyv/gROE2lCd9zzJSFcCD5kmEewHdkoTEJCvIkUAUEEYU7/y0xW43axWV0vB4bKe6VVo12K4E
gdMehJnWElQiplLVoG8jVvYRr46jCejSJWDg67qCCSrbuhp0382QAEjFNM8037GxWr3dk30qBq+5
gjhIW9jWeg3PcEUaN5OIjkBnTSKz3EToI0NyMrPiWjene16lwInBG8035xOJGUz76aXJQ/4bUXD4
IWh2/AhHSXiR17rAG5uPyVZsZwbCblG0oCrT+Rt5I5Z/i+96PO2TAPYZMuXJBFe6IuTBDRFrZYNS
CwUuLVWIY+0Hb7gd7ny0HxeZhQcy4KPoZU/MY/eQAYJvqr2JAtrWRNKeyYMvKZ0z1beXl/1gXwkA
6ZkGrn4diIVvxvug+ORES85AW9GmPRBwet6ZB2jEBeoaQWdyizba/nDjfFXUo9wOtgZKyfcS8ojp
XlpZYtJhs1YV9yp9VGGhukoYjEJ2uQLpw241abkYO8tsj4r8iY9xu+NpoJM3yebvvk4VXZhpkmXF
oRw+ZHdK4M861kFj3QSrI/pR8MdC9ct111GldBi+WPwQT57AFAUdLYuiq7DrBec/jc47ikU3yzK/
MpipY9nruUM+mJRSAQfDsi3RwBrpkRxYxgryRKYeOI1rTSEohuF5LoWlwXvtOKQRTiSOe8Ezb+xH
gJgTrDd28qXqtlIrN3plO4jiHe0FXGzBtlKZCEFLfzr9CLhjmj13PLV7recxqQlLEjKtbWbteDOd
0miqmqPeGGFttAIh9z555h9DfNc5sqGdcWPiB81PPDuF1PYet7eXyD9QW7u29QGNx7+SKuZD3iJD
AVg/cTqWP66CqSV2hbu4TaPF5luqYeVVTYCEmlauQx14OoFt8g12CXQBW5YPCzX39c9lhouaZH+/
qQajJyVh4n62JKiDYbmLgV4MTohXOdfP8+m/VrqxYyWzxAqRVb+4KU+t9TeqaX3iuA0q7GMT6ZxA
BMdmOA6F5CSszRlUfdbA3LkP8F00JN4Uhd1Ra5ZciHFZWAmOB9ALb4VHfu5Wm/ENyhVNxElJvdOg
nd3/TTH9urnEJKGnZxoe+mjwXNXbAMn0sBsJJ6UetZhPp28OeHEA5xOGciJ+Gl+BHH+pDQzUxjbB
2n/PzC4y+UkNdHV4Epb1gopNBudHl6v+14UstGnIC2ds6+BWs4fcZzEDYUHM5jMrReXsHLDKfDL9
IbtDkbd43s+a192Ron1L0OIX2M5u4lcCrt/AyyIYUpDyM7h2+GONchgO7b3HLoY7gs3rYQvA9zYF
HYi3WNz/43ppjkbNzO4UR0VoBnUCszsrNSTpqUZHVP59p3nAhTo73zsK8nzxhJVpNtmcxfCZZRsw
NdKuSGN5OHxu0Ks+6hlgh6R9iv9eXLTDRPS+jTOKrcVaHQcLJeCbUPDcAbT6tNAyoNyPQWHSPzn4
B1ei1aumWgebXOTHB0rO2DLHlrpQbqylgN+nTG8IOG7Q4wLmrglE8dsWFmcl4QeY8GSSdJhm6tJ1
wvJ557hnP0SSltNSQV1eRgYrTty+r+jBh31vw2ZGKz77SIK+sKv8tX6WRyPyJD7chy/OftMjz1I6
DwAR07kqC4E6zrMny5UjDgWD9dbYoRxbKoCB5GpURNM5uI+axw5jLVLCsNsBox7aygU5V6VV9fM2
zUA+KIc4iWO+ou5rH6nqbZwemE2LexDDLbs8aUFqCRyU9TKz1+SlghhIy1vXEsyHay3tHcRcl+wl
XiL3ok6+QvfYWMHJKl503nkxM7QTUKdTiWSBYKP6pvlPG6k2Z0PFPETOcGuSZn9MDU0V/TzZbEc5
pQnLykxkbH1Ptlddv2Kvbm0FwG7kWT+ZWIG6b2tHhwEm7M73xJ+KWRS6Z3woJ5aZcyn4lYszOxQS
6y9PZ+/EpvQWWD+A4ax1ObLyJMxGgPu5sQWkF0mcttIRSrmCPpSzwQcqCMYLcbEMECGAUwV33faH
2PMJzNushZrnQ6JNueHs979vkROqJkuhOktgTbUjHZ6T2SgjKcQNVi6Pgjbajs5M8qUTxJoylfZI
WwxIAB+okdTpwkQnJkCRyPeDSLwwa+66YAtEkJtDQxTnP4BBcG47hs1XJSCMscdnqFN1N43KPv1m
uQ/fI7JLtOcz4QMiD9RWauSx/eqKNRRDasTXbx0GiuE5XrSmk2yKwoRht06S/lhliPdIOpcfxamr
uOQk0tJ6m3MLhlT5njLXECdG/Bh8lGQyrlXfVq1pKAXkA2ipmBgF83E9EP7nSOdM38nnYLzMAyqE
MEz6eCOP6Nmg3I4wN/zORdkV7povyYS1lKyYLztqQ0Vrvk2MxedBM25U79CJoBtS0LBlSa9sBOS/
wi2+qZgKoeBOs03/e6ZR+MdBruLYInlGYBYWjt4opik3yQnPcZvcug8BMTxQpztIKyoA+P+r6+t0
qvs+D3n62kzgVfHOCwRV+S8RmVQ4y4UlanxHH+nycpg6kYzdRbFY7Nz/DcuGdp4UGJSZvlwA6DRQ
Jdk4cVBAGFhTfkMvl7Y+TqS4GOr0L5GZ7p1O4BDypCq7R9GWDkJyTkqj9DtQVLPDs/lPPCDyCzwe
VvtyFuNviJXpeXSx8vYmLlbllnwDu+Ka8+nZwWoZ4YTegm9ovz2v5vGfpoZmYm7tWpkUiKEN4cx8
O4VrJifVtyxHMsBIQG2vUVq6nnx1kCJCfv/35pTM8+8gk+ZghMqBV+TEQhzW9auOmNNjXv1TkleK
Ab9w3n6i78dNd7DIjR0ZxtbPYJ5G5jF09U2Ji5EcjKgdrMOGGGHNvunsXgh5X86BnOr8hwrU1F6o
o0FTpd/xPZ6jFIjOgtnMcP4k13gFPf1+Z6XZ9Qiq1SKzhN2N4mcx+anD3kaV6NN7KvooBfvj6LLJ
HYBoBSMQyXcXq73RcczLGUdPlARAwMoagGwY5rVfMMeHXzqu8swzW8GIkYV2+eAkmY3kuGf3Qc9c
PEIVt8F+GN8LEtFbyd2Aj/pMXpKwAX5qwzcfXihmpb4LYKz6Q08s/mPp7wFF/IbhHg3GGeSm6ANa
UqY3QdXeUhYT4nhgrzd1pGsWwMTv/YFHB3+tR1H7ZtGfDeK4s8oP+Kh9X4VpJRvxkttDtOGr7AuM
R8LnsQUo6oyZb6XoUDqGw0uo4Jk0sHzCUGQATvxd28CFUDvGnTPAkaa2Jew3OrWWxbrM/rz9gPu6
P6ZcbJ8XyAp+LJVSsCC+kxhkPGaCVZNwiuvEfvwUXOQEzhJ/HiKra5Vn5kJvnFZCWydUAETW5+GM
MaJNLOHULSTmEw88FOMn+xBQHuUXFQ9MgQ/Vccb+2Cy1y7syVu5x67jVAJ6E6kDT1w6eGP72nDIc
OwwMQK0J5ceFgEebX5UR7JXYHtlWcmQbXwtv1QsrwFAl3rOCeM+Z9nPTAuw1M1BXawLLTWfWQzov
BrAE7qwRDgaxkU2eVjyr2092wOwiSWxBIHSR5eNXqGeJxTl9ZLNPbdmi16LfNKIZ5SeBB3gQAliG
4s3V8Ly/pSz/Hfql+GJ+kQh4vOPgOERGt1WUOLDJKGVL+GhpsG9wkECtczO8qvQtkDNFovojPC1V
J/e8ldBzqCUD4XPwv6pD1KWR2N6+RE8SXWTtySAHH66chQUhJocjQ/SVdl9fRg0tD2+RIJZJx4My
jjylAsLJpZBlCojIBpw7R7ldPSVGub2oVgpBoSPfgEdo7ereW6RIjUJBwo3hZOyWX+gGGgc66SIN
3I2XzBgcNHxFn+Kh7df1KVcsV0sTvAgU7Y2J1foz86PZ9YnZ1qXPrcutnnspSwKe8xz2MPzPk27D
KOBWrxYAr85KiNmbbgqyMcfaFPqaVZO6XPOkV2xNqDY8LjC5SN6XX7/BIPKDvJrQnVdULYyj7akV
6Dy+reW0RVhLyBlTcBWRuPaKZur0FhmvliJEI2R5hUmf2NMDRSpDMH+Q/fIZg5y64m53d5PQPV5t
/RmNTNmkBALJ7V5zrsljcRDaa6bJWtky3KduBJu9luu3m99tRhSGiNn+4/051b9WmBoBhYN+B5mH
QqhuIIrALwOGGbJV4LaS+I6qMse8DL2yWJ6AYUl6QNJBZhv3Z9ByAkPd5eo0tBtBDaVXjj3DuxXC
X78gRnSxfQF5KWS2I1CkpaUTl08Z6Bna5yGYUYEdsnyYCL7W/pCZaVqdfabcXpbUOecqFt4HN+oY
QUrsFSsyiPk7yHehth7CzG3BrMSPTHbe5jBT1kW3RGUeGJ0vi2YVtRGCdpYMmr4C9mQHEa/41xoZ
EwI3n1qkb3l5r9POx9YXtJcaGJRJ7o/qUGivpOUrXo6FXIooJh2C/i+SgLI1CQ8VMOzYcDKl9idT
MeyG4G/FJMg67ukerxb86PYULlDPgvnZpeEc27EXyqXqrdHq6F9qGL/4Yec/Gntc/FooOpMmT2TE
b85JJGyctJbLHvBIqwunfMry7LCFYpRidR12kr2c/Oz7GXQWnALO7kIDH0EkTO/Iew4S8UbQy9lf
9o+ooYPwHPJAFF+kQJaIu6Gxv8jrEacJkrX1LyV0TmxY59mre1QkegBwFBnVEMMfHGinsSFStQ9W
cPh15u10jUJwNmRRM9yq6/dyIrgSv/oHhob0Io3S+RJHJMxKq7Q2vzUiMwJ/ktYGDhcPGD7i8Qna
ySfmWZxEQfx8xVsCVGA+94/I91an5ROsqLSLxj9l13cYks1KWI7jtG4Gs623sxYUHx0RDNnDKYjA
0Omg5bL6AtUGBcsKVhNLxzyB1UJ6L3cbdv5SjTIf0k6BdX8wlIZHAB/wxeskaccrfI+44bpULgcE
ftps7QeAedAd0Bw4GUtbAvYOhb5i2kRgzbbyutjPv+RE+ial51tDGiEpgmfbTBQkuO1DKymepPXq
847boHlGqbnNgtP6QSKAp6jAiUHCb8w7fiLAJXlmZ1U/NDwI78in7RU74KyWxpBRwwJbT9Pq2dR7
4XUHHT/iMdpKx4XTCvt8rzxnIOW5EoxEfIEhYkrnzcKI4+jmMwBcHc6hQoGtfurP4H+UF+NeNp2W
D3aN11VKy3MHr+RE6tf0nBfFedPkUvUGj0JtdkOr6Nyw1JKc+4G0XnfPSxAmP6WAhUR19AmkG3Qu
/nPzYpOjw2x0nnMcr0+lcKX7UQ1454JA8vQoterL6z1MA9tj9BXNqfsfeOh2h5oTuvhTLYm4xTvR
Mgr1bP+fQuKv6tMa8XfWzhhnLaipFjmaWGioM7U1fktMilJmyca1l8hz9i1JLPh5Qoi4PsQR61zY
1Ta9vGVvy4kO5Ty0kMn0E/IIe/BeJADaPohqvCF7gdthQ67YNK93dphhNnpqaBBvUKg1TElA+Fqo
evVNO6s7rl5cu0+a+SMBxM0g7uV0waEGPtOlgM9522wPtecD0EAjwrwAgHfX/dD0iMcO7Ho6W4+e
M9i5ugaw7NBunt+EutFATysvMjGsR/d75x8xHe1FdCu487remjg8QUwcmZ5nVDGidHzPcw7zpscL
vv5tQ0Z08DfLA/0sao7t3u5Nw22sIdvIWq3Jx6h/lIdqRekT1JFcMt7BuPWFIzsW/hVKhv4Hun/6
81WNwdT6JwaOka+xN7UOythx18XA9oMfY3wfSIuqyldQHQXtWIcUL0jTdiJlvmlyXCdgz2qf34E0
DxIxZEBzkM9jpt/X27VinoP0seGkSdWN/jBLQnd10oebwKYk0nppXTM4iyJZhunoZGBMku/8CMth
4d5K+PSpvfgdb8qh6zbksM/MsObxfLp07h0GLDwHB7DRHpkZG7auIBOOfDPuvURD9sQv/VlJYUn9
gsgnYVtVXnsd0tWtpdJClY5dfGX9NEapzxJ8SzdpGRGA4Hg+cMqm74KlqdEYUtdyoapiQPYXPwTM
Lg5OlkFLvm4z8HlIYWIbe2ds0BxKVJDhA6PHnymvMHPE0u0e39I8BwwD8THt6074ApbcbHG5Hg/X
OMf7/MapB13fSJcbPa/EG/RDjV+uHyJR+jmHgGEsueun9JNrXKv5Crq4offuzstehILQDfDQAAu0
+JmxIDUn9A2PPWuwAF4E/YUT1xKRqgR85ApZU/DmGxhicYLpyr5sNvYJ2tS2SA85wS3lo6nPV5xM
7ZnVmUZ3RTTQgX4ytbyboQEuMQb7I/K8XTYesI9qtUaTYeM5yekRjq9bx3b6W0SZetgmNW86qDlV
eOhDNH/8NF3zHw54JB3jsGodwevrVYkhb/ObQ0GaNVcvVj2yeM1EFtNOPnklwB5VhbAugvEewA5s
Ajf1h+dxo6iJLQRqipWyEyGjX2GpJHJ+9kzr6GwhBi/JL110wRh+dhlXLK0Xc9WfqFkqktzUB23M
XWOGg0DC3f+llhrqRde/UYDkLCIUU39qsW1nzxNtefl4+wK8WsluBg4qqpFQbzWKQeSB18Xc2fAj
FxfArRU6nx/hsTRxj8JXOxKkDWldbEmQh87yUSO1m60vBYfJL7/Os5VOhxC9CQX4I4kuFRI0874Q
wwclE87eOyBd8OBLHZkvGzEMjcI4FBfCsX4vM8H4CpW6/GFw1/PAtUNAhi9UI+mxJB08Mqw99xhC
WcXlewInMJP8tbCXAB0SRz+nadMfEj+oAyqnXOxfFcoxiw6wZrRB1Ent8Whrw34+PU5b9BayTAmW
vkLNg6FAoX2/l5Fov7fuTz0CB/G+4A0+XKlr/r4w4k4Fgc7Gdbhyuc10eIOU4cvOy/d4xq5Mn/Xk
9OuwLhdE/Fb2dLyWICmqlIm/Cg0utS6Lr2uvxBNe5Q6t01PIbkF0dYqb3VEOTnLJZ+k53oWBuTZa
XRz3KIs6zCpniVYt9Lsfvbfri1hVya0+l8d2Rqpta1ieUHJ1YqfB38d3fl8tXMytT9vAWLqZ/pIF
ck90u33Qp4WXIYVZJiRCuCOv6rCAKFniQ52bp/5LCzVxviYZXMcflnWJjngEo0uoOrsKSsiboEna
HXpc14qNytYidCCZRfy8v9j6FBNIwjI1WLoVClB89FBcgXL+4QZDY2n4K26PxF5ibMJ89L7xIHH/
1g8z8xHKSp3lsJF+DsMDTmVyT1wJ4lsYTLNCcWaHy6Cyrd+5neFOhTabGJtWIltIXCTZ3/7O1VQB
GYNii4mybl6MB0qcsum94J/dlV/b8nP4BatTWfHHSp2azfIUoUrzDGHFT4jvZGd6AR7RW711g5X/
uYutEUWH47mAn7bhSBfuAJE9tu0sevYHaWM/zwrDvVJa+1dInLDwz3yfnLmeXhw9EzOH4roZfqV7
kzcNyi+qvCMhIKDKXm69N9rw5eXxSH1FdnD+wyWBhq/ZIe/7q+KEKu+2NS/3+usNwlugI4oZqEmL
Q0qHA5KuBpGGqzQoLm0pklpGVUgy5EDlS9Hi12V5OLsHQK/KSvAsIoZKOJ0/nZMjtK9aRar/+mp0
5XClvO5oA3HAtTYtFawJAtrRtc7SlRO2DF1vpzxB84GOqyLF8PxdFzuzMCJUaaxRazhfI/kS3TPG
4EVry0T1JexciX+/Uy9SxJh8f/6XGw9hNwLghjBj78B/kfTLDNW8BRbGqev7B+2ukV/nSflP6UH2
gRoQvaJy2wnnBmbMFd/0+wJkD2SOd2Tt/N8rTQC4EOt5vt53DxqJcdtJ+mVF3aJUQAGqBT8BdmMT
Tuwsz194UIfkfjbzXurVTAeMNL9mr2w/aMJU6sdXeJOHq2mZ8tFq5gtcG3gz8pG9znuLEJLfLcPl
019frgdrrSGeGkOHTFW6NHfAbAOoeNODo0io47IXmOzKx+xDwmgcKusmaB1Y4ZXI4d7lAvxVHrsj
m12nNwCMQTKdMbE5A5DunDOZuetXAwr2iQ8DdoJpTQJac8DMQ5nkUBMmq5iO2XtiISqk/NtqoeWp
PQ9JK54S5LpYftKnYJsE5W8oX4+2yoxuguEefC+fjHJekzOEI4yU72qrRp+aSFiQowyLiumL+mpw
ob6F9MMc9bBS4fsa3PA96NxT1SKvoQtVvRhGfVWDvPD49WkMLoycjJO3QSnurHu1oOyZs2r0jDNe
4G/b8h8CCj+1yZaGycVgM52c7k6B4MIgMoX4k7e6tdu5QZksNIuy2WUB4jnOehJBugTsRXhbK5yU
v+1QpeeyrC69vLYGU3/7Ai1gqshPolH3SktNaWTq9XUa4epeDGopE2Wnqn4/qefej9cSW/c0WbU/
FM0Lq6eEqPJmnPMmkudlxopFvU7CHPKbB94N/Mh+ir3eiDd5FJp4mcmewxsyFNKL9OLNGmaLqFYL
eG2w9CuvIgXiV5dpSj52Hfr6BzNdrdA3syvx+MAmIDHtZKfAgtM67vbJQMV/ENn4LwGivhVydFAh
AL7uZKhCAgEsK8H2dIXFFVK54eHuLCcGPkxfYd+nKC4O+dXuYjNn78djEUNd/I8kSPyUYzGRxgrr
nCOtqbWT79JWX6d1sKzYcGOP+fKuSLH7ExcUCGx/Yrn8wb50qf6p1aQ5Z5WjvwMV/0ra985KFPZB
z5TvuCiWqOlpftErqf3J6BGMdawNseWMd0Y1pQNzwZhVBcyWMorO66rRU5F4DlGlCtC07LluDAXY
ooOWwRU1UZeeoOz8+/izMXyforOUBQwHDbPY9qdJOt63XVileT840SpjvCrMCBfc2B8/zP64x3Fy
CDUPwdr0Eq2FU18IDOb7iZR1YE8AE2E55EhwFX/GgVxaQAP2fUtLx/aQwD9qMqNL4EtdbDgw0gC7
bMxzjOEfBcdxV+BC/FSmwwifVd/OblAZfgIP4As6BwSjKDR/QGrLDwbH0g77iFfNumFwSnl4hLmA
nbeOo+Ql0ZdNy8b9kPW+oRwUb1oCNawzmyGSkckl2jv2MkXW2SpZNqHBx4+zZ7j0TgN98IGFIPD+
71OH2xTwoI1DnbFS+yqSc/ipTU4bnKmlySsJTcme27bJiZOEkRZJjqqylGmLmSKxIvmC4OcjjNHx
OJLF15H4Bta9KZTr2hFv33WeAGXTQVyXBekU1QQCsPcuk5sGV8Ai1DSMqhExXhiBc/tYeC8eXSz2
HzrNFWOL2TtP6XfIL1XYgSny2s3zQBWbLQwjf24ujdzcQUPjoECUKK5j2sijBhNsXQMzF7K4E4Ak
Z7CrcOs5T07jR1yexdqDt3IvweFS3xUL8A1e/IYfN2xW08ep0b02zMES74oaeLX6I0JgcPy0Dabn
TfWLwc7nYv/RxV36B4N9iKN7PxufJYRH5KIokUxf2u51mCCSCcRAsT/VoK0X/II6eXf/Dk+Ydte1
sz5oFlWz8JPvwJfYNZkEo2tQ+DXThFGumx/tuGi/8np0DXbUSgP6QaAbAUy0ydUXQ73keILkJGHs
UUdib3RNdsLc7DsSsRE7l+2p3tJjML0PhEFv+OOUv9t1hwoWFvJJGg8H6HWImiWJFYj1VkuyLADY
6+CGFeRS1+xpbQR2Djg5/2NuVHwUOUKkQRWySuJNuVPWxD03kyBrtkclkM3/ziZbfvwS88SN/0zP
Gl8Rod+W3qbqaHbFeVizxuaubA96uUjvVZep/z3TJmcMb58g2sXYGq764qSMIBRX8d0PNFPZ/qZr
xOkJ6ifgTUi6pEfwY2qdcHt6pQ2QHyB6kvvujH9in2ywkYZo7wCfiJfrYFfsHK27Htkk/feVR5S6
8Dj81rLgYHtCGzLvWLMSgOXSO82Jnvwnia/izb3QqzUNxXfHlKkJ1rKyRnoaBrMyUlYhLp8c2iYv
gHAJFfd9wBzXyC9d+j9w4yLqCJeDVxiJ1xgQVGRzTp/ofXqW1rJ1UnVuPO4zdzwPRCRqJtvGecCy
uoMBUK1QfVV/DfcMkFj+OtZuFNGBTTrNJ/w5nuOk6YHm/e3QaGr5aH0aPiaxkAD8FR7607J1cXMb
hx5oeMKrNI5vj7UEwi806TKDmTFFUlTWPMEUxC2uxr3pJdcIXG3ebCbA+XChbT9/y0IRtjbEC9gL
0n0e2R5eAEPDbjXGbXNTgyGQKBZxs1q6Q9fQYkfM17Q6zjU12WlX+WYQiXp7AVI8YngvIubBIgsV
cxmA4VAh3WZNxVDG+Iwz51P6dmneLY/UI3mApRF3o9jBQwAPaGzpC4BLbSRLtOmhwpZf/kmU7SOs
Q0L/qDbFNr5LrrP8cbTIEzyKWr5iVnc1M5/kJ2wqZ7RPepbNjAlAjurLagKw3I9tcj2PchbG2B1z
FKiFlYxp+0aRxZFp+3HV2vhnWxNuDmlf06ZUVoxpDU2AIYPDIAsFCzAc21D2aqkp7kUTYZMjtJlQ
Yo63Wq3POC79QQFAUD26pASxH9ph4qMJ/D3BfyTj1zbQUm7Te+t+RbY3+D153WKXVBCIDkuPuqhr
S8GAhQIm8y5skfwo5pHQG6QWJM/cpmJFTgVIX/wY9taUV4G8vr81W8E1Bv5czaOvzN6E9zPUdw+v
OxQxrsBTGlomOSDkwjbuVdF+OIXJLwUig31skPVvvDzmplDveoSqM6XDQdWVn5XeVUNHERiJsltq
VNlJagasVsvdyQ9A3IVxjDnV594pCKvi4pzUhtEGiqNnxfg4uSbWp7D3O0j7Ldd3GdXIzz18KS/T
Xz5VlzQ4FY7uKOwWqwZwDox1i8CUmUr5kNKImo+eKfveF9sRwCji7pVqTIV9QstotLdI9IttAO4B
nyWW1oShrsP6R9M5A9o7HPy7QJfgbWQ1HmTFUUvJBdXVhB+X4g0R/TRbvCTL/NA0/QbRkjCfZUrO
/RLyLfobcOcYDs/4hKwgHbzOALYyHCq0xngy+8lN4kBK9aTVunopK0RtFhZMK+b3Fxsb6I+N8G+4
BZx/jusiAXpuqIocx2PqJrKNWhEyM1yzCDlahokHR8khObHCH1yzBIQoSmY8wiKaG1qmvnpTjzj0
Q5hd5PiNeCzfoRitLM6YisqcIojXaiENu8XmIPjlkSGuKHYmr6vIExvuGp8UtLYTqlnVQHx+OEWO
k1HCwSZ0rPV75GYPa476XPiYW/WNJvXMhx9ECM3DDgDsyN76gtyp7fA1V7dXWbr9oviYOLhh/8qi
jlc1GI73V89fy7eKF/AiKgQSpFmBuJmfAp6bBoJcx9JiamrG5Onj7dbvUoSAsqLZ0yCFzG7VHAkJ
HXMCfJXme3jHmwQMnUvTsEWsp42t1WALCPjblraWDa0cLaaYPTXhqq+h1AuGk8rbtmr4He2aNzi0
/h5LBxnQYW//ObsbrG6iWfajqm/nchO4Eg2I4hODX9AxbXNCJwpAeJiP6T7NedyiIiZd6nrbVwyk
MGVbemwMe/wSGyPAFbe29vbqljXtTJXHUAj8U8Pvq2U6BhX3eWyDsEO4X9slMSisyj0ARSYp/B98
/OfJt7LiAY8pHuGV5ydqVJHqwZx58ha2kwUyrRlsduXoc62E9K9iZefeR9MXQF114Rz3Bh9ZNDUa
6tQ89GTWcw6Eai6Om4w1RJwB6pTuG1CC+g8/agXZrA1OeRSUPUeK/DYsIKgJPDl6lkMTS+Ho9oMs
5vlf7Dl+VrGfqJFXtYREW3QPaW8WOUf0cAxz8gju47eDdR9qF7W6d9byv0ZGJ6HByMcwYJ1tEHA1
3vbYoaseuV57Jlg9ZdffY+jV6EyL2T9A4h54L+ny66a+bBk/t+KRhj+H6cl059qFfFuIk7nqqGYw
bfiEi+XaNx4xkMbzIOmqUXrfTNEj1x5fCmRGwdeLK418jTQmd2ykWn8UutIC+vyeWgYO6FPPGLpN
tlSS+ZUZieqIbxkPT4tfwj9xiENLDIGS5qIVfIrVuHXNQRYyjLwSWEzv0FXhuoT0O9V7hO4hx28z
dOuAkccqKnIC2jhiF2G7NkgbsUe9WheGokj3E3kcISquAL+MmlwyvcJ0f6lZcdwwyHQs2/0a8lhp
ubpb44WLntKdKKOKKr3TqVP71ch9YwG5kuPMT4GRyJwQvvyqaY/JD0OPzKChCS0i9FrqHGlkFknk
H4dGOZKm7x/lTSqxQ090aSO2WN5LHhx38Tjbh5Oj1/ww2dtwwvNgPgLaEEW2Zds4tKJ0IxynDsPY
2kPzKDtR78XSboZfsal/FopJVBaYY1eLgDPQ37/1qgAwuGahahHMUg+wdMJ01WfMxuu/DEFewaml
znRnfRY6HFKiL/n9alqWFfVQO9K97ILKYCfQV/26lGBkeQUhAiSv+Rbq+2WfgFpUbLwMs0/Ot4R8
4o1eCy03uOjG5TILQBzHcqwOus9Va1gexF8U8mSueaX/iOT4ZgzjHdbYXzKovU98esiSof5epCap
oh/lttGY1PTotcLYh/+IOWPLyU6BTxtp/vPv6Rul9lqoT9w5bYsiGa89JpFiUi9rA5AQ90VB4iuo
xd8OwaQ3jJZHCAE009wm4GnjKE0tkOujLVFSteuYfODjifaTB7kl2xBfJw+8QvmcHf3RnjljUKJL
oF0M0TIcQ2e6+mkgVX/MZwCTndWeY0gGgvzfzZ2gN4ymaR+HQwFy/XQDfSqItXK3DuZD1s5iXymE
NHVOBKTLItWEsq4gYIbQI/YnfJsrxai36t43cTggvdbBxG2X9D9XOzeoT6MshNtDbp+y42r3kSvh
6ItXBH2a7UCLYaDJURN4wueDUTRor7CltEjBxcnMqBb9iUyV2XstlEZZtuR+6G5wyqUhczQZhy+X
EMBg30CUOqS2I+4paEjDn7i5Hg2xFV9xLGeiXxzcXh9VScbnNk/uzqMYSBnMTmpc9frk6lT6S+Ie
s2vVZqQ3Ehzf8fExGXf5nu5e9O/2VZmNqgQ8R/3I6QPIUW5zk5oDqevefPyLcBpWsm/GLcFmisVe
WzKYT0nz4uyWmN1ROvdpHZuungHvQSX7wkonJhQZnhzYJoOYyedtE1pGspKv5BYklubVDj2skkr7
TSQlftHvD6ufg1d4pwm2ozCM0m5eHTyvO8cvZbdKH2TscRqIqvlaAyVZptIpFks/1pDZvWRgsalP
+uH7QxYw7G0hlGBEJ9/6R/QNbBhMUKLZQFMfSfBwVCjUfyWzaUXL/CyCR7ZQHKgIaC8PpujX0BTI
HFLU2juhXw2SvJYzu3jYik8xnU7ZboW62rAFewRCWqpZOvaybIv1YosLzwXSTqXRPtDVVs2Eo5CF
wGmjgH8ClpdO0tAi7egXLZD02HoGnwwged6ImwoBIMP3AsJEbP3sTzhRb/dN1jZTxP+dLhmEvIUF
LBCODXCEJULvM+a/rrjzwyRjBIfXCvwGPpBS4cPZ8+BXZZec532THl0J7yxq6f+K6pxUJRlU2xsm
IAwEEgmPPFyj+21s8TxmLqOXmSTe9z/oEvYRHQngTOS+Cp1avHjwMe/wzcVp+TZBSp5f5T9/9ZvX
3zwcES2yCG7mogsRFAnpP2plnmrYXVvtDsvPvc8oz4Nea4xUkiyJjADsHVcHIim1tz6kZzCn8XFi
j6YNMenykSbVI8iaJqMXvHH5/DVpk0Y0R0TxXNo83YJhm2wHCYPdeRWJiruoVrOIdOpY5xWdnp6Z
N6Y2xNfNv56z9WZEJaxcFCONJzEVrl+V3pdIQEu4t9kMYsYqqT62cjqqEeBOKHIHmcp56ICUl3ch
1nVp2Vp13/Twyq3rD5G34SDAAl9UTxb5cIqPXa4GCal40RzcX0788t7YhXpzEhTtq0n0RUiYPT7j
9L4b/eoupVeTxKRkC6kUi3G6rqr+7vBReirULONZT4J7RGHJwReRIyNXUyjYEI7P/YqYnip3MigG
BFah5CzDv65RGZdbixqM8sWI221CuaU8XfJk71MsRdBzd37Os/Yt/nBJ7eZNIF7WG1abIw7j5wNo
6wsZSmCfgxXKXjErbckNwm5OmI1kFXJg6L2XkKe+9JiW0JN8slrscWx0v3xiN75LsdRj3bujzork
la1Qck56xXMXLwkTEE1b2LGcdbw/XclmOhaQD8myELaiTNvodvI7qogpHF9z/idOiQ2Mfzpsm+dx
/6iW7/mbDXZsIkAojp9jdEV10guBZN/I8GIzoreUV8VlzJ1nnYL2hJ8cHbIkT+o1ibzseDdo2wrP
y6S6w6MAPI0g+RIvf3SxToZdsTnjXX+POGZseYsw8FfU6eMN/Qb52GBqCNc/N9v+kJodwd08q2Xy
bNH5+8ahiztUrUzfacwbFToteMRtr8RkonTIbN38YdNQr01rlqP4aH097T4w2igustrVcacTGpWJ
6pFD36rIIpIEbHv6c5ovWm/OOy0OylOZyJk10PSMj1yru7Zag8R1DTEIWdz4jclLfrtLR3aNZLfE
st32a5FUSl/u5Vi1MUTMKhes197JC6oE6oXi9D9N9frZeY85RQ4OQ1P9YVjZ4DwRBaLtboldCHJs
Kez7NuEVWQpNMNUjnl//yhH2UlWigASWRKIPax5HH6lq5lkgIsQmBBNvMWIE/qtArMN2RiZHFgOR
fpLzPx3dY606UqnAtULpKpSWelNu+/Z3YsvoLZW+Mw/w39P94vgaKhN/vbt3QlrIhNdMux1zCfau
E2YFdCXKnXuAx9o3QZ9QP1D/Z6EDo92Xvl1MV6htThayD6yD8mg9pSqaVwfZ4MumcpxV5lDT+ZJF
4NVIkcHH7BAgOCaaHxQ+kfm60lbJi5I++gpzN+WFo1r8QodhMoL/VdyypvL/XV4XAnaFoPOLG+x4
IPScEdBArFnFdLCX5a8klAqbr5dIDpdStPAiXxGIsY0J993OpOWIjRAzfKtyohFC+KKfVwLrMqE3
1HRzS0NbEdg8r1sMYPVQJbe80FhE+xnXjI42s3cznvlQiEFJwexx9KAkPlfH1JzHMhG9j8+v3KXK
IZ29zFu+daL3ovX/MxNWwd2ZxOjr0bwhX1YDz6jNGYqPk4i4b7iscfZtn/Ka/wl6kEhswE7CBDlf
LSKY6VnfogBCsmN8sTg4drf2GS/Ohk6MTVKLCsdX6VgpZwh5pgGu0CZLjm9zh0qeUgmsIOX4LAXc
pzhR0TiQa5DrBF/nCTLhJxFjE+ITu6x18gKzd7aBzxQa6E299w2glP0cQI81oPBnB9rAXVYxMxSO
jjE0BPpP/k+UWj4ZqUvRrL9WUQEC8tX3tn1U6zM7+qaiT6RgWHaACWSqbhmxvIIViHKeeiU/HnVX
EqJBK1EXqlzwPA6dss7Zz5EJPa1OkSRJuhHIQ86HXiYl1J0RnCCSiECRK8tTHkzSe67cDUQRA8Iv
ZO/iHYOZBSx49ce8zwKzXSDHCVQ7pYTEtSCYrSbpNjVLXZ7FbDRVBb+TaALmpHnw6BPcliETXPkG
F7wklAk4OEElS0bd3S0RSJc1549W7tOOJPZjGIZ30AFw2cxBSCTSvZ/6CVNnlAmg7gFP9/ttTF8R
n1EapYOrIWhGhJfrzgF4iRdFJdH8Fi1zCdtuNq8iRi+VlUlMvM8rCk1ZY/rXTPUywdsclC1kL3wM
szLoTA0f/BDlExSGKsLZ9YtmU/ihT6+WPHBHtQ7VP/AvqWvOTdVsl+sCdebFC3ku2tyGUtcRObLY
V3Tv1KI341rD/i/1UObLkScTJikSYymXCky5Uen1ls9YZugP6v3BWEoas9fP5tXnYPsTIJ7Tyftx
oDQKewkkY9xXkDGniFSyWL+1cExV1bA8lHqub3IDPB6lGLXFC+DA8mypv5aE1gVesgkszsDokGAO
Z0Um7GFXlXNSMw1JAeK3NHTUX1Q4B3hiL4/eosfrc3YjEDVNffW0KBmbM5uVme9MOYRR5syn7NCr
e2ajlFT6khKCSZu66LtxKDX4Jj9FSsNVcIwbmFSJZ4vbMP3gOF7eKxW1+XPit8jZqSSO0o6DsPo7
OCHsOfS0sJJcww+5xM/0s3zUq+CG96s7Nom9kQ1VUuBcGeQcQ84Se63k8aRayh+wbY4yWMpRy36a
qxY4drYLFpmAMgqxRRthszA+jDJbwmxho0TSVtftUvO3ftkW8jAjuwpAZlZ7BlDS2eJnSz8jiRIK
4hGf9/li2F52hoRAY1d8v6eH9r4nBwsVbd6DCLUVKOe5KlWVvZoq1AvW9OtkAO3hQRIq/uZGR57r
ZFDkPOoaHLV92B3eMzIOlaw061D9zir98KNgG7qY2iOYwA31xeyUdpLmlthQODhUDJAtzX6UfR30
R9+GASSFghGxXjKW0xP5Nxo2Aceg68ZIe4vLj3STq6HLINcYdj2PWkVD3jTokk6zSNzcBziAtj+h
A1+UO/lcW2xNzdzlm35lu9llz8LQB+HpgEsZ/3BmMgKBadgjXOxzIfZQCjXUgH+MP7L6gdK1Ir9M
MgknE1RcNkVLzYATTPONf4MCsHXC4fN2oeCNv3r8ZuCS2Ua9a7DIMCs76S9WiCWQEDLNYEKnjCR4
K/Ye+dgMOsydpVffEEzr5E0ydw7OYIrr/eZACDCLnxcK8PH6Oe2Rp53k8FRjID0gSHKsh3hOCgAw
XPQnf3vGt7o4Svef2p7dTIA1V9WolyK2BJtvaHjUS4bJdKjA+lEgl4ttWS/9CGdglIYnasvFMFFY
9O1uG1KWTFxHMY/8p8xRYgBWyfZtZoNzcd5FNf1KMLtHY+7pxymVzLHIJc/a712m3QIDGBvpRJt4
OBDUhXy+G8VZEtqibUBojFSqfvKQLG9SBSs5HlrS2o05RN/4X59qDilc/zkFIklmJ3waOJcenYEU
Dr0UL5YKuHnoCkKuIJFlS3pVcPr1RmqrlFSAKj9adx19VPXejPm3mQYZY5CdE/iodsZbqV2llgRg
q4VI34D1/yjpCRkdH7CeuTHHRPN3B4YpggumJXO+ulocguJzECjFec3EBMcI6tmOxFWDCbJAkey2
XqyikdkrtCSjmhrPmeTGb2W9wCpXwHdWL8xJaca/GAo6RCo3iI5hfsMRacePAOz8ZNHKkaDXiOTP
cirF4AjfsHr1ViDHuAEkqB/hSIT+iEEn4dWfJJe7hUUDdOLO8fXx82iCqGxP7a0SQcwNw8IFw4Hr
sXKJaAgp3Xiqd9EyH8iOVsW3bDqfJhOBHBenODNUJu1jEri6Uk3t1lmg0qph9SR6qAC4x7gBN8PO
qZrREviamEv9GJU5ryvJYQmbty9BUfbPXhSeHK6+wM6VWi1m3jDkVG25jB3uGEGIqdNnPt2Hzn1x
d08Vdy8fM0gRDz+Hx3AgSXiXJZXyw5roy4jFvQF/Wl7vkIFz/18jhJczrOX6O2zfyR+mFWzeSEah
otO27CtNelquHB/6fOW3R4/GeEGF9vlbg1+Di/kFJPt/NZMMctNs1yvXEc3j4wCipkcfzlEagidn
s5n6lGewwF7jg/2Wb682DKzdTu7lr+z/+CpRJ7FPwrF0rFkqKhGoXTvuW6tnsHg3P5Sp3QhernY1
2ZtgN1XqQGuMr7cG1MmzBcypi694wkAt11rNMBky2lYqnAbvUMYBxxq1JgZHAypSBqhfMJanNJV9
Vx993S3sqCQh03O7HERyZAQNQg5GRU8JCa400s+qVzA+PlztcAKsgiDyIV8kV7Ud/A5rS6gCy6tq
Nl3SBMzPSzkRQQ6Ah+SzD9kxEF9Rfgspc+2LPZwOyooVM896ppSJ1Jlrn/zlqp305jqG3GtyXGY0
oFkf2qKa+X6ccWd9/PX9WlrPxNMPsUqXfUdisafoq4VmpKI2H9hoKM7JZOBn01wTgrNGXcY6L/EN
5URZnx0I07C8wJT/ll3xjWxyRcvx5kR0K4XGxX/mCcBPg6M/OlUgoP/LOb6fot8MlOKLw9fzPERg
sbZg4P2zTmIQOdm/Q+xD0ttiU+k4jGieD+k02FW8NNwcv/cf+FTD+dyzd5GMB+D7wRM45Zhsn5VW
jtYVmI6roKTVQeNrKdExPbO0JxnynFK2oqp/a7cYiWwkUvpEwroEP0ExZY2wpRCtYuy7EY6BWVCc
zvpJnUkyJ7runy9oT2qjXFZpyRV6zxEGBTc+C/nwqu0C1ZM5rPEQq4nZZsxlXCbK2RsRkDIDenw4
d/+cP2xHlynlgDmK33Ee4XhETvzyh02jysMSzKinUmOeGccnSGgqvQwOXvwrdwrnArpTLEpUV1sn
r4GA1y+NEn0io3we0n9N2TIvTs23yXS2OggAoboPVeBZCTE258z+t2Tf2fvq448Nse9v/RNHYrAG
JbmOfxNZ77vq9Y9bZu5+uJTW0TfDnXQO63V8hcRyAqOh9U52rn30atbwHagBumPnXFtx+KKBypB6
KBjewjewzK3xg5cjnqok6bFZM3eiaQ8q3EnFQJtWQTNh0azKBZ/HPhBmZW9yxHXVehZ4E5ig9nxh
ZPLTc4BVKy0UoTHbP6jy9C5trYh4i/VnGANRjbzIEVoDsHvotld8bwP52wC+UHjUWQ9V/HnMD5il
SP1j7hxZ8VOgrinfYXl95wv9ixtG3fj1oJWaIODj1SktJTidgb/ZUEXatsac0dEZ9p8qhWi5KBVf
UFik+RirJtx60faHKNANlj1ySlZJeDUMz+ii21pnV0SK5EWHcnNAFvLCT094mw3XcsCrZNHbx9uA
azUaaOdPJ3LbBoLhNNF7t5rP0ZIChycaroVF+Ix/iJ4y14Km93RIUI/WBtPGq29KDVy4fe6R8lNr
KCw2rO60+BVRkdjqCwTCiM36PqxdPPQEMJXsFhxmhy99y0eYGRswAo70uiOyL10gMSFwLgcNt9uj
5i3yWDJJ4lRbxfcgUXUWKLQrffK97jRtgVnxSII0HdFllVJyJ+BFsFYixUaM1Ps3u9dcal6k+NCl
1BRBoix9/ktLXKuvZ8UvzIb33hxYjDKJxtcXK9L1dZMTJUwt2BNvVtyDw6D/x844cnjHn5VVHEZ6
NWgqA+yjCj4DCv8AfE+Qs1JwwQ9F9tPEFtjCDecY8wAZQBoMkmGC2xsy2OBoXJgnWShJDhNBVtrO
1YQThOVf1zSHgnIgdNBlC55v+6SvvNyu9LvxdrNSvIMvloihbI99AkewQoX1TngOtaB+y+VG0D0d
NXoV2KFS2unxPVvELBrszltVZe/MMUol997RChiYuW+Bt0BLwW9MztCnxVxZfuxYHdfMOqHf1Jbo
Ol+W8kzkMyyUJ/YEsQR2SlsvGtdAatgfYOyxDbPzHHzyk+CBnnLLtdT/lpQUY1sy3QGhCdQ9lfGM
71Nb2JS3K1rL2BZep314zF1DCRtH11D0Cx84+b/wENHnbO/hkvsZjJC9i53xcM3Uj5ZywGI3NcNC
9YmI53qKougLvMqb+k+l5BBPViwJcSV5r7UeRpbf4l27Q/FzaHI6qpT71lDd/wn5+StFz0S8ufYA
/G50FtfdTD/jjlbcUDv/AzyZ5r2rnuiJ3RDFjzBjuCnNsT7/t6CjB6nrmEQU2nFelXPPQT3/EnVt
LtoZ38F9Buwmt6xYaTEpZn3zSXoUPSQoB+3Nonh8/CYjdad1F6lhfqOp9NQcF3UEq69cFTrO/APf
XpRuqvul/3DTSeEW1XWKRSTarWPp87ieqQ8WSoq4Nz72sutOZJYGPInt4pS78QAMi6oxEkWivhut
KjBId7S700E8EtsDZUChNJ/uNqe07tl0UPqO4OZz0Vlnv78V8hMDIbHO1ICbwrs0ojdSuJRzvCzN
oqhSEFIkjzgQ30E3dHGhJ/D82KHJOyzjaTKQuV4BPXN1tYP25iznlQObf0W5Ertrdje3a/9jwUBl
yUl8E5dL2qnM1rhiBsQE27ttErzJakwOFtv2m6nmurr0N+vpeVESSsZrilhzMAIT0FXoZazZ+3p+
fwsudeRq20no7AUx8RcG41ViMbEhPNqdlP5+PSKvV4pRziUzzNwWS9Q+
`protect end_protected
