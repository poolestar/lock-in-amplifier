`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
lpDxXkCw9L6rcpCJhcWegT8ffQAmMuLBLm2dM4ygDiV5xaID4ZjLvX1gzu2JtxIUgIwwo126DUrv
0Ne+AiNQkA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bI/N/TOD9DQj44ah2pqbNlWUTmcBHenKI4kuZsumOj22FBxyynctRM30nylXtXEFzmnuH/mKbDKR
zZoK/Gf9jizFGhlIThIcXkVA4BeNYQ0wbSNuruSl5QQkKk23LpdjmXoRWZZurr+LUa+KJ29Wn51S
u6ybbKEB35niWPa6qkI=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
epAd4ZL89OR6h1xlL+a8TbQQ68rgtmW1Z52i/8Jzl0H+afm4WE2PEN+8jT+fM/SfycIT3xlmwko3
osnh0nIAAbxFQDXmZ4zJfCrvwW7D7lH2fwurtmoFv3k3hDm5zw/IRtRWkn3dxveGo9Q5cuKLksAA
OsDgJ3QvtQvchFIOFAAfGoKqI7Q5ThBdCRly9HRzLqhNxFOx0FJE3ioJtYjbAG4Ux7wUCpqOhadM
Pp81FP/o/DGPDuKxkBQPxK8DGNabiJBR1x9qV8OeN+pE35kSEJnfIJ9VNwfdZusHOpsks04qCju3
RsADFGePEuEMar9He+ikTzODjqTtNnhdCzJORQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HRTLRZhpl+JkFQwu2nYH+CC+kBCGx9OoDOCgXaAFIa5SlGzFM+jPVC5EC4Q7mT/cinD1GM29xUjs
aTiQZwazBKIMcatYAChoA4sDMwzAiEIccofCp/ZbgxXa8Hr55zzpFp9Cz1Q5aMv6qKjFPtsOYiY5
gTeDLSBIZpUVg0Rm4lU=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cJqzMM6fIBtZ5r0Geyzk5Wawcol/+tlXKLGOPGGayGKwZRqLkoWm9cv0+h6a6w34tAZnlCFosNB7
L4KDQA5XKekRJX6q4LXJlX1GEf1pmP4BeuopY28HAlwtKMjjBkoAdhTIO0vh7hLWr6euhRbVR6cz
AvhstA8JBkl1KDYg0ennxLkHyHgNMRYt/a9WA01I8gqP1YceDCOi0TKf5/JFv1D5xQMHi1vx2gsC
bkzz76oEE9y1xoh8Dx/6lvaaUmcqoEkkvyYncu0QmrBDOljYJsDIez7e4u4NYQt2+yLnz8GGboZE
x15IVyzlInzszRQpO0JSNz0AjXUDKo68YufNjg==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DvDZCz3WiJB+XAZp05gtkTmzsa5eMzZcoF2JxyvIFWaj8L+uZ5frd3azdrYzY74Gn0ypHnKrPTYh
8IKpAYYy7x9TahJc1ccWByl5bLOER35ys8DiZYa0xngQyFSsf/xUYQ/smV4xFMTEJCbfEDtzERuo
ddsf8yi2Z86hkVZbxi6vVFyczCQcOrPTqQE9Dki8zTF2esx9Fc+injScf9767LPQ7ru3lOOobSHR
PMK88nG42T2u256Q6tu+HJG+0Pa6xF3/Gt5Niyf4cFE1qV0SQdIlth0ZaWNcg3ve3w6O/+GjwLlg
Xklus+Loc0D4rzd9Qb4AUioLPMhd5EwxFWpI5A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10688)
`protect data_block
XV2JayWTzSZBAIjqCcm7mDm40Y3z7Ek55cSthfc5miGS0VjFc4sxhx8GueugdDhwWyfPHS7gV+GP
GhGGuBzmsJ2TMrs2zL/b4/viK3Mr38ofOYqRIFrbfd7aeeRPNVzyBEVwS6xDjp7uOow0aI703C/l
06O2WOHMEJh9CdxTPRZtJ1UTYcAi7hRHqKQSuHUsfQ4JbpVnWiN9JYQ/J4Mt1NWuPUHSBxeDxLVR
j5TyNDpm8tHjsoZq8MTgZJUxryYKhmpTItu5ut6qDp5RnFHGxjF+HG+Zpq+9KpEdysDVQV11qiK+
L7gEcgmA0iMgycC6qaAwZnbbxilFVNzXSk/XYOhv4CayKbM9r8OULEwwoIb0ytWzlJx/QL3sz4JM
Z7l9OKTrUW9Mgac45NDV8oBgPfnernQxvHuoLWJmSzYkfNzH+4auAybFzl6Bef/3A95Jv6M6qsuw
o5dcWiA+XA5n8UHp0LSWLkUG2D+ZSqdOWiQmg7t34dAZp6+xCCFEb9rpveu7X/fZ32tKDyNZdQdt
ykAT0v128YvV2usATOw0WUxLipKKeNGKjRdRmvGd2JzrBpPDjmtvOpLeMFsvIecOhTYXxPGV8czG
hs9XxlELLT833wHfeLl41pJNc50DNJwxUoNbSwYiJEpIj8c9S/zduZd2OBMDm14iCna/AJRK2ky6
yWEncTylVodTkAnKSI0nfK5HX2jtbPpVRxM16FZT9tnfLEMc+e3uqFjyqnVrQ0AM5ImFECXmpGru
0J/TAY3Equ7UpkzdaxkvTvR1ukAUwnGKee/MlT29jpLOXgvIeM0wlTrMpCKI5+hGeQXocF8O+Q7K
64Oipy2XzPW+2bRj2hkaItTgklUga481Hg0H/NAvHKmAsfwIoqjL+naKO0QO5yk5qHaEFjpRW6KO
1+3dDJcpaStOh2k1dAE0sLY/Tq3JR6GNh3/lG9HnnHYFonnBgj/aM8KjYj7uBuUCmnMy7oM7wS70
RoQpkpYV1Id5RMDXXLnfaZe1o2lIytxlZhW5cejfkRnlsG49VSUIUTl/V/V8gkUELsCUEL+ur1XS
SBoWSN2KBoXSHBQveaUtIJe6b1ljIC3Xt4VwOGlm71e6p2Fr42kyaeabXqpyQOYPd4A4f32Xp17A
LZmwEutYi2Br4SlxtsntkpPOo1nouzI9Ae5A09jZ5+JIC0a3WTUNEaZ/MbW1PDwadQ12m3oEJaLF
XRcgo2EOARfsnL+sfJaJGiqdroE/uxR9rN+8QUmVBVuV+59psiI0mybhkWbxEhWdL6PZNiuZBtI5
+vtFSuYXTwQ4p3qCRSY2y7le/26n9YRzK1m+7ig3B0xz8xGlDLA8oG0CJ0pgOv4ASKO+3owUDPKL
LJCuHKvoqrNhlup/IiJQUqGRM+aB2u/X/XJOnQjaR6hO6GkkRu15bU2XFybFGUSWzedSGbSDS7ZL
tmvCqG1w+VQ3yHA7rYd86dloALYe3ypd3vt+JYjexrm94bw6VaemGfwL0b8H1qsXAK7YBO507qW4
b+VMplru3IZxFhP5R9Jv5LWb6g7TmPxuX6QSM0DL4vIoumTgDRLcaAxbgYZx81srhyk67goIl2UZ
zDRmMmwEjOMnSvCj5f7t4NYZT8W+f7mve26ejsSlqJxcHDGAjUZP+7y5mDBo5vgGiiwJgo7d0pxv
TXXAQBdZESg2vt8wLJCHSb8A4gUmh6KU/qRUizQL6depNvyG0LA5HxKNacgatG8P0YOHsfba/Akm
G954dnLxb/g3oLUhFAGaV8mXry5c7VTmNY1eMmc9sFmNRAaxsUdkdUYXISHX88yWmWH6rPff8Reb
06o478FWWpeGE9nfl3lu+/Ksc03ZiHF2DkXlpUQAWS6Vt2D4LL2oQo6paoPY2QB0Ayucm/XyA6+u
FQx31PAGhN3R/hvssNT0kp4rqAY/Fm5DAD7VNUHcY2A58Fq9pzNWScSaeBW7WPrQ4NxX6QuOS0du
D408AyjlkgdJXqqDvqTvEkz13l/LI7PKTA3auX54PGm3TUQGJquay4/UCCROuD94TlvmxiDK66cn
2Onw+2liJ5mmdy81j1e3UXtw04Eh5VzrAnXc7L7ELR0vzG4BYcfJ4ThfPxCKSPKbWJl2K0jzkAmG
XiNPoOikXwTOM/hkfsYYG1Nu/tMtXT1BLrZjAxj8Zk9XiH3bdBFNeDMyqk6eBS7oSUMPUB2QVk6N
Kh3YJpo+suzmpxw22h1ejXdDOLjnwBf7QL8L+TJu5k12HaGDPt2KpDtoxOWenoOBSJ2UMGK8mdMZ
WemZWV7sHfzh4CAQocvCOvJI/HvkfbvXiqkvI1nocKuLpyWH9mwa7UyFLyhwR5rADTYCYilduGLf
+O7+NWT/ZzULyyCPJPZDMXb7yLZ2pK5L3nHv5Jw/8c2VW9AROop5F1vL+aPwgoFeInsMvkiD8uRV
2E0TrCtgLUczpwj+eHmbJ85DVV9x7yPmDJ5JIZd7utr7PHdiqwEfGpYJmDGXDL/1icTWrHT9nscy
ocxsMnjoEo31DRZfTn76eVRaN12iiLhP/NCsX8QJo3rG0RA7Qfvy7JUK2HsZkn2ENS0mty7jSPF5
ugemXQpnMLB9Co9t2HmPme8HSHGaFQ6J48qBhASSETLWoO3lqHTmAiOrSw21zbuz+w5EACAULJNy
agukXrwUOgh2uN8edb0oL1gWG7dvh/J8XyTfMYqO+XP47/aNPbb/Kq4dpkcVTP+kSaVeWixgQoU+
D9f5uyJnaKtQ7b1ffCN8LJZYp85pmSQhA1D0gOPJiIgdWTJZL9rce+B3OgVqBf5J349u5pp/HQ7F
wlKCLUAL4P8vTIRs8MbLYuJla1JCH/EtC+ZqhooisDgLLr19Ik9LH58qD33/6z6hWIlyKN40v4+Z
Y3+qSQpxEGIpzebaWy3ZpLVx8/7qseetUCqGurrZbAQ9KdWp6wt7+KFZUiWTBchk/QD2Oyzl9sQn
mIFl+bIs85e9QVWr6zM2xPPRRI11eNDs0UvwEP88ZuCwvY+QX0EPnAfLhaaH2cRkzOOoM0khFbwb
+91vzQ/TAHZUPNXCulFTxm5g+72YvpmSMF1UaRBoVvrwFBbONcbvoRXmZi4zaBQLu0/NXdoFrP5b
+TZ3m1V+giME/1QpBtBCMgwReHONSkYNSBWJy79yVMnNbUikawj8lWBo8k6mEsS2BuFAZRR9QJTZ
+FTQdRhegsl1L4wir5W77/gc2jWfSyGlTUZe4687vmTk9n3P4eSoXhEWGkF+bCV1DrnLaQuaW/T0
3mekRnVUST7AOd1yNzoTh+CFwBIxlMPEghPvLsiw1W9/ffbjjLKhBZrlZ7cpmqCG/zuMFTmMBo1S
JGzCQ0TKdjD08jGMq+tpE3K+1Jw5csIN76iUyh/zWc3JeVVs1A2k2vD+/voHM5YxxR5E3g1d27WA
fX0orOjNPFfJkemo9qInFnp0mYLoSZXFbNdLFwi4tJsupizWgN4FLf7X1HOUYrNLo8bGF53rwkdy
MmernZU/cE2s69XCZwUrGdKgSJxbC0USxDRyHisPDvrljfUqbJVxqR6mw2hO8FqAqyJPAPBf4XKp
WkS8rM/agpKv05LtjhcxZr3sPbUuwLAEiCORfKx/SITRaNyFEDb+3Qm44bQ9YWsiTM4GSab+GyQ0
KJpQvA5kQVJ+Dv074iUaSiAFZzeoDdgtkf8lrzBRx9ArKM3jHfq+nPQMlXGM2o+Ps/KAtjgcjMDA
2ftmn0RZy72ZZBs8u3xZAQi0+S2jdSGM4auxbokU8KgiSE8PsY1RrTP0wurW8w3EIGEMh77xSGwp
2M2ac4plEM5OSWMZwGg/wVOzN1BwGjFMg4lSjwHAh0D/0+IWcuto1s23IAX2d5zdw4h7LIV2L38W
SPQbN9BW3Bait5Aupf0kRmLSillchMIIyzfkch1v4Bc7UeW5ZdRe6J7F3S+1wMZJYpItNXhGHDo8
LbV4yPdL8yqTEheLuSfSHZ0oKpgiLuG9R61n+BRykO4JAdK7GEwyCQqQj42ibh5hjio/P8PJhr/9
C80jV1OwNigKBSw73WIryAZIpbrwl//RXboIiiiEX3P/QHpkkh7GGXU7Mjh30SEO7BLODi/2jWkZ
3xyYlqhAi5vLVlyrTXF8jy8u5puugi7X5J5o4+Z7EFBik5ZF8YSdipQktUKynijPWGGHr9f3/SzH
/uCg4fyncHXT5N7Oqqi0kbx/pVKMkIZ2d3HcyHPkLh5K4zBIHHuY04fkoad+ZIGcVKaRLo1bjl/6
/RwBAtH3vGx6GW0F1anQVfG72ZmEIU/VCF6wyK9naZ46OdF/72Ef61EYlXJ5VNXv2xuBI0x5praN
KuH4hAhLrJD/dCX8dikI89gnEYqdNc07UtKrte1GDitIayFAtooUbpz2ngXKWfQ1x0hnCqiYAqew
qVH1dfnHCmqdIczqQgyAko8Ax5dbFO/pOSjh3oLhVe/1l/yJYVKv+dvX3MNIFuPpzAr3aX5bTnxb
N4O+YdCoVy41jyfyYtZtz+RzRpLcEiEBrDsANviknm3jRZN0pAe8aHy1gICAC6u4T830ko/w7vHO
wpKi8azv6YthFfKQATAZUYq8xDEa4ZZVGMT9SUoo3L3frGMAhmigX6+Cz1bemmi1gertE6kyyHcW
bva0pbvNiMTeHaFqziP1IAwVqkptcMpseC+VTOCGtHnzjdwsodJklRnIQxyZ05d/y/7bSy0Bkf0k
nmsAjdhWrYZpUts78IChAhiRxrJ2x3ZpbLCWApO7qrTK0etqwratx5hLM9UKdfO4sz2aPBSKPQ6l
VfqVC7EznlbAKJdLNAPOYSvpKpXbovVd58LCbjRKaw4IgtH9ZuaU7t0wL4AB/pPvyrfeiqr7J52F
zeWlosQOT7sFsufTjXACg0XzNMrw/bIw03Ps+5EZVbInbhZHKfgH20jU8xMkBy+f0TJDErncJvhw
7KI2WWwtWlS3SN8Dy8FTGpoqhu4VH37LGwCK+/2mk8/Fg8xrImkyPtEWXoLVIhIidVcV1q7r1tii
XVrr7s0fxI9sK4n50wUpjCHvywNgg+TbEVpwo2Anbv1II7jHrrKe1XXzo1UBhZzirDfU4+zDe7pa
NIwBo7KwByPWT4xgy0PzksxURik6JrtMWRZW/zB4c/4ZsyUBtErqRwhJ+cYuSnR4CM82g8YWRN3j
2/b6mUjq5ZKXeVWuPyfq7YXdeWsincTo2MkYdpqm871h88FLHngYFBaxcX7P7kPM8ldcCioEerl6
8gmVtnwnjXrd8teJlHW3YRAM7uTbZL1ckq/l4irpMTvWCrbKhK4HN3vkrcDTICtkJfmB0qEIVf0t
ZEInUSD1MbJixqktrZvnqglFLzE530gwRmV8Loj4Hs0TqAle/n0qarZ85Boz6oTwp0DtMK2BGrHq
v8DSteQvjXVklKruGoLKO0Ak8N0ny+3/GWCCCVB+QWnZoDaii9L5XHACwgm534ScF+jCIAZUOVQM
JXBg4anvPSdN7ClqIIfzsDff9dBNxfMmltg6yUjwVWzH0x+pNSEcglReHVPhb78JkdyT0mDEzF7X
sxKaR646MEkJsuwQGgTTaUY0bJcrGNlmqMGqmBbAZSRni958B4C72h2BmzsW6RgcmJIeQ40twnRY
PGmCq6muO84gyOXtFtiR7vddvcJIwT+PQisSe7+VhOdcO6BzeBYXCqUZmy5V+I5EwvAxBuZnXzKw
xvUnONc965D29lQWmviUFnmB0S5VEw08MSYXUEqVL8dDdqA/lCb6bNGp97bHT6HupnWRp3qmCQwa
UVgxAGGpWBHj2knl9V3G1Au5JN+VLeYjJZRBp8AoTcjiomcYnvvzIDnLDxo0v4/8ZNbKpKUaJES0
i5kKdhUZiC6/GPcTTU7bH2Ol8Ep12E/yCBztrZa832ERx5h7B47P+G8ZN5dIKWClMdbex6LdnbUA
MH8sZUOYbVn5FilFRoonogonNBPHoGTT1PhwoIuArmsfEqu5GUXQS1IjEaWRZipD3wlTZ5dK0V57
LIHuWRpw3gJ86IwnT/XjVWj9lvH9nUZNsj0kEI76Zsx3aZT254Eb9twQ9JnPqKIsQjtiUJ1mfc8+
SKEmBGd1qHDcWwQFKliBx4ALoGpnZRxNdSvXB2Ay0bk3WsR2VeM/WyTkwE1IVhTdmlV9RqWw0iIx
x6z3Va4O46SG2tjFITx7MKmcWGP+R715Q+uzs04uisrc8tsZzfxc7Q2iVHT1FsM81fb9tdO6y/d+
qs4doyioYKYY53b5vsSKkiMhIk0eH75lusa3ln+yIO+JxYQgmReKs3xw+/WWoTn5t/fD3IC9nvWH
O6FerZjfjvPfzo4aSHuqEeTDWlOe+n4M6I/1yU9lRprIRGiXRsCwcuD7icFEQRoFjMR0uG6T9si8
hmX8AdVEp7C/KWnYKBby1pKt8VMoE/DeZcEPwVj+ooGOfxETp5jIW9WxvPvdYNOOmSZoCw0dQGxe
pqvfnDFOujZA49ZJ3okJnrd49nuQbRB2rlAzPNHuhESomo80EFnHYmoAEDJjvSQaH9zuMUgKsD7I
dhE/SYigF0/7NTYdTrYjOqFcn2xakL3JRT4Bmwo1fhWJDKsOhoZqMY4N216Lq/zbyKMZdw1b3lTS
dxWUQ3VRjqO5lalt+uRNPQ/JXzrMks5PQTmDkjGakOsiNsjoFxB0L2rMNtZiwhnwHV5jtpNfZH2V
clyzwzuXCntNZTGNqr4JVvDvKe3jl2uityfYbUH/qswRKOrqMAgYtxPEdy/Ss7et76TSVT277Dlp
aQSARpKnSGD35W5gKy2GsXziSU1+xs0kHZ2FbavL6xf6Dp51Ud3kYjGN98OI+tktLmYvmRB8+3fH
AmVA+8bJ3YQ9PNqZ2XOWhTpk1E/vFk6xaJyyLrfpVrHOl1mN4q79opurMxKewYWA1EEQJxIfhKN8
/kuCXs8/XVDAzbJWJCdk8vCcbpN2wyG3T5kSRPnENSDCUZSEl9AmQzfB/O+uI4fU6GEZNkvKRUgM
UxLx10rpqCumdPIDCTkx6O+T+yv1nnTVjFMk16fxvPodBisuvYOUqGzkBchD46SFp6xKErbAKn02
UBYL2nQvFDbhdKSzGURR6r+PlhqIlHHQ8OJoHmQRr2n7NDcI56I04qE6Cq7WfewnK6WOpun76lLT
R4iWDiSdTgWsi7O69aD9kB6pLopZ0lqvA7ggrxQVRA3E2rp278mIBsP6hNxlIBSop0H2qz+OO+yD
bQGHbCPqryclcelYgbrTKKUaXlYzvfr9TUTMXckVFN/Thi9vcM9aV/0JgLmscToNUTeqyvs+6TBq
n25DxUWv8VH8Vl+I22S0W3Kb2YPmvAjnM1vDsWm50Bj0dJcB5ltxO5NVmLu/C0bF+QZfIDsEk430
Udix3T/7mWH+7zyxnD+f8BFqUUMtCjHx3ro8Zw3/fA8EI0p8yDOZAd2YXz6HIIFrLVszTzZ/qcfD
GZr37ujeYIraps3ZXWvp+5aQCvCI0G55hU8ZXMXFutUempzodfit1N/8zf57oy4Las/ICuCHx73b
EqiJsS20ESsQ6Ki65POsCKYdQmzKzOOrdEBvrQ+8ifxMVv4e8lfu93+wnKMvvv7xp8azlHIhd2hO
5hnEKlMfREr/BcVcA3ZizU6LZ2GxUP1IHkUa2x/81lNa33RGv55PRWPjnSxzE3+aFcP8B39gRKx9
cHB1GP1LMi4AdeetCFfF1ZUGBG16vbpWQPfoXeXoaAqQAQOs6Lwx0IX/Vv4D0FjpIFuaVfnDW9P8
SnnICg5Lhc9OBC7lMzMhtFPu7GgDH7vM4uWpMYVpBqaEAwjPsl7bpa8pAFEVmqKs2nsRZYAbeQ10
Dr10FEv1FS0uuvxO33ce7dF07tPkK46sXYzDIVHt9fhtWNbV4wwOIntjdUN9dg1h9sxEksJpZGOB
dcyBq+GkQzIPRL9bi7QOwK9XpLdGFr2HJwQnhFl6munvyWYKZNP+KfjZb190Gcrm5ySsIvR7ADag
zKn7oBz71+hcKWE7W8pkB6ndnwF+TQVF944tolkd1rzkSmpLHvNWTriC6agZsT3A1Jvdn5gSQW9f
rBy6VROBgGH8BqeEyToGKUb12YH/qnCsK35cnN/+DJbUeff7FsN144KzYxCamAIdZOQdhur9vmtQ
eoZ+hH0mxHQ7jgY7o7QJK/OgGpcEPz/fongIIN7OyRhrOzVgZLGF4AS8OoOd6IkDtCqqunzrVvRT
yg0AtpWVv0gN2J6SWewVPymImm2Gx4YkGIaq8gMJBcyudcpSpx/Lqq+G1iSH803g6ouCpeBgZx0z
riHGXHdc63qh94SXqrLMoEeiTH1QvZOf8VAcTBF0OXFQ5MX+8qxBaw0p+Mz4pGv9ECnDYpNONbD2
lkVDj06cFpTtWhXtS6mBW++stuQKo7ApsQ8xOWcM3j1/A/qRGQAdKbAxCN82F1Bj4t4y2HEm1lRQ
3I1DcqFFhXAioviWYA9FC+9P+2or3JS5lAlDy2itH/vF2v6hQvk+4UY1ckBCI6k9XfQtaFrRf4wi
P2XEQu3v+DPysGn1I/1E/6olNLuc0RcG1xBQx+6nAmJIxYm1wIgcdeTm8lVWAi2Sb7i0XJcWpc0U
oj4TT8QqQV5n1QOvCcNg/SuOLXFacbjzHMk9uZi3isHSQMpo2i/kyaUoQlPQG1agf4C1icLu/ICW
yaQABH1yVjVBb9h1lxSSQOehl3vpLATJ95AytS6sX17RIBb8PhyzyfzRHnt78zEXlgUQxOrvUN7o
g3m8zOfy08Gw2un1rYBrVVY6KMFjiiScPgOutVtJ6PBEc4vLZth9dkyQ3rNYz+tu8bJQKiwTsYOp
Er83C9TrQhsJ4N7elDf5WbN/Q45MauSYbvAzIJokeBzV0dl/M5NnZQqhURPVf3vKb2bZsyGqiwEl
hWIz2SlkVJxe/Zm/6YCHyKaGtw/dbfVzLDLnCbyenHsoxVFtclrtmeggse4NSkawRn6ymN5STvoE
GArFRkgg0XUrCd0PKCJvyEMS6BUQQbWPK+NVKWHcQZ7Gv8D6YO+1nMVqmFCUN+FRA68lVD5PeKUc
0gDvmxFwXGmA/ZYZ2N81GIkwUrl81D7elOiWl3u28XQRcNBRok+pYGSM9CF8hZJDOcZxIcUw3cv5
GLv0XL54Hq3wGftV+ImsNABWpSbFXYAKeCQJDyg0ph+CBIH+k2T9s0O+7bPZA8HyDS9Wzaf0tYLv
U7xdS0Ex1Vyir8G/dtqq9Yw6oAUAVybOROelKgcigo9EBe0EagvGA9VTYkyLRS0WXCuuCQmwI0dG
Ogi1fAaVpiizFGjEEWpxqtSmfMV+vPc9Znt6O9kMaVmwhVf9tRJKl+34DbbQd0iELEYxT04QxlCq
ECKZuX0RikBSP7mDyWmxPBofYqSRqpPLKZTP8A5un/ZREFAo2Fj5n4WewVnsEbMMD6dsMWCME0S8
Rdsw5RbuIgnhCwH7t7w4DtUzTumQiUZc0NdTqowCsev8BEgaGIbt/KxGOJJcnUx2fkVS+J46J6Zo
ST4XUu6qCzkg/+2HFRsRltAdsJxJ7I2CImNC0LZMVNHUjNR3JZ4NoamaME21kgovyQwiW50/Iccr
SiQJ9mz1T3rwq6usdty2p6fjcDuhPpdr6bztz1h46o1UJuJsT4bouKRyTet7xtbnE1o1nvZeXw8K
6VspiXrabV1jrvXLhXQb4Yl9KN4biw9GJIwjyi/vF7cZeU6lrCbx9QvgyuUI4wZuWVQ4V5DUu79f
Rgmyg53D6in+oq8MbRE9FGI6/S+2ULB4PMfKps7/aw1fbeBsqKNqrxLTp+xrBhDxMfdUzhlHFbuv
WC7hf7zGeoWkjBb9+Cib4A6b3SOhRYRssfiSdW51QFF8SMvkYvw6jG8sndtagvXFPpj4rUy8V7F/
pJq+kY+047bfdldzUTcyp5m86726HdJpY0cEvA1lcI1F+UcBF4vZkH7jARyZUW0+uCdp8nXxkwE9
YRz+J5kT1qHn6+vGsiMpfGKnF3xpUoURszJJT0CviJl7XYAm0u53QqBGC2FRBFwpc43kMpJRqTNp
4GfWNPBLmI4naGHCntzt7W29Tlop6IKraOnrzENyFUJd82tqSNH6tyYs1dBdAb3ZnC+GQW9XBAAf
lwBQjGvUpYD5Eq9ukEGJzRCvbvLFBEDwQPs6MKKNX0GPEMOg87nMc5Lrv3L8AuboGQli0iNJnRil
55INl1WbVOLvljS/djMhe5QAZHyaFGVWa+yDjklXmMlVkN9Lk1DJha4y0wK/nx8ycarbffFf5z5U
DBGYgzhfkgVzQ4/UgbZX2yzeP7uN3pCofcDN1PEQDB74kMXtKYFpYezQcWY7tMyvwgvu5v3P82Ta
LFwEu8M0T4tGggRj9a/IFCZwAZ+5d0loLW7BZKzTUQ5GqIL254GyalrGEW6tblU2c0Cb7zodcjAd
/h4WiVx2TaS8LIa9kLtBshFphyPw+gIeptrdaaK+IaX2Dq6J2qub1bMhZg3EC0HIljZAef9np7u9
JyyQrOFHv/fXteCYKe6c/0EN04enpRQGgFe7biD8TJ6qZg1vmdiqgbKo9Ao/wCcZRO9XgDPpQ6l4
btSt1xsS7VvwVdosyrPj42KlCehxjS4ES60b6V82lrnj/ng5rnyaRszKQuKezVlReSKUwNZxQ4+f
4/IoiwPCpqUUEsFfo5ucEDpzZvoBMzxLJ3tBw5fBXSqmHg3c4qDXBFG4HP7XQoNMB92FvxsrpU3M
9hDp8UokSCKbFgGn6GSi69J886JxESjLWE6sQK8pkyTGB7Ipcf2tcRmVX3zLbDFg2tv7m9/3DVd0
lzNL5wD/kzAYB14yob6y+e+kkSfM4fzoQfk2hxNqdvXd3UwvJmF5Tyd5bER2jMl60kTWXoqySuEv
X0KLhe7Yb8UQMfUfTtkLhMHg5V5Wl58Ig9tKntXZ0/CON3SWzqqOfOeSIM2UqUGwmQRrn4a5HIdA
z4z1/ToxNnBTYEafsfOrT1qMjWz7qC8wseOw5jNg+n57pMLUWfG3XgZMAZlp6gnBs7gFHBFRzl3S
1Xwa7ES4n47Fpy1HHJSPNUCYW4PEBnWPNuD6A/+ZwB5qM+8LOQUr6jRR5JEGruyusT3uqseSdr6V
GaJR2xoD+iTN88SyyY47F33WR1EFuUA/OkWwI8WU87+kxmAuZx9Kvl8P7d8cfdEOEx+RbqFYMVIR
epEKdDeORv50cthdwvsruzEI+PlbicdsJyPTsJcsVWtzxnD69tZX+61AsFvUzEdtXmzgGXM4+BLg
wMQBCH9ccXQsZUHVV3SOc5tixjVust+7M8/Ot3nLwxJZ8hQH0L9exrxwtFBosBOlm8/SvfOX7Yfj
G4oKNg9cqCKkXsZwyQtc/dB8GcbKGJYsn6wVhAklpgyAwpajSjSczeYmgyIbkoM9KA2kCmmtjQjo
zBB6f8UNtb39N+R7SmjWEPeDnFeWpXzi2t8bQaEZ9+Pc8ZS3GtnUl88RgjGi0Az0PGbDbyqKPiTZ
ghzMWmCOg9Lp797uOP9pn86vemV2rL75a8TrP4ktGzcjHb32w1vInm8XN+vbW+3YjSHZiuyLbpMn
tydZn87vznudGeAjYuASQdpdPTtGpcoCfU8gVPshl/LQU38TPya67kMaLtZcjh2Tmc0i2/sja11X
Br7oKkoGN/WBmNkRfj4RIfXRK2WSwR+t7N2AC4WP1fSJ/KozeNvNXcPub9jX3eEaG/RQP6aOJi5Y
GO/fB2325mwjbIdLP6HtwK13QEAtbAof6y1xA9d6WnSKN5/1QZTKR3kN1wiWHYbQwmKrm2gWXCjG
vv7fNzcHb0NSl0OFvE5KOwPer7rtTUpGP/S1uzrRd4gWtMhhmR2+Odd7CVLr/4jtS67R1FVFbSfV
nK76UEpIFLHZIrBChAt9Lf2VNNrntD2m/iClonbn4fpHckjnecsWNICCBRz2C9ruNvUZ9ObfKRS9
xDgUwekWQ6ygBlxZRCCQIfcOE0qvmu7hvVGXd1r1m+4iVogHsPvYuOX0zazOHUkj0axXjnxEtdyo
Sjkl+tddXrblnGT0GF3RawwheDEno/dPxA02Wvmczch2vCkggZv5i/h0kHt0mM/ZiqDP2tbH9ZZq
/UGa4LAoA8v7hq7wserpANcVNzE72BF4RSnc7vn9fHKLnwn+ROubnSHU++lhrmOSZGWNwpoHCXH6
qAw4GXJXVTBNeQ2casg5xk+P0Pm14Ok6cHmgdPqteVhBksf5BvRJzad+rHHXAUqj05CLotkxGlux
bfSLUb8m1wGYRIMeaG54kMpxAxsaXAjQyo6Z+q8fRtysVro4tKY7fdY1c+6Rr4cOob4ck8yTpDXb
keJjNzEa6QVpu/TOuwqTFCaEwcXbVbA6iNp9Yn2zoyLflnqtX5j5p8Erbb88/LJ7tUYeUKRZaVb6
r33F68Xv2ruDPAImxndWN0cXQz3ExkDOs8eU1JAvLkpiGtlOPWZTDyAOxki9OnF+k5gliUN79n9k
TesIv4iKD35ueO58/vGBH1Un7bqTxX7sLWheyEkEXSt2YkqAywRxfIWkPS3Xwh/wAX1MpQm0hdw5
oZG2YASF6gPud8P4F6vm4vouD+y4cVbatVal95zapwrVuW9+3FIrvEZQ7kxjxvttRDrkEJM63aOp
CEfrjaPq2hA7xpYGiCyYJnYHWUejo9wsCKCncwfN9HXOkISmasl0K31jxgv93teUGkmfODhAGqFa
lwvaKh4z9XbrHGE6Dp2Dy08/lYMNSqiOk16x7LH9YqF3xyJ92llOwB0gOoN2WHX0ZT6E82xNqqmr
cEW/oouI7tKNQhB4ZGlICowszSK8fvfeP2jfiPinxERORES2Q4ykoRlmep0xrnl1I1jKV1Q/wkAS
d6nRgZQPBDTmZrIoaDKE+nNejWHIhMbiop8/ruG4P9cEdcEKK6b18xiK16L5hn3zjlAqIuRPDQo1
Cso2AmRmwAhO5RYL62IcCEHoTKknUhWkqh8bYMdWqJ+Rw1GmC9/W7vrgJZpYcdO0rqHfHDW3Sqei
xAG3kSCBSTgIRwhUx3laIXp1pTURUOAlNODhhVY+r79B1EM1rM0+7yhYRoOdO0UO9FNgtvGn3mvp
kSiwwcgVhoXk7BQ1Ofs7bz0LhfRTdRv53SGtVm80Hx7cIMn/jaYXsSciOyE1NszIaBvI2U3tyzOA
qjjITHVCrDowimURf5ixly38rW2tblArqtERfktocB1XjcFD1QlqIIidbhdSxjZc/pAFdV547jCz
mBexzBBdW3ZwXjQQvoqGPK5SI0oXf5u3hqPCFleeRfWhbv8hmtJfjbr9bT7GWi8dRPtrZAFnK74S
ZmPLA7HvEEt0P5s3Q4za28Dhael6qWjQvm7E5Yq73qzszr3P9dTzkAhlkvnVx2r8BDP4AnAdthgo
V3pG6ydy+TFKxCTHtGeNb487RfWsjAX+X3gSiIs2W2rzllRXW4Zg4YUklKF+QetvDNtxRwOBtELg
e5zYdCd3wsoIULOWJC7zpUHmwzEs4ZZ4IBCHx1z9eGlttfFEDI+/MHgVDFfPc1RvDRuG4IU4zPZR
CoW08I82E1xeDdbyIfMl4KAdsVIlIjwc1aUueiHqeQxleHmP3mlrJGCuMBY6Aq/SbxFsVyqWC2AS
oI5cWAIPodv440KgOY8rQZYoFeiKZ+mfEjh9J11hIQKUQBjZF6bBgKCynWGa0/Ghkwb3LB3ZDcYM
GfZrufzCHTg/WCRxcdAQmDLeLNmVnlKlcM2smobQhPz+fjlRlox4crZBgP0VgiTX8+L+QLRr+d3q
YeECjG+4fFztW+zd7JcwZmPeeORStU3NjCnGr1RnBtKLFvaNx6K59cs4NY7OdzkmL0KEUMrv3GdO
BtRWvo0nsFo4oJIuoFXZ4Y9vgQBK4mQaK/yTLVIkKECcZyPzEG4AEfTErX5N+4650i2iBJ2F/7vL
ACcNcZizbx6zwM5gx+qbxNn478UREg5KfGxXujx+LWw0Ra8Hee+436d6qxTx7rY/UHTMYdXhzqkc
8MCWGnA1/tlSIVumJT4iBrZ73QrDAKFIG51+mQCSrMh+LYaIhDhaD3xnG9mMzcsaimbdx+h7ts+/
M6Zt6CGgjF6pWzW3V+3h603AwMh3HcsoTJgFPM8xWvZIPWUPU7ynTEl8XPxbwW2PyJ+shbWxkLae
f5Q7AePWvfxPBi3H6v8jpDYnUBWmgxSaSzuO0dlVr9FzjDYCbPq7Ymod85tdYFE4aORhecFO31wD
r9AbxCWryLCVEuGef2Rl1BIC70KrXM4/rZjlr4o=
`protect end_protected
