`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Kx5Auybk0ZnBcBDNLQJ/yyCI2FdsDnK23euP6JS+gndZhQRKha6KCXWhA8+h9T6s5wALNFJHH2zI
wTGtenD1Jw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hrJWZZ3HUyGutlbsoUWN5o1S18XtDKHnUx5XCvkOL3Zi9CP14OIH4CKruKhnJ0ePbQqbYapmIPlP
c0ZPmT5Z3cFIJFlsMfj8xWI2m1ubG6wkxz/9SIR2s1L2tagggnPNJqIp81VPaHOpMe4ocwrblrNL
Agr8XQcGAVSxi+Ic13Y=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
DezIBRrWJn2jQy19r2zBo8NqIsTLUYw4kZ8AyCRv5AFAP7wsyTSXIeYseOHXp7FUB9uWYrYXJcAq
JuJNw6UkOYViTODuCjQr7u9DioHo7+rlAt9J5h9yuVsMC73oRyw/h3jiKsdc6hSWE8eRbXo601Fa
nuTkJnbSEopdZUNQQ5M=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gYflc5EQMCVYCPfL7sHBYv9w8Zjl+W189Ps5G3dCK2JpiLal2ijtpPdWiP1yEeh2Xg6WRDIlIP7A
eyzmkJG7/CdVshIiQCGEOnh3NPNIUrrNbVgxn5Jh1uqaGwTZy9VoKEDhDGnEZhYbVCce6lcur8nn
XdMuks5l3bFKlONIyOXfVsWHfxzCriWx1hx71cX+kjO9l/hDg+bW671p3eOnkgX+IYemiL4IF8VU
RMg5yTQmN7qmnxnR+muaK2sB3kk8X9wAdnXO2tDEqO6OpqYVF8MFNJqOHHjxsSMFfoJUMXBoDXcb
r1kzWn4QCZQcrSLfTg/XS7BOMU3uYNIgJkDf1A==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iz+cnPhtHl73PDX8fq63Lt9oPyB2kN2ZZBchbrH6AUSue3t7S//RouuXi0CPfWpTXHT2gsy8cd/d
mBxCxCkKc6bEnFyNwdVA2/ghMGMQAs/as9Kc/FWFQCnH8W21OwxR1F1KK3pcYyMLHmELp/iwYTVJ
mGhWH6t8mnc/5y4ci+36SV+07yy4+x3FsGFxgQWvuAvQ5AwuxFlPpxvxuUs82DsmJhGp7Wcs4xnC
v5z0yCJV4zY4WYZ6aUiuwR5cu8JUGsxyO+a451HnpDOFBlvfFX/UwAmTNkkH9ZEF8HnJIhqMLCR0
yVosdDD5IYe69tvPwlnA+scWsxHTUE90Lb4urA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
U3hjRUg72Q/gBHpdi1LE524jJ3ZAZGCJbGs9Aq9bzDmWuNVa7AAqN6TcLQI5azwX00El+Jn/pGPk
IFgiZZpmb7n8/XJI/vXo2uqNIbikhvq0f1XJ+6WP9f4I88xQQKMTYmH1+zOpQu9GSwyAu0vKE3PS
bX3jFiMa8yRoo5y0z8L6E5dwDqZDScQl/bqTqKajjpSgxk6YRmnL8MQ0XyPuOvmMQLEnYFg4cvby
//d+ltRB7rhkZXsUZMwwYr/ueifScKkNfNTT7i3D0kunifshgvdDE2pzSK18Gg1yaLGtNbrPjm0e
D58+0bkRPzHCuer02V0b/JWeqptRmYwK2P1cVg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 967856)
`protect data_block
t4cqgYThih/4ybuC73Vg93ihyicKOQZMreJ4/khBDYAZSjdPLMc03/xpCHoIw1o6bIZAg9823iiF
6LY6o/7nkyzEmXBGnwxJl7KC075xXYKb0vYgNUdqpzl0fAVatul2IchJiHCrU3jEvju+H2T1Gv3t
E/XNepPgTRRFJxCMK4l8A9joBd/PRTvAsPRLmWfMOCcdryYGGE5ifPN4afhxGJidriEvLvbeEIaj
qSw1olj2L0SKm9NXthQdEyI/t/TH83k3zSd2c8Q3DRCfzcz5YbfdhAKd+KN+NGPR2fXqMHWH/OnJ
z6j2Pg+0MyyyahTte+4quj4YATwLmVxf76y2bRJ+++Qbzn5JCajGvXPagclcw+qUneTR2plYgl1A
ZeqxH/HaErLNPakEq1SVCRVI94LqFW+6DtZ4LIsNY/7Mr9hbGuVVyoSiu5VdFIxoZECcvvC3zXhu
HgVPSRqnFKUpoBRTXWe3u/41UuQvnf3OHKzrj09H+9eZ1bnf+ZIbhQE5Pv18gIjf7vir0YyjamD8
blYn3uP4EfYt3wXmrjXUJEiVMyhV4r2W3ST2nQM/oMxoUoygr8d/CURUg0CWqvqOrANVaVIlZQC2
jxXXYoTR9JM7ZGcj1QujLbr8z2sNC1IFSUOzElOVsxMyaydlXnqlzUmwItz0CChpedS65uYCF5vm
MKT6S2HOl/5Wb7XNREc93n3hgr58RE9L61fYK07yJcT4Tn1fTVCqviUvHOMWgUCnMW/+BMa8TDF7
BqmtYmRoIgihlFW42HzNpcGsxZxLvyB2VAFTnZgrq0HODZ8Md56TjNafHD2Cb+0IG99wTplkBbrv
djkHhiA6BuucbpFlJLnMHJ7WNTJqQpjhKYK1E6LeS5F4v6Pwszjfz3MiV7LvZJztgu2otKFPJsEZ
mAgAYLDXfHtUxCOzeDgcteQ6VPuq+J5+gIocsnyfoUoRT1Jn9HZOQJZcdhINl1fZ5gvqaFm8jj99
N6iGZhe07n8G0oQmQYSCM6gTezbIwtAuNSgnabcpp6hOi2c9PzrUwrPJkgkgU9p2OqPAh+wIoYEe
h/pRwGOHuc8VVXWsqy8ThegE1oUXq5d5fMAVcYqxeVcQOg/mnybb6wdnteDqYkfzdPQ4+tUwK2FO
7ocbUh2WLsYafx57WoJX6sBxmakIZKIyY1uURaRvg3zJ3zc7qJi9kLE1WMUPlVbeaJg4XjdcL2Mc
CBS451u3T5vFwvp/JPui6rnbgMDLIoTBZE4Y9nrMjF2Qv5Bwj2IDzlr2h7SJI+tQwLUqUBzmQLYD
uRdVavecPf1T23POZGiAss49ZaWcFB+fpNbSKMHqliEbz622hwiSCQ61fKKJ6Nr9sKq4VZF2N+0O
FW1bgkNY2tk2y70PBEbAFG5CB6V2kcnz+31uAZRygImJaMuHMpnLVyTxYoMaxoZs8hegX51hk3V1
jVHTrwvfIHjdOaRXOPggIJIelcvUlGkoC/ULWUCH56ifIvZ6jCEC088NQw88gzGc1DTkj6bh1WKJ
GwUNJ5g9bElAVPHcpdDnDw8gaxkpg+PV85bxc247NQf5lvZxxodiEFtpWPkFlKbW/8Y8qJyPZWos
j1yzCTidiM3BTa50gu5JqaKZTahgkt/0+U/rSQDONg3mW6SadqLFAJ9SOKpHsUMChi1ESRt3RuIc
BqtbrtbIUwAcUgBjD0vK4Gnc8EdLoLZvcYCx7/bdAEz+dD08Doqrd+Ba9zfGsENTiLxVELtVo0Lm
TXS4u4b3B6Q20AKBXMDC/87LFhvmRo/HvVnrU7ccO+el2oYfGk365Ydahq2UAQzKEHyRCYBjyepV
9RZiU/Evv7mqsG3piEKuytqXGNKjbSZSPhsqpaDrBUFpbNFtvY/mQHyaGfilsiu07Vbwh+Zqa2UH
o8zniAxemdUjSVEHCX2z5owVZf0UTJOVY/9XRgmtw1eGPATvPCMiUjG445ZSTnXiBdPgH7Vwi68E
g1jMZopkZJDagQRUP0J52VdxkpiFgmLQxATRPL92sowvsru8rQzZYpfUctZhxyVeSiz4im+PwYVm
c0ZMl8LIYNmf2K+gRXTSQaH97WTGjGVALFN1++WdZMUBg1kQajkgXAXbFqOYV6C03IYyMrKLEktS
m0arZ9U2DmbmJx7m1JqfMK7qREDHCEZF0M3vM8M424obBL3vwqS9U/McDl1nvEQSlTner5bzEvug
A1aISNyazp9SRA4FXr6N82bAh9s5j5mQpdfsqZI8Nc9xX0zHasiIQwQ/LebD5swIg3smMuP5LWbm
06oH0LRzIvbXVKB6QvpVNMeMsNqHU8nNtd5DnqWKcY0MBTTz4Q5eTWkmeanIf6pF0fHPjxlqvALd
2zVI/h29XqiEezXxU3lvX5MRxX8wA8bI6POcRLCb6YhPI2Qe5qIBj/0Gx2EzBhjpd7SBav1atNpL
KED1sbDobuFU7FPZq2OnyDd66ApWXrZRPBBbUSQENVii5Mkku02/zOk5b7DCJ92A4MpOrT9tsiSZ
fl1ZHerPeQLw7DJv4ax8HzKmo/4G+Q+LmF1NEJ+0ZU8oVmeTQmCmlInGBe2HIDazWU4qEP1iHFtD
Iue80yiwSzYnmcv1L4wpUqvgeRGEm0ldPLcvoUqmyD5gKluQO/A6LW0LdMXUTtXLdymrM1bZ63eR
SyWUlQyWYo96+++2Jfx/lQMa9R2WjJm3hrLqTIqO6uMCe9Z/inx+8RG95+rhAcP32YV+ejwOerpI
TUZJBE7V0x+/+on20FEVwls9n8VO3Q3bTyhMXiblYj5t9zYTMDfJUtiAt+3hV7DJ/MihzUjfK85B
V6VWeLGw5bOCmYjkulltQFVdhWX6DodpM/8tsPF6SnSBhN8oxyIqGjgrpvaPkcYCW+pea+6vkKIi
KtYKK2TNDIROVN/4qQoXjxzW1k5DBSviWFJ1RCRaEIvSerobXdRUIOM3TmxCVxxrmFSNCJXZLPSr
f8vemOIU9GZZLic3i81xwR4udaeOanhzaPsqVBte61NAMWv9OARSBpsoSI9XDy+iocK8h6Xwda4h
Iryqw8eeAm+DAgpbYIsKEuWcUXl2LPtafDF5aH7ffQYiT54d8BsXqyL93Rw0qeqXOIz9rS2kONBY
JBvDzill3hN84qsZ28RlveqKCZwbAxSxa9bBSxueG1o02HvF7OdI4W0nQVZvK6vD/yC4QeY7qm+G
pdxAVdmLB0r0pQ7lmEEe6O4MpDl7axJMYX97pCE+A4pby5JplNUVisPBSAahF2w7yCkDohWCdeVV
wkYFHQutczH7sPg1D8w0LhBXMbdOl3f8CTaXoWTXN8OKJIlwEKjFkzp6OgK2rf9pNNSD+fIU5xiq
vc5/3x0AoqhAy/WPOx334k5D4TTF8ARpJTpS/2FPSaJXELSXwsWjKAeP0AxLqzL7YmQv0fihsTK4
TsaFBh/3Txkq3nR1Rw8UWHHUWBFtNNLnGjl50JRmnOWJafxmcr1eyQxXX1CE3h5eqnGQfaNXw8uS
wnDtQIZ8KTFDsvOVHXUJJaNSacVu8/VpdtH6NcVe1M1ZAIekph1GFfKgKXq/4HE6anEfC+aXWMGL
VqM90x1COEWOoq4YsWUbbTGvclUYG5QWzIVxDGmdHb9W0m39Gg1XL0VNlZTSAvMeFV+n84qFU476
hRvDBBD7vZ9dkg7DURQwTaQPoTDTs0eamEZf0ef/ixjH7klcQa9++lQLlsi2BUiDgpGzRS0fLGtr
rP9kQq1Av5mOO9GDpMhi7SVzbDySxRTUDn4SgDEYZ/07FvnxgOmepQizom004OSoLC8//8i+9QRN
w8Ri4pxCi3xrc3DJjx4AT62hSEYSwwQzRdVPcg3c2AcjG3Y2fZyEc034RwbxC1D/oilg42iupcxf
FTuF6AphzRfN3CBVG798rrRY1SvsRTt7W8upri6BGLLfcDv8O8nRt81UlxjHrobM/S+BaVSWvEky
yjgbmQ6VSRE/x1S1KTIwvJrrtdq7je6oGUc7rOGxWV0K11NEGWBrDPZ/F+X09+PLWW40zxzbjpvD
lqflKt4TvkMTqC2yl7+Nc+48bTp3mPoUOZsZsp9ig72LBu/3aMJThXrkyiHHGzLOa/G0KsZx56sn
ITOIv5vw5XMwUhtLY5gX2y1OOdhuS7abe0LB5u1qc54qqEBVtqrlY5rsLMlimxHDoJ5zJCnOYgTS
+uwpWS7tGKJEW5kIOLwxG+3xZf4Iaw7jJmfordON4csFREJygcYxZL7JkPag3wC9yZY4NPEPsI7n
OzqS5uY0eT+k2vskr4vAaSnYD5u4vcMNdHEdT2W28zrppHmu+u2NlVUNCs4yLZx5ZqP8AhpVU7qe
yOhk/zwebtmnoYjsSwNEWYb168618Amde24gt4uBJwDC0o5zfq4DW/WsSutL2HU2yXEFSlplgwJ8
itd44GdEiFzXKtfhu5sD4HplWp7otLiHLY4DwfR2NvXA9btJBcyDvvz3pG6hW5NMIIgytZ/TnMTj
D3SQ94v/kh+lyX5nMBXkUfwJiF2t8UPSUy5lVl6tp0Ep64i69GqihVWiGWOWxp6YngX2vziQ2zQJ
8Vq/7FIHg8GGErMIF7ZiDWqIVcAXIGy2C+eWY85zkzC2MuiSur6mLoQGgh0uE9s7DG8pTe84Dgt7
30/4O2nVOqtpcctxIP+QWs3FhTEyWMoPaLm0cKucJ9xlESFzcA5lLUjKfVlmotHkBvNN96HStbpB
lJROqb1rmkNx+1OEW9jkVaAQ+/NRta4zbXhFcUjMb2lq3VF++nObZDtFevCXkEfYuv9lnp6F9w4q
vNBK6ilhXB/1lNK1GO0PysXCitqfCMrKgA4iw8FNOclHpG3i+AKJL7TG0HenY0YMnhSaw1nhrXuh
jxRuWxwmU7aJQkrzXfMAkpR/C1RgLaiWHhfVQ5Y8RFRGYXELQAXIy5zDZOtx7fNvMjSat6NEYyLx
yBj0FuK+VCGY8+5ejLdgpk8IbxpNYe2mMMcdkuKNXTX+24t9kDPXOiqMy/4QTrk1bSxkqJj05/5F
70ZijPaqmqp26L/gQs620O1pO+Hp81U4MaD8zSZ37W2xveT3MqJ4hh9GG706ZtAF+JwsHHcgIcFB
61SPZMbf+e3blik8ez4/A88vTxUo2Yp+JZTQgT0THDbjjnaxwKFS7Kp8UFr4yrlvP4T3pKi3540K
ckW8nmcVEaDv8HQbk0XnaVhQnSYYmKGdlmIoTlYqR0zqOpZ89apgbtKthlwDgun75aA/kRtmrq3D
l09xYQ5/2SD/P3MmZFoCNNYY8gFX+4V30MYriPmjKyiSAaPsugvby08oQ8fTvzRC5D4bgQyDNw/s
1GV6rA10fECcmYJh1ddK9riN8l5+cT7Tw8mb8q73evyL4HlsseXHdainWpvPwOn42ZVB/4I5nISW
pMox3mMwYvs6RQiXfOfAXk58Ti/FtU1V4+M/QN/+fBNWqszzChuG+atuUyx/syu9iyEzUnOd2h6N
WMo7g6Sog5LhCZwUiLKmmXIe8vKnQKIXswSkdLC9QZJZgYm07xIMy2AAWntlsy5oEONT/7pnSgZm
RJV1FLHIVcjcR+f3NdaIivgqpJg3JxxCCzv5+lZeJo2aY1xt/NWaBnO8gMhvduncUNS9B60KG+dE
CnUX1BHqZd/hPZ7B2Dlj/LfCsjHWvLeXAPHkdXvDNcQ5DZ1Dbdid2Va/rV0h1QJIHPjAjRTz9Iqs
zxVX+ciamWOc4894TgEhMYp1m+Ppzj/gPELRkshTMQLdWzLNvAa5kiyUJ1+mQYfPfOy6X6eO5KoX
lkVI6I+AYcrGuPEPx2AwmpmUcRrGJszVBsStPWyHOOEiO0UvlAwjuVUM2FT0j0bYRE7OZAUth/sJ
pL955tfQ1dz7IFRLHdaZyUZSmX9D1+SdNOTL5unXKy+1DBTOGgK1jKi7WcIcATXP6TJSZeYcbon4
UsmB5bp7S8TmZUXLvS4SiWy7vR5JQUozS2MSUI42rxdhc4EC6onh93fcBPDKAo7na3IbSuYG6Obd
VvHPjdxwGFECIsRkMFjLhyMwLOZV0uHEQjMOWwtp2rnJbFzOJfON6JylMiJ4zUywsz5d3jCm7ONu
IkN3VzBTZUDlgyKC7HPcyOvEEaoWzwCduvlb84961lomazFYK982Ts8RCbxJr/MVlZLYRytz3u0o
v1HuBiibxTfVDQa+uivlEbTuxlVWAXNaHh18hhVQ0I7m7VOQ+JiVki8qljK40HBvfYGA4QxTmdum
Zz1fCDN8adZ85XiSnk6jo38YEm/WB9VYCLTpCBXQlV7CRX6ZvHVtjCIYa+RlEWnLwFQ1CvzeDbxV
cEyoGDiKYeS6GGygxha1ozmzJciaOnQLwZR7Q4vpnzk2eEYyp6tNufX1vhwXSv+V+uBZh9Bl+TTS
XNet3gjcjln2ySjGhzQqdSRnsMx/WQCrKffhdT/FzbGNmfVlXVS1EO5G2Q3T3kb+nxjaMv1ouymG
8YgXns6or6XnYbhSYNDIynuFbWrkfa2KVCqhtR9/jFXjzpX1AgUOnKKBZgeyc2NNHg9nZhu9qHrO
Sf1MK57y7dYE1IT7qsbS7fdQb5tuIFkaTX+vP5pf9gMehxgFsqWMpUY/cE8HrZBd0S68tcq8Du+/
trfyqKhsekpcWIlf6iGWF6nstY/vaBrpoeD9bfCAbQMk47h+Y0EAhDgy5T5b3ynIfRiItff9Vi/L
l2KnOX14G3fYrrgFSy0J8j8j1nZ5uA4oXzH+QiMBzMMSN6zPO02kqbUAvJ+boUeFAlRgqTcJDHR4
4oKywiG0a+cYKJI5dopxLNC82tYxcBI7z74cfVZFdqpxydPwChsAfaHDdqhJNHtU5qKCbvIHcWdy
FEObTtlg+QZSPgkzw8JsPhgXODfiwIZ5MOfu50BqxAkgzpUqxtcGz1/ud8Etc3dMCGwCp8Kq4Wm5
JhEaBDP9I5MxXRNCb0SxwipKLF9toetqoWBbLe6hAcUXMyOoPOKqzM0WS3Vj1hj5JVHqZOyODtKU
IZxM7nx4aWJk7AZdb7j85FgoNs3vYM22XPik/7JbJZsVhgKoxlsdqK96MlturiWGWa2FUwvrmOfU
xQrPfTl/IwY8gYBE89nIK0OeqH+ySu80yKgD5eLaQdbz4vG1eJK725ET/0huEGiUORimT+0TYHU+
DIJUFiqkuXJ3FQv/DlJkVLzgF+Ds8zMI0uuLnRvp79K+iRZvVkLGpgBl+4an50HE4RBTkHtyYlC6
9sWIIONAbx2a0M25TEpimik9NjoTA9+nFzzoHKA8hO227wdJUsJN2Y6fDQ29MBJFZ6X86Qxjbv2I
W8qGC2hQO++07NXgBID2VsM8muuj2pECUAAjWRXG/AbMCyh1016U97LvhDNXjIOwecyNUwT+bpEM
+x2VcbNxTZqkj7CDMOSPLrocqSpczP8YZTKZPluOCuvcij9idxke8Tc5uRH09NjfV8XhO14DRRpf
o0474SxnOV9TDn0rT3kX6Lyoh9d1iFXg900DQ+vGl8IomyEblJFc2d7Rp8KVVVxzNtq4z/OdcyLi
nK6wFAne1VaxA6xvnW0OJbd+mWyDWDkHNCUTMbpOrChsSzZ1wOt0dQQkulvpGPZVNIR1HBuY9ynR
NnvpjhKjtZfoy9l880A0bVwB5Y3uXsz6esuNj7EQROXIR4mmx694vgsPN0LTQP0YFUV0m4VhH2ae
tQLqV/WCNEDJhKhC6peZMnHcs8Is68j62j6y8L1AUj3U3bS3DYWyHxZglmY2eWVUPyviCMgJUMUo
XJkyKKipPJ7BLoWjpJq3pjj8qi+kplUJXLtQpgpr4WT5R2rb9dLJ2NBqpvUbV+4r/m0j8GW/hjnY
Qdob1I/sgbLVWqsQn68XfPmcPJEM8HtjDtD9TzuHBuaUXV7nU+WulBKke2R/f8AgOth4EsvNFE1h
RRYGHQ7WjB80TF12VCWf2q6KPegqwCazEHNsoGz/MF7VV3juzeDNG6APnMZU2XJDxOLQaZ0SsRRu
l8O14r5u1NatxEBXw2Swcti3cD2MfGVXCjxLh9W/LgaN8ZokohFhFVeJmJD2hf7CfaXKt0wIvSog
HIoeeuc18pZIt/o3tSt5LtnqXg4Ll7DP6vt1rusbQ0g0FTkkGRmeGIPpbuK60YHpekO6rmsw1feF
gwfgW2YUbtro1Q+Y4eDP/YV0NZbecR2QvByQzASeG/qMNLW75ws0vm+TOpT2+9i4+1W7oo7Opors
oJpLaT/UbxZNuzzaXg4VcunpIoJRs8qusfuCxUhHTQhac4HNuue/dsBz7MrtGOiDXvBNj7f1fu47
XhQ6/PEN4M9lfiAFH1sRybLBYLT69OtiiYfMIRBNI771SuUUCACeVNlYfQGZ0LkVACAK5hy/SAzL
M++0TEq/N3olZLq3+u+TMEh/MLh8wUel+p3C9otqxSyCDX9WVMuyHqT7pRKsZ+AYdw9hlsf8qF1B
guBtBfA3niwbGQ1VHi5bFTB0tntVhOHXpzEmSUEc/mwmPxphfYmgOesMuetW1yzJVu3NKEWIOiqX
1GsLk4Qk77WeWft3zrbfVw+1EAkOsNKslkxONJpXfl0FaC3qt/1uC9tctEow4sq15Yrdr1sJPUnU
cbmOoBsyEnUS3dGH44cnDTQJ3VJhMikIoxCfRauGz5aukRgBUTjZyUeb4kBgC10M1ezIrY8nuxkE
2cn55aVxJ4GBChciNfMhuWzGsUdiZxabMTrkpXCq08Ih96zzC/ET06u3aiqQDnuQ5QOeHg4YuhGx
Sf2tUET4JxLvzPnSNZ5drV4OBWMPAuwVjj/b84jBNoKceMUpqj8t5cYQUBxDdc/Vn6xxD0/a2tsw
w3r+pWPQbMP+qOsS39c1ip2tdK5592aJpeTKToCkLZoTbhxaeLT3moseC+NUJPT66o0AT9xsQWKB
cL3hrZ0pbchLj7Q8FfpcfX7dmn8namv+OsgY6vfpkP5OxoSQOU5N6/jsx9uKjO6KTR8e+Mi3j0iG
RfgBQHiTXkKGrNPrFUoQTEwEgs7MSaGuAwyDLQ1D4TeQH63Y5Ri3sZ3dnkhgbg//A30qjt4QxCry
DY5innkwAowc2KmV/3kTReLgpPrzGgQ19LVc01lZpCETFvkqh09YTYL9iwj2/LyKDZHbpNQx1o9F
Zgp8ypllpahE25qdfv/3ox/dARCty+4sMq5p5C9qF2u/2SSF/t0tO8gbq+bQHefMpEV5Hen3HbsF
I0WAsqsfa+dfsYjFMkju+VvMw0L3Chmq7FNMRAnuygANAT+Ek1DTKZrF6E7jZqVL7ug7cVNHUtiL
XhB7Am+AQIfXqTvsi8q1kK26Wb69rr1zXu3atRaNdAXVS+xytKwD/ynOXmOqBeVrr1L5TuR/rcbu
FwJKqlDrEUWfJrIlz9IF/LhYYmMSNFgWFSPVEGAziIJtcY6HvIYVHYGdm/H9BV5LBnBsC0eBggYP
SIb3yK5UoL0W4UaskUE9Yu2JZbVil0h5EG00utu2jsXSa1m+xKQv/g6R51K7u35lwCE5lkT7+FUi
VeQNRvS4Lkq4/cICNKpgcROdQcp5s/APrNLDXbQ5b5xVdIjBhJTsgUSp9ptH8ro2RGLl2Zl6Rm3w
friyG561DO1scHq033kCeTCpxSZ6I09NzYkaxMJH5fq58rNMTzNJNl6Rj3v/+9+HmQhToFqgbDFI
zV+UcDHUQKXGXmnUX80ZVlJrgJZzTRBtPrywWN/suaMXVGSbPbilyNobih8GPbeS1oxhdh81iVkl
JpHXUGWMGkCbJQuS+guzQdv6lfO0xYTMh7MsGhpp/lp+PDD2bXComEaBg1UO/yTuSzgrSSD4RbZM
MViVX9t55I166+NG2Q3wRGespDkvz9E7QvNjEdXyAFbtZIM2KmEctz/cI0PxHLJ2ShtxD/2+gdzx
4imx9/ZD42NYkGwga72Hnb+r0xcroBgMDEFjcYQXLvwoewq5YKx6hrk1paQ0/Iv+/U9NfA/Bj4Kn
Ds10u7snvrSY+XjLI+X4ags1JxQFtOMsnoJuCu2XIFGeeJ06sYB4RSjwsQ6Rdd4iErBzjDl9Hswm
2JQmJMo/RFZkz0ThJVkCIYnbWv5IlLG9lXMNgMTec2Fjah1wkiGqRGV8Ipmh1nM9J+GoN9vaTGq6
S0xJmJyR4EBl4b7FKBcFUcpu/1uNAA8XHxTmeB7qTVHM1nsocRd1/sk5kAl5QqmPl+9sAalUIQG1
K0a2bHdUIxTO/n6iJ5/4Olib9kYrYhGXcTcg75nVvXa947uPjrhEXXRoH9QGtz8afo/M5GoM6DvT
A0qcMFEudURGnTH4Z1KF+6XWRXbS14TQ7sgxMGO3UeUzbIu91NqCm3zXahqw09joXx4KvgREWeqd
MjTFnYtylq38NROaYo/yGD2YT38DNmEwYgrxoVf7HL/mBsqESSD9zlTXAvbhR8j4s098vXiRd7RF
3Ushw8KYWHD3FPtdPDQSkhUSuQRuqJK7g/9WuT6OEidZReDG5Hh4MXTjh/7EQMzbJMKpsIq4H0tu
vTbQZiVaTgPjrpjJlHPKrjw2jrzblX/8O/rPfbTEnAe61/Q4vYfiWPqMt4dTcxs83BqV6QalNDL/
nkcu47CbuKK5CQThcMybnHoRhQ44lNfCDkwsmQkcBas5j7Ysx/Njp+nCXbxIitX6tDRrHn0dUBG8
EuAarbaTT/zFnOL8jRcd3m6msBdQLQC+TmD6orfOGBkevXZXrO5pQuZuW6oFT1uSgAB19zeXZJgm
Sxe4HdvlGTQ0qR26bKnWNynPFifUG4V7zTERzs2QgaxAkRxmeF6BpP7NjSG9VAVNsW7vJ6I0PRT1
UKkiK6auwLE9DCpg319Xlq8x0d+O3v2bK0R4Q2xSWXVxpyJE+1pjxIVbfpeBbppndIHEZF0qdYkw
6rfDWdFXijKo0NmoKWTDlY92SAX8dM4zq+i/fB+XMJGMQQ4x1Op/oN/TODv+SRcv8zFDCOMBZIsV
Rw0uxhBK33T2OT73bWn6ZoIJd/DL2kJtw55mBmmAet/2+Az1tfFeFlWGIdUKF8mdy50c89/neZvR
888qklFnzaOIYm5SbVqLadKDokza6e8ceK/mqT+BjIgOoWFlcXEnDcM9Bvvxqbf8/rM5jVepgUYd
cdBmX9iZU+WZLvKu9zImpzXCwBAFwYUHwj8EhUPPIjTAWTRWfty6gj93Qrmf7HkSGnKf5IwmgbDf
SRGelpC9XK8v/EsiFUIWjD7SvFMBmpbTR+0bixLrQS5wzuXXJqEDd7GHRUwNLLcRziTiay+HxmFY
YAB6NxTD+EcyeR0/T5UEJ1FMEmKtnRHd6xBFWsSwTtyRyhJJql4Bx/LHrB983udI1tA/H4izwRTZ
Wgzw1wLKObdPzmsy1oGiPxdMHJH1ZXuZ1bVjC+ahYlhLdKhzWscRGw4Wzton/FCb1GnC/BwContH
7bSPsXCY3o127VH0K5CetC5ahyhlhexV9yC+Z460fPRsxSm3Z/j/DHoJLsxNs1LgO2lB/e7i4ZjE
PsLzrhR7BVYuESrEs8Om1ryBY3/2NzfvEQab/SkQN/V/VKLZRN9o0c3/MkPMjvVpJtpJOuVxA6XO
/drXDi6OMdy/cVp39XwMtj/C463y6ge7xdjUUPRCLoBqdsNmiIBcp1klHmrGX2tVA4D8NFxgfyjh
dC1Dj/cVY11SvL7QsLb7TIBa0JW8CLBrK/lQJN1QF1n8elkS7JYveBEGnRsT5ZCcpVe/oMNSjIwu
83el891sK9hcjhjqEcfhIkXrqGAoAoGd16iXT3+t4K9IzrhWDAOEZRcsxlCULRvJrKMrYVOcO1UA
xNWqlKomX0gK57JV5gAkH7f8WU6VnfO2MBUrMRlnY3CIO44T5hm3ANqXKBTlcyoV+6kLuFB3fT5T
YV20Db/aCsNI1fHWviqsVCsLyJd1Y8aLQ4MUDV9l5niQfUgaa3PCHrVmjCjdwvmk3mSHpwjX+NZg
y4rrQ9UTeVdAcgA/CllpnsS+rNK6JYoAXf/wBHF4HQhY01wNLcW69IVf3xsKd9q+IWkeUNiqOp+4
fS0E8BTj18Mmo0ZY5nkNPnirFvZZiKws4B8ZKunPin6kqvc57fnXz0DuNSP1evnTsiXJdbToa9WI
2l0sJ23NIMCH2Tnr5z3LrvcIW3CUM+pFKb9TIuge5AMPxXhCQWRXk/qYPNs5WbYguAHM120rUYcO
JJzCKDVc599erTUXFB48wv2qRRvtbwNZZz+WLIHywk259/2pwwm5/d2cug+XbwG5WgQ+2qpzHHMo
aZPMTI+ebLqan+KPWZCDlcd9a2V3+GLg7oEF7MqCZUpwHxe9PYL51JoddibDoxQmHVgO5RlYYdPc
0HyhVistMClgdLARLosYh76s7fHIFE6Hr4sPnSq7ZpMoTpEgN4Hqna64Mp6RViibNcB9lZPVgmOm
3bva8N1js1s3J1WV0jV53Mz977FDrsJJ50OlPIAlsUjJQ5/lLIWhLaGwS2/woTGA1rckN+7Jg9w/
gK2DU0LvE2bH0mG8NRg9eEF38U/yS7ylTUxO9n8GMUahgsQBgN0oNcHQYmCzySZNrZd2lf/C+pfs
NvQAg9hwG73wyJ05FY7Y9KujklZkgr8LnRhMoJ2EVJhddaYf6UhozrUG9eDSLZgvNMt2T/3Fc00/
qTYBm7SJnrj2l+MUmS78liQgCjWv8k4o4GnTNTs+bVBwFWH52rQykr/r9upNWj70+tfUSMADH+iB
xWNHoJogfchOR+WTcza5jXTKEfpguQ2GOyIjWvCGMwedcKAk/cjSaKfcJZTAzWhFnSqqpHLlLtjW
NGyMXdkQUwPSIp6OZbZYfoDyYX0H/kemiGpjy/wGwcRXquSy/tehz6wWDwuJZvg54PamKLXQmTkm
8tpmIO74YZcIA/3qh8q97VzC6hzyH/kw22M9I1s1ysMCXur/AoZl1ryAgVAdl8lHFLrVhR1Um8tg
joGv0cYumW17kxo7Z0PbcFe0pY1vw2pKerV/RG+tzJnyBH9Ynxb3RLANz+ValXftjwCk6jgOJZcl
44Dvf6BRMN5MLwL77KDzN8HWauUX9A1dfBHeYpyGVdGXNaYubDdt/d/vsKPJBllKgL4U/Cxgh3Tt
VGav/qwQ6YK2YGEZWjQ8ABlxGiHOtMfFHWmmai/er+fIW5y6PkqXslvyGiFjXGPZE392Fg3/neCk
u8zeWv+JwBz3W3IEDsmSs/vGRto0FhI/O7RcvPPLNIPnNDnpZkq/k2+Dhj0HlxOazxiZr8DijDTO
Op7YhOVGIWSE2DR75iC80mMl6+pWnrqPkxzdhbaqGcOiYAVJmC/dGYPMsaCDE9cendi8zGVw9swO
ocob7+xb/ZmPECvt64LGCjlV7cPBXPtzoHEg/DXxMDmBL3drwCXeST6A+swDNYSc90wQtwsoE9Sm
8i/aC83C2pu6/zCrRot8VIEe59fQTyI9JjF99fBM2tVKX7mQchX/2Df4gDYVpNtEQQXbeQRTrceU
QQAptDeh9uxbwQQ+n1QNtCoqGGXPmBsADwEI5McTh47T/jWjFgkA/4rtStgqsxGcalyesDjEisLE
HCYVZvOx2vBZzQTRhgx4T84yLIVlwVeAEh9V9ZbeCqP/Z6NNrAqvhVV+rg1GPLpy+OqIhCasDc1Y
oBt+El2ormh9jVbZUAEgeT+dEbF0d1OWgworspCZzwvauB/gmQFVo+3pHG+WAwUXi0jY219N/472
xU020s187a9U774MPBSPiKOrCJPSYpK/jUa5k4tMskUlh90Eod9iVuLJ+B61gI/JpqwjGUEVYM2g
qd2xCJV+nK4gIseWTWU5//Ere02n1COpfInCcSzHQZcjNvZ/Zk4DSlbVBjeM68PjFL7YZ7XRmQDl
BtAyiEDvGhoUCiXMzUU/vVNuffMW+TteD7tmbOCt9FWd5uC6j4d+Wjkct+/dUr2sB2MSGfg3lkLw
dnWRF/4KxgknpjB3WnSHTe6oDCPM4LEvXNlAWN4U/xfCkGLm9yOx3O3K7qtAI4lc6vdLh4zi3M8v
vHA51IAIFNHDqZsrCXr84TAT6MTXupIW5jUx0qmLQ1CTFjtHluwPM2iWis89WoPU/8czZxoLCOJ8
er3aSLgIngje5QMz6kW2Z8vynjfkzaSBQi5vdvOrU362HZStP5Co/Hsd0r6XFcpHvtHOMBtnxZMG
oBTzWDSxHrFTIa5y0hXrwNJriiz3f3KOKEfZ11nyqTM1Xn9fpPtd8f1lx/wNLJmxwo3azgSW2cKp
cuk5xWsV3kRBYfMpIXJRyiwemwCwZfn81eJl+pjgAAa3XPf/BAQ5k5p9raJ9Gn4nCc7XOCHpjpRB
woPOsxWQdYyD4YWnmbPJfvPZ0V+Vumsh07MXELMvz5sPytt+ga7AsewSIiOyviCiy3gz9Dao5EOV
pVefL5c+XkAAxPLXQB6UFf5IQ45CaISJR35Sa+vFiyNTIIDbFDYsZsUy74uqKa1AIQn9Hkis+4wY
GjlBX0+lIt/y9fef0QYEpRu+FnjtGxwjpY7S0A81fihNv4OCdO9pWsnnI2FkUNyEQOy4Q40GekP7
+uwKh6ZTEJ3/qb32vm3DIw/o2MBhhgnpASVqNkjnRmzXaiy9bRkCu9+iC9IQQRKF6bhYP9IuihU2
gnMEIaHZP46jfDrHMbmwURHL99EkzdT3ROMuz72loNqpmHCshQozo1qb/9sbR4TONxfPoTgPYIua
bCveIdV+Kimo4wTTgfTeiraw82cRpasKsO4aUkpjfxMZyoWr++k1KzNxYRluwDJYTelN+687P2YY
ofmYnktBaPP8+YoSMglfiay1Nk2rQUKL3ZMsFMBJiPiNAQO1pWbpxys9Q1ckD8yxXKnC/FOh/gy6
4C5NQKj0DUWGLgIP8zhyIvoEsH8mRNi9UzdXBS9tmnhRshoVDnIu2CZuBTPRhzWFqMd0qKeJA0+c
JGwZJCyLzoJKmyUv66i7GQeyDoNGom0FAbKO7ZM/RO3Uoo1WSIZnqXbcmrdNI/tCrL60x2latdnx
rfyZyiEvyjQ2YN3DXbJHYoYyja19BzwQlGQz3hEbF7h4Rxryf1qW7YT4vAW9+dHxZOrr43JwjiXT
5KTPPfviAKf7Oh9/VSi9PJbdqBIPu+z0MN1G1w0+UBHxJm/U0Fi8JNuPWl2iGzXRzZcSTov1OZLv
GKs4Enb3T2pLiBUv+kZOFEnIZFqBr627Zt8NfSF7ByT4cNl9Xxkeq4/cGObaGmWcvmvIcMiqK9F8
u3TTkgCzQZpkxzdlp2sq2I1CnOgN8mLCfnZmFZUN8wO27/pMaxWZz3LYa+cINsZB+IrcDd/pPQLT
qztDv4tZWooVuXMKRmJQtUJw7HQfcD+OUtG0ASNmx52R/m5GFDqN/zpZfqWmNNIleTzJPfQ7j6Gq
X80LdKrr9wsIHqg2Q9aq2Nmn9dwiMYjpCTmKB1H0uiPTQ2GYSTj62Q/CW94URvxiCcgIw/Wc74RH
DeaWRxN2GuYqxv1JGZ6oE+inEYeIsyoSRL5k5XD6UZak8u65BwPdOr9hlJRvNTJEzNzFDsRgAsxE
8te6nU/ZBBR1jtINaipib0A3TZKjghm8NEw/9PAtv7rdoAw75+3eTeINTJJSx8oJddBY3/A0xdsF
XNyTfKolwHJ6LSYekK+UY110nCb6ZqLZ6YNT2osG1NK7F8+MJOwRMqsA6rQmjfZ+MRRlFK04DSiD
JdZWdAnWoxnHRSXQwyVt/QfVJtrhrH5J9s6e8I8NLdDoBYt4kOY5sxogH07dpQW77jyBizH6DSRK
LGy5gaBpgEUOoLsxWiMIYOhi9Snvh2gIAW80l9MO553JhsPA3Jn1qJGyr9/cOUc7PyhVvF2kLZ95
kLxmChK/uLHbu16HtbbEDzvUFWql1c9MUDgqxSNijNlHWtwWcPVEDrL2NFSiZ1b9AUeDeHJQ9H5C
TH9evTFoIMbUzkajCaETZBcz9KhcP+PQQgxY0J3vKU1yIhXwgroB4lM0RmRMhIyuJlJzECbaS99H
U7LNAkOAyoju6KxD5U207JAqxqjpod6gDpBFgKz4+N4/00DlOwKKpY0jfvMcNCqFJi0hlNQr6pPt
ZgEjldAc0lJCNh8EYx+iLvAGHsPAQ3rLP4ejiVL76qUVtB7kOUIINyt5sz4DsiShydH0wh+g3JxB
HTcohhxf+lzOZb1N0pn3QPPjitHJ5dMWgeq2AELIvioN6UUnhH1R6q2ik1qGV0yk9nbLJdhX97cF
TKkDzYBaSOCioyOCAf/YmiNArES/qVON+aHaFqkmFECcj4SyyEQE20XX0AtsNNFGAIW9QQBTaKiU
vGUuuPZlcpdlVRA9NiY5E24xghpIEZRwrCoZndWqpbdph0Sbitq+JDkmpbXl2LGXVB+noqsOdQWn
DHxiVUGN3iMHJiZWvvewEKjltWuK30yPGpmfJEX4cVBr1DTvokmubdgK3xuV3yYSjihAQcUHe5Nk
Hn8VMhWfm4p/2AaJqQuDZ8g/at89SUerf4GD4+HtTt/dh7OiSg8p0sEIQQioSA5rOB6BzvF6kvA7
pgl2kup15hyttJ1eokxO9RnDLY/tcWJA2AwlTpeXPmZ2kXTFA7/ZJnI1Klo8H6aVFBk/QF6n4S9n
ZNYFnpLqsy2jhG0Ptdaq7W0Cmd+R/gHnrT+NmxrUSW/faXfskRPPzswpkk54kjiQn7eRhh1EOtsx
cO2iEpz1Okn5LXyLgeEvk2P24sW8BC2qvYIlM8QG65JxjvUYUS+8DygNTBLTccYUbRiciw1wIgpX
1VezHkR+JuAy17ncKkQxJlnO1d1NV6aj9NVQKJs0xYpNp43mzV1sK+Y8omz2xeyq21Mpg8wT0uI+
eeZ7H55hF71FZb4bhA8bAs4yUF73shwc4UwFrBgmvKTfMijWQn+RgjLQv6EnUbwdn4z/2OaVZ/o8
qzr0nFJdAVuJdZlJ5rr0YR76Nhjq7WWNAMQNGs7FXTGTcsJuxZp4uk/jdJyRGQtcXBpq3AqYVw2M
7qOZKmZG7hexmAp8KFAE2FQ6EJ6L68Qv2KVSegwtA4Ql6Fo0JjyRkZxiuJYgv5mpHcPzDoK0bts3
ynzEK1NqB+Y7KkHmRdNUwCWyJt17z1wlXzhWZtxdoWpj2wjfuMr+puLwSUuEoCfCrqaM6Ap8ijs0
n5+2xBi6HkWJd6EoK7Q/HpbHH6XFfv+54QS88ussTdlP3fM6tbpB69YJ/tEH3GPNY78tkV6lMkAO
rFGNITgg5wCvH7QJmdPEsozmRGVFD3BiIUE+XV11euBvlI4vpiROTIeMVBa6U4m/+AqFc17v53yY
xz4wFZcRbCr3x6+iSVb4nJJWQ9c4H2p8kpvC3qwOVFDoocFs2V6jAihk0tyw/ACH/jxlp2S8WzqZ
zysHIGPgectUWZ4fG0sDQzJhlbvYUErT2LwFAVLSgqMcOC/nGgGE0WG0fKs+R3EQrnoVTcdV0vkV
nejh420Tti0pumduMDh3hkBj4qIhKt9b77W1tgQJ/l7aMHMeVMzt2tvPYupmiYryUDP7ug5RDbWs
wKNBSMBy5zKWCYqAnxDwUnJM/EC6kOiSAwQGjlfV3EMLZOvxuFpR8EcMo3Zf+FzmX9C2ADtpRDjz
BOryV6HnjR9a8LtgRDxLUsJkCdnzLdUM5i9UdRKAB06Wdl+9qrh8aF+zGVf+jw/oybTscgItlPDP
eRn3rokTljAswKGVtrTsUADEfVpomM783IzqoHDzLmKIDxZMov8lzdbx6D0J8KIeYTcfowCPfbJf
kDgVBq477nSkewLzjB8nsYlDv0cLcAg2PGyXS8OYyVxcGp9ZD6A9bXUgb5xk07qiJduWP7ZVYwbn
sEH9Pk2uErIyJ85AbIy/DVcQ2uDBUTYynQ9mA3OTUksHiMtyy/f3UoeY/psSFrL8rha9dXuZz1Ph
d9W/Oik1C5YqFloCjBIle0Wdrl6Xo3f3S3pUmD1fvnx3S1UniTHfeKqlZjWQDm3KxV2g13eW79jS
ZJlKSEPuxdZpRTd5gTn3AXXwHRtS0w0lWXKgE8Z7Zet0vg/SOJZQ4X2HkknXgDFtoNLCkV9cjHTT
NpxBb+ihdQTiXoZiQFijTbUk6K8HpHK78sRg7E9keHsw5Vh1ZwJuNS4AesJItc1HrI31Jl7vuxfR
Ky/hVFF+5A0JNm4R2owoWwH6eh01kZeXe5yE+Rj2zOyA0JYatpAYpbsp4Xik0/TQF9ajRecjJbm2
qbmTcOiP8ll/kEuI5p4TAncTB6iR8au7I08jKlt2ghhMwvx+cEVHyvK/XS1gBiN6UtImbDf3QrGr
PNcnz3wBkmsp36ft3xOTqjgrzdOzi7rUX1NTCDXmH2RGftLChJTLcb0n13sumO/sVIqoi9sCk8Gw
XKqTxMiUgLuozT1NuR5o6m8ox+/B/wz9bamhsixkD+qEZC7m/FKJDQXLKHmBXxeiXc0ifVKuvyD/
16tv0sQ/ONxCnXGGalH6uiZTp4jvLv7pUovC310nAaXHZi+eEzQwdbUfETvMTG5t24vjqCeeT3AX
7Xhy3Q1ieLBmm1onErN6WJbpcsUq7dr8CTXgxSzkvjT+WSHghPOAoTPKXkEL2SGP4vm1FunByBIv
P9m63JIb8EFG3EO9zL12exdNlulkauxsfc4UHR3R7Wth9ULCZQnttKk6TDjKFjWtkKPEw+9nyFu/
TWmnuTy6oJB5+4IdAXtOyaLO0ref767uvnlNQG7yFbD0h6nTvc4OVb3KgYNNr4lJ2+JsKXjn6Au+
8trQc4AWpyuoIOIX7J2fpswQLW5fuA6WByMzHLAd30NkVT6KDyZ+odiDQDjVfDHQUP32pWg1qQQ1
4EuAnxj/IphHK3JpfzBwYvjSiIbr/LlXrGzTDA1h/gkSmPA36vlAEUz1WupNk9UZjF5+pgWjqQVR
GGW3NETm9f7lydeSCB4a3IXg/aLruFsUvBCh7VOk7yvKnuHju/B3vek43Ei5htlkdpezXuK/2jSG
GuJkt7RaIGlWohx8lhfUoJNOOhUiGUasQu2IOWC24GxQ4XAaZ+LUaGMs3VdQK/pmuCqkC+x4Kz7t
/N336RMfsSPVMtjRg/CJSg2TKnMQSoM150X66XaNlBg9AKP+25Drhn73rg1YV4hPhB0zn+z7VfEf
o0i32+nW7MlH6EWlWNEudywW/5ZEVK8iB1C278/iPdCeb2mzlg7SnE4wxLcvp+m+XfpXmpCpFcSV
9BiG9I+ifm4dJAx2nzh5RM5EKbTcRKUpVZ8u4XBW61rTr5XCjSDxWfO4Duv94L7fAn4vhEIkp4xX
nb/InwBfXVL12OupAT5ltfCpA2ZFpXhKjTgs8+HX23ts1Bhzq5HhOVp+Zn9Xon8U8xob39FB1UX7
j/fpNk/pVcDk+yMm55Hs3UE0sY5Q7eHPlmOPdOSShsEZJT/6ygfRyQWy+sJ3x0oE9gRwu61qUsUa
Bt4/K98rfJRqh4SCT7QujEJDMNGvGNdzpGRDE7OZoOVDpLz+BhsrlRRkPCaiUAfE22cRlQAPEadx
eHy/INfve6Du4cs70t8NWY8s+xQQC0IzY5TzasMuw4ci4dwarBQ3Xino0Zldbsl7fL7T9k2hVOq/
SCdhAkjkalcmh8APtLaGZeKGRMB7v9FJC7d9q0V2cZeL9NDylElYg2Z97tf4y70HH3AoXEQQ3kNr
cuhYT4xWktCmJaOmAzoUTNE4WanR2XnNBEFchgxrlolOo1fDlztPEyXqKF2D3Te/HtsOp6y0QJmH
bq4jlWtkPJM+nHEdfv8aX0/BmWQErdUaEm4OiqlcWvvEmVjw8tqma5cICBthXQCNaMARvAr/bhlX
xiPmgSNiDCkTtMp/wtFJEB2RUmXxI/BQPTi7VpkUQZfDgwwKwhJttA6/FYwJWvZEbz/p7gAGWLHd
JImCFvWi1sW4bU12keKusydLbcezWvuBf26pAvQ8t6mwLxp6i9shnQnby0DHe0W0TgKosjFjwKgX
9T3E7e41INz5QYTi8TWL2S+G9J/2NqTmq3CGFQyfqFbAOgXcAQxYZQBMDwODP8+jpvp+HsiQ7j4P
DSmHey+61a1qLw7ro43c3csgn411/dT8529YWPxG0/0tE3/UkPD5KSvXp5QZo8lL8SvxYY4ZADKc
ExO/z4191WNGetUC9uA9aHFeHw0PG7RqRaf3OzCkjx/4Gzwo3rTQ55ZptqiwK4/IIv4cHs/yLOdW
r9KPOjVZd8GkL2xonBTGAKYl51LcXsGHhZY/5GCVE/T6J9mRU1/vnZrcHk8l+hGAyUPppSjgWOrP
a6uKe8WucKhQG2J5QUvYtXINuRWueS5tpN5h85+AsA1gUsIu1e+UD1eKJ7VFKtA4R+H5x/f85lwv
v/7u+yYzQMRJq8lLKOrBYdqAj6X9g+gq3icDyV40z8EdGp2PxDIkg5lUEBcglU1ni0JDMvQFCG1U
+Z7hajn6sBHD1k5X/A1UZY9RXm7hfpU1gSUDSUXpPn2y6WsW9DOAVvv8+cyaz93vwT3/2gxsc7KO
+UeLzxlXC3qMzP2xV6hLyPXv9wpuEL6smBsyFLLBl4QLymDzxwy0hFHNNpwdhFelovXVOOvlxQDB
lYz9xp7EeBXHPtKHG035/apJcMbE6mhrkwNILAOee+vKlyA74B0qlk7FTWA338bpXmM5cDheC7Hs
lZZsrEeYlM5NFTxxKUejonpInrSMGhT9iIOeM0nwHFgIkJQPowdzJ4kpjI/jyeHxpq4LzhA+ngt1
OJfa4MmTNdAddyCfGlQ4f2LyFSY+DuOwNKrqJQ7S2ssVSFE6b08otHjLWIt6+F7VVihXgaSam3kB
0PMZbzEHJkOg/l/3e7YJt853R4eeIvOny21b3yIgk56ITx/eHc4qaw+l0Fsl6g71EYjECnC3HN/i
74d2SftlHHQs3me6jIXQpPdux54+9chVO1WRlLNxPy7R1geGYNk7gcpgtcjjiQKJCSJsJi17pDOA
W0My7oUgMWQ08F1zDePgrU7pgRR2z7g/eZAKjv5YCYlZKAxac9PKAdfi7p7pfuVKyrxoIB0W9UT+
qj1IRAJBmcL/Iq5km9QUFHTbDgxNfkuTzseAZ7Z+WV6DRiV7M02NJw4HsUj13n13EG++j6FuHIh1
hp6vRH0L3AmHQvalOgyou2oViRUjgtTci+TJeE880EYgKOXRrpOzvBXVlpia75+Vkr1s4kp3c4i/
u3apxnhzLy7sRjGbiNEIRJ2M0BRmWruKGea7oYhNusBOXVgTOGoZPInmG2qKmV2XK/ieK6YlzoK4
ieqfZLkzDOVEd+HwJHk2ja2MwfSmlFayf6iIOxePyy35SZRAqkWruNz34BUNuU04AtdUw0Q6qOk2
Ia7r8eOwqulmSthCwNF4o2uKqYpHiZxD9T7YT3XJVKHmm8IGvZdRuH2Zw97S4rGI8Gg/zVEokL+T
87xAOEp6fLy42LG1TbTggWfQGHQRq2jB33gtJencpRWcueCf0cgm8XviCCQ6SkNOlXwQmANXs5TP
z2i47r/puSF2HMpHwMqd5ExnvG2lGpW1e9U2rNgXqZU/HXPic7rGHrNgOv4lqeOHwwpGbu55HD21
ITHfwSAmVgW47rmwgfgSLIrmTPtvbkK4eQMEWSRpxGrY5mB7a02BOogx4ntjTW+uGsVbycXOQT+u
5gFSlQtSCDSbLN03l12+0n0EU/NSILWhkWk9Tojs4IW8Q7+03P97l5rd0Ggr/YjuSaliyKaGIzA3
lT6Sgr8QMMdWemykbxywYl5u6QS540c5/48jUqx+y+Ys3a3Oq8W1V1yyJLn6UEzaytDqJFi+Grqp
wkda0X5Eee61aZwnG1iesMhIQ2quJ9dWnw6JxUjF5XHL0g2DnPx4gGmdNiBV/Ci6vquWFd5FonHv
qX4QS/CzaC2FKNgmY9cKeH20WSuet6pewDGmv6Rer78rD73g97Y3/G8XxRQe57xhthhOhLygJ8n4
olYrxaQegYgs+8Wsb/QQgXQ9TjKObk0ZfIyWPq0G2IvictBucjAT3LWh/i64snNnntpGrFDuDFa7
WyOwmWWC+TToNzWrFpr0xK1JYzW6cNHHq31QhOMo+8JL3oETXcKgkK9tB0Xj7FkSLJMsm0YS1Fkt
SB4iuvnBfsCy1QZzXyLXoTfZdI8zLJXIImOgiAtuNWjHw3iykXW5NrqT4x8RgW1yjhB5+HS5x2Ak
2/tQatrV8b4LrV1bXkBE7GsirZMsgiyYSWh/FPSTMvOYbTkUxa+MNy+u/nmz/IakJMwCCaa6pGuR
tm2UDCIKZ8JMEw/mTbPGJZYAJ8/fHLYIJ+zmAxtjwllsckL0mZ0UlBozL+AexudrbU3x4xQTiYe9
QjhxjemtQokh/4/MUAJSPcm6LbYCT7R2GADRjEVrckI94pzWShH1t/BatfLK+e34gsizZu2CXhGU
g94K2710sOyjg6iARWyXNeqQpoLYZkSJuakM2zdpOdtCpoNJsb3SGy7UNylbdBuk5KjKxIgSpnUE
OTuLW9/7oMdj4+2K3Ha1elZzfVRqZGvWcC5ia4n6U+aLUjyjH+WaZ7wXoXpF3Il4qL3rBhTUFtC5
sJMdX05UGZgYiUK7B37fi4DRLZ0q6UZZH1Ya67nCLFTOlvLhAgJ0I9iUot+cBNvjzP1ZNM1WNa8m
MsjRubz1ejqUzcNtZzrAZ7mgzg4f/jmg69vsnPwPXzolZAF2QLaN19U524+FfyNkgZWtIM1cXR64
tS2eGq02er1Su3U5NE31Cr8PW9lAmuqPQk9FI2dPu7tc5+t9CmtevXGNtYoHXuioMx04KPiAgfrI
8ZFUTC0HVnXt+vQS6uo/DISrhJAeJJ7MFExbF6rmN0VbYfyMcCYuP/IVdP6tJPWRXpM86P0WrJ0F
Eh+xCwdI4oCqOk2sQcD2AiUHqZ8gA9HqQj+E1nKGkF+TSBOkwhpdADjnbThHNkyVNHbfteN4AG0B
g2X2nWC6ODhXy6nxkUWvQH8xBFu9pCiL49UEj0eru4GEroTxJEiEx+HN9fm3BkPApvl2flLf74Gd
E1P8CVZgwPNpnJQbSlB6zFrsVrpMCYlhbrAo3qVxo9lwUjdCrghAZE+UMZ0nkqiHMG9gE9Weulu8
oSVZ/+3lHbrWq0wVTyRKwGy2gzkVzoMy3KlQwEeOxfwPyVwc56g+o/uaFVUFF/BwklnYA8XM8cBC
JKpQbufFFW05Uj0HHYu1DqlNVh7FBGf3G2nUu7YfLYHgaAN6bIBbmcmf0TOVuitCM0Ufa5/I6Ari
VBSvMKB38CmDSI0WJPBd7Fp3nK3uMZTJRHTcbIoI3dVdCxtLtEoqGmnFo0Ef7ygbGjwCyMkAPuAQ
UojMQZO0pMeM7vOL1krhH4Rm94FsjaQGLlm5GT9DZ1nkQZOQd00pHwGUDWZO5eoUU+LYLaQv+7Fk
l5jvX6ny7YVhXFx/ayTCA8EzVaBQNDC+8//rOMVqpcn4TIbhpimY9QPu4egqJCyjML5Wsuh8yYrs
5UgGUV9ZJS+aekZVA31tQUPk4Y4mbiDoKJ50BUpdyQ0Q+5Qi5Li7QvEg6CaMZip5HIaC2xxUtheG
JA6oRsLatbWboLsWCCDXC+XEG5/ypcEhflFC3jSLaTR+hRw+yJV7mqfGThzE4hkmpT2xUWIL3b3J
VQoBSKXas6giPZluNvZWe5kOYMmxBPBnSirP+Chp87v02BflixgDYRqu2bUCXe1uZvZAYmij2h+C
U5OLUIjG5heF7lhBGONbZvcBWDrZiLx227+5qmIOmrbZIuZVpG+JKbkWB+s76omlVwVNioZKgbji
KOMaa7OjkxZUzLREJFL7pREaxt+inL1oJ50lkGIUG5MiDujKNS+N1CHJgwlk4WFikyErOcDyNUxw
toshHyx86OLcgrOzXy40OqehU7Usb1MWG1Re8WCLq6bc6glgTN0LxYdEMXV4MwbftKNkMPCu5XOk
h3SQZUzgPJuaujnnU0avMGXTPULMQYk6QUm5f5W7k3IjQ1A4YYvERThAx51+N/MCyR+bre0D6OX1
pPBehVhkIdQywAeV9bEiJJlTnrUe7TjTYct8IMGFE6AC7oIWKHnJ0vSOxk4a6RkC6IfQuz+qftQJ
OcxALRdwLQVYwIAxarBJC+qM6OpCVtXUJTHER32Xmldmb5Qsqe3/XJtGKaziGXJDv8N1A9/X3+hd
ejp1ycQbnAtQ3RHWOjY2fDEZNBWGS1hEZ87edHSl5GkaehtGEtUXPlfXHEfdEA2J2Zea7YDVS/0h
c+3UBYSygRcUlDrjDf9cTm28FnBCGixuarUlOVNpBz+rXTz/S6Xr5hjyQytycISEcNvGevk7qQ+3
M5gij8z3gSwPgjMHFyPQJyYGaij+qqLn1eJrNT4nDXNqGzJVlqmqHpjMo/34DnEr3Y0Jwer78TgA
J2RXsSTHiobHE11PCimRuXDxoCE2iHg2Vl2h1dBEUZSIspHrT8TOjbSkcWU8k4xe1Nh+npzFq0JR
lL4PYheJ/Uje4xIDyVUvKKYzBjthoNrEvtA1lRQYoKJfCxEX2yOdsIOufI0Aat5hCxAQgHMC/NNa
Sp2a23X5JnXtHfM4aWD7ldSvN6PBKRea+RO13q86rrnz29cU3LcnhDEm8T7MZbZ8yizwbk1TphgJ
ByEQXTak3jbT5cUaOpDRt48P92ueEMNJj9/foTq6nVt3S7Gr50nCIfA4vBmvzh8Wtqt0MgNg0k+5
BSRlZw2OHuaV05pQRvRe2bY8jqv6ZqEAXym7BYDCR8ZmiFWA/qFip1KRhqvHOWNaJQMUmtW/1Zj1
nLSI4sdTheqawwMTriIJCadvd4JBuKNc4fp9EOEC2ljzygfg266HfvMl0D5f2f0245l3aPuphS1y
XicESLz4IsNbhfUVFb8o1DCG5/v2NXqA++2Uocz8h1+RRuCGKfF4Hfr9S4ChZvNt3k3l91B3RTEd
ZRq5aqvoeLh1FhGXaPrMUl1PRPvrFKNwg+Gt1AKRtfMt51F2noldv2EonDef/URMZq4+D5syd8oe
17sBVKupSM/V/GUZp55U8XY/UIyUXS+IF3AXAnFvhToZus4nax+Y7HA1A2Hqn+UteYJOqd3teGBX
58esJYCqsxpbXGBbl3XvriNozk9HUShAo2arbnCP6qaGn4ZTM2MGa0VTcU4Ts4D7d7wH6CB3/RH6
fC5VQ3MtkuPukpob2Vs3QgmL8Koj65cLTyyYS9XFC107Fm2FW8N6trRefO3H6bwa06m2oUNbZiJQ
JaLN4FA4zvfBIUvT6DuObfnADfMsMM7CjmIOO1wLgWirMo71KRiQQQGFsxE3juq4cUtvEjktvRR2
ZKAmzh2DnKu8Edw5s4Xlox6yT1PXJrm5s9JsF8Nt/vVuERD0hxHyYzTrsAfh79f5WqgyiZm9Gdj1
w99ufgZ8HtqT1vHMbwpbQ+0O4QxfIingiHvErSHNTVN0Orfy+ZCmIc7/ZQo1LpWwnG8RbpWBATOf
cW3xOG/MouSn9WKwgbViDvZnyHzYAZ/w2po1GBkwsFcaBuTfW7KEITPJo5DljB/frb2YoEfj9HdO
4aKezkdt4UiVodwpAwFVGRHkbwVGpwsqynm3JG6iH6JUwhgeM3bW1OY0vURgMsZOCid9q1hqgCpj
hB3n32GblogxCqm/5ld5M23W1srwy/ygp/A5ZS3aUG60Nf3d0OJfJvRXOOO1dfW2XkqUfObMxx/c
JHQ+zvy/DqG9FHPiFjc87tcVVZ1PHRZJ58nVXxU6Zm/LiEtCr/d5N/K92jiCTNaik7Hbe+ATXAHY
4IxucVHZw3RFYvhCX1aaOxOltiKfquvQvXVLHZHC/yHWN5aWGHdwwlFdD2g5+5T5bNJQqN7qEsMR
pcbUku9vdQ1N58yP8n/S0LlYepb8tjk6JNzhqgsjPokd4LaCPyb5YeXK2Dv9DiSfrzqGyIp0vG2W
3H182Itk6G1O43nPmc1u2ubGYKr40+2xSmw3upwkLsvcihBKhGxsrT6uNwZwS/i7QEqzsQtkVxvE
7h8N8pOoSkF1MFhuvVdbT0fLv4+U32ySFMHsJa8URROjVRjQ0zQl04Gqz926CBoDBUtDDiekdZQC
3g2W1spdPGa9p8s+hvL5NhhBXUB6kxAVD5pAUXQF+TErGLg3/2+ZiwsClDyd8QQUdPB3k2Pf4glE
ZfV5/DhIYeia4SBX4cegtTfLYsGrXJ9mCpX8Nz0DkeqlIrqJegV9wAR5gYXzWp72vEWSBWylH3Sg
M6G41v9uAiRk3tAJLfni10DHhe+wvqUzSH7sbJHecjMEEyqLR89ka1SpjirNfL5AmCe8h5dtHLH5
Zl4zC6JNo/ZtH/FMGcQuj32MS6ny0o6co+lhyupR821OP8jy3Q99HOOScwbRPTJNT3sBYkRcQfpI
b4NsjC7kzaQfsRVQCagL7VVSSc0JVN0vajx4S3djATrVfgJ4Sj6R07ImzJCc1YEw5LvlzrHyKew8
eHHFf1TSzcvuSgqcfA3eD6DXE+iaYYvEQMF6WdNGI1TIJ3SeJQNnhy8hTzeEvto0ZegfWG06t+G9
++CcmzY4hhRMX2okpZOGNyICHrO8DB39kgmWhIMDe2vVcrnjKy709eQDZqzVCi3Cf8SiB0rlDqbX
Oz99Lq3betpJnjR3W6UDTfaQTv/59Y0By88mhYgaa2tM/DcFnSz66oIWUK312m58lmd7XbCtzGBt
Vvs7ijhZctLrAa6PgBpoKgNquTBPU+/A/KNPVC2LGySY6xpQCoMgsEL30VlaCJ49bn1P5RiCf6Sz
481lCYZazif9OgUxvZtQXpatPa4j/dLxoVJN8axA7YunzxI34qlhjaWO3bkNNTnBaP77b58HylVF
GMfth0hSBXbdOrVqqvwExH4WqYcK1keahWKbffnyZsJQ2sDdIIcIjcngwiDAwYr0+QAdz4c8Nr9z
U/LAJbK+IqN0FaBs8mEtoFlTnioXHYfgJV+OJDKzqJhiSkNk9b0zom6z6/SCnjWkbkB/V6Vatup5
r3dfyrwUI+zHRuz/0+FZtfQRRzAuSzs7BZ+FaDII0mofMCmhMGmPiELNma8+qGM47nngKc6tZMV0
ivI8Gd+l0qrtq8n8m8YWxQ82K4/UlaBycD1ENaJPtm0u6H1xzu1DmciRduPl0wG68eDaR3Gx/F5Q
NqSEMScYQHUKVPXPojuI5nazIoj6RfyVTpQSmpIHMqA9N2JAlsTL+cLA0p8XU7viq1Pi0msClAPF
BIcBrw3VmTh3ijJScooixDXedKdc0DedkTsnrEycCV6jBqnUuqQN9pPj8s/Nf1MLaq0mGO4Nn3w6
n1cke2y/2XObj09bOmUWRvlNL+FetahatDn0rJQHrA5hMVfARngm731dMYqHfB0upOBT2DpR936U
hLvpiwH1JRUezQV2dAo9cqqGq3xQJRGChva7eiRwgTVhWiy3PSUA0yHVN3T8nUL5sWCN6SqeZMDu
tpk5V94yXc9SPE4lVHs42xZlhEDD0lpxy7GVwVtYCt00Isc/nb/CLOV38PBWTzVlVaWc6QYMyuzK
7jsmpwYlHqWCeCkceC8kQCwijOB3QKX01pe09F9cHsKsxPxY8Ww/+xWY2JvsT3GGGVyV2hJgmfWi
rhMX0pJLK+n7WNCgGqrYicAT0NmekAOrEmput8QMO6xRy21mEHvPqjBNiAbBjfUDZqEucWqTYp2Q
x6ssnNxHfnzfPSp2x1DlR1cW8AemiVEHOGSuIHVN5S+jmhSWXeMZYKVh5ZxoD2NvMMohGHvMjS3y
p07Wr8/qeSmbkkKFruI9v7lHQRwd8L7vGywfGWQJ1t8ZbZFHPiAl8s/gNWyjHafFSDrVDOEE2dTY
t4o57W0eT6U1Coh76DYB8p2JsOK2Gx8KlbQU2iOv4qRa7ayZyyUUr5AwQMvY7KX36nQ+jhuk60eQ
H4VwnZ9xL6I0zC+dg++QH2S+3ttcTWgkkVWXqjC74LqFJAUrtVza0j6eEU9a8FCxGO+Hm0K/s7K1
1yhbZmuoLWKr2mtsjc5HZKStNFDPuCmzqvLUC+fOuzWhzCEDbWI5HTnbknI7GvQJIciof6cG4YcV
PN5JJhBsKAbRS3KeYqBLXg9OF4mePKMf6sIvZFKqkI7haWEO7IyJ3xGvxWE9IEqTYpb26lZHcTku
1Tum8uL2RVB6sRqal+VAffCOzMGV6XC/JkjseisXY0C5fbxd/i7CupDqzHgMXUEg76Etf7Yo5ygF
zSK2knG6LRYgN/G8i6qs+1Pk3o4dlCK5aoMs3gZmu9qlt4MWxh16kGo83WTxkLZetrmYGL+fR44N
IrGlkQJPRTR1+24z/IOxr6Od4mt2H8tajAAHZcGXv/MDbRrEnfI2Qc83kCmAxZ5RqSceIoMLEjJ2
G3JmyZ7FOhKRuXr87wvKWRU71G27q+qojiPvijB5JYFmmJjB4ZkajnG0axXoEupytcWlmShXx/oW
eVn09G4xcQ+OGUzG9yVUD+mlLsr0r7uUZMJrDwIRxHNnSAT3sXDZVqBq1BwE6YzvZ4fceqr/+7ch
5zc6WxCD/o8KzSrhixpyT8MpjOntKL883DukwK6n+sg5pSEBtGgCD3lYSsUqO0QGCE5EQSm4Q7LT
hyrl68vaF3ZZxJW3BMgspchIQURbSc/Avn+GNz8UPISv4tpneQ2Jq334nGkyxbt7WPn1MDGMHP2P
CPRk/7Udq+jC9iJpdxYvwlmHIDKYmscAVsK6fzMybEuG2SQ1b3JDpo+2WloFq5c3iXo+6gGVvZdf
bInPijW2OZpCEZyO91jAMuoV/MHx7l740iOXVv7HDbsyNDmSDLPqNWURdryuTk3TZexiaCi3FJWD
oeguuGbLQSITV7Noebu+uRHlQu6sux+hU+/Y2V53HpkXoHMGcDTQ0mi69yDv+RRlwlYf1g/0dAnk
057Ch19U1doXTULY29t8f7bEk8Mu20tWv481EC0NT+ACJZEcJT/qeD3FuBHHin39U8dk7gsL8yl6
Hu+bexHGadY6C159SNDf2tWkt/VDd6NMgcDY7faxbxAKFxAd6NOwhA3Gkk3a4FhhpdRQB4ihr8nP
hp0vSNd9iR+BitJ3RDGGH/txTHZM8IlbLFEZ/CXVZmPFt5yTmAxxxOq2WodP0a8fn9orn2K8Vul7
YZ5lT1r3bOWrYJY6lOTRSA9lyy5OQuW25PUEJzNTnZ6K+nMa+hJRGuMcfWokE175FO3eBdupG0VT
h+MJ+LGJlQmDfmyK9OoNY2pHMCnlmPSR0SrzP/RZNeGO5iPdKAJgHX6PivxpBIpwmhK6dGy7fgZZ
loqqpq8RU2lyiCNJ4/nD6L1LGHYqR9A2hcqWqw9b4ZFoODmxXWr5LYsj8s2MXvSJhs95lxS1AWBI
Izvrx9Ed98JOfkatRBO6hlARdxUf3J+VNGWXWiiL54edBIxZfyx+muu3Lb8UeMySthsZw+g1zL+U
eUREBmDiLQ6QNSCNTB1/pntIShVdSktP7Q+LePYoy4Tc8mNxP+FaS2RbLClm53gPPmYRyS4MWthw
E2L8YxLg24QssuqIAY8Id3mGFbcuru5LRQeN8DpRzMZQDZmDCOaSwDSHCPJChhyaszLxFgGiDEWf
oqnB0ARZ9x8TQU+FZhkX08cxXOFTlrBh72+s8baTlxGBbilMASNu1vr5YkQVMb7FX0PD5VvoYueh
RiF/U2CSL1F9C2bFQWt+rLh/YrXr+/EfA1kKvtZJzi+7Ojasr7OktXvd2J6TOAFPbrE3sDkVOdae
OhUB1u7OFg3h5XxQs3WQDVNZi7e/pqu0Ss2OkB0JUsnBQ+rqIDI+H4r12l+bYZ+8SwTEgyMMoqFB
7MQkFH6COfEmokGo38B/Y8pmslP/VldV3ncuXVEqnt68W5J6OPy10uGYdwsTGEu4Ltuf5Ly7RO9H
KE2JnR6cXCCPE2bxSQj89IjSnTPCTxopziTskV+jkxsgSfwamoTv6CDa8+fxOsWMKKJvjS0h+ro6
LFU4DdiAdVDGgrRie6QkVFtX39QvYcbNr4O8zxXQFJ2Rl80LjV7uKMZqM9nLYlz8BWjXmOkYuULw
/lU2yl0mX0i/0FMDJcatb2Xj2hDbvU/M9fg4sVj/5c/d/BIYKOpt9ViIbtTfQeTfz4qh87B/yhDB
Ei8ZLKJNADaoHz957ooGkC8cI1eK6JnM6Cxks90Y1tgAW+da8c3cWNLgnYypbpkICe8ySVD1YeGx
aaGtbJGX6sfsj4tqHVu2tL60C9jXPsAmfWPvg8/VuWRblutMiyudmEuY9kcaVaVvctsqYJ7OAk5p
XLoiY+U644nvbjN64hDIuc7LRygZ28Ys/5AL9Jbsw+YiWpD4+3bFjaY+UqliutuXRV3tk/NUbIy7
gPQld4K4v7WJD1gx5BXO0U+PONNL25LZOm0Yh4p7EYHhev3DpdRwRZ/AVSq9bQltsB3za3krkVsE
NiALENb56+ZMiPIAkjNFeZPSAnbaWdEmvI4zNRIJpZ18pqguwGYjk5F7rMbwEpJjjYC+hFXqPUui
5QU241g0p1adXjArEe4jDSII/XyahigW12kHkJJHEvVEtBu2Bu5JgoBMUh/CSebv2JKvDPBvcu4v
4kF3fVSK0lw6mYxp6dcGpZ9aGIjUJ2JkNNgJh+GhYRjWMt0zwwNJV3BvuXo62zN8UWAzDn2/Ray1
i2l0W+mcxljmDmJ0cWdHO3fsAjYjDgFdDD86aEd1G2JSekSCn0TOfa+98KLgI696j+0x5wmYdM2Y
fSATZhcQmtaQjUFRFnHiBF5p5OysOZbO+3gyXVOJY7SQRbnP524QEdl8vvz82LsJU5WGnHsOzeeK
hr6TV6tUP0E3Rm1hiApRAWwoTS/LfSBX90C0OWKQlvDRRU6Dops+v3VzudOXQcURUrLxCc3fXi+h
EXpxKuRzW9o2LtA32xwhYkbCXp4dnAX5hxlRynk2UQicqUg1f+biiLe0hUWg7IbwvlbkdqBvhslg
71eVlNsotOGZiQuszlg6cUev7opcqSGe1/f2DiHiTFExzM2f52Z/RS80lrhAyYGrQvBtRUMkHL/o
NJsRLXG6W456wcxRuqHpc//VwMB7NDEtZAT9GhLMWw8lg+DJwEy8+9iQAawBB0ooKQbWjD4DePpi
lA0T4DOkNerkpTu0gti32r7wjB1JQryKZlGi+jLm5Q5gcjDOM3PdLpE1jERG7oX6NrhOUcWkLcTd
nbHZQurFRki+WZ0XQZhjCN8WxWsOoiUwWHUh1NlcBN1Az4acQMfSTR2v0bPqmnCkSTMbfdwJVEuv
7llzhPrVB/kdMWGqIN99bk1MN5NjXnJvJOwYzeeNnfYxkcaAEBItmdsAfwG/Y72n3IuIG8PnuJRY
qpRsnSUIZiLwm01DE/nLXY70ci84wH79RN8qFUHs2GNVzqrPHNEAjrbIbNXxjO6TswyO8+gz8sCS
ACsEdFbtYZofgD2rqMZMUMkvUbUl6GwvWOkgqG7s2Cjf2GEwZ2RnKOGb+ycS0wjiJr2Hgx36BH3F
WLtyqilDu4LfOjIaj/DDlDrOe6Pwc7dVdUr4v77F5lOhIPXwINLJOqLXQxmdOHMY4ckESi5B11PJ
RAqVV2yY0RVYt7WCLVx5ofNvU0/dT5p4loUcuAlFNKIYa9pGzqOLDnb1uDqN6G003uV9gcj+LCKG
859WYARTofjCBi6S80ISsbW7PFofTz+dORyv/fdZUscEVeNZz+2HaoTV2IYw7RqkvXOVXNFB7mOr
9xalILgA3LcdxT75mgBy6oP4qGxKDGDsBuB47YHl/ZImg2np1SZKF+t1VCX87ZNrSQTvOb1hcAK1
mreZnbChWL/JzHLwD0dNbcoG/j/e9ZexQ3KjxgQOiyKqUA/aiwHCg1vlyLEd/X3YPH5CKQP1ZLkX
qi0vlC4HrsKUbnvm9MTjKZdNBy2rKBqym1fCZWOELiLv+xJhie4BvoAB0xCYC0KqbHLOnh1LaOb3
6gyS/eWeOyfZO6UOxNR286939r2AOlznQiwrNDpgI5KRy+0O3yVo8KeK/5DUmwqnKxe8obvO/bL6
8VcVytaQYvoKEdHK3OLXg0z2H1J8XKQu/GB65qnxnJ5/w9DcbWe5rYGavzGXHtD7+wF/hrOQ59q3
sg0Buvs25dhIofRz4O14M4qjvLfe495XzGvzwjUcBCK9FerxwFo7Zqcsw7fMslNdxwTamDPOc4Kf
KGrbXZn8hgeBfsQj8828yl3ved3s/w79wyFLQ464KCJFNBQ0/ZjuIJ/HmICFspg95edsniLwfZqm
tNCkmMqy+PSvBXoyF6OM48zzt+W+DyxJp5kcoLDlPf0+R54vQWbl3+VMtKGzUfGPaevsfLOVyKLl
3JQIyZvI6pqa8ZIdK3oepxOm/cat2eNwGgn++wIuZlKFsRiKCCKC4FiqCJ4wfNEypUSixIwmYjx1
OzBoEsPXx+gUkAI48MBxZxU4fC1qzfaGylaeQEDsP5wrihdTfLcNsdw7O8O0Ob9OLM2wb1AdENyR
p1w6M4CQ5o7CGyvvSWXvoqxCvV1Ijx+FNsw77rUoJSEQviV4a5xR5EkRwSUXGAVKfdy4Tm1ESHaf
aOGBMaoPennTQRR8geuakJTVVhleHeF/cC7pzetyzAawnPkCb3zDTSZgUS1HjhKqC8i7MvO4bS0j
MxoS1i+ehcO5eVQs/pxToU9dKXg1EYvWBeCygEJmSl3Ay9Lp/M1NwMv/o6KXA5U8eGq0fkJT5aS8
8uKxl2CwduO4g9QgDnptf08Xh6T22nTTX40rLagvReQ3kRQkquAPC/YMtfq4R4T7u7rFX1EwDkTY
e829QOqqolRWDpMKk2eR+g2zNa3jIAg+nEbay3l7InEvxwrPRujUPIqj7cZSnGitA/vjGwbC+giS
pL558K0JFGv5EYqTQCJs3mwZ4HTszAhjrdxRl64deRVZLSC2AyhVwgZr1t633cVnqVZPD0mSVqcG
YghjPNxT7DS9Ula2RGpi03iD4ZHjBfhhmq48vvLoeOAIzQ1eAeReORbEdZaPp/4JeXsRTLoVnsVZ
d1y3s1LhKPwNuPbDGx113kYbBb4pVm6WB+ZbNNSOOdGq8f2fCR4Kf91mCjM3ADGPvBym++yA703Z
hxeePexKXiS8cJAQcLDO/xM1RefvcuR5jFdVHeuPwnXPcUNMHcff42fwp0ATQBFhfioetWvVzoqe
5CQHfcfKNak/FR2sBpjlxrDwQSEjgm3x4uA3Mz9CDH4AJXSesV938tblKxOxGqlER6HwzL9f+DPB
TmPJzyG0Iv2QLXQRG5s1LGw5wsHsrCUfuouJ01m0KeuTuoRirMSzyq4TUKFDDPMQCylZXFU0dZTg
p5+UTwPPEu/XpXQGmDP7dIFW7lmy+DwQ2JEpLw4v8u3tmFcqdGDv9J0Z93tXC30hjBp984tjocWe
MiWgWHHbiBNSn1iLDLPlEcUsy9mcpdpAEGvK6aEC5TRv4pM54a6BDoUlx3WyhqbqL32C9/OIVrlZ
jW9pQduJLQ0tSTbtheoKDq4Q7Edt29wwae28wYb3d0oPs+w2otS9ajn8FtQXd9T2ZZ9hKyBy+371
jZFxgdAl2PKpl8FNjhFlI8IYpBI/218hdHiRXE4nxRiDzWQzfaCUqdPnEN5ALN/IJ18AM2FsFxkK
d1zbHD2zgu5/mcU5DRFDv6bv4Ofz6sED3XwiTy8oYxP55+px+PaeL7PYV5T8WgCbcXzQwsHkcqoP
p25JTOTSnkmVe1IFvYeG5gd/ILIdQDiZ771gRpmRpd5HAy6pglBaz4ZWI8m2vGxujx3i8HcZEtBW
xhAQhsYliE+jys35IH8ofhZTRWXbaIm9qhKlqF9ju6ACddnf4ua2s5RyuG3Pn5wap5Kaw7xjqrnc
G78zK143MwTz/rKgHknb/3MNlReer7IIKopRInKZpf0s/QPjex+pJEO6M5M/2PQZaG6g3gVagKq0
RTsh0DJXwlqYCi9oD8nY+5v1whLSCQ8DmkbvuEwNbpXj141l+00QAo7MoskJQmdougut5R/+XeKI
3+0HIEIdV70iJRvMcBSv04ljH6O7CVAOZGl54SqiHbOnDB1Y4KKVcucQEwPDfUfveEkvE8yOtIHw
yxACIWW6G7XDe0A/H9v1EbKCw7SW/5O2+D1Tt9sNuA0gw/rfbGOWtYm+NiCsSs1FboPE5jRwP6x6
x4SWA/H6JypC1w7aXy2xrMUV96C2D/KffXmGDKCVHcYQQc2ejp553ZqW3NDfSfvO1WedTO3Mfrn5
jTuvjr73LLcDcQfZVrZ587DedO9JqTWSQK3v+CiEjaZSMEPOHH9Hs35MWoatrLiNHPsj1DKXGWXm
/FYdZnCkNsRa8ygbiAEfdh4IAOyzY1W/GpfWUTy42yn2x8em0sSiY1IcEjd2+DTNFihmyVeJFGK6
TGgZSeN0mq2FuCj6AjDXbEsrZgQiPQPwdAWZOEEqagJCM0GtxKLHwGPcmuZCdQTDCg06z/eRj8zN
/KDaKYPI/5G2BHlf1zYJDfmgCaDcJK8WEwKOXqgVs0A6WCIwRmzTmdAjloZILMS8rsQPGlZgbmXF
kLdoQOc/RI81oXlK+LNTscI8WoIv95/snlTltEIWWnVG1A7TvIpBkovwMyv+hR/G9SNbVxv+b3Xs
x94Ka9JHfKhxFGffcHyXQYhxQZiA8JUdZwsIBpguxjE906lAgnLDrjgTLHmVeSdjjYKr5nMKQThv
QsuECaoQ9ZBj2Wgs4g8M9ewavDam8Z2r/BdW/xz5lMywHflBMHLjMf36AJKNZaDAvSDekAMLldjg
8Q6V5+LPWDG4CfIeXyrp2rXQ2ocl1Y9AoN0KxTKZwksd92GX60Vn6x/BocGMr1iaD2DshDY1nnw1
N0nYB4b0z2Wry7OBEKnTOHOclY4OHXI9G7qQSIaLTboLoCNwEvY/GYX0XdlYmjeGjOFf0ZMj+2pH
SoAW0U2wndjXj5r11DGPdm0VVPQw83t6qEWJXlVDRFoMr8sWPVATO25kNORhSRHO38hyg2dhgWNl
7mdvKiQPaysH3eJYcgHC4mS6B0ehTtBNUoS5tEl4PlVKju16fhmrV6J41gSn4hKDRSGOoEmZJa3g
2Co/LatInOabkOTvR39b8wXBk8tMoyK1HNPJ2FmoFiuduEF+icGd/lz+TBh7HHgCx25ela4TqHh3
8SnsBorM4cV4IK7CO1KRaKYaefnej+Q3cI8TRfZzOc/fWyzxglEw344MaCC9WA1oA7z6uNZwLO4Z
mXQNdby7AXmRDMOuHUpD1xg/smaH8zEhR7rrLpXUzJgG4r1FQScpW/FbN/sDKyqzceef1eAOvP1k
p8jTofkOVJgJe/yg+zSNjKxvf1ozayOYIeKK3S6dhLFukREbZkIJxpXcF1EIo3hgoh697UOzj0Og
9EBPVzRnkWLD4ITvKTDA7UHRHXAo/7LrBm/VVWjIzbwnhJ+T0UxNHtMeLyLBi7qNItBSBRHr/njK
ms7KwAyp/itq8joME2yI/E6p8blRb8ffDayO7PF1yGW7Puptjr6Dm4kGx9sfwbQAr6l7os3NCwj3
RbbVsv7BABGBaJqn9OQnkj/rJ0BDHxM9GjIaih1xGcBctUVqzAHeJ9TyAUbZ4eyW+v3FHs1jL6QB
LK59wpzhFM6PFhZy1JPHm3h0ivPNdJVAUBOENwmQdjv+aOTVdYrAxyD9BaG38mbFy0xfr3UiN91U
wRW5F1by7feBKR2OgI9XaPbOOU9FsmLhx3pvvNWjxdEVIluYX7GdJBXEyhE/LeQQYn9lG0DT6WQy
DRe1SGswLH10ntthULuQdfjVygypkkqdF8AWTyAJ7zeBbuiYWK8l/4K7QzVj7QBT1NBFPgNDVKAc
tYhF0PP5rPENYuUVzd0Sa72tCaw9w5IpRh3jYAgEpHOdi/45c1OF/Ps8eGJ8TqbyXl5pMB8ISXfj
3dp0FEP4H+zlVgK/yeyxLQ12+ti212U5pl9H+8RaQfTRfZeoTxGbNnHCj/uYt08dXiYUaVPLhH4N
jLCvZH67JT6PDobzb/KwdrWmAb5IyrNniT5V+QlQ3p4PiGQxIWOjPN6noYKV3t0sBHFYLmiAfWQ0
U/10mR++i3TeqEDREZkaK8DfBXAe/ASIo4NLUdWp61+hYJrnkLoOtMRdyUgLRZxS83bFcBZTyDu1
GSCDUTacdimxh8KiwK/qFzFOCDLYArtuwuoBZXry55+ipenf8Y6BotGoMDek31Efjfq0IaWXSWZF
1oWSttXQnE6LlE+kclf8bEMlsfHluU6Vsg2xhkJQ7A7h+A/pPoppF+7nijucptE2J1mdoHzCTTyd
OaaGB9nImF1g15PHlFY7BdXucfOKoupUC0h1iMfvWvdytfpy8YwwtFNiIM+m7Ypf8Ds6vYSB24pV
c5JgbQoA9ZTR1dFsPcpx1wnQ3RiAkBdxVJ40I6gMKXJ8TrcHHDv5Wsbqnx/zt89YA4YgKt6wYrD+
tzfNNA/yhAOjd4V1rappxRX71dry36uzPgz96HT8ppsFk85K1IgoxpNoBPz9nV25EReiHzRPLuYk
TrEBDZZJN4W76ieqJmxRIYaa0hVdJvPbM4VjzSDAZOJ/fDF0YT/n5DdiCNkT2xyqSu2uYvj9D2/5
gk86R4st85TW0nwD1VRbs/AOc8e4qMiLu9VH3BMcpys0giHhfN9OuEAINZu6ValCbTWS2Bv1IgVt
jG0+AymP45l3kv9TEoyanh0LBu8ZnUJhihlVVZ1bsbMwmTOzfoGeXZ+1sKB/DgE6MyAy/BmGIhOj
SzizKFKYXri0GCGTLxx8AsESQ9PknYqfXdjp/EgQ1+K4t+72AsuEslYZgmW/AGxqxOwNPgbPlOGt
BaWtFKhaTaS5opTYCWag81B7aUdh6Qljq8yAcje+7o5kq7TagVvImO//dOIrqFBUvy08P+8n/lSe
k60WBAU6riEoed6+PMi/SfWh8QxHcSDLcBuGe+f5Ru1LX3ejr+dljlGB5cG8Q0C3LfteAEo/VALx
GdTSkTHyqBMaB1/NCo7q3vuHKI2fRGCgIZ5+gDzEXDM2+oeaeUmN1I7wLjhAkxkwAiazbxCmHW8c
Ka1h/CW5u+VmXUnlXEcwMF+ZZQqiCT5xXXkTkD/XSvCckXF0tRsUlxQFwvbYjqNiIS5la+87Lz1Y
9dEYzp192nExBCKzPzr4KsCPhlmnEokWPiEadseP1Mgpn9MnfZO4vuOTNudJMAskfnibMZHp+K9T
2DB+SMH14bDPjR918lvS3GfxnQ4znErCNe7qqLZMwSmmCVgktv3qAvY2p1osPdgHzdL9WyNRMEE1
Y/VQYJe69kTvD2EFD0q9f1LP6fRd23nf/rLn1fA9yzjeGcqvBShuZZehu9POSPAaoJ8mEQ1+WRpA
QM9FN8MtFZOYojqJATjJpAhePklrlY18cNqYkCNY1OmGKV2jMwGtPJspWIk8RexH+4Fcq6Yj1Shv
YGxOFjabaey5fHS+zK1AkLahgBdKzNrM8LmEpI3PsYVJl/u0dyI9IdrQF3e7TKa2lFRJcFv41aTD
1S8lOvTLUvSL8N1ZGHUeY8dtnkX6CfFRSsCgsicI3AMlZ7VgUWMWTkQXT0JS6I8tR79/m6+gWT0k
RJbqoQz211s4zwkt+jJEAbyc/R5wlrAgfZSpHnrl5+aM2e10TrHYDCTA5dq6prn73TE3jtDTI/7u
OWlihG2iBN7u2l52baXXteFZ9ycKbwsUpJuGqWFmZRGLqDNRWCUt0ff2Luk1vUw0jBV0sqef1XO/
JGdmlrlLpzBbNG/vGLILNPyYLz82brbcAkVFHyju7zyYr9dUkOiw2Y1QYjSQlWG97sgLIjHUmyVo
CvUoPq9HEN6/eRIpjNALAbJSUamasgESoKjyVpR6+7Bpr0gqSL+Qay6/t6TeUlytLmhpCgFopWLc
AtBR7ZOoeFHu2UU79SO3bF4m1ohfpC1mC8SgDpOfoMVHjaZKJ57xUQxUKa0J5SlfO+0mSJv9Mhzr
N/f48mLepwpDKbP8z3cj6qnrdv9jiJpWqW8icfAxOPXSWoHPLSp5HQ326OTvcYi7lKnjMKipdXtA
TbjCkYRPaa+GDmT5g3EeDPfCep5UnSIxbMKkgt0IlbP2cdKuL0fNL+hJt8yL28Alm8koFT6fssd1
tvTaJXBKJIg6KNAbWGmyTOfSp71denkOxdqganVhRPXsG8kvSsHug+6+13K/Uqwgv6YvgfOJb6JW
Lo9f956PoEY/dB5WbsoXBsJ8WiE3h7LSIh+8vCxrFKPCKp1tdtR/TAEUjDwUCO0ZFGbkDwUNqbZR
1zFLCykxRmn8n/CljlckZVNzu4yOypWqDFCgDV+oK8SzgLnT67PEU4Dw+/+M9JIB6aFU7gIVhVaN
rn83FkPNxi0f0hmdtZye6QUMUSPF8o31Q9i7M7drSrdQl+vWsBa5axgkIfzDCDsvQrGhfVpJohqB
EAhsG5MnRYeEa2jbI7UkCzbkTGcomH/2ac5ZAbPZFBcDvc6jPGGVMm5OEXXErwSDPCnLnUbzOBNQ
R1IAS5IxeHtWN/HT/DfeXERj4O9zLR9PgkRlOHFoZKqvA7J8gzHCUU1wz6chL0DpSHPRouXE4EM7
qNQJiduDN5XSQzcnxcZomS6fk3py4hbG13SFLE7tPi3zJoe5rzzGCAyAdTz8nAxBrawKeyEVHANg
UMnG3nhX/vvAWLD007cacUzLs0G89uXHL+1qcyx3iLqx4Pk04CBG7Av3QPHWBr6iEN28J0QIZ3x5
0WuMg3zU29n0SgMKEIpodMY14E96XleN/vm1GlgLqyxOqTTCmLtmkwk0gYi+JQXqmp9k+9kpJvaq
YrGzoeYnlaxdLik7PreiBYNSDV2TBltMAYGJorsoSJExCgRDanZFSnJPBLIT+pDnmG4fMw/IwUxh
W8xzYENdTPGC2sGgzg+IrjGbmP+rU6QPuQgtuH9qnNvONkElbCEYm46XT+gfcQIMUvDua78ug2GQ
L0QsFO4wjRFzhSPpMegEmlj05JwHzc1F8xpEgIvIXjk6SJRxSHQf1PVnGEwXJcHTKt26f84vg87c
Gfx5jzwkUoN+VgueX/KcONaK5MBips5AMdaEDtyz8J1IXS53Kx5QTIuAvASvKEm75Wtmo+62TxOj
R1+Lt8ym+i0Or0GIwMz370FAGRVMnoKj5AyzrLS2mjUdgzyoZHG/24tiz7RpBV6XFlsa96W8yabH
5Dx2vD+8H2vBCC0d55AzlFmT6xbAn6JySajYlm2bOPHyCC0l5nDqozUNbL2yNPXt8iZjiAkdoBqm
qxAfNZw14ANTcGqtoC+oSBoG+EDYsKoaEfN7jJ9ZroB/fOi+sszx2Bm4CEQKb8C3XQElA4MFqpdw
2YaWqmlEWHn38tRPG1XE/BA8qV9LeScDYPgwvIClb8JhqyqS0w5sFyG2LA5X0SVVEvaNVAPxQ4TR
abW0OYco7XKhbChnv5Cotpme87tf310dCQ/h7GtzvTn4vyM3IfLFFpYc7pIQimzNgKHy8uny9Dew
13jCArOsfn/flVXPCwz0hsDQPiKi1tqtj1onI7JQCdRnl8Jg1xK5/1uTR3TJpYOclN184YEBIqnW
gr6c4RaoGGwoEn8kF9UA/vaoj28af7XiUtAbAEF2GQfgszhFDp/JUC6lHX7F1YwE03Lse8pakq6f
MU3Y/CZxKOUp8/o4csrP3pRlkJ0YSn6T424aQH62Rl5GPKOHUwKPk+pmuwBUQ7R2TpLNae2+cLv5
/bGFZBd1qwwI99oTgdJm+nwRF1i3mhIhBE+em9T48oJ7mcfRHedYJnqH6MwcXZdrmywh5axU462X
EZ9PH7txQJ4rClLm85qD7yaR700kd+loC4zFM76MWnipaEMMc9iJlpQthIqxGj+enQ0gZa6grIWh
TRR2aVKlf7L0IaHEIub/Sl5OOPBIyJBiDHRy+qtoEV+rWdH7RLHahSPsKsxzlwI3lJ4UF61IHpy/
E/Y908+VmzuLtWhuJEkWPiFC0ferhU9ZvnJ++zdE5V+pK3eB91sFFVijaDtLe3ZQuZsK3tpUaTR8
8fxtjP3qVGkIdWCXM1F7mQbzx6xSxcd6ysnQqPXOVallxrwOn81p+bI8PevYH33Qqn06pGl1Podn
fKnUlbEIxvFxFsRnVXRO4FJAlorV2eyMGq2j8WnJa2dD85Wx6WXkiVXIuwrworcOiOKsG1ZgYjKe
UCCHcpwUJaTCifm0hLFbOY8FH5zC4YEvYq4hw93KQv72mDk88dJYPSsJ3L4BIW4/errnQxtcta5i
svZuG3axsOYxbohmrbkMr56blA/u68ZqRNtvIB3fWJ1K5fVPfjm3h4G67KwC2sJJrwq4IayAiqp3
0tuH5CQLALb5BbsqdmOY0IjfVGUf+FtAmRAlrS4P1DZxupQ513PhZ+5rLAeh64VXeEceCIwti7ON
Tl4YCCUaWh/RlOdB0juaHyJVPNZtzEzqA2NhlricAImx1KK8CXayurjbpjfVwraFRSn70Ji/JCfY
7Rdxo8yJQugutjb30abAca3dC1UDeJvrojwvW/AxtITrSbXi2XIKWd/gyYcihRN704bHl0sSoirV
AljmiDxE/2cFnQr7uygUyaEDutMtug/CWs/lMcL+9l9FuE8VlZ31tzTFVupKusz4WMhbiQBAKVc8
h1MW4CpAsdqLpmb0PUm9XeNiUtCMM9mtAPqDhz6aLdgbk2C4ZBvgis4HQ/F0dd/o3WU1iwZgmxxW
/nrLwLLYWmjwTC47j11cpjozI+NN8AWRzXnUZuI0v2sS6w96qCYcDgc/wTZz5xe6JsqKLeJm86Wl
SW2/7mCEieDhXoDNwi3nOF+3Tsnbrej+yb9Q7Ng0ssBzo8n6wEp7C7A7BUHsudSFYlcq3UV7Lfao
CuhZ6KzhPj11xmhOTMyTuNTfD2TLeBV5wnHlEzlQODqNt4ucBBgUE1Q5dYrEhMYKBPDPi2kpHILW
LaXrp9dczWq7sT9kdGqdvfEqqT8JUBVM+jEjbcOLEbkSJkMBuThnwE5koq1n+k7j/mFHx55bvzHH
/UcFmL0Jr6mqoy2FUob3pQBvj7ndnz7l+dp3Klm71DAYI6+nigjSJ+1bD65KYM0xX4QSaK4g01qV
Lr0DgS75aIXTXrpWnlZGAfk2iKQAMuP/Vig9FBVk8QKXOl/X7vXKZ51399GxXtKFsLz/NZmMDa8/
EKsjqjH0voRaxYiloZYN19pz6hakws6Sd9K7Jyhw5+XA9b6poXxLCLANg7jHYyrd7klxh3DSMPCC
GeBT6P+eo5SzQlBMob2WeGaRKKOz89uQvDCoKssH9pNaNlckWeh19tllzLJmR3Ccqufg69+wsiE4
/h4bfQpe73mwSxBhiC/+8+1qoiB4blzc1D86UEjOA8AUZdwZgGm/iSCjCk2a77j3q6zI9WWcLKm+
HS9xl4Z2xS6Uo4hFytMzWoyIcUCUOWdfVo/QjNF+ntbQbOu40bhD334pJIDkFpZLE6OX/NxK8TC8
uXSAVOOTQb1YurvkoooFarD/a/gi6fZ31hk4W2YA2a18yhcoz57zy1NtPjo3anUO6HU1POQqYdcf
EIw0+He3sfHzKLb2dIxpe1/VtAzetS9r34rrl5QiBLBKw0oiIC4h591370RJ/Iv8WCLbAgaZaE7A
9ALnBnYIG4XiZbqYymgonwPNw7f8qLnbIv9+zLpWxwjbt2Oqm8+MpOrrDVBTjaCUJrMqWYrwuGRb
9+vxmr5yUP6gaOYSlgqOaSn7Z7b/WyWoiiTTps340gcmo3XsJKbah7eI1Zejfp0zYy3LmpkDgYPS
Ir7MxUEtNPDxbuT7aEFI/TlIp+HIF0MQbUrXMHMqzmUooiLMfFi1cfYlUSAE2hXrf9p9wYTJrmqs
HWXtjamGQAPUK9pyUmN9+gXAiy43C1Q1vIRCiujYzYUJ8LKOug9CzC55aa6p3jnX/YO4LsNAD1Mb
zRnqdpdfiaru7tXz7Z3Qhuc/SMI41MRpN4d2GiAqUao8O4u31O+4pAr8yJ7UDVFhxhqtAu9EZxDK
xOH+R09pjSuwvjLl1uEm9J5hORhp9T57qGh0DHsgai81egEnZaKwdJNuscxo80AsDlKjIw7kZ+Jf
lBRXRvPI+CSbd1dObYrd0sckRlUMF4vkpGnznc9aJ6cxO7MYN/yFniPvq0V0bKYOPvqElbcdqK8p
SVV62OQ8hrYeJjIWUnvCsjbQhSZo+tErm7dON7895uYO/fyib8cAlZ9DdSMxOnIcBWWsXs+rVkMU
IwCYDPR36eUMq5F0dtQSlqYfR/DFBkgEdX2qhciNpcYZahDbBbsUUBgItkazSwUOEqoUdY0K4Shc
oMifB/wKX1GsFRfRAffGl/7cmchuedpdq14+tSHqOhPBdfFzz4FGhuQwgOb2n6hv7V/tq8P+YGp+
nVV9AC0zWD0CPFSI753CBVDxgcIWfVQRXnVduDr0G1fEEmUxfFqyZjnWRxBXTyZXYnRQi5ZLWFaf
wv6ajKASjBhHjqfoFI12Ma3T3fMOAHk3S7WB5gGVY07x7wFu0l+3XmzPBUEzwuoF/3glIqP8AqPj
WGXbCUtn41jmeKqcFwuLiU5ClkHInnKR5mo19kGuA/cRk5byKb6Db/HkyoFWEpNckypCiU+Fxu61
yzPF+ceJvbHNeMQ09MICqocj5M/AgQKyZkmXBjtW/Bg9clbnYi4a87bJy/jM5I9punnquqbnjE/m
LLIaARYtr0scNxIwggyHb+9VUoD9MOs31a0lMAqoE1OLrg5eKe9wh0Eov25QlnzbK6a+kzjL2jEH
zfQkAkFeHMRk0f2FCImqUeffeinV9dk7ykGTBjAslz8a0EcGxzkBFdIvjSf7Ztp0jO57ClEw8Jcf
DqrTvV+cJ1w5GdkfnSk2GUmcUAjfXOiCepdd0hOHVt15GTdkpn0StHQ57eSPOi+VmFvd9kiYXJqk
g1qyH6ofr6S9/eKPQ5Lxo9JB9O9u4FWjWnMMqTwKVBy7nsVHKlbmfVCwRJH9eN1KFxLWPONtL3GI
ugh7CwcEeX5lgjlQdvIh+AHRQzZWsAh8QKq56Jvzfs24U/ZS6MFIieVfsm5h17HdZEqXDct5gD0A
8qPqeP9xPkGjzgFy3/X4F9jr64IwULyIRgmQOccq4IUDF+jw6z4+kXAMfYlkJ11vSJFEKNSuu9+E
irk/9r03aAs/03X11sjcDqJDJzDeLZXDiq5jy4YIhXmplrnigTtllQWqnFY1IgdnoYMYFcjBna24
hiT70yAMQf5V5JAf7798UZJk0x74YmEy2ftYOXGRMI/2ncYme0JQ3vl/TKdV52KXmcngnF2Lv3Hz
KP09IwWQhzWbv2WetBILkMFHDnrJvghDTjoRsm/Kpl4gwr/gnvfE/KiCL/l/4T+lBRKuMY3aaLaY
E9fVJn2d5jj/O2wNeT5KQSznIJApYtQhrBxFsw5/EtdgWsb3PSftlNm3GS9g1TKuNm2ysBUqExJL
9Ad7zaa5aFRK8yaz9PCZA5qwuVFycOiYis25isnhXNDR91Mitj+HRG/MWVqkT9c8tjNr9sL9TOSy
cZswbfWOjK2AX2Ksy204NySDMK5Ec76QzewAq2hs8GflH0F8kptLix/O3+4kDF+MhBFBn0DUCAa6
R8jSWPk07K7rjq5leAA+esBAwn0hMulpRtQ5ErC7xWcVbhu0H6affO4InZjfWQpUlws3Fvl6FblG
waACAib0zjecfiyr9rFxFYd2JX6kCqM5dqnmtEz3135wpoNFdYJz1nLgNs2BtwQs8lcQ1L9spHrt
89XKr4JfuHTJ+84swVxkJfPUWM7ABRp0SFowYAuYAGLmxTeV57k1dG+Io8lQJg+IAuF/7g3ZbRQR
aB0QwIzqizhAJBoNSzxc9W+/+yghvUdF4B27d4LYPZJL3rza1dK1LO5z9xksStt9byTa0mwwa0LS
AgjefjUfn/fo0+UHmasp1N6Umhqv09rFLU52rlc8bUXz+9uXtFu8JSbdoINKuyafyxHqg70frMj9
ahrZslw4IN/3tnUPL57YT+512PLtTq2oLU/7/bKkTC7ZsW0mjXYIHBeoRWkUGhsc0KeyHn2x7dJ2
IowN+bhSPXesQZQQbS0Q+J9uRroiOw7UQXYmNewRkP1erEs+K2K+x4mpt+wJ70Cl5LwYV+qeS1LF
iyAZnvp4dB0MGrlqyEFWqJS+sVD+Fe53zEoBpQ8hzCjdPZ2SaQZqPH8yJa921/6fqx37pXfx10fE
s7RIKzdjXmPI0juK3w0KGM2nkuDQGWo3Oq2tIKmO3SVvBBus0giBQiykBJb0bwZBobJm/7y8SnDu
69yy4oGEEzNS0Vb9vN5z+JbLQypOzeEjkwmfVOp3cy2gBrLHnaLI4fFZPxF5nwp/hAd1k2G+oPGf
vhhr0xnJm9O18ryP0VURMJXkN0YEsfZizjEbQGmIDrMmcT3abbJPcmmgeIwMafSzy27DcmBvAPly
ZhFLSMRl5fUEeuEp5S4Bzom+wThaEWuhksK7+rQTV11Xca8UA8KBJqYrGWciLdEMsHr2jx7/X2vC
GHy6h2lwglzE3QqKD8uDXe1UMwLIHgEIm+Uc+R+xmf9cb4hii9gJzI6f7o5gfvjr3v5827b5juMG
35QWyKifXzFx/c8ihzQ6CNIndfJthJr5Q/793K/Q055EsG8+FmJ5aPmTI22esqU0xUS8E97OIHQq
RHQEGGYNJYcQKP12cpntO//sdS6rjKQiWsNLx7jFt9pp4w3uEKC3SqflHZAiWUI8ZSERx97CpH0I
d/idisXdgbkGPQ1eJAazAzFgEzN7w6Im/+WGmTk+EL4jHDrtUk37GbagzQJSd5Gwqm4Od7qDlTdZ
X91nUz+Lm6lGjXtX6L6KuJ8UUhvHdL6csuJDseKUnXUJoMAuAT9jKD3Le6KthheqrRhB+PdIGDng
H+CxB/SglstGnojDzzSA07BsyoMlaUx0uAer6m/FcZNTQD36+Xvz1Z3lqCelOZtRRthhtq2QH+TU
LH5LdMzWEx2cVWM60Y/kyJD0zrcqinlMzo719uv/Z8N92Ca4HCEX59Fct98qQ+ddgg10v+Gb1f+P
/nmFMRPhwAPmZVslfowW8jA7d8ZQ1zcgF8FHTiILiTXfwcwGWAJAKjlpkzknkFigA9UBh4bEAizf
AX+fQxr4L4goQt9eBD9KWR1+R6844YGi9Mmus1VF4kAhEJS0/3MUczA5Z73c+cQeuzGwI0vyLFcC
9XzUdCUu2sbZfa4oxv21+O61PQo2GaeKwd6Hk7lpIxuilIXJX92cpaZhugGxgZXE0B6WALKWAWVr
A5YD3NHkuM1HC8a9i6vJPP9d0MsEDv8HA03V9Bt4780kg12MHeA27rsNvbquhPdhLQgiSiX/eLMi
vOO5ac8FO6oL3q5Ke7nOzvw3g4MD/sr1jIzUvTYP+DJjCjrOUjBbvhk/yMj3iWpq+IJ9KEpewVrm
AcxxJfs8m3mLWqWOd400zBvOqlJW+MzePh+En5rA0+93RZrbPww+8Ls3eS/g3AHtDxc/FEdt/49y
tf5ZKFGdAgtIBz09w70XJ8GDThFPJMdFy5Ccc4T6aXfRTsimI6ZqNz4Na5efEQ7RNb8sZEfeRB8R
Ad0HcyBvuNCI2HehIf+7WFiftoM1TfPxsReZQ4Wd+UmVwWDv0Onew0ClOebkqSdpgT8NrMWs3rvK
GQOxFJxxubivACRPeXTRG0dYUVoI5ZrsPUDDgGmP5hVMk1bXDleB5FbeO3EkFXk6PRwZPBL8+rgr
oKko4JhxNa1y9uJVfI+ouUMj6eHWg90Ytb+1ts8RZC97E1zAbzcbU//X+7OPjdNS9Vt5WGvO3a/b
DzgD42jKIqGXzU2IYZZoAHqSamsHW2ng4rq6xGrgGGcYTjA6u3KLN5doyZiz+BeyVdIEqzGdInMH
HiS+3KfFQwpAqR9Shc17nuB9lz2giqMnZGevwTbKz4+vIeA2KC5Kjhx0iy05q+B7vVKq2zzi631G
65+aJvFfx8LnF/Bhu9vh1dNpwzkhWlBf0vPx8AzJNEC25/WpcIQdAtFA5gd0r6HWfkTNpGlZuEYG
DmUmh2724V44+DDeYL3uzHgs9TgTeMNBmqY61VA/rX3+snQLOenio4u0Ku/8QtPRormMeGVhMPk0
acBT0BnKWZfhWM0mAExSPIdRaeGaaVGWbP6NdXY5ZvH5parFT4GM8jWjF26Ux2PxX96nflt9x+cH
umRXzu8J4w7j2FAe74trr33//qjsx2CmQ+TzU9mXoWid4odjs1JGFeV2VhVMzOsYLUAgFSQ8O872
GHrAUN/Xymgo/nw192k0Cl9vIwLDaZCD5ceXAS7vFHAEKJ65IxLUHPlxobc47ByW5v4y2V/eXFzL
rNzWhWDa5qzbFy/WuRqt2eET8bEMZZX2bqIc1R1luhavu8Wn1SNEdeikj92pwz51sVghLTXZIpWz
u9HYyVPnDNDlqrU/NIxIytPVgDjExTTO/QJ/CTYjHgMC1fjdiqp+r8EtZNZVDpER98khWjaa9r93
abBmTchdL6ehYFT6uxKAJxAodG7SqePAH2IQgrnzcpP4TGE69zLOIxk3gArz+ARwGtiD2/SIJopG
bvlnWCyoxTC5w2PeKd3JflBmWV1QYC42kyEy1fnWZFpS8+vyyeZAxZCB3RnFfxOwUBtsaEQz6Jok
T0ueN5GSCz58gXhBRI/jf3B3HxiyPmfukqZQ2X2ZVNfAxca3By9rqUBKnXV4e97XC/+YebieQ5t+
uvfwoBgtaoCvcbuMXoDC1xgKM6cVgHVwa0VyTLrlBb2EIQHaOXW/eRdyh6zWAqyizZuCT1Uc5Mho
9RocXi5vw9/f4L7hWfrhWGCWqWYa3TKHkVExSFjx4gL7xVIHz6dq7pDAaYWK22Qh7BIubJGm9wxZ
HFLKZdU4McWGdyT2vMjIiJ3HA4LP+apdztUTr0cwNLb76DM3FJSxAVpKHAETDHBaL2xbjVv06LuQ
0qUPZOqHmedViURqKsg2Abc1AizpzSW8hNWTpB/MzfnJ74vml9ZRDqUIXiW43u6ofKo7g8pQ5dEt
Ua4yj3Blx0nWgXz7dyvZtfKgMe5eVzkkmZqlnVHX+Ppckmm1n1Sqi0/T7wtg34ONF74HRLul7112
QGeac3IoahvTHg4RWIcVVPz7DpHftmmJi7rCgYn+Vk8Dxmw4fWkWYVk+6KZYu7Jk80giJpbE7uiG
Xm/Wpi790kpk50roMxRdsqp39akrBWb80l5wUqRck0rebQuXsSrG8QRgKGh12++2nYiAIS9jJRuc
rUyuTEA7mum/hKDVHPulM4wml+zeetW5cvKffBxx7QOWk4mlXq7yW1jW7y1Wjlmvdrz4PuOz63nN
IgNoYoIybYXEA+any9BQNw9U5/GBZHLBxlTjH0gt08lQG7CgZaZU1iOWjGwMGDUu35MdPEQPdHkF
3G4Id4f704Rf8oEHpb1afxSYnrNBne6WedzoWnb42DxrwTSB3XwIg44Hh+66K0Er2yeXd0lqWGSO
+nTdY8JyxHwTqC2tOOjP5iRVIgto10DiXnkDhuqs2fIPJSrlZ+jZxFHhd0m9foR9Ul5KJ0ww+liU
fgK7GLZ95OhzBo17EQUEs6ZN0BCVAAJE+3QR0Nrdgwm5yRPHwWo3/RfvhotHkaPBOtpZdA6GefSv
MhydTxftkq92L+0eEkLe5xkToe+rlYIVwm0+HjUs2uhXgfux7WLQT3+/Oi41tFp1EsvXftl0oOhS
DHd25tNkxnJObcuwOTaA/A7IcKvSjhJTCGfiveFavzVYfoumI8pusCFWOz0XrmtR+fU/9oEo0Gt9
WCPxKFffS9gmDLu996ELMiIsDZFtIZOGZTZx1veRF1N8/Zd9QQMOXMIIIsX/VOFM1Z3KGkhxMPsf
MdUN1kZMDhANvSV1z28s7sRnc1UabM9ec3QV8uUXgyCP8YTI9NmwY3W9DbIN3sgie+srhv7c/w0K
GFZQPFmsvirst7S+uDcImLQuYHQTRp2JrmD0VbwBgkeMc1UVHmcMq06JTy5nmQFWgjSaNc04lV2M
axkq9WS3dmzMjmCNJspDyrLBC8IyCwu5Bqb2bMNrAqqcubRIHwoJixu1CflejtgS8L0lGFTlLtXv
GRREF2Vi9lYcLLH+uyFaCdnJaNi3XJgN1lH0cqrSUURqQaHDAKmrTvVXhb08H3JJIz/R5fPFpX9B
gY9lWw3BzYXfrAmobkPPdxNwuE14wJaCiRHrYMZ+IYmYE853Si1bQJjj2B03Z23I8+Dgf2SrbVXh
Y498YCQP8mqobrS8EWg3cZ5Bc7Hws1BKcHpx+QDmTcQjPdWvWsHXPI47BrBm+Q+il4H1sKTQILnC
x09QRytdXpUbjr8SuYT9Z9upT6/whpJcjsKaoAHlvla9oDqw8Qgq07pGdsmrBMBjadR5p90CLl+O
STx3PkW5qeHms2dBW5iHFtN4c+K7SQbTAoakMHMzctEEQocGXoNcvGNUg+0UfDVRl2H9YRfHI/4D
UTC/zqgh4V1nXOstGzKcirQvuIiMIpRiX6lZTwlVek0gkTrgfww4A/QD72pRId5z4d1jLtKgA5AL
nR2hksLbcnq/O/znnfAxWGDJmO0ASJkY0aHdHjbJLVnuvcsrs2Bs18Eglj5H7DShL5/cohb6RSDV
vDlyU3UmkW9cG31UGsb2NJEJjlAmR9TK5lXoN4DayZZLnexbPS2vwjmXLzhYtGbhv8EW1kTY/4O/
UknhYpLqEOE3B7wO/pQDPm//72TQ6AS5gLbPzP3eUzK+WoGUgDbYbM/1bKx/BwnSGyAwiIqY5DcJ
VBKp8NCXvKeH44bkJG4Ys1UOTesm7USBvPwhzfLgrENLYWhNNM9ZubbDylK0ikN0WekhwuDZGF8q
zD989To1nclnh3I3ENO7uexVw+LzqE57ah5Fbuc2ZjvYeVwVXRUyoF28YoPXdOGUb6Jce+Arw56j
7TDjihz8YyNrqoGNWmQ+is7tZWg6ATfRAOj8w7RDmj7wJMQ2vq40UVw+szc1FBVYBLNfiH/zkVKb
mkoF4SmAK3T1kWZapT0Alty+2qXQzn0Sh8fxgYpmeUa54y8HnvtITgMcn4VrdiVZfKFTv4c3Z44u
eimxPvmM5opN/2WyZFvI+etbDCYrZMrHxCPAH5Ygv6+zXvMJrxdRli6GcFDPmDBrUHV1EM2ainXc
/SD8dfCVSnpKCU+9gcxBPavL/htN0fM+qAzqKnOzGcm7fxSNGppGxlad6xLf/9FVsVnJe1kfB4MN
FlRtyB5p+pBi+LPl+NN1kIXrm2DA58JAyIZTznmR6jW0zRwAZvNbGlA83CYI9DJJPES0XaLj5+Xh
UPw6IJChSLnhW8UJLakbmR4WeeVrTX1UNv26IBotUeqiS4X6uZ8eekz7TRrYa7gsGcet99bxvuBh
MzCFTNgZAm6YYl/7WpJl0CrJiAXng5AjG8Pxpf/WVFOaxkfvWIndII+QRJ1H2T7qVKD9EIGam+lg
f9HenH9641kJgn1y9xHE+jR0GQ1tUSeI9pjA/T5z+BK4grgLjJkoREc25hBx+M9dVaqQtUaDrtrI
0uqeZ2OrDhfEzK1Ww02jpIo4UzrSgMBK6ERsAHicvksg+DovzGC/htBKY6fYbimPXVycX7oqgP2K
Dk9h/+fDkf2WXrONkyyQD9ws7iFA8dS5aZJyyKPGPlf2sFE+aD1e+Mf6D0mNdQH+ziGGs1wLg1+5
CorfpiGbuQHtS2oIaK72J23uTgebajWGtMTrh/KzaTENbtPDqiM01L0u2iUAN6m3TrnYHNU0TbmE
XaXRM06FrZe9PrS/59HCwKVk5PDmOSgjrTU3Krd5JyEaoc+qnI3wG/N/3d2On3khYYc1gfcLWWjD
5ngn2eEVp5pWtFQDrvGmtVEec7c7Kr9Tbrwye3gwkgHcCtPIXNiQnVpQHZj0A7mwYK1CfbCrAc8O
oACfN+ckJ8Qo5WsKI8vgY67r7UzhNlfADvHRcmm7dJEvuwJOzycJYbjN09ASa/kd76Ss9ouohRss
rl+Pcv8zQsfqzvhVE8tfSC1ZpnMS2M/N2aTsmpPFguqT94bbkR9NWJmI3eJXhtBlcSe/Dn2P5gzb
J0ubuwOatHHJxmw73IKOHl7LUVg2uIcnbKj9h0GFml+6WKyYtIcL4CeGdby7TF6Be6R4KT/uXWrY
R+75Ou4dOhIl6s5UNzdBc6wyI78AoQAXwkGA9BvI+xZljtFhu6c5zieY5qZS7bOJuykmNBh2ghcr
Zmdg9+ng7MFVQDU5HhXZE2ca+2WSSz7dJqmBrMDSbZoqSQx1pXEnKWE1OC/e61qhGcYrxGTh3Xbj
+mY7TxMFop1oXA8xY64mrpnBrLEw9OKslK1lGdKTgiFDf6Lb4G1V30xlV5lNpuIoPrCklFRK6giS
d9GCQNsX6NVdpnzLLV/EG6m9o+iHqKoi1OTsIj0INDzj8B86+CbKJoDNTfo5AA3j06bCx5nu9ev2
+oRTn1NrMcysDi5c60K6BE7CvumkuklqRDZpGxO9gXurhEq/VAuMiITU8+sU2jHSV6uuplpNuqbP
NcHHW4wtciA8MHc/+L38iLmSE12/OlrtDtddPxV+I4eL9k3f3HoB9rMU70GaBV8d3F3OMY0hrTAn
vFl2CYEwwEKNRdvlxVbzRnMB1/yYfaAqEa49//LnEbwi72v/xOVTQhqPsxui1gWtGH2FHnzj5uR5
pzTsm7b1VKW4cd/4OHzcgxwWOEhY8c9nvhc5Cxgnhgv/1el5Ocb3U5rwLe12p4FSW58XsialKqRO
te/33Xt/brAU6nXhMMn5/oi49AGiMr2L3Le9MNO3Dp714hxN7Uqo83vuCAr62u5x0z2/i8Y36tFG
0gHs0FWk+PYsXpLGlFTvL4bddrRAZkjwVJAM4tGfPXA+K07fIkj02xD4vCPi1Ghn8efNSrhAB0xY
eZnG7tW+unLdewxzBLBaTLCaaeoycxem+7d33mPWytVroZHFvTeusX36pbthQECH9aRq8dsGTf6f
LAfV8CPaPusmr+hoB2L5j3uPiCAvUT6XpZT2QLKf1fw2JAYLtMtCUNF29aud0QiiHhdPi050Xakb
GkUXFODKzq7iUSvXrHdZ6OnGditP0JIsjO5ZvMa2Kc4t2hlT8CyUwstvwji+V/4vauPM0JWHumV6
WMXRtPbwk5TnwiezzgTihvNOvElDQ1UtXxoCz8mqP3HAegBaHXe0X8QPJNk5mUWQ2Q7+pXc+Fmss
SZh+igXnrGt5dbElk6E4pqJfkXm5kbeQNxJPlQZxa19SlxscMXZYG8acxXjoUtN5xPEfJZ8cSYNa
At5+c4cv6yxrbv1z9YppCiJXcLTW7KjLsXjU+dkIgt21h5ReWQtWLiA+YRsj+R72HIcBiehPv2X6
zMiEY2d1XWy3V4OKDAmSfLuY4kS0zgxMECjEQ3AtiJ85s3J6H2uGreAKAHdSNpTTpor+lM15VBew
9l9ryPQylkvbLzEnOobMTHavyI09LcfHPgMsnuG+J02ZRK7uu8KLSDdYnrZZY0CVHVJaIIN6lgdG
qt6dXDc/ZO5BWghKDyMfnHI39uMKOnQD9ev+9IKRKmea/cr93YvtJdWR6XUyMflAfMn6znMLVuF0
WpT9u3Rq5WDwbMjzEJyI/X1kqc/0+GGt4dmxAyagv3C2o3juSFDL8NXNzEbM77dbQL40jY+G1C5Q
Er5toSzzr1P4DeL1QbvNLC5aQpFqHztlEeSKCibt86R4zhO9pRgFyRzlktfZOkzFKckeNWaLGJsF
mSOoyXnUCEEMvXCPhRwEXmi/bkUC3fvmThzzL8xOddR0FMAwcTO4Gnl1VZzKTCsptA01FwjJ/2Da
h6CHEiMvZkfFh5F6eHNJeZA3kf2qRioTbIbyOhp1zpG1oS9gt2YDga8atSpFR9xuQWp7zZlmmwHJ
YCWw7owvlm7JOYVjpy5xZerhI3WMaQDTv9jWQwMrDHTH8Lxin/Ll1D90iQk0oElIL0TZL9bKhH3m
WbzBlDUhoNVdB3g47nj/aFONCysvHBJ38xCyVDaHRd6BAh74SQ3YiXdxiPcM1ZPdJx+INP/69FJm
Ehn9zKWQlb7fPEMWQvqsm/QYR12AheZWXZRzCz/KAHSiQ25BPfeUJe5UlV3Ly7qZxhgPQ+GeTKqA
7VyNIKNkbi3Iiv+s+75A1IgRfIWaYOOE584j76iDR3H/Gvakdn4A/K7skHQL9m2agKLHtJ2ixifq
/fqJ+KC3HbV/5hfh3ZkAzaYb90p0gLVkP4ExO5RC8czfNyQK1dyEvJG4TrPGi+c8rXchki+3s2NR
EC39vYJaMt2JWdk3JOm0wOMbY6+s3ju9RHJlaRohUQUrAdOW3AFJCctlKJGtbkp+kl2M5KlVStvQ
4+q+APbXiEDqE5mlY3nE5vgaBGIQ41v7DBxI7FyCRCWTwmGBI1SDWULw6Mm3xhBmg7jniIy1MlOC
tTnwAiAFvIADwI+iOm9fqqhmwr0tMaJ0lbNx0Fh4/lLCJXkJ4tS7Kq2TEGNTu7loihnb+As7gFzs
RoOPV906pkinHayR68CUFpHOYA+GjFrbo5ORuMmpaCx2eeR+ITGvKg1tosSWtyg28Ct6SNS0HBO3
NgwXhxBtLmLgrIPFuIhdjpYro1KUgf3lNZAm4lsuyfTG/XCwPfegSdM/X0r97X99ykmRMOVebgle
+oAmC6wXsSqXqfKXDK4/aHanJiPqDNroLc6T2Sgo+2VPjM2m8JgKJ5QWGo72hAg5P8RLTT0PWo32
guLtPr21SVA1YP3g9kfsStCcZCVMPC3F++LUmgoDc5sWzkuNaCuCVMxtETAncqj8s/XKxOSFgym7
4QJGjG2pzVAIYPk51szKULuK3mCCwSFJRTBlQluWJoPTVzOHiAyNCIvCIeahlm3dy1I2q+sz5MQ0
TPcCMVHDb4P02DJA4fGCLQvCODZ38/sB7F+ZXtWSvJk+X7HBJ/MhwPflbATswWSme01Xj31ePBA6
aLTKtw83CzmyBX2RglEBlgpOVYnH5pOPEY11FZuEldcxOpziR9m/dkZHlLpCBX5BgrIsnHrQaVqc
qeR3B+Bq4J1a3UZ2AmKAhIJuYD4JprbgFnIOVqBzeFVNQCHdyXlzFYagSxg8W6FvgHaB2cc63/YC
i++Z09bEuF95TSbHOXxj/oJEgFq1rboNMzq799qNYYrmRi2emtykWgEDqPmWqMXP3193dpK/lVPe
IfPZhDddqI50kincaUIoDV7F4LsJdZsFUAhtqxzmKKRpDnSDoNTpQAK6PjlSvOWxWDt5Ebh798cY
z9GlLxEiWfuNWCwbQLpAVTaW1bx32tSg3ovOsTI1vRn8/joSjWFKMU7kG4wlSF3+SjLsG07uZz52
EIiOfdXnasI/OIOFlo/xmgJqmoUU83CZSoew5jPVXJTdz7cSqgDhkyOzt7gTI4Pu21kwsX6X2e/q
Sg77/l3hima8sX8zo/SNl75TZIe4OY663yaLaKXiWzQnNC6LyhNT5NWntehWFA/huPuT4ODyMPWk
1BdPYwJm6qf19z6kRRulFGcWLSnC4wTSIuNtJ9SUxWArh3iPbVJqHjMy+l8az1qtoOnQikxFk2J9
dPqu2AJdM7RQ8luJuJCmWDefAe80cL+9OGmOFNevD3vjbrPQ8UrRfPgiOfGh6budV5GiFVwSZLR/
bhR0umcYwBBQ3s5cSUwGbJoX4e+urgP4X6uHPLcyDjAVI7Eo3PM29PyKx1sb+P80Hv3AErqARatJ
ivJaSc8EIw508IzTNgJD4IuOyDbf1U+ZHG/PE5LJskW/BeUSLhoDsXpd/rHD2wI86jeyDpXdIUT7
v+NosrhdYYJ95OaGWX6FxBW5i6efE3ayJlcK+tTicgVAUbLPXcMm23sC1bxRQfcn/Lvvl3cBfzET
m0cuMso8+LXlAhJoES1Gy1juPBX+b5gPzImNaV68cBs5JsATYoqmtiWv1CAlYWmQ+O7J1OcDLexB
nx23Bj8OZbGfuTZd2Fpr1Jt5LkmD+0cb7sJrgvP8C9BcS3a8Md246aW2gm5BBV4tYuGfPZmerPoy
+aXlhbH0TeKi9zOYT19EeYW1jd+DSfRE1ohRnk67ZpgVAu2Xh7weyGJso3EigUIA7CKfgv63nBAS
vYbykTEUlPcYCI2BVtSzVKTRe3eR8/owNaM/kh4u14aUF+SU6yB270I04bym53z1xbWR8XEzDoIm
83CqS/RZ9CViTsHdEvzYkHBh6vdJfNFqliyRJif27b3ngit8157ZNV9VYJ4opnbNjc6ETwCxksGq
L1a/aEBrX5aqapWPv6Ll7Ek3BDpcW58dLIX5W7bd0+9gM5WBWvDqLUoxRui9aznY+S3d87DrOtCY
yEq1NV7N2ltPgbSYOI5kbhmx97RCMsWsZRhPnwwSmqi9MLNB0zbm4QBavkV/BWaozyPiA/g7HCfR
zctO5+L/hYa85thQnPZCT/MbiztwjT3REg/7A6eu4Rn4gHWTJpNNcg4pCpNAaOu3VxjpeEs3tU16
qv7lY3069OKOMrgfzo0gs5dB9ChJjJ5MEs1mq/S5pjYo7m3eBfHO2Sio1rEFe9qX6kojqK61S5mR
dUEa9oPwGvgOlJgMc3hcmsTG2mQFHPL3DWPo58QY8dJXNDz7wboJhlLS0eeTPp7ldkrMDsFza5Kr
lSrRjE3hdioFT6rlyJMRgspQwGYcfHRYxBCT8AtX6a+z+c6sgAGXIw9isSZS3iclrqlZi8eenFZ+
mW5J3iQz22zKTdYghfQN1T152caUHkVSoqqS/DST/Zpa/4BS/B6nkJX4H280l/UgCA6DY8lVL3/X
EcKBdrDOnuXFGL8GlyoYN961eodn3PwQJXRw3aygimypDgfl7X4dfHGLEayZYFaYEpgdXG6eKeGA
3Y20tE4n1BibBtFBNcGCKTz1/Ia+WF4wB1kGXHCkux3vpTIPVK41Tn5MkdDOuK70I2CG7l49Hsxz
zoIGHCYWERzRGY5snDq63kHY8WEt2NvzrLCfzS9mAxdLsfkMKEHS0KSG1LgVXBvZXX9FIncW4RBf
+giycakNrLGasdsH5NOQFdjwsiB2lBHbZ5iMs0APYCZdJnLETkA/lXuNQuORjf2HTyYKerlaQiKP
u96mJ2/S1vStKxHARRHDgYtFZYNO9Fw+/usJ2Xfc7L05qdABssXzQZm4Cp0U10sRGmUvLCdYEXsC
k7pUKL/D6f0y+zWlQiAfVMKP2+YPqrx1v8vWeSY608G/CjqcUtAC0+kx482wa1QLLaRRxaEcaGJl
nU6ArM3lIBcQUuVuIJp3hvRfhJQpmAaW7z5R3uqkQWjjSgdtpp4mixB9u8CG2vaAcUD7lRfi1c3N
VBzYXiH8tLO9YZbzAvVKK2ooHPxYZNooMEBFBzdoCjZLdOYrB89TkaSeau0EJfa4SO0EwDYK7/Va
CvMKlwJ9901RPOxh4GZ0o/tcF8Rn4vMIjjrHrlCrR15XzIKiSOycIx8Bvls1t6ouursZk8EMsUjS
WNUA2VR/YEp9Lx2VKRYJfo1C91Ntc/sNjZmZilZRLUPBLJJnKOzL1PcAHhxSf6tw6Utmf8YfCDmK
0ZDiGWAHFxMGwcO8Xk1L6Rk2AwPSD0Issos5+rFF143pwQ1Vo6rxN4KqOhdJT7Aj5UkWm4tGKN5o
5fcSjDEzqBRd1e72M6xg3WmAi5iJByMq+d/gnwzpZyOb+y1A64AJZKS05sRYief5dfo2+UF94QJw
M0EUO2HLh0g4JhhnsNg4BxprtYcBbxnH2pd8zTDexiT/fCD3U4A33joIYriiM+PFZrsfYzDokjMg
HTyDdaPgFlhUvIBTbkdZuo4+uRy/mOja8TirGszn/nKMoVLlMMCjAb1nneykePwXMr/31q4rGIzg
4MAUVLPFJyR1ok4v4q6SWa4k6SngI84CMdr6iafigPEt9F7MFuitC6G8rh/Lki1YHfRoJPEhjGYm
5ys2xwXdz7p/G2+M8g+/NB5DHdwgEgSnOjzF0HyrHSs3FanmpmyM6f5lsN6CanOJWCvAStQ95ipe
RL9kqKBjz3JjDJsquiCnruSctp8YRVsiyBksk0dOglwqWIHn+sfTSj0MxjS+cybb/4N5NRJKC6GI
iBx8oBAkBW/RRC1o0rZzqejnn99SifSeRmV06yFxGuipUDrfj801KW1h/NcrnTNVzcpiNIiN4CH6
0qNY2lCcw/Wd5nqw+344DrneW0HqrkkJCyBVkP26AoBw5Jr+CkGGzXqyiHDlw16Y5towfAii9qyD
gmZ5m/BrkhXevBkVFs2pMSu4+hdKcXfXYMpLPHD7rx72UxYYZAnqObLXGmZ3PzHdu8f7XPcf4NZM
cP3GPArMnF8b4Gehui6uaDiwn86fdLElp1/c1xjUfZGhvAotSUbRbS1e1q2TKHh9FiV4DaIsEPDH
R0plH0S2Tl9hTlODReybvoiM/WFFe8GH7EsMulu3GS8jkhaVJcUOowtfI7StHAKq+SoIHb1doB+k
dqJLo193weRewWpOvSvHDT8hLagP35wI3+KOahBUNQkwYQ78jbRurCe2vR3tHBbKBxi4OX1vZI0I
0rfmpLZVsMWBynfWYJZc9wntd6EJfK84605RZs6EI91BHfj+0pd0hldF7bSCrhsOyQmBA2DDTz5E
zcFCHGUHYMhibxMuCygUwV/5ctl+QgaT2k7T8cTzxWBTQi7WsIhUXJwHcDNN5igMheSsjnySmifp
DdXJGJz3iq/B9UP6LL7M8+MusTydnZglTqkRkzyzfK2n7evgNrNT74lYqxLxGqz1NSz24B4My0L5
g3e2/dhpcRMae1eRuiSY93k/5Jl7asK/37yozRTLug4n8vLbHW8bC41UJTVzkH3YlRX9C4cjQqqe
q3BGlWzVfbOExLFjmCx0kScA+rStwuvuGZsS29v1YJcrMNuVrW418LIhes3h4DYacCTHPYxpol2c
3fvpxmV/KACrV86cEySuZR/mDRDQ881PMTnwgFmd9485NHuLi5jzoemBJN+jvWUsl8FaNeZubTik
HJzAP6b5HdXnfWpdfcOarYj258YqUQhqJfqUGXlVIHiaACSPc2206WUs5PC1E2xGWk1Npy3CTGUP
Il4OMzAh7KkJU23vzTPnzbjjshm8BOFR8IsmgPxTb6d0WcCM7xWfVCr5JnLGgFWBRW7t9WwYBOAl
BIHB1lwjSV3ikKhjU3AO9gQT+tps1MriEb43lFzwKc3HF60K8uA3jJ0+ZbsZ0dB5tHdLiFmq8oTI
GLBK84pSU7GeEEK7Dn4gOq/PtCYjI1Kp6jPsSGKbpQgrjxWRkv7OBS/lyPGZn5EbZpYcBbxVHhdy
Zgw3czNFfWQ+w1zwZAaJ8IeyfYERF3x4S3vFIEIA3rQtowXCwByuq8sJZ6OitvLEflTdrDdZoowN
PNBg8ixtBBs8mrsKjrj0GgMNuors4apUcmP+A7fMuNVXE42CX+0s/dwuZnHIEFzMz8sLFJWYV3cv
KgFNYGlO1fs4dO+e/w4/1OHwT3ldw8eF1iEXnIL15DnX4y+sWkbNbUZ/J+7ILaHGgS0eDFS6+mwK
NEMNm5/4coDV47S2GN7UUvmU/pX458SBCIA3Q87V3ZWC3yTlPZH73au1D0DCBL1nxk2KxgQcQ07B
8XXVo+5TqxwxKz52rOw/o8qOOuGXcKFWBO73iZBFOX1TkrM3WPJhKH+kguJzt2rj9SDKtaQ0F/HE
jhopFMTFy3eFYMMnPcgB/K830o8lhm1Q9QIgHIPI+aLeIcYgE2wo4kQyQIS2DxlMm/k8wq19iK7p
rUSMeOg4sLCVH3CcPno8KJptyjhtTW95LJuGQo5hgwEv7MPMJw7KkTECSzoHeIJstzm+ZUuzddMJ
v4SK6mkrPfqEQpdd1Cl7dg7kX9SVSUqEsXPlaHNchSCmIUs3bD9uDJyNA0JEwjqyOZK0tcVWhiDH
4suSIsPSeIojXsJSe6D12uFQc0p/wB7kpEZFJAf7uWBAoOim0OL9iDLm/+IA2ry686YT9e6PCZQy
q0LEt2FI6BvZXS7DR9EGTdDJLYSi0JrbHUlWzZ+sbIZ1DiK5xl9BqX6FRVW+UJ/iFJvr1yaxNXpt
NAudUOBu0b7gLUqmF1HWT9uKIDsjmcbe3ECNuVaHuv4bE6kWtjNvRcwUQgUOb6HFn2n6fZWIChSN
cepePRGjizizjSdz4uGs1uPl5WszznnVMK4/1VaFJyD+OC9LVSD+8c8aBOe3PmLEZD2XCqYiFTEZ
REli76AgWLh6B/SyBkjaHnzJdmkIi6QGJTPzJFoKN5monVC+tKejgnOi7eHyw8r4muvW9fl+U79D
Voh3BUXo99I4o02ZGpYIb9WUu53qMOwIZGE5x160JjLAJ6Ciu3hBZgOuOnQi3T98SVz7bm31ubDt
WDAnuAbKwZGhLzBG1KO/nQl7WQGuJKJ2sWalLufp/0AAyMOPoHDEiBR7c63aDM+9zc1umLmk2dGi
a1XH3VpUG6R5FWDB3jDJCKA9+Qt7VxLb9j07pizGAGAlaCcJOGRdQRAFMgSP88bxkDaK/7R8lh0b
Kikz4nmWa4pBWG8XcGgyIga6F3+fTyqC5yY87c1p+dKC8jH2qyKU5L35RbfmXMC9kJsCiVofa97R
YFquyj0iyW1V/vzgGQq3n3cHBtxvj1KOLlNcdO8B5twZdNSnHd3062/N7mKK2uuWvuAIkVY8ynqw
G/NftrF96N0sZMnYv36JkuMep68zijAqhQhIihr7H1h7wwqHadbsglSzAa5sx16USu7uDAIED0C1
mkLR5KLkdOn1brLibLOV6D4uo+9cq/8UEhS9k0HYJdNl3zopMzVtiQFuBYkgYsZuh6/RoOANRkil
h7eZKg4EWcIltfAPuPHMW1oslAGRvX3SmvOlO/hy0tVPzEKNDSrlDUdDIdcCVmp8eDW5lP+FblHi
UQ9kGoAZxmVm29sM06gCpnsvfXPn/i6GnvJSE7IlR04cW5/oh+ejEz455fNSJftCwtFvNKbNeD0/
F0LVhr1CTHNvgxVEpBbttnoD5HVqZqutzAxFQGdzjiP4lDq4Xf67vW6ynIrlDxUHxTK7+S5Jxqn3
viV4taImBAx11+tquUi+rbBuQ5HKtClK2E0nnLLbP9csypGp6X0AocN7tgNF8OXIoTmjo8M5o+tX
58Yz1Q2UoBUJlcB14TGfPVinj6jlzvH5XoM4Hn+sub1JLr3UmvfdQjycJ48suCW0wMAdhcLOP0jc
n0rrZxnhnW1XA9vzWnkBNrNltgYnghzXjLAxtOvPQK4njjkn8vnkYg6VhypdssMSthu9N770OhEA
2/g+BRjmDQG3Mrxm/fJ5kySmhPBjF7o3i+05gGT0BKhXtImzvl0g+iq2mIDM7Ta/0Ck7G51ugSLg
Pxx+euRO6DT4PjUXhLQ4VGmMbIDup1xHTgMXOrekUCk3ZF+I4Vjgq4JCEDAaWvoUCB6pSeyyM+3b
1d6pBOPXXSS8CFHvJ7ILiPmE5mWYFXld0G1AECUpIQFEhOufgbikIZeiLJF6S7QSfE1Op3B1cwDZ
P/jkbwFSwQEfXeAEcneWNkmRtQyUaVRwkT1O0XYTb/V8Z+FDJ3glgGA0OV1j71oKGqMXN2XbTwPK
TMBnwJdcS6yVQN+tRTP9vyLMbg46ZctDSHIGrJGUdinZSt6xmMB/Hi2qrjEb/hm3XKDSyPPNs7eL
fkLdeEaASPa4lOPU8YZDaZbbRRRrSXlVNf7WaHYgbGpngBxlt+KKI5KBCme/EO4OGxNaGVSKD+Dm
gIVbsxIpiiAYVSToBeZNVJV02MEah/a+QzSXyhFt7MyYafWYkfsuYJO3f9srz7HtoYIXSHNM8MAX
iVlUdaUJ8O/Exp4WovckrnesQZgLx+EMe5gNyYk/JKnhqdgsVK8RLeHXNheliKgszOU/fQo1mHUn
mgLI2PcJZ9ul94GswLwF8X5qNaIwA1cAhTInim6JqOdq9fNrN8metFKJpBeWxnFE2lD2wdbpjXxR
ARKHwAMyPBv5cAbvK7ruIbgzQbXUD9NsG4OgTynMaFExoArXhN2oJFrbSM6j1MMi9AUyvPGgkfRT
qSk1mNXH4TQEZT87ETzjPTvCb9D/JPbTdEEdZgD7hXfGaDKx/vYsu237xbfzUe8HDYLA4OeF1oSC
DYAYfFhHWO8uvUdnVZZbPOjx2swi2FiFB7Gh2EM7wMrM4GQA//QjwNU1Ff4FjKdEvJA2NEhdNtwZ
x/RObpeOztVQMJ0cedfuGxLgEmPU8WzI62iOJkEEy+/UcOQANOJYssJ/wmyCam0Zi2uE73kB4Fsl
YUafnvcfJVYO7iY3QN4xta5GFBxtvXv3fwCbenzZe+QM+4skopEg6G1rp+1HxLAmUuMXOohl4oud
wLO68yDK1TK8qpHnD23aVPEnpQDWPr3ZCt7bFk1a8uxh1ZcwoR4bnvy/SiCxSewjED2IkVpFvXJd
C2jtb+4KvJrhJ67Zs3y2xXXbhIQKSbtVgwUr6yLN9Q2zK5rvRwZaFC8yeGKExhqI6XpP1/BXAJGf
F3n33kBvjEX+ukYWkLdrF0s0T31CJsPFnRs3NV2R1d/vVh5Gngmz8hid3zGrU4j2HhAOblFTXng/
b27N1hRkOOpaR7VjrWJY38Jy4bgu1rGgAtLKqazI0DjTu8HS4tIdCYQgBFi9E8x3813qoYPViTDg
WilNvOHj7a3V+wivg8/mdCUj3KdUrKf4oyubAJHecw7YsM6t+zbnCZ/RvRmGuqmhqdCUD3a00D6P
J5DD+3KaO+dc8iqIUGQnGgxFBxBZIEV8OqgKLO5KAN38Sf1adjxyv1J0tH3d75+DR5SCCbunVisy
F1qGTTdnVjXUJeVq+9PqVaVbmRc1m0IrVkgGTa6qobcA44yArdd062IhwXgq9Ym9ghdY6cYgUm5Q
Cl9sveO4ShTfBwbWcyMSedmlYKsy89NS2Z1WrehFvkD0M+uVK0WILtqueTS92OX7eTFJ1nFLe9fa
NYQpGmKEcBxiG0/v5u2aDU+z56N4/eXXj8ut/3gIx6QkbY/zuaOr7gKQV87/D/DLM/6G/LBAkpVl
eSHSK/KxTT0AUHNKsl1wr8yyFEBB/7cDetnbmT+6bIegOx2wB5bWA2AfVSLBx7n6HAZD/QOLfnxQ
gN6dUjaG390b1K58YpQHcB4z+Un3h/pWafI2dlKyWa+IiXMnXLOZOMR7/vW8CPQwsKEzcntk2jRQ
YcrBP1u9YtoM1e6mth9MfrsoypKY8zL9kp/sCxlx6g85zGrof/ED9hEZ9CPtNTgvaXqt3FbNGVCj
BTNWjGRL8a1iRJVMRyfT5xCXbDDukVv/rkYvRj73O2NBVyjzK1P/BloyMx+AaNEtLNCCejtdACUW
5yjY3YkOtTlCarhFylprHQ1ef6dRg+dmhOkIf5U0gsfbqWiygS0Mwa5o/0DFcnO+Ie5txNHo7uBz
rfcttHru0rtZt6eoBQOjODJPYLrAFuVpq5GIZ2noehJ5ppufdI7qR6Qo8bXVbSHIvE8VfZlGhHvW
p7p4tDJHpYxQ3zIvfDW2iguxFBm3NbZRDykQ5BTG5zXQmWNtrVXalMIKa9qDF+ioL/lcMtWToQud
FKoDmMd33kgxRnDNgWgsBdYtvBgOEh51B3Cxz103PS9cic6PNoJLKLWG7RT8v04KXDMHGxEuzmYB
1xDxSFEtmjDjUKi/1jGxR06zXkRTGMNp01twJaMEu+uvTIZQLxjkBt7uos4sMqty/JK1FxgAVrQj
Syz8CUXP4qQbca5QTY4z3lYgKhkcQoTNNxYpn60VCv66z7BwaJ85aw+LF9uOg/QsdxwvXPR8LaOI
pXJfsjWbXIrl/03TLM/hHHEyLoZwn7BGjfiLBC6CalfK2Q/osVbbHM2ERHeju4GZI1xb+7mNGe2+
55DicQQVCO5HtzN8c20wNYaFDawqbmo8vDy5AVB+0INRM6BuzrERUg2fK60PIPi6QQonRZRa+ikW
7rdHT6g0TyinT6bLYboBDIkPF6ghDSV6Nb1MiwYIlgArXlILB2f1BAXUWInTSOw+1f+jOELs+cpb
FtM2OtvZdmsYNU7DcI0CE7spaCQbJecO73wnbR2oYlOTOW5zy5ZC4jQPdSQSuTUXib28MwTvHo1z
q0WOsdZXt4iKV8HJk+ulE6uKx++N1Bf8thi/j7IsVz6O7Y1WSh0kuNk5J1kccpcZX6BLp6I89mYM
VMIlB2HCfp7NnP4qkO3el9KLj5yocxhG6PJw8WGR/HmT4gsJ06OrXLehZSX9i+DEt3Tp+3hwXhnh
VlvDdfMGqWVk8O4t39aqu37E4owF0RN6Q1XU6BA1zu+36OgPDEBvbLEgzwVL6dymCJZZE3ATRBTm
5QapqlNkS0kcV/6l6Qu651IVAEgXbe+82g2ZqtpohlaRnuUf+wpfJlUA5bTdiHZFUMT+vc+JyEGy
QzaVsDa47tVSfl1QgeIM9PpXkiDAz78DodCyAx0dMlFqW9VQModZozgjyJLpc3nGjct4ruqmMX6m
hkRs1nNkqAzK61DxKcWE+E/yEKn2hsuhCYrxLxnjaYuHmaBr6qJIL7ZY0/0vqtopp4PqoA740QOV
8LhXcg6zGrWt/8mSpaatQqxE1c+wMuWu3RlzEtYvoBx2wjeeIq/p4PO42O19idFuH8OyQndTkqT2
sJDYv/k6NKC553sOWz87gWhnLX8d5Bs84vYd6wCUGqvEFUuP98WZlQ/6Sic84rUcbzv1ip22Vue8
LEL+gaJu3DbUFwUs8udQGLskZrykwgRyzlZBGFqiO7rvY/yE2V660y7KXd/kiuBAWN//UEt8rApr
0QcVOG8kTXWSONy08m6LWEYgUkaY9qLOCEi+56rt7/HS0U5FCiDDiEmaxhvsXh7VFAPVCIBbbcq9
gCnEdu1+7xNgPhnCJewCQ8CeFlDZD6HPMVCJ53nEI1w2xhNDUPCm5GzK1BKtQEFfO8/a0I4mXWJj
TODX0ZU02PGUarS7ANpuv1hix66qXj3aQhLGgoDu4pBurijISngotP5XIONd/3hBo6b4gLdYOWQ0
IdSU1d+86URhGwwzfWStepdp92BN1Xxu2q58aAvyk9Vn/0bkwnnXfqlblxCnQiE9ColMlAo2bnbh
5ZICcq7z95nNOArbizhzRFzAw0JlCgMtRxyKLiPnCRr0HoW5vKXxLCQoCcmeXgyNK7uZRbrSDHIL
i9GN5lMxDVaSMtugQd6WcWm1OQ/MwmAaTCHKJteojuHoUlDsmSZV8KV92catdfL2vL+8UVF5W3My
OAsNkpgV+/ayCYhT4eAAQDOSbusb1AhdMfftTV7hX3Zoqd+ofUnmTmwah1Z/lEjMULwg5gom2Bl0
olqmbf6D6eCtQ2NwB9Tip0He61zG3wi/CvXs84E2uOvET5AHCEFjjVDwGD1SUQUlV1MHkNkO7Dpe
8Fdamqu480m0hl+ivpB7Xn9eXdk8ODE+wSUuxJaMZXd1znimNQ3a/nfW8bGf08zJzXcznsOJR8nM
IT33xuMCalodh2KVR47UxjVya0gVPZ2DNLokEX8B55aOsUhTMGprlNyf5vc1KBykk+Mgjhu239eG
U8sntcMYR8fP+tb9JjA/6ls9/346u2NdFO4S7Nt7Ij2gV0cFBLE+/xycMqICiOoa4I+X24ZLNSbn
9mMM72K0yllAuBvYJhA2vKgj80xC8QMm7C9IeYmPoIs7DkTkP+pF+1w2v376VU7VOgnQEMEbanJC
thqFKxdZvDkCvDKWNKT7UR6S8jVbNDf+qwEumxDWlctC5OphhUJgYyDe52X3qVMu829y1fjUmidm
hYKI9gmngke8I2hjUnAPClxCG+/cC9KGY0Rxo9qCcV2ZwV4cLVAUQ3PzGq0221Kt6vn6cSTqT1HZ
CSSghve4LRjlLiLSL343uYmGxsFrZ3yOoaKyCFiN1HYCYf9KXxsf9PyDXe88x+1MrlEadRyXLaaF
dwZS7XZ3lD1mDRehH3KqQ3xtyibju3u/vfz8tHtibkjaAx2SK6t/Z5mtx8xX9tyPXi+gbILJRmFi
A9odbuT3cp6zUp6JnWcQAmFuGtycaJ8L2UDMiSBe+LDz3smFevb9ifKBmzwvQSHG5Kco+JxJmBbc
/uWCH0roU8S/e31FaoURVrpw2jjDgLzCKBI87cTf7PJ+Sk7+EtjQUJsjU4ErAWLxP2LvJ+z/FEY3
Tf69nKx/EAyzULm5G0TQlg3lVHDIwnXtF6aIGzg3eKBqaWDYl9/VzaQMlLNAf5R+VjObrZvlTmlc
1FlVMx2UY8xUm9ML4NcsKDnAOTrE2DFSR/FWjX/r3bfmY+oNsMDN78psarollvdK4ekg2wIRDeal
C/m2VbRXZUmzuM0OMODF88X3NP/QbrZTQV7KOj5rtMLjxe03sAta48Sp+3wVKte3iS3e2w+1R1Ka
jKYFgIXNNs186H9fV9YU/89ut5W/HA/I4b63yZ8DLSmcyOJI7symgYUqFa8Gvk5ENFIG6P9HnCro
1tL9PLOGpHr7Oaw6++miAKJ8Rvv5tQtIvlLhV/9NoDOHtSgWbQWEoBvthXjszIFBS3RLfUlf1WN6
/FgtkgqLxYJFXtZhoxBCUPVA7mULqtTIp6lu8P+MKzcgguMH7ULgSFVQja6+K3Qr8sBSzOQfSar3
QFu0xLrSsxWgkWYEo6dHN8J3PbLF/9x9PAgsP/BRhJxTbh6PZZrD5qW0oLozPS4m6/+O1NgHr58P
IhueM2ohsS2wxdNG9qX5OOqsqAMWlDEx6E5UNEFVeiNFCieBUla2Nzyt507cLbup/qRVSoQlGbdP
kqy1N1m25BDuhl+YmpMHka10Ll49GhY55Qd7lq/fT6RNwszxUIMFctJPMiUqOQhEn2EfsrF6EWwS
UZwXWB1zllxygMBu1CqmgAq8+N70zJiBBh6BqjMlXxa83XJTRE0rwqRlUsd0dy7WqGs/YArzNRjM
q8EejUVE7GUGHgaY3rYIL76wb6ebX+JM5VipKTIwXK9NDfch3SfCexwbuNhDuckCBlirCIA8m7kC
QRO7arW6aAf5/8+50BYgS5+SQfRa8ayHBOXMCpTV6+9o9cGWLIYf+vjhzYGdUCF4vP7ZS2PTvVSH
C8xD21aVabY2utcxN+cQWFqqGlJFHCC04bUAntfv0IDSPRvkvYJGdnsS9RCTfcPUot43JN+7v2Sf
hdRh6I+5Lnkj7OvG4/bPqDz8JWY0Z1Z8JBaPWOLMNWwlu5F+nxyvnvhiA56uQ4t9NK4pKOy5g98O
RBwReEZ7hMFKdzXs+mv+nTrgTFgcQuZgZYPGdacE+A0A0CZbt7ZngSF9Ve7Ydw7Kg+E5U6c38E2Y
oVnHuq9ktixDl8lpj+1X86cY03mzVKlvfuPPQdo0bm9AMpuvGiNOJUmzif28SyLj3jEdZWUHP9+8
9zcWqGIwi1ZP4Ja5IdeWajCCxsulo3/yloXKNPaKhu8CS/zqk+n+Y/J41ycqyvlUCuepqwXsLcVV
25wRL9SUQUIeZMa+ah+0hXX4vRPR7IptP6u+r01NTO+ZE5B0Tu4PLQLU6GZi+JxEUqylZV5EZlpX
0yTU9UnbXL/CSncbneKq3R508PtQ7N5k+JvYZbaeCeOZMu+3D9XGaTnBkzWuoDkHS4My4TYoMbG2
3Gpt5yxEzJZDIuLi0drznTibzpM3D9oy77P3QostMKvuRJUQSmgIfFhfPGSHYIN96BJdMO/cazDL
ZYtAvpC+IWQokS0kWrqYZgy51nelE1bPpdJKVBaU7DpVBZakb1FnhYR0ji8wZTdoiwHAn+pJF9JA
Rq8i30MVaGdfNtjzrSl5fcAjOAhDsUZvReiMKGTNgcp4Mxaxh/UUEpbR6ByOM8X2Vyh7XDyqdobd
kG3xGFG1jt3otT44rrW++COtXVxeJQDg67NOnS18EfqM7RryQs8gtOu3aDvn/f+ZFwASq6huMO6G
YBHBCQoUci/6UVVNX9VxMh0DYrogZJFNDma3Zeu653J0Zv1POozDlwQ4V+eZ5WXRAuK8+3/BFmlT
tVxqMIz3tLiAfUQNTJLNLu7Hhziw7w1fePJjcI7aPcK4798Vk6QudKVdnGZJqtQpnw2NykC8h0pw
h/nDCD4x5BH+fBIIRPi8JdT7+SpCfPRIqIjuI0bGA+bbibF4OrcWIG0R8BVGkomU0A8uq3WeDf1S
mpibulMW5tpcp7HrS4FSEPVEwLLJBCRTeDnHzyzzCoJnf4rNAIvtLIQCoauEVp5GEa567Z6+p6Qf
Rux9Vi2Kmvz0O5JKK6kAf72sbI47YvXDh/cHtDTqGzeTPeDgXSsg8XnH/ePEDQVSh/XvOCAf1fQ1
+TjAuCKObpNSW8YLg85pBOS3JZ2PbwuvIBRIGJoAmZk8WuhTSQr1WRFioVEU53U/Gx/EPKMthFsH
RrNLAZPYVmWumcR2nhM2pDAInOaUl5BChUcbzlE3FncK9h94Aj1LTX2mfi5hyWmxaoxvFs03jnkg
GCj337LVzUn9bwG3T5cINgF8Cbec6N+rhBimxKWZuAt22+CzZjaq47bxoP1Uf54xFU/hVbT5RtIq
nc1PwtQEiNi2DTJuH0OgOi8Mh3YMPCsO+FZslMxGwbv08A/4ZQ3IhmM5GP3JSw0zoxjTw2j4KpEj
o9i52oO3s/VLDGuliuaBO/AgeFoO1EXfL+wc5kd7sEw1uLLhL6oN9mlM70tMHIs+bPht0e8X3PLd
MYIk6vo2nXNAaZ4rxr3mIIWIwQEPgbImzKQvW1N/iuNSKWyNK2BmUpZJhw2lLUl9HAFvLeTWeqX2
c6TL3ZmAgGL3bL4r2NVp+MaYvEfHXyxPCEWU357fWjQrIqKnQa4sV3Hsm3gV2zaIeUgVUqqVQZ66
R89Q08puhL8rAzVmzOmdQreVE0hTftZVHadgn66Ye/ea05/tSXBGcNG4cDZrQYHF9AXX6GHls9hK
e1ZeMkrlEQwdiYIecRK2AkGFGDIx7Xe42/kIly6iA1gvaI32RFLih4qijLxzPwdZG6uF3rYeAk+t
8WKR1bpv1CxI4u9YcOY4290qQvL6XnYC+6flIr7CSeyVLP5jVaW10xHnm/A5M9t2/xpIWrT2fZ20
Q9CW/sfixyLCG62Yyh1EPrx9CHkXECUrDgYHw0YNgWdpmMUWTdaO2F36SaA26Nxs78sgWlumqd6L
QMu6dGqUnTe0xRSRIlWXGeR69t8QlJu8eHJG3gtnbN60or0Lbnq5/ZLrI6svkGEQ40xfnuYGiEjl
ewhybKkpF167BtzLkG4/M9lnLk7d7Xt85h+GRC3aLGXffQoJ5E5yAeVjZYYryXLCvfTPY22ni+8s
wBMUXueMGUvgeM0kNgVd8hlNCCWeQ2v9VaXAbpf3yDdV2LfyHCqjPNfkuWtEnmT34LQqKannPynC
TbNC1TeUhjA0EcJbmObqACI1C9A6iag4XymO8G3QM766ooiRz+bAgnv3RwvGEEr0tq/QXGrPmlu3
EyNlim5AOLd691E6hMchWWKaUT6GabKGOmxAH8C6LHJHIm2JatIi5LggKya64ASKz0Zf8oGXG1Z/
ixgyx1JODv0yZVDd38j2gpm497hJG2dLMSavAbGdDWTxErRSm1cOh4370AXswYfgoFVyw2mw4Db7
9Vr4Boj/SrkXBvvkJPJarjca55RgDq7YeDeaMJ42qp8zs/zIA3extJPq1Im1jKuvROb2ndqmzHe7
uUXJkokoEE/y7El77nNmKeiLB4HAnG2rfRuxfbB6ob60R4uTS5qvQp31VmCzM4ka3/8WNSHDqa2w
ws2INNHdtVr0n8cbFKwxjTnkkL6LgLhSagDnUBh0jlcc9J87NtfQh5Svh0QvcUsXS7CGDYj1L1Jt
QJhNRs2Zm01yg2Sd5ZHrln9369QgvDgGS+zP4m1aH6ddSM4SEqVsIozMm0USm4zj/xJNt2sjuvKV
4Mow8lGawsF2Orkmj8hhgUV2wG/cHcvZ89FV7aPVeFEPIQwa/vd2LY9UWXzuSjFDpMord38HSWFa
+xqwREKFRcIUGDm209FcWRAtU8jJM4LB3Ty4pEI++nHej9SloACyyhDUc3+ULDnqURru67qjvEBX
R2UaWOqZWkGtNPnNk2bhwt5TD51HDFeMgQofU0/WDN94iJz/DQJci5AQrkIEkpCjPAb4/WlDR00V
ZRdRbY9J114YEbklYr9NRi9OWgAj1TO8A/3QASfrbgq1BqCuSWmqIHBK45LyyHSo5jdOJ/Gn0S6O
SDO1/hWdkS7PvnTMeRvlNkAEL7G7HaUEA6Z4Orq0oX13RSDVrpWxj4IhWEECTJfbunnO6QHG2iGp
9RqZGgGRf/3OvN9sPuKUTfRamn+YtN7xPi10+aEHtSIDnc7lhV5h7kPOXvmtdcH2nv2XXTqokcdq
JEgnljuP9bEFuIG5qoEiztUiH4V1a/XoDJB032JX2y8Csr0RhSt293bj1pSOnrvc3RAz1/nugjcE
ntfJoyK68iTuUT3j61c+7Tb3yIGdYQ+PtPGNmOXDFfMPR/XT3uIZA/ByCCxzzW0S9BrLhEiZdfo4
upgZAsTMDxIzscBu0HmFJcu8ZcLHvWRcvFdhh8h4++t0yQpZ7sjR86y+2qhpacScDgEjXqkpUAmp
s+pQUMCXS1nFW4ZQ9mP3ZLShQFxRc2+fQ4OHYVeBpzh+ptSPoLL9bpMTwTepOIaz4yxjTAOCLsfT
pdbDdL7Xv7kmuMA9dZnz7ddBpkzXz0PpwQgxxWEAv7QKLam5S/LYgiQ/irbeuoUXKS7rurhvphYa
u3QzNRhUkddd0TsIlBkXfZJmxBZZVOCKKMz1SEpEt1WNRNNxsAQyN7vVKPVtQ8apGsUnDOkA8v1Y
pis8sIqpcFTZUUYRdLML8CABbLzbcbeICPtU71KViw8XgtrVV5w6a82piytpo3RxJvkMemIMTJwx
tBdJjFaHIzhk+OfdJ0uSLKuBAIBoqjWpplDpnjkrxHCLyuvq8mHlYRmvdup5v7pLHAjeQ9eCNksX
jB09Mr0Mksc1OwfkSEub0BkTUN+cUMLQLQLdL9V4tqKQa6HKn3Q2R+/vc8PWONSx/qMAMzzbnCiF
8MYfYndhqHhHuqulk8xQ1MDl7mMc2Q1X1RBdeMRpssnGVGrREfnDfvsFopZ+XItgg1HuUvE7Z1fu
TmmFvgmzVMLOwYQEXjE5ogGxON98CP3yLbnGV3rSSPfwI7Yb4XNEsPaUEU4lcUUqHw9nkuoKUTvK
YlJVKn1zKTne/sEOLj5cUEiH9gNspi7AGz24+dtEdJqMFxMb/knE7NZb8sI/Et6TjL6IRj0ouNmm
sP2+HU2plrRbkpGKQSSwnksWsyjWDw3eq8smAEIpQIZD/2oV2Sn2jETxT1xaZNoIMfd7F7Fodk3f
mPGxxL7Tu1implaRNFHzM4WhcMikZ4ZVKY13JHYnWQH7C4az9RQvmEFitLW+sAzRTtGKlQhoZlex
KgCMByZItHCbTtwdN8a3L4H65tIhCGNVCoR+Z+KCDeHhwUK6FtsybRYJblPIAAeiKUcRkZzaQQ/X
Cisov4qlS8XjwF77z8dsvOJ98OcpO5KrXLWIePuAFpkhSi7fbs7tjFYf2qBqG8EzFbUMei7zgjIb
2BeAp4+xijHKQA0gqSBwyHPdWWA8asLC7tS39dJoJ0mzirZ8NzTaEKuVcr0dvvf6voTWGKTF64S2
foQ4c9QFRkfJC8WJyjj7ZGF6dhoH8WozDWsGgfPMkP3tMv6gd4XrmJGTFJujVZpLqsWqFrHr/eLi
A8JHo+DnNccJ8h+gCSi3gMp29FV0F8bKjpaCr3Hr1cPuPWLCDHG9T16jGampD0IizbbCG0XQyxaJ
Pu3vUEt89GvdXTWH19rZIHTbQFem34DQQrbO4EmX+x+g+Imxyqp+J0kPQDxc+OFVsh1mpVMoRBr8
+GFi+VIeC3m2GlNaBXBuGhIzjAE/bpOf/psGOqQ+F2vNvNNRip+JW/AlpIotdTX75M37RaR/+gLJ
H27Vpqfe5sgfYhSxrDUPeRvdW5sSHI7KyftTNTyihsANLpgOHuCGT7MBizVkv5/FW6tr4yDtGUuL
TVTrqdIc7AaWR41wYYtoZxLSXzMsLyiQrqERlniWclsiiDKVT6jCJlKnnKM9qj7MIRoxpGHFFUUl
kZVO+Af1iL+e+NApFVnS9UhMqfGkKFXm4/5I766iak/mZPXFw+v84wPD2a2/bGZfwNPpnLzXs/Rd
CSc0ILAKFgkjiiL5CyndIj1LE1fIcBD1+jvwIOHNrg33EhHiOuWoYj3zN9Jyq0/BVU6YTv0pusOE
dgo3hiugu7DWUQDGxoa+cnmSAIPvDiSOKXCKlVVbTc7n1M7rIgapu9kczLfjA4rFHe9N6xQqjIqp
nxM/lg1Jb2BtCVnWJgmu6dSZ0jyyo+Y/bwp8bUNIZy/GQ4gKMJG+L4hHP4heTgJ+rYOdJzsg42sm
yF48yWZUdthJSgNA0dgh/oA7PYiO8w0N6JRBxx3Ys6xb7HxTjXh5zxEAqzMdbj9IBrEr6DtmQeDR
kVdkZtTUn10CtGCEio+TK3eCsTdcOOeDleq46xlHyYB9/i7DPhhUe4KxoSs1gLi+B5oi0cpvQb8c
78f8gtMEJoizccHRPJRiVtU0/E8XI2uZAIpZnbIeryzP/VjnOjSfVPmxfNTxdW/tu3HjZtZGPdzo
N2BubUZReNulOHjjQ2a0ZJOS8E71yXnuo6J637TpY92gaGlg+K645QJk4p7DhcsFOM+2vA8mLxXB
zFggbuaJBykHsUNKBquQxEor509ptYERJC0FSn+l3Ejqfd1DcCEcUKG/yI8l9tygYPB3LDGWGR0E
fmjijW5Pwg2r2TU1qaDtf7lFZuGjyhh/YegCbBQMoHS5aKWJnSRHVvrYZdT9GsRYPyZcmUB4KMQh
tXEXV0jYrxaLEE4b9xHpgdr0AooNIlBGR89n5JdfwsJN8soYEeCDLBbPVPdaTzGlndFOIq3jZVcS
/IFty1zuEhi2yq+eMwIF5HXi8LZHBymiVCLCk+C6SEJp/WizPRoWozH2gkNfF3YEa/bczmDWrqX4
HEiKdGb6JjusefHVpO2AvCAKMFEK3lv81SJ+BFAMr/5tu2ePmoxJjQ1HYwWnpBwCOVo4DHByPoNv
ik2YQaBNAinbUIB74iS4h1YBsjKR9/cBSEKyiLOCa8GWnISB6Cx1A4OFiN3qFUkaYCcQbO2I7oKN
OQ8G8CkdgFJr70eIpizT4Bog3WUS93N1pj6bXuW96YipjLZnrMU8bUtZYR4olOe3O4c3/WibKPRh
CmAULznaNSDE8nyrkZEBDdPW8CSwSZKH4z/v+ubj2U2+PV2nxc+fg3F3d/7lBgHsku8HnqV/CMwD
mLWQYGXyodxO2q5zpaKTy2dxKfRerWt3k4mlqVhi7/+7elXMGZGMK4MoqtH61WElaniKvyyoftlp
R91vjyJBkYu3O5y/XAR4f358QWF1/8Q83sSd1z5T2vpPhQ0r6IopAOUxNidJdLUwuQLsk2/W1VYb
VC7rk4JfNkJTqTAdXDd8CIlW1CJyM6MnFMl/8ZPq1eztaqwqBtsaYT08CZsIxKxBshRlk+F9o2Ql
9gHAp2rmB/mDInyh5/FfJpg/GAg9O1zEJ5OQ2oXmWwSdPyWSg4IgP170eLn9y6QAXst0huUV6axa
XcBsR4pfQnrpC8HLrlTbnx+xxxID6bWaOPl+UGoUWy5+v2iUFArPA8+YN74OIAUFa12BshPQDfAb
RqJhzvbAZ1p6A6/mF78CyUZDxD6YZ5luqAzvE8H5vhWD2JZuhTPCzoE1fBOIiFlySXE8sxG7Akha
DSXymFNJpXdcQBIHt0h/n5bVs1aWQeKSKqqg3d+mJr9wIlXPlzfJvZIOtcS6J3FT6aVO6qQMxfL9
zJs4MjdMpdWfQ7xa8erQoPfVNXK49JdSXF3k6gTCdcA+jNqfO6vcl0XH4jaEVE7zk1NCgKh4sBz3
B1krYSvo50u+1mPT5bN871rv3fEkQb1KvcLUpCu6loi8UF8oPz1Gwk3Mk9RSHlszn1kla2+VR+PD
22sgv+1e9ilrYmyF84CmXVimZmxyUjuIAsuYr34rS8OsEznQaU+QhTu2ahZr1DWdkh18iY4E0j0s
TUkNHAA/fgHrR6iFJHA/lmM5eg7bWfFfYd8s8QsCEugjNWa2MfvBFk1LNK7QR6fOnDDlXUA2i+0J
+6JgARBa+0gTg1kxB3Yl27VHVRXSGQhAfQNDNr1JEBlImidD3nVXm6rs/j/q/Az2OA2EQEUo8Jpn
bwhDCjbQk+cFvKRAGfYNvAKM9J1eR+odq8grQ2XF+JpedVHLx1Cic2fq2EQiC2H6lNpshuYyzaxD
Oo8ARefsm5QOozfiKGHKZkz7pBSCrK1CfMJLNL7VKdPdErtIsIsqGs70ItwEpR8vYTLSI91KtPZa
Hfi3BEP+PVI32zoFYhems2DXSgqJJI/mKbkexsd5hT1w8N+gO5rhLvBVxniHYCnu5xCUvQmJYCC4
3SKCfIhlAInQk8SNIq3Mw58f1ZOLyEBqeHtvRHPNUewKUi4bHOSsyFi1n2gTuJCAL+Yy7vQkgpq1
r8TXHIqFmP0CuuKlQ0EsgGDTykW9sKUDkb/gQKymdY2IcilV2DBaXw+Yi2yAwJSMlRlJKy0ewe55
p6mzwew85ICTIBAfR/PojHqWdo/OYLxrf1/OpXFdzvdejVNFXZLdm8GdVIDMALMjdqgqWzVnSio9
S2lkV2HtSU8BiGtsjv0uubo9LP2FTZMYRLAPGgYYDEYG9uu0QABnoB+mzvDatkLbdy+cLg0DdLoh
zLZqVLywhqln3xgDJ6DwMC1vbccEPpcCenAhdrFNBN71G9p/DultXcvXb2EYcmgRgxsG0xmy1SkO
epguU5pDgdy8SfEOc5QB341wzKyQUc+rFEcSM6T52SbUI5YexyQ2I28895wFskFa3whBgG/lUlwK
1d4dtCArhNpeH8xC4h/y3JE3rLR2ezC+gMLJvGK3HPFALThROK2mGzADmUNsq1RZBi8N9L8QLwGb
Qb9VXfW34s6viH8NBqHW7iLnmkbZCA83ccDRCLsUKjBUMWLSlQWUXDdn0AdEzJz8cQpfGA9TsqBZ
0jo/zZVwz1+hPs3Xi8Y8ydYQqGaEz0xLvGr2KxlMuHhWdrR0Xm9VXor2s8wpWzreyYNeuuHg5nER
7pOCco8W0kBwXToa9O2s/7ODS5J+nl0KR14R90jFvmXAjVYU9QXqr+WzFOwCqX9GZ1yYTnGOPZ1s
m3JL2yKMjsaSuCx5mw3gzyECqifx4+JRn3nCPyXycffoC+XhIo57SH46WjIutpYY5q4W6S84lW0W
Htoip2eeVEhhCZU4apnLPl0Ir12GMJM8uWWl/gmVdYwr1ywKaV9wtseLhaV0S5ryNoKN7DiIl+gp
pyeLgH4J6Bzb7A37pGVylTIt/ZZKklgHeyISkPNvIMd4qTa32R0sXPolkUgMFIkQsXzQsjNYfTW8
08bkPjlIvD6OGCx/Aok+MB/Pc6WLOfqWVttzvA//b7kegifw7MrLEPdb+idFocMlyzHt466f64zl
LhRk4gPxwBqO5Dq64N/mYUOEewfxrVdk6u6vFHFMJUFgfE3s0DXmXaO+XJM4tzj6vonw9kYPDR4J
UIR3yXdn1qAS9cD2UK67zN1rz1wUKCLGR71npSUbzpJTdQpjZjHa0jvlqtmAjEcS2jzLmEwqoRVY
79HBAw6WZf9d9bgDM7hQ07TARtJK9dl5I2GDe2Bi6Z6lzGHIo7Tsxu6oAxFhjRb/qspVczh6LPQy
qChiU6vF9q3jtiAjWeisUs2u2kMjbPTlBjaCiSitYzEehbcpODK88P8LzphOYVdQzNq5+siAhsUh
j0uUxhaRIDsoGJ/O96FFju2pleAEGxPEw3bxciekVS4YCIkpdczaCTl3m0WyDstlMI5x7p/71O4m
e+E0LcZ8kH9iQuhDf4pvlVEBQDtVuFaho5CJqFQjuOaMXVEFikITwTmxArLrM9NM11zO2wiqnCVw
DaI0SctdIS3ImJTkaF9xKlZu7YXKPCo/c9jow/f12f70Imr0rq2WcyfkSpP/slIywqV7YaYcWPdW
rFVDCoKTVts41qNdVqTvIh3Sq7z6YRwGV0MrDhKiK6qEOYKYgYIpgjiHtMGubnVSwQ9jMXhYA6A4
JExfqE7DhemKUCTlO3CbeDa3c+3Ga5lk7lCBWTr+n3ndFOYtp9sEMeEi7LxPy/ZLWnL130n64ejF
97xVKyomWMnc09fkHN0byqrd4asf/kyxzXtWNvQd2htAQi0455gvUNdCBLjQkDWX2Mj5PVH7tz2w
PbopSOcBxvupjJjPQrywr4LIpp1HmNw7D1YI8YAN9TYFFuLPVWH00f94MJKAE70JHmBDuZYt9rw8
eXeEdYjTihT8cb8YIH0+Td8UlA7Aa8fs8yIzzxszOWyhmrDFjyRvQ6qnC3qLY2Sh4iAVZFPNjPPb
6SvfdKF3XyGgGLcZ4areyS7Y2mA+XyoS3FmSdsU3FY7xtpQRUnAJ+l6fVyod3RVeOOpSX/10+GXf
fBwROpD5UEcKGZnGXxXgSpVbmYBTUn+zuyN+o0E+OD0xG3saL4b9BAUESnnPPcvDRwNFsBpncYeY
8vaMIGV8mon/OP/7+NaO9hv7xV0/UtVkmGcvYN8so2/m8EvyW5FXxveCt23lDuRDh5guvMZyjXW+
TW6gpGSvfCuHL1IzQOzLFY+ILG2gkOG50FRmU9gkbfMcianDXnjZTgFQOT+C4liqn2fUWsYNUrQw
OOFI8p0K4kEIKdLC5/HT+GZdxEzA2vhHBsBWoRW+j4dma0Tg0nmhcc3+cDohE6TCtAoUsEgLJmcD
vBBt2pBM3qdjx/S9Ez71sqWmVAGN/vnxCnozQu9Gd8Qj/Zpnlm1rcUI45StntXNbmDRVRHpR0k7W
vZCEN1OVuzDmD3HXGuADnF5/BLZLsrh2BkzJOqF/GxDAdxVj/sqn4atl6TccqPfEiyjjnwIyYo1e
rd1FkWNgEqsAzkuZ5RpyMfoaltF62/q9kVBCrd2Iw0uIiirphTmw13ET4Wte+sc8kcJtH7LkTAmk
tkRjO/PqekDTmUY3sDMykDIKKR2RtKXqTBk2eNUn42D+6zP4qA3O84+ctMflF3e+mbGwGScXBTJE
ecKW5s0zT5VVqrUTAbegDLmWK2Try2CbwNqY9vOSgtiBBqsr7IwBFjhDp0ijDx7lEviCfg9tMr8O
AquDQOmU1zp2gxW03C6cRW8F4IlO7WYqdPTizbzKPKK/9KqbrKFh0oJZH4VzZ20dYUjtlSniczrs
G2PU5QopPmn79z8lSGwV1UuiX1bwfYrde2Y4rkFXRlOerSaQjCLDfkqVaUjLGuLzUJH6NZHPUiLL
dFsHvcqV4XchW4Clnig7cMVBT8molaVRa3+DzIlXlgZvNErBM+19CpoPIARU05wFor00FPWdkcYv
YhvSeTOT2LuV7OgNe+xNqEKshB4oVBtSb6QabQ0ZpbJTt2biZzjgeLgxGKXtAEEKDhNJetEweC6w
FwnsFjRE+V74S6EQjRB2QRyKli6CaVGYgdFczu1wO8ZPwC73S+RK+PPqAh8Nx4Jd9jMQE3NxwADy
cdQ+TWyP8oNyQCsp42shYQRGmstGWfwTV7zSaUbg7ATQNl1OIBB7Y0V3wNf8e9/eZIg3rC0/rUKZ
5M1CVUjhG9yvVN4s8i+yI8lfrK1U5P5j9iT3CfwHS5LDfqTAgl7jv8qTri+zFkAw9aAnBbYmi2ob
TTu6bKpaWdYTkEt51AikJ9anJRNnW8ZVNFlL3m3vUf88eJC9+PktOf5U3frTnw9gl3lDMm3s8ev+
d7X/VPOkpPjGL6J7eIP3FOeJbyXtLO0IvvQiVF8ySVZPwgBYf+uJ3gOnC3wPZkxvwrK9KkG1DgDa
JHA/gYMq3oaZB0Jidu7osg/i03aEZr51rzgSxmSq0TtQAtkxhmon0j+aGbhPqktzfzv3Hv36Glp4
/CkFHoyUf7jJP6vk4HXltCZNEReFpeUzpIwBJkWP8/AyYA2boQD55tmDieS3m+C+u1+pgkJeBUON
ETTsiGod+ZTKmZSpUJiou9+BDKR/4GPliVPAriV9QTRmUJl4HAAxOfllj6B35sDAsbMfRkG2XJ3w
qQDwDwmNv4UIcrGnM1rEvBuateycOzeOM9C+zIPKjJGtN7zklbr9vFmfh5RyoUzA3t8P9kVrJ6I+
KFBLjxOXQCClAVWqaraFwO1HPXNtfg1OtpWTIdjUr65V7afOp7+SEN38+ZHZDi57FvzYP5K+rnKC
f1XeYqdRryeRkQJpkkjM++uRyslS42E9Xa+VMh252gxmh3H1upoM7wi16zQH3M7vlWsbtmVC95+/
0spbv1DGhq/qtcwJEjAdHLZ0SbBS0FKWZ134N6SkxKityNWGWYV7HguhHpuPdUKP9x5K9IpC+Ykj
y1jrz1Z8hY4grGGcOyXxqeAa/RUkWBNEHebnuBFB+7Y2zFJzZHKKCphEzkWqCAjv8qleybxgX0uE
QmZPpvIy5BRpOp0Vs3wUxK4kp3XJNv6gU5+Mjsn065ThVF2B5nisfuXMan4fcpTn0K2oBGWZ+27R
FjbdTH6Sunx1gpzSI1b9AAp/owoLvl7IdZRW5gkrn+LDAFzb+ZVAlffa2aefs0PqeOh1lI54MIh3
KElh/YJTSfaAZ3k40RSsesyzBUrs4VFrY1T+TdOsUlR2LdT/eZey5XeHNPp4Y9jLze0d5bp1u/rN
L4fTLpytDdDQWjY+zjdGglXcVj9+jMGAGV0LrzQlVKVNF/QSazbqeU72zKkJ/TggEFeFua+8OZRJ
CXjcsEQH28+D1A5lifWvQjUaIo1Cn6MQkwpHGwdfGMu/J8S85ObQ3Ggqmr9ygJuzNRzLSxubUDga
zMsGySoRRcvPUO96UgPqkaSo8oEYKka3nvpuwB6SfK/JBtFLwZeRWzHVVDscWf7yQD76a+3Gk+sy
NWy73pcocRNSdUDtPQlGqhuPthGOyvAuVBqzLk9txRZdG9DQNBZIuuebnH7WUe9JBE6mB3RujBsU
WOF2H5PhkCdTejr+YscgBwUY+ZYOcq/nIVuXjqxx2sUzojQesJPJVEUHmIrY6OdNTFZMBAWfeMYF
cT4w9oa6yog3lo+2fZ45qQ6/vK6BJPNxZI75UCbw7hw3XxrFrCqFCHmzeryoyylXYoNsQajHji5I
TtqT6tUIJbv9gq87DfgelUFZQVJcHehvfsAK5f2Dx3p+9AqlZ2MmXregLWAZcdq4mKePeOVRTCjy
ARkXtMi4qxTzE6QSNyul18ZdGYYYYU+26AY1NuLmkds4eIDh0HmYNGk/L4fWuaQlRigZeS8GelVH
L5SAy7951j9s4/Sk3IO6kqv0w64BQ3CHLdgdo/JuAR2DtFjELxew6M0pF9ODlvn9QOsaFKhrimjH
66YU4BKmtqZNDEMf+4LNGGHsBVWBWND2a6z1Heq5fbDfpxTvJg9eMd3+YFKreMUdGKYPpkI+abbF
gqU49KSPIk3KlECYvTqGdUIUqhDM+nHIbmxnXDtd1AdMWa5HwbSjqhoICQ8bGQzIgCysw4mhQLoR
HfEoh4XVwEjutazl5LT6eO0PNrVQlLmVQ7EEL/i3LaZp+KPgTd8RzRnioaUbVL6/N72f4lV3XzOi
rh3ooa/IzhEEmwYAqczda0KRE216vaYZocHkLr2GYuhWlDzgfCqM0ag9kA2FapNmh9vnHuVnQ47e
6pyvXuLs9nJBPUe1uc0zIbX9K6smHv6N/Gbn9rI5qQm9eRjp/4a+zZzHIju4rYFD4u6MYP7zXqh8
nKXgk2hy/P9MHoKD9YPeZPyL9wILfd72VHXrxzcJMnvgW9nPr0ATd0+h0wXUMdW6ibINWFsn+CT1
7EVgPE+NkuPY0VpqIITwytuRbLVulZqV72C3clPnxmys6sbehMcyXQ9QSCp8rQP7FIsrhc74vMAH
BbyY3Nrpq1fNylESWj21YG6wdIkFyHqwEzqAn1Zf3Z4jL0O8tIA9wmad0cFbRRchv3iZl5BGHo0y
8u5AsbrB3r+HZ3tBiZmK6Xz0L7WaFL3jLlLCRv5bQanWctp3D19HJk4LTXQlNQHqFLfZPD3SaE8j
CRTFSaFYZRVVCg2oa2XmHSkiOH/0KfMo//R2tBaC6hx8dCVGF98N3OKvz0378qlV1/PAsQzt4c3m
8tOPlBWgLDCMw/v3allle2a9mByjaWcu4L+Ycvto3RQxIPDGw2mvMlNNKZ9cbWgZSofSt8yaAMxK
ou9VvfgMYGnBkxMrm4zRNTfL2oE9wZMCv39H7MF1KAKjQ3WxSOh6EiSqULHy0S5JFEorDQoT6GcL
cf5M0Gb5mQL7P9/O23KfBW/ufTgYPv6EpCgNBg2LVtGGu2YldoIhrt/J2dArby4M/0cODOpzCBrg
YSy4o6F6VM9+zBmU2b4R5Ybtp6RBEctDEdebBIVvDkEmsgBPSx3kXrWQzqwHo6lttRYZvdLH3Km4
CW5VZs5LVyuxFclGlocHK5xDXdyDJ0UKdVgteJ93JflIJAf2M7uhf7TcShKlfRyZciBD7eyTB3D9
NLtij5QfjLL+yLF8mGYYtYuKVUTGDJaPAV4vm8fDBmz2E8kQpU/fxaYmrHOSawGZProOShiyChFg
5j8lvULFUk48nhFm4I0zMQPWCoy2vCLP9ERXZIhcnwMHCwSQAsMITWxbwFbEjwWG0zISHiAkMNRx
kAPquCmxBwDfN23BleY2L3m2BI8KyD/7Dglho1bsBnEU3c6ufVnl2IyFxHxi4H5yIjszZorMrhUJ
SplFXuEASF9uRjPm9JvCLymf3OngJ1fB56LpnwpIaTdPm1EC8DcJap2RsvdloAd9DZ0RNIG8TSXb
yR6htB8tZSZipa0FUFP81rHZzFSj1Ic5w3QWFvLR7WKS39+vMJLkTwCI0ykx2htT0AacWP7TqPXu
V6dW0lMw8ow80X0HbcXyNXt9iXosISc8EB4GbtX19GQqMnXzuSLjyjRqWZ8/5ZdzrVqntOW2NsW2
1RyHoJPdrlUrNn/UMabpoGnu7FpnxruC0PtB5ZyjbEg40Q6VaBMUlrPj6oB6rKt47fxrzikgj6eN
iuQhYQQJk5UApxF7WVVhoGaB7XQjKpOD/4tiyFIWTutDefbuXblolGVBDffh/BLfUX5lgVNxc0yd
OE8H/uEvyZcLM2R/N/EkZfrwGu5v9Lu7j/fAa29j0fEpzhx9wtWXkXs7lWZBbFeU2LfXP/QKjEGa
ateNWbO2HigQsomBYdLq/UQxmKbRMwYQNWcYGi24loNG3WSU4HsVDMcIjei902wqSeuGS8oYevFU
Lvk079YVq5aM3rG7RvE+ebuVchXlpf2VVQ7tuYyr0AmTL4y2l1ORLGn3Jhd3oeiJyZUr8TyaaGEK
oLSbJRw21TDCzM5FvM+V35mCykitqNRLaF2P+ibh+q1l2MinOFRrM38DA401sp3lKgfLdFuHOiYZ
65oFGbwDwJHJnO+WUSIYSDDnZAPaMVy/wSFgMF1hIad1th1rptAoTyTbNyB7XbTyW5OkwYCzpHck
nif2TUlCGGqGpdimOc+IiY0eC42uf2rk4XRmW6ec9VdGhkvBQyHd4lODg8C4IKTHP4UPZHdo3ZOj
Yk25WIDSt/FqOPelITsN1jV+Et6rLpYQ4i4elA+ZyPaPqcIj1AuYhc+/uqiAl60SzZ7hd2+nu/y4
5tMQkgA5hg6vbx3CdFCHrZeeVO1H1vs2axYlPg5+jokPY1G0YJ+oGcbFpP+1JgbLAOurJMUTgXcy
og2R2kqsXMntFPQdG7pYCVHyqOtdkSYg0NwUHAMhM5/zzKwfgdKoOGmg7b1gXBEjAHg4XHoqf0Od
TjdddZaejKecXYy/6A91oBmAowutejzzptH4Sj3hHDl5A8ULFIs93yE9sOzcowA+2e1pf5+7yd5O
oD1doo+I+P4b6Iu6i36QsLF0rKiEm88B6KPgOnKx10hBgCkKi365+40O2jy+Y484Rk4QzHhtwDcJ
woy9t+bNhgBh6p/TOJIdqe8SQgo3onIBRCQiTxHTWPtX128mvx09vjz//SJrRlYS1AaNa0bs9X6r
P3A4MX1a9rTx2gVnshjia1MPmjDMY+6mchO8HMOXjHNyhqqY/r4j4Yn7lzOz9TNlT3mp1PHDHeWg
mGfA2OlRENJwBMbX91AzalrYm9sbAtFPKFG5WLuqMBXr/NyCVTFkqokkBgWlwf/W0m7awLBqOlGH
DeMDkcaha0ikX4h/gJyL2rNN45KX1rAEXFc9xl5kAq5b7/8pmVpizPAcfC8o6cKbC00SAmnxoSNN
RIfBbc+rOTfo2wVN3K9sc+zi5nhzHwqHLCVQ7mUgnuXZsAhSd4epUHSp4duV7OOZ6kb7DPKCDxmX
fhwZbvULBXBilfr7jbd7Bx4EtxRcrtZy9kTyOVgvNBOLKQVN0sFDPMstWdPq3rQOSpCELjXh8Bbu
+qDXXyWHmB/K6oRP++VeA/3CWRQ/Mw93rq0J+eTTNB2JfVUaDpj8gExKWIzuopDUvYx4YbrBzJwp
1Eo2x9K7b3wycup+a0aIt1Iwa5B8lZPedyNORZxQAA3CuJ8N+ajFMiJvJsyXXOatsa7pnt7HqmJL
b56ygz9jAz31w47+UsusV/sdcZFN2t5gBhuqO8U51d7b3PCuTT48PQIlpfYy34diwvUd2lQ4zPmu
mTBdXlRVHyEsxpe7ItgPZTuCDE93plqVZm1znXMJccDI+PZomyIwrzliK5ShJiJtUvrRNHcxcyAA
6Cml3SyXkeI8BtNH8Ts0wgdyzMEKfyaE3ovTmluGPkbro7jbjeB6nBjnDtuDM8gE6Crj/fMrgTsm
vcwk1fn7IPWi3PqnH31mZaFlBUvlWqycDnbMF1U9eneHnsXQFZRWruIlVKh0GN22EqpkO2V/0NdI
BobzJqlEpPw7kWdEDmpgyC1bFN+AoKvwHZfiNIwVxPhXslxIOp6Kwd8wd4UPo8+SOZWhgcDUj2Q8
UvJBWQus0qzKxYLyQlaXeJ43RKGslw+JvWS8/DVExcgkQ46JXLv0ajd0ynn9iooJCIPyqRjuQerJ
a0VUDjwpi0NW6Q5Fv1k0Y1O1FpYoOQUo8i5uhh6sqB6Q4Rm+yLvczCND1NWrRHs5vRajT0Ta+ASl
QZh2JwxmjnipNVQCXvTcP6ifyl3xyNByfX576Eq8cS1uvMvOzb8UeI1z5Q7zaG3Q/ZTFioikFxiO
ZNSr1Tp21N0/ONM2nJ46LD/UOmE9W+wNH1i1oomv8hvTMoh+nGv/1KubRFCS7AeiahRcd7ykN5T8
By8Jto+V6OkToCx491455sE2Odt/tyIYJDnCO8o554cIoO9c7mDrthO4TBtD0vR20S19V8G08ni9
lusmwRgppsOWjk7fzbcAEaOcye2d2Hu+U82849Xnp5faTGus4jR1Y9vLfBSG91G4jRuc9e7eXvMR
+m/1EY4rJ2ULoSXTk9Fjf8knxP5vPHKK05ut87zOSHira2PAcI+I0J1EKPe+BbRJydYZAq/vZQzV
26t0/WPBfn+9K5u5ii7cL289sYUzHdLlQMxUh3L1ceuPGg8EM2IS02py14v4Ubj9a1vQ4mpY8IdW
7tsghPwNUyrNxBh0rXtalywsij3kK8jy7snIanUPQA7zZIpUHRcafo2w7faEAws4R+QR1/vp3fp2
ZGgUbnoboDdp/kQXz4sHH7VFXZXL4VME4Ororb3Dj/WfMxxgRZq58CyfpXgnSW4p1dmiGV/7aYDO
X3yO3othsgR1VhPcFfHdiWIZlRZMya11MqrDcM79RwFB7IjmHVSWNrAyqAeEmEOo06TiuLtD9njO
8RHA08F88vxs0Jjm5Case2Zqc5XMzqtokUNSfg4Wkjz7It1OLxDJVWnuSC5332E9J+0VpVUq8hMv
etQtIFXFOr4XDm0V/WYBqkN4wgwJ4Um4ZuHq9grrBCha1kZCnxk54Lf0QkwJBorNCkQzChcWa1MS
u9KJseBLNmIYfUkP6dzd/nm5vHPvu+Emw9N3ZVbzwQjBzH8sh0Re8f6S5dzDyKah31RLQmRpCkdR
yYU/9MYZn0zjo3jqQOl8Hc5mZ4TmN/ZUUQCj5x94TgDEwRSnKsOV5XeYH7+D1s2ojIgvI+XlTx/K
rYz5/oRDPEKaloMnw5H0IovPnNeD8BJdvRLeMK6FtABc9ti70HMKdqkQKeiNTOV0P+z2l45hcRVd
vaxSiIRpL8gNNxejc5y/ZTxzcGhUbxVHUCBC30y8rG0lEwhGOymS4uxjrNqAX5yEwafsVowyQV7i
3QJ/hry1yzgHO8Socxj9jqGCA7tZpraJM0z9bRl/6QAX0jCL7pkW2Iwhg2mh10c42yB1aU5DCs6E
O83nsN1VDoASnLrpvDcMnlwuG3btAkdUNRKph7qMCNT+b2um/+90Luxk8HshhF2mn0YBBhZe9cNY
PzfFdB3ajG58ZdVpz47m8e3UFl5duE6HM/zVUR0OMV+vFPg105YClk15BmuGa7MlWYA4RtcoPMR9
eSYt0CE1mB5tNII6wSRkUf49REIag0c+oqsYOsZiwbRioKp+7agXRLtY0+bdJLb8rstw9h95Pb6t
6jQtyJZP2gzunHj642G6XhBY4Z6Z3cqFJaePMtJacEDSZuqTBW1AFgujoBVhYq0aDEHByETUeuU/
ADyA3nP3RD1EsZ5XGfJIpzFFiIO3e3BZ3FJm7ix543FthnypaxJGChE9nxTPxgVwGs9yLlpP+jCM
drTBNz505+e6ijISruQm5rbNT0PNVxi4T5CvLVqnrGtd7ooR2zq3+9fZi/MiGEgJ2PSqesZ94QVf
AOY0y/4bGsagdmj8mwwpBx2RdKU/acx7Bcpt07hEhSFh4B9oEHH3JAu7V8cqY7kytVktWJsaxuuC
/UW2zgVWMepcAjUCAyIdxEM8ehbPnch4tFTumIFZKc1pTXhLmohzpKDYYpinXHpc32YBCk092O6p
ba05lp4QFCS/HmOM3Otnooph2zuNJoeSZ47jMIQ8wdOA3DebZ6J8Ylqz8AX76rxoTs5zCiG0+8df
hjgwvllOnR74U4PBo3ungYFNSVaGry6gltn78ZXTlIBImBcXst6pt3+bfKPJLLULHN+OiB8lutuB
HNGjUGEPl3dCU5wgxrd/tFhOZKobnytGjZTqBvlGFfnyBv5HM79Oa5yoUfdY3Qsw2YqEGH2YWBpi
Zbtej05LkpC6hKbg51zkuA22fVbwnku2SbwgAWz0pQHJvR7b7uCWx1ieqHz2cFxL8Tcn8hctS18M
xm8CpbWUR6boLxx/qdo53jyKsXiPRxeL0CGJ5Fb2Ll8AKhAQ2OpnHjnlXcBWrQN8ruU3wexycpAA
GgpmjR2HbdoK7gJzwZr09TnytfcgZClu9zxGsY36jbOrhzZlOFaj2WrB28xYx7HlQVYFKcOsDOL4
AkbfAHK6idEn2w5mfFbyBr3GIoKR7ErM+uJrKpKRJtbu7H0fB4USV/6hMibsB1rYJ8EGFZBQ5b4n
AjF3GHGO3r4xjOAnUoMsZFIz/vm+0EEKbyzzPXz/9Rtw7J5sJEH5Pd2Ds/WRxfTbAlD5Q+0nKIcN
xAGng8xJWhz8f3Ke+5raxtm3vjycKjcJj/gfpyPszT9/hGPyPsKzEzn6oKpGwCN5E8D4GLjACmed
D5hm1YDZZeNR4uQ1dEOJciwn433XDJIKD2y17KsMS8leD1+O1b28mlbAlySRHJ6bYEeGifkSl7x0
rGNzrjGqjN6R274rZw7jRk4nNWkgUxOXU7jcsrxo0a4gVmmJgCXX4xoont1e2YJyhk4UzDnI9CRs
SQq595F3er9qnt+jewzY1nGBrI/HSCwT36tEG0PghRoGnoXXfx3unPzJcPlbraySvTYReRSmJ78w
Pj65HMfiNx2CFkzNhje3chmP792TFOZwiD4ZZ6x+nWtzkYVjDBJgzJNUqJ8MsMo17NIL7GQ5i+iK
ptnfirTfxNeg+ZGdy3xFxQlF2V/0LQHStmoqpfR6dVRlTXhUjotmBLXr4t6DntWg1GAqr6XE3L56
Z6xxg16PbXpDXvs7uZNRrHNlAESGdJK8+WXNjeLhUQQ5eITXpXWxEWUt4PlzXpoprCzHFw+1H3Le
jl7aB4gblklBUOUUCrBpNTfaN/Sjf0b2DZEEfK9vNR1Pd8RNk3rH9E+9M9u9DlTE+OhdsJTmebkH
wFCAhE69eJUXfibzGp+qmwXfT590/iDLLD25ZNzNyFKu4QV7/VlNEo2DkypdQgqbEfXk/huYqYzu
lquMqWbvPopP55Yas/rvXH9BLlSx3CVRVFAa37OjOxvoOQulHzxaSjMXbzBUxRC9jhBVD1GGSuJQ
QbRPcO21UowLoI3WtKw/etgWyeeK49odwaC3g3+cPA4j3Gi1qZbZrf9S3In9eYxNozKU5+eceZe1
ExhqvwyAFHh7xoYAuOkY2d7JV/BU3KZxosEFSVhtwT2ZCbAm4PuEyIdIqQRD10KzXIPVPedVmHPg
pwwY8rEAm0clFtqlA0QJXMT2a+n5gbHw8VQCqMZ1X08D/nYJCrj7PJjz2Oygd6ZguQpmQ3OWz8ao
jq6SXvoFYccaPq4iLsggAmLo9vvbyTllf3s47xwjX+OXlv9UJ0cruauaO6VLQpgyXAzPOrmgW4wr
kQ82T0z7daXDl+RubG7RXlKXt4foFZIE8tspakzFlGr0D13z4vI8I68qLfV+lJMhoPcD7vBEg8oW
FofGnDNqGALX5q7ukpkljyEu4AKDW1hyVsl/H8s3ViWkNUDp9b40oppWrgYfih3FAyHEXYu0t0hH
E/vyqJvDkfmaolKCXee0zeMv1oUINeAlf22RZBiH0xPt0QaUC2iN1+RK2dMT491nC9Ke4I/aS32v
l/LfxIOZIsmHxdwSoOZAncgYWm3e3zlOS/LVbZ1CIJA5z8QNtsaNBcY4wL1dWjSth+par/ne6WY9
rHceIxA5lMPz1Me0iaPY4HebarLOIQiZ0H0o9+/sqYbK9q6dz2ofA6fU6lQbd2gHsIOxqomNMMC2
gzvWJtj/GSaUBlEvlzmWcErodWRxSQQCe0bu+PjVrHG0uT9BNoQN2lwfVuuuuu6ivJhsEQQgfbsa
4iHt1UzmR9+fw62/34GPndwFmw1lY4ddEEpcACS9cpHtYBNAIoWPUfr25Dx35J0qV/7ZHbBS/LGA
+ozDiiLAZskmxa5ceCW5IDPpVpX/1I5ejWH1BqAqpl3i04m7m9fyH/p7KMZ+5PrDvHNI3YmVipCL
otfU/cMwN54aVarwpjFDSBLmtzhCmFvwTnwK9RDlsLAdc8N4Y/w69O7QDiJunfi7rvykHp7Ofdlr
JNlS6Ou+p6hKJJXnJ3f3fNVG9oPbHEUWtD/pHvhuCju/tAgNo3maIJRoTv83y/qeul5KTGihNZKN
aOvUQzjosFXUUxnfVRtCqCIHjxmxtAb9BY2rzwVuBDi7Z2aJawURVLpxKtK9vfNmWlGhx5egOK5B
IjWHXDsbgTwce0KUJ62ZJIA64PBfkQPwzBWanEvAO65faWD/tEfeuDozgGKm8kVL0ok0j74oigc3
6Iho3GiswSfy0dzM5SaWzd+LK/PM4dvu3HKFopF5Nops2EwVkP5k5XoFNqFiBcjltQ9lnYfhLvtD
DIWFueT+34z1KITkEtY82SZX1XSUdRLnmeVriv0+SW306lNxyJXG4priZgvDMqn214XtVlRjWUbR
HV/RFRIIFPGsy2zZMAYWySm9SRGiCm7qrZCOU2/Id/NZ6CSzzX8KUurg6g3BQW5SZn3yX4Ucj9kk
Qryf6xqO6yMMjueriWRnOt/V9FMLg79Dpi3H+yWsbSCpnVyJz5UasdjEPuLjT5HsmTfmonqWMhIT
sm+cWJY6zrmVL8ycxu+rvjuVGlsyr6fe7BD+k3PtLb6/fxlD5RDKiAba+ZXy9qJQ3ma8BTPndeJU
ASb+uxGSQRcNuREig+QalFziIA5rz5PDu+TWEInk2rpDQ0JS16qapJvwoPDzvXGQoZZWKSO/Vv2k
1qmJ0j8VkU6uq2TNAfqWEU/NEPRDSEg+yQLNkk3oKH7J4o74f4M7KpiVW4EtPQYQiViERXrYzbQv
YEmh9AmVaZn/UTQSXtqNcuYvhNENGC9wqqAUJMfOyO1V4FxcEacbtoG603cdgr00nPJrbHEDy24B
FdAREdQxy1FuLB4Cb2rnCn+ELeeSi8O8QXULUlf0AZIKnIoMF4y/Mg9ZuVVkCSJGpVXrtRwoGPYZ
MikQT2xLJKgq2COhINg11K74XmC1B5fcc/gULO+azcOReE+dX4aqHrm/2ZD+8sYuFzWKxp9V6CFQ
e5POZd6z9GCRBpG0qivCtwWZJoAb4wwD9pGpd8yk7PkMLkABDnTe+T7Kt6s0VN02uO/MkAPg73ul
xYq5Szfq/PGTzWt3u4PVy/9qTX2yEmmgzgdXc6Dm71ouDycjxKHtD1IbWKrud1Z40CSipp+1lvjj
RNXkb7uKp29qIxbZLpG1N/Pm1bNf+SMQTFVccC5c+g796p9DPMxAIVjkWWCou/HMScyjQo8Gyv22
yVoM36NTONxQmuCsl6Q/6orvxgjr3nMXVDmEnYS1dfIZQJdmkqTRZ3hnoFFFYL+esHZ6QSUa1y+6
f4gIBdk7bFQnr2cqfvdXzauPTQBGQVnzcLzYgc7Fkw8t86bUo8a3xaN1DJ35lfzbh/YINyDF6o+1
p3pqZDajVZ3sObKsDuqNWJGXqbxQaQNrnHis5sPsw9Ok4KV9J+CbptzzBPEEHYqi1XPmY0U1/kuH
9rvwjEPn8NxFvFeJNufm1ypmhNEvxh3ejdpstimyxe0qevwOeV3QJfnuFuFMIV5nNH1vbyqeDIUd
cdHrQ77ydZXTmnAKlCJD8ZIpxhC4xiQ9GpxohfpkEGN9LcesohS8gIhriN349sIKxuy2WEm1sSQK
5GeHUKIIkZjEmSovWdegab8MJHWjuyD6y4xEVtlLvfpdJjhnXME+AGexbEes9oYJnU28cR25dK08
YBQyBwLL+qkGTS+cplNuPNiwfpXXgy/hCeYCbtjEoaewC0J88yAO11dzT50LRjn5TQomq4HyHLMK
UlcpmdO8UbxtLAtyCWJXC5ut7O98/DcyBhMblHJmGw1bcqSRogirjYf7TN8tf49NxDzFnPIIJHYr
weDKR1sNCdRc9M+qT/jQ6WcVV72eOjesxlOGQ7UlpdTuA0StNINbvCcvOD/ZSPJg4R6pg4QwqQ4A
1KXj2WMKPKC9XyAUqfrgv+3OVCe7lnh9S4fFEQXd3ZnaB+LQxVGvID69T+2zT5v4aNvtIzgi5OhT
y1aQ+kofMq4sRXFQwR92eli+QrtY4pY1dCADhjQOKenw+78SDnCeZsOij0qsPT7tkF4Z2FdwvTeI
oMkwLlPJuTelmi21W+RgGxcHo60yZaQ7IhgHpLU2Tvs+Ko/JrJTnfx5Z+uTXEVITbsSGsmnUui3G
vh9wNcrayAhMHm50nV4jGhMPMtH945WT/ohKbRRHCpP0TLOzN98k4apLpXlICBP35WzTx65eI5R6
nXvFTRejw9/5lUkcE+xcHWw2Mhp9MgLhaSbaQRAqhqqF3fJ9X2onfWrWdy2KQbFfroUGa5L1YD/l
TBZs87auZD9JIYOqgdcybDvkuFlsBGPbdihEZDij3PVzsz2uO7jQNMT9qK1OIZ3pC0YC672l5vxF
VL23/Mrxg/CLobBnNKDbGnEoiIlS8ByvzM0VawvU4u4IEemLu/R06za484tYLmt9E/wwi4h31kF4
Hkg9MSvGmu5CVRF2p3Ev+pEko9dPCudxjpwxfBNCYoEBonX8Fp3Bun5TRhSo8KwHiRJE7OTa3i8j
sdZjOMBRwSsiWtsfcOtyjj1hNhO++VqQQYXhkj77wRpwaW3SZAIedY0BynxrocBjAi34FIIsHd0N
eIH9VFWdxwM9TtygNso0Y2NNnPJxe+NXvcS+/HYxJn1BADFw6W2cnnNkL9sO8wEULhNPs50Kd7KB
uymK3X7/0zvDoHiaH6rkMB62tkoq2qatI/jvGdJUh6CwUJfr0FSCtAo/nnpIgbMSb2LxW5EVQy1N
hp8PlWcm7PujLXVzwNUU3mHshOjRP9vN90XPyWbaC0I7pawksmYU9FyBJFcTTZ3/L4YyBgGYLfbJ
9VKkd2zfP2rVbqDhyyJ5HGO00kJysnJaOXjownsJlAGsxi+duu8rEyP2KWtbU6NcAjqA5wWuSOpF
SSjl/hdKaj27nGmVVkd0grCmuBZOJDHrlctgogP0FNbOLUjC24vlytO73WYwzuWPQD3tMVHMFeOn
AOf4m8LiyGL9nBVitPV22WySCf8m7RcHOrI+pi41BD+45ntAtgiRdyAPgnyp9ix8V9ty3n6RlAmN
Ff/zyH2UA2ySFttU+S8XGesq1uBY5VxXwNqnfV1oEEFBFR7KyRgkRzjl7IQ6PXh7TMnlFIz/98Pd
zq4SC7BndYh/Sy0NMI56zi5FzDq70c84wu0mvTrpF4RvRiFWKXVygYGcYKirDDZmA1xgHhOiLaAr
kp0bISxs9e2ZiLwQtTVP8X3KVQJ16cDCQnShnNHDmNuhRWUaY0f6DJ+UTyp944qYrgr568YjgQ8L
QQmAgZuf2oRFfamuy3fH4ujGRGQJn8KKki1D92Kilw/dl1Jq6LXVT7lbNqbhjXLja7vrxGtjAaMw
4uMYn0RkHy1XFW9KOfI5AyBzlw1lxiogxuVQyChfvEYygJF67emLD5bYSiVAqrepPSzCn6mkWmMF
tdXaRvs29aid70/oJhQMq8r5yirTMEecNdVfwOpsQ4C63t0QmyBW6nNJRT56N8KWjPsiD/hO0w/s
fXKuwQG5h17KpwzXB+B2x5NYj6p6OW29nFPUwiMjLE/Ynsjee4/qT0neu6TxBXeHoB1o3+dYw4MN
3Vz3lEhfEnM3TBDpVbjDCrD68Wsayzhv0P6yMdHfEJwar8MjEEBe8Q/gYmiuEzUdjaj8intu+ZC3
lSEEkM9Hbpv/zqEtcIpY9JRicGuZ5RXlCyhz90tTkJTTt29TNtQXym/AxSEVVoz7E6H1YjSy7ALq
HrQ4eAlnp/LtNg6Iz8t5bZw3lSLizXR+fJIKmyQ7dltzzd7G1UHmKTDyj/2JCKtItH0XXZHYNasl
X2vqIVgVpPPV+GQ8WbQtDaWjttzFZpZdPtcPocJ+8aZ1clcLrlTqas2CA6X3RR008OfmL3covV1u
XmuiLhzW7cnSjARkBm5yN2L6LafRAU8Lb0xMH2lVnuywvb9X/+fYUBIcNx0YqTOnZucI6yDsBtn1
VEr3wxpD946aLZghlJ0VL3ChhLr+82SFPXpsHlWeyWcBc96i+7lZBNmBYBydvfr1oTbyWZwQ9fXB
0E3OtpPfSzmo5n8CtNPoQY8FIPVnegr1rX5LiqFiHPXwB+YQDSP+TyoK67qDBi6WLof7h9vD8pI3
hbXqm8U9gcL2uooa1+LSnZcBy9ETtTr1Q7ydgmmStxCqtrVVne3x0d6wGIkAnt54JsUUE3RzbHII
ZJIYcZN0suoS9Vhwpcs6MZAqFusOhIwdPaQnIr9g3ABfprYbELGEg4qVYC5bhIl/ismWm0DBVlFQ
LDL9yTT5CKgNjyMHJn29PRspOjSvagmPYxEeevAShaXh9Q5urs4Q3yZlMlOHRLUSTwaO/HAX2adR
9YkVkBUduojbiutAQuksp7QXSVqk1bb2PEUdzA1d8MYWj9rGw/XcTcPqfs/2sWxGJdm9N3yJOPqN
HUpPd1TylQS6GjMU57rLUQtJIoNbGypojqe3kiBJsUB+r2c6XhICIhUD2dqMESqPnZxV0QVKfYn3
7LATnWuKze623h1QabD2V84Q76wCz7BEaDLgbsNFUgFHKhL3OambVLjJvaCctqWG1av+xDV4wlaP
oFA/yinusxKLNYIM/3Nn78XgLnJeGOch5JP0syaSP6J2xg/NcYLAHzl2hrQLhpDteUEHJ5w1uPlU
CDq5+i22w92dTiJae+Y94VlnEN/6T7ACN4JG+VTXWJ1qi9do+3udcDzhzS1ep0HsoikEqb1pqP/A
d3/hXmy/mxf7G4POm574rFP3KEBeckaWCZZscJXwnSWRbIP/uiqCtFIOovpzb/GANBJiGI787ynR
oNuUvVhANUCkwEZis0n71YflxGiDHXvjn/K/eWcGD2C95955Rl/4la5WKVXMDqY1afkma2/W24hB
s54G9wEdX1nbbLLnXQpOQimAowZ3GxLUQEZpO8sRQnPeF8/DE4WgAfB1zgvWmaJjZWxFtn+mvP8h
W55dhqh8/PBZ8qpN4TBdla2hQ4sWgUP/i8a7vCKqxmztEf0c2vD36S8D4s+7CM2uWqZJ+6S8a4nA
0wtmcyYXqNU42OAckkW4AyG5QlULt8wRh4+5cSpZlu3j7jbqKCa+RS+wjCNJckhF3i5nVpprHXnZ
jYB/S2A/eJokmssv7XNCrdqpy9FYroLSID2Sksu+/cHge+IWQjGHTEOA39LORNCPBfjKGh+ZmhX+
9Cfp/kgQK3r9HLtblFJPyJJNtheTK0ANXobdoymcFaKDx8jHRe1AL5TypuCY51+zj04NFvfmX+ql
cVoVQ61nNgVUJjt88KW4Ap90gUwE50flcFoRIAyDLbu6MAsA8XD1cvpW2sVQ9J0QND4dqqsaRfGU
b8iXZ9Cj6v41FCuJtl5T3gf3oZ0J++lVrbOLFbWnytSUxsdm8cTvZJj8DPPcCf1cwHZS7DToicFx
Wj+rrqNYxhZmT0xUlNW9C6EYHEDsi9dt1a7HmgB7UrvJPLzHdi/5JmdyNmyaE22DHG2cNVxl9ZTi
L1NCg/4O5MEKQpMdaIWtcRyI0Ye8gWrr9tq/4l79QawT1SxhyJLwhlVWRzwgOKkAh+h+Bldtv0l2
Ds8uhZUn2stg6S5ZLKdr4fmoRKNLz3HfiELriKEZi/ps6ppnxy5hDGXCCYG4wACtZwb6oHwzpcxm
jncxtpv0SeE/zbRQWufn1bkpWj6BwYXczIWXrSs5GqjxozN1L8e9H463vjzKz/mPuhCoduuXURTm
ykTFCEIhcFaVyNzZczZ+0VGps5NUVDwQa+4k6bDoMa/WQdd7Tv32RKHzcmJTzbOXOV1fXeRdo9rW
8LFmoASg5db0kF9+uzfmX+ukDM+t84cHobw978nmpFAYyMRD12a3oWQdnODg1tU0wI9pIZ8KAIej
MuURDle/xpyZwNVFmUolJMh1uKO2Si9eBiRsABLe0HoWWTS5ZVtho1RKDOQa9uQMc2z3eHco97wO
q4pKmjva08DP3dv5y0GwfdGO2Lb5C4NiW+fxkGEjCPtYiUC3Nz23sPpoxrAu9JIE6+ksI/1JjtVk
UFFEtBj5dkru7DtBKpnYwUavPlbJonh1BbJHQiriIc2PCYniecjKr3ib9XrNnyJ8wf6ypO3Pku9o
FmFSfMNQFM75PDzU6EGcjyy097DT4pK4/whayt14jpZa2V/K72JAusDgwdEdU7/OqFlgkuL1oRxH
U2HwOna0qPE82m3u5UjaLTZrKafnkQ+NVdNURnXtyUtQ3WAX8GM5mNkKPzaSqupfmo+C2QWo6uyG
OKTPy61LjGnomg6eOqDlDuCwWdMiLP9TQ7LUC9VszCCGddfDHOCKujKJKWFoFIL+C15y07Nj2MnB
OdRTQd/hdlqhsqzhBrTdoPB0RtgB1Y6e8bJbjHi5zGPWx3JCo7ZUmjkcDMJRI6xq5lj1oAFi7pIz
63otcnr8g55xBJP+DkAH0mztsUUegKlB2qqu0X+5qNHKEAK6W8VL73+v09TuXMfYl+tAYHRAkjQB
+t+ptlQtTkl8ZMoQb98x+2he1DaUDLkASlD0USDGDdGxDZ/rLQysq6FTEqTDvzSTERO3UmGC3TYd
O7+py/7jOuAMR4BEWIvuZ2retISLuo5aF4xu1NjMKUN0qxfcGBTi9xRlR8dNlC2RpIm8OHLKIE3n
ap+im8UtOiqH6DitSBCXUwm9SeXQvEUbbCXl5qgx7KcTRJWjSKBr6ROSMTBQeVnCymCndf5MHq/R
Suy9oOL4dvOt4xVneOOtPGh8Ovoscet0k9/PQhfKXcQ5W0Ur9718BNa4T0tXLgPScRsrqFOLi2c6
uf8/vBOFV8sy94wIIIwn6O+0gMMLgyaJkd0ty/MJzDu3XGsmAzIQAA6s6mtbMtPzuyk/GNsimxFS
mgN+CuCBaNqT60KGE9h5orycFxDhWlHFaLUXA3xtcsUURjDtYTXaNkC3jSR7mGdt6sjb7spYpfFB
dotbv3OE1p2E8Q0AlqPFpjaoUjQWrZh1sYU10veqUAPLevDwGVL4rp4CmaRiCgIwMGJgm2fzUMFw
jOqxOB/a7lzkP5AHR+XSCrcrRLpLjS5+Z+Dt/HnOhoTfk+GdOSaFxdaggs4laK6SEqnWf2oHlcuL
3NsDIUlaga8khFT5f7loxcs1z0h9QD8V2CkuqCI4V5eSkCEgF6Rtw62hFuR5dVz2kCtkHk59MQ7J
IuEOKuMozqEkz1npHkNwZfzQD9Nnym8wCMciHO7eARrkb5HwoyX/C4O4sTcTLOHiBjmjeAX4e/PK
S0S7BvqLtTgjZbSF0T8/6Rq0I7gqB4CRowGEb2k7QZFbg3WD+lwY+54jDRrDYI0gel6+QITYSHqi
Zq4ACiFRGZhrSWZqHGA1i6bet4N8hyl+RrLb8ti2IaaKgRq2YQKJGo8nl+RmB0fGNJE6sEUk0W/C
CHb0a9sDb+2srrHwgHVo/Gjt7pYmnnRyTG3Azigf+V4rvObDiW/nqFgYupBF3loU23ZwDsWxDRKg
lJJfauXPKSn6vcTvAGPaI0F2F8ghLLEWBrIuIxbCs5edkMP9UCsfYelxFRfpLRhEjrlwlN/8HXm1
M5NIbAQmKsBWVbiLp8Uxee7hUYMGQtFwaM+ZxjVd/hJIEypWht6PzIlPa1a5pxKKaO0qXFsp7EUd
uMEXUdzHm1TwfxCeTO5KAbWcbRdg7krvSTsiqwrVI9glmU/veWtXQR5qgu8cpl8GXSOIiMylqcP9
SYfNVUXJkJ+x8qPZZFLyKf2ioBZ1tk0TJz8+w8N27+qiXsQXYMA0tDs1LZN/cdWL8+0ybr3kT6OK
6heFKxBfkGeTD2yqvL2hTayC7cs5ceRQbv820lnJFQK8vTWxFYLKmFBOtTAdyXHjtmgjtSz9CAqY
5bdTiUmpOM1VlU/hkrmfBkneSQ41kYLKDOm5zFd/VVjAXUlEnP8VwJJMh3HJqEulHcZwv11lekTv
DFgaJfp6gP5YB/1WGfcjewr+wnv7iG1e3Upkw4e/ydWqnHrSC7L+3S3qy4n+GH1UnedJDTzMCmYo
rDcht+AdojPs/9TgkX0jpmBpCZz2uX2COiUy+V3LBqwc5NC9OgKtzDkfAxgBJ9s61+Takq3k1hfH
wEPQFpwePFoGH3VnmLc11T/cj2l7wbWRKLtHTeqq3cV6TqhoLwCMmO1Snepte+lZyk3IuVxCGsiM
Y6oWf2r0V4AAr/dgcowURzbYf7YPIACthe4VNa+EGMAiWw9/a0naLQ4f1Ccv4oliRuuwxPJR+b5y
Im83uHxAtrTCbyH/LImWe2eu7jEyxS0KgJLBUyZ4xkovAudlJJ6jKfh9hdidkxO6Nrjoajf2rGCa
xbQjddvDgNuNydtGQEuqGGXD8Be40cLKt3vbnr8v+oaTmZORLU6sQ9mxTEJggrZA+8RdgEk0cfVn
CZsyvzy6a+Np746Qu4kL32TkVgYcfAgrJ76kyyCWYQpi5i2T+Mj/0E7gDOsqEZJorlqA5Iri/TE/
X3bfaeXwi7H//1vMSA3lWkFGrGugdmlhrOqbNZy6jFIxJpoDU6S3jd/PIVhQU4ZkvyUrW+eJQ/FC
9dLpTOh5s2sNJskjrK2ItFoDlazIaLyoXmpxwrJeTnSLmzBZbRbmzcc3MNTpk2jd4bKaSzQvPS6H
FpXmMNIfzVn1ZGlf7r3deOpzFnGX4r9UHMxiUeHZHJMFqlZBQXHbHnJxJk6c6CNSCjOFWLeErEPn
jdX6PGM/3Ou3DD0+6XQU0mLuEpfpyF2yTqdJMS6gL+OfPUfnK0vGyGxrU7oiIKsEoJgnDBIwwiZF
CCiS2TP4S9vM/JGUM0apksJogigt+pfqi1PGarciNrkJ+mLS6G9Ylr6uIBSe5wp4Ah9vXe+iNu0z
PZ0eoFruX++u5s7YhRy5PvTiOPTtgLhsySb4u/0oSmu6EqMrDife0Kz/ou1VLJQW8DzGgr9rcZ6b
//fKipDihkvvpPfImrUXKiIjJZ3QamkbT2heePPx1y9KRdCBLuEkBUVuQvMP3uo8EmdD9VPvY9ts
Y0SZigKpw/8XGkg8y3KB0DOWvcG9b0+AeLckDnJKgp7/Wy9WYuxw/HO7j5OL3Q4RWwatI4OhWSYi
wYgODTUB2FbbgPayq6alCG3z5n78tyxBPC1oEWXJNAMYBNpfjWBBpdAOg21NNrk+EymDUTCc54Xe
WUbX61BjzSt2fOkssmfGZPEmIYIj2Mr6eezEY/HMsu/BAUbu5Zi3uBbLsrBVDIjuBOfTLlnjnJow
hpUNx/qHOyf1cM2t0EQD89edyQ6bBAgXCTjBMWUJPjud0DOIauHUyM1j5BAYAwFHXRfB9lldp7OC
KACZOgBnsblARqvUT1Jd3Q5DiTFPy+mQxDUJ1ixkYJ70j2WZeexZJdOJagrZOUR7pYHOW89hQ3v3
sMpWD2p+E/n4RoKTAX6Y+RLBtbTGL6rDJyxqC9MP9SfnABmQRgXf8n+Nrm1Cv+TnitOJu7zS1a59
hHt20nHkm3pR1xCU4JBD+i0Wf4MVAzgJarovg+fXX24gCwwC98z5Vthz2W1ejVDx9dB719/4D2Xh
kHRNJqUI1G+J28nWyRnBM+RkXGybV036sM06nspWFTbC1fOTdW84XJUJZOL99ATtmzNlPTthJQM/
fAQJYU/rtxGW3ZGcecMbi62ZF+FBFwO4uvHheaH83Ye5znun64FoEplgwas6cAUbV/Ry6uiDqPGz
kf7xRian1/i/HNLXhXSe7QYZIDkDZa3nKwHpFwTVPqZsVWfTtW1BsxEC0FxLPmDuSLd7Qi61SqFU
ZJqjd5+YAAAUoq6EqzD2D33qmCiVAtQxvgrvn+wIKyBHtb0HmKXoYwvo2ZTXFM6cz2SgLWn+p5fx
IeNq4Y7Xhv/u9+5lmDJy++fY/LH5gAi9d6hAQAk40ymAfzTq4NK0wVagGHYiOmAMo36PT27WMTTW
vKOVzk/f2mlxTu87Ix7EOIpnXVzwtIaRgg9YQnpZsVg+xZJEUrbyvy9Xgrswp1FpKpD/sZbfq5Oj
nMh901i4CLVUTIjPQhcSmaBJu8UbFghhQgzub3W69GQXFt/Cv+G/D+tfxyHQjXQAS826sebsigV5
1MyYQRQPlfrBUVadk9OdIsAF40Rc5HxUtkFb2pMvX6B73Vhso9jgAMQozVL/0sHfwdZ3ipDFj8ns
xxwv3qgjQcqiJN3JLkn7Vln3IIRAuHqwS2P3vMwQ6Tnue74vGPJg8NQ8inG/PVgp3fdWJfNFJIQj
lnBB8IzgCnun3mKIy/DHlqZQV2uLY6Jab90qIoLqqZ0q/XX7/cgEX0Ss2xkeQIeBpD4TCqhxAE7N
Da7FeuFSpEROHtkfQrMHBKeVqmuIDmzqwBqaBPF55xHTV+g8g/uDrWU6XwIlpFRRqzsdWOQHQiSh
nqvznA1F+1liRg3CDvEbnSWlhfncrg6j098gdpPVco+nMLM5bLBuqlQBaZtPQuqT5/FrfQeGjMrA
COvsMDRQUhCdR9grhKUpYKHSvvrkLl/Z3P1lGFcwtheyno8vYNilSa0GeSeTurZTsvea2c8T4aeB
UWVd+nY4E1iTyCkm300xfGpcOYZ6qQoAVz1tf6f6FKmeY08nB848p6vqYb9uOPYNZA0YwEoMK6Ht
haqXpL/ub9PUlfCYffIjYg3KJIHyOgP1QGDtE2R8ZAbL3XnfGFOrJFevbO/XTPKKWBJIYv3okqu8
+g+zrBSMvB0c9rTecJ3BDqRh4laUZ4MgyXllP3XIjaPc30Kg5Dj2SNXwN+GrMv8VeshGAxcxSVP8
LDzWIYjlu2p1petN7T53xXxwGXlvjWJK3eSYb8Mt65OUZqYCLtJn25VskH519dmcNLYWP8rkLMQp
13f6BiXd+ZSaCJCgADyrg8+2xZWMYdOlYTaRALSp8boFNng078NGgHTmkZMuJ7kDhLDI6rV8gKMa
rNUpbxWbGl/NjzsSnrWCsRYiJVOHudYTaI6loo7LVlGZLsQKg/N/+FFWZvH31cfX+zg5QaTAWCMB
Ne01jKquETkFN6gwzOiVl0sV8X4fYiK6ZAO5TAXCpbQ2R3aPmAM+9DLRxYewpaI/hBPYUIg+XK1w
nI54lxjTxYai99I4BiYO7AUB9bpoSTM5pjWwU+MA+bhdgxuzgdRktSkoaSNXYAWPnLvFYok3J4rw
POIdJLvVulr4LuSrET5dJZmItgW1cbb70LAJ5zTN9EmWR64tYFdg8UJq7WZNKdW1lUz66CUJmbJN
Ar+zD7ZWTw1K7chQ40uMHDL1vfchKnBjs6mpw33M+Ued9zsRa2kpvahOweDuJZxJ886erqVOkW3F
zAOTrqgAG6mHbhHrJQUNQkDAxrFCA6it2P9OPKaiV4q/j9kekaw42IMPx/H9yIno6hN4DopI4yxZ
KDvbJ7nX+iFuEaH8pFQ4ekcVDAZmgwhyfWStS9T5w1pgjl8jPj7dVOvp/EZVJvcSB0kdn5jDjaFM
5A79rP6E4l8jXqL2kdN5CziMfpUHUJbMy0lJGl0BY6j/YT5ifbmLojNFHZX70Sfd9sJZyITXhm1O
Y46a/cxxyKIG6bLO4ccn2Hw0qrf2iuHTljd4iWTSKXBcaF7hyRc8frYsiab2htFOVD4TIdvgqq+0
e3HiATMzAF1RkkxU7seMiR3xj8cghzNe1AccqaUql6nIbWyCksmSG2+N815RXUpB1BpgEcQDFw/n
MWCkAwSUPRqem1a4o56ScfBUwWlpHfj0DLqTaaG4kKGzjNvsFv6/aQRIEJHYy/GPY1R43Q680YPV
36suLJ6XN0K58TNhH5Fpu3W9V/fm641rm1VejTB2wVGWS6lYDbQ7vwxGHT1eT+nxbO14u7Yy0QjO
ZdVQ6qJu4wbg2UpnohDp9q2PVC1K1ncfIX9gkfbT8oimk5nN+JOgeuqtlJXeHNcFk0Me4pf4xft0
3uEy/Q1kUv2ZsmEdxj6x3Rh7aVDjm3tYkr/2ZpVfsAvspk0dpqYkZQg6z0rSSFQRPGcRLMpAdmZA
PQg18d/GpePMjrIBT/9ly/bMR7eKiFIku1MbLzdW9cskKV2cDO58V3ZwavSgG1vyEyoYLJBfZnK1
o4b4ihPjbf6+iGtJ/CuIff4IEe5fNRob0OhxZbQH7sCyrAu1v6UbIgiSKWEANs77YtCGRXR2NhO+
wYAZTErDglPgIO4xbX7HI082XF07UXMA2wWclSf4tRDYrsF35pfm6LlZGMW6gc7jZh9Z3QlmmB9n
JhsBLRfb7jwSfN/YLQ+5h8Nkv3U6nClnbvwOureW1vZVSxZYJhNrABc8mEPgI719yk67YbMvhoQQ
NrE3mxKolL+L5mjXcftiIOjtUWTd/Y8tyeFXUxgfk2pACRpCrZ9orQOl1+L/72L5RLY+5t7xsFeA
3TSOYTb3AvTNrElMWUyXCTunL7O9kQhEye6KuyKM9eFi27Yl5UMCYL8lCc2tdsf104mMiQWjOjvs
S4vOmr9W5GHdxe/ehJfQyRkI7IlBrjYLhd/Khhsxzg63ZldRvHLgQcQCRJ2fxwj6BGKFb5CMMuSS
e60KTAfRHfrbfbq39gt+ZXYBT4WcZ7liFZEfwNXy4Zm65zri6KvK9cVh7eSPj9YNuMqP6txR8RM1
+ysZrX4mmyFJ96IG2zo2be9ZfYLljLg5EDX+BR0yh7faJaPGmaTv75tkPpEMKqBqvRB3aOEkbBer
NTXMvA/bCfiMYd/kOyAZPOV5JvhTjU6JlCiECX+q4N3YlRVVjgxcfL/AasGolomnsK4Ao+B2xGRn
oVk5JPRbGMExDBQcvZjcZvNmBv4j4otoCugVaS0oSKe7g8jK9BzlnWpPMWmUF4muwvocBB8Am6GY
0hpxj3EcemmAZvBOR5GPqBkDqaA3xpgsXiqcxy7a2kqwuS5T39JPNPY72i/uz0RA3eovQuzdcuaD
IurHwtptMrIsc2KPOfHxpbLdL/CcZrAYCAMAE+SKusJRKHilzMFK1AoqA8HadBXw/J+gfIOgh1vS
aorZmCfOYh3rdw5peEptMRrfhOxOeo8roURS9s4TEvpaYUakrSJztaPOl1/E3szvI4JIpz/x72FP
tP1V/t+09Ua9v3zV4CsaNEPer2iMiPxnZHC1NrtyJiaQHzle63WIEfYYT3rb6Bz5AnAERytyF5PG
FeD4pdtZW+p/AUZSyCMdwV5U3Ii5+yRkhPtJO4wDbh+omhPdahp2cBJVrAxjLrdUqLfM3HrzoguJ
Y6tREyNoYskleI6Ad/+lJ4vY8KYBdHCFEq9MMyrTk+k56Awh0/tkJb5K3MwqfQQZVSkGkKcvgycJ
9M1AQrHe0uRgr0zKU6UIULGzobLCVMQzML2jtSBDI4I9hiX20gEVPnhykuXYo/7LbdkCQ3gwTpWr
cykHWk/F/jiusUw6D7H9Y6rzsaNlh766fhPNagluQqW82Vo1zapXf7KqnWVY3VD7l3XjRaumcMnc
Uqk7n8vy6bBMZ4TpzJ5tGp4yXQDR4tBPDSFtIktRw5l+6VNx41jLfj9/RbkSPK6GytC0hhB6ee4i
XSNMtWsNaCT8HlLQXaC6+R9ydmWZDj2zqQ3wTq30o70imfKyPfPyw3UQhO4Aa9rUxpaMxwRwWaM3
ZojSkSzOMa47R0Ndo65VDNZ2lGl9IlXnxevDLTeuwNMuObYFb67ZZ2CvKrbe99JqBshk3Zp/pqXs
vnnYztDjbiOozlHVoQOpNqMaVvYSNkPRkg34xjhxoiAoh7ZHbE7SfUN73sIYNhK14g21UcH8Cd21
f6uUT+3ELD8MlF34u4Yc+WmIlhuddoxxvu5giaHzywdF2jO8NlFXAv5TPVO5GTCjKZvIfe6B6G2N
bqz4+qQeQf/kG1xVZrodOx9JIdZcXy29U8MdZcamfKW5wHX6ok/y+oexWgtqXx7Axab5EYxm6T0I
VwHVj9DLcyhyfhv7xHy2jZsp6xAdhA0ElqngoSYgWPusrC1v4a5Orq7I3f9MsI/66D+pqJANA9vW
JtiRbpXdm2c6NKOFCQRJKAxfqU98rU9V9DQR9qr2KsSilOsA8AEuqoHP5mmJzN+592Wk9YNX0Zrm
xODRnti40gpeTQNT073Len9bUGc4xkQuxW1nbbUgtQOAaWxHekN3YXFRlitd8bCwKB0ASkg2d2bg
D2eXloCIAUJB2hZB6+zVd5HgkM95Pk2BeJQhiw+UvDOGznk80c9vxVizl0tULtS6B+2uK93mSfKV
6+Jax/UlqyszM2mHd8+fZfieEV/UZ9fyVPzuJDmQurKhF0Vtm9kfmMIkTfIRo1J2XEt7fhW+zhq/
qrd1bswwW0zn+EiZZDFXOKWdLOF7XD2QVRF8EyMjTo/JV60tsCFlkpUgGEoxoIXkg08B5EhRAxpB
PR8AV0DhPZnSICnYIg34myeDjLmZG1vuD0pI9SANrcGOMnDw33R81RqGtOdXYJn9XneVh5tW5B5R
wP3lTYeQG5inuZ0XahySYPcy2OYXzHDJm8BjzST0lzHASWzDJW6QEJ+RZ2TGqrjftPq479kHX5EI
q41irYU4XS9W/WsK3uJJ7iZYZ98enRq2j0J0vbmsrNoS+a0mTZmi6Z1vYFDIu7+zX2x9FgyyukaS
lHiENvTUGfcqsEet+N3JxhOgm9P1gbuQumcoBME/wIe79iu6m8cQFcczYbNNoobrf5kO/XIaP/ce
H9CwDpXgPXjPqX65xw8nhVaAE+8TIudYCGv/kNXzKOcvUE7W+VAeg3V3UjIJHF97x7eSzHmT4XL0
4uTKra1WQvyGa/xsB+zpTn0eJENQaHzDOawSHJFSvfCRySK77jieSMLUtdgTzV9rm7PvLJEDy5QH
k6BHgCPwq0aV7nVDtn4/B9QxyqUy096UYz3MmI7UQrciBZBoCCd2/mlHFRzr7zAXptXCsjFVsaZA
TFpwH5QZcBeq2wkdMGp4ysAsec3BlPyL1MnWFvDU90dxLNOC4caY5gKPfxOrkZCQYcjH0dI58nRF
CsKcfgsW+bDTgWQ2+aGcwhOr1P3CF1U8LoFEuqHELky4lXpbA0CDsmwlzm+wU6F2sI2oTel52eIC
Vjh45dbnnY0c1VDsArwb1wEtkdCZMimLnqByQknI7m8StJJZ+lvWwzfj+sgtWJXYJSS85uaEJbXd
QgXem+4n2PwKmLSNbZzC76nlcvpyiJw4PpxedlWEH1VYOYKJpJo2/IeL/C+1xCxdnpwP6k4NFRZf
LfFArcaSdJelsikucpv5vEtzHDciuuB1XcblRBdaOy18VL4r2earRQYQ/cS1zQGbAKl76FA/z5h6
qvx3HzGAZwcUDqNcUAflJwFJkfKQNzJZaGBiu/xTqbfAsPIJrRuvk38vz6zdPy2FPLLGE5LCFh0K
5gjxE5uTAMeEdw3NKtY6Rs8gElsmW+8SxEQr/RkbBM2Kv2V8pwPnjfA29q/pzzXEqxDttXe2W9zL
HTDQ1hZuz+BfYjoBQsRPXGZsM6FYVZGYHYKbdgTF9UuulZxMwq1lyBwvhgiZyQhkPGlckTH2VR7X
Y9jUhVv75yKM0h9Xk/lfIUnjsGCZWqAkMsADviwHENsLysiQGgYWGRZPRMPgCWw/i35TnNMFXtkE
mdgD+ooJwZb93tPtZMqQqtfL9Y66Jl99nIFlsTS2OLUX7rFem3OlTxwzcBfQ5pdyLLPzotj+01Lc
ZCt1KLTyFLD0VfIIjgcmS+GbxHQ2LOigocKJMwTC6F9geJZRazGEbTnzY6T9Ye8YCmTvj+1JpX0E
dC24FmPivKG166B8oiR+nejP6Guwj9LKVpEA5UZIPEj+hODSPR6KO1fPtfLSa3F5+p/+/F7gVBdk
+GgJYh/v9zyfk5NvxcfYi8Rr/59nnPoCj6FDw3YpGNcZ4CdklKewQIrwgujoyPNkr2JuWpKlgHyy
dVwg9M3gt6UnlZYfxUngUcUCzyVpKSlqjhI/BMig1+/P4/Fi/IxgPWQCTXT0MmcTOlEGK9hpJaU7
1N+gyI1PQgGWXFoMIl9XlUoSUruMgVnrwkAXqecCqPTPmGc/R7STkS8Leq/4uJXHERDVT2wSlxgP
ct+L2to+HKHm4FTpYtsH1K+wooZzFG/gCEeuOqiJIGiUm7WyM2X+hfqp98Rke69dJ5Mz2aaJkONY
l+C+OKLsYyeCMIPMkwkGXFy+8aD1EoqrNWmropKPvnHY+XmV6fABKGBInoYaQ5S3D8pLtkkvSXZL
fZLcryASZlYnDl6QpcOCNCIuEr4HtZmu1O9FXrg7KqhNfWtWbfwmtv568KH/UVqXDHYWfs60ZCob
dY1wJs9lSYQwWlgVgDtflz4ICAgFKbius0HKwG6a/EUZYqxxgxb+Usd5TEM4OQ/b5DRrmyyTjEFe
wDh+F/5wrpJGfTnm+iz0KNWVwW1DoLI8oUOs/12MluQjgr78cIlXHc62HDLRxs3O0fgX/kyBwIDB
cEmgLeuFkmzcSAgISntjVRUvnoqCzpPU0pIvsrcZU1TZLbafD8aan0onNhomVKYXrVKaYkZtimbE
lWmvk96Pc9zVTIGX2QWxvYqFYj3mnExypd6gFa+u63Ynd9vsOIZQHLu1K0/SF40z+1b+ciXe8WwP
GB/R5aNrIauzT6EBqTUXVzt/ah7UmVE1VnbCqi2szuIOhLQ2riydhZkJFWSZ0Jr5SrJzZu3roaUO
K7VS11AmIt4CFOkS7/qu3du834tMuKZ3G07UsYZK+5XMKn7DWppGpwIJH1Q+Fi6DVBkpoJuomxGd
+1Snpzn3eT8sbBFN3hb9wabe79CrRN5L5mSK3o77iWhgFjCH0hUexTdC+1vIR4LSFyUVUm/kCaxJ
fCd/Z3Hh8p0cjm69VcI2mP8lf5AoyFb6kD+MYOHs4wEpAD5TIAUsj7TwX2sTEX2tS5T4V7zc5Lly
vRfL2UpxbOcyrb8xNqBCfxS4SEjhaufUMECNl+QyjCRbSMmdcWLlaULI45W+TSYiQP1aAy0o+2ak
oBXkGkKp0t99rI1p7Jx/2P1f6sc2Iti0P7yAX+CN0t9C5d3dsuDVIE0MzCRudE9iGp1ptEIMWxZ4
HrbHQ+FHzJDbgQZvg8ADw9FQpdqme1BF47yX4+It9OH/z5lEZj8R+A1DGSS3nlhRhil6FrA7ALDF
Q+NUOZQv40dap6+2XPEtniLSb2jNNt/wTVU5r4v0uu8HM8igGU6TopIDsi6S7C9OYcRXiu7y2/J1
BG/tc+92INL6JQZFRDhD2Thvz820XccL+i42xna9lDOrDtLEYHgT7oPo4V9yBuP0D/cLBe2XjiCx
scuxv+zIiKKbdtSAZXhpkxX0neQOPDODz6hgAC6cN00YfE2sxiw0PADfJa16doXVHV+id7vsLsBz
16yQGyVlHCUjQOQ0ipsTLbdRkEowDbpdLTxHdZaCx4TnzMtQUr3c6Rt50+hNph4sHP/iP3YW9Ong
l1kZ5fRUpOuZL4aJ8tIZzCwDGeG/CSPMcDpUmTG0veEfnQgMjMBVk7q/oW4n6sEpWHvCTH0Xr0bv
wSkB++3w2qCtr2LNBHevBrnT2/XQkld5JRJa4MZ7vO4L615ZAAyT7rx+ZBYrq067ax8iwlrf+GHg
P7Gor1TG8pnmBjqbLnzEmhvPCloaWgN6c0T6J4f5FipSm0SK5e9bMNPbXPtYiDeuht2gxtMdcBNb
ja/5Le0lVzLFR9ocLPlmwgFeiGPMYfHER/uOxGNIU6nSrCgdpc9siKfyEo3OqX2Zmf2j5WsKUIs5
ussBK1SjicGymemF/9TzVps+Ti9GUsnXOk8jT1vkB7S0lXEfijdxi/FezNVgsOP6jWdLBiNpR73S
3YGxC6Jz1xtvQ33M6WDoV9Lhb2L6WBu5yzD+PoaPq8IY7VB/Uhihwj0VCcSBHWho2afsMihmXwXr
rgkyMHhR4utzZZMFNYgbjtPkT+522bAiwhjjBVtKt+EfS07pqIxRNcXaiwOfZJPGINzOcgCUtWhy
XDAbc6r1g/rXvh486yHiN/uXIHp3+N6XzgwNwptoNkqoIkNrdhUIvkIVs2PhHPdus0nN1gYPr4K0
IveSOIRJCNFiQNWpwqwEtKzk/VXDHKaKQ+cwpPxjcENA8yIBT4PL8t9LJ78VZyDNhPW7L/D/R9iP
RBZRYt9Al+lIgf5yUeggXrDZn+ui9EeA0ZjJG2vC9zgnZ1u+70zsExQezsoh75YZ34G6TZ11AUZg
XvNAZUSe6MW4wX6UodZcf1lTCAyLqTrtTY3Ay7DgowJ349jPd9J+F+vC0YVPBnc91lVmCxshDXhW
v4Eou5HGzDSODPJ0QG4HGiA+Sy3vn90hkgWp1cOBRThH823yvhXnrqD5OXnd6AHvmdYldFrn0B1z
MORhTYh+OulM0DrRv2w1jkN261M0Vq3Mk9aChnJ+FlKrO8+jgiMiD3DMcxC60QpCU9XSQAAGFiF3
cTPE4KTsQVA+vKrC0t6Qq5AdvBksUx4pkK1bBVpBOSqc0U7GBwIpnk+lT5g7F6VO9Qf7YSLHMW+K
D86P1r34zRCrHCrBXETLt+TWIgEKonl24Ds4qZIpmLh9K0WtBwqVmzyr2oaZu9chSPxzy6eNqXvj
BrQZwaBEeXt108tXCw8ArygRXRmJloFesQQHz+lapXvgq2L0Glbr8ZpisehWIUu7g6ErJglaP7Um
YHvB7EBlmO2+zOB5D28TaScg+hLpEgN+l50p1pyItHqq8BD+qaD5fDHLyxSii2rusG3lhtd4zJv2
7IHY7VF7zk5Yqk/NgMw2v4X/E7ohPphLx+e8L50RIW3a8Nzl+OLyRGvm46Ab/btwaGu6A5dfw/5j
sS2O2W+eds3KBu6sjrmicKRBLazg6Y0p6HMjZo2olmbh50TEiq7msO3rM5XN+VBOCxnMzydaTOR5
TSMBB7cjvUmG3Qk5aglKwpxJKlCmCHZ13teRAQgmA5hVn4IpSyhQKvW8iiJqNpep0Zb1MUlqy76e
tcRG1hadaPJo6N0JZE+ALr73b+IhL4Z93FWuoHrq6NbJzs0GBJeRvL3I3Qq1y9a0aVJqiQ1m3duy
nbNnuW3NonblkWxriCd0rhzVfLufQUIywZvBHQ1zw4FF2IofCNenqPlD7mYvW706EWfDGevhPQm2
XnYCVbgdghnPlCe5PIUDpf2XoFHSjBO4dm+pEsLeuqd7024T17X1+8fzS41T8sF7KYa1TtgOExgh
ZMRDerZt/7fznWM6hVhe9SW0kd9AaUuLDL3qPSkiNtEVCsXvw/xr8kx8aV//no68JWAfmZdZ5RhT
CNi4cP4a9AMRRm92eMzg5eHoFS1TXcjGzdy8hVHOayNMF6BrwuIZmuNC3gcrJSx/j0jS1HGWxe4U
vUzBPTWVJUQqHJzLHDSMFgiaepjn5N1YsV7QE/n96hMoaMEKXdK65AbNS6bXWDvVg9nb8KEQ6Vhl
nYSlSs/+6eG9x4lMLfcYf5HKObuo1C7K1RSwGq/yqwbiTsOXoxUqK4SIcaWfZm201XD8rNlXHGSc
bf8IrJVOrhFLUbm9gb8H4U3+mvG8RuX4EAxhQwWRt1McXhqeQk5ElrY102bfwi1NlgiMhfUF2/Ka
Zmn0fHfUWQ37wl2TdnNVZlXob4uXqky3Blx7Bm4zisLOZye75sTcqogWwqzNzzvEsXSHbJfG7VLZ
j7wCDvc/i4qgByCoLp3+d2kzEXBXj4vbhx7PdQayWh2zDoqhJKfE5NfAyRb7l/N15/3vhktkku1a
W7bpKIBKhFS2NJ7G21iqPmj1MbL1n1yIeZe8UtXk9xLHHuQtji3Tj3jfvUaVgS52Och0aJjOpbJN
uSWm7JdN6zBXByDw7Zm+q4xceJ9w8obNCjmSOpjzmGpSPG0Afb5E+G8gaZUL+4Wg9ibB0+gmTckT
ZghdqmD+coLhdq+7tXi6BERfp2nTXhvCP2fRLszYBPhO7UlKZTo1zyhobj/lEVGQooqpC54AdBPb
b1n0Pr/VwEtWbzezNRc3gT28GfV76OiwCpixJXlgUDNc+bZnOUuH2LCWCEmbOFvSIrI02CoS+8Tj
Eo3BgB51FN668F1cPBLU9+MrMp8ar5M20BUn/khOSIFtPjQnbkJUruj8oxE2Adk1rhnAP7qeBoLw
NaTKTp3yXAv0XDh94hSknPt30XplMUBkJaH68YuuZFaQ0UkFqWzTULxaCur8Ox1GIfEIuAXHjh7a
fYBbyZi2ln36MXd8KBcNFDzlX3RMQJlEiKr+1eOD0h+P1/1nEKcTYPmhlzaNHRmIjswsoyQge80D
0VYdwZyKnJD9eyA2eZSXYMuhSi2O2xCAdaq+5JzgjdTQ6NWGeTo+1vjuveHef+CfhoZuzWuG5F1H
brDGuq7VEjGqK3MZgmngJnWNGytnbcaygYsg/sELMmx8s7Ez/b3rJ6rkfJoIT3BcSn5XiajTeeZm
PFzAhzYMGLpI/CXHk+Bv/I+MHdq/qHgg1CB1wtt5hwfN936PeVSt/OsvS4xACakwgfwFMZo+g0Y+
nrV5pIiMQgSRVdmKe9Y6/bpRkF6wApGOr/duT0i1t+F1CJ3p2VfX8ff1YxmzbIqNtz10etKqSsuO
Wm6emFNu9cUpKDsRYUGGXbN+dhfA/+gU2+6UNi7bCFfyPwjae4/a0Yb9a7mW7zxzjCRFv9vNAb3c
1lbkyMm4lxUpl2z8kAaI300vdNGWNY40Q4gAnbAifHUYmgHOp5mUoReUMZwikZTP0UizJhpfxKcy
ixFYE5hzdMhmmSz4dz0NhVQpht9csLZuoD5c9Vdj7q5clv0AwdVRsGPPDnfQKTCbHTNer9RJEenb
CqHgfX/Gz+i0+XlJ8iaj+sG7ok6r3m6GBJffwJt/L2KztZ7lW5T2xZUum5SzHAiL/d9T22lyTeka
bl0zZ78LmYLd62yp/DKhE1d7Iz3f7wofkryBdld8VcWU5WUbmFSrpOg7GQbZFvwlhGQuda2QntAL
w8ujKJCN+ZpjSlx8ODBQLpzX7Jmb7GFTW25SvPGtiCtOoTq2S4NdvIn9PxRqFXomacVei9JA8ndZ
5uztW2Cbpx1sdm80pPUBKgb5TQ8TjUZ390ZAxJarMcPbaAHUi8evG3m0maxlZlgGMfLParAT8Ey8
O/BM6rxs7LE9Y+8fHg306kbYjvl3lDJtrnxpPoolKEFXGvN+rETIEXpjKnZ3W8n3ShX1JlZTLYXg
EEnngwZycmCqgNQ+ndSAZ5G3rAZS65VKcxOoSIOTeLuWVl0cNuemZ8JSmb0f1rU4Cz9BPAUBL6dI
Bu62oz6LJ88+y7rpzJ4YeG47/+IAnouk3tY5/z1sWuL+93c3WnfAwJAASQ8PCUlDWAPRshC5OODl
5hmWA8X7Iy0xbgrQflrSS9lT+MUfi5xkNSqw8aT1hJy75ZKmMFBciw4+x3kUDI+5ktZHPNHuQgRF
q/5rSJ5yYYPK9LOiiFv82kR6TKhdDYCVWwkSGGn/SQE7iCErStBr+KRQxLueV1X2iQe2BPOwTbVk
pB0a6pyx9DgVgb0ahAyJIKOGWKy6psyyo+TBcqBZ1AixM1dRN0qxx6uUlZHc0Um86rVzpqx46Pwn
PrBvUAlW9f2jW6VKbxQf8exFx66d9RRCudrwkSnvBEO//15R91Od/Y0y7Z+9DDBdAQ3W/ePsiPZR
2zbFDDj+HVC5+3nVlh0gYzZCyQh6pw8Vk4FL0frqHeR//CEkU4AOFgc+sfKBZPNG/qsgBgPgX51e
Rhl9lCaftuXkki5MVitD56UFCGFRAZixg6CZQOffA5531EGdN1sMlB/Lp8Ly+T8gxeG1RYVB1fb0
SO/m+KKlj6jUKDj/OlHf7YdVra9XGpyHPPxu11kTJIARWgCiuz9pAOeoOsxZYurE53gxdn2RuI3U
48vXK4rwpFG6iiQLU76uLwTY7i7xvjaeguOR06mcbsL6rmLSCP+zLV4n7sLk9Scg0h6ZaHyQd0Z5
ORBPjG+ozGpiew2bwvcyu+9VU9/iDouz40XOvABNlJ4PTF9RLweCWij9QuTBfAr255X/HqJzq+uE
JcANA18jhOSezLhE52gi01louC7cKGyvGwOfwyb7rElp+MPDdhHh8PRQOlATh/m2ithYdoPSDi6D
geXOJL4Fe+IrQ4NAPPM/vhdV2jzrASX/hLs9sWvidqHV99W0FVVSgGHBhthhEeTHB1ElPVHP8ffl
bnHmzpo6mPGI1y2f2YKSkF9oL1zPcqAehqeycjnD2pzTJimDsOKW+WMSFYYSVBgffyJX8vMeSZPZ
8vjcSSD7wPr2rWPHhksrb6QwbIvLf52XgnQ52NCS6LHl9dLZO/XJURksN45mxWF4+YECkkR/8C+f
A5H1jV4KjWe4R4R4PPzhCC1wOYNTdB6O2P4ZSzlYvZZamHMBXq1foSgJiwJr9VnGVvEjvGA5B0K+
jmwiXCcqQc1wdihgd6sYVXwFQi8psfxUVANE1s5maoG6Tb0NuN8av05767Xhg5zADtS5VP9gyCRR
0WggLNvJD0DiF547xp6wKyajOnjsIeEGlxoMcaxVRxWLgJm/0lhkaDivqN8SvDsE0yg5Z8qOqacd
frNKZIqvn3FCtfiwYEJBC9C567FScM1iYtcUqemGEGfN3SNb7OoUuMdpqYU53QwR+Vs9XY/TZ0Fz
I/EbiyUZphHOaTKKJgyIEEvbdGH9X28I2iXENZ2QyHkE53rYrpklHQlhkXivfsFV5cPNZlwQ0p0q
QEe1IyH1krzmiT34bEZtJgy4iglGAV6MzKwdhSPoJrp4oZNKx925MZ1oD6fpQcF5GIpBEFvvZaRO
3HixGbW5+xYjs8PNINk4Y5XeH4juxKTUezkFuGpkl00o0CGxbtZF+w3S4LCMWKw9SA5MSKzfbCXt
kqzpF3EcB2JgnkZxsWlw3a50ZbYa60TPH7Zh9jPlWLVY76m3CqPAHcME+9e8SkqcfVuTzbv+Sk/r
oBb/F7bi/4bZNYjcOj3HqR3cJsG73YdkVzyRCk4aKK4idFGwwlD2fgBeWtqsTQ3Wyd8nzipa/o8n
RAO4HWkA6+XT/UlGejghiiWdZ6eUko0W4DrhUc+o+os2f2ljTfLF8GWEGkExPZ4eRML5K34ae1OU
3Mq4wHWOM3RJpGGBsRmVGm50cjmgCL7yK85PG1U71/X9CGgctk+n4O1y6craHTRLQR4TOCWwX+xh
mLJRTKr4lnQW/37621aTUXmXkFdLdvbb49C9xoYbzUYmvTfJx8MIV3BzFeg50fDYzwW6iQjF3VEq
/b60D7pRfZsPFVwGs5rm1UQFXJGUHd6P8NZ/BF9WYcruWdJYgfV3QpeWZHdd6VQbNAB9KnGu4Sv4
81yBv0kXiNnNO9bvevSViiTebv7xJMaqFIU5qu85Q2POYXh8v3skAQG07a7qvgBJPnNGywdDp0t/
AszT9RRI+dfM0gVUojSSbyjvBdBOu5WycTrs51vetMyUq6Rvub2uY7orQ6Wd17mby8cbK6e9t21o
ivDdWqkjN1e3UsVNHpaZeBKBPU0wZjsT2uPmk8Bh1rW2WrNI6UR7/Ca6MeAhoBl45C4Mpea90ZSl
DTsuQ+QQBHkyeWFxruvBj58j/J2IVr4JD9LSShU5bIf7JgOTh0mjRDRYeGCGWMSSMKxpTLoZEser
gIZLg/ld+VOYD6wjqRQSKLuR4mHSP0M6mF1ZDqgiaJcXUjpnVxcT9TMCPBf1wqlTwrueMimhlN9H
Agx/nEI4PMjckrxQl9OO22HK4l1E0gEuWoNEes33njT+zZ5Y8dREsbm07ym1D3xIK+i7kUZDmahk
gK+4TaD9zC7u1FhlMK3LsyZKd+EdAR+UXWWLbPNFYNviygY3VnW1xIx0leFS/e7bJfQ6VK3aYXBc
XFPO4+92zQf9VNXgWh8thL8abf3sLHtASMc7WSOj1hSQumwAdHzAYf68AqB7UeZ2VBdqL1CezQ4V
uniT7x6KwGVNhIDU10twXE8I571yQJaEwc/4OiKK04vM9fhweoBHLfATQ67DOGiDQrIJxi4agS42
TQukkNKu+Oe0xuBbMOTCmJEKgTqwmb5IQOsiQC+QkheF0FoH82KGhKd47j3nI/mlVNcjr4r2+6PA
m/WJ1bOnJudSkQbrXQXK+kroY36VAi3NpnS99jm38xbquwlu13PuefK6dRRzMIF4yls8T6cDorVE
MYZTA+BHlUwhSPSr3FlWF0ZPRgVR5ds3aO4znVNz0f7irc0EaC2mS6bdHABL4qbuNt10CURBph/r
W8iliggSCd2mign4fVbEOUncjQXxwFdtGC0CQcFXZ17NJJ1YQVAjsW8bvWdYTWMXnkG2JwAJfRxn
5BsGOEYX114zaaSiEGQPZ9eyNj23gY0hqCqYg10VjweKypPre4gTDoDLxUHT7FbY8WakWCeAYt48
IMAYulif2P6pqdIoYz1Ov/Yk6gX3vdK5n2rYglj0MH62cSIbl1OJphVGXYc51H8opuQRIIRWhvay
H8u0RaeTLneSkRTcnuQ8oraC4iwv3tLftyzSdUyW9r0lZz7ijPH4ub2wkHBwx7Ws/QdMsU8H0o2+
RBpV+KcmrNDOxmfyuI6dJK3N7g/5TNGzqzKzHuLnMgvzR+nKZYnVxF7LAqBjKv1gLcq2uIP3UZqK
0PnMXTX9tREnzQQf8RYn5nTGIfqBEXbtfSNM+pgDlyj+0psOamyVfU/Rn2Ixxi0236zHSSSI4ACY
agpMqb2ysBK08U523/qucCZcx63NwUendGv8r2ubA1IKYozUllUsx1ojGoAMnXIZPaXQfaXG3CXY
8ifKURF80xqymezOosVOP+ieCGbEYdSFtGr4rLVNBDhnZG1PPATts52FKgCW1nIkUF8cW7QL4fOc
qNI7+Tl4elVRYKE2Yq4IHx7yVw1rz1UL2tQ6endFPztay/8s+3tXTnMJ7UGhNN/uREsz68w7yjNu
GEOdseQBYdIEXWFGDs6cClZeZuqinm8ZG2PUaSZYfsVnZjhrCPMcY0T3QaR9ei07xloF1N3ibSwU
fYpbbgYcQuuwN9gFLXYwOAZ5YVFBfi4edq26lAl3Qj+zIgH3UIQNBv20qVXrAm23r9h3giay4v3P
ubfwPDNlhEgYH95wpxWdHjRtW7lishi12bBHuAPWcJoNe7ZrpIR/RnBk4a4bR19/qt71nVMIJeI0
bwxB6cQHuZluFudbIqF1D/JZzgI2m6JzNz4+um1/XlaZHexJEW7n8Gm1J0lXmh2zz5xMPy+pXBag
gcLlj/0W8KhySKWgkgt21IktlRFZOV6e0ymIHlb3x970llMrhNpJIMMfV3NTr5A3MPRifs52TfNH
4NcvtxbfYZXVsXvL1fz5QABnpJLTAmb5J/sK/NG7X891cHYecZNwF+a5T43o78tfFGLbHoFZgfax
kyNqLHTfAZPnBZ28RLRIbmWu+fLriQgkzBt71kcHE9CHDW7V3N3rVNMQoM5SKvLS8MJiHXp/SmOy
YFiQT+KDgmy2ANoQn8HikEQd2tQgrLtQF5/CQ/TEPDrL7+CwBXigLARTYTahWzJUN8sj4jTKA2Tz
8BzwJNtDTC4CbWHSBOY1f0f8cRTEIl/YYrzUCHbRs990YQQ+BkOI6HNRtyPoV8/LymKkyVwakz9i
6n6gdiS7wgzxn1JnA1qrjTakDH+TrCuSA5tjlU6Z5zJ51kpZBh6WYiOGeFo6Y1N376F1cOsl8npT
GT3diFyQ6ufXO1MJs2M/sTuWE/echWfNmUyFT2mH7rIeZZ4xVwU8loW8BEwbz2zuL+cszDFqwHLa
gtaXvyUjVe2pWXUsWieghG2MofiMws3yVDib4SflACGDNJR3WO8De587+owA/bE7fBmc5bmAT05t
JB6QJ0gyFtrA6ZTdJ61vv8/hFI8w/hrIyILPmNDHLHfvnPf0oFpmGzbKVoYLphJc0Eouy9RPl5Eu
n4agkz4cnrTlrtIx3e7dY16gtVR29E0pk8ibz/gLCWAQUWDLHxF08tXdOZlowRI58280acpkS5IW
VxjXawUzbmYNL2swKiK2WDZE3NVLT4O/1QDuk1UtS8IX8fXWD+zLenG/icd6gvg9/6W0mQmY26bu
rL6LfqCBQJvk5TFtz7i4AJSnBuNH0RfuL4QLy9KHgNsYa3iSVuCMKmH7N4KN5VViayXlXIezYkYW
oTNtLrCf7l82F8dpy5bAjH8uo8puK3XP4jINtF5zCCVlTZAAlUjyGXB5Qm1B8qNLBzLrxefpjWeO
9vr0jI86mnPnMfuqVI6ZJEYLgNWaGHZlLYsAJ71AphLv9wHWIKaNWcTGIr2XeYSlOyDv+9dPOTy3
e/a5/boYhVYXSm0nlvMUNApy9CnPRFWrkwZuDoBqiKCTUzCMBthpnFrHZHh0yJF+yoYqCOIw0QGE
0UXoz9oxu9SCHNqFCWURt2j58S4xCIQsN60XoQKZAw8QyB+osoiwAtXEmAHxc4NQpJPpEN2PZT96
+KOVmC/KmJuQI4M+0e0cKiK7JlOE4mKiRVjXOt+IHJFCNvVeZAWMuudRfG5flQpFkm9QLtEI7Y2l
SfXrRET+ozvfIyxzfQbvu6ZFyt1B/r/YmDMV2Q0joBN1n/eYlWhAKVTCV7f01o+G2TMo8PYE1lVw
I9e69bckdYhhanziNby0zZkPkJzbJ8c+7iLBBLYUREOv5pQdfbWkzQj4Kohciktd1qskWvoFKiu1
YztmP4h9n/IQaNb2xeN7EttL5sjaNYgqqV2FKOs11X8BNU9nVb8rqgGJTBiwwRKKqBMj+sZjcU/5
nGpCYsKz436U3mQPDeToI+Xiy3JgCAHH1RW3jCVlJkS4N0SZdD1R4BM5jJPTaBOvmK4JLBZuHMiZ
UWDck4PXN+NQuLj/PmhDmmDinHFho6lQBuFaVLUPO7AOJVs4m9pITu9pqPvVB4+cpLY7OTLpc10d
q+VQTs3t0O8nDtfnikgLJkRRE+9EG3q2YC93uiQF7cXpi+LpH2jCfS5no/QzHmNKz7EarJrKpjmA
OFshmqLoXf3S4vMjb5UDpe/0Cxa0uk7iAvk89J65xWduDXg3IPLYvCkBZzGRaMpwjJfC64I00Wwv
pc9b/SrA9Lp8O0gp34Z2p/PpIFxUNGBFfvmj6fjWX1SwAFb55yZx9kPsu2ApzZrxRU7Axgl7iMCy
hISkoTj7BsWZvzU2QftpHBqbsHZYPgiSq09G02+W9Nt5pFUc2IAtms3Qve1SLknD6b/fTPUdHb0h
DwnBpUaASSI+OBSzi63kvYu0Vb04kbx5yx6zEb9uZ9m4/HN5JXjlNqu6ke9VXIq+eVptuyUIhmvF
bqFbUmxK0ETIeKvnQk+tWXZiPj0ATe3jFaI6Rt+ucJ0sluAWlZPfdk8PWkqD/2lokmwPNT4nwilc
w6UOzr/MTuNJK1P1fU6m9AY8/tqXESpHT3p5jRrppb10wcZqJL/x+GLMo9KALQDPsmSYTlo8YCTD
VOAenTw6kzMbAOys9IPye1wZXpdc7V6KlSup8wJ2Dzu3UpLwiBMo2QhgDDGT+/xqPjRJEmcGd6dl
zcTltokS3dr9mbKGRjKzFmfy4gkKu/8Q5/qkykOA76wKUwq2RXeqxtFXLrqaV/NuWDA/blFiJEDF
+NxqBwyNon9iHGM2AphYDwejmIAy2LcV59IrzFGn5MvoNG/a/jjRwirDEh3n/3UEphc8tHBoSvr4
esIj8sqgbr67yklpRtkaZr1BlRptfgofqT+R74CL6i2ZPKBlNuo8WomPyC8PahrVoldFyCu24xUU
1nJm1sIPRnBAJLdyJI7m6S52JW19tN9jDcdLaIm/D+tA1NQpcCY+wJYuB6KU+hncjVzDw+59iFZ0
lw4WJ6CkpTuhZZMCZnKSmuyQIQpX+TyU5FjEZZ50nEQCZ5NmL3+EN9rwFo2lIvrlXBjVVscG/kNx
xM2KNeVKixf5Nysu49Ggc4/az6SE07GtJV3JaMB430+w2DsySOjQ0UoffTO3bd4124V0ltWuskJU
xErT/izbQIx9p7I1AoMzrZmCx+VDvRxdgiZKcsQ0RJIJHdJ/EbKhsXQrtSy5vPsjufIKe9yjzqkd
KBc4N5UUHmGLMHZ6r+jyI4pLEjSswo6LyxDb8ckEfCB52GAPo4NSXuWK1/YOBVJsMOX6d2vlapBy
12gWPScUji/aO1WDRe+9q3yDUfIuuebYh0IioaX0m6ooMyPxJrFPelCyG9sX/2+QF2+SD+j/n5wX
Vv/kdkqnGeNmAZIWwxw82h4rQsQodKuJpohPnBRt8//Flq/piSSL4ckS3xlF4tlm8NvDVg2U2T2Y
p+8oiLtixUsQHNyzqJAgVZDW9yNYWxmr/J9G++HMz5vRkLISHht/D9CTcNZZO8nQFskYSs4VFYZz
VPJjh2GB3oKvoniARl8LukhrV/nlzTWEuGTWZH1RlXd+h4mz7YEhRUiO9C/uEJ11CW6qHuXVSJYT
mM1952MJ/Crp0Q4yBlTYU//YA65OFJgW37ba+SUFbYwNggHwXWLw5KBl9aZiPulIp1BBn5blL0mf
DhnvEkpodlOa8wE8H+Vr0/oRhlVm+e9ZNy+l98veAeXgZ8efP7j1Xlcmkonf3LpjJOrEeTD6babv
1i1ItFH6n0IdJJFkcAlXL/kxutFSr0uDSm1gdgq6p7PZDu6wNowcBZC37mo5y7CZJFZPN3+685Lh
wVvwEIlP15pHqB++w3DvbVk9vaA1sJKm9MB+6gru34QHzgHoHs6pCdLW6XsSiSU4Cj+aSC1oebz/
xDUl5q8iF3ET2X/BKWoGX/LVENZPi1kLdWBX5EcTQG2qyEVT91H+Mn+VrZwWsrgBBIgT1exZygPA
/Yoq3kbJNj7yyEzyY/M19YAaex9aWNO1BhiTk48G9GOQXmgFz87e5oz90k3icZrAXuQ1vdfwXZ8T
B9b5JTb8KN6PzxMEHU3ShPNWg8Mr/Gww6bRAtkDVNW0tp21vhlimxisWiBvxMBNiLeWFuqQcBHtT
ivB9CEXFCgKL4OZQEpvsF7KDk+01IthN7lF96nicT3KIEsC5ylShEiQfvqWlh801py0H3LQmFyAo
aEBwNljVyziVvG+c7jjacu0tQZC62JP4KAUcyh6BTIkPIrO6Nli6fE89jCXyF5B3FP5Dp16vxibW
Of0ooEkw9w5/k84sgGtjPC0FG/Br4ZwTHUS5fIEvVQVO1sD/b0QN7zVMDdm8yiPrPfziaP34rR0m
ohQyhYypcUx/dyOIpz5mRx0Wqluc4o3W4d5fFpSvn7aZzPH1g0CP/sSSflY6CGAh72tFAzspXv8z
XDLE6YwcKkaeSwN6e4H8Yy4oKpuE4TEY/dYI9CbsNWITXzQszacUsIEi6KZIaVW4sFIEWe7Xnd9z
ge7Vxm08jrZf6zfLL5/zszGWXAwtdfSSpyeoI/r/AI72gScSNqRg+w6+uxFAi3nyV6p12dx6FgTR
201fkSYhM8C9NEs5jTlWOeK/nLlrZUkRzjWQwVPRqQuRMY6p0bTfCO73/2b3WmbJ0cZQod2gvWdg
YzAAyxKL9JVzaXBD9YuQdEF5hPApENTx8sDRowJnkQYPgcZb3fn/9hKldM6iKiUHw75n0Bs8JCDE
6d2+UeXsDqnzE3r8L8XygtTQVaFzMZZnan+KdRocDd27SthyOhdd+3OZB/oZwIFkYSi3NR3PSAPP
3h6rBHn1OKIxuXCTYN3K8ifddgWBtKNVPmrWRwUU8PSyBo0Ba+J+C9oAz2RfILJPD1/DngB8/7UW
/3rJxJGt1B6X5oX0qQzgbcyxaIgDIs8Ztxu59JQaM0WuLKM8HVeSnT7femiSg1i9dDiU8uYi49OC
1ZfwxLx00RM9/Y8Tu/bQIYrs8AF+5FbmEUK3UDbTpi8I9NPSzZoAnFGCgDKaACi9Dy53LQOFZCuo
6ZdE2TY+W12KaXremnMaZWtWvGNiKoVYFc+EgiNi2gagwAPzmaAbbkFCOw5qLUGGe9YoIbLoxUhW
IneIX7YNGrqdut2XGe5II/d/wbqfXk4JNABUJV1h3+owLhJrjG9c8EptzCqKFVtJtadfZ9IVIm6N
GA1Cc74gw89SeAcqgvQnod2lXML+6aPm0DKxTKvTPfLNLR0a5JwTxWKXG4yjYXPfxxeK3z9UMJ2A
FXzgjfXZQtQ+bcIjTCOl/1m9IYSeKIhKh/03bFladb/C8UUoOIloARJm7XWvxKlgtx/by/PliD6R
AqZ+3w/4bd+V91rEelWtld3KCrLwDIZIlAXyY9wX/vkdzp3sP6VneqDOXkVKDRHVqj7KF8ZYZJ3R
njT8Sl35UJEtMhQ0Yq9HFR7VEiHma6+nIy29nxCmzikKnhExTjGfWce7Bndog5GmJERyyli+OxTL
R+wMMstFAl2fZl/l4OSghSreo5NVAlxkjEMnIUwyxCtWpgnYcC68jn5xPOzO1yy4MmYFXvb+C2lc
A//cwkVV6rzqwrdpBA89itjz2x36M/UzCLCKiOccFiaQW2Zx09TSBXgxdnt80EhgAH/xpHtKDr/u
g6kSiKvG5duAsEvTx4kFLqLHtomveLOHrVvYG7g45T8uqDVrTB15kwFOk3NRQKnYhPERVHQMLJyY
Kp4gfeXr+jrNehr0BWk4cOwDFZFWmakYgNmU8IRG/ywtrZhBxlTp0EJ43bAKVNQWmdTDWRxk3pPw
JZrnza+sCVNsY34MA95UZyPING5sVn4DKkaSNtLn5x4FSmlpcU6LB7jiY626hfGAbHDKXR3qTW+G
SwuonqDgTrPuLkVy2RogQh/DoFYT5RrU44BO3vX54RqT+z0q3UYk2L0pJOm3SaQpmwmzoRY2TGa7
LySVaZovuNbUpr0h4ZnmozLYEaIpWSHe5rW5Smyi/SA6Un4ca0fWr2L8adsfGL6s2Db8eECzfpda
OpD9VVRhaM3jpVE4m4ivZianMNOut9ferrAGM9+ePIRS5o9M5ViX9FTkmbuA5Nm6haWq9r2+1YBa
jgxNsJzg9UwWpxULpsk5UuCEbvt8mUdUkSDS2Gs/c22VFPZyOBK+KA6GvPu8IXB+KpZX96z+Akq2
ZttNDFYwr8LU3g4NMCG4SIYS08vr4junulWrNXVZYLH+EZBthcX2OS4876goRBCmwlQghTINYeWl
nn5TZGQJrzMYxjpTSkVK35xDLN51ft3tD7YmrJ9SnapIzwtNts/2Td322yV3Ww46JTYywBfpFaUJ
Sx3e/8jGb8gOGhvu5exn+OG3i8grfxMfGRUN2e7Emxp9yyFU8uJxFGGIIFVlKqaxmP30psWlFLl1
p8l2iE4GqCkbiO03awX2wa9ZpizEkNVOLu2S6uA/tQ++DvKycGvcQpyIZUbAbnO8Bvib5rpcIMaZ
2pa/uuI8lLgWG3aYa3hiZayXDAGaEBAO7dsK0oDR6M28f7YYmRUVgbIH6Y98VL/DSp5+1JNnALoK
i+l2oymXJpZnIMSCcs0jXySeqn9SsUBzH07IdJtPhtVUWC+TZLN6gvC44CDBtjpoUqwSGlZ63+Lr
XizJynX9zSutJIk+9yU8DT52klB7cikqOaaeUOrAzfcc7iTol2BjKU+dRxEeW37x3cfJgNdi0FS9
AMenrj1RxakS+v6G8+lrJ8RmiSoBCjSYfkc5mT4beBQ9UMyE+di1HlyCINC9sn7LdXsq2KjhHLiq
TKo/XAbrE3gp3+5L7cNmxcXLIwVNtqBvWfxoim12heTlBJij3/E8/zqc5Xy7u4K9szBjPfQAtitS
3ytoY8O8/mWUKhAMkyDHH4kyMgDP6UqVUghbdPqPQBafM2JKSESoNGVoa2OcIO8fWVpNEgRiihut
3o6lAX/y6Q83Agz2K1LdJ/xy1fd4wcjR+YDYbRdThUXLNuQDOkLDTaNbhs89QAqbUoCMYD0Tx5pb
Uw2kwayCaNHR70htyMRfxzmme3GJrMgHKXJjyffn7fGvEg3zKnFO+9fHq8mxmFieRAqeVzZ+3cYM
ktfFYo8utnS4W/nyQK+xCP6Pi9gMTFp5OeIkNKxwTtRLabMgQIEf9zmnrBGvkGpprY8JBRA0IqNl
iAPV9UyA0Q3kA7Wew5bH2TKbDmIh5sQVPUxwTnZ4L9BD8gxpEhjLH4+lbAnjw89GJTqxx6b36d2v
BNXXYfVRwCcztvFNGHb/ie43iyXIkW5Rb7JzA95WlQZ6v/JOkVmsX/NC8dcfp9NTJOYnGECbKnQI
941PbeCJsfWhPuEqnyd/r14nH1pPD2Y1tE8a3rsEobvou4rIEQgyg4LrJTApVrNLK/vGsCANYqQQ
P7FuuKiD1Db7JKIG4BmHMgYR3qkrjz6vXioKR2Dk6qLifaRzjHZ4PAdVnyYJ5BnykI7q4tzX9/BL
IxWnkxrofqELlJ8dvKtxbaCW7Nj9VG1Bcr80XgfyDwAVosHuwoG2FtaA+V1tUcgi3yoBv/fXF/0U
CPNa2ln837Sg0Mj9VUZJC+rTVzrkSXvzQnerjZdR9odbZgytkDe+bs3HIm2rPqvtt2XB5kB/Jmix
JbqBT9GWvZveQQt/V3bJ64Mfmkc/m3eIOMKceZMzZlwOBaKDdt3RvNTLT7g7sRQOOxsJoPpniX2F
osqZznruhIoBzETfOmsTqTautpLxBwGQtU4CwDwJ1HC3ZRy9GlTG4pEPRD4MlooSI6UwqziS6DKr
+3XnVitp+xUJAUB7vvcVdJXSVax0xOIZf+NNFbTRK7oamUCWW/C1ZMKUQoQN/caLWZfR1LcVpwGm
sozLAzouUutt7APIu5EHrmFNrhGtIGHRe/Do6K6FhNx6F2DVJ/eX7FGXxY3UZEyb6cnT2Mk8oKMm
bTk1lmOTPjlk5qxkJAWUf51QFau96hjszTuSYAD4ucpcr8gchj8ZhrrpJRpUfBD3qrsUqk3b/+5z
UBXuebdD3sBsMavx6ynqpR3U17PNRDidFILQXeLBgyWq5NWFSdYXhWfPs8FuGmf8rizUa2OplULU
gmPGryFWJIUsG8PKC5o10BIi/CIaQQ5QSpfOP0tY5u67iHwXbtaVHsEJda5uWa+d8tj1nYsT2ZPH
DuN+QDlhOS2mVIPftifzafNB0Re9Me13WSeJ56o5QKWRXG1sUuXEJTUTIM3zmClDLbFqFOvVS+YW
EQQiwUPgL4fuwgiGpApO3+vAGeDPwwDDUUgwCdjXjehZcWocp6RbqSh9KmnnRiPIS3uLl/LYjZr8
i1Gdy/I95nBBKxgJa46I2kEljOcnvqGeHrlhdXQpOLsv7KNI81UvQCp1NuQsGGWo5YYNda4Zt0eh
LNUiEA7mUnm16VnU0OuP5tyoX5M45rIfhmW6FXmY0g63tQ5jbUIiv60Z5GJ8jh5CcvEWRoopHRPp
lcbKsRzK/1J18Lngd9Q5pNDmXlJlCFmCULCJ8Rp7b83+lEuaAmFtuv8GUCCSjl3hNr1eq8wLVM4Y
8zOpYNgqWYdGhVK/aZ1DSl1blJFDAMnJuo0+C++CI+e/sV4Z+vo2wnTAohaJ9xEdLcvLyevVgWfT
8MWjwsi0zWdET1EdWRxjgtIl7FzfCJ7PPLXFoCLmrlzbToB4OUWow4BzJjF2C79Z5E2pMq5wI1zd
ekMD1fCf3Sv3PLtjvLLp/lv6CQtfq/PtdPV4SoDuYT2XWWJtpq+lGIoEVRvxwCg2vyxiedehvJBd
R9TpqgOv7DpziQyRliQCzchXUHqWiIg2RR3pyBQcp1x7TLTgLjIkejlflYlBij+urzfz8rzQVR8x
r4bteT/FeXiDn7J0/f/i/Y3c5GNTlQ2oAERmq4KosKVi9ilPmkrVHFDG1VribfYRf55crohexcDH
TYd5BXHFdEk+B4iU3AAZS1QF+9cO6X2zDoaDcmcDspU02Gm+l9P4EOwqlWEqRMD63FIR3V0CbUIP
Twf+lVZBTOiDIUbyfKgRNeL1Fv9E3/MD8lIFE765QuLIVgrTLaq4/FHsYy4sPWD1XrnA2Jog2RVz
AK7KnTlYJI/zugv8tZ8g0T5llFn1paP2ZM7X9fwCyjV1yy5vMkiAgGG/MAS16L9DbejTdbfYN2O4
TI9Da8hrEUK+qZNy8vAzrX4lO3zG+BG22gvKCKyV8nZTL6l9s+53ypWKQwLi1fsX7LjLd7SRjP7x
0Hgm03BcaltZMVBDay3ewceI1YJjOuAl9+tm5wfS7QkcE9oZKDxQChDAMavnhp7m8062Sw4UloNT
5FzrlkiIxxHoktvgp5PmFAIsSPbM9gcXF7JAImJ0f5V184ssVEGkXoFdjNNNfE4oqr4SxUYo60Up
e6FDNKDr2O63jW0yB1DIrTB0r3yODvQXFgBjBypChS+mkOYTkS8XLnCDlOsnoHiQ3JZkvd00HogW
vWY2tU7kp+TDaf+fvb1VFppmWA/qRT/qqRpHBOCZPattcc6CvHflwNJu80ILCK15tmbQJmRPmMW/
feqQlRadY5J+LvwAOYVe+ZfoNbHICNJlRUym3GAdFKFU66MvqYwpw4ZqhgSHy1nr5Tc9qXspxFcS
fDmOoVrh9lLL/FtU+lRkZ52IJgiBjVzJdxxiibt7qFfDuuG9HxLcyHtGEytH4i+7+bhQazN3/ok7
BKrxzxdZSAMQav3dVvQtkW7sotEU6rBxMNrUS8YHAL9zcFYjpVvE+AkD6bDL9kuhJA55t0TmX9xV
XyM+BUokMuOpIM2XunR4qsd9p1q6XXcwbIzeZHtOQ77AercHQHN1S+khEid9KEj73KZCFThR1G+K
H9NMrrpubbv2EfRIllS8036dINCZuJUG/vGZB1dDxiCTVpzfgS7LDhtbDwz4R29GwoHXnCBCc+kI
x4hnLbWS+86lpfeS4w+F3syDRXb28oEEAm8jrn5SjcpCYjkOQuxBBADErx5r/YPangcNM+2P67KR
eUIQvIJDjcUkTxguObdfxc4eR+YicvnahrU+zsUuyx4cqpMk/1cVJVg/XQk6BMkKqax2MRHytPZV
u1nzFESksOsMk+MXBombUPA+AfxKjDqR6o5cGowRvSkFcXN/2FkxFfZFQmQuOxYKlLecanX0S6Tu
L74ff/PiDjWBljMCo5D3xZ6Rp0fBy7fvNQQUQwUagCo9ASVqn8evxH6hPhyQr9u/jpEFVKPxmSMj
19Pg+YcAk6DRcb0224STII+NG0mP+WYL5lacCKdlcy7I4a/SblAS815DgEtK5iuROFZBUhR7QVfU
VJlJBAVLitX7KnI6ThjeouqgiTlGxKqieDz9y7k/HFdDIencrh1t7AWDltv4xgo2Zec/wZYnxUmS
Lbpkh/unqnk0onB40mBLrRMRTdsQn6BN9iS+tIEiF5c0cw/WKqBFC4ceZlbZPTlBVImYIOj5uH/W
0A7woxgr5DRITjsQ78qwYaj0ft4aj0DWUKBRzBU8neKRhCnT12QDTv3kXLFkcNs1zWeFQjoZOOgI
l6nc3xUanARdWm5vIFEAyJB7Zcg1j9jcGXL+rKoAYCbhOGVEwXPTINFLOaAGAQudDjghFUjEZpOM
cDXAMBDoD3d2KuoYqLhkqGMCwpYCayQ4MyHYWgjv8H6ejWGbpGdDMgUXbSTCalu/7CP0S/7u/F6D
MRa4EMHLdZSP7F7j6fJF0UYj2xcozF8bVltpSdOwkyBzmewuowoO2YK8JgeKTF47ApsZZY1r7rJ1
xeZjXQXUx4SYNBrp0i9calOL1+ehxtEQ/KAUIhMuuPO/N7LeZwyk0rvh+H4y4MXVSysYAukiNuM+
eRbZBDPn9wJzoJEMk42qTe3UXFiKZytAhF3YQZRqdsgk1eI8hli/M99zleUCGssIgMyGWcI44npl
R3AAD2hjw4kobtg/aAK80jVq7PVpZWS7/fvrytbc+/vI5sNawomTqi8AeLwrpAhncWOHiekAOS61
Gl3t9pp5/1A/3cSGxDHOjTiotMV1ZOsdDOQB3lx1eN5TRBDLViudmMYtQZq+Hpr0XpM9DLWGN7Z8
A7sqypTQ0D+sMglumpXbAxGZVYxHWAcuuTI8LUtPpLXsufICWD6Jel4SA2y/3k+agrVE1kxmSSRZ
VEBMa3c4pdKw5QMFOBaSihEU3OXH8NN/bL3vS9IYU6le1Y3nJHGSZCs54mHx5+MP5+RYRcJiXKrk
TmViYwCdlA19Dk78pctxNdjXLtWzVDdKEBWMhxtRElcXehHeGvAE8neCxWDELi5iia0+QPwL6bJ8
2HAVCAVlQO/MeZ7FNdfcRwWCXbTgcwIzgJTMVAlv0WmRGFRTVPklx5Ipa09yyIhglhkPtW7C4tZj
J1E2J1fsq39rLAhM6sYyaMFSXWZcRapUFxQsK7oadTh7CpGmGbDgxOYnLUoL3MbXiviWnI9h2WmV
MsCRCPsiz/bPEKAMvaQ/nopPYFEXsb/pXYOLP1NzILVBxg0pUTnZameBJXI9brBFwUfp355m/Te9
gOOVn/LlfKQeC3j/ZWzF3xrSe5e14VS63mE3lXjaT5rZN2UbseDdhpZto21PgVIrL9VXegimJ1v2
BSh91iaLydzwrgoR+eBLtR7k/ONW+LnnJyHU7gtKCNdb21v8Y8KCUWrbt2J55+0ayNLCdjKapGdO
WyF5AIUnCJZL0m7lAfX033upXNovch1SnLd1HZVtl/u+S9xp748FVc3PU4OXSqUgrdBlXSq9rvT0
AZcw5SSg5u2WLbxVD/f0P7IdkmrAE84PxqfpKSA8Sk8GXg8ga3ARYZL9/dsSjTFCKAdTQD4KnyeG
gC9/0Bx28TNpUnW4Y36mMqsec/WXeMniplR1xuRmo6PCsMZVJWLn948jgYopjZqSbirhmzUIf1yd
s/a/bO9itZx86eJoy3ArmmanFBJ3N281ucdU6GOtAQ/85ly9FI6B+FxBS2Fk9P636+DiuI2PvZ1c
UAiJPuRwAoiZ7mVoSWuQB90HYxh381Y2PxdvElpfLLvk0iG/praDr3vmEHrCUgErAsOmeMQ0dLyg
yMQWgQZ/t6vvdFxg5fxlH02wWR1nAh0RI0FzG3t3lBfrdzkFv/34bLWzcNw6QiwIdFPCUm5R1qgV
/iSVj+HSAXzEcyQJihPJuThEeBDX7T2CteqG1YvFmHMWRcjmk3mDBYBK/5euoE2qqd+nPVI5YZYh
20H3azPrDC+MNFz/YTgInlNXrI8dB+aqjyeG9YhnaqD2+GjVG3Du8SyLTJzGzUe+ycDwwZiifjBX
E6LXS993PVYQW/suZ8ns7J3yKcOBJUA6rZqDHTUdj9DsbtH53zq3kftQvXnt8J3dtvTMRGPAJZQt
G5etA3BVNz7P63/r+Ulp5c1f0gj60tjEfcLHx9NpyVrPhFB12L9d+PlhUkNU08U/ikIOACipwC3g
cgbkXPqxce1IIkMKkErgdWEt4R90QXf250rW9i9ResM+dH9HtG2cNEIH3rU8L3BPAWSOlpuIcYMc
NB9G1qwwbMyjTCeZej7ErdK108p7d2ZOW+gSnZIerqwkOj1lHByKHUK3sQ4UcWrMS+EsgXoCXC5X
zYMk/wL2hz7Dt54OViUAcSPkOqrYXE9KhLW41QvPYlspR0J0HQ7kw3DEjkAxlzNsjEy794xrOtrQ
BGwhVBQXcSe//nUTdJEhFMfprrb2GHFIFFxYKURopUWn4o86zgHLwyMivxTm9tvCJPiEx1RFhaVS
PteNJAzHdhd17lfNsHoRu2LnflA6u8xCl5mwYe5kzpla8PTjkCxF39rDF0HNN24PSETjTWtbaohv
gmp+XusNCoOaiIOXTltRIdsMMFwoPFxrTzUyihXjXOzGNPb6tspGZZ0yXET7OQXTWkE5404bey1L
5jrwuBfvlMPpx5LN3osQofrcvRfQpuFYx/8fLTydP+WS4OKZZGsXXVTyEa/3jki8VMhx0Cm1O5Lu
D+r7o8OrvHHvsgTKRcns7crxPPgiT/mbKZHxDOgcb/3Zo2sndtDDiLZ16c2zhgx0PGLmPRyWSUfo
ow/+vZlUG700GgP9OmhUs2inm/YY20+ufY2mBZPp6RZL251Oy5pXRCM+W/Vg+OCoazDsZy+lsJ4O
w8Y/nCZVb/ggjQdrxQR8wjGDxWlQEdUNZn0N4qo2A3D0z/kZNCcwsBOAW+ypZeJsvWY9VT3Kyijw
o6dgL6ShPvJe+nSn3r/IshVBTZu28CmsIYChA4Y1Axzf6Dsb4frwxZibb2wiistDyoug9YH/suyN
JCJlmU2LBB+eZZSEwIJ7fdBWdKwCGJA26vSL9/MPPTz2nDjcd6B2giScpg9OrTVXUrugkeJjvn6U
uccJBUTmuJB8eJfBx1b1qRInz774A0uV4cCXg1CVofyiu8dV5CdN2fOmbmzmd9a13QuxqjSA1krh
jl5+zhC5FBOQbkpBBn3MYsvC8sAxF6AiD2wJ6g/XEmPIgNXGOuxzfiJKI6ViLhaR40Wmm0UsNNSY
Zm5HFCeFh3KRYvv/V0+psvhbHRc05pDoBGDruIeF8FtD8WhuByWq84WbuFDMaWOPj0JTcQ4y9TEd
Thc5eHDpho79zkB8RxwxwkndbmOyKPCemXlVMdqZmnAetVkHkYQSNAl2SUkFxiMpD+a4jzwjw4/y
d8ZeFzJAihllIx5rMp4O0cadoZzt0S0ezcodFKwkP+HHWlzB0x5s3juEU4Cuh3rcD9Y0elFT9lZc
G+OE2An6qA9fDluOhwfPZoaHGqqhiXUJo1bQBNg8Cng1qlWCkr3+ucqT6MmV6PVzBrXkULWflrRc
Ex//3VEWqP+5MYJC3/aqKKAQaA/ktyjcOHg+iTAOhOhOwYUx5b7/Dq7VNaDueJ/cFa8G3N5yBHxD
zvTdCUyv/yRS1lvzP/3PksnO5PH36WKKh7NHf+0wbpgJLXOCzP1PE3voEy9vRXxgBdo8hjTPj50B
tfow4sGnHeanE6R8d0DWIzWsKQsn9/IP9dWMPNtBB/aWsXDTassxKYvF160QDT9heJjqTV3mie/l
a66rJqAacq0bMF5zJvFmv5e2bUIzkNL+sqUHXleIUgqNJ5tULdZWK1EW2omLp2E0EvutTh54NDjR
WZ/815PtCa5i/Dhht7p7q6Z4fYPOHhVLWonk92ML1ADMoCyVH8F2Zj7A7ZV7uDAAwt9jyS2XeU8i
tfawhPXKCxtoiHfgFBfLkwFfmqE6X/WJX7S6gVOTGfEW4NGFHewF71Vm+WnL5FyT+TayCPD56KOQ
9v7cd9S9zNSwTdKK8mwugyuLtepxKZ+7RTrRteD8VV5cK8OzgomPWsxUydWhEEp7mdGJZV71jjvV
umyGwFY/3qMJznSJJzFkolcZBC2DXMPQQYPPKD9oNo87/o/3QJeA/Ixom2g6WZ57HwpPy3b8oa7x
F/UcY1ApVaGEFomHeXsSTYbaL+PDOmPpTxow1tW6gPvhapeJaSIRucJZwo/PzXbzw6kCcWyl2PUe
Vr8ofk66WPITy52piuR0fbusqnO1+I3PYnShG3g2BmBHL/Yom6X/V1cd/5ATmNlCCY9/2MiOmNBf
wWEVlF9bJdndjnJ7UTY1nSPqwyaK9QAaJJEmtl0R1Kx6QnsIeBwjrNs/MfpAcKL/5tU/fMF0HuWh
C1eQ5U2Wms6/EECl6nVvwjtnCRRUIkir8FLyvE2B0ciYh+6jL1NVBBJBUIYw4E9usGMgqRX8Y8j9
ogjgCMY1y4BOBycyfKdaeOfixpW2YjjdvtGutYxZbY1FHRegAmzNSCpWn0dPY1FpLz4WaDfY6OHU
Zj3+iBfcERSMO6UH88pn0kgYIfJ6VEbtlQrYMGYy6GpCnfCTI0DSBDota5+koAGena/kfb7MfV9G
1JQ+RayhdHyCbwNX8nLGjNvT3LbVTTa1JDQ2dVu+IMC37gEmJV/jONpaxHmSA65w0+m6GvyfLpgL
p4brT2RU2qxF02NbOAI88EkU1V2EboUqOrFdqnWPG7t2CNu7uKe3sZSkh5XdQ8DO8wKzwVAXSLhS
dWki4l9Zsf44U2PeoWYdjOm3gaVDUG7k1+B+867bBrE5z9EpwT4cegdWY4HyLuuy4nA3bXp7vMFj
qQYJY1VoPcm3m5BUBW9bQzoCgVKFXe8muO5JwPrejib9qLC5vRierE4uc0NWuQvs0fZDNRyWszKY
RFOg9cDJhJb5UqqS+scz2vHOCSagrK1zPK3VKd4bp834ZRn3MHpOXwfqYN0ql77KSqy5Ae421EmO
88d8TI+IfUBOvK3AgH7/YlxzWzzhHahKLDl/MlNlKSKiguxomC8QHGESFj+SltQnJ5l4zMeBg29/
M7jR01dAGcu2FY0wl7UTw9QGiiKPoq8lbO4YSncOWwxogYgsNadjsm3oMOpn6RLPvjUDsNKzVeZP
UacKs98LCraTZQ7xiku7fn11iKo8WtHHNNTfvsQ/9+l+C6rN1JZUrGVBC1ktrsgiQqufQRra4gLY
M2JiFxjqzI364Jku8eUDiSHixHQYAtCI2yBXicFkbhmEUvjaIevF7bAFreM/iXZ0HzATQhqQ3tE/
cdmtyZjEw08AmIKm+Exi87Mco4A+aNAczCgcoM5BmepyGpqruw6Jq0yU7dFtnnZ0cdN5eEcHxZV1
TWSjwl+bs/ODEQY2qnIFX/Vup7sIemOb0DbDzpNWs8qGJNPSOFjByST6u+4EC6NXy1sY0VlQSps5
c0cwYr3GCQYxkiCqMRKDP86OLEvlcXaT/nOzwnadAb1e1L5/4tgzF2GGcZGYkjoOX6ZAo4KgDUSX
ofgLrSnsP4x44Hq5zpL/foraCLX2BCR9gkL8DAmNdKJeS5ZQvBTYT65Wuf+y/cGnEzZglWIfmm0d
w4XqIHgGSs9uyXUiglSpauMo77oA46Fx3KIaHvKtHtkUKjEFj3Sh+ZqRJ3SpizFslQbdbRqfRMvR
SiQikFbBwACCdu8iOVJVEuesYh33TkcQ7d0xUlys6rC8Mf6BIvNMh0KIrWiciw3+h9qkGuofME0a
vFeIt2LZx+uTbvCroj/pqzk5Afd5d3RfqiEVWTQbZUUtl3jJhlOQZALWwXay2NXO6H8Bjmtbf5yf
xapFJL+Q6BiKZpHkSFH4oHi0BcLz7GaTGZJuRLJpzlOimaTDSqj9TvbrcIb3PLP6a/AS7trGIiyD
4O/c1Q56mW+2/rAlQE6msbo7weEkK7EbdqNw2Mvr9k4eI1ROPIwd/wTH2ElfLW0G3asv7+gY/0pr
aDRr8Gec4UxBuAon+3dcxRTTW8P3Qg1C2SQ7cqy+bUghiULqvNdlPFXUakiCem+2NbAjd2iQBxHa
QfDNQB5fkvkYVYuZXz40V5NxIygiHcZUYNjFTvqv+TFq2Z86O6DgEOtykZ8ghhr6QVSMOsr37+Is
Y1xxeJ0LTKVQMCTWh7YmddlXusJn3fwHhV/cSiYoAPBR8+kRN8PzRapSETUAk6+ics7Ysggd6jKn
HWPB4aDQyTw9EVwjeC1LkLFm7KA16n935LV6m3nN3MDO04otKtu4Rn0pLF5BleINP/liYjAFep7p
QH8xzKol8TFJSha+PNEspC7GApUpk1IQQ9VWD6rQgzsTMHSd7pcl7qAV88z8qlnGSg9kEvdI2iNM
mjfrrQyLALKJlOFMIuMh8q2Mei6Agw1wHlo4PH8jI+TlA99IZtwPdfhyH3WaBUQ5WMQs7VGjACDg
csumQDwSSvf7AT6bsee+tLZUcNjrhjjMraRT5vP8IgNxp2WQFIDuCxmnqcm/g+zcJXVrWz76vbbR
c0SpRGONUr7YYLOjdv7fNq4Ng6XFx4ggttsEj21v0QPQGggOENbEmi9NWK7gI7zMrekCXDnPXK7P
Q78IgyaQGokRBNu8yjCx/SIGnJ6/e1NYHb4XbzTGjXMh2u5bBVO7l743IpXUsXUyhsNL6814gB59
Tf5xsrUJE5NkSQ+Il+fXJvW92lC0guW/sBiIvEzpvBeeDJvPgZAOueeXu7qGjUt2e7dah/sqbTrc
BIwjEpjFcAb+6AsYW8e1QOUNFwgGeAFKhB0xi3xFq4Il/yrh7aBJwI9JuPjEC/zyCo1zDvbvNiPx
vtfKQvu6M2qkDwAde7/07ezgXP33Bu8Qilc17Ls/tMAP1W73QD6uUL3vFREXYsGxd9Y5zaQGpeM/
khTSZl4SeFZiY+YiIDFy7HxfUPrtlROY7f1O2IirlQ5eqfDUFaUMHkbPCiOlt6mCzuKhxru2pdf7
A7wzQaOJqQyalBsez/HVtGKgB33zyzJwm6HWXidfmfgo7G1ggQnWBY6T0v89h3e9oFSFSTOUTbh0
UmSsWNb48CgatZTSPCat7K2RA+1cKB5Erphco/+V22cHY/FepSLU+3nswmc3AmGj/yGceLiTvLl3
SZolJ31AbGzBTxJZGMTqz4jRf6+00vYionqovfE+ehm1VWzKSdbFdf2nPP8/DG/Icf3ANZXf+uz8
cNtftfkuKjmGObvOm42XkD6PJnT6kgjNPU5z6ZhiN+Sm/o8SssDiCbErLpeeXctVhpZ2WueR8+YI
euYfffmVlrymzALB5pREMNgq40DamNLl+i6L4LgyJTECe0ZDNu/02yTX1XvtbWme+P9xlMpitqoO
+QHfhI48OKUL6aDOWfjA3HnAZP8FVfMHoq1D18NajG+kcYbiQN86J6HLJrp+6wGpjW1lHwn9tjoc
nZcR4KELLndVUA8BnFU6Z9kEDxCymws3NtSxT0oKEQD/sIcYtvvIlPayBSNvYM91335qaHDA48Eg
CGWHHe545MMNLNiX3UNmfPEF2pgGbMESDqkm7U0EB7U/EjTe0y/cubPq6c1ikLXZQSAokD0RnAq9
DsZ/fkAbDNll49OW82vt8oYxho/cMpE8Um3RnIcjQfRwyuCbNkiGpeMWf/RloagCIRA/eCqDCAI+
KDxWJ5lPKcPxhhsS3cd3nVfbdRMSeQFr0SCRMQ+7fKZTcdjObg4INLJHTZez29469CTvI/6r8VFS
2JJoDXP3uulNsPemlbT0Jfk7gnrsn29VVqmariC8l1NdbZBC0rGOcJy8Sy4xJI9dEOyFMJZV6WD0
tgGSvj2NenifdVj4Tl7C4mtCI1MNMnYA5AjRbDLZtTEOQz1RPKGQUvy1acoVTDJsdGgBviL0X/3m
RtUP/DdPdkmNzAia8WPxCmdSKNiraIumuFST1Mx0Op+Bzp8Lc36N28a0q7gdJe4pDCt8xx3iT9X3
feXWocGfTh9Ms+bfc20q4rHNwby/VNQ29kOEBRR266vuISrSmwCofj+F2sJVp4GRFLYt490a0P5L
gsu+lHzHyn5S5HYnWNRajeQePdqB/Uu6a1ujUj09VpRD8pzFB+/c79bKBxM/uRGJhk/MDjQUEW1k
ssj0OFVkN80C0ym2mEjOmGjMGzXyb0WNMb8tjgnLguAZFhW+iJfPZEsfkfSSH4aWPE/vIolb2pvl
dD2Hht7s1XY6WsMtd9cTvWjmGS77B12TNQolQtsTDtRlmvh5Br4+6di6HoYy1DQhkcMdTRJDLS/L
6ENwczkx8vWnAeseIZQmfNcyFxUmynB3PQCjIx3X5JVasAiJRi+S/KvNqBVMBp6nP5JjEAcFrXux
MTS5CZrMKeTWhkgOWkxN9RhR9zFCDzIopwCvKNCuEL197nZDYSTM0Bp6nB0B8uuWF5Afjz2bixs/
YqDIqKLVqy+QiFsijG4uHY/+XaUWrq8uuhNHzrF/5yO/Vh50CPbnSZWGT5Qvs8mtZzVo0xvRvWs3
Y9s+JyRuEZom/HRbVDW3b+o3Jgn7DLfIYInEmzrS1OWVNU4pngBF/oMpLMFGTVGWSMetRH2Gh97z
wD93b7PfyZwcNfiSyXSSIvSipHiTUOSwQ51Z7GwPC8XbyMQnn6m+9Gi/Xyg7cMUQ2s/QtayGCUAx
AMmWEICQutq/yeKqNLAgmZKzB2pXC/vURyBX4wHVJJ1WMF36bx6N8m5yYqLkIm2Nz9UQWzm4u0oV
Ld3CljJLLKStlNXBheMY8BRFNn6cKyJpRNEfnoEjsT8KyjKHi1SBto7mnxQ5UtSBick3pwRQT+En
BR2H5D7JQ1QO8VEBvLHvdytTZUDUB9yEuDsPBTO8R3T6dag4kRpzdJTSDtm+dOZ7X6tatvHKzDN7
2ua5pnYtWnXh7h+hQbIjo8jexIl1CY6WUsu1C7a4a7x5tSCU/2wub3IFgUVXYTaArir5Qq4ZQkWD
rqVJThgjKHyqQCaVWV5jd/72jRFCa43tOgrT62v3fyYPtC5S4BCCCG5WQyWxGl714oSs9I7mMEcC
MxHO71JzrrB/UPVENnUGrCtr6/unrqUaT757nn+4l+DbIwnr64khOP1RZrQSGP8K87BIprTqR81a
31memoOHG0rl/ZJPS0qJim4+krcZk9FBGF75UVNJ82kmxJs1DRXMU8bZYw0/JGqoodvkJeyElfzL
fRldEkydW7L3M+ZggFb0nsgB8+0FLygfbLtAUIs8IJH9OjmuSf9wUnJoHgwJ8PQk2ka2LFAz4G2S
Tv8wudjO9ylQeWKaXV6KEkegPKeJNSOcKWV4jb31HAsinXg6hhAlLYCX5AZy7LcGpQgt8Ls2pfpZ
muHLw1M1O+kanN4s9UyOxW0RGeLEAT3yiiwqKp/mLxCi9YMvp5FwNh9nmEM6/EvBoEUVtJAgT0k5
8Ys0b9gV3mE/4spmHQ1hpJxsUoKRQlO14cqDS69jsePsCYSmLYlD/gxXprfiGaFUpBkWCNYWYDBW
wcJFLJWxfVEi3QTB+LJNDzlXJU2wfLXRAe1zp3PRorh2z28+zEDcax4KEvZr2i5Y9g8sxVJwAGBl
p8+ukcuv60YFxw5n/5yznefli0dnxcbLl5j7fU0PwSKq4N2rUDw884sVTc4SvxsTXAGun7NgtfdW
GgF2AJ0M9uCnKJqrK5OE3BDmtAF19VvlDyQN6I8fK2iPD8x6khA3NWPygFWF9OF7Z8rFrvQYybgv
ZEHWdmBSTxdGkAgpu/Osj3MgfiuNGp0Ag44rWcK64XDnA11SWkjrSw7dAavfbcoRQHYIrIeBKnPi
ZO6JVoZcxttMvLags54Who4F5oWwWpG5lFIBRvbBS3BQNDRU+Q1pkpZEPsjRxWVNs6L8bXl1Y2Bx
qqfySvGIf9XXxlARhN6IutujRsPutaaTXOtiX629Nnd1VOkEb4HPL4EJd6ANsdL5/VbE5n7EQIjM
lpNmElLV6XcqbnCmQEhduZKRiIqVMx6BbQ8OUBA75fPWb2HGaNeAfDVwPXli0Pu0WkrINyUxofdH
2O8JpvcyyHdAEApDxXzeBmorrQKCspleg4c4in70rcGv85wGl4YnDFa1l9wyAmGvBZatI3iDQLfG
TLScVaXcTDwd5m81RH3/zOL9vWO6MlcEIGWjo3eaQAN+H9UO1u1qZvGLta2pKVu4Q8dKafltZBL2
pNCZswuPsIovPNQqgShXgzPwL+30XPaRSui893kK9oy/38QUJL+6ImjIhQ5oTWYW/ss77tsAhjzG
kHtTNjs8lQVHB6ujIAiMAHliXz8gUR8GgvQHff3wu1yIwVKVLdB87gxXfN+Ls71sXC2wG/BEItjG
Tyju2uP43ir2aa9lPaWcH7Wr4M2638xForrYtY3WfAYOVTkxClTftv5zoy1jPTWmv3lGjJoaYdFS
nDcbFLF3Cr7ECeE7Ht5R0KaPQTmA9WZ+quYHxZVl/L98D1ypX/4z9K7HFos4RtHKHW5iQPu1OaPX
ZLACwOs8g55xhroewbnrVvdb1AGa8dy4xmSr6rEZPujJ0KS8CBQMoWAaHVKFBeL4n7AihXl0XX0Q
TqdiowTckELQX8HkaGMykHJdpzMhyigFEagMYTxopeeWL8/eTJAoCM6Xs+V9p713DheN0z6ux0hl
ZgIqL5lEbQG2+W3pAmzQ+3O+SjB0cU2SrZvvK/TNENLVA3ZgQiCvfGfS9GURod6HvZCd9VWj0oSQ
AvolFAXkaiEtslAtFU4kpRoULqk/G7AaT7ftSRIM5vtPs31sSm8n/iqKP1Bfn1ZJ/WGejgnakINE
Eheg1/ld5dzJzw0hX2yD5RbDCLWYDpSFX+q0AczOsd91lmBu+PIkcZteX/JfSslQBE7jLZ5dLJbg
BrLliQIWXAziFo+FSWBPp/UhFO6IJaiPAwYtUH6XkJjiG9b1EYl/t0vdpIasSI+5xjXpUop0Dps+
CmfJCq3n5E1l8YtmLkniUt4Tt6ENtwQVfYtl2/9+2TISfuMAxSo6TqoJdxIVUv33BWv+3mR64ut2
PYUdBFrkAeHAA9XTgzuIxVMJCmUBWkxcm7xmtyzf50nbWe+aC/4LvMO4UUxAxeMDmCBhgZAA79vI
v5deA4o4sZSaow4l8oaqocoGPlHM/kCytzrf6SZmF/Knrql+u+Vfv4JehOqoDG4TA+kPdpi0teoz
hqKO28WibNlWdI50E9tbqJVyIp19ORIyuKUnoDJVC/nl+hOcLKFW8cfNX7TV0jW5i5Sqv6p/rxhH
4eEnX0iEAe0yjgxmY8o91bRz4k6TdtNH8N8kjGRo3+M6/sfhQjIaR0x0H8Ddc7uGZlRJHhSnWt05
DlBMUuNym5LLDBVIXrG/F62NytmqmrxBaX0M0JGxtiaETpaC+NESto8Kqw+GLOPC/doyXXHhsO4c
AO2PBAlWZfdIevJ2CqF12t7FHI3C+zBJyINFSN/Y0NQlYJo7NBDDMbD39YoBRkicACEkbrlJWjhI
sGzL8TEe2nXJ8n0WcutJXJYEuOHhHl5XBNCKssTe36336t1lWhhHO4A7SDLhqbMTeA3WMZtXA+0h
x+QpoFDDVGKQkZNHRcRHSKxEADdQjXL0hFdnP1v/lUzRUwVxGi5WfwkaIQ2ygk7Syz+NSvzVmcj6
Ze5YyimtsViTmTK8ZUr+h5dZcQzhW8NOCY1tNLilInKB5bMUtfhq9XV5enJapJql4Z2cHgSdmCG/
PxCyClkhimcJo/UfubfOD/xAqYDUqzFcVbeYNYn6dEP/4JQsPpG23eKdxcxJ1nT8IHTHQLm7Yum/
wLRJFk6uxtmjva0lO5eQ5F6tujnShtikPnjqaQmIp2bvdjBeTjyZqJ2Gno/y4I4IEgO+yXRHRQ7l
IgI+nnLOveEKYUuk305XyKB/Ji33WoyljJvJe7TrsnfKgBqnJHJkU8kt7ZZ+v0yGRL4t8JMCnYIh
/JSGdnDhwaaI30OYQC5n628lxRyKTvAWP2ebdDSm6fpsO8tBf3lX/dcU/PFiEDfSSOUH15hkZz09
nREp7gkri1wsngtTpgQJzqAJUZOcALiuNk8ivUTQ2SyphntAsYNef7qHQ76Zdo3lo87f8iVhh4hR
jZ4svh7xSE/fE720aYMTk+67jdQWQV8yR7R2d+cYfTO7PNf6AGwNlg/z6tbhwCpaZ3t9EsXXUtFf
X610SwvIPFv/q5qFpkA4eAOEwcfTObp5OtTqSmLDDdl5sFfTPmbDsLwg7QtMRcus8OrJiIbAT2yo
Mw1CQNEHkS+Jg/Z9uLFfEQhwQ5BfyahLaVGZ85BvRmImierDW65mJHP/jRpAIEdNb4ngkcIf28bG
+JwvLWHzXCXpAXvtGOikolt973sqZPwcS3aZXe66IgVnaAsnarnDP8+xrxMTR9TW97BbrNT8/W7J
xKRuyO8LXG/1r9BzHaJHI2kSjXvyi9z9rp4Lhg7gYci2Na9fhYZs1ugvgpZBswRQmG7Q5YTDrxXZ
AFXFC4W8n/Z6QVqnmeD14I8s1NtMqlMcI1Tnpi59CXmv0hEpju2ZwHKVRyBzwAb0YXPGnCu1aGzD
bpLQsn01MWJgW2HqC75LuYoX+9qniisw03zt1LL3BD0wkvkPcMOqXVOzG+HjJYx3H6GBkjUfO4LS
/d3KoEd6iHdv/c0WoVwGcYqUyCR6gPGTRv8su3aat55eNAGTzb985ElCtXzsIMIOFSLsEguSasPE
4LgDembtv94u0cbzt9i1I631zYNvv+RJEF4Du7elmSZWM+0MpU2xv1ECMUJ8McPFa6VMBTiEs2Cc
5JlS7d65uVOHp4slvpWTzc3mJuIg4cc7ISaDMHNnpWhB+lBPe+g8XAmfH1ekTeSOrzEi5cJGAunu
5FB8L2VogIfg0Sj3AzcK4KARs7yQv/OV+qMPNLFjRXQ32rQvcG5W1A5oPP9mTBTaVPLKeq0bgdgy
9+/UmRiaTkFH8D1ByLnlb/p6A3csB4uFzLhIKOamujUoi/2YiFlBhC9V77YvioLGmVMtxasyMaM1
vs932WVg9Lh3rv542yWDpbHd8Gfm9v3NimZ9ZWgH0hIneI7CWiNKUUMae9EtRWn1VdF476UsfyS+
SRHNO32MJhENQP/sJ8/wuyw39mZaCWlRujA5+77nCHUUkINwl2BhZpEmKCj+rEJgaHNL5n3a2U13
ZPOgCXCC0B+FaALY/7skPXeaT5wvJHlAmtOtGQ9VMrKx/y8Q00OCnHTaa6ODCx89466/5V8x0tEj
g+bDUwjnF+jx0SCY1VjKb882Pxmv606WpCPZdyeK4IuzWgP/hJsRBVrC+1nFuQ59bXzg13XKDhsA
FcB9YC830xs1Qrv2PdswWLC7RQXiEC4ioCO/9ilOb4dd4N/9zfkj0AaqV29DCzEcAmNblV6BoHFk
Csh5igh+i+EvJpqZzdETVBhaP/3TIXq4U/i6bRBh3X4wf+gOh93x1dTE4Vgk4r9Tl+nBREMi9nQn
PVOqO+/mihvK/y36yaEUaj8nPK9BWMgbzkA/5pLj6yzHMqEJXzjW0eXVx/L7XwOzPcZNl3qvmOMy
pIK56CMeR1oaY+HTWvjrRke+hHBslbi/kdcMMo9qzgFf8cDapz6QiSUPiblWgUCENPkTE0XRqUJV
1tkcVewvlf1ABasz3FA+2iYWFcPtEHo/Xb9Zk8SknhkzT87S9qAEnKz7LrdrazQu3fq7kWHtTNxl
cTO/QA6UeGUQmmVx0IEobv/yLraJ9+d7KhWkutqXWEtT/dk5UbduAU5IRVpMiMkzAjS9qG7cGmAA
A7eNEExJ5u3d/qh083IdLkCxxyzFSy2uKfDaTQIloKoWvnpjfZSjhP2Z/3WZ9g9BpWSNBYrZrcBc
rfa9b0kiPYxFMABAYocyl6QFxif29aXY0uPVHJJswE3C8xLlndkkOyHEfR8z10A36WPzncP75TdV
5WUqBUIVwDitoDoB/eztC3uP8hpcLykS0rzf/83uJ5zFCQt/YngAT5lw1wIon7FA4sKmMAdHs8uD
QT/91eqyRtsTlDFx3BZUIvHo+QXs8fGLaqFGSSK6DnVOZbD0c4vqEA2TpztjvfwU+3S8/OOxpgs3
UChPeaktebFDgBRonxGX/MGbnr6zCFt7dD0JyMkEyXr8+Cd/bTB2on65bKVoIXM+5Xpf9g6W6QmX
RhRp89ux2O/T6Yk5aFwIqGnIsXtmnPkFvPfL+ZwIMlkdhZcc2BjtosWauHhW2syiv9wEeHgU2Gzv
fziqntt9xgmWF7wbrv5IGa5XmMKWiDmOYP9m6pSS2YxihqQramPJwpQfXZlcgi+oO3xqS2d5HWUi
3Q+7k0nTgOpRuxcDLUgu6c8DSLK0ZhF8YGn3djwjHEeYEU5q7a5liSEXUybNSEKD3ZB5ygVwLYc/
i0XckYzR3luGwDlkzl1TwmtrpfjJEyb+fE/SjqURedhIuEIB8lqSjdNM4HzoZ/+exx3fexQavata
Rxh95Os/8uvwBvBrYJqZPhgXIhdR8gBvjsBzdlHexvUtz2ndJyHblt+CFRgQyEYQYKhNaNWA/6Fp
27r/HKcFqB0eCif0wRQGslzIZhXVRpqq/orannwy2RcvAbFuld6qPVtRqbqf6Flz7sW48H34ihqm
IoWvMwHj01ReROIxEB+l30bB7aBk3wI3HCwn+6bmKI603ChXWz4JZgNCTJlthCgZgKVXKeTWZQWM
B9OsRzi6VqqlBDtTGsiJUWFjIl5T0BRx+mnX+gG1IK7jQrEkFvJeBnNVZmeFsfIuP1u10V/MVowK
ng9GVBMJdjUdBM68rtA0pVwbDkTViVtGqB5SRLJ5Rgrk8/f/aYis8M2ynqhwwb3+Yw1qdCDD5dkU
pna+rfHES6ybeeRITChSvDogdnRNIVthSBScIEtDXMLGEPOgoeCnPiRf6VL0wEmHTLov/PjOYqEh
4Xvv/rPvx9sLcRcbsc22ib8aN1SUus1xSvE2ss8tY+xA+CGXY+Gps8JtGvmgTDBbDhNi5isVMNqF
boULBRCEKwAK8G9Gi07OUj2xYTECghhUQGUjbf7qxuvzCeWmo7P2FNAbDYhMEYt5ltHkohtKcrGn
RRohLRjaXWT+CxbRXmYtUcuYbUANQl1ENKdbHU4k1go0DcxL7UAXhn7bxfqQoHI5pk5VKgAvb8XA
wICOB1A3O+fV/C43GaLzdUm2psf+0NT2pTAG+XW/nusuXW5VSlFgWONEwt6x4I3Nh8+sEIJGPFZI
KUZZL51sOkSPXEIvUsni/BL3FBdunXEyzW5o38jz70C96DnjSphwkXYhQCzZNKpgUhn4HJ+rWUW9
mahxG6E728ML+dD50eF7f7LpudIZzufvAcxKTfjMq8ZKtv+ejnXlVoI3RgSPcJ3MIcj17D7HFDaq
k+9Vg8iDpxNvyLX6Nxytq7DbV7S72JgkjKDTfgIFaf+zN51S5ALwIf9RkP6u5dJKP8Fu774zViY7
YM7Vo7Vhspk4e1Ti/NzPAhJf174gYKIFbtS9iBL3PRlLa0NSNW1UjaTfCQxBBB9edYpwAB4vjlQg
szQPrep2SJGeGEmd6/HDtvbyboEm522cecfXIYkYn0pNAOnXUpQuOhuHPNar07kk6SI7RUS4kUPb
9xaG5LS3n3iQj5qG0oLSm2fRDSFCMhaU3RuZoBA9jOH+ATS3Areh8Pr+gp/yRqcRvRd++Q3s0fYp
c4PzaAMbIp2XBZ6CMghs8zNwHocMKrI7WVSKePYNSN0py8lxJXGnGqGNiYe9kldd9NsU9P78l8dG
ZbUGu5tk4MeqrgakL9CvN70VJfRjl85dg5B7HrRJfuaKuThfeD3lgFdWs2omfUf6DSLbcOCxrkcc
jsffO8YKaf0Lzm/BQsYvIUfZH1/xgUpUs4puifuLm8sbIa2e1cmY9o3B9lAOGaC3hWYoNbNaEaGt
uiWrse7U53RRfTQkTi1fZP+YRY8Dq7WDCqy2TgZR+aetDgrALK2Qy2tFhFDjx/yntJ7DHWJ2i46z
R6GF/bE4uCb11A/o3chY4lZeRJ84BiBMoM8tYMqQPTsMtPTlFPwy9H96M+b182odzcs7xH9lnI7C
GU8GtFyySWnGJLwvPN5lpaMrt6nObI9EXomHj3EbEWqrhsLPaHzXTqNv1cxqJcI6MoY2X8G7+aFw
M4npPJRylJv56GEwpGwUmeYnX6POFbtyl6bAqNlsnnfz4eVf+E47cfTF4eBxmEM4cF92eI/D5Fv0
BRbndM8yh2U58ah7zJgphsVV406py/2VtP4DSCpme3uGx0YeQsq4rJtr1UgEUUNvYLWBNnY5Cq1a
77Bf5C3PekuT9H/EngEZyTogIknXcFVkHPkefcJKEQ5zvUQ9s5GYkyDeFCo7FgMg3uldbzgLGGnB
n/7q61t7vOJ3ythA0tC+g9QVErxM1d/8nqbd2W6N0lVSVKjFyeNgxZpJwgxaT1pTduT+MTA+LpLr
Tw04v/UAr83A5LkJUHLoD8jso0Dc1qcs2BlrKxeEDnrjSLSqcVR9RlfHxjLSPam0KktS0CAk9zBx
MOUBMUewBv+dywCUoDkdyqP8yN+hD2flZ5ss1VuPLxFI5D5GvzGxzYjTVPo2leLu0f5fwrpZZZhy
+mPQ7b+vGV/Rs5jmuRy9G0f0sngBGIghWZOGkbN00hSaLTVRRM1vOnU6LjCQtWcXw957mhjOSTsC
aT9Vjodrbkcywfrw+AwlAbTLygkqR9VJoBZHkN83imT5Ra1ZGVv6hgTzNYdWPd+y94TTIOCUnhjY
2W1xzkhsZe4b4ngR70EU00H4Hpy2D922AlWu4sPNYV6s9pWcJgJAa39QUtcJ2BA+CzCIMrbuCfwO
+7Qs723/1jBepowZAQY7CsRu8neU8QSKvSfJjVkon5q3QjH9XjdQJQh6CFjRSjk1K2NZOWKBzEM4
auFS7UGssuP9pnetBEtdNCqieilDVYljSJ/q01ii3/ukNae+NXHlCWY9fDjOqtdEUsLPFA7t+g2/
w8R05QVKJ7LpD1OQko+ZCPF0qkYdhdzGYmAZayr9c74m4FWRSwOQDI72ervYDBC81o7UqOzXvMvK
gaEYUDa3BwyxFnuW1psXHhuoOYtgqe8JBwWg7a2GcB8jUOkzS6GYkNEKt/NT/yotd3mrk4qqHq09
BXXBsbxQ8HmRhCkXJjl9LtsCrIwDx6gal86eTNa2Dr5ki1BxaASJZohRTSwnOCXHZXrMZZ+aXM5P
K6LWfv3dfhHy+7iE9fNH/YEr9u2gp3qsXFTPUx5ezY1lM4tIAZYoMcZZtmdt0MVm1xTLZAK1BBrF
OZo3TaBhDzWOQDbZDqX47SAxaPPCY9DXlZBFbUtO4tZ58Hb9hKVGvZPP6l82fdhftK8r4aOYUkiT
LnpK7o4tSzgjVK3dnp7aF3dWNBZNJnMQhCNqK/uOyoQ/sTaWw/A+Ec7OpL5s8kG/piqa/K7Ovpm1
71yi5VjfAC9thAbfxhxDXN9Vy+Ud7BhUZI4ECnQAmNpJddsd42xoPVnHNVk+sqoovHq184/s3yRr
ATU6OV7C/H6edwKQn6UIejqxI5voZ4tr7+XHpzgvTbqCNO5d7R0GFEp4OWLB6AjsCo/6sULlyCos
WZ2Ny0cIRzHwAXgWFrhkrOaZgpsMNmwLwFlig/5PaTKajL8rMWPoYupVel9vjwhP+lS/InhDQrQ9
4U0/zgeBaI7SNP5Q2bRQkLoK5jnkWQzO4Y4ioiJiHj3/ZKn6c6OIiuXUxcducb07LA3FII2NI2u/
Ofn+U/9UY57y3QnyrH9hM3ugyo2F5s9ZwWLg2xeY4zGZ8iRI09Bm8L+jYF2wvhvTx/j2NYZM6zFr
GvzfOepD+BOapP+umsWt+fF7wIKcjZ1wc77kB8EquOQT2K6WMOgg9HH9zZCnmej96B1HnVmeW3hQ
7Yz89JCI0V1oMvTePl6fnl3rIAMRenRLvbgEkteRUkUO5KvDUEqqu4QHwHCwO8tJct7dgY7xM8Zj
fqkIKSfWEeskiTbpAin42XTYqw1VBfp7K5uVI109Aj2SbbfEUJIPTBOS1Uyb54L0TISLsipdG60k
6pE5OHdTDGhPqavWS7e65VunSGhf7j1gcs2yCdKawEF3Kf7G4AuoGgfITuvU65XbN4M9ZYNNjsNS
ijM927DhYkUWJ52oAtGCSG0QiALPienr78H9LfCDSBeGL5+e58PgxVH77JKvUexX1n/7chD5815N
uHEOnEDDb/rsTilsWdm9cABTDCB9LmBan9z+bMFdabmvXKb1cePoo3J6gVl7YTJoO0GoIDVv7r8g
rjZl4GQXY+ljgePn3MdU5382x2O/S/wiuYce9PZ4gSjXEPI5HM4ObEqChBZ777p/GpPz5lIK5rCB
9HVG7mvBJu416AcskEFbyoDC7+MpqpND2pb/XD83l9wvu2IKZD8Qcd7uGZuL+DSjMYhgyqPrqI7Q
3Y3NgG4TBDCaiRUkCn4K8UEXjmojWHDCBA1y36Y5IzmK3ZCgSgC3skztuQ20CUrT8JqQZ3zQ8eLM
Q9DJO3mo7rqhdfv0wzZ1TausFCuIpZI9mypJKSptX4S1LEiBO8rxS+j0VgKKVIN+GWuLFWAs5Nf9
mOTKZrGgjplVhOXQ92VC95OiPph/ZNvRffjsCtUGctEdq7VamA362EvG/MNAbhvXryNRS5qH5rYX
azLz+dt//psykTL0n+CAOY908YGB39Jy0g5Wz49v4AxPYt4sMI81zZ2MurxY3kr4V4/pzoj3nx8G
3wnFKQqb9ITwmB9L/z5liIs33NlmugE8z+uyyQyxw5AFzQfBEb6rb9djYy3J29NSH3uRU8URFqtu
x7Y4ynaxao7S9lVCZhTEMqwhp3a57PgSTHPBqrpwYSnsAicc40yLaP/HTY34lmFREr277QkjP4Vc
O9wnov4FZJq2p6orKpXGrQWfzqOOY3x7kouqCICeegrB2ZZpIEbl1Odg4LAwGKl8+m+Gj91fz2jy
zh7sfupeq5N978QO5PVZPczqeqDVbZAec4Z9zjOcqzIYqzLeGODfLikYTDx8+OVM21q6IL+wDwQ1
RYsQB94KffTIkN+4Lm7D9lvdbNTquYj8DI/Nx3rbVhmC/E8xx68aWqQ+xzgJrI3jFbExCWc07eas
cj/yKyHce5KEe7lBbXjhX7tcqpB52iZ5+JYORgwgWbRQlpHeSYJi/jRC/Caye2wyMQX1dLFVnjIz
t3ImvTQCAAtN36Wqc+yZeeyo278CO7yfe7ChWfeEtwSxDYh0mu3OLUVy7BkEL4NhQ0pi1yRRp0nM
gHLWL0z1fbYpXC2SxnevB2CDzIGLmGchpCgOjmoZg0gUvJUdnn4Ia9WZJj9d5cG6hMdCyx9hJL6H
G3ytidPBSQFkR2HZQJ+YarPfIY965ms/ceoF+w6C/tlMY8Jql2TjsZ8JrUvyjAfOmvigFqS2Hc2E
xV3HYyQCqD2jhJGbQD4LbDzMUpWiFwScZIZ5X/P1ZDn4eKSRioHAF9iwuyXfnX8Qn5wl2MJaRScL
xLR2QHSuLEekBe052TXFG2+D+p+JziJF7bShqsJsBYhfPWhYczSxKJ6uy4CkElpr5D5LFfmhpo6g
YrUk/Lz1xWow8TRGHNLt/LnKg5eU5Xo41IjEnBIi9doVaXOdZtizLXdeSxHlBKNgjjXvKFtciA0U
XqqqtckonF4oBDyKyukSxadUFPNZbHV764U2ticnW1vep0JLYSRI8m9LtFfLW3BMHRgVU+7nQK9a
ltYzk4H5o8OmUDQDwjMGVGIwgP99rHW/go+LDG3n/AviAbbR9bbNpKIWBziCOQ+k8S65FbmYO2qN
UomT2bovky/2dzllJIZMVyrj8Z9DiBcsJF6B+CSD+B4n4eZJd92U5BQE1odddoOfGjXO3PK5UiG6
wdgcbFWz+FWRK6wPZeVUyLmQZXHp63CeFyc14JvZ/IJJLbI/O2nwZ/ywEy5TqE8D5tN2pO2zF7p1
3cWbkKn7GgFDj4CTXLNum5e6QG/4D7mDFVXkc+W3X+ZWYJOJkPhVr7dy7g7+oytMouJIcSDSXK6l
lmw9fF+F6F1ytM66NglNEwlF3QBGntpE7OzTc702Q+JW5HceMd9EMPJniIsHe/a2fG2rY+Gq8QU5
taTNtuv4Uvsy8QKc2mhwv8uC11BvRgpmZC+g76NrTnPoB0j1W/ZJGeJ7hue0KZVu7G2+liKq1pXb
h9/5TIUUeNBx6QnpILblGhrysY4TUVEvye7L33+hwu1LmB1EB2U5WIOA2dF3IscC/nu1Sp+BlZ9U
asZyPpQ/E4+Zq4cGydCrkHCWd46w7/IG72ccjTJzybBNYTkEqHrkVZKybIcrtm/WIy5jBnVCrOrQ
6Lw+xzsjMhvbrRdibAMkwmnFPovog/l87+y/Ii+4dYoZ7/gbiRkoeraJOAtey8UQeOsiRKG6mfxq
lYpeMZKZdCNB/8JR7uPAtLj69NPfRofzBJjmCkzE9p02apHVI36d7ecOwzcTUBLCbFUhu5MggBWG
u6FJAyJXlnU2App3XdUh36yOATa0N2NaKWzIE3kUjC5HRf/SNOE1s/n1a3CaGGLUKVTFsk/wQgzV
ul6kxP6CWs2KBup8xWlNmOm/RnEsxMB/rNgmX0wUXK4Ez3znhmvMtCo3AATu5yMPpUvCAzVrbGNm
bfBRcgq01Vi7VAZH1Yk9j0LK/Kts8SBiDRtGOhaeU6tSWas6SW/hYeY+bKQH+2SL0om3h/zhg0Up
FsY3hcM/y9G1an3IppZ7waNL/3/icDFiXziqfWti1+0J7G+0Fom6ocLfzHkMbDulAP7pAo3TmaDr
xhk2ISuOqUFKcxaiGZeuVDqZXAJhpSrTBSYcEFYl2TDUV6oRrVE2HswCjbyFnLyEG+N9hiSCClSI
oC5Y50szHT2iZrlx8EyagBh9JpK1FO+X43hJbsviJCImKxB6fQ3BIYuV8TyHZRZXf+2CerzHe8IH
LEw3v+pIgaD3NPjut7tuSxy6umBmhOtK4RJPlTt7FZqTh5uN6nKyWsu5BbysGFdBxjda6UmPUP9J
BzrVOKiMned6So8qZGNEQf9NXJWbLYBPwOAUmr+JzKvKBvMut69cULprpxN34VQO7lnAKv6MkT7O
LUkiQiVhim7m4U7wfCMF0h3H45Wq1NTPvUchRnSWGBGoybkXYjlCwvnqSVsIzcySlaEo91IIWesN
1YYrDwt+bNVrba2avSRYvyG8821unQjVrkBHwemf6e7S89WzRACw5DgDohVMdmguSpcQf8Qm8c5G
T2nceYhaGY0g1XVKlLF0v0dxqAM/mTkayWOr9zHBcyGzO0jvouWKNtL70oc1GvqBYophx9ZyZaAB
/OvsN8zbuJuQWjYQIzxjwtdr3toNS+38NS2ze6YN0u688Xo67sWM9DeB3xKFVdCEy5StN5VEpZ6p
87X71lrVlQU2A+S3kMj/4Rbl8oV31D/sCFQsd8jG+XvmC+1TYs/6yDCKxiGZU0Wj8VXZGBl+RMAh
iyqqcN6shiJpzu9w1nAa5TrvlE4fHxd7a9YZwhNXBDpMfnQCq4Jyzl4phTppUqcZGmM2TtrqSZM/
r6CnY3I17GYGZyNBouc+i2uE8WWmFG1Zc7elkrklEKZC18D7cxtZOrhgFLl45kP+QbRRULjx3sd2
KfjkEGMBpjRhc1C5gm3olPYM/IgA8ua82oidNM8JrsP2CpVy38fMECB1+Of8hjyC+dZHhw4CCkQ2
JQEqY/+UhtcQU++YoadZAjhgIrtrMzF+ucXDKGCMCulJnz1TpOZkRWVv4ct/QQXOKrGYAypxfhAS
LzFH7YAOIJEOvA5nBDc0KfyuRkQ0li+7svgftRjfFJN4LUkUPtLC5bfLA2AylIK+SiwoygOAaOVn
mDT9y05CX7JcmAFtgTXk9ChOky/51TfX2p3nce7GWtNM45vfaZ0+KBQwDnpiAK6tTDzDxs+w9wIp
EoyJdk6pFm6U6LmGVTEuHbtivJ2LH0g8UApWKIqKT8Gb4WnFXR2eYwU/90vRwBFlcluF1fQ0x0GC
wCONF7Hw3KolqIHfKh4ktb+DsqWgH+EICybWQSleXkjfnVKhVglGAGQqN5rPOFMGNQ1bXT/i17WT
ogpdLcCRkrPu68LYY8nWepU/efrSnQddPmEE3iudPFXHDKaidCSxTG5BS9uACPZ2Si1hHse11s6u
AwN82ZaUDm3PxMdQKuWcQZUm906ctTgV8ojp20Ac7J8s/ifcFrils138HZKcmmvvgfTBIhihJJtr
TJNrNYyj3IjTJIXCIVPc0z/ewRDq1zK09vrUAbQywRit402RoVzjWqe11d/GC1dHuXlj5E3/Euul
1OpwL1ZhdcCbPRsU5X9E/O6n6TknODLrbY+YPuDe7V0ovcSCG4AgAZIn9aQP16QgJUQmBM5WGcsW
einfGyPOPgnCDhJjaT5q/8hLLIP1R9SmY/fq6Ka3GOkbOoh+9zG4HlKtbs4tcqKgwOs0ZixkpD42
FAdlXIeeQOj9Pt1kALxCqVxZsLtU512n3BJwPn3I+dy1ef4/698WT9u7VCF7FJQij+o3DdyjGUpe
AHkKKPkTE9NnWB0f3LuGxawOR8q7PWnHipF5S/a3G2MVuXl5ETP1vUGfCxBiunqrxYbBaWV0Vzse
DaZIwVJqBmrIhMriG4Aclw0kgGsXCMyERXRAjagrecHDfAqmZZfhj5Ng9R7aFWeyWuWz1YIiudTV
nw0QBETiUCgnZa4/XT6jcH0S53OHGT3rZJT8ckOFjJ7kvhr+j0sRLmfgjAyVuVVGe1qW3HniKt10
agSRMi/05wteql5U1F1S3X0m0MYVnpFmmSwvDmZXwXlxI7fFf9qj0wlWkap9A9TyEGQEQ4QvNHU5
TFqinG+AN0Dkd3B6pZffXR8SJ2GolyNMvMQ2muLGqcL16cROjdcEDQTcE7dphqbrLQfcKOqko0PJ
w7gfNxCf+t8sA3JnJ+ShVj7mLROvYteY19GoG3sXS4qlQLnKNYd8jPMZ3Y4VwB0Z3F1hvTmVuSMx
Fs6JIBvTUKFqSk/MpvPSmfUqPYMcw9AglR1U2Lv4kuHbBt+Laxnx6QXGzeCZBBpFbr9FXOevkfhb
/Q8ubYElla8soVzsboX3p3Ywjq+krjq39zudlJ6JagypVRZLCupzSYAxkHqS2KcEugEsjBCN/B3A
+CXmDlk+Gc1Nr5dR1mI7ZP1ULlo27ozvo91p+rF0PgxbtxG97172k4mfX2gj6qyf14ax+Xvrfr+Y
sS8Wn+lvkzzQaf9wDl1pCz9xZmZCwzomyADJ4oHqGIbygAwX1bbnybcFGn3Zk6TmfSf247UtqA7I
Xsi3bFesk9O7POeL5XjKP7flYyOP9ddeHiAb2TTCW/P7gocyCO0s1RviI/xEsPK8rh1jKlUbl0dl
5evCtJXGfnFhFndvzrZ3kqTPKG7bvdkgSYu9bdB4167iyg1QQ3rmjsRNRVh/I0nbB0eqfoC9NWQP
i+5Ym5CjvEufO0VjMc/GGDsSMK/5cBuz3S7aEG9FZnCVUM9phdWVPVw/OK+l63YyomY4Mti1zoRz
HsYylp8Mn3D9x9pxYOlhFMKp1MVPhGR0xaVDO8kh/sk2C8OrBaQuEtdT29FzCCr7P9N4/jRyMm8V
TkLsAzg/lXSWJNVcJ758x3M5p7x5Ob9V4sfMqlDtKGICwn7lArQsPEbVQpEKnJ3Jfqw7mXz/SHj7
twhL1GGiF5RQDk/qNRbyLvcD2LvTAC7MnNBETtCqBqETJvEeKjZVpADxADkpdNGZpZNAo62icLc0
q2LLgUQWI7apZbvh6afwNm6D6i+ty8cgaAMto/i0JthB5rpP0sKX+6FBwZcGz2uOc5trxHuIooX/
tv/fE+KKFq/GONLQ6Xu4PSXxgRhueo6PLwRikLNbCxDFBOEYeG2vyexr5n5iNinJegSfqkKMg9T8
+JhdOd2pCfXIyE6h6/JQ28LKalOav/oU8myiNIMyb2hBxrfKECmkCFNXqahhN7YkUz0WaIHRS/e/
Jc6rwCD3vlUiKXu5dztgkHpLEnTwUuu1SV+nbFMWqTSnw4/2+9HqxpdT3PtJ9VwLeNA7FtkirvoN
SaHLjB5V1kEPP2HDW75nxcepQa2opO7H5lkmgzrSBmg8WjUYm7XIkECWMeYOtzYd/JPBpuSPocGl
v+QoR98KCTgjIGa6i7sB6E96ipF+8O/ceNN+Fgtp2Ojuh+i6N4nG9t3pCeyozC3C9NmxD8+tTutc
kAgPZh7jkJm94hKfaSK2YrN5ITNLblAN2ALbiuJ1BEkSPKmzRLJ4objWewHu/QB1x+3GD7ohAH1Q
cn4Y2moxTgomzdWy4QgjL8zn8YCVR6co1LAJ8OaBATbWWT+rkU83bh79AEo/LJrhcZPjJJ6dmUkU
itjOhnvWDiuxmq5g+c2b3zkZ7fSbGkOgIUlW9cYmOU5/jlOR+HpaDP/aavh22LszMOva4yFNeTeX
PaHrcEls3T/ZHcHoQE7VaJ6n0HLE73/p6nD+qXZsBiRLe0cTrVd7LJTNL4t7RQMdGie0/nNoUsQ+
yBPHMRAGSEAyFZ1LJWGFwB0THboxnb4ycGGy+09iPGy28bhwy6ozf2AwHs/kd42xdhqhJJvCGjWC
1MupGB9cTOH3fu1+oYs/fuKX7aA7tClxynAKnHKSMop+VTAGMv8NubZoiD86/ZR6ZLYVYU0tLQub
0QK7h3nGr5W2h/BzPOmLb10ePKLjH4fSQLp+FgdEHxjYB/+gv5zuJ4GqZCAvcjJPKorx9DZuPN8W
hJupkpX2/BSvg7wOed6eKvCsEvmwSLSas66i/knVhRA2WPD1bDLIJkMKKGxEvz4Flnh64k0A/uhD
88TI24Gn8l077XoDob7JT3ITb3Az2CjsQM2TMRfVsF9iZN+hRHTPgvXifhLXLxEmsuw5Fjefa+d/
RaX+4lrF9AtaQCm0O3n1MbbTWCtD34E6daq2ha32uq13zVqNzaavcLH9cowDAyEtrErxyGGUuv8x
roh7WswszVdQdmW/XE6Hsowh2ynqPKkLPJlLc2AErsd9oRMYps/4ARP4HJ/DE3H3UVfM7LKR8Ugu
6+dz7xVmaX4f73/2A5uRAuuu3GhJHC2MwjXaNsus3uQndT9TsghLld31RBAzgHs+lafwCyfDNg4A
KzrUgTfLvkvHKJX5Xw7KQK5V2LMJCATcR60dItMbMPzzT/67wC004KDfQkSwTUvG/9s6wdrXZzBN
PBpn6eRi+MYWVF3NDIV0TQci+Af06+5QVkmimhU77R96yeRgarFF6G7wMTo6AGeTtOo1tpfgSV2D
v07F2ZwlnRkUhvo9DvPDE3W83L072DbSLK1mrDKTjaK0XuXdlEuDUaaLAyc8ZHWZfp5lbduMjrpu
GCT3VO3z/GoFQcPEgO2Qm0UAFaBDrqgJzqtcG1aAzADTiskuiIlwo8kj+FmjYxj25fYXZDLmwXRs
fqqPfoDWk3znpE3vL/rJVMwWdyHCCngGK2/EEQOtPHKHvBDmY3/c2K1nm6pjIzeVXL7iTuDTELBT
fBQI3azskVm6n+09fSnGFJ50c55pVVTPi8JnOHOMpou8vpvKJCUSs1YzSM1o965SStE7QqtovN/Q
9wkubVptp1k5TRTiRa+cQ3xoohDVHHd3katRJ0ghneNPgb41jd4dFU8Uus4W0IqTH2dA87VY+kxi
Fs868DyVYKC0RHWJeMJpascURpj24jkQn5IVhSshcdcwBLmxNMq4xcjpSqtR6ATz7BbJpkGYCeE3
T/kQAuIOdgEzi7QqDV6tkwABprWP54mZ/t42TunGqjCqk/y/IC8DTaMyOsqbpRWzlfiz3GX9BQqZ
WbNBiOnW5QeqEUzOcGtsdYKLzxl5ApSP0+UGEgELg9kWRBvY2GJsbffBG8i2VICatspjVUVP4pgX
pLSDqOIw7N6mb8/VAgD9h6zMp4sW3U1DrHJ8+/fejuA6wC810E+v77GHbNrgTmgY6jVVW6dxbYRo
11YC8DQSy4Q03p+JQWrQ0aji5nHD74vKuwj/8+VYj3mYVihRH52+XaLnN8HRiQAFvZmGiGn2MFdO
RwHK6ZtYtZmSeB199q7JtXqiPxRWUHZINnGI4rijCXD1/LYJorlvjisEGWnIZJ0c/in1M56GCrmz
xFlY/K7kyXYelBZW5r1kPdMUzlGI/DH+4H+vUtdwATj3nx32ZBNr1a+tJ8q9YP9F0oq5+eCjDCMX
IsCq+CmK/qQ3LDSL+xil80g2XmVpR4nX4XWlU1ENJUV/44cwNmHB0UTUVRjVsj7mnt3Hu6rqrjEC
5v94UwpD1qtZi4VuPlmBmrsRPP96RxVqZ8Aht4vjL4j7BONyQS5Uu4pRKqDwtQraI5ea6VXs/mBM
KJJUCQ3FT/WOpCrrQESMqYHhTIeDnsmPPuu54KlY5vePrVQgL0rsE21O5tfx3nlV75D9y5rFpbz0
USlkv1LvMqVsTNBRZd96E2aJeA3oaND5dM+UVa0dZUdQpPD8906wNGNWZz1MFfzwjSL78MgGSNXO
JLCXPk0O9aWKUh4xJE4stdvZFvNiAIPWpbkpLd/5MIhmLV6oduiP+XAo3tmnXXcxe8jgFdc7o3CB
1OfM8+YEzfQ9M4WAuFCgZtUedmuE3ozxVedc09jVej1D32NhHwZYrhTRiJV5N5z/Rva98gbvQN6H
1wQVGgybeBsa8y/LL+EnuVbaPFFZMvMKJZqLsTzcy/q7rIYCN7NHRN78N3cIYX6n5wLlcm5h9ptY
b3VdJUCyBnDkOww/kTr/rsiR3tQ0TxfL/JY0b5EmnYnJQ7s+onmxVBHwKl2mfwHedIIzzktPA5WZ
wMdMliTd4P+L8P0hIbVupYk8QNg0eI2Jw8VwaYkB/Yuq1B8rYYemQE5MopQ11qxw41mnmamm3aO/
9Lyvr6gy2KQDc8P2H+PDC5OUQA/P1QDRS3w2u+Rh8cXyHYND7dUR80kl6Vog+VJ4fbKRVGQQccub
Ce3C+naWMvU4t97pyl5UsTUwSolIJybgRWdltZrrQCaz/THEHHJ6Fvjbn+mf0bQxBMA/gHkjILjN
0SdMI3Ty7xqLBA05aWWiChtaHCGajTZlgXReeZmy6A+MvwVUrg8HN+cw6G7CEjNeuduPKD7ra55S
tYTqhKq0zsGkSeXloLJ/vQohYamVXK8QCvBGqOkmC3jD0mOV2ZwjOCO85yx38UnBObjNQh7W0/7M
8gAzac3HAfYoZ3dp+ULsDrqri4xy/BpF8s4DfGlH6niKkCzG/L2s+U4ty1bHY8YoANNxerEs6Sqt
C+3t1flfD2ZBC8s0NVZvMMEArcNCul5xO6Qho7Hj3ntiCd5bnY37Z6HjIPU58rW85TA4pdAuTYTy
4Nt9mF02BWdsHUXx9p/bWN7Wvn5YfFJ3WELQCGyHlZBh4UKQlEK6pDh8Zt2xua5lMjqBUasiEwHM
KrXvv5JZ+jcvT2bCgdCGRT+G5iq2weZ5me+DgGQ7x+z3qmNr1R/9lPSlkeJX8jUZkWI6mYG7Y3sg
7bBctCUp8Gm4KflgrRQxSmeUFhzAyXn4ellnNjXNJ3+lir5ny8maD5GnkOBG8Fi9QRRHk5MYYViT
jLwGLFtLy1GyvggQoE6zk8t+Lh4kOQXPK9AQihb7UdYtE+qyrCGkF7ohdPjZMzLNrfyHj+4R+jy3
pUfEDQe02eelZ8/BPh6JohGg7WNRBVBBqW6/dVOYcpBqMuqwVZ636bkw0jTcZ2Ko+iP+1WIkv8f5
bYFXVPgkgFq/IERB0eEfLAkZpDNpohfVHcZecpVwdvfxteji+gnqfGNqSS+fKaqNabqYVlFwANw8
bc4s57Gx04BNWs2+5zA3uKn8tXYI0in6fJY/Zg0QzUYk6+0dh9m+wLywgn2G1bEiv7MoUeTg2czU
aQ1HxpoPLwZnvFmrzXdcALUARVyoQbMROya8VoH0q/IkYXS2nP5S/c7jTUUzVj0d7PwBTV2TiHQk
YI6vGYapb1hpnapspLqO53TSd7pKwQ8j81SyMG4uzISBC43OJtNJ5/1mz+S57+xJPgZ9udYFjB6z
waWy2LuvlifVHjKFNx4SXPDB4YHwVH1lQ+CjG7Umr7dflA8w1ZpaeaMraQ0iiVeqZwPO1s8zca4z
7gmV6TNS2s43xrKO7Cyh03LyXC3uFgRMt3zQEefIYVGbQ1KcRecOpMflSJOz1p0D/XdKdPxMe3t7
Xn2XV4zPEvpN6xr9XsK4n06LRotzYsucsa6j/RZNOGDI6C9TNXt5u0iqck/iB6DOKnlGsFr4T6Ax
R81YWTk7RoCjd7WiPkfmHTux+dhovgZhqlCQ/4pAX9ETY4luIykbnfRsxX99ZA+Z1WN75nhDRFT5
ylvpvgRescmDfNXVAYr0jubzSSm/ySi37Ne1tQhOi5mrZ539VTcppmfmwVlOH3g4Lp3a5im4JKLu
R3atfD8zBM0rdZFro8+3CU3zp6EHbjubvpMADNd8hXKFeCaWvYeDLC5esIWPcwthjr/LsHUHehto
hWzVZ+pVb+k5pqZP3j8SndDDlzWpOX+h5g7QyyOYvLwdcHnzWTqyAGFhvsRNxiRdG4buYTzjGnwG
x8HzzTbOHoqLt5kWvbv8i/CI3b8EjZuZSe27P+A5NseEH/ynWrfbs4diGlKAupScyaFcqPFR+PBG
6ewxKGZtGWvmDL2fzcT/4g5BcEScfjh97eaGPcGTGapq/TA6ooCDX9WxrQBAv/4QtQE0PK3V0uWP
K3Ou3djFKLcCBcpuMfIGC/MaZC1TLZwpBtU/mDCPPggEVf/cpBCVQ0yZFdQ8RQu+Lym6cnXvrl+q
FWs3WKci3ILq3UakKIZUF2W6mvhRo9MItnPoMeegqzo+uJdsbO8Ai5RmS3SMFXUS1o9nQfXA0oPh
svhT1575Mkt88ERsxlFhjZczD6gs7r80MhhC2AiDPeq7/JxMxcOE7wPr/8GmB+PhMWbTKeNn+jir
drtcZ+HHKD9qbYxb5ncRwO+sIfR+jRE//sjE1C5mhfNo/mlY6rKbxiJJL8mMgsM6cQEsOmGw6pPv
jwUp58vjDEuYL/6SmL8EfG8KODNBQ5wEtpPTliBBc9B6B91FoWQO3ckQvOMfEowyK2WgBtk1vECi
8dfUDWPAGZ/8wbpc2NKFrKo1H7oRIwOizOSK0DoCj8O0Q6d/Hk3zBRvc9CtG5YJfIiChf7IYGpt/
6H/uo9zTPlC5Q03S/W2S228vzWSvlSaklyl4DNaFdd5S5OcatEtxktVLcD7h2tj2QBEnBEAl1RBd
GpOBHxgboiJykhukzaqzcq0kyNmf752JAmAIApc+5IQAVH+IYWT4HL3bQNPKpQuqbo7MpGBp9U5B
CbGEYGgrpUoj6hoCfJIka4siSl4fbEJgXKFxitd9i4xlUlY7QYRHltCayGvAAVxm98xaoZ3E4Clf
SIaF/5PUElfqqyGDI4SdDdCREVbEZQddZoOyySWi8BEKL9wZTi22tATiBtwf4QvwpgDzqLFEGDe/
RbvHrAMAKRR2/b8WQTUi+ARHrfE6apntkt1iRDiB1n8tMRSl3tE+WiJyxauUDrov4hyhZHWbkhsp
3ZiKP0v6tbgHUp4slILZr/vVlKdLYnBiY5LwYJ4SN/wesiR0PqyoRah26e9dPRhZx13v63paPdfk
ORLsLejoV2jRrAIrJI7z5Pm15UyLeIsSMd2lik8Za47FrstsQJKmorRorX0JuJHbWDhLLWMR9R65
taqHvcLBcu70+1vYzBRttSwFRhoKRRtIYVVFeJ+3mBEXA4PnYx+n+b0eKZ/Tz7niEUMDin/99/XE
s4ec9uhIeEeB17F99sL98203tz6hiGLIUUQj/LbD8v0NUIBD3qrQ6tlESj1RV8b90JHq75ul1IWh
yuH2I9Fg+3XM0bUxd0TsyRtF+RM52+/9zVyMMwr4/pugP5rUn6n4hFZ81tcB7Fb7bzd0GlPXIJ7I
7Pd6RaeWLLmBUhTXNbwwjG3TZgObALoMmcHF6zS/0NozullDo84cbUd+hmdcYdrEUOF0E5QhdyiA
rgw58V8gjvrreKhav9FRVyEMgixq35NrKjQPHKz3Z2TftW2Z1Jn4Wvpq4rM7JiYTTaOMWZoIHAUx
MmZErRHrEog5jB8PAbM8er9AVTOkJOOn9Mz9Zjp9nrL9THrcIfIYhD8jcehrQVDSC325eJiWlCYT
UMR6f0AR+4yRgVQUwiiLzyPeS046wMyDKB+oZLtThGLM9KaqlOAysyFZDPPgSYW3ZygG+Hby3Bnj
tc/V6/Fro7g3GXj0LoCgH2vEljMVEJqakQ1z+1YsT0tPZj0kNymyDdR6ABEYqQmqlPtUHFTZ5kEm
Mfp8O1/Lrw9GPTeTG+1FKiZk+04qjEvfq2Koot30xZEzKWlyXnltcJsaWUVXm+Ej5EsLl+a3PKru
NRaPZe+NZ1WkL/r8GMJKbFWjduucIrmw/TWvHHGzqqdkwacN1ydwb73XH4n2U3wTNu66VYSWid4s
rWFx+Lj9U1TQsrHobKV1TZIX1aITAoozZv6racENvDvoy1XL4dqXi83YS5Y+bC+tcXvu3Gj7oUnX
NrR/Si4r8eQ1zIQILNyQf3NYCBqPgZ97YV8HZwKNz66aQ4iXuO/RMxgyglYdx3swNIbHBAQCXcsQ
+7G2WXf6kcrdx6at5qD1IC4ZUINypyXuUDqakJsmPwUpG26aNWaRYxsmDDM1lm4LhiwACgSWT9Vb
LSZmxFtFArbC7SN9CU/Dm+37lon2IjamcUsF298TT3quncbWfuL+8eKL1UldDAj53Pp0IzqS8X5i
mH4F9/eVI8taUYMwQ+B6ysPvmKKnsv+qwrnzW+c8bkBWslaoXpg9I9XuKL9yumvxxLw3KJ90iLoG
CA1papCULzjHMjZ5v45cEmtnEt7Iw52GTZx+LlPljka4Qsfrey999rnYUZw72bZIXIVpvN3axZaU
BBu2ICd5yNN0GkUyI8+vF4b8rVUsnYsBpxmVw+FomQ5pMP8JTAJociETvJnuUMHpoVkUdJDll8lp
vb829nLIQomE7dXgwQeyQRu+NcuJvu5zOQ6Rg8UeM+OruCfapgQxipcTk41KeSGfcDwjhS0tz135
ZmQkmt5cUgvJ1oo0/1v1eqwmxjxOCPfjD4aqfLXn9PbEWnIP/cNxl1DdFh/djhAISYYNIiCYMs8N
I//BWVBw/5GafYxarM/V7i80UEpmEe/OQO+ngf986HbffHtm87sCpREUxVnh5VhbRb6GwuJJbzzK
rnVvFx2ffIMjwucE/Ji8/hsIaPnU35ROTqKnOswbxtZKDhuFI2NSjiY+/Z7Yt0v1lAM29Nay6X8g
9gOYxxkbi0KOdsBvf3rCkl1hdyTS3qsjNQwx1v+ulmtL7lvGzMHo+gh8xTocd2gMyFY1EaOP6Gl5
sHnU/E2rJ4LmcpSZLHk7FSgIu0K744jQjYTd5x+ZFsGHoSd8t26i7HgZwEavvk+GJM9oeKT49vAq
OwRY2kZYmYG5J1zar4CrH0Avto8nCBkOpHVg0Kb9gv/FHXjg2wqFrfNTM6xnY9L4NsYtXGwIzJVX
AQJdlDr7O1bFRXFhCk2nd65scSRnl30RedCuVdOT8aKq8Wu6Dz4mUXbrPj2+6TeTG7zE99aoJKEd
iwlEm8pAqxIbYGbMP9vDYndf/awMiHzQgnWCWO0gk834USszvRultwOJldLLd+55BTeacv2pE0wy
7u/YfrIKhBs81P0Y8HCtIj8RANcfSwEqzDRAJd79ffehxzCC4i1UNzsoOJPiYb1wRUhCT6DAvh9e
Kyg4+PJ6xuk5E4MtZJl29sxCrFMLfe+BNLk9xrcAyzSZ9kaAhwAUKCbcTUM1Cr+iX56yAT+WlW7r
h5bm/EyuDhPsA5zGZQMN/c4sw1GJITcVnwwU2qlcZ8wfahyEeJGyog+ccdyqP5QGznsd8Tbt4wmp
qQdr2aKDvbp6IblEW3QY1H36NQsCyCKk4ntwhOUqauRCnROQIUFrfzuZdb4/ACtxMAeLPZopzbD+
jJ8dWdRhFgABwEi2rJFAwPc/U5u+m4PbgGUyNW+J4c+2DIpPDlMvh+vcpPqX3YJ8BZnFNKvT0Nn8
n2I79aXXI3FVnU4CDfXJnnDMi/OmtPULB5PPwS6NINJ0Tmdgwt/1pZEvFk79Cne3tnwbTU9fdVuD
NUdUUrBBlClFumA8z0YwlVCkXWQx/VZSSKsgTkmu7MTT+TWcrPgtfIAl8Yp1+WOcg1IY4RbdAs+9
HDNf2SYreRzAHzjdZsul8ljixKVhSXAxpha2/x7W8pp6ajDXnwPgbhMDSPRUB6q2ae723Xw1krgP
Y+R5xRh+2cA+HCJtlHEHRhNGCzndpJwW46xttBOwl3FEHjS3V76GkMZFvXPvS70aKqzgUjMR4VmX
poQzGvZjrru/YWiYPBsyVx8zT2KHb7CYyceLS5K9fJ2ThA9B0xvM+rkxqjVQd/Wi4gcGJ2QuLo+7
35w3TN+gsQk5z+wNby7UDN312Qt1WRHBLFlyPcqXYcUJ9xsH/uONHbb9rTFOk/KWZ1LacAinxCKj
W0Fr00WfOv6ft9xwOhDMQfqtcUyr1W1yKDOFojv/5D9350vUb0ynkPKEtGHbFHTVkkBBvHwYvCzk
JuF6hQ6/6/EqHpiD76H0XoqrrwnkYCZCJWx0UPWpw8stJ4jFK9K0iPVk0A6QDVPzuytqhEjgQ3Cs
StmPVmuWieH4B5dIN9c9ezZ9nDaajIqdOT7rmLBxj+ZhwfNzA9PoajaIY9hXSzexFYwn7AnFKIdo
dzMsoUu68gCZh9PXJmSGa9xDFiRmU4PH5oHJDo8/WINW1XET8xKdLyT8H4m4Sgf4nSHmAvYE32D9
mu+/D+Pk76T76ZOvxxmuI2LJWcBJKQYCe7vwonvvI2tuzQdXiRi/+DeJ/3uE4w0suDs13FkOMJse
Lmz6MfNSbaj5A2b3khGrJFwzIKpTnsXNoMB3BhNHy8sOjx7oFZne6BO/zgPF45lAkaWZ/j8Pl8GR
aR2ABT9Lka0jgQB8I3fwilI6lfPzONnxPLQyjojW1luXUUKDkXvJcmtEM03Y1mgWIw7pgwVaIVkC
VQvGVJosBGmBOTFJX5zEj5Y+P+ifQl4HQpSfBYzXN2FigBT+5WvB6+YGHOuEKD7x6d6+q07Ci4Cf
sQrOmkHHnv/tkN+OUnN/w0/T9HAVXJZEgcvPpsNT8CLIUrqnVoCGZN7h5F6PHj3/jAtmZa66vmot
5zV/x80AELz8hay9MhutCjac0JN9b7sWolSMstLiVsSkpkMIit5G5d/Zyey1RWxiEteZ24wnTueN
7RCLz6ZTrtj3/gplWgGCRH52KQqqKzM0l3pAi98iZY76RGp24hQ8nxyQ+iMNfvQTTwXWPfsxsnNm
BcpmyS1y1k2/QwqdIarbq6Jyub+t8+X4G73vh3disyJfFJmp6rnWiggq4CCMcMXrRiaX3JgIImr4
GbofnLQRqnmjmbOKubwg9LzZO1kIzXIRdt61SG7e6UnMNpQPkaGDArjkZZvso1TV8/Z2/OfczY0O
1jiDo1KaObcBYvCgQjCebOsMFfoDoe0t7WeXpc+ziS3nKrdm7rXZWHcbjwvEJzvZl4JycpDnMJfl
gpqOiKfOYV9+36UCv404zjtbeXFYsPPYRkFg3HfSQfi1G3YhhG9+brH60firB6EzIx4MP/cgM03N
rLsCe7MN31UeetRkVHxtIAy2xP5vClEsCGBUXnOnA9ZavigXwzPkIOgOBgTsSQ8aAXyart38sVfy
WSbNv5Mu2pGo7FzuSmxSlb51aSf+PvFXM9gfyqTMfq2NnL+laJXnvxbjNcGD8eOe09OEOaEY90ag
lhflTp7zcJqnYo1PZ2U3U1k2hzheskFtwJv5W3ugv9WJrwOlk6H1ijbl1cH0UUkFJayUFBICGcUE
Joxms0wnUUz5NkgK1pEQuvJgn4wlmetNeITFPFap9mhxG2hm/96r8ljyrcCS0JK1f6UZcSiLwjaO
eJi2cZkvLMPB4bLHcrpQ7PpRWKG26QxojTbKYFXEMG2oWZPYW9izhvahzVK1HdrHb3TSqlTKCeIE
SsWq+jlPBXWGzbjNsls4uWneLtrSln7gAK3rRU4bRnxA2Yh1PeoPNfblh9JwdWxbnw3uQy/zA1ee
NsMQhebsZqcCrTzBFmG0sm3Dja21Y/2GHhfQG6U/dsGw6iVgV18smbL6zA3al6P8FMY3BHUm+0Ga
XYb3dOpKoFNPK6qfGq0cDnAYnzkHYxEQrRH2w6SlP/BIYneEdsLMMXPj4aM/zoPRgF9YukZT4V7Q
PNyxQoLusS/CN7CMFT7s2QeUmFL0u3bfF/XcdhxvjE94zQ8mLsbJSaXDHZvyX8FsJg4GkBvgHUKm
E8UFRoY0ww4pNpxxlj151UvvAJ8ZgqSstjNvDqdQ3t/FBikPHmv15Qgmp5RMdmLrPXgcvx1zvySJ
icHwkh7XCFaJDYVF7HP9fV+V2jd9xtpbVbSomIyK5f786akkHV7r7LCi5hER5KfCgJG86fUfhnX4
hF3+zdPvjErTYfrc8yzqhYrvcCMXzgn4Qqb1NeOMcB8HkSTuspTC9a4e7qIlRS3GDMXDpH39Jz9W
eSsOhmPHb68w28/TvOVG9VYh555YdSKGkVQ8qTLPhdgHI0aTet7EccC63nQ9iBA79bY8/4mrnB4H
UprXvkfb2ATlcIhwyrSj+QKTQEQ+BGk1hmYMC35dsIU2R4VL4b6paHxff6DCmAuMMIG7/b7ZRUk6
e3GFwKw4P4JT2YhN7poNyLQ4qTxoU5/tq+/o9m+sfmy+u75rq8pmTy/Wl4QLzhNF8/9TDgf2g/t+
4/eEikxjE+F+pQfjpT1mYyiXbXViR4fvDHL3sWI4GkFvI1sDqdfgTjRb8dpFATJXPsL3qGwRpst5
+jTvh+lzx4XsRbnSZs33lyzAnSjqihv+eJ9Ah3LyQcyWTNZXHVygh+jStUrXYp/Jnobrx+ZH+957
wLZkr7P96KHJbg521VcSbptoA20oioyI9kiZionzDzhMTI0I2EPc7XLFjNtv/uSz2O9W/XZSqOuu
FIXT/9FDkg+I9vPLH4w+cF0emdpjyyUqktzRVnjUKdtN1Uh1IsYD+henWVEDXrlEffxfIM9FhELL
3WcRPXA/f5xmCYD6gwp2oiKGuG6DBMVVqHWaTdzb8+U3iuyurK8PSE12ngnjpA//Jmg4R23IrHJ2
/bLgruBRANMua4kJOW/UscHu4k3s+iQoYb9HQ1a7VqjRRcJUwF0S7F7GEbauOFKx/2KZp/tG+/7t
xO6ehWfWKlAKd1iMzY/0gBiOMfcVLDfGAL1MbakbJWCdw0+tXVvn3i+7k0s87u4oNgeULByfSZl8
k21PM2MGPs941Z5T6n10oFx8t0GgYqrhe4b6aAo+GiLW96GVtIGqCM2qhspugjRuq/qFoipQihxT
NQU5xGlYu89Oen7aq3jS9SZSo+douWknQR9zkbEpku9qIE5Taej6qeEIIA+1eAjsI0VtC7QNl/RA
bUXEbxhSXOpQzTUJavOHiF3wc7afRQc8YxRJg/yp97CLBsb9ANNRg7ynOD9HTVSHurIHzjOp/2k2
XMizjGF3VIPoHB8NHjuOK6GNXbobkD7eFqVBp/X2SkTLbbWG6SWAAeuv/wnBixkWc6skNIHuIBSc
RwdGNtN07Y8saWQIz7PKXyHsjRFNRxfazd3wcDB0CmPEMUitjfpMm5vg8M1njSQ6unvbgwKdPl/y
f4ISUizDesy9AuBESh/KiSLu1iSs4o2PNuXLE/ngzwJAzOk+lCyb782XzpbefFTzgeWweN5Q36z7
PDJOuAjJ7wUmMDnoNtsA0ky+Ux5K+6CfHThbSotygx++3wTk0E4q6hyvIxcqCVZjD60hIEQvAzoZ
48LtYyiRYJKGMgTBK93OCnaEzkdEDDjy9L4NDLvwoqB76Hxzwa46h6hxnrb0Wxmf13AhHB0QU3/S
EGBd2/Q7WJEUr8DZMvU5YMKiM2getu+GVwvSv+OJYrm7wwhkAAZSQzurc402bBuD2Q6t6Xl0V9Op
U0yGN5ezjgDdQf8LU9b/xi3V7Hmgz39kqmaYR3bwqyWK2wUyTQIYwqF9NRriGbm1NRewNbjqwefg
bXR0SSLeVywH6b1scAGjSMwdqiz1JRXp5R3J95/xDPt1RWm4Mu2l7oN+GxKpBwqSxs39vJp2+4dp
kXNhEi9teZ8eBCQkkaa5qM6/0eb3X+c71GhKtvo61fFb/G7DsR/HvJEqsrYXsVD9+yzwJrdF85qm
CMbwNXERSK3OaAGla95ZF6VO1IddklAoFFW+5LnfbvXIeZ4u+gfHJ0tNE1tWl4LhCU8v7BsOo9ti
UL/NUKMPDrp2djyG3t7PX5+iRZVXo5wwrvoBAXaP5Ci0OT0XDO1wG7nVcM7fkRpCu5MII661VftY
f4eRuy+cdU5lRIkqiWl32W4wWBsdXWjGU65kzBZbwdlTlxMrQ8vxmcTmCKPlBjzHnD9XTg18C4Ee
sLSgJWBtRUrz80SKuMCUG61IGaSeO03EpaW7OI1To7Agox+bEQ5aihDLun8Qrx17zUn7GzVgVrGg
pXNuMd4+5iFBf6M25a5IHaDDzm+etqnxpn5S1hN/4vPXCb6ZkYYE6EiDiRsHN7Oy906wDhPMpzoL
NyMTtizbEfoW8jcvop0t+kp/GQ5i+jnyMsHxf9fjVV4l2Lek9+0cuiuGmZTgIvIgsWBmwmRmO1XW
a77fQ6v67T8mAw4PmyKFhoBT75dQkiF9gBR6/ZRtGr4PssJ7gxIqHTYzBo9sw69qcpmUfeU8n73H
vE8iFeQA86tAkUfJ73iouh+KPB7lLubYzGehQUYyeQ6yDV/w7Wfrloa03/h+khq7r9h7aS1ai4L8
1C1vWyx1lGAM1/d/zlqph8eyDlwfmjpEz4WlqlPfgDle//psQZW+tY6JZskyTHbA/FNQDeYBR4VI
OnwG0iycPDOvBk1MV0+1hEvqEiFZHVzz/IvuyOlP9utsneJGFxiFN9Gnlu9iDWzoVVjgH5xlsCVR
1RSR7LQfkg9YLJmkRPedRtbqR08zea4PPDeMxZREtyjdstD5afjZi98iiBz+6bW1l0uzBzl4FIQo
hn3xHbZCCWGBxurrI5KM+wH00Ig9ebSmr/FbCROUnrrLWoZqvGXJ/Pz3f3AOBBlCuHpvKyuxrqJl
PMKKALr6+iNWVu9Ab/A8tim5BeNn9DDE3svj2Z9rfS3ojHqdKHmbI8JLCPj0PusLCS4YZNG5BEsL
ATk6Wc84SRo6KpGDYQ8uNb/il69JT/4yiKz3xHr2oxuY/LT4LkBbCHTpvfulEA8DaUzneoYMtL+U
vrdxbVG+/UFTuYtE95XvBwh1VuImYt0YROFEBdB6NKWRKgL3R+ODvGeD1TlUNsjT/nTLcb1oU7dj
tW3RAbcVwMcqppzdr5pB4kky1NiC5Aotjn9yzovKyAs2CF6pk8i4qYYWIoggRHYa5QRceyYZHyQW
H4aymLDwrabgbR0soFW9QAeyznBvOlc11eMnXvdYSuKey3ZpwC+3jVYNOhD7Pm6BT1shDEGwb+oW
1oW381Xk9DnEKGT9ZS2LDcRE8vZtrfhyIC53SodokTK55UppArX7ET9ralR+34B12P/Sp4W4lStA
83QEbc/6DuOSYET9PfZvPXGV6mM17RRgk9oF1aHQRsTToSSMADRos5B5yhvoRIHB5GPhBvs0viEB
G/p8XXaQXt2nlxpakvd25x8GqeqlerLJbf3nG5yyA5h09v57ZrXuKXs2xPu5HBu7rLNHj5JA2Byl
+FrH13U5pkE3Pd9/nE0L8EdeSf0/7sCBUE74wyWbhkoOkmQJZ285qyl0Fro8wJ1cBeR2l3WJEKek
8zBCKpPYo0AL1V+p9RbQ0fc1ya4uBGC8LBWv8m1USu5R3qTWdyDOwoMoAGsYBdQEtVWFruPudVgQ
235JpLlCvYfxwBylZrwFmXpJUpnMM6dGFUi1Gr7xM7Nq78e/KGfgLTnYSuyug+54yAFGGIaKawh3
lMkscYPIC4cMntFYOwdChC7g/XJCH8eJ6ASESB7ZstcQ4HUM9Cu1Wee2/aGo8wmUL9GyPnzASGPT
F4cdnNnp1ACIgM5pJafJT/hR4bzWqvZLMSsLH47GXhvyonHZZAmLEzMqyyNeCrjVaZ1SHN7YXkg7
D6dLbswCZP5l0mUXuHMW4xaDW0cyZpNHUMx6D1Zk3osm+bik31p3sLISGi2hYv1pVJli09QDLXLX
Y0KZwjoEX8fhINe1Ea7RtGtqxR6KuJjl2ZqmSiCrMVM/6sNRis+scoEAZt6F7p2dOdcZbtCV08Lb
s7WYGtjjB4LdycXih5nOyU4VyCwV1Yd1NFgYK+/oIZHZyEfw6jmrZ4gbdVshi8jgChUQaMUFzESX
ZLZQuyaZd67IxEPeo0XSEKryyxx2YRwDMpTk4eH+YaSu7qGqYC0GnBorj1dP4fJHyid6CcsGoRvT
+3Uw7jmf/21o4rEXPkg027enOB8jdVQPexhh32efPlhdpKja7v28fjDEE6xORVlquqlU8lDZWKVj
S4zo/bIZgF+hvZgZJKia3pe/au/dhf6InC6815O2KVcKfQAt/dgfeGFlUhWiyGSGEUpEDNQ2iQnM
lVYz3e/FWS6QN+ulhlxKG0b15ljFubJq0Ar/wisSo11zunhMVBB0MMaEthgnyveaPVBBPFK1gi/6
xNUROe0MEPnCDJIrBmQCNi7R2R7z2x4eAFt3EjUjP2jvKdq6DUH3R9pu85Pt2A10IbLqeaWf1O4a
EReHUG3471HCW9x8xbgR5q3Sr4Iz+ixsRFP8BEZWBAOKky38OBXa5OxYJI9fDGLo8yuRjSfP9gPN
FN6dCC/MruSbcjZ+Sv66VHNJa6ij9Ue6fNWHT6rM1YG7H19nIbCkKaY59TtNbDfxXj4XbAEkyR1q
Rn1kFdrGFebmmFXi8GViStQ1X+hnVAYGyeTIQdfFtGwUn0Q6uPFFb4m5wE8V1D7Is38OnqUXT+AY
tMk0BD7oBX7Surhu6sbxDfbkN1vE9CqKzY1hZoY0a+5e6vtY2qUKRnFyTyf2kvsdCe7XBLuP5HTI
jusOJ9GcOnrKDTdSA1F3HZaRGTv72j3YHJhkVRge9/D5RtuCve/JaiBisM8/9ZyCKyDWexab2LES
+XtW4tbU3T1QEJTyTh45ktLO5vthNE1vZ6iPR+tocYU064Pr+NwoBLusjPybqnclUX+XGHGpMAY6
X4CPO1Mgx9buEs8vo5X+asnYuTT6eCumCahcynvkYOmUKIuMApZCscrFJIPkia4tcGlwnSU/g1Vk
xJ+aBHoixg7yN0dMZpXxPUx68oV58GdCZraMapwETPN1QbiUuTnmYuu5TYYZzoMzzPJFL79vAIDx
lHC3MFhzFrD+Ba9dr29yzPA3KXVSE23gg8s0ZW2pf3y+w4r6zwJEtddY51X9h38BPq5ms5dq3pb0
ty2o1LEhoHVFCEh5Up0aqPGPHvRiFRTMA7CCGD4ZRuZpRoPFk6psyI+hiBzgceyVdnVZiQPhOHfJ
tLrTjyQ8yrKnHD7vfrle7FcFcUJn6u21srkcfL/0p+EXeZyp4zBGuQEOLYCnV2iKvhqLTTBuWdP4
9ojmPIyOIEzeYeWb+usAynpCxVPWvXpTmPt4ZbrY2/YK+FX1ufwQHG502QkG5gviukdVbI5llh+i
F1roMA23DQCnIvwjcgFpWv8ohORWS+yAszAnOMRYdwHsFm9hCg2HN3Uaz+ReUS1H7mlmTHHJi5FM
SW/lQhCx2gP6GcXkKYC6Rs84qB0/1VuGxd/1YhpYor0d6nbDZgQgKVigQ+x0mKfqXDTXb+IbzKI0
K/mJ1UsVsBVpeWnjd2GMbmGq1yo3SBUE19MhUnO6VUnTpZF3yF38VrAJ1Xr/dP6SRptnBUAUD6Mi
c9QFtdGTeZeFNK3UirTnENCm+OjBLnylZw8HUpwOrDPe4/1kMDfFeZFOUIuJmpTwqLOad05CThu3
4TTF+fMRBFmJHcK/lIkW+jY1H5vB4qdOp8fOp0wEYRxePXxyA4leKwV3kncpRSqHxSYPex3mwKdk
43+SP8nwzRSGJOqv986M27eEn8XAW89jvlRCcieSgUECw2YxPos0v6xeNPbwXgxK+S6BE4jnFpCa
1PmtA3dtOGU/2cdG7IMNx+zVtxTjm6jGSvRr6wFMkqh/04VoyWnd+ero5p3vAHpPLfJYWBx9+5ga
mhUJl8gKPA4Iyr4eP4AC1UtEy9mX/8dacSJ6zrqPnEIhir7mZDsaSGhSy5Vb47Lgpnn+SrPl4AhI
Rp3YdFyFiCBAlc7xfwmnKpC0VXNCfPxVXdvg/jpD1a14D6aFNqUEGQwB4xS+YrIXn5vI+zMY4sNh
c8KoY84Qp5GMsvAkZDg3hgWKQWZpPzAfr+DAGHxoqGDiACeC5mcgH/lPQ6QHaj3A4COoCS7wQVu8
UQLpiWRfoNYkJpwxVjkSsReTm2u4Ts08J+O9hwSKK8YeN/zmxzuYpCWfwglBLRQu7cX34xEuLKQs
dOE4GHykibPaz9STmbDpWb1qy5TrsRNUFaOkqHRc2rYrjDcvZe0cCIVQIPg5McRDcEHODIlEAHKT
36v3nG3RrTW5B7Nt19POXdcjY8Gu7JKdvU5TP7Ed4zuTgQo5R6+ABZlEQDkDLFEM3JU54iamGCHp
hx3VxrYNrj60HaQ2vW9FxA+0qn+cMsARUPR+aE6Fw2S/m5RikF7/sQzVEc1II4fl8Lu4c7BO+za4
msmaRZID4RSe0dgkIIvEZTTh8Mzy1A5yL0c5Jvl+X0W7q3JBI6LsAlvPeSfzO9XsV8gnteRBe4al
IVz4iOuUt2h94fICJgWwYGF8jXmep1JpD8071UvaXBgtV3/a5B9PB/1g9PI1J/Afp6cCyFHB7ztW
p+J00trIUsFNMCP2/QGBDhoFsfH49tIl/aiEmFJVtbw0llWmz3LhLlc+ZSHOJjlD4kbM2eoOkCDn
G1goC7w3wo/YTx6Xvt8jpisc7rfXXtxD0oMpMghRLKO/8BtFWbbv3dWn9bc9ad0t1+8S2o0p5VRG
ExWRhLLynrNoLU/OBY6IDvxplQdr0wLRFFpD3YiW81nnppLjheRJeiLywwFB8j9uMu2A3GcEq6F4
XuiFIUEB+UCZcdyVVXIVrQiFS+dWR+ZEKvYF4yX3U8xfMJhk0BIGDjw7yz+kgu1A8i+PyHWBG2UE
ltp58GpFnzWL+vQbRQMHV0GxlmHdwdSNBqgZFn7MQSVLy4xS7z775DSMZ+cQ9DdueQxdCVq4CtV5
zhZ4rs7RQm9LiDEDt1XrbvYuzr9drBL+xAK/uR240+2yKHwG7h28Es7PaGh6CUdmuCoQCAosf/H9
xPmEmhq28yGDImztdHnCbwJc2ven0sII/6CRRkZuQVQA12gi8+l9E2PJ/lcceNiqC6HIzFzVkTUK
o6k+oRNJs0iab2/u1JEwnptTZ7Vhlq8MVjj/Ft9dZ37BaWmdKo7ZSa789v5MSqCfbVnHo36Wo24K
9pXhmv7hEkw/E4+cz1uGQ0vCQkx1vrnLPuWTBUvh2gPCfRsmvn9MFLwY7Lzaq5EnVO963KwGxxaP
9RMyJpVPFK7m/y+ddNIW0gZZ6rTl2Xen95vZNItgbKAmjZklV5fEuk6CQperVEcvMW1ICr6/mS3i
7euS/ok3b69ZY7+vfe9mrKUd0isqNR4/74pW/FZ8WnMs912HYB1ZJoPBrW+50RpcIi1X9Qk2sruD
zxDHYwthpQ3Emcne5aIwlk8esRei1YmudNEygHECvujt3sm2eEgU72rpP+kNEY3pw7d2ppJSuv1x
i+5buHsbn9E4VKOa7ZVX03NbxThzWfFWErC4btRY76wUKxAL/MDxo1It1+xaHf4Fv8ZIvmCpM0bb
pQm58LwZzSID+e4gyZ5HpKW/nG29iGiqw9agWHZ10PNA2fJPy2cP+qgPlpcYpoqkE1dyk7h7YQsy
QrhSyCeR2/0VjwN3tnR53rOpMrW18KEZwSUrIPTjn0G0GbybiCy+KLARzwwkH1VbjcH3J0QGdMXd
XoETLvzOhms4RSvh8MnbnBmWC+JQbROGuu9LOpY/kO+4QU6kSOwTyU82ndlH7yMMxh//ERg6iJDx
H4ipcUH6HOBQ/XusmynVa2gBo0ZFDXD1zDIdoJBkd5SVblPmk80GH8HRoply6TImOjk8Kd/S0+h2
9Hti46v1XLgDM1qPYt79ISwPTtA0JKE9oBG1tzP7gIAAPPbkfIswZkfxUrpyVgMnrRHf5oOPp5jj
bvTHRnZt25m8l6PEzf2X8278rDxlaj0Aq2yGLKqobrklGjIkzlD8/Ou4ryvB5OqHKHN7h5hTiMWQ
f6tQm6MEd6F14tg/ooa+EAo53AabLSKM2qoa4UaaMEBzMKwwiWP3hOLWi7lBAzBSwU6wgDnE4LWB
zy7YxKXXuR54MzDm6/8wMEV8vq19xZCxkUbVRw8ggJrHoq/dCyv5oAh+7i7Op236BcqbMSeeX1Xf
PjFOvAv8GD4FTvs9tIcEqizPEnJirwBEKd5OQEuyAIZUOTpgN+ZhFdVa9NFJthv+gxqRZNNdhfwV
pP1ogaIXrQ2ocCueCA0vgBk+S1+VRdTRrBsySx5sSdcnf2Qj2MghVyWuNXEgPyuK0j8X4sECIgJs
jUYAI2uCdzsXh3zm7zpS+POTaFmdRKMg4JYcTkPWQVsN2jFRPtlUMswv4202ucSvaH0R2wohkXcW
OYp0tlhQkh1RnvZSxZGeg5Fzk0hisuqtclhTAQhXWZg8/k0usc+z44IM46pSWnv8xPi0t23ogPF9
nSkH3P0ZQluJKT4NE6Emd7fVtbY/f5NDju2Mq4Egmyxtsr5FhyDqkYdpdmpcJ68fgy2LFuxH4BUc
HSu8TxO9L3EQVcVndYvRGzgsfQHbmCyMMy8q2LSlhtuvi0ejTyc3wAMVWEQZggImUWBSEP1ZtOxu
TkJCNILnUXdS8UHqp++IVzYAA0A78UjZg03Z1Q1uxJsEJwQ8aB1Q18X57w9Nu8cnZX5WXwG7TTcK
16Hv1bO9bUm7P7nrdSILVbWh6f560Xpx10ypW7aN4rRLBQZD5eH4TIMvSvZgD4Gv78KJ+RBoJbVE
gXuz8set//yuL37+vYAUb5PylxHCBzOb7lEPGaM1CdKpatm9w1Bbsk5hnEXD66IGZ6BgpziNEhTP
d+QOnb2QjuWYNkV7z248O40ir3MC8q3r3nNeVaSek3fZr9lnXLYC6d6P92/24mpYD9cMej9ZccUD
T3mzz+wNfkq03DmGucRxnGjRx2wl/249lUA8EWw/VozYKSZfsuXO8NauwiLbuOHdRTuADueIVHCs
uDKjNGzmG43N6fpx2R0i6sVqtYh8CrLidhm15lCVxYVc57e8NJeQEogr0a/Fxq1qnNE1XdcFisKI
idgmPq1PIDoj1LrhjIMj+gUGLCc4LlAqlK1x6//tAZip0UQknB2YyfJFNpYn1VLGmNgQNbwJxhSL
Trutncgp+0AJfz6CbFJHYgV1WzSnerJfR6+BVoS3tWvAgYnZ/B9DXGUMWjamIkvNjWO0D2Wrmd4S
zprCpHFudWMb5hbF3CO1zyklahpx66FzrDw9Ii9qmwaPJ+957BtzZltr6+cbXuB9QYOcjk2/Wi2j
9+qy14hGx5s0Cqj3Y8lRgl4IJ9C6JZvYiO6CKrN+11IWFRTp5pE6ycf2Voyy2JoKLS+Oy5yvhjrA
tASehwj+4GtN22eHZJ75TEZOOCq8geYFRQmK2FP4QmkHjtQ2rcrkQR87prdRAnVPcXZBVncpWe+j
MNhbAuIpBJxNOk1KJfml0g8I0l/6+wybr0OdItc4z/j21eti+qsLMSWrj12/Hl9BDZh8NQ+yyFcb
cALWGqsiO3QTz7DQ2p5mgU1LUx/vL2x4K/nFlTixGoQuaMAYzGahJy19KZ3Zzf2FHeMZEpaUqT1O
tUtoJUaHJpYGxRT7qjf55myj+c2XUlKP9Q/Q7mIj+fBWNzHrHO+RvSTZW0C3z3Be0DkZpI3C4u2m
9MDVjVN+QPICep/zz0gGiFZpRh6nyIYe2MqYykUGbI4wOxTPE7MlNG5ufIypQGsy8tI+L6BeTPQZ
i7qAxlWmYxvgyX0Ll9oz+Asl8obvAquOvXHbYfiUhcDuRUKdSmDVacSF9akI/SJIsREsywzWmNUD
vqUHIFZQuvSOeXkAZsgcZhqyoJg7IBaq3A8o+/1gifDLX1FYFbePXD7XDOa5q8vRFCt1O2PjZR9U
NDRp+kGSqu16TEjq+eTMD7r+f2vCBfNdBL0uNO01fA+8IgmitkU4vjHMzdfyqsknSgyBf+ZbPsro
VCjt6p2gt9/JhR/9UfUko0y3nNZgHhdJTDuf9QfrIuQWqSvUc2sqJt+R0LVTZNrwjP/0aVbk7KH8
oAulCMvequYRRRMdTl2Eop9YAE7i56tQ5idE7vJxC3RqBcKMCEgja9XX4eg62hhCkmK5jLWvF7iS
8GPC4d69rE6bNuq3mkdlZZrlncbqbvIRdgVHmmGQUwmd04fDgz5rUgZg4kqfeG0/8c4KlZ28Gskc
qGQDmrtZs0TLby0KlkBir0oF1aJt6rGcbIN7g0RD86TSlqIm4ewB4zYmDqS+k5SjueRfUWSQu2/d
jSKk1PD6sw8FvVHGbnELcBs0QIVeLX8cjajysVigu2Eyl7rgaRLO+4z5HnAzIcJif/QwvuWp8R8U
qHkr9ijAhGTN4nb985EQy3nBI4B8gztT8OgiQ3QTJLYryn8Rsb1QSPf4PvxBGtacorKmeQWLXxXg
uh4pWFyKyWxbBe65pAaUwYmODf48CWEmqBVUo+JYL6mNVA6CNRV5mmzVssXSd1o2L2Zz4jH9N62M
LDCd60iJV7u30MikRNKubDa8DwrW/5xVOPmwXjIuth4sed7Qaz6Uwbgl7KKrzTSgPPgvN4YghDAI
tPEFDxol164JrKOWsktCwrVA7pHGVXEWg6PqeDyT9yCc2rMmiN1xw4qJJmQFO1nhJeFr/BattLX3
EnG5XjshZH23al1QNgsRqXni/fTDjc2XZVeYLfiX0sETjoKNvSIIow/k5XyO7p2odU9pghQWJScc
F6BJ5uiG+G0Ww8baX0A8ycHv7CnhAdOwmb+Fa+qQOQHcCMyjYMbLhE99nMt91yJazQdK92UNTVNu
OEa0mIN3R1XIxhwXyLGfNVqzGfbVF1CjUodoXvQ3x23OPienw/kjS7rFBavtAXQNgx8qTgBY7aNE
2Gv4G495u6A9JZuOuzqJIPGDLQecEEzkwE//B18n/YjsNjLc7Y/GhqG0clSmabej9N6g1T0GQTlq
dycTEKSIbY0fN9bgTpvjP+OIlKTc8+tB34xTBR7ZT1xHErole0S4kYVjZTG6IArdvYfm+moJlodA
yHSVcdzAInBOtGrc2tll3bflcjrlYPnFGFoJ9JLlJDSGJ+7Vlwhq+k14UJfucyXNkTtXMdIgRO9U
oc6VWupwkeD3f4AU8LJrfhQaH2pWYYFy4jsyMsx3Af7DlVe7TxzdZreqQ6DkWvx9LIB5nwtQXHNL
r9nh7OCsy3U5GCD2H67cM7naIk6Zp6v42sxn2w2beOHkj6xwW4xHIMfEpK7BvMed1oiSB92zh+5n
GfeuK8ufrLpSXWWsbpxWoNnpg35Rfxc+QLm7YgkqHPjfbD6tWP6OQZWfbuC+o1m5t8F/OIqSAgYe
lBi7qXv9ggo+v1iZ2xhj/NZ4xgcZfHoIeo20ukM6Qs0P89pg/HaKnVkwcXqaqomiebUAfCbZJcfO
3h+alWboYfelkocxNGlRDJOYk5t92swTRpNuOj5BVG7Vm3FsK19NupLdlzlM9akdZIOkkx+NtluE
3VyKAso8llcnNj+r5tvGq/k5ZxWyrmwAoL0IwEIzflWcReR6h+PhbIu/Wlqci6qwjdPNAadP5MMD
4490jGqw9/XqThhjp1/eq00iP3nmqlsV80uByz7e0MIlLgn8Zg8LTx31VD1IQZxtualGIGasgRL6
CXZ0PgZIUQ0a1WCONcu95iNvupujJMjY2vbFCkSuh9VOMmE1IhYsuFI7b6TH4b+xayGExU2zy1M/
MFmJPu7urUOkLOGb/8pq9lDTHY/9TiV4RR7VvYEb9DLrHpYsqSMckzH/Rd9Z3yCv6F5BCLf9GEdM
zK8QGkn/gSynmiCcOgKyjpjSwC//vSfpQFyUQQodv4st+Tcz3MbOaKVL5AgzvaxKCFrk+cj+tnxZ
1mQKm9EnKgcz4ylvIyEdkQNZQth2uEogso28uv7JSyIdBoUPykASDOZJGofjh4k/IYHijynUqRnj
OPQFDjVHI3mQoipCDna8VmothNIpve/t2WmIL18XWMOHKgCTOOWX+QfW34dGjVC7E0lBBBbixBy3
fLttv/z6g+ZYSZoYW9uzU9sI5M4uP+q+cVH+yafuulHK9tNSQFzKOH/YpqR4r16CpVxowWK+g2Hd
A5n8I6hXBuBCGN297iTpmvONXSmsf/Kwany+TAopNbeJJ7IRch+0hl5ghLeULp3AvkXOOdwcZTor
Zr+JdgWsUmN7C/tmZtUR2jzs7qWopGv7T7JOy13ui9g54uUItA6Nr3OJXedPfkKgflZ0M2MAFomv
4LsKpnh2sWuJmQwAKsLs1TErxLF1BcQmv5tMiM1VxBodJqrcXOhGNUv3YiHzYv0Qf6/mx+0H8tww
UhPV4vu6ROPGGz+GNcOVSx4hAbD9dcRJB4Osfwc4+CKfxjPa6oXsrcUUhMhGVBS85tcrEM7Ye/lL
zKMuc1pDxVOEGxMVQooyvMSpiDy4HRC+gHptZ3VYe2j8TStbUabsdwo15s2g4s8tJFG7YF1xTU2f
iL2lsSXXPaNKX/3pazJrHoUJrUCIMY4WjcvJovagjgjA6jMufoTn2mALbJ++OuKWJ4QHIsU9Tq8A
vbbd5P26BTVVyCW4GIMJjsaSVQJjEYKvdFaZx7eNW9QGTjZk+cYTjZ8PVgIwmYO2G64zypLHEJZK
Q9RtAFkKuB51vwcB7AXiL2zzW0dJCwO1sC+CuIj9R4G9aWZ3kxW5BV/cUkzEAJ6rK2QnR3Hu6rsG
uYtAXwMubc50HX8MBTr1JeVm097EAJnLwn9YAIZV4DPM4NURvNfLvHEDbSfuAwvguLCMY0LyEOuS
E86Jeqa/f2WnkkckKTeWmXIv+xXIqb8QNnYMBmfBRBARbufMJVVKYauUlVO25kEPo8CasSHKiVKK
Gwo7ToOAXn3Yb8QBZQGb31V+fxI0GE3jtVqNOzFszYZjX0yrX9MhLWIxvO+Kqc3xSc4byoeqKVlU
gMw+htc6sWfH0JYAeL9xtWQJGjgmfTiE/RQ8vsNbMvZM/zse2hqmomL59LZh+smbxl3ZkZpXJlwZ
uhBqGRObd64xfOQlze2bx3EDpbZDaAIruAXp1xM1GNr+65+dBjNloYM4OR4CzhfpiDdGjmRt5Exm
p0Bm4OYKxcO53SQMy9SIK22l7SvSEaT+EH6MNT4PMhQKtaNag7grxRgzDUEc3N6gmAC2bZQlOqAg
4fI66ueOXcdrKQG/5vMKvQH439dP5iGABMVhWbyFlpWLSzQTKn+qX2IC0tUgbHGNOUTW0bSu+rCw
8g1TGjlxXxINJxUNt4CyyzlJtOLZFBHs6no91/izL6CIr6SAM6FsCeHgDhVXUHiIw/wnIPIVLEal
/JhACUzfVc57MG5NsLIlp9XHTMf/cxuQPjUb9t49/Cf+oSd2Wq7nuUib2rwfKBMomSh16q9nB1WM
SvG9m6AfgNo2RCLhoruUo2HrAS8yh00EBtxYi/OUFjqZjA9y8L+QWJkvejSxItHDAAwQJndX60J1
/JCtq7pUt0jAsTaMCxj4FYvKi7IHk6RcvQefzO49VjEgs6LJzIss0lk7VQmARI1TGLBoblKrHajX
BymlY/c/mNrNzctZJ0twAe+NEObCxU0p4icGYOSXrCRW1hRnDFygO8LXv4ByEZY0jeMGGFbE5Vnu
Pq1lZuhmuHHhk/tBq7iXnP3Ds1PEUAICAaVENVmp8dCJbD6AUrRTIuWMNyo6zcNYrnfYYNKKPovc
RPhWT9WOVYfyxMf5J/BWyUJ9eXDdXFXKA2zKrXFQ9GWVPX+moTq1nrMfMnJrXot87XuZOY+chxc8
haW9m4In6OOiGUgTe0h5HrZqxyKgwMPMmCIpOnH/IwQDKAI8HodqQn0GD6qg0nnbm2nHtaRsbUu6
Yls+GFrOOtupKnu7rTKE2PxC8KRUukXhao+fsK/YJVo2IWpHPxQalc1Axbd2Xf7OnbjauKq6nu4d
evSEJ6VsXcnWCaABUHu3rC3rVlOoda97D4SKX4jHxNkVRTzGS3uHRbsEP9/3q3HXpsC76aKj1b6W
A0gLa6PnLoYB6JmfJbJPFqecz3scGrQEDOlRWJes1Va0qxuJVNK6cOYkP00HMUWpylO7zUdYvBJf
eRxO8kEMI3WBgV0PMALn1Jm8PaQuqEsSBXm8cT5oXoJhsK6jx/4GMepJqSp4unf3Sk9XCR2rHx9a
Q1R8WuPC5SworJrnfSZClZIU1+QVySUhH6yf1D4HNVej/Ukh/tRiTeJ6Mtk2/rsibu1GajICQ/xP
tH4u/XgkMmhI4vImQIPkfEfQA2jJ39+UdlSaLyMWMPYYV1B2rhovVGx5pKaOgJpMqUbozsWYhCaK
bmFPs/ZlqB6pli4znAy5OYk6eKJmFAxjC82PkCQ3MOzD6epE/P+aAexmB05Ojoedq/7BYpqey7pS
+D+skwcYPRdZWMg9s8OGPkDgVKCTDcxkigEDJorFAcd3awr7Xbmn+IW1fdmdiKXvNqkdcFDTh0YR
6gKA2bvzVvPp0v5O2Dk0RvilOlSXLSlItgMHbeGbLIfNzE7LDB8/NHbLgzxTBVglEGlZBU5achi+
B9fdf3nMbmBpRnHQhbUlLQ78FjZT691Pu2Wbneex/KEY14ahATCrpe15ozhRbmNhUYD9sUXKp4kW
gve2+EjjjIDnoqfrqLyeP4BVjG/Dek2i8mZZchlKY9PEvcLV1/iTDYqiseDj3rKJ6Pdalb8vbtj1
TrcczbRvSVvW0Ao33xjPKzuoCoUknXdrTaRygOLY8RRBAfcf71CvQ5Jek4uPRKI86w7aGuzCM1EU
i9DENmRpvTh9TeLFg6/jUy3g3xroMUgeP3aRzFtV/d8xMx+uZjE0WVf3cVlJP442PHm5pcMolJ6P
xt6Z5wDhXGDG80nGaJJIo7BKIbEX7Th12fZL5AjdZtx+BOVFozU8cWNlGZ3/uvY7eCvLTE71q/IM
6eHKrmW1S2/8OSa9+W70MNJKO7EsW5y79n1tkjp18qNtlrGJlXzMNmrpJxEc/0afQoGPSFbQjJPU
D5Q2Taw7K/C+UUxlYLUV5fAow0eZSdtmjM9wvQbyPmL7ZhEhjv9zCPJBOL1i0+cq/ZmB7ryEJCY0
UvMet5G/1Awcx5nm7SAhc9HROzUw789ks2QAG/FZRG/pKkUpvE49TkqZt6kOMxnVPDaeP7rvrDan
+oXYi4x8b/NPIBhtwS3Uk8QaKnz4OaODtBDj0qYJ6axrr3f6rKhpxAh829BGsIq/RNZewXVqsf6K
BXrOW9e990TqPTDDHhgcpvdd/p5AxA7lU6BztrPhvK+oyKeap7IUxqmxQpWUJpGn4asuDL2be/Vg
snQgmQ2vVn2MR1Gsp5bhjqMBSlbars2tESSzuJ6wSWeEQEHT0PPYGrSRqs6+Iw61quM/eidh8/UG
8PXeCyYgZS/EbHMJNvtUvr8hEyyw2gFUehDnEF/rRWzPvXM/PGk3Vcf/SEoRKBLpdmcSwn13wQq3
TO1EHTCN+AER/coR3ngUD8Cubkl3fimUBoVVlto5hy09uffEDAJILEBpsfJvX/Xq/YMEJSmI7w5A
O+VAPCi5hJxTEIM2RS71I40xC204ScETIzTF98RelIn+GEnZ4vDWN83SlpTybN3YdTDTbAQ5AMlq
MHPbbnYRSsUjdBkK4er4DQljY52JA+tafHr2IZQO2EOLeUlqCDTSzPI7/r1Wbt5uB4eDWYuVlfRm
+Xk8hsOvrLwuBLxRiUWaQlKQnLopv3zaxh25JuKnAUH69lbveeIJfHq/cbY1VtKgQiSFqYTePrr7
/f7bLaKHuc2MsT627AvTcWC6b6F6kN0ltwbjgpSFdvimwXC63jMZX5aFl+/Xd0kiktoA48LGcqPB
nmlujOn/a3aDyWIQptRxvPzMx4lkKF2YCQLOneMwuTNJA59rhbXeOOW8uQpDm34RMUVYmffjcq4g
K7wbat++xMTD5U9Sqw1IafRtp7brGyqW0NKkX5W9knfKIH4HpqHS7rpdLrGR7tYr2n3vAKMHoqf2
zAiX/c0Sq77IXqLgANEZ8mk7Rzq13SgVwwSwtFQ3n8lPuWgeHHo7GsKal3cvxEnssGssYbGM7Hic
H2Sxa3DwzDnqxOIwizlklF0gUf88glSI75hrWqPEMVdEK4XGtD+Lx8xXo3+GDREJE951VgcvUD7V
pPtHD/gLsezLbQk46t+VWYW4EkMTqnszZOXD7/LiNN9Xd3IJdrl2WC0uMz7fnJJAYum+LdkLYiaJ
qugqsSrEWrU7o0y++KIDiXz+6X2pDoOdKQc2VmATNHzYYFH44vqPt671DN/x3TpgA277o1rdDd7P
uM9CqR7k1cjI16LivMorEl98azUnDpZ9R9YOauLu0bOnDS/to/0wWp8szGuzZUEJa+Zjd8oVtIe6
32H+WPrPd4+/2w8nfTGbcL/WAeFxAvp610pl4RDd+9aeYl5N6y2M7HVDZz60hOtgVc6W4/E+hOZA
Sy+7VN9H2kyDs9leo8CgN4ZvXc1dYUsfynRfbvqHU/jO2mOaDf+9GhcXQ6z/DxvXh8mMvhOv9q18
374CjrXZ0p49LAUP/oJHD0L0TZ06LTtTXzJgXN0nKTkrUIe+L4DhiNvfDpIc3QwA0Drc6UAgyBhd
mcns0DncypbkXatqktieA+y7Wgmaf0zoQomFIGmVCBjIrSisKEcAA4vIOHjv9DmYFgaNvc2GFFtn
RLtoBkr+Cfq12S2U1LiDoEPy/R2nEW4YB1xDBqwnKYGeBCCKs0eqm8NzGtXA/L0UR/6H5bizFUfk
Fy3IlCBKRrVH7PNf2BGUETH3AOQn69hyVhFBAu5aaB5oSwaW3jIjaCl7JS3Vy6/+f1j6DTzfw3UY
Y+dic43ZwXQswQ1AkW8IiXqqS1A2vy6ER6vNOLEVqdSBJ7Zhm96pbrIONhafIh/+hnXLJ3rZFY5/
mjhVjeYlTyp6uqOT0xn57/TOiJ7pBFv/AXRUwUpaoh6xcOzhaPfbRyQKm6l4Eehz/IqJzZvYawKh
98Z3Bh9w4iJstt0Wp8f8eraPv83JzZQuvTiyhLARU2Edw92s1EvU2Jjdzc0n1r0VAq2p12PIWDM6
PKoFkYSzMV79+UX+KuLrwVwoRrMwhFR9VJbY2oFj4hJsrGdk9nx/C+cqx4zzge03ZmBCpa8JioAU
4baz8T2jkSjtszh6rXU9lZi3WkF2BSHtbCzkJadPrh1Exc3YnrOIajMGNtyjJC9es5ZiJ9KgBLmI
0XbujeHIM8qTgxlBlkedLMq5eOX3RrOWoWF1fftoAbWMP1hL9ysjHoQI2DssRdVmOJsx0H1ItvEn
T2ef9wplPOmC2Wz46MlmWFssaJnYsqgRAhLDkzQ0J10nRvY0qsyB1rIuInnY2CsW/vlfE/yBSH0M
Dc93BXF9uxD4bGvi2uiiUbNQucexgDw5Is9iNHpYXm5VTHY81wY/gMKANYVbKafaXihW8dwXszsy
+x8sxwjMdos4ejnJrmGtvhvwbhDWfCQ7ESR5cA7qVd+QZsCIS3QRoydn8stq7am4i7Umkwjp1NJ+
KnQ4950Bzy3D3wjFLMA+4jXW4mg8HIZYDBtkaEFahjwXbJTETm1fDZry0QEBdMnQNIXSfyvzvAH2
0MhOAz3jeICKbiEIXmew/nkFF1d4+UIb3KbxcAPifIuwaAkhKYbquIzQ2hV6SiXgv1B/9NwglTKB
q18Vcn3M5Kisz4jXn2ihh+9nUG2ch5c8Qgux83/ARSDJTV64HYwrDQhqyzx/ZUqum+IMdnshFcpc
ncUYDXN1Z8p7AKjrY9dHmcsgAe4E1Cw0L3myrnYPP52PpMJsHtZuTYuV67edg6Wyj3EPIO2h27eC
cqRPKbKldW8C/sHCtnQnKIeYw7NjljhWO/hNEwqe0cN3wW1re8TwsAx74wlfvkHdmZca1W4Ioqv5
m+zhAST6g3sUgR+KZf12IYzsNeFKVG1Z7BdSauR2qQqwSGFkzmKnw32riPP5lhL+/dBrozl9H6qd
jJiIJK2m2zSOIgMUbyy1S+t9n/aj7+KIFhIPAwvSmbPitAvP+k6kk1kv1F5Rc5XRiLYnF1E3R3xj
j4wC2kmsiGoGd3FS70LtcNBDUV46bpNzUJoqgSQKqazELHKkHKJHQaYIh8WrB/uB6goDyxPNCuPf
uYPM763lsxVNCqAUxVR2YDgmt7zzpgaynyBjTgU0fv+jzahMBIWH4K94WElY6wvbIjaaWokNqUmg
JiDsqk2IJgZwUtghGkVnk787VEenZmW/MhyhhqBV2TR2kDiVp40P7H0jYtVc1uVldFyijgAedSe+
AmAUrnDP12F0MvSOb3JaKnjBTQtmTItlYBD51XW0cMwWNvgeQlguLtpzE2sEY+g299BzKRy4a/Np
YSD6nCYstIrw8epnbN1Bg8DH+c0xCrXw8qKdLSJvSpJTLaN8K4qWRSRIjyYIP4neQnWd/fDi5WIc
Jr6oLtHmtXQGNr/CkcxKkfKMGzPP/R0dNxlYvhsY6dqLDoSvk7pF4SFxfvpw3P2QHTyWKI6f7fAn
ij+HSMNggNElR/OEcgdoYRALBiZmmwj+Nb2j3SK8C3JfQnAUYgD3ZDMp/7uoGeUNATagit2aVznE
AaJNUkUPHo4cOTfJy+hbBNEz23400qoVsOcfnNIkeN0C2sdjICp/3DVutJPf221k2FKVwXTgEtKS
tvnvBBpE4pWtpf9mWVT7+Qaik0GNkfVWYwSCcGdnOmzdMwumNwuIc1QWeLLfgFej6P8bIaSy+xTx
x5h6MKBj4QrjwGD7i9BioY56RzW/jXqheUlM0v8kZiPv7RKxy14oEcGJfBgB0rBre8QRwoQoXIOz
09l3Sv4H70DRJy4w7f/yh5TSLLw9p+31nLYI0qncqPeirUPWekY+vCvomM2nzGJHzW4RWW3gmxeT
5Hz16cJj4MXx8mKnFXlPChp/8hkGAWqUfM3AT0DSJGThdCpup1UgZ7tV4Bq1X3X7AM3GUUKVorik
Z/0dtLiZ/bV5mZXBPWKhi203GFwkwNvGyy/KQ3/POW9dQf1+EBu7i/4aBFYPC6kP2KPBF88c111o
R3aBEJ3HA0jWI4Czik9JV77eeFHmGaXeJJnaFnT0/BadLcIaqHMxnpTrKbxyee4h7LWLLP1briR9
CDmxPxh238PbXz56r9uwrzzhNPSsEsVa/F+7pUSlhIi5XWrOyaOmAX9ObkXr4QWIMO6cKCBFkjRY
aWnonBPolIohpFmmLGm7YhCTjAUAlPcvfL5c/NSBrnnGDdnLEqByBgt3X+5cub96JjztDVN9ofTc
/edgpWwoeBD8a01+W6fgEEV+M7AdLzfFE+3Fc019PWrTOuJ7eSnW/HMWWpe3Hp71WNID91+li7GJ
YFq5d5huvL39yxtqvmVWBsf0MNwcK8/CeDE3n5pqT9niIp87o2rEHwHRsoX2hl7LRSwmZHh0P3+/
leqNqI86CaleQUt/QEo5i0uuUBfAxOPtnKv4MXQqEeY9WSKMZHLr9cqKt2iD7I1js0/pSj0btMSs
G+M4IVGQj3bMaOpzNdiQkJ+7/Ukya822hCBGssaDTaXQpXg5b6XRtwczRq7MNnFuVxCKfkoWCjR1
AUWH/b6AXSU15htmNguvaVj3a6Ia5JoP+P57VQHxwdkxqIEhXCDWhCSPNbbNl/MDjzc88A8PBDLg
oVBxFWvuZgxjvKzcsbBppZ844WWHNdKV+uv/e6e5xgQVdS9sO9G+HMnoALnYOIZa1wOyHmbwdMDl
U+5XgIKwYC04bkCJVF7pqyYS6wdv6J6ruIzSS8wc9QYdGJW2cS8r4leJNiciKkIn/5zp3c1oj72/
51z3Vckc0tw311ixV77FlDYsN9vXVNQ603c+L4ZGicg/+IB0erB0jxvMgJ4ULEhBqZ02knDnlZ9G
o5+4uSMUM9wR1cAFjYAGTP5SY2gY+0Ax642leC4orUzM2qcM0pYqr1zgm5YEBndvScQl2U3gzI5M
ff2pfqKklnzjhxBZVUXv9QosKnvdzei6Wdgncu4WjTaMdUfnHfSceCnVlGEYlHt84V03/YehhSxN
ZLTKd1GgHT1f4XvzKyyLGnQEOBOh2ixboNsAtuAwQWQ8hBzZfDPej6YiSTrv7EIOJJv107VXotE9
0X6M3FYtCj4VJVURmojHHSmPBbdy+iEKFrE5kNAHLc80tA3LH7S0e5aHP7P4F4RSfZY2iI9k3IUH
Wy4jOLwFAmPYkbAogXTsgLuMLKvhCy3RkPDaT7IBKSJlCVTi3vUgWKM+2ryC//QVP+HP/WMLckrg
uky/RLBphXGV6GbWnHwH7Yz0eTzSTYs7kCP76cCL++gtm12ODcRSWVX5aGqzca3kW1u5KxSIMwYP
6ltYtJIXHGwoPSUGldIrAbnfx6l7c61WwCGZLyK+wjxU6SLqsGGuZPnKskgrA4EbHwJQAWsoPQ8+
jp0a4ms9O2y366SKBETm6XcWOD7+epBJfSNnVPGP+8QmBZvChdk+gZKj4O/Il+Yb6rC0Gy/wgdc/
D9w4WlXPTyXdHXVPR56WgIKEemzbaf4AoOgUgcWiGvwVEIEYXjfzdkMgKuypWy+3M/l5Wc5DimUA
4cQ07X+8o6JPNQ4fpSboHF5jws2yKnq57TMXbX1Zy+Gv7mte1IjxwBWieEITYg2+9XsRtIbiNm1u
8AVpL5JyAVt9Rn/WZXI80fWmFbMartVK4cDC8x+sqPNKIhCn+Ymu2GWbHN07wcwxjU+feJ5zUGSQ
SijMGRUNMvOG+SAAlWHwpazTSbDtGDBQtCsXDAGVV/GIrLCTe9vNKkrfBXLMqPrPkqAbZ/CWrtbw
YG80lkkn4IeuJCg4n5Lit2YWlM1AskLUTKmWFUgsxR2ihrOTd9aEe3mOUsP93h6xPUUfJsX3ymFB
ynNy86kzHA8EmfyIqALouI/Lv/tX7vXSQcWSjw3SYWX5LoGXq+vt6iLPgmq3t1BzUBFQU7RDTUOD
VOXlyZLYqHGcXQVq5Kz56csGI1Wwqcr+1+7JkGlTCbq3dq8vM20om11kMus0uhnQyoUZJcgCLcXh
EyDpc+h7FDzBmE9i1dp4wyOI3JtprGoV/qkBMa3Kf7nqj3MM+dtGF9tdPjOM92/9sbv7DzbaSUR/
QjTNMgodQ3nqHHraRAPiuD/TZ6hQ340IVrBVuhb05d5r0DfdpyUt/XU9/GF+yAn+yb2SNztOyvOI
RX685+ukdYg5ZVyMNRsV8h7flK6vX3M6k+Qdr9GIcxcGVW6jMn9O2BRCP+48QcYGOsm5OZQQe6V7
5qlY3Eechf9bhicWAacg5FEXz72rXOHV7GsL4i/jyB6ESZUX1dKdo/Qff7SHytuKSl4FnmtQgsrP
FktJRwREpV6hBeKZDgkLctldFVEUlu7s16XJGMFMkiNUKFX+R2tLel9w3n4DC8NTt92qz9bzWHnE
0Sv9G5mv/egxjG45AnJ5xVlSXU+nzLpAjkOANiE69NmwLo31gqjj0BJfu46u2vl+Qrhf9+8+8bew
xdhYgHUG5Z9wn9u46kS6ECrdMzflkzTir1emMBdOnMWe9wRDhyLK/w2BlhYEqtRokywJPFQk6S/f
MKF0sFx/PF4gOx2yRE0mIMGrqRwiIpEfpWAZFJf45NxSMYm/cK/Ms0ozE61j29GDKxYJQG2fvaNO
cCwdSunKEjzp+3tl0sDw+rR5aPcsBgWd8f7inF0M85Iy6ZFqPtFLt666LA0LNhs/q87nv2t3JYEx
TDQfGwBPJ6JNGeu7PwQh/GqUDlzH7F2VIzezEEZzwms2cMDsLyCU+w3QgKiXE2XuGOsPa7hI0+bh
EGRqfxOy6puDfkXTA2CkZ1idOxZOrz7DC15B+ttkuzZtZpzuakCNUNgz4umA8FGMma8m8zk0bOqT
p8j0gxNKJYI+nBOk7kJti4VQ8S/TNXkXvWv1zMMNPI4mNEGXajWOX55xtijjT7Zu0NXTq4h5hgQZ
8PyDBmf821hEx2/+Oo1ULVTsr6zpJzrU+w/aMO0cvRdj3a9a87v5E/v+IEeL0aTm/TFqvdUuzlc/
QZ88ioj/ci2lN4SZzk9GZxBgq0pSEaSKSt9ksuoYlJxnT37oO29k8rnPDKOACRAJdUUhvq8wyjUs
N8HGV+i/RBj+gdb03ohUmukVWcw8M2s3iKzK6lniaTMJkyAYkdBlJ1ZhCXf2P0cEBIwQAxsSrRJk
QdGOBoY+AMMD8buQVXsiRe9uDuJKCnVzDEIDd2aqK1d5T8/FiKJAYwxpsuyrtRM6zGCbxtrzvR2v
/2S4sEkKMtj/90s56psWXkU0sVof4deMMnDJyGghgodjEYkvqLRx/GPzKmZtpu64Bj2qkkKO1qtW
4vmcl0eLtR+Uyq4lw1nsFV0BNrHYu+3JaVaIMKqHP1YhDRiHjl4w3i6cHJmcf+CBUsBW/3DkrcLY
ozjAncwMhwb1FVTqS5mbkZV6k3kP1x3RpDQ3eMKvI26bSfScL15YmvZMw+lvFZBfLS6pJGgcfUgj
kyo3XAoMxPyspruGnTPPM3snc5ZXnskliD0faVG39dKn6oSnA3n7gQNacxdChwWAXpZVy6RQ/ICv
jv/rbCbXdHncjtgB0aPhMzDPyuixm57MBksafPgoSECGSSD35tUbPG4FGYuNGT9tbUx5zCcWlegZ
qErf7UrhQ6Ebwd15jfBlo//JoJNwFvMLUdSycJKzukQS9P9cOneqxxINxgaCwNuJcQHG1teogbgD
FgCPpt+w9FVyl4J70ywx9wB3X7lgMgxOtfnn+Td/E4dRfUWNbTXZATgypAZWJyaQmm4W+cZw3pIx
XdyToL+819eLplTj55k2WMtRoekvtz3mJLhg1IfCSI21RUoj/HCPVj9jx8wEv8v3eQmRcWGOn1jU
XBH0nD6kS50rco0aMdQoTOszNy+IQz/gjxEuMYctjc5qzxM+EUEJaTNKOyO+t9sI6f3ns/uW1lOY
UprsxE7KMlUTA7oBznXfWszGMd8ZXnEizE62+6uIKCXxzJxzXRym0a81ALgVN8XvHFJ3OdemVwll
X7Ckgaav7npwMRA7Vszob66cEAdu7jUvHnkfvRfV8T0SOaCQNJ3xoxqIb463ZRGE+o67UeSPuolb
00Ox3smAPT0Y1sfo8BMS4gdB0yJMzskkIvBGe3Xi0Lp2SH9XhakFigc+Z8NJeUN92iEWi9Cq27MM
cJ/HmXdePIlYW3/f8zpJpj4zaV+Br/W1b1iQQqxspMQEN16Uv1OGhNC7p3spRD+YYkfVhdGRVK9P
BqWmUFi6v8dMxdRjboZrKR9qZj4VQiBAgYzR6bdJdEtg5kdHxZIUsBa63Rw6kzZCuq/EEJcfI4Lt
BGBQVHjh1UuN7EPGNoZZDqPhvUoHARseQwfI1G09jwNgVqvxagfpr0hWwb9vwyMRY0K7QS0rWF/X
MjQ4OuuLuRACHyT2NkGyisHG48E9SUpyI/T+k4qRjkG3eCxiqV15sqffbuusoNQ8mQNefWh0gYiP
IM/euxr6770vBgIaMkFg8lXoz9YY4xVYbyFpw90sEnze6KfVudrBNwe43n6t6MaX1HqloLoA+pxt
QGybRY271C7r/ptPUktR8XozXdt0ZDrZTdfdLwuHUgT6dcGchqYqQHII1OTvlSDN4aZWctuInmYK
dOodp1rOAypa6cjOQzj6gWRt79tRORwMtnZXKrzhf5TZQK54bYWEEyQmc/UtqtxtH2hOqCHbj8kE
gt9cwGrEtnBXlZ+M23ONIfBjGR5jEEXvDwOWx/hqF2svvX7t1zQCM38+iv989kAeZxkkXdKQhlFn
QEA5nIRdcLU8sW+Utm7sL40hVVnBgkyx/flbdvGW6LpDr4cGV+p+LCSXoEZsaATmzNYWHDvtl5Jm
F+kZLFs4IMKwnpgGCvZ0CE1tLJ4VBM721V+dX4cPFhRxBpyqxv0IgolokSVVtHNGi5xIkMUcQbgp
Q5TBi7DrDHMTrVeR3KR6G0sjtXsTeBbfqWfYJQ/b8BmiDZjMcgPIm/cwkgbmr74E+pK9PHarXeJy
0WABg4aNlxB/gb7YW7A9eFVgXcN0LollkDVSmOGly35pcRA6ApYwlljhuSuIdk3gh079faanLHJR
xFMqLOYtZWoU72yrDyxfB62gsNm1iQU+JSISW8Dhjrhho5T8A3+/gXyFNKpkSMG34xx+B7BO4A0d
anjC7/kkSRTIvfS3rZhZs/A7iQCrCzlZwvNsZX1yJCJRkIiccDbwbNhhXyubFNSTAmqg/JPRrNyJ
amq4LpkTwa5tFfPVFHcxH+i5AztiMKRr4+V4P/f+c2117Vo+INBNTW7MHbojVHVFsDrnFRo86Pgh
xuwBe3+wcUekLbEpoN3FjHe5QlXRzq8KlhQ9dhc02e+KwcABsjigKywCr0CB01Z1+5AcRZYzggrs
sYXISxXC/izK4eBHsghUblmVA9bWHqt8V8s40HeEQAGDzk5fsUMgmF9eaaSSGC9mIxmob5hyxyN8
oXsy7ib1EGNOd3hnFxQr9L33Exlag/Q7cQv38cWWjoDISZTm9InAOfs/ddqJ9hWjc6gdJv4C2YZ+
644/TD8iJj4ozfG4zxyIki45TrtdgoZDisS/wdlCHAfBc0fYE83jryNrVqxs+aHUhOlCQhI6pOEe
znsYuC61d7ybd0sRyXS57pvHLW6tRf/4Ymqtsp9eDEy5zFla66D6Ncdh9EqDl29LLLUsyQua6n6e
+4F+PfCZEjsrv8wyu2arPSk59IOpgGtoEZZ2WNCEQQXrk3tTOTZSqLKSMW/weea84mjhTlP/d80W
FUdHrd7So7a7Va3EWRNnR78ToCm/nUxYugpj+hSpz6ddPOW5XUgfQsfbsia4rwYWR0TBvO9qhQC2
+QIb63FRcAUoRNAtza5dbegGEvi46DYBiw0vpaFolAJ9Qus8OG/9FTKWbNNFEIbCw29G2TrmyfSP
X7fGpe906+lDD0tal0rNAhj75ZN+v9do82NAzaAMCANTPexfMCyoCV11hkcQe2z7D/WwDlT1uzg5
aHYQ9bnO9aMO7rD8mmi3rkSoVz8S+MxEp7QFr58hofIX0gk3AF4Ygjlt2m+ilcGOqUpLPqT7NIB4
8FVTsyrE6K7HWK8vvp+3QVOv27cavknytSWOqsmvRaxMpJygTnNlcLIsWibwQZA1CyzUg0bzX0ZO
bGjbr1J3Z4qDzRdp9gOg6WyqlzkSBcQSOv8B9iq9/ScQib+2YkxMKeH7w9wcazMudMbdbajZVjIU
sSlP/D9HUJT99NC5swQO1fbZrF5PGHb3o4drd1tRyo2N5SXeqL3UdjVUmpZ+Bv0wImmOHFODRqyo
gk4ZskeRLWISPPBKOQnglvywV/rYaBEPkuYj6bEHzEcnGUrF9l2g9H4FczZ3qA0+Mlleo75jb8LE
j3AuRgt/NliRIW+Oy1nbmngCMkebyDEC8J7nYjmMVbDyhGY5cduEgPAraXSnPl6qaVF5gUHiXbrT
bgn9Cz9oKQjHaJav3EPbqnG1dKY/gq01NEsTYb/2Ya9W/u4pEW7ciiR5tJhKyu5GcSpaZPPpIoRD
ohtXR0thkG4Ps1hgcYtutOppHKsLbQ6nFW7E453Z02vTxaGzQyN6H3KPGgZq4diUCJjGY7WGRdG5
Y7jemqfe1m5bAzmYlkdgmet1B+BYSpTKwSSCo/CmT/SeLSjG06RARDHE6X7CDDU1kmaUGKbBsQNM
JZoRx5nZeItuPy/FutN34Jz5zGQ3fIB9kcQXjEGbFZk5PWE8A57pTPaWFSOGUo2yXj/bCZoKXl6T
fwwLpNZBFq6ad2JoKk9y0MYj4d1R5DUF3NU9iWZxHK9xJqN31dD5fIwl/VbLIr6bhiP1y5vZ5v3D
gyXznK5VIPuq49nw+2luQ8U36fQKp8ocHNPKngkkUc8mzjjxgNrcQH1EZgO22KjDWs+RlBaH+W3w
T6bp1TLgkq39eINPoaqkQ+hDTc426+JjLZzRov/lhIDpxqxqaSji2ZhlNPVcL8EUUPmnwCPoC5RH
a57z7wsO6nFHeDLCRPkhmDNkN/R15HhMPRkl3PJY+m4S0Rb7IbOvN77EitojdcCq1i2v2qYZ6k2s
r6CWU5HhLCE4Gr4aGJrA0F2I+Nn6OWWaqzm9Ejqbu/8Isn8zoVmT8evt5O7u21skXn7pWz6HUEYd
ZbwaJ0cnxbBvCiFOGpjMwhpUoFoqwbqM4tNpYKN4kAq9L8uP8yvSNh8SNOT4H/68ihS8rsmKE5SB
pfXCA5StXm7Bh+2egz5vDSuVEBbyYnbAHp8Zg3pDn3k2zE98C6rda4Vz4ohByCrkYQqYUsOgS5M4
DqodUVtLu3wdpHwHhxZ72FEJ3MtGPab0dUc88DPQuqjJcd+NFKl/EhRM3hJmJCWEQiGaFW4Fn1y7
t/yLg+Df3Q86po7CM7VqMiP4/ZLTsIKKzBMHd7WxJLkyI2uDiHTHtgwXAFcILphHl3VhJH8FXQhE
Sc22af3A9BhNNg28TX7kh0MEzF+Xn6ooofJE5SKK7tPukvDMFswSQpoUByiFYCDvNRZEpxUAxG+O
Pr+GhoW3IVuqm95OLHtheGgITYc21LEowqXfY83Lv6IOYydUkq/p7lwHtQfLQHoFnpnOR3fdEOWx
/Ccl6CjbuUCBGdshsB0g9wi2kfjH77mRztK0/VJ8hRVn6Y7v8wsXol49khryqH2/+5KwvP8agxPH
ZIJKfp716DwNddO7cwhHNrTRODkelcrBjo5lPHH3MpV2/UT6sz/7mps/jsBeu64oCkTWOa/2uZmi
y/clcfezwPgY+Tv7If7C/pDp1lHalvyJK1B9GCCGLEwe9gOvTXdGnEQncjLBOUZ4rAb5BG0cIjML
o1qRtpVGimSrzxCiG+sb02yLeN1mUM7Nu/jBmhNNGOtRsF0lSJyzXNuPJoSl9BCh9MG5lOQTF6zF
BzTyDSxW5RutC7tnO6f7EACBcprlC6XfQsOCIlAL9rFQIj8KPQWveBO1S5GWRRqI63pP0+uI0Ov8
LTByH57laZaPxMq9qYqNMjgaijj7nGJ0x0m8uJD6CjaT6jnJM//YzXyDeQ6HdV7uazlVyqzVrel0
m0T65eiSZd9vdep7y5XrjW4/lu0tfyX9XHxSX5gBdkCUaES9woChO2fWzXYxF8JctKkIcvWh3iup
St1JRe+PmzfUUBFdu47Gr3VPkqWxXJOMX+gcU+WuaGB+nZOal3RiFID937Z3YMlBsW0P+WCEGr/i
hHArYhgc+Cg06SiVYTDCUagp/34q8xIURl21p0zeRs1nkqayclCVlZNp0bY9YA4upBtyanxj/kXh
3dkx2wAe/iJ4jKnWzvdifftnv6bb72MXti102bqg8tMkPgSY2h6yPzCAZ8AHczZo1mweCGlYcaFm
EKArvi90565yJbi0h3knlXg+vzq3/RFJjhanfecLYP269ztuLRI2ffNXpeRtg4AXx6HwEpnrMstG
gnuIramOM8iP5reOw1RiM4UgB0xXgbwHE4n8+nPzMuvco/kL6dnHBSdym211BM12usp8Zhc5MiG4
ji4lw3w8shv/b97IMaI5c9h6sDF/5XZdEm9hAZyPk2YC8VtOLd0+70HWOyPvxyYVbbHW1MBzZHxm
0A9m9JaSGk6ae4lYDtFQPBks/ejjgVxKrCfW7+L8RRlnt6YnIxeM0DY4/cejESvWjyzUzdg56KrN
2QLiX8vEkhI70CqylUiyJK/uE+U9O9U8JV9nzbIj2wUTo7+z7hzTBFI9wMFYmp0iqFkhq1JRsiHs
aXD+TSBP68+Nmlp6U1fPzu33swFxOiiU7UxdnuXI57vaedWbqbQukmiwyCDKOtyKPjyDTRupTyPF
TdAzjnouEZTGhmuWhb5gXqSzYwYO473PT49gQVEPXzX2cc0cVPoWVJRYeaN+AkjVRlHV10wLiQ5h
WfPg3shdulbIvSAkID33GbIS/9xrL84C3JzEEoUT1dc8b9jCni00NpgMym2rxDpMqPbKy8uzHe9o
K50zfSM/3953Dl1dT9nyw8Bgs7gEDUGhKGe3B/meLiG7ZJoD04SQzs4+54+jejAmrl9NBXYxwv0k
FfXs70qH0SDbLRWKmLft5x1maBM3EDK1maPSksvxtY5xKhAsv3y49LaS9k7jhdZHa+VlMya3R6tb
LH2UzlzzOYidY442JgLHBNhsjgrlvvtb1VOwFrtMLo7DDL3H/i+z5mPFug8+OK5O4Vy6lYFN/NG9
ilRYfvWgmiMSvDKYtSiJK8xMKNKEx6YK7pLDQN/Yvn4vMlWI4WxN4YBxtbRut/1IFn+hsf2bzwjw
/0sdDd4htn8IYNuCAMhsHu+WO0cQdFavr1CRIv15yCSuemQP0hKDnQ0tqINVXHSjgRf2QVPwma18
eJzGGYTGTcHVMbbieE1PVfoJB/1IrzXB5Z8RGayOk+TDD+O6jsbwbSJUeq8bBpzNSKmzDqkwhS7G
cBorhnuDg36bDmb9gTd70bxm+/0PuAvBKEsCkpe3Cqz/1T+Ig80uB7tx6Y2a2lRK0rwmoZNGRBBQ
VV60RWNGxpF3glvFTDo4kcfmCyGEhAgFu8RTC8x8wXToReYj096mxrS2+clledEwPIX7mYQugHbt
4xMfk5zErjCqdy020CZ275FSJwYq8NQ71FG7XEbaTYAp6dldO30nJjKBEToxrc+Nuzy7Ci81RTxW
+KuygHpE/19L9DMAugPyz7KVVfmsYTZnlfxItb/KWmV9Epw8JfibI4zokHrgxJIhPmzNwwdZUlK/
sHWShw2LnZIBxHIPMouuS3vinmYTGPTcHcoPqEBr21SsnQCnWUL00rDWKR+yxUWSwja6R3mPuNRR
iYO4Fcp3STTKo2jvildVQInnaOA7JFIfs4g0HY9mtSknrzM7fG5KKqUXvMnPm77eTpKOlC7UaGHo
1NB0++E3FuRNxuqqbFhqk9c94gOEkvPhv6JEzI6lzqBXuYMzNFgPqHhrfoxi2PntU1kVfGjJTk91
oMuS0mEGPbeIEs20F1ZI+sGnFlF/vLImY0shMWMR4PcZ9FuC/9KiNM6bE7HeIwLwCGD1tXnLm8z/
yYcxAA9dOQ2loXAR0jvtFBNWeYAm+7UG+Ijwk3LDEdJCeYkHAx/PAVaw3sewDYJrvYwo7GoACbIZ
U0ykV0Wi4IlMrrEEkgLTrxAt4xt5VU1E2UJ8O9aXEnTep7pUS5fiUwpJ/t51f66nYXGObSL8e8q6
eAtvLWBRtwGuSTLwsgIPvrBSWcTEXbIuarFOUpK4SftIOQ1P3m5lrbD7vN0xI0wZKgXHKldC9Q9a
IHtPVJ7IP4TY60OnjRpdOW//jc/6JQjzkeimk6vZneuV9ezY3jXIffue0SbRG8hgyZtuS5ecUf1V
krhpugDcM18EQ7wo4TyFDnQmFC+hgwSyyF4BrmHi68jsxZUGuuPN/KsCeLNeAS4lCUA33ZAbBq+2
Hd0pyiyWOyU0cESLGyJeX6kA+hm6WRB7s4uEcXq13O9gb62hmotPtbLNMEP/40dulvDbDlWk41h4
bcRf5/Z7HsgVTFVen3u63rCvxKOG9F25GXlRJlwaVzh5iujp9e5MIxV8uc98hGwZfKNlkk8KSHtt
0YItC+eesXN4f+L3jF3V5C4gKjW/nOZtWq+XuEiMj12UyWdS7iCWyB/3Vn1/XGzb6/9JnZDUDwIE
00EA9QGBj2AdD6T6QmRzZOYSEbp1LqUKqHGHRSZh+7qq+uFAyppXfWH6rZmo39m4cpGsbUaeWhEA
QAIvawak2KIYrGz8QqU5nTg2iRv+kmAN/fPQCSaURZBg2A22NV/cLiqnu1kgYcVvyfONn2hK6GER
Qh8IzVP5Jyr1WWjw9Kz29C/SnP6LfNlJupDt208eXjdOgji1JryPKKgeaTrQZB4xy2t8WErt7rV+
Js5PH4eD4Whe6LNlfz1wzS/QA2tQ2PJwtpm5gbjWJayBEz1gT3r89i1UaJBzWrkmjXnPlFHN6AxK
CEo5wd0qRmd9VzpCA7jPA2511dCypFZ357X/ny7hZMKpVwU2ikv5xP0rNLb/iH2eP9KNNu26VGbK
cEJ77s73mnzfgrdRpRqnSuXnidHFZwkpO9ta2w8dX2aEdE/da6ZmxNMownz9yBvL6q/PpqIPW/M4
vKjDgbJLBtyo4T5hgZ29Gmv5B6cYyqtNwVIjjXdq3/hfQxRNerFUTjMezCv7Ucx+PhZKnwr9O4M9
HmwpInkpj+hskRdXBicKz0ajaaeeplUquR+zuaIeWdLPaOAaeRBH7NJ4dU8Q0PLsvnZsAw7btP46
Nfc2FVhaoFST+JfQn3qVnAMT8iuZXElNBBKmMshWkkM7p4I5uPaupa411tZyT/Qd2gbDkWqf9h2a
2tAuXA4Hy3RqqAKB/TW2fpTNEAqHSgY6M+f7/I6SEGenBZ6amVRpbB4tdcF3z825uJeZBvfaRsvy
gFD2U7ub6n7PMtPCQ3lzX9QfFQ06P3wBACcQ/nnXxyfCLGVtQ8q1RxBRWh95oHv7kb1EBHzOXe3R
cscZcBxOHQylhmDdBUWysmLxQs3zsIKP6Sy8i1XjiKcM2JA0w6ab2ZjWAzixDP4I4m8T7ZYmim1D
Go+XbTfkwTz8MVhWjbpAAvmLx4/AYweA9bhcPMW9i4tXL5d/pnXDcv6LDggpIwm9s9Lphhm+6D5N
Bz9FITrZZPCAVlHiYeL2gLxbsVCpIQSvax8wawnxYTOj6s6BNVQVuUxAQrnfZNx2ddZ2FdR82W70
yhWvibaXR4tV2WupMWSxSvCqNLdLujFF34DKASUUoLqPcVyVMvmgZ0kXkYssY6p5YZZbp5/tgxxR
yNT0HTh9jpLcoGLGPpdrl+CqzVhtKJhD/6L0X0IHUbjvpodLg70okdXnoYfm93SpfcOVTNGlK5qA
w6vMtMsshyQSLbvBfV2+a7K2gzaPHArvMMXgFNfER4/sHuVDU/chlUkWKK60D7itQPiPsv+kRsfa
5C0pih/6Q96+XSIGrsQu1jGZx2/ulb3fCuimxyREmiTo+GFSGJStEV/6jKWFqpGmKfpulK/7OjWu
eeHmJQ441wna7Iw+8WXSEFY9gtI+FcGOxqmagPTzc+cK74M9Rui/HmZMTc2Xu090tZfQENmWrAJI
qpzHM2aIbebYyCP7G8Rt7Lu410pdmTJv0vPbkp0PUscP00kh9zflpouTEDLybPatR3B74mXQJCkf
nd6X9vBEKjKfJl6PdXtpE8wtZ6r/vFG8sINmwwP7n0AO4BSeYqlH/PqnYlwg4YdIHu4yHkppzUOU
pLfr21A/bapqmprT3AVgO9SH+ajkT6GX04aW5bOt6VUJ6yeB7soI628RSMKeP2DBf60fUP45FFsy
aFLMp9QQ76H1yG0HV43p9HFOsMcwNE/9j5tcO+y362wjR4lLnchsakZ68RpxUG/+5h9AacTTPxnC
o872OUbjiXyK1fCCmZlu+9wF0hHXAa/DhmqvgmAgK6eqOLWz2cvTLZXsk5WMsTMY91Ztnmjx3+Xw
9f02x43mQyerN56euEo/5drrdOMs+f7brSM5/jexWoqChi96GPMoIxQHDtmCwr1FSbd2o1Y16s42
9DQyVtn/mb0gObIfmxmImbLnYZQRhzQq8MGdDFyNi2PN9GGEe2A3Az3RyPunHAXuG+40XLpUaP5X
eKB82Y6KLlxUn6AhtN9O/uZRHIxGUVrgpbxGGkgl32L4OPncrYDjdTKLmpMFNwYe1ON6CX1OvC+3
AgBdcIIPgyM5sbNpiOMr49OAVsnmPyR9sUuLGbqPTi7mG6PBofOUCJ9GthNl0aN2Dn6k+a4wvlzJ
OVn84Bv3I9QCGyKc3/w6lNuWGwDtjTLB1P7KPm1+0XqU7z7uVPfYr1F5+giP1PnQKbaIc9gIdggu
mObPSR5DRSXj4ew/08TWjC+7M16sugcSX4fOsQuJ0t5bvvN0E+8Pym1qvMoiZcyhPRRvs/aov1L/
HP2fxHGFCq/MYk1dDBo+xko2DhG/NoscFJ5BEKBYl5vuQwc8CN6WWlN14qJmSKO6zTdtIgAwYiFb
v4mfS019dW/UItw3UetBq9xX+ZBybUWAIfKhw9X5HptPQPKDEBO7lYc2L6t7Qaq3WUfO2C8nQ9hP
OQlsj2s/JBx/XEikhKo2eQwycusMWlnO1c6j7otPUwc67uiVIBlMZ3afYUmBAwMUtlZliYBZWWED
ysal14tawMu8f4oF5Z7lPadYJl39hxIRz7P6zMf6xn/vIl+TgNuORuUy4UliUtRjWQxsbfKGQG5r
RQNrHa8y871umbVKI8+9y1JkMsfIlZIWJI88I8y5lnOugjbV6taAUvdEttUSRsKI52RzrCP2dNVn
Hqc6U0VVs1LyZ1mmqUmeOBPrPooQ3nzEdUeo94Z4GNUvngv70gZRE5OBCT0KLMPdIDNoUlJD5V59
VhQlrIwpJ7zipBpUyCnfhTmzejIpaWWxvZKVj4TyYvdujxUcvQ/mmgCBh9JDDGE7ypkfaP7rYdF6
5Nb2NKZ3v9E2mFGI4PLobJQgCtYyDxi1xJe0aQmWWS71tLrfXmOlQNPG+zdmWfdgURoGT0kXbk24
pYEyvPyDCtEL1oFao3AT4+WDcR2UV7FpFSDnzd9vi6kFsxoeVUAe8dj9LAgMo0XoS9AVzAFxzftR
2GlwjwduV49G/XLvMsrxgfd7tFMtLry5PUpnGu+9JwxAIXLIMzu3gSw5FMHbc3N7NwzZ6PoU4+8i
jkXx9+VsstlHTRJmFy86pzwcIVbSBSKda09vvdBJye+Cisu9iyuIz6Mtbh+yc0dhK48WP6T0aJ8x
z+Je2PLSv/sU62eRfxJMQmvcVKc/Gxr8/XnxLdZ1HtGWInhTMYvFG4BTYPDfeCweWzCfA59loDZV
AXA0fyNGMBR8JABtkRKPjbRZbYuc33m6UNipzoSt9CSQE8BdQn49ofTIO9nc0ONspVxCve7RJgbW
sCpypFg+uYPW2nm8nS7nY4Uy+/XBBjgciIokNieDngAtokxvWLvddYtIhM7bMhRC1jW8shPK8if4
2CAUyaZJqKMbXndypVkbt7zaUdabQm5INhfz69QbalhRzD9LNO6YKT0gFXTcmimIUUBdwfUjaxDC
log8L1zHoZ3zelOYzxGM2zLuxtZ2IdH6EAtbQgDBRH54w0uqCuY4lo/ndjR2pZUDm6krdazfQ6aE
ZU2RcFvUdJxqNwDBmviUWoymqzMg2UMvZ7t/oUzZJC4nX22lVOmunstjJuWT7Kb/KQ4IgME1NWPS
4Q2w0C8IS1l65HHJVeAegANXMRpnmGI8koU69CiKmnTvEkmvyHAcRFYMOyGXa7HC9LXo1cYSyiRg
CrBlRC46TSRkbJ6csUYoU+GSB+CyJ6bUBSGPf6wjwNdwyg49oG67rZ5HLKE8eoSfPoyDavt0tt1C
ly+nDdVj4XTPEKiZbZaraQNEkzcUdXYv5wPU1oFOtkemfv6UaXHCYAV2jsvBxidtttyxtbH6ODqK
JpWbDuJKE89lGBGqPbt2l1yjN2K3EPX4RqoKqMI56dEF17KaGFOBbhQQ8nj4+RJ6sZSEa/YoZmR2
IwBA1HQRGyh8n1ig7Yfni/VW+QrvteVP7wVg7zIorrBEMaMO6nOLCRfQnwPnK0ePbFCCZivzfHO5
aMNVMLy4DxFUScB/e8mDgmfnjEbrgPs+Q+EmlnOpx/EwyUBK66RWg3lnCwSEjOstQCNt+znrA6H6
p291eLbdNql6gnpCVGAt3M0jINrZcDT2UPOgjodCPfwAMtpkCUjCtYGPDRzJXzrdgVqkVZ5hnXZh
fxb97RKQ6qnf1O8y/tSivpLLR1yW3wN080ftMijgrM8Lgnhg1ZNAGAE0Z8gLeyzuCDciCNLgnvY0
dNDOKcKK8N7tJswWprcYc8FCaaX6cxGYf32PedhfVBEp8HDBVJf/0uSidcvWrGLtsqyuii4YhMbC
FVnUCZcWBT5SvcLpZ0MnlY6nVjXbJLZfjMx9U48Y/V0K+8vH23eVdN4yoNvNzy5E4v6pbTuT7nGu
cXvqmwFRi4F4D/gxrn6pRgGoxhiI1veyapTMYiKKNDdIMRyxZJa21ruZB8FNHVnaQ+FjxM3bQiWy
5eEBvhOKWroyklIWbmME8PcS+i9FGjzW2DYTi7LPpLU82wHz6HFmpy8DGha/pXeq/svZ84CUa8NR
zgwntavuoRETSSWKLRk8vrsuxAgp41iHaBR+18K+rj104RQUioafnGJitAjt5nO2guR+DkHLnwFp
bmYd5qRPaLI67lTjRCVBHYV0IyYw0rNooo0JCDja1eCP6zly4lM3CSY5SXYXTUd81EMTgJKn/NNl
nCv/gfrXIFG1In35WMI+ZiqITM27UZfdmcnISgPtr76MfRu1EnW8o27Tvy4Pz5sjYGqShD+EI71B
NtgYINDKJj5VfBHlPJ7GfZ1L5NOmoGBUxcwh87mTejJTuqKYWPrWPeJ7AV/aMs2oT3FKgSSxoQbc
nQL2GcfyC8seZD4GPbz4M7geY7fRnSpGJACY0ryo7IHeZCowaElHUZIObpk9d8CzMcrtjJxkjiPQ
FBGnoHpgVQkxl1dO1IcMYkJ1BeltIZcF5iEvV3aCHuhrM8tbto9MeOqwdst1/ABIkyF2rQM7KceF
5TVWUQy+Vli3tlm26+G1h36/LeuXmmHoKe5yz52DeukSWtNvJsu/6UtW6Wh4FhXOroNgrX85lCQZ
+yVyknVI02fP2wcMi2/EfhyiOLoJqEXB/42ha9DjZTKjGj7XBA96WwmNFYlTgKgE8605QsqimXq7
MlQEy4xJuj4NBXN3CpK4HSXyJFaRwC44FCa6zh6qV/QJ/VTLxWfemUKbtKgFr0h4jdvRGCOcnp4a
/76cImCuxwwT1qtqWNLw1UaGuQHq9ln88em8OfMOJNmDFXG4WN88e2EZcT83Krj7SLTvF9THinip
s1hpwBZwEmwFU5r32n6Tm6EsjJU0iEkl5BFiU0QTzMBnu34eRTB8dYHEmVdh67IUxUNVxpVic2MU
LS1um/BBupJLpwRVJO4R9+oapIptWHIvZBI0TyOa82R1+0Ym9zO2P61N4NDkstXNvQHSR4QsbuNV
g13Ib9Cb4bdebbPln3VLOziDs+Yuj2C6vF90gDR8kQF/AWo+3nXkLBzHc5IQzhfvt/QZgaNJAtWa
y2YioZAyqJlHl9Wp+m4Ek80OoXZeZsA1Kv/eclTJDwsFwcxbp86EJ0/Z8Lf4winKTA5Fv6ES2DUJ
uoU0OAKMIef51ZphkD1cXq7L+5txiXEg/vplSBJGxvjdIuSc1x0fGBLhLrSqT599NDxm1iod77Cb
ktaOh092d9oKzDEXTG2LZZLy7WZdyuxmLkfpg73AC2nse/SRIos21shDmbWfd0NGgchdl9okzHpZ
2lBBAGGBMXVITzxYGonsbMbVYu3YIjEAgF3BTpgr7y3xK63rP2whxssu9TLsIPWnwc8pzdaICNO+
YfKuEOmZGR9LXOOpHwtIPIt86EOm+7db+S058IQh0S5VeORdj9ra/hNy15MBMlmaVADjV8tl11D1
m3jNx/j/z8EoMizc8gADunou6L7F/Gdce/cfxLOXI7/PiFUD2/zkkDL09E+1XwbuHrDs2ERxdTOj
scCcJOZr5zZEfVilugrJmJezwig512/hKf7F6Cl/VvXeTcz/eL1KWYPgjb6m3XSXUrQInXUhnhj+
nQbvkO4Bp/gUSPpNjei2Ms7n4LHfDxLIFLy/YoBe/03q13T5ruycehiYdvW33Ja/XrX4Zj37RoAY
zch+b3tu9SPjTflRXQ0xiYvoubFBBErmRivRIuVZN1CUb7YpJD1Zn4GB45gDT/U1PIrDOkhKq0u5
9UpR0bFuw0/V0Zn1fVGku1tebprKGV/RmzPyVUMS44xUTaZEmrX4Z/IRObOK1beeRP3QembB5SfF
AzW+GFkoiVAdjyEuTMPxSMoOO+ofPJBNj0iNNqbQfnqjvyL58l+aRC9s3Gyu81A7SfZDTqn1Tbv2
LxFa4gAB+fNCidSS0R230TCL38NPUAyDPa9bEDBIUvSB2I1wDnjBKYdGqHhG2us6ZTZ47vKvNf04
1SusQCRnC0acM3L/IbJ0ccB/zK3iKsdmL6Or18Mf3EXWRpp0uKB66d7C4ZYz5uN/ffBtQD4M4l64
zRzftKBroAxtVCdbn3dG1J9GTt+QY82GcAjbBcJclYHyb8lmBDfHI/TR1Ud5PZyEzDSMvkrGJypE
gaZgEqu5fYjKHhLioXUl3jgZwWwgGvQAuCD0mHW2WoPDax+VanfWZ8kF9n34Clw3ttF6T+C96Ijg
6HalhjT6Nlr8orz3F/bhMIcx5ELfb+W+yFwjlUlpNEdzUUqj2Na0EqxOH/6ksdX6elc6eD+ejF19
kekiD/DOEIWvgNO1pEBVg4MYF25tUPLwXK0cmkVNMS8UENOSJz1I4sYq8jrJNUGT1BtBeQHNoj0h
lfh4LcRPeLU/E1ScKoSJmW9a12kboOOc4gH74Ie9kyTDF3rPkczx0MCy9YLXbhkzsi43T3+aUYEI
adva9iHXmCDvIuwTtP4f84KWBMG+Iu4DFFQs6RVoHJtFUuDc4J2ZPf1aa3shfTg6DQTKppFjn4/S
62Ar/GPnel1zNxguh4xnKBGTLQnJ0LVR/Q1f9xZ/NYtQ9lKRGYWnh0sjqGqQie0nKa87pQ2kdxIz
6yAg9WN4RjXE0XLOeizarhk4EzjcC6vk1Hacs2lj8tte76zDqabm1YGv+J2jEfv67TxVRo2BGSkS
oHewIhaQUXUzjHhazG+MdVrBlEaGOBOaVrNZB/vNTXdyvOzE+8L/o6gblJGvOruFjAlqVQxaeIUb
LehcoaWYCWBIeZqg8xOPCs8pQQCmzQgBisk9jZWl8JhGeSU2UTJ6rDqqoxIkhWqdope1+NuObXzc
fmX96O7hsIrfMs80DnpWAY3QQ3uigyKuT0aZV+lu0/28n0Ib+T8UkDXNbJRM8GVKlY26olZqrJIr
TNiAGNKIDcVXV9uJJCHQ57LefijuN9OsBvqbfFxDCnHc8LZMp4GmsAOac91sP0DweTP3PZxKutA+
b/91CdYltVAXmBF8vzgom5lhJ1xOYQXrBY4mf7avxrZrptd33BlDuDuEa3ab4M66hbuuO7pPnETE
utbKwAlEmX6VPwp3WewlBHOFaEJFTgAG92vNzZ4rnSvP46IHixC0DfwSaxjc2cQrtDgeUHaqG+8Z
wOYGnO5vMH+1/yE9Tq8AT8+tqL2yjm5ub0J+xq1uBlij5lZHMWz2uQt0BPcMVHBhR7kcPjUPL7V8
9LSkjS36knr4izOBiJYKlZD8kZbHLkW3VDlOpwPypIvVLsnu2WA2c78mHX3XWdI7tcGWGj+YNqeX
/O+khw+UZC5O9vEa76zBQXJtIiiTuANII1FByVDdkHJp079DfUvE5hFqZYLpQENPlGx/jZ50fjsI
Fco2qO9trpR5seeNTRQIustfpDh1p38rB2dN3ybcznnIERUQOWhfi/ZhxzKLGkFkzlJfDtyCokqX
JYJsITAwmFsHSMF4eeg+YvaLBomQhhuuJdpsTL9Q/Au5HWEGXncfN5xgITCjDHMyFBZF8Gyp8t8u
EbK9zMrYGVRfkUzdOc/ZQlMyliPx4tfBaFj00rdl2k7jbAFIpaOUQRPFd0pN83/6Gkg/ELCPKyxx
mR5A9jz5yTWvQ6Y7Ho47FTzPp3wyW5xohZlXD4ytK7qIVFzcQSgsccclHOr5x66DgWwRXOVt+g9c
j5txpTdxMlBD+FyxtTcNEw43NUxntQAogM8G0b8g23r0ECFfTZvdmiwU/hjChF6TXIGvOzTZS5Vg
k5VXywFHBKKHerVQ20NMhrxzIsRt02I/T28M/gXXrt5YbqFTVbz8BmbAOhOdgw+p2bSpUJIg7VW9
KV1qXklmrEMdLwryXRH0iHlTqFcd/h0d74g8LKoPI9v6XZdq96XIGGS4E7LrVJPkKYrynzQC2XaL
G2RPtaK2znW/oO8QLC7U+55J3Qv3FM0pa+1+wKjwjTc6FVyYh2slEbTKziQFujfIszfViFWrBWC5
7cxVPU4bC5OW5pCVSyGo7Mb5TWTL+sSWzRPvk6rA5xGi6lJmXPxWCBhqZOJXnSpGX/Wu3sHHs2JG
IWWuYQqRs9Vb0WRKIGWfm3GK5FR9hxBvD4HFoIKGV4GKljB/7KVMFrPYVt5Lps4CCqziuoSHShf4
kk0FgwO2gmSCXpn6bTVn3MSvgJSNJRDN4/rs7vZaR4VhJUXSzDvTWwkFjnGUG9wLjYvWVJunIwXX
KTNdTIl6/e03PIIDuIcABIb88bgOvzTeafq/Y/SAuMeNzzKJfoWBpyvUNtUgOeTsahTQZojaBzXW
2CDzgo+TRAV5rGQL67eQqIx1o2i37zEuq+goCK4i51GErQSfTrF8RZp7vCUE2e2Kf6RqNebwy7Tr
Bvv5Nk3riWbosCdzufwQHAtfsyfR4ZcP+Q6sZZBq/2qhWvMMH7Ev51uDJohK6pr92tDb4aevq6Pa
r+D/FZ+dSoNKwqQOHgno3Mi+tanI7azSK+xi9FZ5SfRz4LeZ79mjoBxxScj06CVR8uZt5/eeRaJJ
hS2gjCJgQ35/99eta6xyuGBt8TdoDlKiDu2rf+cKzgAJjNm6eAbRGANQk0SE/8qrZ2p2fwIUVmqZ
N2fSHi6sdgVsz9M9Yb5IZBaHgvgqtGuFP5pzOqySMPkNlVHJR1UnXm8+rv47KPNkDoLBZKdhr4Bm
IrJY2aHp7WUA9dKmt9+CE8nEEZpCv3f7Bu3dl0fFiJJaqA/H54bdG4qhZkxAWARD/PPcOaf8YaQI
8f5iIYvlDVKhcUcMEHfUyudgGyuHVpEG36Zyf19NeTzmfJqgisV1A6KxBUX84VD9TPmcQANthW+l
f9J6w4XPVRylGdRKn/vrvz0p0zAuwpV3mwAFrUAGBEYUG1AXhzZb0pgrvlw/8wCa5WXfRbSJN/TM
OTGy180gXqlzCxaYEXPzDQSALCIkkvZqbU3cEgLB/NmhPPrc7aF6PGUuPFcA1OX6gNvmqxULzWaj
5Zk+VGCMIAGOpgKKy/GidHYoo6RQVtNooG3CrT2TQ/MiAigGI0L0g8QlaU+PydSODwaoTBCkxFZM
s61GyUhn7/5HdO9X+q4CC8yxWQCSu04l8JbiJ9a9YyST4dRW0Jr0pNxVvn4pOBgXBd1NWJnVVPAq
BnyXC4aXu0rI/Nrb/vMHTOMOE73QbUibO+OD3tvc8fZ7ZzUJ8rgWrgIJCqduYqnvXNTH+BoPTzfm
smgVc71gz9pxIRBfS3IuHvxE4FjHCvvXRupRls5Gh1Aqn1a0kHE/lG0jmELXdS5ET41YQLRge4To
t+KdkQteX1gUXUOuKK8XMKnGADbJ8U7GxqxI2Fm8U4NWrFBKfFLM47vkaot6L78zrgrPqHh6422w
+U7dhw+/S+lOqn1yDXDqDcagPGuM/v9guFwx2HhNilz3VjP4DddMD1J67inv9bnva8N8Xk9IHVFV
WhJAuxbgcQu1cy3TgbTJfSBO6VyXM9gvIl9uALaWhnCgMQZ3Z1o5XRpLz/N0Kx2sLJX2ivDkLTq4
AX3tLKWg2sxTkc/gzM81+qJHmAv80iKULA3cjvUWAYHBdfBscYi08DKXWGYNq9hC3DUszQDxo9dg
jpjShnYBxw2TxnoYOaS1rzjcD8TTf9fmd+HTuohzxtXJjVINbi9r8KxMfqvJXt3rStVuHFQmwJy1
WPs/uDQKw1GwDPAC43jm6T+sZDfLBVpmhGfoyhz57LEgrQUeQkMUMPMbTlLWaAkyySaaHjDuUTa4
VnAchyOZoVugldWchtDGEQjISzDkFNt13NYj8pYSpMd0Wz2PwpzIQD/NQ8jj404XN9NaDGeUcEDC
6rK0dwQGVP98PMIr5F4u5x+kR6JZIDvpuZ0m9mrQ1He/Fbixh+TEM7i3eP4KCO3TA03qF4+1emgz
vPdJgcwLAXCbGJwDEmtBcLnRbv95dPutjjaihCpKhAxwWcZwq9qk3FRPmg9MaS0gIUM5QTiLY2xS
6eusaxp3bxV0/FFkp8orAo0AJ12B775GLvnGpo4rpce4tL2Hc/A5bpIsIXA0rYs7a/3zdTr6RFPG
AH+rBQxZu2IMDRhc3QNPBPM1k9NW9u8WGgZJvHJFWcl2/5bp3wlrUDoNVLwzw8zv2DBMyKOsMRtr
/F1rH1sKkO2WdobgjOQImsELRZlQ/Usf3U15ccCJRCoVg5ZB0Q7EWMWMiukzqiAf3FKDUw7QSKzT
TyHedzuoKuRjtJBJ3VShyG4fwJKjEu7QTBqJcCYlfQE36wS/rgS5f5BMPx/OHq1KQioo48ZP0b7r
BkW/Q5t9a/jwivJYPjsBMT2GhrQHa5sHiiF/un9byLaPQw16XNEazDJ3s1pLgIh1+nIcHt377kuG
M+Hi8yu4rpx1MC5pDKDD4049N9v+yNPy/yntCDv0Tc4xkPGtD0pNqosvpOgVvn623g0ROhJHDY8r
jA+5hfQr1wvbJ1BHDR9vmtFXUrcB26Q5UsavaWisKfJOCu6V6iYio3Cvk2KWdrhr4U8O90qwxIbW
uOT7nn3J2asaVY9dJ/27VZAq13JMsKbMoyJfanq/3Ka/1x/IS1sRM1lfwOG77LyuODM1xJ8rRRTr
DqQ4pRhbpaT4MT2k63mpU6c8N8Pln++l/m3MKoU/7vRQY00D97QRvwLTDWpsGfL9RQw9RGo/rv05
KaG55VMEJrHHqYo5jZeELKOhD9j56NlpKEGb41EG48500KUH+3VsUCPf4TrVWpYDu4eME5OUM02O
TssAb7KHAto33BhLwjZluIzI8nd564uV143xfyDqKGGIdLnZf7vc22iD0RRUSFcrAoVayVfuzYVU
gK5eXRQ7hizjai2Tc+tjXPbNM1FVF3QNW9Uob/ZfOL3p7pSNdxNyB6GMA0PXG06a6B66EP6Q1gor
NhFHAdQd+YPk3gu64ko0m+LZxRmuXHPtMoFQAIstSGFBBEeQLr8t3UG+0C1KNFZsEJ2ZXoHaOBM8
f4W+TOLu6D2XbjILo4epZm3wIVFySL5BDRpB0bp3+oF3Z25xtF/7n6vvxkUVkkSQAyHzFvO/ipKJ
ao/UNqITP+bzyUmwEkfcZsDhNA0c7LlMGXHQ7tzfsl4hfjamHxxsnmTOL8cn3VfPcWDafJQdcDo3
2WgflvSrk0KXyowZTaeEU7kumddJJGsNBdqNEdD+MmwSaKy3dITf5dv06p88RIREaVe/khQ8L1qm
Rs2znU61rKg59R8VtZ4Q2SSacuRl9dTt2N0L8tVK/R7NVMaOdfnD0RGet+P49VaLHBI84eQD9oCv
pi+L/Gpd81C4CHEk7dF0SzzMrqN6c32ujjYoDL6SFox9nE6rAASQ/dJ70fRSKINV7p/mfR/QJmHA
pKjrp3ld+IZV/HnYY7BXuxOoEsJku9VUTL1oTKfvMB/JsMt9Q+DmJIAhKjcAH79uXXRin4CB/ua6
IOuEiMmoqSXSns/xyGi+Oz558VvtrMk0ecXr5dY6W8LmC84QeZ4dJdXu7t8zFNPfK1zEUQtrr1j6
rVKA0QRx5rBx/8TxmgbMJt2CKrdzUbWZZgGoEfGS+67kBqWk+C4aCfpTnAEUHunPamjoBvBY9nb7
FrLs4lwbqIx7xr9NDiF8jC0OXahrojPobgTTewAWQtn5cRM92vtyWmeKNEzTz7zMc+4uQviQGflt
AQrji1BfRuLxncTkB9RI5pThLgHqEpcCRglnu/Hmk2LuimzpFf8Wfkn8yiYpay+hQDckrmhOjMjo
1MlKbB5n5HJL0SHSK740am/j6Bd1DWobxO1d0eKPAK4PqF+VD0pXSIEbMXvjd0zbkLJWN7O7X9nm
WECZnbfdgREE5cvow9LjVly71cXHNOAR5LSGa30Kq7JeK707dROwxL3VzvVIZzocGto/k2F2MzgF
mijODL2Vq52Ueu1K9OR1J02l6QAaGfRx7/Esi5Ks/4ZtZH/5JXrZKB0DEOQXC7VUvVXXFs6RfLo9
vspQH1Hv3ty4y7UBVhzG39qnNt2paA7bHFW9g9O+8fjZCDsSFAZjb/gWzlGGWikDeqPJt7Pq4B2o
42wNGYw68Ej/mSE4RKzGwphH52/9wfW9IwTfNXSHibFJR4ie/TtJvVLC6uxNOGvgUg2AvRBBnDqu
SN6RV3CvFNy1+6dYJobZva0SSb1G+xTNKhMgTQPaXV7PX5b7FmG4f/oELtPL5ypUuNHWvE0bNp6T
RzTN8bHBCSnW9I3Ks9kyDmQ1Fuc1+Rctaw1cOg8BzHGSox3F3nbFoLbIqjyemMaKvFekAoenGE9R
HxkpILX73osfojPVdRBa8JCFX4u7gurewLgdDCD7CGYPcckoycAyc6uWvWafyBflP3oN4s3v6e+A
dBB456AoCaLTEn74qNQw2ZsCsPODlGLgt9jCS34zXH12SWc/uejXG8UjihZZ744KvrhwaJMTeMee
OiQe2gP4959IhPSnDEu0OJM2IPe9n2FlIxdbayh+bXoCuTT4S5qjS6261rQvPUNkMbZqsyegxgJv
oxCGhD+0uXeROltl4uGSnW3EUB15kEGRicJ85rtLazMhKx836yhWiKn9MFhy3pufbZsAKR5svl8m
m5Jsm+0+3kLgSd0yW6hGvtUHo0bLx74P2Ub4mQ/gWSEqZRwqwEKL4Tknn84FgAApfHZlLFC4HkLC
Ypu4rWMInyQxZocnCg4pFrYRCaQqYN0DQl9nE/3noukhheIIqWPycLZ3tqqJroQA90n3LiFZDFv2
6qkoyXn0714xxpbL4FiFYV9blF7gMfYcL19ofjfEp7GTcInfPoZCgBnsTnYfeW8drhBORXrBY5nJ
aDtj69TiyshCTBd6dh/QiuVdrmYfF9mzx5WBW0C996rnCdzyTj4cpz5LQz4e0fqWhI5N7VX/2+9n
l3bRdd89VGMFWM4amth3nIs1+yoHkV0Enuh3u3Dml4vu1rFhbL+/DVVXZTOnCWXA59VG/M4YyQ2X
zTo2r+I1OZRaZOBpSQBlhW2jU2deIB9ptG5kzIggoHPZau0unbAxHOK4ie8uvrYMpEhh7OGzzO9Y
eHwDdJ3eb+V3hK+oq7/yxUOkOiz32hvVAXtLJQ0Kl+0TqrR3RI5a9bINByLxgMd6SNXp5FPSo+7p
zUVUZcihIj807w+0f6h3lanAm0UoJIGEfmTpCNXIfk+1Ko7/jHupkWuuq8SkZhXtqp512Usf4AgV
xwrldkbStxUepn7YFwHJbH3k1sbjut1Z22/pOgzVX/YX0epaWaTDqLly5hrTOH2GMFul5GjqitAw
PPxChZo/ikitGLq7YknUpg6svOqwS7cZxwwbUBbR+leDQLBTTteLZeUMdI3XoXV4aW7aE+gQK94f
pB5lo8vFx5N5ZM2vcTPg6y7FSwKQAK+oSaE8K/X5SANWKqS4kHsyQxuK7uVqXx54VFXcDIKZz8Xs
2uYNRK0Yyr055FxWBRi8RSQ/qtkC7Cp0LRrhdj/JSqIswoTAfuhf4KP1SI5QNMfUrnSR0Y3Jx9IJ
1rTE5yPQSJ0fDcqTEhwfNDVANxnaWK6iyoZpFJge0YMY4cW1wndclHUWoMF/XNJZOS9qzOY4xDxK
8YeHnRjV5x7M5i3K2hPBibyVNNTyzKEC5QIaCQuvCaQqv3Fh/fGoOvjOzTDg4ulswuocNNZHm5Wp
JAmue++zbvhAa2B3p0OVMe+lbj9AlFAF3L+Qgj9C2EaTfmCN1c1ZDtfkuYd0D0KChz5M8KQwmTzs
9f9wtV+V6zBUZiuoKjG3oGNFDhtdHmF/14DovilVZ7SkqZOUZG2YtjcXZplNlTg+s5TgWznesNC7
t33Xq7bIJ5487dQRmj8PmL8oT7vCsDSavmyuiGKmXCvrsx5zUUkU4jFDk22/gn4VU10+sLx3zxqI
/F63VavV/IWSIW1Hd+BPIaGNB8dDzM4BznlIYhiCdQcolAV9pySRsmvScaN2Jl3TEQmaqa+NRd8x
UEi+txsIsOO5z9oDgtU1JGuUKokxXfr90FZXtWg+zWKyA3waBglQiwSuFPxUulFNn1F76PWM/bhP
d3XN9sCikSJNpSquxDblyF2kq6j78aRXvir3ooZ+PrQe2hTnxUEzEj16EPHdLAfFOGz8mM1b9h5B
fT2q+erwFzGBtgDi7qK6rkQct+PmBJ+dnbCuC4sGEZ62rQZ4W1wet5Jqin1/1hsUsyh+ZqJ0Q1Iz
ZzTdM24Fe6viFWHtBGVCSOUBfqIZdk4H4rzKKev1zroZY8qNlRnq75tvOWycgIIMSFgVeV12+pVz
xrRADDv6BPALPLnB3fehgDz7XsrqHa++HlkeD10ecPbid1Xx+0TLsZpsYKJHOJILthYk0Fr0/1di
oJ862JHrJmlIMAcPdlArFjpnd1ipRzpEHerInmptObPMBNTFro9yOBwvnKwtp/LnMOwR+vPyIaVe
DJc01y0EmqaxdpCqjyHxlK/X+RMykfRHA3A/p+hF64tihptDRhNtLEL2sVoP50bDW9GY/KR5vbpu
42Qrqdas/cCDi2qXMHznPJgvbXTBhNIzQR+tL4SFn+FeTuE/GTcr5/eMF0+kx95t7YKzIj/7DBQF
Y6dnyuWD4ehNQ4/t/Aqgz9b0WiCpI89C9BFXaDnZh6NnehL7Y+QiDQf0cDFL6QUl/jh4W4X451bx
iSG0c2ngUbcYXLygya2uZ9ePhsNKu6ZR14Kr+uMUA1N9WLCIZIQkv/WnazBBZzVw4hv6ABmLLbJr
Vy+YW2XFi0MGTWZz4znD8SeKxDpWdrScoY7O9ZjVdxNm2Ud/U7A6u/SEtFgWzITEQYVVlQewL2b9
A+042iZmKLkSTMqhUeTQgRxExGatQ9xeAgIRDrO0OD88I01Qv/edJntPRJZbGurtEnGK+PadIpZj
oSJjsQgeQZjHrNqhM2R4PpXXKVj89SkcRNngdVsuxYo+mUgX8j1Qk6R5xEygVr0jg3ueR62D04l1
UTexPyM1R4rZTIBzIQVtWlMv+K0xPCFPNEMnfKK6hFRrkEIXyObT94fzhpXtnww3grFgdyUpRHiG
PmQ2UU1qtHl+efB0VsbKMXXUstcTGsDig5fYnRdCw/YEs78IN057xuivkwO7dLHHPexty3UFpLTD
pS5egjS0ZllCSbaHqWdOHZnF8n+1k9SRSHpDFzHLl2HppBWgGCtEeUHdxS9Htn98vPo6ChSyKy7P
+RXfh6TeqNyrPAlZgzUKzcYYmPhaTDPqLgc5NzbAcP9ZDPm0gM/uu4zCebkSJrYSqjX7cPJjJJEp
NQDO/M+09V1wkAyec4OshFNk4pNOTEj1AnS4gmunBbZ0CS9qQlq2GpRRV/d/NR3r7s3ecPNYLTg7
oHLf5OJk52s1R3TGh7lKWP38jjdTRm7H85WMSIVi8HiWzQ34zVLG+EYR66a2uipAdXVhZtHj/13w
8/d1dLbUIhALKVq/GSHpo4Okg7+8xBgZb6kklqSu02g97nHuCwmwT5wukqYymPNEmKuazBwUssik
n1ixcdgt3n1mqFdN8f11xIVDuhixCPa4rzxrvw0h0ZsqLwHSEC7KFq6qTYZTwlNZLO5AoIOZr5ck
r4FI7cqFJwdvXQo589Ps7XlaZn2w3Vu1jRo61vJEOlLom0QB/FIgaI5lg86fDQBlmBKrsTo6BIov
t20uS6CHUtOnT38a51/6rezD8r3AyXf0yq04ps1ZhR+1g9K+kAVFK1TBMGdQ/LwGo93Zu55HjOYK
VCbjQQCD+iWl9y/gT+ROtGKyr+ecpWbOKzZPOk2GKOP5nlKFAd8ruY/XoLw4MUIVJPngKbRNSTKQ
fZsrAfjAH2rH6GYxbY/SNvFFWZG3DIdBtX+jZ/3uRCF4+BzFwOcEDkhZ7F+YbcwKFl0gTATGKz75
ZrqJfkBtcJ16uNaNnwVsTEXHGkgnaccZWnceZS4BzA/ZhfH8OA9nqunUNJP+jvXnNQ78ghCcZMXe
DWoeTh3rcarsdTOjTQngWY5pV20S2uUIve1qm8ktzgfIjeUFIIldw2U8uGVGw2o39J19Bl9uYD6y
45RlJqFuyiXNVEUwQo3IELm99Wdt23AXoiITcmY/afJxqm/i6I34X8k/1lqY19gXGpQAJ0ApJpke
5Dg1izP30+oSd9E5LG+i7jnTLGrFUSxGMkehVx+xcq43S3+9aZgPi9oOBarYUrf+Iaf8yKkZsjZH
6ivT0xWb/3/xzuV5jjZRG7d5FfIk6qTHojc6r4NHNAJgBASSHqTN7FQh+1jn4bWO0pGxefUEoM3X
Y/vpL0r6c7YthuHABpq4v5DSoZQzrAG2n16e7y5wdfFrr6V1Hzr2YYRB2B/qwwjw4fsTeW17EmS/
mM5au30rgZJY7jqoFhZJ+PhoOlwh8IihlfagfCmueBFF8rTxKAEk6Nr3bHrqRrO1EiKc7iOvoztt
8cLqitdT/2FtJwe3I1aFnPprjSA5aFHSDmAxFzE25zEaxP3cp6/gvHmUexZe7fsSxHl2RWwyuyLG
n1ItaGiiaWs+6dwjJryU0ZfhUbDsu1SMuN8nZleADQuWGHPdi4k5QKkvZYDWgU/r0rWvWNWx+ZW8
Ti6CBYG55Aom13dxlPHjQdpjn4BQ2DqEn8Z//GuQLIMIkt/oRldYTAMByPXu9bioPbJs1Q7Hchz1
nmPUz2lqjrYksljOKqAikVKYiT82A8P1Qw2ZeC8jgjJYqZKDyjND0T7HgEiYd+G6lFXjM7LZCOyn
EZblHcDp+Y5+cPGtSWyRjRTrCqLiknXzK0SDrcGwA1lcaidVxQfsT2oiXS+aAPnypAwAHfoGMFWS
0yAbH0aTDZUUC7e67uyROzmOSKMtXa0sML7FFA9Wo/VPTm1fcui5l7SQHmRIMhuR5qWNFZ6m8OHe
1tAMd2iioO3Tzbf2CDUJzRGKOKfUeXmFM7QZDZEl7uqYkrwIlkp90o+FP/Ywkomzv/Y1jXi7ql3c
pwSNlpyIK1rxGpjwjHilMkMROUPdk3IOMutMSGkV2Foixc5enTUrmbapUsPYEf3nwZvaDcQQIN4j
ImWgc1bQBvxPcaeCMHapmXjghpnzB2siYRUGR7qNleqfAFnFztFQRzImUyJh/bb5z9RF+Qn4NySZ
zbh4wv5s6Zvcdr3qs7Hx/di1IPNJJGdqQPcHgaBaB8mn+N+cxI8YoGE6WcH7s13zfuBkr0S2g70T
zZgOaeXVM/aiKOUEH26GcJqWP88tevJs7dG2ZHfFdk7lY0DCfsFx7KS/nX6Io6E2kmaYkpqfPT5I
zJSTSwIWiLob3oL/E0XxvcE1HPXODiFcaxy67NhcyqZw8lMg6/XiNHysLvrJw+FxCYOo1VcB3LSW
3KKClklwzno9pfSE6mw7GBevZIJ4SBcxpnx/iWNLTPGBhg387zRoWIib5rY6lbdeR1rbd4y8KG4+
UbM6DNm9ZiJVA2f9a+4ewy8JGQLTHNWYGtC04nDy6bH+5nOt/N7bcI0K9CE9Dm5PJfKT6onsVh/3
edoaDj6evuAJBlNNN7JbRd0PTiU4XGd/7ySDplzgObIg+SCwrhsbkhiHvmmJnd6YFEH1lToaPJam
0LYfCU+3cJgfSSgvzXR/GQ9dTDrbye68eM1VCPZCrkXbw4mduvV8dJkmeAdOf3N3e9snJkLWXieh
udN3bHLZotSXFlJQQPwtHhrOGxuz8zmljkj7WMejYHtvZTebOhqHMQmU/188jsrVvTHpx1F+D5xV
yFrGH7gNKf8hosnoBcdX+LLF/1PqlVNeJqws1ahqBIViDKaOp3sazH2FxMoteYRauIXz3Kmc1qpt
BhgeESuHOvf0sbgzmG1nlO8q/TIrlNy5S3RcJCw9YGaXxgoi/i4tQ8e17Pysv1H1Z28FPOdaqql9
xDXa0afShja2NQIr1VlQnWg1uEODZtcNVuw87URXfMUogjPZocTfkxKBjVUxy5b26ewJhuFyJ3Ds
2qG5V/+q45VavqPpL2uLO3bWpacHbuwWcxG7VENLthw7aiN7iCIPkJd8k96/G3SoinW/zGu9LTbp
M21trwnNhJClM7VZKFdObbgiakX/yyF/cGpzr4cB18ZZXX95JmPNvQS5o8fnumbZKdJQL4QwzBrm
0prci0k5z5wX/Mn128ueCkBdj7cbJYtqsKQ/bw1gZz5gS8l8HbcIxV8tO50jcRMDUgF17mhsYfJy
tjPeNo+3QBiyfJMPjvkEVmsy8RjbCtMKuJ0u0dD6IDwSjHfSMrQ10G5S01lCRxfISnfEOKafkPnq
FW9mP7N3BTY1dhhflqb2X4FA3XwTqSKCJyI0AiqKetVvyauK+APkb0F33TKdiUpBScy3ElEpFdo/
ZZVY3ZUza+7sGnPst1G2sxwsYNCqor9Uj6Dsdppo7blU/iLzNrp+WQAwYo3mgOK4F33RrqTmEhuB
cmlxpNSRpBn7z0MThaeZuoG0Hb4nMu3FCfkgMVvQXe8AEYeI9UJpOtnSJknss64rpqENAHRdrP2f
cl6+sG/ZAYdoHj4UafQkfdCumzJcs+c5N66x9s/EY1VoyGJj0Kdz3QjA5txQnFlPpIj9GjDlKJCQ
MxaX+YuxJL2Cz1C0oMzucFpBmzXdGjMkS7jLR6+BEAjF8lUL5fxfyTY1X13RnOfS09LoIQQiui/P
v5+2dvTLPAJOcvBv1XszE9Tm+cQ/Jl1yHrPDfpEVNG6zdPUw3TjA3NwfHrdeMxYn79wHaQN372xh
PUsswe11xLG+IMnHknuMz+7wu68sxYIL9kgcNij8LTbTXnVpX6IRBpam4Zq5FiMxyoJV/VnBPpUn
NNyoPEwnqYCZDnL/p7xdTo7ObZ37Qtc3R8FqHuYPkvzrQGWqaPNrwLN2A9fjnsXG4cZ7IDBEDpgD
rmFdBJoLRWWLft/hdy/YM5C2ligje6y81zs2oSMbYVWa+23m4AujVG7PYWe6jLkzbsGJB8jlouob
fnZP3T9Wx+d6hYOr23EQ9yv09rhDVsTPbPwuKRHwidaoi9fgxa5wvMV5lSj18/2/7FRc1KqGTpGA
27j04TKHBPhqaoKoex/OgOKGEAVb9wS1evA+stq/dtRzUw2hFA0Q877N6AIF88QotFZn3uFlIPuz
UrxKEGQCrT83LZeSnwm34dujZX5thTYEFpii2lv0sBB7/RvHRL4etXHRzsJFQEaOeXzNwyEh0ofC
feNPIuQBFOFKxqJiuu+CK1mBaz49CaJW1FwKxjqRMqCGgJJneadnTXrqQpWncwAKTLKwVpdwpeWC
levh7JceDsRjFW3Ovhml/OKmGAafO6lMeXi1wbEq0MK7eoc0OCJszxPc9aISSlkCxMYTOYv9WjPF
Oy6qOFEh+tm5TtGaR4MIZfbI58Ahk9+nsjrDxXKZ07KxGZQqr5omhBA0ucs6Erz35XeH3wCFy5XD
P+Daaq0IbKUzKv2t76q1oJs93dNhkWHNUNjfoQGUW7J4zH/9fSdBB/d9gXxcNTxNYFQG2mrALYCw
PD9bnF7hD7NqR5fUgKL3BXWfa/G0ls2DOZeOwADfQtENlBEKDiGvjnclY75zZGhgRaFIMp5Qz+OZ
SVn5ypOg2bd1vTE3qzQrHhzch4jYtpdPlzjuwfvWizQm/E5p1NBqy6PliHIrwDMs33W8w1Q7BhoO
jM3gEwaK81rPeNCqG1N8xGYbrFPyRJaAmiXRnjCO88r2iF6skFJE2zZaGiERzH97OhJN/G28eb5U
kKEMgB+1wLEFviZPt0ZaR3jbhWIof6wrMO2OkBmuIzyUM/ImJNyNkbj6jx6LG+ZUtv+/tBrW6pUd
DidzGRxkHI9lp6twszzv9+WeUF/sbWuenoaQQIolPwQey12hXRNcViLHoEMGHSBXWrI8tsrM8eiM
8sAbC8IFRswIznhXztotLudsXX3QCkXGFZ16G9zxjDQ+ztF4v++FlJlJS9M2h0K7qublEJSuoGPK
+U4H5hc4lU7cER6xXv4eZmuxrRCqTQpZHpFt5zPveioZ2xPXd2qCyXmiqs/pDxBtNpL7yLYNc7bP
NM9Nzx6FK6xmUYprMM5GMFUNfgkWt34GwSZfjYx5ZvZf1OkICQhSuZF3hJ6qbOWF44vqA8WlTbSa
Pw07ac/rzSSauQlOFqvfevHm+U1dZE3t0D4sZYk6VD2dXPBQ3YNH2T119CJUJI+KrCbsEBDJu4G/
sCya2HCouj69DuEkd2mWUD8BVb4Y0vBJ1fK6Qa4yxK1AqpONj/fLmRXxtv5nTnNj2B2N5blvqMoW
/8N2mEV7PzQM0tczosPwNYrOdm/ccikXH8zBsud5O7SIwCUYdWah0SIKUEMh9/FVVMlcZyyFXHSC
3af8fLjT9J0VrGcmQ595o2zKTbVzR11irBmUO0BUdn1yzc4stJNnjIWV0123hmCTeOOJFCHSE3Qx
qoZsvWij+DFsZf+JrY5GVAR6SYfOUPTCnU+ibWHfKJLuwZCcbaYikjUjbWyTRWVGjdmC5MpJFOQN
kAteATik2FiqQnDc4bw7j3xpPxqrRe8IpuGzxcAh8y2dFHT7UrVPUUPANyWe3ebAfyGJyIsdAAsF
8ftLKWZTlhF89qloObG4tLTXl5dAxqdj9fmfcHzuUeJ2npE6OJMa7Rp15nraBbPJjX0Avlf1Eh8w
KhtJsqieebe2c1TuYYlN/le84FQUTWQ7kYfPuAbQHsbZ7V8VyJmNVHD9NTtcA90JMdyWcLNAi5je
IHR5BOP7lv0OpyGaTMa+2X0rjSPVgiYqHaO3g9DF71DsMYykGqbdzAhsh1NChUBpl/JeoOtn76zY
UaIW7NqWe9/ysJfpv23O4ufby1uKsBci7jE7L4VVatBUDYI2S50XF5LrkEWMcKRo0+WO2E7o7RV2
hUfro2ZqD4vZt/eK+IJJpr+5uv1tV6V/bN4uvnni40bZZJR+vtV/0go/300W+oF5uzqRa7RD9opN
hivhein/hFl9Rvb1zT/VCxN8k95W2Zs/QDcPPl42eE8KhDmqppxDLkF3TfeVfanAMX64MFBe+eU7
7v8oZ4wMkzolBzUO78G6WcWINbCYXgEkSLcW5LQ9910i+8WxVeQWg4aHkU4rUWkH5PaDb0J8ZxrX
+DNhJ/cOAQllS41VGJU+do74uDOGHgnsl3fHkg4tBLxuTCprPCeePTipbDMVFpubPbJiLD60bdCs
9canJ7UW8gm+WRSPpo+gZMMLdCEL5nHsIAiTMBfKTUmRk16xKX2B5fhX4SJYKzIhdc/FybWwkC7u
w88CHdUzXwwTzPgei3NYn1H58KNWvoERxC6BVQJTOHu8LKGorMJNk2s5cfvfd7+ygLIfl3HA6fEW
N2kOcSATDol9Cs27/8KhYlNGICYd6W0WNtApooFGIXPLqL8zYZGqkW8sNBerSAKWXwaKE0lw4SyT
iYGPmtDOfn85EtrjFq9f2BszwDyH6pYvF6bWKkZmIrV6JthKPmnzMKpFWf3lcMV0NSnhZLoY7+se
5CZpLZw1/TaipMiSQtIkQFWz+LhXPbrHtsgtn9Z4ii8IZhjsZpkf1//0OvGtx2KCHt5KLCafMfBd
dGn489JOjD63ZIELhjGO17cWqXNVUGCzaf2yH4cx4r4SBp+bX6DzWDJC7l1Ly3+c3h3mlCnrq0uR
4c0dgACsgsQnj5HmHP4Rs+svL21g3uXMxWvBbT/v2v5OWdRlfdeWKHy8YZTDDBaSZ9YkOg2rqd7p
uyGuKgYcz/ijFgfsuiqeWfJ44HCiLUjyNw6jbJUyzALiU26HcuQCBDq+Gr7R1v+I6kAKzKT6sq9h
uuXjvESl/jDJ4QqeDuhl6rLihme1dMFGvpSAjILxnyl0Zl8wb7+M+rpJx195AW99+B6nNmcinJ71
Qsl4bIQoqiScr4kybSlowg1JTDMBcCqwBw/43UZhRiaqccf4qDK159q/mM30Y450LyiPJ3reFWIi
BDCf/+b2yh0lzH1FFmfwMOGruqv5Qctvhq5IYfYeuTsiaMt4DBUWz0NiGZ6TsR5CUFZ8pQhxdQt7
z6elQhg4QxtIHdtbSVLcbGqqwNMuTU35yr5Xy8mJYxKUaFLxPCz4McsW0iEFfBKs8PSE70sXENRp
JbhF30iAbw3qq/+9y7GTk0Dy3lWAz4VIpvZitIgJJBToAZ4zzd0NuyLG3XiarkzV+N8pqQruHByU
1N0Nv9ApvKpS7BfMnV2BWiias67Ck+1T86UenrBwL2akFEZt9yBUM6hU1iY++DefsS2LS3vfjf1s
sbmaTibKokoQcebYJdGWu0EqqhkkA01OT4CFarpiGzBrtSUX5Kbpo7Z1ddkL7vieFEkkwygOF4bn
hPVr5kuePFmVTy5bhj/MKDrRV/fxDfMQyzxw2yIC2TQ8A+W75Anggbn1pv/+uc9j+W9D7RUuCVwO
IQdc8PyVkbxVvOTA4ml3Dhzz1raZwejz1+FFenQkhJuoRNgmsxB7p04mV7DRRiaByjyhmyIXRHJF
V3lb9WZtWXDzHfi046EjDi9ldKAOpu1jEDjHHWqQ3vyvW7hIbglT9HfjMDmMnMKykmav1NYncaYV
B36HIC/LRfkpAQIwzZ0+iJGrPPkFUpk78dyFlsnOFpzIm4lbRCOtFkGzmM7BpB2/lcAYJ8EE/qo9
eZ0e6iRafx5myY4+kS3OpMXVqQcY4Bl7r+G4O4EmMg/Vdz73wQMHY7P3cguuJ1WXPy5rEIEJHyHS
GGUbFcdN67Ntyb9t6whvL1KRGHYsVPinleo42GS4+S4QdYzZCncbbPABR7ttnbaLLescmLv75Fjy
fPR48NjYKQThcCLRRW8pnaoa5kLb1REHau4RhwsvfCIPulcQPIVmcYC0Rv4feerlae3mbRNCxkSZ
NL9/M1ld0sa56ixFmwZrLraKPJD561FZk3iwvK87VymTPYj9AMZRpWIub0SAaNE/KpOtRz44+Cx1
UPT2NKxlw289ENva9kmMwqxXvUDIpziB6yFZDl3PiFyMqsLQbnRfR5ORsUGQwVi8difraNS/hKy+
aMoDAEoMab48IK/6NP33KcU7WjRkg4GP//CLz9lWdYatZsZgoi+Tgu2C/+oCVecJN9SD7J3SlbVt
UFoHyXGbv8GQH/IBtWZU2gxR7i1jWZ5EAdilTgBPDQ+5w+CO6zY9B4Ox7YIQUrS7U+b5FQKEMC0k
FjlvILoFWd5DvJThTLh5d5xrVpgvkOTGgOvF9OCov9T5W4rOZyXW0e8VzCBOLNBWB0jTI/IEnVgf
arCcChTfXHP/HDLYSRllZ2ywg79khflBrGgi8/cXEJyuJ2D8nX0BLyW7+j9lo1Q/5/bb3D/FqvjG
3+mrsctv+XcDF3COy3BYGxW9lKwGKSEJkxH/TuRyCxfKsqpmS9VOW/t17g88E5/EkpuOukMQQkys
lybkFPHwxKt5tjIvcfieu7sdf2jNaz7p3CD6eDeCT4PEDiAIfWO0X4w4mFcgii+zgwE7m8s8kK6N
oww2GZ+rGVyxbELYiQ/9byhmK9dH7UcHYqLkSa+TzxsrHmVCGZqrvZU3FhInoJYECnWHPS3Gefks
WVmPWdOjwPGfKZYztKJsW54jY0gcJZEPiSTKLEWukdej/yHJWd6BHvb7SsV6O3Pn08J8IsFG0ID6
6a7g+IsS6kJPdoybLOTz4+wHCHdSTNH9svYOQJo1TbDHbuFqkILWfWL4yXt/tzomutvD30+t/ddx
wv/j1QwaWdyI8lYG3m4P24q8FpFt4p2/qdV9kgap9tltb0QVjZOiWOaLI98CRnD/93uJUDpvogeD
VozXaBEZDE65QMZKkOWKTLQn8EVpwP9nCAV6ZdHZ20FZcjjVt/YcfKrdN75Qwt+AwwhW061XTJOP
XJRCH01+iWvdPGoAhCz1YGuU5s3MltIsocfiMZ4tDFsVBUc2R/wevGCKM4rrJjzYx/nQdwznZ3+k
urjPPRYI3M0Rwj4gj/Prryt7y7bqnKnXz2bhk0d1ej+afahDkRSxCBNE/09Y67397fuJlFbsFUI6
K3iGI4zM8MujrBJBNvOCa+X91HWfxh/Pod/bQsMATwgdIvjOygKQlLwwlp7ulk1Gz4YWkvFgR7qW
8P8kmf2x8OUMR+9/CVQQ9u1oO3tIEdHRxibv26wrnpecZqZFIrVW4vndoEgbfkJF87r30V8pWwMr
/YNaAzMk1SrJSVsQbcV9mhulrwJfCdhnG7VnQsfXXwoAsJV+u+rDRkLGL3ELFZWOZpmzaEVMxjJz
a/r91qTnAFh0AiVDVpiNO3Fai5q3nmnw4ef4nEkNo6mg2/Purziqjhr4Hw6IL7SSb4TYRUKTHVcD
LjFf7NbpN77pCq/gSS9Rle+CrdClKm0QvnP1fofzvoiTAcWCzWwu05XXIgS3dpVdbkPG3pVdBqrJ
HthxfPdqtMZKGqas9/iC6b7xsaRRTtwObfE0IH9uWiaaS4R7qD0mgy31wl7BN+I8oUG97swOrdg6
EFIDRZZBF5ZZgG4jjNKKbitzGFMa3mp5DfBx78rpePbH+oKxv34LTh9nfRv//4FaQuwfqB4nGmR0
7RNuo0h7O/lpwrKV07rfLzQvXqzGq5BlK6a7NDxsMLihbAU3zR+5Ha2+t89iLNMpLH60EAeq2RLS
3AzCWdw5dvjGU9UM1I4I/kqeyJk2iCyMKUfAUhdPzDbK633XDVvv5pxQmFUiJybMQcg1M3+OH6V5
wC0HR3xYiyxBbsuYoTiGClyDBRLerFQRLTJXjVBFH8UsSI9rSeSAg7BASwwOiC/X4u9s2nkxT3Ps
FuPwH+G+zKFZ5fchpHZcYWuL9KUUaft3T3/nch6MYXAzO2UB8ObhrJNowit638tC/xfdQ9X5Bqst
U7CeEU1QZGmzOcakW6cyQ0Fdh/ntcj5dX/mi8Pg5/jHwExkD3ZydbyrL6jsDgbJzFcuyoBkgdFQ6
0FWYAPgXnun2KZlehy/GYevLedsCv/MWtKHZOE9MDNAB0TLmHs4z0FCquizmx6THiFlYEBIlYoAZ
4IDwPh58mvBWd/s0zlZ5vE0wf9gKzWFW0Z5n35fnnZaLPv7wajTTyZ6FAimuyUc+yKC9Um64gDWx
XXpsbXphRBMi/Nvw1LW7hqqlMhL1CMdKYLL5+O+VsF/mEcSGdPT5+mGzzXgSFevt+QTuKzig2OqC
+Q9h4afH548cyD8AQhhJNrgHyp9JaDHZu/8DoZQ8eC8y/zXdp5Wax+pELy7KTAFUXkl1aGhEnDyt
HyTNN/NVxS4iOKDmAv1uTuXWNtgBxmZ2rbahmfj3cKHvLvNdZkeTNMp2KVOkiATwa8plGo2/uyOq
k75U3Z7j2GzxKCVkqKUWomm8+sP6rMUUU+tla4nev7L2dOklxtdY1kXCovwPp5gESF7lsVL57etF
fiDJeKf/LDAoAlK9YbAYnrbmpRIT4QxgTZJdQYsN4lSbtLxiRhvPamEVvcsScyZ0PYTrR2JcV4mB
jOBgpc/sYP6l57JC7xqDh66HqEE8VwfB82ASRsNMONHGKQfUWTZGucMNrD1uzymLVWExJn3CuXgs
xxYDJrUFwJ2NUCfrPR1+obe2Iwfl/gEvsbJ8ddOzyQaFTWMuNHLXWZ1urMuVCs6jR2ji9FMZMDom
lMOFa8XqOUaF0KrIh6LzZ12JL8elp6VyqB1isEALcj9i0UKz/RM93PE5S+PQrjAYWz0TKXapAgUi
v/RhKmkeM9m88GAuy7emoXs54S6vlvwx2A61cFevFLiAGpzx8sSwMevTEQzD2oz3UNoYeyQpbGH+
0Yr/4gNJ6/q4c48TXKs0YqR7UsAmj34LaX1iH0kCkNUskgly7AIyDhFif/zUdjsuiP+QH83QwLur
HDExS1tyReu8QDhCt8snZb9b5BtWsR0039Vsz14Vwk5nQyM7m+cdHLdbcv1O4cBhVa5LpqPr8VH9
mAMsCIcRHB1PoZRVgGHQwNwbMIlcg9GebLFDQYdGaJeShCqQl8DcKyoAYZdPZIgDkIhPfpCEZ8XN
J01vP6vlzHDf+2t/jkyZlF+i+GifzYXjPfmM7JLR/es5sX25X339iGR9OeBnNhugbE/01yAiK8lK
ZoeAd4bAizYc2LaJURKw7zt64bSYdji6WCM0XQthMkPvfzbNyP+fhYYb0im0uLX2/i+f76UZIerC
Z/L0DNc4sPL0GFn3dapFSkCSTeQdaE8WxhUwandlKIqBj0ekHb4sOoT40dyx+tb3e+xz8FwJttPz
j9gYnW+R5A+sgTWdevKZlNOEnFBQhIe3dcxIKowFERthiN1vfI73shmmwOe1o190CfZFZTL5ShOa
zo2TpwcUxUTNDr1FzEtcPDSxoetZiGrfs4+UBP5DRcCnS5lTmHIWYfqy2/Ht72T1FPVhmffWQM0R
Cy6MrZADWqQxXwA+vHOlG6tMNkA/tA8pJEtE82Z1SPx2BrjJzNJKVfs4x1Y6xcWB5HhtA4M68lVf
3fTRYk4YKX68GHFQz5ewXOlyVEQ9aTs6neQMRzypDDEcyKsseA1PM6Ly9VrCpygTP8XIrlPhD5BH
4eehVfmQgVIbINRSSvFm6scCDgci4wdG2Rkjt5fePxGJbpxOPiBFQ8XcnLvTJOhHDfkUkNf+Z7jg
QUKs4en3BxVyqxsa46KYn6xGn2uMVWbLEOt+XXvTkdkm36Pp9izKKcia6H8p+E9zqDRBMf8/50wo
Nu4K0KXqkJd1jXpYEb/24yaErRyOTRIyKMJ9efrcMGG3wcCGdBB/t7GgqEpJuDPiasjfNh/CCSND
hoYXjpmkPXUA8Yu07dldHhjJpuqzma8WRHo9/KsZKkEg3M35yOsIRcf+5ZUcW6uuGqOREjsLFdx8
CanG5oeiLjYn7UfBBHO6im7OfzrIJCzTUPEhmWp5+ARL9/yhu/tyVAwpt9Cg/Bo/svdEbPnXsEay
3Xxktq7x7lvvBl+Gl7aHj+vZBC9XkQe4oXPyHTc4Rn2uTsb+bMRZQYCPcO2R5SlD29luF1uole4K
pqC9QFA9xy4najTMsmRT8hJCYyGz6RcKjDNZVjWA5FhnIR7WouJxG2glDClQNDAXQb5hTbRDlRNc
s+ZZXQBEKZjz5XofeHoUsQSykgqdEyiphEiC554TQeNh657HYiLKtEQIUskuRo2cmMKx2bePcJpd
cWbEbnI/NUVoHc9PW1NkBVXeswouYOqayQcmurCUdvSXpMMRQ3nEhDfcHCgyY9bQKg8yjXvj30bz
NaeQNRVhfEK1un/xo5fgSheR0v3hucMhd9kDItzdP4mhdXcHrex76YyjPnG5r+LOs4gcczaprry3
cX6UAo+vOgbqOkWUzEsPq2KM+DoY9e4SmeDD/VWYykAovAZgqov4mn8kVgwzkxFjTfaGsAAgB8Of
Gkt3gGZsfAnMLNMRebLRpfzWvai37a7HS6dj0iJwfUySl/dwcDe50Ohas1MX/v9qbjDioRuFCjHW
EC1DW7Nf9U1WSiWUIFyASP0u2YMIUOqiKC3hxP1BG9PGoW04G1Cyitli0o8hjSSRfSn0P3JyIvTq
l5aIySeYAWyrqgjNjFuTbmHq9S+2nkXAIdhAo3Cmb2AyPWaDvegDn+u4E/wQgChjToNwqF13N1Rr
mwqdyOzBrjILovCP/gy2RZU7CljRupKmRIf1e7svtOmTztW7Osnufwzx1N/7VsDWz+5iJhN6CX8v
ckWXgCC3sWdd6dw9JVnqlcN/zmZRjNOwNugKd0AMfkY7DmMcE8ScwaXFY2stIzJ5qeR2pKvUpgEi
WBRl7LZ9JBNpnxCopzGXtGls/fegj+MyoF/itr19FTqA1WU4TlUlhvYQcGNHwBkqCefrrP8XJpHn
sQrMafX7HkmR9toXZ+SU1CHx95T38dFmmrBQqbptLN0S8KpA7EdiPNGltofSxwMduBPeOsTBmqc3
GPoHBmPrSm/E4MIRk5pc8kkLDIkd9+m7u0dSZOqpLr/oc7De1As5vqllsFppumoPTnuxrXEC+Eo0
TfbJhTS5ldpPtoj8lgAG9waZNa2Nd5Wgk+H/hkDhpyJtf09Df4FFMt8xJB4vmVIuy/P59AWAVV3j
/kFnVTmeIusPV5lWoZvjpafAng6nIQcMCJgHWZJe+vlgJPGenq5BG0/UHgJkPnJAFDg/GRjDkNGM
eYvYn/6J3guTZRq/h0rEAqKVpIlusagplsMEq8IAWjYLGhDD2ravXmaxqKee+fQAFgNCodJ2dQtN
vs7ZLyxI2XgSlazH9YcNpwUrGJ4yFyKnjaFkJmO5arLy2+m6Rh3OgliS4gXCo2J8Xz8J36VXFfDi
De7MCWHnfyHeObeFsrYoV7M8dd8WNO0m2CQTmQ/KFEECOpVWHpTolVQb9gWiCJPDbODeVc/DQz0a
Pz5xEgpi43bXlxVqp98HJw0vdwscvAnEHAo52EMH1VNPe36d3Wj0FytK5Ac4bNjBDQgBKa3q4r2v
FpIYhD/MNwnkdVeyNcoUI8/6BaZx1IFD5Mav38H0g8kfpYZahaVGr7lsShwOYDO5xLjcBKai9v5O
GuvNBaXe5HDIxsVT1VKBRNSyy4IxdkIoTX+cQHv/epqqNTuZz50llP/5PBfso5birkWhTw6XGxGp
tvl2nyn6fXr8Ulxn83a8eW6ubbqboXl4tT6dpX3jK8nTg8zbeFfcTZxRxAxcj4zsCQcDFPb0mT51
+TBn7z0lYp4dITySkl26WgeQd23Ha6dvejCc/c9Md2UY1+afR4S6SF/J6W1q76rrGjGJueNC4jNA
70ao85lJygG0rCIniuKqX6aInFB2fFWQdyRn+yzWWbrdTf7pYMWqNY7TR/7N68Rn/l06ftxHWG5Z
u80q36bSbgRkaILXcPdL89AeB9j3978FQDNVpYXdVglBjfDCBwUfr7edUpZEvmoSTyW5Raf2H9+Y
8oiVMXLNZbqasw1NeiCthuUnoZgFdxc0Cug5rMM4pweoZWsmSriWMgfDPLpoxOHNwklmCozYqpqE
ATbBX+/9ylva62YfsIT2DUEFwNabYj0UW1ArOQt3ArGPIrkG36BTaU4yLEU27XVTPSki1YS1ebsL
LeeFrBzczHreMJK6WWM0K9jSlL7DnQDPkF/QKaZiO0SA5ksNTG3p5SdpSS6ak+ONA3jXmbWGitsr
WBeQtFDQVKmnyK1wkhMOJVK9jc7mkUkHtpTYdGfUz53S16oC27exMeyZwoolYC1WPBgWqWwJ6DlS
dd2+Kx/pHWhhcSljJ0mmEaR9kBZl4ztI5/Ol/u/ik1FsF+V5ULxZ/4T5ZXf6LHmyoXRwVlYlUBNq
6zIBkUQt/HETfBhs409okoGC51FwbZBFw8f6BK+CZPGcJMWwW6xX1hsFDJdvTBhYXZins5YYdPFG
JrfKynDGu8j2wlChEGJ7wGCHxw0KY9hYrkxXxO+Ib4AHNzidZodI2GSEcYc4GLit+oon297C0vQ7
jQ5dlTVg+f09btJrPFJBayCwEWd3zrKXeO4xvZ00IsESSq4j2Iz3VFGoUMqh3Ccwx2ZhBkKDhhxi
tiyoDZRydCcgWuZ6SsHF/nyYkVZDPfef0sCyRRYO12bL6GpNh5Sx01X8MRcbt6naOBUtTQp/oBXY
AqX96il92pbVziXvMDa1pwFvZgsc8KkRoFWh0HJxTte5xyng4d9FW9/UxRnYf75mskjjEIgTM6Nu
jdb8kmvZ3JWH1J1rB80jqUTZaJKhtpMdrwX3bVKIEnS3V1iQdEWdaB6NnoduJ4oy1el6sEh6VaP6
3Q5iZ9XsSc3M8LYjKIm/JAljQvdkpl+A7Ic6iWtJapfPKNM6T6J2P2D+cH7OTNtEcTDv7ihcHq2K
6Vb33iAfYN3KIMTgCOZhD4BdUl9uwBW3toFQmwdGpi+hwZ+KwJl1GwRBrExOw8TrxC+Rs6i5PIvK
b1/INm9zvodUR4eLGE97Zxh/5saiWhuHQFFF79I4B01XB2Dafm4PUtAyCCEbxKSctwhzR1xGgWTG
Q4Wh0uf9MegOP7go+YkVk95gVloM3N3t6hdEHpHzuNA46sH+WwC/qjcGrXd9xo1vClk6k1M5DIGJ
cV8KEdq/NxkKB2eMT0b2QeXDjDRjVTi0RulEQx6/Ff4XkR7JAEmDAKrU7i/78tp4H3q/znwoWC+k
HXyLO5l0BZYchWRQFlKcjXbUej1FdTiYIaPZMgchcZu+bW3iJg+aPJUPxmy1S6SmUPsrg86RfQlN
OnsqxB7f6Lu+C/1J5hsVLgrLnUveYctzHUfs9Tx7YnEgX8Wwc4KpIWzuUxY/9FU87OYlhGsD4isy
8pHy2PENoMYfkJh4bJGVAv4Xx3KVQXMd0owH4GYnPpSnOAgvrfg1lfFKp6shCtr724idm3sTfWj7
06cmuABYvqwRIVB43aQyytIfTqrPSt0V3crB5UEcEisqkenqKOdxhqreYKnXLQBu3dLNwnK2Y7Z4
/oiEq6Mvy8O0xJ71L9xOYBtDpHsNmWCYSgnX5Rgl/vYuxYJ9dtfpy2zYru4yvzJ98ufWYdQT9DQ2
FhMkXuckHGUcq1V3I2hHLBoFIE8taeSIZTH3hnzNpuJvXSQWNFPtovzEzJaNHPHkmGvmcbpkxhVL
LsDjb5xik5WdSPJ/ygPdbHamA78R69PfzHNTDSD/5WQGsGZ15fsEbwEv2/4zrbBeSWwwkVqCXfcR
UMa27L/Odmlezx/yXbLhd9fjYgrcWXGjRHeRPHfpRW5upBKjPfmP0ac2z2hZOOqDz1JHTF2ozTm6
uJ7Yh9HD426+2HdB7uCTuriTWbAME85Vw9RLmKSYaUmBP/8ekm5ElwSbxXjsEZnF2zyCXV8Bt/qx
a1yESi54MpKdiqk3yCvwEZa+gxU8qgH3/pO7slWX8t91YOQ3lpnrU8DrS4zssNECvdGypwkDKPJL
y3ynuzyk23be7KOHLoqcuDUv/SSzZhJlWhi5dZeq0sjDPehRDUka1L8xudVJTJrP2gvuGq5cba0Q
wHd1c1LhkMQoYpT4NfeEgku1W5S5XlZW0HS9WYPjl1y+9g+agLftp/9QW3byJAz5ZxiWDJ0xvr++
iK8HR0ZZHpSauROGElKeqPZgHlVCQiyF+n9a5qhNkt08ERX88AF3QagpnfYZhDPNhT4xuAzCDEY4
NRv/+AvRfVACgcU2POZUPLqaxMx4sKBGMa6Gp+Vzt+ZsgZghvok8H8fFt7pRnAXlFkSsfauY7MWR
A8LiTg3t1TPrLF+Kb/6n2kJxqOlVo1Fd+vrdG5IYWTj3vWNkppYT7fTlCBcOTMM2mnINsomlOI3R
2A8kfbLqw3OImizVXsWd3Afot/sX7JBEnrwKLkxoFV5Ll1ZLnxlt+xu9J4EcAuHk5DUjWYBzoG3n
TDNjo3Jg+RElh8v0xE7HWONuIke3q0OrGHRhsUlL54T44VDzTBm5YC/jduLp2Z0ABfZJUcUq+KYj
q8dbC6UvQEIioKe5CfqvkGgY61vYIlcrcVtobmgpvGxCzPZequ8TgcZPt0+PGaeAa8uv3dZbWSkY
KXviUdoAHnhtBPzglyKXZcwH1LBkP0P/nExaijx9WhXda4YYXt4YKA0O6bhshDDHP97/krUTtCI6
Ec4WEGR8jYmT4GlhDWlQ/tGCfWvQE2XyhKhJCZgQcA9gdjajXR7Dhtcav3qh+pBUAbkyyVAByAYg
6IkmDRs9fqFx4b8LrjWUgBlePPbDcGA5e19xMUzrh0BFdvWKFakhmdj1BWLYnmWuE4fsaN0DOKwe
gs34LcZofieFJ+d7BDBkpUfq1c8IthCXjozCk1LgZ7LWPh1U9Bslr5zV19/VZcwDAhoKlbnip/fq
z+nMSSh3XDCbVyZsquZwDFD7C5I3APjWm3qDG/+RNUNUVx3WGUZHX/l8s/1DJXWIsXFuRdAI39se
JuDvok3Sl2JAKm38XqwqAC+QM3Sk2UkyoB8KKdy6VEFFK7zosIMRhIHrvf1/yHPzC8y/5qFznxnl
YUqp6wRw4KYWjHPnFlWQSjX/OwgIhJALPJ1bbH/61dLfI570Nk/rjpRHRA4k5oXKb2we/2Nn0llc
GDHSXNbWvkSNzPzCHIsvFct18Lf3QBtBZfrpAvbxcrt5nCI1a5fTOt8xzsHL8kaCDo9EMMpu/Rpj
Lu0f2lE/G4XjX8dCY4178e9w1mxMJsM54gQYCixvySlJEYNUhI2NHXFuQqld6eow2bVNEjFu66c7
TprWuGQt1dt7rM5oZabBoTfTRT5pdVXeq/ks0eJQPqlY7Rnb+Ob1gXW5S1RbifvxGDuEVQbiaUYy
C+SKqUkRS44t+JJwxSqKNYqEvLxR0/DAASA2QcCAf3vws0MhUaAqWkGQJ56FCpqJl/AJNAWaDV5k
M7JA1X9YLwHdgad81Skaa0/mVb+AFrwRM0g129VbAPk3rV4EZVQ2dFNEDIJ+cFQoltQPbdAqve43
kGqFjzut3q+3pcxX98tXAYleBeYI1lzxerLzHRAGh24cYtKTtIUw3eAyL8BBtVXCMJeZ8Y6XBR52
2LffCQvJAqjYf/nT8DbFyNglsl+sbnfJLns7NxPfY6divIWCipNF4XfavPVlSiMz4scyrtTbgcso
TOfJev3tXm97UTXY28UIrG0JUBC4P9AUbaFClCEhNdzfIialsln3724+GoV9DGojic+kOZrd1vSm
sTwaIwhXatqZ+QF8IX0Eko0iBSh+Ava6j6uEN7+aC8Id5xRgFCf7GkVoRqOyiLixnXELvQwgvkTo
ZqyAOrDiBmSQkQkK6kaNtIAhMPXXWYcu/mY7DXGvLVrpWPRKhLVoDQr9l46kP1QI3bpzuJUFlw+t
3BycpzHMxjUCFDmgHlqkpsIlqQlYeM/PeMwkDlieAEzfgzkRD1WWxhte9rb+uaBTfXtkAPsFxemu
tghmyyzTI+ub38II4kGu5Q4kta2D89c+mn2tTs/W8xvj9iubNmOjK5WmwaFbHW2CUeX6c6nw8Mmo
JSbnDFIvKSr03HHXgsH+AWhp+Qt3x5M2pK/4IF24brA8W2tZbdJOyTkCF5tmJ0ICyLdyPoegA8UC
xdFJlo+K+9p+76r3g6Zro1n+ZjSfiOJjiSwuA8bxNMNUm3hSobbul8QWPzD8qw0LDsNrL5oA1FZC
MQXE6uu5UTShW6+kUbw3YXJdywCAAVBGhPMSJxiODvtprFNx3kOQrOhnyJq+A5Yw5jW0fhSoiROr
nOxhV1/IlEvJwiEsCdXI5fICHwmGWnNlc4hVx4/8qFDV42cSzDod1l1+GQ0jBP2ErCF+gHI5H45a
8DeNeNDzT1iTVi9iKj7NngUFy+QYK+YbIGqKQW0p9A+g2B1jqR9WfdFR8Fw2Yiv9LRFmAXD7sXdx
F+sk9yMqXxSPf3ziXuDFlo/D0JhEWrwemxT7DArZYINSLOQjj0pPBrshUi2OucyY5VGmuV2VDq/N
vMvoV9Hf01aFTuWjBSiJU/XJ141ZWHpqOk/TKhdLRi0BHhdMaGDBT5ttzLrYamO4IZvSWgOLDqkh
qi9ukYATKHFiLQoRpQRGsvch7OiWsNAAkj4lWKCHjr4T4uUumrkIwWhENm6P0vbnJiLLLBUVFrkY
uDb+9l6FxLgfsOeHyaoFF10ZVtTi97zHcfzmWgUJ+1GKDkutwvm+f4kpXrf9e74nOeBQJvZs67UH
c0lWYwrgpFDs7Wfay+0/ySAxXvi6g2GSJCGGWPzt5dLV2DTF2bCzdTi2kZ+k2w4uKImLKVItiJXv
w8HeIuR8nGbG6DMdLRnkx9CJIR6eqOd2ZrAF9WjtSb0AeFB4EbDEtnFw4NyDNtwnKj0WZweOOTZU
GvyS0aGoYCH4dr2e6NuChqBtaF3OROGmYKNxbFIC8dDE+s/DAxdLTifG5yVR8DYczs1ZpwM09zwp
A5S9e5V4wtFtPlrVhlY5jGqdloe7WiU7eiDzD2seOTj/VTGJsBQl+XxWBxvMNOQ/A8jTk/0OehAl
yCGiLWSSxZ/OOd1QeJWpmLof+gjpYuv3kky8ptrw/xVOchSw1Hz2ENztoznnIzODZ8rmTTpn9Fya
b0xku4Guu8BZ/YjQTFL4ly96kTxwzmj8QseoKgnXCpulKnIMo3f9skjqm9q39PPGnyGljBlfUspc
SG3KNesrvew5WUHR6I3AQDJ5SuBKpzPc1qvAK1yIpSXNScf/KCz20NtJoCKaIrhAgTlz/QKKdrJ9
j2o6toqAQpXTkmWMymswpYbAa+LxYy1vNJ0PAnqR3Oc8VUiwoE1CoXaRJWkNWRwdQUDkFOQZ4pJM
ytbAjacobeXeJKJzx7o/mr6JKdGpHKsgZjwgPwgjr9xdG/uc1jBiZegeMILKRSt3zuVs5duSlV01
wAGjhTjKRpIQsK+EZibI3M2FIz4M3FbhtvcVzXm1fI49h8Sdq4HGLSWuUwC4L07uV3H2541fSrAi
KHCyJfvb55WezdRGQ7L9ZED4LmnOzTKtDCJb07lcSIwx0Gg1bzuQM5ercEqipfJlWnL/ebcwdgj1
uBgE4URTv2c3txzbEI3r0AednJjVwtGIiwVcWp0HPZUm2+vCH9+ofJKxi5VFMyD6OpuQVedwotaE
NiKNaNB4gMM6+Gok+RgyEfhXALPi6G6Zz8zgVmgQifBjZOwAYEGdJiBOAofk/peF/PIUFxdKlNWd
wJSXthtOaP5YPtzvjpzzBI2K3tW6PAOn3q3y5HCEwGWYkKBadno+Lwv1GXAElDTZoF0m2N8lwbQz
JJsnLloI5v31WbQHWzjXV6sr2Z/drnpb5e33ty8IQyh/rVTMMGhkm08tgUsrCk7qXO+Ud0slWFy7
s39RzR+U58FEu0Nw/mX+JRGxWYtrex2V+PSSpASJjSR2kHw0JONcPorGMSfLPip5js0F5kVU+aZP
T2Dig1UoDaBjvgm3ymNTY3KqMSRWu9DS1uDZw7NUfEJgWdURVXOZzBbksQI36mOsT54e2EXlUke9
Art5q8M4leDxbVbHSeBQk2UunEWleImJyrGij4O9/akcPKvqke+iTinQfYCwWVsQqsQym4e44jcT
C3JOqSUoWmh1YcY4YyI8tQl12X15fy8HeT/CCqlMrrlkkyrz3vFRzXZWj3oWgwBJa5D8Y9CslifL
xWOP9uYnZhof1XtHleN6pKMldLKiD8iHV91xhgX+rcnkSZym/RZY7lV9BfBfD3kXTKKWHVJkDsZP
bc6IMvYBlxs+UdsC2f1FNRRMIGKQqORDGW6MggS79REFSilsh+s5yATQ0LdC5XGAXTmUW10CH06c
XpXCjJ4/PtjaUV6mYZv1zOO1XnNiqKppB4VG/yi08dhSKww+t9NCsT4tdfoSJtuMi1iaNvAU4Hqi
DbXx6/GBJI54Ff81CzfMOON76XA78cxVFSsHXrdxccEYxJkEWAAaCCidXj1c9Vjb/DWGA2/21pNC
IKFk+BqE0miocw5OF2PT2fOE0irke5I8xQgZw/Ey3XwJw0LAXsva1FaYX9AjowsHn7FAQ7Q/Z0oi
lpIs1TpeSAFS+163wOiDdznnRPa4e9tp9p9Pjz1nt1K2wUWgBAETaZ0tHrhyuHnd4W7hKsAxH3K3
e0N9T6a0kWfzW33opj7NgWFU4TEfdKM20cyOHe4omDP4w9XP4abgUo/y+NRq9vMOugytzaF4H0mJ
TKKtzZfsfSMm+lA7SyrZzlCtCge62Fyb6ytPo3V4tIirxSWdEKT6ztgtS5mVYfqGOdrEDsjD52dv
XBVm/rTwNW1Lol55MEm8EYki0m92kt4BW07IrfRx12r43CPVID3GxDhl6jBQyF6tlzB0L0IIMiUb
/T4fxA98N56x7mIVc9s9VPymcCGVER+x6Jvh1+Dp/DgaHO9DJbfrmXgzpCikBYJSoDfgFlDBfPbm
QmfgWiuwI9vT1Ta1pNx5aD/0dSID3nSin069kDyfP//MdA3leOFmHc8OM2P6byg8gh9qBVEW3Pn7
BCOtoU+vMI/eRSeMP2xN5mYy5RoAN7CNxc3HFAj8oH9MKNFXxBneIXcwhtGSPyFlkuVzKqmGLGUX
Xxa5KNxh0EwNUAQiLkZQhldLDnWE+t0ABoydQ/S6NewkkuQh/ACBbKQuZk15RDH+Rg2nVNqWAupM
rxXLZhuTwq4aNkNWReI0+TmJSKdu14cvxY4iXvctQACmSjZIOOaoeeNMEllWqjzzrlCLbxIQn6Yi
RlolgMKieOpftNAlw/WiGdq3RSwH/7VcJMtuSg86gs/wlE2UWgSiG39ERYtLkFXfbDtsgLkdM0y4
Su2CkNQJrtswmiBjvHtKoHaisTW/gf8WPb0yN8hjZd0Kj0bRsAOFaSTMV9bsvq2esWO6stKH13BJ
G9ITLAhR8sY+UxxncPNFiv/Mo+GLnnbSSGgs3yhv4q69Oda1L/5x2uV1BX1TjuTh0uNMugDWQVkC
GISmJAF8cO95iR0k+H4wN4F4v4vXM8AQw1m1PIGwpIjMh6/XeyucERtYVU739CJNclr8t7gJ1vVe
ldhltO3dxZlor7BBpbaOeD3kIOncyx7hOFA+LRGcLQQi0lIIv8EseXuY0lsMrRfx0xGXRNxJtCQh
EsyIXdmopQD2uQV8NLfps+B2IrmPCIX4wLsX5+u3ZZUAr/23hFsgbVMOrnTH5sZumRa+jDr6+QDS
slViIb6muCyPZF24CJwG1bfCM4bdtXbhUQRUHE7xAdukBs+49MdjwrOwlyiEOFtipOD29mIYZaNH
FM/+ISg+g4z+NLPd8tBLZNw0zKPyEzKH0q5TTV/Oo8b0fXPa1I1p2gpplXKyHaVT3mcVZS8y7MPU
xD1etn8rHhpbngu/SfOfMPWygrm94WzL5t4XVCCmZoKxRlAWft33TUvIM3ncClV29jdtz9X9kz6h
MxashnmaAC0AookqrXTt4MLZ0KqNY1/kDvTE5ogBKy0a8qg2kcdMPmrnxeqHYQCoYtYf48Gwcr8O
rUWJ8F1lTqSKCYYwdbzaHm0kgbZEh83uoqoB7cgZMah+6XQOqO1RKm6N1KrRUvRGMjAThyoz0SyL
UpZrI6x6hzZXbLlXNv8lZ56TJPjYziH9JCvQVyJPuocNq9QUPoWm6+0p5EUBGdjVuyHAhJr9mXKU
n9fKvgfuPRDqgXs783AFYRcKkzgg057KLOh3LR0bBnZCxTHf3MbLWGXiM1KTON+0Hz680UmkpoJv
eABoE2ff7mqeIG7BdsiGIOqrvOJDIIlw+j2g7yAsxU34QfiZPllqzB75zMKINZqezYG/ZdEOtRA3
/e45Ku/OLt7ylSYSk5nkInwghSfolf4pBswWfPJ71xqjuu8Me38rwv6+MG5+U1h+P2uBZBl/ia8s
PQE0IKc1wn/0YC2mi1jmuNQaj6ZteFI51Zs3SGyPapeiv+bW2DfLBVZZu/3vndakwtbnyaEtV8Uq
aVJa5RSMD8jixAqETXsAiTr0ERdoVIP4y+8NXJX/3oH7EQrQDX8Rqiv5HMdoIRNaZOmfMvuYvL4Z
wuBDGiPn60LcIC70kXDwQmhNvfMcYNwEwlI0Oga7fz9JiPaktnHCr/AMf86WUwsd2UXlCKpGJtBq
VOKaL9zNxo9J5E5EbaLzj+2PcBm8c9UxLXHSrLD7Xbk/UgMVO5eF89it5h3wqfR8YHogK+UNdWK1
DfpiXqtFGKXy6+Pydb1mV3MPsG4UkQButciosZGM/YEFxWPwRbrH87G78x/0QB8TmlQkAghyh2cd
KIMLWr6lRQH0fLrGLtKgs9Qc3kcEJBM0vXkD87UgJuassfsgbjjorYctACyrJuoui09H7G9I7DC/
DHXWHtRHy6lPdy0Bx78dwP1VHtaRNOd6kw87jXtxsdGb1iwYU1AKH1LufmjtaYHYzUTkKGMdTPcK
4xqNWWGoxOe2WqtsRUYLZiiuG4pA3oTrWb98zxl7ish4IH8TLalYSYZtrn5OsC+Ny1PVrTQTpBXX
W8CjR8cwmFJ+v4hGkbD1/aA6V1dmGWnlFdBUC5wc+i8w0G31V4HH2ACerP2IYApRUqqhYgrrLg8u
Bqp5bvw9MhWBLpGNi8vXBoWnuRYybf7VVeZqJ1pSA3UJL6DoRalX/tEFF58FlgsHafjL0EJuVgsv
plkhCGmxifcEQ1AZM83Nm1AeYosxCmvimDPM1AuAnM0ytwmDgEeih2fj67NC3yqli3IsMc0PP39u
5/sTqZpz4kZ0t0TnHDhPMllLz9HMMZ3VNMTNmtQWZqd04JUyMNtP016deGm8RAYY4No22b6teVrT
aZ6DZDWWYccrUKnQOQNa1fouN+GOnnFdTVwOtifBpp+DwZQ7K6PDgmCm1F0zyq4lCo/337tbv0+5
097q6niauhR8mYnMlRGqnJNA/n0h3HC3YzmjeWTJXjyzw97a0q1eDh+BEAAGZHFGStnDRyiMWJ6T
QBYYLNnrd45lzT2FG7amyJTKiqbFoLmYz3JmggE0rb+A9c8cUmNaq2raalPkxNtFedhZ8pdKvvng
bj5e26sRkh4Q5d3tpLz19ESIoKS4KbbVyalcLLgc/mL/qoSZpvgNiurXjL0n7h6RsGjSNlvA239q
EF1PLYZCgKWCEGuCA6n8aWPXTJ53QNwvtgnXZRyeWWfrUgXvVLQahy/UqWJAcS3AMCmUEhEXE/Eg
2Dy4P1tkH72mL5vDIEVA/wC8dQvP8FBzR9nEeJX4+Xpgob4QreqnnvagtYwWLiDbTwIgdqWigmmz
4junmyzAZOAJ7RG+aX1AMChRnVHyCZzuEhQxM/NO1d5mZOlyA0HQfYKQf36Q23VMp0pHwR0PIB6s
TMo+w4NEQ1oj0+09OfiyG1asP33WVbbX+XwE7adNZUDfGrgJD9BYpQVucGrzxsQ4kcItLMWnzBRN
GqZ8j8d5kCNufbTJ1IIYT/bKS91f5JZmFKGLPOA2BQUzR1pHpKtC8D1ZdXeppgaXh1bKyayL4TiW
pz+PfcB5YJVV9+6yfqMZNIOoBohC4/3gh6zqRbJWxwH4p3CEtP4azq+PAFDsqtHSBzQsEndwWQSC
t7GeYZdYe004PEbixBhgl6L6hNlYSyJG14buOnY7VsniwW7SWSrIFsuhof/KCOUEl7bitFSMSUIh
pQN33RQGPFG4kdYMXoodXMtILVJ1iOn9xGquMdfTqOh72Iq6asNsnTLMzKV7u2NHRy5fTOzQH1ju
5W3bRVSgK+uPyiWve4P8dIIm++5s34V1FPz6V80LGZbPt2ejo08YGuBD0SMfpN5OTGh/RXK4OlD1
wkqdml61Mp3/JKb/fkr2TkW8FVzIqllYFTZd3yeA7AO2qDUOhIykX/bCtSBnaXrPqUumjTIMHTgj
7ph2YfKYlFy9hrPgn57Nc3o81A5OfTjWWfGccHUg5+DF8FtQYU7chlVqyTqYaM3t5MXnIld4IxxZ
E7TKQT8Mr4VmvYhPZhwTVxkRj82aTYRaEZ+xyzJ6ezGRBtya3/8XXxDJX7BdM5Wr8wX7PI9y7KlS
j4Pa8aKaT6+z0ThWajFyRBnXrUS7xpdTPTnXC1je1PowdECDj6s4cI3VgM7ZUwepublJkQoUjHXQ
/+sHZUTszk006yFg+p99DBQLbq3fDifERzrbKO6h5FNydasp9mBP9m9jDnHOCatrtktiZZi5QBWU
FmAb9JobnA75cymIedjXIZcHncfpZcnEy5RVLo39JVT2qAz48W7TPuuyGjIhWqOBldS+7LZrF2/A
c1p3Cq0ttkr+utY+opfjaMn1illgX3s/qY+Ed8ZPGxChdrxJHz2SQV1aztvXlzzL70M+xjLFF1Dp
fh/EmkscKee9aiRKQoOT9cvW+sQfIhXTgP51cvzE6DmZxJpZm9LNr9AdDuUGaXFXr7oXz4GCMHqn
tYV39GTPnbkn91e3hO17n1hmRbHQD9Kg40ff7SRlifNqStBnUCF5/7NcizXBrkZffbqZdwpRY37t
tEmb6OXZKXJXAsbAHL8VE1txTWHubxR2LEh9/5IODNwH79T4bCyPRzM5aUeR0FbtQeAGFkrOyj4k
AbSO/Z8wjxrh9CjqBBSRtpZfPpuC1oSkTqWUDMlf/hzFfQoXBqguolzxJEBy1CLYjSD06ZCrSBHn
g6WItHwVFji4QWqSsEUQiyDR1ar3iZsoNL2Qv4IglqLbOTOKATZK6qoGdPLsFziREO13FYZXBBuU
+ePJqCz/woJXF6oABmWHLb+NrQEGvcigbkhU9eQ14q4GDEJPIGtkTIIaf5ZMnB2pZWQWqLaYcdAV
BCeavrpyL7uPI7lOWYz3wiao6Ic5cHZUKGbG1kS8IzcHu8pavsAONNsmaZSws/mhaDz/TaehsL80
SYlUPzDVcIMPQJYLdkiJs+kA9jor4bgyDIE1pbN9ublTw064W2Ss7Er4XWZy6XatZKVzhE0ZmIiW
kgnx2lq+PcnfISH9TUGcwpdVfKuwxZ56PSfFm7pE8Ohedpi5NDQmflTmLu7nRoqXRmJaJupEHl87
7WJzKBwmtBGH8C61Uwg9MTkUty1tXGGZbYt891+4S9nf7BuM7WNbCvBeRmI+TqJTvZXJKE6VQ3W4
ymumuEIiB7yptSj1b6w6SnkOtRkyC41AbKBrneXnwnMO6Kd7yk8aXl+sn+pf2Oyl/30NlQhK2Fwu
tdW8kjIg1Q2tbl75cgYuS9e7lFFSik+yaOdotuB5bQRnR2HxovlaGHngTMQ+IFUI/J2/TUAsd0cC
xJAMhKXm+nqpR9Zr8vMXnubPSeIycry/UzexMj0lT4ACxtUPXNcyKlkNY6h6bwtxvhvNODhCUiv+
FXHSz70sdb0dUOmJt/BRrdXVbD99T5shDx917OjdB3QNvfMWtZSEi8nSapvsgTHe9LcFXHqtQuz6
wbAfzGXdB5+A2j1N54vMmRMgGK+MpJUlceNtWfILIdrRfhzDFh/Dv4DMDopDh622UUyFT2q1vclM
F6VhJ8sPOY8zsLBcMkyGIid+XyozD8x6mOdJarpAKhUsWqDXjhCKM4XNZo+KaIZOZ7O+3qsSzLwa
TbWBR46YtOQBu5xNanLxSeTtgPPe0/GBDX+BRT3a+juDFc7Nq2aNxFRdLec7edBsjl8lRN6wTI2A
gF711Dv292Mryd3POYV9au0qxn07OCRSqC/AYOS/QDei47RhPNPcM315x3xNMDXiG+pvsbyb9lYT
fqYDe0kUAq8fqmlTQSWE5FqoiXYSYq/s4czh/Jn6vNidjjhCCRCs0nzRt1oHWUse4aDPKl0Gd/7P
N5Chd1OdG4fAyPHnUSXYfOqxIEtvlnhsy5WS82hcQQXzsczSyg71tTlQ4/UFE/NU8SfhZA0nboN8
Mx1Le+nwcWKvA0TAsFa7N5lGULgnQfTpW0/KPq8cPsOozjtzruoBZyYjlD28Q9w+T8SVEIe1j0V/
7pn2njNu2vCE9E2uL4fhbRNHXkWVM6mt5acJt2bovhN7UULgXrMyBqdV8FspDlMdPFZrQK3cFvAL
dU6/iPxlbr5yqmE2FKoBs+7RSK+EAVOLV12+UdfgrhVX0kPDvY/XfeKqEoognmVFSbmuh/+MARxv
MwUJzQ+LmvKd3zkzaWw1xxmtcu8fxMjtm+r8DCgtY9kWKZ3k9SR+rF+jPVnDDKE89hCLFA/BZWJJ
JS0EV6AYFXsaS3gtOjowQyoJ9cvZnnITlvLPERu6iXhz/Zt0aaxvySBA5rTPt8UAWpxSzDgAGo9r
/FXY3vmc/q9lmLpazGXolF1vtY9ziEamTKLgu3x7YDiffRdFZaUbL5Yy6r3eVNM3GBvzaM+J54HG
ChJ68zErsHymkEAmO0CAQtgyrPxF5a4GqjUIeBX+Oa2U5i2T2nIr7gmzudq94yu48+LkCoVJ/eVY
UvNKNKgW274fdt+ou2i9qSPTfBIO+Bd221vKV0dIXcomnBKDGzPEUtjxty3/eYLOqTsE+0FUgvyd
1Z5Jl9JnrT0/MXdBmTHfkUN3uva3/OWKl2n/wqQm3Mt5WrwPsz3ZTMnKwot+SMTZHP4LZJIb+gYY
6UnIhYniG2aenEwPI7tSfLH/fD/IUkpo3MEW39En86t6UGPK3SlMN5gYIYgUyzeNQUm+WrG4YADo
Kk30tdYK8nv6z3edXYfpSXbXGcJRId4mGyR+sREsaV6SkFvB1TXoVT5u7UdZ0segSPkkc7RGZiL7
BiSw3Xu0qQY3znVykd3KtCzDtdYxfmIsQiwKLCpGKLBz305hjAki0ZWteFBwY1dRmt9tEy7OfUtt
TpxMSuTcI/ayEceG22OPX3XsEdZ1HhHc4Ku201XwpsmlvYV4iJ/tKJrWm26fqWjvuYSeU2wSaElU
2Vhexjs5aK5uriyyM3RZd4tI7Mv/D5UMA11lP62xAmqr0VUdMyyu7/mb6D3yicF5Zu5sQ9LKTTeO
wTqzenzno0vODip2D9svVT12oX5FkKe25GpAjgBDo1RqQ8Q47wcS9PTzV0iFZxuNofB71zjmI/Zh
LR+RPHrKbWmRKaAEjqrakA0aQSMTB0oH4JLRyuH+Z6ElTvilIzFSQksmAnKwlYT9d5Ccuq/I30Ui
EpXvh4aizNl/SDRm575HrzG663axqmF7/KRqgFMbw9FiTgE4hFjmeMy88donYT/HXjqa4mdK4+Ek
ih78u/qHWWxaA57/KyLlKPeUCc/3xy/ib9pDglmZ8Y2ZfjURxjjwrjLiMxhoKzZOWYTETOY9OVZJ
URiRGPeMGSk+cnH8e7DqSLxcuK1Hk1lcG1WfHRNTn5YmUfJcGXTdPMCNuNGNnBEB4tlhfsuoQUkh
Cw2PcC738goAGHkauyx6hXDL698KbEWDwo+MxU3Al2q5/ZWO2adG34y9gaPTj10NUsNo4n/hKY2C
3j7O5dXc6AvWVVnuJgHkBSxym2a73XbVivbsNpHldjgtJEOgI6tWoBPVxjMgkVkPEbwZQkfaL/Ht
JLqbAU7+LGVafa2mjYkMV8qYUVbMUAPCxkfuSti/C+rd2TcZflGlb7XFkaVPnvSQFTRgJext7Y5e
LN0mvjIZwVr5gRV9lVgLzXN5lU5YYMiRlzMTf8aX/PiO91aCwfPtzhju8S1B16Ips1R8ZUMblfa9
BrO/8OCgXL/pgr3AePajocOGtxH1GyY+jJK2e8KlqZCnfhhb2Mg9XgeTHqAuMEwAIMjerFFyHHTn
TgcPQulTVX9RLl6g54fXMTMGOI1zPV3K5DZhrNONtOeqRl6LA15Fwx0nY/Owlv/W+Db53FVsI8Wo
YSff80n02q2ViaGA3Z+57UKX82ktl+o7bXFY6xQLZN1jeJ/2E1AEkcdB6LvhEhqbonAyLtC4/Hlv
mbdfKNBXNsynEshyuQYeEqSIiEEjS2VEgf03vgySXVqniFfhbInfix592hxPY1PU0EVAgO4R6YRc
2bb/A4tftNWxW8u52LIbU4yC4DqpnWKyrancq3ywoehYIXBxPZVIjBncfiqPommgoL92ZfzrSOPS
80fHQAONwURJyr1fckCBBqq8BBcxrxvUD5bYWshljQ0DrOMOYVU0NI2pmcB76rT9DS4A5Kc2GVUy
xKrPGypw0BJGpKT8lJRVY0RKlE6nT3gRmsW5Mlol246gvcdDlTwAV9MiRSPGAYcsSHabrHckaSkX
kcg1GkkvK78uVOLW2fm5Ct4BEhFljuffd6UrMKfYjUlYfKVcgg+ZI9MPa/PCNO10hatGo/dag5xC
4CWAeFgbmnkOb5y5iOPQkJ9qwNCdLUatagxLnI3NMs1JrkVQhZNHzw1bvKptVyZiJOV9JjUlNhn1
0/53Fl2QxkQOEwS47VttqnQx2kTNYZdq7+fJ6jSSibf/GGrdRh7KL8VoeDGvMoE6rdtd+akuc9d0
6ri2LYMAZ0J5v0ee924Pwi42sLgltyB+7jYaMj/2S7+zrYf2Bz0UtwqYdKPDxF+MJaIj+J5Yf24q
HI++A0vlNcaYCAyBHiWhlmR5awsateUUcB94PAA5P7tRXEOPASrZC/qO1HOTkd5SqevK5E5C1+WT
nYFNWoyGnh5FFPGpaXbVHEg7F4xYhUJM7mfSViz1iPyKFE0vfkp+y3i4qEXdFRDBD55Rmrf4dA6z
hnrlRdEz3kIgK1zFY6ATuSYNqyvrEJQA6hPWE71VvzIODorM+0bZ1TeBp2vj4cmawdKULj22+r7b
zR8D5aubLUOCxZqe9IdStv8WqOF0gfH/k0GnW98TWC3VFxOWhifDHCDwbm1weo6TfwkvDG7uEjLA
5MAb/tXdolwOgO85bcniQmO8yUfBOSBRUhK43GFfKLkRsgk+9EkVOaJROOvEQ2sNkXWYz0rBsl7q
4/jpvMxoG7GGDRAdK3SLnNkRmFouQ8ogOgJppVa+XbiCAPs3MRK06JPmzq9icSHBC5GzpSOJoLk+
KjPPck6RKgWpTUIGzj6G2HqOvve30l2kGj7pqYdiRk2MWF8w/0J/08ng2weQC6kp9ytHgewOOXv+
Fee5DAjetjIksUTxTCY+frc8Uvu5yaijKSc5f6DNhsr0gUVDSPixiZsZdEy2dCC0Y3vTcOSC42tK
eTlH+3EIMOUzt54TLcYlWmJtSxMZvJ7mLwEGSuC/mDlKPqBxwGUnht8Ynkz9es2qjcZHISI7+zjy
O0u6y1mgObYRF1OPV9hr5iwmRdsFi5iprOR9OBnwEj0ImYbRvZBe82QJYgNBkZxD0fmKA0S6HM8g
B4YMM2snG7QYskSmbSB57xitUhvuBew1S2Dw2LQyUlEIW+i6BQNgF12Y4jhKpr5taxAijzDO6lNE
YSJYiaEdCNGQmzEK/kJarRUBDSSZGu5gNgb5pqMqt5KpnFD/5Jz+Ttt3/Wk7F55oStlq5eXJEA1H
hhqxYyDT7rmvzAXJOnO3iY33qDyRb9WTnkM4qm2GJjDLNKe+yVzYd9D+gK2McupsYUGeGbiFxCl6
8I8qGhvyLYGqjLiUGdvzwwxRZHX4MdXwDeotYcIrm3fi1a64wo8SOrztbYPnheONF8wDfdlldAMS
owpPrHv/2/tFws4unoqxI7apH2voPtmWL3eUNaxyX9OfiFFYVatYisZTChabjPIu8vP46Tu7Jok0
6mWVBYvg446hYlRRg3/6fn5o44rMqh5sY4W7XEf+iOwE+sVLzX0nDqWYNwzcG+ZLa+8WTmv5xoRQ
ROsdZn2Cj0HEgL2vkRrvnScElWcGDOkQWYICpVY+OBAxDmWJP35usEJdEBD6edXACCQJBiZcuJS+
rbsu+E3lagDsQLHtsx3OUpBNVbpZwR05xZpDzt8czP/FpHm1/fE83OwHW6rSF5ZPf57P1+pTY7BN
Jd0csVsVHlCgBTj2N7FZ9bSKTl+DSmsRAujDUPjmyHF6kR1LUaKKcvOVSPXjjIZawpY7EMXGmjLG
s+llBY7UZuSPxNDtuzsgJnuBav2tYpE0v9G0oAAz+2LJLAawAYb7mjVj+XKbyiTN1/m2KXJsWG9b
eBeOoV0yh7YRBu3F2gtUNjjq70aC900PaE8OZiR/MJhp8dcSamgCUxcQHp4zD8UuLrI56AEJpNNH
r1fCx3WtWiq8QneJYeVDZ51C0KnTPhtKpiGlp3IUIyAiXlHMMYbMcPiRzr6eUmqKUYuiaqixCpfU
ebc+X6nQFvZiy/vzWB4CEW2Mu+QQ6moixgXsLOf2dB1z/+TLUS8pYAiviUo4lKJXqLa9JoHgtv5j
0OGEWe3F8+2TJyXKP6MenK365YmKGu/CnpW+UflLur9QObYyfGxB9/ZctzohLlEqet4iWvPi58L/
DdpecJ3frB9GdDP3iTlWL9o5jkVKx2wVV6tRN5sCTTU7iBkBB9qr014PNB2CZ2TcSRJIxEi/YpDG
5rv7JSxLyBKsd/xCV991EvDseoUsVy9HOEdz+iTMG1skPtW9kJ0xvDkVcLooY3QMoC6a2rmtXFKO
/htotPC0zwuxomw6a6U2eLNoGZ9jZuQyRXz0dX1vrwF4ga2hxeo3vEef4O41HqZG/wJtHr95zS9T
kSjLo3zl8OJ6Smbjmamga2YUOyku6T7+WZ9SqRBaVuzwNYkIXQFHV1Lz7Kn6esBImD8FnfuWoYUT
uy633MbD/qajs5I6it+j0xdGjLXRoApFXjLDMnin5356rJOEKo/Tq4sOrEJw3j+NRLDZs8SAqf15
bijWue/wDgNRSb69WofTuxsyaSF48zPvoHLNShpzA+YTOP/KjrKvOTusbYwmfIXyhmWyRebUbvTJ
00VlxS24XmQZ+IwYqKRTKJ9QHRdbZ1Ii0LsOyznKakDMmFiMOB0A4D8WErmg+AXZRXBjvznj6PDZ
cCvG9rsXAZVvdpMoqHJ3JZstTwbR6YT+0MTH2efsXTtDBeyezP+2tc5TruscAAbpu/qLiVXQkeCA
YoKYoSWdvW3s55pBbX4MMv+1z6vDmxZ28ED45W9lwtwWoytqXC0i6+A1eG//iGWEY+JZ04qouhoj
+AX68cMrhxM4t8jzgaui6KlAz3Qs0JrldY5WkyL2pY9mPweAqEQDmN2sIzAiln25dKFbYnOR7vtP
ScHo1mPxpABSlum+6eGznaDXRdTx1gqBq74TB7MYUyFNwxi9T0JDZ/tPcd+LEi+9L6NcYKzOBV01
MPydxKs/klhG+UHIj4cireIl7gcdUeuoK5+JmwkSdhp8L32wCQbM1w+eASrDffjQDM/C3rSkfBzf
BZqmQPCaa4sY67uDpq4M78Gy8W9fKa1B3GlEf5fRHbSO/fSVqjJ/5UUexe4tEfjPAtJG+FLamR8e
ORA7JaioxvIwfQA7XCoJ4eRgoBKvhiBe/Jqopr//1B83DBjndX0bSFFKCGwUrvYEUHI+I1GYg+iS
kivqa7xoME8MRkL7gOJPGzGw3Xe/BA4vAzaTv8lMwopvEO4+lh1uNcA+zu6oRRjyW2Lu3dTbd2kG
iijZYNt+ky1EBXOWShAuyASjXPBrez3Ew77t62PaATHFU6q1cw3iM4GapzD4C5DhUkQSCOu9AZ1A
8AnAH+bgSCslizeG5C562mJA+2TC7/KCjzrcdeBGmZJtH5mazuJ08sMunYSDw4oUH1G1HTKoG4yL
wZfAebJWPetcM8XSOH3hnkGWe65d1O+TyDFXibIoeBZszY3f3XsMcTBqvD2Bbpytwabwvw+vdCgU
dSOs8iGv0gtJweg235fQDg99irFt6/mouEablI2rtGdeyhJCY/iH2kdxDPygVs+Irk8QCBfOeh+B
14DLnzPoDB7gWb3h0COMsr73aExCnfp+wHJ5Bii6UXFKWooJBwjMl6X0fH7ariMZa6620huvfFtR
aX8iVXvtdWIlM9DNq1GMgD+lGtjo47btiwCocv2FGCsl6yezp3qbdYum6dIkC+2VAy1WPXlvXE2p
bcwG/o5S2YRMVHZm0mhKb9EFEEtPMy8sybMPVqL+Bk84UPL3l0Jd1IOA7gVu+9sLjH0nFoP64cj7
If6HTt5ljFbpDSihXIJo3cckXcO99p2g7XiwgL0fFQFVQ0mX9utLf3fX/+oWvuRX1Kjk1pYO523o
014sY4tHEYDb3nvsKah2G3NNRvcL20pLwT3FK9e8StlYTCEUEij8j13ja4HSOdsvOW74mJMe52A7
mrsimMry90VfESNtJ+ltyKzWowuQTv27XHkAcVW9lW/5gCq1jwKXXjcgMEqm33m11qiLxrhjgans
+ia+OpZ5B7iMFaLljsHFzIu4QPnRCz/uZhYfin4JPOvKLmjfStV6Iyz0oSNMn1AtwFu4x7uxq40b
azbexGpMs/gtXbM8Nnod4LwPeojhQRQ4HYfpN6m5Qi9NrlXOeL35f+2EpZzW9o3jkTX/qWH9t5Ig
MGUPJjO/YNcBAfM3QBeCd4q1hUZgSUP4s+vI9+sfduJ0sAw8qninJpiTB5vjy9SvZ+Zjz365OBMc
otdQ/He9SeYIUzX7uBz10xU7i/1ly8omhEAaNduS7/F5wahGLawY19jP+IezdFkTiRSNEU/sl4z/
Onnrd+QvITO5As4ELuMUFmGUftgLX9EH//ypyoHSZmUzmP7LSMDMb/JBYLv0bjNs7ZxuJdCq/E0+
PRHYLJne81TO9LXXqItixl891+OfXexl2PdX//kkSan5FSkPhbWCG7KtcLYNXDfnUtwliqyzyy0S
NFs9NBatyBLpVtF/mD3mWWGvJ9gu6BbWgu+Pt8V5WY9qhoZfm/pQZxtRHQEVTYLwLo6gal2hoLSX
TEcDAvko4YvotsuZNXwgJFWwooJ3Up/uth7GkymMxBwvbU+idV8hgJCx+sVbCsKyJB3RFKmDQ48j
5ErTzqsDNzXAkhc4HEsSW2PxhwPcp/ue/uA+qGqdvO85pb+l9awsxUuqiTmU9VDPCGxr+iSpfYBT
hnFctVwq6P/S3g+rKzLjF+2bQh/rpBrmVO0dAdj0F4h+6DM0WWOyP3qjT6n2RigZ+pJ2gfBMNow0
+u78ICCOCZTEylnSXrJ3Tw4da3zK/dvOk8VgVA8veahSwyu/60hEEMitw4+88mcNXqNG6WrzxFHl
XbKgwk1bjF4PMdBfVZWSnLipra6dy5X51x1mvETS4Adhvcynd6K22qZR/N2JqX7Nos5DL37I6znS
wbgeQjhVYKwdzYcIPLDopbuB/CyNS2nj2oBL8gHSv0tXZelg/SYNKQK3Gg8dFCFOrorjalci/ipA
Rj1E026HfPhXm8RQruKW0iUtzV1ocS6HlDbh9wpcxnyjlTeziT1Wl16hKaS//GwOh5Ub/5AgaUB0
bDGdR2Xvm173B0qa/p9ns/j/ZiILSnqverta/01v3lHCBhLsUFAv9a/0PBB3ZxwUMaU7A6lrw9ik
wzl37UQxD/PqYDEF2QUkK2aMNI1kM9wc7G3KItl2AVcXYcAaNqF0s4b7QEywP4L1NCUpUpF/Erft
XWLDzc9eMye4m/2N06EovsQCzQ6W4w8e+6g0bSRn19QpS8pUfMlM60CexCoasrjD18eReaheIzoc
OleqfluGAHGebwXr8EzBzxMp5wxPIAFfNdOuYB0SJNwN1QMk6X4MafG0fULfb5n3OJ1ZHtSj6qRS
wQ2NVV/avQMoFb1xqCHoy5cK8IDX+uzgdRdRIPfQdXsT6CTPMjoCS2K8aiCwJh/gEiHmkZwYz3QL
p0mjHfOymQ3RjqHvj5+pRslXWM8CJlfK++qYbMHwj5LjzGqKe1p+KytmiG3+dBSJLy5g0ODk8xNM
IOsnyDNgsDQBMo0JUwv3KeOubuuW/jjREmvbQd8g6RdVLBRRnkdQtY1oiG5YIs5VPG4ggCqwEdC7
cvQw74sb12vAl26LR9GqK3B2hhKxbiy0IBZfgN776tnznrqCXQzXoMmQHGnduGFket/nhtFPjTH1
TUrum+QX/iYSLGXiwi+1JPbPLRKdlNekJzG4VusEZrIcHzLYcZ7Xk+hxKhQfNVhn11JAXtX33XhZ
66IrXHHaqts+I1b0kwYQqSAZ+duWTNKz/AksIwSwL4F+YsDFUpJJKvZmQ3QOE0JFvZXBnBF7hiSX
jYQvnCPSra/M8Rc2TLbpWxBfMFRAgzwalxesxCXDko2kXpZ9yy3e7Uo5R2tH5cWkmNFxEpm/IySf
Bc64DPO6+T2IwXqTyJdtjPsCRBa6/pmgvIFSFkWRhvGofHW6SUyc6vivPlVPNkcodtOZcVmIQXPz
N9IO2eWxbJx6ikRnue8GX3L+faf2nH62NT0M2T6c52eI14A3vnTSULd9ngMiXxUWWzcjxZgz26kI
2DDZIst4euASKVE2nyzuqcDMoViqETd8ed1deu5zuCtsJYZQ3CC2TkNzA4ChSNuvjgkY/1I11jj8
8RiQk0NLQunlvB7trvKfRpRvvL1GmN9b4Oyqp0jfy1xoE+rn7sHBGqlqy52Itod+AOJ7OcMzEUMO
/zsdviqBmhXR1cY01N+6H8ZnArYeW4Ew8Spo4mWeGcbQojnGUEu9XG88GvLJ+bCvFFStIhFSbI3O
EBua0V2rmwnd43txQ6AclkCt12MNGK/HR+/BdqPr8Dvx7dpY5HAmEHV39N3E30s3OFcF2zTl++FV
9Dg7+pg3FuwOmrVcEw/729GWN93PgZoXNevFp0dG/xLWT2EXNCAU7spDieeArHYmxbEQM/yFBVic
yhMh6g4eXi+6nkJLCWe4h2S1bRVrHzKYGfcvcsVnJfojOiASiPTLLU0Zy2hHYxWpCwjt3imZJACl
SqDO59qavzIktBzXrd65uLQn4uj+pZAl4dB5LcbnfL8/UWO0xdezlL87veX/+wTfknT3faR+NgSt
SgLyunb0jFMNmnwgX5i12tdeBIG4N4BtFq/AMuHAeWbn6V1zmk04wXqEKJpYpdo1fWhPrxtrZgQk
fJ4/O9u5furJXYVk4YNlxqAqj+8otLoW8pGBKMl1CoRwqHUVLEtZ+C+X9DQ9ilfXznt+jUOjSvHW
NgWAO9Hapr9q51EPzbC+fkEJ++MmdBtb+6nOlFwcr6EtF6bdb6CY0zX5V1llGCMgu3LTpIxn6Iv9
/pWb9cWHa8da7dPMlt1fjTYynG/c8aZJEfgEMfXv6GqOwuspY4KojQMst0gkaxIz/eua5PGhm4c8
11egksIlXRXUsBLnbGI7QVZXrWkVVPyDersHjpHFV6yzNBGv/Kr6PzlNTANFOvXvFg8we/N5/Cpm
HZF/hk8S7aeEN2R79OohxSB0mpARIkQZI+5d/dMv/NOUYtx751P5cQtEoyA5we9LCuhzJoEogbgn
b/wRnZI19L5WMmM57EYWAwO7SHBfR0DA+bOdrypMnSh8u4ha40KLEfnaytmuvbUgYlmEGe82E5Hs
vrT8RIWUuCYqhkAH6EHksNt3Pbx2eVWNOKF7Oe3Wx40t9im06XtkOKFYZ4UmzFKAn+oFg/xfAmgF
wlxWszvQnpFbN0VcIXxE4gQR29DvExicLcIjs1aB6LdFMz7ls3F5+DJ7hkhQMdRWRwZTt4gQcAlO
+Sqmxor6SGNMoVlZm695N13IT0log5Mm4/KHpgQbhaZc9hsslz8ysC5QuF0AAjBMcBamYwf7vj4e
OJSmzRZm4lrZ8nunmw1HidH3owvHHEGnezHiCGjzW/hhnYriUVqHTev5iiZk7ypYGSycK+Sg9LcM
N/yg1RgvMeLRfTkaXFBXLLuVn+AqNJPmoivmvYaih8n+xHLPyWoX3q7xihQXDkaw8O4EvLALyDPr
L2+3q+VrA/PfcK0y7/buJvPV4SMw2sj78NZDAOSolNSM9tX96nmvuRPQQOWp3qFVJYDgwRlrxpEz
xkc4jKnATLt40PURSrRnAozG5ovlbiLGF56FXIhg2aEWRd2BH1jhWWGUp6f9CorDAkx9yYSlxAVv
3K46eqVd8+G+IFuZkLgYHoXpphlP/LUkHf4qFsFdxWviGw3epv+qUJeAsphWEdCm8cWVMEpP5knK
XSw/sBMTioBkuYg0hhOnKJLKrDy1Pp+dNy3Sofbzu/Zi/2JOenmZ2sqE0etAo05BPHJC60qcfK+I
I/aN5F6UKwk/XYorIxAHH8RFALaO5ZhrcHk1xMpSVlT4oJZwF4tbVLwTd5vcoSEByFpH6n/eahBm
LQWI3KQpPQyMJgmeWoYY7gmz5LRhL1iACpKMOsQtnA2w8xcUO4jHkZAQ4AFjkQhUNgnWGQ3C8Rlx
spFRAkylapHFf8c2tdPihduUACI8v6RfJAorhVCu2bBn2kN27hYcKqpLMQ4iP7At2OTre4BZFENc
kNAeMFX/2Vyj9bg+fE3LuAg8ft3nKF4Y2QCqnC/GR4vN5mv+W3VA4iw3ynygR+Uyiv3L23UcGY4G
4dR0e27dULR9x2YxRzNYICgK9C9iAZKTB+kvkootBxm5On+5A+tMOXpLibdKv1FPheZFpzt/Cwap
Z6k0L/GJfgaLY5Pu3sIaQKxtNHRCAZs4b74GDjY15RvNnxJb3olB6RZ7HPeUaklPThLHHMmoZrv8
kpuomEE4lkaB/sTszLMtcB0gxgWmeO5wgCvjBjIvtSF2Cg9MFmSO4YJ+Hx0hxBLI1uXHUPaNJoev
9/mmAWpotmROrSyDLuuQDj03SDlc0MLLWSgHazcUws2J7ijnCdJ4Xm/2fwkrkS5aP0dxwITlylj3
J9aG26s8I52ReJS32boYNy2J1AP5uh/CHV/4+cYndB5UoFxQ0IP2xTqriazOONq8JX/rptVtBTRR
flnE/yu72a4+zEBT6eaM/ksNpZxzVFr4SM1j0kS+LxJsNJGKGrwNgtTBZvVNR6rHaaHTY/xQsqc8
Lj7CCx1qYXIEUGVpAaMDlLqybjTgBkp8ELZ7nhImepfYNiePI9mO9pYfy0X7hAJfICrrzb1UWdx3
9aVfqJtL9zTu5f/C/ddCaowdZrBtudqdNm4gFgN1d+vWiBiopwDnEJ3uvIn1LjXB5qkoeS5mGDr2
XtjUKG/iv1kVVPinQJcfSRu5dPa1B6CsU9JCU3WBSCDZlfMXuCZN9exg85TuFBFdqXClI9XhLYUv
w0vChmUiPQKBO1XRqZpl+4wAgbTpatB+sPfzsJ8KpRmt2TnW3K8GLKzmm+blDmlXU8K7Y32CfL4a
DWhidWKIjniWjMTwQMf3b6LgkJbLOHc6I92d+ZZErj0vbP+E+2HMP7zeWlchP3CT5DPJ/0wLEgFy
dWBBkHBHVc7g7OlHUNQbGQnQMu+JG/VIRsifDp3zefWV1nCdAI59XxsGTuPuV4xjbxMTf1vgEIIJ
SnNXD4k1tfuVJ4ILzGXpuaWOP2p0zlV1bkCf+9QVBwD3QXwjj4jnH47VF2WuvbVF0jpFOTjwTBGG
N+HrkbadchBFUhILuHVqA+x946ku4vd4+GinDQ0PM5vHhc0S+gjs3u2yQOHbuJfrIvp1HYLOYTXa
5r1A0ufSNHK5rTQ2mB18GAFT7Icc1spXckgL0RoUb9ogzsXCb4V0iFEbz0N7nOCjoojTDVmCnjwD
EhWdew1gbMi5Sr1olF3OA2u9NE+rAh78XWA6k8q9tLi1CM0R1u31PDsVU8HsKGpJ8x83KjM3j+t6
60OmoCb7s3+tGdLPl1IX0Rf5VZC/NHA5xvLw9GdI+zd2A/3gVV8wMqin/3rl4gZKIMMPsGhxs+v0
eQ1sScC93f5r4brmj+NOoCb1pus+2OwLaxe+VyTQqoeyKR8UxOuD1yH+U7KoR7wvdsraNTKPgF0l
iSNZhMex/Ebvh3ijQdSu0uSSGdRo0+5gibiysNnK2y7zDLDbVp+YG3I+uF8hVHI/U9M7UwX6OU9E
OsGzDW/EFkuz3gG4eAxMjxs/7jr8Fe58BsgnRUmWglsZsoKXhlU9ihnLyRXuQVw8Sax/EeWi2uJJ
0gdnpneD+59P0BZ/8YntUa6oA7VoRWnzVrHExZvNqLhRG6MpRgs+dYMG530opvtqs9WvMmlNsIkA
s5N6e/z09V1JtJFBY/8T3NcvCAsHBHMg+MBYFGzBiZVz6rl8rTgNPWpFlulBLWhmPa8PBdA9HlBz
lFSdCLe3fb2f3sPgWpekp/Lx42ABwn6E5F31lhwUrp/BNXpHHDSRK/hNZhNXCeCiyNpaY5NJ3I1s
MLinEA3hbgS3cMcx2RN5bYK6xFIObDbzoUQ/cR+JsPSdan9vAKov2TGFl3Y3qwoA/AYXCXi+c+h+
hVFx436hmrIjZMz1HMncSxqJ5Q9W3D5pkbnmV5mHbPQMiXu+C1/I1HSnqdCgAOo+wYuVkB2LCI+o
c1+TXeO9a/5UBIzfpXFM/A5JbhQpPemhgT7DfRn0z4PYBC807UNpp2GzUKb9GFvy2npdIUjgK4im
8gtih/xFt9u3ZaYXcjpuXbClvGk3I6TLC1Az/vguCsAhMFg4iORss/KT0Cu2N91q3LMvc3CEmeUJ
CLe9yXuurvg3MQ8p381/HeO/AikC0Noy3wglqSuf33ZHy+SuQK1m0tVxd+NKgdluGY71wZbGVHou
C2ZsWFK0xRULhc9HvemnhTHUo5DAmsF9Lm/iMN0K02iMDj8x8GJ1iSgY8C4TQvaOjjmBYDzzOSJ/
jfQl3+al2XecwQZcWlQqFCPvKY5Z5T+t2S+Tp55tjUvlLQkOY+WqgUl2GOlq0nki3310e+SM+V5s
1iTtDP0Q41lZasYhQQWLa1mqeiz9Rm/DyEmNcXsH8hvDoVNCiNuCLRoa55QqA9nc7ZfEtXp2hEli
QUEtYJzVwN3jOhrnPSmXq5j3M6QG6XRqKBCMP5QptTmrnDjUCICxP6GNAF0z9gqtfkdXfZsszmUg
VrhASf3Z7hdqHao7syUOTH5Lcy8834DOfoUEXvRiRQkxoKPZr6Tazb7XwpdchRFEcXMTgrMaiI0K
TaNwttmhs4W70+GBZLwxzEe6OqgXqyYWLUQ/forohAb1nCJyd5m7pf9WLybQvJPvSlshyuLynXmP
dS9PuSVcbKl5hVWmwHQBI0AT01O1tn585rGama6k56KjBUlTynL5jYxnXb5oqSFLAXC7PiINB6/Z
RaOzKMxp1txr8tRE5NwdrUCqELl4fnBnA60CgGfjblZX39IkbSMr3HzxA47ARqDYSnz3egVsLylq
FutYTvwZ0VfyuQw5raQXq8uvQ1e0qingXV90uNREaBap4qRFR5Mw9VPOb4yZ1MfJD3IOdX/xlPIz
8w1XLOFGooW0hU+8736EJuHvJX5MglpjAn1EZjoC31QOFXLpG0xu+LzjB3KvTJlwpFp0z5w2mF9K
fyDOj65IsnRECexKo8+6XPTEpn+Uj/+c4VNEI6+4vVheqceieWIz05fV0KlA8Yfn+f/b8gzz7VQa
MLpASMYhHB9aVcaDpIAJyH4OSANW8nRzpDm49Pv6AIwEnQYMt6fbjgzFD4ljepXjUPQF4Z/bSSDj
7EXiUKJFXGYZtLMvROUQdsRjRXrql8GlEBoCloI1v1E1+YOqAaO13T64WiCyhUXatw+52B+TS9Op
G0+4CHlLZ6FkF1xYQ5fmG05rkNtoR3FLOtQk3+rFa6hVhXqBufpDJ1hQYStZjLILHy7zqo6jBHjJ
qpUhJve+k92ozF9jt9PL9bb9r0sJ1vDMNp3Xb6gqkEnbUPJg98w7Vge1zz3pC/W4k9YgI88cXvk6
k9Yn22bFi+rVkmSd7zmfUWrBWEJJgpYtkwuSsPZCVG6a7gEHeqgQbP/0XKG6aZivYBlQjln1I5C5
pB3Ja6YGW+9/NbeDlgmGKtB8HKzEYjDfqKGpBMvjtH0QhqdK0JhlMc2oLQZXfPpgZn/NzgfaDmyk
FZpV5Hh4EJ/QtxxhXI8Wk7789FUQnpAmSeG+UDmZ2l8I0pRnQKLgv3jvYwdcxp8Xh15v4rcMbPLq
QiU6E7rKI3OI+ZlaAzY050B0jAKfqhQrAgZoEnaL0ytBzfjuKViP515PBcWzgtpyzPY9xE5bp5rk
ZVRACDHitgY0bQgdv5LC9NXwy+c4HMPXrk17hbrV5fHw4D49WpQCIsT5nKiC5OkYToXMpMAq6FV3
ule7wX/QC+zEzXsGrV/Pxql7lOC3WsV4U0d2uNusvqzNqQWkgaRzwJLOAq0DrKvFusgN6F9++qRs
yBEMysjZctqKQx6jpIpz1XMNKkDWLtM3TcrGAkodVDRmJah0O48QMxtjoamTxjc7FFXBtklDYXCD
n3bmrMCLsPKhnnjvSyLTVEcXm3n4jA9eF39Rbq0VnwjjMSoFDI6xFANFgFDNoe+qOA6DixMGXnoP
VnvaWHm/NolK8UiZCHv0YM80pPZVi8Um4Yv7jXJdE6vhzT01vlP9yXtZEBV5ZyXF/XtKSVjn+6Kr
SV6jKZqmSD666XLPp52y1qvga0Y5/7NDeSTzCh/OFSbdta/iD7/nevSRzcE5WNApNTlAAuresK2F
AlFWT6gmx+fsnyPru2LiiOunGqsvUmMq7MCpJkAP4wgNSUdC79DWZPvSB8LWM7xZVcf1ZHEUVRJG
ItXYZaAPBRiYiIPKAbrkj2ZTHFdcvnnPiGuO8DpPeOOKtuOt+wkLonOJUfStE54KkoXYDg4X9FaL
pckkSkAzF3+I/TqHKGIeXffeopzn4djN1oDb1JOhBianzB4a2BY3DI412tcS2TI668FE71b0n6e8
TTxZINbBVCZOsgB81dyh8nILg4JU9RTRIdwB7quBEPXpC2063YfzF0chcpG2YjUxM8uaiZhZgCGE
gDNVjiNmxtORbeUyHVowDXBBFc0D9U7aBKrS+RH9Bx9nCCnNkAk5vlbhmxaBdMS8JKjfTyGaf/lX
Yc9Pmo8nU3smj8VdbpFQiFEKGSqnrqy6/ZCK+7ZnnMHKUqmkLbBFQ3FYewQS5wWpNZWyGrSWEuz4
WO9IkqTJRRf1oDFnVR9yiLX0VRXK7dF0TIk/bVKVM9iStLpjhdJnFzWgSzRAM+r4TRZnXyvaZyb0
mbmVLl7NhJ2WbZ39n5FaRG5E/RzcquWBcxnXcb0jd62gc2tpSA4606x61ULBJyg7IXUzdkXp4PPs
risliH6L9wcg0AITjBuzjfOKTtDn+uwCkm0nbmaASFYH5qCWmo+UN8LddJoDVwPOQnONuwTlvomi
FrNGkLtZbCcjXFsiyk+rYjhx4vtG9G5QfhR23776VxBDLXmNULGM9auNu3AuTeW2G94u7Zx98Ejt
d+FEhJ3HJ2MchEkcun2aHAh7xqHZggMqBDRxVF4MbP7yWXsT2zcAWnJEQyEZ7dpEmGoQqpQFR5C8
fFCNz7DpaHwGt2wkrPc4ftnrV3AQV79nlV2RkcMLQd3EA+pLKODdf/0AjSWkYjMe02796+E5SGbG
lLUwqiBzpaZ5aTLXBhIVXfJu3IZjjHIuixSsngk8+O1ux9kzLdo8omxx2epdTx2wAUsubuZ50BnR
UBNFov/xYDyuYxOZ1b30edFTC4IiIL/8x2iBx6EeJ3yj20fwf1e1uvaA6ozmVJM10wSOJB0qoxTz
bx/Q5MTU96yeGK8t0DvN1o6bclXsjBozHi72dzRPxDaZlzBNIw5Y3fwFsqqeGJgQjRsvB7Xw836f
u6njizGLpvwiiGAGPu+xon61MmXjIaS0Fyc5vPd0fAdnIcFLYBS0PuBmL/O+BluWnvwmAIvl2q8v
iUb6BWu8LuV2GXZ5f70nn6dXjtLcVhJKEhRATQMDV8KmR77VpKzCSFy2KzfJro3jsDKL8poDQmV+
6A40gf5bz0hjH49eMErxdnORBBitOFvrqPAT2b/ArZdMn3RrlKsgVeEggP9zN2lnDSBuec0QZLS3
+HvrvHVIUNq5nJ4ACeksdN+xVgrG8rc0dN02i4ScHKZo0TaDsrWT4sJqF5mKiApRAVWgezo9rMlY
ATw5zMliY2U5O8dC1gFFDehODtgLwywpCXEPYfJeu01omoRSq/KosJb5l8xMQ2up0dApaArIPYck
KpcQFCoalKXoxPy/mLZtG8Rl8fMjjk2h5XFjE+egEec0+LCclnyVHHL2LR+4X5/m4U6gBbIHPiaf
QcTaQNnkjSBOHAFUlf8vlO8mmnbTBPRJG25b7Kj50wu0uGBEZd6nGKfJ5FXN2nDd3CIQFCS5ABkk
W6Ea+xxQ983klE8l9y72lVvVE4MMh3J6g0HdfGLCqm5XsOLymXNULVpF6sEE6L/zOMknEWPBHW9W
bdlV8mNk0yzuICqywJh0FcBYeDZFznB09YmfjxREBYFjX4DHMhfHp7+OvYeg2W/TsXcnh5s+U9bw
vdELJMPLArQxq8kNSZRa/5toVg3SKiu+c/41a8GcMteXYc0xVPMOsv2qCGz7h7cOaOQmQyVOPfXM
oYYUpcYfz+acEnO8AiVEEMFHxfmbu+liJbP//VZfx+CoZmreRMCj1vO3o8+nFO26Y9LhSG7NtTGs
oWw2s3Exby+WnrW0sRd2GiaLDN73/d4lfsYE6ZQS7PiAe4zDB1mj5xmhxi4sxqAIafOHeLIFVDGR
K6ylgjgll5cssOowELeLrhnMhuRovBQsjN+WBkgWVTCsVWOPR9GjGTz44Yf6iSFn53tl4ZU88+VW
i07OhdAyHQvIbEleS34iU8Hbfrtg8BMz+btMdFDf3yNav7RaEPAq0lMwX9lwSxQA2Syh9ZDMKWeW
mGElfjLhmSjjcWtV7KpUUl+HSACiJ74DrwFsvOHAG8FLHs+iqMAY6sV6VvvGMnsG64c7iEzRf/HC
W50obOM2QlbIRfkZYHH4kJ2NMgSiLE7M42aO2vWFOGNHCLArbketVnya/yaPsbj0EDBbUguChCWZ
N5I9L2tM5KMEn+8dGLKnnahaFK7Mh+FaJqvCpKAnjKJVPIeGP0owd2YhaqTacBGha8qaCl5GOM3c
07i6NoP4L0J7L4Y99dEumcFyTi0McYvJiaBJldiy3ds20+YDuZd7yxCp99DP7VhFkTtMH2eJ2YIX
nUFkHqPxfbHLVwrBkTw/79ABfRu2l5C1V0DhEXxYsplnZJzQR8QUpFKwWntp1s/g6SVZ3KXZLM6E
JJB+GqU8IfymPO38fDGb0JtFPhK+4Uarc6uaeDgiL7k8cWJ6KI7KEfpZANouHvedqXJ1wb5RU0E9
dM/iWwvRZ2xrS8/ixE1VGq/XaP9xwb9nFgjc5czIh+2A006QxF9EmjnlRwaF4EFqTdFpdSw1ug97
xkVKImlYfJc1wVNzggwfk3kHc8ipCcIylD9HXiibV1A3AlO8fpEI2hgsTpcjOUAPj/fH4xNRbRp6
ptIvFAQ0I+g5yvD7yhisFcsUyKR6+Xkbc7oOJAyf2H0mX5ohFjJ0nr8mlmztRTHnGt0mtHfO2Blo
AC4SgtRQfpBbVT4WNTFLZ2UKYs3jlhZxlqLFZ7GAuM7OqNo90byMrjGdGtZnDAR5N9uvtd2ix8Gt
zBLQ2mF1oiQBplUSxAxXRzkZfWISzZ4nsXLuHlmnnmsuP06PJKHWcB76pvyK6YibY5RuddH4o1aT
NDmrw8O5AKUnnwa4dFRkLGwKFajTxgY39tgGUk1HBiDUGzFb0wLpzstFDo4FFLVlBCyL7GToeHAC
kGOvAN+r1hhb1or57Zb6qxNSrW3/OcrHgfhaXtaVjIpjgx9Sk1+QN0zKUkqBZjLQ7GrhY/ywgLz0
kK55mWwEDcgp9t7p0e97ILhB/SWA9tVIZAN14X8dqgBvjuy6LWWdj0EiUQIVZMSg/soOl51a3e9A
Amb5MitMnt/3VOUb+0GwZVhIuii38ftHc+lpapr64LoWroP5rJSubmlOuj0tBxlmoqAqtBAJuMxq
o9f6OyP/uYPwCQpQDIohYEN2Ijy6a1dzW+YamIfI2G1+a1XAFRqejx8f7G4sOM7OKICJFmTmTqOs
nEQ7Tgj6ukRxkuCoJ6MR0qPf/4Fuj91WBf8QgkBVDu2itL40iyZG1KavvrRo1EjWE+wae+MUYwdZ
oZ6a38PQSD+ypbNyhti498eo3Iezjn9t1EXoEOl7jIzqkZJvSXHuJ06HKwqJyqACXP8NZRzLixII
aKHsRoI0b7v8DSYvasUyvq7zWPIuJgdjlKFM12n0CeYkobXNh/y7QEmMvLEl9JfRN032emNJ0QLu
ACRdTZWsi1QRQHSVwMVc+Uxh0bUp4sDgdcu9JDt1m94Z3EftAMEflFwa6/7RES6eG5nNP3OHXMAR
Z4bBzA5NK7DBLfTOQdT8nB7TxJ54UI5CPi5aeuEe3JISNOy3mgBRg6E4/vbu6fGum6rNxOIAVe8D
X3S/gFlqOaS4Ihr3d+k+6lWDvQ2wiBz0en9bSy6YyVlFzNjXIFGfBeL0kovCFDD+6G36fNyAR5xO
Ff4EN8sRsi1OPO44GOB/0t0jnt/JbTPNyW8Bmwsgm0INQrQyEufCvRNpqD3IpD4UUw7TfZ2Gef+c
Mx5dQjs8hrySH20mZRrn8qTnnE43295pDAHARPzcKUF6InUYNHXLUm6NDiYVPgDrRoy8iKMlQb0X
vWqX0FW7Rxfsm/TyuB6Ek6TZgOohUjkCJjJDYQtC1vV0Zaqm4Jd8BV4Ayi9KDDZt/wn6dnAaTRUg
2mU6voXfb3bziXUeWYz9uD/Lmy4EZuhdCaYiEz94N3RA2sjJKH8LQHMcjD1GBw0/Z8p5Kezx5t0c
Vgpp9YvWGXYC3kZjQZvn4P0gFwqZCqKrumTnLfhZPw8T0A4kcDJKSaRq/8qanhcpfFtBS864D9w8
ySeLfM+q/3nUqhzjo89Jsp/GCk1M51o/r6SOUcDJqDKInXWpPnvNC/UDcIHXVl0eERdLmXnaa1mX
HAqum5QoNH9Hyz51yDgtKN9FuMrUi2EOMF+sSnkj2nvSwhWF87ZdYCL+2NGXPBYzLoTzo2xrVWvJ
96QwvOg5xyRuvN+ax5+HK/3G5k3c6I4Z/V9EcwbiUxDVPfzodjxdcLKvNxJdhtyQwxEk/waH7B55
CNx6kwYlyWtAaH4CGAwqCPzgT/APPgVPq4JL7U2fY9gGklLVmLnKDh6f79g94Jm2TLWn0TcUghBb
Mxwam86GzYKhvXOCX6WXWlOdoQJSmHWW63vdwoohtchztRD8ATTrIvmmAFG/eSNPgjRXs91PpScv
aJ129z30ZzTJt5K8229EPHgCV7iPh14rRfz+SQl9MwGdOYg63uaFH1O86gozgBiEdi+kj1KJ27ki
mKTTKuT226IOkqNNEUTO5kGzu2QuLlAkCp726PUmCaDRFNVatlpEuCA+lHXPExCLl/tX5J3fTiiy
1zuqQXp+xewJfrCeWTPguM3Os3zKFdQhw2lxkdUVA4dSZCWYEO9zeWZeREI/TZTxBvBSKZHYuSGt
R7XrbzsnljXF2w4Ir2/2KICIegU3xr0arTt52Wlkh++ZHiAz6koTO5GpeJnBhUSbSlu5cIZZReFs
vGJdfEdZAP3SOEwySiNC6t9mQKKi8LdrmIVOZmalkut1vTmVmhWMlinbe4tUoVwBC0BQPjRNugrk
Bzsqqo7dTVKIJ7OY7B1iOXwddUEaGoc1VatVhptBZzpYU9f9Wc5pfeQIMXsbYL5BdtaO33xI08/T
/L24ZJWdyflPLQnXVrc9Ag7oGc3vWIJXkeoFlprMjgSg84NqikAqhxgorep6ReWVWlPwR5OlOPzf
PS/t7JKacXnsZysfYLOjRB0r1CScHEwCB9U9XyktgfVwWs2lYdHJAFMM42lhAHv7QpZ6NaZhs5FR
ajdRD7QrNga6Suhnc2l8K0LVZilEUpv87YlWQu+ROLDFTalKutRUbnZFHEkstvxMtVUYNgde/lv9
teTRg9yk9PHa2AU2Hkl5MU7rnekp//0TABeHoUZUlrcyXt8b1JQivy576GlpYVTYJh62SXNc6wEG
UftuWbaR2ZTfJNIXXdgbvu2/7A5vGl5BofoJ3ITAuXh5JLekOhSBcXXUqPLc3TFCGV5ZH8GVmpiW
FXkEoiIXjqGR4GcTxRgdcALADqGTrBHr9FBmO4N4KLPFoBcgTMZwmwOJVqOjMSyLHPKXdpk0TsTj
FCeYh4NJMkagvVf14oLvYOTPmmcKPM2NmEbZTB9NJM2kZFD0gl+2/pOxikvKOpCW/81yTl5eeVzx
hhgEZc+x2b60NjZPNU6jfjtXAfY6BHO150RFPevS0xGbySAAijSe/TanssS/Af6O0Dfg0OEsZsv9
NeUjXr2G/E9F6MU8GMvpgeDylQ/3NGM+SC3j7yVWco0bj/vf9WcwCNg3w6jhek/ArhdNiwECMiZw
pnuHSVj4W3l5eNuhsuVABs4TUsE11DiIpaAMubI2DY3CVvnOjRM3vHp6/Uw88knsuF0tcpET5AsX
NCER9d+Y8ecZE414GqnwfZEV8tZIu3qeIND/nSmNHD2DCe8FwI70ipBMruu61k2+1euKlv/l3WUn
nj7WTYVG6+9icdOQ5NOeCdpJjl6cjlQ0gRoS4hlTkdUxFVnhD5Zv4Otn1Hj4q7oNDI/wG7A+jodc
4uePzzJx+7GqWI1ldPEmNZc1bP/yXbD6en/KNBGNszhqAwXpQ+u3qgQ5zTfgp2z93uD8IqAl5dW/
Cfs56EBU0M1fc2D3i2VF5rWxgOhzwZCYETgbwi057Nefric4jcdzmLKhIALxDit9bjmZevfLsGQc
Sdt7qUOQrfGZvA3IH22epHjIYPt5o1zdIdAncxb/JpbTp0dVQiIzIQGy1CoEHuYTnsZhZygm3lqj
V7LEBzLpDgkC1XSgKuOgolodpdDiJvdY6Sbbjk8hYbv5j5tWMzU8ZmznF6cFPJw0LxBgl6syIs4m
njbcHIAseBCEQwB1HbqNrj8j7EXa5NK2vaQ7F4jOf98Y/hTyy9Al7cDCZpD3Lz+4FKOZUfQTCQz1
Z0b1/nQS31zuvf8aGFUx+XOAv07rXJyMUG7QPg7RZ5BQEtc2do1edohi7XUccHSdJXV38tCF77f9
yJg04mFxowd+qsh4d1uhE1ZeQ7V43W1vgMxmRsxZHSiNyxyxupv6lUzqpk1r4KLJxDvb5Mz79z8d
17bYQNKAm2eT/hkIUUQSl/kRLE2WcuVccN2AcBpf2AzFMyQOjs+URy0swAHhbW1MAhGtYlLTyy7q
2M7LOIF6NsYkDM3u509gygHZitNWEMJrZ6DLHrCFuZz8cVcf/kLf8/BnfKF6MQwlrE8nmUapqpDG
+8IQvqUUhAGbn0zmfXa4cxtHxIlNX+6HkPotcwdCjEfB7P/jVOrxptNQH6YKbc5uq+4qWb/XWcDR
is0PVPEmod5ENfY61ZPY37PgYjKxfM7J1xKiRVxxmFTqMG+34G7oF8fCW5PSXwX7p8x4AutCdbjg
BNqQeVFlude3KSkxFMcK2niH+iA2+Z9pQnscpp1DOlfdqET7iazEbgqFoHnqyyJMJuX+kdQPDZhM
CtwSdomDo0ugVlkvgcWFnoWfnQr6x4C7QgXifnp9pXDwO9bSViGUSdxUeWGabJOKcy5sNF/fmc2G
UAxJ9VAs1WZHe2+KWAYbNNck1Tcoc0+ZgCzkQwDcz434cjoBB2qAc71nUJTVctxDz7SGpFb01/Dq
wSuq8Bro4ancVFY/mOTQju7/8jZm23uu253SYmOb/J7F0NFrovOr9ILKhCHDkm9SKEZHu8yGfvbk
PUykQEeI0+yf0eW7dGW3z3jqYrJyEXAlwAnqulFzG9pgnwlKz+NYstYUNuLJCvCBZCzQSPj7T+O3
Y2nCFiu5yP4SmuGJSvDyZ8r7lFi7ApmmxMds7hyGo+CFgecknSCRNrxenmx04CSgWs9+nAaJqUky
2uhXv+v5dm/4/M6eKzoyyQihTn500V7cWodjlsSqsHxIB1fEy4sQLb4aZCO7JA4H7zFKuWPd8UzW
HRvL0JmOlKmMwPRY83pcKxglNY31/w1DmJQh8PL3+EX0wVQSqT8IDyVv9jm64bcCU23REMTmUVIM
Z4vgxDsIQ/stvPfGSD4tBLG5pm6l8R7dMmoF27zxhi90EBb8x0TUo1jX78xF+EiEYCm735tKHpD/
Q/1tBey7RA4uJYrEr1u4c8+UNyuuJ+W7Sk85/Y0Wy2zEWOHhNs9bPh/bmXR8Eb4jHv1MQ2WeWA2g
kQHCaQo+ZU/eqFVlRZsqCkECs9wflYipQapd616xJoWWo1Z7F5uTl9gfWX2C/LOGSIxdlHHS7rRL
oPwLNvow/c/MoH0eO2XTkLpjqRnIx7bf4vXG3uVHYoK1mQlT2j9oIwbXtOgOPshYfdAY13DJ2Mf5
CzaQUAApSE4aahMpWi8H1YU7fZZBN7iMMImfmsP4F0DrxKMfzk5wR2miudecoLiTQ+c1U35l6iQA
KAYeP69BJX70NnT/W/+q2IjE8VXLtlFx2cML8ssdyjnb1NvrwMhpjHo839KjondpuKfrJti4mImu
wbuxhMx9z2jX7b50sZWBH36h+ExjNieSAeBnWiLxvkVVJ38Zz2QMtSzTh4/1rr9yL+Q7upBrommy
+kOLylqg7z7N7E2N1Esq3aFJxkRcvqhzl4oFzzQiWesm/j5ylAR++6RwcRK/SADeaZt9HoXnWl7F
WIK6w2vXDvBUX8fO07ZTI1gDeUuU1/RAziFGQXW0plokMkfr6QG8x0VWSswjAV9MdOWfkUaWE3ku
xsLBbJ/H7eLzd/A6r9L3iUa3t9dwv3Sbr63n6sAfzoYlpZkEIwuNMZQh1BE5z9DhLb0RgaMRPp3m
e3iLXkyCXLZlm4e9JlpsUAl/XRs/QpVcJ8dXCX4eVn4lk1breQUtE7R7G0svq4ZVDz/UYaoeo9k5
fALiDGqF5YXGve4csA5PDxNCg4wR7Tz1pLBI6/9JDvpYaIECCVhX/GLWianQSTq80PmDd8Ilr7mj
PFwjtahlWgB1TXdpi24YVZzUt28lYvx9VYfTRjL2FEx48L1sGM6hYbhHtirT3714YaKOmGZ79mjm
r9b069IiZfIBLsoVaittpukTlOwAkCTM54Y3hG28Y92vw+3UimaFQrmy3J5wNvTq+8rSLwslBXTT
pjLU8G5tVAeIEQLCbEfPuJ8VhY3u/yXjtuEmPh1VkBOWVfpNXYoN9HVl1xx09tAKs2/VtNN6Z3eC
F44z5VI4SvfVeOpFh5H1WdX2+r+gMmu/Lcs/hzy6QMUQ9BRIvv+a4Z604gFFlxsT4AzrnkBf85tt
RWKJo9v6SlBNOkje+huLX/wcPnDKZThN7UGZKRfy65Am49rQUWyJsNaCWWm2m0DgJ3MKzOQcmIT1
pRV+n5CGOtnxMTtBw/bxEjStbQs1LCU2rXR3cAjLho1VhbnMUB36KK1LwPHYuU/9LyFchZ+1tTm9
+1fGFfQXruEj3Frju329NZY26b1daH1ygl/pDSfnl6LnpxK17CNV4KlIp1BvJBUQG//aRSfEwMfv
t21R0FFOuAVIsiOwLI5K9q03FWMQyAwND/BsJU/2v7fqUk0S2It8ICY2Pkdiw9kntHdlgsR6p/o0
EM4pzV2eR6cSJot3EXAJTz+nOFeg5z1dirL7nJVtcYDu1pVK2+clu6FmJelFDDe/2Ky1guCwlzSJ
bsaelJG9IN55KwZ1ezehQjFhEkY8elXPqeqhwaf8nTzL9Dh2YAWWbWho6XyjpcpiPcLnUcZ39dnl
6wbw/a1hjZIIllJSQfwBhPDu0DVQizcuj93BCrjvCAdVmeFPSVrX1M1Vq8Lyu1vMJLlhhB2/NxSI
V3AakcjZS7jGklDHtmbXBfKJ7fRd0/h6l8lrcd2ldMigf22g+5vor2BWF5obfmzrAugmHJbMLs31
Uvv2noil3h4wt5WXzL6A8lb0a9AqBQcT6/vtK7iwp3KwQnyhUKrxnntgY1wEVZMV0v4Pe6XNJGcc
RpuRFahSzzqPKrTy/ykE8ikx5MuzrvtYWsfqCHm8mRaSjxo1WN6PVVFB1N7D9OyOc8dHhxC958Nm
oI/wOThT4HrTECaA/axBc1msSanhnjMlk+nsdqH+OH0H9Xnn/KqPyD6fvrGj4qkz2zkUH+iMftZ3
WLkxTlQm+y9wVPJPCeQdRSCR4muc+mToqCfTSxM6ZpXfPnj+qd6TwDrqQjhdef9JhB7ktb+t6dz9
rFTjANaLdD4pXRnzMpXEue889WDpR+kdioxY5HrNO3hKzdh+PP2rTQJqJ/nz74Y73R+qyqE3ijfU
hpCVkWMpVaWpjELqvJoYPj2WfYaI7J5L2WxM1+1bbfJU6gcbv7AuH/ExRU3qGBiWVKSBPS3TSPqb
9ts3Of1Rj5BIoa83Sk/8+EC22WwgpS+FszCZaITpngb0iSutqAzDOtaULb6hy+ilXQQ0/feNVYXS
ptgvzU5tR1BIYDtvVJbi/DQY8zWrnbcE7FT3r5/kElyCkC9pmyvFa98tb2Y8a1SRNwj79wIMrCC6
wN73xBhGIGO7txRzCAH02lxYTxy+ej4YJxYrivtQeC6/5V/rE2pOi7nS68CwUJ/xnL9ZJJWzyG7n
e7n0i+ovxXbbht1BurKxk9Hv3txuDxHivD/YVdSdcZca+P5mqoJ76XiYEDuZ4BziG4IsMyn7iHbi
O4avszW/FprunOny0pPyJOlaPIQq7g1kGP6pqDNTCCSy2LRMJ2pZhV/FUEWREqFb0RPUgN63mDFI
uOD3JRDNZhjBBk+URFZwhS7BFupRDUinJp+oCmhqvY4QawL3B7DUTVB9oiCzwer0CHW/hbh4aUgg
oWO/RSMTCsMSmlUbk8pM6CI9sdNqsW40zXqhK25LUbISG+IT6n9eoUZEstZWMDVJuk5y7O7C23jt
h9zayqjsakVizbKA+I5u+FdSMI35A+h0xfwzJ6RfbvB0ljXkqn6ZRYGGHJlfgrVcucz0+eCmBovT
iEtzkcY4HjB/b597B1t+sGuylGN2oLCI7Oootki1gDgPAkkGqy7Av8Ye9MtX1dFQ/Rm1lWVTZfgA
BeGPzv1i99hBCL2L0yplOnysBaRMLcJUYt+GVR4g1g0dTIjCDcySzrGbBeJ6zfxIaIkYwNdLNAPj
t/W8eeA3Yui9u9Aeosqy/sIIqJs/Se5OuOyImamgEfOpDOUdG+QwfrF07RKA9ddNuavSw6OZOsG4
qysxybaEOccM6YOeHrqrOZv8ozF+L4z7RUodIi5Lx1PQRlqYjH0O4jv53g+/rR2QweTsXirvdulP
NlN2RlAaWad9A+g3p/pVPnt95DB6/iLccovwYsxrCtJthkoidfM9i92MoqFSfC1qz7VoF5N6xwxk
TzZurTSAXUUYWC3PsZLB2HKHibIHybsi1Bg0Wi0SP/ncFJe4VRkeEKzWVeJlHEeFxqhTZY6dikM3
AO2ia97cYc/QOnSov18BKkD7WEEQUzqkFqjHYc59m+BgT5j/g3GHEMN06/cV8T1uArN9QdMmyW25
prj/gvVALsi/L4fS+g2axy/JCqO2stijBTs9/0w/LYqFjEUm12vFA2PIdhwtRCPzxB92VAA1PZ22
0hbMjOJzP7fMjDHTko/IBZVakx2vRIl/lvx6dDdnm5QIC+SGCcynbIAEbRyNUE1EHE7tYhyQy/gD
7Q3T+rSayKBHKP3EOOYb9zHHtVeciG0ArK/DvnRd0oCtDi/9MGkV3BfMcQ5tEMfm0WobyTpJ0ZHE
hBPBbbLu2l5gU9C00KefzsYJk0NgzL2Gwf6pNT0wk2lruberQyKzuYCdDiLK3wvfBOrFoXWd09ly
b5x1X7hoKXvSs6eg7Ow9XaPgqUJMocyC3aY9TLHAIgNuvl+uiMpaYxVdxbwEsl7wel8LwesL6C3D
wFg0Z7913svnKGBuWWeKcQ7/tvqz5idxQQscsgd6JYmX9FtH57OiOOCF2X2kmSpJ0ennrDYYJsjT
mQpTvqpZ2bgMLZKp3X7eIr6cIRpICnFVFcmGCS9MkXDzZdM5+linIkBtyBanRaLI9PK0VdfSK/hZ
TbEv54cxenMnvE1EqD9mT18yW39jfIzGkkKe+V8scvYDFZJg2VNrfz8AZ8W+QKf+QXcfPMi2BowF
o0/U2SjZI8CTFdXxTZWeeK0Eah+ZNcJrEf/CK7KxFgBK3MY70NxVdhZHXR5ij3OTSmwoDD8iXT++
fgLER++yDoRpoa87ViNKGSB7TcXCTd0tjw2TBNhj9+Y4qiZXq/uXSKUlhUE52+Z/gmVRkDNrGEml
JwRaolw7gBmUM1pouM7zYWwu6/KjLsnIWZWk6RXbYKhItlvJDZl3RyoqOA8M5ag2ZvHMBGi8mroj
DKXUQ0wjx41H/fQgloRF54zmwi5/y0jvWVrlEfOtw1uRvj/B4z433dCd9gYsAScvMa2g4S7gsZZp
9eYX09pMH32FEA08k9B9Ef6Q5nTA3vzDvdXdHW/1gSRCtWd8GOI4qNO9agj4IbCqf+7dQ5lBXxfh
H4yaxNAxdncIC5LVBlUURW4/NIr8o17AT4FmP6LVaSL9GxIgcOuBXp0cqdHtfiOoEFkJBTSiOclA
ZMAo7xs+khSfWxQE5m9hlZhj4XtskhA2jLMbsfQZu3Gt88xtOGhAB3bJApc7fLjrMs/AidWZ6IsL
OE/MgUUf9b87p2Sb+X7qT3io1tQ0T5oeL7NfyJs8VDdalp4qRLhNNBsK3rHEJZIjn89axkG2rdGb
HIbgYZziDkALMN5Qla6AOF4ABt3APRqoPSoLzQ0s5v5s8BGRASPaHPYsNIV8Hjuv8zi6tqhiUGN+
2jKfv+WCNUU4S2SeyCL8P8BNV8hj8JRVe6uLaPMdrtPLbt+TCgIDVzl8oZFTJ23BK3xflZPDr2eD
PfAP/Sy3m2c0SuvTvLyoFEHauIM7P9cygkfdNdBJBH/9cOLNrDUG9OxDMSakcdzmCuYtQLwvdLIt
mkCAwQr3vVqgtsQ02bafRixZL8UxRHWVe8j2D1ZY98NYIxO6U5NVosoAEAhCVAfHB4Hph4jgyeIY
VnP0e5hgJb7JIhtJ/6wkj3zD7E0YPdjkYIWjWpuwnB129ipr0+4P8KA+mSTPFPOxy0o/g9r4P6r8
kocKFp8e5fX5qPKGAvxxbQYl0EZ7l1Hd5iDIA9GZg/TuxRcMBVb5vOxkKf1dvrnuJbsKPOUyhpOo
mZV3TbSzvF3n44UZkE+LR38PbvLEclK7Ue4e9nXGQ5kVNTdJ8F2Sxg5Bx2KRc4xUY+e6+XINxY5q
kVadPToInuCTCc4BioywvAVYKC2BXbPK5LDGh26vW6ta5Tg1BLfrbPTrhFxVH6ilZkUPZnk3c6eq
XF/kZsimQ99sH/1Pf7pQhI0Z4kaTNiDvebYIYzR+fxF2MSAEdFjdeqhbXkm627Ii1oLISmvpzQd5
AfCpH6f9imee5nvwuTi560svqwjIOTn7HGAsHuRaRrMcFp5qvq8O2DllZbcwfsG54o1fcfzG3ngi
nRfzjPXlesIy2POyIffMtpDK++Oc8UeEHHlMfEhjJsW/jb8Uo1LpYv38UczrTptRfzETqll34PmM
0p/Ry66QW2zTEcSuYLxyGTAPdettip5jmWzwSOziLZ4gEwdPmhiEq666qKA+IurGTN8cqX84E+zQ
Ap7mmf34laniKXTKNBNiMFxKJ7GvciNf1wdErkYHjBRGy/RoJOW5g8MCOpgma6gVsNxc+qsdkTiz
fC1PVSI1xIg7o1+q6J9hnYyT9+wBBVUbmwrUkKZS9Q8QQzMLiR11KDovoqIbVq4XConRmrTyPAJw
OOFaBAugh4qUmhgN7kvhYGFgYWbDgpUq1yJ8gHjJDJJUiWIGXhq/DQ5tePBOVpJ/PD0mxN+2odxJ
EtsuJE5JGCSkjWi3SXF0CkeKDRlo4YjBK8b9NC9Jyfe1FgTUm+QqE2ZP1ustxeX+13saHlIGP5Xq
PrABajQO6/iVt/2Wr/J6qdu0CO57NcBgJ329gS3ZXQMUC5kho+SbMBA/b8737fgW1K8VydH084TG
XjRL01rrbSfcPTUPQQv4mXJ4nNDQE9ANA0XAlNvvvk0MEUGwF0O6gLQcz8pANV//0V8FHW+nbS51
2PxzZ6MB4GMgj94PuQhLQJgjoAurAtWB+LAjpy1sLwoo3ghlhK9dtO1NtoIhlaB7/DjJ4Km9APAF
kN1ZR+jWMN2W7GhP2XBnJoByX3ED7Nz0C29cK0cvTom8u05HgSzxBz8mZ8by138QKeQ22Ylb1o6V
mokhVWltw31XiTQv3Bo/+Q3/bnfgssyO2okxMXkyyYVfMe9ALeumN8LG9zqsKG/6UuS9oEPZhTlc
PNX87a+mD8D2cvFI6JZb0I9M8JpaxdMuHIO5UmsajnGkmiBnp16bjEkWFc/48wuaXScNeZshVSQR
reHaiCPRkXdbiAN/yXRb8WwCvWimJLV0WUgIeeimcqtzBAph9fDY64lVH+PgB/yNNZY933LWqc6m
frl6LOqwoVTYRXdTJknY1TWpeiv5zIKPsa/uxXrJo0KBKvHmWsXdaRu/2MHeGKcB5v6kTblPDl5l
+aImISm64PKrmk0DUxMEChYrEl5xSJWDyxk8wP39lrhgMfy7oJjFyi8GMm9ZkqI1oyqeUfJBzFd/
S1iyC1ov8V4JYo7Uik3xxRT9Z7zKsnbf7c45B6sXhMdlEbG6+boVZ07REy29mOvdKFpXyGbTBiXu
2h6srQczp7zWobdtilAzXk3hlUeCxyGv0PgjZGKJNR3snbdHMw3TbVyeAR3SnYiFd+vXdCwHAJWJ
I3UqVRpQdO8LhvFpcmAv4aQ4khLQ/9bz1oh+yV7FKvhgmGp8GRxTi9Vma4B6i1MkJOAzWjbuIKo5
7O8hKO0SUTOkDClwORT6G27n+zGQSp90+1Umns0eUenmwMIRFV9JnLaWrgYGwnZ+w7YGvfClvCDj
KQg10dbPp+AmWqGh3uqvCy9i4QNEC3IfXzwlzMLJljlxNuNI7i3zHAol/fbdF7cd7ezVNxStK3va
sF4vPBggz0iQpbXsZi6V+dQd5VKEruB+VBlj7SuMJhNhswTCbGyRQ8lEaXNSkIiVBQYtPt5kGoOO
2OFgBilpjAI+MZqSCj5KssR+9AvYWwdfymPIoKX+N1y9NN7sH0Igt9W2xiDOCCKE83j/exKgg2jl
dbdXDleiAtrZoHdYid62rQ92qYb0HjfLuLV2+6dc6Frv8Ng2igWtDraIKltUhh0SHsgCjHfLQYzK
co8NYfoQbf28bmBIVRXErc26+Ohq04rx3rkQuT2Nfj0d2XIZ4Kit7bbTuMtzKFBAUBkx9T90p5au
7qTUu1U/uvKD3XT8/s0h99HmjkIXPmFqpmo9yMFnvdICDjI61DCdyObBe5yo6b1bCWjuz1Nullbe
poyXPv+xOXnHYQjVCjnI1gJ6x8fiYvEFLi3pWvZ2yhkO9PIHUZn9bDZ0m2uIoNRVJUdPB2RirHvG
1pyDmyVlJUI7UZy4T5eA5fYyIt+HQ2j9CKeGUsJAmW3wHoyK9Lj+7nzy+ZcJcSSYINoOYMAOKLOD
OoH4nx/3BndLjmyG3a9sjcPXGkK78GmKcZxGYvpHUAXmI1eyka4Uv034dD57MtEnhzOHnl4Z7KQk
pBf3RWPfk+EfGZAqmysTm7oUdiZjorEg6+T9YEcyKaXZEKGuItY/bzV3YrSo6EOjQwIxjKv+Bsj2
OU+E/31ZpoJK8rlmeMcJPhPgp+aANI0xvZ0CItmK9y/B8gJI+5W731FW+7cbj4xefgq9P3Q0yZr8
BdbhWAEpVfLusP42xU97AeiaSpk7EnA2va65y5KNonDh1YTj29qJATK5cGAM1Zw0AuBRM6yGfdKO
AiFxJiqX0ig6Emod7Cbfy7mB92S+3QuAdofJxFnXPvME/RGsmlQ5vMnvXqTcRey+hZ4eJiZPfiNy
sdVopPdS0JXPzzae3UTlBxObf8J5heuDBWmU6u9I5AUKCCF/xlJExiB7nWXGq8Hq6J7PH+1fwsSn
EW60w7Ps6AI6dQthejUcRp348woGzMPslo8tYALxuZ4Nlt0Cd2y5N8W3CSR1wP5L/aAq1qAC+jdj
1qbNK1nYOhvbKUTQI3377eU2477TJw5YgIu2hz6XUugeZIeojHC0eTsDBwR7pY+DRweMfA6gPOlb
SdjrvTG52dGzpXPZ9q4/iCRLbVUAyBS2TznUTDXCvijcJzF4wUFz3qCh0uBwE3Xm3sa+IL2OyQKS
YiIIOmLNRJQW4ZA1eaVYpoh4j6OEsBkAoJdR3Kj+9DemX0UG1NaRmBkatpXnqV1FOygWYYk7UQAc
7oRHlCQdT8FLk2ozGK28xKPB8iKnG8DTZA4RaEoxPycHuAmEfo0ngcxmyBZWFSPcIIVxgylnpGLd
D3rsKsC9rHgetBawaPesdJFzTNlmo6aYMRzam1JdHPCcWcLcA5Axexj2LfguIR9tXQ8bS4PMJbmG
PUOBKbHSgvOSbLPXg8XvKgod4etXG7XvPEpXPhWFySWguXziaFm/hRsm0heEtjm/IgqP95iCjPiv
aW91ulpieb26uZYEWW4TCERqHqTsJwJERPyYegJuTsBPdFI/JibxFFTiDdYRtd98TjF6PYqH4hVk
jUYLJIJdsHKpCZ/vQZIeCzFwn3S9LWNUjpjNJGxKuulsQMUeQaFaNxctSNA5g9/NVYViewBlf4zy
XNy6635gbmB/Vkpnk8uJ3X0H+Os7makzpuIZsY3ssqLmeKRmUAvX/awhBWSE0wPzCQOWuAn8Rpfz
NzaC1K69GezmAmsv0aSMcg/IUy4DVvf7XXpi0BIVnpc8QVliBAF97XHYRjqlv41Tcq74TmgXL7hF
jb3n3sllj2pPtQW6+4xBmG7y7ovlayzQtupiKR0y/mifVSMVCHsG5fJMJbyp68JtLgna4aV6dTFN
q26QVbT4Y+krQ2PFPbN+Z08ghe69ul2S6lEx5RPjZd9KcpAsqURaL2mn8pY+IbapJpS15M+VYjUE
VtiLKhhQyizHqcQ7HtbB9XSYIB7J+0pZXCnwDQYSiBLeopjDewVe1DDqw7aVPsiGTZfrg0/+w0vk
CGmKY1nV8evw2Cjv8Koalot5Bw+F7KHacW8Qe6qtdNJedUQZRfqUZNSPWpID3b5rWTOp+zn7yMIk
m1E95l9vos8CNm8FZRroC/XkfnbnEHs8rqX+rtLlOsTYcEAsv3nFgH/gAjHOIE15unyBvfiMNItB
8RhU+YBLC1C7TKrwt9dWIpe1Mm8ODXcSwSbbtj5/1sDMKSTLBMBFfh8ZbuUuIYbouRBay+VUPPTV
uKTzB8YFpZcODEW1ukXgQglUqAt8GyQHTeqAV6rDKvxershDkG0FpUu6TPWWYSnB5tUKPXpg4WWk
j+Z9+t+9F1jyQVA0W35a3mBYd9AJbqpdYi5ymzlV3eiDkRq4WNg5D0Oh8QA24W+WbINpEe1tb3f8
C9CweIE+kxQgbIEFJ51oI9TK0eXGrW/CNwslaY/Q4B1JDxvRZw+QmfLpkEEK5lqYW2WqIEKqa8WF
VvLfNsJexDGnQFSimHMKD5Ztgz5ljQ6aYcMbmUEJF85aH+gelPA+fGOwxzkrA1+pP+JWx1kytARs
ou9PPr8ByZizWZmk2TPbJ0cJYk3u/AmsagO/2bqTQbjFo5kxhnynQtXxG2+WS/y/juLB1ZsATsb5
z7stfsvQqiwP81hRcUr9SAd7tlekAYtURrn2EY81YlJyLywFMpAkjZ81MgwEtpS/EnMAzj6TOGkN
XRbWokqLjT/t8iK9vES5un6bjoSN/BuObKLTIytr3vOBFr3yhSpBvImk7sYdXt/TcZsO1y/YuJTg
JTH+ICVgAhlimJMf2cpm/0ipp+CpqDSSVnTndkfgfPxCpk2Xy5Ohnz1SuDTRsZRTBXyijuMCT5k+
QQD1AQtaiQobSvq5QgKRbuUqpjfIqj1Dg7GgEmKz8Wk0oTc4sWOK614OnkW3XpCMTWSgVDVmfRIo
3kQaDgpLaMfezkaPuHW80vW+cVfYxz/VbrGbvYkSI3c/LwXw3ngaHUr4EWi0cOzZeg7oA+Q6Js3Q
6BL0dV4h1QJwokvUgRq52Wgq6QRGpjqLZ6y323/40BU/LGMW598iJSh1yHSDFwTayX7xoIXPNjbw
f4GaxRQWzbBTpX8gaEhMDrVfVBpu9dJ6S5XJs6OYrXUuV47CNYo6uU122NhhsvQmzZE+XaC5sgkA
m7Kf/2iZio2EkhKh/SoEYdGYMo4vgqiLfb5zk1KsmQdSv+inpK2maUoXbqDlrCSkDE589Vh55gUN
yuZx3k91KIUrgF/vFqccAU0fDunV8rR9dSYHWB0khlAGoapfIZF6xFpk7Q80vaO2i3sHCDqOM8zL
osP+z5ZdrIn8GFVrtfgjGu6elTbO1ApeBi2H31WhbvY1mXuefLEXY3jXiIAsAhFi0TwVfQMrjpp6
fcpGbOVb4qZY3kmem5lk0bAIbLsSu6tEfblKCtLIOBDB/9NsMGDzLFCOMfqrM46MZdPJKgWXvV7d
KOYdVw1jDoJEbYbsFF+OmMl12WLhBmV2pW29P9FhVt9P5aK01HaRX2SSvG6Y/wDiZsQeZ+6ShmwS
If+ciLSvEFqxAgeLrvvVD2enGD+uhylvUOW7ml99AH3/vd+PT4XBF0bR2IRnePb0LL4rZVVSdTKZ
NFGjk4XlD8tViYHPv1xuP4RRpCL/XfS3uMjLg58fNbPNOsydxU5nVLbs+nZL69el+w9rHpULy630
eHPEsRpBBtHYe2Y0wVJUO/XuYLLEj0PQVAWR5O2xG+wLoWe5TdVIrlJ61dcB5W97rCTpVUJuKzm2
F6ouyjtyR2UmPEpBtWDWOlE9WOo366TtGzgRwhGtE0p2z0D+Y5TIZCwgXzEpGuUrA9FHtmayFczw
bfK496SoBNd8uVPab5VsPNPy83RViATak3ZIyZXV/TOrG0Dt2UOzm4rUzhuvwe/zwcJ9oGc0PwNj
D3FH8NQYyAlBM3SONollzsblQow7ergOuFjoiaTEq3oSjGFDlwpbm/2Un7HJ/kPYcd22EDqTOYVJ
pifC6DXxFgxWnq3/ipe/zEnk98AaIG3rHOsY/0Z3DcShyK4N18894wuQh4/eCdSgI6K0ElgCNdPM
3hGuKnlN4zHTyt1D1gO03OH8j+SP+nxhYnIku9Mwu7x7aldn+FOvGgDcGokLU8xhuZbvrxU9uve1
gPvtfETQfGHm60RrxhPDnG0ZJWOW9rD3BQBkTDemRzFeOfTBoRceQeL+U2FYZg/e7TMJWPjR0d07
NBM5bOgK0a6vD5HU42ejq4m7PDqhBuRLWV68bHXKnL+8ez9VQXDHzb09IEXKuzN8rAcXI4TyNISH
e2P7fWfNXj1pxii1DpKPWiYxFUMoM2NkYBQZEiP7SVioMYTsRgNtJAx7/0bUZWJQ/2wtUVD96y3Y
/uflOLnMA5VhJUBmRwWfzYF9kxxEhytTfG7Q9K0zWLIiY/q8xVbhb50JPhP/zyyDPLd2l989Plc0
2/iXlmicaRYj4GrZd4Tn4ymxhUzTkl1vXXXiR1rXbffPSWg4zhSkRltMHdHLiGCZgOHJ6PltagXt
hJ0yKX8IDRaxWe9MkXzwiF2Loh93WSAcCk7r5nXrC2l/zWEMT4XRU6/ecNV6nRcgxq/3fFIkZ2Zt
/11XgT3MH/Ng4OitBqUk/St/JDzuqZIn6laP/aF2dUQ3gP2+lymYNpBzEORrqGMJKivT5kzd6eoY
LyUBUmtuR48F1DxU3wLvykWL7IcOOdJ/Dw81LXTQqj2PRmWcJbCj1Um2RtWIV7qwb8RS2zydo1C3
n8DK1wH2MBU73gfgPkMtA7jURf7pqP8SqF4N3bWKxPyK/ci+O3ZYTHhkkyiNOr4uqRqUfOXJDSz9
UHdChxKEUL7n/0/EUU/RsiOsSWRQq/yi/TuTjZ3+Pgi3Q8OCi8xdLbxIXMyVilwr5QzA5aS5PV1y
W6l7elIjYaAR1YnTvmEL8rxZMiyeD9YZMHmmg/kls+LtGUUOOjK75aXNYQamL97QUyXLt+LSUEA9
pjBTtpLlfpyPCph3+K62jtF2SoTqcfWhXi7CeCN0O12I7mFdIxtCgiNC/DiHeb5W8SZ1+tee5akv
//dWfGxU4LqgfkjpkZtKLUMSq6TUZXqVh/GNXXrBrI/lX8nSaOpamExIhBh3R0TZVOQjKBbv01u9
JuzZVTgGY0QXpOPaarNxbv2DqWxiGKySRRH07Jlpn12VRUxjDgD0PPzgdVRBwJ+LoWT59g9vDpGr
odlsEC05EwlCfZIpRcXloV/Tr82EJSYJcTLe9NPH5jzeL68Cj5Smuilq8xo7MbJZpw5Udhnct2OR
ZlNey8FdKUd4IarXDg8VvFbz2XAUJkAsffXVVrMkoKfvPfG9MUlT9tX0Po8gq6d2AwnBeReEs76W
RJIFLmi/UaPrlBfDDVFxyR4NHcliiT28egwMpxHF5gSliq3ZX84JGxsttWCGy96ecTldhfLEFTIM
fRuHcxSoIVm2afgAWC/PBVbGALG8D9GHhF/FqwvcSWuA1Dxb/liwqpPCc9gRrY5Urv90hqHDJhPG
UdAs8DUzZSgZrGu7la2GMryPjgkf1puHcBwhislKfK7zHwXM0Cm7ZSS6qvvv0GOpVWUDmVUaXzXy
tSNxNjSMEOfJBqzH4U+DxM4yHTazgUWJmW63ohWPsBcipDUj+DxukRxVYkyIUuK7nD+eSI3RjyDz
LpMDMVXcJlPquylpsZQqQs56Wks1FIzuFi4NIH2uSqzaKgMBHHU97HqWq0dNthVEQJeKhz0boPPv
gmabZ9fQSpOe4ZFgDifgYHbReiaVMNFskwEzEM6kBRCv9qXRkFJAUAh7WRlJ+e7OoRlQMPNLskU0
oWNzn3zszaSeWCjt6LdWwKAEEqKmAUVr1EmYxT8x6bULCtiyaa0fK723jKkjTZjPy96Kz8M4Xmmo
dZn+NB8Skn+CnNmIbg6a4QilBuVAPB5+STzbOkSoSGXcPV7grlSbgJqZYhAdwgu44wC+OZv3CJD/
i5hwqfxTQO6Qzu/HavTtutY2NnW7vVC//je9Y9V/XC3SaagkWnHSWP51BqcQhyqMANyyDQcH9j6J
RpDpb8GbzNQw+asE/VgUe5IQqPnOBnDcAXFyXsHAJ9S9MHQJCOmuqLQwhmXXP4ma1lunyT6zc3dD
4xsjSbDcFtiPpJAo7XusMUeLx/yXsoMX89NgTbZqfB4VLiAnHIM6U32n0bpkVWWq3UG6XbYuJOIo
6ntDseiVR2CFtPilFpZQw+U/1/PixxBNKLHUXNKC5cEVm15Jf2GGZFf7IAacjxZIyzx9fKnslhp9
nOlayjaTNaPWeHUCxzAZtQ0iUHioiAyi4Ugp9NKrt3j6qMbVakWWaeDr8s7PzxSaIhV70iR5cYMl
c3IRGRF1TPI904lp5iIsZiVesAZJM9KzLVfL6zoROX+UBnyGxQpjcVG73Pa1iwvYkMQ0REmfH3bx
nabR8JBxkj9zAx4/O+U3ckbxUawfKJUKWhCqTp9f6QKnXJX1b+sGT+pa7jGPsMxJbNo8+1QadxU9
dBeGWbGNuwrwevhRxIq0V58bKTmWrWzsrN8JYExm2lIVO1IwTYpK6XeQBEkd18O2dULH7ujoMOkw
L2wzO7gfWCBEtwxl6py0W7FDprPj+mkX2E+pm2qZ1C2O/jdzu+zQ5hitFv+sVC69LWHZNYuVhfiG
m0aNySF5g1Ju9S8mxk6aUKJ9Fj3zlsEF54fTT7VzrY8wjn9UGDMnDB5i9Rv2M6j6ujbdghj6DHpN
3jnZ0ujsuLlhcyFb0HCHKBJVQaR5onHiWMErPDwcwGmGviOPXTRw+nReC6I+QB87OsvBe/CQdcw7
24IyAPZG7tLkYu07Wv5FU+AKH9Wv/eUbWjwOH6ENBGXnwJDDNH6xhbARadymd6tQwywbJZtPjjLO
u67VDuJA/m8asTCesp6H74MoHBr03JPtZPcxIE2AJTioLOblhTzl5VAp7QHDf4R7bwq9AYh2rsHK
tmYqhYfGwj51i78aP4+PPUV7V/K2g5hB9Pl5PJr8r0PLRpZGrtIdWG/94fOlq6HKO0wutbJ3DdOR
V7mF0gmB4hdtJ6WBzhifpqlvvSfehNioatNsFi7/ZOPZA80TwHDZjYesgs+5FiOjpKrB86y6unOY
B8v4195Pr2NsWGmVi497EK+GuspJSsbRPOjApjCEWqVPtSeO6orw52FwrYdI/z/pQ6kicAPnE8Qp
pvxUCEsJ6aoj9MdOJX6Lb+qsLK5WEA1bSZtuhZXCWVD92LNDIyxXRNyQGFUwtI3PgP/ax2eamtIB
WT8efxPzLn9H+v4JYmkmPDRIbhRtnK8FSEWa+LowgoMNGBmFGJYTqJvVd5r4z63JPMvxSYY/B1hI
XvEpkfZxBTiwEn6Q0Ruf2lPb2GrJsuyYVLDjLVMcE3WmvxInGGcpkQqiybicUiRvAZafm0RKj09e
+moPEIUpLsgZObbaQhr2OSnx2rsMmpxLETSGS1KQ2k5RPB4qTsvw+6VPA9SiPBQb/mWzCIehCMlo
l9aPxG441eYK/lVbYRxCuOMrsk9Q/EaLBPgkqghioG22FZv/C3lhw8qeHE7VsjQMrC46igvxDAAX
k3cTxziweLNqixXsf/zy2ZJGB62DhZpF+uBGsWlg5j+xbLBfGaS7eJxDuG8WLiYlC+LjO76oPigP
d1dT+I5JeIDTm5NGz11ddIKZ1A90c4N0B9GhbT3NYskp13XoprRJ6ZsROYai8Y+nADhfrUwCh/O5
RITBiRyUDSmfSGA+BXifEwLi7rNPHiwcdjJdVSIE+6GdBpAK21Y6lzILg2myCEycNkVg5BU64Tte
2QMW+5N2kMsSgDzY/1X18vOBzR23By3FsXlOizapILHXqywPNZrxx3gpi6iCbMBplP1I5EJpE0Au
V0pNyAFmAJsj8VsEACZwFXAwuHtciucOaQfdt4+ejD+srtUZ+AvXgJgK3jgXYUZjFmEnCUsajZOj
5aocVWNWo0zSmnZde9HjhKSgqc8LQ85WDjtTvmilKxvgiGcXJvvNSCDWLNltdjSiO1jZkkYJcFx+
8iTlF/xFB6x9yWl8UgPID2j3cv077e1qy89irev5mA0cQAfYHO0tcdupxrooMcegHEsmSFKBiLjA
q4gKkuJlePOPmcUul+ClZMA27HcCwciPLr1WynvvKt29WeAJFv0gg2lTCB56IbePX3hUI26Mqt4g
bxQlYjqzgDHwhgh71+Us3J0XOmkC1gNHfW/NaPgSNRxTRVDzGBy7d6GKRnCOkHkphHtYqBTy+FcP
k82hwk4rfS1JJfCp1H+Y2R96ngrqsVAz3MMqzmOSfomgn841CTjoT+BSIi4mMM5bplfpGQ094+Wt
MEYNB5HinnuFIsfF5BC+9EcArajilwvfJMzfjkkRwhzgtoGvLDlxNHm8ZsLvtvero4sbXIcbGU48
N+mzf4ByBLXjcSdPAyXhVPBjoJXrssZE88c2oFTUIFlLIhTyHVkG2D8B5ZclcMWB6U9aql+epHQ4
nyX85pguI/5c8nrD7bqf1y3p+p/s978/R4eIkdan3xtLxrMoVu8Vd5CrqM+GSJ8d7i4Y2ray8Brr
1LjCT5qXvbxjkKLOhZxOwyEAXuBf6pr2qQVECXt3gwu12Rk3jNke/oSju+6Jo8YR1IUPh1RCndBa
eMlLNcpCgsbSoRu7rsSFClu+vzg5b8n9BzKHDKpN8nXfHgC24w3iMFGs7noGUx7XtqZuWUCIENSy
pbtxAGjx8/JC9msuWkoSOdCOIhIaGjTkoGFl4wyclu58JMoSKYObrUuMn5b6wVP8QsQm/n/nJK69
ZB2GPXb3TP7t2Uqk3IruO4RlYs9FTWtjvW5q5fuqIG8GHjpW65iO5X8jBdY+jVZJpvlRFfccm4Nu
Meq/zocBhWqdRzfGakgwoQzQEfnoouHncGc526OIZnGMQK33xSjgGXzcyfOpYaNOPILybm1SO7DT
doK2yr2DlEB/DHltx//szZBwQyyg5ESgBC9dlBBjYi+DvDigoFKDU1j5DT8gjswZueUeCU4Td2XN
RtdGuFbaACQr/QEgdh8kCg8xAkKDhF8r66A28RJJmsqE0ACfz9/ICoA0o99FHc2S+FWAMBi3cmn0
LwM9Ty0pspl2Y+s8aYaUiHsi52RwczPH9BX8J0YTj5FQAMtUpfeiVnuh1bdp8X4VGELJ0o4EIunl
qBf0k0WAnABUhyXdjPUm+iCT3Xp6WVLJbSQfBQqNo9aGQhwv9To4viu2zG6jkdXR4gROc5C8MfJD
4mgGjTBWR40kNtOEOvNSBYNbMBA2MkFHU+lOXGaDlRT6HUNff8oZBhAYyf/IPSYYY8l+u0GWzgvC
H4un5uTfHSUE7ZWtPTABEv6kMSZfvwWsFl8+A+kBb2rCSy32D77lYmpoZAtgeyP9sD+HaceXsWu+
kYduWbjGA4WBk0Iy8CeKTzADpF7kuLnJXOcdmPioxp2stFJybBKNGjdlk0N4FoWLCYq3c9kyb6iZ
tpuYJBbmMF7+6Pcsn5QL82kxfr3QO/cvCs9LDjAdidMuQ5l6oqrjEhuwiL+Br3+RNecqGrtuAzqC
2zAPwfQgw4Ak2HKCW9RyBh9AlIX7a+QXWmj4/N0oLajW2uv3MrbqGUPUlcuY+ymzubFhJj59zuWk
mkeyyhbWE8HWHVB8YNb6eQsSx6usP2679gS7dWDShjWEuhglqcYmIPUac+JcS/CMU66CKFLv1ufO
l06+yEuwCf5XMNtUCoG4YQzwpsv1wbz+As+KU74RfGo6VOcSRMJt1CcPmUy1a+Yd8WtVKj2q6U4f
GzfqeQ1EB+4JCHJXoP7h9TUDAZ00twLT7uxix3R55AOChR7GVYY2NhhekkuxP96QlmFTNKrB4v9e
pfLfh+f8PXOG8Bx7qucnvhEluZgW2t189vkyP193zpf5ELFHJQ+HoaTO3DJuUOaAbXhgFpbsiu9U
bUJdpg3jMmFnMdTM+Dbcex1FSOQKhkaBwBRfj47jDqnCJouZm3WIM3Su2xAMMHtK1KKGPkpw7AeV
8OVeflZMS49BZFOnWcbpNnUSGUnL0g0xTjHsmPMYZdJWUs0uToNAQ3rD7xrdoyryWqPeSFBa/O8I
aunifbhGkMKeTL0+QZO2N15KTGPG370xM8qebha+O3RsaW7C5iWiSn6AuSMTRYJcz19fUTgu8fFL
nmxKnAgNTcYWmU5wK0zthDdkMi2hDNLlkFoX1kVpnitR9Uul4QZnyTOcGKcLdwBMcnKBEaN0aWZI
5/lhg5aNPmVaboWn3FomS1+/wAqQQcUxqCg5eAIUVAW0+IScBec8xPH+t+xuf3TanDiC5KVicL6q
UlSYI/vrO0QZN5FCL9Yf3mCSkyHSvLCTwU0ql382Jm3rq8ibJQGOe5Acy/umgl38MIvHCkYyDbJJ
u09kYg8HPOLRMadTRwllCBpBGfqc79JJzcCc8zhIkKL8sbBOVSHJU5oIIgxBj/1826KL2IpUglNi
iOAdLvDywITMMDKDk+ru948IiWIbWX3ItgdWXsdv09XRcGHGONMrjWSaUeRVqDd/dXFY9tNeYnFD
dsz9tRd0+fx9BdErVAW0fEvkgdwkN38WicZM8UL9tqglqrP+K0+bId8/FTCzdYEly3tKU6aFi3tK
ohBe7qa73kt82n0CTNydTV+4RY4yPOPlnvmmuR6Ml9+OGYjTFcxsUTlRhNgiCfJY3PdUttxUKdiI
J/4VXHdaijTRA7JUpRo6zRKIfgLRVj5rOunx3kgkAW5P6k08wUqXt+7z1ldwvMdob0G0vlLZzksV
KtNF1gptPTasqtzfgmJWoWUjHUasFOSXY1P4WzJHEIMCsCtFQyrEW9bvXXtxD3FkzVuWcqS+nYP4
xlfdRtK5mr+YKkdUQ+BfVfnXW4xEippgM4X0ThdjdqHmJvck22CCdnpVWfzCdnUKoXTFJfURGXg9
rD13u0xUDiCJ/69ga7v2U6NNqZXBSeQ9JIfprxiueBhh32L4XMdkuQY87hwyUptBYqy+9Lr4YdNU
rJBDa1gt6lZv1PUEYOPt7NqUcbUyESy/JytvXWK9FHXT33DCtewgeG7WzRi6l/weEJ25KtV9gT5o
5J8M7udKkxQhfA9+wwdt4ZnA1pUPvRTpXjgiNlFVtpGjxcivfgrCWDYC3oy7Qvwyo9zB9Nadtq5v
cQ+3DPDSAzMH3F2hGqN8sU0TwSPciEqQf0rt/95vczoJQobk8ATffepO6rprlYP7UcAW8vLW3yd5
lYdG7tDxyEviLD7CZMCWsTL9QF8BoBJwwUVjSJf1FBZcdI42tmtu08bsAsgvixXKTp7KUlhkU2hH
VNHxTch0DT8iQlHBW9AT0jBi+NUOBnGbLuIQdKI131L05GhvVUCO7IGmG+Rj4+Ud4rx7THJOSTHZ
vv9rL4qnfJxUZ3SjfD4yJIcl3y0gQCXKJRTO4IF3y0mVvgTd8hfhTpHaajcd/j0m+5kxwqGSNeW+
DuXmgDEZkrz9A+XneZZuMh6uNDeKf3StEViaX7griH4GquR3Z60e3GdvgWzDVCfju0VYv6eSBH4Q
3dne4Kgou+cDT5ZaLiTt2PCSPdnQyKQ3FeyzownsrsM8ALI9CCVGOaCjTuZZvoG8V7K+m/T9wzAf
vIl3zidFbwMy/4/1SgcCwUa9HgV2YtpEQRfFaSiVXi0XwdSq/weZyh2N/4jCo5SP1MvRgkmYUyGA
bVW+VRoWIA1JDDOH/J/wdwKR4MkPNqjuSYCiTbZrbyI+6sWbvkRepGSNsvDVhpiw2PaRNsGROqQF
WUf1zE4t5lX0bylOGLe+KQDebcFzv1NwdV0V00jNB1qF/ua/Wp9SJTGF4jM43m9eSfN2ll5aqRsF
Yfh7vHcc2lDmTGr6BE6Hnb7+LeRv5ReRqLMelRBPBcW8bR0d4b+a0efU4TXOtcX7V3VdWbsHhxsn
kpugK/iW99SV5HNmhamHGaShT4kOLTx2rjS3Xjt70dkcD/BxTK++mgE63k/lMd44E+cqRg67RqwU
2DxR1uMBFg2m9UCbc5/YGpu3xejqBSuKCFkf0333MkLDwoRj6MGWjBUpYiQp9P8s8IgaXATfzbdO
CV3mvhR9nmf107U0jKuqpT9tkrM2I2GFm9+6eKYgH7it+Uf+7M2fD2Sz3A31bSuw8IW9I+0C+FgF
Vq30Ro3OqnLJ/tffhOOzYMfEu9QEFjNs1KUaTkXOhoPC2Z3lQJa71aXwksumPKwjDP5X3f1WEV48
9E01mmOGwiw+U0AcQyNqleuJfKHWZjXrXeHnR8OePWXn7gVBxo889pndYiHp9xtq/Y6eKvN7aVlA
kb8Q5k5URHWBaeiKa5/oW1fau5SgPv8XGfKDWWnCN410EYtdYpV8HSY1JOOwLyZENIG4VPjEWEMw
QXjIDpgqwnLRf3LO3v8+Kip79GVkjND6YUjjOjKnaLEYYarGR9e1EGEHEjuM+IeVItxvn2jvWV1g
NIGFbKo3Azz8yqzwLKZg9TgyYQeWmZm/xFfkx46eDu/PPjAN+cOx/a9Bube2M6eem9HbBSrHgvdD
y0hq70AX7HxF1NgG+y7SRIhjmWnbfIncK0gQeeeGwm/4gCCXANXElB5vDUEAcOLHbw7mJbLIzHQe
hv927r9sKQUQuP8/rR0aEknouty1OIwErKeIGCVAvj4hxtS4BQ5eVhnXI3eVA1/n9Q3zFqWzM6jK
Ggv3b+0wWKiVuRFVhGArEuPlS9IcnIHLqJ6m3NDgOfffenOJWIBI426NfQYeuXoKpxrvsunjep5S
CLPDW19ajH2U9y36sTbZmmK+tsE107WjJO3veXCI838gQksmSyuKArso4RDIEF41OICuhpTLv8j2
a6k8g4gOTbP3G+MZmBbGDQbqOAn8rQr9naaj4KbPfNZs62ESUH2rmswxPf4TwKEeu2bvNta0Z8U7
Q30BO/0eIz68gcDq2Cfm7HL4XCfYcgAyXOgZQAmDyR7I3Xpy0SHMCarAOGrNj3oBcpzfxtiYNYtv
VV3+i6a+Qo4EmYuN42yBn0/2YgH7Xx6rvsUlPW3fY2WVMggLfM0xAniioBPQdFjKU7jYwWngzWxF
JZn5ITrS7QyBNyu0EqaeRwPFpmPCg28IuJKCqp6zUmot05oEKmUw22+MROfon1CQdKuBJKkGimOn
SswXFZi3G6gD5FbntpY5I5VC8ul9jfVny4qu+T/uHoP339cjcHGFveWdcBs2xH5vxy9DrJhfpYJ0
9SY+cCa1fcQ7ozgc3kdGoNEjWmLDFPZqphEnUeGGhH4Dr+7fElSGFSmofghh9oL264dZL2dpPx0P
vM6eIGPmO1amKzWrz0wZsEwTQ3rks4quUejUF7cjDkdZbkdC64THmUkG7IxhhzcdXK4OmlPf7pYQ
PUjMC4IugYxULPmImvmIOLNX2BJV8bZvpUrhFEH3+Gx2yhkRPjoag1pXliQnfjdjNqXbgnxLKm6G
w2inJAazytprB8E+LWDMYnFmaDK9YWhJ3Dur/HxqpKEAEypo2fukLEMB5MNbKEbR4YleZur3XX+4
ixakzDd+sKsrSMTk/X2EPGFF7cqtQ/nbF5PdiPbm5os4xW4jKW8nliQozGfJuSYUYOHC5nofsZhr
E1U2TcQxyiEtyJVT2Cq0QPUQfslG6cy5RuqImIcuG8d5rZgDUpQxmDOxu02uMQXPWSOWeGHGNfJp
X8WX3St30iLouELgVok/kR/w8QMnW0JkGzxrOpTl35F50dVzB8D0GJNyAqbhMqk4EqD33HvvGzwA
XXRmmuda/ZyAJ7ixUNghKq78wvwRmoYbAQNgj655815QCvFmu31ifWCwiHKGIQ00FYIQ409siOlO
HW4mek3HU/PpmXQH6TYr3o5ZnAtFK0aOTazk74Na1CEFQygGuWfAyDZoY4IYoIK60+U+9lkjSa3R
9as50XFiqGXfrYs1LIgNNBil0Ow5oqlNH1xkIBY0ZoUvRPShA/0hGBxwtXIkPcgezzzV/gO+yvi2
n9Oeg3CF+wsr7d2jsUxM5ULs9i8QBVSqQKJN4FPxHUdXNa3PKVSsoipKoHBoSJX5CEebjavxfT7x
RYH+oehux+3Z/8D8f+FrEawSabeuzyKT9aOep+hMUCz6DadqrGuZkvAdrn4MABamkr3on23uBq7w
3EmOK/PhuMtcVpgxsck3022zxnq/NDAho3tLoU6DAutS3ehI1oqq465phuI4BtL7pN8FVaoX3aYU
D5oCeFMJ1sJ0bgaqqt/A5m/H/UpV+A+HhOhYCUYgcVZ/aplylHQBXBKB9beJ91FEJFyNH4GEDeHI
VvHG3yQPOkSYj71ENTdFL6ARY/efEAl1zhyipA1fVQxuphxCTaElkfQHdhOdDYRjzaZBFxPpa0Gb
TtPMChK4gbOIgx42ZGx2AuQMvqL2gfozNmASElVBma5jctjyspvdUvYjTNMEAFkQmU9XjC9H4Izw
ri2xHmrW7F4wdNCLPpyv5gRWjTeA1q8tVP1aDCnE7bIvQGRuMKZ7NJNnuZPGcCk3b4ykjqKfsrh1
7pI9P3FGbJciPclF43mOOWJWCJNH5E4hejC6vwqj9sEh9hW8Wr8ZzLQyUx7buFLUGMtA4E1+ecYE
JnQVo5vBnPSsdNRTn+begDZGpNd6s3j9FlvZ6DqoFmD19+SdBrfVEpgV1M3ByfbsWj8DRErIPmm3
CVhuKNMhLZeLV7+RKMaA8P0zfJFZnAdLN8X+YY2DZnGncOVIVfQrxEvZ0vNiDLcLSdZkyF7IEIh8
r4jqoeMuq+OWmsvmNhuvOHugJDYwwDKpy/MVmqvIKgMNhSqTbbWh8pgat13dFzBAkqGH1I+Tdstf
fOkDiCgBs2YTtD5WQnShVpUe8VwVTaFNpnS5UMGy/SPQvNnh7tCPqnCTKrew0Iz2dq30hoYp5MGH
TF6U/YoJjMYLajaZAQ7xl7XP9U2hGfzfpdpvxWZ7JLidhhji/R8ksBFcgtuPBYgUQ0emjc69vbaI
5ZVEKXJZPzxzmfJ55uJ4omy3F0pI+IgmJsbDII7hmETycJJRM5sI3KUBuw3iZjWboXBTLtwS9IDM
Rfj2dw7Zjoxl8JUOlsrJfFGMkgzHPjHtwNepBsAGWsyJBr0N+oDVqqnGzqvhoPQJ62QlRhNGJm8q
LmnhI+DeexSgBBAp0JWwAqV7VOCUp6/AlAWNK5V16wTCSPlJD0+m011w6rnKg1ULjCu9aMsTPhUy
U/7hO/pORQYDEkb1GOUBeDOtVcEf6LjP03M+5zGRfVLgrAF+vcEUP5JuCJgzWZSx6+im6imoeI0G
LzA3uT9fzfIiMQzqHzKFUzs1euYATltGwdK9ef9oW0YAolZ0BpvF0h7o1jAJXFFNKVDFEnVaXT3R
PDI+KFnHb/mFj+YDqyRv2ss9x/yB50n0kI82piW/FILG0KTN+SGRDoK2LZXzP3II7dIr81mlw6AX
0b3/jWyHBTBj6kGkFwY5qBSXqDoGmvM8Rtxlg6vva96kTv0DPSz9US3eUJAaoQ3uMucTOywfWUnh
9Mz50MoB1DjDlseDEDwXssGqQK0wqXO/yPKFHoEDIjRwn8/o6KE+Tq+v99a/WGOUBuHQ/GXVn9M1
WIVyAlSM8XcGVd3iH5b6ccbKyBT7lfX57vKVWX1Mj3yIOBLcLDX8jGEOU0xiK+BExnbh2nS9lBd/
a44oof+pxJ4JtuNX1V6X+sNdA5exKvdu9U3QUyfozm1hGWJJwfsCMb5XEuCtKc13ZG12Kcw98K31
kQ5OR4Lp1m+3qqxoPUtEDS1BLuEuxUnOVd+4DgGHECggmhxZadTjv6OE+ddoytnRBpBi1Plcrw9S
oVtWJ9+pVFBzwntZyIMwpcvU2dIIKjLhoYLh5tbnNgdiww2el5cHERy6nbW64VCsSWB/Tb0uqFmx
Fh9dIdcxH2gPRTAzjOEw6vLIVvM1REmP7eVe6FgVWRirvtBSCBeZeGwo/MDGNb7CtTVLp+3AqN26
hs7/WyulyZPXH+kpkrbxx2bSDtsUGkRovYrNDZ2W/ltiUqTKgdkK7YDpQBVrK/T0QToCXHqEn63l
R0E6VP40J1+UMuL4dqCVYf0czib5MPnhX4I7RSL/qkBGOxzghe9drEn0vLYEWiqkSuzI76+FBi53
DXQhuWtLJVklNBEsnlTJQBr0DhSuUI6Jz4TiGTkFq1Kgk1syBSn03SLIzCwqXS0qSWSftVyMuDC7
ePhNB7X3HFyuZDDw31dKeUaLcBwUV5tfd6wpN2JD6d1JZYXceCTdpoXW64UBsiqHtCyf1NGYid4v
qQBNFCUdy3+eVY9r5mF2NvQt1WrGAWYO/cTsuMQUvWPnz+Gawu0FQm3LtvKymezXiNG/rBCg8GpV
h7z7C08jbtV1Tfae8cOxK3F7UP4cuUl3RVJ8N3lHm932D3W5HIxH9nQzBNKd+HgL5Od2MbUJmtJU
wi+wI1L/dHs49+4VflD3oASpp/cL/SmFt8joBIjIhdPpwfv5Shj2dr81wesm+zIDwbYMN7iKjBzI
h/f1031RjPo1ufeC53si0c9qIYyKQE89UMRKmb8Z1B8LRqjb7QqLw7BC2z4T3k6t1jGncdPSlxC4
qSc4Nhxy0RRcLPJhKUANQtSsrCeJgZRwhMmhFhHMElpNzsxXk+ak4bUBbJf0A4jta7IbASfWFfst
sEzuU7uWErxJf3TECPMF58syYQCvkrPcPL4Fc5YUb1zpzFKMZUz03eErIkK1De7Kte3+D4BGRo4a
Sdi7DyxHXzvRLR/FS8nISwWK5lEymBiDg7kVf1u7ZWvRe7BI1Eofa3d07lotpOak1VVi0+l9K66V
yb7MnhaArr1gZvPs5UymkgTbztNr/l8+zO8jBJvYDZZ9aJoiRiBcxz49J/6jQuHb1os7EJCtwFk6
yYg2sPdUM3azfLLHndWpcBVbd/HtpzOFZhnFpYJ52rE/ohsA0JiBpepvE2Ae9IpVb4gokQPQM5/Y
Y473WFjW8PHBRXAMLPm8KFCQO1KfzT0GFHYyYWUK6kgibpJp8HNI4vMPo4CKWfHPlNwkG5uCqMvN
EVIo4uLRyQ1BFOgxX/t1tX8zssLzKafsIKxo/OMHIpl34aSEr3uatqTGESStt1BiuT1GMQik52LE
zBZwGX6lql1jVdmd7/7fOIENT3wKMk13ukYd3SVe1qr29Q8CpCQgYp8Tly6zk3rf3dc7MimrLkz4
BOyy2YWWaYm5U6zB8PcglBX6hYuIQd0MBdObqBmmGtA3KkzZP0Av5FlqbeJDzVpLSLoMgd5hgS0V
WQ9STV3CG484Yw7wF56fYsc7kPSCA7I0lho7/CPbhEExEuUYZOgIpsUjDNjTuHEbbplgksn/qYwa
QEXH2G/5x4dVQKOwbhrI5NucNdxXcrVJm6B1TzpNazY34RXFATNhsVcjgmlauazeKVSUrEFeDseL
V/NETC1+2ZO+Vtq9bnSE6kMGmuWR/9Xl5DXMwfu5FEvevEDr8WzyfudA4Fsqe0YfwG7P2ENHQD+o
/ifL6oEKpSox60rlFWkYoq6QrW01uDl/JfOqfsClYFejLaoAeZEKROEXJBDVBNhrIPRHfhLhUi8w
l9DAFbbgnUU5kQ7RbO3JDm5I3EH05M4kYyUNCijfA3HPaKt7hmTsgPQpER07YphKI2qGu9i07mWP
8CVypwAaV7GL7zF1at+loFpLg70bGI3MA9ty05haDEgMxJ2Glssxn/t1hJO+DIqVAhrNDxNl1lu6
wal2UEIdURbM2YaCEjWvCHlqmbexnjfLI+vczWhlVcLxD9s/O4pzo4K4Yc9G1+fBlM7gPezmVudY
86gjxGOmXDEPBiCMzOmlL0s0hFYTQtToHUlF+pXEm494H6VDOmYDKK8Ezl/ACylwBRP+Lkyh5Byd
+FR1mydVM6g2XEmAadkquePeotM+j7IMZtVNgktCFVUhE8xB8ldxjSSsH76xeExVcMnXizQ5UqjX
EhTdO5JBNkmiPYYwOtOWWimE9ztE9nFVeHQKuAU8Zz1mMDljG/ZytZQ0gyoKsi6ctrcw3QfbLR5F
EfoNsaskERp9iJ8xNinOZK0/ZnKR2oSFRNdInO6/wvTARGFSy8j8hTeJw41GLBVqiSNAp0gmRBe8
LO6mgEo+BrsxJhvWsVrAxI/CF+3JXzCEzCENBZoRkJqtVwHphbNITjLgKVsbKxwfqb9TZmXJRUkk
/mg/UQ3zoPHCy1/ns/3q34rfIvAdGfsdPNhNL330reZqXLxh5LbSNggRKGaQf1yfACOuYvc0MM1g
WZUQu6QrrJYq1mw5Fc8HP7xRITZ2dG9myjkPN7i0TmZXsWch2txJqiGCJWQIbmvHOyjcwb/e3stF
uFOCtk5QmZ3jF//UHUAVPoGCJvijA7dL/c59WmO4bApxYMWTahcX95Jm5vRa+n/0Nam87syw9hHR
VCksI0C2KqtdLQJn8SwRkzAr4KSyj8BPecUKUxxKhZ0Z5YObRErK6jy6VhaRw77hnVM47sZL1JoE
+fq8gCzB5mUJGlg/yybMrSho8iVbYQHOcrWpivvcuTwdra68NDsqvx1lhNlf9d+of7MxIk/Fd+6+
uBBvSPWzKR1PzUPa6UDfWO/9NV4Sk++IxJYKnSd7Z4fwwH0Hs+yS5BPLqwNJegrgwOvJtfVvlr4b
NvI8SmZpRd/LKyEZIj6cT2vbDuJkntR+xDsybaZcJdnoKBqdbG0pT7t554PijklGgCMrv0xhxHEc
8QvqmH74zeQBuj69WjHonHdhLpd6B2t3CFTsCrmbvzLfk9QbPoxzlKnokugA6gFqsqt5KYPiu7OJ
tAAre4xDWomjDF9OmCEokYA5K//DfzEssadB1UPuhqK6TW9JoWbk8DiiZJiEazLo+EyUCOb5PC66
dhGRwyAHtFTC6wMSIkJGnaOHO/GX0RUkvzgDCgOW+GUYFY7YO+YlnK1IcF0Vz8KBo/kGpvD8oXv2
sipLssNWaZz9rycb2A6SDteSvfRVt+lVQsDaV2eY29dZ3k46yzLxCOrYktKT/TBkrEbWy/JvSrJF
97Ac6w0no1pNoO0rEek64QCoYa3uOJP9nQKTiQhCwhT2gyKeD7SUhSpt2x3AxoZ3fyg3rEped6pL
ndipOk4VjNuUeLxPnOXsqFqUa90kEBKVkgp8HTRqeOBwUPJ3UQKi+uIyqQ3g1ItsLygHXh3jwP3S
jwffxrcWt3hHIWuHc0NiLV0h2eGTzV7jWJkq74a24Sh6sNw6vC+hZb9O+boyessj/mbggxSxqItL
sJ0g4z/lKiQbsPN2mIQp6WquplsG2qo5W7CnZ3B5x55fQYFbt8Q7GhqMxOTR+Q6264p4JY/u1eQv
9TesKuP1nZNOaG6hDRWYdyi0lR7Dhu7MHtmlUsl5dg+qXX8n9EKquj7pb4bTdPYUtIvNAXJaW4rB
5ysRzom8vcmbMDwKfzAL/ljsnd4lds1x970Srr1CDjjTufVVrjZhHAvUn8ZU9W6HWpsOEIHpvI0D
MpbbKPPGmOarVOqg5+2Xh+MtC1PcQYpo73rAsBL5PE7gB5w2h6VqF6dHFDZ8Qh8V8zUOcl0Fpq2U
7ffbDzk7ZKA2chh890kMHCbwL1CSa6DYME+ZLwZ+hTps63GDvJn/Oabgm6dxw7qg6x7V+Re1w223
+sQ3nNbJALW2Z6VIbcG4cwimj0hpI1WVqatAFEnIIm3UsKbmJtLX+/Z935cdcemdylrYum0X294X
BCkBkVmwfGbCiq8Ejz+8URPEHa3VIW8uBqZy6b/LDuHuAUkea9I+8kk/ePUmBxjKh57mr/wgRVRC
sv5/EhqSqnGUWGEh+jzMvYMEWLq5wNiK4X/lt4S95G87DQNyW0QPtYyLbcf1WXhvoFpER+rFJuWY
ZjFC6MHdgTxr+1pnro2uqjCHIjwohKv/OCU9NLQLll+AHck/KsJMw4I2Q9gjx2YDT+kqYzpRCUXU
gPFf1eCuoefRbqphBZTsNr+5ZLW6m2pN3BZ/Id34HxuOCoR3rqzjaVPf2J2o0AZE38jGb4SLjQ1M
Os+ZGtTGx8rml5GBW3uHbrCOOqai0qExvZw/2T+vb8n6YUqibcO8AWKHrSgTBE96eAZhwv94zcZk
EDhmPZHZ5YMuv4tXI5l4dO1V9OUeoksdadI+BfMR1jFO26OjI/+7fi8JudBHEzH06L+5To+gFHe8
WKtJEACOph80JIeKt+NSgZFLGTg6E7ZcVsCClPw4KNFXra2r77frc8xFSmGog1Osj2GxV/x3p8BJ
R7igza2x0B+Oun0j34wCyylHWiFh65PJiwMmb27JSbm7bUdxksCf5p3JohSqLojnYGj4+AdJbegX
zqt5U8II3DVxQ+hl5+qxau/1QR7/Bwfhijr5cB92IuqYgYAWd+EKsum6Ky4YxdLN7WvwVflFkHeX
PyxUrxJsckKNqO1cUjLtRdlRWxDpWML98ONSqHJBMdQ/iPSzR6zSGY2lYXTpR5HgGP1Ti1i59S8e
X9D6WGpan8HF366mYC2HnoVehDlfhOFd34xNRPKdJjjiNNcpwMrjT2BYtvc4AGtGDOEBvkCtmwvX
YPKMII1ImOTZPnRL0a9dv56VypkaNa0DrlVuYFY27WOw7dGq+tsU1XMwHkendhSkOL07+p/OjC3V
6y+zP2uZ4CNytCKKz0SytTN9JYLhVFi0dSXNAgIDZ3mDm1EJEx6s4LznK6yPKy2yTRcEYWj+HN/q
Wl9jkHjxJwCiqIWstedsa26rHLPLzEYell4Y2zOt4HYp5FxF3Zrdm+sQZT7KY7fwlTbhBDcL4s00
Roui5Nm5cIIJuysrX9L1IRT9DZ5j0Gu0+y62fTxBhSYZwwqKoJtJ2O+/TQ6WdXcwrNBIQGTcBlF4
s9lJN+o6QaxEdsuQ/KoOfkZVpJ2ioNVnIMtUdK6sB1t1UQflGAIELDIX9CovTJUT2f1+aD8oicA3
aCO0XLsTxyviw7cbfP4gtA0EFBM7OTCkY3wWqkslbJpKCKSIEq0Yv/zs4dHrdIidx9Yx+OAVzk/d
dhBQOcy1izsuCMDR4KXJ+i3JeXkHkz1z/5+cCWCL3+S0YKEBasH4OB+w0xf902Drqnj/F1H00Lyu
5BqzbvFk2+qt50CAWcwcn6SLGT2OmztDcWpxJa/LqPeVPxN2Y5zpvwNN3EqmVTMShYXoIbQSTWjQ
FE0vaxjKcBfgD2Hkig+Gqoy6E8vijaTvuohNJ/VFOE+S/qflqNz/v5vw7TIn0luEd3rqLBs27fMu
86bLtce4QzMW26vjSgW4d5a79ug42AUPQF/FNg6V3u6ClspblsPqfynFD06smoTOsMHUBH2ZK+3/
qymLKxu69UyT714MEwpMpPtI6iMY3FASY8xpZoZFGJh/0Tyoj7BnO0P9ZFqCAG9uE6VqRwphsjUQ
mcQuranpmevwWXOK/WwWexvtC2uXLUzRmJEa+i+N7VV8qmnlRSfIuMcsKbyJmMg3m5mHOpuMQGft
zW3+peJ1GNa8R/nTk3JhMPRw6FF5pUT3KzP8JeGpmlUdYIwFPoOW9jw7DSoiV7ib12+CR/0THgTw
fxczk8ALnFtJiTxG8xzxLuSAsKir/lrj83juBKls6/4g3j7nTfkiyMEFr2SlQJM5i+rLvh6GKsJ/
r2otTOcYJle0dL2xYdLY6lkdAj7HGL+KDF6sLgQgRVVbDFhqa7YeqSNJACJJx3zDiy0gH19TPuEf
wJMEpt75DWLh+AnyDmOMPd4Oz2/cuaJnxTyc5rCjNrAI/EfjrqJoipEWCk5VU/NxnofnWiC+OVOG
d3MH3orZ6/mHCkRQ/v6Eg/loyW9M2jpqDaJBn5fT17cmhgWdqquiwjHAkmX6HgGe+84F+rUvf/JN
UQon5L8OJeazIQVxrx0pEkkKW0OiwqvkF5vL2iW89ueziuNSEPwsx81m3fDWCgan9D0PDxIyeMdd
gcYzTG0nIpFbVjTW9DTnf3jG/7GhO0HNXYyp4SEQTHFBab6lp9epm6Y1J8aIJ5s08kheg7jDXCXE
/+mmTITO45Ygyytmag9D3f43kWxsKuCyKi+hBAVoltQ4qYAdK4cYkBqp3Mx3vtTzEz4OlfftjFBv
L81DKGZhPVkTqrhwjSQsQC0zsh0YEkmWkNBjlTYVeAW/rvwWF43+NC4n9VaTqwG8r+3QbSRETe4p
WOIk5pJGnj/mWD9WiN42fezWH1FG55jFlIQx6mfjwFTFgpeNQs0SHDI67zJTcCYLDxKzbmVK0n9h
o6OZojj3fVFRTiyD3oFnGhdVQynsdgq5XaFAIrJtSbF38ZfiIQJ0DPmtOiwgMP9SG99NN6kVq9tR
6CCAu23Pnmp/ldDrLzF1abz/c8euhgAjPjjPMYFAHJPhIaga1jVDLpRtszAgSDKmhYBFPhMJKtYo
t02RmSdi0daC8/JUW039a0D9KxAQoahnaH3Q+s3QfQLDQv2MmLzFy0BYzXTvfLQM9jGD4aZmBqir
GK4otT/MQtVkgZS3UbQ9r7Z9vQm0J2piSuljGy4kCQVQXn9joCAVDRe6qapmQ8vBTox6i0BWJCYg
2ujc96hNvpKQT6R4JGjxhglam0p5TtvLPbmG88+9CmRkyAnegwGYZj50z+F6cDmJUXPm4hvdTQ8j
7QhBJ5xnGUqup9ey9mvCdG7sl5hfV4KpgbQElq2Jf9jteCW43AdGGJV1Uo3SLidA5BlKbA58D4Ex
Z/lbHErup8lcLvMlOH5FihQ9kp9Y0YpEI/NFI3at+LaGD74vFWWwq1nAneY5QXhWkFiWm0D3P1+S
ndTkSBFzedHsuU3t1xBvBTOKhf3HMoHYlgG5D9rL2RxqfMLD4bLeqRmiXam0Gd3ege6O4eHw/J+w
jkfXEsq/M4U7GLcIdw2DDNsCg0XqFdxt7mRGuXvbvCDKuV4dXbH764uNek2tyJ4E2a2HDCpFyw9I
2UpzWo0HzF286ZFBvfsZooLnoSeBOptZZGjR843aGY3S8+ir60jgkB5KJgqw7CjMU/EMwWp301qv
oja1rikZ5y9lHoc345K4ST8TrDpFWPX6BaMxzY4BSy4Nsad++QZKNbGs1Y5KXN8a3pOwQ//pNRMB
NhYalwpjJrUQuHWkskTjbGfNhQpf/IJH46R9X/g/2BOjSLYb4reP7F6qbYKZrTmDPH5f6TsAaEbN
T1JBcw1hY2r0VS+EAxL+XGMvGkYsYluwL+f0jcdjRA7x4VNf6he2Nq8nIy+HlspXJ9NLjMHCdJ3t
2enjMSkMV0RgS4izcVBVcKpFSjBBAUv45624M/GL8Jvff9GVjL/PLNRWjKLx4786JiUN47J6fZYc
VnjWTkdfHy/Pv1qpZna5NXMGovvTqzlQXdwTEm+AnfoAQdzyuoxUI+aFNi7+M+TDaDjoZ+jH45ta
mr+om2pq3y35g8sNbUpKu/tDvmm0MHvdMRZdllAQQFQw9AcAHu045S+sD+zfwnRbj52jUQJNEvPc
5etHyI87lvWyGN+u9gjfMPqsZ+enAUTrsT3W4TknzU3zbSWAZkzVBvhJRHZbHDAKt+yu1+v87iZS
ZwZ6LbvOz3I3LolEKUWcG79YwR4o2gyPbVnziCOog/IFZsGKYu4fMcTMGD8We8HxnnQF1O8MN0Kx
4MDWv3uipVrXFntjxpXDaH/aaXxTNn/IBORSTQWsGB6xcPMY4uq/OQkolXTdeNlXfeXh8YEYSU+9
XshLr9tEzf8jrpTbW90H66fPgY1nF5rjQht0uCH8MFusMQyq35EamcWCHI8EbbGQSeO4T/Dhex7k
GP02irFy1KWXPtVvdSbGJfWvkqGH7azl8GcevP8i49DgNoXW6biot4TnpVUpr1V8njPXDSGzbxQr
I4AaYmpoIPbsQoP8TaF1hu0Jzd8aJ0aEpXyNkOVw7drDk0/7NJBEQZLYN1edIZBLt+scdj09ZLkc
GJ+oIesEcwF+aOpNPx6GEGNXK4s7VdsLalP/8SeMELlfhqk3IECtw9T6BhWvaY/evASythmE2eOo
wmpRvbl60PPO9++tO0Hh3Wh1am3uGOlYRO0AMlrBLN2pcCqX4bMt7yX3Ie9tqtz1D+XJMnKY1XWF
G51yE9zkrrT0931C/TjHGKfmyKzWcYN3qab2SEOwGP039bqJv7fN5XBoRH+eksleYmt3yS1Z7bbr
xusxr+szHZP57DcR21NoMHeav1gyoeYIJCA+pyvXKzksJYN9zTR5YrdXdGjfPkPIJ28KfpbJiszt
uQWqbtAxyMoMC6DiFnuHLIIJK+MS/qyhz2DG0R4b9CKR3CBUqpuvGsqdXswLen8eA0/H9Nm2AgW2
lvF2qmzW3xIdyW7AiX5QLVgBO49fv5I/nbhginc5+aquuZKnfa8mcDXb1RoOG8zPpbKJaJ/SMLGY
iwLre6jva2XL9wC83gDangqoofXffwws9iQ8bcjFK2TL8EgTHACo45MGj4K27BBU3wlrpFQ71HKR
H4Hq4AORbmRt40kDHL6PDmKF9QJV68nqh2PKFHHNxvtCiAllB/7/liLwFx2lUULFCCk05auCL8xK
Rk/OesZsluXFc6WDmNVT6Putzq1NwK+zo4bc9Xt4POjf3PUuPX7IiXPAOhen8w8e3a2AMn37cX9N
NTC2ka8/ZwllEy2jA50u8PVjOixxBbO/6eKqINxha7z83sp07PLfUN12yT+Qbii3NElKGygvcotQ
5ginZIYG/OSmIvFa6vUx1KhCSSbo1iic7+kMd//DSqgwvdtvZ5zAZyghf8f9YwdrpNHGn35YJk17
r5Udvm8uqfyYpMgxwbUtJmBhnYU4M6cIiTV/W9Uhx0Igu5xVSaVGZx92fAdVE33wYDF2zx0GT2vD
j1niYdcCacfwXt/L38+m8ySCHW8AOXSkPc/Yp3GrY43q8qS8wiHoAocv2mvWa6ckeQNc0w9IuNOT
iB9uoXQcp9Co+5yt2IvsJ8DkTf75LitLWJfTqa0PoaKq/vNj9YkrevJwr8um5ebZk2Ups5t7bntq
FB0fQOdzdhQW5tHXAzeP4r/RCNkgfjlJWblzsG+93HJNCdQSgwhdjpHfzapNJJ2Il061byNkKQlV
4PVTWN1SqzR1n7x/NuiInXnU3N+Ik343CRpZLC5hOFgEgP4/mNELISlaLY67glgDjpVMI2iBVp8P
rIJsoFrO4au349TCJfA6h8Y3Dza1Qm34eHIQFNI0mhFPwToa+DmKosfFxwkX81vM6t1gb10r7Z74
iPoNNuiw2+9lvQzBR35LyGQ+E+hpc9ciDIxFppKJZEAXsVYByc3BGzlog7f8UrtvoQBQSCkWMUcj
+yM4Dm+EVnL8arqr5H9RhxYLNMg8HermelhVvSO2hiJuv1jM6PNS+62YGvfZ5FkUBHqi5uXQpprn
HXrk15hGiSC6Ttfs9+Z2Ooh10L0XdtcNYn38e2cT7oohjQlx8Ew/kQ+CemGdFPRDWSd/n4pEG7LH
HuLdzFEuU+CYpQUtGImkEC0qd7Ncl1ViUq1CMSJHspfk5NrJwut3fNAbAlNU2kcYLMGWkFxpk7rM
mKMNg14QtaALyU+nKHDMcSnKzjxrOIXsyn24rgmIHaXihoHqUi73cUWOa/FyhHRhTcJMSmSFjiYi
A7NZ6/ieDcITDgVo21+5k6p9SzEtR0/tAPdpqAyXVyYTqtISJUunjpLGOEY6XPySxUAtLoy1CCMf
SCVK3KSoR/1arl2yZaNpocDHwWFrFx7mrdd0mBg+6zkjEI+FSDt5MMftQ238GmYys46JjgJIg7Xg
856yxxxbzlk0haoRha9NzubbCnVS9biK80zQsHUqyujKjHYCh6xHpryqLwIOWfDEWcVr8kBm2Wy8
hn6xAzeS6cca4/KhRK5jrjT+rjtv3JbWJtPi8n3pjuePEbkJIKKgx7lA/m9x5uYP84+2nZDZi+g4
SgEcG50XIwe2d7rrCp07yoAAA40ced/IrVlJFaHcVXst3v9kka3AHR78oqw8gKfAKR2xkuWiIJBW
c5tuqLjsgc06/RemCyvbwxV+ojtfKzwQlgp+ETccaY74BBrRkz8uAUxBhGprdski4yL4iedLg8A5
Zv/O2Jb5QPDiSqtQoCjDTegCwF7xHBd41JO7hH3+RpvEmVXdBeBGQp4Rza4KTPQv3Xw7djUwDh5j
hVZ3ZVDJkYapUaX7WA5wbWQWmKxQ7EDHo7NhMG5tRnRTtt/4ZIc+Zchf9BQBRaNVs5HB4EnUBgdT
f4tzUqAD2UWc8AYzxhT2ELg++Cq4mGw0BU0v/66e3xbu/3cuEjb2ch4M+hTg/8QEHGh/y82MVSjV
2OVg0sUNNZm/W4WyyLM2gPAHD6NwFf57diVrh2wHnDV319p/x/hDucc7D/0NOGqVlQU6KOT/PBX3
3bqr57j+2arhh4oYwJ2mYk2pCV0lZwNlm9qzWu0ajWjCR3P4+WkJkyM7ghzfxBvScnV8f2jtkTby
+RyGUnvJhTmfkdCv4ywN0ygyxxmvzsu+YtRT1n0hksZsI0PvwOmOsP8sEoK5s3CXM41ON/Z834kq
XS+QcGwXxefoznSr8mOPOs1b2pa4I4B+cIIQtGBFJNqgDpqm9eJnk9F5VkAwCmoQNK9XeHcKe1n7
TVautb4EwN6drkOIiM5rm+yPXZc0flHxgOssdhGPnL72LyMGggGQZHm+CAjQ7FES/N9clkeylwIu
zvUzVk87UrWioDMrCyAC1izIYNMGwudhZCSs2rKEQETIiEqZmNBNI+O8T2Z4hBnqP/oAw8uqPt/f
nFn5sLTLZ3N2aGU9vkDTXNsfAI3JN5I6doq5uEq90bQAIjsZdeawR5DWJihFQ7PQABbc1W0C8Qvd
yCFe+xBTCedrj8lNIvCHwKyS76YBuU9wA/ke+S0HmiJk3YJ0dTmqxmVX+zzpUoTGWGJxOj80k4+a
12/EkPsxhM96wgBSpOoRb9sL3Y8zHB1b3nlTBJBj5H8CjQi1VMyvfaOQ8FPNPvYOGh9sJ8i3ltzd
VDgOkaLrNkVGJzNzr1/qL9NQE+sDT9onubqPr4ZP1zOcL6L+M/BQPz+XekOwgXwjmlXV5vVm347I
UBQOXS8lCdf18EgqL3o8Aq5EOme9eTkah0cLtDJWRhyYGPy7CMYGON0GWT6Ot4wof1g8UR8VL9er
aT/RXk2vgIVn94tEMMoDsrtaZvhjhmJIcLlzmKhs8mEKKalix8aj6KNk5BiiUZktUOzPFzDwzJqE
cCxNKz9NN0q+JBj5j5HVRDmfqkxKfd3QDZzWwBF1Fxdbs+2usSBVT9hducw9LMNv/c3D3tCBexhm
uLYn3Gt+SLKpn66SrlTuBWVqCP1bNC8kQOZqME+JYIgXfEsTzaSbYLxBWUdjKHN8l9nwto1cLcqw
NW55SAOA9fpTSlZ8lpd2WzSHjTRwneUc1ZKhIsCxAg/MhCtGPespPqCrXTY9+IfcL8M04Ioa0BHl
A3uXkaw+iEg5VRJaTL8QZSkTI8Af3U0GaU4sJ9bGU6sBkUT/Agb4A246cZnvXwkuwek92s42sMKP
fQg5XO5phtH9v0KGy03dX4NuentwLfknsvVtVvzK8rdH3JV754+TiWsXp+a5WJlZzOt1f82Ns0r3
X0/szJLWdnZ4OpHZmqNLCWNQ2K+CK/K6uGU3mcvT7Upiu5XYI6mSh3HzSxxr21gLjM7d4DIohxCt
JJAh8m/VYp9gXYahGSSVbd0/danOyKYV9vEdWdg6e4YWWdCLjP5lXwzvGe6p5q3OAZ3X6ZgHzIUs
Z3YFChyT5ZQaLVgoca9/ZUxBhLXdGBiV4nIK0HOnN+OYxjaXE/yl4bGu/7+dHEQVJcGt7sDS6KX6
lnzLakiiSCVAqS7xBpRk+zSfLGda7ecdSQnfw+4jD4dHs93Kz/Ce9U0sVfqXBO4eLYeOHp9ukjjP
iFFMWBzyDUts8/7AE3PHo/iXfs/Kdwv4EKJ7z/6/sOwVvijL84A27QqDVkLsSHSEEN1ngf8Xq2f2
G2Ize41T9vkfPqmZgN4+6pIVqNppHR7MdenYlaX9NUFcb/Mmi3Kqmrd1+MO5E3MF3XgGFVuK8/rG
YBeK1JqbCDS7qEuNUtvaLIUS0SWF6eBBDGoPDPcH2fSSN1ISR80cd5AQOElDfOc+Bi5aFOyn+H1i
s8t25MWiy0wBvSpE4p06qJC1ccewWo1VgpMbqCcqXMDTg7lPOdcDyOsymZjBeiLL/lJcOm+i8FL8
+PxnHaNqtEylO/wqNT7zE+lXeEVaQAVv12yYukLojOS3VELTUpbbnbfi8amlksi6NBUx5GpTBfKC
G7nOzCK3p7nO+2kh6QtxnxHAmForC7O8TjQahx00vUIPZHmGDWGe4e7fjwOoTqVQP272it8G447z
UOZyVWwx/hnWawmu6AqHWaUTEx2LvURqlzaCbaCLaP2KyFLjkm7w0jK2CNlPVi7j5zWxrNjESb9J
JaD/0hGZHZAaWOy7/ZDsVncoaopc6AeM9ZXzgtyOIo04Jwl8G2J0JERbs6iIcWwTBQeSpt+5CYCP
r661yjxPYXjLEh+Nk/925o97D3zAUCTcdCJlpRUMiATP9QxQchm0v/l+xw5f+dQTONeTIGHptshu
d/k0nmI5N+kMobeTaUb9cbL+w3SC1pzHpdYVU79lNJ0x/fXvW86JkXNMsv5tldkSVVdebqY841rU
BuTe8Waom43JBBjG/sSF+odTM3vi+j9SmlKVxxG/s1R+VxcZmupRXq15dUkeAT8xsxBMla2o1El0
OMxPu4QJwkTnB1o/1Fg50PlTUyNq6Doq/pRZ9m5llUrT/0OG8k0luOAIdWhpKrylLkOwJdupBncq
UYSuZFKaaYoEE8HG5Oa9QHjDbZahk0OZnlkq7GaNCw1G9JoLvMeI4SInUVQXV9Zw3jKPttOk59ZF
ZhpD+gq5FBJDYWLXVQKEC/07nKOZeBCXsWaKGWvDSQloMNhYzTf5TlmuSk8u0FsV5QRkYtKutW95
/Y83PjTVI6M5JFxxqcPqxLwPYw39z5AT9rwI414RTLkZ5OuNF75zlhIrBPiy7+KAo1tf+LcurBc4
Tzb0HelEc/tLF8Pq1BUxjZcsS0nvPtKmYusIi2i67FnNP6UxxyDT9JZ5qHRcU8iv262prZV9k2l6
t1k2X7jTljwQpZKW2Ua2ztnD9EzZivcBNc6H8uIeFPKKznQwXUwJp13zPrOB8K9WcsRdsnLYsfst
9q7pgWhucbvIn2AII8Sxyz0ZvH/NRPfLOF+Dmaz/rSCKxxagrNewe1etsDu5tPkfQDDH0c5bjp22
Hua22be9M/Ar7ed+13vQqThbhWMog6l/XwhhgYK+JpW5XevmGf+II6yJk2dIIYo/oBNDmhEOb/OR
FYMibABuFcPsSys/dcCr1hgrfgKshFnlmRKXCCF36Fh1tWHaxvjyvC0kInR7DP48PeXOeVqhnW1T
c7wghKgJoqpGu07GjQQW9j8BfI1xF+1ftQl6kyujWH5Uf5kj2aPtCxIoS/0HusFMJjmH6+KfYWwO
Nm28I8t7brwNEcwl3PTJeoyof+N6uVTQverL96EN644bYOGz6vu0be/if+VYaJayLSl1ss1HD5Rr
DtOyQDZ99QVyrco2OCpHRM6X/0De3JtubmVzeUNPFXUbgSBdJOA8Bk4vll9t5uhE2rdAv7M6oyrb
cmeIH5+mqOVDVrg+e6TKLrXC1NYFvi5O37zbg2/dhoPOVToByFd4HwusfoYYxCej1AUha9pCCT68
5JRvnNuzgge2vzxkphhxxaG1clBTJCK7hBQjFFMnHTvZNjyCF4bhJDD7IUE5g6avJUQTOcs3rWGC
1Y7h+BhoP497qnjg57zlbYJJ8HOxNny6HuONPnIRPAqTy/21wZ3htVodhADdG2rEcaZtT0o8VeRp
KgMDXclfRFhsYiG6pbN7/9KgCqLlFXNSj4k9QfyNeXS/JE9okTjNgqDobcN1PbmTrLIadsMDO8Ph
TaEGcLCgXcygFkrWYzPpF2FXRHaBj0lvu3BrYVDjNiHl/fyih+wBjRmKc4ByNgPWbrThwcBePhcC
Smfs7HxmONx/L2OCvM6fdiX5uOqlH9spGj7veMeD5KOkQoqlPj4nUn1t4f+EeE7CeiHYQnz4kp/T
Qnd6bxDeOi63krSudRsd3ktHzd05vheKgl0mCNjbM15bVNnBMcn90jpJzwxD/NlLXsCsY45qbw8l
zie2cGdO58Xs7RHqTXAbAMin4pAhV5u2X//431kYlvWGkRdDrLwOuUdluVnmEZvamP+xpNggih5e
jPwJm99vi7jfzL7Tv5H7wjYdP0/gCGf6EdHyEnscMsNFYCQz4nQ/SbX/SK3at0J+v4GsBUyKqAoK
dT7HION4AEvQDbKrc/bfYAy068Lnpsk/AxF/kkZ+KGmoZ1E5fb8jTo05ns1/JlfK1tsUQBgwHiSH
R6PA0fDGeTMCLDVfVpNcPMEDrD6aYEh9N19UHyzS86uaMtjNVDJaUJMFWXitFkS8ZiyNxNUOx4NT
6Kcw5AXwVDIKEi+H39frNm4JsE37MYeSJEHF84x6CBdNGuDXRHx6oaJS06Cx3ETWUz7923id/Xhe
PDhVlypb4OxuSAFw+4Gq5/adaj2+PqJii2QiND8WG/uiImS2n42/0iz3S6yEdZ1gKJ0Pq1PaLuJM
DYYVn0qKyrCw8+nBqDeodEPPQpRkvdFi8rdif3qGbUKLTVX8H1mdotuz9sBn9Yud80iJTYg1b7pN
9EsmPKV3V3xsxspIe27WgR2MtA5r2WbG6g26qou7o1PrxvZvwbDi0j7mmVRst579QSww1dDgh4iw
Lo+D3WGlRA1SEWtP+doOglE9z+C928RYGVVpQLDMapDBYvpxxs2nHUsuUD0R9yWy/I5QVahtQ/2h
At+5EzNY1o2hXZ0+wEZEQ8Uf+Gc8TOT3G5A2lqAy9CjZTPs8dg/QD68YK+IbkItiJbCYe9a1frXy
2z9NIYSLNM+ibJvPZqy3RSF8D/RMkQ4p8LLowF/oBAPXMSSxg6652H5SZfIRArKUdDIaLaHNvIvN
ycRnmCP5ssoA5pOOvTOpZLRx/EW3xLyp5nl3GIJY5lb9hLSaHq5EefRGRx7F8fegfvj382+DhgcP
TkzR8edzeap2J/WDIIqEosa463kD6XPihVkxo5vIOdYGQ0WsR9eTURGjCkuEKIh7jl9WFRIV19AW
upNfdqVGCTu7MOac85s57iahZA5cG5MyP5M8OvXF3yB4iiEXtZpcNWmUjfKnFqFmrlvFDKWu92nn
xIUcgXQvbOgtIrQsCQdYsts3WwHQoHkz8+Uhy6vng1zLillph8ZCH8XAw9/h/yTIc5+iqjlyXuNZ
26ZeNM3ClOTt44bqfnGClO+wMTVfJ/E+FqcWs8aVduTYgYCNlAv2aCTI2vxs3nsUYJ+R1RXcIYPY
zmIyIGw7Z2pL6rltTHC3Aobn+Nthbwb/Pr/0NhsIKKb75OA3X2VzzGe2yrbNVVEU1G1Ong1g/3qd
iXueVRKrel25HFxbxRKxKTtJ0yfYXacv6nDAat3l+j/ZjSr03qovU/taNdx+nJb7Y6zpsnDE8xwF
f33zrvnN/roNPTmG0m1tXVNHHnqnherNQQQFxqerhWCwOnwHaA5NuvZ9bpEpAn5igwMDx1DaLZgS
iqVtUpURxc+dvdtV4QGIkyYcEqUH+rUTFsyvRZQloUsfdCfwhHKBYvLCtrYeQPL/2eQfvSjxKuFe
vJWdpvmRSy3N/wCChKX+FkRozGQHBu9P1MXC7WEXvNq4y77y3idx0mFjZX5Qw5M+uBz3NKaI6B+t
mc4ox9u6c6LX2d9DtvX7a/Og/bGN/qfl9FMpfRHkKp6jNIAoqJguYSQ7RFrIRZPkgDAWoNz1XbL9
VE2ymOuIcY3INDX9nx6OCYcHQR0lsSillWqjs/MvPNSDhbtUzdv/85HuGnGQtDMCDmZBHs8zy2Ga
CPauE5WGwjA+apkndV0GWmBA199fyu+TRADhR5ffLLXRMrpM+3AgGaZzYnnW/oApAsOWddH2+IZt
H7qlTD3Ye+MWvE3YAiWG+LzLeOSju7/WbdEh2MpceF4LNRVpBYkCoRxMdsvvLw+Q6dOTkhuHaZqD
2LGWFNOsEwfi54iFKZlts8nY6/QViK26gjotaTc4sAmKa5I69ECK9P5jmF3DLlGB6pt7lg8oGG9Q
kXTnX8kXhXMEcZvqGjnejSPavkAVzNMD6E1STCLObcPzwd9E7f3I3JIQBnr7buaX/1seL3Yi5PwZ
s92anGbcc33GlgRS+8aQvUSmPWxwzHmfHraWAzf7rYCdYjl+SAyOfKEkd3Qg3YUeUnwCUKVUUiRP
8Pv7qkt2iLikUx/VcNE5FSGiMDUW/S+RAqBTzNIUuuzJDdDQK8+zOiz1sw00dqKQzP4qVOEzeHW4
XnHpp215I8o+oK+FPElb97aBlbj0wEZ97XnCYdryRIiQH54mxRHK5zHZCJmqYPnCONchI3hlRDN3
UrrCWjoMyBbXuSibG0hMZQaflbZVTbcYrWAVg9NJ8pW3FW32BPVG8BsGNzc1CbW5teDWI6qCfvLA
HpADFV8lQTEg8v5XXBruCcErz3+KC5hWquLCZRBhP+lCAX+pNlMa0qVNjj0R383R5hs5kHDSdvxH
SsYJcM+GFw6vp1/4LZSb40hjY3B362IyRGtaKGRByAUZv1jtiT43EuxJD8pZ941hfS83eCan27ka
+9HT7NTe4uXrFqWiTFqaH3b5mONTMbiINSZhrtjlSv2mcdWGSicT+ivpej8NXjeEEzg9WTnCZbae
y1MIOg6P/gfuq06uKwFHL6YpYFNIFvBdvYvqobo6Lvcct66H92zOraprwu4bM638kJI7cECnO8Gf
d+8hV4bLAvt1JCB07taWg03hrn6iDYxojwaDvwZtUG4gZ4268VnAyhfmKQok/YtU2L3L8p38xc1s
pDR4pPHD/UoF4LNrWouwPX/+1V8PzLmHY/uTft4mpSM2sWmA0DV5d+qkd4WYkeJqYsj++VVT0E6T
rXAbcsVoQjFbDo9eSlTvU2HPMCi2DIhXJIzBi+x3z1Xe2uMKpVvNTPlncL9E0w2M4eMCPlpDfFbm
cWXhDYqh5WTWAp3QjiC5uHlgqJc4tzLiZfdsAss4CzIlwDRUp1YpytZJRfy4c0OIEk/JCe06kIax
suUrRye3TgyD4M0hCfA4C66wDfNs13JUxRrG3gaWz2N9yi4Jk/3k+/1ErDIe0gSxmufHO7kLJsq2
Pzz0h9mbgEbP1cr9W8BV14+fNT+M7M/7T07Imo0zhzf8gUKaQZcyibgWSshDX9I5oU2WDa1AUY3w
uR8xC6PPFGVjgJQfd1PZ+e5ckHjDqlCq4nJN8KvVqXZVdfp2TlZS+jx2vWrPHQNF7JtAZeko/+49
R78wsGDdMHXtmsW5Hvv7Cb3BvlZQ1YhMp5uSf/Svbg0JLkEgmIjbc9ziVSjUpJYG10+B3wCyGKJG
D2khLBbRDjmPC8XQqEc+xKuIGGNVF0ar3t8UXo9GxOabLtUvOCHWRc2drngeUUYfIIKxlYu6L6MY
XwoORU5r51hv5tME/ejGFEJhjXeXOLwqC2++KuUE/4A6XKQIWjffUlNDrCtlkK1lgNIdf5aTmnEb
IrtcyUcqmzY3V6HlkI90hEFBMjq6PF7+cKwW3rPHAZ2j0rxTEpzBbRcGL5jsvsOJ5puPIO11BwRq
wztJASz+YYJ355oYPrqHPh2Yxr0+mCQLSf4EF3lm+Ktg2Ok5Pgm5tucqyWMsD1ptF8xkM1hLF+Hd
opkDfhBEDyRspmTb1Iq/I0d0BA4THDgcjEV4hSTx8NCWFi+pupxennLnKfXiIHh5Z1iIGH5s3Uc1
13miRC43QtmxMSOWUhWcTEfOsJ/Qg4/XYyS/k2Uy/blRDHpkeGRg4bJdONvQWU5bwMrlXkYwo8zu
c0gJLhO6J/D7aM8WtT5+eQ4BinW/FA5uWqOdtHl9QcICfVTRh1nDWRqQvKBmPaSDT8wo6Q/QudBV
fEqi5uhnsArTe1bhOH3Ki3sOjAEMXaod+Fsk58YQ3Ph6kQhahCAZrIEIi03el3QnmoY5Ie8Gtswd
rVk1uWFEtpAecSD9Pg4fX8PjSlEJNMzBw/5EIV07ecJcaE90aARCDYK37AUEWQBvp+HCzrdt26Ch
fbiIGHvIYPbx/P2JVbfaMBAH4xqXoDU8hPsbNs0CBr15bVjeI2hOybYcPPNOwTLc2UW0t+gQdqTw
chBYk/SjqdmZPS8JhC6O5UQHuUJajwmvNcItVZZgK6oQuJ9vIANB9T+Ig0y3GLGG/wF7VhyAfVyj
AG+UvTF9N+WHAIfbvJlzKjejYsnu9GdthB3sGpWvvHkiBfHlmQHf7ULiYEMjsLe/sSYKckknb91t
nCtAvDs/iKvefVxwUrTNnWPZIJ6nNdvayng0Pm5lWzHpXQ18uxuZu/0HPHtkbpb4xQeIBoxb40Wi
20TCLaYQEYpiI9JFlTSPCP9V6j/L6BYc/JIasxX+ksJrYgy9xlSU7UBc8Y/0h8cWhjti5T0gvGrr
2D0rxQWh0Ad4WDEXL+Xz3m9NaTRTcwaZIZEHELCXGuhqQKNAZSvXVaWUHuXpJZWoJJuGet0ud94R
8w+qBwqqflpcWDjSFHGpia4KO4jdy/bU1HC5RkVYx7S5OpyUpuBXmPYgRU3jO/Y8oD0ZcrcOO9zV
K36OiAR4JI0FMi0fkcB9Qg8/PlRi7z9Hd5dWcQUTm62zfYkm0YIKeyPYT33QPp/imV/jSH14NY9y
u2Tv93bsS+VHdSezqtZEvTG+ey0sLoLkEpv0TzPRqkRGgpFCDFzpjN/OYGHL+ud7tYg1Vbrpl25f
62Thr97Ju6lfsPGFJ/utEuh7OMnp68Dz3QGljGIkEanT60d/90V9icnmuJ4B0WKtTfa1GX7EuUL3
IxkSBS6m9pB4bKGAJvKyCIBeCIoms0Ak50dw4e9ziKF82cTnlGU7vhtEOB++MVOse5H8wuL5Fa33
gXNj9/AOZAY2jVcAXiRj+BROkvdGFrsZ0teOzwAbpzi3+rozY3PIZENs+75ov9MSaFIszC+KCsrp
P5Rz8DbQOSXpoX6KoYoNaLe/lBBDFHV+l7LB+ko6sMmcw4Ha+epv9SwIg6Dl+SkK9DWhMwRmdzRM
GM8PbqjCMDCRqAoZdlCuhIQSHmS4xqZHs+zWXj6BlfFcWjKmq/TpVFb/alrwE9s2yGZprTcGpK+D
HZfPFhxM5RGssywRNu/APVHYOHg/h+i4GCu1pI4j12jU1nR1jvKy7U4b1sc8/kZlq4hLcHEjgNJq
rmJ4EEodSncxdS9VqDt2GHLTWjS9PN8arImwePs+8as2VQ0W1eF5slOVgqzqSU5/02kYLNJ4r6uM
xjQMuYCdtDTTUKIFDPCRZZc7QLYqQjOmezMUVYX1HGv+Ye0wZMItxAJ4xA3scSVQ0zAbDbZKN6+L
5g6IfvTu6EI9UV2HmGW1CcB9ap4rArP4H+uCrM5C1va0FkgRgk1NVwtfUaL90qCEEpexGytMZhxX
P2t+GpkEsym70FanhG/X2D9MgZU04BCSqGWtYcGkku6UCIUgIBcXOBioxrxEEz5vmy6lLW+HgK/7
TYEkSVVIY2s+uH/GhHsw2hiAxjb3oRcSrNLSbbuARYtqzPP9uWM157mkzBWzvcGzIqzlYlkK1Wwz
3+WYYf0D7OM6UBsoWOchBAdPYuFp9isDMOPhh1BUO2/i7WMJC//MbKlqWFuDFPTQudPl57beEQKK
Y5ioYhlsAh/xFOYFlixo7bywxZ7K8EFcxDbcLfbTKWRdHIVLgboWGq8DtHuj3RQ08tqspQkV1B7E
oog11+gtYX3PXoSKw8agLFcjo+1CUK5+ZLEaKZ6v4ie5FIoVvo6EtulBn5Xjo45GF8AjH64yh55W
2L+GDDw1vb77kOjypq7Yvl/B0phUmiXQ4wQJ3dysjgKFeD7YF20XCGKASoP7vRBh6B+JGTUDbs9P
C7jxKDJW4Luy5QP6DyZLGYGiNATlM1A2uJ8MgZnR2n3aiqB5omdFd7LIv8q6TZPviFZXGkUlAI20
gwIVjZ1iiXbK3Sfie8N1nOSePgyGOzDZFai/TFFq4c0MBaQhhgKYYJfWh4xwaoFdsydR68kF9Vj/
9g7bjcrUx4wlAfEECqocojLQ7DJLOOLJ/4+tayLP00PIFXaClu5tpFIh4jfon8WbC8JpXl/FcQkt
5Ats4kw3SXSVeVI/NNjlZGJXD8m6iFFNqQ57Lp0WzGHay7ESBwi5w0pt0ObwWMwIeQVC/i9nYwnr
J3Pilvj/5CdAXo/wxEc7hnCJvtWI5DxQW6ilgaSXjS1JEd8jDMr9FXt7Ry6TDfnRYo3o4kRWQUjo
74U1mEgCYgG3z20Ut14TQ+kvJPzPxZSjoPQhjuGil+He8aeQmqGIXYyZp40gbPmKD6KwucvNjaaw
b+NG2WCXo13etU7pq62HEiY1IkiFjcoSwv39eI6fdU1ARGG6Pv8bE54ON5mdQ6UJD2fcHUnwixX/
75dmnklVhlMr4QMMEPGR5ECuG8Im//PN0ADQq1L8z2cYPFhc6k2gNPTxAQWAOUy7eXLinscn/jNs
sS1Hk/mzcY8wCUa+p470aYdFVgdeXXMQecta/9vzEaNCJZsI0AFG5lnh3Vgh4MzKWSa+Lk6dqSPS
skt1M7cE9W7vzc71g0uismivrfmyuhrHKpaNu90iTbm/rEmgG72VlNJwDbWRIEK8LFsCE800Dbfj
lrUoGrdKzVWQkjHsIrj7spIJBX3wQjP657EnojS9va6a+jjostJAKQY174qAPNKCnfJ/hbGx5aEK
JHi1WqLE2dkJ2xT2YHzzi6F1cvI7PufY624XE8Q/x50LcUEby5+H87zlRf6kdKQspcN5CXdcj1GV
8zxzemMi0Wi5QG8dPKyqJvBcwA5uwc36/VFLI4m3QRjJ6QQXjpk87U3Crq6guQyigOmASuaTQoeC
f3/dcDug5Ia+jkJv85gXHrvsSEk5fISSq+VF0Ih97Hou4JM6nEZUlJpA9jAEb142ex9fT/CnnP1q
iC12u5uv/Rie81eHkBoaMciDtrdSeBr8CbD22IvLBnMtKPMNRWXq7hvtAFZD+SOSuNwoSf3q7DCq
zVYqfe+Two1kDV0Ift0WKS6sjWzNQqCd5Cjq/qMwLEj1gTvFsxmXpFNNml2mWp2NYpKso9+YYrdL
7YKJXaPfviEJwa9tx2zNAXLoqP0akocFLLD7OXcFklcqnb9SSZOG+B0i8g29mzbZ3PffdHzYQZz+
JEuBfqv0gXzowwzpe84hPPq/RxL4otEhwomAFH/GFXBbibCc1ms+UXtuKEsYsMBNSHPEsqEYb1uT
YL1eHNPaK1IGWYZFzGbjZ+JJoP3eEFWHzMEugs0xVzzicEEq3WykZLni0uPvcHq0RfBBk8SxuFnC
Drr/M+3CtfoLM0bdyUhssnJQbqvHpSGglQKpjSvtWR1iTDhIqcf/5aG9XiJqjkcJIqx7VTLlpr2d
iEdDOqJtQaE3DB2qiT5GtZrn0eodGPy/20sAGYDwl2/n9NNr2LiaqTrhkHEOPrOQ/iDkLBBqc0Zz
OkJaBfJCTQVfAP4MQlH+c3u+DE42vHBJReNOXr4vnMOGpJeQBIJEO5yxIcST9+yUCEafqMm36j21
49CgZwKu+zCzDXfwL8fY+LMl+kS9nkyFM2jFY/JUKi+T+MuzV67zbaoTQxVwZx8GR9jw9eUTZJuK
2JO4hV/0Ng09DQWAry61sVnFg0qbWG/Dm6ffUU/fLx2XXd5c48J47pzTYm6ev6ZQRHbwqeeUApea
3KStGkxc9bNxunhYh0xR1hroZCqepUuI6+uekLOpFHZOWLensNvSU6Y4lYT3tKEoiHHUBc/s6t6M
HQWS+T4DOvZfDWDjvYq8wbaSTvj2PMnq32bfqYWA63ld/jsBPmHIqpasdi6BfjlYww7kgV4LpnWl
chdOemhPDGJoVaixQKd2I4wYh4mjECqFFdTUNtuXVUFY1SyBorG1lBNrf+fHGSTwmC54oyOC23DI
xq7Q+pfzROI4kwG8acCH6Fc4+efv1M6PmtIZ9X6l75cISJHXcZVOGDhoEKpvRtPQqrP50SVumEDW
Qy581MzURX9T/LS10VL2oLPNBhwwTQD7RjI2eI/r+4Agp6Yx6mn4He0qQFU/veLdr0KbNo1cj2jK
o9ZXpYsTxGdGpgLXIbFauBcga99bbpM16NbBaf/w+P7ifKx2At9ILT9PfN6dj3z4/d3gYRdG139r
rrKGl4R4Uue/atfJve0rA8Vt2AIttD+wH2rbinl2cgSdxezh8dMBMoLdFARz/XeoGEMHeT8t6X9C
054ODb+X5QOfqTLbThgaLAglFgmwowcEVh96GFKyV/PzHT4qTzF1V/iapfQesatxU5YPxbZE8pb3
P7JVo4cCCYNnslTpc7lbAAd77DekNiHZrrL+mlYiuWHw8jWhWngmBHUQ7rQry8hjgstSNmhxnWTb
JSCbJD4s8df3Vd6MQmeSs9BGpFjjxAscNpGB8y+ktaim2kx5pKdkohMsrGSgbYHERYZ6dNJVAH4d
SSp1vHmkhrN44IsuJ0c32A9wLzc+4/VDSx5JsMf33IYxAHIxzay/R5/e53FMWFbuJoWkFCDN/K7U
zj1iS53N2XEkb4q20HAP22mwNDRauUAaM2NO6Jt6Xf/thVPjB9He1/M/fPhHkAbHr7fzDRnNxBgf
fv48K8sVgzmOEE7YD+Bu9C2upERbCihPHF6aGmD7qRIXEsm1ACfOdjX4nTxGJV1ZNezeKE9qxn3V
QTySinRgox9neMlZiI7LLzZgqSpC/gvAtuBR8HECMdEJKlOPdI6q8HYJYLBbiLLCQCXWUqoIL8+h
9HJ4qlNKeqNI9BJGiYbd1wYngFYYdag1nGFQFuvfsbAEe5rd1/9BUpsj7uSVGEiSD/1Z9jt+5yx9
p3qAI7h04KGSBmrjCABzCVsTfbA/LP/KqZ+XbJ7ZacnFPgz/uZqOVn/CXBPdjpo/zaKMpg9iuGcA
7ONABHvx8Ho/oQh9HT1MktDMf/ztpNy8Tn/5yfM2OzX/UalB0KgWl9DQ2U+ZTSySvR0t+D+rXZea
Tfmm56u4Yhd2Q/Mf7mud5AWYOAQqsk8LxhfPBGUi8cMHXGannIiGS86uP24CDvzDtaBUeRf0qJMO
PGvD4MQdsCNKNqRv3xXOuuKilM30eqlnqdg8NsNpchY5dpG95e4INjSKXm0+ZOEjPteRwaoMCZCn
EMchu/k7+gAayLfOb3x75pvrlmmXvZxHwdZLbx9kQIV88ciz2DDH7Kdc9+cvD+FIT+yufaGNz5iU
vseQ/NUljbo290RTLA2vTprg6H4C9W51ZC/y4NtKy4EbEjpAjSvKnLzp6X/ZWRHoqmygi9ecj4IO
lFw92ZwmY44n4nLidB1PU71SWQDJcW8Ua3szTRYKsEQqBQkiN/jxVpo7BLENnInH+wUSjwPwbmr7
MkvoTG5rmHZCCNoJl+oXnDhKirFZEcwnt2HGjZuABhTaFntOgMdzGTQkvVwVLxO3P+95MYKyTLfc
7N24k6wntXLJoovIBYuuxbs2wL4+2XddoTxbfH4kpv0YKrjVBQhXxoUp8hi+mC4fE7UU7IZDI6Ky
cBWsARWbvAgS9Z3hlo3htDKTCC2bFXZaqMajzVtBiAd3tZ2fsxcdWWBkiJxTf8Gdg86cHxiYOTBD
bCd3A+KM3lNB8uJUu5i3p7AGj+liQE4zjRbwP35Gih1kivV96plpNWLHxoC1QisS0SvifQIuX/bD
Ygh/VsD3HhC1F/uZjSn4Qf8vGhxh/qPKtZwnBbPfs/dvgnOqUSlyrOqVEdrvnsyC/uGZXM7LIa92
immzmn1/XY/K6lQGXdP6KNX5q//q2FS6R6GArmhemf2tMnbn/waikUaVw6Ida7ZajmnsRigbUbaJ
CajPfCLQi1IC4cCAlc/tGg82B3NMIGbVyZUg5fvcnaLrIKSWQqSMGd7mh1WiD3e4wkLO4ptWxDOz
ywcQ+QCA03j53yqpS0iFVXjHywnP9BH0npNMW07vfI+b7Xm4NGRReoeGnSKav1AznVzx7IGu4CKb
hS6blbPpDCGMvuRtc/86zbYenC9Hs3zYga3OlmxtozPmd68N1XGIOwY3+eydNCcYR+a+dAzpci/+
eJ6Tl4KkDuQEuB1yTi0OL5EMPdmh3LGEr0PPm3E5x8SOl+72b2+M2t9YLiU9hemZDIXySap7XGer
gG/DHlVI6Pilxdrg5b5hmyAbiCstqbcWYDacCvbUaGUU3rPBv46VrDx5FYFRqTrKC+K5JJu9zMbi
E33+Z8WTm84iXDRHXBR3wTZP3lGhKqLJlHMdPWadNtmgF0ugmM8mba8/0GxzhuqUf8X+qdvqOUhy
qAO8Jwus3npBptSncw6EEkLoPSF7PGwhUO18yCZ4FsYSuAkMS65J6lSjIaPeNiAXxsp2784ZDmZc
bHmGdkb6jeQCtAtfIIYG1HIevEH8Xvlx28czDaK2cZ4PTT9syoRr402VK2jQRr4qTGSFDU48WP0I
upr6g4oZlxUgXnSkOlRADVdmg8RmuWJDneG6isLE1+cWbyeB1CfHPKlCV3Zx7gDbW+xE7+s/RDEK
IWQsFXMMXuB3hX6EoGjH1jG6Qtz05JWElYXfu7kqFBNmBd8H7U8ou/AT+VCKM/nKauLmYZtwu1Fu
0JtJvM4hvr/yc3BoQwerJJEzwDaTxwcM02Hu0Ixj7UDv1MTJQuHsxTSbjC3aBNnc0EKt8nZj5Nfa
eaJBPSyM8RX0CDRK/d0pLPk0R77LbnthoR1PhehRUvMwDJ0PkaiPe8+LrXUbE00YzXFXyR0Ak4rN
6AUgk0elaMttDIzqW4F1y2ZLNXDu8q1UNTK/7Pu4bpuPPJf2Cfwru+LBgVYhBmvpJ+GP7pDH/Bx3
SDXC0hNYqX9fuRQN4KKXfEB2l1ppuoOoCvKgdDsC9U2oVoqEzqTE+27blzX/lUZu0x1wTJxr0TzW
hdCSYiKFcgi/hUlCPvVo4RVXNhs/7KAUkz3QJi00m+hfLHTQL/7sb+oMu5PLpNGfGUzKjzF45Ump
FNbTv6pm3b+rct/7tSInJ2lT2pVJRB1rvWW2uA9lUIC1vx2wgGrMaIAH3JChiwjl4gedeLQ+5aXq
XFwC8pgT0JBC97Sg/MaeKijAkR+oMSvEDNwPjLSQsdV6oY3amNp0xwBsNydUxy1fI7PFI6JlvvZo
9MGh29vHp8dGYIkOLIFYiSNkUKNkc3Tl88U5z2YYTAg5UJo35BvuAW5c1zxTvxZR44cbokX80pqR
DaxxhUakngigRoy46DlQ1a0HVaLcClUjJcqCaEiudJiUR2ULFBNloEmz6bPi+M2/wSkjzjn71VV0
nXJfsPFYZRWgSMXBWD1Kl2/F8yvvY/Tq1dX6sdnU2QgyQuUMWx7u9Nu5oNIe4S0YMWiLcRZrAuXp
N+vp4q5L5GT0MaNTsylDH8h4yBf+WROcnK7kpG9YLTuvpYfh2vxD0FmwIelN0mjwbdyl+onsdDSv
WWYAvXQfmqW1M8MJqemiw2EUGw2WpqPRzHZk7iH5ysTU23QFBL1owtUjj13gWeGm+LLKrz8PQBq5
yNoC+4WX8yoScWlX0BfcdXOGZUUm47Ddy3WUlApZU8oTtO5Xx79heb/GKRnqzHu8By4fQ91H/9YN
ysVygxnGkS6MKFl21BfXBQ0CVFyW7sblU956kO1/OF8RmnAKUCPhRuIz0sDgr8uKnBK7ciWwKAd8
fOvZOStyMnKwL4AGPrJuC3IlRfRPJSd59N9IhZ1A7vxC4rA9J5recU5PsiszGZ2mol9opjpZ3kBE
7GuBmu71CASgnN3vv06rmqqNKVDHsWzmNl4Gb3GhSBU3QNNjK+zZlJR1fAAHokyOxS1l89wSHShV
7FUyEMPg4WecC1qVhT6DUzRZ6Oq5/DBcr0DC9c7ck5kOkuLNJljydrWy8SNoyxKE1bmlmd8McvAG
wgiEaf0fKVN7pDTgDoIol24+MmQkcE7dmbWrIKSbhTxl1j/ZMof+BKpHxCVxK9RgMuCObC4hS4/t
CKCMHtHcGxYm65UFCHgQIls9SnXln6Sk9RiT8gBTwJxCdKoArT+c5nyA+Z/vx7hZ8kMirXkOmepc
2ndpWkn/kz3uOGmhKEgUzC/XABW+ETa23aNFgg3UdqNRl/cMivMEbt99SN6QefN7ry/Qp22lubsD
7E4MnxY0GyCzWMViJjBSZ08y/obJXsUXaU5YvaHLpxDuZkBJ9FcTUz2IUnAoiNEvDMk+kT/3sOxM
QoHF5rDuCKOPj2AYSYZ4TH7i8zMN8g8WeNTX0Eij5XkEVLZxKnJzd/0cHIw8XK5jY04jkZiun+qW
NelHSboLFzShZrpaT4mDk+h+WA//E0CVVHA7MH/Us3C/wkJf31kdvqR/QBT4z2NihtwFgU2zPi4I
bk37MTpA9ZKc7R9c9G9bO5WhQKWxSyr/STFUzCw73JvWHpclw/Ep65l7Am0HRdYRG1GJ8Ha8JSdy
TwW20N6Or/Uu52Fmwwjf+OiLoWTm8KJW52Qg4xO1oBJVfGUZd5oSdm6c9rB7nqHcUwOBXxGTBbwE
OZJfbAJyqNhCxtUTGZsxo7TwzUkOaCoJPx8KmppdPxuwKEqg3lIhcwLmirTO2+XxR8N8wt/hhiAq
fh6SlCy9gYxcBK7C8WNpT5MXZUw8vE1k1dJD/UoCHATTXutZMOpMLDCOZKEJ14P3utlwAdJIHxx1
orn6CfEIwaiOC3bObuQMUqH5wILQaxJ2Mwp3zE5lFs2XoC1/ycz+1j6oLZPmvGXdwxRF2vl51nNi
fJ4YCR+NIAyb4btLK3twNC1euLmRAM+jeNGU5znhjv4TRI5RqSwiLjIVKspK2JBJV+fDaZS2HZF7
JS/Pw51jJKmLuHe5pL7DaTi4lkPP0MxufbK8McJwBIWLI7arLHgdJTpNheaXh6TwseZVkqtVj2dJ
28Ipz2yoq6XbskJg3KEUU74QkF3r+1HuUXCf/qyF5RxK6+hvb7dgRdgR337gSdJ6sewtq6AieAy8
/TfXp5jZ82/y5vDy2fXST3CudUuEgZ4wXwSWBNM993UUdGs5wogjjWf0fFl2N3tcdM5y/8DiX2Zz
y0NlRdIbVeRbp/GPlQPrjmlc+vf1u/DIgkekHzlx98kWIq0P2VEQHwNdDeGROXR2VMXB+j7G2VRa
7fh+3S5tOXdJxdK87z/zKGH8u5sw4/BZcj7ujztaCtn2N83GzBrlG+LLO/AVC5asZRp5iaaa3lLf
Udd+4WWceXi/DMXmQe1f9yWnNY09gfyewEP8Gut0P7edxLVvZ5iR7tgUOgaHmjeM8Aq9X1jpk5BV
NKkL8kmP1AmBD9+obB3J7p7C7N3UnsESbY9iOYwRydeIVRfK+scMoYsF4bn5yfPGdQ3lCxSoXFiH
6jvu/k4kkJ+RmVpk3ViTnWC2ttHnx2hs5QdzLGtQKveJoQMLzUhLRdFYB4vTizI6Gge+2Ee+h35Q
aR5pRT8nkbDnsYy+7Wde+SHGOOVxpbKMqgFKQ95qO7EQIC3xGh/u9Y8G/RJsbYAKLnErfLCfpzPB
lda6XqR6FeSkpUqcWQbVu4SUoY4oyjyAqo+VhQVXQDei9q6eB7pP2tToJwMibk0AoN2UHIexh2o6
OMz80wwOQK4SgqWkhAgmJ3rTn02YEX9i0tsyVn2CQmsPnYrW6N6AbG/OW33fMhoVNmEk6FAUUMZd
LWdXhXbCdt/THqq428i0gZXTFuXPJq5Q1UvxzNDDTBr73VkOnWZI6lwZwyO+8f4fFb1rXqKwYTBZ
ByfT7k853rEZwiBJ3gcgD6T4zTCSy+CGmyzOeqPAuaRtmwjavmPHV64Nd2EU0snvUVEOM53ajNWI
MLWUr0zJ0G5Nw3gajLh6qqD2YhQKSOXGPv0VqScOG//rTXR9zxkSORyrRBoN1RVO4eip4Alsd+/X
NLz36MLWwirL7Sz5iKBdkq625JB+5KlGz92DWWmjGPG3Bvl5Mz+o4Z/WrQl7J/4CIMc1pyCzctCi
fucVw88KyeuJLsZorN5Tm6DRjnJBT3U/xPiSe3GBrwxv+ICJ011Qj8D7Ma8qPKP6JXvTuq/l1Yf0
cLx8zRA8Aeo1a0FoNf8JK9adeWE7KGr1TPfrMXYYTKa5y5mGd32m6dy4O5oaZQpzxYdvYj12Ou9v
6l39AtrsYchWkC9b5sur7zeuCBVU8EHT9leNKFWPwu/qZ/qlRlk9kJhx/385kw/4S38rdUfYZh+/
HjfQYfnsfr3O0Z0wD3vtC4YqbkuF3FA0JC9iU0EfRgUe1v8kTYeasa1MawCxzZwVoVpRqHy46PeZ
XQM825k1OymagjvaLyul1huUVQ76x6A5qDVDVVBAlNLvqQ4PLx0Yl+Wx0lMhY4FQAHJbkjFRvX8w
M/eRNYUe8FYi+SfvMjnElv/OokLZx8t2mGWUuE4qE4AmFvGAii6D90F7CiqmXpp6MDmVkcIbOV0l
aY5X166RZLajTYqCFt3lGN05jPDYZbNe9rXOeV6gaHGoIf2Gn2dY7L96XCN7/wmnhJ6zpLDtk59b
AVGQjQVNNnfTUEvdkfrp2x+A602BoVso1EV2N2y57vffs0m+oac1DJRaOSId1kwK1vRgIquFMmPB
m4EQz+Da08ULGL0JZoeGzp8CLSeOt0Rk+dp60VIoqKQjVya9YH1DnhVKv1Pzm+qNJ6sUVZ15uQ0K
bkrjLcgTueSelAeL0S4zOhExiTJtMv72CGI8n5flq9X5xZ7f526PbTwWW3GazSlrFVgdZ3rG05ss
4iW2QCgt0fuqsWeqiYpUK6eN/7/IZ6lo8yB95tPzTouyK/Oi4FVtpBAfO28EI9BX2lZUDP5o7GNP
MEn/PXBi7BqymX2UyD4cb+SSoKTvCoxBe+iJSiiQKKoF2lOWs21kZ8I6TYVNT7Iwbw5+biXYhUfM
i/cSqD8TPLmlc6PCna3XapZYuXUDrRDvxEX8aMf5zl0PRcYjzfqVTmNE4Wds81jh5L3w7FKZWs3M
eMey5cqY88rUSUTHsjkF7yWsCeBwXw9IhPegJ2RW8rast1YfY8F8TMwPGln57XJwe5kJ6R+9QIKI
Zi2Ig9ZoNYFVhyOfwbmqCKgwRsKyEyaY6JPQy+qeYBX3etKEy1hILZEzFlp3KABsSm5ojh4eksrA
beWw4rMKTiWFeNbAa7W/y0V1d0wNMKKxzIhEQeYmIFtXRHPGnULsT4Z+u3u1/KqNNAqcHphgS2XT
gFzpk3ZdsGJAgA/LJrwg2vEPS0shw38N9hPHSNfmaORqDzfJfl/6ZI5QxQKo9zHRrsVXLK/OJX9T
+v0WbgD0Q55b68/SCEtF2+Tqy243Er0rqGYQHzhpIlZxpxDsxRzvd6BUCOqWb2lG3umVHsWl5Ynh
RQAU6nc0lj9Xdk48Ct4LAV28Rl3JD4kDMTNZgRVpxzxm9PJ/stnts2rxnB6svi2WGYr9IG4Sdyy1
p1P1E9mah1PLAVJhYprUgCb+7j2VbTsXdzqNgS+1EifYnjWoa6cUgM0PjHUFuFsgntrEl7NC4hRI
ZCAu/cJtiHuh9500mjkUa57D4DRRWAkWa2pqiRfyObsQ+M/mx4QFOik7qdHGhEBC2yaYMi+wX/Mm
XqPGfcUopC+cjEUeGsDUiFi2LME/buSjzWutihV/PY2rrjv9VZro+iKTF63CjOOirJn6apmQ/o0h
tjTurbr6EdKIVaLXJUzVwSnYwou2jctKgGdiS+tWjje29fDYK1AVgUHoTEz2TG57AJWQHFgXPZoX
9QfdM9xmzI+/y7QpCif8UDS7uE6IlSRbo4omOmOVLN1/ALRzPIHpHmnK4CPEdTUQpqmQHVCjDCHZ
7S1JeRve3ojXxmVJnwOm94YxyPm0zpYSQO/zPct6BwPxGHW8FwHhwADFBDuFj/PSBhOJHfLpfuRd
dc/8UJuRMXHNRy+dt6NR4Bup75BMYjZBx78kMMTr95NIrc3BMmMv8iqYmJlAwkI3UU0TcdMigmsz
IMMf2FfomlMRkbsdHLdjftOaB13dJpoFeMzr5YpN1uXC5hpvdcfGBD0zd9o03Z4fpurw1zvF5v4Q
3umMG5wKWuSjUjcydkBfRN4GmH9xDGENdwurIh9XSEVId7pH6VE8Zvi3IylA/zxBH7kwOsKY4oH9
fIjPXOPZc1lLgsUqwnsEsPe0A5fqwaksWziTwWWeh40aJ+XRoKvQwn4GuNehP+rrD1HYESRCswE8
bFcLCNtNLvwC/so9+sCM8GxKfSsOih0naEDODaGfIINi80NQzlG3bXv2gwat17eyjg0Vonwf9aEn
zP+JZNXOu2w+HjrvylMUkKvldjsSF8eFqxUkzvvEv5s/u2GEt0fxU8oJqOnbsdc+wVqwUVCvM7YT
d+H0K4jwzI41H98Ps+X1B0c8R8MWx65npOQTh4EMv5t5ocMKVm3KrpIkljDKgTM8eeNWXAdQM2Lu
zuXkcehfeJ1y4+OdJTBBDCwFcQlGYpmiLt+LvQ2Jy9N7EN2vvJd8DQ11aAZtt33c06kUOBRUKQAZ
JTeszGcdHaliCTMDfyRXXdywJd6VQHF6AyKkc73cZTgnYABp4oAXAdhkke5yIkLDSs9LcK35XdvH
1PT5QQ3nWPuHiIGfilFIGNLtYuQDCDHcWNC+GL8yYfQCiF5aHrkzlayU4iNQfHoJEiuKjPcFxKO1
yuY40eRbMfkXC60I0+Qp5PUc4dBO9XOgxzaqJ8jKAJ/VyTZ6cwugqJ2l9t36GiB0flBAdEQjIVLF
Tnwtd/ZaF3EkbsLryv2OopRO7YVsIm4PJ0NpGyzkiM6nGNHAIyk0VfhZ46xw1Q1c50AgTPQVvkD1
tNCsxuP4gNvAmO6d2ZLQu9BjWF+0hj1/+FIqT5DgTcMq+NDIN3zyLihHzsW+pTJ1HBJw/AfLqhGa
+JlXuIvj2xpIM7LNH4SsOBEPpZBlkxS+7ENffz54WkxrGDqcnDVsHECZ0zucJbD26uu1UMK/xE0r
mzN0zzJW8ay6V6bKTSlD9D0PqmTEVil3Oa8VnHknpLlN4+8FUzxNtKfXpZE+ZXgNcviwNBNg5EEU
5apgAP0SAt+Ykq/JMLuRro9yicRz/0WnL+U2ZANTck14kcs6gaiPuyPRDkT6lsqWDOmK1m3opArK
6ONtq0Fbx6pynYVJ9DfuM6anuYPx23knqnHrr3poHsVm6ggS/iT0s/zwUipz3ESOE4aG8Dm2Hp4q
yGMdzPpKQtT4mSbwLwRHyNudA5aJQ3TTzm+KtxvYxExl5wWGEFuueA0ElhanzSmBvConWQnAwXpX
oFWwq2f0oculqbZBlrierblOfSHGviUFy7B7n8MHFo7EJJtba7KWgUfv0sDXjhsEwjZ8hm4dtgIy
GWqTQ+1DOgUsk18Lr4up4GwSE00oNSRJdQyE13X3lhKOM8B9dDz2+0xirCU7yxzFDpEgFtL9QZWf
EGilMmtNshsZa4GgGZSZnlNDEJsVwgID1C+yPGUm3xzDop2GWmOROEFX2ukg/5Ljcm0XmaQN6XB6
hdngV12c8d47OREihABVRKAb7hfyYQ5ZkKq85EuV6b4uriYSt/MeDNV9vfIUvK7garVUJSeuCcXC
F8r6i5tWFUvHRnebIBMXUCLlFqDtzRM6IGft9dcEB7g2q7G6ybD8YkSiB8NsGFMAmCSbj/G4ljPa
yORL9DJ0yE10rLvMAf/OaYM57wbt+q8Nf8ZNWQx0rlhU/qtu177jCJI1rCHZTlLQGgykZpuJzgzJ
r5kQKW1JRByPkpcclpCp08kyk4GKiqLj9pEBjFIg7RhJ3fJDTdJuTzNm1UKSzm03B8XVrYz4FkeB
GwXhPHNhTCaOjZg4nyotnrJJEuJellcmRCdxncHNHc2WSrw1guXw1FtLK3MYHaFhUQuJCgrmd1ci
+1LOjM6TkhdPn1fE6qUpVcau4EE8XH1YKsz2F8M0zq2AaNatfAOXSA+Hjg95O+s8dUIBirkuSUd/
aiXluIhNHCw/MI9QRHRIncvUIcwZwUCc8ejA2F/P86OG7V2GCtmq1uPCLk6h6GuqEavEQtbgnHMU
PiNvjbWC1MPotjgI/EMpxZq94au1O0Waw7x700Mzfj/Q91iZ4jQ7jr3AmNOYH6x1onrUW/JBBnmS
2X2JDZnc5n3wHqUYGfZthaFJaqQnyfWv6ebATe7AsowljTYRel2dmb5c9hwgfOR8DMx79H9/ezPt
Drcxxsgkc8FYxHXNJBBmGMrGdBYzDj/961N0FEXCCbDnj6ta+Td9yX+bdbf8m9bcWHHW33tl30Jg
yp7H3B/CUDp2OPxkP63C2vK3fW1C6Ztf7tvjyLBupMgrxfI3oiP8AkRugSnstQBecyMO/gTszUkQ
LpD49PSSfsL4WOf2WrFjCiJlDx9+54erRfuQyccbXe/ZRqR8JeNDAP/gaiXOE/ADUa/LyJ1GcPev
yX0clivB2BUPTH/tqfGztxqCmHa3lLa0wnsgLEHtu8Ojpiu79gnt9AGo/mjHkaHBT1eWOgpW1fc/
DMlMZsdFbJvLa4O96orii5MUEkiJvOE2MtqWAMOLRDbfaBKNXPSqnJZLSnvwot38JMMjGS2YHIFh
yw+a4MPOkFHOzz/YhJgbOjBnvcBvTlIycLJrNfNobCjFfmC3oqzgQYlcBqdcEGM/C8RmO79Qhz00
kCZpciSYmyl/TJWt1Z/VlQtA/5mFcuvaRwmawHgBDR5mdvadVgoippggXes6owIuI6ePGG4wUurI
peH4Qp5XeVZ9tReVMTd3WtXidS0DkcXrvQnPcsouzdisn/A3mviIOfIFLVsp6F8t5EMAC1cceqYY
WSgVUGOM3FpsjRIgQjmn4kovFoAe9TVbxv9BxDkxz+xryNqvm1BYr3wYlJoL/kXpv6lfIO5e2o0+
ygHSiAOgk7HskOEu6tDmf7llIBnGv7ai7Hgt8dhwVFffMr9k/pGUxrJEFqRi1E6C0H/PtrHeeQlr
IToQbeE6Xd5YOGEaLtfZPwVJRuURwa6/p3lVkmQ1vWl4lZGkxblgoNR19k/53R9E4YSXX7AldVDJ
qyfaw4NEQ70j3zIVDFCsIzhxna3bPW36bFa/i+kLn1SmFXCf4l3ZDHzTGked6/UnYUlUjYgXFBzH
EuifrxsEkowg7iJ4MBOEkI9uN3xNxt+4zMVgynd2KDekhZxKusCpgoAlgf0aH6I8+byk8jSiy/rC
b3ObKwRQH3zQ9WKEBc1N7onOKzYqQk5/8ThzAUScwvopPz9zNbhY7P5bGLcXuvBun0duvTBvjYkv
8tjYgdkchIaJp4c8witYuovDcfBUQO8Cuv0mueZI4HlMTeH6gI/TgEqxc59ZuSXIYegGT0hpfEtn
G4mu+fYe6rPF7EhCzqrAc5uel+1k+0+iOuP+zBxwp9qxgPqKZmDa7PoqgbVAvpVKk/+P49JO5Vqa
wFDpv6DP2imwJl2mLoBr4etsNEMrOL1XoEt+hewfUH7lGlfEnbOIQi7eXwRIMR1MntMbUGh6tlqR
E2HW5DPYrDjE4ycZyJBzkuJVkI+1gfjaeh3BQDAwt/qeSfiWQZDzwxO5xCqv98j0a1HFBZSbU+NJ
Mt6u1K5B2duEeA9ebdVbjitf6HaHoORosLV18X4k0r9f7MYLYPmok+7mDeXhNcj9Kk/8WDfhN/5n
tXHgECKL9ZObPFtTh4nFM5Sj8ILDwv9lkcxVm96xyktFdFxGRmW8aP9TCkLBxlgY0g9RWYlXjKwS
ZwuQbZ9KTdrKpOPq63E0HTQ0+Jei/VB8dsK/EPFL1UpBOMXY0wTTpm9f9MQSPi9a25tDt5Vp4raw
YaIuebIlhD+rLjWJIZoRDtuTOsSPUwMJ0NN1tDr9SI/BlIXfsKB2oPESFI9b51EyV2KgrLdbwPAM
Fny/izcrezAJm9N17l0y6NDAiG430eWDASPfQV+fLYBpq8iLXWTnFPInpElh0sUi1lMIFjaFo+eZ
CsywwIgcbyG2qbMEb0yEeYiP/zMuyDkQ3pxEjE4uP1Qj0ot0YPuD3FrDSVmdIljPEIV5+VULo8A2
Z2JDbGCne9bVilibuwilrNf1g7KoXByeUrLrR+LbuM7R76HsSu8R0XpnVNxzcHoHxzK/W62WMZbk
h4jjmR6E7fDlY9JLg/JDgNjYv3zKIFXlVZdII6/BP0ZMIOt0QtpH6kTI772/CpWc1L5AO/GNoFpw
rkhbNLOBxnmOM9xQ7hq/ZJjBHfVk2Dii/hSGUGXs9RwBZZ+5NPp4VutN1QFH1uiBjZwBCu8XkTsi
+tGQ4QztuWR5j2k/wwU2W08Hu4nfIcSOpT9tbG+tU5Rh68TH7hNSy5mJRbF4ta0b18UoEs32neqt
GZQY8W6tlHMONae177MIBfWPVxJrsa87SR26XnRg30vuyqGxTgG3OULS+UkfNRLji6vj+OKrcEbR
MIit7HNEvoaQvDI7eSgTv5agGtEhl42jDRluOzlMky1Vqj9mXUZIsMES1ajVRulBe5ti2vLLruXd
ruUl9qod6YxgQwZAwqYKkcQj7rTRQeSPUUsUr1PgXvD+4F1fe/E+LQBUPjlljTDLwWvMlZOCKY6w
qlnpnWPa+tIQzW7KtemTkW/FO6Odc+Y/wGlZ/diS2ZwjISoFuHCGItdYmaEVSi4qO226jXuWiqUb
o6TrNvAmXxPEwVL4ifvwuNoi+MJ+DFWvzyo078bKwr/2PJ6Q61nLUMYgicDcxIJNV5kr3AYcy/FN
Im1xWniJeoCsrRkp9VE0GL9EY/g/11hFpgZlsXjUx7ki535ENXUd0IZI2QSO6igfYm3mgWS2SlDT
CYo6GFavYSB71dmE1i7LEoVnaa7A1As7zTdvx75B/g1eCrMLCBW6fveHMoVJjZ5GGW/ubhMYTyEO
8woOWQlsTu53GSIRHwtzC8XAX12C6UdBPk0pguBDdUkKOilQeZ5Aq/KpdnzAHjMCw+cJHExaTG81
2vKWmll7ZX6lHtE/ZxgihAlPvqC6jCh64Ppv5Bfnzqb2G4fbjtdYWDF9NppbHH+bpUAsVZ7rZrsa
7CrHz0e2KIcnP8dWyFocOCyKC1VZvHZOaQVKBNI5JpinVSMtVjWdoOcgtu50R0WMS7lIADGYfS/0
MWcxIL9jd4kNtSX/pjBvi4/e5wEV0FfvF/tNKcqNJqnGEn+Th7kF69UaStn0KYps+dEt7eFjDflu
PBVN6hncP9Zx5bLI/Jwah6N3v7dN1r0dGd0VqrAES6z3Jdc8xwP0u+W0HjxdUlY1/k/Qqw0rJW4P
7ZxPJxc2YtMhJOEWRI5TiQhDOyX9i624a+bxaFvcFk6D7+MKKaAu3laTOLZuRV1+gVw0HeKqo5Jq
3uPq6VdP+0PQ5A9RfbsB4cdDeNVZrmXae4GGr0cvu2Uqj22okf3q0d+PhPaww/Xyluv8ZY6Gp9fl
l8HnywF8v1ewhKu+qZlG7fM1UU5AIU8bWf2Q9A5gcdxSv3PXzQm1ySd95pAizpneJ3QZaoKhOTv8
NsN2aUIdmFzUBh/3lKrpWjFsSskxoFf634XSaFXCCNun4teqVljOY7p0D6Xdb3fef+/SuFQV7Bom
63VhN70DHwLRMI00Ax73QfqbtnBgZiddAv2IJLGWYS7/pQs3kx1ePvpIgIPGO+AGOB/A9D67jVrx
XsS8GWBECYen29YTX+doULjTku3ZysXKKmAdbd6y/C2Cgj+M4Cvl1RzEPRxwIOYzu2cqZIyr+w+T
49yzXXiXg1m6uwANKw8RmMjNjk5BvppVr71QL+cLSdLh11bhslTNbFpMn9lIJpY3dJK4dp+efCgm
kv/Bs1gGaSxH0KDpgd4jNzU1XzD/OCJHFBzdUCPq5jUNN0uuXcLCOyHrKmTc/CFIZRWxGv4kzUnQ
vGwslr38d5ORSHZnA+hHpyZjH9/dDY+tu8fyrjgxrmv6DSBNalMkN4XF/SpcpUTxyyeW+Kkb9r6z
B5kJGtkuLxV5Iks9PwC9gOQcC0lQ8S26DtPyy6RN4102QTdVaA+LtmjF2+dEojQAPe1s42a8HssG
jauxB+MeY9/P4QveZs7Piezd+G7zhXk02b3LCEu+SLENS0bWQelp+NXM4nejkCLnyNn1NUxkBnkT
JjEImqdXmSce4oMjKMY47b9m/JAPXr15/4rNKrkej8AgqIvA9hofzEVTp5Sa517PChjZ/IPidrd0
sBP8CcKMhIoErEbpnK+ej34gmG9ja24qFGTHXA7L081pvRfUvPogYPysOdysdhdwxDekfBRifsTL
QuxrtvFrvLXUu1CASvnUB9mGrCReuxV9qrG2CV0Fr9FVCPLZk0WlSqEoDo7uxhfX8miHprd0GgKo
KQAU+aw1wuRirB+gc7CsYzklH4f9MMjDXmyGegqRVCikWFbhio/F/kUhCCfDl45iOdJfW191s+CJ
I/xdf5t9cg+r7W4FAcrAv88iPpS43mVCymxieSpiKkiD6QyqSmLc15gFhXda+KwVs238MycRRSJ9
WjH7j0aYzjh3UFvEw4xcXs3CvVbqdl3P4YTzGjaZGhjBXH5TfyMV3Zewt7PFaXFFuoMlCkIcMmOX
chcYjq4jNoXD1xqRDByYwERY8KURQaHaRcbR0Pefk5Ib9+UizP9yFcLngHBsqO3UkmbPY1Z2quqc
qjuHRzMrGzjAZW5oC6UzhM6+dJ+r1XDyV1ceP0ym4RhUGF/cjatO5FcgdKwJlgX+9wPx1zrjGquq
KVuulVg/MeL7Q98BTEy4KOryo6ZYt48bJ85BmOyZc3Wv5gYl0Tv+vKoWFKEf3QOlU5hgDo7e4pFr
GHrVkok+Tqti/6shF2orl/qfj+Uf7PkH/uA2DRgJLueH1igICFAvRdtrCkSD+u76hRskTStOo5MR
RakcI1+cVWz6XEREj3cVnBK+cTISxQ4wfje9NMwuYDFypb3yi8Hgxkw13xG9VMKp1TnuQTiHxI7V
Ax1tTmjNOWvffmp0bpEZwLWnRmwjJ6I92KhvBVZfjH4ZV0mnslJrq83zoR98VlNWIlFBXw9DQS/A
9U7MMvQs4qzBJIsfErXh785ycarzCEP8sgH4k0/2oeyRRc+bIG6MxdDY5e7FmCImpafmdHLzN43x
O26vMpwi3Sgx1fdvmXiBs+yVvQF8sVaqs/9OujGigwz6bB6Pckvw1Ys/w2W8soj+uwl9OyPYMz+6
NkiE3pa48enlHnkWalQMmp8y5+2vEYR2FT8kmvywWLr4Pbtng0QPVWOc0ELuXZTXQK+utZDQT+MN
iKQvD2R1G/uMYopagAeBtgVS0Am2ItQMjk8eDCdTgJDzhrVrXWJFu+l80P/cuwFL6x8i1z3luPRh
IXmXc82vB/74iU/wv1P4c3mCOcYCSxleeUFUDG3YtpGs2ufYTmsqGriIaKzeP2wJJgkVDp+P6oNB
EtDMc9Wip8D71fqKGVnidvjUDlkCW2KhRSgSg72ChJwPs+EyXNA43xUdgdPvxp5AzdIyOAPYnE0p
cOjpQ/ZCSpdRvGVkQTj2Z8cnM+SkwDqsI3+lr8jbV3ujiL6EIeGXjUADv9UW7shwqgedrCa2DKXo
N5pC6qIKRaYq6FqctgCqGirwnIS9HTz9DDu8slaMSr7VdNhNn6hbwm5WNstO+TbLAcOZTlju3jBX
4cCp9zdM5lGdA8/ZblmiHq2aTXjTcnNSBKSyZWMiEJ/by1Us97BX8n6N739MX8x61TsCkDlUeLT4
f6rj1b1BZN2dGhaYzOP4rPRNzCsFZ9fnqHlFm57t5nFSK9xge1Nvfs+Dr8+RUNGSITweU9sd0LVD
C8dDHCeBkpOLWDnum6wAZkWZ794rtGZDSVMA3gG2z/msDV5AjM6t1Zg4UQa146fM6CM0JnsNGblN
sJyuOuqG+4hwJaP2lRe13f+eg6J4AFJtXKhLVR17mODT/bpok/vhj0Ri2epklVwY7StIYl69ybyI
wkyNLac+VRoTlvKmol28OSY93sUxyTmou8UyE4Feu+Ibg3gZqiW9zlitd9EZgb2MVov79Y3CVXVp
Qk38kHYRaCmiNiKEujmyaygS/7EiCC0aRl64FH+AWj0a+IlcOwOVB7fVU0Hgw0XURKNs/1siMPCS
4Oe3jhZTTrwtglHg59NJ+Z66u1SZhp1lMrO2SUmj/LSYChQojQG3PcfKTGFzX8Vx652R2d73Fmg/
rvHwgBWtmkfp35UzOFIaz1QcfzHZHCVbm7KNuQdhEinqsbzWex4QmIUcvvCjVzsLvgnn0WaflAy3
7LaP1IyEozbEd8Zjmx1uTxBlUarCQV2BGUh6S0sKNQbevflm5/jxqGCp/7+xTQLZ5pNc5e4Xa78d
Jps+rFZTj+f7/orfKHvX68LPATfMfqVsB2nA2uo1E2ITtplTIn/hVhGuqzBFGtDyk8KStPo4HbNs
7VLLd5x0+N9QSyENLh2siGxtQjVT3uELWmQOKRKkgz52qj9GdUl1KhqNXrg7Meo+ZCtKuEvZoIBe
zNRlYt6wP2PERFHBWXhPU/Mu9guXB1zTUnXuzmL9eHCkeLfckfaVMRq+ZTD7uyy7QtTL7pUAtoRR
Sveq3Ib9uN5TiEfkhxRaCiO3c5tmshq+jDNPwgvGNNvgoFJ9My+65KiikhtUmp0KT/Ra9PufS+lM
8TcgSevIKp6dNEI9c6KZvMVbK6QcI2YpV7rnjaBZ+AWtyqE9f+YugFOQnnVwflvbK319Uo2h6W+T
jGGe6evC1uM4ydM41s7jnXuKt8hoyj0nKG7SkBcBreVCP50p1TP6U+E8xiyGuBQ8bhNrCq70Exg1
UTOraARaJaab/9RZ0ehuXam/vuB9hdzrw0u4W1ryGLe1veYIug5yJdVa6SaO+pMMN4m1D2y0Nx7n
oS0xIbRXEnZKOU8NrciptWdIb6mqO8dAMZjpqikghBGCQNvQQzRko78Zhj47w7Ljqo41Gy//OIEz
AzBHl78du9MPd8buSVMO6k6HPoV5Yrxqrz9eUGJWqA22++LH94C8Tq16F0GILxyI7yoqUOmyUCXq
7L9K9HmhzTLFelupZ8y3rV3yukPt23GNj2jkYIMeA5uUqX3OaHW3iVe279g7Sl6abPdUAKGd8v0y
vmNx6DngbR5qoUGKo//HCROOUDbEKf/cuo3gyOg7H7+KamjChZdIoCUUW8RrJl+3CqYtL9h0kEY6
/93UGD3M0ny7prunRcdC9L4IHx+5KuWx4DUzcMHlX7+Cw2fuzXXu1f0gRbAEG9hUiGVFpPz2yPJT
899ir86isp9yqTM4jK/l1F96TfV+LS8lc/0ooYYE0c2VmIiFg9Aavro70tfFRWz+sMrWG5E2G5ci
sqmxOx6epekxlTqal8uo+HfVydIW1SqGsaEffiBUySremR8X3a3dAIH9BulYMDuNQStq2F1NWa3/
yg9m5C7P/avjbs52cFimvTM3jEpC/o5asu7YxEDqyQPV7oNkHzE5CvxA5bfJ1S82mT7JV0BOmXuL
qlJ6qFs2uXpz/qDdK9k0Ei5VNQws8pCtyFhCQRfrIeKtgS4JSOu7+tMsHBh2ccna3XIYsZSrtmEE
kyyT+S3WsxY4sENI/lUvsCLIsCnHMkU1nIi30GnZmu+yh4+TZR/vFu2VGz/XPD7Eeuse8S/sNucj
rLeLWH6A8jVmOcVV0Tc/bn1CYzBCc3d9WVUaeXmiCsGzasrpCAi0RuuEfbOZK7rdDYwuA/Dfs546
lLJybEa5UIRLVVwxFQNLacvH//+efJUhVS93mDeCXw901sKjsBjiPAppVZPHYFGqae2IOsTP0aGu
8ba8WrmfqQVkuoJtvewDKzIyxNlEkdGzLTf/jolxTgozaCaTKDJqLMn1jXxTioljdu5iEVkkXqCo
M3Bj0s+uZjM3ak3JpAtB7+wqjtElirTO1ZDHddOk99qiTpJNm7zIHs+2RmW5YGisZ40dvmFsjf5T
L2cg9ePdN02dvsY6yEVemcAas4YpIFCUnreipaTawLCa3xsVQUxwR7GXooO9xiIw7btwLRVhdloU
u0WANXucTv5lFnMvT7oh8EBiiJrVDFNQTejLqSwAPEHsqG2x3XWGSMxpy7jMwRJn0InqzHiTWBUb
45vMMKLw4M81CGVuydZFrwXvv9AVY1uQ1zpFsikmu/DGlnj86UPu/RwnXDmElEi5T0VUuhRK+8DD
v9GYNPhbSjZLb0HiAL9rNOdNWyjPadNoJyvfxlV7x+wUVgGu8zChaTsc38AX2cQB0E4whQzhtHFm
wyMhFW+1art+Xj+2FhpfzewInCFjcayFUiRNOTxoD+uMYtrHe3QUcps1aRfNsEj0hx9z0oFpwglG
idrrkmrJXzu80qpeV3kXtKIzMlbGzUrSBL9LIC4HrWqnmuDSjv2W3RDcMTQUOf4sXwYVMbjO8rgW
MXULQqedE/CD/nh7IsxDweJrqpy6LF6nfYIAd/M/9x1rl8gxSIxBfU9H47W98DleClqSkqhWL+2+
KAv0jD0QJe3SVSIPW78lIC0mQnSBSuyDJuNXAlJx/pXTojl5nWgVplw+EOVC6xw5tkdhzAt752gY
7/n2XAfEQ0gpJ4+Ys/fHBkM7ClnCmAv6d1py17WbgL7k6aIMfb56I2pP1LPdP0xDrmo5tb58n8sF
Rs+uHPEzzQq6pVQOEVznuPkbUNhvA4YvagsYPRslmc9Vc5Yey+PwsnO6WVyikT5n7rosjbGuNyyP
l0qnwKryeqSp8zMeyu4vUG6QhbTH25poBMXNQNwoGgpkBbwmvrp1j3atnbDGelB/guS8pOsdAfSh
wBXq6RGnPMTaTT0OI5iBdCHQWOJLut5EkQMK3ZL7FH0w0oth+LC/7cEJQuuowxd/HUcCGFvWPiqk
pW3H5IxOheXfkOJWp4zj6E228INzdRjeHPbX+EcT93H5kP3DDklJm5LUiW5SZZv9mMKO65AmWO0h
V2zLwRGiQ7d2OZe5/Y/7EJdcodqJyBxmvqK3MaS+tBF09vs6hhZ4sD946ydQi3AnRxxWw5bBUrls
3zHc+Yg1mpqNxZRu6Y3/9BXZDdd+hg3drBMwLtplKMCmygVBYVqLPqdDuv8kvlFGJ3DyTU8N6Y4x
SJ/tG7a6ABdteeffop9CLNpmZVJlazam5kI7jq4rOEXJpi8LTbje/X6F+jBrn7JHN/KWuUwSZt5g
mepP+EcJsOJjykl+OtEkPoi+FOy0bXIQ+8gHPiSdplHN1ulVHCKX1U+LUu7dr67w3WAzSHpVzBjH
b8j+S+907Z/IJJuWbsF1vEtvQcXBmR0oZuLyNFH0btvUkRu735qztALZP1TAhlg9dgHGJHTDTbig
O/NUJ8x2xYtBWO66U6tEU0i1R1kxJwewjPls9AHfEDh0yWSsiFCJLz9hSJobxQ8EoLdro0un69NN
pV6sHBypaSLDDks8MwvqMZErOBVV3e/KEqvNwEdyqbXeyc3tTqXVp6x3IfaZjUSEDANTe3ATkhC3
nTx8mlu3SBqDSYwJ58dtar4HqPe+zU6rxOu+JO/1qBvgcF4eakyESa7hlcl5R0FLbsqVOnrImSp8
bZ3vahc53UcnC/7k9TkWVPzTyl91hoHv6q8NDLpjfpQS74H1GXJOidAF/fW0tw22+YtE9Rg+hKce
MjDhk08KgvRiADgLQiOWvzLQw0HdpAsZhWxr1fku3grth0EYAXEtluAdA4x24SwS+HInEdvBIW8J
Pdf8+Shwx6R+hSdM+KCEVL/oSIqNmGVGfthWTUrwUPfl6fMmXHXnnFOWHJneuWEQdMQt1pwyTdj4
FMg5axXAAksq0W5fnVLS3wDkEBMV4eCBqZnVIku2OpeWcjAXGQHNqSjXvrfmX91zdKJGWa404DXg
m4R2mPSVtavzGXykwDp7WDAE3JkBqC99X0DldUw44aZ8064V0EwZVS8YYiTweUeTT2osGqsWWLE8
yPoU3EUXjlew1KWfv/IPU/Vd4WH7o35QlH+ylpDfQishefxqGkhNAoP1ORFkwL4YfYrtA2wK+0Y+
iWsgK8asRb+EisNo0icOTgmkAVpeWbnB0yrV2MmMLU1CqVlrzBkW75/CJSoWpHio7sUJ/HjAChzJ
uTHbrGv4xPnDo7c4xD73Jr4zUUv1RQ9NjqabihM+BpCoFZFDgFP7196SO72M8DRVbkcaNa3u5v8j
UC3YdHKiaEoOJzoVzkOGpbhEOf3OTIzYiCuifGQ+x0YNcbuMpv6SD1ifmB5EZbthreUXxFIybUxZ
3yTf1oNzqOVUSyiNGaiA6aayPqE0zDXlNAAuYzj+7TUJdqmP7vlhhfHgtiLL+SHqymqByusq67U1
vx66CpktSdMUYAStnUTYep8y+01557sldww+cw81NuXQ+XZddGvkYfbC1u+d7esZ+zPHF2mIX0kO
YPRVK7cnFwJ0hlXMtQV45VouyDy4jh5eXkU0tPUunZYlBrisGNbru3rK8HieqLyqtxeNy58f0LDw
5BTXZLWCJQqKiF4Owj1C4RmaeaTMDUuQ0U46GGdlrXlrA7/VeyD80ScFmNwHrz2UIHKsP0dlHCKB
zh3xOHajIdaPy0QN3/q43RInRXapntzQS+3yX1NnTfrjCeA0aG2uIkTvHR0SYKvYiGhTR9jqbdLz
bqHGgoA3CXcp2lT26wZr+MdH2XAL4WjPnJCteXClDDoPn1IotlQJlLobVBMOsl4xcHycOrD06Piv
y+QfqYqLGM8Eyuu9Iyk00uucImt1NIsd5jet2UHcT0xmgqhk5cQj2q/BY9xzbCwGQkv58oJDCTLg
fRxSG4LjGKZ81ACWKmVKoQj2rEcIqDaFnNRGHIaz1WqG1UK6hsOec8fdaITyHLwMq0PZKjrjKSR+
JQ2Ls49l//YM8U0ha9Cai3zRU7NmynsQ/VrEeIq3lRzQ/45W1Sdo5HVxa/RT64KySWy8CwxXEGt5
d9xt7TeLTonXexh5fnYHLHyH44sm97qQ1SXU8nj85CKw1AbnWQL/6xYxlAOkNUtiwsgL0tu2JMGf
PmwnSTKtx3hkwgK/Z5ZKVl2OOIAdD5Gmz/QMMnjIQyyvwumGqYwFs04n00lE0pNIzxXFJPdztfqB
KYaC1xz916T9DwEm2YP5wisUKRZc7YW4aL/Puq/q0hy89G+JDjsxLndawhTQspj4J1KkWLQwfo3Y
+rV0wxEo7jpa261Zq9HuZ4ZXudxzqRCGi3fi1HLG6qjNjfp5AcBLAerZDslr5FbA4lnzjXkxhgQp
JcEBmC5rW/0ZL0XDmTYvVeoWCFAqmR7sPRMCgSgbDmpLXziyi6xLhDmIxVHPbHlv7B/jnilRJ/Tn
Yl0HHaLy+O+3/SZuf8lru2kfXL0OVU+xRx9zntJJNGLt0AcDi4fFGLjPpH2t6Sk5dguqB/nKzXlZ
/KNAPgZfoIAat0TYVDmD8uQU8+LrtH++Z6ChygIpsuCvydnvt0Q8aehB4SA1UbjdRc88j9mbc3TP
0NyO7awtgShCS3YH1Jp3qDn78To73ADAzq3+GXDgJb9pacJEvU9ts5MMta5IPDT71hXn6QBhfzLE
GXeNFMjEWc1hG4dBf+UQNYwE7Fgws4gJKGp3TSdk4gkUhM9kTzLZxYm0m1Qu+DaUwkgG8JOS6l0L
L/XOWLANf5IJprW+NYiSwK7p1uiSYjtdnKGikToUraQ5BFr8bARNwwlZfdc4N6huBkA+4uGetsXV
NiTid0Q2e+LXTDI7Q8wpvIp85iXonLNkn4un9PEiPzy8FDER3gt5gQHS0BI8kTf0cmZvoh5icgud
hqXpRMP7yNSBp2vNwiuiIUuFIimxYycEa5ZdjeH96Nkc7nH5rXOBkbR0zp8NPTAfNqWTgf01eSxM
PNIpbHE3AQD8tHNYC24xMfjN4xySLhcdfMcKW2cDdwzFJg48woI17e79cbfB+mfc7IviZfrBU6Fz
bgoni8ZRUf9CAaJRjDsbd1cVDNFrwYM8n5a7ty/NAIuFcyVWV2D92c8Txn+EWTkSmM9f/zjpXEqn
zIlUzE2bMDraR01D6K/+ok53FMEN6n4pAUWnLUiZPLBJPMX4fbW0QGCl06PtB1IkBHCwm7tEWm8F
CdakXLbcZpBOhZQwQ++B0wV6YhFttKSiJWzHN/EobDIyr8E70TrWOwKcVIjUHlahoYadMTiKTdIw
h888mS4QqY/2iFOkIsA3BqAlwMQHKLUf+lPQ6UBfpEOCoGlcjJlgZ4UY0x6YSgIpa0P/cth343EV
u/1GfTg9HVzO2pwYxHJa381pNNH4IvkGAMA7oWIHSGLE0466jBLWc+h534i36Tn5NiYL75+fReUE
miciEViBE5Slb2SW7v4K6i+nUibohte0ssjocwlYGjdVmt7UVXW9jLDgFZihvuKQEagPWpXxs2zW
7J3qgGdNJUnDKwsCHh/5CftP58qgpSQUq5dzXMToHSEr7W3Bh1wTCRTRVJz8l9L+nlx+Y6/r1bfU
i24t+Gvk0ZpH2vp88dwDlD0qave7dHU0sE2jJEVskJ3uzoBCNK+nFKQ4UIRt6cCPbIl/Fr/QZ7YJ
USQU7RsKVM/33EoeuG3CB5uKQb0fFm2UHw5AiAAjnme69DX9RmATjR/ONsfDLzowu2buridzLi0U
1vYGHgc4x3mfgkbN0vG96VJqAjwvAeihL2nRT8VEVkgsfAvFd0G3wRQg9RQzQ8Wq7OjgpWhKc/D1
Q1aoL32drLdKUTdm2fklPa3R+FWUiBV8L9jYpCG676YTVhBfOJjeCThaSBxyRVdVS9yrl4/OPBjn
krWauxXbe5mRcx2Dzor9XoxNbX3/CVqQIIiKdr8BDsCmbrD2LtJRrUqwYiy8XiTbotcqCQTer9gY
WBwycgN6dhvAanKAjFnK57Ep4UJfndj5o5KM157HVmc+azOdRAssEd8SAojuqf2/X7kKnlgV1UMG
ytROvlNYoIFhqaVFUushHYXjEzqJ9EsMxpdX16Wn2GWWFW+lXg6FDMv6M6398sssNSSsdu4XqJhb
vuNbUyxFw3Y+VGfvUcXIsqTRsEIBUdUIuB/6s7Pz7RqoN7uE8+yqzU7LICvY8YjFHoRhfy+AD4Ec
4SHHyfTUlmrrkVVQTbgHhTVsVDsGGfHyCa7ZWQnxyHb0nzNOvaZE9N+PdfyCGKgESwVnCY8lzWt3
B8f2BHu756vnIQyCo45s1mGVLP8nrIWQy0luH6G5dU1+2ly5NkpR4fRM8BU/VDsJG1p4Bez8q1qK
orSjkyzZBaMEjZNYrygTU/xJQxBN05uBUohm//bJfzUXW5vog8gepKj6OzAHIpGxDXpExI0BXM8D
/txM2QXxDCXLcutYBTFjrQDgyLX+YPwkMA16DA5tOCkeOKBPKI7KJ7Do2/oJKf6Z4WCwN0rDrD1V
ddNIlLw+Iw9s/aeSGik7zNwffnxdgCevzY1HyiMVKRejBLcEtakf11dixlL8jXDGuw2+xzI5UA/S
6aWn/0RV+Re7tmOc7abg3EV2E284wdhLm/rUD+DIXbJBeHIkNFBFRIp9t0/nXFo7QOIOemk6OVGK
aA62RDWWkgUhNh/P5uPGYkHvsD90G3xO7Ug1uLOrtnXs8pHS5i4C2mNdNBGDDGc4U/G7XTasDVNZ
GMPOeB/V9UcWL33huPa5pvZqrYg15wWi06qpEfKdBOQdtM/CJB9PGJt402HQiJNGpsseQXW4ovbi
JVq+Ov3MdM4FhE/fL1PX3oQegTZ3LtOVWAphTtJxU0YxtzBwOdfcRsrj4Bw00/v+Ps+JBQTcp7SX
5eiDS5MULOtkNQDM8UPKf7y1Nr1Uumum7BxZtRfMNoeBGS/TDeirpx57zr6Z7ciqTDOR/cs4pbpO
NzY/vGJetaWN/e7cLzU8XG2YvTc+AL5v0O5FmgH5sZ2jXOE0yJ0IWeve06LPLOWWbJnPDITmmx4g
V5DERgaH6AXFdRNXybXmNQZN8bB3Tq23r+fhyg3uqd+UDdMcZFq9027X8Rt9b/QT8rHa83pskJu6
xF53VbejvAiFIxV0QMQRaEBJcW/tqH/4D18JfZEOwKV3f5iReiM9ZYaJvfRxfBluWNVNIjrrO1Oz
j71FpTE7L09AC1N88Jcm02oUpy6kI8LM6NZk9EUvbOG2ib2BdPMCqeIzAYrEX+3R8axubTKonkBD
SgU2BvDfW1NCeXNa+aCSva8i0keDwb+zzR07Xx+Vu0LwRpBf1Rk3BFzf3FU1E8Jrt5sho+ljSNZq
5//CImRU1DJuLsoreHMK4DqSjnORTvwgpRGfGjMrdKEbEQW6XfkvbkND+Eai+SDhlVFDELNbZLIB
y6ChHyPFktDImxqK7MHPYudD6uMIapNF5Z0mMdlqNj/CJCvi7t+cHjoYeaTpJuzy5GzgZFwtzy+Y
Pv59oYMgK6G//qSIAzXDbXAANhR2A8TeLJgmlsgGSs/TU2eJ5i9U3mMuZ6hVRWgvSJkHReanXtC/
Od+lbGopN7hQdhz3diD/H8nhGnWRk/nLTa43p1mJRYLaESMx6W5J4txiubTyS1c6FLfYndNBrpNA
Q5R/maupCrRRrMUHqC4BNU4QBcd8jJA2vyMrbfRUgqE3jiKrAME1tQ1+k+AILp4i2ZdN9vd1tTFf
u+HZsLovp2dtnQ/l7C4PrNkElZDwIfvj3eD9I7PIyR+trTQqw3osrR2oTealwWL+BhnLihcyE+GM
Vho1OqNY5lAFnuTiCgdo0wc5qaQj08S2dLNKvKNpWlhtslkn+iJ0PzqHWoqQf2ngOGGDx/JxbN4y
5TOv36o8NOj7JOzfj16yeduSr42LiDBOODild47hqRtSx+HgCLDi/ReVABFNvDMm2vifw35SD+eF
szn6N9A7tkBcCufpeP8LYeSLgLJyyIE87AStzB8Q/OIARsjP5xcn/p2Ki1SeSeIAcEAidX/Zj5l8
j1CdsqNVWhrq3a8NIQbvWh4bNjtNsX/mgoA2Aux/f2M40rxIH8DAqKSHtaalH0c+uNmq3P8QXw+R
pb5VjorHEhzpN9C9b0EyqYFUQY8/ymnBWl/I1O37VUI96NgWbXDfusQMpm7wY2PglUG1m/pfuoUG
UC2Xcdvz+ha8ZaeAJnt9auXuUp6B6qjuNwiVOt3CNHg1ys9K0RYHK4YEyxzLRYYMmj0V0nzxJUe5
lX1/L/+fh7SQCT42nyU2t9hWuPVfbQAmJrvkekeKJ9vGXSMLhBYPVj5aXhNwM4elUcVfj/VAGsAB
iPo7GAoBRLc6M6uinMsglk+HaiSAWcRw5x7OgPJNU6+1JpFfalIB7HHaZOh8gP7AmqttLlrP7EEf
HF1DCUKMjULnQ6LX2V16syUBo+1mqBKyxq+ql4hP8YikT/gVmTm5TnhScIGyWitAbgC6o7Wtxfpt
pL51t2+HXv9c9pYuzrFzTkwNZ3Uo3T/ZqVVjfGOlqLyA9j3kNipmI+G6I/IRUvdX/zM9lT0y615/
btVvxSK2TtfAMJhdi1fRQbaTrnHgbytBxiS3M4uCpIl6E5GvDM5wj7QHuNXrDiCutgzTgzTfjgrh
BJDQKCTUSS6A400i0k/m3guYEITgRul6SdF8oBcpDXZ84dfu6zn2Qi2H5LQpf1h5GRq78eH+3uBg
5kkfumC8HNI/7+reqegzbLUY7FgojlC9FsF3dllyj5/VULsbI9/tJvuArWAeljx/iPWurHDP+vvd
xpqbxSJ9jZizBtXO3SSsVgfPJ5CgIEYyJl8Cwn1POZhsSEeafPwFW9nBTXRognmKu8Hbn2gtCxtQ
bVgUGl3rfnQuHB4H94bxKfV0aENbo2ZygVjLa0fDX7z7+rlosmMz9fJ5egJW6V8kLVdEuY5kr8/K
5idloZi0QSA1cBbTHZSqqrNtc25SMiAd4JKZPAyXBR0kSqe1LNOz46pmF/WA7dkydJxzcl3y9Qmg
UhXkwxLncdSU+w4sATxmnVx62BfY25t6TPQImYlMPs2gvaRUfUB2yCNswRuTuABUnTlGRYeOn0ed
6rNXXtRQGdLMzwhfDDbrx1p0uUj9DGoXdTV510vcIso1VYUY3PAKBV8CRQlm6zsVTaOzbaaSTk7w
CNCuekeGB7Jblsd+rn1V67sQMGIhIMTP3NnOTnSLtEnP+nOfzFDTrdcMkzLILewzcXF/58fgvRow
fzqDFR8XETKYB8zIPBJCOQUZ6J2PHhOTs+crUOt8+t+Qu3SmvEe6xBpVSoTtMyYIfmWehlQlUVPc
CAExfToB50ST6G1qg1cQyZH8twU+fXSaQa8bwDD2nFXSPF514riGwYYb45fVs5fEvXen0eeynDxC
BnKKwto30EOLGdfT7fRLOa6VryVuhN9gEKRFPvLxRlaO5nDGentVx4Ji0VtWqnhkJgWsgVtYJ7AD
Z8CEeTmkxpQe7iviV4/buaefYusMsHlQu8MRovq1l6I+IDCzOZadhsGq0sRvfT6gGLvNi0S8kRhV
ZoS/MYXeExmNGhMlDguhir52xhIjaUE18+0hw5gyxmu260de9rkZyVt7yz7EL1wzBftS3XN2mk1H
zTL6XcBYgdoUnk1/wwuXsNvGVlX0X+DYdTL8mNE8FW2Nkld9vLBrfD1nwxtk1lVe2GuUG2Y6zE2n
mR0JPOdo4gfB3X1plj27xUv5mFDxyz6GVJ6mabvH6hesaesKWiO1agQcBfgvWUEkq6F+yJ6tpsDW
wMX44tS83mszWmAh8s8p3xadYSELB9tSkZKPdJzUEod73f7PEcOIznu0bIsHvJ3P+Hro46v/LXFZ
rJu2IdAFtosSxflOnl/K/e5XIMnsSxeO98mlT00dqX2RTqURHkJEjVamUmxo+nt8p7k6WoQB+/iE
mzC42X4BS7T8VCXHMLZUab/xc/mLGm5zUuJJrbDa1HXinHhFsIH+wACsQv++KvK/qpfv26jCdibL
wNQaYxPdnILx91WQv3xd4Q8nEgB/NvyirPBWmonui3TtFqvubBMTMAN9+EXQ2/0RQiqQEBOPiK2L
6iHTcnooVDcQ9ZWanARzhHROJsy/H3aMqxDwR99K3pVQ4ciJ0nHDDQUsv9Qo3yDT1xW9O2BWItjz
097meip7a/Vi7Wj4e8gei8ATBKIM5xadQk6Wo5xSRnjk8kVxu0JnphcULF0YJODo0b2CZu59nUfp
Fb7m/14/eSV1AUnmOjB0xx8vm1LTFjCdkcvBz1qJdW69qQiLV/Ju6BITIpUcBFi/NN3v69XQAskp
nEshVdk3ITc6US4mGdsZTiR5OMQtogCuDavi/fNxwuzR3MEAQ37vSmayCLHq7Z1a3mw5kPpB4WzW
qsEa6CdeoXV+FvxeCnQtI5zSMNY7Yc7p1nAbI/axMwLVpPmLHLZPc0ZOemFB/XkWjK/gi8VWnIDo
7O6730T/hIa6HdZZrRLrq+5OafYSFD/0HEuhPmws+BBel9h/FAs1rMIol6Es2wdM4D3O4kV/op/z
zLK+tN9dkzTDMaE4l2AEaPpJuqyqeNKgdhvMLR9SkUGbc37ODZsR/Iw6K3cFFK9iM30HCgyacviE
kvmN7zFFV0IS1g3rST4pmz9+CpfvIt20L1/f9EsgbRqgooeJRIVummuIxXG8r+DYD/pB6q7EJ9HW
ieWhQXFEHbg2G7WRvbtRxpC5OkIXa8/5j3U1PiEmBe0csg1Dc7T0QKS9ZOn0HU5J0p4n6OLLsZiV
XBrcSy1ATLVS9CGJmMWA67GCASjhExR1TgHJGU4uIkLpUdaT78q7iXkmw5MY+zACtJkSvXoBu4MX
9p53I6e9oiaYnCAGBKogs2JFkx7t69Kvf0EI241MdDkR6k4dVaxTIERnS5NGYHpzkXO4DIo8SmkD
P5RIsLrpLgdasv8KFYO1X4CAXccYQu2QLVj/ekrMZLSdKaq0nmmoJk9sIakW/gEIp+7FblDkFB2N
XkQ/8uXUJSXhTxtgKRGJmT/Mj123U6pz3twFQKWImIR1zksxgajkSO3vPmtgDk3Vgw0xHJzTD/hz
wBn+s8jRsadVC5lql0Gp9233ssj3UBbls5HC78XLU6m99vxl3d1jJQlHsQOcRjl8JFLHpGGODNzv
RMhQhWF7vBBzgazMBRgz7wRIB06UBZfQcVxgf+bp+3Jhqz3SfmasE+0wTKLAt4St4mbaK8soHF8a
tRvoBNaIDzHe2IBuL/32vZkIbTonTYy6VAGCJWS7kl5Ho9weJGkGiy74XcgA5NX4d5y21hSIyyEI
4oUTPYeP45OWgSDmZKybCVyLLIIiIi4UVgQJHVo9fQeLf/wjT5rplp4evbkYkaIqUeJEAx/8EbSx
9X/oajD/aLg1DxfAr2dWA5mVJJrJuO4E6feGB02rC+TQegKUENSQSDXliCa5zvgdMN3hn9C4NftG
l+u2Yl0GlQtN+VX6x9g0/7iBJF5nTAPv3tHzLZQNLLy4mI7dnjCFaKi7AGWcVCU2gOugAV8s21Oo
GKm4d7Qb0OtasSbuGzXiOVuJfmIDyYUDO9dxJB4AvZ6C8x6BT+oZjHrPxRNCgH1LNYb+PVN/r2lK
NapT++ZqtTa7loJkuk/uV0tomXK3OXCPZzOmf8bQTmQmFkdUtHxfInA39rB5O9VRpUSqlu78JLSi
5Zaz0UkQuK1qNuz+2fiGEiWeTl3T5WqxE0pRw7nxSDpdW+59OJ/uqwU+4ytB5UOLTPnhVb8pTkq2
orWLTySyLQ3kLIW/l3kbpbbp2l6+9TI/7xSfCxBGlUZ28eyGZMM2kyMvd9fwAgS4EejJwIEgf7XE
1h93no7+FRU/63OMLOOWS4f6ITeMFSQOKdniDTM9l4GRZbNnTOW6N/0GNc3OoMzNMWroSa8YbgnK
gPlQAsu8nTnFridzjACc4mRyhR8c348X/Tj3zWoOpQnrIsIK3a+oa32gd2xGZJd2sFx3zJMzyiEY
//Cmq2DMHCm948Dpg9SpbPgtD1rC67NvNnh99SzD7hYBgSlPS9ms7zGavEX8rW6rUAN4ZfCy2F06
2eCA6uZP4EOUgtctQ/UiLgj4oIWd6sT2DKQlgqKpFIUvfBkH4SssBDoJVW1j1n5SYIhT2E0aYZDj
+aiuwjMPVsB+zPPT0xTYk9VS25cKaNAKdseAq2CgHXTSQ7eZHkkmsXJEqvmSLuGYde/d6hLjaKkJ
rRL9qPvwn+QmvfCqyjjjS5dqsz+9fgEzyxjZD7tWPd29gRNomGyyD8l+dmvMXqnRVY2oi4/PcCmc
0EgSkJf6Dor8cUJ8NnPyJsS3wpEQUoCM8Uf+yeBL9iD8H/hZiTJb+MzE2N/RnFqFK2O0wLWJDkI6
ot1PrzxFBAiZyLhH5Y4uOIdKFM8dKvIuMAejWfOnlUdfJLTsCSQrtad3+7omGdLO6/WiHbfjdXPb
1wfll/FPGjXUmt3c3SojaWKzNkh8JrMl+myJ2ufNuFjayPj9jto1fPWlHeDjQ1Fwrd1YAJgQLj1J
wOXwtRBPQgbBabdRLo4ZaCH7JeI8+Eb1LK6HOo7QwXCzpY9DBj/tW+bNHBanbZ4dejQl/dWA+7oU
2a7eMyTcLt4jYe5CZOACYNni+0x67qPPr1pCh6if21b89jbgkwEg8xwpk97lDY4cpzLFf+Vl6X64
HWrCtRt/1xNlp+i1+kdUblnW6IOzwyxUAkVb67Z7qNf5PrDEN8T0tO+xAl481yoycRq0RuwIoCrZ
A5oxIL+GgBD6TcH8njDuxW6DBmYqHJZdyJYBVZ+Y68Y982peaoK26RUTZD1SspgVVR0zHb7uho2F
xIlvZZbf8LXoAw6NGTPSHeuG9CSWYq1L+Vjab8Ias3YbVuoXqcma5EYxRII1ENtQD8t3wxCQ9/QP
B/DunxoKtTiiUjTnEVhwG/do9U0Kz8IpTD9gyGrTdruckD775OSbU7oDtDsWC3DnZ6/X/aTkhytF
udi09nVPSvNGYJ9AlfmLxSqTr1IrILNZInbG+nfW69NNb45r04oMeOC2r8Rf7+mJlCWcsaeH86MU
susHQz124W4ur/8DR7HQ3eCVxNstDrhySNv8ohoib3Rb9oDS30fcPhR4dS2VQDvSpVvsZXdZ5Kod
30SWqIlftc+WzVem64u/I1dMJvdq8MhO1Xc6oLGNqw+VUQYsXIn6eE4yJECpbw3Lv7X+uN+MGc0d
DYyGiXBPBLzh+UkQtWpBJHqvHq0ckAclalpEZiyWSZvq6MKPsBz+U7MZef752vuIOLxQJCDsUFYM
L+azeLLm+ckxYanfmXvQdCCTR1UwfcMHu+Zplwz11ancCUKIso3pdmh6RmeXaFgK72iaB8JkCChk
bz1gX9nYSaZV+ymk3kBMyrvrcT3SeFZLHf/7VSaO2CcY6ILQyicFXJbmRwv0MBkKcO0fUNx6fSwl
ZYSHQ/9ryEy75dhwh/GydYEA0wU383kI5oNELCzar57IkoxX4ksXexciPE9WUBaMOxh2he2zJXZ2
r3bev34FgoCE4Tpp8yHP+uQ3bVs8jckOmtGG+J3mJITxfYMoAPA9F1bzZdwgq7NoTnthHZmWPUjR
bDyJESBbR28E1UylCXLCK7so18Yf3gjuDxwp9pKP0pOUtTQblbIorz3lOeB/eyHy0puem5/x2GH3
XtUX11ogjPsIew1eX5ljkVeiyhHCAgMQWlTZGa72jFz69T34Zfrki7IxFpHfCqPaCyTmfcj2hKbq
CnXync6D6MRPwEDcpyuD6lHV3vbiCeiU7yxdzxUJH4t4P2wL1a+FNrhaAC6rFpnPvgDAjyITDZ7M
xH38Lby64IgesEu7dkRvrfJHFLcRvUT75+a/gNdO/H921RwU32Nj0/tX+pYWdpWuVLloQ50R9KSN
nFikJni5DQGwxv7rtIHmRgprlGKxp7qwE4lyw65WmMvLmD2SiPatZrpctFyJ+GqGXuGU0f65jdKz
150WfAlhg0FTn5DZOOZFyJq+BOnLEagnPYYWTHdqxi35N9Bj9GXn2TQjcG57789hhRVAgBmHTPHR
FaoPak11n5zP+RWTgeYXEeIQeRPzlh8DYofwcpLwAsIrrYv3YB+ElofT08e8FL3dLEAV1EQzNbsj
gVXMGtAPs2gy+CX8XkA3BG2Kdox1uvPS918hIOia+CEm8Y4++2lgTCP5l3wvKAc0p4bt8RVq2k4J
O5jt85oyQMdosL4Bt3YVyCPdTweaA53rdx5I7WoYlJVrjY4pzomVygLL+lGfzwC4IAqceaJglpZO
LC/KLZdO3r6wIr94iVfBIKkcLEYaCC3S6SLttIoyy6Dx/IdhJnUoNxLhF5O4vjWFnpDwQ7DW78di
MDtJPq7+KzZhkLhHcX7smEu8y7PrmUx53AOypOeSvLqKRYTPX9PQWE/C+1v4icVFbZkSYQG4UrK8
U0AZyscVIvW7F4wvaRRo7k215f7/T5zSbJ1rL3yZcu8hlQCZjKjdMH4FN/ypDZKl75KHGg1KY/vu
RVoW15SkKa9OTGOQn9rRlYY6csCMey0XsS/XVyrMM0T7ZHnpYa9EwY8G0ZdrU6LLX6ZYmhVsJd9P
3TGUAavyACM5unJfjG9yxD5Zicx0WB8rq94HHMkdtVAZ6VvzfqmpzP6wBaqFT7EnhfDVJOfd2yEj
c+BjzbBdp/c+BrVQrLaEd/VzpuDc6lpx27BAvy+V48K7sTKjSZDcyp9gbq1Eq/FiiChklA9RtFaJ
L75qFXWWZYNZ2kWgO93OJDMO5NtpgRUxEBrbWPl987RBWYK4eizHZondSFDXOCWGgJhOzqTaaRpB
C/hUarshsHoqZmcm33qXJf+6RF5BsUIcjKejWCQ0eKefLxgtfGqZQIJMbu8yZS5Z6Ip9BLj2warw
zCifHlq1L7wkNwZHnoMoajdQKI/LfDmJxoxU1yYjtwpYDTpMpko/WO4fHY2lXUpR/cMhDT2cqTHl
4+/uDFVhbYXPENaB01z58DsbfQ9Q4EkfiiSnWKmOAgVPDR4bl/WcC3ttOdwf27LTfOIN9ALiyNpS
QFUNOIS+xOLSTcT5F7YCmgjwVT0yzOFKZnE9WF3DeZuOyGQ/8qfLuLO1iN8X7IzTSyLKeLoGqx1l
rZgxT0PBXcJQXv5VGyYWYT/iP5q5RSUKMbshuHzYZ9ShIYoAIcIrt5v98draExZV8rgsvfCB4OmQ
0YqmAGmk5q353ctHK3XU204/sBUqRipDBso+24Jdbv8WibCeybvBB6XljX7GuktLVrszbnFb7c2E
LR7ZYkO4axow5OjPRRjofrHvSFl55XXf6+G+S3elB6mHxeKh6JH/6JiiI2YXWcfVWZrcdDo7lqmu
cVWubg6jOKnN1QGFAred3cZaBKJEuaMaQwMNhK7UYjlwrid7jFYBpfHeeiCJN/Y6Vj/YWc++40Vy
/X3qI5fziqDtnuRUGXrgoR8IDygZgLLwP5iXCnq2LEl42FLR3Zb91T/MVKbZsX/MDlfi54sJNR4v
M05urQPltXBJz746GE+hUxtmQF4d0DZOSaqeySCjP5o3Nxs7HnFBDTO+gHtFady0i+CkhqvSeVJI
W7CAtI5uI6T5y42T4W4juH7qxyagblHxcK41NaDlBXnJ83YBdFSZXYPTlBe00QF75WhkS5lLsXrk
z/nfgCADVsGkGLFKCKgUjl9P7U9RDZ5BCa/wBImQgnfn4hx7oDvzzOEroLWU2nOY7PM6R++X9uau
IVGiNuvmW4+i+bqNiRkkgz2ob3ZdrwuYkEhg0aruCor6eO/te06QkCLUnKqZ04LOTpfdEN3/1mze
jEF9MX0dI72qZSv04G9GOqiXcxrEXJrTlbQQYHBD1YH6gxJlXseIWNC9htQ+jU59iNYc4I7WAaZi
htHRwkb5OJoiEXHstcjvbFoB2ssXVmTuXfvxtquMdCmuAwRtwAE9I7HQkCBn/yDfjrkJJp4XzWgG
8ajXvMYCZVXaovfSnYSa8el+TdI6x+RfeRXDVByOkDZylg0Rdt5D4DtG1oD/l1mZey04UJEQDfTe
wlL6i1qEaTY22KRftasjEgwuJGYzPZlgZUU8IXGK/5WaPABXZd+tG0BNNBP/cusDl/FfMU7tDW5X
+KVeVZExGaTRVRbANHKVoPPAKiF3FbAnWwNkvNt994tne+FLK03BQha+7tyjFz6h+CjMOLJJLj5M
OPttLPsBynUmcfUOHW/EqRXohHYi1ISw5Ku9nm25ZJv9GEGeXLQX94uIqBMccga2CycGbjquxt+r
4ADVo/mwNdYB2X41fvyOOZwh5iZUrtly2Rtg5K5hc4Ihik33/eQsCddNWB3TT6IxeHxXVdgSuYU8
kAHJEO62bGQp4u7l0DRK8AqmTP6KWdRESGij+36Ps45JO2Un5ZvveLLuJMoachjnaQuYaCysXaCE
YQWAdTeDqHiur6pXz9lomLoGzHNNDCIfqKNr5q7Uat0xXrQmWeZnkjgZSec/eq+gfOV/FxfFSCnv
jwEzsw+s9tBmmHKwzwVMJBUrebsczRb8EIEZ73LFQxHUPyvKXVEa1GVV+LS99qm0VHcRqqnbVApX
0mu+6JIyZdIgmMFyJe4xHsJoN3eNeWEpX09I7zNjJYwMZCv09tLaWSUhL+QKW6NHKm1RXMdTu69J
t9qyouDvTzCTlx7Njgnlo0PUWmo1JyRk3JJ0B/CWdFDnnOfAXoBkw+fqUdgxm6fJbNtU1WnqiOgW
6Gl+g4WB+/MvO5fWTfTwAgb7GwgMb9Hxyo6gvbZ00WRSYqeZgn8UA9ukHd2L9NjfS99zhk0bh/D1
gspAwr99bbzc8v0S+WGowcDmGJgD98Evw9rAtQyAg+P59PLnO2DKD+F8kHSP8fdDxT3JhMAXeNFd
3ezEZF2Bx2N0ZvXNsunRV1Ugv0i48MgWjd+/0vM3ToehcorWw10svoaY7Uhli1bdxeenpL1BRaW6
QdZK3eixAq9RN8git7qQiz4KL/DqeBjuDGeXoMMCHm4wWrWXlwIHNXvTwXfnqnjwozbMbAVyq5hg
ECfLouUmKQy0PW/sqccBHlUCnMbXQgwqjvMMpAtB9sz0w+YK8+OeldtAQSE6e+/ErEBjyGWVtCqM
3qPmKiGK9mGhjCIMZTO4/IFmckGHeMDQqq3sEDe7RbjKoBfCPtkfZbZCSVnHxSYaqD2MzZfS6u5r
xKSgudGjYScJcKoLyc9GHM64a2Jgpp8Z9Du8KWZwV2V0O0Jl2eLQhjwph1wbSraWW4dpEwpdEuPM
QAvRgX/8YS6S8NxGaSaWppKbwJc9LR5klU+rg58RrutivYwM3vqcujpoH3VZF420sUNgQVC744dp
5lkk5/jT8MqBjXuM45pJIkr1jGb/+VHmf7H4gvcXRgG/DkfBO+0bESw2MA3ocGMGZahHeAgzqcgM
CHp1NQ/zMHnwcgMH1QIM2N55YcYhF2E0beV0TrPGG5mTZ5S8kGhmURjb8ZS1mLF74hOSu02L0kku
XSqUqCjHtToeXV4dnaU3bEtkqXP+6T9G4rR4cZHApshElCMm0BPAdRqm50QH02pcR0o+WD1yjPKR
4GgNHl4rhX36D81LGG1wsBZWlue4XWjIrpTjfMQosbm0yqYnUv8xi4rnCbEtzfcNmgtePY5fURU3
ksvmwFcnQvtM4rnkhEnqsLX4awWEieX7b7BrAEvi9BD72niWitApwtL4kkV1ZKDlIJLxI1TE6FxV
ONX1SrHP7jmSddwAH1VecZUqHc48H4l1bQIJ9n0v7JKm8eba2t69AxMOlbyOStXdifHqxLiH2LqG
G2VBjjdVK6kMiwflF0bT7NVf+8pVOqYPyv0dkDVxViva9C2XGwD+GKjDLw0Im+HmDJAHFgkWN0NW
0Hyadz7IKvklbYSrrtrHO/SFs05ukTmN8rv+uSG/aH9ttnBqXWuqDMqT5DwETS0FU3svL0y9p+uf
hRCRC0ntphZSWMncqBU8IZyfhxv3KWwyOrVR8oKk+0dVosfxcBGWSt92mbT66WAjih1EhNyHkGTs
FUdvcXjt+nk0+66vq/G+a2fjH8bbXBE1DpSSDFbYqqvDij2P881aXUqNvlo3a/7gJonq1r/g3oZX
8gDEo54oJJ2A6QyQT4W/OS6hQYHpBPyxBGg/1d2gXVPJpSm4zplaZj0p9ceh6m3aa8tquCsqesdw
DJ2LGHDo8RhX25ENM5TrTRp4hAW8VSgXCbLqSO5612QbdhVOiRQ0sscRd7WUisOW9G30Bu7d3RtJ
Fna3vzIlA2nZBpnMhMm1xuyVrPEVstWUdfcz4ZkoWoRxO6ajs15mR5y1Wj01nkbr0E9HoOLSkOe4
UKnhjS6EafkHNYuoFbwTwlrAB+R4d3z+9fXuAlMKNVPvJpTIw+udagx+CYtpxXCGLyQhUur2u1u4
lXwgGHNfp+JgZHbSLNE248U7PJKVVFQ6rJhBGyu2PjZL+2ZxVIx1gHCPIVzIIvf2rkrJiyGPOzNL
y/DmG6nPR09eH08t7ewNAVXtFAcsY4mPUmvYy4g0L6YLlvgBSTdYNIrnS/v1Q3GmFBJUgEF6aXIt
2K6WQH9qE/3WwV3BaeocOx/iukIK7hk8dytxfF84+nNUpb3lB2kGmKDPSVVeUCxMzpQq+2pzr03C
noAYVf9qm20h/OMg/cyW/bkN1lACDYx7Q4Tqe8Ihe9lYmMfQmZpbQ1Mk1FBFnPJBWhFqjWy6RN0k
+cUJSwd9phTEO9O6Nht/chI1DiF8TNST3YsDAvepXII2HpV4Hn+Oazpnn/8Blp7T3s2yO/JubaCB
3RijTuXSXM+Zvc650s3WaSb7yJHjHHLTqjOiFPKsPu+4UGQT/TxPv5vnVi3XyXs3bGvdSMXQU9Xu
RYBcPSlKe20CWZ1JBEkhn6Q2vqPk87rz4JVHsPrCaWCrk+2ZNvLqunzuuk19gfntLHWFrKVC2GaO
7IZDfHr4ZkUAZq79VIrkjM5n3ASB/m10kJgJriIcha4rNHn+AeQwUVWnfFpGhUCKpCKaReYFGenR
zgrsF2am3TNZ0lmscMn7nMv+psi6tkEQf0SMv2vEJEn0I/mbl4wA22JoL3mqBe2uvCte2nJBUYZT
P9mnxqZgKsSj5OFri9nLEAZNZGPee7qd5Qne8TkdhG2WsW2C4EXlUoQeCz/IuGAW60KMJyaMdm+w
rZtXbwi0oQITzO41HyVOnM0Tb1Yem49SPUkdoDd6xFGO0gnTG9gJ1hKeWuglgw/Sgf4MJ5Awq8Rj
keEZ2cXO4Y+k0IAz6t+3Kz9B4fHhZgV+5JnFG0HYujYK7iDfU0BuTiH47dom67kdEWmajGim0+sY
zF5rlPVp1dOttXzS4SbIAuAZLzu5jm8N6YQzcpZ+VwrrjNYsRWmJmxb/Gu+rp4uLjY54oG1SwjLg
Mhua3UTRF1ac1SKIFvs+QeyM2jF5zmvUwC0V63rBh/qiHivIvxeiuIi5OpwvS7xhJvJmDKC69/yf
qDQR83Sf7a1rs00jDrwiCzYlqzvpNjX6O6zwZ3vSVNa/kBlyeaXJGHGVSr3fBNjPoenVbxNfR8Gg
Yjw/6FyfaJs/Dt8yt3z6gTNZXrDgQEjxhB3W1HVSAwLFAaayUCaAcyMWteNSRjzvLOu0fGZh5T1g
lPrbi0O47UgplnEB4tiYTRDhjYAFI3tcCYaW2TLU/7WJnNIewD6pqE9sviUKdLopJ/tWGw4EfPhY
XLJL44ksmCSblkcmVDd+jMTSDPbW8ItRcoGyU0QnOBqJUXHdCnF8OxeqRkbPFVvNDkaB/SNBR//y
JubvmpQO3e+drdNc4nrvKNmK6Bl99YOfKopU1ARwvkR2k0mcQKt0EC9PL8iUTkRpSTnAYx0vhQNC
Q6EFdUhS2wsGcWeQqRh/sIqn/9YCbz6bEMWsrNbUNvj+hH6RNWM0yPkofE+9j9v/5d2wvU6Tu0OY
jdOP7NUX68J6goPHipDZYPjK80may5PeqXKhsw6fdrHdXD8uUC1xpIbhCRLNU5eIChhbPJsvxq6z
8bz9z3LWknziDHtHkfhOJSzLBelQPIVXhsYgCHK5fcmxFjKXpFHuZXvAU2lJ3cIFqhjw6E2wmSis
l31wi02k9iUJQKWMx/gtZmd3h22lOw94xjSWIC6EnSAUzZr1EWeE5Ro5t5lBXUrjzy4XLE5ZtHCx
e9zx/gESLFq43JYWntFolTTYjgx1PaG8LSgrk5sMd8xEyr6FmJeMUjWmCsmlOVY0oFzcGg3fYhTa
5AbLJ+5NLe8xKR5cCh44P10rgAGOIZOxXxLl+51DgQCv/0wDEivzC7m+7LtozWmVnn0zfhc2gfR/
7MCggzMngG0sITT0nA1EfzJHgShoJBmV6cQoJurOdkJn1DtjcNYS2ZBMlvEnsJ98qF9HkpBh5Twp
UK+KD+b/aKG3cEXGZJsZiZI6vadrEzaZB3b9MAl0dz4UcoFb+OuZcVJSTtw5ECInuLW2DObWW0ue
w85lSx1zTV+k+xwjKAH2HKHKMI6rvyehrladlvUt4vPh6J+QYotPI7mkuC3Ro7ZZwaHOabFgDBAx
IVK37jjopxDmJPGi7eL9DVbjRyM3zuoPlZk9w4PNdyvPeWGChzELxa+YWcqfYmx+e7XmWszTLLsm
SS8mC2zcc0B0PnwwKPnIP0NO1eROBbUdWpDubBlYxLFOslrcP4eigJY4N06VbMwTxK/tKNBhI/Xh
fGV+14V4mYvXYCdCERNh59cc4FHMzfLjT83YLDUVp9OStwqMLyb4JPu7uOxZR2NOo8XLGNSqhu9H
WkJmuNXPcMoKfSNwNANrQigtKnyJ1PL1WxoeypCh0e+yKLWyCNMyEy6c10SwAK6vjkakfXEbHKwl
a5CCQqEbYB4deJLYHcY01w25bcLkD4w2dyg0SQCSufgEleYwKxkj8uPZ8kty7kWqItcKzye1hwoR
+QCF2KRySuYTphD6etnUqAUmP8KIRGNaXf+4czM7fa3T1cnCEBc0VlzC7nUgAsNx0VG0C5R5wXkU
a2hLeY/D5b0ppue7SuRQGbouwbf8kWu1PeVE4OaWrlXYiFTlKor+xyKI8i8jmElTU+UDJZ+GCzl9
DPvTyYzW56atwqktOPd1W1l1BhKU1bdcJ/QZKkVUEimTO5mkDR8DUMeSX35DrfGPw/iaxE7cNBdQ
48MXCkJ7RpJVOB0x5HorSt5A41N67o7L29y+RU9FX9q8TSwatfXjVkQB+09xax7om7zQp1cBOPqj
RWKhcemWDifJ2SFeIQ+jlNmCDxV5zf1VYwclw3kG40OUtGLj4LssFmRs2n1cKGO4644PJCpnympb
ojqT9IzGNI2q9/LqVwXSDFLSEKZZKKEs3vnjjRTXR0jsSQ6Yxn1puI3G95QWopVuz8aSOFWhVpsh
EThtOR22saCrUNWD2AueWjvFdT3354ZWSMocmBRWSKuQsWoymIyxRp3/wvAGVSkkd6tWtE4MBo0f
ew3UCoGmGImGinjr7D39GcJG4IpkeQ+4WnV+wx9ZX+95JbBHEGVLEB6JcP5SuVBUtpJkhmkYmteY
KTQVlALazwFR9V8PlGECzQal8IFmahikfvrNI3shxMlTx+G9akB2gtmb27pkNhei7WSSt0oegVLK
HdZwd04IKx6rKx2YIuP7BF+p3Cvyuya3eDfvQF34GWZu6J7w/O3hFYxSpuaUXuJJd3A+u380Y5Nk
pfqQN3S3W1l1f20bGeHKWebQkrcEebcVEanFMGyfCvFM2p/TORZB5XFcelYwefPQ7/vEd/rZF4AR
uMzIw6tmRQAtt9LoHFkCcb2qCj6dbpdkKFFXIpQ+ZXitn+pN0ZSCzfWV9qDtfdyjTC9qBwEo3fMg
uoYRRzka/xwhtI2Am6shnRmaO8vXIrpk02EnQhTAK6ZOakkUD8BpEITN4PXJLoMeSLUX3Oio+Bu3
T+SIjt5TSt2iSBF162mbbUpMLR1f9AOtvq05Boycsr3h10FD1KmI/ZZLTHKScXOQMya+cjNBykIg
w5ZvNssfvmwhX6asPWKPl7aa0RMwWFtTH8Xsk3RFHy3SzMEhJ3E8N5fbv6LGg+eRDDMJALlT4+jO
lhbTC7SLhvMVzWikTTlxixiLJyTW8/g9w299htnSp+v/m2Uc2BxKveX7IzOoJ0XYi/6pwkyX3uLP
XOW3UPojB5XgqNje/GWznm1VHptAN1e6mcJN4rsTOtt4v92aM0r2YIl98BetS4rh2lXJjALcF7hc
UkirpoRB7oO7pnXM/fgToZjVJ/cH0fnyscOwYSXajYmrNMsWz7C2np0N/nJ5VdGdIYWq5UnE+pFd
KGbkvNn/T0zg485a3v7Ns/ng6LOcRJ/9TCnUJbH8YIjwF9fq5fAEAgQZAVnasdQlP2xzsYKkOeRZ
OD7vF8VmQ/zMcxLHBekMkBBVLeyoTKZtysoDQypbyn4tGZUaqZRk4dFAykXivQs3LIuqihbJsdCw
kVeohZx/n2brpb0gO9sssUOVFrD4A8SL3UcoC46Lhe4Xp2v9Ywoz0BEk6KjD3+Eo9pOvJxtf1vnF
5QYZLAGMNuemUI7t4tO3bJb8ThsTeGFij8LkE777A9rxcqE/yen4g8lAvVRsIbJVOFeHG8LgHSuX
GCFUPUftviRB5HGVcF0nhRN2IEOAb9Cr900qa/Unz9jlbYZedcuFG2liwxkx+dqTp74kYI9jZYgv
ffGvvW3wSEErEa0dfsUcX87g6Q7vZbkAvQrTB3tneR9itcIPsrolhYeNeLge1DS/tmQrdT+toPLm
JKrdYeEgtj1q3kUkpx11H2bHvhyEAEmLEKeq2zTrr6laKKjvByjmrBSNRljvgeXBIk0Z0PraHHaZ
B5ckHhY8b7I9tVlA/N+1LumRNSm7W/0e9AiuR3GU1q17Pkz2DiL4vf5fD2oGcCWYRzh6UwH00Pg3
uprGCGDKe4qCw3tS999TkOUpZBbaW7moh2i+lsPsygveimZH+3gJdV2jZAdGfPzrhyVJlbvpdihq
/UzJW/Gqm4Ef13OYIp7zaGHrLkAVvgHKuPWNOxAWFKKk0XPycC59MBJTXHQdKTICmbLboNgFFgcu
rrAD+FGam6gC2Zs1/G+5PUrETMxblw8xKcaagS57UxRb7ruEoWxFTr5ddWYrS2pv5+Zb6bfXuWuI
LrO7lTga7rJLQEAIRTuGo5aSFCGX53es30A2BiJ4UsSYWkR775KvCnTm8A+LBykXgztUbjPOkx5m
e3Xhx8L26iZsG0LuQszEdU0I+qOeq2D7NNMTa8tLNBcHUVQbL8POm8uAR4M/I4z64i9xr1gbXiLk
4k5CMv9Rhy6870c/+l2GdqgizKLFqW+ukjPszhVXeVXLTLCypVwMmfWxETC2DC7EiW3TS0LRdnWL
V0oYKypCMJm/2sRsV86wJjsOnvM1vwjfgA+RLhilhUyU/Lz7Rs+IRkFmZg7356lfIzci3o7hp7Fw
E+9xe/V7MomoGqZz5GpTrn23xdZauCroArTKStjEp4tpH8pyfa3NjXDHWjnVJ20o+zjXmPz5XsfJ
VNs3Wr0MsVV7OKJLcGsbqe+/4AWFpzswHCVOdB52Ahgu2tKh5OWUe4wZm7mt1uvp/TWHoZEMC8eC
MmWPmUNlt1w/Tl76H57jG9i9wMp3Y15aZg8o66sQeHlYp7/DAWR+trYf9OMwTxLk70iT9Xf7fYFV
+TuP2VAmQi3gUgO0yWmEFZuEPQV/NBEPw6z7BPXDbXGVG6yF24BvZ8DU+Ld4cpYAdOdnmX/AZaWF
TEUodsuy4vOZUhsyNDmLEcjHs/jbFsslxFWMbU/w7bx241iYgYqzl71+7Hoy56RcB3hYGpmzvys8
dznjnK/Iaap/dTnJzJ9joPhh95U4vzy2V/Q2bzlt+AfIvAE69o4JyDMy0pzkTe3NQRYNQ1Prlx3t
c+iUhqYmrB9HCTUvTrdkyE9Amq+455/EMzHAwrOrlRKZX+sxiJ4wIt0YPRhwK4swae7P6cWfiLP7
WJTdZiLOHDQegmnVY2hX8jlVzTjifSvDPNMbh1oZRsu5olTLegKwwfEHgdMZZa8NrQc+1JNOj/OR
fvzlsiEGnFerG4unVOipVKTb4etbogvvLCQBAuIreM9mYX8q44anqTZ1PTiT4duct4J21cIQhO5D
0TDuGpPsEWJDaKUCTgLg6z+ZlrJnE/g23DoJ7CgeYNef4X82aSX7OoMG0/WHnb7dTWSH2zPfToh2
hExQRU64N2AqaU0hYLogAEZxUCG4dwDsCK/pcDk4pYMBXpuMMoJbcjGS63AeuYhKS9pI/0WyGEOF
NdP+VLweaE4gISNxZ9FwZEpT1WwDNfRj5QF7PBt0NxcuG2KwhzCanF0J8SBbIiiGFLhIVhEcspwW
v4hPh8bGXNGRsJKRQyZpIfD9BGedqbA+QBUQDOkGuzDBggDkq3RkzLulecyt3NgLm6/HeRC+U5T2
cPCzjt3bdlNEdcENdEjjT7NXsBUIY39Tcoph53d/PbXfuuE37EbvbMxrtM6Pj6i53o87aJac/sPy
/jOK0E7ZEcareBduhxvF1RfDiqWG8QH6UOJzVAigcZ8oChjio9OM30ooz5ztROlnqJPDnyq43DlU
DJqNu4D0H3R+zQ1R8Oe/whViIfL0v2DJ6bs0MfyIcTww4vackZ6vlIZkNxWr7rGVjSkcVjfF8yCg
rWjtqrR8MQCLC8haxKhiy+L6q9WOWdd039mNXQ/+0R3ZU++Bte34Ob0NucUOZ2lJnV0Wg+OyP+ft
iRts7/FhhRVtMbtvYPGupVqlu0PCPnB31D8HyekKjlTwJAlQ320c5G6Z8FH0M+of3EGEV8nB51xo
VPBb3u6fh+xO7d4Eh9FkBZ2Qt0qzc/aEWsKD4M5rKxYLZYmvWji8yJwm7Sv1UgjAa1yL73dHV95B
GGXNYD1Z2+wsXTg5qlDnEEU6uZMsZtxjT76CfZEWYCmKbLEUJNB21DzV8FlGdVFwG6h8nxdVh49p
4zwRJcu3RrOY7imtXVhnaTSy5gwG1Rq5EeJc81ae7YW3SNtkVJq+dbngz+S/NE1xjJ+NC7LNjS/+
UHjZP/N64SHNzvAPw4Fv9FZN1ElehCSEnxYsbXLK1/sREcbppduxCkhnH1Z2/uQudFx4I4FFxFJF
gbPfwbeLNGh633T1EqBqzgf1YuM/eZuR3MOfjjfGYdrpaJ6OWcJcqghAWyVJ4udFh8t2sxoF1Euc
y2TtRRhbzSPWNm5eaVuo/JMeqwkTgaEZ4zgZx2MhE809YBU3M/kxClfVZdf/pekLBiwSuo1Nshue
BSTTD5pPke5tJ88QPokU5MEcrtvil7EQGqO9DtidkQeHdeE2msv8YhriuphRXehqKFc0VxJb+KBl
tceDBvpllMYpfNxhI7NC6PHQYQoybXLhpq6P/NyDE+v/nB4whZFW90YoJV7lfxL13LkHcyKEtu6R
M5NyJnwvuwtBsNL1nW0g6EWD8pZN5KPPnUR9YpNF0WeDFwvimAD9ykxbUl+pehbspT3UI2bxhSSi
ZlDFH0omT/TfJVM1M4H7EnFNlCwzF0Zlv50Wa9hkfKeXzIPFJ5ZmrwnP7raXUCRt/JmZRkSpifBP
VrZ6sZ4CKkvRHc3Z+YPr4Zp0X1HbHB98dTUNi3PgaIIC25S+IAwRjkXOIaOYHHaSNwPT/sCG/Vez
hAPiQDOEZslyhD8b3P2Grk/VjhV6npMVlkVHYHP4mcCQ5ReJ0pIrvNJMiuNDoyKHosw9iheV0h1t
c2VNzxM6mJHeR0ec8AOWKOMpau6i1RWsX6SPO2KMOjXQwvDnf8KtHznAMmLsmrsksUexW69vGsh+
JUA2M4OND32himS19h/7cqQ2ytfwnaFkoV7fBpqGk3/HJik4m7xX5wfeLiNQ5bjMhvy0Av/oAmqe
bl8Y2GIRlbfy+XodkTxx5VwwwRc4rdsUFdy6LoidHJqwKa/ouJZdHioybICDf8kXmUpx2g1UK+tW
2Jn7YJzrfSxs93R5hzHGbTbBZHQt/mOnpWxZuflLNksM3tziiDdZNMSKXZHM2UUpitSUe+i9LLUX
sLLDvvWSpEUmyr+U2u7C1g9VyUxqSM497S+69G+09jK8NXwpFyGxwaznqIShKjN5/ySwGxVnnrtB
jPCWbOtVsZdghVmPsDHEM0MvWF0ZsWtcsdWlFJTE+vnmOAelHVugozJMtM8USuOIy8erPvS9ZLAk
K302wWdxLz84l65vcDX/yi/e+skbjWs4YmYPZezm8G+R0p7H5C9wlpTqbAbCvdj975twigvbMQoa
j0RTHdVPCPJ+OM7Dx4itGiY8W+HgjQ/TYBZYU4GLiEJk9vGE4FrC1OqrpexEkKto7Zr2F5KnfiIF
DZR7WoYNNNOKWvMaVPMC9Ciw23AbUMj39X3mPTmgZ1kcWf6zXInbK4CeFYgsGN+QCw89kgvlwM1x
UK+SrkgAr8ApEEGg3f2eUEWQohg01H4zAS6JbaXJf75kmXWfzMtkpL6EnqF6I4KSOsK+q9Qq/U/i
YOPwGBF/HqnaM9dzj6cHCSxxjRk6HYCrHbg+M7piOw5ffxFTNAvhlJGd+khqqfB4kD0TMQ5m3UOA
LXcqj8kYKhpA8L/havepDnE/otYDR3+JBdgB35J13+x/HNPe2QuxluNbwjn0lULS7nWiWMJYMrrl
N/ey//pBaJtg3UWAgvZ8Ec6PF3MfXX+1Mf4LJ9GCPbJywHgAAEpzPjRV/Nz9uWd5lUlSUHKmmAxr
8zY5mkHXXThi6DK9lBlnmwKDHzVRr9U5ZaPc1/WuenGvycgMGLtH9OQhTJpSb99CD0mBcQxumvfc
LozKl+a0+LTcguz+X6A+0uF5yM0HyxbnEu16WI/rn46vB7ZyLomxf9Zdsmy8rqZYJzx0vSrM/itU
AvIax7To2GevqO5tQ1kiB3Yo/7rIs0Tjc9hGDqABXY+IaieruvOFLSmIJXsRN+Opg6Y/KOllCC6U
skPMt7iia3gLJSO8GW1tiNpsYaKgsADJGa6TbzLf7oHZK1qSsjFvYh3YuYTW5Fo2GXEXx/I0/T7d
Wcfb4rcCb2DIW3C1UFPQID3/rcUj+suctqECmM6G0QlL2Ln98q/mW32pviGWhoF1MYs5/KVk1CfM
LEJbr6ua4UGLTMn/Nou39oSD8wRh3pr7OonGoIoHfhiLMV/VUS54nX9ysMzg80s82pxxK6sAgc3h
Xsc0GQVCU5AmnMsEWt4nD7QTYQtWVPdNCk9qg/9h9/5tSkRRrhFVUfdjQiE4rGvDsmSFTE4M1+2a
RHa890gRfAkvnjZlwOUi8IL3+LXoeCSw9Yt9b3r0vULejlgALxf/SDTSpUtz8ivA/dQiPjGijT8h
aAH6oiw8hn5m7iWLj5Dn8iHAwhmILJk72HClmlwn+BbJP+1dZx2DPlKaKFA5vj8hkaZzBnRJDaj/
p6YQ9H2a5zcFuHp7cpnLk/F5Kn2DludATV6klA8C/kmrMlKO8R+PRCma4nZXPTMBZcBNhOFDaUTy
bUDCAHGJvVGEiIuFuxp+TU/BOkB3X9cOEe/sG07h7xOHii8bbgf4aO03o9U1ytZAdILnA8om3HBj
H7carAdfPfeNkfLM400n84iI1jQR1PASf+YaqeS/Sd+s6S9pyDvsOpOn3qHD6TZYv9bbbu06CRuM
rV8/h70IXxfRaLEYUoczp7zEbpcwvimLexMouZUXmc/n9jB/Pe5Vz+7Tg4saPM9y3CC+yb3kw6T/
ihx7UEB5JJaYiXhyHoMRJu5H+4K5DABmQXNRxE5LAJcfJxjF08L7wGKsOYVcsYpoS6Ky1XQrmIUg
cacdzHdQhqG7B+kl8Vh4viTLYMdFciAlvuOpWOGEjZOWGx84LyCeYR7gCnj4M+NO7n+wZpSNayNa
bT+cjw93hcsqxg8dUCFpXRwKeRnXlmO1m95LdBkdaLxWUGJymT40ZEgCBCEbLiDgdBpj+JZtN6Fi
PT7gZGK30AKAY/usAQ58g6XaBsrUoJz7DckuccXCxW5RqDHA7Oi6thG2IWV3mjq0KoRYVWlI8fbf
7mYihVDL8/zJrFsOi5SAz+n5lVQ3zABXnNoY1YGW7wFEww7xlliiK0blR0QSlzwZkFt3leYMH5BB
zowbaFFfHnnL4izyg1Kjh9TM08HIJfSx1JOkY+gDxbLS+f02W+FHZJbw3CCuaEmMW3CFbOgN+ArQ
I7KfMsE+dU7rNZq0oY1pvlF236/6IsmwAAnjcGGzZ/nA4xXRFlGQleI2hape6yS2yRiVEvKM3m/4
7h9q+YKjlXMUTeQ+ZG9q6G/rT/z2OeWeUNV8c5ptq8wXkcKEVrIcnpFm9ikA7GNuy/6nb8dusQdf
vtAjkhPQTk+q5jHv0EGOX8a9oC2KL32nOmHDUDni7C81eVdCgn6p4xo/gYeFWRbKdx2ey+FpzQ3P
8Fydf3FFc51Y55CjzGoc5B0Dy69tCCedB6v1Otx7JuXNlV3L72zYwx/84hdy5o3qCVswzPtjd8Nv
Ypw1wdLjJLywxeNS6WwNJlwU5Oyv5z4LJ8wiCgdkPwRCI5k8ueFrrlZBInWXzusddTif0jWG61H6
V967D9U0Jh7/biePY9oSSfsBnM46jJ8Vu3iRKJvuwlsLEjeBhyOSqr1K/i12sLLGv3S0CEmfw+KL
v4IKoKnAx8mOhWvDAwvy3avbOQfxW2me1mQ0KjsTd1QyssalcMheRfOL/Nc1QEy97DhcVx1h9zYp
5OOH9bEJvzLFgiJL9Wp71Z741fvhcxbNWq2wrc6xXefy6ob3lwcsuYtKSO4glv1Er97fpJRPloee
5NNwd7qgZ5Nq6oezhpN2HXeD12dcouuQP8t5is4bQXQQWxgY/t1liXCRyLuj1Pzf87U54yTwoLII
aUTiJ0XMxTNx0D8iq9cmZuhurRJKqycrQqikpbNWPNODI590iLRDZUiD3PJvCOOXpzm7e7LwntaB
H1BANFMkPlUdvdpDSGDqAd3Jt1mZu4WYzfs4neoWPWf1It9hEwggkL6wz6AyER55V9fUHJHQk2lC
YNz9CjCLGYKr932oTVaQTxPzmEzYZLjLIrLhDtRfDV+PiPddI2nuFr8gd7FWgkhCPgiltZIFiIvI
AjQll0F4Cfvyydz7bkh6QVGBrGE4NFAi/7AnoCBwzy+/QiIAj8jWhGsTBX+NMTPlUOdCUP70ISPV
vSBnxCNISQRSpvMReILav/SNnOlL80aloG2r6uy8NqpZuePGDHlqt43OFey1bHzLgvyPBi+gvRS8
SvJOxUrODt6Ar1+Kb6/LoxfAapjahhhARdxddfLXSMouDcPrRbMY6Y6ouIi+VzHrx1wSKejYRZgf
ddzBZ8/jHuHJSzoDApImMr//PjnAmVDeIy5weJzqMvqtMQCNVnt9/TXrfEUklFmVRRQnC5sn4WFR
tu7jzZRD3yEzEUc4RIiKA4bZz2QWVM1ubzrJZ+eNvj5FfYNJvCSUrp3Q9UJP816AUPNkMVhyYxmz
XRKGVy1a+RCa4+jRaubUEZEEsb7a3iJ3sTWiXPH95kJmPk1jKBa+jV1m/WvWSWhieDblVKfBVOBT
v7HZ7CIZmdFokJNMIIGNDhJyTZeHwzgZzyR0qmFFzoqw5LoKTvaecWxeAHZObvoYhPJkdk2925Oo
1wOP1vusBNA2urWBd1aWTSz/8ntX2Eu1ienKtPOZt/aAtBqFNM954+CUpk+zxUXVyOdIWLiIPtHn
hb8ytdfFhokYv6sSiBLiJyRkMalWwr5I7YUDOnUgCBaZg6lhqJ4DcpBGIgniSTEdf3aD83K5PYSg
SYxP7R2nDWlvcURQ2bP5v9GIaRXxf/T9ew/lylkC+tbhmaiXpUOod4cM4tGo+jn8YUCHmKTIPsIp
YDRgxMC3JZYKaqhzbLf9NZFY/X8hi6kB9c35lfhwzPYoT7SlghR2oD3NF6PV0ptNP1iekMu4rl0O
GPZUXvmjydB05Lw8X+hpUtWpacq0iEc6HGR1BNHRS2SR2VXGbrQOX3xwMQaLpjz9BtoKgOSy2kUU
f8ghAnIoVflPp41FwgdqcNgMLYzMZONgrbsSlhRjNUlhCtfACXo0BhTZH9CckFzv2upN32N3FzK6
FmZD2kSNTWzh5HZi796H4PTauGadajyUkyozU7caDvw8HevKXNxAALEiPM28MTyFHdwmh4QB9qYO
knDDrqHxhxB/5KeOWpBFxlCweEBIC6lmaz5yuF2jKsTFG83yljt0H8FZVg9sGXirr+59QSgXHQQT
yTXk4apBO4AabQ0izxVLEGVvIhAN8UebH9XAkHEDLzAMtKbChJ+ig6AU6+ArBb8UMc2ETiIsZgg0
Pm5gZP6+fOsYYmoVIkIbW0bRfeNBhC0gAufFoSH8Wj/LftFSogYX677Tk3/xNn6TzoeliyDamVTx
K5y4yur2kKG8VLNOfWLohhxE9KkxKJA63xG9ArtwIqrgalHk0sJxtsGUw+vxcXFicwNyhfT4IL7V
wq5+RnOfl8dvCYnsvUi/uf15lX5sWmRF82XbmTKzZeOI8Xuqqv3UqCzbBclRhQkQcSJggmJMPovF
x7hl164H9rVooExrdCsZz6uax82o8bLGwE4FAlYuv6l3E0nN/IGhYoTRDYIly3COyCDfej25NPlT
Q9fLMl9soJJ5X+rRT1Y3MwPRt4abn42VCcLy5bQLFOc5odb4CpLU5dD3NgkDq6kAYh5yJWKhTyp9
ekNz9Djw9EJM23qpPhcKuW+Uz1xex+vXRMgXmjehhtPF6l9zBwzMxfuW7RuHORMZFGIcRTOR3n3R
598F5Qu4L/L3SH7igt2k6ApiCiFafKdRcFHIJ1GAHqgUaFl6K/GwzHdJ8tY51aeNzzEocQqp8N7H
h8W3wt1n36dMJcFjeMuEnDiq8VFapIz6zrHfJxoGj5kgO2HSAHbLuC5Rdj4CaeMM72/xwDg/MZBJ
kzJ0+RmsWNyX8K/iM10GfkU6eiDe8zwC7RLMicgsAajen/dVTA1XsnWJ0p0Z5f9hOr8cP9Ool85v
vUf8c8yenW4454B+nOT1HU+YkxRRcZVP9pFqUJFE+ArXMraQHSndQDx7TEFkUOiDQ3cfXcVebduU
nbHoOgP/yO4j/aYh/xcrS4NFlHLHcW0M/nAapYBccPbmfhf8dVQyAcHmHodQZS5+pSOEsGMHywW6
g0Gxfizfe4FMsqEhRQRCH4N7MssWUJg/hK9SKwVMVSr2M3xNE/ixOECw+n1deof0gJg6hWdXBPcd
nMNt3VSz7uXqTAb/9azAsYaZJjup0ua3sIQDXTN8xBiXd+VYKgKFoO1JdzmXHehJ7mpTAN8wi/3x
D7cBZu7ok51EAgKMkKosgUw75TRNY2+Vs32zh3Mdf1FRraIas1EtHqsf1zcaKn6UEA7XwOVqbA5w
JuBK7oiMf3QSJkdpBdl9Lt5d/lf/rOhaXdM94fC1dV4SbjfIhC12QeTRP5EnzFaZTcwkzZ65djK0
NZp628uOQY46ThQMoH/6RrC2TeRxQ6h2h50VrAiJhTExvOwsuh9izVkaU6vpRTZeBgVjjq34Govp
J2PJl32Q+slq0P7QtqkWBiiLvv/gnUi+yXst5OHzilusLTkhTpbIPYV2Y6LJpTjHDXpXfPsJpXDH
CpCr67UfTdscrH8xyCG/Ncmt++R8tL8NltkLW1udMz84R3jwrliDtTA/xvDry31CmVAP8Dl53gH+
FtzjDjr45M6KpfX7o4YtJIsCsS2MsOlcVSitj3onzQn4Ih/FkieQ8VOlguUqUQrMUNWS7azMt+Nf
2pxAcGcxKjZqAE0QEWdkhvMy7kynMTWu+x6+Sf1j1cojHNL6ATanoswUI5+lNV0RaAjWXnlKLFyj
vTc1KsPLM3LKmoenouY61Vz9+vp4BkEvCS1l54j3dV0XDh69mexVmNZ/WGgLsPBz69jolzQWOaN8
SLETVPX7NUXo11SMlvcohDMjrvB/99Hr/nKPgKAY7o5+OVyj1G4djLdPl1XDIZrNA9+VLwiPXQkb
j3EdwLXPQbx6SG3skwLvwcerFf28TY26PaJGd4yzapdY8EvZ5rCzjDK3TKCQ3Vb1BLs0FeNKO4HE
Dnh6ZTx6htLBh4FV7j4nnCyu768wwU6vbwLUvI2fuWo0sDGgkVr9pVF/Oq3b3GbfBb2c0eQ1VV14
YJPx0Zj5vf8LM8LUZy3DhAuyTMKel3LjFqHvxM0J+VyFVVfx1xL62bbPD8d+Yi0bjcHqml3zhW5t
GAJu8Jodxmjcdw1PqdZNZ2GYE5gIjLP4VEMj4099rNTT9bO7V9Ggm7NtsNxdX6k0GMYN837ZzGbe
G2FeWRgMfIrK+1deFdURGvKE91YDXTJsJ8h/MNvrIw7tcXE6E0RFAODm25+IcKpTPDNwP0csn4Tc
aFJtfdrHgPs3SHTAZJ02voq5Omg0BxPYHWJrhiatizW4JtneOBr8vC6MpkrZ8gy/IEIIriA7ZN/a
mjGNAw/0aaYOiWdFcF5cpkNbZ8xMKraCLZfBnKYufQrOCLMvStZpoKWJYcU7QCiNMwr1xpJUpH/X
ikw5ce50Yzl4Dgj2bN8212IVU5JM7co6OnpiFAkynX/hobSjNoK6HPyWqTxXHVVIGvmzZygxNqut
fgXVcOuMUnPZinlU6uV67qK7gZTKe6IqqQZ197hRmKta5Np45jITCwft8Jz4/xzdPYxMxBUwy6of
uJqpI2/GoCGThl4OSY4QlJvFUyztRwuV/iQSIcLyc+oujDxN0ZzEOA4MS6shJCxpUT4IDRrqkLYc
6k53J8ekxJhwVLT6pvAErhStrvq7k4DjgLlAoRk8ZpTZ4vs5tbWqqflT0XNS9i+npg1ASpoJX8S9
lw0ZqVjwsmY9B7zBoCFVhUR5qCM1Lia0TEyd55Cj68hXzBjKwdbItbYuc/TEoUXKFCvT40QML5K9
dZ2Hqln4j9wIadQ2/1SnCHF8DAO9PmZl7870ei1RUEXk0ZK0+L7l/GOUHn7SUVKCyg8kzl7S8whu
31TxZ9dp5PG28CkOAB6Pjc4V4gdSDkoUcj7y8vTNLZOUQil64sg1fLdrYfZzLDmFN16fXsab7pbK
DP3WwTMeCIv5DQS7YseXwRPejn+mdeRqy8Sp60rix+luNwYyBn4DdiPxbwPLZKBnQlVqlDpUoS7i
2/1S4JNMX4ODYdvQX/dxCWDOMCA8k0oWDdqV3aCJelOa12mDbAvZu42aW6CXZzsJxhxFN1fwRdjl
nCW22P3cCCKjY8PB12cj/mnR1pkzbwg/hZuvx9E8QVFr2bKM9sdim3qYXDVyjJP6pa4YvVJZZCu8
TzFZb+5v95rk+FMAGPuE/gqdAE4NqyhEQhCUVPwbglHsMWYRRTYdazNszasy0e9WZH+/u3Fuetun
hHaDjFDr3q/VC8JHlpeUfkpGF5CVtWdXLfR0E9lLY6tc4uIxjmMBXbrYsJEUeBko6JLRRtBy3Fc7
kNWCiZHz0OR+TEpUhTJWq8XLC30OhBNF53YMdT8P5Wu/jg+jvl1rMbyRPeI7aYw48r0uCVjXvaGK
u1vY5AWOzhbJpa9AYhRp6SfoS40YgnGHikw6EUm2ehGsQ0DCrXn2dhfK/pGFYhTMxkVE6QFxMWGC
2UtMnZI+dU9yLOQKbYX3lhtx2fr8Hrt2+sWBL0n3bz7OdfoGoWMOiaUQ/xBIdSNDch8ZhXBxVTiK
dRayXRGQy+OBCm9d4mpNN/DdCxKDnMwkesKRNeSkDEdC16P1GxVeYt/h/l791TgEnFU96vYNFH3i
wguvBoO919ExufNDQo/GfMwkQDPV3cKfrqsOXn62KUMSiqLp3InsB83FiTkWXtkPSqhfh0DgSR3n
jTypAhI6cWYy8OiIm6Zdvb4ZAeVLB2K91gJWWv8Qhk6Wltl/T5d+NRPVPpz/35S/xrUW5oXVX2Nh
KT+wL6JHey6oo5usy+mjoXo+cSNCWzoEwqoRPPigGvs7P62aRw4bRz82NVBkJlz7/Y6n1kA8hFKJ
blB5WW1eEi0k2r07cCyq2blZ1jdzJR4Y1azD0HqJt5TpmSz96ccl4QwsJL4fdN/IiMzE5HjwmlqM
sB5pLwsZibFrNX0iKvmOZBTyfdY8rwZw3gmbaKhsWhIuptz5XJV3V9gSeK4/m7pKK+I0HahEeGdd
pzRPobZqWq5GnhEtTYCL4ThTw4lYJoN7KzUf/yc0KaFs9o3cI2g4js1EK212PNpCgBcj/B5c+ytp
Y3k37/h6WpjJg5FWv+1sDZnW9YLi5mKeIvabs0ewAw//rX4y4mXrN3ljUmzvf3F5s9RgBEnB/ALx
phasbSRUQJoaLqGteE4mdnA7h0rhugizV7hs8zWHTRKsJID1vFAomfLwfDiGdgYl/f/2i9O8JUnJ
De0OMZ3lokK32UxTlJzbpLgqCkfORVxDrw3dZ5pBssnwucG4ubWxPTZ8OJ5UFN/v2BMsy2ks/i0d
Q/ld1itSxK1q71gKAilBYLra+RO6+OAjx4D/1Gp6EWbqGLS4Ek8Q4DFRSOgKLgJVsQWoicfaHjM7
bE4cCoceZKF/HIKZ2voIlxZWJTCXuT2d6PwphBUdsceI5IqB6Oe2JpuGoGQBOJqlPW1V/GQ2ubfB
dd26lhxAMa/Y+cGezUsg8zo22szSyXt+12XmvD3V3LgaPtKq6/+eloU6h9f8JGa81m8IbyjWVgIM
kRhohGUSYR+WNM8E78qPIhqr0W1FkidAHRfEEVO7QE9kvLOCFhXUtvZQvw3LDp9lUmEX2dwepaGx
WbiQYs8m9YmOjpIgHIaSuuTxCFBWmykpfD0dSVaXIIfNy4IRIcmsTfIIVGqC/FJiy5aQtd7AePHo
HZAhbYSgWkQ01jaPz3W0sN2SelQ3nXM0AhGUhVQj8dLN01d0g2qvQ2p37J+wsIGupRrePIau9lTp
aNWt59Uo5OhrInyT+CGgxAzftAhQTkbs9KVmvCZrefqtIMTW4sK7yjWsF9VpW+51sPBligPCEj5U
S0L/yjj8A47XzLzzuqUJdvHSxQRsnbNVxKoRqeEPUFfxJpmsSiuVqx8lmx/czO75yKykkR2+Lc4N
j9O0CFA1AT8aUHZMzeecieZntNhmmdpZpjeP6d4lMO69SisialPy4oQsPFy1LOJdjfy18xdcBJaB
nbdim35NE4U4g9Jj4/D/ibm/jw4qHmiWQiGGmLHUi+Fykq0z5a8WgvA+HViFSZIiiBNIbjSdQwlR
ifXXZD9PIYmFAZrAANmy28h7vfF/Es2uZ1XBjdMg/ZbfXpkIbvN1xn4BVpIJstvQq5pcQP0pJRyR
/DIDEXmJ0nAguZqBq83TpLqFcLltqrdhCgwYOy1M0cECC+zgn0J/C8gNO6j5FMm9U9tESei1Amoy
FFjJn72wlCkSFYxpzoNDUvEeuLk5tRGDk6hde5fdPhN1gMX2GB3YAceslOyMWxsbBaOpObCrGj9S
dSPmyCpQHLH2VSgsOR7FytVT6Gb4N4WglYj5MmLGOKYeG1rsBab+TomCYUvKiZYXBGqDekVIwlLE
FX4NVxcI66sGpGHTy8IgFfiJhVzwwBIoByLhvjtFKT+HsHNzd9WCZwrZk00edcap/NXzSdiPGREt
tcAAIFNgZekal+arqQHOBdrXkug43Ejl6ENSmlisfp36w7HnY/PPZlgG7DZGlD5JteAf62JeRf7g
mNp3AMDdFD+stA8JjyHttQ0Sp/3FdIeD1oBuYCQa1t5B0PZTCtYPil+l1agkHIodSKJPP5KYsihb
fr02IfjeWIvpl9IJSwPhtEE3QrxBmytHBoFr1xxRxEXasRgZ1RybWHZh1Uyq4JE1PQ8iy0gEoHqZ
BnJe6zN8xC35s7+VXdQX82J3b9UHVcN9HMBqF1wM2AmLQ67d4TYSIdrQSeu6BFRt/NjqdGXUWdcV
byaHAQomNahQ+RGYxyy0C7n2EPkYHX324/6fQUb3Xn9ia+5/lk7ruzGXa8E2oCN8O7tCEhvyZ3Al
FBoK+KgEpAvNnoWwp3IrgOLiIQGKpCPZ5p6Cn4uyH0WkywqWIfXa3IKKMBnBq8prklPljrzTWeR6
IJQ3jXsJpKjU7yrEGwRRThqJH1HD3A25dcuiFzWb9gMFq89GcvEonDaq/lgZg5wFdQCfIxyAsNbd
+iO/h9rACZ2GCvnIWbQU8zeF8icJWSG8pef9amOMgaiiyxRxkBNcSjsIGRQjjsWW8t3JObHD0gMo
AOHafoqCqGxjMGF5LSJHEohYge//I39Z59vidVEa/XxevAvtLPapdNOWgQ0CzjInXwZwSPqEoQ2e
/ZNDT5c5iQh8KFCNiSip6ZpmXh5PJh/sEfGiCYPTbN4bUwWAWBOM31LcfLdaUJvI4/3Hc/Ey9edP
p7fHEaVF4aZnCun4V3QMKCI2Kvg8HofCoxNaPePH6Je236TAtwFv+RYZzvaFnCqF0jVRjBba0Yfg
7xyGaIzMUikFwdQ2BUWxfjZZ/BL801CtXoL0+4rayUx2oYmXu4WATguQ6zopE0l7UDMaQIREbzFd
PaHHO5spveiJOFppS3L4Gglvf4nyQ/cxEyrSFfZNLkwp2Bh7oNN8qMehNmjB+XwOSB6p18CSLPtU
j70cZebkbaLwySBGqOzjV9vjZgqiQLsq3yBScKv8Sr/mEY55+yj4LIE/VnynudPh8cBE9fPUs8p1
e+s2Bn6jDIrzJo5B411kPscZBSQS3viGSc6SzGRf1kyb4rKDEia0Mq9gzemNO5NpPNSgqiQBL73F
kcS4tZ4yQ8YiPUbqdP1nN2O5xaQQEj3nrUbJspFg9HnAz1VTmhDks5ZHnchM66bSQ+4/krTgpTsG
iCffZAGYVSenR/T6sYHKZU0E7CDZiqVPZeC1aqlTC1SI3u5uTi16gB9VisVowc63GsTRp6GHsK8q
vf104R4g3/zOZbfP+4b84R1dkyLcbNI3HoKGoCxh2ljXE+o2kGrRpJteZ8uNlI6VZDTZyxhSVlE1
x45xl0TLPN/ABr9tozj7If1TFBXOCKarTwZZeVr7pOBygbIrxTw4imHkNqNt+dGrDVptuUErIbR5
V1HCdYz6SGtcOOqTkwAONvof6Xk5NXKomB2ssjsLQ9F9GigfRXqSsGqOX8NQuW3wzYjs8ma5DRrp
fJ8voq5wl6kWRu8z93rWM8XldIRNxl1zBIbEETAGO4v91ZD0plfiw2fbYKeVa7EimXyvphSOqAWj
pHdooz3hil4SCSH/9juxt06KCkIAmZ32JpX6v9bs7/ns0VU8jmlLiqbtxr+DDJ0MEAur/TPHVXUo
KIOxhbdIu+GMxUCaRpRlbC9LLkSjLGItvYCTwXpEnaJRrP52c58boY3cyHWDUEm1j6zXyZrl3YZf
fIQr3oGsg67T1V0RzJh68h3rNZP0qIlqGFNXMTjsN2zunviR7LS6otO9Zmc+uWEfNMg6ZpFxfn0t
MV0EkXzBKre8/ohLvr5w9cPUYAaWLDE9pazOmMIGSjqGmHRNoqrF2cCimPRtqsaAcqbYY4wnVB9K
80GAa1oBtxt5otBoMjTXHMUXeJfYRgt39fCV9xFm7DWiaWy3ZHs6HPwuqgJlFvXNCKnHDVyDxGIb
7g7qgjHNriVARQTKz4P6gIafcaZEPVvH7nLzVj5S58vyIExXRy3QKII+hwIfHUFyyOZjkaj0l0Oj
wtowFrRtZuyizuAXx5cfgGx1OhVXKvgWho5xqTBRMqhU2X5ClP0qGcW2rSODNnqFXE6ZYnVjeA/y
ghYjdEaAjBcvkZkrw050Z/A2xGiLSWDiduwMpj7D+gvrdiTGOQX5m4hZ55l/ccP+0Jx6sS3xPMzs
PpmHZmAjOsIZKLehFFZ0bLCFEBe+ty8uHxu4tPa+fUpBPNKlZIFiOEwssOca5QqnWSwVPU4fUUDt
38mmOc3kwQKnwtJGSq1/Jtv3hZuTvimrbtMkW8l/KKDgi3rgyJ+6NwE0z+2dj9fjOe4h2GqAL44N
2QbONGIURlBIQ2OeqkMDsbSlnBBFJIr5GrLFDOD5S+6Sv1S/I3x62z5nG4YLcmbb9HtI2fvdeD9m
HA1e9364sxxr98IM98LJbcAKOlnvzpe4VbMjOihcP/0zzsPvpveDmorsKSURx2Lb9SHI8FbjbaPF
2T3Lu44YEnHbjRZzB13RkhzMGTTCOvGWHXQTmjI3Jvuvprq56T/ExcE1Pq2gPy77QfWU+LNtMbTN
iMV6AWO+h8Uq7BlsLYvbyRGmPLnRSrHA94r6ep6gQtL3WzrC5EfVQ74mIlqBvQ+fLkzxX6tKK+rp
XrMhNwJgXtOx+NS1leQsCj3j+TBDJsLA7QRHh+UAb48R8jPjl5KqOpixIboAhDlRYF5yDlqBQUYw
FNa4ucUvLz/mjDvDwDKsq+YN9etJuXfkZdAFcTeouMeAk7SbwGxMK0nKES/Ctdqqpd1ys23kzEdB
ktvzgxzt06qhmo9WaV+zaZka2/cUHaC5SViMW3V9bfyfWgC7lzjNOA+Cdq5+V6nidxGN9WVqgMCX
3vpj81r7ZPhCtpNab0Kz9/bU/nFD523BicjfoBBRuoxlo91E6U1T3nEk8XGwn8iALPGJo4GNcmak
pn1AbIas+REpRyxddrJ2MUNNrTn9RpLSMwTCc9dmM50sWaE3q0vHwip+wD5qpNw9+oxl2Ym1PHXh
yaIU5HoVVqi8ULmQBkILnHA9KACcym4dcEc+FT8EfbGz5HZocFEufY0I89CcpOPWqczuktcYDJqL
4GC33QXPw+xW+DUS2XRhC9C2OmG5wTClqcHjKBqD5Tyq1hsqYNJIbsGvjE7NOTv73EFTk71bnq4J
TWt+K4v7bIQT+UZPHiUpBipG7pdjo6cKArFI6Mk6E+LSeRLzgUi2IEw/u2YEaqVwwANjzEgfeh1k
dYIf01XSBjpA/WZ6cLJO8KDJGtLpOv/Oyu5/iRUpk1j3Ya4SIBF2IpWgipKjSG0h3eZHO1q5QspZ
ZC/WbbOE1QEIxePXJagWvOc/9eqFVwM4RqcbZBsHRaSAS0W88wYBWgHxAhhkuJCsvxYK9v1ppQyU
FBSdg/g6JLTRsty0IQfrRkTSbGqDxrvHeSjk5xQ7DosuuwckfU/ACN1pmwhyVH+Hk+9tr2uPBrp9
U8XjyWhQRZRgb3fqcO88ZTh3GmQdR/JvWgFyPWKQBDigBTswm/nrEWpS85otjaju4RQxQStIsATU
/YTvMFntsPtdJlKR4ihsCoEv+hELngDlZR4WhjtcKhzpffulEeo8UjgdBSbg2k7AAGy12Qx0Nc0l
N1kSP01k/65drYlvM/uE4JqJ6EiAVT8axwgsxhHLs6gE3W0hKKYpFhHEI+x5pbJa5/oHpptSz3Xi
hsnBuYaJIA9ZmL0skmd+IyzHTZxu0dQMwv8ZN3ptMRyEZiEQp+H5COkrUj8IvobELJxZOvuIRXbW
8FGyMlt9lj213OuzTljK8qclYMFtGYwW7234vWxVf+murZX3JlXBJIbMzi8Ro6zayW5ibamWf5F9
TbVRVtcIvFXbo+LiJ5hxpdu1Zy7DX4IV6pbYwkUlboTGEU1iepOzQAj0SbREI8c9gLbMt1aq2U4N
W/DIrdKjoT3rwhqNFctUULAfEdKSOHf0TGVr4mbMMxtMebnyQsI6KtjAlfknaeQTspEbyzhgltLR
55qYPNOtNs9p8+450ksMhoU2vrJuiNV9eoW6eT5Oky/6Pmekqn4TkvVtRaNb0oaHXK7gwKi4AJ7X
RWu8gctAqnJ1/K5Rg+eobRGsD2o7iEc2UW1URq2pLp+/oHwiptKItnOwwy7hxcExI+xeaz2kjb3p
PMAjtkbr1EvD1ygCtTh2OWhDCmXfbb1t4ibCNsF1+nKqxkcPtVrKRl9SfHAhDmCRycBKJWSqiviQ
OplIdMCn5ChP0WvfoBKIaWfEkZuXvGxeOyzprrVSnosbzKBKV6rUuGdlGClmWWkSkLLiWTGCRZtN
e4KtZNq53fB0YHdoBOA7W5lzK+3HORJlfnPIvji3cUgu7d7xDCyvmx52ChClmw720SmTFlsxiF6k
zFzvlKn+utBy5VTBVX5/48e8Rx2RI0MwSWOsgKoZWRoPNTEf8vjANH5MDbTUAAkGe7nOv0PIm8Tr
mkJTYjo4CJSTitf6ltVsRaf3+p8iqXq29kwf/wU4rFNTDNyS119i02+dLxvr241FB9pct0pF/eC1
Vfit4BsQHY35xXVcJGnKUOyTc9Vt6t9fy1TbECgH4K3p13mWpw2WokypV5A8qhwuuNFKBs5pmJXx
crbqRXYrFiNfkk9tCiCdHvCzrynH5msrKJo09+DxFDX9vTyeJGMIkbFffEopPe9jsItfN9F593Dp
svv8Mn/nXuHM+diYGbw/uGgsp+sH/4B+d08N9ATTAtYREJvW62tbwx9Uoeu/hqvjz5y1tZg+9kLa
MD0ueCYo89DgI9jPNQx5OTXMPGvgBt1JFktJuxn1dpugqtGDVdpJaHEqtQS8V8ZsvkzIisCBWeIg
TVUtNEbgBI1OM9HLWDjlkwyk30iCN/ewIKu3NPpsjSvlxQ9fcNcAE8y/lSU6Q9kTkNViu4J7/kkm
sdXidRR3LFbZmu2wgsT8dLRkC2YtmKA5ZtNxa1q4Xv2za5KJbgJ7yQbxFteEXjMQrz4ta6wKewTC
TidOxfFFKmSG8Fi9qTQkbXcmbME1nkUYUfuOlwQCk8hMxYScbVJLv3QFpVuLfCpkdIHDNXuuVDeC
aTlNvO6vtC7pwUW0isdB2YN2D1yL/FR74CX/isfueKSu2aml0/Fox3OlBFbxiGZZBON1KGbZW2z4
DOhmAjYkiwkViY7voLbeNtSj3CGVT3h1NBDyHTx63yOjIx5WbVeIlP/48bJa5iXWBjPYGz7WDN/Y
GGqVGNLz72GXAxpmR0blF4+Mxso7Va2FElgI8UPX9Cs0BCTKxWecBKm6JDTYrXWlc0Qi3IfE4sp+
YLinfAQrO0lx1ofL2YLSbfIYe5DAJD+XADehiKotdHVp2tjFrvcdBsz1assBTbxHOLM+EbNlyI6P
td9iv/lwT+bpAWDqq27bnl6SvWVEAvIW5RhTygbgS4Wb38Biib4WR0c94LFGmtidP7+aDkjqFU9v
etPmDtTsIRhV3sFNlqJbVnJ+yg7wPIxIpJCww1rP+Zsh5TgUdrl1Mi6OFak2OpJvpS9oabQ/GPVF
KSVO+g/ZUGdVziFpBuDcHdQJzAPbF+4kvRXxZqiXC6z9qN0IT/W6Z47L+JfNtHyCGND4M9DP0u70
O6tPD7J+cX+Li1q+cFgnHVCoquW6aidFNPNSxu8QLNdvpXADhs9bxsqGTOGHWPaR8ejf3LpW3Wgb
Iki7NszG/7TwlUW0cm+No/MqkN5P8c0XE1eC5KGDKonPMNMQIH73mO7naTPfySpCl805BS3yVQPw
nuIVF60zHPXnZCxPIYBA2VTOE9LdQswr09uXyt0epEJhp46PrcjWlO0md6GLOjjyu60glNkdzB1c
F0QGkSdHoCojdJJ9ZvyhUS1IvmvlxndOe5IMBlhwlnz0aK1RC6QBfU+K/a5PjrbXSp+XSmOIEyOG
TwQTEJ+SPiJlyuAo7cTWWyp1KX9ATxYP2yjL4+rwNia1v9JHsG3NAXkwkLr9Mlmx/K8mR85ewIe8
IwPfHBRY5pQuayeQrGztC9JtZC+sRyie3gc7uSAmvH3nFjSJ5luYmFs7ScRyLeCIdfCW1Y7utMbr
RThlb1GtE30/o9Oijv4psVVm4Q3elFrI4zoyRG3MsxSiF0FGdt9Gmy8U85soTYYdTTZ/8ACwDSmw
+RAjZfa8FLsVf3f9ja6ptA6JztvyQuI64ppCYXx4k5VXPbUyNgr+kQgIohdG5Rg/wymlki0xpCq/
6TP2eiZ9g0vwakzFKtIelCBB4fmNLcNh9zK7b1iWBKmnQSQJATEpi820vj+i79pKt6Z5sSvO3koQ
J+snSTjr52k6cLsimtzDfua8EN0mAzW4AiRc4tAeOzI0H7La4yeXhuXIds1AbG2VodzVVKT+Gp3G
Oj1TB8C7awTEDalQoyPHcYrAU8zUdwQc4qP8DFHthrSVye9QIqKjEuzF+NiMv4QOthBgi3KWQ/Yy
Qe5Trq2nXVKjo9gL1CPEG5YX3dOjsKoRWEPxq55z1I1VzmBlIG46G9/+LsK+OnFBvbK42u/v7plc
muOGZMKoI33FT7wM1wPSNwjVAbP/iP6LHIDQFReaiYtUwbGKg2g/tn1PjTeBrEj31sy8xexLrD/W
fWnTP7j5jPZ2ckY4gjIGGD95hp9MNm2jzW7nTAcUkxl1M1F0fK6XGOfTi7BG7KGHF3qVVBAAfYrb
vN8SBPV00e9ikgz+ploVSUgafKvr7uwMoIjM5RAYSAXbrqkPLtOU5A1qVgxXgAncct+t4+TB30BV
KJpdNOPEaKZd//xSD7GwIuH/WgTsFrdDCZCEEjHtJlHvTK4DRaQOE122/emilaaqMEBBXRfMExi5
7puw2geoe9d0cMnJAcW1bkhZvD5zu89iUkTJcTYr656ZlCYhQ7iFBePx4JYMPty4m+eXPmZYj/Mp
673NsJWAyGRgo184coRX1N7MpA9dDIber1HsrCINC8pCDXnslscP4xrM3LGgxVlda2A0CYTWeSpv
gKmCHF1YtwJaZul12uaq0O26kapp5eq4UiAalNy7rR/lNescVJzj97ikGp62h8PWgw4lqAx+FomQ
w5QKMFyMP+5VeKxOPWcwcXlvejiIdV6ADPBMooIrE0r97XquR5tVvXmoQKGVDPOL9MPNU/QPRONC
Tx8qO7UZCvWb33LZstPsRHuIQhAsCFU9Tp7K0MQYuYcCnMxSOuiWdj3VgwuaBALcYo6qVGlXcTuH
41ZuZxFoKOMwH3TgrmCPHSZbrzRApTxTTCsKct099yqEHFupIR/49/3dyC4LCnMgb76LY1axExxQ
o9BmCuH3x5T74Z6Q+lpktf5q5QhWVigxYTOwKn2p5xWPcu575X52TWSY7S6lA7fqg/Gg0JoYRk49
V5MIRou5iIVg5nFyAEPmBysAhqjyB3oJCVKG8TdGWmmJpzH+tdwS7UB5GBPlawp6vt4wYeZ1o0tI
yrtmECtrt6wHC5oxuVcJ4PAl8B1ATSrNtKNqyTdPWBkPSWcsBoOP5evTNNT1hzOVGPfIQn3MNj2a
TyriJZ4kTE4CVa46fudvymSPDviGgA1khggP/W4bLtYTMYRUe3gklEzLM2qgxE0vP4ezfStnr4zz
pFfrR1q2v2dqQ3mumlwko1biDNmkqotUeuPUP7H+C+JhMi42WVmM9VpuCiF/5h4L84qHqHksqA1c
LZh2yAxcGLX5y2lXvlFaq44nT3SujGBVxIsAMdKaLDANYj9SXaYK62PF47ZzkxFclkrhP/oCvwyd
aJ319SdizEfKQI0pnRoOQ5iNF3bGF1uxv3penEhvawrQuJxmQaMIG+rk5f0dgudLUkuwk9nV2qla
p7OH0kRrVZm62ssLOfquhssCv9u9yHqIGTLdo71Lq7IKvLkDKgN9vrioMpJizTvPmvvr13RyM1y/
IBVSrJZMBq9D83ExgmMMmtV1dPS8wj8bQVCeKnRcJPH16nkETc3dcVd4k+9HIg1xL/QNZU5fzfbx
KeU2eEftsl+yG05+q2X+e4V8jjt+6S4EMJ4Z2jiGb/sSkA05nWZMsmVFAfTrXpdweTYqE6IYgDZW
TH3zGP2u/pq19OiqO7K8//9wrpaFHskAXM3xbk6CBKMDBYCLnee9Wd7//6R2LGeS2xSUDjZ+LNw8
Gc9GH0lgOsN3Rj3445+6jy9OpG27Dn5pwnctg43+6WrrT6tqU10cTCmpmAS9NHmR1pxJINexjdBk
ivBLUdmtnDOpNbGFPKdZaGnSDzu/iQeeKixdw1Z3+b8pMKrQDlJ87x943dGWDEY6rFoGV/BLomCO
0OzXpUHCy/763hKlwkvPibQg46+vv+Ug3/UKnhpLF+Qr7VHu1ETwahbvoEsXyIcI2uO4c1nS22+/
fDLrhmSalFdQcYxSfcYt0Uh6hQMkI8Nc7n5DEQwDbB54GF1ESDMrMOS9S4ve1uAAxN8xgFZJjvWK
zft5YKj0QTa446SacC82EUFU0Rr3PMzes1UyyeCrA27z3nEvw3tqXGJ0/n4VLr2UbO5X1cknGAgT
Icoz8weJtvuSWdW9o0wDIX3zNryE5IloqEE6fCOBSLUPrNg0TNe6Y93HDP9rdfTK2J+fshLO6BTr
rgE1Lr5axbvbzOu1BMpC6Kb+IzxmupCkBZ1DodYFkhA4uUaea0leGyOPxjCbeeD26OT25sZSDbDS
YkzY7yjXXETpMM3yl96Fmb57102a8poR/7ieiTQAI+tlYNKsrYFfaRyQ13MPNxcRLiKj7DpsIYPj
K1ApNyG4h6rprlBHsEejey+Kkz0OXHmhcIQv0JQsRQWdqaiJvKTP+zOPl0dq7BjWjTOJOOQ4eOZK
rjFSqsOTKKqfHCjqrYNTucBhcjS5aS1D8EWVOpdpJPpLF0Iz0Qm54C2NYcLWdTBTbGyH+btYan5i
mlK05CeiS4TQEv+U1Je/+Nkcita0F4DDSQszKYpGWGRuOeG1S6oEroChYCBuUo1ZCCFup/Bn2sdL
TfaYYxX0D+DETJZ/9VfxIgRbWTWVZYmsDthiOkUplylGaJInzdaZ0Wc3H6d0hCzQFdnlATzDAvgR
qIfmreMCgZNHTXCQJ+8L9R5QjKyM0fghQE3k5AL7MWlAN1MhhNNSYXCez3JS2ag3qmJw0tW9b+7U
DNR9KCtMOeSpkGJRKLvaHgiZrlLAiSXDLlgQs8VZrCkzVenKN3ET9qnARXsd/fiYD7NMs944Nax6
xzaMkqBNeF1Tle/WrW/cT/HVWiDfqHKlvineDtpSehGQuBo6+cpQBD0c6M2lfDv6cH/iT10kZKR+
udnUJ+eUWReOq/cu/q5NfwA5BZN+PMHSESmNnGgwyh+NUa3/j+vFS/VlS+REcSC8x47TfCZ4P1O8
XZC89QAazlZR52mz+LbT7CzDqniYZajlB403tKI5OCaDE9xUiwUm0+qRFPAsTK1Py9hdbZ1M8jtu
+GWk+A4tO/yILrdIiU05+0iFdQP6+gv/HIda1n/POtdJ3WkEMepHr0mbA/hDfXtxAZ5nJIxAMYgO
aDN+Es8LZxVVXm4GGM5Y0JUyV+P5bxvYHDloa6CDAj6uE4kHaVUFETLd/DFAhi2bcmqHiFqvJF8O
mu6QbggYNjp3QQG+KOC75erMLLo9mskcKf3h1doy2WPz6raCITpkO+KqR55MDhBVFVWik3mkt3cz
5liCQWD3/l8q+AZEZ5PKk6A6VEAxNd4tMyoLPgPvCMwbkfSyXuvMoMkK4u6xF+tdVuL27Jl1vS9P
3uuPiYJK4FDhacKQsAwVqOu5KZ7s9sng91gluJYxp5k/hdIneFwTi/3VjfPuA7kyrnKlFWLS+oCm
Uhqz0z2LFqypIJ+gDRSFyLK0b444JvkgWVmUjQJ4RmwRI7IaCaVyYWyAgFhNnClA/mE8EzXWvmR+
jiK8zBD1iq6+mA5K0/f6rp9cMdDoDDiKrU8DvhxotGjyAQGjDEd3F0U2QsQFz6nskLl/AMNkWAO+
PYbnP4Z/T7wLSgBqvi8AYWS62RqTyI2z9WavP5Q4A16uWyAjWeEObuD+C6Ta82gPsrZmJQIDtXMs
dwzuBSlpnrdImrl8HPXRi+tPgo6BxrveDIg7MdzyIqzC96zvjZKJEURmZb38tFTJalbKVebsyk5Y
XEMdVYwBKyODFGZY7HWVCC54K59gHTzm1q7EJvirdiFjn6MPo/1QBcEpHGQ3IvdpmFiKn02gvTKt
Fcg1FQKLkR8UPcM13e7xs1PrF4DEbkO/LKdnmKzDQUyqi0HFO68vS+IZVhHxv1cC0wcvticz5Wp0
FRRK633a9+FILxKO954I7q/wp84FMQfyGgxD4doVYErT94OWacmxN+pnWCoNEuaTODCNba/mKJk8
q5zhCAemU4yxzjt+Oo95A2Mri6WPnn/TNZJTEnklIwCqVfNT49ugkWtwPUgodPj4iNF63pSBqyFZ
9hcfckCo4ojd/uVRZ38PuSESJ+Wbu5lWHV0nM0EQ4O/RNT5xbvfJrTFPXZ45Re7Yx81gA+IM4GbY
eTF5G7RrtSMeqF2aEd/Tt1oIGeQ9KpjJZPo1B5/Dw93S8Yr94Z9Erdn+QxxX2gLgF536Qu+bq/nO
28ydBQPLSGaFAVoF5R4SVpjhGqoV/e1QGZLJXc/TY6gESaOMn9gy1PjaXhymSPIJBLh2+kJfYzrC
VNYZsCHRkKt5WbTxCjMJoHbpfFJiSse83y6+6PCrGwTqgh2FgEYpcpMFyjXeWQEmco8sl9VJBHmL
wkErZx14pwINeddF3Q5MCbgYT+24mq+jOGGzev/fz30+ICipO72+JByegWzWB44abnXdHNdAOLrg
EawGsZUy3J80S+MDf9ystHXQiIMKOwZkdFLKui39H+p/KFSLIcEA2WjNDToZR6Ig/+Bbsij4AV/S
3FTlioJOkTczHKwluF8oG5l2cXj8JSie6ZZqDwuICFmG8pDeOu8FhVs03qm2h2D0YIOXmgsv5oKT
7R4VpR7sbQo8lu3Z4XKjsNI8zgvmgGjyRf5OCqxGlMt01bI6xyr8xZ/Y1cbSH7NUeroaanYoqcoH
SXaOeIS+/hZ+WB1CdgjN9j/EBWNkquXWBdTWKPeYBtcLDKcsuR57muiie1oFmSXw7mYlRucYfxd4
33RYavUTgeRyQXhnguhuDMpW3D5ioK9vpt1nTpfH8Ywi+ISBclskil53k10QTgh0wIFHZM/dyorZ
1559A6MEwE87HjoSB6uEO29sgeM6dFqBDma8lLDcJLmKpkR5+T6W5zcBqwXjZLqvWrTKGYydx+vY
z7Sp7td4PDBkPrpbP+/wWFDpqOSRPQcBEvNUYdnifg9gkNgciZg+uaw1nBNn4gGNLbDrGGNzGG9j
GDfF6N/XdFWijMSZu/Up0EoWhc8GL0RGQb+xjAyz/NCR8SqGaZNC6qLFlGaNn1hEZFh58oPNx4uo
4oolrPUuLixx26rUOeNEvVt+cXfTbw3l7JRhwqqmRkmdGT1EuDMjMDvyFRB18OhFXIuqUWGeUbku
USPTZPk/qvLyeVJfUOEH+zOqXbN7dCC0I3epH5RpoAzVbePMip40yUnvAINJyapFtx++rgWG1pzI
tzmKgoQS/71t6WWGjbeIcBi1+UgYAjRvrYuFLeV6DEilk0wXZbAUk6/eL3nd9QOaco47bHJw6f63
rb0Tu+O6EBcIA/DHuOiT35WZfIUfKVw1BB4iGHbBjAv2rgx/OW53tcfz9jUxJ1rjJUxCbo3ryhD3
ZNgEObdcFzh9xNqa96NLJ+B/+BDXgF1oLfcMc9PEVl1lnsmQX744lnQ9VbMEMRaahnY8MbM3IA0w
Fh2v/tGy6JTrBNiJdSLAE+GfSCIy3KB75pmy0LfKcXgE1jMIwFaic9r12msgQnnqKwhEDAOWDbJ7
M5NWV4x6dMBCvfiTjtzVZE1XzJL2iPqgmXo1NTrSkMsGUHln7ysVQadlOw0Ou6Rgrvay7WTmzZv7
i/tm8EU/6peoB9yi55HFJyF+Q0zrg8rmVYDwgv+m8mpijBblVBFUHdpGw3OQgdMNAuPPQf6/N2KL
gqpZ2H9OmkEjz/r/qqeXyv0EnYGTFtUsCXA2ERCy5vA4W+N/Lyze6qjIavurGECXJfe2e+SKcTVA
M+JrXt5yjpOyg9AqmFu2Cuhi4IOG41yhiKfJdsAou+Nz1EeToKE2fvfwOwdS5g307lVOIw8vtjCe
5uFzN0h0F+zIFPnBY9zs8U3U7mBJl/izrVEOSipZTW1/EN8Fgbqm47ZwQWpmtxk+6VmHnSMD5k3z
VcJ9MMrwZb2mqT4MxkGG42ld4vOknv3JLtu2tE0ACdre86RW7/WIGP+OAWMZs0Xti5Y8rL/ld2aq
mtwLyP3JIOGb7vAnYNvC1X6zEjxrLssKTPLEib3CwuHQUy9n/dAPI0nq0GQjJGT/iNpoSGNoUoZh
FZfnseFD7yB3trMEfcUDMIJB+l+sXqqq62GWkmQCrCzKiloMJbwWtdzYAwHcsYf0PDRD2aklYZBV
JnqfeWIWamwJyiFluFSj9UXpSEnd9/dSKNjcfC16kzCMG8PZsvvaLaGkZjCYJ5Eu+ATuB/ERf3N8
YfpxIDpMHuKbWNfjdvmyFKQ3bvErgZ97uHe3Myau7TpdesW6lwuDvlyl6ut0xCXxJv8OuUAK8Bhm
iz93IqOZbsYM+vGHlA7Zbn8soD8SUFcGf+VodzO2HLoM+zoezYYR5YxmkvHccpiDI/gwKigN8qOO
AY2QxuX5U48vggxs3ZgWYlQtbYrncxKYoC0JJpZYHS4MCwy9rNimjaiyyYg+MLebh7XIDrAHs6An
bj0VBsOOv907uzttHUhK8lvunx1Nisp0nmIccZDw8IRwONTHgrmAJpUnOgMbwEMXBH6aMf/WV5Qs
6o106Z4JDc0GFXzCNSK9sbRHCHFCCgoEo0G8FgDehSVpNFoRfxVdH2vKOttz5Cnpcu+f6FAMzZsr
O4MzvlIdmAa5eyn0NmQ+PjDjW7eiI0xciP3TBFu4rdEcWPX50hMhLpPYRM++Yw3oPAIqx4Pp1wW6
lb3ZBmyO0FF8KjBheUxwe7n3kt4+Cn5TuOU/CndXH8o8TmIu6aJ3ViPOk0QyFskgPhJj66xfqkop
rfBmDCtPXq+YEqAS0JczHs6b+Q+yU1Klxm5FmG98clwS7IbFOpjcLD/6tsWy4ufynJMsYq956HWQ
EDNpJfek2lxT3shxduFM1sDidbROxcOJbpFpcoLNVlYJmv8kNhdakjvpxMkPpAvbW2CNf7MZhy8X
sMAMHmxquU+5yxNlLUVs2lUFUHfJkYMNF0A++tjV2t3tmPDA5cu7M8YJ30/OXTRaYf5LVn0QQPDI
SZ/LCkHml6w5aqQCo9eyacYgNJw8gURIh18V+aDYqFBBOBX/Qg0nNVe+I3ZYN4H3p+M2DT2ySFtT
9fDyknJVLQjt4yt6oI0YmKkQ5alMa2acLu2KTx8SdhBHCz1oSFXWJKwBkvUTxwvZOacTM9R7O9p0
RCru5RLhP+F7tUrlHKTceP2DwIMaQ1pmgoiWknkW8Cty3Y4bGJXovzjqqwZpbyx69Q+47WQwhrm4
xFwtQbjZrxps/koLKvXnpGEaXE87p6Pchb9lpkRADtxMB869FFjWviBbaZAD83tPDYLm0woQnba0
6iK0N13XO+0ziEu5Ba9zEWuUQgR7iPqSaE4Y7oJSKu7voM1xRq4MVgKkuhDS8d8KfFStv08OFUpw
aJGY4YdlX9KsEW26qDYrjWEq+KHuODEV7BGzbLXph+C14lLusPZ/bbsLohZZJYECOZZ0jwI17Z6T
gwyuIqgqoCUe9xwd3F4RwZ7n5EAWpWcOhBdx6UG407eKHN1xgwn03gdyW/9suqLYcUT+GkV7owsW
d5nhg0Dg9jelDpBGzFQWZS01bVhIU5TC5Do4VlMnQasxkCuWqycjYUf3anLjSQMqla5DwFoEoSxG
IzZiz+bABAQ5Xq8hmsCrUYx/FydPenUg6TbjxxjkGFz1tiIDwniUt59jktlKu+i6Yw3vKCDGBwGO
RO7I3WgJbyburV53lPNb+God7GigBUonAaZ2r91ttJaOpEvzTtdE1uXWojdfQr6kxWBMkK1QE733
Cnlkg7O9pVk5bzBoaH0LgZi2tMFO3CwAHss5HuXsGkp85oeBHcccrKhoZ/Z6lpd5kgpekden4OKf
Q1E56mTmuBunwPLlE8jgqBliaVuZdHX/1iJfRQSJzDPDJ62QOBkDy4Q/FQqMYTXa+RAv4pPRzA21
ZejgOUoQ0tgNsruSiS96eOZZh+1mC2/9G6ILvdQ9ywtc2yZ3Onoj1ZinplE+hDJuftNSaqoUPXhs
+Ha74NuDTfJXXZtc0kPZYK0EwrnQQ9DLYbXjwSEYkZ6vtZMb+l1iGbwek2+Z7pMzBd7lolzis/xj
sdmcELOpOZnc6HWf6ZTv2105JbXFLMDmMssyJFSJn0Qa6PaCiDXsdjJuhv/cMQWepEWVIaSN8pJG
CPZtTqMEkKGXarF3L1LGUIiPw53oStOgmmtDy084rHEnVHgt7T7aqC1LaZgi9FclQIgKKmYxlXVs
Ofk8O22cN1Qx5zYsq0mAoStxX31VTH2na3Ujz2Yxitc47ItMVSV6sy+uvcIFB71MuAl1SpmyVpGU
w0stIWYKThJ1Czul69mpp2nDdMHRTNkKc2/R4LuaOD141baIJnuMFiFw+UWmJ7wZUsKB1KTGK0tk
yAnf2yYOACro/OxgFVuX/hE+62A1jww7BXB52eg962SYFTVVH1n8j/3wR0M7WGc7/yY1Bv6CprXE
bglpBYz7UFuvsNc9fKLbyVDOoJrI6ULaCj28si2X54VojmvDNTCEzgcte55FiAlzZL7iPIejxPwa
vLc57lYIYFzKcSOFP2JRvOKW9z6s+P1RmWS8Neeg/pIIU6zl62DyKNhu1HmgOQnwkRwl/ZZT+eUI
eqrgx9YrAupSBaAeg77bcgprsn9SXc8qoeXef4ei/6KrX3X+QtIU4lT8MdPJDg2pXbbQUyEvpxaf
P/BzHZLRgh5b9WX8tqd3WM9sZSyJWFFQ8YXbmn1wfs6Z0yq+2tMe/3Qb8Z5QZL9jEdI53RUPd4zI
aKrRXBvjHH5X83X6hNUEXZYxjCiuEXAoSkeLNcOfzyLI6S3RVJ/JSTkXpcxa24Ro1DOawqtqL9xD
bLqDWnx+wXjYzOzAXDAcGLKY+NsL8CkJakmuiWPHkN6BRbzKpPa2E3OZtEcSui/XuFqNSfR+4T+y
1AuvZQnQmmOy+RDefTLITOjqlw3wL9SNBF84vlZB7VFcO26tbIgGYRCjo2igUS11IeZ3KqRO4S+T
kay4ky1VkyOFeiXUz8vVTVyk+Rdx5OW7wMcrJSFBhQwUaIsfJG6CwoVvs3GqrxHcDteGbNfjOmmu
jZVsx5Kr1brgnpVfg54c5VMvhun3OD/0U68BVV0kGecvm8uwA9p9BTudz6KPC+UzkI0zE83NA/YL
BNXVF/BE+N8A+jO14wLj7/e090Q5Kfxr8GwyQEfnLqmJirpLwKfaVFy1X/0AUCsfV/kDfgrrfer3
b4mocF0q/WsfYgzIuNljHxyekvJR9ZY184HPuYU0S2tZ3fO/ZkUQia91/uuQXPTIi/alpv6PbPSs
LE6Mcp/oaQWNKqd8JqvXMD9+RvbMESyFkKGppppGVK620FB9yrSLlznwFd9ktq5w92bFTZK2ntlo
8jI5NvEdX5S2FqIVWt5Eb1E1qDhuo9WC+AMJxysRnGtWz20GXSX8XqxpPq9TSID4Np41hk4bUBxf
oDWxBbNXBfznv6v3rGKuTynKcFPlw0ISyAcALTSsYpY4u5tPmakF5pCsCOsDalLGUK1BDx4XAIXA
y94BnAST+yMpj+/4sXqCGUyEWhRhil/Ku0ivFKfkuilgwsfJ6oHLQEuEh82O48rnmRbp3tR75Gzn
+h+CMmnj9V1yetponhvBVM75UHgCDfGLu0LgJ8t72W9vV0pxmkQpEvpFhrr1ZxpeIdAE+9VG/GED
9oO9bs6bmwaHtTpeK9U4jm2UGWa2eM7iKwhGsQYSOMCEOwnb4MIOu6tLbgG0k42wkIKWJQvbgxgB
5gNIe4YDlgHYuOcNTJ6WDnXBzj+JWFuVaQlEw5gYjB58j6V4fO4i9rjB5efeYg7PKfL2p+56G16N
d1YhEZhrM0nVwvd3GPJliGL23ZdmovxUz2Ex/eSl0mIImC3g5x+x+6R2+sgb6nzBgZCxQVbqLJwD
yofv5D5bM4uPSxg2XpDDzAisJ8Yxm8L0yA+hEUoh+UxCmwkp1h7z00AtGlTasVYY94V5r8YfgTlp
HbvZpnTo3V01iNgeM07TRtELVKmuJEmMDKeRuvQLKNarr+13KBpMIQeCCQ2nuj7k43+0S43jr49d
lqBnr5B6QJ0XtRYfPL2Hgmp2eqkyVaLDMlMuQZ8HW7g4Il8xykrKzmHHsMrRCCB9pnEHO0tPXaCG
/sXQkw3fDrJWPcLAcbU+t2H5cosB5gYvcy1bSB7MotsSaaT5MHddc042DrZ7Xi/v3JINQolUjreS
DarQ2fipJ/vNGF1z5Zz52bpBP2y9Cq2kUHzj30NZbcuIDP47J8yBtD0s1gy+EeppHqL5hCzFobXo
OvFIAYZ4IK2nwKtU9YloJ2BBOx8sC0vSiG1hKXFvtY5WY3UEF7smDVHcIFZuzPbH043R9QZDx9j+
9AfJNg5SkKdgsZQuxs3c59VzB+MPDdvTh6M4H51NHooOdNnk8mHL9J+QljkVZs8dtmKC6x2IzgMS
jFhcz4oosrjcujWgCof+uqWbJowOIL26K/ggwL4K0dCFx6jZBsRZg3RdnFjteFRofrYqfH6MsHTN
E8zi5BvvuJsysR5GlrhSgDNj5FFZnmVYDg3W5g9vpcU/tqJUsS8XZsX5ecbjrZSsMwmqdXoe+HZJ
70vYYlol2Rmo199+OaoOacWIHTEGYybVEdn1DejkpxBKdzYupsJ3TIMi8TRU24ddHCY5uqMyb4eH
Fw8Myd1OxUAPj97G17A78ETktQxGkGhJ0L1CFxKV3J2OxQ1xTXkHhYUGPt91iRmikEW0I7PnEldA
0nrkYKkZQJxtGW5PQYH99s8hy2v0dhz38NK1ZimxCjVFuY/tw+mhBIycLWMVDwoIVg9QJEa0TCj7
kQlMSTOtQ6FN0LpCLNqHmmDvadmLeGID9b/y0Hz5QMGTx/fHAdbj8NP66C3ekY4z5XScza6hjwKM
XV5I/1ky0odsTLEYlefKWTGh4kIEn+IRZvjhG0YjAyR43BOoN99dsjA5Z/UMtuyhw8AgukWvx5lJ
kQjXm6hPtBfj5lnvl6ELV6eHP9O1iUSJzJ5lCZ/93tTtBeNtilEGC7MfQ/U9QyT4/ZzilCJnzMPR
wryr3pQoN3ER1BCoGS7QWwAoVXWIQLm8z0ICtksAPlk+VfPg5+PzArTHsn5wLshaQvrv9bdZLeny
NmcQKYqTWJC+BybFOSaJeBvL39seCZ0CIfNNTfH6ObXm/RlOkT8aXLdDzaaaDSQQ4EJCixw++5mn
1/tVNsSwphadV3wHmQH8IzF+3Te4IztHHcE6NPcbtR0aF5XNW7py8Fv2RDyA2/zWBqdC1XebnDQ3
ijLgIX8TIdkFHVNeVhyNCIfHhIMgg35PpAmZ0TIoo1ZDkGgPIzYjv3SSgJQOzHvwG31B3835MYLI
7miWtlobnHSHecsI2GtPzJIhQuBGRchkqGQhq9vOJhcvWV+V+Mx+ubQncI0p96cV1ohTaPlWwG7b
vj6cL3byq6KpAXOc+X38lHt6eE9Q3JsdfgMiNh6e+wS50BlQJtiZDGIovQQIks10+1CM67ZQ0PRh
B7i3h3O71DGMFv2DWi3ArrXVPegYQ8FEkKPXCZPhjeq0r9XyPrF8HQ8rmd69Q6wHh+cyaN/qhdKR
174LF3D2ERaYzjpO17/zvIgjM1ldm0Z/Z7s+8Pb2wWOyzlWSmsWImPiUSIv87Tx7Zn7BTYJLMbrX
GLC1FIzeS/eQpkdzTXoDhg8hePA7YWcT7CtEUqwzTHomNVhipiAWDZePHvPw8amLFInOJhfLRZHh
TxV3OpuCDepfQ78rIz2/MfxfqaKcxtewSt2WYR87m4jsHFfJGHq6h+S7ukUNpuarhG91fm3mBwtB
Bk/6kUX3Cuo7kcxO0txyTNfqRRqJaT3IQp2Pv7xmIswRQrbOKkC8m6vjw2iW6XXgBPu/kZ+/NNij
/QimMLvBVUevxFesihmvHTSlZadJ8VNpL6MgrRmE6dc++yopQ8vpH4+PYe5bGmkyX9gu/ff6+qL2
Rb28jRp4bUJhUX2KdvvMs/1dnti97GZOI9UlJ5WyIWysC6l5+KCQGa58M5Ei71OQtq6cCKMDdGtL
B3BYf8MkkVOFaN9V/vXEOzf/SE4Ld3FovYpW6TRnZ4AlTivYqU5SVBjiSFUrgZoibjf6LSI6IFXf
9hfJlUK6/Zxh/jea30muJ5bphh/AnP65POlr3uDOmiHpZzmZmltd5xKxX5PpXmXnXVJgpgRC6qd5
YC1WHsx2lYHwSvLZ7zmIL6YwCG6hdcItkdnalvy3LDLMMhOo6mwADzmakebt9JO7HcfQ/WK1mROk
2qHLCAbszBFYNUq/pSdmKruqkxw0uzrPyh5Dbwby9bEESKYsatCresxpI5isAcVLM83Z1mYhzTUW
BmTHXkhGCGS7oU7ADAcsnDKszvsBykbwqKZTUTMwBuu9SMA2s2FOuz4XKc5svVBi81/PQKScREWP
legf3oMt7dtR/r5E41pTXaUDOtIp/UhkTr1zLo5EYE0eGFZkC9swQ+OLkzad4tv+8vP4iaZFF6S6
O1Ys6BcKSGoj9xEtJe4e8+cexCLmIt1DFk5PFhFCcltJlhpWPiuPsaE2+2rq5aN05IWHYqrxIAfB
Y9/FoYXD3PdD/diAe6WnKLX7GKGTCLjbNI61EGuJJUMtQ3Ly0rGMQ7KMYKV5ZTidU6tvl2E/zhWz
7o9nm8FOil2QP90WxX+uIBBUUZ/XF3VUvaWEC8DBzDRE6ZdbEFRU4LXMYeXybhbnbkDo1hv/UKU7
vCPWcvZQZOrDHdONtInYwzgnyoVVItT+rjvLF7/G+Np7hwDdbKwAuQhSfteE7lulx2xXgcKqltqK
KNhC0KWFH85HGUVSdA9zSqHAG5qLuQoxsLnXBxecXRFs+iD50XVYtaUzxS8wECHCcCu5bzzXVkLv
CF90TOs8xmDMo5f8VcwUZMnHv5xCYnMIBUJO0l86INrbJsf1IqSc7+DaasiGPxlBCHR2YFfUrTAm
3XUJ4Xm66SmpRuwuUZdZ7ua//709R00C3kzBz4iu0yatw5NL5in7ta5tV1Ek26UyRA8mf82vQx3F
yEdYUVeKjZFv0Br3l4QP0lsMBPOE9/KBZ4TIiDqKx4wiMMSqxkq0aPJOMnQHknHR16RRIA+GQVGH
vcEsDyiM+LhfOHNGvRykFwWWDzwEpCfkrUkLOgIESw1x0FCLlYadQbzVP4LTgAwsVe1Ku+JQKSUc
Ss8hFHADNq4HRlYcd+8NC5XPaQfA0lCZfDV6rllicJ3ma1zEZV9L4XWzDfdpbFuuJKWzC8X71Bn/
tDodQ6V4CbUo7uAG1If0L4LPUeAyGb3AqYdxpQJ8mJtXRTlvKbw4ydl8eoaUk3npPKDFhbAGxPoN
HeIyUqGkdFzeJg+AkFvN3dtlagJLuHqU+Sgup4d97+q2pbgNO0/XnVHrJ/6Zt7IKDdzcdcN4TZh7
4pafmiMqyUxgVgzoJKn/uH2vx9HVyprvRqgfadM26ZDzbIXNoBnX5FKKDbk8AxojQaEXSHiuFS2u
2RmIqrCBCKF0jBwriFayVic0VBMFlU4W6wmFbC2Bikss/d3HA8X1ZYTx3FGd3fQaXYySsNIycKNW
Ew+r3hGhM7qj20hGE0/yK6lB8GoQRqGNUyarLr8cvq6idriBgD78TO1mjRDDK7CQmJxgAlLUAaUK
nIyQvl2wtXdcrXWayWMA8tWxYcmqcd4eIIKhKPBv8pE90KhdfLJuKRn/9/1DNZ86BixOxRr0IR9n
vD49HCrUY2mhJgWqaY2ANyqXXfdhZnjwuME+YXtF7AY21p/H8SEdRXt2ih6ar6nYS08uN1rqVaoC
LienhBdiBzf6mOlYgx2UabUOjVoX2Q2fKJ9R7bAWyBxzdXNhZlJ3/H5NXSgE6EgyjJJbWqw30VL5
7YUucdwSkOFkKCQis3aXV4GwIHpp7ADVcXEFg5qR4N4ucSd/DAvLGczT1014aFij7gGPmSa1sE9z
w8hscK7Oazrs4q/46dd7CTgldH+liTfU+6rBzt/Xbqh/GjCWmHcbkC6L6eRiA2Qk6kH90xTzDn8v
OkMA5Tu8QJXG51t8t/8UW10RQKPzFYBFZddtKsDpQJjOBHSIcSRikO1kOPjG50IHl87Q+2pvXeEY
+UQ1zKBaWMaf1roku2vMJevStYdWC4IO/uXNgYY/ZFY331FOGfHlKyQd1iSN3pAJBzzzR77bvr+/
yRrc62PZ/U/LnockqFqlXs4B6+Q+gevCZTq6sGwRFd+XnCk+WBPe6vULcpNiAKivY1jgLwsCt2l3
YS1iXMEzEEhgM27Gk1U5JvXRI+hfXxG5ePMR5dk+ns4OxeROqPgi5DLQ5nhZzzE42P8VwLPdeHzF
8JNUYjtY2y0TCOBKIh1SkofUrMeSqqJWI+KYMIPwbl0630DRXxXIaW5elJi30m6rMlvA3j0wZEgc
WcVAfAdsTsGUd1xZBgtcQlSwS4FdveGaM8DxmWjdtFF7sEnIpTiJ+ohW62ehI2Z9gu5tXm0Dyp2v
m1ME3LR8rWUHNOiu8437/JH3wRIMiCLNI+r+n3MuTXnVkUxmtV4DPIjnLDP4cLUU+wgdDBopJD3U
U3anOwTa5ULaCj6qrO0EeoarpfmCy7BYrqJhAyvaS1twrPBBtkO9ilMd3M/AZDwO6XRUm3xtjxnG
gsLosMO0oyl2WbkosikAzCtMJsMhLWtwu4bTpRLOCzK+NmaTKWmORgZw3Mg0ReF8qorYrL7k43va
wdI1YPBzLxyAL0UhodKpyTtJ9ChxEU+Vd80XnENLL3y5iumongqK+yz988uSGW43mByir+Dab0zQ
uPKruflWwinqhy/gx+JYpFjss5UopYyBzhmZrWjq+lxlC7kh53hGQtIlNVN84xqhpbsyva+FVZAD
PLuVMsyIQ42tePnH3P1lFSgL00fOAetDI7XwOozqqMQgNzvGBR5oZVczj7tfnlEiOwQRxEk1NKn2
YVScokoFH5bZZZ0YVpTlDCbuZvABCsisw5ysitO38JuGdLoRGPJahX0mpJaBqljhWKX1MKZBaCzr
t5shlQfb+R0SozliP4p/zsUHwv1cveMz1+Tg80gIy5iQpjeV2dmyFYkLz3fcGPM6SuPi7ZqfxiWQ
xJH0/MrQxqwkRaECN1HoTL9+M2ir7arFdxRFieIM5J6nxjUOjaCJGFjAYvdnFlv2Bslp+iRUUlFJ
vuvPYZniHT4dyV/6Okpe0BqEyy/RjMmxWvdS9OqDHYx/rVPTiX7npzRPIwQyYbw5Nzl9dK9D35Dp
8oWGdUSGTc5PUCckrySHDmyJtcpvJ1FWuJoXrvuccrrKMi5CjDJTWG8j0d/PkVJocAiliU7el2z4
UTOTlQ7lXRHM77GwaWa5RFTPZkLshR5I1/XDmat8RkqLExNrifkdezkHwkYBvkvW4pe2o2g8Jf4+
q1ahemSI6jYsHPPDqELBzRYjCVAYlG3fIK435cUO6AQTTgwi1YyM6PBw0irRzCVs7EMAYFdgtJxW
8JRUHhrQXjnAcGv0iyhy67DeCxQb42rky8OKkP5FzauaFuVUaHgPHfV0UZXCHZsX/blIvfxC7BGT
uYQ3ajb1dZO8b/kw0LrSsQD/lY4o0pM29FOR0IjBuIbrj9i/6AtEM7HwENSDee+Iz6bDI2ZjxQuf
Nv64dumb8FjwOiYnsmvc4UX96HPhhRAN8qE9lvyGkQgvlcMVWOMfjXktCZILIAeIyDuLOwVyCQB2
ju8HLa3OZlkpIaQ/yJaGzoUbTB0uN30+wsyR6+4k4WDbEs5fggpPFOz/PgcKWEX6jeb4mvKKYT1C
9K9FOH1BRlOsd4y0YqaWeRxK4Kvsu+fCfFxtZCLsQT4rGZQEj/9Yd4OB+0/3rX1xP9nt+5YLxqK4
0LQjiqgPdvbApZOuNCQXuU5ZzVnYkKYluVXioYAQ/zOg63/zyE3d6WQo9Jg7fObDvo1L+qDniOyC
fv71FOScDR+mQ1UNxJsxcaA5Hu3/apIVzmIUskncCMrTf+Ww7xSSWWUVRtb4xq6GWVuHNSmfU6UL
H3SIriRQgpfUUV4RDjH/c+23enN5pxn0/ZBk4C/1nNChcC0LZWh25SA5qqsplsXyvr/CZAUnATEj
AbNY1NA0uYqz7WVR3gUs4f166mg/Qte1mk/KWhdl30gqJYLyt9ekfrshbwypIseYDazJFHbBsACm
R9lx8yCPi1r85FH8zhCYB9WEgB0qxfeISEI4DHOrj1azdCAIkMTfxa9eAvlzOaDe+G/7z89m/5MS
7OUG6ctjHoYL9HOFHKWQ9H77XK3PQDxwywO3rCSNwiNUb1JPQMmxkZ8xCtYluLb3CK2Gb6tiPTcx
5vd9HuC1+jqrNh4HNdAiXe5wqiVRje7UxjTkZSnWVGHujCnoH3DkpvF+3VLJOjuUEwI54yYID3XS
HvHkgRiFtusp74goiP8pIStveiApS/YBx8G57j3CpVtse4cZw7SxgTYnafu06uidXXyFeLHBrxaQ
hDsqiL7TadZqqYi7BGiEaxVdwlil4gBkGn+slmw36zkJ9AOj4i8acf64BfWDAY6dI4NsYqSicIzr
RNA8Q8bbqrDLIfsULFoGhgT+OGcRLyL2zMxOHzD0HUB1Uxtoe9/+wFJ5lNOIcEXUBGwejMsP/JtV
WEer+bo9okSUoCEjwQNM48Td5cgZ3agIWkpHUKK42Xucs/RmP+eXvArKldZi1jhBAn9Q/V5bDr8l
isVUG81jFB4GhzeRPKgCef0Qk4DNMAhSeYnPqAwBq5607N5cc5IyMwBwOEEQDoumMpKOZUuP5nO6
+TEA+I7LhhKDzVc62Q2K5RLb0r8Vadzw4v78MmR8lP4iaqt8ps8VyYgXD541uvAZZdu4UfbBgOZz
s/Oj/L6r0fXJ9Yc0lDvCoFn8rhYqhUyDSFwqN1etNoSF/PyEACy9BtFdkm1RBbRu0OuS/nN80IUi
27wygbqviuZQSFtMD0b/bW0I8x4Uxp3Q1WRnCi8e2JEqi1Wy3nNYozIO36UkO32QDf0Mgd9wo4HP
VtC2w/ZWZnp86SRLqtCxOn7WUOa/JXY8xQZ5j/C7MC9an2VzD7VUzpiF/3+VBi+vkBQFxe/64erj
LKjtuh/YjkodsM7FA5Th7KGTBv/NdIaF6EOCVPaMVFvzSjx1Xgrf0Cf6vUE4opuGqv3dO+1PE9I5
FPVdkAMILz0KpnqaoIOowU9/7HjzMSnKxQiefH7v8Q/ZvzJEL7vhXfox1NeyiugEekBtP+JP395B
7mDr9TO21GurQXIDUSOzEwETrsjePQe4fgB9CvLmvqmWH0YKNGWLQP0yjSZzogGafdUYA9+1ijxD
5ulFNP7QusgScHXa4Aj7Xottx7z3cV2pBOmTFuKNhmXxEtVgEVmRRPI97Gj5oYWAI6cUnw3kw0jK
OY4z417RNSHnqHIgi9zo95pq6DfIgK6m8+1EwOCyNJiNGk4mgBAQvFS+pu39xtoQrMj7OmazjLFI
l4Fu0LNeJh13q4c/COk7pTTo/g7oeeci58zMhJEoSCDt5TaDO9IssjfoljkYdkcKnSy7APBU5EWz
EQh27D0nHFJvVsgmcQ9Gt18wTWpIrsWdvgLwBj9Ev5Bh41ltp6lj0XYjDmTJIDX3R89L1C5Pg8xq
Zl90zBlYoFHrah1XKF9r7H8iZWHAeR7IAWGFLRNiPIH+PTO6jmIt+f+TImyoEAv6wTFW21/1myLN
AcEHcpwfCryGQjgPEmNQmqub6GPzfkdOInhMPOj16FB0AmhQ3iiIEWgE2fmadOou54Y9SqghJGj6
9NtQgrTxr03eGVFvTyrXknkengk0w164kfomGqHq3n17yyIyb6WVo7sgo/1n0syoMsvuuWQ1V+vn
sUV4e2lgN6Y7o8B1ekzYCBXkn/OnFM79G9BEsdwhz2MoZWwumdS8OQoo/RkoYmxxjOat2F4xe9cF
aufEpx89XgvEg2WsjibRfsSmRmtRpFIg0g1JSUIHh4mUuMDTZ9dbHxkil6S526o9QEQcurXBH2eH
N2ok88GrBjPuhgEJbFX8wzcmGM4BeYLCa0mMmBUGkNtZVHNxC7zTh7iDveztyaYWXMhwPZFqFDNN
WXl7qAmgCYQkDt1vnVGuwT/e2GRzQNuyCsTCMAuVcTh+rO9pnA4O9ToNSlx8PRIECouxZrEKTN49
rNUZ17MjgOvTq2xhik7jCy0iOlfPs5MllGRYXWr0miJ5ZVUs1xJuYWx5DjdF7Ic61w16HPEOUUZ5
lBp+G0bWBH7596yoHgOgA8tNaVM+GxLvx5y9logIZljZi2Zmgf4ZE/3SoSd0lW9KCjy7vbeonLx3
8FoC+eNUCabSf57wc19EOb7AzaoyoUXGNtFUPh7ZERw+Fkt7qmBNY8BXBQCTBHflkv5UbhpHjfPt
admmsRWpePO3smJrvKkh5STq1QihqrYKePxLfPVZ3shF2zNyLqgxsA/Q29/mE5dEB68O3DL4mXk2
jEzfAFxfVteL0m7RT4G5WkLhmBxwKvcj4hW6tfQtdYDml9p2uMyfIYF+TVH0gLBFO9+mkVQ0oyZp
A8w/Wk3KSCPz1Gtlvd4utTYFuO7QjNAqWIRk95/McrM6uOsj9LbzDzt+4NP5zG3pXUZk7HmjhFdL
MzOFzF4/a0VLGsQjeJuVKTtpRnJAPcvsVDkJxwzFNj/cTPSqY8f5uOvh6QVpMw169VfBFIVIb6Yl
6GIJA4eIurno7MOCIhIBPUP4TeC3Cy4F0Nvlj09tAmOWJthX7tCXbGmUqmzwQBSQuB/PuQnOS9uJ
xMKY0dO1G7PQIP26grNdqOqhHHk5yIZ5uJYs/RPK+BNqvCy0SCp01Z+sDaZDqSF7DHgjULbbHNSh
DiepNzu0UEPD8f8D4A7kvVZX9GehIt6otGSgJq/tvWedZZ/p6qgDTSQy1jd27040nRJwKH13szhN
BeBBBrA9fbqwT3sYSqLAn+suAfXIfRNoDLENkQpRV85ek4gUxvB9dizMEZ0DVgdm6eC/tCD9Zwv3
zz2LaI46Cux04HOqOkOXZ5qOfWKYLyAGHxNR+Vn0r68B/svMcRhXKANy95yF19GQ5+9E7+9uTAWP
Qj73Itj6zpznc7SNtKJZQzJ05vfi5e53c4sJZhNU6+ZEPSm+9sUghfZEp5xZ4RTSViu3RDGTKdtY
/EzUF+3B5FLV4U967yFRWqtP5EpXYtXrwb2zH+JqSU2qPYHu11xISc70set5+QO3kr+f9rrGoImr
fubRFu5uAiI7qDGIzGkY6JlkpSMkGRg/CBDMOGAkxFieM/dZNDG3HdqkOJhtsarkOH7CEdnTUUrJ
Wq0kW1Bzw3dX5EqWlG4pSTMpsV+ZKGr0cUrSb0iADylbUfK8vZVV6EFvKSJYM0q+RN9cSpLX0Fln
j05gy4siwp+VCFSyhm0Uh4S35UXpV8TT6dJPQZZOBEuKdMWMegHdc5xZufhXu/YsUqghQGHnuTDj
Uvsn4X3UMfehiIykSxAfIRAvGmzlcSWBo8RnwlBFywpyTbhkbil9vpXb0d3GPKHg3oYfSCtL5O3r
IJwy3Mr0GAyByBpf1OI25CfQSiJtpW4xgIumGlAv4sGhSBLWjF0Iov4lzhgoZsHNCKOxYwfA3dHq
CmkknY4MuytKch+MPkSlkdBpi2TiDBz5Ro/SEY7Vh+ku6TH1hckPZJg9bsVRN2o1GxS42iVkUwcp
LMsokVwkIriHRsrA43BN9jaAwJg6YmJcVKtmSxc+FNPEvjkklMYlHhWnjkK4kAjtcOztiw0rlzps
M78VWnHK3q5TMC0IpRL/TLciuOZjg89aR6KhxiJSg/MQ0IF96BNZHrxgfMKYN2GZKsCpJflFHEVJ
o/mV844U0A3MCXN3SGT2vqlyanmv3Oy6qIjeSoDRxQ98qQ6zIemHzKvz8FhNkUm/DZo2KY7Sqgnd
vndv1t/KjYS2EB87zsYa047zCWM1M5+Q/PrFkCTIcbxRsGhcODdgVLtlymzoz4sVJForY2ZB5q+L
gn4b9Sj3cjppgGg/srRIoM0Rp9q0taSoe0DTqNzgqv2GjpNA6Bb9piJEDqIiuQjzFVRV7lQLR6pv
50WBfkImnelIZTdM1D8C50jZvByDjJDRqllILOElv/0itANqVxDKjxeoJQUN5LtcUUYJcUSw8Mg9
rDSUdZXSSuJd6BRMujIL7YaugiO0TT60gi8yx9ObIOGB3IhR9uhPbtswdDZVICzBceTlnBqKu+M+
w7uDbHAuwpWTAZ6trHnEsggHSvvruWcgavZKIPMV630yQKl4WxHGv4wpzw90LIVzir1dGxX771By
jS9DMxI2dQmCIAQso5Yv0ExYscoQe+SgD60bqDPMy31acz9RVY65phvdSy+G58jbdnFGtGKE95WY
SGhib2b8vnBAgOllHga+hLoLJK2LsP1Ur7XLIWZG0nbKon/kxZfOX3Qq/0UYczkZmatkm8p7XDF3
G6QhKT4nh+XtavIxKnq1qdsMFgdYGLUdhEHGSdKrC3kdC0nzpEXwqU7QQ/r7UCYsokEvekzzPKZ2
GLEd1SmGnHb400Bsqea6uDhJo1T8jk8a3UHU4be5PvM7huYDMJ2WKyI3vgEMKHvm+3ByN5+Vqr/r
JmWmHuFtMAKXkORetPzbYy7QKTbqxkV4YXDa2959SyELaGXzWPaazR5z7atIWdu901PN3jIXOPZM
DXVkTs/IHWpDzrBUXgMeYj66phMxG4GwM3B1d5wMCxcP+mysUCnE6hpZHrkb8XMFAtdMXvWvTvDh
SIrz2rUUJojqTKwTtRjAoM9ymZ7IQMUry7LaXMg6ct1ki5sSyr+khbuqeM8QIt0pCqAlqP6I1QaB
ILM8/RI6wqXARdHRPOxOt78sStCLsrE2muSIOSydEqeWIV/Ir3ekn5MydWWDpdl83j5DuL7CTeRJ
jBGq/apOiNeVy0FDw1hOD9p/jg47zBRU26buhosgwGW4lsqXCbHQrNswhue3XcC7MT6nwzjOcylY
g0IyIBCAAtctq87qHV21p4gs8yL1vf5ZwY1DI8XGWRir6bsa/GkLtKHoK5h8FdCFq9nxoD+YsPVu
G/Yi0XmrbLZgKP5hqBA5TGoy3Fi9E4PEgo+ROHVRgtE9F3d7LWiGnIzp4+XHG8abmTcA0BI2YBNt
cJgQlxYG65+XP74hh1a/xqdEqkEAEN3cjFZFgh01CLuv/Dq/IprdXMU2AMi+U2A+iAp5VcUn7mVh
inlFEOyEhGFYOblpImE7aa2c5RHS2ExS7LfdgpdRIA4BJ8xmUdkbyBcYRmHGjNbz5x2oypCVKIDU
nfKIkbhmIWFQH4thwHO9YWolxtMzo1XM1hB1N+wzB3xjzDJ7IL1o45pT9G63GuYaSDl6y0Mh6ShO
hEV731pIiSGwLkxxNPtGtPi4HDeWeSJtX+mYBJ7G4hZPbZuN0IMgTjwjGnbku09nWDSltdUX4aN2
RDucUt5oikGkYdfwR+vZm4uBS5hcpqENjq6p9NsTKqZ/7uFo7vbR1G+N15CVtOCusviWcKBxZyBd
MRIIeCQXhJmWT+ENlniWm+MiUVpvoyyakC+xNChR/Gy/5W1auM1k51IcVSSeNJi+VjdIDitAzIMX
SvWxWpzhJdeHrxL/x4MXbHqGo1aucPJKIkCuYbm+aVEaa0J/TC3j8ht9nJSGcfs1S6FXqRzF7nbd
QQ0otYTx8JvTSW/XTRwlLBwN818qQKHwagow75cK3gNgxdLSkJYJPqwF4DhHIRYegHLQKdfnQsay
caFttliyPQDQZivHvvaEasuI70qZiUmHD+N+vyccW7CCORlzxnSdACgEZSKgPW+FFdAvjAb5oaLI
DWIJTtBJ8OKYoVUZekLDMsbz/gXzMgVM3zKEzHz5fKSO1qnfgql3m35FyETFjlve/nx29NFGerog
K93YgOZwz4b0EV8DNNW6WH7GFH+rSDZPYVtS1UDz4jEifpD0Pn/kY3e/eO7naMyJDQsmjgP3LDaK
9KrawtZcce139yXguSAuCpC3upXeQiPDOwpofUn1b1XKvULdAZ3P3VR9R0GpnnrPRzOS02LVK1UB
hxMDnRiwInQj5sGERDBdUuYpw+8bOgmD1gnaTme7KP4+ASReApwvAaJMoCumBvHJKB/5X0ezXWSX
yEiLC0LnbA8gum6NlFv2M0ZBE+P7V7yg8y0uG2cSNEjA7r6lc/OEXiztWRZDBlz2uMfgdnZ181+z
E9U88ePac1MxKQUfuqEvIoId2PflCNXFGoG54StEsd2gy4FjazCjwii2rKe/34GNVx6OlCpRwcs+
vQbIKLdydqyHyvMRvQ0q5R2/+0gP+yexCrcHjA8Vqc6dbBGc5tTCeu5C0/PusSJ0zaiZC9OKZn4U
ZvVTYH11BI4S88xMeZuS9vT2P1lBz+uY2odOasZgzP6qbscYAU1bDnhfAb+4NgqcFe8PnqUEDhU1
H6RBL/6QtA94I0K6faLjTIolL3brGwAiSRqyoq8ask29SI0b1aQRvlavG0ian/VcrFtUaXZ5LO4D
eVutFgsuo9PprOEIFdYP7zz8rsHafGP0f3OQMM6+KPP50c8MMCzqBByga2hB/B6ijM/vc2ibVEYL
PrMsOG8ChvkhK2LRAX04ZEQAK238S68BtXCHRGzkGyf/SnEGMaf3d3HwUC7mUxePzMpeV1mv6zzp
bo62Y9O4yWjA9BPrgGlqVXC9b/75M/kn+nBP3IZ58W+FoYyDzQqd9K/Phnj/0wPtNJmaL/zlpRkj
lKUkyYoTzIqemRz8Pdn5yjS762aarviRkWc2tBncuncaskkzHLYOCF/PX72XUchaw7fQCTEY+QZn
VIJ9JFZjTW7ei25OucT++SOIXDUKMKD+feng6LgtrxjxMsSM6T5yv+mZG1WBsyBCTFytSFaboLiG
TViCkecIkKSIPmAFJP7THDqifDkDGHGqk5uTTvPk4GVEE0l9eSlZT5k698UxnEhzrWEp5lBk+hH+
LlPxF0xmWnVVM23dYPrLmfKa+hycsxdg5R1H7+bM8XzJqtvFAaAgno9ESSgOfW8kSnjksmC4w3oi
Nwgi/BdlRmRNdARGB0ZntU9Hhg4gTNgtYhAtW6kETfnNLUR8mEkH/iHV2QOiBnvXyxKTdqcq0Izl
Bp/5Dij9vVz1OYRVHRf6ikNnko8CofW2sOZaNomuDuMxI4KDI+M0V+jErFW40/Ppgfpr0iOzcSvt
YRj6yr2UB36hOwsIjPlX6rNsketghlE3ld8Ofbvg+wU21G3GHrbbeDNoQQunIhwuqWJqADI5eEYt
EH3NJloP+e3mPZzBMIoVgfIrjy8JBJ8cSXpMa51y8zpSUPuJvoFnZWuPioW6cAvunEde52reW+Ih
yjtgNXkBKkalkav97lb13Q7HolCy58MC/FAf4NpmtH1AH0kb6puGhoUY7avlHxWA7YS+He9Njr4j
QDiUTmk6ZZpep5qi7OvLdqCUk8Ripj1t8EaOXPima6Xr9/oNJVN1G13ApbykiYoqngu8XXJ+CJQV
UhWyQXZAREWZkJklpOccYpv19chvmGHVXDSJKpNyWzA0270iCeAWxXgS4uWPqzrpZdWOF/jaOCIR
mXKQgA8Ek9UnQickWwmE/MPyHx2NvsmnuxVPnEeb9DJEoksYNSRRSdfPPEY4vyy2WOFgWroQ3C69
IGmkqzJ5QYz929UCy0CeVa6NUGrSAa7oPXGjYFfmfD9SIfOCKr0g5h9VqiPj2NAkMBJdzMPuP2kr
ttThxvwRTVX+O6m1U0KX9tN2r8QBETUQ6i70R6RIX+ldi0ze00hj8Uo5R3+NYq3Fpl86TAZv84p8
9cw1/Wqjf76qvOj6Vz1iKWchOo9jDM2kAg+bCxPmeRrqBaPskHOlAczFKcsRCdDrV3aBTpwOexCK
Mab4OzZdvAOyMWjvOFFrLIjlg5P2wHIvIMtaves0stTDxx13nQjen55EKsZ4UzgPTt7LPkBtCaey
sICX7GI/DqN45eXR8BOkdFdsoC7ZMK9+shR85+5Uq1bPlX1JlKEpPe6/StaPg797sxJVpBGkb0YJ
/t3hBrIfyul8FMjrplo0o1strGpBQo36dUVitHYDXRBqsD4TX0A/qyOSYdH9bRxv9ZJL96lTNWCg
DOcFwRnFenY3S60lW8SYqHA1Nx4jhrBoO7SlPgD+4ZMiBB+BajWN3kphrBMzVGgEzRe19sDlahhi
IlGWEYHtLVh9Rp6GjkQxg9m3y0m8K4/Ge59QCOyj/Uk3L+kOJKvtOsFl7V0CxvB2+Xp13uRXQ0xR
bpMXStSsGOXmWSp5kCYV/i/id70FBW4wj1GaU9Uw0pFMI2uSsOyrNmdZgxbVUbRYaLHmsRTJ/jXO
jzkC7C1gJYE2tBdastyHwLMeH0xjsEnGZfgsPeqXlmCiJTZ9ZRKDn7esFffUghMaU2nyvQq8F5iU
r003O3K62J8ZIZiv/Ly4PsdAeyNrRVnlO++K18qRusnfb/p2lVoDIYTFdVaiM691aZtViWCDox5D
TrsirC8jdo6oK/iB0m+rSNaAJ28rwgqjFQz1N7ihWXld9Dsh9kSlNIwyZvuNr8R3k4URRR0Snac3
uqus6DVUisAd47TZZZDTmXjDVHBSVKtLNudrQZ0xCo9+PNkGoanG/8xqcQ/JjCiQeEixnOqerk/m
G3cviDgevncwHn34+3DUemsFbnx2gVFHa4ORBrcmV8oYwAwJcvj9ME6Yn5oI7Oy9W+bRaaIMtXoI
YQ48sh8PGiFWN4ncRHRh+1mcvvVpzkyqBjwuUhzHUcyMAp3neVKjheHqzM7/wTcYMHr9OgoOKX2l
CD65p7NB49BhKpRl7nxhtEir2Ni+Fl604Pu+p0kfEpEyMljD+Os4WvvAQ66Vh9VGuIxTeIWwUFLS
je32TMhPSEyXTJ0HzeunlDLrz1gMGz1C/1mBKyEr9AZIyyOoTPnZfS04SVk3yWMF0vzeqjJBuYiX
LsmRwt3ux7vsjk48/4ZakVxbgiTLkGENPSgxx7+Jlo9mcI/DypV37wqUFcQWJMvOwo+dYnh69O1P
5FylQSvlI+jrlA/1pQDkkNQDeHi6Sd23a2KT8OLUvLmazYqPgM9GcABUdH8MkBU+4ePAQPXB6av/
fT+s/r4bkvyx8RxR7XEcm9GKHIFUzSRTiD+LT0xXpMBAPThuwJ51r1hdD1Xi0ILwsqwr8AaLlVc8
3vmQZXs3YhrO+65UWFz/5HRxWSNFKaNKQmWlfiLuGAen06lU9z0AxyFFRE0FzG8RJJ1j9IvkDARv
hIPYaKlDr4GRl9h+Y1lYxwVcuHKWz0zWrcy+2b66V94wpJQ/ahja1ENr2g0+Dt8gXV+/3mpJOWgx
cI63k8Feo/6FGso6iexS1+ZCGWyhrEmP/VSoYy/KiXiSG7pmr17stAUytUwkeS4vKPzSHIL4JuFc
YD/BcN/EfB5FYnKM47Z6+s+Fi4A0+cabS7px5L+My3AvwOkju54rvUPso9VKEMUHx4JnLni/4pS7
v1nbOePRl225y0PPr4TWX2e1yLRgLotJkEpHMTNWKrAoGECCLyOGXItSOb/2eSqTUhh6hTSAlb5c
9ey036xnR3SjYfJZtP8WN0+9gu53n4waXKk5A4UTF5AjWZjoEahlBbeT+G09tvbTdHLPAe+SjrJD
CP04mvuS3xFCX4vZ5BvgqWS15Uh8rtCHwT5KImp4gN7TClL9hJTEOrtG5JjfNSxVljiwli/l0zib
b8Ir4Up4ujaqFQBr9jH+JswAjg0o4TfR94OTF/I/SqBvXMb/KULDeyuJG1CXgkKLkqiWhhtvGGnT
xqdCmDbvprEICaNJ5UITQLt4Lf5QO7p1pcGHE0hJjFG2Q7XRbKSB06A4S6LO970CJ6bu9ZA8dYYP
hlhjVcHSeFJ5oeuChQ2sNV0ANb3ztR587Btdv3tnrbry0hIqVrMeFCmZT04UCj3ONEZcvv/DcXd2
T00qNJhhS3vZBDFnr+RRYqcprnOBG+R4T5nErK9IskzMX6zIvDJ6OcREVg8+gUt/oHeOi7E0DtQ2
kT68qLjleBIAF8wSmyFJGaVMyAD03bcoR5ap6kLXtoqMilJZw0GgOdCKJjKVEukae5uk3rILI/wQ
YhtVU3vQ21PC4X5B24/rTskh2y/TPsPatB+SVirpcWJEcC+EBOeKYpmT9pcB94HNHLDgccjuXNY6
rCSEu2NOSE1Js/U92UUvvVAwFG242vMmBN9ZREKwteOrQ3VzZrJQXTzUcvaA6csNxOONr+7/TXYa
a3V814WCZF6S/Njfw67kJYWHHUeUvfeKBfH8KMw0omkS5Kxrcjei7ON6q2DAurhOXVoT9dimGxya
CCGgqvCnnNUQiWq4rkZawxUr+NVe6Kjhnwsfy3dy3luO+dsDn+QdkLLZV7goLAZpeEmUIZj3CXYJ
imNy8GEoRNhTuZFW3skW222xTNrCyEN6OqvPOFfnjeFNU8eF/AqjmdZTSaYvC99CblxEk6Fg8L0U
Z/J8eKCQv8pr1KXzsz2R3OZefR+/WHvyElWp/TCkC9rigjBMDp08H67tasm2HIk74Aboi3cHmtxM
T3VL3OMzNiY+aKwn92lCQ2DuDLGUN+o0ED1adXaULe3X4QeseAl1WPjHYHeQizz0i6e8TilQvlt3
ZlhcHrVOan/r5sgSvg8WntTJ15kGME2cm22+U9MdsGhzvb5XvdvDcbk0y5RTO4DLl6+X6fWhxYQP
c2apXFc9BgWYYRXBT3YmxgEulkv386aXje15j3OvQ+ARz9fX0WPto0X7CrsAj0Br4zDTJT0KpL0l
8Lm61IjzY9Cd7Kxkc882h/k3oaK2XyTKQfmJF2/OPU6/3wJDW2eiiEnIVj282mu8zP+/JNGmbTOb
3RYc6zToacLgIXuaNkXXDD7Mu+UopUiIRFUsTigNlMT8J51fHxr/6ndzhjE63LOlLJsyNLmMVeRD
KF+oJKboTaI8EtgjEoAaSUh4prXr+1ZFhJzHbj5wfleDqNuJkodzJrBMYL7JfJolvx0d4limc1vh
zwW30y3pDgR+TbA3tbgGaEeT+vrjmNwDBWD+Nr3mR4X4Ei2nSKhpiqHQCajDH8dXbE5PbMESi7x5
yHvj/HLDVSsCr48KyCZ0Je97/D0wfDV3E8fDA3fHilk3SYiQwRQRbs4Sg/BSa/7PtugDH7KN780o
6wrTLAjkpCXG71NAbxM3gCORHGzpdU+ckds6prNNG7vhRhMffXzd/8l9FjPUrsqJYhzUJr+rkBop
StbY9F/XyE2/BGi3OS48Z7gK+tx57TrHXynGxhJehBpGVmP1yt+1nIR52t/Uk8Qs8dVEZmROnB6r
nhinucQ4z65aaDSxawGC4C8mqczkmbQcg5SIaVrix3UbVfSnOzoDQd3hKseoiC91CFmVw4NzFuzv
SC/41Hd8C8WU2Y+XdTOJzg1HqzoPQ4VOX+fsPiMjA52qJIeJfJVAXg91rYeD6+Ayg7LDmnCM75qk
AGsdj80bw1jOj3CbSNeljqQxx4At5TfjOWh1Z4xDGLvnTyU4QUSGCeBJtTd8g3Eb4FC9ELhQLMBb
D1NL9ZiypmUwHq3MwDBixCTTPf2z7rJ6Mg0OfFy8eFxVA3N/TOpDJ4lveh/kE7TmDfNiA6bPEYRt
Xj9zj4sgmnSXRKIhn5pe/y0MskVZjFummE952KsgSYRIyaqFqNn0FGgr3Cy1OqsPI1iRYiK3N3pI
QmBPE/lfonahqW9lRuqMv3hh0WoW590z9sT7FdGQPz2AiVntOxBkvBV0zob497O/73Up/D5ZtAmH
QEGvA568RuN54e0FqZG3A6D3+vbl7YPqWH5kfQQvld+mZDdoHblMmNaCV5fcdtPhU82PjfzTdlMs
+M5k5n2EYzD8JB2eb0fi9tSixTZM//wTBD8XkTTKqctKnbJ6F9g/TSpt62NC9OsWsGmICtLJMCs7
grg/PNOJGMBSUxxmV2uDs3qU9lWul94zpI9PFPK+1862M/+4WDwlkpRaTLhE+kkbTM8U7YDiPKvQ
+FEtpfPjtX54uBy2UB7uuIptkPtS+e+sxqBPJHdzf6ZFboy2PIAkN5tjNkiUC6Gpi0d3kWWLDsud
rZL364FSk88u5WPUUH13bsnn9gIbbw90enVl6Q8U5w+8KgZ+hFBqLR7JjQA8upXSmZn1VsXKxgvK
X69GADdapZqb1kyqWRHbq5yLHDlZtyNPZ6bBxCc/FSyMqpc/HeSZkJ0jVPxWT9Y+YNURfRWOKkCY
zyBIGioys2Xd5eDqJ3kUmh/7EiZhNHWTvvXkPYPcmijPDeXqzz2DaMyDxudt7rmToQ1G2gH1dQ3O
EF2jfKP5UrZMsI4CGetZNhFsKZ9c6CNXlAMf9o6D7NnElhNGoLVoEHYN3qakF5I03d/Y3Gej9FxU
sSi+OJ2Rd2BnuedT2kIsIy5OGbrseIyqhBBF1dHVfURnMip5X7gjm/Zbkdx1nT/n3P6ahtZO2SjR
R/2fkloFOp02/Haz6kpfh7l4Wday4znl0I9/4txlh3hcRHqK1NTjNP7qtFlLxG/JeY+hMwhqRDVe
PUoyPmZ3S+4SCdg3RMUr+aq57dVLtqVXLB2DG8Wf6df83LMDNwxDGKLq66pdiyl7iS4YeLRE94Rb
GMqAhuwIwH3L83402pm+jmqfLkDbNFl+crFuRZIRTo2Tuf6uywN5rI/GC35KEb4D2wnLBcnDO36C
5wjljeXRXUJbR6Uknoov93+Pfswa91/0x0FqcFF5SMwv4Gr1LlS9aKD3n2iLHxt/KFJOMcza0Lh1
fgBL1Mt0KmUkJ6XTAriathCJRTcWDjBGoVEwrlZwTu8a/rdQ1NELoQjBOsnXx2pnHiN1xielnXFf
mhqTBiuZ/PWIavv/p3fF/0sAARReHTGIdmmvZVvTpQ3PoqjHDe+MoCcAyOyNjvLvmKZTpOh3/EAx
XB8Dab3M4qCyeeReMRbqA+aR8j6TKOsUNC8NQJGIzZw3BVYFBrJZjHSDWlLbzJTYpTmrYDxnWou5
OovhrD5Dfd3lxtbeA0hbCbQeQg9cNRPijMJ8I8re1+Akhjpslzky4324OluvYt2CRZ4lTvQ9pz0j
uVY1RvP3uJ9mTQEWIn1CI9hhcIakIRnEcvn2KFtqtPZbGOa48ZqQSxv681TfuE42xSPw/XXKcib/
v06LxhvpLbpX2C0oLllxn6Nh7Hxg+ECabhLsrXI+crsQwaBay+OV2sctqGhppsTOS0Q+XWSQOBJ8
d2R0KcLHwEg2J8niWhMJkQMYXf4Qh0WTq97GdmailB/6SWmAJ17cyfKgo4ml5/tWY2EQXFB85dnE
gVDOLyqJyV3/cQzU+S4a7Sj9zBgZpofj0h37G7FVxyDwf6h91Ya1UXbCpkseDPyFHIlvTDziomtL
hSH/cu/RYueRUCOj2OIfSxbeW99h3golCsbABqu7g6aOk4cicBVdk2sUZU5VMoDACGWOmCcjXyGz
37IssLLVW4IKcNb2GAQY3yGow2CoNuWc/CjaVWnXGhotUc0omqbmuTUhK5+QkJgxcEIdiq+LInrr
01mQco7f4QV/rHso4nuY78r7oJsqxEcFHpQNxhF26h735/a276AVeRV5kxyVV3sgtNMnvzfbZmFF
pcYmBgMWxoukvXSko6ii3vCJ0bJ+CeDNSFrVK+g681zHZoeCttPqt6KN6urlcawbK9kk1UFf/wtq
nSr/9sndEt+c0O1nlktjg+hHoMumav8DPXYtmzZcgvoh/2rabez39aXDAzXxza4T/MqBxrNaxOpv
a+RQlx2fzkLC5iSo6dZo0QRZh2qHhvE/4iMcK/CIaYM8T6s+y39rt495XvTJ5kVTK6t2ZxJtc0b8
PElLnsr3oEWl6pFDnWzkiPCINlC1KiS8XH2pPwUdAbA5+zo3wi7RcPDjmERi8mPQYdvim5k++xpY
clyVr6NI39sLQqEdNoQ1TLZRcH7ZdTh7C2JXwtmXOwBBnawp0CnLi0UG0JypWBmEjE1iMU850Xac
UipHa6V39GMEO9C6G918WiYgxIsg2S4fdSVf7sF+Knib1fvWhnoxPOsN9DiwcIAgZ72hRPtkLjhb
y7YtmXU+SmND70LjeT2ueUaw9O2AH6sJ/QT+r5GYpOuRo7ylYrbs+I82pd0325+832BKoJVcBCAM
MdmLxG9kNL7OI8qS3sabawnfHmFwTKbX0P6ggd6wlleMvd+NhAMn33nc8AliTIeapaOBOK+aFuzG
JB79WfXnvQMxj6jaT9mmauurY+fFGDC8zjeyZNdWNruIpcVCxBa0cUERQ3tr+MItAPBhGM3J8dY9
tRGgf84M7JZG4RlzM9c1ebHLqWddQ59MPr7AFTIpGgNfHj2cqj35TBaRkEnowYr92h2nA3X/CeIr
TGZg60key0Cvx4wocSSsNxVzo4Fqm2JVkuBlX1X3DJCredQNpvVy0y2ZTeH2Xq0jYVByxgTdwu3u
gcOIeT0CdUGZhouM3jSBDQAxpJOcND7Yz/tt5gcf3kAU83xI5Exy88nhHHtQ3IrmAFRWIFEpQ1nk
R6G+zgiWYfsLdh6K2lZRAf5niBJD07xmQ7bKcrduEeRfLBpDAlhU9TRdJ4AOL43UnBYAoSS1eQsg
oJnTUzaUjXt204fBs3IuNYxl2UTtSEqbGyRV/4QlIjZjRov0zLgZjhGG3n5XkPeGtsTvaXCah+KD
KOnFZESlUwt6dcV9nyrt1dkIo52Z8qExgYdJlYdBdaxm4RW4symzgJjvGSSGOIa6v+ZrUBKzU54i
mTWapBmyN+U7nNIadP4nFPmKQNW4pO40CE/Sl6sp6jzAiC4ACQih8kJ+GS6iggzZ1hCV8cOi+FLa
MFveCNe4CK6ohBBchTFPzW6NfrA1XkH19Inz/lHqH80ElqxOSKW+HDFa5fc7qH5g2j1+iQLdCGII
5apOy6J5m3zFKDbii4DOg8h0qBPf7iEbxLasMfGqxEYnH3U099TROUOQDXlme0Wf8VJCVB6SopGq
mzA/G2nBFMTBc0qbyEckxnjHpLEPcUtQ7ee1I4Fen9dLKShE+AQIbs+PXjyLepE433TntfI9Fdan
Arf0qCabNFG8FYwx52XRqSr45/MVke1895BrMZ3rfhJhuZ60fnF+KQ8jTeTtKWz/swgSql4/Sho1
Klj7vFAlPXmoKMweptuRBzFI9OYUnHbTJac2jvzGoiakdxyLkdXaWnxHU+lSvJZawGI48xKk1hWb
G7udolYKEy6g+/QUeRkrN01nh74zjH5YPc1J/jDsjriAZqH43RcIExTQS+F/SE3Ep5H1tCeYjeWz
RCu5odM0hkGGQEbS5OjvWqYZBtlA2Q/sHl+R2nmgDEQ+r0SgzcebLqHEiKduWte3wqsaCYIcMNU0
mGg1/02dCQ4ED6lZ80DFx8MHY/S1iD8KiTkQ57N+qhHT+fdyBdCh5JoX1FIfQsIhYgkJmYg+GG8+
DHdaanXmICQwKqPqkEZUUUvLgvHHeFahS0gGJ+qdefULXooSFtPmfaenrsBuiMphgyLdSri0GBkJ
CpBJP6KIecCB39JIaMbjtcJdaoKKCN+vX3WbY0j2D+4uR/21iGiRAhoGDsosNY9ykZ58Lvr1tRnM
MDww248NjfPl9MfZuP5vLw32T1Kwuo9V3Pu20pEnqXNZdvLYno2iyIOR2BjTOkXcAacRF1GTkety
weClbfY8IVZBmW5YzqWgRJuayuays/NYzpDqFEbiSxYVREyUC08QCOfDfKDUa7SvzhegL4UlVxk2
DWCK6n8SQho7RgZGuSDMAkm/uIS0ePaKJQ9vjEqE7jd/K66bA69Yqm7pg9HPcisqZpjRIH2A3opa
PAqzZJKjWcvWACWeiWSw5gpS0Yv1QvZNkweyfRZEOW1IRaeVnzDiBsTdaRLtYFceFGK3Ict/Ewkr
Pd0mm3VQUQuSgyLo5Q+HASRrrDdacGvUf/2nwg5DgfcDBMzJSMQhOae8qKWyj+MIcKSFcCX4Sm5X
4gNxk4PbeLSzM4r2y6ZAJBks/sqn/K998gt0sA8M+bSKfGWHWsD0i9m9YnmPcdfknFPl2RIFnaTS
rsHMZWtTagraTP80/MHy7vnMxaStwckAW5WQ+44yoaNcqb7ta6/rTEkcoq6JwiEM9RmRv4bLYWGX
7I+8V+G0Hir3aZMPHqZdfLO8aG+BZp8dmcdeeIxIhyYcy2P7HDN+tZTqyZZLOt9ycG1WjiR8E4nO
lSFbb4D/pZjCXgKjS5oNZEWRiAsbXk4MSYdbhvU4AjUmJQt1pwELCT7v706b4y0xCX7YaRaqY6O/
A+3FFfD8jFlK470F6iNaHwcOrgtteXVMGsE6iUwa8eGINIXij7PIE+NMzs1+GyDlEzhq7PDPVLQB
a4wUUXq6fN4chqJyUSPnLUxWeeBG52KPiDdinNXZ2u29HqagDyD8T0Unp8wo0FSjiEmSVJDHUO+z
VrfEjcJ4Z9xvF5NkeRvCaQlVuytMzvYxuGcVHrPp3L2/lZfDircZWXcgofA6loACyu1+5ME0ZxAh
Uk0D8iVJeyHu3FkouMqQaPq0w/fHR2bYD6TVBt7GN3CNnTr6b/C4Ne+x9KX7IM9H7h9xZKxiOQUw
Y0UJLt63nnpX7jgQhEdrEjnE9Tk+cx4CcaHWTWK/SSiOxZOEmzduG0lwMGakK3cwKxThDCs+ENPj
EAr/slYugISZsrLJn/u+F4dhH8g18eMggjE0Q8IlYdDbsZSAgehOke+Kz70qnPjUXS9zExM4qDYx
/hPWCZSVx/E8JpkZZLVxKIh2exfSDKwwarAuPrTPzZO3PclmGBQdhAsCK7hYQqfDeQgOhUnjD/UM
h52MRuWM53OmCiyyDSkwWt7L+AroHavAmqMVc8U9Fwn0w6Luk6vIefJbGofjL00eM8kGmMD+S5cp
uZgYkCUsATiQM+2hxVxQNSzoHR4nccoDeRDaFS2Zx28tFSccgPHtFudMDTCwkVGIOaMxmgH49k79
iNSq4f4284ibxPbowwLiWT/YFA3R+pp+IfEkgUvk6SajmQaVSQcj9YUeYUVSPtpOMIT83xF0gA1X
vptQ7efuxifXSTVWYRDPMhPwBqwc+PZctJyL3lxXQo9EcPlae3Luig3YKRUSB6GjgMzGFTsLbK/v
sUfrn4WzFe4PrUwenRxELUHk6TzGHEpJat1YW7UO0fgwiGC6JJKs/Km18uozfvd51wcPyG4iiWQH
vZO2NaYxbNile/T3d+lDknnwWHMYEJIQk4qxRpeArFZR2fFxvucyOg1LIzts0NWiuA4mCr7rYqIp
gZii0KNEYelJH05V3lzEVeusO2a2l+VIj1Rx2WfSSOEDefOH6fKaLOit1J/H4Op+HhE1y2G0V34R
gdGIylTzVirvWVfxGSPfEELSZtOX7CsVrLbspBZ24rn+tc4DdVcUDzsQLowEQUBQPFz0WZbovvgM
w8MEgw+AC55UCJkp8+Iel6v96xRzkLHosuDoSP67nNFVXY0S4IkOvOsezg9SxHNSZfRnNNq11pi8
qiWQIZU9X2Y93vz2VXvzABXP09kylZi3QaFwlUMymEaZ6R8tKr54irMyEIki81MgjvL4C3DanwnB
GjqVs50ixnWcUd+A6X4zgp06bLhZtiMQyMU30mxSyaK8Xyvig7sCMxEmcBH4mbY6RyO+Iauqp4Hi
GQVaLLRIQtHcraH/XdN2VMhOKHSST8iWmFSuVL8FEQvZkT4WxL0tWHb0kgPNJ7vQlVGZvmOo6AGa
oH8lQ+HuF+hTJNm/UKlW8sfhsWSwgsa9i91TRr5Zdarj/vsBMuo64rYM70WWg01BTflCezaSf6KU
qdMYZI3mPpkFWPQXlek4wsncfu3o5kQGtlFbFg4rECCOsPR9PgnLYL6KfZAKDcI7e22DNtu4WiUF
QoOVvfrwlxPx9d5liN5xeLqbw77lpCgU/ujdvXSQ55spMWF1fnV2UG6LS1FPXldGPVveYPvmL0LI
e2K1mNttEYKhClMlIAS5hEJqvpi+scojhbYNlNC9hOv5g4NTk3fMgDMVZZIktRQMy68qcs2cTjRE
TKnN+L6GBC1TcE8ftYrcgWLRfOz4fr8imhwIKGslZuFjX3XHYIXyrCtoOKj/+lm+JZhGeHKLNMRH
wK20z/tG7d5ThOPlqYeJWqImdCybIXXRiCWdSTk7scgqG3Z0JW2FuS1UERFCmbRIbhXV6RA4RHbu
w5mUb0Jhq+Q1fqYaV+vEi2yCevSBwirHymYcllOYmOdI/mmrQnRKKJylC+/JJUml7SQrRhL8xU4R
lvY1I+9bKQJd2E5jcnOklIB3fw/sEQYbNfS8o1ZhV5sY1c6OWY4iDqCE1HlQyxF7QZi9qhCDhCLf
pV4HEMpt0YaHuY+K6t0Sc2vU+RkLbcXUoXPE6oyv5DRxghQs5pBihx/q/uzqlWzAfAZ2n1nlLqab
FcSsPCiw7NVlCotBZSLZi7tB2woEyxq7eS3vWgRf8w32Eg0QZ5DgFfsscgwKGlpP1USptUGwhbdZ
mMqkuciwmgJxNSBy309IsFZNF8pEndMUCpSZVnhhSAfZ5H/eldP+LrJjhRHwtrpXU2QgE2Eadb+k
dyBrYTsy70I2shd1DF/2QsK/fUErdqeP776OfREA9495jydJ+dDfE9HqTtznb9TcRUewmE+FZABb
Pbrxn59CX6lN4/9CdQe3FkVVk5Cto4ZNxbnKb3TJgYCgOdZ6nCERPKU3/537tdCDhBTbpcWTVFq0
0rRSmf2T1us+cIBRr/9mqr/bNv97L5h+w8XxQotcsmp0vTgrV3uEvdCzr0lFgaQfw1MHSZ8bnZIo
9sgmi+2MhVJ62ZKbejH/Vfhz2ggLpi6BleAZnsUgelLjPIzPZ70VvGPohZgh2z6BrWywv3HdEZCe
xYyUwj+xjdCBB7PsGCAzvmX5vkLw8m0jplF6MDuuQGlYvWFNak+RR4kOft2j2z2/MQFFNzKDNqbU
oQwB6XOR7BZ7bNFCV/esesa+xxL2R5ecAM41cHn8w4klrJMNJXdXRUyeVKLDlx3VJ/8wXESGL/dO
oFEKIFZxF2LnvsVOvm/1xdnDvJ1hO9T8abYNO54QcYcfr8UqE4MYQkx88+BQI9GBeDQkuK/f3jAo
qZq1ozJFACENVOf1ixt67zT/jgNpgIyuX7BDdG8nzaBhRqayGjezdP7tx7EMtG4Gw5xvLSa3iTf/
HiEvJon4iydsXmC2nSG7UBG1niRYPzEB76ZPg3h9HbcQHLrSNP1VnktdBGK8WpAq67jKdcNuAN9j
soIVAyMG9bjRW4oaNX/8MYUDWf1wBFUwWi9j9vf47GdFqp9UnL7w5uVLjv7uXIU3yeBvDWM/Aixh
LRjvxVmZF18e+moyYOx4uJ3f2vc2zpRXnj+UoWzEzRXSeCets49/DDJtqA78Bis2Paw7tQUyeLn7
Vp2IBbV/rnBzNARN8fZulVy3JVVaE/5RdWq5SrAuCc+TBYmP/hVaHlivQYUfNKMdbR0caPyJtkvS
/u99gVPygGtUmSCJyUyEiRUagL9rQM6QSVY8jvza/J8rmP911pmduysA1RRj1J4hwXpO2Q22Ahto
X1oEcfJ/PxqLJajdQEJomL9ayDDQ2J4dflN/PeMRBBxtaz8JyNp2x8Bff5T8KwYMbCFabMDzg9z6
RaoremsnyRX3y3DU5r1QNWpXi8Sn+2GExf8m6hOm1R7UhmlmeFHPvYcrO/eatpiz0mNVd1JG6JDe
/W7uuel5sxQ4/3QJ7Rphly4iXbs2S9DjluEUYxgxBvFCVZo8h6PCFlR5mmZi739xLNleziXTD/OJ
dknD3y71BaBSBCXUizw51QLf7X6KyN483y3ngOX5DeGUWMUAVlxpgsUcUYi9Lf7WrvNo7C2DDvlo
x4bYhyA685/5qbSvD0up8HrS80dEyiUQtpTJs9CrTX94/nY3InV1a5v9kppYTO7SDXPYLaxTAlhE
6MoROPltonyvr+11Hwnhk8ReEQFDNgFTq1XUImu/KBvdRM7+TVCfsPhTq//u76HlnhGazboy3gfa
mYHpdT5naKVdMxhk7bs85U452h6nI0wflkQqifKp1gcHse3fq0upf346NUtdPYQZP4mfs2TP0qDy
TBIfYcfVCphl9Fpb9tzcd3po7vKP35jqMA7zqTPjJlbRQvzavO28tHFSPtkgnQw9qNfKYKzJjwN8
qM4EYHZGQJ+5mY9OmZEydt2MLdcaST8NCVHiVWSQgORtvvJaU4S+wAMwgW0Lzelm/Vhx68JFRMUE
bX12YV+HADTemwZttHPXhU9bijZzXQzvF0J9MFw1+fHRP3lrGcEPY/yW1E6UbC4irMuQreIHOu18
vc1bDTFkafW82ulF7l3SkwUYMBNH/S8fmSX4IjQIGsXx1PoSZi4GvKiUayvA7UkTIMUn5Dg8+B1s
UO8SP1Jo+38vaISR54YcgxoFRBYT/4B6n37eHa5yDbuuEE2h8n+hAd3wM90TiVMshX8eHdS/YQm+
tjSKQ6MpeKM+FmmDilVZ18kOdJd/cRhFGq3hCY7Uc5IhdJMP2QOZRTQ/IFzvao+ZIulHF3iCeMVA
WIeiivQ1iiFukTtv4AZp9xcQ3aqqvEWzmFciVdX1YGVLE8o5xPUlq9VfKJNy3gtMLtZh2fVsoJFE
gkpM8MSz1wLT5umanhPruamrDCknvx9PZF/9rUpzIlkgoEb82sF6m8LgVLQ6Y+2t4lILxP0Pg1z/
ZOCyf6DLRE7yBuJVklY0EDGuuw5nsLZHmbvUwXc2FBTyUORFXF4CxQsjblpYDY9J2Z+ujpfYt9aK
MWIDKblQC9LL5t5Ktx3ayedz1O0LTMpHKQUJ7lSsWJakUfuUjcbAvEdbdxd2aQ30m/SUcAFwgQPL
sDq2IE4IeQu5usTPjj8gVgRh/zavF4N+FRUBMxfi1mscEWJs2ZWq/4q9IW0k+/24Xa/lTan9djRF
cjFD1lzyOozk1wcXchDabjHBNXtBSx9n6YN5F/zCXy+aGPpkEl1IR7P+2+G8WxHrVpCGYvYUEEJU
AmJkW3FqcazKjTbQG4tlyWoJ0Ck6c2pHsCHJ8+Tm8hDg/C5JGoipOQiGRgh6/mIvarihpcMxtcDZ
d4vMt6i/jVGh0QyOPLGRcBPbRf7kPCi0YwelTldvVpNXOD9yigbuLygpcitcEHzqNxKIWemhMEFM
Gi5NnYP1HGM1HIbnzRxIUD4xCflY0l11zarlO6rp/LsPynPilhta1njnvcJ5m6oVTmkVz6FXRkm+
1vjs9p1RuO18tR4RWj531Evhet9opUcrPzeReeQY65bQfKY7JlyD6rlhYI35nd9ioo+vve/CnbLW
MacrnlPvF8a2OPPF3WN1jvB0le6dxlkv+3hwvnTLofZPOSVD0kTb3eIaP8c+Jkqph7QAfyVxsmO/
+YTm6Zne7Bk+QYtwKp1R1m+exriqenVbbOvt4mEHDUNYZc938sVTr9KM/c28u+nuB+xcIZ539h+Q
8mj9sXE2svEpu3RK+4cOsqZwSQyt3731pbZxrSqLosAVWvqc4ju9sHCDEpxutNY5vRSgNUJa+vM1
rJVjlGGBFvfb8G8nEdLr9HTQlFWlZeU1+aTNxVIZsLc8boUx4GaSnSRi0/6z62vhKNbNhQTrCv2v
IFDjnqDb0SjNz7BoOukrDAQfgTrtsmthQI9fNG/YQOcCbA5bClvk2D5LdJZpScQmKduF3Lfk9ifB
XxiXYuqxq8KuJh7bSIYbHT0GK0E2Fgo1HMf4vINSAugtFUwoAKmTxbKkqzgFzS5NOT1/6SjGyru6
T7UnxWtBgZJPWJOxupEmvSDGI9floyLXbqGUemitlYYs9bgmljwiZXenkEgyCWry2NYFKJGKkNz5
n5DsILBNAXj5Wv7Jb7BZt4Ph/ObrX7ZnvfQhrLMGk5LY7hfx4gr31OphDRegcPuL054IrOZfoWFS
Pf6goxODYqoB8nzoW+peoO4UxCQWR3wrR1woYtm8bJ/lnuBHv0ibvSzDcoFKR0hT/7BXsikYxKos
ykF3CDYNu9F/EECVhpxdNEV+ZytDHFXTzN5w31zZSyehZ/RAf6xG2F4Qxu+CfOeas+xVvPm2iQtn
dfzO73hSqigkvScbq7ZTM2XJBcbNJsXZj+rPCaVNtRENbmZ0Ks53Ffm9cw+UeRF5D9V4xkqO2svk
Kq/ADLEoN3oVxBYVvCMvjzmiBXsxbgf3rX67CGLRYf+0t98zs1B8G4TmKhMfytYoekThOfX2dB32
9yTeWdW1+tzskEopsk1pes0PUTU9ojuhjNmIpUcM1xPtE8/gao84rHLmesFn/CfPPf99FEmiJoR3
8HOiszGvbgLgjiiMu0g8F0A2BTtcBFWDLTxaVArLbFAOeUuMazZTXZ8K6RbcQizPmahYL4il7DNK
Jk+Kr7pe8SqsctFuBBSKYpv/ezEFMoiq/fEKdXTUlNxhho00tCKQThq+MuWuRTKGoJbRnMVXeolz
Rk/qLDIaB0YEhlV/xjaxg9dXSy4fyZSOZLRbLFTC1VWdpC5ICPHjtCNPILEboke4y3qoiEARnVaW
MFwRGpmCNHvlBpsOHdS69u5nQ3sIIFHCZvsAXK8kPLsYTv47AbZW6N3M5IwzWxxf8lFarjD1r/ME
Ef9yd2uNM6lnfynziMNwYgh4Lyo20+ILPK6btFS8o3rFQWOkK/fZLkHDeZldb8A6aWhwLnztp+If
Uq5fq4mF0BGSEPD3sZVIsm+y5X6ZM+7NEcvpga+epZBTVHFOmqWNPbCq2qY8AJrWTctNWX1Fup+M
AYjaaS2TOw2WLm8zrGuW5SP9BLuxwFLNDAAbAp/idY3otudRIzbO0oulLIfdFGGrVQ2vFOwm+95C
/OJiQhz/MpTt+ydJM5pHMT4Dm1K9rQyydb7vFFiWZEjg9wkUxppKyL+wMfzo2Toq/u5tc7m8166Y
HwRj+yymSZq1Gfif83evbFVSPwQTNBTxMptF4MvYbqSX2yYrbFv0BBMNBhRDjMnW06bvkcPprFhQ
XKAf613lDetkDG1VrJL23oUwEfvhDCwYZ30oW4h5FRtZH8SLFxnCSYH8S/JwCd7yUVsJanIAD0Vi
0foqGPszR+ifSm/GLhxA7e8tPgHwoDk15UO2AN1+3rCKB+Pr4+xzGSsmUcq8ZIesEQTbJIaTFt/A
jPmy+znajQrK7n1lStnMYx3UkUX/iJor+oUPcgqs9lmUOzcxCYXyMENU1JJyPMEpi6PNXsTmggDp
oxJO/tV/bzA+Hxev7bs0zgGhhKnyQLHzbN2aLF2PNCBemLv9eAcRxEDT+t9mjP6QIZCJi1ZMq9MG
aIPR1DiV74x0XIssaJOd/wYGHo26Juf5F0mjv7YyyysNkFlofzfTU1uYdHvQO7pB+V5rPiXwUiWX
lXRLfiMspS8crsrIMrK3jyv3gQSktJwlpRklJsZhJe6TFi1Ibc1C+lRAEhtndaAey6xQFWXz5wy+
t3nUg3N38eQ1vRfP3UO9aM5ccM46UuucapTGspnBP5QnkcwdSXxUt6PO4+qZlrlNVvWucOltY5xi
p1Qji+GEIEdPmtBwcb1JPAT98gDownkiWs0jkJyrCsAYvZLZ6adVbtwOzaS9zd+UaDETgASqqlqm
f6VIkc00sx/cK/iACEcKFtVvXSSQWXGH0ueN0vD1oBh9PrenQzME7pjGzMwNZlgcMHpHXaa5Z7yC
XgGMM1n7rweBLGMHPbxl2j5Yl2ZSD7mOeCQnLp3YTUMO3R8793LqN6cvCzDYDTs99DgRob16Wv9r
q0FsKPuDQBRfkLc758DLDYHO2lHlPdBohGRiaN7rEsiy6hmVFg/H3JHx3BDmIJY+77/2hpxleGRH
IGoUr31BeKoxVOL/S6hRRQdxMvYRxFzeTZkr/pBU5LutyMhRuUDzxiI5NdNx9Ih18SHZ51ey0SU+
dEbrCB9j7zFFYHyB2RuLnMVbJ6JOs3RMGrlmLVCRI8PA8QO5sMBBiBCJEMbnzINwmjX/CHtT6yRD
BFjyX4O0qCv1WFfg3agKTXd8W5NiX7Tn/rlBWINWvWQu3w1943ASiIo+/7kmqh++Ayj8Y4HHecv/
1ajzfsa31Zq/csc10nyHRQzDIiokoSMYFCb/LM8Wr14n7j1CoCLfm/s/65RMy+PJgyZ26xWV+twl
aE9HYU5tvBotbIsUlctma9tvX7GTv7OYgD/ArQRhhRrFSlLGZwaf2Qs+OTBfJ7OqxeU5EjsUcLl4
gKIVO0rRcgztWWk8MEOgTLWjYOicy31T6t9/eJv4iHPz28YmQysGWOHBTIRrDg3a26U/Ry9rSGZs
F1yXKzW7Y9N+K3xne69bjNozzDUdOCtauOmscq6vlXBPL32pdSpm9o5EinXaVbyrq5941OSLpNUK
brdQ+H/B6Xfyxz+fPxOfSOR5GdajkqX159mMMuJBj9ccUITpZBQrzKI33A4infIg3XOjXYM0bTtk
angkQ/N9wT5fdK4ps7wVSm1b5KN6/tw7u7bCEm+B9+sEe6VHeHk+icsyf4ynfZr3NGGZt0PTsuef
oEQ+oOzN9mvvi38ILFjPgZukE5erHoRCZlQxqYU1zfnr9B+1ovv1P8CWtp5shh0oH+fFuo9G3Ve7
WC7W4lHMUsLjociaci0stOcCp3tUKa/La8ow5O3IK1NiLZKeEzRjjp8ravD6GU2O2g1RbLRmrLkB
MxfuKzoAvBw0RLPdKmno8q9WWc+GAuL10rI/sw/egPFFvVFA9jxlA5sRWy2iFcGby/aRnRUZ8cZN
opl/lGL1nJ29tHnpoEw7BW9G7QpZQqqeVvkmzkY2zhU1itZ7QVJcCRkZPHw1oDIopUtQhJDfbQnw
6M309a8up0gA9en8qfXNTrTm10ayb/+uG4BiWTVifa4hQshS1IMKKykt5Yo1MaITcbqzaKlqrtqz
/A2J4RB6VXaKYZIw0YNAb4OJe94lp9tu0lCLU87mx5I/GuzRe1ndlQVZOv7IjH0FOJX2DDk5B5b1
F8pqk5i8aUGbOPL6tTpzs1wsGTJjF6v3wwgU+7Yy9V2QMQ1IgXfoDElYVA6eiD8Knq5pmAB57/qG
3dlvTvQ1NZX0y56ZAR64J+NFDliBJykyTARMTGisbvI3Xod6rVrhfx+Z6eDFC9BdOlWhmPzxNh59
ckVLu8K/N8X1cjqRjU6/Dwn8DxagzkW1BJbp1S+vmGWdxbSdsiLgthVXahbacBQ3vC98CltkX8ol
nO5vC/BJwJrUOcQT7vUTY88I/Nokz8eW2RsuqTFBlI0dBlKxstWYSjbc2euZTrTMsFbHfzSCfaG3
bODLBui91I16lFk73ADLYjji8iXCspntlttN8LWsrOfyUF0u9wbhDt+trmaVfaDOIlcseCWwXFO4
8ujm+YMXd4+EhxB2X3qGQVWpj8d52/pKFEljRa9Sn2Xv5Nh5L30eP2aY0wyNRKr7/jGjTU4lKitN
4nIbSWpZjrAZmWBtVo8X3z7OU+fhqYavpS8b94AY/EZoJmtLTX9SgdFTufh2lCVQG7OC/ldZpFTP
6l28qr8JerMOk+ITN6iRGbrS4kf2hh2mW4aPt6gxdUTOAp4EHuiC9QH1cD/TLPykjG+kQmGcj4He
IhIfOor3c4ViW+UXFfvVbsF9Ej4Im06mCe9laEqVJ43ytgo+u1KPH5rVCwU0V2Gb77rrIg+zOFCe
pB9roggAVVEBNd7Lqe9Ij8rttIi+lP9yssahTWJ/pOBsgEb6mP8wcWR3Tq+1aO9CPdpmi/eVq8dT
X8y440CRFhbZWJOb5BdoVQ0aXJyuvxb30F8P+bHKsn4cPXY1LARNoO3P6SzkER6tjH7yowv9iihm
IEVk2U8o1N6qLLH3rCjXWnamBqejJnvxdJC9rYlDLz2Qcngmn2xifXCOjR5lJbmjEHUw/HNYL41T
dt5mRB2HaJ306DfdweLc0vBv3WI2aBkK/j5X6JG+0UqEdXxbzVz35PmErxiR0dZYleJelu8UquOA
Sc6YLW/KGqqvhLaPlShihtkILijUmKw9NvDRCreX1MQVNopL6BQZfTi04YvAVEYmrITQwnuRdgRU
X/Qo9WdnObZMf8FqrkpWT4QvbwKDRHWPTvTzbJAmYf4GwYcE5gAseKZ7weJ6aztOpPvWXO6DeIbY
zyjaTWfQzFIwViTJueOH5RFejD9U6Q8hHXY9fjGbjESVMMEMQ7NH6pCWpEjzEb6tiUt9YqonCPTp
sIq9JW2NAJFOLtz9KhFc4NiW8FlD7tWQRFTb3flrqUhj26MNDBmjIHhdkXKZMl46tzdcQsgLo2nq
fOt89ZXJvrUVFtW/S6pLh4BixGdm1v/9nL8FhM9+xSOQlFZEmmRo6Oidx/uDv+90xFVGOHkb6gme
EkctBadeO/s59D5op66JxwyTgq66entVQl0RVXSMY3RP8jbXRZzSG7f8q105R8gO3bp91G7flF/x
DApxAPT3LxfRsFpbYVUtNjRjBqx2USdtjBVb6oBEEMqmieShoMGG7UQ1mFznQvrUWrfb2Ik+c4cn
SXwkR2FPHlLHo1BjEq0QR6hdJlPx+2/uFtR5GPyXDSugvYVnF3U17/b6zfe16tGuN2h2bzly2lXn
eeMVyArfJYlV8bbtjKpcXdd/YEhXmeOp2aa6stLEoea3KbmzbgxX5fMD7EpSZYCSaFVjKvX8vlAf
g08/7YDP3O7i3FAndwxARtT7Zbi/m1v3CkBJlJr3CfVE9trja5zO0G8O6Dk0R3BvQw39tjjFQn78
MZ51kY2rnWrLuP5c4/bDB0EuJ2WINaQ8WvZG6Ab2egzlpytRr1b39OvvxgTHoqtiCkgiKPqkT2Gx
RZ1nEWNxcC4PofJR6X7OiYuDf9UbBUI4atSkSMZrRdbRWEft6qjuTbOxGj/kakLBeAbaJcjGcAnU
uxD859HOj1ZK3NXrEpuPdd62TVLSBNo8xzL7/ONkc8UKbeNOhZf4g0VGsW8frdkBeuBno6DNpDwX
r03d6t9EIak+cop9Agfy+7jwXz7Xc2G0VvoHgm8If1jGTQ1qLVBAAcnqqDMmt5NOhbQPA26V3r6r
K+aP7fEWYYy19uStZoEOm9/3X2r+7Kjb4EFTUTLNtJeTefTbxGlic8sRkR1kwdceOJw0fUyyt5P4
lDInmoFUadmf4mx/BGXr0Z4mX+TjbZfl/H/npLpkLgUAkz4kP6zXJ59M6d7syQ5X27ngchawRXcV
6xcUuYXE46g40//YBl2qSGdkdyEY6dyE5iZ/PM5uRa1LkC95s5l8lpp4eF7UFDZCdau59KtYxh/K
6XyrLZV1Qhelxw7wvau6lrQRfaQOLGA5M5qZ6BFQOGcIzzQKIw1ULKzerWl5p4CkTMMwVZyRP27l
shDAikJswQf9JJRlIK/9IfmXpheBlv/MxbqkEIVS/dMRltNcgbLdVLvky+aa1xbYPFmR+WM8REr7
aO/faXmPHzfmGp7zDExmU+rhYIJ9V7FN8/dDdMG4HKrka4h3rX/kmm/feWeh3nfkfOA8ErDmlFYm
vj1b1Swbs52uJ/Ehy5jLh6l9COTJCQQm76d4scFgVCWM7hkTNbUUDIwuu5dY6J/gJPAQ9hHOF2AE
OrngM+RfvtHuV+nvJ276yhA3nrVckZSrkAtwWvdyy+wu7EK4hNdDw9dIjck5dF99PJr9ToO8int8
m1lyRxLyr0gt7BGhCx/D3R8466b998ge9fI3Qo8JpOTudD9cLoS+R2UL9mTAL0nIJlpX3essQ5Yw
Meamy7XLiJbJKcsm6dAek4F1Z/JCX77uasTqCpNnzUnH1UWbwhw81X/E7RRGveTltqLPyBTZ8vT1
fx0rZyQ5KWAguQldUqUA31nZhbmS0p7gsqbeVOWq+YOGuh9zkF1ayfovwClcBmjm1aF+AONL5zU6
fsLcR4P/FnOQwHRS/uLz31FdFeiS8cdDS/nD2rILTKC4TYxSAgHC29SU2dWoWVfTVztDRuOsFbBM
uLyMoIKM6xcfIWnnU9iLqK6d27xRhWeVOZfZ2HA28yEFuLJJKRXKlpq4rE5dvP9DGZWLd+DAqmKR
Vs7OryfBenmFqnhVKZNX9gE0FAGmJ6mbLWxkVKh3CjcrCCAPWedonGGk/XLnI+w+1UFFt5Fft+Q4
y33KazZY9tNB1r3YSL/F32cPCIV/WmVQjHCpbFZqWUAzxqcv3nXMgrpMmUBx1fqMsGgSGqY4wMDQ
SDos83k4tR40rslclpy1MhD3b7lLxnknvho/3Ioj3h9aSzdzdvcBBlO9H3gqavvGYg1l7UEJhZaj
D+be+z1Es8L1OUkIWxbT7amw9Myl8pLDmOdXqvG8Y5jHf+TQYMwohvtGpNX0sWmKbkFg1D1uV/Ys
mA+wftF+aja9KsKlOfQqjUrlSbQ0LDvKXYDHt/+WeaErK4xR1x1FxSLCPV6OOvAl4X7lf3xrAuXP
/5jxMRi3t/h3AVDXe45GkMRZkunbgo1EMK91xyaQKcJ8LPSsX/r803CEJ+m23SEc5y3rTnILqEi9
KFI5MqYCYFi7vGDW52N8Vey6Zui+iYCvJcJhSuhxu6VWXYHj9hCRmCsdp0JQrkGMZMsJ+TYBkNyS
iKyiAHmLWb72z/c2mk/7O99fZGKK9Pvl0pa5uAtwjdxjSQCFyIgXiICxDzKdhwzE+yDcnciKlG61
Ui/xS6mk+53kXsiaJzh9aXhfWkRPmRU0d4agHAtPyPqt8NlpwVTQGpew3FDoeTVLK4ncZ1OGZyC8
Dxfgjxk+vkxBmqmlrZKMTJK4WJFBND6d/WRmpefwh8GelFUuN+d9xnZgtBK23zSa0k7gPDzlW6uc
WVsap38bzqeNYIbsCGZBsH5WqZmbTNhoOft+vj43RcipsOBJEMN/gVicAZ3ueZ0nBe5yhnqVkdmm
SopqL9ChN7ZIRiPqN4LEOHJ1cnxk7kRBrAwtoYm2gk6zKEkT8/cvK8GRQKI43kbXNQ4dEdBNy05m
kvd0oGv07VOfofArv/XbF3Qba1g8MbcYqvzJeWRMWPI6BQysEAniuBfB0U3Kc6tkOh8lESkRhgjF
bCp1ITsKjcpwjlUdIVaIt7vist9SdOkAxvJ2WixEWZSxhkj46Wv/CL0C7uxBnVZ4j5fABGLUz/dP
mHM4cuYiFiEJfegK8ViukZ87ux8xs638U/w+X5tsb4mg5KOsy7d4yfjhvfD3Hs/Fyv00VIcJc0Hw
bcdsPsVJl1Tm7xZ8SDl78Tebbe7dxFacunQTs5HKeWZfJ/v3p9GbOn9hfe5WnpM6BjIPgOE3Glh2
bqvW8GCkzfXjiiWKxQMktNsDwFzO5SFpbLsQFFg8FHTMbVJ95ddwo9aKrg5FBFBF7EuShlfX2nTG
/3yIxKmYYQkFcGtXTjfXqp2sIygsNnxWHtbad06llxlc7ba1WYvyGBX9kB1vYtCHeA/kjZeuc/sz
tS9/8PQRQqStY+lTQzpEf0HXoljkt6+l+unStj6abQJNVPX0EkRn/gSogsk5G4OS3atRua/prKlN
Y67wDHg5J5Vybn1Fj571AluMlFQGr+4KuBJXuNekBPepy7srgwx/MfBgADwCLp2jwz8NnPLFMspD
S/ngTeoU6J8lxRvCx7t04KOeNm8vrHIlqI2337OeCK0BD7aTUL2/3MZbE8PgCnGXiBqn9ZHGv+Lw
nHkiPJ061+lui0tgvuOrwlcA5kWmgZLGpTPsRIxGhMB9YtIKLCy1pLMFlaxBVk536g/pfrivEgkb
eurIFlLA2BVggw/D3D9AqdebeJ7bSwJKwatPZQspYg/py8N/OSTjO160TImQmAEG4ZK+Wj3WXtjA
XJ4kR+gF/CTsNwjpE0BmbQfrbediP5O+el55nXmv/BY9bHwT7kCnrGM+Mvs3UnCFC+j6YZ0hJ0pI
921mpKKCRg4dacQ6E2egROvMR6bzro25HzN0oXVqtvT8SJvy+5vBq34ULcHiZndW8Zcnks5i6XBL
odZDY8fSfHGmXC7I3i15WtFW4or+Ts7GCT9r2+V9FbFwbm+1PGi7b1tjZuEnn148bAYr8DETMQf0
pKx+PWCwYtv1cfX3HAqIGZaTcgSpnSSAFSLTI18qdAI1X6Y/PStvMclTmvBvcpqwFBbz9vQXGgz2
qGsy/HLQtqAzvHKH4jhv9nrmid+VaML5KqmcNCnWw9cFKrH/wttVwttaSH6nJMmFxZWRuF5CTt5o
zFHZIl9kNafatkE9auRaDdk8x6/xOFIl6q2gkveVPcA0Wh8bp/BosN6noz98D06eSytE99ecg8D8
fyjNHKPhrNNQDzrC+xb7eo2himEzbYcwvHMGNJo+Vm9k2JDzItx3CGxamz3ZGyki113ObO6yhdQq
PkaiP6DuRKj0LUOyY9vNO8pd+KONNfzGpBrpQiCvVUDegXIhAXqJkxWpeSL0msazxXhmQ8QVqLw4
GcTvbxgQTedsolpnWgZuEtG7KPbMV+65QqYsVIt87jULVOTt0wP9vBix+Ire0njZcALErwVAxcid
YfjglGOmPxb7XOOyJZlmR6fbj1/L6XV1X4sFF4wSKhuWLPF2I3aO5BqimvvOoi42ENZQr9NMmK6C
3yTi2D5548Mmwrsykwepo8ggDLgECzsap2nCVAIcN3MG1x6IVm7VNSdlqjICgmCEzPuW3vPlWFAf
BaD4CXclkXfVhWcr5+CMLwJyg1OohLBizunb7TdA4WTpQlFMk8yTqOyPAHsx7eXh93z3mO0QxtrL
HrFCq0/pJKzG2A63KlFSKFtTexnI6ItiFZrukQvTYjYYDH/JD9zZMo1fLoFn7wJU3j6I/qWHLpHk
8ntK5cqSsLJnQQ2QFSreRJo9GY6dbKoHSkk2aMLTWF8WK+Uq4kmtfYKiZKqWWeLwUKtphIIPEgLu
X4olrHzSPiZhTp0Rgce+CmY1ZbY2dmPVijFEEUa3GF0ehab6Hk1BF6ipH4//DDG3K99WT52YQtfQ
5PnLNn41eHt/frcRe/hvpH8dd5U7Kax0AyqQUA8sLLZx73LJOQDiCmdLQ/rPpQUMT9/N9Oq+d1q1
YzVjZ6DjojCwsV2X1pYclkIbFIzjNgoID+WKMpFiSnKwGAUUfwyRgNIonrCLUFVQmO5p7Ivt/17x
4DpWdzUSoKKq+URZ5zfy5k/YTPYYfbiqSMsJnNKKVn8Y2hT1HGlsQBog2isrFAM9uTEPhOINxIlb
vP/s9ESaTPS3xUpfvXI8Lxsa6hv3CJn2vuhu/AAQaB3PPh/qDTAhbytSL658113OFF8Jq+/VaMgR
FeueOEiBhGDvfK0LOJ1zeN8rY14GrewFNSlBZTU/phu9W7SI2C+shxpctay4gKA4sFfu1uMxrWb6
OShhE1boXGk4BLhfi69N+OlwhhKtzSuZxWpS1Kr0BhPR+S4sNIf6prk5z9A/JOp0k37bJAnlbFCY
+pOA1bWyiNjxMCX7g/jAHBUcQ0MpOH2L0jC94ttyjvBFtDulm3l4MoKpblTrSzwxJs73js/iGMC/
vmHjSJiqIw/1df08bs0v8/6P057ptKVICZEqzTpbeInPa2mCWIjA1y2/JN9rUGR9Nqc4UofyxtH8
XoFXnedw+/dbmS5p4npNm6p4IF8WYoWf9PjhVZwbWfkG0ZqnLgxO0dsTr2vJv0HVboKmheR9Gb/m
yvoQjHPd4Vn0/a3A+INP8GP14m07Z6oLe5b0KF9bLPxx5LwS/M5CI5fj8NbiwiPxpmsSOb2NYSQn
MUsNutt8Qcjodvz50QxWJwKhAZ51z/e70IoUsHXJ0NRYVXFOBdEuUZY151cBq1Hn5mj0oEs58AOF
SHWHaPGlP9wF2g1Sm5HLHMqoAAk/dZbqINDrTnwBvggQkqsR7dT2IXuJHz16qRPvARtrxt4tNoud
omfHdZJTGhAWy7xI5ULlRhYMXQstS+8nO0dndJYghc8vLCg1EtaDccx0FflFwj+7r2SdsqIEaEPf
Q9d6RzlOsqH3xxkw6gpfawr1b9VRW/lOTHQFApPTqw2nt8qdmwHJSi7tzlLNbnhuvTcUcSxdIYAK
wl6YZ6LcsktHPA1gjMqb0Of/j18OU3ON/n6QaVtFKj7mUlmeF/XsAEbqR+66jqsMe5llev7i1HR1
buHQxI6KTWRSSMfHKLkTt4iv4jkSpNMJhFc+AmM1SubBYPkKvSyjioNYJyonxenU08AhTAd8hFaF
7gJ01kR+T31cC+yRmtzw/YZJ8BiWDBbAPEiXaYnwrgN5YHdANb9EtBXMDYr+sB/mH8z1T3qr8bKV
gCKQAHNoAIwenVeKhEE9D4ZI+WJFiFTYjmUEkcLQ2rVW5MY/VNVlDW8aIL6PobczmGm+3lLcTpOg
Wd3HAw8mWNW2gDGf2YIfLxRRQ1Z8rRrmt0fJuJ4geboST/cmpRWQurM/rtTmFXSYH1DShB+8Dv60
5mlg6M8zvnBpGJzM2/KkDA44Op8HMsDXee7xVbLgcDsdqmjdoKsK80ruJx0GstJ0SYEK7rU1iMjG
fyD7nGN4sO+aTfnGJlIGQC/k56Ay879zzADFTtiylcAxOSKl+BPP3JAPFjzLa1ZohEuQgUr9pLhL
FJiqrPLu0w1zdlmy00ErPE/pl9XY3lh7SOv+crlMEOtpPgFH6LOk8HOq0orfldfAGE6bvqJmCfYr
cHT1V+kOnDMtIQqAkBYZH8Qq2NJlwfq/jA2nrfTv4WAk7koq6l1TptGh7VoFsVb8SA/0njDHHNSy
OWq+qHprBVlpFTtWxcl0imzDIRvcjFCizCi1yZb1jDNQEtm80Iwa907IjkRIfbAePZ3cTq2hdZWp
JXIhmNcfbg6REMX0GJWzvpuIAUXjWvrcjRFktldTsUzSCSUp2gy9MkxLURxwkZQMS/aO63w0eiUQ
xKhQLA/Nq9hvrmxLwHMY8LqKD91jJTlhk19DTi8sIb7Ge1Qc4dwfsTj1HR8RcwT2Oktz95s/pPPC
cgwGQz+dEecb9ugvSXIelcUJoAcD/rh43f5U6+NZuY55lQdFrt7p/T+Qz9UzSFy3zw0zHZneBXTd
eGnBIAvvatoppRwmNhNl+GpLVe0CE625jOO0JZl3fPpcs54XNY3M0o6MZy1mGCqZ9hKi4TFNzEuk
K0pz8NPsNcLWVGi3eWtvEr7KFDwQPdVG5LthBweXIDbw0RgPslK4EX8K3gwu4W/Yk7CC/smC21GX
308IKAxVabQzHpjrG/w2A9tm4iQ9v7bl/zlkOFlVPjqxpT5+gBg8b7qA9hU3X4DtJHF5+JVHYAD2
l56fF1J0XHQ4Cpbv5iNH1v+Oi5+HQoUHLNep23QaF+EWFqEmz9D4EPFgL071NpU09Y7DMjPyWbRB
tzYYEYDCwyYJKpm3D1OKrFkfn/NMFSKVztlbl6uwmOejREHj1HGNHpX8d7nrefDrHVrSM6ehrsJy
IZVADxARzwndPHtkmhyNvPnCEdy6bP6983VZ0X/alvl3i2JWU3SBe8brrlzalLcqo6+tvx4lJX2x
94/+wFG3PGw4ZyC6adLcfpCh08B63HZxU30WQTf+oCvB+vznCQj7E6MuFYj1+lotHRlJQnWB0evR
aUH53WK6bfPYoKODSio2/5eUC/Aty8GQP0z+0zKvBlvKi9iRsH3nyKWyRHJ4XN3tE/AHoTeBnDX8
bDjgO96Qso7pje+alWOwWz5Kk4/DLr7BQhE/sVX7gEBzrvIIkf9JYWDyxWFvkkjfqnreQZCPafrr
VWjZ3v761XNTca0VLPhSROCeVZwespsXQrbAqOU49NFcuV+FTKNkDvUQsIVLj/vfyDjn0GMedRVr
YuDI0ji7VDSmf1aCabhaK3Cpr/zBDQlpvouECKLKPnC7i6fFad1KKtRZ2/PDP0lw/0kLPxigIyV4
jqF3PEY7H+dnO8vJGNKkAFmWCc97p06MkF8e4ynnutfytFzsJc+DwtDUj5j51p776ZrUoL3Lriiz
k4lk49GkzE5hOLYqd8Du5pZZzGwJtTQpG0fgt5sxutft5hhqhM+eMolD/soMy5Jx5TlNYCxMdHZZ
bbShOD+rXmjFQD8qJ1/ecEwo8TuCJRC0FwvlTXlhUGxlqn1iQL+bEvXIgYlegZ/KYV/OHSFiB2H8
3i3B3bUzBglf5ucrcFwo1FzoRbwYl6JlxFGPk7kGG8obYPssiaDmZq/iTJzAh7nLHVZC6ytIhPfK
zvVqmzF2E/gm2+PbuZEjwNg6YBml9teCOlomb3ZOrdVjpl80w2x+Qbvh74t8M8OsacjXD6OKmcPX
wt5SBD/4/awved06yXj3KtzyUkFHVyrfGOZrM1OHyw5Mkcuvc1/wCRwQ6pTrY7Y+wflb4W7SbJmT
YURBxIR4QLBaLIzkSanylvG9oTV2fEHL3Ww088PV75PLFTqsk8hi72CgG82BLjIQExnsGaeyxIdn
UcHQ5YlffXfFgKByWHlWNkEBYTqH6hbMpwbhfgmXN/nikUCkm6yw3z5uIxvqWbT9KxQk8lphqhd2
MW5XjoI8+aJwh/M0aJsAITqIzMOqjfmM2x1dShC9HYpgtXTJRL5RtZSsDc2pVLX8t+PISEBHfzWS
4ZHtF9VPOGygsy+vBZHSdtBNLvTRj7tulvmEcAVr6P4VX6SmSncm/gKnNKy483J9YvkMBRyXbcQe
B0oBlUiNlKIj6W66xci0OHuPg46aTzpNrr1Z6gM8dM/PG/kVcq06Pi6qg8SJgbD2U2oycxANcuCj
fDks9D5RtDayDfMU7dOq0cV+LDWkTXQeHod4CQXXaeaLIau0q+uTJUpUt3/5YsSkpyAsK+u/iWO5
NoSeL3f5eCT+B7tQPec5iOL5/2nOxw6S8QVj5hks8zX1ObZ0arLJbbbFB/3M7YSi3VnvIvqZfD2m
8fZbWqA4hNsQYHUcT0dAosIXzbkAjU5ft3o48VYzmRkt0/8SMpQ0hOB/MlT0fV85murdqzAgDgeQ
I/lEkFRFi0Dr8aYM1Gx4hC4G7p9tJoTsbwLorjxDzFwhyMACa1s3YnK52QnKjkfR5idMuLE0Uf/K
e9WXu5grUIUk9szvXZkdihCkWWm11lY9HFn8JrwKbA5x4bGceff/fYFtCEKX7EE/h8rqL92V9ib4
GwVibxQJdqmdiozPaz7867QI4JPs6UDvvHgAnbH61OdfevqjF4RnNFryCH5gzZZuqBAjDB9/wMDb
MLezfg+eTf2wIbMkVLNciD4ls36NRksfg8eyi4q+6EABqTK6fsw8a2foDre7maNFNe1bBH8Sg9op
PHwojCiDZYLLWijeBTEc8PPHzR70QTx1t+fYNzIu9iXWTrYRUTYl0TRak9jRuYaDvc8ji6m1tFBs
SZFG5qKVmzLKXT4L0NfnZf8MiSTgQeid2wEg3JRBoXlJABEVp6mutGyF1jf/X9OI3vvnxxpHkUBi
YkoJX4tE1jL9+jnzRK6jc016+MeuxATZxJBhU2ZUtc+k0cDz5IRwM2kruHTvmni7eBQiUz7BTOQs
LatUNoyRZKiAs7QuOyfrm0VeYyBd+p4309Zc0wa1/vuIOfjqBw8cskCL//A8trCYMvPavbIoLjv0
Gl8tfPOlNtLJ7QWPziu/ILcwbmAkrlJfVq3ZUW6a2KiLJkaeW3RYTwF+fCUzM3F0vwZqZycYuAjP
dvkBzHcEdqfdpsCD22tFX9L1+nIbtnuRm3Ukdkwju5rhRLXvTqEv/H51qe4tkNJ8A9soNTuXjvPw
F5+ydk5oMbATpAm9m5NncXeYJ3X3XwCzV+1iymOX5EpJZEpfqp0SQ9KPDInIR1vll3Y7tJwY8fpy
Fhjnwb7TRV/AhsJay9kS8K06zbukKCoVopLYIzX28sR2D+8eKDGzVd0eGvomTQV+96wjQfukGZB/
YR9ADkA9xSzrMPkFA9+eLnnl+YHwAl9VgwgGWFa/jkW+oRJMO5YcWW0F+MEqFicOjOKO88HNprjh
UdmbXd5XlK8B+eX/nbeGWPr6cyCBAU/KNhmWcvREls2BzbqIfqml/0LVvTCuXK8OlaJyf2fc8UTq
phjQCjKsffYMhrX+u692Xxq0I4BoxVAx2rMhCCfwgPTw2JbdqC9EfZL9tqB7SR1fcjEN6GsXvFIb
T+75+VhI55r+GyTbe89ho6rO6MuqoPhBQjiTGjDyKODJsTWEiXihr2uTqL/SaPL/avVYVAVkHRvq
C3rTaeubIefCFa9645yFtehbyE/GbRXFtU6vZmAQfSK34t91qTGmVLYmvDfu8ELdGilnSRe76U/L
C0rMqObE05iFyUnKzuXpRlrz+Q21/5+BTTO+fTn68upN7y2XdWHaP5IN+wexbxjo0KaPfNrhwSdw
3UrHBxU7Z0nCgk5zjYH3Xl4pKN5r6kBX8yZfzOWxMl3GQ1aDjF6qOZRVljjw0VzgqfYVAmSf2ad5
rDWEUTq5sGAUhSv0Aqs787vakWhtnFzJxwPeY9bbKkhF8nWPxEFw2KwfHl0BsrIr3TRIaJbryNV/
EIo88dP8aT2mcknmAPr2t3/PdK3r8k9OTu5rFQElVCXwnM7s4v1YUTWrXLEJ0XQdqngOf+AvdPbW
XLIMH/RY9Mxk+paangWF5d6r1vPUsAlK40ikP/2ZDJZKieOa2wYxCgY4EYGAatLlrrpgbVhQrutZ
1NowDFh9Nd8xTh12RGG+R65tm1iKoQfsEvJbBNk/CT5gBvbJ3Dh17saN49zzPhQKKIKI1nmX+CjI
HjuY/1G3qQU73jMtIxAXU7pZYj6w3cQp4FIC6O0EccMIP9lKFbL3TbBOMO8nY6xC1E2GNEilBdxV
jXkS7ciOTtkzp7Wwn7Y5xfje4vo76QAYFcsyMZ4LQzb/03l8eOZup/omWB9BVjku1zCmBR3N5AQB
kSGJpqclqamGxuJnFv4CXn+AFTA/7lxVpIdV9bt/yvuowWkkakSXM93KCo8IxdozlSq+6xaS98K+
V3EHZyj1o+DXFTMC0dJfHlk/1t1KnkRqsEt1S2c1P008QX2PoZTwksYoP807uy/b0xhjOASKFq2C
uBzQrZtpTZjgsu9GGxYZ8yBCzpiIPE3N3reMz5uKI2R1LWnxf3OLafqV03PxKjv1HooCMpE3ElPf
VIYTQSFHiDbFSLsdzPm9DdZcFjRGdstU5k8JiKBH6HhOLbQ1TqhtgwFiY2Ch1QSX/TSV04k00zKF
CcXtJ8WEMiXEhx7OhBNU74kWGJXYB0kRsFjTKaGy00lVs6CA/SCsEnqBoIzThru+p9wMC3TrpQ/W
gDRJcSOJ2SX2eq3+kq4lbj8z0QijuRBFZeebDV7DLsxwlCqWPHMnA2iIcPe/Mf3SkCV8EWtWPdrT
OObti4W2+07wK9D6vyhqNk9oY6+6CPhdae//6s30rrAYYnijZjzpdptkWc1RsQQXQqclpUdAflMK
5CypKFZeWZ98J8tU/gUmbkntDqR8OfNzKsx7cCG9IBOvHYnJXEPjC+dRwsm2+0BFvqfbXaM8Ht+F
tUyX3mCkcvx18ngreGfweITxtl1cZVC/mgqggqQCS/k0Hcc7/Bmv8nFrNyJA8fxmHqVzquAYTYvd
o2KE7WDxpcz89aL48v3vKdN0e8sg/00o0Q3E8DNuhsMjdfZQYCk2JHvNQoVEZubqCRjSTEIU3Sax
Qo45FNlaa53K7e0y16d0OpagfHYSYKH0E7F9H+/R/4ORnf1sZbnflrO59Fo7MOrZbklhUg+1mzXV
bP9OHbMntxZ9f3Rn0HpJhIzKxCX9nUQqne0sHfBOn3PnSKBCR0adQWgM6fh8y7XpP+N0v0dDsOYB
gdMHeWHBRUawoQG4R90mprihNJfKv/D5KEKw+NblaijgTRIZ4o1jlaUC7+dxArNG2K9bpENOR4m5
1JhLPsNa8cPgNOEMtH6L/JxdGVrNGqxSpA0721Ie9wEIMw4iZq2S5q1GW8cNR9+QKdN+TxzzcoZc
poja7ZVtNkDO8Eu9GhDCBci+aVjf4hLM6JmRFiQgTv8uyYYv8dP0ofJAqLA+ZBCmqIEwTcsxLgsv
W21tf3AH9iALaCxG9Q32MOC6oqtt2FV+4p2OGapBLqaPCecJZu7vWOhqD9OpLtQeHuE1nP4i++0k
SVE2F+RPdrcsFLn9/ymwphHOD31cxsEHgeecW6yAZ90BAYrPpw8UIUs8tY8cFXkbw1WN5HoA7QvP
93aQMTiSNODavcyOsnMK65+v2+Bj76uDqI2temuntEG2dHnETZAKXeQ7Y9Os+NXKPptA043Oe8kI
6sZNFrTOmuqxp7GtLVlZnR3F5e4VB4wlwPsZKlpKyMYmo1Tpby3BeIt199KaSbmu4IL+FWhAI8Gl
lcPsZw1EA8/22Yec2PCJFYMFdZid1l0VkYFMxFQIwCuW15NbAcTQFpTfPgUaW4uSpxOkgyKygLDl
GqDs+faJp5tbkxnxcdsuCavE3AdaJvPAAoVfGKmoqzHrGW3y9zy34bNq0tX/kpGUN+E2e0xH623W
lI+8lXvbp6kOMdYupmeh7rRCxdeaNfcHgGMYEgO6qccOW8blPZDJZRpOCbIkizCWgOWd5U5dN4vG
9lULdqApSndc4XhxK0U2xc0EADiyi1r4KEB2a9jvOdmnTTi/O9+u1sIccP9Yv8hBRrNV4ogM1Ubb
h/841CwUqbvSaq8PTv5Mic2OTgtGlcNpZjbQyXtva5AnpzF+86KoZlSdTL/Yhj/i5bEBhHlHw6Gw
QL71dYdmJ2qhrfUOk+cGRKJZn2a79i+Yg9mrwJiNzNPaQuqFYwHQ4t30RjU4zbqsecyA3sFEhamk
NGAHEnHYO2Dljxdoq1oS5/+A33mWyEAnzObkw0MVNbWRVgenlhif8SI05k6mFn9PCDV2NFxX228J
Ea8spVQ+Uu3woRoRV7C7UItbU9N563CosImAnTSwJ++FvyfvCxpOgFYEv+Dqk+TbK205pFOCEiD2
oh+BRo/CrsOamSiF3OiGh1lemacOIYBQ9Eowu8NUrauLvEtu0/iMHdbRiTx4eD+TusHtB3/rhq2O
d2qpTTFKbMeA44ESSgmVVVygd/MYZf/RXL/wmnWFawcZl2rbm5IsADq/pptPMmSAX9ODWqPRS8zH
W638RPxuLoCS4+fExGIcSvvUcvyJwsACTSonLB86psRlg6XHk5MT8PaPo2wkFpRA/ev1eCadBCdY
Xeal8gluLKpfDCzzxmINyFbSioBKGH9m1yDA8AlOmoIulKsQgEhCvgrL482tnEXEzc9GhvSR3Oq8
VMhGd2FXrH5HOv5OWoqPpkCd3AP4Y4LTiVAFSHXrOh4p7UqVKLZbYpeRCzElbr9W1fJ/tDuW3Z5c
ePLVw8aqi9/OWxymyV6ENCrwcasxZ4b5mZT31q/1MAkIa8HFvpG+NiU6/tZvIJkkr+3c/pl1S+9U
dpQAtXm0EHxcBRoLyXP7NRRRshuxYqZMS8eWXjuZ+ozGDITkPMXNR+19M19vjm0Y5bBAyDaiMcQx
A8vm11qBDnZrQaT4t9DJdL6nNwzT9mM6rk/qGzEOiPWRv882Bgc5alve1WRc5KputiY7lVZTUFAS
AJ5mn1zSMXXF5IT9qIHWuELLu+W1xSC8E3hVFuItQxZBkFcJ5eV4pP/L2rZG81UoeA63/kyxm4S4
fFBK2B2p2JDs6OirfxwuydJnLbg7ll5Puj6wzC8HPEzzSG48YxM0iFBiZJK6gYTFdKT82RDSHCtq
l5hUikrQPIoiegKnozmCOOWPAa3q/pNZPSDZHUNy6XtPjIH9HIpWUfC296pknr6rflGbDagqc9kv
EkkmfWcOwjw0VZBitGE70sgufQYucnAOhaaQ5oUBs2+QC9fz4MuKkNUOOYkjF5+RjFqwwUyiO+rg
bX2aMw6DJYH2cX0c1e2dpcsUEzP1OyP0Wgx6vSRpjzTTSuSYQ0S376O4uuPBHYQK2LbEjifQX1aY
CJ5kN3NN/R2SmTNn9n38Zsmbwu0j0Jw7tRHKvXMOR/L9wpyii/WuUygX9NPSN6xpeHLkxwR+8slM
ZDVEm4QaWfAjD5ksnVKImLrmNnVAquaJrclKYOCcxS30jmtcZhALC11+KVfGjx75g0TOUbCpmruz
vA9ZwMn/h3iFY8zMcpr/fD5vayjUu0Uw+TDPKsFLXa2CpYJqiIPm9m1Lf9IrhiGHkJyUAKg4pXnT
Bn1U1mFj+sD3zRl7xIyWpTw85LodBhasaurVdJltc4a0kWeZblV/VudjFqAx1qTvZqX6sLqEuCSQ
fCjkin7TJOi6n+QQAFP8I5O0Cy4T2FqGnZPvgUAui58TPoMDSPGgQmq3/f8DaOmze7YaNFteFSjj
W9LVLCQQ86BbWWUfb1Hm9uAD9Y4vX7douJ/bWTCC5OLclANkxC+u7hbhCzvwArp+ccbnJUQFTp8W
Cb71iW5c19jhU566cc0slfVKcyHNg8laLAdyOnSLc+dDNvRG9XRU7YawIUa1cTaIGlT83aWkZ7Sb
D49Gx4cT/Yvm8Xv/V7FBq8Uwj0nIW4xlu/4f73PwJWKAQwMpHKfJFVLf9oDwCOFe6+Bo2Fqc5XMt
2y7C/XDglwbOjpFY4YU+vOoKQBaXSbYKT4yKhpa2vC3R+C5JLcVCNzQHJlwd2BiN9G41b59ipzs7
ua9wLDTHTg1tK+zAoFLdVToBQyv20fnAwdGG3A+O7YGIIHIM/bkSkdxZHZwTebHgNwjyU8kyu+1E
0y/vMqZf6h3AoPU7JAxDvq9cg85W3+Ndlt+BAyCDiKzhRcrJ6MI9BpD3N3ZpIl/kfJO5NPkLzL1A
S+vQwteC2wp77Wi1NFErut7BuD7VuJCceSrqMYTXUg5YVDT/rCWVV52oyU1bYRR3IIY1R5cHtVAF
CnW2jhWbnfqlHTvXHi+UJAYpItvUnyvi6jPEJ16Jvhy3MeaKvrBPNlgXxPXQ2SAghn9o4nHbwNZK
TbRDGc2loTRBJ00t4Xw0mpG4wtb+tnP6V8++mIxMSau0dc2wa8Jfy/aIj9H30iJ6aSMbaa2r4LzZ
9YXL+aU1uX+3NnPcnBfaV8G94drQySjkSbbhLuDVLjZCHhjKqSj3lcTn3l1UEe83Z4fgYURJd1GL
fygtEJ5b4icG8e7qv8d7Fo0nGvLC+S11Wa6PmhCNGtbEZ9urJkf2y4C8C4OmGhKJlwojYXJANNMO
AMhAiL9CT9/7yp1+OqRp01sXCTwFHyWRVmwakS5TuoTeXusHqsroiOzdj1xUvsS9xOhoe9YTRw88
jd53ZJwh2uMXECvAB/MmETiyPfEgTAtUsOmUGlh+gVUnLKyhUgPpOLTwKKQmnzd5wOMLmrgYUMjF
hB3TYHx/PkvU4HvhH12hgaxIFBlSIDKAeo3ytz21A50U5XDLXFd+Gd2nnaQ38No1+EMzPzwmu19D
E16yG3JSu+MVKYq7CqMz0EdYdVKGuyblG4qWQE/+0eLg+R4IGVqOSaxp9Hs2NlPLQaFi2ySWFHb9
Se7J7xoNldGyhKiUMYCkgqx3Gn9PAcKhyN9EMw718HAOEoIFq7A6tFniAG3tkCyEOv+zHjzVSnrg
88WA2UsPY6mTlzwYOsSOSB8KUuFzAjm0De0IuN3OOyUw2WeaeZP38tiCJB1CAiRYyhnLE5xn1SME
IqVZ4xe6AgAi8FaKdx9zXqMdDkowQWup/jBL+uFitB6i2yPmSIiO4r0tRK5mCcjuzYGvRdYjosz/
M+oGypPu8EpRyFrR6Js27bMcEnVk6FOtuxBUSHas/bIQXxm2CPf3ArjvL5xmnFF30RDCCzKsIcTm
deXCGfHQBShJFXtJn8HKLKguvvU2qIM4deGbqpgxM5yo9zkBhxI9HxfXVcGkMnKDfoFhKsOH8AEc
rWINStmCybbh7k99VLA/giskBXMzcUekT/Ei+15d6ndQzko3ltLuCaB9EC/YUaM/3UVhCeZessOY
OX+BJKqFQLpVHfrFicKSsh/iriy38u3R2TbCCUG0p81k9fCo7NmxGhV5zy/Zt7fnSEK41NKIagEz
aUCOFCHWQSOJxugIXfIoQmyRHw0oDSjkxQI8ajoBTZshiCZqFaZfeGXx1ExgCMn+YJsOIxCNt7cY
3ydfd4SH2eAaeips6f5UWFMeMBkboQ4fx/SRYXt/Tz0SAXJ58LUbeyd3n70qffsn82xgZtJ0Pvad
r8xxA/TjG/k0AFSh3QsU5aaLcFD5p4XkzL+h1zT85PNrsZIh6wi075X3K8EntrToZXWjdsZ7J9LF
vDFO59qb2O2p449h+bQGFnXhRDE2HniDveUFCBX4nG0b19u70gvkGyIsmPTyXX+3hilYK6qWCy6H
bc1Ev6xcwFZ6rS77tbS5OoKPOP0dbefrTzZljpCoEWRea1KcA0FJ4U7ZHln+wZBa7ipCnWzq5FwG
WvRtEPm2FAtfQmXe/Ufe3D3r0pTHw+FLR55rDQ/hA6cHc9DqSVGX7ehrlYfnlgPI1GHXgXoX5Fo1
S/4nOYTz7FaTEiF3oeKwvEl+PuLDa6ut8Eh8hNFM5bhSer6dpWfP9UgHpDtLmFDF5KRx6a2221qo
/+BH0NuEpELXX4nT2NI77rgy4k92318vsA1+D9gpkukkLBbUeSmUWfhf6qOmw3FWP28pLj8O0RGP
/toyCzvdTmGqzfgB7pXwHbVmfKaRJrQIH0WzzTSyAx6P3FMNlTfEAy7XfxGggmVf+htP6obaR2yW
BHbWTSuPcnVRMaRth9qpID+/1Mb7RNOqsTkh4p3tXxqI/wfsHfL9DkZl50u+IHbhC5oRwNZOaQu7
/jFUOL5WqF/jmc58bKJtonSNH4fa9NZ73bNkOh7p6WcHmvlj7jMY/pOmwj2rzxVTxkVYDFkCs2U2
8ZzMx/K/OIIDPxTRpyd//K2xO4J2W7wRoIbbzvJcY1PQ6kOI/CvjLmYsWnbiGjeJRx8qtJlPeLCU
NVbpKrFiHhoxlrNxxmSOIuDCdzIYppmOSRV9EKjl3mRdAG9adi/N4uXmCKh11vmuZ6TXlyHpJ4bu
IGNB2LlX1cBLGWan4HiuwSBd5/I3A13TJsekXsoYcunACZpLuaYUr4LmS/DQtTLrXDSFVUj9DCVK
/wyzrKx88lErMoMsv7DVEdXQYbjk0gle3ARqoPs4uRoG3tfVf6czTaVDyOf+p8ZLLsMnx7nXQaww
WaizjWDcAQUDJViNFyE22wTmmkyFao4oom04OsnkA0oWid+B+0sIS+6b1HsMvDnDMvWRUr4+7TD1
sDGcaDfCcUM6Pp3iD9Nf8l0mEdDX+ZxGctSUXaX0H/zZJozt86VVkYKZYWvxmpzlbHeh7t3HGAR+
BOdEYG93X+OmWNHkoTKT8FcWdJ6YMSS6aAaUTbA2/ZidK4koQUvB23C85xmSrwaT+jHKQ8MrHiKC
DbEUiV4V6PvFq2V0W0+FAFW6DYwdkew6nSJpFvf/L6xYNHQPkKtrBcDUBD0fOaZVbYfUCMKbkyvm
bukn3mjlFuTQ5z9oZg1fmNm6u0Gsuc3xtJOjhWv7uhWh00KiKcK93uqWHSub+TZeEj7PsruTvoUw
+xKdACjcij8Sf00yc/mWwU936kEtZoIq97xt9d8h25hxJVCByvMOZ8R1KEeJAlekfSYwUdynKT61
wYGl93opauObbNaLqZ54BhuGnu11erxbZPjuycNR3SdcgFVUeqqi1gT5hvHWbWpksvIOQzyETKa9
W0WWOmEidyB6iGkXI860TYLW35zQ5QSFxS7+rkS0r4IS+e1a1b3J9h0iwgG9vpqEusI2iNUtVbr1
gojUlWRi75s37p/aEGa3gIjcknlr3qsUbdjNUlph1/4f4EqdOfslDfhhV1CYeKT8EHMpVBOiaTUW
Pcgd1Xomx8w7zQDeKFSP3vzsb4KTOPPvi06D80NhoP1xhJI0JIsaN3mFD1rZT9Aobq8Im/V8P3hQ
GG2S75ujrLBSJ4z5laCTAEIEXIF3oiWh5ZFscsqIBE3iuKgSvHUsORIzaC3oYBlDqf9tO/DpYvoC
OgKBQtVHnbQlooNJQWYtLKtti/8BDjh/4WjxBEcYrU3fnQ8mjO79XpWwcxq3+3KYq1OUuE9kgHSb
iCP/GsuxCiMQRlC3HsaBawhHfW5Rko+tGXip/GD5mOrjekJC1vwI1i2emA8r59pTroQfHrxZY+R/
rxPP5b/tMjjT7Oug95gWgYgKF7svVMKqac/o133SVggVn7C9iIFkHUEqJLRH0jKYJJh97cU5ElnU
21f93VOLevJi/Cqa8IXY49khSEuph6BwEQ2fWRDFu3uh0I7bbb33aEy53EqoEIfy0dITZILJRDYz
IEFW9pcZMIG5CCcFHIumTrAFi5+lupIUMQMUCIHk6Oz7zycXQYxaxiRKiJlWi2SJrkSY1kaREkLD
zQj6sSArPg0b5l+mBJ3HfGggk21IbRo/JEo8Aaet4kyH+v5AAxwhEOsyX/+ZC0WOcWe1O6oKjV2K
t6jmn0zIBEVZJo1908P8WRPBzX8GARFwbkc4qZKYLDk3SABcFwuqpiSRrWTrVfEnqVPDK/qgZD/y
UIWpFeWiNOWrYZHMjmQyCbZVEAP7ueSzkgDPG6fBCcX3uHEPPngnbfCxxDGwHHhPbVPRbb4enoga
nA0oQRylE+0nzDT4PSlBxYE8TD1jb41T16k/O2oa8vl/35M3s0bt2iCgpOhpXPmoa+1C6m0RcETs
AX8M/dZVktjpYrkvE7H30GSv1mW1poP8JFUdGoTbDO5frvovJYI5xg1nirP1QWghPR2y1PMe1ity
JAQQJyL9ixgXKQtBQLJ2U5v31TBA+MxmntZ9ns9j2oZ+HLzrWsm0XTDAve9p8jHm1aB3bnyLp9dN
ji22renZAhNOek0uZuQSfmxJOVltJtxX4/AuZSJPVjiUthIcKJlPnZfznuxJj/x1rESCoOTQy+ND
YVVJtIwwgPI3Tp2dXidR2+7FNSK2Krvr8VntAH5WZZdjHtv5k3XbTvzP9fpDEX27qCOuPPWdcXeL
F5g7QTXnFtjedo1uSsBb9o84BeXApPE3xbWtmzpgShOGkpSSS71aLRj67jDzYB60WaF1yrkvYN1H
jJKDc0SOCdUeoSdK11+PJGtPnj6s6Z8xF9jna9hq64lA0N5nCU+lH5qKkVXqaNXVGd7kt4ga12Dg
ICX6zxsXj2x0hyW2yktd666wAF2p6pbN5hIuz9DC19cXE8o2EuytAI/RZD7xgsHW9P0vCXrbfca4
VrT7UQRw1mcKFBfWu8D47Ee/onKmAd3FA9QOG5JZIO4wBd75WmWO2iEpGB4Idt9opk1fMMIhrSiQ
jX/jq5tYpYqYA86nuS6Uy+9mAaMAvYlxHgvWtA1+tgG99G3VjiYX77DsKxx3JW0Fn+/cvMKZ4vu4
XH5brgpq4f7q824Xw8UqmKmlERKXjTtpQMqkaiWgvusFPzjFJS82K/jy9L1JdpGSTNwV++Mtci6D
UwWdX4j5TmHy0i5KVGzu4HCj4dYlEZwm62IRT+Lu+veYXEzz4AQ8EJp4GtzzWjn/WWYvV0szjwEU
3o2MmVutKVJHvqi0c/Tv0j44/r+Fg1mJv/BLogYVVx7mxi7Au2E+rXK68AnFiB8EkfslD02WR0V6
vJ3bDnn+SjeKD8KL2Wzeqsn3zty5KnkjdiaLxKck3uh2bWgyN1C4lZFMYV7vcKHGaQnJLfKADgxJ
8xbrrQuO9c9lQwq/f+0RvDgb1and2Ci18Q7CCkJc2tBmN5z5Pf5y3c2CCcXQHqxTmjdjuPLS/y0z
xsqXJSufvcwQEcSqQWPJJbcB73ucVscJYOAWdi1tgHSCKXriGuEuurTq/Ipmukn49QLoh/hUirrN
2NkH7le5R5aFgMAl5j7/W9mHMFlTGoAMfpQYiYdqiQNawcUBVt3zosgt5A83A396R+G7qEL5Pq9K
X/KBEcFeIyyaOhJ9jUlemy1X8Rx0NDKXmg/Ou3A0JsASjpqxfP4zeCFRmpP+x2X8RmOLj40w5oq7
c868vS3fvooPTkWe3tF/Ac9VuZ1sZ3Q4BgwxJdQ/E3ZFBExBHl4fxbxkqhIUOqjbPxD9ucyCZSSk
vJdDHZt7UH3EA7ztW+1xRmS+U2XalNHTLhN5y2vIq7iN2G80rFFmsjHuBDcV3dZrtfTfaML9dPqR
FBhxRqHMJw03cpxE6l7vzzuJAs/VHTimy0+6bsrhiUmp46MsqFGn45b41Q0FrNXSQH+azqo1tAV7
3MWMUlINgSED2dGu1KOxb51mO1+l94aFjzt5OrrKFLBe9SVYxkHt8Wy4i/Sf9m/oTlAOBDJzjG/K
hKupUS9kN6KTeQfUpH7lqksfhM7XE17czcroVZBnruaNWu6q1n3g2jyMuDlTdsYCDMuef6/rqQgo
G0sGiWdb9ydpR1wCf3/ErZvEVKhZR2mGufWqfy9O6s8nxxIgII5OHmI8hXudxnCrX6o86z5+Zkov
hE7cHiMX1/AFhF19fuyz2w2eHtrQeRbkL9t7LQeuRCljTfJJghMm9/ZUrKJ8Er16kP1tUgO+r8q9
wg56WXNBfUm50VWjaWKDwae4ogYbOEvZZCz3foAh1rHLZ/sdsyQlmn4P0kw8+1YQkgqnp6U1pQfj
YqOSpNeSMsFRGVABM81fV6APBZiNX0RK9Of+wZIwuCGklI6k1zUaqJvf+AroyOuzfaKq2/qkI4Kn
grPp2b0so6GOwwqUyBviUTxfJeI2oIO+7Y8J8BT+6xRY8VWthvObanVa+xSCTCmO3s97vzFUP/vX
L9J7//jWIdLhD14lP06cA7s9Tk0xfmw9UC/ycT2msBnE7JfbqSGlGvrq1z8Y82ew9tU4sTdCG4+i
vk77IBIYYgjyA7rv6yP/pLb0ZyGVAvBckoSG4AicaQyQLRyCRoQlzYgOnuUF5V+16fYeIKsB4+eL
EPhZMiCFHYh/lpaNhydzcAN0M5K7Jxm73rTXfqBvB996rA/tcU6CO4YEUFtAjDBZ956D6Ivx8o/Z
6WXw2kZfdC4F7NrcNB2H/KpcaqnYJXHwturvTT0i7oii/HTQ/4dDkcVtE+baQIXGTjVtodYsVKcT
87zSIE/ASwvBYVNDaLkHLdV3w/HKa41OPKUHuQ0Gh/6hz/iPoCduDf0AOQGTSE9AUWXnm3B8+paM
xDADk9oeoeiyrrJqoSt/yoJSk/xVqqcbszlCkJ7qp6WAw03Bc2BiM7MaW7FKdFrYfv1liVOApP22
uVeZu7j5R63rCQegGIZjBcbuU8HytmfNTvRwUuYzs4lVYYSjwG88FdQKfghMHt3ll/tI2FsB++9H
Mj9sCuGBOZUjwj2CI5fcJ2Li5wTXqAUYiB3tE+liRKPxfkHwOkG/H7JzcXyAEinIDkTIHhw12MNE
QQS8mizrRDRJmPvMKHKpUoa83yrqELjaF+6eFvRjmsbi2lcH3DfnVdqKnAt6O1C+CA0XuV3iNxdJ
u5plCM7LEC/2UxzNs7YmokKzzFqWNf4ZnNXB0Dt01eNU28DdZ+UUk++kopQdugYRInvCGW9dlcI5
M4UHk0djuEMuD14pLHS/DFItI+w3qw8QXHrJzSHoKcpIErJB43eIj0+rV5NX1/2HgLBcBUCJKszL
uSEyEIxgX5AUXJ2qk61HADdk5KEDWTpW5ZwBVxIvYVmPQm+VSAz0/YyH52qLq+vS2Lb3wepIBVhB
4kbENU77uW46KUSHzuEDWlfN3W3u7T6NgifWnQw36flACIb64J1vQzGDJpTyTXX0AM8JmByigPLa
LCoAl/BHworhnPqrxk1p0qvWqJMWmK3XjZMg85EGP2TP/9STXUxv5SW6aUe8My9+Alr4obBSxnHh
QnkWYBDcLjzIAmkqFoewiQVkDI857Az0ryfxwQ/o8V+jkCmgPE2L3RWMa15hFrJGMvWoP7Zd7RA7
hkk0WEv83sPDP9hZ+Ev1Xsw3nhkyR6iIMO3HUamDbztC2L34m7mtia2bm0Ws/05GspVLdzfzKFhI
qWg/IsKexapKH/fp6dQpuvXwep3kE8IGQKmyNtTygOpHdMB3wcB4hP+spAfmEQKDcfKh+K6lMQ55
w+yqe0cH9Y5x3IU0iRQULQRZb+acLook2BWhZ4scAx+X1y8BBGrz1ozh/buJEiXMO1BclIcJVutS
qDUrnKVONO9AFj8LB5B73Ps1paHHCv6TEyoyWb39Vfh6SfCk6bDhoWqgPalcT8vuQRLKvA9wd7Ln
IIwW1gRn9n0CjZ5uSAcSY4oehqCP6l9KSgMdhmLRvL2/PqpWmtAgIwISIyDd2nF1t4VSQhJ9sSbj
gmMJopR5vc13jPea0fbMARwBHalq2ey5Aj7/9wZ9eJofZypQwGGJzNp3gjflRBkYmXJi37PcBt1j
jeSg58lTYO6alSfRPzCZ3+VniLLqFaOJGQRd9DZuJBV6uSYQEg/HAnyySfYzlwQvPLZ951kxZo8J
HDVI48SFJNf4SSyI4HcP932Pc/fVIvxOP1tzOMbcNGpq9f0SxGTirTMX8fa4jyPmOO+4bE9VpxdC
8Yc7U6QOMXZDJGJDpu4TogeLu2GzUGbDp9zmkTZ/bh59ruh3FXWX1edAq2UW4AWKPP5VBC3iy/8f
htN4nQxHgTvVfVcLypqiGG3TSqTEySc7MNvj9Tts0q15t/t/geXRRiM4ZczEFsj7vVC09+/Z/1+z
nqOEc7aFUMM5ISIMaY8nKmqVqTzAR9qQN/TlcRX6cTfk//Yy2bG69CobJiBK/SqF26P5xTuz08Pw
9mVx/xtib5X1r7jzVuF4eg00WOPE5oP2PlqyJf0vGzDCOrw9BMs6e6t26ImwKSjV8qxaH7W7ka7q
WqB5fhL0CcEhw6M3B0wc+C07z2hJQrP1SOlazWaN5KCxzFtGzCtgen61gg4MjaqQPryZpamqxCKH
CpROq2g283iHi6Om1N4L1tr0sis/UlHWFOJOaa324mfUkT/v2sKYPqzBkBOf9dGIZk2+h8fv5li0
Pe0rUF3pnfewE1F0R1VpgfiXEPsL4wBYUL2RPIn5pMYHAOdnHJKZUQI20PuAKnmGp9qe1MhcHOpz
b92piHkdTL7psSbPAQ2jfKgysjmRPk5AylE6zaihyDAKb6DNpJKAf51r/4krVDokwiOjcKGXbYoQ
akJa85m8uYWPJgsyMmGqSNvn56UYJEXNrU9AyW/RUFvg/kc6rp0yWjvtAm7yq9unl/RhQ4DlDAK+
xyHLH9fqKv7FLmA17lh72S5ZLfQvyhxTMfcCyw69wNkPQaMcn+f3PZMi8SCZaIVDji8bRfT+gdoY
GtJ6MGnw1SepjvrfHfDfkp4Ks6P6LUGJeuZV2UkvWwwplVhm71oamL9kLKSfgOEBT+BeuZotQLy1
TYG79hx9XOK9SyzVON+O38+esEK64x1WZh0XDH6GCQPAVgXPI8JGAb68EBD/WMY1+FHktuyUApcP
ljYtaqPFHTvbdGnqzR5skXYP25ZGUCO5TVDy1jNDy1JL7yxZKIEAkzRze2PFMoKdd26f1ZltDKmi
Str5Oc0DMgCKXAKLxb7zr2ihOI87c6tROBa14PHP3ScPFdZAaaruvAEiH900NKVJTQhTPFAtgbEI
ktGqmRXRsa2WNUjejBl/qFeqsoTV74Q/HFWobSYT6TK7ikO7qwQChodYHkVBnZiPTsSP5Lb/Nrzb
JNX4+GFelj54B5aMiEzUPiaUHdhB5ZZggYi02DRvDl7XM6eYe/SpdxGVwoVWY+eI7Z1o0zFCyijr
wTnMsm4E90puVRzDptgFCK3qN9GKChj13iNIz0Lh89ePEhbi99Sgxq1XVFXSMEnGFWWC2ev7akz2
h2+rTdFsJ3WXPSxCK4fVzlzh6WDCACrCCFt+kQ+4PXBfYUAxxnmHPdrF/XmNqQKa45sotJdnJk0J
97wpEbnPHg/QPY/TmsibM4svMm1eEwMA+PgEnxSZugIB6gxLesRJjDRz0b6e/ZVECNCzXTwqiB6w
BPDc11HoG9k+WOEU3oJvcb6y5BnhjnNBdnqjcH/1wFlS4uu02uR8UhfVjaIytUnZqjsm9pGB5kg2
VIXNxfLNkm/gOoy/TJiULlqeXA7q0XzJgSc7tKfFRFKSAWWUfTMOZmGZ02IbTXWvzi4gFKjwH/mc
QtvOBx6uc40C+PEgh7GDWaMQGrll+SlCQPz8Tz8Jkkt790/DU4OilyyXxpqt3AtPgVNHeg3HSdHw
LbNk7Oi56GGb05zQDZrvrKHvMbfrW67SHayc8lXkzTthIDw5nZ/bZhsbMTsPgA/vTFlXMsACJhjY
dGsYUDuaYV3YIxSU8/VRYQ94zFQ1TslyTrKhDkym4BqD6yS5zCpDOiiW12wXsmZ28JGj0VWWS9V2
a7yzv8kdOJB+FrgOVVdNIqn4TJeQ7pE0YjigTXj4bCS6vYAf8GU5uluRph1Uqh8rkbk4/Zm45C40
07iYR8ghQLsfXs84bSbLZCGBfOBLZVpZLr691oQzYRjjHtqfLDjXedb+VGGJNHaef/LM6upM2NQt
sZDVFDBzs+AWzSZfmyFpcE1HyUjEIgi0V6Mb+fWmM/a9wHNk6wMoDZvBPmET/Wn0GpNevcw93i4/
3hKp+b22MZoF09ri8wh3ZMUBgk1yQg0epHIF3vavRX9oqBQbpsYBlICVFwpPLx1+bwCFZwVD+e36
Gx73dgumYNChjAn1HHTULrr52/y54fj9HITs9pC51ShhsVJcoDmyrYk4dfzglIv/z51acb/X2upz
DcVYucpoeJEfZUlThJymV0eGuGRMvkscaoq18KNMTgWhLsc8tI/CSkK4lptTBV3tkFUXbwLX3khf
O4C9j/criC3w5ZD55c6G59ufAY21IjViWJ1J3pD8TRSBXWGryrgW1ld5QhhFApPlZIqhOLfW0Ofq
7NzlBoTGmMKFHYDFOeSPs9ulx7WfeY6LwvjT+hu3DxF/ZjR3wfqFdgoZXnqh3zt7nAvhAi/3ha0s
7Q5CBTFCTAvvFESNtSNPdLE6lkn3xlnWs93/74iRyKuCE4tqHz2N+ZQp2VAZCwfntuvDZt5ZOkkU
tuW+aGGTihXxAwzyxKy7KxotJ5iqZCW76oOZGiqSXhvE/dpQP4V1qSEcAd1L9wfZamLNT21IBu4v
C+OWcVKrvU0xUvGHCETiHclsqaMcgY6oGVQCdjp8JMDl1mRhrNihvHD8r9ulNRjx4dDZrLqmFeRh
WsOL3VMqO6/Pyg7zfeNH4jNOXVUAMriZyKVmmZ0/fEZWor7D8twu8e4TVWJnJE420KUhYFt0GKi7
vRlZlueVLKiXMivg8RRKTrEpFFvxWoJ/eO158lsN9qv47YJZnBuaSrH/BOvAiLCorrMuYLW2KSwG
RSQ0Xd1bub8cjuEMZWnitoFSJXuzDyjOx50ZJKe4NxLIk12ZFv1wKjh1n7/a7YiOuJoRBN5MSPpt
cewJYmfELCv9gaBEkRrgaAcbcbv6IJ3SmFsXzjFJMOj62azAVGo3EpiwSOdl+uOu0vUnKDOMi1el
C43HAb71hd8hIFxPIQ/SDdz3lajn11Xg+xh+H0qrska5p8HezEvdftm+gZrUwTG+spkjnHSxmUQa
H/47RnHSjoyAQjnWinUC/r1TT5NrdkeuetOdR771OLZiTWEeVaJ87IAFWow/eUfDaUf0b8G2GfxV
zIU6YMqrJXe225w/5Eg+Ec8uVZnTGy682ji9Gk1xXCQ62YOJ50ppsMs1KC8rE40jHW9W2vvtmZss
DDqAXXr6hQJGF7b6HD4TYt3GS9q9kNC1VoDJ5zV6sU1zwrTKFM4iUTMCIORZZsAe1gRRqgPxu4qi
XGgmYw+v9Ss9sC5GxPCzXEkuELnoKpqDHetsEYjueZWzdUhMZgfWyBHgRl20n9uPWlJZrMQfEEN6
CExwO0p3in1KJloLQYIHB5nlApinlwmoJeENXUwY5rrseM8S5glpp5SmhkuiA32suuY0MoMIIend
qTlxyqcYWDBAvBKHqEVlu2YASYeIo1L3qOJlq0Eax97SI7JxMqnkH74jrvZgLmplLxdbmZ9reVwv
xSqqo7QKMoe4R4532lUfJStQiLUrYKlBZ3xPdbTKdvvgVqnSphlpkg7xWGnv9SVbPhIe2mEBwf0R
pgusAY4wgAnGUODnu/nJ4SJDj/LLUDvUf1+b2YlaP9+kV+ehElV3FfV/YWHaNYcddLYyPljOfVw8
2Iar1w5vSVdu18RvLMeVYkft56p0ACtpi0DjIihojNdLrIbm4rZEp/VhvgCYW/fKGBnDLAWXI+OZ
sDu528BjwqSodGrYWVDYJ+a+IQl5+910iRaubCTN1I2o8nsLjcmWTzHp83hfUcMIsWG8WyVHCbKF
v5Tl1CldmQTxolR/V9me/r4Cyk3gZU6O27FlCpdRLUgxe8RY+r3k9QoU/XSxWwaPr/4sB0WHvhYR
LyaqTODfp5llIIGgoqKxMLHBSEx/VxQ6GlXN9VIDUdVpqJ9X1BW24fa88eaZIwQzaObHZjEQ9ff7
PdJ0nFMTux/3Dr4cv9C7OIghvyzsR57Nv2Jo1ngMBPap4mDOHt9WgAcfYkgIUUpi6Be0fousYU1D
6SdefHnCwbzd3W8JiyiJ6HPXNQ1uYNa9IXm2PLBQZSX/GcROktvOMsp/wMr+lRzhaP69GZ/KXmqD
qNKiNYVXaLxH3eYo7M3/BRzKyaSlDKtXIBgcSBGfi0v+oYO+2qyCbwpW3yZFFVpBD+CNu1X/B58b
eLEO32MzOsQVryupEIXpzFzNOj+0d/W8XXdWpx9zAnJsBGbkal/A+oUdN7OQGC0WT4LghlCDM71h
+Gs0GXH7lPZE6OqGO+NKxy1xJizr2lkh6vCUoebywKXIYqlGQlHhv7jxRrVC3S00s8a6YgJauF/h
SdE6v8q1iy8qt4xzHN9wUeYIHDKyWdDk+ckYyR3PYGZSMUWtPaq2aeCxuX8RiDbzq89MwXF4al4W
bVggFsAUBHze9Uo4D8I1LaAO6jLm1dNcWiVryY/fJhK6lLBuwBTaUWDGTQGG2Aky3+tBvrmVO0O6
m44Yq9B20RXiER+ZbCbl2vA7OB62E3P0BHNR/iNzD+xaLMwyMSDxGJbGvCcA6wRaOM3B4L8UYeON
ohTJOwmQvHdsixvLIjMRHSMoLM5lzsD26ydiebRsSBJkaHwC///lK10OcVWSCri3UMrJGPHHsORW
ILoOhGI9yiZ69T9YsR/oVYZD4OtWyXgi7/JkMUH/V2uukaUG0ISU9NQIvPrmy2BdPQZ5UH2jQcTP
tW8eeInYEkfzF/yCiY5kuB5VeZ95V/DldwavK05Y8rCj9l9wsGJ1Rr9reVS1T4b/MFfU4DiwV3IV
IiiIPz174RHwU2nrOFixZDKl3t810at3BxIU4gO3MtLMlRLCXzwibtCrWQX9Iyku75PVx3v2Uaxn
LzsaKMXzLQf8WMm9uRTxhlEOeC4+VXWBgtPwm6OP63Oh8lEnbmnQ0FVHDn7K0uywxmR3OlTrEDvd
Xj+tpa2ncdJ66ckeiNZIZl8sbgV0lfLom+lHik7U4kpERHKAQdAg8FkjOjsUdgCGxzTFq5wgjADS
SZqLc7iNgJMcIDCzVVe9b0WORprMG7qz8qGAI1eZO0qXY1P23GmtGDRImJ8F0Bhgeq+89Z/+MdXK
G9PKjJXEH9U7Xov4t5e0PNleX53AjX8uP1blk3VyFIYaxQ9yyPzJu8l8BtKjG6WeQgJukhAOHoOC
3x1SjZ0Ir7YNKsniDHds7PBNO9Eio1AQ2oCbs1kadpy/iXCjXTUK/T64hKMdABzxsRaK77HikFnn
IjAH6y4+W8aLtuPs+JftU7Ls7CHktwI4MZMQBd8EBVRP/4rQ2iOSgepjAoybfeCEWnqMj7gL22Tn
kc+XItrKQa+tWrmSP5GR3WwQD8Hs+eWtogHcYITj0DASd8kEZ++k4Qryh6GI/syrrZnOadXOL7NI
CqXJ7yLBD+alvA0GVWNLr/1ymwEod2v/HKZ25CW1zuTcdkb5jA14nYdnCvDsFRmslKuzFRfMRC4c
4ulIqkd+9hnx71FBDoO+OBPeuWR49eZUlpmZLDNlai0IQW9K6xPuypEW5wVr0z7/wr8krY90bCs4
bsenq3D1GQY1H+Jy6TJJOsGGbX9ZOrFY7y14C9yFSZPCvjmylidOKVCZoxMUd+UvkU5LTCdMRXYE
Kab+f0dSmNC/EBo86A/HiGwwWSnqWAVEaGtgbESctXIAHRn0SLoz9Nf3lMHj86iBCDNCa9T9NpDR
oxlMnOnbx+EDrpyNzPmxt7n6QpMxxpf1jZOCZCABVg1YI/AP8fPLyZdHbYZVLopIT2K9NDUxapl5
YXrGaxVMJUp+CVozfng9HBZUDAFYCi/Xj+6l4HVIv2ZWBm5e2ULa6YmLgvzcEE1afaSHQFBWf3Hf
9LZMnRVlA7tD+fePqHwFZnE6L2LsB2Ql/YfNjRdP3DHAWuAEqo2K0BYVify5WLDdreaRtFuRmaBl
ju2eZMEWIW8vICqvUqTKZrUbpY8frYttwQdrr7fxyJ/cYsBwo9natygiyIjLGNaxZtZKupG5Fp9l
i9TJCHLiOAZ6M9OtfsOsEXO2dWWGQtf3XlxWV2Vu4Jx+PKm/1+dAfreko9bpNX/3Sqrhj7ffXHCz
k9C/pkdZVkKVMJvNIDhiYqpBbFR0RKA+fdos9KMhE+8bmlWKPxY7Qa6CJW6+8R3704j2iaLgQmsY
tG+E4IfQ3VpM0/SagAC43WwANDCTHN5J5241+J6iZyLcRvcowY1vuseRv+a/SSAo1PC6exmf+03C
hm/JXvXA/+/cNqI7vl6Mbkz+ubIREhikLucVgKT6R+Ozs2tTj70RCN3yAVA8nIvhNfM36dOCj8Ty
ium8VChVY8hFbxz9pVK4ZZFW+ff9Jgt79TTiY34mt7VdR4yA/f+C7+UWXALgQ1Da+ZlwqFqIMQF/
Z1Fwk6mYYtx9O8XGMh2wV70QJUEbXMhqW4KM76LBvtNYAMAK36lu7sTUeTQNuoBp0O6betmUN7u9
QObUQSn+E9Cjz75JKXPa5p05QB8TzBeEqTKrfouZ6R8a3WzNyixHCvVftdV/lB10OCjNdzDmbL8j
opTQcL+9DIkpPQGC+/c5hdzHVNgxyloLuAR+udqqFhaVEWgU5tRv96S4ie6skwaX+GdKsElkhZi2
htZ8omHe1CeUMiHRJH/gFLWmaVpH4hLaIur+qNRLqyXNY4XV/ZHozUTnZfV9zD6Qg5tzPRqCrMpC
4oVE2P/WE1L3b9uITYjU1cr1L186qPnIp+wYLewu09iaFG5AMiXkbauc81XnlOqWuOwBkrj+O4Vk
d+koGVmjJVy8eqehqyPzQEKZ/QJiD7fqg1fXJgck8vLSSyzzqgpBfifMubit2nLpajUTr1gYlwEh
QXSr+i0RMcCiK/GkuRAxDzfeAu87AEfxPadbMg0Cm5L+UakwoDpK1AbEvrvd3ZQeGxHsRP7Q8lsT
z/lRDFqbY8aqUpMsXCsVi4rsiPl3Iv0G1tZsoqANM5zPzxixqbuiTT1qwACpQ2rbFA3JWrlOwSOn
iEapnSU70357QxtvPS0ILx/Kl8sGz3ABBibdQHRabNPCVSn/GUq4vzSOJcN52gzbrqvmrEcFr2Mk
aD3fjUlqXXiRwwAgvMf7PFmbQRj8cLcsyhhpA1wknxMB5pyxMED2e5ib07sdY7m4k0tDm5qNibjD
t+M5BOhKpNzs1Qy5GpHohrAkNji5cWYfUYIwNWrC28YQhlIALdysyxW9qChbUhT2YfoRcyGU8V+u
PO97EsyWmolFUwYLxjVDbz02kugTgg7mhF6NYdX30fJjXL/03Lg19S/VcYwcFi0UtwWgS4YaCHR0
OoOqCocikZnej5WVSREviEY1i8XxbSgs6zSDCVHfg8In6bsNfVT9fmGb5TYSviEz57YZfmC4ciRN
galReMoqORa0rTKFlTn/ItyUE2R8Qh+MCd5A2jh0buXlosNk82JQxoBO5mBHmNle2UV0cZEa7NHl
6NIzDzDSfBeWNLOglsINnTlwHLTWHI9OBLaKJi/CbxVioCDDfuZ57HwTzNm5ho5pMzwuE1FbWa5y
o8RPfrkTcS6GX0GgVqMjjULGBnOktACb1FrAYp/IkfXiK2czJRP83bfqg3emRQM/a04+znAAMu7g
hur5psUzApgoH/TzPBeGkS3qJ2DDiY3qTgVxmqj20La5Juj5atNDmmxLjUqBg53JCr4MvvOICp+U
lJCKLITM6yZEzfBdVxJ2yptHC/Xa0/2TIMN8IIomjOvkJ6e6OOubivmvXiGMIccawFfT/JzNg44J
KnXIG37V17rz/xw3H8AWLvY+YngcQYfQBEfyOCHbovQgDdazu9VhrWXq3w1ZIEKKjXU1g2EmMkvE
BGxFKf+Eu4LaPsnk9f3oqdNC3R+3V9NNG2uI2IFD8xMPpli2yhW65P7EXXKMt8Wr6pD0r2Awfr4p
hAOL37DhGqV08WT98kavUS+TwsO1p0NcfvJ+//8FGQtfCzaawteVLQAd0AsNwH6hpDojoRZOh0V+
ecub5zuUXfmYi12VTQcmlvZCUX3sTWeylwEGXVRgX3BYfknZ/dbBZ8Ayf6WaN+YLNHjBL/byg2PD
4jq/lgVsBEVST8pzcrgKEREJ3oqZHRKf3662NrkMjO9DJHznVfHj/WVSvVfz4kV51LCiNVhy+S+4
GakBNZmierlMVzOTDdSwrYHEg3s6LL2EwXGHgvgcYouF4nFkBmzpmLDrLUfiEkXUeA1cC7jrubDi
QQrfbKF3XNpSqR+CpsLfPcxKq26vki5DWHksuXhXOhdFy1uTWmo/f6WZqLk5PBixzvOHLGj11sh8
nmfq8JL5N1DADRjehAy/Bb0YErQGBkU6twnam5hHX3SAFVcFhi4EgQ1+Z9HY7EEi/EGTcxYaMry0
3bJLXDqiHDdFHcOLYtMTmv6jBcpCwVayqLU5IEbkUg3gby56kC4sjPeQIWBHAMt/+bY4CnTyQ2sH
EnWapdWV//+hd2+hN4RPhv37us4UyqT3b9U6rBUnhWsrt9mL3wfvq/Eh9ztbBvH8F40PNwBtn14G
BnFhDHJnAy7h0a6Wh8TcdOuIwOpXyrAwA1IZEk7JojCCM/AHQxCsDp8HzrQht6jGRmT6wTYlAO+k
Vk0Sriu9b/y7dwDwcibpDrX9DstNbgm2G4l5BGx1j3QYg83nILqa/X8Ih/Hp0TYAdzKcnMP4FBni
9GpyB9yxG1saaRabyUW/pi+8gnCcth94vc4SUV/uCD3uNHLiwbq+xxZHkNogQO1JqX3NVysft2k1
QGnJWFQbLXLpLjUpzXF64VBgrVZHuV+CfFuzlcgCh0nh3i4qO1GpyWCZ+5ahC9xbE8zwyc6I3uPr
8HgnxL0XjI4MXAXD0vBPEKxHs1B3CmdU9BUJtr4o6ELr2U/+h6UwRr0arNMr1pk82YrkgSCMVNkL
najXYJtNninFPw0zVXbhOri6qtvysOxTMbc28/tkEZA+170NmvkJpuHps28QX4Qr6TlfRJXpHT6m
P3iuTuGkmXna3eWvkR5A0g9dvcqrEhx5cE1gLsvmbwhS/nT9/LcrGP9MeRrlWT7bF2N9aZbrpASN
8Rm2ogq7V7z39s01HtrDDDcnVijT4ICrTUZu22aZBgWGDrE9bOK9F0tIz20YuWHkURX6ei0BfYB0
30AHlTY1ouQw1R/U5/xlLNXEP4Khf0XWfRkVV1Jhb+Z5VYcoMGWA8bGZMW0aT0sy9D2M3hEwYRF6
4fgemXWuF4BFPlsSL4azlANX1nWQ7JhjmJfhz4jliMMsPOhUzd/DoYVBOPf2QQhoX1B8B6X6ixpB
88VqX20purREHOe5Q5yieR+MNlXY581pZil9j6nnZbBiSSej4rl+x5OdsjAyjUtxag4dUURrOKmj
qe5b9bMxeCtcKa2LClXvh3OH9dkJTviBoBuwgQdfUlAd3/bYlYOL1EKlrQX+Gf9gtfYlv9lPyk6Q
/0lrYN2DXUSBE+/aDCuDnfYCmLiJ63BuO3IGJTAhijlSv5e7Kd5PiI7/yRHWTZcKCSj13mPxsl9c
D+MjY201+OhEYCSYMK2rpD84KM3JRujrEhFZIMEoKZxt5c3heTfr3MbUGCyilMYIVbVhEnHheZzI
OAj+U6STsyXxQap2KBUm+IJDvMaIyLEwBMRQEoIYlnJjiwBsw519Oh2LRb82pKApzvWscHFNXKw0
BWeKgFnIq0M4tHcfOl7UJhzZ+rmgqY9kiEvW51uGF/Iry0XhkY/Cyb/8v+9rAQSOoTts6zyejymD
WCctFACMj+Q4sScBewzjsZjZgbFhIOtwFADRdLGL1a4mQfHVFQP81165pPKR2z8HoNvpqreDsNtb
BzaQcUusEIbnSn0+XSI0MLy7w/CYPPpZDU4RPNUTtRHPM0VxqIiFKC314RgiLhlC18tZ8Uo8hxXO
rsI6KlhIO5orJTMyHJv87AWrjrAF4Ea+ILgV6b4nMkIzR4UqzKzRyetIiZNojsUL6f7FOAKhJd2k
f0sOWuAjdli52EVcB3m7hzUDvmhc8z6xTQenF/UBsv3Cy5fp1iOxUpjT1KXByJn4HHZkkxjjF5Z4
L8805MqA3+1Hk0T7A6GlzKv+ALwDGqbu2I4R3l3plLxv2L2B+7SPHf9mnoj1YX1MBSEAUFyX6rmn
eP3fSfHR2DQ1u1IZ0kpGTK7U/Ka1sKZgMe23jraeHPKxes6jhBQ4J71PqrrX088L5AwEacbpqzU4
prXsWpbI2fUk+HuI/2NHVdjLxR+LdaseyEaU/z3wevbd8bNuTxoriQYoczjtxJ30iH5J6k6/+mEE
J9eObHf+WnUv41oswiEZaSBCRlV5xFojfloms5v/1fOVUTghyFcwyfh4HJs20q4/2MavQyGVy2GF
xeD92td2IRqMKcmbLh4x+e1tMm+oxY5wd09gHgwA0CVinb8ORnzoug9poxUbDZXzeG+s4R+cVT7k
ZfRt4YiH8ICOlTUN9sJlQDAqAFzkaBdAF/y2d+ZJZJ+Css93G9K1H5LoI1ugfpNQHWmdjnlGiQk/
6J65rUh0fN+3J+Jvfsnoii67Aj8/b2HdAxgnEPfd450ugi1QUSO5WzraMy+XLmz7RP3FAgdm/qIC
KQlfGzi+3Lr7UDzCTz4TC+hARTDDJUt+P5UQg0jNhiXLGgCVT7mlodxs/Z0XsM7mVo0IbymCFvn8
u5/ENgVNcMdDsyopGiqBV7gQe6moWgJG3kBI2itvmZTsaxMGpPjRTI67sbZhGDTy8JzET10XNK0K
qdNAtOao2RWok9Cg50Kv9RoxNqreNlUChjwFIiMdvBwyf77Dz5lsCuXSRpb3Y+B2+AzXPgzVPM/Y
q+n803Pjb26JZLsQ5vlrDgfcB4wvw6z3l4ksS/YtGlfDVX/Z6dmqIVFF5T0H3Tj5wepyCHW4a8hR
Y1FdHJpGvN3s6/J+Sde842uE/nToheO0LrAeHjrGxUkQkAh5maB4xajT6ZLBei+uWgPOMB8Nfcpc
Kh0fn2oin+U2CMV9g4K+ItUpDE4ZGJvmkleE4SP5G6ArMURG6EronTr8PQTT5kDXIqTLKC3UROSp
JvpGmr6th4ltuqsH7+DoGWe26XYvKnIVxnWo/l+AfKf2c3Skc4stmhQXkdHG+SoijYLjA9aoUh4m
vDSw+paLRD/kqs9giVQ3Byp42rT472Aymb4+pa9pJD7JhXbdWs5sUzRO+Fs3Ouh5o+RRSNOPTAxv
hX8/Ya29ML6/vgur3BsVpJfzKjx5NsXhGkdx8Y7C2oONdhqRo9iL7z1B0Ex9xC+R8W1iRfPpscoZ
qUPo/jrwKIPRTW1UljNI7lODCAfEBAIBk0Ww4QBcqgmJFx8I2mHzGxRXN+D+d3qkxqibrgwSfYle
FbKrs/LjI1vDmmXC41t11ZciGIB2xw/t62T4LeJ5a1SJQfS+zVYYaT5yFwPQuUWph/YO8aPd7mXZ
tVEjymcj/AiS+U0/ZAqwecHPenSzR2iSC+RhyejcdR6uhnjpT3k2yT/r5vGzFVTRZwqHkTrckHkh
FbHvj+tAEhvLliEHRxDBZbuWRFMkxqPZTlZjIvgqSH81kHZAldDFOBsnbspTR5evMgoBooL6vzAr
0UAr+rW/Zn+RUgHvXpJWQY3QIshBEqP8wNSDOcIRgOcFhbVV2boTMint1PWa3V2TZ9wRuRsCI1He
7t0cbYpWCs3mXEaP2Di1cXSJBBz1Ash8xtm8BQbwvPbFmPUpunQddjKHzuAte6tATvSxoLusLF4R
WQ/B6OwfonxIcytXQZrD1R1kIcLE2H5bM0JvvZRkoBxeFcl62TBhjZ8XoZy3RzcjPXJhbnzmGRjk
+QZWonFbgA0zENKtk37fesxUn1oVfKeXv4fZduJhIzyAcFChhqPH1jGNKm2rvBksjnhzh/CfqQcB
z94Uoh18PS70hVV9UMkBWgt3dCl1GXGsfFxKqMz1FqsH9YF5s2eWlBy+SGMgBvANYdPcBtKQY66S
xrKJu9hNX0hkAodwycJLvEMRH1W58NlRVHRDcuWQQJJbbBxDxzwEnnVhG+v4R5epLM/oGTrtk++c
/A7coHseMRtWxirQdcTrxvAoU6jyU6oEEzfxFHrCPZoQhDHgs5WTLs6h0D9BASXyTdIN2a7yrEc2
RSjaXqHm539M3LD8p3otuqWP76bVKYP04v5Fd0WtqWlhne8q20EPoC+RyUrclg+s8hRA0nd47Y48
+RfajB3lkX0RDpMdF6q25S+W+C7pEJc0e1Kz5L9nivQhj9WxKJr3DWMxFbRXKrWS83bXr5LeodMd
5rdUVyq2ASeg4NusDf3L1DEXH+Xz7PVAXzyVeb2r0zD2GZnWttZX3AAT6kC32S4VSS3z3NjN6Rzc
oNsYoBmAuDlQpV0cJl7tm1ct6TKAcDpRvAgFynKsVHDE3syxK/M+F5Wa9x2zeoGFckNpkwEv4vJV
3n8avLR9A2dTjP2nd3QWQZQ6vceOXi/UlMaDTFvlf8RDwc+B/EjLW1dox8fnQm/xwnt7GgDD6xaU
ynnoM8BKFL9T5D7QDz5fnrDPr/aikqR8HnKBwTpFN5bTTFs/u5y0Ocd/mroL6E5L/Rcidjw/zfhG
NEQai9//R1Amyjf43v8YzBiPNH3KXFKN0f8Y3+4UwaISOHD8mjl5QT6pPXdPTaSPYNTF5Mmd9b8y
9ZTkAs/9wJFQwSsC3VVfvhlBo6csBg53ZOGYH5YAfyAtmFmipENXN18ja1W1YBXp35M+kWqXW0i4
1+nKGk7XzrZvYFq5d5Ki8QIsqiX3e731zHzCLzk+K8zEULscH464NW7TGk1rVDv50ZTWpLlxbMHZ
sglFSNKoSN8swKwNQ4iI8dei9RHH0VKDJYndg77Jaah1jfuAxiEjUA/5+SUfl5JriCzPDVkn2J8t
YvhI84tAQQT3KKUY60O7m4dP+7Atyt78F/ez757vJH9Jw1UfseETk0iG/JP8psrDiQYgwe4tuDpF
iRDwMhuDnYQheQl57xV3erO3etNtAqX0hnoqiNlKMhPYv9AZG/sGhboqGOIT84SBrWgeSsVTY2ra
EBj/iUeSXIXv8hCnjVKrQV7KpdINJ7Xt+MxvVr1J3YvhHJodvln+zCm6E+zIt+s6ddCnfI4dvEzJ
akTMtncJqj+zeN9XONwgtlAQ5MqQ31YucQwVA7KisSFnRmMXi1wiEapt37XcaOUuMP+D8mgqcrYa
S7+V/aUcZTuQ/Em/ImHlGn3rN8UmbMN/9aqw/LVmVNG9B1EIo515gas0gik2CDS8MR2MUZN1ERde
u1Mw8Jnl1TuT8MBhpc8iNtANwsBGIopPmxtgiTYNBpvV/5is3i6dS1I9HchGKB3UgusMKkBqK3MX
7Bf4ma8A2LXe++GyIeU5ZnR4+qgrbMjnGAuK7XqKMoYlmuWUbwUcFMlPkEGtGP2Kb/WnjqAh6Pxu
s8ELSA6ZL/pWlh5rNZZnTifL4Cqx3l+WWsIVpklqo34Wa+9rUjJjZPU9IGel/x1lB97sCahqLKNU
KAMcZ4jjTb9TXhCJYtCfNde2Gnd5+2OU4lXb0SfcOejvplR1ubAWjZ2x9tGzUtDGXvS5lL5FdIXN
FFSC27cocIgp7fn+SVA3hA8PY0N6Vgc22M0eBv69eeY9QFg3i/nPQH6kOYHjRCYbw62YwgI3s7KC
v0C9mi5pgYSdhDUaJzRSFOfMO1oEYECuF3TSq8kOmxC8+TE3jcFsEzzu9+WZbE/1/EdGy16TNpPh
pHuAi8G+i33pr/9WfnpomGPeqm0ahP1hFo5/rkuuRWY3OpU3W0RcbQFOW36FQxK/9OerKwGZzekU
qxKoYjun9s2nLcpF9NVBdTH0RUg6F8Catus5hoqfD8yKTlQWlUrkB9gfjcsOLIHI/722u2PkyBRi
Jxd5h5VJ7diUKYmEaZoiSVAvRuNCk/aIJfdeDLALmVh37WREj2JfxBrHfIlveSYxu/JUoGrc1PWg
oX1bF8FS1M8zIaIjPe0D97G9zWdH76HshLfKed6d6mY5uk1jYPXREOr0uxQyt+YO147ZspB5AeY3
QOHDnbZfjOIBy1dJvIav2orv2oeGjoB3ZLPHTzR+BZfIhVdJgMxWMXQyZwqTGHGtN7rX+KpZRzSL
VxTp5k+6TAu86sbEbqXATuONeM++oxTDNL9S2b5hHXNyt/spk8YF/6rD4bR9yviZWQpsQQDQ13Tb
W5KtI1b+lKn42fmu1M/XYT4BceIPi52qAdH2aEDxDmxskBEsQfqEPuxBW0rrxGw/PUf43+1AOHyu
OVE9LgqsMyE3IbPzRQUivP7MAp8DzK6WoUeRptvDm8sWAZKoaEY4eo9mrn4euaac18gmbDeGZm4j
WdkXuaeTla+tuz+lh764dN1JLNIoLARGKalbHSzdw/rxsYuKqHJWQzcy7qfPiCQVkjZrwVNVM4xX
72l5Qs0CM3VRgjD1u73dWx1IeC2776TGoCpaDErQ6Wb2ZczorHLvGstZP7TgFpRm2Js7jmm8O24+
QaUoUa3Sj+l0TG90o3rPrF4OtkvCcKHQakIE05wfKnc/arttZ2FSvH+VZTjOfkT+xachC6LIU4Zg
e83/kWKBgfy3Qo+e67vzQ/+Q6q7IOcE2XKOcRStJvZ/f+ugIcrq2sg38ChiDwbq4YPVnJbjh5O2Q
kNylLg7jGvn91K3QFabVEs5oQLZytvsYbpMYRywy+w7rXNoaOeFvbC5XHP1BI0HHXOZJJO51NNeS
jG2EeUx4Qing3X+5iNc2GNosBR1tATe7S9NXh/vSWWhL9RXwPrkd0CDBDOC6VBjuDnP3Wz9/8FpC
N7AUt4g65puaJAtyAL0R0Ls/4klAKW9w6XRZ3ImkEttwheI/u6en8k5Q3V640pg74EIfg9mZy9tU
j9knem6NBJaCCTGFrZHQhj5WnXYyFjSk/QznAx2MM4SOAFyVSItLgxHkYLTIzNYJ5gnD3nv1gCFm
gHPE+DIJTyMQvoAuV1I8MOyxBKWi7ENYqX2WZJNA+wpUox1EU7oxZ2HDOaHKLBIcf4FS9cNrxLa7
VbNCk4fknOMCpLhVnlAVQML7V1aMQesyNuQcvgLDwtlHCD84xeVpc1HPBHyBSQYMzw69ZAQK+vNk
2vTbS7AfKcxAqA/gBFJ2wL7ucxLwDZSsRm9Coqdsx749sFm4o+2aRe3RLfiViag72q+NAFoyWZ+x
0s5dOlYylDezu8XnOr+eQlX3kMQr9YkyfyIuRy27F72szlltDZcOKGgMLGaMtayPOfozRG96BIKL
NRevlgotvRIrPj8qJvU595lnIdHquf6L84CLFv6HW4/Id0C9MPmjhy6VEKhy7SS4c36iSJO9bgsW
IEYY8dQrvUkR8PYzYXaTBZD2HJBj0NBzQBaJTg854l0zjig+V2XxFliIkUXND7Bq4+YMGRnJgZaX
bwhuFASRHYAi9bQkU0DvF5I9CBCwfQULupLZ6Z6aXJIYF0EBDO9wXhfTDwfhzryOmuQ54Flx4fH0
O1J896+t6iO8KGHD+uRi3Hil5Q/w/G1WiIjd0407cZjlPxz+jv/49JMVklIMdgcHHe8U1NFlUOJm
zaPAuy1oJsF/pwyIARjeJaPz8esTXNhAz9B+T0R0FBXnNzWFX/pG3QAacWr3LdsmUXNd1K6kHcNM
x9qiy1/ieRAz/FCj+CiJy9r6y/HIYsprCQmg3UQ0LsvKSlr1EDa1kr85LCUlfMfr0aloATXbaGdH
eTwLJi/1MZeR4JfPo6BiQsdDhNhoOyXaIVeKzBiR33dYAjkbzaLDFtn93ZArOy/+7t4GV+J+hLm4
DJWXDkEMS0sN+5YaAuqOh+vAqsz20reioOVooqwO8mGo7Q5JdlH7vEgL3DoRgz7/8SCKpZ9i+/3f
OdlCVPQHO9W8AgjRYBWw715sd/MUpueC9WnWfV5JVewo+3NizqgXjXMLoc0I6w39SVds5Ow28hzl
aSxA9bbktnmO/pjp0P5Wjd7bU+m5BdV+2/f6ooShJcG5tz2nDL7WYGLjJD21gozilTpztUcW8YEg
Zr0L1J1hXNei2ZItoPVvGpDSL2Izbf0b+gkkWJtDpYH6Iu/jiav0mo7X6DzcPQB9ulLJdxjYLHmE
Y1ThRpbZASBMqEtrJG/PTdmiRZzsKHagdJyFzHU+JqEu4kVOA4YlPo8eunwjr2m0R/mfWLSzXiie
QekcJkh5iGJNKxTDhaPZfwCYw8C081Soq1irl4fOb55OQzlY3FYSPTF0XlixybjkOqUpl5AFiPIX
zJP+FqxZoelu+BZjuZ2yaDjMJMw7x1E5xD/KNaYvphZ3zBBBC6VHmlnt7QUwKSsab0AX9r9/l17H
gsdV4Wq8jjwpVZ2i5uNcnaKrYrc/k5PZLigjvheDGDzrJBp67W353YRzqwey75YghVvr3S7g16IR
mC3kxpUn1HJ+DYNUrw2cgU+Ven2U0PHC7+1wQAKOBm0Vm7DA1GRodDTRh+ejsMNonF3mJm+FhA93
qwoThMTu5XgSXz7hD2H6/0do1iYL9tT1wwiHUAlXcx7zUTFPxsGIQDLQqcQmOt7Od6kKrargjICb
RVOOtZLF3Uqx9zEmRHrw7t8jDdK0nCMhdHW4XZpM+vVzagjtNTFCxGo28HVlEFD6M5lxVMn5jNTq
tOjmdSxe8j3JHJclwmSwEyTRNRFneENRXB20jAME+7gDwZaCRQlVM0h/cilnp0gzmigVOVvrWXFA
t+q/8F+lT6cyK+w+O2yYF8baD46bd5Ohqi9o+CqTFa3INPwWY/SNX8l1cKj2OoH6h5IRkVDdokka
m+biyKDnoCf/ZxX+epUZjKITfhdZQ4d/DphhdALtIo8CLYP0UoP/lnEdY0nG4hweWg/vc42usxtp
5gq2WIE9G8JOSue1xkO/etJyR7froUyZ1w4lDencdzfw3ssCXPCzE7Aw8rGfpFqxe/7s52qOr7sS
h6yJswGENu4abeG8Z8jh3Mm71Wqzcgcg1j9VzCMJHZI7namnfdhN1hi5M0evqEhzIGktJ7Vh5yUr
uMu7uODUAx6yRKH4GtWrbN5LmfrfH5mOn6HhNlE5DokcvdARpXB27UThc/HAaN5XZW1UExm6Nhtd
e8/xKeFuv3KbnBrCkLthNWAwlEcGdA6J6znG+mD+QK9FAyYkOO1iTLjclxk9iN80KuNrxoRKTnFf
F4BuSGYpYbulAqSKNNfr1Agt5lZUpIAJ61WYsMQGr40oO7WJ4Y9vj5ma2QszlokLyzFZkMmhg4yi
CB+E8jeWVQRkcUcVOqWHH9UqJUJeozhEMwq5XVvI1+xbayMI81Yb/Y7AYjPA4fUBjhlsU0kfI1p3
5tcvI8+myNGGzYxXumyjX+3B0RhQ/ua+vG6hoNHQeYOR3HMmQ8Pijtgy2E2c5bCjIVacVghLZU/e
v1CDU31rtk99GIWmsQCE2lnLz2LMrphuiDYeq9xkofoQ9uvXfoM6budvM2QnK6lRpMX07UkpCTL7
dts9qK0k9u/EzPsCRZQ3uozOfR56CJ2YDZ88SOFbEOWGVONlWxOa36YrWB83zV+T+yeQYCihLK3f
M8HKvIMsR4Xm4iV+0efcmYrYWCneVF3OzskOOc0PA/V7bqFm/R2YEb9EMBaFTQsEyvbNv0hedvBi
2Ewxm61SqB6V1W4023kSHJzZHfFES+3bbBCPIerzaKpYiTg6eoNlKCzcVzqHVncajj85ZPzF0XUQ
IABH+gG2d1Pvi2WpA2F/10OQzmPDL03JdaQmqxKiLMWpkxIjqssiMNcpY/5+J9FQUE5RMeoH99eO
TEgYNEj/adWX0Fh1tFtvRYO8ZbqVU/Fq8TZnRVNuPvpaB2FTQ5lpyctVFVHjuRmH7i9uHISh43uB
MtX0APK4iqA0EAzbd0nfWCiS+mwujU6jScSUV4sAKDUHGx6JY5M/35C7Io8p0wd5YxK2s+VMro2O
+3VExIawQ4WsPI1cHAxZTT8rRUAdSIzJEbLScjvQNnrPs4inXnGWssPPXGT2sneJmCe0dpWLjt9H
6cFOqNEsk1XbNCHJpOpeljJSZe9Xb19laPUoig0CoHm8y+ApElZUQ4hbunWMqZTewV6WixVIMfiA
ohppP1zrA5Z/oXwKv8JgDYVdrgZAV2eMmVWN2uyFzcyhueFs6pcOOZStJxo/xPniDhrZizDVNRek
qP7uhicBF9WWQdIkMyZ1CCfQoowvidCrtxY1PMpCExjayMlTaKP0Yawef9HzqbazYknhpHPVbNqB
s/LMiGxq9WuxZFQZHJy8AtySefrTmaUacX2iQ4eNmGHEDeGOPYh6NIBirT5schdkFyn4KRPQkTm/
2fzhTVBCoyQ/m/A89NetvedCNhZ9K299+/z+wSR5VEIgUzsksrRek8HA0f5ZZcvm0IVgdFlWv86u
mqiiUGK2dJKoGZqo1qsV42b3Zdt77452ESKAKqRPfX3xlWrCDMsSEf7tmjRRSZHydumx08gPK7rO
+IkXByhyMsrRX8FoDwW/w+QRKwCqqmON9H0uLGV1NBiwwDEvLUf3hICQRkgo9K/dIiS7AiVviXrU
O6HPXyfUqY1I9zWqtXb107s1/wywBaHtuuDyZZKYGIy/KZdsucVAQgcmSmt4RXwILcn42XZSboxH
8C14rmafYA/iAtrpXXDtWshQ22kIEVe+dEj96H+z+8fbM0muhUAe4l1gCnV5Cjuc/yF3vB9Joowu
RV3y/h7gbtkksuy2Rd4OUlQVMce5FPDmaGAujdsn/6OQ1jRzg+If9jlPRss/oaXLe9shVuMToerh
aEt97I0xh4aQ8fmbOH49lSmBpzMB/zAkTzMst3lVNEd69nhK7HP0jpV4TKgONhsgRmz2VpoldeuG
UYASQ4UkEGACVixhwHkj2cmAO8xfxunaepu0TBgXQuSmbd4t9xFoTd5p+c1nTEZInj4EWFnYOKKt
OxgcPcrSvnpjQEUcYinKJqBO+kRuhFpVIPcQsdUR1y1pWSJaofTKSN5SFFbsnAmGtfmdqHFtbgEk
Hrve6ux8ViHVyBYMXtX7TH0cQeMCv+091Ez7HNOY1CrhjXlLotKaxoKljD+VmjWRMeDnQklQoysw
EOmkg1QGZaT4LzCXC3s5PTIAgvPilVTL3cqfaaKoxOVX3LedQUud3YA0x0G1YPcXpxnbp/WPUPWA
T+GgwClJlwILeVbplVbYgTRhq/r0vJZXyDDciKkvC250iq5HALNf3LAoYGCNgO2A70QLdU4XIBeP
MrsuVTw+C6Tu3Jq/WrKXgu7T0X4AsZZfED/Y1osiNWJyQ95ekbfFXMa5VW3IEVSffbcWv2fGieQY
dIkunbD1em3/1Cyfe8Gqnz+wcjT5LrHpy3Fr/Zlt/0+3Jq0I+nJg8ecjbKPxqE9RvuJ2Dd5zvDHO
J/hIyj+tXJTJbe6fldkVoeQQvMHDSh0gIfIRcSy7ECgQbRAy1PGUpeDlY2pRLiARfdkUHIEBu0YK
v8Mep010U6rE55V+wUTCQwJUTyqpxWd9VBizsA62dyRZJ3v2IJJ0P7INvf2ODiLf3wxkX24eMPTP
NhHW4Vc+tHtCBC+X0ZsB6AH3P8nSXXdBQp0mDTllffKqR4187BGlMZBc78lVe/DgtbdRz9MNhCaF
apKqnhCnPRBBBpXIXNcH5QslDSonjsM371zxbGiYcx7mfG7of/9argkgqHmHc7z4GOMODkcvYE+V
kqAk5FcoQ+E77ha3ZK9a5QcoSUHd9P7OHfkz0Hrn6WW0tRCBoy6ARlZcBUnGvPT1zMrrLK5BK1y9
e2PvfrhDhQrHYtUMro99CG1dqqBr8dNKB9ga9XY2OBASdmqcydAs4EyOEzPzFK6YgZaPnJI4wWyR
xEDaXlqSDIBc83SqKZutV2xVkxbjE3M0R5Q2Tk+uZN+0N+Dk00goJxz3Pj8vIPqeKO40KRfkWB5F
twn2EqBxjs3FqWZIme5K8aa7nsB++NFkPURHKvZW9fS+HW6ivtY0+gH9rePH/4bxJ/ZLawp4M+tz
o2rZfPVR16IB2YCTV9hF6V+lM/vA3xP5Si8CwK7g2U4tebE8xMl99YLcok+HYNNjH0UoqZXQ4Zmn
gog77bNzfmRQ+kHMeCPW8gu10EblZHZ7cC5xdB2UhV/OZqx65oz4qSjDvASV4q43y9Kx2qqZlIeJ
+M+PU3PVMPnio68Mb1qCi8BFDYD9udzMlNHXiEnt7rLD6K7vy09lqPe/oX1A33bqkOpuLTTAP9Pk
V2WF6DPBXGLqIycyinGw/8TGbBAfx//0Eo9Md3GAkt1cgSJ+AvRG7zC7u21SQCLWUvgSy5E4fVka
Vo1ZTPiGo9tNsUpgrZD63/snlRUZg9/DNNW7Yl9v+CwHeNmG8an0lXMnq9tdUFDzVIqJJ9K9gZYP
D8MKaGtzp/9y1EgmOhq0aYX0el8xNfsGqfviA0W5qdrZjBB1bvK/XW0ldad3J/vnfO7zaR+sNn5u
wt1o8L6SYbozp9w8Wa0+00HdMMEpxyaG8B+M4c81WVK0nUsk3zBlJ8i/Rh0BSUtoSuAtcdu6qHL3
HSXEKTrAO3pM1S0Haqj4ttwGUTu/qOFTZ19btO1+3rjAJ4k3bhQJWvmynYLA2KB3KscY4LnKxS45
peKFsahR+RTphoIiouj5/9ClmDadTNC0jX81JSiKJATsds/T7g/+lmN5OX5oGgS0t6KiLcUTP+mV
7UF+eAt6KnZ6UNbKYvpKguO5N9eoztI3KbiQ3oU0zflahyOBLA0DNn/bJ1dft98Rz/PqbAbv8Mey
Jc1gMrlhvNl5zVtapaIdp4Zg0fo1gfMe9RInPDaYIsDgoAj/ppKfa1azPXK9hohyLw5nMFwfvNT/
JzIjgqNIWtASXUiYhNDXwK2SjnMj44bH7PT7IEhBPGU4Yg4rwuDyeaCXWzvfE6G79IAnVVQP2tl8
Z/mDSS9iiTMaUeDSg45Q8Y3PBJqW6pEKpeBNMVwHFSo2OaCyv347Qi9xv0nfEXI1PgfyUOTGwsGL
WXgOrH6PzT2hBGR09MCpdZl8140PMzF3Mf9GM+tMuKa3gRHN3xe/5rOMWNfMTwUZNLFV0eADzVNW
ZMD1Om5JL+4Hjfzp9K6ETypWfq9yYFA6Nj7tCexAebLYyTluGNTIlehGPJqycMnZfcvk8idpGHNX
IeRz1X40W7hOg0/NduLPGqS5rOwJRm4aulJQVUeMQLttyq/8SJMfXCEZVva5C+OFjTUzeeibnOz+
HgIYTBKZFZeHMl8vPPG6c4r5dCVBdBBe9t0sYI4NXBZsL5TLCadmZXcssUhS8ANGsZx+Jtk/prUe
QKd8Xi6A5B29isLoUDwjLKDcKZ+MO8ZAf4JH14iKq3sOjfrfoLhSsaI89BlmQS0Amye+GHOrtYSn
cCD/QUB4o7cKZ6bBTOmOtBe51Q5CJeAT32WdY/YKh6uOcEvAs7JqZvMlJyIrEEnmSsjfFOJECu26
TGAE63ffOHtF0A9vUn6f+5kL974HEfh4NmQ6arL92xBO3DPpFPvEB3ZqSzfpsRDiEmCu/BJYXR9X
+0vvxmWM++g9luKoDuuTtkFEfpfX1YLNrpIZHrjEX9PS+SOWIrdTDR/p38p2I9pEqqZBsBIYUdDn
qX5Kp1oC0oFVtH/5NqcWnf0HscrNfS/5eoYotvQP+Bsc82bsGlj2bwrDwUh0munJdKKbFt0bcQWk
E13ubfZsTsYpOLnLSHditSPbD9B9kWHKNALXknFogR66p53kdkeTHzPgOrvEMgbd9zEccZ9O7e56
sadQDYIbi9XhOPeM/7GX4q8SZIP9Za+lJ5Q/ZIHd+6UtbJBpBVN6ABXj67GtAJaXR0WcEYDx/GEx
faFW5wWosbrZEUOABsOfyPbhkcE+sklmPQ7JnWHd4lqmlTixCq6V1/ELgwYmVIYFcQgYbT7273XA
I/BXEB8b5qp8lASX+oFZAvHOy+ckOXHM05hVGmtJQiGyJAkJXua7yBxiVNVkFXlkBMNmTIf6+ay8
WY1BOLlufEfw+CxqAnO0Czs56FtZ8spxn3qatwnkVijstjOvZG8CeIImoDnblZb5Gsj5KbLAuh8/
THc7HHlIjJ/PfBvIqgcl6Ob5cua0ZFqkCwWImJwz4iw1LH2tGaE8ANMmaC4h5CdWnOE1SBJtbegk
pNCFDTWzojzFLL14BhM7frMfMwzBxjluMT2Z3g3Bv2p5OquPob01Auwx1Vyxg+vn4UYtjLWKvQy9
Ee/hYiVIQI29hAzweFvNRfKgf/t7R1zBZeQiTgVMZeq9E5dJVcLddJKDz194c+yGY7+oB8nafUcZ
so4dbRsSOdTMLzPCPVPyXjZHMJbc5VS/UJqWQjYXuA5OtiYAEVFp5nDkmntiTCPpYTfPFJVIpAWl
6dvKX4hXFjljS/WriEBGuVcwMGGTzdBVNfdyNzfRFgqtCPvwaEZG8jqz1NHB7cEtlKhWi4RNN+ke
qlLyKYXGOhLthOYmLP913JLXn0ZsfU9z7bs47XGWII2yyOif+5o49AKCBI56/CXmaKccnyNS52Fx
Z233E04Dndu5c8ZuEDVX1EYJmroP1my2cdptMzrHk25YW+G+ZcTnqcxungrs1H2xTseNwX67Op5r
BRx2nZykCbq2S3WhV+ODLPcHU6VfzaYUzyLg4r8zm7GbKsAkWhGy8BuEzjuAHQVIPGyDCn5gyhVM
PY+yLeWBwwkCyFgBoLQOcojYwaWvnCLNXu5MfevsnEy+JVqFveSd/cv0cRQxtMTBjJns1oNam6Pd
FYkMgMm6Clj6KSPi0Wf9xwSqUJbf+V6OE/OnnaR7yggJRGnd/17kqS8nLccxL53bj6M1oVZeD4WM
kGLISK65SC/AYlo5NnTBO0YUKuh3sv99szV5PDgHUvTefMjjPVjddDkcl2GbGgazmqdxOatuWr9A
QILhsfOAFXnqWB0IsVRSFqvbQJ5GrD6MyxqKwS+2n+1GAuExkN83z4WpXblpB0evWCNmMr61+N0t
7puH+n8FRk+yayB4L+wSQ2GpKo/FkJt0ydtyp0ulVIpLsbe7w9V8xvtuif3DkQIxQpvVR6+7aZYU
8tjf3OI8KPgHcCKfOTzG6QeFZV4Q7NS1/SVQGRY8gzFVPNlMR/m+02CxUMrtDKRg8XjUOMPXff6A
LMH3updG2+yz3BSPwDcxFsOfdWbVl4+91qoB8stlxEvTvzimQDaNPvHUXBJ1Kr8U6YbZvYDK9U2t
gkP9LIT7fgDWzYoWoMxJ5y1Ew76kNlPBMngfKziTqR5DqLML5cQElcPF83Loca5vZunX9jA+fYoj
T46/Y7PY3kLLlwhSUgB8R8Xx4tOEMXZ+rq2Hqbyfq+sdKRxOXo3TKxrjsA+4NCuwBfcusXEcFdID
zLlyOwua7gd3PK5LFfVfEz4HeHjDa5NZpovdJYc/nNZ+x1DQ3y2+nAYDq3ulvISQxWzgaaVZMKZo
l/o1446ck4RudbJMLNFbnxpMM05QpVHptZQdZ2RIaLUin/8gZA47ZYy0q++tx9Bdd5GmyduT+RYr
b7FFYiu/7vC+CUxWPtRQatd1+k8/O1mtPEp2wsicYP9JQ/dcXCXfpF9G4wYokA9qeQie1Z8VOlMk
dPPovFlnPRNiG12PwzMklJKbiJosEYexzlF78p/MuYHCMeaaRIzNCkXz+8G47KtvIeo7tEbXolr7
Z/ZcPsRMo5ErLZ14n5k/PoBC/NgBv2lmOi3uUdgXUiYjL8OX8ycbXbbJsvJIJapQ7vP7wqDdzM0n
X0quTdV5lcrxrSscsnl8+hTdT6/vfcR/ooSf5uVHVye9QTUpmZbfbqPeYPmTkGvqTdIoecNtPv0t
WuMPMxmlXnUAwzmeYQWwOx6gezvCDgUl9a4QQjVAAn8HUnLf3PJYV85WslfuITVBjrsvphcMWRmS
iXfkvEU12m8aEx9RRIIwUsYjKu1m3AlRo0VC07M6eTGQSpverluVCTQysl6lK+GolN+xie1JjnHj
l6h2GO3ec4kJDSXjD7FlGNFoUwsOMLrfhDZ5mqZ5EpGsGg6zGa8+CLc5WAAmv4RrwnMjEGDNa0yH
cH+ql0IyvLSyktgzm8i/YKYHiLvBbS0RZVf5sM6Aed2c72Xi4cPdMFf0SRxhfo+a07/zyeLfFZR2
fX5TKY943T3DXoBRMaAGEyAQLeHyyv9oVjxO6cfO1UZoQfIW2I3bCjD68rKwkX05IyJAA+ue8F+a
Y4pwjJMT+XOYNt60sw0vogs+xFFXTpFxsuPCoDZXrrIbcxo4i7R2Bx250SsvuYL8MxFjuWoI7rRh
teRtQEwYnGh/xY9YOq0+FAuKTocdNXeNjmrwf4DfPRS6iyLgeGktKVJmcrp049I4ELkUflrhMPZq
uNuiK98BKbGkI+mYMce6JysJXEv/LjXRzXQqNl4MVDVt9AAKbcm4aTRUkKvZBMFjbMFh3dS72xZz
TU7g1gxfDN6IwWgH9zgjHRvHML2zytg1eRyJm2zTVJPdoT0bJzbPA+AhX1wUSylxgEVIaKqEeNSz
7jH1BtwdvzqwkCt1nL6fdnk3OGz3MRBH8785760UKeQE93q+vLHiYBAEmV68ozSkvRQWBxdLWCIw
sauTTVgg0zr8RTrgo901/EucithP8cqu9o1k3mwXC3NczC5wWCRhG38elyXNjvV5Gi4PbDn4t/yk
XqNlSsr1D87YHWCud0IaenErzDyCKEN2L/tLbUMC88WJ8d3vGTpEHiS7ajKaWNh9+KcqDj42U2bN
ooqtS9H6pwn5thw+aKRjLnWHCg2NGPg8Dm/JNzWsLlFAbT3/rmOoPIor/eo9gP0mN5Y/MO9RaXXB
KkN5KWe/vWbV9mSya/4eJ3D45ChqYoEaucAYlTh5aGereiTILt9m+e2SDhA3yjE2Th+ebY71sBFf
7OwuBw7Zm7IiCArDDj1jw0QGjJkt6ziSu7E9Q7x9mleqVjF8KgLGoT7v3w/K5sQr18Vx7TXwEybK
Dgaq8fViUjCarAsYRUsxAIN+7Nq7bugdUfBFTNtGGGgfhUtVQ238CwNp7J8Rc5FGh2tI5Fw7GU4s
MCw0CinlXhJJEyLjbFhPNji2kmHOaGI8A5XqOkeXSmStUJhmbppEQNKJteuQ8APmuYkOcI5YeUwW
+h7hGtmeB0hbeKFqOzye6I12rVkwYg688N/59qZzG+tVYd9Apqor65hLjkFp4G3Y1wCwsrinPZUM
eh0f4OHuksB3XtSTKhnGVRZTKMBpB2AZJJvsYC90lgfejAFd2is56gmUp9hsLqkuuHRWBr8Xj8e6
LON93i8fArCYo4TgZAWgu1AirSUyoJDsMwQ2IosOSj+hGsZFoYlNydltlJfpqaw5gMLEPv1A/3So
HLt62xuF81lK1QUo9zG/Sy9HxFLhpTrn/VxCM+uDN3rJNTPf5dLhG85CYHUW+12aTwDvI7ea7HQt
FIBed9rhDiFo216lrLZ+1lQ6I4OMMRizd7pSZnPgZSqx+kpuYuQv3Mui3uhNGXzmP5iq/+Og+Dgz
s2Gmmv3WPXHkOWzOgYoSGDD3UXfkPMwOTM8lXKXv5g8zQUfsi7oWlP2TDb7XwZ957gEkZiqvpv3M
xbdATWy+0IrGFILDhNWYA4ag5Q3vOeIlcHbeZ3uX7e4KfHuhI3b0ABJmElLcb6gvjGSQjvYTDzaj
eno2oMHUjZHjYez3PGE899FuxnVWUWXT4GFI2HLj5GGh43+T5OPyaqr14T5imIISM3koFU9SLeGP
lIDSwglWKwCPM9TiwKLRboRXe3Z6SzVHT8WphMwiBqHzFvMQzihtJx23jcXkcyrLPLjrgIne2yDA
aBQWRF99FL/qCxrrea9H39wYt8O3/I0B7nX7q3EqEqtko1R+TScYw1lNjKQQCZDi65ALZ0kLe9G0
fgXoS8F0Txxz24fdYh7rf3RdRyBaRVtGFakBH3huyCXfC/ND7iRQQO+hu0qcU/aif1cRdhVAF7LZ
PRAXPc435EQYD1phivU7Cl2yhbVd8uVSghRuZMFMHXPxpGBL2vvMfDgQKUyP4CncHNKwMUTdPCcH
Epd1ZjWXpbA46sQGDC+uU0ufAJ7QEyLPhhxQwEkwSMbrtNuK/kn7knE+goJMmm17WMfpypQ+2zSV
Ysh1ATJerbx6ruv7fF+vDt5824eq0tWjEDHMMdf0qlS98xsjHdraF1DuJQyRbPlY7dAHPqw3Ybm0
GC+GjcXlWXqnfYlfNi8/H1KR2521tz5AgwlJ9XZK62MPXWFlAvylj5TY7yzN2CNyIBz02eLaxE1V
dTMYsa/Hb6X6l5ajoXTSH5nj5xOkPMpAJIsdVQgeZtgEVTOWb0MS8y62g1dKzaMhPUfTGENYJ5xe
TB+1BtFe+z9k3ooA8or6+C5ooDY2s/ztD2K5POLtus/hhodtOMXAwEOY1cKGWFe1To3Ct6N/C95G
mCIe2dwNCO3gMQTusfs7f/4FAZBtUf5xd6WBRLevmQSBFamMXkc3imnZq33ekSvBgppja2IVWv+T
l0JAsy27G8RkcPOYSGZyX8046Tu1BDH91tfFp01lbS2tF2zTUI3dvaenI7/NkJ1rNf+pIBcJafBZ
ErD+2PIIIdPKbQY5pbjkWMW/xRGJ9UovYKaKaILNtSeRE1O/I3c77GFWQ1RNMENHA/EH830T9mOC
yKz/qyDE7tC2rczOh7pY7b7oZhNfwAyR4qXfiEvdtT6cFTB4O67zfaypAgFx4uHs7xKzZM1YhIE3
27AvtWFR5M4hNm4d+eOf+6t2BJh+cptROwVBqASx02FVlJDarp7ZfbMAZW2hZuaJrZw5YKrFzuKs
d1Axzd3Ufqc49pEFM8D5AdgX8nwlm/xcO8JjPchDooS3O92vrB4pRKP7QeXWnWrd6lRovtncHnBW
JOaHvYbVYtOBYxQTp4DXMNwzlU+S21LFtX7HXcVxDt8Ql7K6O5G8qAnUzztRi7PtOOGyoNf7P3lP
AHyI2r+TMz8X1r4CLbDSnq85+mzBArhDOyqYUd0qFTGRaE+0rxCZpGLj3DmgcukyOjiW6Kg2jvbS
USVL59+++/0HLhU2s0FCt0ddRA33eG+jd/PBToopxb5BgoJBoOK+GG+/6wZc3ighwpFXY1rWrV72
ePN7gK33Ap9F2KKQ8lLMmdZbP+jrrNkvZ4Uu0/+mk4MlCX5T6ZOUJlR8B6MbZS/KWhuUU1LDgy+I
TUBCKBJ3JG7fVzbo0n0vcSGs3+U2i9wCUELbAcJlvaK2M6CcaytXM3d47I5DiknTVZqHtgUTN0Qc
KO0afjfDSoYEOLRGwvDMDX8T/Kj6ubI9wG/CbZZ98Q6K+xqxLuyP5Vj2a71r6LFhmDWV7oalx3X1
GwkaotrQo/e/GkzKTziLJatuG0ldZNmvipObsDl4pZ2iK/7TGGJYu417j2CNyr+uMoIHIKdgjtpr
GniIvzNm+WoNcNPfe4a11yqLDHHsmJJWmet6Yiny/VhM78uFMhDMamuu6arf6N62mudXMPOApPu5
3cPehVshQj4Wxr75FsSBC+KMEQ4W4qiWMbdho7BcE7efQboOBYU/FSH8q8fcXZ1dTxmG/W92zrCr
zsuyFAgrHKno9AoUvXazwSzYxLCGvarVbWwXIkwJTk4LO84gV5IWvMWwHjCENJ5T4mSw5i6PoiNZ
Ts2luHyLtrzX+QrT21DgjUsCFtKNX+PkHCKSPVcW4kIOpBEfasm++6oPcfsedNeoHeG8A1Tnk/zX
3VVjRo7CSwo8CuXn8J1r5QvYCuBAVCAqQOJU1EgUTfUBA/EqSVnbQeGMqLAdtTyArToeTWtUF0Cx
ygg1MVv8n3eLK5m4bVPb6JX85HSWr+WIqikk2ZJQmn9IHYbqzG/qQmKHHiK91KSi39bEz2IAO9mK
3CYV9QpHEpamvKHsd35SH24u/cVFXWg4Exk6HqvkezalYVZZJl1GW4l74iE6xvYLyAPLhezDJ1EM
J48JHHBR9GsjzOFyKDoojxEyTplfI7FjZCw6xru3xK6dPFmCk3SlT0nUi+mxdX55xpNtkLpwVfvK
FdM2H0rTbqAxG+CvLj4b09FvEQ72FxAeWXU76VDQamTNjQCjYQOjRlJljPfk5WmwPBwfY+N4cfq3
oVG/zfO+NCQIO91hdZDl1PexttYex7vpbYSE13hvWmkgCDyV/a/ZVXiDfopOfBwWJOrKLNeA1Nhu
CvU0b4BvTo3NHVlnkKs8ctVH2Snak2Izb6yKQI1sY7URD6Aupfzvy04H55KEd5t3CDYojUN2X+yG
9BGWmTEmvJlQ5dYE6QqhBuXkcDul5MfBz7Lyfkcf7P2+FoGmSlXHquxs7QeIhUs/IUIA8umiQ5iw
mCnmkG98am91iomZ4EHfy8F4ZvQwqhOnxmVLVVg9F7iJHSr933kUUC5NVjPmNmQNuKFYZlbD5JDc
/6umLKH9D87mMk91z4Px50etm55U4MZ7VxkljhealhQGxl2CdbJrca4R5HHsEPOzzrflYNuQtzXJ
CoU6Hk2SjGWj6+9DM4AVfNYBj8ETDl33BIA+4qgYXHbtQJRybCTNXJ9b02+TQIGso7Jk3O9JIESb
zkmgAVTcGiE3M09+OrapSjmnX7vHt36YnVtpUruIChsWT0KW1xxGisCWQwhHdiHs3Ty4gwjJQGGU
CIG5Qi7B+Du/+SjwgpkRSvF01b63v/6UZAnDlbQvLhCGvQ58VLjrrW3URDBXh42VemVo0pQRjiJc
iomnv98996dCdDlrMvvenfelV0V9NArojLkH3NvlkVjhKyL4qPXh52x33RG45Q8TIKcZ8N1WA3gE
mPbSkQOn760dTJtKPmrxyTnwL79xE3rKg6JEiCn/86u5Qk6fIPr5FUg0iuSzMcTGjDFZuTRA4RTF
VHSngA+ks0GK5Aj1Kc6407UV83X7lhxMWoAEH7PwmNsvHWOMUYIn/UKDhwuYqsrGYQgyFeX6etCU
aNfjQ/OrcTocSIWCFgByOckslRFwbsFQ0EoZFlVltHp83n59vyFIwJ/GeRZYrzdCvCC7ua8Zt/jT
lHekHIg70UaReh10yRdVJkFnCAmvuGVDID+Jsxs0hzLa8tawxf+BcrWDTqdq9XDmyDb3FyIcOmLU
7Z2m+VKZCFL4s7HhhqtwlzF1/jypRxqQs8pA5VMIn4T1XhQdzVf0gBs0d+W1MrUNmFVsN398K2p8
DEX3+O9THcWeaqKcoImkJNEy18dnsuXJJjTV+sxCxrx8h+vkfhW1ohf+UelD3TfjHpMbUj5KJzTz
Jz6Rto8nNiSQCLXnlK4Rj7S0j5MHW5Tc8t2TQTg2uH0WgqkKBaJPJ5gB+f/JyMCBiEvCQG84UWVu
hCPOIPX/BFmu1xrh54N9xi3ZX2onr1THkY1fblTHRno8K5mrUW8mvkRxQBtvIMOc6QXgkPPv17dW
E8BY7o/BQA4xfUPkS3tqtnqmkizvjDJ9PsgXBhPYknsP3YR7NQEdBVGaYCgxm48qPoAYtdQXSepV
BaZjMESbITo1Qqsa1kZYzdHq7HSYsC+O7JMIqxf+84ydX/FyICZUA5jW38IA/vdwS7xsSf0aVyty
8M1ZpSepFmWETzoc1nYqRFrML2+8gs0JJZ+BPd2vl2mFvlyiDWT3IZc3jX3JsDiH8t9voPUHyVey
M829NdvRs326JBdG4UIq7ZEIJ8tGYORzQVsE82UaDwCmrV2C5Hx3RlASt8ZVZBlMgaIItYNBCAvp
kTkP9vq9eXDeUOobLOALaZb/99yEqVOrx01uhUI+XBz85cC/69aLsjSo2BJeSTQai7L6IwrHzZoq
QEIruN5G3AA8lXp6pmjB919FiDLbkr2szPzHZzqp9V4etA2VN2zz1OvYUd8ITnEHTRkaVMYv7Aoy
co00vYZZLreZfGwfsBLBZhUCiPx11g8K0kiU7f/5A7UldPwzOdwe0M25SXbEdiFch9DbItALVp26
rn00NX5eWvY8vMU6Lcl1zTs+/RJKhFPAufW3L9z9pJXBvyZOHiub8mIPsRPdrwDNZ9ED0MQh0ze2
HtUN+cprtO3rJNqQ76duBLt0ZDFPpx0oi8xvUkeIWrZg7kcS0gzIJqG6LF1E3Et2Xr23sf8NLk9r
KdihDtkLKn9CCG17dtibMypO1NexGMiPRQUoM/xZxpysISVM57HaWeYfndqhgRha/8089/sryOWk
uNg4ZQgIjTkTa6/48MH+d0Rq02DRd0vHVVGF6ifO2EPUfTZ8ZZ154Ev6rZUe42ehP3ciue5iDVqV
LSvEdfcndWVcDCXTAXBpcd+DSI+ZkBSxOSU3dmMlc91qdEnvqeT0/yhzf9FHjlq6wAhU5nQmQogI
gI9f0GvH7axhBrZxQCktUY9tTpQkuH1tDI3mxHyP6xCg8WKmwFZ2YDh0MEM1LiPN3kd5OGJ2DXnU
0QP/CUPt3GBjae5HAk0vR5rwmRQDNvd6YfO4l6YS0Do5ylcQB49hkf10lg3nCE9OEQoJjYFAS2pb
TGkKqw/2kWkOL/OucoGq23vKAYSNfK0BpGHgw+OCMSHB80c0pXr0lQwViwjeVmNXx56n/oOB8G5V
ANWnW3d7R40kEcK+hEI5LfUtiVxlfPJDSqKffGjV8V9U5Oxw61UV5TGIx3Je/8J+4M2RoZXgYSvU
7fGll4eD1qqUMkxqiCvTAKEy+fJ66Faftta3Wxsc296ijqCz7bwQLewgJk9velm6yZISDASWqKYa
h1vqOUpcxSZwhlAvemKI7F7CfhKuvbiiYO4/oK2rWmS4QigtpJNAICnLbel/lVU4E17AFpOaCQaJ
b7IksxUUxMaG6EaFb+ysXApApFtxsPX+gTp8OzL5140Ky7g9vGaQQ31+ykSaH/8UJEW/hp2NTzc7
K71qXp6qbCW6A4uRykyKQryhXAekCZGJVZ/zrb+aYfXEHeoZFwiaHvJYxyjTyUq9rSVGHFXSQjO8
oFeJ5eRjPcd7gWl2OKVurfQdz7/91N7DA94hV/Zq4U1lv7bOmrKWagyoR5eGQkFc+MgBpZno2iwr
clVCHrSwBGtgPNthMbBx4kepnzpTM5HuoC64ULjGHb/k85kBrneHATvfwPsxsw75KPdQcKX42hzV
SE060GCjT+GxCIp53SgJfpOqSJL8f8QSMzOez1yia5sw+VdBR745E1417r7ZN7k7EQOc3Sng9exP
vJeUegO0j282IkuPBEVs4nPi2d/bLhRjSz21LdQg7RYKFO34euQ+f/ebPgoJAQNUVcEWXYx9I5xh
7Gu7tb7GVbNaAnFkCPoKVnj1iafK3B8GJVM3ex7ARYw70k2ZZ+jE/L7tZfWy9iV52wWza1/Y78Ao
e71+vatycNFKLRAryZ56TZ3roqTV7igjoBuiZUJ/Cn6fC8NnGNau6BZWIpYGDWTSkm8OE2wsNLi2
EiUtT/vXbUO+K3O6MKobv20yjU8xXLsDn7kdEqyn9YOB6XDd5d3cVXsKo8AUkWj0xqih83YAOmKH
liY/lZlN80m8oo0K1EwLXp1yiE4No41WLuiZWU0cBlTGv6gJUlB2Zn2vKoyqfbpkTl2oXd9owKkj
gEAiObc7Yl9jkrpucCrZuckpvZfUYg8SwUwXrJIIZXviH+E0KNlTGMLqXzTZ+Zb8/bhl75io+9SQ
hHHSGhKnUGoa/nnvji1UrlxnZkJ4lQR5tYBX4YzLGOIfEt7GIu4OxmtSQstVEqVnDW+2ZGZ82Nyg
7CUkfJG8FO3NI0YV5/0ETvpzAbb+MtfNwfee2fG2BhmF+leYlZ07FZKRWAU1+m8YMfo/kLQZgtjH
Nr7bmwVDaHmr4337nOijlVVvWVck9ITGegxziTEVXqdEOtqa7aERc67x4Hh/baMZdrT/ld0hNbbl
WVg6RNDObf2OC9cApn0VFuoVJ2bInm2KoazJrS9lPXIlIgoAJ39S88MoXgXJumGfQsIJ1n/yCGzY
HwtQV0YQDmy9eMlJjbzJH1xD0KBMuBP0GlkZ91KqiEoAdhCUlwKXQQfH5iGyDePmI/k+R5ZBvzhc
Dgve2/mvFyj6Cj7io4T8kzZyzd7ftaW4w+KFNoi5L+u6sA1NXYITQwuAei4FkWasuzJ18k0d5jLh
SMd3P51LJihYsyrv75Reaw+QS+MCrJffJ8uKM3RlVhz6qh2M2gip79MmPVAfOlPblqKr3N2T3Wp3
jdpgTjmb4mVXdvoJez2EJ2LNbCn+M5NnYD8uBLsyAeUOH7q/VM06pd85kxiPQt2E9+eZoP77S3jp
s39ehDaLBNmQ4/XL5zezzxOWxEFV+otMWK+McBiqxN7CGgRkHEZkZS5RXoXw0FSk5uP1Ch4GYx3B
ZFwSIGXqXUibxlhQMDJUURNUb+pgtOhyvHxJFzFsKzOpoKe4uwoV6gHmUkmXMZqEIKEelxJ6qSak
QRKN2lVd3vOVjykyh69VhvsfI3oacA2Iw85DNq99pP8sKFzeazYCB6Iyu3sZYeRbdx65lG71IKf/
J2HbzfXYnyNppQ4yjXM03xaAoVSN1iiiIkRfnIPrZmBzFF1nmljLVfRxYiKzASO1juyVnbhXwBgb
sq6f7gA1DX5vkDOTAoSTVuH81IQdvRxEYL7G8H6Vjr+A4Igod1w4ucaEMABjXneLGywATeEhY6ZT
d5k4QS0DVid/c8T4TWv5TDqWM1CCOdjTd/uRPnbW3PmvwQ0kOLmJat0/e/fi7C9a67SkIrgKpqNU
cW7E3rNhfSzvfrQN7lnf+QtBDnL2RhY93XmkuEu32MjoA99926HIsyeCUfZnXloKmY6HkKFb/pCg
FhEss5Tjq+/m3x6Rh45B3R9eyzqQ6dlHcLINtqJFAdg4vcSrFvozg4cH1HpsLjMPWLq8l1n00pJG
vA+IJgXRpu5Gp1pi4J1ZukJxWn+KErazmQoEDNqsbosPw7itDQVMjnZfrH4Z6gbzQjLLOAjhOqPZ
FVodpqt1fJIDqO3W4LqX2/EDV25MmPPbB1KQa/+86UubLoSXCbvJr2+M43NHTI8NItC2mGOl4tWA
7dq2O6BwbF3TmVIALBhJaAcO93VmMF48r8T6b12/FlKZ+F/COdgfMPnzCk5REjE8RLQhHJnu2Mat
bpEb3AmT/CbHs8L8RUV+9WpBTOhgjuxR2AXeFh9M+9aK2D0g/R8cuJxZb5GlaJLQLtImvGO6+tSJ
oz7SNnW9/jmw+7Ybn+WZyMFpRnboQLkPmqSktHvAlEINOodn119XThF6VD5Auor/ijgLosTAhNmi
zIKOgioSD4scnNIZl1q4qbcAkYpUpqPQog8bn2BMGc0g+PZ+yFzT8n7PFYmZj5RriDDaIgVJX3Xy
Cl9km8vNmmbiCkpJLojik5d8nYXHVpyri9J1IcegVLLVJcm9EIKCPgb0vH5hnZy2hIS44nNEEc1m
SB/0yvK43VAapyUn5ggIrCn6RytgwVQWUk793P+37XZNaDtt4FrwYjpzV4rz9REFLoPMb1FGUQ/N
YJy+uAMleHNxTQ5bnG/nqQ7ABCd9V3c2ZvbDy3z6neeIi9egnkuqzuaJJUR/h3Yk6WNUivCz485x
UlPOWcgftaFZ/qD1/pjg1m2RJF34MkPH+r+v1EMcAJYWIeeIWJrZBiMTjGR+sTET3497wRmAgDCg
gTzAYMN5Eqz7JdcA3/F8OWhfFYdIS1UtLexsb8fmKfld85MPZDJdHEMIe6CFI8tlXlJQek7d3S+/
15WLzfyNx0AO2omsZ+QAqctC1Lrj2Jonis7qOzWafGlpMLJJsSmj6GTqKXhPpQLhJTr2sQn0V+4W
R9Wc1h+Wa0M0lpqkPIbj95LtGlGocwKHfOsewTSCzq17llAEIs/gVFWeeh3/EMf5hJgjsQyZg3wl
GW78RqdAYGNiXvBg6ZSJLOV0GgajANU8NG7Kh6ixEmn6XT3/Zsnb9lRDMFgAblPWPcFgmWb+y8YG
JJIHeak49VOtM6SWly6rizR4alNDHU0vd1w3J4fGc89gjU4yl8M4vMUZYXvQwX/i6ak5ac6iGh35
uxgiB787bF/c5WXY0ENn3pxj+dbGD6wzTz4qXo9trHltjk/bfqy4nJItJyvNlS+7Lp/cPVEtMk91
UHra1sMo18Mr0QGV51qu6r8LLsbK7LNE5dLmT64oR1PRYcAJ3HP/vlY7ms+pXBcwwOyxlW1yAddA
bRoeTPkIOljquHx+Jxs3/RdWjBtB/PA6ufzjJZX8PbGiOrBaSRPJAxrGfbb5bLofFLlpXlDPMAzI
O4KJqy2Lonyy+2DOMNmeUjFYGlrR0nKtT92TTZtxwyPqL6kBNQT5n8S1euxqukKrDpjesz8C1aj3
ROc41TCvuc77liahOBUCAG47go1Na4oV/fddoHoFlrM6pr2hFNh2FgFd6JAFjDfOE7BJgQvR+84F
QQjdGIXhj7FXopHs9aIPwPpOVScdfHvEgs0EdMLmJ35f8gs/2q2RMoobBTzK38gWYKPzcGfH7SSP
i6kE39X0nmAGIT89oIeukHSInum4ZUzeUUjqkCZcZGDp55dGLzBn8Ky0Ze8iWZcow1r2H0ZKCD1g
qYdJHqI/fg5tWlMbjUbwZDVIpwKqgQvjevdk0BUll5JdcIShXU3pbwtrrojCvVO6pK/zPkbHK50o
S4aq4ZdiDLkJoRBu39Vd/2hxLmayPO3RNI1AYBs8voEwZvjTfU2hEeE5e+iCkQUib1ZRfzdyQu00
rkZDmuNSXyyGuFiN/crjAkD2sn2XrR1devOG2CcrebPSGcIz96m/F6PHfLehH9Bum/phkpZn5c8L
y+yKYqEDYHpmu6jW4fltilGakV6pDhLYN3zo4PbogjLfpzqtx6oxayZ/5IJ/ueU4J4WToWbh6B0m
n/ahqZcxcgQQzcF3ForlP5a1N1v/uoUzGX4hLaC6oReZlKaSOF4+JchEaYTk7H4w7IR4kjGT1XC7
0Tme0r5uzwhINYCQc3CH8egATRtnems+jxICTk8swSJZpZ+fOkhIJNiYddI+X9uiQJwCMkOA9A9I
sTVNbhf1KN2X7JJFJlFowQWpb5bk7yttwoTxGmFpEoiW6KcYCmhWskKlWqHWBvNnMuJV9Xt93p3I
lZ6d/QdC5BQyYNXHxijy40dBmVzcK1FCtrbqKM8vQ6YuR5ddsRiHGtnfYDYxpAMbgqdBpvveJl4B
Ek5MwehoSxvX5mhA1+Wi1qr69UIcFD7uvW6n1YsrbZDb7MZcf710zGpYyGxI59Qn6G2iviI2V2PO
UFtfTBz3jdjIFVVrmB7BrIgAZMn2ki68XqSeh/1uLBWF3s6M2grcuf/Jzuv0J2xX6HLUanVxXLEp
VtoBhJkRWMYEUJLq4bKEan70EOyZpgZt0uViuiBQI+0DbOpPLwpb6BpPgBFROWcEfQWmH0VMrFnJ
Kg9Fw3CMjL+bnSR/CwzglGMEBVCyYLMt0yKmV8rwWlx4azjfxbUss3JUSBjxlasGYjmDh8bjWNON
qinKUSlMuhCvnT1SSQEek0DDrzLkCtKIcxK1VC7B6UudwvsK5KC7LBhHOpYvDIsJ3/+LXKNHHKTk
eok+6br+BrM/Yt8wpEgQgkyzXD9oDZwurs4360GLlsTGI/2ipkPzHyI1jdHe5h1AWuR8sWwBogqq
BtGC8iJ/fl5EuOryIQgKg91aje5Rta/vHgUa2qprqe4aNVipuErrDmhOlnUN8LyfwmYmBX1aNSM9
vFRUsJpjT3HpH5Hjqq1PHFLnDuE6iUzjGIwlzAoM+XeeIKI5D41YP2y4UnFfHxtpxhaQt4ucD+Ok
ocATqoEyI2NBccrMr1pkyk843xWDI7dtXEeywh5tg7ttSPrSP5tCJoKslOCOTI6ABhY8xYRRIqMX
D9eHdWisUqylM1gL4lV8cBGQHv02TyXkSoA84qLXWJhoCgatyDTHsAEuera1RlGuhCNzbvNIeakz
kuBpwek0RFBw2WpS7WhuCuZkn6GEPtI+RmcbK39qlneWuT3Lb0+dLvFHRzK5FX/OQmhXG0dbAvl1
rUWzaUEZuy0r54qHgKnXy4MwQ4BxRImXwO25bBxYBg7/fk1gatxyVdbx4tbWr5BGGVaXF3CbehNy
unsh54dYRsLMfQfEaSKcFV835AbdeC24j/VyFpDsNYg5+xZ0IKt5p6173ykt9fWQsDeoUORddXil
7snzekGsldpFjaDbHZpqUNhbcTUOXfv7aWNJR1IyWtdzEXE+YlQKR1/Bo/wgJZYpE0S2SS3NatyO
CpzjD19dsKi2/OWNtoM09PliHHkhkQP2fb1sa4NLr8EY2SpMpO5yGCEmCOFmSebhIb9rY++lDW9Z
Nrzf6tH9JR2lzYo17XpaZfK0yL9QTWSGUwjsnNTdT+Vnuc2OWOeuIXlg8b0uVeCNYIfv9r8kfyzW
ZrvWI0LvUUhB2HVqkkJm97zTpat2MndA32wum3rLwTFnRzrGrh+EjNC+pzbMBirs+cG9tp1KYaZI
8cFd+qoUzv622NbOz4qL1Uw7747VG6M6wj+4g0jeysD2SVEYh2CCy7r0ETPGSgCzVpo3iLDsgBwp
DzVga3F1P5Y34iN+7EhBrXBTnccyV6kSB6ZzxsEErrVj6+iF+64VRiMEsxePXAUX8hfsqCfXHDQA
1f+Xe+sI1CViO8ReUob1mJrYGn/95/7Ldokkh6QdCBx4ACkT1KpJy1XMSBA1Jmjo/la8RE7KWg3p
k5QtGTR9y/UYc7uTZjtL/NAGkYlwvhTteczJQCpgCzFewxKFjGsUFDBd0bmbwKW4LNrC1gpaPKJI
Rx5acRsy9TMGY1ah9PKJiZ1jHHVGE3mshtP8QTqm97lFCnLdGmvjj15AHCu7QIla3cMfmc/LSzi2
KAvJF+906KvwZwsXWPUxUwOtizNZ66bg6eUigSm/6XH0IVbObdNPuI1G24uTNc6ZrO+Y6NVhtcNP
kQLkF/ZwL1IpjEIpDJFZLm8hq6GhF3a2LK8tS58dqmdXTXiFZGxcAqzSduzSfrjWtXzFz5t5vkQd
JbSKgT3CphqX5ojTf2pn/wmIURRgMS4Yt1TCQqc4N4VAosRUZlewhdm2LpwShlxAnPkk3AijKw/7
YUWUeyLjuyvPWr5MkAuLj9iev0y9zlf5rrXLOqjpEwuG40eHPNsfnk0LtZRsvfAP2PFgLEpoRoRC
zvAm3e5Q3YBa66RK7/wSbko5eVJecTUbfhqfJwIcI4LSZ7CT2jAPJ7mcHJiwoeOtjhDSxhdnw/WJ
LP3teDDdAytFZNNO3en5y31fHqgtxMylueZg0KDrepq0rbWi0sYhRaykuW1CC7Nsiy+Dn7rZRgRO
uPLI1QntBUq7oWLHEioh/WFUfxiPBEgDFfZO2WnU4ig2MBe0dCNx+vCXQ+3+y/NYjkp+EwsDv1aB
poORjK1EMxw+PYA2OVpBnOmxUPCS2aQvJyQlEQ21cOTd2G+XewPGY+YMUBuR4l8L1G+tm9f7hilP
53K52QlZj/eJTBS+XPeVO/xQZSSyNUGXz4UxT8tbKhdmF76UMgTICDzHEATSq+mfezeAmDvBaTuO
cA4a65IuXjjEfeXqeE+7IFasSixG/UQw6b+E+B16qsiMav73lLbiibSaX6md2rdxW43WY8pEsGf2
+A73hvXF6TDC7ZtMIN0mDtT528fgDqCRoeLP4YlZkAlfx9ui0gTOAIK0NkUlH+7whgR60kaq6EYv
HepuSY2u7iu3MzKEMgduO+oizSj1LkB9jwuF3oJkCWLPFrw0SKulXDDBDUx+/DHSB3PiaYOT1vnv
C3ipwdzNYWc8SsZVvyjSzYF/bwDKiZeObMEj54kzG4MkvGaXl1lYv6xaEUMuglupfGG2V8HLwpqx
ej7w8+xBVptagWe7dpwXi5L97IK3neNbX0hNjSK+gDQuzCWl2IgL4KfpbReJpjTL2Uf9lsbzbtoA
MoKohDH1zbVu9cW/gRY6aCU0gTUmw9wjJe+eg0xlAEyee35/kebs2QZehw2vtJtIndhGxt7QfsOq
claER0HxPB+s/vnFI4Mwe8KjbCBupYX4Genphyt2JKEQtjzsFoj5GbA4yTzabTC92G14qigi6gs4
uuKnYizk8ly0bQM5m7T2mlKlGC55ose3b8jAZS+rGagW+qoY82NkCIiFArmYWqqsJdDQyM1Y7vjL
zQ9P8ihLV3Nj+u1Ked63PyFo6ZYEDVW6x/BC4mqrBgau+g7q74PVlRvx5AuFIl+8zeQRibthMkxA
zv9o3qnXFMecCgAYQoqyMSEcZZHQW9vgoq7FawA2OFWNVKd5oCvMEcwEgCdFTAOQiTCNeY0cIbBa
izGu4MNjYnojOLiUN7NurLWBqHq3alzgNPbQflO9NBSE29p6sbL6bQq94z+RhROviLdKPH+J4KKL
yejXzmfsFyS9YDo2Rz9f7PE0eCgi3h8kPQOm0sfxeNMIgIxWRfux85l4G4e7BsswHH/HApIQUemN
0FGnrY1g5gGXle7o2hp+qBUP4JeLs4iOfcu5qjiTvQ3PjTOhhEatYR+E3aB0hiVNhnCnI87VpC/y
03O0FgSH37JQnCgpUOkNOH78PPH9OfPi/9/162fyF3ktgZZUDPVIlJ0S5tv+roQS1vsYPjGNUF2C
JlH9CN4kgDVmUPxKbmZPcYGFCCAHKSTfYeM6yXuaJAaquhMDSWf0opSkwGGSTc3P0+LRJKzurs18
M0JQQjvANhVFlM5cQM7qNLFDuIP5epbj/3/e5iR4OrjHqE9mg0/M9fuF2hpKgBZQs5CBi9zkhjRB
MmyJtdOOkkomYay3dTvIM+cP8VcHE1QSl2VAk4MbLBsAsn4u1sZ50XDwjwOqIaOTNWgp18GFW3xU
FBgXKHeeU5uRCJaB3s8Z8ZriCJ0iyk1INBt/sg3p1xBUaDyN+IDUlL8BV+IV0g9+6im4UzupTxr8
Jv1IVGEt8c5D+uUJOeXf3uQJKEbLg0QTc0qcGP37yxzmv7S40ofUdAWR/1duL9LVhA7+vW3XGTfu
3FhyYrwo1NW0lhNGo6uA0OIwzpCkPKVS1BC6bePQKja74zos7cvjOYrJdpJpG2PZOX0cWcRUbf2+
xn7gv+BxqhPV8vE72A2oTVVRTk/v2Xz2pXTINpR9McxK9skMO6n1qo/qfDWz8Sw54aWsGGGsBtLF
PKjOShCPzUWbugg5lbE0gFknNDoGgWAxoAQOP45L/bfunaz2NgN70jC5BIIvp9+hFNzAIyn7kkJC
D+Gtaw5h7TtKlS+uztkWaDlbMYPArgStxA9gbtDVRGjaSyCHX0ucN6M1ugYLdjdW608e/Bi9sDGb
6It89BO48L/lSc+f9E9u88iFWPUyr/sf/xbnZw94BXYot4B2dWXjMHJ4QDpzYNNJrU8n18MBFeW5
WqeKdRgC8iNGBIlnfG9/inWW1XzUq7RXuoFluKTS0DEU6e9nCprY/byQpehF3AM2U7pkJnMD2uTv
2GDDj+JlJu8Cw5Zb+Bslx8zw4vvr6mpPWfG43hUKWcLTXRWFRn23z+iCJG3E4k6xo+eYiPr3CL+Z
vx/fycoAwrmdYkcQ/AoMPE2x8H24AZ1qnEEbREJI78odpv6qshKHbFZ6a5OUKjSeURfo7TXknPGn
KR5jNFVsNM/U7eTH9NzTsTx6VUJFiRqffVRq9xD8+bw6FrpJoVWngfjhUhc12skoDPLYPVCoK4HI
PVwt3DLLVjIsEVLqciMT1BHbQHc2bWEH3MbouNqKynsCFQKqYAB8cd5/DZRHeUAcALIBnDOkKUAZ
1vPXp7C5Om4yqy80RF6hiuXr7hSHdDBcMqL/kwdx4ZVomcdGTZ2hwo0MvQd/14gftvO1AgtFeNT4
HsW4fR+zN7kzhnMs4KWPLYiRr4YoEjfZY4jn0v3TR44PCaqJlq8akduTezF617ikUy2XIHXTth9+
thHtsw27sZGpfDgMNtliKvumkcuyBD+jxk6etgZqhmG1hrVFBcQ0ZaLGePwfn9Nw7Zz4VOuGXD6F
rhxz4IsDIfkeWGkuijFTSeU9YpS6rL510REbpUlcYXjr+mzxY+sqyveuJby1i/6KpSb0q3QaKaj6
OR6h7ZJ4LqUxKSzcn0LcxG1G4POURdkCG1GgNrsosb6tADGktFMm51rUVMeMJa3JYiBwbEoGHX99
yi7Zz8Pd676vaLVSoLMX1QXy2meieXl3HmoEQge5fckj5avyQ3iA+P3Hw5Gpgf1Wjmv5iu0Fn9Po
rwIfJ9KtldLJHaykc0PmNV8gsKes9kxVfa38vAVXB5xCboFTIySDFwS23BtrmTSxMJZTFZQ1TWdZ
R5ddHhiWryyDnQhw2ZYmaWf4GwkkqtlJP2zfu5x3FQLov+1GPF+8WhtV59O+eUbdAsIGwgjguq4O
A4OF8ilfYy3z4hMOnxIFKxSR3yfxnxUQG5quvp/m7Vd52+ocxEJyglg3gwuGsC8Qu25tm3BTjO9X
18FLLoJxurF45LBGwgtJXPXfEBL8lKzyvs6f7ac8hHaUcz5WLdEwFeOW6yXUpy7VeyWrDkhpqHPg
481UZhk398RSeejMWo0VG89FxEUmv7hqJx1eXqF3XQMNKhlscESMM6Sjwv53W3hglastTFyBKBYG
Gx4NTj+UH9WCLdHxGqftzir8ex+kQe+LVg0CFIQneks6r2pGa0ffn2bJ9PrQWIDIhbgijkvy9ZPN
H6XAMdbNl686ctmkSww4rHxkDkHyK4gCbA0YJKRQWJPOFzInG/0WkD5Qn85Uj7fnkfwQ45LXfjq/
Ev2Pvwpu6WtR3r6hpKcircp1av+s4zfwIXRenvOBlbbJNrC2aBwwAgw3IiKRlBXWAANKyY6b93tj
TmxwcyA4ExZ93J5/XQbSlVD75kt/mfwWXgUD4mgJfTIOtxgZsQw7W/jRHh2Zncmf+D8PQqjv52/n
8tTehEHXPHy5GuDzlDiP8WEtLpUOMoMRxRKxHhLEcnKAEpiAWvz7RbmPJoHdw8obm/ORf3k5RgiF
K8DOt9A04yhXMefsI58Gg9mcGNP+C79VYRPyNGWj3FNqQYS4gjcaS7kpAtVfQb6E819b0A3chqP7
2KidXORacbEEsC6Woiy52Y/4cqeFEy0znN5ATp517urjzk5RlLbeHVFq2oLud8NrylMcOSkCwIK6
RDtvh/MeuhO/hwdTqzIDKqousJiG1uudsuXnimn5Vulg9/I0A6m8Mt0jIQV4Js85Rrgq5MlecdqE
Tq9jpw/fXYgmNlv9/JY9dGtvt8o+6RAL/5WmXLS6NPQiXRrCu7ij776+q0oKxN6tXFikSu9O+VV3
0osaigfWG2XzdQ5wFZOMbYPEo5iuiY0Zgr2XNUDYmvdIYsX6h4sOCmJGTh3edQitkLETZEK5GR2A
Ug356SJePIoA8VOYBi592/03kSFtnU2ufw7a68tnLRTcPf9ZngiSTEI0rnX2oK39wwbza0oibCtj
eM/VG5TVgNrNWsOJqJs/Lieo8Ic4EoLS+9L1eHfck4TM8ZUWWVkalWCD1X04vFagFEOzlQ2seb81
rNqgffA645Xi5HHqnh03hlgbcryMncPr+ft6LUT+TagwJXHSIqH9SVQ68UnfOnHRCmn2iC1agyLE
OHDHzWWyNJa7z9lb3yQaMpexyysbFg38Hxk5Hha83+tJfN3zdc2hRabb46JzCCbxS/PR/aon2gNM
OAk+UZxhJ2AOl7kbQ9s+vVp2PNRYdu8oYaJtmxkA0FdSAtssfNdFtVXeiKv8vJU0G3zEXwNq7kf7
isWg14n67r0KSsHhTuYU2WvcYnUbdcbNubu94oJ9ZUi2uXA8mrfsnF3tXW5zfNTvs9Klgr3FB7Q6
J0s2IEgLDqhBphmH/tdwvWeWiPO1iwXPntcQIazaTOa1VihW6mynWbxNRBJ0Eq4S03Ce8WN3/GLV
YH3/F7Fee74e2x1ybanKsV4T8SW9srIx1/hKU33X6BdemLqFI0fIov8havKx3Bf5Cl5KDVYOJ4au
vL0GuhgqhxhMI7qvh8y2UlaYpoZa08TcjcZLECBtDb3PhFp0qbv9c6rSCuOYjo+fcESM7lkjzft6
yzDE9ISWE2rAvkKOyQms9iJzhCU7vEg6eMI8r2GmKodxc4Xgk2o9ytakSbR+DONal3o7WJU5kQm1
6p1LY9Y9uO1jT8L1G+VrIeIUv+hzd3w633LY/nWVuzzgLFGAII7xvXkxAw4vP3UvWUDyU1mocyE/
f8EV0IeLfW4EPtB/zf+zfYmXhvue4LXwi3GgDoBry54ILlAIQWUC1FHzBtzHW7YUX5NpJgFt3kst
w6pyA6FsNm8b2X2uv4W5l3I8fivSPgVrvW4uOfanaQ84rOOfARBTgYeH8d7BXHn5M/JM9SEjDmQt
iLp+Srmt3cMN4G4bqAwzECRl8Y49HcA5oSB6rS3ewqHEdwo6Ro+nNWV6AoK6fFn7xoI5eBWQ59HD
52u639oPQr/1x8o65f78W4w2Qx0aBqr8dHnRm6KrQgiZToQIPoRqUX2kRtQy8TLZGX8eXI0emJdV
LW4TaobIl2Y5Io0RBJcwtjGB69D29NKvRPiczZvBhjRVpgGXDG2LrWjH1oCtfn3dYYYpCeIDWPOy
sqjP83wA5rKMwGMh1Yor8nLCUWnnPoHR+7Y72D+EiGfdRV3GNrWVTvaBjNJFgHqX+oPgiCuD7yrz
Zo31GbNliVJnL9HE6VqxujzQQRwrJevtwFF9jrApvf+rt6hw4JLULD14OSDB8fnQJpQZOuy/Svku
YFB5rPvV78+iTHDGPfnBDqGy+VssxXxX/Ka5ZLmDqCfLcomCpIqpXy5P8ihFBxLEky9joyQy1xka
Xu2UPja1AuffU02Q4+WDyz+bv91i2LuWLk2annFHFCqeFX+n/q1D3rPLKR2Xe9F2G3qr8oxJwynP
c3lP7SR+33Da/fJ3/xeRBdZUxeu0kT8yIaN1SUuT5inZQTD21r5xKRq/P+8PZYRvLC+Id29rbNfN
rPjYBQF5CsgCkaBVKXZj1TbELjcs+UyQ91owTFOB/DJfypXK+WCyQJWLTdlK5urXQmc6CipbrUTz
oTXH6SvdHjnsBdPLJBs+54cKPL58J1KuMrLBjn3iWNBz6mSBtjNGaRbWkvGx5C2bH2230fYkCgH2
ZFZ0ZAQ8A+rcqN3MEomiocFpXIs+82gOVOnlilpVlTRXTXrNeLkvvZi3nIEVezM7ZUiczaHpueZx
879HEpON5SfqV/8ezxNWV9x2VFl+dvo+GAL+TbwS9Zm+aA4n+UWsnXH7tsHJdpMZf7n4TneFs9Bi
xGGlRS5xq0g8fvVEI0L80psQ5lB2Lhf5DkCn52AQu3TI83ziZ3Fs9+1aCmfv+6RzcSCz962BNl+d
pk6rKgyVv02NeStfSvIxT+pfxeWx07sVQQLTTVvFaf1//zSz5TqDqoZIWX+bRj0cYftM+AY8rgba
3A1zW3NpzBCGXxcqlNzA9YTtGJcZ2mEU/6vKxMF0npV2X90YTYsYsFnpLt+sqXpUVPHptMh6KT77
/lBXcOn3Muhn9OJzN1xv9hkPmVXBoMlsIAYisPQkqk26brOd8e0vLrKHnBu9VSYWSArs09KxVv22
kYkVYG36H/AD9kcs/UT1zUnp9yMD6KML+L6rY7pBIu/0f5wp9w61EqWc2IAUuIpfzcuTk65w1b6y
+tzlNUoTU9xp/oMZHNN4AOpFKr17vGsvx+LIrmk5ldlV0VQWwuIKclj7pl5qydNIDUoOMSmmytEf
0E2XoeIXXH344j/GtZ4tb8S3D1NqHN+40KiJDx0KA5Nv3sWAUXkdooqgLBD44h4a8xpzPxU9AFT0
hUBYXKjm8ITiPpdOOcHQeUbjRpyGT3z5Xtxtqv+Oz2iv22DgpGD0KzVtjWfXyVgdKjLkRdYDCVLy
ULy0SSgy7TB3zpPbmZ1V/SapjZhCg7lfDdLjpUpOGbTtCmS9j/YQLDWTYjllkpJaF6QZIU1bsPfy
jUODFr0k+omnF7QFMBYg/c2i5cXtvhYRMnrELvQSM8wBBR/lIhQIFJTAH/eaqnODiNgLr9G5P1QN
TwKKhzJHlpWXXC0vpv2USQy4zWiBocAhgn044FehRXUaD6Gra9QXAGhgnUxMHpIRqpNCHG8RBGii
dQLwE70fm+9KSleBjyCH2oiFrlIDakA7omWx46T/y7wSfmaIGmTdFjA5s0c4rprQ2gked+mEnZO2
0rcKBvIPIKHX2EC4eWMUZCVC7bHpM84sKW1S0oo2ABvKCiXnd/7tbIDvygOJokLq6r9yz8o+AD2N
rjCVYUW7YF3OktswRcbF4dAWttF8Dt9oW6CkXVNmz05DoQzyHMvceLC6wfEDB3WirOqyAIwoj9Vw
M3WU3iYZhpMnQm2bP0F+96a6Lti4pOlxccs3p5kHc1ybAhsdOCVvunWHQLzG7M3c4x6m1/KU/pz0
Hk1Wo4Efrb3GQ7gt0mo85Y4OJvU82/3/cJGXI1mTL9YGIluzLIIg+NK0JXodqZND1NaHp/AiKGb5
uhtA8B75tIqE0L/mjvTlXPubODqJZqshr9KHnG3ty2ZstrCUCGNdA1yVyeleArGNwi3hOU7P7J7d
BmoZhiKL6ApRvc5WXdLGXSBEjIUtEZn027/FMPH1E7+7BDPSDXHQh9VAcx3PHnIiv972jXyCHnSA
7ZTBrJHSuZqqpMGSVU6bmg9lZr/PomxaGtEkF9TNjBc7fzk/VpSQfJ3gQmc8CCoF6beiTXSdSjE6
16MSw0gMqeniSTGyJIg94tDsGEjllqA6ho3LeRSOHSBPKKsVSqqM8r3r69sSYHH8x79ZUmBViDBi
kPS664YRKuJfwAVpd8eQgAn/asvRAgmQnlPOBpy2HpYM7IdcKW8LO1z+usvIgkH6kVL3+8QzPoHv
geUfqjwbEgMoJFN3T8QDfjz2GjwwPhepqKGmp5nY80l5wgJW/RNUSDr3jIMQbBb9i4okuoSeBD5A
COespoDynNMM7Ll0tjmkOtj1Gf0ySbBnTJgBzhzTzGYQpad5JP7fluLVyGRm7YsFYKr7OJ5NcwrS
kHnK5P7xETuQ0p9k4cUsC6LUBcrCPdFHUzubh+fLlXJ3U8eIDI67QWvkTg6aHyPf807DOuJ+am1j
3DXWPskA0TRW+Ia6UEqQi0eHE9OncAxtUY9pLKyTZ2fZDYaZZ4zB9ju8ZkmzsJdgpujOmoo2lJKw
mm8OvSLpk5stXtMcjay6Hw57/9rEVmwjFXmV/eJLpECklfvYdLfzpOaiAreH83CsjNVAZVxnnOCY
u4E83Gv0rc2hygHWP+vckLF5VP9kaubpUw3awZL1Pvdj2fhjpqSBVhO/hSYKzyaUZugxz6O1+Oqz
FUDMaNX9j1yPsohAicgWHskixfoMP/eoBiHCP1ztTg5LBN5YofX6NEsgd1yBMOR1yLYLfMZUOPBn
GvW1DQi28tbSRqoxma6Ou9GKQ1jJhG31moyR43aiPLhxkf6PVacFVI06E9TZeGt5Lrgf38WGahI2
99ZLpbBEa2z10fmJTTvLKO/3ZI9RvsXV/gC28sRgQQMPyqHm+ViqWC220oI/HFguR1AClsagpkyK
kPz4GE4xzEPDk4MMism6CwTKH0CkoN0BNkltcyiAjeLcqsv1XCk7a1uj0Wa3kWA9sudUvDqSnrRV
r091WcmvfVqQlC54jrbPOwXpjeMxmrbV9kdbn2TErGaLy7CHqVci3kRiaSTT+tSXLvBJiRAgup7x
/rq/m5+m0uVTjAPZgnPD/eLY6nWJcCxyCTKoAkAv0p6H1K5pFAGSu5eIpiGCiNA8n4h6EXv19zGS
qoPPYBNgb/XZZSg+cgCC9uxKdbi6C5p4GiHe6/SpnJsUY6rjSIvQE+4eO6sxTew59fUBRzHxAeL8
+EW56HWiOW117LsGRlvnmIfoZVCj60/0izogZt2P31I5JxrRAdNCFAs8i9kTsoUp2fbl5LnwXXyQ
fftuhVBhvOMULlE1xmyr8OBfaD1CIvaqf4a5FB1gWrWAhzYVCy9VGihwcAf8XXSQER34oVQff2iN
VBFuaEaotu+7yvmsz7YiY1amR3UA5ejgWMEBLwuUsdxYIixmu6/ShpNARigqD06fbjokXqOYAhgj
0UlWWFa2u4/4VEM6FS3OZ6q7GvhAU2XKLLF/xare4/eT8cEmOekSZUch7NLc83BnNYSJmqOkQt2B
+lW/+CdoXZHWfvIaRBymLnhXeja+E7VnqPWzphyTnKGud90exASE4JJgn8g5giiaNFjelBkw+zHn
AskHkH1df+9loVBnu1MrsE8gpwXXa864vYohABHoGF7bqmcPyVRBwppMLe3g50y3HsX4/vkw2a+5
XTYRCpogZzK41SQI6HrExPdA5TB0+Hu44Y4U7MJ+m8whJa/VFRIJNUfzpr0rH8NKSeRFzy7rhasu
WnjB/8E4h7b6gNOClciYrYqvZH6Fw4IQocCKhnMxkxas9S1f3eQrAf0Vrq61RYqfeAuzM4obaRD5
F255FszrFoQU6anWzNdz6eB/fPI7+0JtmVgP76ljdH8nSzKvRMt9JVpEYpD72i8SZIe+KDZJqu5V
FsthCMPN/eygtUKwvfyFU1ZISqfs8hI4lDIBVjjYw/KDYE501AGc+pVcXeuOcODv26HRU5dpOfwA
zCKfiFSlfCQGHWq/opQKYXjU1MbZIWl0KzJ32esG8dVF5YG9TVmYf0PoHnqiAYhvUSHx3MvRFNWx
t/l3ItgHEzvoNK9ohAbkTjv1KBpxyz0kxphhYF7tKEPqGcsCXkcW11iyyCokvnsHbL4QuYdjCE4B
wAdZn2wja3r91XJTc7S3HkGajFxuOh6BaXHzb/L2VcpCpdXv054nDYx44h1bz3wN37UxszDZgLOd
c6wsBQdOLk+syFRaoV6wZJeXn5evIFftwALFGulzv16RdfIZ3zdXiY4p4whP0N0a0TlhadzzKpSE
6brvvC6/M955CRwjGZlYavgdj4lqBb0qoP0jaNYPrpH+jrzAHqDVapKYNhzW/3ujxaTDcEOuCfyL
Kj08uCfNdkVwS8gPT5IpHx+hJIx9+4VkWCgqE6rhRUhxWRrn3D7T974+0CfsZcxPapR7gJOMznbu
sD4GTKGJvdcw2QsYKQLALq4AlYOB8R/63OLyKzY07hYWxgwPxfUs8jZZoDEp4yAmekYXRV2NeNrC
Y9Mw9ogxGvBbRLtAVTJBcQJ+kpm0LgZGPLy363h7coQdx5AzxtEuMeDcFvsfMQvyOhZuO6DIvDxc
YbvIyccJxklsb91TFvADNWNoMF5nWJuZeaLOhcoo+ajBMJOq9JJZSWhSOfLYaVt88kX31unSLGBo
3xOSONui8cDAnr2IGCG1/LhSGsiW5CCHqikseIpwkPHER1/WH/bNrp3OHyNlXT0cgALJgRpOfEba
nEoGFsL2zppwrGrg4U409WGZ7PqrFvVkYCx7BTuqVuqzhgp2cideGC1/W27Z14HVhf10BjesoQAn
kmcdNF3iDm+K7T+8BEe5dhkrG63T4oLl5yOQFY1MKL8UA6dd5AsQuyPLUKYRudaY6c1NkDh5bQSN
JZUlmxizz1OtgjoWMxl+pjd4KVZG90SPWYLyNzoSnlTucGifMbRsFzqQs6TrLU36DqJANdZCQ+r3
A0BGF3vmhUnWW0vJgWo6Gb9Xvkx1kwqo5ePTnCNs69zHK8R/GwwQVnGrlApFeyetGqMlI8byWGlt
FgjqbKaGP9fe5AUYSlY3tSeW8HULcmC7lxAds+paD7KgvOrbjre/aSzd02ca04n7Jcpna1ungMLP
LnOvheoxao5SrHVizM1lDC96B0pKKGgCwoRpT+qa3DNurGwRw4+/9DQGvdmEZnbqjLl3Cz288eZB
7fMSCaFCrpHYfQR2OJOgr4pywrbMbgtZ217OpWw27yRj3wns3cCFUqJsFT3sZvMPKwG+i1x1aaDQ
Vyg0GQjQMDAkFUr6CaJWA+2NBLvC4n70xos/mHiYporlzOKAH59eN6/M8JsedrRzNGjHNAbVXpuv
rSF0/NKbBc4RUgM7WGIAvcoQQZd6N997M7B8s+SfVa6MXXzIPDebCG268+X338xFrT/Z0EEGyH+4
sFNz66MXzouzldClDrh586siqPnk9v9f0d29rXn2SXCXgO0fTdIhv9nR7jtkO3K8b/J6V5vP4rul
bVauGe8kdu4+FnoLvXkl0Tj/LhHmCogsDUtVGYH+sw/hollTw8pE+BbX+4x30LpSBx5yKPUoqBQF
9AsZ5M3FXoZPZfaQF7xOVJNMRF0ahY2eCQJdgfeZEs1XhVS/QwhzDPMKYutzad2TKQHrPoZjyfb1
MZyVSkedi1VPZDRc49riLWIF93A274zdTsX1yxFOR6kLDOsU2t7HC3EG3ZmkrqgolgW+5bX/sOLa
ZkQ1il2d1oFYNeRNMnPEWV4jSVPt2Y5E1ji29HPgo5H9nXdEdxBYi9+um7PO/mLXCjH295q3KeuR
2FZSbDlMwecYJuRp4N7sCV9qgxjTP1tIXoBc7dVKojizNSaHPlwI4nZn7Z6SQfyW0zg3QMiUSyBz
aVhdi11YQoS2UcXcrpk6cZSj0xYp7ZswkHtZkBy/tibxA6SPd5u8rS+kVjSEnnc9tiPHFBubnqIu
6JfB7/mOVDpEiv7UHQEYrZg4iHRH10RDd8nzNKvtpj4ERS6jDAtLyvLlUJYurwO1yvO+jwL0uaX2
/ZdSGHq1ZmKTNr5l9CIaMrg+YjHvuyFmZrzK0NpOAtbJLLSbakZdqYYo27Yjrbuyn8XcRj5sohzf
7vxG3IL/Jvofe/WnR7PXzcNLoYVCUCFWJqMXWU5RtZkrY64d4/r5UvN6cbRdwDJMz8PlCFx2DkBT
8mH6acjIRfYzM7mB/XL03hYGur4YkN9C2WMOCCh0kMprJ4i2P7GUt5zTUa9tqJtKQBNWcOYNTYNi
snvgMi6VP2Y1aGeTnWLWvKKOju+dey+U5R746k8wjwuPQydkzVMlm2TTl+RzwumQJP9QF3YXgye0
nA2uePyItdB71uYTmgLUOQC/Anh2WFnqlldYkCQPIoNd548FLJkS0+IdYRChd2Sl+kqeauWYU/B5
aFPyIFY7IMZMMa47uSLsxgjMvOWrJiR9i1xwMkYGw+rKD2r3lE4pGSisfU0fDm7IH6RADDSlN+Nv
O+ND76ZKMj2Slyvr5RIBh8he6xxdqbYwRUsznC/LUFsYpTOSdjrAUlW/P3wz5Yp3D7K776jgU3zX
DYoZiFhzWTKvieCNvrj2V1467LOfitjvonzrggWQWN2B5VWhyjicY8/X367ZFk/fyR6i3Ikbk5r8
br4BOqhYxa3JF0x0wEXgkC7ARA3+SQgycaZSZCiVarlxJSSy45LDCh9ptWqa9Jl4RTTwE99ITR2o
YlOxioPY9b7FL4vQlUIGFY24dOVl4gdZ/WvuRnLgei/qU7HDsf+c5WUNbJ1QCuooU9DA2obdbYAw
S6OiS8T7jKQg/9DA+OFoT/sz5xi56VL762mK8g+sQPwq5kfh+yxkSU/NIC64SZwLHhQQChi+J3OW
eK/rKGd2sN+MzKeITGLjwNwa9I+ywzPWik8PM0xVDLzWfosgwRULKMzTNDKzXLe5ZA+n6oOt5hpr
0tsvGqPJBnk8I7K+eBPkm3OWJlJv9OPJelNMGX+hoBO3XBea4OAiNukPZ1r5YCF2OzyMiX4xWxDX
RCPB4/O+UgErJ/QrpGDkzcL/c/Uc3H+3+QAUwypbwn+DOiOr1aG011l/6mDPfO4iPJCYBY7qPpUa
WB/Xrm/lmrz5EcdaLFxPtdAGzSm7z+xaabhQnd5TpJ7q7TgXKozJBBbdruL+zHFBaah7nsqF9GoZ
WDMhS5bqDJzJHkRd+WGnLQ3jGI349TfB4AheL6cGNb0A1vAZe02WE55HXJwdCOSmXIF2mqMeb6H4
KsdumLbbt60RcoUmQNGn0wu0nagO4+8G/gl2eo3E5N0unKA908DkxOWeXfXDsu8ra3t5bOsXAO/e
RI8O7KaRSNyCuKHc7sLQdtrzShseFL9hw6Noxcu+FZxmCRDxTog0jGTwWXo0+3g0L8tG5P5bqFOT
n4UcMjLzrW2qoVBq8LrEgsfofTEyHeo17by9D+1fLUb5M5vmb+DlexuiuJGMOdBNmGUOZ0bT7Gfy
EQITc35ZxRqhIqrZCilnCJgp4V1E7/yuu8B+GjMg9bJwfpxgX1sJW3QUptenuDTAXamdN7Hehnyh
M2mLI5lPsXg973oHteiQz/9xXQKaWMHZ1DEnsQrRXoM0V4LHmB4DiAmp4idaqm8ArDGJOwimTi79
3OMw5eYW/l8HYGC2vtPqnvhPoHcBv8xuSFzhwHCUmoYJk2KE8GHRTV327zo0EnsqA/catvrSHM7C
EioLr9h7wPNYg69D8YDG1d7dckbtafO86gD13VKCKmz0jpJHnq7IXXIsCDZI+oAFNhLJXDTaw/H7
sy2SH42u7o8N+PqAcMahxXYfOfkcnweLz+CXaZ+cxcKfalPJNBt56YRjdAaFuognlXrjsslEa3f0
azoZ/jk6COuZK7BD9IFGPQKPYKj37bHHnHPXZQpnzxlVckeu3RiPjNBzMvsDZYrVNh5FRZbQajnN
Zb63N4pu+n6mv8Qc+hFQGlh3ywTV2+sBUW0jwjoSmvrdnDt++Y+eY9WwOoJYoIneHrIRKHmZbjWN
hWtIQrqwigTi+UBEfU60cZRTxzAbDCZOjnowVrQySRw2KQuimGHxd8P8ruc6lTK6rq1vOFbrNtKi
WHruoge2TE5k+BLT/5uQZsu9NcOJnLHcovuEDkgqZ7tYvLdtbL9EznnzwqE1207NO3L4SE+IlBx2
3c8xOWWae/hYDrkVK1faIOgnuXzY/evhEXRHUlrrvgw0i8gTvwFDyHpct3xzGyt3Oadk8OyDKBYE
M6EtfdWxDDSiITHkRxg717Xgov0f+ZzLnax3AxGQWFQDasN8YxdcDC94UDRDAhTdztuvWPGObKjc
EkRmcwUeTHUy12aicLC6rGRtpR6eJf9H7C8vPn5N/OacKBLGmOLXIVwQYYIjuTevM31GasfcwkdT
KhgLWn4SFBu8vpegFZGInocB0OgsC3sXNFVS4dap7UPhuNTdZyhdHUXEud2IbuMZfi/LPKyccybF
dw2LDwdqHRSyDZly9pwDavaV5Ku4TOf5/+Qa1HmKBhpFSEPRGAr3vO5z8l1O7TponDs9XWv8xWtI
a1qg7VYyWy8L44r875O0aa9PvrM79JY4oZD0bjri296fysJbbI1SnLoZHaoR0dF98YHSprBefoqx
E4Z+ebXMvrXKWckergstuGVzyijXe6h8q2mPlpZ1hkcgxxRvGlRZVSFgJ7Aqax7qOpwEqH+8r4Ja
7n/VeHyJGqPyARHqHhGO9k/O+RLfIHnMywYHt2Y5nQ+uD96LGg5P2w/tcnwSDqLw9UkeMSFxbM6V
JTJgHeBmO3W8fYcz8bQ+U+LS/uCwNJupFoDVoCYxRBM75f8ZeEgdD77jHtxBv01oE1ijOWilE6Ut
oF2TE1tsS+6HrYL9tvz7GBwokDAJ88pGoZE6Z6qxhokkk1k9bDLardGV0KwpMTJOsEvbXwd03pxn
a5UD8wvYlYEnGptBqQUtwCm/iJAAfqP0pc7Q04i/G5L5dw8WD1he0rhZzesMbKR+0uuK3JUp5kuR
TmwaEjlA1ZZB5DY7+BXnkxJ4rSJP8/vaYMSgyfdqJfpqrM//d5lH8k9tKMl0bjapAMjzw02X4QE1
LWYZItJXc1mmLnT8EkdJ053Vh9MEJ5K2erCadCzbQ8bGbXt8/tIUty3hX6d9RH+EqRJ0JYP8uTys
DXwNNwT3P78ijYaFEt6KSpUFoPVsh1UUItzivhcjjjp98EHtfRAM3awfAFgA8L5g7zAz1W6eiqQg
zlXeNufA88REXGsPX4rvQwpxO19dqsUuxEgNxVFqqS0KBba/hPgQe+AxNf5ghConLPQOoHO1rkf2
sslS1n5Wb/2spB5b1XCkbipLvjWxgdhtSRU6JQUqRThbXdxeF0GVkHLCoGqwNcEfSEOnBPivaJ/L
a/GT+TT9picnOLn5xBOwxbUEv37D33JnOS82I5LijCAtjbMQAlnZepJnh63SOobhHBAkXvjAdzg8
qy4EMtXKi/G5gEzYmgpHC1t5VDbhH7Z1RhmN3YSDWh2EotEhgF7d0G4uEftFZNrSQqfvHhmmvHvM
F/dCD+INwx4ZOwegZDDtsYf5Ih/FE/aBl+BrtzRmJD4ZJ6V8rE2kEIIjJFLh6lJllenLWjZ+CKN1
YAZ3cPlOQY12yAH8sIf9IIezEW+AW8gwq5WHwJAeUz0UiFkfDItuOSofXS3NEIA7jm0PZZm4zlPM
HkyAqgTgDocbhh8w8LJlqYgrPGIW+EmSYi05sMSgi2XBKiEu/aCT86y7uGZeeGkrKFfOchcEx+d7
/O/6r8N+Zsc9/Drpmutk07EEHwjMdeuVziM87qqJCus1Gq/x4dQAYHRItbnaM7nNNk86elzKge2P
RpXOSdWvTL8cjXmABdRf8rdg1YJpD6tNgcWUXSRgDl5ij58erliFvsKr1zU4At1RzM/UX9haLxhu
ECl+HOZNM9BH5UpFyRAbP4lIqCIyPEyPuUiaHcCJFCkwqQHsPMIqesdBzNGpKKZMIe1Tvkjpzj5w
iJDK9kxJihaVQ+T0t2lHcdXt59xDHNDOiuB+vfqWMlLdZeT2YAMQ+5maM94UmeycuamK0vFPuLIf
k26AWyd15bMITp9RByOTf0F5DnnWo2oJFvALVkqqTonGVnHKyiTtL50POIY5tS9OSueyivJ+uaEc
0Bc26DH0ajCfs/2rpmJsRhhrWov11/HTiax+MZb4QLoXRBKYds8uFCQ+f/8I879TwSdvzUTiTRQ6
dezFKELgHSahFjG8QPeHZpCSLeC0MOi+qlrMBgzH+WJu1EOqImk5KLZwqD3vB5fLkSQ58+leXT4r
/aflvY1Pe7GRbgABS7VeO/Lmv5wcBDrcOc2eVvGusF2Ew34TDkMWGNyLUwIshxkx9Bj/GHZ6UnAQ
ZV0WQT1sRvmXgJWcbPvtwlTPgmZcFSy1WEYEByvl5i3C6Sib0LxQ4DimskLwKDAL5cUfD72hND/y
cUr5iBsK0pir7V9NIWU47Fkb0fLzw9BKxqVyrZj3bJdtSstcuBsdFS1riX+l/ArYJR2wz4OOW6M6
2IftLtC5G8qpPAuy4zE/Ynfdd+Cs14/Oew/+aQlK6tus8nN5CrXOM4NrjUQ6wu73aKqOc9AK+Scs
aC8XePX7cgjg9K0f5LhTzive52VpomgL9RoDkGi/dC+zOLB4kETME45CBL93+/a6nXzw5GMZ4psE
57AZp7RxZVByFiDygGaKzaj8wY8YKIBUp4Yn17MnlAeMLKgebFjhgxOHhXXRJg0lxE2JMDwx7TKp
Y4EdSBnKNJE43RnFi0b/ymXfwhIYoCyVkKfD2zLFyX8CyD2+9qC8mgG9Yfl17imd0rxuOeeITcdy
DcKzW9HsndN/FuSP9KYC+9poXiJ0JVhExfxTTYDZ4IaxImggj20/qXX8dusbF2x974w6pP7H8ag4
h0/Dgntm/+g3PImG+9/VPmgIyZksXCJP7qgPFBUEEziUvqu0RQyEcOjDoVBh8TN0Y6oyTbkSGsJK
Fm6tXjrWojA/zV+Ji047pL1f3Y5NnN7C6dAG1yqjSVGPzmeDwaoOYg6tzfmHg26fu5SBtFPHOtec
pH9PdITtJzzM6HEvDEVYrPaMN2id3O+ZwOah1HJO6ZKS884NoG3LtGhsszLVZ1Z6NHykNUI0lNZp
eRsSQmYwDSB30l1akmPd9AB8TdQeqVq6T28MAdL8mQUJXvImNqXTk7g+JdYIpuYm3d27d2Lufigc
hppdhYlX2zRGMNkhw3XQmshdiInSyY6MTRwjUOc/97DBFWOucYGkd8+q18E4RzTXOt8ZSCKdj5Ys
B3O/UpopG2xsNH0OE4aJGGnE3kE/HwCDuHZs9IBVxusRBJYN40YDZnKzRp5mVg/DABx9fMm/GVLY
iVoMvJPw7ygZlAF5jNr79OWKvMePgPf6nvOopFP5L4eIzewrnqbg6YaMnhcHpZzVMhJsCnHDOZgR
VIywRaYJlVHoXU7gBdNdEpE7S3l/STdwqgM0Fu+nYlthWRTZvDEVZIK2LRNZnQjMfIDYECX/MNPc
k8IJybL8nflvMz+PPeBZOJXT1txJxevJ+gfmte91AHJR80FdM1cWeOx/YUs30AQHdv+X7ODJiCRn
nuUn5AkoVMH0ElZ9G6+qdclpCGypzilh5PraHS+p5pSe8FP3pgqZDGthLKDHWtG6Vment+fBq8gt
8rs8wHLEXkQDOZk21hlWVnU5ZPm6/NAM+fXemGE776vTRAw8vAfOs4qVcsoavFZGbv1U7NxWxMhF
BmCmlhfYxavEE9MrvKbFWQ+G5ebue3DYCwk3VbDMMtWtzoxefG/y+IRRYq1ddfjg1FyPo2zXcY9e
RSGTOPeAhrAH19SZuvkkAyUI0z/r+/p2sT4khisGlVym0PjAzi/PeDtt05TfvHF4NRpQvubsdQhv
BGwQnsJ8dyd0eB9WGmpmAJmgaBnUHZzLspPXYmKUAVRGaIX6siBkwP++VwUvUlwcOMYlkFN6Ub2/
fc99qwdSSPonCjONqeMMODiJuKcJbg0Koe+RKcLSJb4Bd0i+rDOK9VC4qhsQl8okNgnSkuAc9gse
E0eiQ/0JE+p4vu9+oIFB0xDngsfs0n18nXDnZrjW9EvNN7enzu/T97nU0uTQ3HXHcagtdpGL+mmQ
H/kAqzY9q+s4zqRfWCiuZcwgjDpW5HjWc0pKI38wwe3qUFVvk1fL82UOX8OqkFwX9TiZQxCssdig
yVVy7ghienmK3TOehVWdzziykDYCbOdzcBOii2PXxot/tvbKY0U5W7Ch3fD6Kh4LHo/o/edwjhE3
5oyIVkKo5WNdz9fPBhTAJhEjjbDZ3Rb0krYKnG/CntopUA9RlRT/c+jJn5R2XQqTnBrpsEo0pe/o
3njbyII8CqG7DWGa5Vk/HDoJq7xAl6MkXB4Hq31VEpPz/oZYylWtstNK/u3Rt/eez1slp7mVIjOL
uuhMglZSzdxLvdZ2yNFsoy5FmFqcjDFWYq+Ix+8JeCAEMCNIO03O/xiDszPlzNeZBug05oLVnT4/
e/MiTsYEMGEijpv529f8ILwy8cP+UWbKSYsJHXi0Ad0J3MO5NTDNolvFEeJQDTrSFqQUpjcbAWAr
jEUjSPQb4sacBHquqr04DlkMUfPmMSLDBsttFs4g9UQ2jvwKznv0T5ml+kEe27VOPe8Ei2/1WPjY
gxtN0v+B6EFF9kQNoBKIwFyaVs6kWhBkWYLqejgrd5qaR89Pj+gdRuidjFOkvbQ6aYs8bUtCH3TR
Cvq9S3CU5y/HPugfQ5xKGmZacubXLPSVj/eYDZvR7ma6OhOmOrzWyNqn1/m7nm/ZnW9Ry0iANZ5l
cMyKYGZgldOxDP/s8zObxtZAgVKhhm4SQ5X4bLJEsMUVh4HGbpmzLdBk/QDPXi1IWwM1KHufUH91
z6D0JgmsI/BmLlChMV8ZA4Yq7i2Cckn+ID1jzDygnBq3uj/nyhf/z9iF1YrZQvVIbouDjjFjoW5q
MKsrI/KR9fC1kVMgxSdtZDfvo02DBnLaxumbtx6ofj+507b9x6bPdglg3+bRrDkUbcArmBRCvH8x
lPFFe5H4/M3UekN4a/wXKbijq2ztjAAw1pkkOtjOBedfsKEu7SuvfJTUsYfnW5vYhN1iCtScbpYt
+j7vK0nAfS3Is0RyxiZA7+U2A/BuVAcl4zD9D2evtJL1MqAMKD/w3FIXPd+0Ii6pl9W3U2J3MtwR
Aq94VMzQ8CA7T/SnR8gZ2uSmLMaZ/ga4UqgSjWKiL4LY/6LxGIMQWdZ2rZuxU/BQCgkF8FfJq1qE
NhAeEPjE0efT4tssu27lm0XysxhEIzSPLwY64xlNzDDgeBVxBFxSaIRflHAdia8PSk0eqLyq1NWf
+rVNtarBwQzW0nP4XorzzutJHwOTE5ZmYmWDaS6XwCiBYQ8wZbyLVvVEgX1b62gKGo95Et5pW7aq
fPAQW0xRBkntJpLKjyjRenbVADe5NoH6mVOhhVbZcRsH3BkMdJDpOpbv2fHLI1bmU+vPapu9fBEf
X/+uqey/NUpXWBvCgcO6v0WP13dUegpE0/kHkHSEPvyNG4Chh1wbB6LJOTwLKQCwjtO7qdRlly6A
8SqT0OS+5t9vIxWAvUTffVLU0h+PG3O9rSOPf1o6UcfSLQ8+eMyhvABr5quZczc+gQss/7bcI0N1
dwXYtmxpRCWTdTD4TKrir8OX1RcZixK0NA2QOUphBNhdF6peFyEYE/JSwpBXrY4XocZVsFoIHKZV
Z6AW/UEQOZ5edgfsG86GKrFDkDa4DHw56/cQGiklUi5rRFpE/Z+qxA3Hgjpi2Clt5RpH00k/+rDa
7CRpbPhWOk8aG3RBcLH7aN4dHLgTShoyfnGWjJlwO2S826ZQQ4dPk4gDuAKQ3xXsFfWXcrQpt0h9
LQqW6hZ0Txg694HelpO/8Ptkx4eb+lbTp/27U3JEPQVAjeBdG3+RmwJnkQpE0kwnEQjxkeyrKyCv
8sS3T+9PYPmPVAHvptw66ncsWIYi8RAIUtLk0rbKjaNZNf57bP3BH9ez+y0caszwJy+q/zttyJkZ
++0uYnGjxHQP3e1q87I7H5dwPiy1B458XxlzsAvbi3YfkphVW5g7/EmOc8YqyhvGbAfSuAV3oqWP
RSbcuJZMcN0fmKJHyeIsrGsCwkBtcG6B0jjk/L+7br47leJxyMleT9QsELQfuYEi1/Zqknunrurl
be8am2N5NYKW4CXeCEwScCs0om1bB82llYbAD7lID4kvousk0l26bTiZq97K4ck2hHNAEgMmoT8S
10tM5otAtRyalxYJijUvw/w9cT1IXgnPzCI6twUSpjLlaZpqcXuntHRePue8FmzZUxTovf39QzET
O0IRWFAe2yzdyynD6wOC0t9cvkdovbf5rZ6mP90k5OkycDPisvDguzm7NY+ifQCFsa4L5a/4vxJI
1kkcRUjOu03qhujB+vNqYckzlORktLB7hLrBBWIeMBwEJbAxyK+jgpWln9Yr1izy6KOVNq1mwSwJ
HaNo60Wgm9B/QQHM+KIO/EvjrzOXMbqrsCyZ21i/QM4Be284lJp2o1Ma3be04Xx1f8dQSASA78V3
ugHIzb1QEEKRXSv0RWGYogzIKtshYoFGVC3lcEHGGTE0TZmOUBpx7s/Zg1tcPW/Hqa9ZR/5+iUEe
MPottidF0TaQzMozQSG+rBI93jgUgWsmwFxXlZ8DGfUJQVj7sUhNnw9QMkf4sLhUT09wD3gkTpko
99T0vrHdOgK8Dvx8pf50pmDX+As3q1dManLsMvNTfVB9eZXoBIzxygj6XCVfLCojsUPVj5NXUa1N
cZhjdNhZfCVCKV1vo8pUy7YwAKttfbhtBvBzGDDp5cNEiA7VcAgyFAb3ttBB6DPL6nP1yFrdjkY3
Cq23Tg2is6PMZSv5DyM92TA/GYxfp+e575wISIlnkoBIuArkfxi4DZri6euHFrEIG3FQ5fSbtt/t
4T5j3PzfzUJRi/1689kModOgwJswiwZD1D+eCkSVcIxPFr98IgIYirSyu/XP8FOOkemyBn2VvIki
p1YVCpbCFdVoh3qxfKarPEl8ZHDOAJNweQj9rPsQKzmoP3S8O2V/uxrvjMcFZxM4WUBWm2bVqCYB
vqchE1x39zwAJTnMr6nQ1luVta3+V/BbObWpK+n3l5zJbbtRsVfhpK1cHp1hTaKXW5LhVdPq6eLA
cUHaq0MBwXeNuV91E4H4cefD9yC/GZ8obmlycPWGP/fVWpizPJhe3kRDYtwQJ2/ui5EE4jYMsCcI
0xE/M5fraqIKcg269J0r/wc9D5RD/mq89eQ4Ohs5IVvyDbqO8qXxrw3llbv7bv+ZJDfmmzkbhqSR
1r3+gPHXRO4izi2UFuXe33MIT15E45y8Gg885ve6HR2N0qA2BDgRpEBAkTCKfbd4o54KypK2bSAQ
2QZrP+5cnT8feuwQ1rYTt9eFoGn9sRr6qoxZqs//9zuMJrp36NZjACyTJ5sTYWsuWt6U0MG5SYYy
Kei77+rMc2Tv3yGNctarlBtGycR+rAK8qu8ccFcuz/sZu6StzTYrm6xXZIFbYjB49WhewprnwxcE
odvn9D6GU3w9JswGmu9CxkZPnYyoPa+WSjdfereLeaOWmL7zq+/mJSthoUjSczaVJx2rWJrSG4wn
pbyf5VmSi9kjcsokYj0lwBWEIwlH/xz35hFi6RhjewqjwFvt1E+F5fMr4l4xzaFb4cEFm83xt7jr
ulzQHuNAosncMzkEOd5N4m3a4uta0UOGzsonfetH2LSTNEyJU8V55D5qWTK4+PmLClSfoh+tlM4e
I0YV0HpGK6I9Ua/GTD8p53lyIz66wqZ41AeNbxvfuhPvLo4+ck+nLqidpihaMllUWDHwOWkuBVP3
UdangMwqYusSRgzSSnIxpElOTd6OWT731e8XMowrnQ74m/j6m2zlhEW8bRCV7j/NE9cv++ZxwVro
qm5W9GY+2EHWrcbxsVkqPW4CHp5FZ9PJVgxNx3/Z+mnJBHUE/2dB2iyZYTosb4O6Inw9gJPlvZsP
7B4j4y10s2gkkJDLzlE0cJksh95Eh1eK+5Tnn4kfZB13/F9LMhLxRU0/+RnDtI9K43xx6Hv7hSLa
QHEpfvZeAAXu/H9MXEFmTGSKTR/OfwbIGq40BXh1PyI9s8NZcFDSFGqUEnpvnfpdqZIlhMEbaJRS
vFyXLikUqaWSMf6tdUVInvzUvoVtw7GDnDaSylrzzIDPvFYjtmmM5/8guxxywXHmc+ViTARQyPNV
B7s0p5C7dFYuyGOWNZHeB2vCSLNntnss/NxpqS3ABACHBKJi0whto3EDWI7Cy3r8uriuq+WdRUaE
C+AeVgG1KCyKxZIvBOTM9eKyHLVYtjKanldia8t4JHy0RujA8I6EF8GtLOwcnWPBWpb76Wj3L5oE
/sVF8IIajJRnkvmPUnkktzKpB/ng8TXg40nTglXr/sOmgiTup72QBlNVPtNj+qflfDsCHqJABPg4
mDBf56vKFoZl0PhCln1b2ZiWaH+SGeB4Zxk4+M3vngaICL5t8JpAXUByUUgvfp1MUxiutyqhXu2Y
/+ZFDZ09FFbMgVvpRRTBdGtf5T1cdBW3IPEHMSoWAAKADF15NB6VoUfmkRdI8WzlP1BWV4vGjyK3
CIKKDKQTLZX0T4iYisKLLCf5Yhgo9QUtStSs6S7vd1zqxFMQePMZfySJ7qw0gfZZq+H1XQxr55Fx
gqOTX7FkGM/pdEJ/Ry2HzX+ziYhcZFhQRZhC3g3QtIJuAOCkPxBxJz1S0X5mYZHcCvsb8LHzEOTP
5KhIzaHfZUqNdhk4WMlVmh5B+xJTHnzjHZPXcl5z/pbUs6C1vGL1s7C2fwXTK60UP7/L5R3UvXsU
poXjOoE+djQN0kXMOTt9zu5Ko5Dhi8ArrBSZCs5CYAkhuXobBqNIf1iWH8zwtcIW4v1WjrFipSk3
bVE7kMn5sPZC43QPph6vHDPHe7/aYB3BBbqstwaYKrmnNELJ/6gleJi6ypPMWKSsKBHLwwRBgPbW
WAz7pORO+jOamcysJ72H5GC2x7idPqTW3xOyACwS3PmfoaoJqC+MWsYdxicEUxam2SAaG4OTX5xm
n0QQlOZbGAN4Cqz4NAwrjAYbwS5F0CgPz1hHadB8cZVtrmEE1L3zTXn45XRzSFEZKt4MTf58I2zf
Se2AzPA5gg2lpk4ZzDfhpn7+qNR8Bi8U4lV//lxUMdZRJxuw/l0R05wLnBO9XQ3MLmKci5YePl6m
Z/KEu/0646/2RYKyx0tzOlhpid1OnKj20RDRb47rhbzJgQ2ut/DQJ0YS0LFZNNMSEf8MehfEVPQr
45N+fStWWHMRhmJAH+ZPDMpMWauBG4TtEqXRD2fTTDdI9LHQeaV1sBw7Od4piiR8yIMgpzmcIYwF
DZXlZSfKxAqwFf2xz6Yw7BVBC+OHoT713FKKC0yyWLoXJYLKHAwOArzlfNoRTxcEd6CSJZ19Tk5F
ilnJDyBwNofcgQogvWNn81oFtRYoq7wpbHSqow4Z6SNaWniWk0RmaRgwRpiEfyO5/YtKZk++9TU+
9VUH6rdXn6h1XYgwwfDcjnv32szmmzkhNccItRFxkBlU/qMQr6BauvHYKflsBRG4SI7uCID8CYOP
dnipS1LiceI4BJI75sI5dhZTxPpncp1a4Uyn6kA9wz80BUOG8KN0LdR5iVeqturBVOSpsYiGjPV4
XPURqvDstrMWmekHb76wzQOFgaHvagY8b1mPswLTlKOGmW+FY2GUKyQssPm5rLzxIUWasRxWY/X3
+IcbhhpEKeCJn+4SpOB6AyX/36eqUXiTEJl+e2uw9sAdglZHXYnBoSn/Jkw7wtnK9bM5u8frfOR/
LjFhMYSg9BlKUnWpDiiom4ub4FHYuyof20GnsLrtRiC1QKITpNFR84hHZ8lQ+Q57IuQk5e/g7Xmh
mnC03PessFzUn7TBiVs6qNi2ECHJVH8ad8XAmjzDWXT63ccipxU1c77aRKlTxz9Qp61q2LGuaKur
Nxf4GcjB8jIAmdJjgdwpSElfyIYotEisfgI8YTkXQMiTMFZSCGvxh+hOOFPN5VgSqnRnbhymglAc
eCjj71xt9Ssio7FQ7c7caDTGKgi175Ke73s2cWL9lP5soYaoYxUFHzLPs8kfJdJf+YnQlfsX3Fym
pfCMIVz83NrO11aATwWR9Bmy77OEAg0dkD/r3U//F1tz89VpvxYAzNsBETfnMkZvUachQ3AQI/zi
w9b5x0x+pPvEhb7Du5WytgcIFU+ZyWfauul1ofKnwYWm2bdM4wVOIXvMDr35/DhAgiQM/iOajI/O
3DmfOjC6Qi0OnPp6EUOdF61BVHZl10hqZBmge2sDuTWQY6RcSJvi6PkFVW3AAgFoMInS4pjwLxW7
F/yXfdiaR85oBglR7KdsluxucIPDF3Y42rm6hrhn5IfO4LunFT4q/SpF9zuvZFAH+qjsBaT1LQke
53nz2Pr3WhUY1Nob8y4YA40TRPhkqkK9gv86uUPki1p3auFFL4Ajq9cUJ/FnH5C5rh8RmZorFKk7
g1YyMjflpkhDj8N5ScYsmKT0XyyLGgqA404F06E6cy98Xql5Vud6Y242h3UGpJkZFS+HgF+mffNP
KDrKZAMe3HcPIyQIYW0yOUygdsLzPwTAdBdjcs/BSqvmTVFNHb16zThPv+lKNuwZI3L9Y2C0eOc/
CpanaeH5p6zvAEVsnF6gwjWM7crQBPL6O/onMXTPwP/d0uprpOpxdK5dGNX1J//qEXHFlrbVz7kZ
KWd6fNQ7HHgPR/++zho09rvveYSeliegsBhaOaO08L7NILHgG31aiqZzyAMzezmDcT6QDg8R4wJn
ggbMd21/xahMCQdYDZFVKQj+2EfLfKd6HH4jjxg42lFIuxRtUVQtmm8LuFZhntr4VCbT7m2uG95F
4iXe4EfHd+ZQx5TUWAGapm+Q1Mybs8k4bw38KBwcDTygV29bPhFqT8b5kH+yln5RuLG/INUClPzm
loWENK+XEI3ANIPIyUgdG+t2OKAW955Wsq4t0B/nWLFIDgRsXM6O/JlU8av9lDTaiAehk0JHEA8J
EsS3GCDmtaDqVs2qMakzHx3UwJaPliREjxsSiTeO4PwHTzJFRersG+nDK1XUSvfSW+yYjTFpkgiO
8SFWNoBS7kFaA/dQc46G29byd/oh3JHbiXBpvze8v/sghBLFRSLCxhYGIAfuvrNRBr5+nbQb7VGA
z29fKNIeUYGCRCYnx0iWMWk36YjF6OkxDvC0m9xFEPnz7fxs1r22OauX2N3W0lnIar6+OO4764Z3
hQbC/3Loojl565RLuDDsy+es/0jE5uRDKReV4xTWtVvbHrvyjaVyFQjd2WVDqufhB87e8tjtxPjx
WxkHFtteoptZfZAv9WkwsLI2SOy+PlaD/IaSKZ03lI13qQk+LGlMUUYla1DsJs/Fh0p+Rg/tR9Ku
7LV+SoaLJHpSsVhQ0BbIwMKkF9DBzJ8U0/bFl6LEPXcGLK5iduQDFRwTznIRZe6M8vNFZYCHm4OI
VGawYz3i98wYzfCa7tQttD8aRdN/rLTY5+AqI7NFs2fEFCz9VAfXSsT2SmYdfVo3QsjwD3G7wEMX
NHs7NwM1ctqgNg87kXfwMLwD7UY35TLtiE12mOD+NurSO30IZAAMreD/fTgXcoMWyQWowkqhuC+z
aaV9oTR0YOjBs24fLf/S/1V2K+LO8MDjgMAmPeHjRx+YsEh++BCTgMT5SlFKnuZ1FiW9pvgY1Zt9
h4AVDTFMO2TSZbYohtqJQrHk61eAqGF6P/tvdpbYR6Zwfj+Bz91nMw2FLXDVdPb7Unx7AgEJufnv
1RBBH6b8MUr1kLGkBd1oZRC4wFrB/RLjwgI6Ykd41TmLzh1o/nEe2KZPxIaWfeUGn8zFvSxX+CdL
Iid4uAap1yk3xPmvQlLEG1FxTBA42hmM4Pp1ErO+P1jMZgs8ktO3KxaOrc7VcY9Y3w9rYgTT8h8F
sEZfEeY9KrEXjElrDbj1cO9X3RLqJhCOcruAV7jediHGNNRbYJGXr3mP/qgDbPHFWTOIGrt5AntZ
X2W8jJMuGR8F9cQd8xG9PXB/zDCFsn3jEWNy9xHvQfG/b3KKmfOZG5tsoT2XMuLHfTbk+A9wjSQM
MiEVZC5GbpOLKo8VmVEyEspoVjriO2kIaIFD/9AlBg/W7gu3KSgQ7a3G4IEebmDmeDkgNGQg5MJT
9nrQU8V8ydCQY+AK2SqCBNRBvd8s8qvF79dt2niIpyHzCpJwx80og4SjVpJqmvauXBoK9kZRq4Fh
15ZhJOwNtDBmXV5YByLlzzM4nOfWC4hfW8T/Fuqt9y0UudXW1jIEWWXJbHpYvod1jYkI9jdMOoL9
HAnxtXnNry0p9FVzekJd5OluAJh/maiuLKI2wJ+LHHcNDXw1bvHgH4FwLw4eCHMFCaQiqTf1zHql
Q/Ea7AAQOdYpE+TasPZ5CtuHVDuEb/exUfj+43Bg1JLoDlR1qCb7VNTg46Z8JUJ8atdUTHaJFbTq
EcnMKjSxNlYDV5e8o/NR25Xm/HsQJzvujaOuKcjTr9iA4qw34+38tbiVnTfuWlYxqHArx6Ldn5bR
MbKHgS9fDkLtpSImJqwYL3wJ3BLMvBpxcwmGyYaAP7V4QRzlJc2FtcsMKdup6eIvZmVUexixgY35
3e1yzznUJCeUtfdvbLtxHcEztTwmdB8ryzdqiHvE/202wWrakexvqAq01ILI+hAu0nDlyofCySk6
alicUjGe1cDa8U3HKf42zkdnFlsHhdRM66A+tT2OkOpDhtKdnAtTGpQOrEnstUjpqkbftq72FZaG
cmSSxFxKvmzAPGTGBuAL38LDs7jgNyDo2BgBPD3jHLpOiPZZlAfgILYv0dIhSsKGNNEGNZLkzWHx
qQFbZO3okeCUcLhD0iUu570JOBZzWIabTMODhromB9iQ6bEvU1zYvkMo+opQ56h4Yo9euBlbF/4R
8sbyNmX3Dk9sKfBnFpWv4t6ZFsRRSforyxIHEI5eWPivjd/GtRQ2qarIt26hoJfjA9PcF/EUmv1i
ymSMTcLREkKKF1BqgFvv22t9iJ3jiCPnQMKKdcvgeMd9N6KdSPv1sj8p+jTQwMjXOD4FTUFJOKwW
zdcEXouoed9+xviqozEljbIwBjIfqPgvZw47uxchd9aHn+dJrKj2lcbY6/lROIuNp6okQIBv52m+
Yu9vSf4LyggazSpL8/1AsLhaSl5TenwgAMVCCp2+TnlMWrRsGb5e6XkZOuIq+kdpXNVML4SQ6K3c
+QQNxxWHtjY3VRtFzjPQWs9uQLTb0AnlO+8FcPLCeDqAT4bglpJpjrYXcMT7sA5GhU8YfsvOPl1O
WzDhn5FWin4QwbIOvTy+sMLSyDPmopnwKEaskrlQmAYNIav2ucpubbjeXW/6Ngt73rAAi1zQ6qbE
eR/+/92nmJ5bBjhGFGHIAtWqkSdWl7Lo87rSzOi8UgGdWO4T+akRx09JT2kxX4pqE2C+c7dgRD30
G8uasNQHAFgUUv5bvjm89ASWx7U18ZV3hSSUgZ1gSjmtAAM7+/2YBMyjNbVjtJ5eTlpbuO5Srv3C
71XOksyQ/SMPQRXkIx44xjdgxtKjvXPs99Rk4sL+2/1tdHZtZyzLz6wOz+L0C4EaLB0NFt0h6XN+
iBjyr9CArepPFQWICCrrZAWoPbBw4LFrWJKAcUTCMNewfOXfnku4GQvmdz1OOWngg6GOtZR8lUQm
pl1/imVMbPumNQy9d2LirlGPW5vL1j9+ga7hxw8ApmoXr13R0zzmiauKJ9V7m8rsqdBNirLk1jy0
wk51odJBXAHqx/w/wIjCNh2y/rVpcwtwBKj/EeAoZ1lEaSf6WBktbwFHjKIVTyxz4fDAuw8bajYw
KzbrLgGLNcDkqfsMNmBuVLXkGaJnbNT6rzPNhTewN3hfYnCXqJn2cwWeEvzEUGrcvp6NDJ7EedLU
AYZjfwWG8YwIFGkBUxZ0x1mBAtx1zc9PgFLEA0RrOyMQ4bPlLuh5hiB5HiE60dkQMQI8l7KYnW/y
gX2gueKeyj8JNxFiJ2Zo59nC1BrMHV/xUySqSEYs1dBBv8xLNLkD1B4cwLv7SocCGo2pfM53KJJc
PziMSVZrP7RB0Cf6T9L3pvNMQDvC/sETWz3aTmJW4h9mtNDrG40TgITsVtCMc7B/waY/tIi7cGlA
WV2Hf/JRw/DjF0XO4wJvCyOfg3mxyp41Jn2iV0pbzM21TopZokiPO/3c+0qD9ZEldkJ2u9HyLNkS
LWGMelRTc27xsQ13T8oKkUzjyrlnHM42OdIFrE7zrvkrqR/OY15mTpj98n8xLnM4rj01MCdnQK3k
O02B+T+Njd1oB14+MnttQv3CUZCL1uddTvBnXVDSYb8oglVao0WQzFodv3w3evudWLsNAoU6JJEw
Yoyxq0YOYrhGzyqPK5B6Vng1iIvEP0JfSLeKSTaaqBc4nLyb0sYX0Np8dfk6sg+hlXs506WmQIDH
g6eGMJ0lY52fr5Q2cDRMdb/sxRjofm8+rtrNdks3mnyaJQ5CjfF1udGu9WC7KdhyMZPUK8nHHvll
34CgycepZQHSx34aDuGJj33CzGGM3EzvYVZiPcQpzcxUrIjwrZGE10e3iDrMZgs4vWcH93kCnthg
GEBLQ12lnOKugQa5yX/K/34PiTx0jFsipCTS6aMuSF3heR4rvOR0/nSb1bDDdpq1jcB4RojGewwQ
kKO0FC2aeA+VgOGnKi9z2PgC58w+U85HnyAsu5AYiWhpqHUPEpfVx/iHn2MsYmMDfy55pBMnFdwl
3H+lJXKIw8L3c+JJN1hJloPAl5CjuYRT7ckZuXmX5nAfDbYUDIR4STlAcSJW/aPSV4dPuhrNxg7S
kbzGvzoGccbYtwxLxulp+L7TvnPLCFN2rdZcfst9fCBO9solaKcLuyQcFxdMYObamZnZ/yYSE/Ay
w0oaULTr3teAPG++74HpG0FVMJn4z9Y7ADE78nnJ6sfRKaov+Poa7JAZhGNGMqqICZZTBAFhr8wc
FqC6Hj9Bu5F8crk4uj2uFK0gqDG8FOzAV/ctBEu72DINZc9pW3W79aj7n/U4uvNk59lVIrwEropa
p8Wlj/M3fOcDkxh6dH4hCDhp0iLscOwmMIBjbpdj0pIRDQE7h7/UVaOqJXhAxYwRQ6SRCM9B+AbF
cws6FFMx56ChnLF/a9zctJuH/YJpN/sE9iMFcW2PkZDNNixrgx9fCXCZLWEm0OgwgWonFQWNUnqx
NQNKpzOwwME9APNglTGpJv7p8hC+UpSyQnQ/vbUYZvsNAMNcTmnbe8aqDGyUa5GVWbcMFJtP1cb3
6KI8Fwnuu/aAHJcTZcxzXEYZrf+57WV6Ym07BNAzwVdtPRM0hEcshjYJ1AP3GITidEPfxjeXITVs
fMGvnb8adXB57kHKwOwWR8Umkew4iQxTy7bLvyqmGCbl0zoAd/ST185IcB9VOQK95rk2OTOTIu8J
U7/4/TAk4JG0u2vVZO6ltLi8iD8j9EYiMPNg7s/mWXty3jgMrBNjFI/I/MX1x6appKdMaY1jWmwm
MDlLi/r7+ZjxRt3R/Fb6NUc03OPH9wMy50IpavfrwcdYkb5i/DVGnLjFuB/oNQqz2B1JXtDaoDoD
z5HY4rbVX0cWAFExPKGQTGQg4EI4WXb9gCkiChEZlmqwALjnYwxQ7mPVwLgRsHz8hA7MF0e8+mao
1ejcKlhIDnSiWDmhZuLbU4xEigYj1GX6NYq4HnHPMCaSmv/oK9ZwRJ52RUhAU6WevPC/hBJNJajf
2pHNZLGruXZig7ptHkHiWJ/8IE4lxjjQd9JA2BgNL3HeI5vfk2A5JZEGKCOoyJ7kpkVqcpMBiYGF
NgUIgaljcBQ52KNwAcHfeuBOqxVVyND326lwkHYOVv0JDbqbaCsPlf4OEGvewXHAETHclcGMlB/x
NcVyheLrVaP6Cd4qzbdZV0IW6WJMnblG2O6BZeXjANrfaPRrZrVaLNyM8DA+xf6Hokr1jbseTLBa
KqHGsFRfGSAKCf2bEwvKjHovJmgcVLjAke7AYvj9CXHSk/TT5RNMJM1UqiAvuok3MlX3IykHDTZv
5twDqhgzUVNroRN9ff6QnZGF5ACdzlsiSc4BiBIdSf2331I4y35yn3V1zuWCwABfHEB7Vyp0Vg5E
OoTO6gLnA1D7VpJGQZHbNXmbilnDRrSpa3L143dGZtdZJWbYB8BY7jx34OLn02Ntc/gFXGpHz2Js
54uo4prSn1kJV0wZJOIgyRAaAYk2K0C9F7fZ+vZOVVNeQ3RDjE5/Wecv5+Z/WPtGuBxoGKSer9jf
ZMs8+x5y8XDSZDKqLTFcZO3IyMfu9fdE+5kZXQ6Godj5vTADK0Z71zXG4+1ADIEc3hs1B0VW+3qT
bjG9jg822Y8CLzF/kwt8IVFNixcMNOfrmwwezUX/2QuA8+0hCC+qeSQkLgCQApU/NdFXMwvo1Y6v
BLHEfFOUp0qzim8oqRslrST/0FN5MIBY/DcTkU0YrwtwblYE6SM9Zo3kFdznJizfyMEB4ggMVLkp
YTwrvEAQRpbCxC2WR2mhFKWrtzaIp97XdOI0K/zx9MiKwc0tlGfaXxxDvq1mKrcxJOIyb4J5c4XN
/rsCkCk2zhehlHTMeSxJzrSzzfQZrKoFNHC77Bhbn6CfPZu3FWXDjM2iIfpJtsxiKJkZzQgHvD23
Bw5CAtqeLEvb7cch7nsSmxY7bafc2ml3jaLDVgko/EqWonGqmi2G9KxFpFny1Xs3uaRnTY/VAiXM
t4LgiEsbtcZBdMuRS7BvkDvOnze+2K/jxaaJNlyv1hY8tJ9fyVcVCuXKxSJVz+em60Go2OSgHH00
vNJzsCliYZcqFCRuRNGBq99cVBVBy3PxVOcAgNoz33r4FVINq9ZYhTA+jNlcYoZlBx825bDDE0Cn
FpFlYzyi7+1cFWxibKZS6Zx4AGCs4hRLz1UivF6CRlAPb5B7oDUTaeEoK/Cg0TngLkZxw7OxPCpa
KlpvlCAOsE69g/6KnUHMBifP6aIMePMxXKJs/hfR1vrkwM3g3/vrouvi3ajsSw4LqF0kep+JNRXz
1TVLUTpPDAgi3bfPLgqoxJhV3SRR1O+75yus2y0LhXXFk8dkDpW8j+ukQgOPbGLliJzK9lOTrEmu
eR6BDzzbuNhAJC+ZSJcxFIXdCSSSjNvcGB3PcXvRNZp/pdwE0vMIuOj422/mZ8HDus+Fb4lovfU0
xfpXPqY6wfhyED3NTPIZ/Y/RpWQe37sBG0g7j2SNLvUsxP1KGdSc7RW7u3or0Z7qguvmrkBobGMR
+ZxepVMNqG+3NisuuDZQYDYUZqZ+pYWcmGVrKTS9X4aYAj6UZYximRAZ3wdGMpoAV4RuoihdXYoi
pEdqSCCOr1G69Vs4FckjDiXUGJRKsTAqnv21kQ9SzsJstQJlk8zRirl3sjJwEwZnMiSP0aC8gCaS
j5qN6tCxMekdDEpZu+MnskyqFShvPqESw6+KS1mOlevewSQolDA3f1Pq0mKPqsDOAO7eT5cJUDRD
aos9MBVE6ViBWpDRQZpdIpE7fuvE0CF/WHNLBeEBP4ZUl3d17RVZysL05sklrOFUXqSQItveiw7p
0lJ3Xg23ZMwHgrbBAY6o9YJjikeuWkY8rnSupQ3yyycIKC6n64ipnPHlTUWhXyBWDPktXRt3v53h
ISuFuXKIIvAKFmDhJk4oyH3o667Gk7vrKNI9P32OTfF8WesOHlEUBt4GRRlkCDxyxBjgHKuxbrPD
BzOm8WYSAtlPFZlTTZBy9xxKjO7OD4p5wvEIKxLFNwRpkZ9L6gNkBF+a8W0KqUC3fSp1ZptsqGK7
pVfw/ZCXmj5VMPUBKLXpOcGAzN7m5a4UaATAxqqaM0Anq+jD4pwJM/3RAhuRaZFWi5WfF8sKPoh+
KTy9cUOdQc4UMXNKkc+FI8yGQXlWXb/ex7BHxdO9KHfkaeiwMhOPy9YLPtcbw9mo/pxBg0dwJ3WS
5W8zm9BWnlnj71SBVzMBDme9QcVS+ZdMSFRL3Mebqs1B+l4KKNYWbNduY6wrPC9BmAYHWP6mbx6C
GqTRLXoWhSFegk9CIWq8e9KGfOHUGo4saiySr02xNsFDjxsRU86QD9/dIxnf/3WfwtBjmZu/4BXV
k1HJwxpJgqMEbsh+ibnANDzsTas9woOXRv/xaBJ0EjpY4GEnQplBOchBGKOkag8Hsh7RFo2mvqLU
Bk2Kdk7M4O3BuUF2Qklbp8mGePUL8C8aC+HENIhy40wgbPD3wxKSXOPB4cNR7mYdFscvt7F2A2cZ
kf5zvMY386q7NG7ZP7cYJZUXcj/UgBxD/dO//bIt3RMTkBYyyy4BiUmcNJpQgayvmK6nhXIiIj7V
PasugDAWGjeBv96M2adTGhKJb7s/UqLSdZQZ5XYBw/afm9G0aP9xs5eQFtB7CSbqNlN84pt6mELW
4Cl7VPepbWe2XFFp4gaPkpf/kql4H2QKxNkYIlhDnQQzYHPoXKcGQ0S/g3wY+oOlP7ciEDj2Ic3o
WDppRQa231P915egP3QWZEHukhYsUdCFETXSqDBCpSyG1GRH9fQwq8PzL/mS0NQe4dKG1wdaZGbR
Q//l4zRUb42J3em9LdhPWdD9xUlHcLIixPKMBt+X59oYEacXh7dw+aZlhkG+xxIOBuU03w2WjGJC
IbJ3wZwOh4YVamATbh4B1GknJcZX9BbgU14ctPZkXvPa4+sABddddJbPt8uAvTKVLCKkufRkoBrC
8cgk6YKBS48D2CuNgCNJqFCEn2X/M9+zfM1SH3iUwOZs7t0J8+A/av877+KwemfS+Wvh0ETEVK7p
vXuLutsK8Q4LLgB3hjSwz0IIWcbn+CHYiuxP8KiHAt1PIBnaKnZ2WfBPogX0mhslDm85/zXW2zXs
a7GOC0Vl/++qv4Z+4DtmJtGR3Cq5NHEm0fd9oqw6wIIxgtb/MiUV/9pRG6PPeZBO7zGOh593CE8E
mRAoTUQxCFhrMhys4eTnWJB7+5VORA2IeDqOZ+ZXYmmtVn4eLoqfPh17bJjBzHY+mLpBmnMZTbXx
LYy4yTl0M+tWOB9X5XYCf6SoYf/MfSF8/Hq7FGV5iJuZYZxjPUELbdzCVkkZppxdM44ee7bq/G4L
ieqvz/TNseh1R/ElMcD17N7JEnWxWoOv0a9I7ZrYTsa0RZ+MG15p0b5Yo8yRsgzUXq9zr5Uz6uQG
GCrThJPQNsRzkp2tCEVPkXjpKMlJosM2aIAGEJImnVu5vbZe0JY4skFuSqEmSrT+vgvfxkBEnHyZ
0Ig2QnbxZtHIasDCHZN2kvzZnwhaybVsjrVnBr7GJxgZYECavOzbWCf2/TiSRWEBxKXB5n7mg5EU
Vf9G6VQl3LliSNe3JMBIv3qXyP7l2kJBuYzw2l/7mbVEvUm3PtrOoUazhkTwkqCMoYRH20PuJQfL
oqWeg6UAUkzpaHeZEARaWDEAGFOJ92rgpEhL2WwTnma1lC3Pk080sL1+dJkz/hdZCoYMQMMdJ6Dk
wB7+E6NGBKxEHgqtJIAGmGFqL1L/zLu0mKC4FtdHAewc5Z9v98doSCgngT5CZZwg80JNe6oXx/lO
YBvwWho1jXmA5BkxDp5XYBpgM2loFgZqjBcNslz3/e729mR5qWjel2kqoBKDcariqRL1ug+WsWkE
BVbXhABGOIuzwu9j6KEa9foJPnEOHPSF0jFazZE9xfJLs+GaEQv1X/fa6w0Sqn3nJeUmbeK5Qa6/
Xud1Rfuv2n7dNeE8vpKcYCEqousWUiLGTHOCSQGHNPNXPdBwJ0PdLXi/dlIjY9GPBHE1+j01aDa6
aGxukAGfChqdtRwqrJItTDQbar7aHKlqgOFZfqLrI8KBELjX2bc82Cz0CK+A8RtB7VWM+wK3J6Qs
Uch3I8TDn6dBHtxkR3qn9Bl290yV2qWTSaRYWKO+H1hLZMZ7l4PS7J9sSG+/JuWcmwbaP83arBB+
XHVgfIo+98xInbKnEBnc8mIXF8vWKlDS2PGzu1BXvNrXm/tOl7yq3A5aceRQW7fQ0A7Y1ygeCAhM
HOgD2q6lzFIUlWWxs0QbBqfuqjDw1tLgab/EqeqSXVlXtp0BIQCYdwwHvdhhUqg8izQcHI3PiXVv
2MgyiKayV0SD9czv10P77g7T+zmDKHTB2UM9rgOp0ptiaXVDmhWPQ5de7PceuWNedBC37/WVBTmv
hyzdKigMQQI0bm62JJRrN8xPqFWrZGZ4r6oppt0cyTh2Y8Nhp3djCBMU4YD0YPfaEb0pAK2AFa3U
otWeEjfejUIVC1r78ZPKm6k7flxCeT3mZ7vFvQIAoa6qZPGgZWE0f1s+e+eEqlvnIk3mqtZofdvt
a2MzYOlPtkV4obLvThe1rEIn3K9Oa+abA4lIm5GdFomQnH+YmI2TayJ9UREV45iWVjdKpaTu5sGM
zeYaPUUbjZqThfpqjhszWjmOVg7kDKNCSyr3Ijm3D1CvMxZFKd+RuOHDQsSloGzyNfPfGFSfubug
eS4h0IsJcMbB4aupcY6vJ53XvnGm1Obwfued4vUmIkTwy+SOcA/nVYgrxdOOH31hHcbQrLRRXBak
KxPQ+/3w8hFevAOi6E7dqReNICJdCmpOC23FOiP2YEh5x0mqhKj4bneHMksJj5pQX1MsxYsQLWCY
PnwZQZmKV6GLnjxh3mpLGt5tEmg4V8p4YT7bzSItyKGp/ZxuaVZ8wDW2lEk3A6Ximz7geZUev4J1
fXeYnB59/apRPYI5fx1XvwUBg03Br8cIuA5nu1zVT/4pFqC9IjW/oJMM+V58E7lbFaEVoF6rOW25
ci9wYqvYp2RRx52vSflOwUCgCHgoyCBzx4Ur3N5aVMGXN/tDNmur8ypXGg/kfQVeeZwSI1YPYnHk
wfmmlGA/UqgNtMv1101dwfPxvLFNdVQwc33uEG8m9wbqD7piIEUjx27Kp7Wms5vrxfjHXGe6QDtZ
3VFXfD2MEUcr9f2/RhxjhWwmZgsNk8hcliGEQD8UzDVv1SDgw80seYC0Iu0swM2lgIyg6U+VkAS9
ZAJ7GtZcmHqfCePMBvw+9BzQ0edsZIMtqA5EvFqjJv66mmn8NjhR6b8TCvoMtXuyxsWo7HsuWR0q
ShRMLaSiI2smfkLtBr+Gu6d13D5Sfln45+ta1aOYobwcO4qDBlGFt8mnUSbIXW28TUUlgqprPoZv
GZE9j5g65TaWuLHry3vYMbzQE81Bg2pndl9NVLOQ/iSLgjNCRuX8oseWhr7o5KJU6uz5O/tyja79
Gn/ejJSDePkG+kMhn+2bOqwatSGTCOMNThfOnjqfi3YUQxeahKI6T/KSEbMUInMKlcbvOlchfyQX
smj+fZ83j605hXf6NHgB/BpurWPrxekSc8uz+OuXFLg+a2S00F27KhqC112fOAY9HJ5MIAPhUIpi
+/d7eWkJJ1YlQJVci+FgacFZyCaqmV+8O7WoFabd7PB8Keqyea6Bn1CVAUITsCQgYKaIKD5ygErl
PxF21IfTWp6pQaAyOlMIuGtgnMnhVJSHLW4IialTsIwU+1bFyK9dfoQQp3Gux6bY3vxPXYrfPY7U
bXQ0amCsS8bYlXNhZaEH8qVzH/opl/IUS5lUKgfFd4iG+tVkCbw2MKUwTnJvFX9EtsjH8cLRNnL6
36qJkeMIfH2IqOlkHiyGc5YvKIZkYd5qZxQFSrkTNABhfhPEd+MWhaCb2zpCXQU1eBwTTMXkmaN9
4YFazRUN2xplzEA30XbSe9Xk5Fo6b0gHNdzZJby65uHSYPzNNL3WPSUmJdo3yvknkucZhMee6oG9
b+9sNWA4gE70o1gDX7Ytdxh4BhNw18abmr+Up0beVPHvybzqa/q3d1X8jxesGt+XJVdebDS3RMki
/N1qwFa0ifRTzMP12XHNR041D1vkqJy+Qhyu7RHdA9eva3HmoRvlh2qCN3t+zuk9wmg8eH0zKbuJ
eNApXMFnfzYOiAN8gcQQmOHgkhw0WnJxxKQNIGHk2pJ2pbjfFvZ0KRZligqGEtlnu26PZO1/x+8Q
vfs+RmMTmyuQDeDen7tKUB+7GmR2UiV4BZz8+GY2RO9Fwnc7tTYRfhv8EDp5gFNzEAy6jGIE4jQd
M4t4fh6hKPyLyRC0Mlt4050rUbesAc/3CxI5IxgMECNG2j/mtR9GGaQSmtFsXaHUoieHIPC8wx6Z
auzRi05s0yREE3gYuEG9zokaFHgoA97Vdu7yq+dHiN4G36TvdYLOrHFBooq9IHntJru4J9nuJh/e
gAJnwtUND6SzcraZ5lZocpKtD2Ry/pUh5wuoiAUVmLOYQhKHE4cMwZUT6THzXie92GyVwKv1DI7T
WXO8dAEnVMu2tkCW1NUg0YKQa4hTFkLB/32AvI1d4ZYLnNXZJxHJ3WyrgrIGb1frqEz0IK4tn39H
8SGv7NgybXG3Yx1c8ufW6Tpo/tTg0xhaHmsZooRC8t3mEnbViJEqobkur0eebx/gNs8fVPoXqwIP
Tcb+v6MJm4XIJD18MgZLVgtTXolkEgsW/duPV1ByKqnOH6UJ7/jHsQruNdxXxgb8qvcv0MfTpapv
cviPpgnWhmKP5OoG25EJD6G4+vUFJM4BDfM2t8uB7PSz3nE9m63dHkyJlchy3ZagCU6CeLzTMzH2
XPdewDDcNzxDzirGcT8qNpl1dKwaa/4TbJaTBe48ZRVNyJ6bWLVFKKSB+HVEh9d7N7zingfmikye
P5Rs3GKfAEuORBe4/wuvQIwVrPi8zwq4r6kHFVYcNv/ikaDwUXUObANs5yQPUVTwnvr9Lbvizocb
osE+Q78C9pLpG5aiFQZo4BUrk9U6fYIhjZoZE9Va5vR+a0KBp2/KA803U2rBKZLhyYQCo0+K+ygy
loyihPE+1V3a1mwbyjfh/HuV9oSB8OXIM8/GDKT53kms4lamNahVVkJ9SJ1SgMzDATFqKpRCz7zh
dUcrh1M1bQeutFxqDmYN+XwPt77/qIAJOwAQhnf/afbNIVxRhWpTGayO85jLPE+YbrKG8c6r0gu7
79kfsGNoziJA9D/6hsuNJfJot/stZUdyMebGc39mOEf18ncZev0FdR1IvqHIZpZ5psFU9PMT+8d6
vjVhQAG4Tu7I9lk7sMsHU8AYwXsDR6c6/Y8SIKpy3HReScwDnriy+dIuSKsRu2a8toGcwddo9dZ2
XfNFQnAmh+SzmcSTT05MnVWBVvOE/a8G1h2zWC5l0EUbyJzWYSLcERbviPMXqARYJGL/ZQswn6MA
YUz056MyQYI8FTiDzKFhFYa35mnL6eBK4NoG2Ou1Go/LlSRZ2DTFxG8KOaQ33xduY2Vhoy8pmAyr
tXdOjTFnMKkD8WxDs9XFe97qv9Wf2VRz6DSUEC2t8IAZmdbTp9xfFlKuHXC0isMx+IRCY2QtlAmI
nuuOOqLkrVKBuhhgg6Q81lWEGHL/OfUpWz3+6WnfJ/yp/gsZ6elXQ8LhWyeY4fdvytLOCKzOpvKX
0O6ekl0UrotB52O+5T+6cfhp9FuQKmhPgvRFA0wtRwmTRrcnUFpbWJwa5/EzqSo9aeGvSQs3zDV7
3cA99B8oYrbQe60a7BVw6IpdbzS6jKJJKn7qLoAgC6FPACWHuIWgjnkf+sLMQ5/NFhc7bH+uxWZp
hg0Y5LoC81U4x9dWprH+TUPt4YGsebO5BA4hr5aMzh23WIlfAgvtoBOBD39K8srrYBMKwz+TDL77
bUC93Bsx6/8wKpaoi7AQZelg01mDFZGHzyBacSMohfEaMwoKdtyGnVS0O5iZrwbYbBPv1bd0Urg2
lRcA9sQsAOdZZdN4xpMM7yjytYljvOS7+mi3WQZayCon3Tg9Vbfl6EWaPsxqQQXM02vd6ObJ2RVy
i15Zpi9lWVj6yfor4rMcm2OUnTyhM3psc60/sIwPWVdeC3+wM8VB+O+UI16GVsQk4DCvcq9DkpsM
yaUB9rvbqP6pQc8VMeN+vZzpf3fZ8y5ImDo5at3HsfHHsImqmf58dOw6VfEKcCiqPj/maBg5Oy+j
8B/eL9BkGphpgGjODsGcmA5RC/KcXfUKWGvD1yiEJDrmBATv5idqawEn3VofXh5JuP6C8Z34R05d
9smJkQJBBNWbpp+QNroKDrOx99YMRR0uIOuDzWmDaJnKO5D1Y1oDM2/2Aoe3dB9kA0n2saZep+sC
va/HNaFN0cFNcmxNQIbYicQ82o4/1QOPp4CpYG5icMb1pAMhn/U5ul1iHzLBTmGyST55MSrilQKM
3uaMiBEd9teOiV041JiPm11Gn3r6I74kiLiUaiZM/erjMOnbCWqv6fehPPDyOUxU4nq/zzqAvYIV
j90/yU0UJFbDsRbqUtVEjBtvrrC7Eh3tV5p191WJP9aLWD3hquh3AOLr3r1mp8yZ+k5V/ihwPhqs
mdFs2grum+ICUC1+f+5qHpS6aaCeUbkLBEhe9s1Wx9Ioea8/2euDs7Dka5hkBw21PWywZWA54iyf
DQjTyk5xkaKLYYC6TxCaWopOYW4Gsv5vumoqnnKgR5F78ZNX4PCI0VBzveLoi28Kvqf3OH4XGGh8
Z9NPE27FbaxhnAADJUZdTKnwTryA0bzF9NW03Uh4p8WACmp8ReKpC13m9TMz/v5WLvQwvqJ/6qsQ
TBuFc3PK8BQa241V0weYzgrA00BFhbcBri/nqzcs6ZnGoYuzC5VbYaqkUuaGiMujz7mTG1pkMb12
fOorSqSPDQHwW7VSnnxW/c7xVvYSzAcJx1gdDwqMuCppBq/Jza4tbTfvxprGkloacKsOvv9eEEM1
MSJYUiJ2F0s2rV2c8IMWDqDW4MYMebTVmkKInU/mYFmlYVMxgkY504hLJCI3wA3OWY0woD3AZv/n
hlruIagLGTlt9kkI9WIFSpoWIGVpn74Qnp4EYvC06loKvlPO4RmniIHhthd/rsxYr3wnDPhtHhib
JvA6SfM/VYdqkFr8q7G/LvpYtgWZ1nNXYRXvv43AyVkjE0fQM1jUQZ3swxWZddFe0CEJ65jnyDCi
0U/PA6+X/va/+sOy3WTARdVQD3lT7OigXQXpVJ+X+Q9z98ppEGi6uOXetmq/s8Uy+IemvnGd2MDy
/3QgAyL06wIevohsWm/Mi6gXrjnWV9D8L2pGYZ/u3ySJ/teLZMBA4bACnGTGnsH67aZYoCXTLrJn
8POu7F5AqaD16qNIbR15scrS+2swblkKgbWFyDAtggUrotilD304TTOfL+P8zZtD+rkbVDQugKPg
qpANztwNszK12w6x1PdH5mOVOqRqPIKTuT76P0xqBoiMQjsvcwTUy7WgIZXh+HJZaWF+Z8keL2gZ
A0vJ7b+uxxGNx95wNqbw0OrY1eGp4WTFTu3H5dTkw8XXQapMJuPCqwb3eiqzzJAMdx5axak4F3NW
Go5jb+53af1rBhZIKnY7t8dcyEq5iqowMf8oJvYocwQy0dvvVEUbtzqABh9a2Vv/JdMXVoBDtopR
ngFcY419H+gWbhiqU9OkkYu7IBgzLGVI3iZNSpj5v2NzOSbOEoLuBJLhj3P4qHFpFnmvPJTiNVFU
CFgElJBwhnP9kmVpfx8Tu0XJaOT6wUlVF7Pxp+htGHmK/3DQlnqANVK5EaymC3yfNequEU7IXQfc
NB4WFA7fVA/ZpEkATXhXxwK3UgdbqkEW2gR0G5cQNRhs9onK5LqEkgaK7p3laukKzpibGodkUm8q
96dQiee03j6KkacWeIRd6uVV0VyHUNkeWFeQEbx0DfxN6rfnAS3bpMVA/Wv46GhvjKpynbUbCk/U
DCCsJ/W9xSU6VF+leFePTgN4PKnnjNrTCnKpCKRQ8s0WaMzRTAX1yRDRXy/j9FdjdfFkpGU/XgaG
u9wIhBZm2NppJESRuZXSeoErCYm21WGpj6VVH9pYjxoqW49yjXsMmVymCg4kSocN9a11tRmusNTc
/L3tniAg4N6ZZhlEGXu/voMpTd7QR72Kf8//yj22rpJ9ndUvdxqNq7NU3/ulj6+/CgAPVMDOz8IP
F1fuosL5Ud06odAR4CdiZuiwSnwF+2JMYmWd4vIeDNFJwPKSh2bf/ArSsO2P9r37xjGgx0XAYqeB
VbngUv9owFEF/N5gVk8Mnho8rQH8unplfmSyCweA3SkYI1y/O6YM/VDrDXW6QDo0iQ48lj8RUmR3
sCG0pYyGQgwWs0fnBGYI7vjhCSEwaKNDD2mwt4t657tMyEULO0s7dLtVgp+/n68ATV5N85w8DCmk
T1+GfwTxPa0wOmkz/C2s2eVDddsQah2bqqQww/IKewsD19r5LlQbc3PglOOzq77TJIHFOizDU3ke
vyUciroGSzl4W9jOjRTscDUqNJREIqQWSLcSGfObIa7Vo1bl0Gb4MMA8wY0gLfwOUq3D35CL6QJG
fEhlnsJcarEpOxEbVUH+wXW3NBKO5Qk0S5ncuLFS1gxoPvjfnYLw2Lbza0S7aQyFmnNJrKV4M5ks
p5Z2qlRkOpxIKr1Jf/vsRl6nImQcLKJUzbjeKSrXrK/LOL8cOcLaQ7wTpkHfPwBaVSiS4R2yu2WE
VFigtmbz5U3ZetjB5ywOGGfE1suFKdlyc0NMae73SOtKdGehrr4Pmpxf0/JRyCeB5yfy+lIq5X+J
8c1R1acG7oOUPRN6MvKq7woPDbyEWHq1I/NQjplW86EaF99B+bPBqLwG4fqEEElpGVrVmNerGApM
weBPmv+KXAf3KChMPbVgS0m9OYHpgtbVd10VMrR9wl+f5ocuwLqleXZIUU3I1zJMWhyshn1El+p3
doUHb5xvESbleQER3ExkRIEMCLOG7R5c5926EGi/20tpq3+Eqd5WZYLMWKFfHEADTpshWZ1Fsvk4
mJXeIoj0cMPeP2myE7UTuUYnizuU92UNAWwa3Rb/K2z3FkI5w2BvB8eTxZfKDwwlfnIW5kEkt5EW
1DIbZdeljKrlWNRu12XNustHeDoA95tnB2GLgvtWSp5Zk9aMsGU7umfmCKUtcNXjDY1WWAvROAL5
Fyri+3Q3v+/+biFhDSruKfeg4mIpkXe6Ms+hyOd5nPkAdHXKob111YEsuhwQ7gLcgPlotwYnzKxo
whdZ6np3aPSyAXylsNpj636n2my0VhXyLuGNoL9sTJoTAHEaR9uMF9u+FJqEwXTi03Zpxtmv8JaX
KmqGq2Ys00UT9RgFn4EW4iNwe7xQOTSiv0AnaB/VNmwsdLgmzl0QahUdp4QY5MBcOKcImARqJQG9
335UCQAJV9UgHNNVw9smeLWRZDmx1gkCq+DVm64I9yLt0/aPV9RM5Oy4Ui19N2OzIReIudOdEdH2
5nAeeI7LG7ZWUXfqTboCAl948mA9himqLUv6sWfaIf/0ij0cg8XLNqsMdXB/nfn8PN8/s28qmixJ
yaj2dJRScFawdQMF47TkoYs/gJeYXQPposF2T7x6k65JyX2FIsOI0UFLSzTP3k9wiq23ntQwFLam
ZP4i+A6YRXyns6HDH80KMZBziftSUGflMyRQ4V2/gQ0JgchyKFngpdE8IXPTcB/gJZTtpgN/GyeY
FWQmgVkrZb8uXdYMFjD5vgISgcUEdQzZRjqQJshuYvVChttL9/WiDez/OliFdCVODTR/2a9BmXug
H8xeIlIYHlAda2EC6riqKY1ZZhoEhv0UwUxuCT1aAzjXQf8dl92AthpJFIeHgvqV16U/RYQyILEP
MX7s74nw0NAB9fbGM60nN3DuB3hhtFJDNEDjdhxa75/1JY+5waK8b5BUs8VTvK1BxiPnbtuCxRsq
DBUskvEZwvKkQVzKstf5MrJjMi7w2r1SK6ko15Iyb4eF8taIFlZB3a9OrtKhGO75adiDnTr5brOZ
ikC6ZXct/b2t1zWdezImC+5zVsODbYDz8P/lTMa+qztE8PXMGM++tDxiqOaQ482FnMexlfnF8yWQ
yuiNmo0VNyl3OS91n6VSw1vxsYnZZoSMVrt9ShSDXEX7Azn+ifgRZSZHr8p2OSUT2hsoZ2+gpjBo
6LDgT8FQzxXajeMhSqfCdLKsUImFiXkrivfMH6ZG+Xp405zTwLrzaH0qr558EiSA8dUdN3+zH+R2
uEcW2MNGN7a7LCv5r6CCrjku7Nom7FRyEPk7vPWAmhI8SB56D8h2jKkcIw9ImkbUi7hBXE4N39I9
oEZ2kq8ZNJ64UVjTSTWIB0dG1lYb08koOQKTrJs6JRlusDkCLhfdXzBh+VDvOtv5eGBZ40KWFO2M
bn9VkzoWI97Gc5/hIi9yGDY+2IR6+RIR23Jk4RDhLI+VBFYLMa53/By5738rL4OCN8ZJpRcuisUU
+RsW2+bect7421AZQbwSQCcOkydYN6LpybzsoykUY8v2Yo1321xgJVns2bfnDOz3PXe/K2JLAoU+
LLvTUfCXezicEnz7Tan5xarvHvT19h3PGVz7atpm347mIYnzjE8du/XlNU2H5Lxb8KEGOv0Xkcx8
0DOH42TAbTMxLOzi64FgCoFgRi3jv63Me1fyw+OuOHMDRDlEthGqZz3GNX8eTKyvto8AT9bB4W21
jFr/+be7KSHyGjnICNq8dPW9vAhgTLqKqiEYbx9IpsMVyKlAv/nTys5NcryO+FpNGL5qj1PxdoKo
CA8Q+jrf3b77t+jWy64IxXSzRBhn29e7xLr0bVXN3sU4EnNU13I0yMpO4b8mvdhVJ/Hw9Fv7Rz8Q
Llif3mdDxQM4VFOg6hG1QulLkANjqdA/vBYWDjftM/5Z/6WJIrgGOtVEP2QsXT8oS7sWjMq5sktX
ceGvInMGUe3NCA5N4dsLuS9fbTkdwoNrR+mQFNMGJMzhr+nI/c8ztrlJe89lBKwxhZF4PRaao/SI
yaTfrRc9w/Rp2pee9vODi9wYv94ttygPE/JmrcI8Qd/vyXkR5FU1f5woZqLbJbApiX2uWwscnVk9
uTzwPtsiNCjL7l3aEeTQIh+ICGDbTTJnGLOdI3fOe3RNNFJTFlwcQf2RS1RqUzJao/mzICSR94b7
3N0Q5/dhfbvRB/c7fhsxb5zZ/5ArqGWWe3gHrX7xR51Cte1JKIHgSqcLCtJkr5XF9A/pn0JUhWqU
BAqJ7RgoY8mDuzcpdMKqsoQ3HvDTuGoRCQ3oweilolApwwZeI7c57JS6viG7QLIaMM+WSQwvYUfg
6N+FoKPJibb1tLss92ejuJMUk7EUsgQhrVuf8GOLQkNnjKnsQYjKOVbzq48aI1v1r67tbDqbf83k
ouoCG0MKs4cjl0qitB92kE/l+0u2ChIiwyHZfe/Kmu7axSdSwlYfUHQxytmG7usQQlitAitic57f
Ykq1Nb+wMwOrkg9CfxkPcDY73GGDx3anC8vKHh81w6Qfu9HDTca5olaq/qsuRbhBrEld/fRndfLS
wgH0MCmKpLpoFUsxD3MbQkcainUe08OOfru+O4kyXOd/VfAxXy2EyOORhoDOpNPlZ2ZGxQqypTMZ
SOPOMndhl0X2vqUg+uK8GbCVD9eMuJPx9itdkBpuVOxMTolcuvr/WqgiTIMCJhENp1HecRvcmbza
BGrCU8diWIIp8OgxLlX3YMKhZLBFwuP3/88G6AozRBBdABRPYIkAu0wzaJsJHiMoKCzS4vpXJIwQ
b5ZDxzKuKsZ3rk2YK+Nnj5h+2rwsuJvh4sHS8/xRPmvpO0ynb8kMVr4Dsf7CPVMxVQ6zC8nlI4Qa
9WmqdFxn64w5givik3hhNHB0/hJ3182v8NRp3/ID/YegbuAdIg68A7vlzINdLCjIfEIxl/syEDcS
3dTr7G3CbT3lMGemEzzF+crcYG7HSXE7lo/rWE7JlScCZmABQL8ueKCxitSbAIH+TTBNOkD6qgyd
Ypms7CDWwopYy5sqLSt6VDlq3dUUa3SsaMq2dDA/QEWnxtPzfm0yL8bx0Vgn2VlZKoCFSE7Pn0Xq
ndTR9J/Ka6yWfdRQSbiIhm9TsA+UPYNvoj8/l4o5Qq0Albb+ou0QV7/zWteT4l+Un8gcyWiA/PBD
zenr73AEJQfqs/bxHWKBqBm2Jpld5B9E9JadHIShuYlYuAMnM4D61tQyEksC3yso8MzYNcns7bgh
4dqmQSZDBUOLe2XV1lSCOBuUzID4/yMG4WeJ+HSV14TOk4ZRCwotzx+OsLGUNGHSZ6aYcilW7lJX
eVNHeEojrPTZ1XStabgY5zjm1vKpQNBG+7nLW5QJHnD1619jBLseJ0r/V+3zNp5baVUVa9PTVE7i
lsN/DxCHIjelO9gFK2W8Li2E2Q6QZo0b/47kshBKxPVWLuhLpctxmJ8zIWDTAgizkDGb3YTzbmVP
SqNA1DD4NvuPHZL8fAtpiK5S0UovSEd1wWp5yjh0OQvg4VwX+VHvvGuEWTkGyljDG56C9U8cra90
FCybkp8805NjXPSwKmetfnF+k5Ua5oCVV/dtpJCOUrVaBEcwUpH2eBUOXkuLgTW1EJrxkzMFKtvX
rlrI+u+ZWCvn4ACr74xpuy4juYAAydK546L5yaKtr7V/LpiyyYLV05O1ITzd0HlZA6goD403BtOv
iHvYQWm3PfriF8FfqJDfsUobeMkjKFpxrc5LYF50mlT4/OS1ezMrOqyftjohlp3SBg1gqR5g5uwX
1Lg8zwHt1Jla9RS4NTUIwcridAq4dIm+rDZZcSFbgg1MwJp9M9jZJsGTivqCns7WKYKm9bdp36N/
LhkPVOeH0FNJUl0rCKVtxHRswARlUdBRNm1AZycXxhTXb1VVy5ksGNkfin4S9eFLmYCFkXbxFS++
60o0KeH2ojp9F6bk4mXVyw5vGq3R6oT2rq7Y4QnJV7MtWH/2rIBwaGReXPjA6dwBAgx7agj7xvIh
SL02qa5Pcv7eUskMEXjam9ykvH6gG8RRIJxlhDeFbO6HdJlcjlWp2UmLW3bObzTMgPSwD4N1B8yz
HV25Q3f3z1Kor3mKC4t+6B8JPxxTWB885falwOU3Dw4hJs8HSIejcPUNAALKb7QEAn8Zbb4MuYLt
UnaoWbc/xjYV5i/35SBTtk+xPoPBzbCFW2xaRwBEzz3ij8DjtDBqjboOjPmtMgCXdBwpg6Dlm7Ox
j50wn9325oZuVZJF5izwLrqrTWT3IbAxkmZELc344pFcJ01BhS/13o/YlDMN5njSMSV5BD2qcy2O
4atlC8ZWbabid4Lk69BQGxrPiUuDkvvS2wt1kMgKGkdpgrBR+4hzjJpCTnB3Wi7+C+VFjAwcD95O
WR+qotAnaDdo6JG8cOrBvGHFMZh5wrtkR3VhpZM7wGGPC37ZgXzqtlKDzaxdOuo4pBrhNPF9O4Zu
Ec/I+LkG0kOi/LchVuYLMlJYfrtIn6y68oC0VPH+dzZ++dI6NqNkoeC7jXCvR4zsCVTEa4DAkIct
WmljvmN9XSO6wMXvVCHO5oItPuOK4acP1jrRrGX58F9pMNp2gYj7p4uEofOvr2JkH0FjUAI0LNh7
vjpYsFhFugg4mh478zokJsq2ujJPNyomuWPn4lAvPYb9+gzQDeuTmzptbHDSPhuwexCK6wXgRPG+
AVXkBE3jXrMXUH7Nirbsk7nd99hELzgC+FfuC1yI+U1XgMEHQrur+PpP9FKNpPGG/3uin57s/hXi
MZ23HwlCoKrM82Td0oZZhuRS1hQpb1kc4gDuWQGhPaUuRHQgY+kEgDOQ9tfiMpzXBIcmvrxEKqqC
5kenAVCmPMipCFb097arFT0y7syUWBIPa0WPETkn+7wD/wNGjoSiQ+5GHlMQHwECC4E0VdfdlHeB
WZrLBAnpJeSy8Cvd7gJLrj84JesbQzxoDawtGBLwif4JRe2V9tTJkCQDCDR41/ebGPmfRm547iTk
ivRdtfuto2NhWBpqBkgjNaT1PSTdrXS2SZmh8twt3eXwu970QpVhlt6cUkMKLwo7usupDB1sOdcm
kV+3UB6/7cB5UoaBskokAjumudiPO4AR2jXUVicZQax2GzW//aeH0pFT3D4rxf1Bas+A9GpB5LCH
ROhAr3UDvnDZyh8LPr/c1bizvNeAxtPlL0GH0zaQUjP+CketzWLS/oX/3B70uzW+oQsPVngYGY2E
j2murKIRA/Dqauv9WrG+EHB50G23aVuVbENNOGz3+v3R2u8xY89PiZPK+fGrHkn31j8lrIaXY32p
fxDeAZmbWPXW4hYILSI4tV0Pkig+oR2vRljlhCLNC9RNLZNJHX7Gde45V7A3rOLMCN1htZntaKox
VAiZU0gJdsXi9EdqwGxl9KHA+tL5RPReDrcqypaKa8bdYwSUp5lCRt3jAKi92t9gU9nrKeQnQ1QN
T88sxucKFFrhuxNMnGMYKU/gTiGEvoWLJMhfs1BdUMfgrOld8R4Cf9MxbLT/+t+U70H33/aND2vg
zxvD/3vAHxeomzFVLlBFWGp1z23wyrX5Rng7X9MNdCITtBS5389oXXoVC+C6C7jA12M/+7V0JTIN
9IGHdLC1ljC2N7IPzfY7Kt93IqhXfjGIS0NlLdsEc3MJy7i0r2Icin4307+76dRRu9atUh2cwrEV
22NqGTqby7ahQs2JKHS2QrGtjqs63R12k2SKswMfGd1+NykpIMNSqQrW85z1lhHoiH46BUOB/TX0
Bx2HbO+YgtsEzW6kCRHboBYIVJ8aG5cutJbpnzbPswVxWDF0y9vZ4tqOnBoXO73Kl0nlqMKUZMT1
dOi2IhadEqt5rq0FRetx5fAm74B2g7JHNKafiFj50042s1nQ4oBqCNbxOKkA30xAtDIhU/IM9Dde
Kt3CKMQY1aim8Hxew8ziBaPSCeKuNTHIJALywdwKZtJuEVff8FyZvRp4BfkQmLJRzqOlJ80FFU9b
B1CsoN+JSoV3xfjRQrUfEXiWc5BDz6QO36lkg5PTavLGhytMaFBXY65ItEvkADx91gGzkm8hSpyl
bScnwZ+mM2f/oQ/XoyrelreBumVamJXwKwTVGAdHj91D8x3VZ4FqTlDdayFm+bVFbwL/zPhMyecJ
qCZip+0A2JyZifrB6bQyZhgIF5u2wECsD53t7itbDgf6q+EnDpKqW6oPp4Gm5Ebq9/iPwTXrLrTw
73HWtpWn2GBI4+jynRZoqmGC1chWwD83seazYagBZ/mvCDcr0Iul1+QjI9AyzV8Dgz+O03z7ViuE
nZ9/t/HjaZYqxQWsbH9rb6BjCw7CY72tPkk8imPNCk5xKMPMZkT6CqmrLeNK2V4EwCZzGCAUHGRW
qDsb0ZHFEE6ntZ1GNtDnbbCVlAp2dDEKtMNTngNsDEdnkriEKrJe4JQdJGNEjiD3CkgQQmK1nMlv
iviTn/MRA8aHY7DSh7VCyDP4MXqskrEQSHVMdGwVX+pxH9HQyGZ6Kormqg9PEIburft8dLAHfnot
IK+n9F75nE/a/zR9q3Wr8Kw4v7qIBFBRm5kPkmLk1QXYqIOfOHaXzjQUpMCWZ45BDgN+izzC0riK
75NuYPlG26a+sovanaKVNkzfaoxiruFqEIbGolW4tZ/MvZ//K6A8XkhzivPFHXDRcfCBA3u1Norw
x9Fk41jt5s7pRRr5CnOHj7wRS6oYbpaN9KTANJ/HTU1oEBke03QFfcPAWpZEub1dq2Y22h0DklR+
+E5AkkOj95q44ZPclTCy9vAnmbwX/d32hx5N0Is7jEVqlrpz2I9oLqT/TRAhgA0BqTclfcjirYGR
E+vW99GJ2WL+eA0Y+MJyGng1hI1/qDYsC2XxGpFYa9Qy3lAPArVWfa8O0NZJ5MXIlpIno1ZrGCzK
MEl9TpFxdSSr3je5L28gD3efXcivNNQHTkNepHhJoxnhs3VT9HJjy7QhfwAO/aih4T8enU9oYygj
LEsLSXyKHzu7CU6lVY6SOXGwdbdlv4AqGUOUFzwwoif2PU6hdLD/wqSZMZLRMQT1rJz7JU9BcZ0p
/YN9rCn6AGgfAcIx5X4YzWTPFgQpqn8FWv6DkGdw0a1UcS9xftWz7xfYaE5ffUaeIHeUhMgLv+1V
vn4RX/z0je6aMDJLfJ8VJc0hekiQjgt4k5jYGkAp66YhIz2rK09ySbvgb9b87g6Qb7TdaT2MeKY4
LfnN13fQWtCtOIYkPExb4Hjm2ZTYBUT4P1RJs9OJrbVqTEWVV4tzWnBYRJow9u7iAKeQX9Mtz3XT
C2k6060WP1Q9ZWue1bYBXYNHcfzDY0/F8uZisS71IiUo/XmKmxLk4O+j0sy1mVv1N6nNy/U8Z4EP
mFuQNmTdKmVlym4082cK6GXvU0p7PMYEYaWUPh1Sy5H0gCheBgNt8cYqob3z9UGO3TQFz6G63Sit
If5ytgpUdUgHlK9w7kCrUnzYgKcHF8lGhMdShg5jH/dkS55BMgzeNrqDE06h0vh/i0oDgB1AVlrW
UuO/J2amB88YSjg/w+40B9fD09k/T6ZGE9KLf8gqy9JjXv150NGCMvp9vkoESHoh4oOV0vltwZ19
0DAghPASH9IqL358z49x4CMfTSFG/l/4fypg/qdxZ9HkOEKsae1F8z3SFxLHLfliAJz/eKZH9seO
LNnQ1Poi7sdb9KogT5mhrTUXqUxvYfh3dRDeGhgp1nvcqVjHQRhI9+KiVqQVHZT5XVJjpDBATiiP
dHhtD2k3CGpAD2HKLTH+AXl/1/VVIDC+HGdZtUhleKKrdTcwTXy+2OujMIzvRPGsZEibYHoSCiQd
LLczO0U9b2Tzi9C4fgVDLpWcWPCJMeV7UPd4vB75AhueXYm3a5M5VFuZITU1I2oQb5Kmw2itIqG/
Z/E2lDDHF7umtt2CFsR4/B8SYhy/J8zv1jguSXuDzYrfOP5U5YFUtrBBtfHJOBBYZp+ZcYOq4PxG
79Cf1TmCwknZteoq/0iKfcUyA3rR0IilIOhgarg/Kt1WEnqY8RfR0GFABbjOA9cXrwMcdacWXoUS
S3SJFxvAn9IlsMM2kj8rQzIQ65pccxI7J20eJS39SE06NEb9eUaI6NRWM4BTpId+/ndL4eBIj22j
GeEKFPYMoYMVBe23Pi+i01lVWwHcVbUC1GvqwLlkkSVj8K6XJFz0484akJY8dhpeVkl44Kx5fsk8
FYrtlCKJwu0qwEtE6LX5uYQeFNKojdjr8c8THcmSAIfFcYrkeh564BAAmAiQuL93xLIWm0Y23JKm
zxclzW2FkpJtX8gQ77Jn8p/n8eWgw7OQdgY3SqyXicU8RCdXXl33wYyiOmKAzQ1xb1owhRdnWC48
ffUpT7oZravqIxHTkPkASkazSmRkRjO6U/95UjSXnElebNNpwKtjYhq/NX0cgQi8SEZHfky2xdqH
1d9oR4KuYGrEIyuC+zBwoCt3bfMGQEnbucw8N2tef+l7cCKy5fVloLmoAZa5+EE0xYhUPXwDLwr1
9xggcOt3jlRE57MDRzaQUhFJ05R3Pap5FH8e1SXvDVBmREx+FAdzE8odXBXvnjPu3xnH9MCcdMEF
fceZAKslbwtvt78w07/T7uCBA31gXBJczzU7pLBuBmtnHBdPkPEVTvaA6ZQfayIwJU9gM9iWuCIA
fmaCRj3n74f/7JTbN1ws6RWGmlEvwDS5OcJOh4hGlHSp0+SjP6wU1UKuqAbLhSa1zVoHC6IgmPUY
cbUYKPisqE2CFrrtnclDmxmXqfTURPqC4EdhljSiaqdez3iwhhNfrlmP1Jnph468To3ppwDrzDnh
L0ZvVKx6Mj2PVK6Lk7Xm0rx1RSaJP63+d5Pko931aoDPOCTWXgHbbKC6X9ECqdtiH+W2OqDjXipH
CfeHdgNXxtk8XNTqYPG3XBZGjbrLmxxZ/uSnVQYRJswn353EvIGVSbUG1N9GGhWsS+9InHQDhkBK
/VYtVJ5U1q8R/Wd/aopgTNG7pT6dy13YT80pOxKwegWrr/SidOQCyVUEoEKvAowSw7YjZEU13Yhg
hpAsWlxGUhraF6PWGgljxU9yjmf9FBS+41V3BS8uDt2o9NK1QjYB2rw8fO6/csdgWraKvDg3kXtL
izqsSIqSr4Jke9NrT6qgjBRiIvgs+pzXZO5Fu6+NpqWEbIXqYD7ZradHF8y5qJbjQsTZdTkch9C1
PuOiG7bN+6WpBiRY0MdNRE+mu1J11OeF/k9xzda+IcFD63LdBFiOXH651i3jo1yFqHpa0K1WLoMQ
T8ubWt6FxUfJmM/jcc3vf7mwH3RJnfOvDwc44clASHN7hXcQXw8UJItwp61OLtacBdaTt5aJFWQV
AxMoEseSuWqEFTV0dsQpmE+evigNvkmlWQPEHbLIb0NnFiGXoKt3CfMjTV1UDApfbFnGa12dS/Ek
XBENtx9wvIxKsevKhurEEgCxQGJfWu60rerN79OSFOFvui0erdeSEG0e3IOZmqPCKIw+NC4aW3cX
ePSjUb8z1SXUjxwvFEsq0lpczd1qmEX9JCBNdKCitA3lZiMzPmjPVL52E8JYc5p/l7KbtEvspg5f
7Kx2pSbIylbqxeZhEZKky45BdhvADJJDNIcEGPE+gEs9g+Hl3RSMepFju8DAVJBrohFowMuF7T2v
J5ESVPdzgEDgW9oyT2bP5cTJ+ugakmg+pJR5f5eNnl+sJdhjMo1WtCysPQnU293tKAsx1YLbmnUg
Y0Mt8dhj1/jjr5grnvMRJupuF8jdmDqdLluPShrfCHrVryEX9jTp1nH11G5AoQtgrIyBk870Y8+Z
n335j0vt7C0p5cH6czw+BSY4osqvrL5JPQVLpTNawS4YbxoDEZdcIirwgLiYj5scNGm8o9/zP5ME
fb5r0Y8lDVEoJsn4QgRF1qrYsL79qrkb5xvubKTgEfDEJ3NKBU/rfpMjhHeXqMSlewEs2caoWzeC
HTRwHOOi4VMaEnWqI/LtXc+4rsHkJrPoRE9pgVjZCw9rai1WLZRJWZj1aAfvqGvKadFxAnljmN7v
iHFhxdIgpwmL4mwH+hIZjXHfv4vDjS5LSHYml94loJy9C/Q/AwP9pZ/nd+IAa+buyYuh3V149v4I
FYbRhPbL6+8wEnOaFLMrzyoNwlLtaJAyHiwMgGxwBDafNzjAgyJd5WZEkt0vI09GxlsNYiSiozCG
4GBmGd6uIn2PlYO1VH1VMouXeocy+DG5nnEew+5nOuhdWrRJ2mzn5W4ZVCP3bXIghN9nUek0/n1D
Jqnik/SMrSMm0mDBLLMjbDRODYanSQfYlKZiAkJI/4oBhPLP8YonbW5IdISaANVJgUdrvplnLCca
t06GO1687+l+AAu+jmhlk8KA8eRxm7igOhU37l+u0DYHoy4dTADGa3ONvVoN9OKMkWyeebkUCY6T
GJ6C0SMMJZdF6AWC5iv+QMbHxIhRH2dNo5DnDSJkO/eDc5rEiiZ9ZXCwoRxPipvEvOBYJPtRTGCh
jEF+fiXUq/Qir6ypbhAsjydFVfXzb2USihGfVbBLZJKQ7ZbEHvi7+92f2NjzpiE9Gun0kDvbAlfW
806UhzsEsmVcd/WS+Sp0W/R37UayBdGSakUeHlxV55T3fKX88mx+MTqgKUrbKTuCLPdayLth0oRl
HJtxwIwHO0aSfUyakhOJj0sPKM31oixiFTvM++HYq7uAEnvGpkqQOmHcXs15+8yeuDC9KEpvCrJn
iopIrcUtUlp9pfHqRxtB3KiWHYE0rignLZon+8WO0Sh4lcvJPpPAIBATNXJe669GGX42e//PVof9
YWHa68B3nqHvn8eGpdLUBbqYrCgNsg4a4MtxrWlVXg1kcKLZw/jisjQBDPOqB2KgfTJiC2ov51Un
vzx8yBortgMkUiL8XeasLpZI8mbumxedAcXZcEUUgZglPcSMlVSQOOgKv44DaYwOmYspma41KMuO
p9hbXKsgRvtODQLkRqTO6XnXpVsxxSA70kI/5WOOJaWXdPczFK94Vm8MZfpISfmuybDLYCC+Trtk
lAHHtpQ9PoC2VxKlKyp2qMI+9UMXgXwQQHNssQKj3UWoWhkF54zPMYrJPHuU9YaDD4LCKrmkWxQX
plRikdGct1ApBNnyhEY7Uh1TPjuzJnqFrSWlWqSYvfnxdCwy1UgF0XLH/jHvixUE3CytWe0NZPui
X5Uh8HgEhDt6gw5u0E4OXriSBowIR0j1Si/r8omCPj9sdpwxGP+zZnQmbJ+ja5deooplTkR8mebI
K0Ttr500mxh/Aus0iSN+wcOv+QQurDuzZtgz7nwQ7T+ADlmqMmgrkGsDQZkZ34DXxDCsrnMtPyOm
6VDsRmWvdHsZl2Jqci40WOOylqV9maRHRu1LjUgwIhbPP/7Nacp/j7MplbqBeYvrfyN1XuqvrG54
Kx3AZaBRvf4AX4cGq09fXEyy35ejxjHlr/ZiNE3Qh2FvjDei9AJJLAVOofSueFGbjTBNchTMM261
PDYP+owyK8XNpPJ+TsJST0ZxLVwn2V8SjpS4w9jMKkLngr09s77iPophQgf7T8frjqyAp5oO7QZd
5tH7916MXp44lMXl6XJB0FrN7uh6AbcvXZ0CSEan7UDcBEmGDGIKH61l0Az/kek4zoTWLr0cjN/K
CtnHlqE59ewq4Yck8h8G8IhslbVTEk31bv3Urfg7q6jCM1/RSEtTzWBQaFIhAqGZJXPufzETcXcD
WjSdYnxqRrfQkY1uWrUfQgfvAWlUbNzCUNBviNM92xO2DhzJ+cy1iEJV8R4Jla2oKp5YMSKzZUgU
0tRfyZ/lAjN8tM28zRqPhjqrk0AJZteHeSF0vz8dq17TMU6DV/rKUg45wo10r/bsoHBZwdLIqQWH
qHdOIZEZWvj8NfvKT94Ne/DQt8ggv3YrBVBe9598am23Ai+s9HHY5F3WpuPwfC/zYxvSYoJnrqA5
Y/Lp7qf4LMuReFiUj8JVRZLq4/SBYxz58NnprfO2AakyfjRsdvitrTpudwpkE7MP3aqWOFmsKPzZ
j8bS1CBVvF7FIa+Y5NntATM61a/CERF3dAZwJpZAO/V9JOM4NUkkMi2EqLHFm3lD+YvCyKkegNca
Gc1PMJSNg71kPL3DLVlHqsm1JlCAkLKcT4vftAwEjS5PAR27O3wfkhkOO46ZNo91h4g/6/hevtyB
YXETROiVg58Im45kEWJz9xu12zNNP+WwnIiqpBpnPBcrie8mzjJetDaxkjB0DFVr0maa+n6xYMPM
ExW8noT4rDughUEew2bzfuYwkfIN20jlLkqRgMPuHdACTm+pIbcQ1s8c/21bLTRgEhsSOF8RKRpH
oc/CCsvF/SmTusf2R5mk4UPuLR5BYGjvVgiwGUcF7QB2/+YgTgOpnNqd7mG8R/C6/+vHORbKpo8P
Zfsgq2vTY6boaJvbb1CmQju4brZUSDY0X23Jfqpqpu1TDfkML5pC6WpLNQPJAg/Vtk+A9edATngz
c+xWwMe0hJqwn+NaJ9WoAS/IGeF66onFrGdcJd7rtL8PKdP5sf6RWO2siQHczhqNMoMuuWjsNTW/
SSPsmvCnTV0SjM71XM6oJ1ALJ+LhKbLdovxMWBkVvg5+FIMmReKWhBrGCTrkfxS0DheccPMd/QrS
Q9tWwN3/OCpUWWu/02qXXwA3rDqF0RLQVbL5/f5GSNMZW7LqTAHyWgAFv1h9xhDrDvtX/deixdMX
06TA7S9exNkKjV1AZpGFTybMIpO2OP7g//6350xzm2fS3kfC7aokY+lfcEm1+bysN7VXyH0jiOOz
effNZDNvfEBWZZLZ8blDaQoobS73QiCfEpm7tCiWrp+iDYmqZHoiFphNsNwSdL9G/4rWpxgXfRyx
KLE2HO7MODxjls/ewPEUk35GOW1/6HTwwXKoMoTMLX/YB3Ff558FGE3S96dzXZaE1wn08jwyFiuN
KVAdHJNH7X+Vp5W/4BWu+po+UWOuskq+Qx5OfL8QelFurZE6nK5kYx5kD5+5h3FtlszQFSrOI6iw
yPS8OGXSaA+f6tnITLgtiHZjqk2XziMLXgilwHlGlPbwDs0b6VRKZ07LRSGQ52xn7o2SWqqW6BtA
Q+2EtbiRJNT+1TqunFh33DCRID5tOVMyVSDqfcaV+Ts4JIZvEJyqz2KVZJxrhoE7KVbjR0hhfX4Z
X8WUiYix7zgT6B7aB590pBkSFA9mNp4yfoCBb/ubyz2x8lxYEWuy4fFZ3sWppIuF8e9hbs9/Ttwu
8h26JOP1rqdnQMK81hEBIS+Xj8flv9iRKWSv7dokL9RUPLMJqR2OryHvHXn0k8oRe1Oj/8fBYFau
j4f2SduSJ42vHeODCmuBDtGs3NzADYwyHMDccgoU6gwhn07kgkhDdMAf2CafPOKEV1IJ8wvFhuQV
XW63bW/ao9B9lFJaJnhr4hsfYl4Qrlva1N9/Ll+zRRUnxEz2nNr96IIVXm95aREMUBfUd9mFE0bU
9e6/3TShbS8R4Z3KeT302KYEFvhMl9xi1dNoJNW4rLjimZkPwXMy78SGqTkKadDtBFH21j0P9SKU
gnCowbfQwaKhWU2WeJux4Fs73BKDIDxUVRLga7PpH0wT9WvuO6651RIDSa2GVH2rxH3vQx+uNZzc
BIM09IXw6DlqrVwcZ8TVjnFRUdyaCsX75gCscd7+e3MKbebcZRqdYuSFRn7OCrDMF63FG2M00Z+E
78GOzb8EVMJ68umfqmhPEaFPe304UGAFR97R7eyGOYzZJRAwna8ExLe/iYDVwyD+B6quwGwh9g81
6TjB31IHWG5s7C7KFjEPT5rQCwhQIZTO/5sPQm4/Qc/snReHPD1xIA+TY+DJ2JHOd9uM/WeA9Qx9
GsrumWanBAIrrrL6C69VL/MKrpzU+lYA7ZXWY53W6gTb7tMswBsGBPbi5ZfWTE+W9jFgb/J4q/jG
v6NwldC3bibGHd01hz0cbl1W0Pz80bAqjjU05y4Jc48+vE0oJjIcfo0CNNm3P/4l1SF4lrlPQljF
QLW/rRdDOyCPV7CAWebiQB6vPIqGWpW85CkFJs6ShWbgCcLsP4UT5eMa1MWZdtTcLCFZF5Dh8LJ1
qxnmmL3CEsXut0wkAKD6Jhxv3Lb3OZ/Xgr/JDOtCaOYaZ2/NIEDVIpIHt9gqUkJFHp4fvdHMKJ0u
vVMC6L+wcaYW6+xx/XMMqz+ADJkTgD5uLWQTgCHKfuudI9UUtFvwrNj+yFaownq60vn/IrYx94mL
OhozuQmWm0txhGAnLV41jxm7Smp+8busem3R8DWvibD15Sact+j8dPCLr933ALN7U8GmjJqgBX1e
NW0vsObqSamqv6TpCbXDawG/KPr9gk1kru+YKdxOe2kdOH6932PTPEKgCHfLg37IHRoSeRqZL615
WjzZKaPzck6ElgqwseoChdagrAIUZAyu0QuRC1tS22RCIZ3vvtjqrowZFzf2X6fhOibIaMSdn4OD
2XkCzjjB0GKFqLLNcUNvNd+fJaWk8QU2+MByVZAH3xTj328ehhGfFPbzMuvKVEM6cXJccY3VXuyn
yIHJWf4zOZKD5RvYWspZ9Bh96dSYiDnCpPKeeajVG9hAHZaBxqGjqvhXtLgHSg9TY1+kMjEu6zhb
6Vol3cBzvCyhhfhvtZrc0jjqXw+9XuMkFv+RQlNYXrGUCdjlmlSU4cfcZhd5US5PFII1qr9HCerI
FOguDfOjtA4BVWEsOZqF9bGUIn8p4uYb01kr4eybcSewUj1VebMLwc62u0zWKpfzaujkx+9GRzkb
sXxZNoenXCa+Kz2w/4OTGjhmT9wDML88ItVaNygm8ba07fhEPe68JSRtgWV2mQnqqfP17Lqi4dFG
FHNvYeDPT6MQylgpIrOoBbCjp4RQFdfojhF/jH8bcyvuAzO5Xjr+p1Y8TqHoGwvXTtGpJBL9x0e6
j4rngIYwkc3jL2XpJ/k39udkOTZ9SIIbkBHqhXsH13HGzPEa97k7EQtM++VKIXGsgeey0kY1QFRw
LsMFNCFh5G24ROdW1nj1qC39OLaGQeTrIUmVbh7zn5CmijMIHs126SDyk/7/tfuxn60TLabWCWXv
TBn+12lcTb1Y2hFeOCCNpUsI7nQBDegc/KQwhdGT658Q0or73f6XVzUnnSSjHAq/XjRElFxpTjM1
VySC/QMrF47gF0NiGGQ/FSLjyShETlg9jMY0h+9xJj+af1PldfA8j/kdIPXh3Y56U/bxzZ/GYV2o
75uxILBHqkTaL6ZV42MDk8Czr/Mp9DkHXsbr0ymK3SKbRuPaeH+6yLAcbT+xQXdW//oHq1xyZGnT
Ki1nzqMkZvmuJ4YwL6Lub/3b6w16bgYkqhEmImuzDxcidHBtHkZ1DJkLQ8xIFNZHOJVDwNIulWXY
kSOAg4RBRXmG80Gg2AqFaomy32GaqlJm1qPcCLw2rzRs1KNdJ37l2JSkjPG1GtPktc2UJdo7hqc8
16lvaEMXi4rtYQxrJJqeSETrapaVZlW5e4OxWtr/3QwH5Ec40HrIthitU/4YSZ8Nth7RoMmKDbm0
ZjqpuS0BQy9kg1UNY3maLby8YzAorWd4ddXSK3GmuNlbnl6+xpeeqk4/3zN+XpPyj+tkwbGmae/z
aZd/MUgMPlduC5EWDKK7oSqmSauUdS/lTHLH+jjkiguGNhsUaW4SrJGanVWFlcJve1PSMMJsflh4
1tgA+tw6FHsj3yt+Bb2uwAs2W9U9i4u4goLXsamCb8myXcBT74UO0M6n5t6mKT31smiQDk8iy6rg
IYuzTMRTJHNc2ac4dOHX45YG06vXbozKMpGOe3GZxvhhii2IsfcL6Hhjaz8OmQDAARV9hrHBE79T
Xt2d4OwFjZlrCgVvcCSSHErhscbHhe+mFMLTcGqWTnViFuvLjNOlxHi1gAOd2xyC8u8zUovtWsan
mfxq89xAYqAqI1W8xR68nHMb1sIjvzOh92GQt2uw3jUQz+H4zrccvXXgY6sU7W8u90+QtUSIlG6O
lLuL0bXAP4VyCnPVI6n5aOhF93LmPFcvpogES3MUnZGx3mZNIdPmX7cAlHoEh/b94BB7b5dUkYO5
lY4sVARKr+eilKZ1yAf+iTjAwoHP48UnTiO3qbTp/TDVIelE0tsZ8oGLBCJSK2yQSSwRB+ErYl7n
Ta2Zw45NNhikTwy97HNCSVAExuwIuIr8DFuhMxBVfyLflVKIilZH8t2nZBuj7cwdvbNgooERzb9f
1i41zQm1FjGhPdYAgGJYfOqZSSlIJgl9VS4AYGC4WqE6/QHED3cHBfZeoiSB/hJz6CCFPwEzY1qh
Ge4xcjP9CXvpYAksEuEIJf0FT+We6kzjFlQ5F/3dq71hJJCIDVJ0TQ0syhMoeQ1Fvxycibu22ae6
uqMSGX42e0DPkOJ+LeEet884xgsWVWfDM8imR09xSnaaDJzhYFbufE+R5+9fuxdSeJPrK5HdhCXo
DML6YCj00TDyUr8w6ezAZwusWlaU9CAqd/td/rD9SX3Uilp5Te0IvlDg+Qo9EHA1ulVUx7AxkGII
dacjw37/geeR2OAUdSx1fBZSaKzkFIgMdXDnlUX6k38Qn7tXxMVKyV0caWNXSF5A/jPn8dA4/jMw
iNTwflf5W4fv0qCMCOJcI3HeKEp2ta1x1DJ2C+Vpu7vjMP4eZA5ohSGutGgCyof5tZqcxIIV+j2T
nHmZsTr+FGMqqqCtfGn/E4r6Kw2UQD5gkCrx1Jg+63yHYmpNqrTgbLdu+FusdjlhA5u/L/HKw3MV
BJkOQhJHM/no658s3orAn7/z/vfoouuhYUV5Udpzc2eDcVtSYQpIpya+VV+ZV4xpHmCZuxAtCm3C
AJLWeSl/p/23Oxrb5egblA2rx31pmWqmnjf3ciAxcISdbr2HowXxST/1/xFoNYw41hVPG4cE8nIT
9v0qvLSa4vpgXG3ppNMWbQ0tOm0TvvI0lpup5tYXWjkmKvTOauZXvlD0V8MjshN2pNOFqoLVftw5
yP8a1W4OzsEhdNUF6Q/nYpbeeUU8t7No77iB85wArZMYZSzI02P4wCIAhSiGwe5pUlGTUgXMcVQI
eTvFSBaQy6nE1Gn7BQeu/AD0G5C6anKjwEj1Oy9/0a8jLCquhsBojkEXXEd9o1DVL43J528HgNOJ
BVcyYx9sww5OYTIlp0XutAEHg4x3xeFJejn13depXp0xZjlD+aryc6DBgp7gRlP3JI16s8NjAl6h
SrNNJLL+EXb1EroruboQhWxqkmY5DikS/1Dzevsk1GOJ8+MWo6kk9z5a1Fxj0rlZy9CCM3nWJ6d2
8ZxUdDVbBLVQJnCK0GFZe/sXPPnYvrYnsmUjfh6KUx1t+swseBlI+Fpu/Y/gSSK4rgEkzTHx7LHT
fmTsu9nT+dGmqYrwlkBcsb2tgGe52tlVVFgHN2XBz0AljSTZkY9Lgxtr2ORbYNIm3aslVyZP9UZJ
2jLGhJ5vNSsvLwWrAReXTs3MAwLoTy8Jiw6xwSRADxSGdqzmDsd3Uzr5jLc8jqUwFG/wX0/GtrCU
n5McmDZFfb70hAeTUzy2NAPod+x9yuq3JvEeB4T/0zmjOhinCik2soE8y9KR1rWo5Uvr8NCEUmg7
KiRSo6JXny7Tc5Xk3QzbUQr215qIBdoPIZ9cvF+VgKW7mg4ZqpvmMO/mx8VwUdVedt7POT6g0t6I
+u9gylfmNPZlLxgToGfXpeQs/8Fc09RdnX6o2ycPk3bsY9aFWI8Y3lmubAgStn/HnaFO7JGSwP88
Z7G2CWWnEFv7Eniw8Hq7Vu1q/SOLv0OT+1DDKDzssiORHPNUF224Xggp426oHdBhWz4Hsvd9IbHg
RJ3PTWuRrbyTW2XtSfBKoLy8q6YK9xujjTEzsa/90vj5E5G0RGwBf8uXr8m6pftp68rnWOTAyQk8
crKZJk12A5M1ECwnMApYEw4/eN0MLtq5iwEeNrGVVoj+KDf4kK37/X6cUFFNDbSoeC5EiQYqCJ51
/WekOpIrX+Jx6f/Qbklb59fD5tiBynOyb/QFxhTB65moZiPDKoe1Gs+Ai5hUpq7zHGk2gIwp3Tpc
VQKVw90ampqF51/lff4jnZIRi+3/3ftAQdtN6F5K0d+tEnoRrZcAEh4KqUn9vHMMUeKhqeBBmlRn
er6/T8nuYI+SONFsuyqjAQKTPd7RPTKSqFCoBkuK2c+VEntSoWeYIhirwyfz9rkX/ozT9D8V6bj2
FF+F1b0zTHCwaMD/U50rhdcJYEfMAKrcuX7fY3cgnL3aeQegoW5OBSAjZdydU2XegY37cdB8Nxol
6nAXa2HWF8KDI4zixZMv2Eluwx8ou6fQTe1wtvXQMMzEtbTHMsdwQVoUfsQVg2ffwJMIzalrts31
7i/YkdxNEba4v0xvwNp9zWWNBuLVWDl8QPXDLWro7NMMSYmpHaw25A6bLFuw10W1LxJfNLcIQIDI
ygMBhsTB/hMlulsFgyHFgnzCQYohVAK0a6Vgugau4+lX5T1KjXNGUgSihOD31wAI3ej/wvOzEFXM
ExSz344jIyBnvcsgT80lg9U8GtgNgHR/kwv7jn/h1OCsLhhk4anQhaXxb40720jMDqPgKqYEaAlf
sUByx8huEqTj3DMxGNv3kgw1s/TThgcBn9JRETwop4/6pttsAVM0xHjm9cpEVAmScM0JbgX+z5lL
y/07sTPBdhC+zIZNHUjLuQKJ1scGqwrXzjflFLHJG9upgmVEOCVjzBK9PQvako6ovK7LwQbsiGOC
I0ItTza273bJP8OT68Hcq0Pl4XnA2lN5x31ZZ7x5fzzS1EUdXQZLHARlbiCJ1lwjJ91VTiTlJ1b6
ENDMw+KFWiRDlSE9Nb0huPs8aVtwkErDPX6XpHaeVXcT1itjdAjBu08hEkbEu8faFb9ljZhRZpio
X9oszr+zreFnsGnT099ptsE4Wk9vrRIneiz2j0Jwf85P8/S0lBpO5vzbWrXdryN/mNigmsixMqG+
7Cw35rdfxenA+ZAcUrvuvGKuDao02lo7s+8WJnGOQHgnD3f9s9MWM3OIzj+wmPHjLJQ9ynSslKDJ
4wT1w8urvLA62kh3s4YNrj/JQL7mGq28snEyEzJsUW/OKo9x2xQWdhDUDpQ5OtrB4jSsuFaYWFcm
SHzhQm+jjT7AFcHNLNLjLaTx+4EWyQL2QA1anBD6znZ5axzu1LNH1WQ2J/fpPYFpBQ3ptejISIIb
32mrEk1jdTfLkJXLVR09toK2HIXFOyTFp9v0sHe7y59KQXwkxUmU4aE10R7fm5+ZhhZKSwpPru1M
PXd54dDA9gPsYHy+ZwRXCLUk9fi+wPynLgrvRPbYHJ4WZ8PpBAQKCxwMnQEPwkA2OTaZih4wZA+c
lIkp2refFpItYT82EXJO7QjTq2z3wbtt0FTXQhssNsfCcpn4+pQEfo3fVtwT7fgdyDEO6HbQt16D
NlOuKxRYR39nSUSkUEdfJ1hSxnnf/X8Nw/O489X2fG5yoGNNUbVve0CmHZxUXAAwaadL7ygjcJAz
kUzry2oZMCZSz2Qg+/k/kNPPQra9GZYRPxwtP+nM5qVq6rPGKQsvHp6nJUvyhUJvUsiJCb0tKg0M
wR2gUXDiKg+CpQgNBTtc3B2FHc/F/Pqp0t8rNaU3ikQpFsLu3Uaw0i4NQxYBdP/3YIsy8+uHEasO
o0590w4vphdYL6NOobDNUrtkybIHJgBjcSxe49ZmsmKyWzJYg19S0jHZ8mSSli2pjkxfkLhjyeDo
lOms0akv3EuF/ETWfZEzBBdEr7HEkvfI/1CzxN6ckndrWHvEz+ov7+gC6C8VpESbhliqqyyCn2QZ
bRK3rCXzl4dl+eKd90IQPtEi06qLmoJjt10A/YrP51U+C9K5TI2pG5GMpvVdixtqhWFzHlBkxoTk
hlYSDacBEAAg5Dqu1RS8Qqf5gvloRQeDMcxpNV7unVtzGzeGo0Ccc0hGlMNZKqTb+su28tFQ8C8G
Vxxo//rmNWakN8ncDymWfTER2j4HrI8BJZv7/zO3HWeTaeescZkD/nEJq4DUaKmJbEq+57TaH0zU
ncw5fomTBg5DVdG8ZePQjmwIFgLn3joMbMoGr2jkJ2LRgCB5vdTUafqpQo4lRawZfDyuGI+18bgi
8cStfk+RDIAKfvoEcPlBVZLNShWBNztf3drrilj5R7J77zRccofuWtB4wtODqk0RR+CsBri19iVB
f3sKqO0l3LUVSAxmE5EYgakXNCnbGbsRQz+LHTrfA/LwbqmGG5hjMl9I7w1pjaVp8KuG8daP+TcU
olVy9mdbyyO0K4ouoMTz0dJM45NszOS0E2he0nm/3mqGdzYoCo3av3NJ6JUdwJ5Je3o51DK+WVLv
WE2aCQmAoxHietyJHsI2wHjj6cY63klmNl3qkrXefhYg9JgQHXEBYshU4b+sHD/N8R6B1otfMQrI
+ET61B2YInB7kPw6WqR3/aXHeR6CZrd0pdIGxHYM6mKop44pgdgq/NCInXxcIAN5+f7If0Yjte15
gerZ1zt6gp4Iv9JwIhlZhhOEgG2ulcvh2zoo/BnMZ3x5jI2i1tq4KIg89TW7Ucufuynyrts7qPEf
Gw4TpA+KPVZqmHk+Rj2uvnv+VJ+6m4GP13CB8BpSWppMIxmRUVl14cgz/oTRaA1xhlWsqiV3Tccq
Q0Wwuk7L7+4d9CFSB0pzKg7YH1f2gJ4sUQmYPh4tptHvXZI0nSo3pXY4oMdeMq1rU0PGFQKG4hAw
b+/jWWktYZaGm2yN9fjD/hgsQK7WQwF9brTcYvf2NY4wH6RgKV0iJfC2t7cf2BRefO4l+NpMIvma
VKmHNUSVQdf1rLpeL8KQL+kPInqL3WcdPm3rKvyoEbNF+ipQdavjAHH1hbRxl7IQBOMQPzLp/lCL
EuFj9trnQaMAH8l1QPASSiQVdA35wc54SAw6FpO+AIq4pzywfNvufzUwUAjqnK6XzKjKnr79eevA
29NvL0INzQ/88O2ITUBukHtEwwgwjjvzATCFEM1MGkJv+h+ZRX3TO1bDiTdwR8d/lmiMSLQ0WltV
AxPla7cGlqdN5dfIjc8OBHOwG4kILG8AR3vKw2KrDmjkLprqxXMmfsXUcFdpWrj56xT3V1x+YDfy
OZGcBwCfo3IqHsFd5hlCsbtsAlc2fhfOPisLdPwrSfHp5BJTb1s0hgwAua56Yft2Wd1mPmq8O3wC
9cEQS2ro99m/cQ9YQbMp3SIru4b5RWFyP1pgiJmp0Fri3S5ES0Is2CVFWoXH9Be9Dl5z9jMfHty/
GaUf+Xwr3omUSX2feRwYOxM9xb0WEwqwKplddiFg0ULIOIPxLxTFnv0Xkseh1waRb5SllEjOZuFq
9U4pVKJInu5JCbBOq732R7vnkutZYNc4WMhJBQOupQM8beY/flCC10cptKBg7LgP3RFOEefMv2H7
MTWbQ6FdN528FytqBVIAaasyzsleJ9E8BT61Wtqp7eEmTT2LFdPfX1uKN6McZwZ6LpW8qMpKiOYY
gLCPH+M8/l16gU8yyPj84l9qAqOXSEMzhj+PLy//eUoqhJ2hXrPTyqDKSQwnhe7i+VLA++REP3dJ
cjcucDLa/GZnIZ2/kRno7bo2mZIJqSlf5irNDULjbbgMOaOPyJuauFVerEYUt9wIgPrS4Em/X0dv
/fXdm0wBCy9bkrokSUKJTRJCMFqz4yJFAqfTed8EIZl/Ryy2JasmhuJ6Fpmfl8yHU1m/4u/XROuJ
zQr9f+8n4QzKA4vTB9jubAmPBCRYmQ05zr5X71fzxEJW1HwDNknuxrFlsOkNC4hipK7CYhwg7ki2
+ZzdD5hXmt8vzKID2bdR9GEs1rhoiKiUTAMQAKvW+H9atQ7vVm5bmwVtdWXLo6vxPhZHS/jQRgjK
xdoTJC/CupexqcMJm/IC6+O1aLdNMuV9c4vkfYlAkIdXVjuyMtOlbeyXJbo1IFIRZtENGIZwhmeI
Gd6b0Z7vKyHFusvqa56R/QvWz32ugLAVTwMJyN2Ozx40w0ijduupS7NoiKRInDJdyT/UZmEilcwA
/2QXFk/YvV2WQ9iH9YGj4wmn2GlTSpKl4hYs2sDf/AbeE6+cGfdU+LIo90tnNCiPZM7nbDCEivG/
aSy5qnOtvQtkHGT4ArTZsOQBtYeT32Cm8xCoVsFHRrNf2Coefm5TovP8PfX/szMXvKN2DoBkUN08
vtateDCf8lcF71dkeUpYLuUWWgVGj8y6w0Q0bfbw6LzMb6Ub5e0RhIqUNTe9J49cmP++a7ozQw1Z
coNUFOCPYxpeEPidV0HVEOpfk58rfk2TytJvkR/scEk/rsHG7aPRgC46aiEhW2cDGkPlBIGncmGy
7G44XSd5UPkdtpPOktqNrJIqc8SZSyTX2o8VXPUi6lyCS3WhUEtQgAA5eJ1g+XYaHtX0ucYgXteY
HqHjtzRlbFvm2bQaY36/E7G1sPzs0BiSjmEMKfSyb9deb419NFOGzL/wV2sNIXch8xfYDmPXR6MA
0hthI0NE+zvyoEuTrD/2d4tQG3uA8R0HKo4G5/Tb0sECbU+WiSgWLkDTPNH5z7G+69h/F/nS4nGF
CwuU4Yotin/47jFRO6ZehXrugd1rCse7JOddQkwp0sfA5m8uwYDTEW1/N8o02AvuWxRT9zW+0N9n
OqM1VpswiLBgkM038JsQO8UR8CApVnNJ/Og5yk0xtPEW4ru4fWyKcHjMLgGMQT685EQ/fXpc5xbH
typuPjIrJI91sN0o/uDf9tkN5wWGEsgYLm6mpXYGwKTWFqYMA6XDdKttqMb0dPq73v9Gxk+EhnXE
ShhoAKjuFkiRI+39iIS8T1QRohotrimp/ddf5GxRoWujr26qY2boI/8tmZrKvEJy7jBC73iWmAG1
sfrWxrcg+8fJMtgAKlybcbRkBDK5SLNUG6NwjA0mY6goLz5XEtHhJk85JbVWadaOaB8E4VoN1xug
hlDmX/OuZNiVDU4GAuRDN/Ar7YzQHzFHkvTdHjN7ul14OlS2K05efZlW6ZzKYYHW5h32SzeXGioC
x1/zEKBn3G6vDEdjTZtZazRH0efyXAmWt8Vp3rbBG7NlCuZFaeoUPG0EO3fuVDXyMPAIiQfKWWaZ
BFSw+dWsVNNw57q79mVA/+KUctD0LgtKdaf3fN03qlF5AgEl/PWth8Ty8lAe2zOkoKYSJzykIp+I
kSeb5+12oH3qYahl8h25hh4SZauCMsL+4YjSbukOpfzixaIrQ5Q/ELm3J32Vo8Bfl2tRj2Z5G1rq
p3CeV27vuqopS/kNzckfeuoLlQWmTQ6qGnFsQ9+MIJOwjB/bORMHc8yBr0RgGCWNfusifEIMbTIh
fzF4xq68YWcH0j4uXvmKave5ZKhJK3zi/NZhOAxo9jGUVikL4EmiaZ1eryRVfGY/IJJFEXdy3agg
VyCBwn1oY2udxFuW3WT6UkcbPENbxEkOz4O02su/46/t9N9wlhhw0UaIzScJE0obrIV9Mjsk5d46
LE20L/Eqp5dTxY+zPwoSF+65iLlWMfjCJMuh6v7UVRVCXba2ZKO0AnCaN5tkjYle5+9svhGZrD/N
ug7rRJ5y2NvIO4yVG6dgBkFaw+2pNNnp105gGZIA2/wXZtcv+hZJs2kbbdntmUeFnVOBFA9DlDTA
2W0/uLkG9h0dy7kaikyzhV12i4Dw3alylmXv06d7tOcxDNA6+pDqD9G5cGftdVWvNZXJKtReT2jL
uIkktDQlGr/zBQozJjlH1AxijjFDaytkPQnWuaobV1eBnBmEhLUYNE4Q3K5JjsrfLRhtOmFgzkeg
NeYbCik2q0gahIkg6r/mMWqB9zKQXnupxb9zPTUCjIfSIkyIqHXlxgZeV+SmMLIcyhmN1zEPpp93
gTAJ9JWgf+IXuQROgjAThrhCEtMVKfKf2hZLbaqvy1vlCxdU8fP8c28EHHOrEcjU1ldAFa0hkAa9
5USqAbCvQkbc15XCSjNFlaM7ebyDIQrjG1gubxQtnvLRqRD0gVu0xq3oUB/tvr7tbc9jniaUA8A+
Zqmy9VlnCqDbB9xleIGoCH/45QkYBZqfQvLBucIN+L9NIDhrXWokNdZds1dv5UFu6UBhg90X3pH8
RTdb3INBhn18k4oWzsz91ddRGrIqBTKukGWpBlFGIaLgarQPu3p6Q+T/lSnrKQrHPRBLyV8B745V
b7K6bqdvc3MSKYJ/HZCYt78ct8DSRx9E6msXX6yOlg7rheMjcut5yLxRsYdi+LK5/umlsJVS4nDf
FZKjW921Z1kwiV03mND/uOU3OQ2hNrEGLC/lgup8PFfnQAdXsI015yv00ZL+WSwLEY1pObCYsE0N
8A6m85Un3lkvO2bM7/aiH3UoEoWBtaqtL5YN4XIJgdbos6lA3uNrrJktOkvmJFMtbnZRAdadq84O
ryLgqfiESIIKBjBXLQpkvsF0X6DKl/iC61Jo8OuvE/FxCeuSEd5lwoFaJ/DryaOAvBm2Cx6olsDp
zreqPGRNXcmtFJ7nmvy0RnJlwoTlOZdGvvwR/fS33V2E7hBj3yOr1PbciBxC2ce3Rx3lkw/PSxQ/
3+6ckaZ8EpaAj9GJS+a3CKq7oTGikfQEcI9D7sfyb6RBEsxiv0nF7W76kTiyyvEbpZp8joyMXU8c
EUdD4AR98GlNX54i2l+pAwY7GHdI2bMPD2RfKLgSSptIbicmRmDvHteHKy9Buytna1gFCBnnz6WW
MaHjF+9X4eKCQNu+96VRxTJhzb0vR6X4nO18IoI4VaOJeUFSvf7T1DERxcSq2bRBlx/pwcVS7WqW
xN8kGMt5UT9MSmmuz+ywEps4cQzfO63hJPocuP8WlKHQ+5pFJlP2sifKkNLECOUV3L5GLqLwC8Zg
Albwgix6wqFEzX0UJjHwpZinWb0x5hi1GNYWI7oSW4gBn9ktuoVTQLrl7coHwBzJ96UpmkYwRDWy
wCA9tjeNvns0YB3+v9avddgSlDBVWqWrXYUaDdUi4Kc9yM1YrCtkMRqr6Z9Nm16JX6tx9934CzzZ
zrHm4NR55wPRFNOIPKquC81yxAb1dS9VJjh7Zl3ruEr+zAUJhKPHq1RX+I1UaLS29X+UcXiEkW5D
3dfx7kMwMesVI0LYu//CN7CM8ylXmdgh9SlQ7FiPmIdNjXxU6RRypzr8OJ+FgVyWo9DajOGz6r+4
217cliW/doWJoNvZAqMma+IYqBfDFKprbkDel3qeb98ffVMJlpphIzAPmHmqLUrqgNDTDzz0yvgA
eK+cOigFTgN6gnWAlzgs08K7MoMR51a2vtR8AVSS6WDuv+LmZf4QPnbxBeK8UPARyKnUBWfAZTOx
h4xRSSc0TJmtz3KiuYihZMTbVwFjYiX60VXccwhi/dNr+wtO51YuoJbvcaQvK8OkzOquNWbimmpE
H2kjLvkQq3gvZ1lznkIyAo5k0x5+ITyDiNLHfJzS7KTR6zHHogMc//33zrKS50jKC840Q+JGx1Wf
6m0Facjj+iimiATpubdNzFjtzTeGnVwXRoDIgvXPc8YsN0xDyCixBpsT1+TaP4L7PXDOlMDDIyGk
x1iJ5FOOnvoirvvA4UZsTB4pNPUrx1UmiC1DF0/U81EVNFZg65M5dqs6cBhriwYQegNvFVINmlXR
flPhMCk1RgE3oCdiDJRlTXFOv2NO99ow0o/GyA/7uGkMYLz/jxQFoyg6+wbgG6oiIU1Ef5AA+o5X
BbV69mRZbKAfkCwOUMDUNKLxKEqQrWEVLiJ3rgYVwV6PNie7dOhr2I6SkTwbZqXLRpGoRxv559Hx
3GB2DJldb8WwrD/2YVLs2fRAT2Yzahx4Ma7R6IALu8lVqyPT00CHW4k0S944Xz/8QU6vHsLm2DF5
VvcUjUaAEgM/JTUu9zBtYomGhjqVevTAe0RXANRbwb1ASFnfkzmL6vZHn5zK5pyMTr/tuAkEh8tZ
1ez4dzj6uG56Y702lEOIxjowqZBb1OFSHL3hy7W1Ik9//3fPZbgPOO0NXHOe1n7jghfEHxjHpJYP
JDoT/l7Winrz2b9uOgpfdKdCr4jq7KVXEEJPUEIGUdPFUEeHausJBrMcpRUNaBOSkwrEayrgBU4d
rsZ3VDnlIeeUJNGWvpsep2VS9F/FST2C1fEekiNpDKK1bgjxc43dkRq5Ow857F4fb81X5LzwWweb
gcZcZr7ecXl39bSQmiftz3hSbQy20jb6yzL2csUhjpqUYNxq0UCA0S1WbYsiiQ5UIqqaERv//8ti
319KPcdesrDo2bcDv4hP+GmQ7Ln9pdzMpb5dJ/D1MbU/kD6B6f0Wiaeg/eCMWCvm2Gwvf5BOrRbT
Zl7aQ2wIOEnnvLs8GRiCRkZ5SJDg2r6/g8Iab1FRxYmbb8hl7UNVGRIqczuFeqG/TukpsbwwhOlD
hqTFU+r+lN5yY6+o78rCpbbKD43KuOCYTyFpt9fV9w+0Zqm4H+JMI6nDx/OagrCXBcz72U5Ch7cD
SZXGDUqb9r3EAyZ9bZ0v57vpkjTe8ZO9mHe/jC/nSNsCnZHUsCNMoSIhxaAZSi1ALSk0B4MAK4D+
L53mHT2NqzIw9rv3wFJ9KagKerSpQcRnq0Ax7ippMkxcqFW55snlzXac8l9t8BI/CyXMoj1cfwM4
HmkmxJY5LEZFpCakVXYAdZVOc3mE/akIGF2tFBrFEspU4Hja6Q9K4o/v9AYisA2bDpeP8Yi9mfPg
45UtGcHYh5HEByCua09MYAfRUEfLJMK/A1F59RBQZAfHF90Uy4Arobs/SOZFRWnaTn3bgJe4oHzA
kbk+b/NC8JWMYD881o0pEU8GgBggHvaK+yKrBobM6P4zY/QhhUa6qt9qHgT1Fn8Ws7woi1g1iEMR
XFAjW4vo0EuOujnZIO2otU7bOGe3HqUJcXhk9OIb34TUfGQv90DsPsw1p0ahj7pB7C7iNPEqBwpm
8stvAhOR0GFLUkT3a6GONW4cQKXrAOnO0AuAvt6GjHwmHjkeTxyVaxRKzg5wmgJh7cOekhGjj+ub
OtT5alTeOpKXAiJk7DAZPIUaQR3krRlFG9Vlt8mAMA7x1bmk4OmEHcCxgZwrec6WnVuaKBzwGnjr
bQdAiJTGTSweI19D2mQsNgDsnIWIM99Zs4yzB1Rh0V0vNgYnKEXrZ6wIQTo5ZDdGJG2dkt29pFou
0vTWBrvI/dL9ehazNGrffdV4iXliULyee6orQuupnQP7dY6LqmnG0MDsrGFsWy81RCc6Xb6VFDD3
b2nAD+NQ5pI1mWp0GHa/40dxSnBLg4PXrXH/XA5yhLklK/DX9kaiGs6xh0wakVFYYHXvKQO72m5T
Bop322lRTv4vCz5KbS6ZQJGrpGFFXAoqwB+qlVs1pV82SoG+PEWiP9mZ5Dq0AVCNL7ppvQ6+OxNF
aFNL/Mnde4lkMScr+ce8q57cENLVuGoOmVYMywxlNyGuCTXrVAg/vpVHLJQwlHlHYmzA2dGLVrMW
QMjB+MDCKfSKQXZT95jibGSqSUFxIo0RG5yBzIfB/CZgarFEqE60/2mvAHM1Rrtwp4NIgeBR5yX7
9N8gMKqXMAPg68R9pBNFat4ALDtrZB5tH/qOyTAU27qCNGnPDAK9vyent82VCtruRuyd70ZX03P4
mkZMUsA/Fy7Iju5iVbBGezWtsA9v1++U40HkWg8TRgsK4ehkr6RIryXGdqV4aywOVVbV/d1Jl+jV
Qg/AeDSoYD1r8S4u2zmUO6xgusgcWHO8VbBrjcKyqW8g/WO1SK6IdBUx0VOZVk1eXr3mrn+xAemJ
0beWbSYvx7wxhCywxkZPXnSlBxV1GUaUYQtB2S9+0bvyGgW3XySXnHeu0a9vFXYYgnSWO83v93Z0
ond8/eGVJtH5TxQRVPuD62FbL9F1x5pVK5DwnhKIafDi/5IMvvF24eRQSmsmN7TYSyfoA49jvoqS
4yYmytH02qYNEqXDr9dQI8uH7McgXNaZq2tu6PU4dIDT3s2uFcpbvZNemq8I802hwvh0Si1FOl3K
EbXkcp6wyZDT0D2TPXx0g74icyV+kOx/gTwUewRfhaEQFXRBjPlVrqG2jMR+sl0iTLgejIz+E2FW
OVR8EQ7qowuBJlb/EjWZVv1xkaZ63tBoGyHCYlX/3+chUrNnBuCkrBcsFzUscuLJbAXzQEslfpx1
ThI49VQCpZ7Q4N4h/we/W2yvR/nYvp2Q2GpfOA8qGtxKFjRHjtX6/IChKjHk9VCxaRvvTe8wrgr8
5qiTF+6jWfLhB7Yp1wRPLzRlTCItUav6AaQh2WmcKst9YSVwAsslK6e68kh6MupAxkVuwAhAGxFi
gGIsJbKEs9bhAzLalVVvmGLsAu3CSuAlPLubyV/i8SkBRm0WvDzNiwMtUa12R/rsJ8vl/f2zMogB
AG0L3jaIXgVHUwLF/0WPJ7kqEChRS2euLYvoe0B8Agw5bucanoEoZEgDlDCkGRyQ2GKrigJSK9VU
TpW9eOHT32VrHBnkKCAIZxGBLFj/PpRoLGBZXdMiii0mjBy+i+zLlPUCHb+Zj4WfFIc4tHHJjs+r
rSr3RlxlNz6owz9ICylmkpuugLRUriNa+rPydjHFV96m3IvL0UeZCPLXtuCRkJ/qBtxQEcfAxG/0
PRA3aay5w1zweQA+X1xi4DoYYssCqYB84pVB6KKwz/gE51yEqD+Cv5NizogL5dmcXYRYEvhvt8gA
PPeXHfUS11Ek7QixEyp6R+pcFT+5yNoN4xYAbHSFZlkWduYKSBiSId7Nxi8Ly9Ue+Q3EncdL3s6Z
hHRNntC3CH32H+QiWjjc0icwAjqPFpRj974yPDWcTNH2lOSMNv7K+8CqvAeHiKf9NEUtzHRLDiUz
EV98SrqgTwnrVPGfsVT6AgW/qFbbwqVsulNDgZU6mO+QrrQ+QsUfRfF1IO5kcBi1wtXCDpa4qDAn
zbNZYl4JrZ9ljsS0HT8yr/wXks0sYcZrGqcUIQnR5NJ/NCO9i1HNhsVLp76BWUiXUjaJDNh36WGy
eIqe0YLalR6KX/Bq8stGdYrMYR25Nao2PIWhfjWZkETSs6vihAHCVOxFEVyGrINtMVlURLZECTDw
6WNuZvrFSbk/Qfc+BzL7dWSxZARglWypP7JnLvIE4cL7T+l1KBgNlpAhrt42D9+xdBlni4rfzmiC
p/j7hjVf/OTxwciIz3UTOIwn1PAqM7wKcMR7HO7P2qj21P+r6Q5fS6rEzmAPtgF4n4VQpSi0WMQ+
J1vc6DJ69DmRap49Q5K2kdz51Li0LC97royp+Fpiog2w+OAyzYOZL1Zahxst5XKaTExaQ4jd4Juj
77pcrTrNSJ1wQwR1YxStNOTAOC8UwgkMCfmacuF9SvdIT0uDfBWeY+x/bn/9GSj9nxKq2VgSWJli
t4EODZx5T/AokAQy2vHgqassvg70n+PLCJ5PMIo8+x5JXZW8giPenIw85iXdwWQNC8tsTxD5lvdK
8mABU5+du/qO+HWiQGzp9k/kZOOa1AIV8zBssg+O9p9qOceu62sR6qT1FasCvzm7q4zq2s6p8cyc
Zvqlu37dqjDb7HFyG5qcn1a2wzln0xTbcCCUYEHjBnkIezGTCmsUwSmmLifP9cQ9niMUu/NLkcM/
dO8AfqNfySiaFtjJI42N0vQy7fUUThGXEXgDu9QpbPR/Nvfxhk5gSMSdU6gLurk3samwnw3pCAVh
lAQ9MZEtIUAltdbAR8uL+d4i5YA0DQ/evgg8+kLNqPaxTvCndF64+5X4Rq9WeVD84SOwstyMuOKe
Zgsl6p+DWYC0eqOqNyi/TqBjLTQlo4y22t/wbFBWA19/eKkAMIzJW8DJvjLvIMmzSeM7Cz4GQPqT
5rZGRlUcpEhBiT5Fm/9Amh06rhOrXs0ne1w/qYVRqO5AncVTHevdTLUtYUys+keuI27L4lMLaxYK
gC27apNek+F1p4zRXI8ntg39S8jrr/72hnE6RmJV7/eA6PDtggrWXDQeArChf7p/ag7hhZwXj2AK
LIy7itwUn6fafV375MZzCIPlRMxVa0pf52lUZ/kk2d62D+R+pnL5AP0VYu2Zf+mN8s6+1i4nqlrc
cqznY0SW5ShdBRsybRAwDArQPnAz4cxZHD1bhr99E+11D0kOQj9IBnZNZU75bDr685eIs6naL6lD
8vgo8tKW4sn418vGUfa3F3Ww+npaOyfSr0oQ1z7L1vyyIGPpcOPA+He/dpWWRnqSEy2ncq4LfRA4
G3uZ3L1gn8ukzC58lx3U0LCX0OY7ILnQ/+nxAIGRgdWdrX291GqVprrALuCOf9IPLg9ZyOayVaAZ
0WxWBMciHCNHd+rkqEfQ9GYXwJ7t5PEG3GzA/HbPUZ/LYys9dS+pl890wivtJdASrrXrvPz6Gzzn
mvztnuT/rc2fbKnEDKrdOO99kIkxRMo0upFb/KtZJ5JTnYxYp3n8Fpa6r675ERN9FF1BURJ/rgLl
XsjxfhdUQiVjmG5XLO9l/yWk+DUyO0iV63etYkW/CrvqhnY9pNMaVyX2NAXnbxGR9ZnA00Vosr2r
xO5LLnPXAebiFKuNxlipI84DKXZE4khY1hZUSC+SHEv5kUoyFrQ5utwvZjwXVeEM7fhpY4zDpqiq
qcLSVpL+MyPGGzAUaDjDmRHZkqFDFSjYw83aa56mbLIyPqx9UWy7d2I+YOTJEuRKLRc7SwO4x/Kl
0y/nsjRB8q6SRl06FKTbPCFjB447kJ6lPuHv78dIke1EVrEIlxM9zdp+lu2hpAwUpwMNY6ukVsA7
0En0ayJV5n4IdUYZLRac9iZXkmUmMq7KzzHovMA+GesL936dnLVtIXfn/qGO4fjqAs0QDVDQhY1c
1pKXKv2WAN5hHFiEz6nIv56xrp1f1GOwrSw+ip9AA4OIJtiDEmQ5zjOnqlsyXIi4YShwl4ENoLKe
/AezCyfzo7R3Qtq6yL8MPg0VXZ681ZLknx4A7vfWWMNon9mhPl8PJ9/xugWaZyqy30AoXdsgW0uL
hyLD8dBH+FypOPhbkCd1W6tsl4lPL4XbDBoZoCHQhvSbg1xRBVJHnt1SjirWh0gQEMl7p/S48FwE
7eSKvuMGb9+gQ727QAWcgH1iD717fyBgzqsctDiuIlNsvK4QkblxjUyfA+RYEQKRN29ciGjwRKix
khdKnoZbvmcKwrx+MP+Fo9xIqqmMn7NU0os86Q6CPMCKjnsd9dsnodfjvpYl2GlqL7Ly9hfHYVS0
W9+X5DevHZjCEO2O1ZUEUNTaeTod2hivycjYJCukTb2EGQ0vBYbEvVaTyGW26pobEIqK78BnN4un
bHb/kFp5scRobLFNtD7KiitnxhErt2ceANZ12bRGpVNtkwIhVIfIUzoMlzp4Y1Pv4Nj7orVJKyuh
e8jVlNJ0jOmMjzNFErA+ORbkOoXvSIXPbYo0A/lAhrrxGHvfagE9CNjMMR9hRD3Xm/QmTrO0bU7x
normqTdSsOcJTQCtBrCxPejDf9BEI6GmP08KVhF8ZLcGE4Zplt8UbkDXLw152h6K4RGtU4QGKul9
UbsuKJAowhX8wMH9dnhR7oCH5v17JvZj9PHMEcyPlawFHEEJ56pnSPx23oygm0D4P2iu0OHK07tm
ZuiI4sEDS5d7YtAi6KLgUy45+/HTHXMM1Jx73uS1sutr5bQb8UgyJagKSnMkpRXXA0Z9+BqsltEZ
jIColy5v0BYQraglqO2r9eC7Svjo0Vac3wM5Lns+T82YuovD6zj+VSgY1BWj9DXGb+c2mCyB+0ZR
1jgDm2rmw6ojgQQOlfUWDCrMdBu3mjjSiRJvYsOHZ8wsV8B7+EIAqlBfSu0OhFqMhQGBtusiHbSU
UinNzH9YYw/IXnNzpV7hUup9qDJsBN/rezkBh0BTRTo2fa/bISZ4Bb5Tr1pWkMkOJatAa98fgzhI
4q8pxeJ26kcSNSV3Vj5MuQAObBCs7jPIZ1z9Wa2o48EcWRW/+5VKV6J+Ufs5CRAsKrPV5FMMnCzD
YbYrtumveIgf7W7ptYkigxozVZUj33S8Qie9/nDNzal24/4OS5u9AqvEq1SRqVCiAhYeflu53YTH
0jmQpcfNTkU+BeNwHdzgIX1by6SwBPoYm+zeQdndpgfemuGEHY7roAgUyb7nFwZUnRqvelE8SWYg
C/ImVVT/UT1onz9WwqGjlLnIedZDUSdGr0ONkbmP2JIluBFkx/uO+QL+bKmqVzMKxyw9gLeXLFT7
pZeY342ppxgAl+46Xo0CSWl6nu9HqtKurdSpuzdkpExvLMsRwrUkNE1G1GJdZNg32XVJWhI2Dc6h
HfW/WVWpN784rcyrGKRg/JPvk5ZYAN+rJbCQgfEvVGL8AVz2BBSsbZ4lv+du3ru646knYYKp3Han
1/YAVZLxdsolKYkEAYlICD4/wknYOd7MGItcrB0M26snXvmxbEIwxS7X40sIHIRISi2oveIYTq3a
O1JYIRiHoOS29KbgFUCcxPHvbV1A12YkFsVI2S9HXFAPugvlR/8CBjDLVQI78v6Z0989M2Q6Ixb8
qvJ1KjUljCJTNwOZ43PqkmCpzBrjjv2uKRRAW1Z59WX+Ws+PZ0xXg/dwcbNULFFG+LMoXTUQOZOP
VGOcgfuuemDLOgpqrar4NXFBARV19IHu3XHGhw/CRPgTqwMz2V5GQlPOdqMDZ1hCDrZFoBhR+UBt
gbDD+bU+sNtGSlO1L0tImpxBYpl8sAuHIPW/3+izqt+7SgCOcDdusXTNfpmS5GsCDYnd5lVPL/Z7
F0uSPn3hrUajoWGqDGx3jhan4i3p5TKuPcFymhMdSB27yhA6B+2DWmNnNsZx2cBAp4an6yPdyK35
mErIo7aGk+NXFMHfbXhMTX+haI4ERE99RihG02hTGUU3loIlgvYw3euHYydJ75nweISjy8GVKpa6
K5yajATLxF4RjxPVF+j+2zE1b1OnH9anmHmYO2cbTPFqlWWYY0Q+9PFt8qIbwZeJcyArw8nOIT99
aQmBzew6Shu0r99jn39brcieJXSN54RCU5C7h7Z/oy2o/hGa2CsyMytYMlzLS1QHPwQX6Nq2sgnb
q3xE7jY8eWe5kmECTJGrHhq9zuBQGndRfQs75tkNsFev4qWgn4BJDpDrnvPDcJx6NZIeScjv/iy7
f04hd4i7XZR7/xhRLAm1zcnxBfL9imEXXEmg6QtyMVq01HjrP3n69mmanuufiT+PeYO4ugnKmOhJ
Xv5Wdn95UkfI81utpwxBKr9iP03OSCJ0eZReqegLUeT3k8j4oQh7k8FSFAsITtK2q1uPBv9kdcUC
uRbW/s+bCy6sU1MZkEQYDoGyugqghuAPtam93thc+3AKfS9CFW+qivLJQlsEw6GGTNUNDpxeUb0O
Qy3DBV/yuQu18qjI3lgAW6dc/uE2E6v/QqA3VpJzIT8S1JgBKRYvIB33/63N6wjD/4bc51H6avWY
xhGpavu6aKjcDSh5gj229EsOKzdmzmlqDAzYOH8BiqG7KqG297OgBq9UmXheHVZbZgTaTqKfOq7I
k733UpxPdy3bU615h7dcXJ9uQRcbyoGwSyxiSEOvfI/q/Wxj3IxqFK543Z3XsYpILlsFZA5HvUkp
KooWTVru57zhyew8flozKvMS0I8EIG/CxuJKXdUyJGKHapmpapr2B59CQUEq9bqZUFbn0cS9mrSk
caag33M+51YDQYqBMvkehTQ54B3tRMCumjRADRl/aUEdE45byG67th8PANPXD9Cskc5+9wMfVujx
jy7JJgYLV1BBA4grYOFq+mTfBnt1KzuCgII5jxImOTxBEEm+Pkviz95GoTlyPFEIl9Mj1VNVl7O3
tT4R5mJjljUPA0JrEbza9tFsQGyqU5Pc6GQP25GwdpEB3n3YKD+U+kPJeIQ/7xuor49HOY5uQxSE
AZUx5kaN8NYb9mrY+cBJQ4GSGxEWU7bM2uLce6jPP1vuDCbm5hIOto0YsPwY0Gn0nmklagDKz8ti
+v+surZGoFc6V1qkY2xbbB22iCvJoMRDGukHkxeAxbCVk2/8D6NaDpqTMIIOVt5m8MB4pLy9vOBZ
d8F2SziESyEpPRag3X4veynPxFClQFkqCKQ1sBXlsp3Ec1cJT6iFcP9SAu4fExGCHd0CrzEcsDOc
NLQwC4v5eqpSlQn/QPkE/pg2DmdVwwdOERRYJqmWFbgKjIM3WEq4KOA5DiaZ47GR7W0yI3Dm0sUd
lV/XogC7PLaZNs7XiaIOiTwdYNtNRQ28pixNeO6TJPl1zlcr3yzee+jwYyp86isWN97DrJB0oceV
eIL8DLXbzK3edvNXIg2GO/XTJh+u7IJT9QUM/xaUYora0ssU+X70YBJ0vyYDVNj36oEae8ie4QwK
ou/ou6fnIFXGzXB2l6whwOXUyBSJROzPlSoh2Jg7B1K2hbwOstsso7Ubdh39T+8fB/apOFip6VGk
gXY0RywF4XCJeEIoi6FaEhTFytYgZmRSmntAH7Uta3zOEwlHsGm0cS1H1ZMSLcuW6fX7GGR/j7qt
IAuutfkHJ0gegqdNUwSqYw5juWtnheKWeMV2rIf3zDJFsf8uCD0s5B53dlzmTYvIUHGKrWQAPhZt
TTqWKc33zhp7o6u27CGIYS94dxN2W2fPlwzIXABnQhPe6u2n5aBtVyHO8n2l3iWboY1Ar1DVi0TO
SrTaa8RHDrP9jUo7BamFVjiqeLxkj4KutSkSdCm61N+o/IrRpYwyuDmvvX8hDCvYDtn3uZxwyGoY
+q4cEIq6bJKOGNDYyEsVH78XfwdF7AgpovefGuMW8FbmewLNKBSfkxtkFBzSAnhKWJ8ztxVU0rae
TUwRdxDvn2AhT8gpv7C8M2CvmZTA8fefEfZUZHT9up4dmnhZRkRXr/07PWLnyc9kqWeUYLKfzQsd
AV8gtYMT5+CpliUo4cwbFB9eW2yzayb1PUI7sZkngmRyTkZojdQrTLCUBtXS1+0XFI84//mSVg8j
+ZAiQdq4W39DAXuzDXUBcDsuu9VBP4/bpUMbeV8UuKR7wxfKQXCvFYUH4Rp8cAXUUywBmp62oPxN
yBPh0aFeeAXA+LCgEW2tjXLQR6puqcZSsIsw/qhM9rhFMx6q7y1Y2NOfiw5gc/WDyFY3ZjQtiyaW
9XveY7rEHTqgkqPzLSZ0o5NRHBUJiNi95ZlSr3nzPk7SmtiZaCZ5xPCTkB9zDQfPeomKZjWHKl8w
RNVrpJLyKLy/uTkiXtH80Okg8XpuPZ+9RmCbBSgogfITjjcnDJPauRRJ4rOtiJL12WryxSpOyshJ
8g9E+bMKVg/QrSXJv1xqgIsFzOVQAKBZbU6zvmFxNiMC8fBKp2RwWRpyqaWHnb3qHYDeho4UO200
3cRIizN8GcG88NJljKjnFHYdrcGmlx6pGyLJUsT0bQLtd5hCoFGN0j0DnU3/pzlM/SHDO9sNF24S
CpKEZiTyT8XzXVGmI3/kWqSH0XlKXQGe8GqhdUnw4JL3stvCm6MPxcZFJAVsf2NimeQGSHkv6oL7
3STx+JNBDpFI+6hdye11wI/+zCqkozxScox4EiUOSgJgNY4GdcnAMqZUWMIFyejpd7l//iwWPjgY
1WpwsegQ0rBJTvSj5NHUEKtQll1J+pFDySwfadym3/fHDUFAyvxlwZJi7GkvYSayrOOv1O9J1WmZ
9ZM1z8gSPAtBqm458YXsXnxsr43RUXfcAMSwtqBY6Iq6tSPQqSd5PyyOAPKGVAd1WMidnUKfs55R
Z1iMmkwmpdLWQLxFwD9WOg37AcQW7jlfW8V1x8TFdNfCoUEfWYIwfAaBW2NuLXg8vDs8OadDebvQ
o9utdpYjK//R66wtG6p3v3lAwXGmCpZ1NxsgKyiqnYD8NN5l+YDKmVLaQSuW/zfy1512pVgVJ1dV
HAhE3BHyAKFMkg7LE2QCKmL5BnlY5sBEgAI/luQV3tuRp4wzV5bHdCZF1iyQnuI/dY2qwQsAigec
87bZXUbjdWCSX5YJhG+aM5aiJoFhusFdDr1Bmsmgf4yeLldDGLDWBCjqKB7UQbZOWKgzlwFMUEH7
3uyFPgM1ksLXW0usCBq5Y424f1nxWDNrr7eZP3dtlQzgPwNivgqBbOHt5nW+RvTbv2jS1+o6YMCE
Z4sJaqibE3LqwDhK7vNETvp+9d9ygMTOyjaf8cqPUPheVHAZ7F8jsnRgDpf7PpWyN9y7DuqlffEF
2Oe+Vks5tPStPk3AqeSxMioQd7CTVwKkNLPghFkAbpL8ereSkvL3FavPxlqWsw+0bp40AVYDo2BP
JAKCBQT5mrciTVqtu5kGWtDsWn8sChXtq0Zohl0UMTx53uHLkCbxO8FFxHcRyTyEbyBLovIIT9IM
1UAfDqxXOEXnRQQ+YAkHm4rQluyrhtLAUO27uHAqN/Qep0vhsl1ki1/AkSXcEUJv6lfw3B+ftk6a
M1sYNLZNjUladknLTxXJEAV7jQaqR0hZU0CYmxTcl4IgBHDt9PkNzElBCbhGYRkodYvVgonkxp9l
TK3p59YCdhdbZbYWa+iXFgCvmaN3i8nhrOkHQAjYivkzHoIPu6W87wQxNXqwnwPgVSZDztoOd9YA
MTClD0BLAWgVlmd1ora7d60+nhBNxah9JJfPDhZ33Z2u1pzLEreMP85wow2f6TVBWXEYmauq5xs1
vMjpZLrKuBk2W+TKwSWsGReWTxOf1YUKGoSuMMerfzLOfgsS3MpIX/hUi+2zZdal0i0dKZlRx8PU
ni4zt0bU6R1/q9dpclQYLyyBtLIG9Gqj6nMaELV+H00HMKgqbov/kmD13QyU0vw4/U/5Us1Vpj0b
BYiYuEZce0RwyOLYYqaGQ1LASpgeWQyb7WV8dP11CPuLcq3h3EKIn7s0fQ7JveidfwVscovVYFvH
cP8C88CkkpgFXsBWlp9BmJrNN6qTjtr0f7z6KIQM9SXt15BRcRqPy+GRb98J9PKgNa3+aHvvvoJM
1SYmrlL6R54IJLNlL5CG5fIGVW+Vo03ozahvQVRgUChnVpI5Sju9EUkL3T7vxZ3Ms1Aq6iwajpG9
o2pgdWuMt9Nd++O1QL3PhwDjZbgY9an9P/UUrt9clUvrswoFrmdwWr2tz2t8D3Iz/yWdutHF79HF
1vexRSdw2S1ZfE34qOwymbU0Fh2lKKCXMRCvlXIpEqRaMY42GxlvmbGznJBs8PtAID7SmVz2mZsK
6q55tOO2h8rmctfVaBxHXOcYNgkPc99dYEDepOUFq/e68JPB5ECtr767oEkB6D9VBBV4JveywFCn
GVjHXHbBln0htyjmnu6JvXfJijX7gS+RLgQV3lPMaxOdTY4y3sDZ12ui1x69VdEbI77Q+qSx9maR
NYaStZYfHO8o7W8pOyU7A4dRaR1eowWS2Q5OkfrXrumo36SuZKhY+4UlV1W/yfHmoYDMcXr0k0fL
nkuZlgFJkxXlDSGBiHZexNw0x+CVhbC/6mjJrW+y5blW2XxhuZz1RRGSgJ2vi42IoSAohUSe2iq0
ho0PDo1SgfTC7QHf241V08/7LqcCNLtaKOseN2kDRCQPcW0jEjx9yuSkm70IFICPWZlRR8ANC5L+
JB5KybpZM7zRrTzN2sZpRLlHdV92iKrUJm1Vi9DjS/4ZhITyNsIMXdcmJAQUf+C3qKZo0SLuTQwH
4CD0BrNYqqt3ECP94vcUlSXfmlHL6lNLEZryqjJ2c5DknSfemzGuuEQrq5h11I4RHYGM+M08A9qG
6CvfOwJeySXFzZGgUrmexw6nWsmXhy0o7ftqkalD6+xwMSQvBlnZRcARskzpvnFU/0fV+O2bK+GN
EcMBXKbh9AAEVDh1BTsze71ILgcTJE0wzIhgYYSWeqaoZM2bBypct7O0lIG+Lw9oLY9ULWzyqSvr
oRgkvFzdfcTC/daP8kbmR+e/PnG1frjLmRkfzxuQGa2y+krRAD+Y6xbz8tcpPW8QesG+sBgwELxh
klfy0jcAYU9WebqrqxS+7OIs2d9ZXNVqhnAccsoKzO7OnoxHq55WK4WMWNjD5ozG0dS0qUvPrILu
j/iUIS1qjivmryNQqWC7kmdaRp0ZRNdhV2krgH2swW0zMlbuvSccgSLN31zMmGNWhLovoC9cpSfD
FuBUKqnYj52PK+wyjMbF1r2gnsf9zzDsscQcJhjHEblFad2if/bRT4MKxXcWjJPzN1uVRJHkdzAV
iNBV73ILNLGikaq70+HkS+maksBNNODK7xNy4Ykw62iIDW4XwuTBN1SGn+aOucQhQUFSpAVV87we
OM118aa5PtHOXe9rp04ibRa5EVh7egGYyEbJRe8XsDMeNOO+32e/tISjEU1K4weZJliKcf15tv2r
yohrgcp8E/VFATHRO+KCn8e4LyKp5x/e+M9PMaEzVaPzoOCte1gXBxRabocA04h+LMfxSH2UHUBI
z9tTnjydNfYnXi7nnP9PrWW9R6DxHLwW1Fzj1vsKdg6Q8R5l/yJg+kNaRkrJ0/8PSmZG4nf5ASY4
ZAuFmlDksjrqcpxO+iemUfO2mFns8i2U1gVN03CDboxJgZwqlqABVcZkIwzAi7v3TlQKIX9tsqE/
LUaLNNPCGY5ahPtkR0pE4Rx/mIXfh17daT2jbXjq62EIy+I/6Szo0BZS2UuoOYBUrKG9KRR7Cjto
39dKmuH/s9mgGBxOE3Ok41DFRFlc6SvHUv3S4flFgmF1ezuNtzUlt6x2HKYKJg+Wn6cL3wbz9HUr
8kMaR4fHrr2OBnhbStFUapmUnfWNZfB04Amm5ELbRSCIIshedTqqN5/vZrR7IOUfhysANCWp70Qq
G2wL7lxRoY9GqxEU31zU9j+83y6QztbAyd3Gx6MpZOQ5ajCGDANVkrK572awNJME6W2A6DnxiUSZ
DPC9Og/QrlaYtHfRHnccvt4IBEjfp3W7EWzej7s3zAFCwBE17cHJSe12uvk11oVaUcxyeG2BiLji
Fl7gRofwrDc/Vfy2MNntpP1vehEk/+zT+y8TUyXmGwNb6kayWM5R+bmWNYanzvtH9ab4x8t9itCy
o5vNf4gvMuDvHjhGxYlI3rlZ1HEZhlDQD8vEUKnsut2hh8pwe+io2OfJCFhWiZWz9/kNbnF9oq5i
pTcuXIOQuqiQC/hgrjIg3qa5706lz7agx5Oh2vr8PrRlG7/JbH0iurICVjtD8FNoQsJYp4Jux42U
AkMBRKCOZZbc2XL06tbZ7wJAqOfoqI+dbJfDVGNgJYcl1+UfG0w891zzNulPTqfxonwYzrh39Kdq
rvMyNfeYGYDYqyr6hwX9SD78rBEA2JTaLJt+rZ3qVPGAVJswjzlJjeno/cI8TiZVlHkMV88S1xuE
TpJwNIpEvhaO9vJ1vGbd/Hc0xdC4JCNBNYspFiMcY0LuBvqQYv8u6kE8ximQ2OG/RPsmjyqOaXv2
7e2Zzm8sH1epOtXY08FtbP9DScAC9Ip1aKZ+krbb9ZzPE+TXahNsmDHW3/2ha3Y/RFI3MobNYgaL
RUIyrpdP5FOv1+2rpAmmRWFqRdJy5bdCyZ765UMKiTmXwzGxAM3fJmWas8oIYvgXWi34lt/6STwo
LTea0LDk1OrySNoqCBviueYNw9eEWjbDCSFMTrQVGe88HnbmGhc0Jy6cBR60OYF6VxJWRZOnF1PO
4CXqPgGd0NDSHZbNdWYoIgi41/UU/ko39GIQ7S8mODAWVRtj6+mU4JCJkaEVspc+egekR79w6CRN
68yI1Gnh48Jw6QVUxWzsfcgj126SN2vgcpoDPDIi/f8iOm8djb9ctQVkp5XOQFjSK6jouW1DP0l7
9VV47u3yt3ADbzyoVlNOLGCQ/G0NmKeqXHXaMvgIdxL4r05m0S9lZ/Va9SoNUFv0AufZhj9wsXJk
rfNlan//IDoSLogrLwitFXGwnkh/I+9bKnpWkDqwUwV0a7XbgouDNeTuHhF01uKADZF+mA8LesNP
w+oRHaICyNA6QJV+kvNIZEPNpRxatOeCB2sh/VSCZjdnIM38A4AyPI/nAla0yuEjlwIVl9Y5FJy5
WYYCQhtRQUVAVWYkxyToi+uCXOkeLKq5L0bK3oX0Qgg2XHYh7xlNymp8Ki8PXLgKR6jhzj3bUYFf
7gLtQA7hkKvZ5x62x2cLH444AaNHquecNxm373Hu8+aEAYdSqDh8G/y3BkXaw6Raod+xB8nrzoSl
bTeOzhLCU+Hl67O54s3oU0Qe+p8f4rFZSYs7rgY2ORfxzjGxHBN/Nx67W8/XDY2L9LSOm4aUrOoH
Ab2msa+4KL9o6PEwaw7vjujCHATcL/lGa+mSiNtqks1c057PmybLZWpSYL9eeWOIF9PDUovBrrzH
ulL/MPR5JCCfLXuWFbO3EO03tfa+q/8Kbbk29H2geT6CSrotdp7hy+HSXA5KLqneia9pkTX+Xfny
nws2t/5cN/7rg2lklhvlqPw0II8cxdSFlm60/5mWUjk4z8+P9j+k7PzK8govvhGnR9nkytJw9tYw
O8PvP7hcEa+mku5dX0bbtCjORhFKxzC2lv6vSRRVHE3JB6CQeODXw33UA3K+Z/08FJuF882HFc5J
hxrxrVCD1xcYw6wC7ZMPRu7VSf0CibiDOhEsboMhZzJbq5eYQ5uD1IOuR4xSIU/e+Ir+5SWTu26c
bp0bQqMFL08a6feG0iu1mMSSsfiXlLRQ3mJbdBYmtVh7IwBmTmtSaZ/bJbAFtmHXdxjLX9UQ+5ci
Pex65gbV/d2u1r4Xnsb54p71jr4Sgq5VMfSzfudIycreCxJUdfY/18PutBxrnairZxhzpmk4tLOt
+a/EFo+iQ0sMaN/XdcF6MDrc0bhaW4dVWiywmvSfZ85sPVnCtBhEKoguWZJhAa6e54W6U6qKF5Ju
Hd/qKgChluqBp1VnBawlDGu/bbbONxM7QoU102C7Vu8sFfAaFHnm4v1dGwAusQk0XOp1d69XICE3
tz7OjFxY2MAxs7/UAb0oBDy7eIRajKRXPCSTObQBuG2c03ONYIfBRbxy1swiPRhAS7lbwAxIsz3/
KVcHCOLu89TEl26+VCa63EMwEIvvcwcPZEGsqiINXT2cx4EMG4i/DpfUhuv2AD6l92jst5AwWfd1
NJBxf4iEnIpxJXxS1KCBr/XjSYLk8I5jNuroPp7UlfGBHMvkDe3EgwuEaTI4vgbzQMuFqMERo4Ob
q+/AJV0LdTfDJXIt6Vq/bN5Wl9T3qQbpV30Qnd/r9uU2pJwVq72IDEVSMjHZEMtvkOCwFrheVMCj
AanflSX1ehzsgqy3QMZfe8HsP9SyIzq3BrppvHCTZRQJiiuO/pl82grsYpWakeq8nYwgXE17Xhct
gGnUxMhpwclG/h0TQy5yT08aLPngK0QYKt5BiwAQOxmKCBelA8LobONHsbJnOuZMyyksaroFWXdC
p6/Yeh19r5Cha04TWoJ2VYlmkVKkYKcKhg37/RJKeitpWQL7ICZLzy9mMiz5JKnsAavbmSwtGBeY
N6TYeOx6tzBP/vg/goPZ1jcYEJ6r6ruPCsso1XrGRQ8WJSthOphhURMzufhbzX0eiGOpn+1G3cbB
xq06/cP20QOS/Qc7zPHmAK4X3A5Pp+8C9uDzHscG2H3furcvfzqRAKoFFC/5KFvQhTcdSIJHqDZg
A4oUX7d2PfzwmPwIkAAJqIv0Vz/7T+iSskxcRxMQ9Ie4NKIGrrbOcauXt8abnZjv0SaFYqVCrmtn
abAaJKVbYzpPqvNTvduQcQah40ZjqGfn/3KbA2zRoxX1tP/SthHKFC35UgSXpnyXSj8F5tOHJue9
j6ITSm0mEJ38RcucvCjQ7g6j3Cw1JB0RVh2Zo/CBaKktPiYoBoOidps+iWOLe4gHCGeoYTBZPXOI
y6wauhynQ8rzbmYEpxzuAPAeUaTE2zjOuL3yeVZUXTHQtICTsoellOiac7bz0YOSqyBzsPjk9R+D
7/cwlSrtr9xwqLwLCiPLqTeA0nQIxHrgZbUZB+W1dWE2J9o1vldhVcWz2JpMzUgF83GDOMtLFqxz
PJdVU32af5zE4jQNQVm73gAs3vuAD0GKx5nzwsghFa+gaTnhQ/qkmgIRTySYclFlKLb20MGFWHI0
Iu5gGQgEHOGO12W2l20SZlTNGjO3UO/VISTCI77lyxXQ9i5PAGVmkc6uHl8+ZeSHxo3isAxhIHnL
CwxpVz0BjQtRfQ8XkZkjVXwI0y8jrGhL7zp/s+2O3Xl4owcbAn7N368TAf2EmM/sCw3YoGBljQZF
so5W/oTNAJ5EPG3O8TmQzzgW22cmhW7hbyKBPsBlUp81pRnler/5A7jqi6itKf17asueiCONKuF7
ttLN33dU8vA5JvW/SxfisqOaLgt+8TzS3s4aX58NcX+o8l0sX6HZrJQ/oAgsNDjgKoHY8vPnwTeV
6NVWCFvInIKD1Eii5MwF3v/YVKQvYCg2tfCWx2jdC3iQwuJRKHvNci/+KFz+o2kGVwiukTL279UZ
lrsMoPVRC3SKCoJSA0hCMZtkr3XYcWWc8aePT2tdniVlXf7rgDhmR9rShic6Nt1c8iJw66E36dtl
7de6Hu0M5B9JNinmmmDjazCwkJKlzgZB7/sPVtdZJcWh2T0xqJSnDLd75G+fBClOiK+WCYfYN8IF
xCUMGEtvrAjC0SgD01MFKwJhgvhCBvx26m9+/WgUHt4ByW/MDZycxg94V7N6VW7hy8uXG9kr/eBu
v16iPtxZQRuZzpSclBSM7ViHx+Qc9GkEuhOw1LKd+WW+TRDHG9dBzEDQAXyVEmkVP3MWPMyY4NsK
EGb6SesFqO2sQGh/ed2cfSBMji8nSsegL78Dp6JUBYvc++dn/IqkaZ8JoMZ47RsfuuEqdMyJlWnj
3qN+wfmnJm1qOM3vSSN/9AhtDS2VQNp8pllzh6kV4mLRzwSoqsf1ecOC//8v/vizqmRoxv/ZYmTU
7cGWLrF6rXpmmYfpW8zfxX2CvYtRSRS060k0s05Y49Xo6gpO3uYpR5VqDR+T2OE2ljPhp02Bcs6V
IDjCurSHb/aJJ7ANZp4DgZbUZ6SNgVNlXBGcbhBRkPEB+7460LcVdXD45ZufQMGlmAyvrOkqGVS5
U/58FUpwTzE1Yd6zMtMra8n5OgNGbEhxWleVm9cGtfzU69ohgMuwtMoJeljFM4x8ElOBMrhqe5nB
LbpXIsH1NPBTQxllrIx+01nSJl3hMVJeTeWVI1K4BggjVFeZ7woVZOBGh6DA5lfIA5+CcmKQeQTx
IRgo99/BKWOeJaZ5u18lnnrZdI2YsfyKipAVYmD1ay0ciwrvSFbXNjVcPNoRXoTVJBkNQPfJaJSa
1iq3YN6mBqr5JXbNTLGCynaM16Y11yXhlTcaF8xnWl20R11R+Vb3Qeu3ZWmTzvbIrSoJrwZ0eSFx
web4UbTEUJboeotFq9cEkkEeGS7BSgMbho/bIiZt9C921lsm+3wWKWXmVPppnma3HEGD2GVCFwQu
/GV5wx/LD7hGSDjBEzqvgCJPQiFpQrB5foKEAD4RgLHzFFLkyL/Ndo9jFVidwc9R6U3ne032LcGg
jnDfv+Lm4kEFV8qeq1KU0A114bMC3zkBUYv221MGiVT4i1FVDAwJW4FqGXcmE6AREYVIF8c8DkQV
Fpfu1WtljPWHkB1b/TpwyV9JcZen5Vm1FKjsBo8YW9CQUmzqq3n3kQkz0ppinFbBue5ow/2zTNe8
PGRoWrctINOQb12xYeu9RwWW0bMmMZ/bUPZOovxL6ikaM42wRy/xzudYqhjcJkhlGB1u+A8XqREo
Xjhc5hC5aT1ifzaQhqKSB5FhZ54DDFJRWr7u0A1+nzT+qCSBbA6T4XIg3ZmIR7OGHB3NoNnuCT2U
uQg1qDUNpeMEUn1TbDH0cE4fuXafG2X3pPumbSmozzoc8TPipKZS9xW+0o5to48YtwU7FZPdcpt4
Ng1LwSGUPAF0pMdPCvPNO1jZMWiJ4p7pl5P4K2XXVEYzrBco1dPYiqjoi/ZMiKKKs+yJyOxMrBI0
0wyMjqkujeoBSZpc6bLsk1quAccZH2syUC5Boc9R9tOUpuwxBSvtS9A/hVJqyhYRsSXsbQLObXQd
NqE0hY2RQm4lE9juqpAFDUPbfKfTLIfOiH0R7l9G84twOQF/DeGIIpuvQDsYqSuGeBSQFNrYYbRa
qmF7pI5pBUtzIr5cpae3eVZzPH+GaYNsQKH1qDDPuyIeNXh6m0943vlhgUWTfFJj7Vkh1Pd8QHEN
lsh+NxFAICDN+0KbfHsY4XXlz6rbyGtLrWNe8aWsskg8TaCvK+jbHqAYc5KzFYxWmpiqo2NRndZT
ot6ThEgtt4tiodp35LkshSi6aM8VKroAVCXPXuHuXM+WiCJBCgSO/zE5EjCN42w91juT24vg14QH
B4aahy3u0tDXBi6dw3RuMMYoEwYC5QNv2fPfWhTBJOfx9pcXTyWl4ryaGTlFl0eFWw67shJkZ3VL
4MvQ4gkczlXNtcB42ucw1iCNJIvnrTk8VIPeRnnpdxVq9Mp/h72tN3WVJcrtVCp3a40wVOmZ7YWY
le4zJsDTWl6ote4UuIx3DD2eKiSMhJNd+WoIgY94Nqsr9i+SmQ8liXfAfNKJz6n0WK5ZRqGwpNnw
yRsVfhTNDdGx/1GQbK/Ibnbx59CP4STZnGHP5lnMrGYTYsoCq/hRUAnPkMpYBEbWyIzsmEHoMHUx
X29NIxv+9Hn1Sxkpxe7oxIg/gTmOK2XRP2X1SA3fNOYM/G/fcr774I95dc6FuAamxtqwfn3auLzU
kK0Y4wMkUKTWggOxHN6zuWD+luRjKYTH7j737GvJKIH3c/QgOpWgBSaxfFfogIlnWUMYabX4tevY
/CfDbYPKJ4WyzCl41y2LaJfGliGYVveWV/YM6qTDkb1R0mTNmiAUOSaiJWfWT56f4CIXCgT/5G0G
JALvJPCJBdUPVWkWxC4bUM39BlpDm5AoZSoJkUoPI6PphsRoLXm5xLofU5Xz2WYMirrW3mZzgpQd
krWSn5s8ZAhilDB94cwJJaBZTeGU2nRcaOD22tqRSnQwrXK80XuB6D3NlNdIDYtniBs8vZ+/2aF1
dpOxHEhFB1V3x/l1zIXUG1yCUW+VTnOdAijnX8q90c5oYVC57LTGSR6GphsCmf/8LMXqOJP1uG43
S4eTJwMQbi9k+Zz94A3oUCpFbVNhooKs8kY5ISc4/L6v33QqKho7WgSIEBKVx912XuYyPdyWGt+c
fOw0eIadP0a+nd3eA1GKyyR2jEVJ8Ei0mJPbsWLSzR6yo1CNlX7waKauqYyxxZ+7lNTHr6A/yDFI
Z8gyQTUAyontj7xsAhNRiXqKZW8jgQbwC01O3c6AKn5U9DLa2GogomXoycagK4cs0vK4g2fC1ZOo
wpOXBssaS6XMp83ohwaBWo1Rs5rJSb7Lf3shhGH97Ne32te4xTMfB/IBc5t32M2v4BfUelVKGs1m
9ECWPANZ9RlDPmEEO+4hBSxs1fvt18dgbTrBAW8JcTsjiRiXL7E4YTlLlCuDO12k+NXO0jbsa6qB
5xTybm1Skr81FVHX+3P5E/rL4gPLOlHe28guSqBihHlDAAI2Zu1BzkxMROegVTPOaJQW1CEt9it2
dVMtiS5m+2AusG92/shctQT28E4Lf/WxcDfao/7VnFB3lkK18uPH+r1o8E7ckYWm7w6oeE8c2qhZ
MNcdZ15UJ4rJdDJRLCbATIjFFUjwUHATZqak6qVjeGrAcneBH5SIBUeBmTwHhrxKE7rGV6sTn2rk
3bmbCtHjliSs85k2S26bSm2/G4jG+lnzJ4DdLIh1beYNlbaerPTvkvpP/wZGXAH0yJY3DHiTGYLk
/Ubm8FTGe2yG2EgVbG/As6Q2ZxruR2V8P5227Qq/ptskw3cQ4LqqWl1yRTRTzehG/PnXoYijxMRb
0XcIUyR974pJzEjpzI+xTz3Pg1Zx2WQG12R/EMhh5wHb+7u9mMYhMD3LGJSNzUwcO68hLT+zsg97
fezvbKMz6SpDALExSBXknllxtSfrkMmVPnO3Ll+dQ+Wb5IFF+MmUeBliGHTDLiu/jGd15znNN3rR
cGS3WknqqJTdUAZ/mzDu6JRvc5hNhqVZb6XwxyuXj0YJ3DUL8DTNv+RYbiafjGueVL8I4ArkEukf
+qYq1ITc2F87XLoejKYkmoDn4V9hsye0jVANjx5XUKGQIOGicWVD3rbDZji7bCuwUaowSBJk3aO7
TwQwN6Y+a4w13Y/7MyBjoxAswCSboyTCHOZ8Lrhg79mFhnQOlBW4Gy8aoWz320/3ys80dPnuoKlr
DxxC4yTPJJojFYHnZPEWpnLmJDV76iViDblfJ6sTKiyUtYcgXH5qc1Si+gH4uk+sSBnyvqHIUaU9
uo6Sz+mn1QZ+cfmPspA+w8Xn6U5ZdCAT4yMnFyS2/gre85Bcn//zZDV+NIDhC5e6GHV1Z6SPSoQm
CgULdxUwvX9I1XgcCqqLyvzzxCUXyPytyeOww6i2LCFVhqMHaXQGaYijP9ftZZvexy+YczSyfeyL
Ysp9eWIHb/MeckTb8gaLV/n5G94OTO/PAk2Kc6UhesECTm905EenxqcWyuImUtla0zMqKeJkNxWC
4kcFMnFsrQZnFqfgrnbl7QU5DnRQi5t7E7idkD3LUHUvrJsSQEY8yz5ruzwGcif+y8uJzDmamNGi
fMTevb6u3B9C83oXEghmOwBjwYLFwjv9NNBydgr9rAVHqMDA/5rB+OaG3NVv/T7QG3VFwCR82Nsv
a9J31viYsWfJSY1zjIvqItafKG0/SCz066OpwYfl1V16dcJ85knd8dxwRaDWUD+DZu7kUuuHAgkN
58DRIOBkgsmiBoMSSyal3bG0lrJTwnDVSUFiPE2UZI146DKqy8ctVplbUs+Q85rAt7DJOjCBXXnx
sQR0afQNqR/NeD4h6mxOHzKvQ68HzSd1KCu09rSwWM0aLomn4jWSoQoyedsojgH5myjjfeUzSG6s
+S4S6JkLvpopWdU7N+f93BGbVvlw+JfFrOijHB5+N6GqVJVADKsJX6J9KU4gZ/pN0RFf0axClqmL
U4XFxII0L8srSS/+nojlxPzjiZJOZ+f2F/dDZYmQUYplqco32IDhagC/B8zYIu0Ug0c2Dw+0lmo9
idvuAb5MQBgNzoGhSMyS2DIyojUAbzyEIsotgmU7ck0Jd4cWFue6Ok6fmDtb2Pf3oRItnE58OTG5
MpNx1s4kKZu38NoEmiGA3vFI8i8Kbb7K0LfUvsHeIq9DwvVuQ6EVJK59agqUgfb+GyW47BH1k/v9
ZaNaNFpFIxOEYRRIleKY71eOW/q8RH1OCUoj30uTAGXgjlI22cGirT2ZfQxNoZcoAMBT7VDChBEw
pALdxSd6J/GsJt97cE/qChRj09o31Y0yQafDMb/pTmCYcmw20q84m6EEHVh61wPjGcIZ1NDvF0Xr
7HNOLHRj+nbaYNJ7guYeoFR9HVY6FFVllehvBxBtV5hMtBb8uLxrRiT/V955jPbXaHCgzn0kREIu
7PBOT4nPwFNexb3bREVLeykhVd87gbhP9W4oE/CWkSmW22EfGu3u1AVF5Dz4QgK+s0karcf/KLSx
gaZLsBYf6fUdcSJIys89kh9m6cxjjDDkVZIu4hMNpI6k9FS/QUYuSDPDLWrrBcTsTiv8YPgn+uwz
oGTxts+2mvE+SSP89nKBglL0Q2SSryiJ94i/90n5gWpFlLngf9kNOVjgUzT6JKd1jHjtxlFhs1re
vuvbW7TCiahG8hiDbeAXVNnVznrRbjCW7DQOEprDrNkjupwS2tQc0eCCetWkiMI8qE+rpPPcLwoB
/ZBOoMnfPGvORtPsF7lNxeEcsuSSAOX5/bOVnBphEVl8tfNX84phkobmG3so6c5+r66ceGgd5iYp
YC+9lyKa03WYhQkREBO+LZGqHwtHCAk+a5FPKbZzFmW6xZYuYfLOZdSr5Eo9wDKqYDA5sFKzTOBY
yAbxRxD7g955tpJ4Og/STGWAFhSieWDYPvKuVC/q8yDW292NjUEFwPRj/rkj3f9ay3ctTTU8ACuD
s6E+6gdSFp0TahbFAAAaDArZDa9gOmwmKjGv+gwNT4xTiZJxTz48e8m7BdUGR3/6VwbBmc8lL8PV
3S4ACIoeqRr4YXvUcldkcZwWC/iUG6+UwPcHyWnkNagO+yCtkhbJrRisPfRV9orssXNxrB0fQ05f
mrPGozyg7AsZm3zW1UrhcwFgHpRnGf2+snrBTpqxk3/jmYGHh8rIzyNKcuI9o8NK0OxiNIRAE3dN
s8v9+E+Q/5tkuFcIglOu32Uoa6+W/cO269Nb6iNOHeIDJDpCHgjCWxUwbvT2H9dwIYLUZlA/gOHY
sGeAVBK/dXwF2/y8u597KH+QihpE71BJR8siUmRax19VC6KtUFVLkn+0FBFxVfTQF2BWRV6pEeU2
XlJEBS5Kex+0djJlQgqz7RBdHc9Hq71He0jaL42P3tbay7oUVBxQjk8AUwOGx9xgzoBg/yU4O6pS
OPWdhSle4s9ObE95QAxQAoY2mhxHqmmlCR8sy37A4oa5WD3F/RSvrRbT1+auf4QmShN+/NJXBONx
KAC3ezSwmLYqemJCI/px8+VPk45LnjOyHjOnHMK4e4dniW6IIdBXwkftQrs4NOWct66mB/qhDDqU
FdHTmQCuqLVnjWaw/iK+MWvpGE2IiMeFNeS5sNX6bo1g11p5e1TSe1nbYL3g+DMC0ekruo71pQux
ZyjS7VDaazWoIZT1NrDzSyKe/DqX2RScRRQywgAomJ8PAnu9MKnRUwXWSeuS9UkwDTJHyp0dnNxp
d5GIa8t1f5Qj5hrmYyn+fl1gEZTnqBoHH/XVk5gmz9rWac/KkiCZ9eHWh0BKoS5dYpmlQ9UCp7ql
NykOdfMqecXyUUO8PFry3APLCM1tZT4qvF6Ux0wAV1UjruQPMiYzY8U+RO336PmMMupQv61JxVw/
PBzyIWfr5pOwkrua6bsqQh92ZEHmq2l88dH5adJaQFETaTpjMDG2PFP/yLS8djNmVsG/V9n7lVZi
q0gwGVQ93rH2t2IAxd3Ad8L42mQ46YZkvVPQ/t7fqN5YoZ+xWt5YtXRIQtpV/qkhZ8/wKX4NJJ9l
Y5tFpWdvDpiOlQqpPhrnkud1MkNMRDgl+7bSTJ6xYc+8g9qqt6aLvjXB823litTUZPdOukf+HTxy
QWzGReXrLrNBVBF5dckRUXdVQcznhHqTDrjr61kNCP4izFvof4ivN47iJ0/gsAC1zXbDVElEpQi1
jYwW2a5BfMSBA8c5QbZpmCqWy+CSJtPvUpNYDGLjDJj54zu8vKADdMsR7HaEIE/EIL5kk+6/03A7
Dd943/rfkZrOEN+xwwdxgTQOJsEoyYW9MbjDTryPy4yDiVkW2+klu5nzD3Etp1t/PVGMsrIehK36
cCEZQ/qxQXnEOENcIr4Wzv/kpXI46KZt7SgfdOr6Fwo4k+Ua6z6AnRw/BH9fx29sBJy9OzDHM/kt
tVYHv1SlMAjstmzOL8YqCZq6AhMErWWXUvwgdbztBOK5HdB+Vb4T+nzaEDcpNpHvEKT/+rK7Tg92
O2o8noDN/mwBI9dEBYnW8PFQhoyJ00m3NMj/9CWfEbJMiFIL/71i9UbxkcYRGbbSyWKBgxCfPatJ
EZT1RMKyooU9w3BE1KuY6LKOgcEdwzRm+2E/+q7GfD3UNSpsi0PVfCJM8cMFkYDaZbNkNSedMCtS
2CvOU1Yui8f1EyMwcWkRspnp4u7WApfHvKNqRuDN8tNyd9P1HWHZS+0iWi/GtYu2an80PgkEniFp
TX7fwujwpah1MGtZkDBOnZvfctot5eOR5j+FHWmfLUXg0KMrg9AXE6d8/izMS/axi4IFs6MWe4IV
eV8LFYh4EfuJlYoUr8wrmLAQrg1q7hBmaEU9TXLv+7A/KlR/hWFOUKfQOmnBAxNnkR6Rt+GyIw62
Yvf49UNM1IbxZ1B2LqsKgFmqYWNKHZJ4MzaUdi/1Z9xE19cBN3vAn7eUs4HSr11kvxZHFjXZXEdH
Tp/fgr2Kn+iKfelreRe1S5O/YDpHEyXPYkpml1e7yCgyrG97eZ47qCVoaApD2wRiJ3kZ5B6stEfB
iC2MOBP8sfICOU4aNszRPG0dbCiGgB40pYFGjYYNVjU6IuCD/aIrKP/ofRMd+zisWf61dM4p0B2Z
Km4lXV8QuImAtuUZJynVmvJoYIoWUI0wPna2jYW/J2jghSG8kjJSB30xvHulYcL+Wl2UkQFJYOaN
euGOHAVhk7SEkIQXWTUurmV4f8KYBUaF2qBAc0e86RJLRhIL9YDXP9I9jVJ1dZW9dV3Wo/g07+KF
Vc9vbwVD6aUn9wrhiC0eX2sauTwWUjAtjud+9tiKcjdxgFmk3XGhj8AYb/tSjxjm+O32W2ZgCC3K
0N1isbe/w+Uqheku3iZ0ma0DnJiZ+oksXbT4AgsPTkfEQL+h53wXHOaJcH1FYt0aA4dITlOsK56r
bJDD3KNiR0UJ308/wa4gnutp7XndXeKk5ipvWSdjZTw2bfuuUJuz6o6QC7pwyhpjgq7KANoAtFkw
Yoqo5IkURDFSw1Xl612DUDgr0t4jIfSUycpHU5cP7qZlOyD90dyVI17E+6CrTF4KXokqESpPiuqX
vIGwpRpO1tk2EXUpv2sLMQcpiMwziQ3b/Pdz83JNtkwETrK3kiw3ilGaK7g0svBRs0LSa8DrS3Dp
Y0ZJs0LT+VpGgXO7YldrW5qKCLpwWf/6Wtb0bd1kgFKAzR8fFwPS32dDJCIepQO3aALRnCAK6XRo
lmFwiZoNzV+NuPFCpZMKoFmHoXMqUEzDeo8EFdbvIXBY8LIFL7wEaxbSbtvo76SsPtgwB3AvICWe
/Xs7Qz5k4v0Oy4DokxqLKfO+9ChExv+OIUF0qu80uEgB1W3PmIh0keE/jI3AEiEw4VNm4X46LmzI
PKySxK9MVcRhbaV3cBhJ/V3AvojfIUVt3WZ0oxFyCfuRptoBP0+l+YaJOHbH48C2x8D6mH/O5UU+
/QhZ/PVGfchfOFzXa7a+KTFbhZHM3/9jt8hM5wPiCzupTHkO0MtUpqbIZBEzHl/Q8cXdHEuVIm42
VZTLPJg/sQSuqM+WgVnbJclBGWqORUdTLsU2LhZze9v+mccw3CO05HkexH0ypTfOLCxoHfLEPXbC
H9Ey1VnG9UEhD2sbRyjjEiEb9DdC6VSz+n3aZs8jNxkQdSA3UJWEge9RpeosLKi7GiMaDfLt2ZKr
kP3W41n/rI9Nurkp7EYfUETULrt90j0K/vvpNs07rQp6Pk1QKU6zmHnoRveJNEdmyf8PjGkwCuV+
4vaPP8X1y1DG79qv/31IMqj605QtyorLrZ++3aEio68dgt3/bblBbOdq3DKnkvy5noAhJBsw1Ehz
DJ9mETqlJqUpSH0VDSgEfn6E7bkdkf7p0yyeN4qg0Z9JLs9yW0y+fl8lVv232FnCzFobWIq8nyHd
QHCBPSqn6bzs8tcz8WgGG4nExO4PfiamsdZIV6Af+DBHeQ1aBK/rl6C5MI18mweDl2TaE1bh9Nk3
mwHpzgxlbDQ0A1n3HMj9pxAYuUfUDoRkI9x8q3YAHYnp8iikFQhhdeJzm78BIQZiSjzDvXmzZyuD
bqj5dOW08rfwaAcknPX26WYjJ2WWtxF07EFmOCp2vUmGhcwp5aI7PFXsWBBTNZGHTXTBR38wjZhf
wTshRjDLWh8H/gNUgdfK79Zbwnv7DdVnU6j9tmnfpBnwZyzvW5wQ7gJ2sHea9p/Yv/ZY0dOJRjyS
RnusFdnq8LEm8T2qM/yF7pfigfQc3w2UPFAEYAhP8RzeTQ4MVxVhJbrdIfMP1iwI++ulyf1Q7/D/
yFJgeyQt+E26M9fq8zcqe7vWA90stEWpe3Fs/PLWM62UiQbDkxwVkIP/cPn1Su1Nn3CnfE5PHxds
7Nhn/DowfWY/e8veqXYSoXbwuG+7CBou5/Z1EPJLEXnUU+I+w0LlSbnXz0q5rTmB7xPqmokrx4D9
LKaUfzeQGfNaI0N2linl9qaZdAUx1ormWAzBWPmnM1AXQPK/l6fJPbe7q+DQ7aHbLxKyUaPC5m5l
zPCkRzqNJom9EcKDqxSrvxNlEIFCHbBHF1yi7qrGFlOYc1baYvNpfgrc87yKd085I+FISyRVJBgB
H4ryIqW93XCzMUxbnlJybrOS/Hgi1ptZP2UeT/Sd38Vf9M9lUZMrX2ee67IU2qAUhJf8F+peMatS
Bq0tA2ZptQYxjVdoWanFCFhRSmqW+d4SHHW9yX2l8r8k8rj9T/5i1KO4Phb6D1aB+HQhXOn2lhmr
77A3I9hlqudGwW+pML06pdTlWfU3/TaimVbwXfJouz03uuhV4Lf2VtLbIM56b+p8/pCtgpHJbLWC
gim896O44FhLosaIGhnhUl7kXEVbFGi5hrGhmb8U6+U69fpm6dRLSm3UITNXB2xO4hGpdDco/sh0
z9N2Y3r678vKgRfd/e0S6Ky2cYrCdTgRuxc68xfCMxVIa20PfIkok5ZnhRzEcWs1WgTgBVGrhv6A
hN3hQqsU/ZC3tRLZxHIbZVjYxuor8j6s/n3J3RTo8K+2SQ7oVvE1qj4QZy+jqDzr5/MTIBqIMr9B
lMS3TULWSOpYEVxu/d3OSYU0vnW8uI2wdFWKkZNRq11Nh5RrXpMHIW84PlYjNlKdlVkWVdskmty6
HZ0LqP61l+CJ7ncxZB0R881fSJVlxGrJcM3D/VtIy8PKNBdZvOw4mBoSWcMcqw6nSHaTXR135Hop
oekhM8AJKBBB34oP9MPZu3HRgX0gVmL1Hicyvh0KFOdiMdODQhBauI6PM+rn/IxukRXSvTR1nWt4
Ajf6cKf16Ios0Fa1mXjFpKot1lsBOsv7xjQaHCkAoqTZ8OtxqOT4KCqaJYbd+xovSBmOHomjay/1
2BbLuvs57F5BkTenTbpltWzkyhEl33EEB3bvKXJMBE3XRiAN1+jLtI84KCISRZKKgaPp9JlWbKLZ
YmNxpvbohAvkvq1UD8mRHh+7TbdlFQ4iilASp39a8ePdBLPIMMuz1UU49piACCbEGbSG2XRoaMtD
jKq31ZaqRJscWIfMT1mpK5iC1wqs2peztjU8J8L5ZK44zZlMxfHDZfm/3hEj1w4rJ3nfCnY6DXEH
fw7qbwaJ9/59mFrn7ld3kda0pJJ0Ugr7zZOXzKPFH2eZxeLniKjE+bHZffm2jVbn2jh2kdcgZqP4
zAwqsl3jljsF5H83CAoLZS4rhaPN15sMN7qXPn0sQjtUU83EHeqT5YUZaWlDoCMrFWrvyYlVHCn/
GyO77lJrh6kGH2gI/Hr/imAciNe30xPzJKRn17cfgZlkRcUkNvwqc0C6+ybqy6qOfvnqKtnZJjeh
cG1f2r+FNEZJdxvr5RNznLwhVA7YePoeS22NHL64jP8ANGkuxaQgAGpX7oQHSVSY1fP8xuBbOz73
FTwVRX6KAi9/Zx/jEJiOMKXS4uZsU8fUqqKnpe3FgDcvCRZFL8MeARKYJG7Jl9ECMNZCH1azTLXY
nl7OZZoZum7PzFC+FzcyYM3taT2928G8xmj4vvBKMHFHUVbqxyV4wXmJa5tiuM9Kfwm6yB+gjYU8
RgGzYG/KNF5eePkmtjyodvYOaqvInh+7710JIhOqNzTImagncXvW8TpPZTOr6yQNMl2xQSg4pkqt
DAyXJOMeYAuGMTZUQRBaHOwltl5+hcUyRA5QBcnkU+LTV3ILHHzhoFV2mRTcf1chKdc6arcNOh8j
1XxEkS8fkAJ9f1RqoSvwbXRxJZGSlWW1MBXw99P90O1dAKCcSNUVg7e8WJeqCQEgFK1sxrfwYQaD
2dxJCrwM3LNgaW8Nufzd6SS9Xw3dKXze8SmP4FXvamRNLh7NGLTiL2dJ3mW+CnbZCGrfcHe51igi
pKCJu4OFjlaOGT6xBLpj703C3Xjd6L3jahib+iYqfx2Y0stbjVr4oDgdhTcYmJFbZpUMak3aGN6e
d9e8HChi0mdz2GyVoclv46VAxt2+ZrX89ArKr4lAgbybcDL2B8+GW8PB6Ce3H3YhU4vy8g+4uUwu
2KA/5UL3Mya0cKAccVJLWsqnP6TTSzezBan7Lp6+3lQt72LRULrzeWtJbvLcAc6A9Flyl6iMV0Q/
33I7A+29fK041Z1idwbZQAMHfVwiraRTF1YGFo/PbLeI/cAKAg5Ly8oemkGYUr4/wZ+AHgINuzZ8
44ul3NOsitZvLv/FyblPaLldh4fkjyjFV58BWl7Fix44yhVp50+0sNE1nB/oxvBscj4IAG+fKp+W
MxpJZ33OzVxBq1Dqd8YOxn79Hg+S2qNptxECTR+Kl2BH52p/lIAKtlmCTRrE2aov4+gtgM3866GL
/9OCIm52kXAtMdGtZ8tIDRuhj2uY7MYcKxOumJnyrQPCokX/Oo6Bh35w6njgSzvTKJwgSj4jfqZI
7jD2mvIKfIN6NsdItZNaBcFoExwPDCEIWL4WZ6LhhPWkmCa5t3TjNkPTTYe+ohiB2xMgydbsQSNB
jXhlzSZlABN5ochchbj56bbKR7w/grJxJE8+LQyPtWSIjErPQwUutbH7YMZdRXjbHUtXC41e9Tnj
b5+Jfn8BnXy3Ni2bj/lY3XEjRyMCRuF7ahy1hQfXs721nWe8HIrSlciJ0975VtSZqwhriMph8I7D
iim0+pMSCN1gIk3bQc5akx1gefmwSTn0EWgEUfStiJDmlkvc6RnkhBXetv5VdhBnFTYl2r5qb5RG
rtqCDE+DA0KbSqeJFrhZxynZXNjrfHPI5s/difPrC/FKjOhmBuaurrho2WwBdUlFZyM5THEGjDqq
qbyzSE4/MfMhfqHZsambCyZT/J1oQ1wcmvKeohQNLVwy2FIaGLaDkU4ATFEwf8Vgz3EXWO4KwBP6
JRVSV9F0drDkJyTKzMxUz6YB7cUquYPU3ErlsNibfJvz+h/Lz03o92Ryo/fhZ4BA8Q7eeaV8YUqF
UlD9/CJ7cmfm7Q75nIW4SmR9gDXoGJiQiyMk0KTJ1xQyeQYEcaUBGthAHGI4rYJfxxqyi8+A3N+A
ff5eoDKlHC+hvQlU9zv2gf+UbO6IYqUauMabYdg7cf0Zr2VJmLdlavT2WepE0cZK4u+6To3iONnA
Sr9tYLoQLigRrx4xOq0OO6SnbUorArt6ejrUblozlrbfmFDopSshccH0Rx3S6AT6W90T7EF5gEWo
NT4XuRlUeY2VDb/dCQUXnjXSuPQ1s/NZI4i0RWPmBisNfea6o68SOX7i7ol3rtpCoyVDVNrlJB/t
ZCJZ1U52pkfgP3IEFUBvw3EwXiIHasv2VZYDxIi3SJBNMDGo0WvmILNRQWqgqTFcWFvp69rBYz7j
kv/+V5IF4cCpJdiy3jDcPUSk2im5KDCbYhVEdf6WIB173UZWf1e2aahJ4u+CDtdJ6xjBZgjfUVHH
6qT9piXX7+9xbek2gj6uqckz1K1YtIqukGMc5euNy6Kri3Ma005vPmAt2PhNBpgj47HK8jH04lLy
ZzMKrBz59v5b1TJHZUnp655ukvs2wqxTdgPuKB4phvPTPqRH/rd4bjlppH1Bva3tdGiXXQTVqTFN
l3ZlCGXO/Q1pZWI+ciMojokA8mafKKo0Wqkset+KORFRGVSMAdLjl0Sr/+NpBCCDX+GdnUiL4hna
I4lWHRG0cySio+hkAlf1AN8f5Ag7DCXQ1c/fr5fS/LkEMBZLEybiEtGiW+LzmIQ2jzUHmZ7u66O+
PCeC6XMpzeVnJKccm+sjKsAXOme1YnLifjWLYtoMZYy4fNsqXXJIvxyUZN/mvyEKcEsmLaAreGg3
Z+nRxcZqMDKZB1nheApCTziSVMkTiQLa+3Gzu2SxhYPQKt2DkrGTKuwupwgiy/LNVQKFYqiU6oq7
yCIa1zJd3E3aLolVtAPQ4GS21rug6d0IaW7LELmBNXWTc/cXy59Jd49EDUqInuIQufLOfypmHS2J
9ViDq8hZG0n8pRlWeW+MfgsBQnp9NjBgtFWhASFZUv3cbZqUCfUSup/J2Ho3wjQpWlm1F0gd74Et
NVzt7VKeOK7bCmP35MblGXzgPen3CBgR4J2eYazKQsqUSUyA7HNP31+1gFWIeCBzho1UuH7d7wwB
2HUnDnn5z3XZkYqwem0Mnae4N2/DUzrkmxwUtK1KpdRN8Qu4d9eY4yZIg3ss6mRN9ngNvN7xqmlJ
/nvaWNbdqTpLzG1lbhmvYUQqES7MYlyj+OJVBh6frxc5/+QW3KXnKFqz29lmD/E2wv2C3QNQo8RJ
QCC8hzGyKwjdO/DjOAG7Z8oa0Mlo6C2W74i7g8XQ+/pd2+OaROqVZAytjs27+KLSFHnFRcUVTE6V
iJK5aLAlH9iiF+Z2SP1GxIXMtM6vgOOgk3uIZZmbEfMOcVKHUvw8SbgKxhOHuUoaQIEhjr38EXa+
sFmtZ+yVzp3JelRQRV+Okhw+BacAw+Avp2QdF/lJklC5cCdF5WaUvInxRc8ulZjD+SJPAzAgNKBS
sGbxWUXPAO7BOlpn1Uj+tTUauhusyAtNl3cZun9OBshC4alp1dCUzlc1Ul4DVm7jS8XFK7qx+niE
nhtGgNI+TulLnJOJj4kWs5/vwUqWRqtDttsDb6OBZHBLfDQcksy4SxDHklbbC1KcWo5wPcHh5epB
+0chaRzG/sE4TN72LToSNv/sx8kSvVKWe0dKnCgK0FjN1FIrOvvxVmNoJJbxoxrjXsJJmNu0Tomc
Pnj0bFRpcDb7d5hdkJW+Yjad+TGVCPptNFauX/+xgmF/h4GPEx4u82DJymlbHbc2S0do5rJ4Oym2
sx7d7wNBSLDv3Gez1aKWmVS1EklnbggUjTdGaz68f2bssisZ76X51N3XokG4QrRFlqkcBkFGm2lm
WXyKd8C34W2Cu2dVsPmmXuH9l0WA8qlsvc6SCikcnkJa6OZdnAI8eqqT5YmqsfCIJa6FiFc9pSLY
e8VYPLbmnfFj/ORnEUE3zfmEgk6wcIGEKvow2kf9M+kw1nLaasilkR0m9ijBKPw02O9kaxJRh/nW
WIKOAd4T7ZNS2lL4TFAUMO5g1vfAvTMNWXMU4MpmYJfzfFhm6WLI7swCw5PfCbF+nCNmWEO+mVep
u5Q4GP7vx/BcpZScGN5XNaLFs2LEumQcMvxGIWlRGxrkEmtAG+gqMA7gu2224dn3m1wbPW3wlKVo
c8PtcaZCuM2KSIpdOtYJEu73w1a9xnwWT0jqrySEclzr+t4Gav9bREecbam5G6RIRZs4UMGLC6wP
XT5G0psRE3cT3Y9hBoMGWoFJEQRqEeE+s3bdL90ENpBAxrhhZQcl/7UxKM3JS6WPr2wlFS95+Ze6
U5TAOIdiYC4Pa/cEJOVMBH7e25n8+CoaFzAFlbDOwkzCVz2hoVydT5jJ8xwL9AGyNOi+FIcAubFF
DmSJuHbNUa35ehdmN2x1KZx0plaAki9SZ0BX5qKfzax5/4lLZQObYapwjj9H4xmPUPvdt62lHVvU
6WydnOpDhqI1GiFO0FDxXQliXECwnShPm+wjsFZfywgmYWiyRNUuI3OhyqVeb7r43hJ92PYJYNGC
JNwypJvEqU3q57WyYF0zpM57G/UV6depI42Xwgsf3DsXxOdOvPE9IXRlUtN4m64dexgW/yTUc3mx
lPYwRD+vqLA78ji5MZ53IHoDkHnSfgVcDxT4jnx3UOS8aZFAeLwRROj4fmSdwp7H5lvnwQWtIpWu
nwd5e8X1TxuXOP678NUbjCbfmPSZTF1sje0OYzPb/e1u8rYrhwyhD76NHQCQuezedNXkQ9DaVZ1f
OMC+QfGr6esbd8Ur+hIMIsqWetio9CxNvxUIlraG5tG5aVaFwio03PcBy/CtYMDACqwZq6026+Yj
zWNT+xGyTGjt4sZg+w0Itefzk5nmr/xM5OphUB76UgddDw2GY80qe15qmq1bvGE5n/vD6UF0gTeC
bD9JRrzwje78fZCxKR+efD5JmQUbGJ8iq/l1Zw1JdSXwiIdSLedui1kSYrfQUL4DdIJrKhvRUbhu
HUcxuyuJSxnI/3c8xEzYjDHjApeoc9sBMVeLgl5Z96eEcUIABgbz3YQ10VqY7Fk4y2J4drgheiJv
k8Hl98k9K7WR/gKRpyhedRD14o78W0/RrcWlflsKjQe0N4o+5vVKOv786oHzXJPZCgMa/p5i06XE
4wZRcKE/LWQE/El+1ycroHvVUir0B/BTQkFyJwXSCw91orjz2SxRU7RBd3ekG8eYxOAxXN0Xf/Re
VyDcIxOD602yq77sGVls6VQzOJBmqDh+JGQ+h09NXiCyKoJac/rpravvmP8mv6kQ0W/6NDpZy1rw
Kem0zy0JXDe/2zLwGEAJUBSWK7+nAPFOajgYRdB9PONPrid64iW7vMYsqt6lcAEiEPumNMVGn0DF
Vd7we+/+e/tEFex7i1VRlMQwHaj42Rc7GnFqQG2gzZSzK70Wfb0rZqof02+FVGPVfhTN5iEUOf6D
lVXDBC1wx0+2BbWnA+dHydUAvp7izrN00Hu30B54BE9RInkFUetSperuazWeQbqtRCihm9CQboLj
E5u0BrBbieHbESV+nImZCXrboWA+8EzHtmxeHMz8lpFyXsMCzxAp92h/vJIKgaYTEcsIxz9jafs0
aLoWUiAxxCeivq60GGzt6CT+120owbVUgwhRjl7GYV7PJ70L715byuvdX0GXdS29l48h+tif0GjF
GT0G+woOz0edtPhVSmT1AnWnDfaT4qRWzWi2dNwsvHfC7ZzvYN4OpflyXIc6NchN7eJUkpUZu7C3
VHZCo1orO+HFV/3c5Kv02LpVb1XnCOrkO7fBSbe0ppxKOGionGBc4SiwyC0iMOUHzo3XpppI+6VU
zE8LtGcrjSxRrwtZd5WGHKMrL/5H2WwnwUR259fQziBhWlCBDiaPcZAPig4Nft3BIvM9gNetdVuu
fYj7fmn/iqkcdNdtxHaxsBHmGq70hIJSoSkyzrj10/T78NjXNYs6GTfJq8PHpEwvtJxMM/r1MQTj
mcNrSmC2Y5PDVuQDCeBIQG0rCxw+eseNuaovxNw1236nJDaxZFerm5l5QsLmwe7NIRc1DybRvtJS
3IoFN7WW64RBOWM2oQ5QoN6KFYFqKLm9PBtSvv9u22Uo6BFpt25GrPBhN45+6UjgLDY07sJ8gj/d
mmWcbkP1nI/+S0jRUDdWuWXOhB2r8BalHb1uuoPwPP34/PDOm1kNWhaoI8aAZ4BgEn9NWHHDo915
SFaZZagG7FmG4093pFnfJee/nw2jrtawOndr1zMj0jwnqcPl5tVWUtI9XvirUDBulo93p1whpA/g
0VP0eiCwraLXTTcC8yfJjh5IU2VhrZMeNKZJT/8YjaF2svkKvGjGiZ6NRl8Q0UC44JeTuXaTqsne
8EciK+l6f201hr9V4Fq+p16fI4yRFt+zCdHGPFaQ7VdBIZl5z9OCiCwTy8Y6k8V2OxZaCHQCzATv
SsIB/EGbljdSjyzKg6oK9XtrBKJpz42f0Wqf9+kH7AZ8FGCxoETlOnMxz0Q3h+H23wc+8BX4sUj/
XGqJ/i2Hop5yVWrOzOjQ70/5Il5++58y1SMxsEarnye2HX27pontqbCg5zTB/NXDXFtqBWuwRsvK
CDSBoJxwxoE6X+jH+uR62s+m4fP5eaRHbMkKg1142yYOyOEtVYFCU5k3sNnF5NNOqjiKfQTVhOJE
bqYrGMHjgVDqgGapmwgL8jAM2igPIuRradwH8cIfB9Uumw94zGN7I1Tw9KhoXbwt/tb3HZ84uJrH
bJRMy/VN6/99YnCsIUwONsrH2faX7ZsdbChx3OqltZXyGi8qJEVZ7nVDcDsUmF52Opf0yFSa4wRc
/gNaUMDUzCJ8UQflSl0YD4QC2OtdBVdZQGocrnLoKxiyz1hNQtl5slbBayChfjLP6j5BwlkVLzyL
3PJf6bl34CRTAW115jdGpUg/AihUBcnNfxBdyENm47KTXzdKA3AKkI0u7O3+IRD1vGwBMjX0Grf7
XwkHR9jm+elLLMj82Z2SgY7PDsS+a+FcHDOtlr8OPA275FifLxZWkFs6Hr5KltoBj1m2mkOsBM2w
5UbI4dVgdQYgOZKNOZ9jtDcsoMR5SnRuuquKmm4xm39QZEntCPUA5JWnzx/nWgjPqrOPZBeT4BZd
PN9N/9uw8YNN3kCddTWtFyzquEFUL9dlPZ3OT4cX2zJqI2B8k9OUA0K0uXU7+mgPdrm3ZUzqCsP8
+tROkEX8a9NcXxXtwg7VYzNfatYWXvuZ773XTzBzwXaTUDHoIeJLP28Qd8Ezi5Hr1zcAOjNEMCNa
VxfGFSc7noRKtl1EpJCt4ivVON2PzCmvx9BH42COrq+BwJSz3tcHLvTxk4av1EzEKt5lpAymt2xs
x1rgJay41PN+YheIyrx2Ee3oQRrtvToOj5+r60CozTc8nyHV5u5MhutQgtifjDy4NmcosFH1tF54
5Z/yqfzIylGtZ7QmaTo+tcUb/9VFucG5ql0Ppqz5torihRs44u6jDw6hfAiBq2QHBdf9h/yYYJn+
JqSZxGtTqQnbQvWO/pp+i70kMPCHbQMmR0sDpFWgV8NHTEkHg4xpNJnun+4aebs7EOKFrVmrsvAg
ADZN417s5izwPeKaDo8Wp37X6FY626VndVpVuQNS8hbZRHFK4cFSXpUIvdHg1OskNhRJ5RNTrQjq
UIMGzxoMkdoF9/alOaeEI+5nAObo7oDg5gqoVcNDiT+2RAigATSQk1VrobOhEXlBPlA/xzO7IuV6
niuiYOLizuek9rVtvmqUbnpvPAV4KNWjye8L73aNBbotTD0wsDP9B+6ZkMYHWeoP9xaJTAHAUdji
GCc8+/1vkjzvZ4jSf2YvNTLtyzS/1QqLxf5cukhaTZvPQa5Y/XW2VbzMK7kIuABRcus7f7V4uliG
ViqbVUt/SrE2FZIPwNbdRu+KiqiSTXpxITy5sakuzAZoaR6+0frLoGeiQhYWvVFWw/HLAZyyL6TY
JinPOpb87zwBclComKYxUzufAdunQIdp78kiilwIbLgJJfBv9Tk/0cOZRjVCLG4C7vF1AYB8bJcs
PBKh2htVI+OuXO+jzE0UD8iTVpHwnlDXYuwtx7wiKneab/9dAz06fGlUqBjTeeGucc7scqu3I8LH
Wf5tNe9qOl5gWm2ho58DShKKWHG6q+O5fr7g8edmjyFTEbMnVsJ+pef4Hy9HSlSBHgpolpQIGjzM
ZULbUBILmx4SL6ZQStopmDjLcRyMAb6R9Ee5gUH8xakdG1lcl7JbIK3DCNru/jRyzXg6W4qUO/0w
7f0QG66fas9Nrxvb30wpIbF9AjHodjTEg7TlB/p4GCTwxXCQpScd78PTcbF0gV+4+16ADTGpbWS9
EpSieUVf+UMAlIpwg4Jkt81yLFIlmyVZthsP8juMn9cjvHF2M8F/TeSIFdwpWjz6Yz4w8S/YMIT6
w0y688X2QD3n09YAUyIioprzO3IWOo3CYYHmhINFE32gNI3UKiFYGn6VoFxGWzX9Bxok8zCSojlN
EGNDOeHJ2a+elA0wD5ta4iKikeTd3j+X4s+xyhaVf4RuCo3SKuw4iQuFa7IvbsQhbDmiDzzFBZix
tSUdeqdfLtl1yasyNG3KUy4gTlgrdjCxVLG241diblkgVKdHmrMBLeOEo2oHQ+T7HpdgxCymjL/b
MtD8n7KsbGT3WlRMCob0EGHR40setS1xcppfTfoaD+RF7hsibPnFY1pjcNGIM66/g6MzWoZbgjAM
aIAUO9S3ywWgk0D24lNCiWdEz4cvN0MA17YjQHIF8eYM74fvEoZq2U4eA4j38temblQ+nBSNpCLD
NuzSav50hf2fMjpdobbGVZfSFx0ldEppJ35C21WYKjso2nPphFHKLPdxmy6w6WvnbENt38L5LxaZ
O1AJnKeMAKQKn+x75PBpKnQ0HgpO2rBiyYsyRWayLFkcpxOiZ8Rah+jsKERW7MFEg9Djf0bT8P3I
Q7JXUzGJeO5W6WTPqihEM6qvsxTRfpVsc/6XVVOSvPr5D7WUPF6YkSit0kycZE8sRvApm6K2RlCf
Yei8QFpC89erbII9tnviwGyafxNk3PeRyGJVvhTGE8z5+iW0TJs/M/6EGZ6chiG0Gio21NvsnUO0
1cJfn5pdlZe+Vykj1o7WVDxgoYeHZnSN0k8gj/FJQNVAs1BBk3pJUkCxJXuS7s6tg9AgozWNoYbj
9OflXCI9KgCL2/pI8rPHo84LV5ly0HtI0olAJOdUTYEw6al79R4dMMiGXCeRI5MNi71pihNq0F8z
FATFXyEZDHQ3Wel8xbTHZke33tmLWn86piSbLdHsALwpR7vihOnt+EW4zqnWXYf8YcbT6ggYgYFC
aFC1dRcxgq64wpoUCIjLwuGZftN6+skDqdPAG1v83plRQV+J5tS8E5X1pw7r59kB6OpiIyY4Q/iH
OkJ8SgdA2JBhZfMC3RVFj7hOr6Z8C6zxXSfYTyhmqekAVumvoR9LeLeWHlDIQjowfrXQ3MzrTCC1
gfwHttaz0eepg8d/5s3ab0e26yc8iLrqYLDCx92NBVUJ6Ss5/xpFgfg3VTbyk6MwCX4xzzM1a2pk
hvaf6LJoh3TE3RrwkVqtcSiNbTWQ+lqCWlKZzU+fW8nznkN+8M0W75ZHPPXdyok2f1U48l+SA8hQ
JXA5xqSmmy+6oDeY9ZowY5wQxPpFbSjrSSdYTuziTJc4l2CfkikhX86sqAXlVDgFOPqxgCLMCgLV
6zQrZWE8DYgaoMUY6nfmNznaoR7fNht1bSAhKJBA15+Znj8EdD38lKmFnhae/nOG7dNrO5SKjiQu
NCKCdqZiWyQlidQc0Akp1zEdWkY2G+d4rJ+wOhrO8gqf1yoachUJ0zgCZv+PtB8sA3mJA7VPxU9K
2/ueFFOLxIWoKFvclTiYBFmP14mQ8Zlx8vXSP6t7w9Mzo1AGMTTqyj3R9v/zn/6u1p5H+w2zKJNz
8JrhCYMpA0XVrhIzoUKFfSXN50FYQwDmmnh+HCKK339HRcOFMsP5HwkQrzK5oxTb6XWqX9HtwgTM
LlRJqXTHddeudjlcKWHDPQ4xd2gj/p6qxaNouPjgZPfSMiHZMiU/0WD97X8A9jiLU6li7OLqzema
wor2fwCvbylv6/ycUEEeMSvsimnkBIHkvP/t7HmlHVZigJXnxveY9HihkuOWZB5r23QRnI4omITh
RZ08tz/Zm6DzsQZ6tOSAWvXvjGcHKmscxsoAzKaNpN8ep5yEXC/pXRp/g/FeFO2zaSAMpycMOe9e
SCjLFPOTuk+fwRICKd/kB5PHrXcTluMUVwbdFF3M2lABbnePv4dbS3glRxuvS9PGbFB/eMwcUFK1
1oo/yvEbVo9zARgGubTNKdcZ7yPRP7u0YlPaWBcVM2x8Iholk5Y5JOMa6vTtdqj0VWNqYB6kfGKl
ApJ1j6Y6Me+fKvIyYJDCSyzl/I9N/Bqh9MsSqa455exwBLRQILD2kzQ1pCZPN2iGP/7UGYGhr08X
oCGZXe5ekTxWI6UnsU2AVMsb4b/dlsWZufBUkjpGZOL+IAxOXYI8281LcJhrSoF4KS+4vWESRH0n
ORPAgO7TdkC/fkxVhnY9a3g30a0HNuHl+eJJlpkFYSoyZM2tsmLpomnSQPJmdr0oOYf7URGAcC0M
yAGlrAmC9WdNOtegEE6FPrNMlJ+1zbVevQ1bxcsGJP5/z4amqSrFKfbGDqnU1Mcpr8g+lWecujMQ
Yqd7ag1GC2znJjiTgSaSuuU2qTbcQFVEGzsJjdDteHVtBAAdApSfnZDXa6U1DGFIhPmbAXNq5ipS
Yt65bBjZjLepdGJQOpFdIo2diCLy79mp5IVOpn04V+w258Xa1pdZF8bHnls4yscVED1rXPAz2U0i
AzzuI42d/791k4MlbujR4NUxjGuY69zVmbTHU8t6OxPhsiD+K5X9L9YtGGfeouGT8+fIhyUWkZE0
RSyjlkh0o+GiUGR057Rak1krwfdy9FVH7uoFtlbbcgKEMHyr6Re7/kyKNnhWpr3/UU21VP9tiIlJ
P8dYXSaAMclw8udRhmDLjda/Gi85/5HYsZjQ7YtuFJdRebcdL37D4r4vaurzPwbRL/QFGs4SpDun
rPeBpbv6cjh8S7ug2tagDRFPHMaUgC7SxiiWI1aZJ1FRpeWyVuh46gQUIUS5bEU9aRSX3tUTInYw
2XoHSs/wvOng6gxFpKLSmPAffElR5ojX/AVVv9Ye5BCxqK40BwTkMJUrf2XE5zBCgG5bK8OWOGN7
1ku69BJ5Wz8y63E7G+k//BIHgsAYVlrPhOOYFG61Jqhx9HSIxiNKnHdE+SZpHkOxH8QvtbM77HJA
gcy2lQMi6N0Jt7nxPUv88kR25RacjebAPWu3QWq81vXUF++cOI6K8wdq2wtzIDQcI63P80j2Iimg
QcZKRCcNpMEIyuDdh3uNOSc6pCVcNgil5Fq3oPCp1sYXtkII7OaZTg0jvd8LaGeVP0g84qz/GE6b
xvVwI95HUCiPDOmwdbzRk1gOpntssM1iM3l3YZghwAhP52DaSE1TCxLWErACrajp98rAc3Wd1N3C
iGomuGqiAJDjQNMEbSjqoPlJycu+hGdrNPz1hyPTkoynLEB2pkSn2ULjkhcQlD1f0eHBThG7gvha
YYpl6fz5X7hvL/TWobIiUAvcId0Jptklr8onedFRaT/xdXWmBkS/HTUfqD8oc7FtbwbSW82Y3C3x
e2tj/R47lalcw4y9umYamNwxgQZQPzjX370S7OMLUGzIGrfauKnJveyfr/W7QsLVkGkj914woKen
5IX47vIh9ScwMMg9BMwCmdBME+6N0xoPdwhJMqQBVqBmNFl/DDPnNkek0Ki5tW2fBi+ja8e/ITjp
FeEID7n3B9dlrdzFmvqkm0CFKbWbYvvk1XmVM5Q4eD1uR9GCwQnOWgKa2kq+77MaHxZnL1c902zT
y/OvXAwVpMiBwsz6DhS6CNIdCW0TOmJu7xweO9FIDNc0dKYxQFkUofBW4g0JhC6wN5lfuAYq/owg
H9ckuL3jfgWkClX6bceiJ5nFo7B082/klr2+vFSZHAYylMKmuHFYlPt2oql57XwdDkANq6c19JhX
CNOfHbOo+Dk6befmjgs87aR1ZFFDg7mo1mogWuoMDjA91N/p8dI3B9uN/eMFv2ROXBn82tlbFSS5
ESjZdN03n+9CLyM92W1eSNFBVDubhndXX5BeAjk1pYUApIYraATlFEwYNPqCxMW3jzCD3o/XlVHw
tT9WD/TtR225P8cjN48+WVeXTiOubI6yKvpuNfWW/B3hM07nk99XO2j4oY1HzZZZaSd2HxuGw17E
IsMopRI4/yGHSaD+aWcqv3fL6zTh1vmEOM57lAhz7hMW55kNgUvts9o18O9Qwt8T26Hro3Fzje6n
Kkx49nmA1I0jxZKpFB4aSonjVnj72QMGym4HE7k+rLO13SkllYi6rQUFJF12kMYS9Ux1IyhGoU7F
dy7YokFQjPzWcCz3LAiw8msgHhT+zmFMT9MIkE79HLwibWB9e2Plh6Kf/WHJblo2al9wOkMzu8ga
1RE/3LohbLwU+j0bMaV7Ad8WqHdPHjS10MRbvaIz3KOpID5uCFfObmykZ/is1+KUNuBXDcv1j7A1
Jcwgxj+reIGo+8G98dsFtcb7KPLf0dp+GSsu7Ja+5KFWhjQ0ngI/sjSKbGNq2DEqqXX9CuXTzRL7
VVut4EhC6nighnl++/hfZTFofaPYCeaeqWpjtYFhgm2leSWJF4Wrh57w9W3kPUrUeKU9q3249gdV
hysqQD/dO7AgghjgppU0CiEpecfVzsKHbDR6u5VUh15bWVq5sFeT1nwfbNj7OYBsB9lMRyV7mJ24
9EIthsA4jkIdFFb3YRNbU38DxC4N/liOVXJPfkd9Z0E10iTzBQBtXlxs6R6X2+3Usyw5adbzPj7Y
4Su71H3530KzLEt3tDVVDw61E9z2MHqmMqx7AIR1rFp2ZB0CGdir8Tgq//4dKEYHNqmI2CKU+cE0
eVeTRjWoeyZDbbpmRSRjZ9+rjr+Bxe/riq4KtnaZkwmJe9PfROJPOjgdYxytugvjqs8ITvHYcybf
bvRzcDWLh2JGw04PIsWXv7FeFQqOE8M5iJ9HrtN9zp+inNvmGobCvZlT+VSoxBcgLdLAXku/pLUV
b/neRXuc+vfpKelMXkpkrhXvPzM7uPf8A80h7E8f/hVxjJXPlVwFAzk0EGwoAJyn54ubrfnM0Yqv
vq/OcRfR7qfAJVJbFWBX0yEHFiwn7XX/rUDyUiiLCi9hVjU5WdkGFroAIasDz4sg5qH4j+rrwDaT
Xh+qXEJhnxssg6m0kG1CRWXxkFYQt6ZkjItfVmIYU3/DG/eAY0H79foctqJxLrOhd2L4iQwVFGch
B5Dv2HeigUOSnJHMFJKKzMtnwX8LoQMlw6wAqCCpk40t2MKCQVwJnynoemMR84FS8VGc2ZSQBpCQ
gepMIQTbka5OG67s3ZiSdfBhoZNWOYxQuIeBRDwr5qv9FamyITziWXY5e1bOuvQaeQWR0vjESc5K
01hxhSZ11tgapdiWSPabLZxwXefCJsk7Ln08D2bZL+bcapjsCCl33gah04nh5MYWmeq0sq4YxDkP
uRgAy9to3gLJmj9VEO1pKkvPCFoYTaKhU8x7KTnauS2w6sdAeMNk3QuHfwt+6mYsNYQFxo4AjJn6
xn10sR5QcZHl6IN03KiQ0ldEnujEuZ//0MYK/lv23zbbKisW4C88JYSHD0FJsEycX1JnapvNXOBb
6BV051QI9YxgVH+0y73Sbrcz5JTw7gEKVjHFFXsDGdJtgA4QZzv1F0wS+oC49alPAEBsD76StMsE
2QH3WOudH2TNU3Q/8U5wlv+DLFA+If16BYv1YgqCic459V163JZULptrl6aN2nLFaA5Mc49Nhxze
SNt71gSFfq1ZnDHW3GGiV40J9k1/j4WYUNjdYJt7sCUluqLjpX3YtzpoVFGvptSfCZm9lSyfsDMH
NqYwF7HQpQaw0ldHv2rDVeGbKJSGVvtmQ85RyJBEc8VumGei8DwbaK23oFlw5xuj4rrdChs29AsT
n6FrgZywNqE/wrHU8PsjLTQ0JIATFXaHJLgdjdjwvZb9Q6l1xvipq8zpDsrEHFPDh++048+JnjWi
usOIjF8oRDjvp/EnRk9apCoa6Y3zhBxumj3JJeIM9UU7krgeopnUzZoI3E5AMuNdlwAsdZXb1Nts
ofNFVn2EXK/h8kP1AWdW31UwB7/45LIJBRB4gvG9OZaZWZrDBb7jcBP5lmN/wgJ5y7u0FX5lnXRd
nYb3xX2VFkOtEsWR4U9rIyT+BOULn2bTatgoJYoWEC5JL41vBDMyyJBtg3o4F8xTOQOWTtXRzAzS
zkCuXdOc3h8MtjdexsqZtNfS8O26oiBwpAS5Ndi6+AYiNoR52NMGle9s34A5aMyBFo36Lx21mtD2
IqqTSlIWkf/EJkwYjuIGn6O6y5ov3XXN8Ark9+O9GAT2rB9phVza2UEQHIIZnSdCQyq1C9HYFX7y
kR40wwkhk/e2jms5WbNuOAObjB7/Smx98Hud0ix7c+xjsdhfbsS6P+6VaHch7A3JpFCqAYUzAkMe
/KDNNjyZry6u+lKRMYuDmnoxx08Ieau/FUbiFkLzsgTQ4k5RuiKz0rVhjsXNyjJjeQKw0MB/iJ94
t2IoJxo3WKil2+eZ040mpnjX/dQTaYXnZ98ZY9bKmvZzb5cIdE6+vOXHGAZWiu8+xPazgZbtPvDN
0jPic/leZStRqTjKOK2a4iKnFgX89WjsMboZCt/jVz9lp57gehZlPuqXTV0v38c1rIMxcAYcEZcA
xpsAoAHxoA3wdn6Yq7nl7vfm7tV2I99hqgFu2Gb1+LOcneN5LM3qq6EsZy2a+YI9RC7QdggWS5IN
7e+U+gOAA7t6OQGLsCrWzq2H/naC2flB0kU/X6MO1LZJ6sWX7pP8I7JJ9FW9729lS62+qxCNRdMW
R7AB3JWR7xx613lSo5/jwA3/bMFiDZIukRw/ATY5RVHdvFTgeC8F7e6xTdhaNAqazV+4D0pqKS/A
hpCe6VxLhJ6eTIb3fTAzqn5k0IQRhFNQT7LbjHwCXkOVlxCjqDn1sloemtaJe7ROx8xF+oQ+NdXV
hGxSJ/8eilQ9GaxShpiBGTjxsTRm24Cg3JJjNtYEOB+oPXpcbCYdbfBbVHbuGgjE7hNuj3l1Bt8n
qL01h1YazWCgMJ3uhMOrQvfwrle2frGdMI25ylGIyEC09CwacCqEPKH9+CjdOkwHBA72SaFMGXS/
1gSKio5lFEP/VvM7RdW7GbdKqXpPzXHKtHx8VarAF/+i7+wLhDMR+MQMUmCIzyoeSlkK9l1HQtJV
mKLgKWNdSSn/UGZJBEHxxxe1J5RFlPIiCnuXKZaMv6F5n6GhbEAfesb3MKNI4rbCquSaKwA0E2+/
SK4ggBCse5uNQY/OBpPuh5wpOYgtWJq0gu8jmQ2ONgOhxBPZcvP4Lop9PA9InHlRo1QWPAGTWEkr
UN9JpRLwDnKfcjGynvyLAsb1ONubYgcsSaFrIHr5vVUJqvj9I2VxIrd1yGcVY01KOPu4zOPRMAQZ
KMbs2zwC6E9tKBPo1qeasPYciJM4wqibSrIKbxzB/kLuDe1gqAsCZjuZJzCrnYsrJ6YPtLmlpzi/
YXffmiJOTByJ/GRQMBDSt0PoVcl9C2O30YweX9bAdL83jurcb/kRGWrmwQHFth6PcqU2Fe3bK/YQ
gH1a8ldX5H3nfQvi2RUzkgzbamBLzQveTXMREZFe22fMMsfQ1O3eg5oiMZVdnXjc+eTK3CnsFncI
vCGH4TobVi8aKGgFRXdhUlbJL9tF8xhLHrf/OagoTzs6vCtDVombM7FTy5OZHVqFopsJmgcWRxpJ
/cERlxDss0jKTC5QNZ2bMZhn7pwVDS58sgO9L0pEAf18ovEpRNf5Z+3zSirfvXTITOXPlzCIOEh1
sS6GyVNeCA/LRkgBu6dqF15yNYdwkxGlgNi9D+9hVnJO+My5zxldRb2F/AIhSTr6C8H1XPiUuOS3
Aw1avBmgROOyp90TuNveb2APS2hiFReDWwd+THG++q3nmb2ZcdMR3O1meeSqgivCKvFHZ/xLCp5v
V7LuN6ZH3wT7EJ5H7wp8H+CiYufTr2PtRG46Bt6lSO90YWsXkE+hnHPVHy5FO8JXKq3NlE2ZNfFI
kYxtIuYPEUFeOJ8iEAYZ+40aauD/79A/dFu1WVIlRUVyXGkiq2IPvvRPRkg3UVgZlv5jC2DwALMu
5AC6eYXjXpXLYrz2BZJkS66tZVuqaUdC8V0tFyhEJKuZiU33KBBLx7S/t32cWcCGorUXp2zhkhgJ
2xTkx5r6gJKvBAsALz8rKKCc2XAmITt01rwVxV2Gd4pgAV2yJpDS3HxOSCmUhyX+9MhxiAAbmPUO
sKyKSzW8ukTOSxwLfk69Vf4MVLrG2kVBw+Cosq2uTvKYPBoGlgXpiQ5Hj6RZuEgULwWITEwiwXu/
We8ImBvkXAeVEoVMDN6aVa4CcqB9T3FlPBnW1G2LXqlKz0Fn8HuIQRr+Vk0AlPlfYLeeNYmy0b/S
L2QGk9Ftz/WWeTpgKqwOYuKgp22XNo9ZCmZPZ4nHGKanRCt6++114Dggfux6VoLlPKenad3rUNEa
bHCqDXUkS1mG8qIc5qzdLSeKejoJAtwobiWBWpDJmliGp6GtqsjJzdkSGsA60kTSYpR2xiqx2tD2
zfwxcb+3VwCWYxVgr+bZsjrEJRGM8zskXiI77lqN/ex8yZ2H/oqVUgaSexfj1vau0dvJX/a2oLhR
KKFiGH3v/mX2XqBctUnclTClvrjaQnPuqs5c/+wcsQ6aOloq6PjqssrWQG9RblM3+jfeEBoNQl2s
V1kKFA/Cx00oSagzm9lbCcFBYSF6PcNGi7/M/OSjBWOnghiWr+X+iyJ4/E8ZIvZJlFkzByLyFXkF
kVsOF95q/eipWAULU02jD4bHpoHP0c7512b5EhYGmrKKbQrDLkw6iVwoOJjSWfWWFb8897xT51Fo
Hr8eZHWs6N1LVEg6s9cP7eDeI483+W2eNPWyjUUaZA87/7J2Fw7iNoDlNz/hMwyrIWoOa7LPaHwv
j8PRIxq2l6jXo2GnX493ggz1r+dUdr8nL8Se9NLNSj2xmQajUjMsTDLS+zw6LUBDuSZwmgPcqygp
fc7ffld6VHMBCjOQndhrdV5MJXqS6kFEVEZMayowgYnG+mMnH2qDNN2v50XfwNZSK9IWdz4aDN6g
Xq+iX98OMO4UCoI281qbvaP5fEMoqLcwx7ltcrsh4PFijSB5/dDagchOzHwvg7jrZEnVhsMpOL5D
Kl+YdWEcPYMKwBc8i09B4kSrm+NGgzAOaZUPZp6s6v6sdpHoTwki3OsLCAp+HWcnAeSLAyMnUw7b
c2RQOsC6LzJXpB/kH9205/qGQbK1/sPMIYN8Tex6NMqAbJJoO+jqD3uWTtbsrrMSAGURVEN45B1Y
fqL1ARpPwDACwpSAnyRLhbEvb9lHzS+2cyPywizApyiJvQWTO69hjc8gIA3VQqYyUP5rXYWR+UVu
RBvs2IiTKRfZ/oQxUyw9BhzCs1yrncgPyPzQlQIKfZvRKVXYXvutFo9GFWiIokKxsdPjykGkGBeX
ckyHHFSD7kpUYeDZTVSudKpz3IeMs2RPIeWi31+7oFdlbnffvSgaW0ElQPPpa0gYiQCR8rCq231k
FlTNWLZizQFYf8tkxSse1npGGtnq6y2SMiYz8ygk32AezvjD9RY003wzRmd1IHUXBRNHuTB6vSGT
4wF7K4k8Qa1d0rdInTSZ76kMRkjQFLqlo45luvoBBrrztqYDZrp1heglCfN1SJ+t3o6Y0pZHeigv
82SLSHgxx1Fh8nV3to9PNi6vaiOWeoUvHEAuf/P+w+aLJtojLDwxlyHrsFEYId0bdhrtz6YuLg5L
J8Ee3ABCsoixyt9H/XG55ip9DhrUEKbtH90XDF+Q4dDMfZralClXJvTw9uryoQf5zY3qKSa/u0KF
E8bWBljcxWK8NbQLmjcEoMjUZo8XAwPK6eau0mMv2ivB4zf3PJICb55+FRrehXJRj25ekaKSZwaj
tAmPFL1KBSKDh3GSoDtSElFcrojq9g7Ju+Zz8YFbQeSSpZdKKas+MOaH5gwLER7mo1uGkCXf2aPR
iq0RQT9UduB9nXHrQ/WwRJbNGpeXu1McUsRTZzIwb+SjLK++wnxuv88vPLSLEB2xsWWHduocS4OF
yAeGA7JdekVBi2BpPV/33JiNATA9rANLmD8V7KimPkjbxzJUFndpODucpQgqZug1zSFhhOYSQR41
nSmJ+pp4JSBmvwe/qN88mVGQsHlY0dnLIktO0V0C9vTThmhivOKzKOD3XFUFwmezezGXnyGw3iS+
SUWWZdy6DYiuNYaDe0Rz15NrCyMn22JZ3ZcUibWIwssSi3MV36xZ+wKlbgP6cOirpmxBSfk/oteH
bMQU3sdAYFPbzbYWQRND43GSlGItYHme9ZOW8MKzZa6TyCwY3fGULGxhAhr4jBia2mtFISlNePbl
vWVM6pcppfr8f6srdWI1B1oC+JV759lEMUd/g1HfGV5sTjmVjKevYygHC2SfWKWCex6/oXkbnq8F
eCilTaqey1atfBd+SLslF3BrIu4kXA+lNKZbSzw+UyiG8ss3wIw5hI+MPi7//us0yI+TgfLdWmWE
3LmlO4eDptlmqeWci6VmsxgxVnzO5JByAuNypFO+iMDnNz8Tf5UhPeFpUho0Sd3Q522ewQphzNFM
T8VwLu/d+T29YMPflrYQZBXbE4nCEm6vQNhL46y5J9vqwXZWoSJ5UqG0HxnR+Tad48ASoo2WZhT5
zXfhi21UxRccjDXNWAfQA+bwRnEtGK3r/s5l1PyWKIrgG++BhdAvfWWMLMni6YP/IXgH13PY+ofL
Vym5Kkq/HO7nV8TeeijRyPcBbKpXWNTTx3Iw9EdYkYEGZMlimNfDmWDYUm7NF72V1GI+94RzwfUa
Gc7C0MD40BYo98YIEHDgOvuej4QmDCk9TJJAUL3lpiaI+LCTO37y5szeZ7ZUR6PfIFP5niuUnrto
bKcXh1v9DsPRLlh6dAiUamJDfFOtS4GCrAoLaLXaoUj9pCXSjZjy8bldBXTiQQxw1JQLLKu9yIFv
gHOZlAcVzwdA0tP6unkzQlWnO1t6S0tH5hFaAj8e0ZknBSTTZJbkMYUpzHK/4tQVIrvpN4Anse2n
f5AeLC3jlwoSl7RUF4e/m+Xv5M1oypsMLv82qBVxMUD2ahHvfTqZIsNlDo1PJQbvgZtPM3xVsLWy
C++WxdnbF6BHWbVc28QdKD7OCUwzB6T/CFLWSHGLggncMAYr56q0/b4C/TR4gcIkCmtqV0SViYVO
vbc41Axs9N5UQy7OLlLhmywF3GiepLMIrRZ5y4c5L5E/L0iJEDuNns5Cftjgf7vlUMvHiPg20lkJ
ey7vXxpoT9k7Gojh18dKaZI+2AKNO/0ynuDdN8CAhzHs1Xkn4gBwaF90sHwpMfq0xU0iuPUYIqYE
L9Ha8ImXZvT+Da8R4LRkaj1823DWsupbIiojh/GCm4knpW5RM583LoiHALBG0xm63ROaImQAQdWR
mK3HYcqfxzcIw3qflAk4M+Au1PT0TN686+pSI1BPX93METMbMyUZ5olgSzY+nf2i4intGP2VkN/K
0zcJ1kSBwTad1U2lXvp7e+YQLvRmMWXveL6JOTSzULTQhGG7hUAEoiJ14up5B7UOarevUCft5U0S
OG78LN4+lOVqNDvZxdMH6uEAgjCVOxfqMSyLuBo3BjgQn0CKjH4JIhs3q50UJiFtsigDvCz+trjj
VT+Z6MWXST8z1gz2YcLiMXPFzyc9YeWh2/4cFKx9zv1Hcdb3cE6QxqIpDp9IeRtWW1klSofvcV3i
Uq3iUsh+mx36cBi1gyW1F4Kxk6l6dV6X9XbY5OBmcMRPsnbrH81NZLn36Wf8CSUWj8zcAXIBartC
sgwCDS6q1Hk3vUgHdMaQ0kVWM4yn7LLM15ZOtudY86Pq05K4v4trLrPzQof83kNPqvIJQxF2XSMj
jR11UGlEi91HGUFF0VqK7NDkf0DTexEia4JS+1fKibU56o+6mcGOZfl5NP6zA1vmukVj5y2aAD1d
2cQYUJUa0Id8cnopEdt9sDvJotQ86yLRjmTGCOzAlZnlIMwpmqmPNNIOnTpJzmIZin537ZKSuDm5
nM/2HvNvJW7vcvha0CYv84kV9stUQ0N2g0Aqszt0RWf+y946NUeC8ncIUW/2jG3OwleJse30sGTU
SO8ftGlx9IZnMTv6PcS7B9FICStw7l2xe9WFZsfLKsAIqb2nmYmdFnKTGv0YMQlJz5Bi67JjrFio
3JBSZwyZ2qb6p7lGgw6F07WOqVmsE2G6WtoRXq31SYfpGyzaAjYznW2iuPdaNloPmrkgy8l8KT15
y2jcMkHiuZnYRq5NIpLVlqXGw8hPG8zG9PnA+JMod7FEcIKrUZO9664SAJeDAHY3YnS90j3vl0m2
r8WA5h/NgU2DFUgKNve1psfUXd3qfTHFqqdxoQ1cakIhhgI+XaZ767CskP/AITpuT66Fxthv+z52
zOgQRVuvZySPKc1lmLduhznxWA6eVMn2ECc0Om1kSRLelmR+C8M5OH+gm/tn0dRRQrO/3P1hBGbe
kCgu/FztZ3XyI+OQSyYi/Rmsw1xjeFUytydHTuPjxBQ3/eyqVcQ5Uqb9DnS4VE/Tc6kwySeujYEI
m9VJuitV40ZNPlcloTyJqNgAqi+wueMxULZmFMOuw2+elHzeORVp9yZX/LiipZKO27cGoNlT7VCH
S5lDpA46NddcBCOc6CPeOGcpnTHuDv21JwoVy9XB8OfeO4Ke/xV2nmWc5lZhpaSGL8VzoXNEDIR/
EUQ3oAVqFm/wj93CH3j7N78OKwLbY5LrU3L9xUHNPmMJdv09zE+Ehdk/ln8iaF6oERNeExEspqB4
fUhweQiJZx2DVM+ZMwYoFHCegepZWd2746EiQqvoG4QR1n18kR80+oHnCbDCwr90fXYlVVY8O7Fp
2pAJgh/bcayXotI4HTnqPuFbdBP5EcPt52hcQgL6H/KczqSmiioOGWPDeP2dnwiC2/wCq4Zb0iZE
xMowSn0MICXWiuELhIhq3BJ05J2ryWnCCCpzVxyRvGEq4CtG73JYdbB+wwPR6gxzmD/s0PC4LxiL
/6wt954rIxaUzZT6E466E2nE6f671coccHNhQEPuac1oF0xXHCXRrgnFmLXY02hKF6vKW+TSqxOz
1/E5t8AOi8BJToNzO2OfPYHPfBzNfzaCgmk0xr1HnUgMc8hRspeA1nBOI9Dk8BQrpa2fbBsTpMoY
95o118nrWpVeY5GkwtoQvqHnZNAe7oQuG8Ae2GyC1UTKp9lkaU+FgAnTQaXfd4JNUPQ0Le1SHYuj
yuMdhXQSvVGbYxqiyY78TjqER+fN3qXVXQcFVmmIjAhU3NXRNGvby3n1VX8KgTf64NdtmKxqKFm2
AjTeGYfdY3IUSeMCplG5jjdeRlzrQVIIN9L29hveGeRGS0bm/xQkaxjxL4W9iDWWis5i/O4AQdJD
0cdq/13a+5Tg5hHTdSyWC9N9RPArta12oP3ryX4LD9QprMvqklSDi7lX2crvMB04A8JOtSPNeIQs
rbsh7R7G8Cv6Vrn73qxtNZnbATpIus3PisfI7FlVgHEST58HRVTYIHvviLHIJ7gNcdmoYXqKv/Lj
vljBuwamPPDulasp9RPeJdTxUM7K+ZvOHIpUKr33bWSGC/LQ/LY2KxhHKGME5pE3KFST0c5jagOr
6ntClDhPxtNs+unUv63F0pGbmhTHI/2rb/lhnUF5618LNQExki4UMDsHtOpinjrHMzFPPE793r+m
yQRL7vyvs1RESlvq7exCJQx4JkfHbM0XkpO0uUKWOkDfqMppIWmG9gCuGemYznjFBJIKr5rndC1h
VffdFaPGz3KTGygeOtsoiGNRwveuLt2usqg6R2aPbPW+Qr7MoiVzvKg8XGIeF4wK6YHXuKMHnoaa
GznOmtsKhRfcxmiv+sWg8TBQ9BYc2E4DGxSAvivtWESFxyGE489XWfAZwEdGJlUR0rrxmy9j+Tj4
qSkygscm1CZhgK8PT+2VSue+fTathCcXBqGh3SnnY2CPzEhjjJn44cJNrTdx5dGRs1vkY66MNmbN
L1Z8LiCqogtdQ/eVfeauZq9dlMljwijPWXE0/9a2Z0pu1B6Xtg6K+scpwJKGx8xuSxoVaNGtWCtu
JMspd5tWkJlzU+e3p1EO7/tkQ747QqYY11ICHZYY1oUWWrezqAlLjpDaIYQVTXEH1ppVrxavd5AP
aoSn3emU9vfZnKSpT2Xptv/A610meZh9UqjtRyHF/izEfWKA5ROhGk253COXfV2/ej2y8LCQVXu/
TrYaA74+UEsXx3END+ruvsP4SqJBmf4egadOUB2PPSpf3iWo7lLY7wje9M0Y5NVe8sjdlrzLIOyZ
Gg8i36Etk5H/asibV3Z7AWaPFbK0rHL8GI44NCOiG91T+w9qyhH7ViqZARKu91vw7VHwwXtiDN5P
EhCPU3+SdMII7aE+xVgvs4cX7JcPzvYJ67Ok+7ynuDz1Q+0hrCvUeD+goaoayAtZUDCXTKZYn94N
5aEGPo8oPOn8NqH+lnOnSTeYpE6nURw/n168BFjyU5W7HyKDdbu//Pi0szP18qR+fS4XegBxFmea
stea3LEat1eMuESiRpOmDiUYzdXi5DH8wO3cWZmXdLU2apdR8b3SuWyarvKiNmlOVcGC3FznSPL3
/wlVAgAksv4xb2VMV53h5gxBZgflEabbQeqbMYlYohOZy9i8HwROsEMqTcXa3/cvIlsKjSMkMR3W
WPyuXalubkr225Z2zUNBt0qqbbvvuPD17mxgRLaMkRYr57XnEHPL8KTbNUwBoknvtMY+kTEYqTbQ
N3UJwTkKL/FkqtHfWygpqYxmni7hqEQsDde7NLiYsnZP6dNqe5SRKQkLhXWJ8Re4hJgPiHnPuszx
+FDta92o/dNYAEZTPYAPg1OtkJGs5fSAXCCsc3UqlGA9mIWB7b5+ykZqTIXB+2e6c5xKhBD8i80h
pyHOdm5p+jZPcBSh77byy+f8WDt3S6rZXeHCeF7jywvrKzxzm6ED3ruWrWvgwbF3UaAk013iDV0N
Y+esnoob46vu6RhFk0LOffD3eSdx77Jcba9WOns/lzMy9RlhURbFIJH/hF1Ex08HjHyW6mUDWXtF
kNDP40wNt8VaQmf57qKn/qd7tmp94HnqhEpxeQTBlJjn1FeFUlKns0vahe1KKBaDRQkhkgmQRMAw
8x//hdq90E/vjOkJBBTA6748KGJECUqUHtbclM2v0sxcDZvqXJm3gK/WN63E9sXSGoxEpBHCqbJG
SCNeVMiSWGa6fuzvxsbiINB5uN6CA9Dz/ig3ZsoRRWyqmCbYYuEerBs2umM2RBCYm8HNF39guAGn
kFdQ6Z6wd/M6kwoVY/N1IVXFh4h2Ghr2JGNX/hkE1zx6zGjpePsT2ZdbyqlQ8Ec6fu0OLJETg5vl
2+dckGzGre3CZ/5fHrQUS+rQ0IXo22hwDH4UovyM0o2zu11VFM72oHLZCjStBbKBr4hpSNzCeW2t
fDR6e/XNzw9IzHBQVbHjikwwLJ4jGHT6OKno0jUTaBOl7OfbNzjQMWQkkFW6jb3R17kOvgLsoBWw
ryXd+jgY1F91Dj9MGZp448vsgRAoGNA6dlBrLGAjZkgVN5rFvAmCFZ6v06mG239s4TmxBEXnzdBz
TY2A2A/Z1ke5G1Edq7EMUfniNcw6LWJG4dz0u6Ea00fPgGRIHOW1axfz+1vtF5wy9BiHGjF5ljJy
H3Oy+Twjk8YKp0GMQ+OpXXUFLyrhGlcSHJj2OKq3R/56OW9UUg4+DXoDO78l1dBZG/in+3bheTeb
ESK7RV/Yjt9/g4K2vVV3kS1B3BSt4Om4OEtd5n06B/WZS/wkUMp2M/sJB8nXWI5oAEoxLOZ+bK7z
WAOnPVcZYQtq+JL0HTTxaQqSS29CdSeXgXPPg7MCHdBpKWkiugsmWsHbiEeA02cXvcil8uBvraqd
SjWqtAr205lgZnN683tGE5Qyn42daNOMFqD3IKev0t6TuqCtoV5O+NM31zoWqxXu+/MunssEZVMD
HV8xmVaj7W4oa5JA8RlpWyMy71k1qzQMKZjGaqgAueQJp0jL90pfCPQHp51VZTc60rLkW0XRX0PE
uBGize3XtA6jHphIQvHPQf2FlXD6Y7tdEo/H8ZejjsUc2JsK1xWqjufZRV80TBUbaZrb4vr3FC8v
tcCVM/bWa4rudVvDa2cdOPIlYvSVdtwW7YDL62Eu0kK4tvUfHQ1yn9ixV48Wn2NSPfuRmXJgU92s
jsLbqjFzpW1TsoZulDvEeOlb2Su8Uo3lD19zapKMXYRWeCKHECY1H8Jb7JIT7yAWu/fZFtTZeWvF
k+aPtMe8wgctD6SqeSVaPQI2zy9hxxEnzJaXewHjcNZrL+pOIrLZbj6Fh+cp/5ZCKhRVwjjO1Ljc
/D51cIHPi4EPQHlO6CzVKJeiliFjhooSCrRqkfhGT7EFLaocrxc3wtZNt4taCH0m/lfthL/9pP1u
G9kMzCqzlvGJR43bgELGMl8FWsH9uwOA/paCtlHZodi0YvqEzqP8YJUsS06RBjdVyZRBEapbeG2r
DRiempuXHHFmGsdp98NNZ3oF7UAQUZGJpHgTnnDVJrxgFpff+R9rrU0WdC5WXU7ld1vaeEk2S6BB
Rakh9g4rNK5lXU+4DYfJaWYf6RwCVq215FWgpu4jQToaLJagRb4IuzW9YH1U/BQcjFSXZ3fbZKn9
RAdEQ4bb7RsO0NAql9NBM8qaUkK2cAGgf9L8Ef+v1GpfHbVehnXDbFOOJj+SmZeM7y8WxEidRLnn
U2wTGV9DetjQe218aD6XnXWDV+G06uV3Iki5sjVeQl+ziOSelFYhZvKGyd8cskJNG9ZzSCtkxz+T
WJTwv0xcj6kHCWxvU9aG9VTrBtCDng2FpyQuze08USR3Sa2OMRKUhFK4rvXkxXevyZW2Jrgi6OwL
A/BHlg6n07qGTK2GH3PvVqv5WJ7phdk0jNc9cHyeduFCaGHzqML9FJwaYJddK224ON9BVEHXxUoz
bo+ZAba+hwrFDucV3K54k4FY1hbqOTbCFV9kEcmq2a0ZKVpEjbaorAP+wBc1ASANFjCN+1UrBuM4
GRl9Y+5xmLLsbtq8XFhMGPkb5Mwj8BROEccmVkxwIsAVlUqqUWOwxqENk70kZqwXOyD3KpLxq1jZ
24mqZ1NOQ6YzbAUCwtlepw9xBQ79/KydxQBXWEPCOsEhnS60HnQrhz56Glz8G9VA4GCPxUrUUQ5J
HYZrCHW0FAFUX4OvVNd6Ai8l2xBl4aPFUEsUn/weHDfcO7DPZ1gopbNRDwWE9G28VA8QG5wZE2ge
LpBQ4CDbrLvgPO39oC8Qx3OT3DKpX0RTdGNfcRhAiyGnINZbmku/YRrOnT49n9U8FdTDHNK8WcFF
soXfetcb93GAg8Hmdqgv+DVOcj2V88KQM1/TJlrjgUulyp2yWCzwHhRRzvWbvNuSTpVpvdC1vJ3Y
Q0DA5yS03JaOBDmzL7ekCAD1lI/p4nqvzIsqVRVdqS/TmXlM7xVNGdDjGJ/pALALaXYmBkXL6/AR
DfgGd8q0gZMvQoKefcJDfLZFlTNcrRgmNljkX0ZqNZDvKlm+gQuH3FfNFE4eR7o8tYC3S28M9kkc
zC8tsIysNiI7AxLdr7xZ8zYJ5LUa0eGiOfie8Arnp4rOF84gV/izCwJjLq45UThYWffGqid8gwDu
aEgW809+TM8CKds+ATjacBko/6dkNjW2+1W9E2SmRRlcVXO2ExrDq4jd1zPxFpwrPlCxmAcZF8gV
sZrCR4/sh187BM1TrhMrvky3wPTRnfV6hvuvSLrdxSZdcv0PTqUJYYnJZafkVdRtOPzesJP7GB2s
TdV9Uj9uOrvwdHmpCk15H1jI0Sy+M6vGWqq/jN6YS/gmRFwIll67erAnIyVxlxi9Ni1coi5rVUbD
g5UyfCJzOZRfhnLut9GZ9LKVRz2fiTyW/o3jz9W6ddfc76k4Bw8coLiWuLuuWqAWjZikLi6iR0PG
0OHJdwaJj1x7+v0rDBvN/xU5bkP2XDQ9naFPcq2v6EIhJsgs+LB0GzdpxgtizIsMaJk1BFyQQyWg
X3wO4XkElgxKX8nkSpnNa6GEKPrhEbCT8JHmZWcnJIEUMnmw6SgsNNPQRq+6aCgMZU5r4ax9WmoE
tkk+Tax+Vx+gbBmz5f5ZZcln0BegoKA2xK6xQTJOgfrQsOjLAoWlRx6V2kv8+socJKZic6xWkOPt
ZTJyS4P/dgDtybEvISdZ+7/NP1hzzv6wnoEt9wG/g96bHXcJa5VBCh1yl4J0o7JlTPKQBIyx9LmC
gNGvJxUJaZKCrht7hUBMuo/WelzbpeP8V69G2N3Ya9+0ptVq/k2CdfO2lx1hPRFnW3/xeDUAjGJe
cLrIF3XLlsj6gljokd7FMmooyc9FSPe1O6naVPfDUBwMtrvqtLc4brj8lbGQIsnxVhTMKY4nHBBd
mOkCQOtxvezk1hYmOMSxChNVisuWRog44zcWJqCzLJC5YE20zC7Tpc6GTuiy1lRZG2y2QHrQ7ufe
WqISt1ORYSLDwS4kMn3xdQp1qq6kP7x/fFxpNAehzT3xkdMGkaM8+WGKgBicHKsg8VC/eHlwTuWH
lEwW9G1/0LonP6PqLEP3+8n8Vyw/cGiF69UqNNi2naA6/2vaAayWSrKWnxkiy5FCDV2OfJV8Pq22
VOyQbi/Bay6aBdint7ZIs1GAUyGsbCE9e0IFNgNKCapMLnGAYkwsIUwys5yTkYhfoLtgQOVE9i0P
XJeMrKuPZATiQwCahUgI7BLwQx/nhDkfJKFxGTrzSPaz4bJ9LQjh5byXtev2UTGz6RQOZ5soqzHO
UYqYjuMasEDkw032F7UZGOGxp7fBI/2KLJ6UfjY/KybK3qacMV8c7yGq+GyWurV+yzJ0bozJ5oxj
6p+qqostFXLXHT+eYfDJRtj2pm2LXMHhohW76sRR9rSOdTL8GO/KgqUZq23mBh8c7P1HVSmPGxJ9
oSwOnBMUQ+K02387UkljN3uPcVUylFHW0B0wlIn9iW84AbReEVsdRwugnsIRZYe23o6tCNLQ0By8
W+Ktse1C5hpeiWWoQrJJtuSoIkbdonHn7LXtmxufFrp50xhG8mI4LOgFrExAj/ftmMfMywhZ9KWK
CzIbKT03fNOo+HPaj0qZBSROLij4axEgaytYyaoz1r9DIjp2FcSoHlorh4WFCgZwhgegRyRVLdG/
1hKVApfg6YidDmgzdYipqx8P0V4/5JcmNy7Thpp3ctlNl6BICjJzrzl6vemrtbPtQw/i7ndwcRGV
CeiZP7fhp1Km6oGD3XBimD8zZLRGIDXH3UvuMIdLTokLUI2yK7zf9x7Yjbiia2HfEFSaVcnz5+Q7
D7ijSQbM8qv2c6uBIgP8ynTqa67W/GziSPp+D7cR+UiJHsstsU0XzXBSGxiDsXyd1hhbp310wLRC
cKfP1GGq1yrLmMSo6/0MYxXyKZExNaDpj8FCJQX9/17bpDr1ER6pLRSRmOSApxkWCDpHZ/oyltu/
s5gNTvq3yLhIrYgDt5UL5veomcpqBs7raH957aPKyDlpgRk00w5utMB2JRB5r86epkEBTM2QZtqB
bDh2J+xYZ6k9mB0zbfvkGokRmlfzif+KWOx2+2khY6WvwEe15+dT/v1nRxWcS8/bjujlKpWc4QjS
XcjCqKP0bCgFFAfh93MTRFYstnAF3G177C6meRtV+fcFANjgHXDEjdr1Vh3pyqsrlR7SQ0jOEgWd
qg8bNAdfbOFlLIve9RNISEQta9RKZp7kWl78K5zZjnz5G2ixKKzhjt53zOyj8gLcN5OuZ2xuPJOz
M5GTPHLMkxlbb3xaw4Dtwq5w8vr1NMVx1uitDoiwBk8ZwvVAmLMJZXx5WELFDEX8kybsB4NCI8LO
sG0BxyKeYsJIt0jdLa/oX0iRI5wvyqtpMaxc2Fz69gD0ttbq5SI4Sb3nbPejpYtFdCqYZZx7JxPP
sJ0cq//0vitzHoYvY9QwaI99Tl0KgpUYxqypNw26pVJnuzSXF4xC4pqauEeWkb7dKtGailbv3s0G
lJ55qIUZ/zR7kIv9JxoiRE/gTrS2i+5h6QWViiYimKOt/gDB4Dwp1W8RHXOF/oeRJO79YWA2IT2a
xWYpm0bKx9j1E3+DtJIGEqNl55bHgNgzOaOtjXTp+1wO6BDRNiHwuI1uu7U65X3ZoMvFx0hFgwiW
wXOIP8j6qO9UnWKrvpyk1vG7ce3mR78DUEVx/ZAByo/dDYayu1lkZJoD82BXak78+ZvQ6r65qgWK
MddynbSBsvh4C2OqSXubZNrr+d3IqgHcE+T39TMaG+eVUDQeesV3WihgO84rccEhbDOmWZ3n0QVm
GDwJI0RZcKD73E63iV0ExF54kPhQia9uPrfKtJAEUoOlQaudG6xqTXoHl/7p2V/jQ8A1OIm3xG2a
D9nc4KrkfP59co0FJI5ZWrVW+LO5+9Vzjq6BUqFQnl6+pRnho+XZueH8wvMbnyTnwqEF99wNxPJY
zaN0uVcEgfoL+Rh0BAm7+ErWokHEA8mU92t4KqeqCJa1pwy2IlEqG/oDKERW91S7uMBpLGG3ZOu9
EW6Lx6l6MA6z5X1GuIuRF2PNNUG5iIQzAWeUs7W/58ktsGtcgCFSkzX53jepV3JmPkUemv8ZLFR+
yjPk7Wug7QFIEEYhTVYaDJXjo97wD3CcVV6PQr2rU+b9IuB/DaSl+2F/lrpCGuGyf3EqIs4Cg6Em
2cTdMWoZDVsJoQq2GAusQqr15m4/1k3LH3/dFv6ZAD9XSTmXPqplEVI4PgLiB8Wt8ZukTEBSE5vJ
O6Nwwb3Jnfg0yFbyqxxiZZx0qdlCE5n5jHsGdE0V166xgHOnUUTK9XLAuLXabmb3JBmVt4qc0yVT
I8O+LxCDCKy0sRTAYS1s2E++v6wS0h+Ahb+Ly8/VVf9aePYvV6E6NPjz+9V4SokQOYyH/6pGY36j
3Q7zyrfSaQD9V5/lBNr5wBMfdAuO7X6NpT0gEWhJulG+xS6y6qjPK9BuFfS2HPmNgL6ZHciA3ila
Q1ekblp6kIG9yPCB7y0iBytoqeJzaMkphlqsZT2zbqfghNnUA5gC0zxY22PVPzSOnr46k8yLmJWl
eQgyNKnGXpyhJR0te16CRJWK3eVH7E/LMo28b0tEJCg3pzAWJWowNqda3aqtMXzafTDWfjYxjez3
hRMujd/oFZrUgaJFkpQScvBSxJfhb4qrAVzYDDN1WsuToo6j2d17z0nJC+sZttfyDAACv0mV7cE7
ZFYxmZZ5AdeOV7h3qeq4Q9BxrYKXuKIhktnVtudF4/UAAiSN8ujLun/smrl8TONLkZlXJyiXNk8W
M6I1YcwpKA+vWEeUmvkjfHJri17A/72ehSbGwmCd+9JHtuj9iQQFgQz2ZuogOcOMiXqnKUwSQqfy
5e+hcMyrnFIcfJLX5c72iPF/gAge4LRFaR55nj56lP61PImPW1j3uTK1AxWYAl6owMl4ZCF2iVtn
xLa5tEydK1Zp4DW+pXcTGWWhFkrtzzaQcHcpb5dBoGqYA7Ris2Ehyl4YNN2wOED6QxVvENzhtj9T
AQaYBnj5i+4dhzw8H3Vi2Lns8f3qe1xulZOfmmFHw9RWNC2GrNos1BkFQ/FPMbjqCsgVHAMoTILL
mApkqwfKLSGfIVcPWzRf3+g+VAbHYVxwgVktDYG2E/fdiKKxN8s0U6c2mgADuEdY70ECuoflB8t0
CN9kNyNoETINZJb3KrDxvf619gjWiE38y0oUL/rdhftWTIMFOCHELB8TCS5b2XGZKu7o9TxWS9v6
2Yr8r5SiNBc4jWNMEicc/vO9u6sTtOMM76l7N0cwtYjwEfUv8Z/asl2OsMfZa0wFubcQoBHSlR/L
uFniCfedV4Cnv3BjtJoU0UFpRiI2Yib/u/KuLX61tIluNgUabTt+0+I7u/XYasit8DSX3Y20xMPk
LHP28DZ3FKQrsZxQLeArRUdyhACAu2K0nQRLUh49Pgogs6mck7RfkeFChnBqrQamsbNJXwUhV4EE
iXK/OguKYB9VPqu2gw36TcR2DUpRTuJhhvUtbAQdlStJIwUyDUPZFolQ289m/Eer6NWTDBSqcLQu
ZX5r68SWJvf987jOxbMbkKAQG4jFsfMhrZHahtsxVoNkj/aDl1LdGOLqtk85hTfsh0usBzpNtceE
nWr2xuy2J47nibv87AztvGBKZVtR/HLzEOP25koWnYXvK58k4pGJvBYdtTx9GXmByUty2Hlbji0e
ZEeyM2gzjUiYqmbU7caGAtBBOnTRmYlwjFWWZClVnsK1DryuDQgXjLwLqFr9twkcnsbXCVR+np2I
AgRkAxb+kpClT4qNqXc+YPB1PvRhD9Ru+SBIJAj4YiM9B8FGrBrNHVNAFhSDxwmGIg13K9Gy4SjJ
1zpCapQuM6mbZV0YgQgB4uJLnQtFiO6Egfzis9F6tbAibcD0hQAaJo25C2sVRkOj6HEvr6JlDoDX
wOPZp715H91Zl1WxTzg3Pk5HKM4QganhsxTkhimvSvy3nD5ojv/H/spLYjDGaoAdtcYC9D502DLs
Zer29mBHJo9OEaiBmlmuyWHyRbCnRyqUxtswnlcLqORRLKTyYK0L66r6ldahsUnsV3lSpC9YFPhw
CwuXqWMZNl+oonRtH6++Cw/kx9qmZZiz3bvOQqF16oG1n8fNOSBHePFBH3x6Uy24n+bEUTZ9HAof
1b1R2rYWjQFE0cZmUnd8i7GQWdnMLocbNE5uaqG59yg//yl/3htXsubw/P7cm1BtAXCkcyp7aqzk
ROoc5b93zegBbXKURro7adx3f7iaFC0+V/RP50n+rFlp/U7r1j1Q3nMwip5K0pW7y+1kdHWjrYjB
5TmQ+HZS99eZukNLCBVrgl89CP3EqavoJWcKlZn0GBaFMsmG/q5uPZ+32JpbJPLqZnoghMc6+ng3
M8J7KTLs5YVpUeGLF6J8uPbZ3KttyXgLwZGSIYaMDdaf0D592j8FcGdTN7wZxd9xCK8zfzlcqfAl
0/i9vv70qhtOPyvot+q3ddVSSiQHkU9W1jYjlKBDsWbegqLkQuBvLBOJM2vDKpj2IhU5qCqP31qR
tsUVaD0M/qvdRMDlKQASmW4hlIh30KjDMYPt/4uWXuRQGiDBMcxAk80xVTTanlHdaBYMiOBey+C7
BG434o6vekDNvkNcCfgws1jSiR7qCFyEWn0YgE27XjhRsWs4EFUGvvn6lhwal4aAGfsXQtA44naH
hdYNC8IMtZkzSztlswMTN07HNtqxxDWNWrOC4D893aCN6qLJKPXH142Qh2FcklVK6i+uq8qErfe0
Ccw9VxHVB40sbYxTghZjY8ar5K+eWXdv09UH9FYzFZRbjLjaoArSzUDhA4ZFOz5XYpZNEKLhfr4P
J4PxAmX+fF6u7NUUX3KfStUleTOsTSn3tOmq2GCp2lUtM2iQxQUJcdjZnoGoq2Cdr/DxV4Y2VE3q
+EfVEwyLKTzZQC6DP092s3Oq0RlUHghOKDor5OmGa/GcGlwnrNbtByoQTTH5BXpVLqbxs0/1CAtD
pNVm36mBSEQ9Vghc9ttnAC7manucfHSbrIIQPffL0RXSxM5/wmPi4G0fAvC4F4Gpbm/3BKdjOw47
BQi2Rtr3QB5h7jzQDN4weqZp1xfGqWs39K9Cj17zAau+JtN8p8qHhI52V7oGliIQzwsutFsvjUrc
2ADXYydIq0zlM+Vj5iStV/SUg4kFcC3i/3lQrWINrFEBBqFxcZIMfJ7+DTsccel6TBl8HNsvFrmJ
5giI9Lk5mNeELzHp50bH2ZlLBJochm0PXAhxFG7Yn/HNOTf5m9VXF/iBOdNzqc0kwRBq0PUwsE8N
uTRuW4e6byGPH2757dRpiZf/ixqEvrRURRvJb6GpHo1gGFNRxJa1VgbkQusLwWTawyKyQEQu44CY
5LlVHWg3FbqzlPZ/HzHN2R6FVAfZTgUUz9/DpnTa2donkuDatoPzc+R/+i5H74lH35vBknBAy9HI
axFaIsbJ23Gr7VyyytWrz8O3skFpY6rdnfu4ujBqMZJulohW44nlb6UxX9SFe3euns1VvzS2+tiN
IAr+GHUgGUw9HGA/UdINWXBHh9h7sNTQ/tZGcKLn5xDVuQs/1aNwHNR5mgh6QzyBuWElNDDNHJQ6
FrlwfGaJ05dHj9GaDuPPWKcarsKMG5tsc4MKf1CEG5WAEq/2AEqb7KTQNzU4txVAl0qnxLFsrY27
O28cyWER34nBsbYvnFgNytwTvhDAvTuPJN4LLOc2m9bEozTNNMDzp8CoQSVvpjdSAmq8c7J7RP5Y
3enauUP6qiS7gnKePyqbtN3ueYXt95F6qSEY/2RSPfJbvQcigrmJ/lRZhPJzQmzTdkEQSlf7dhx1
tWqSN9V92IdDkq2jlxIZKuRl6Dwxkex1Ff8ALKo2JiX94s+gUyJopnQGAKxbQaIKrs3uXDpskzZ9
+GU1OhXbgrVs41KfEIc5CpmfLMjwMqHrYFQP26s48q2+WtKvZOQYz59vQZNXHL33kI62ZqjQxY6Y
p/0DoDcRAaWUfJLTqAhSIHMn4UlCMQN+pX8v8X9DVS0+vppJjenXHm+Oc41zDVWBR1QfLIaOsIqr
DFNUAHnFkSWPv5AZkWnwTmPnQgKi2fwtd6HT2TaWmBlu9OWT3vWzFA2K6SA+k9pI6HuSOhThXOdh
46J1Ma04KraOZkvuZLp4q81QuAJG8KtdtNgyqlNuEdSiarNITekPlXW76sYHgrofnuotAmFcWvcT
wFxqM+iGVzSJmxWiJYaQymmdupajYT26tq1HqGXmRyXGcPqipQV/ROJu5SIv4QkBgDIOetylghzm
3fkU72hOE6EK+09akcv/LmUP1qYKQjaZM3fSItphl5qz93zu2KSQYEVHqWAb0x404OIrOs0+2NCC
bzMFy80oIKm25CxehFPJe1aj+BjFSx9tc2Zyd+4dWZFSIfb/jTf9v+Ar/DhZS2ligosupvTL4uih
hx2PxcWLadrJWU+6EuWNV4AmLAKbFGZV5P/TcUoHZOLtydwVSnV6aN4pE3MPh2OD/nWF0W2q+n+1
/RCQF8RaD0RNRgykEZ1vA39hvBd8UuEurcRM+I39b2vealtOzrp+IT05RVHtXZzwOf2qYuKjonh9
sUnOWj2upxWPffQT54T/HSIQ0+ELneeWOa+YjalSbCFywRgTHcYDZsi+CLuoTgc38l9hgvj0GRMt
Gul4O4O1KFRZ6BpXs5KCYp6j7emjuIcO6FLjOk6MJ4H4LynLsAwafVZgNSrknkxaxVqd06f/4Ehg
Mt7K1xnSTv4Sh5rKHQdr/efsNqveOX3/bUz3kbmSkE3WF1KsG2WKXfu3DPMP/fzSzfQwxQ7GffaW
LkEDKH4pXL42l/7NnTAivntp9ERNQz7Oj9BslKZ74VQGfjFnb4kD9QJW8O+ZS+qnaIoV4mh3g7y4
fzNmlBYv2+86ZDlWi56SLiemNXP10jV/o11flXs4qchg2NQY1FiKYYsZMAyL8PytH9HzChNiLkGA
HfboBNjv7kRUZtHVvF8AGUAeVccDF76VUMvsW89dmkXav6mYAEcIYP4hENRIvqNLu46d7jApCXGu
F1Np8jz9qhAoRbOnQoq3YL1voNxCko9133/SdGms1vUnBWUnfepN6hWisuJCb2EfpiKgQx9MAuGh
sK0nNbmJni3QjIMHzfI9Sj6wE0L8Pw4Ros9n/Doyd/Vbv6FwQw2vjWGiLhf/pC4Hy21SDmu7ZZbw
lH/1dWqIhyviHK87l2D70V/3Vrva5dZPSc8tOfP/oniFlMtWdyo2vIDJMV78Imx4y3054GPPuhpz
tdaJHcEzMVQl04txlsVUBxB1y2pzfAXSTIiJk9GL55los+ngFzh5niTP+W8G0JWrpb13y+OCKx1E
miBXmCAIIWNxW6+Z3gP63/+lHALwV3dMhP3RyFmthJgOK9OPFA9j4JBtP4+wq1nUgHffLvL8BdFD
LdbCCteuv/ODKntKap+jygYTNy1YugMafis80TZBX0Aa862Tgu6dHb1Xa8BQCzhGO6JX4d5v8m4n
ApaLxJoednbOBJ9K7VGFuOot8wBDePLKP2amNQjsuFOssHU3q/saNVc551SHMKTpZntuUUQoQFG3
I5FmvWpQOBV1NVrDuDwlSuiIMI79eZjJpBbO42taa4g8N4EtYzjrGvuFr/bs2ofUnMTd6T/9Y8MD
eCHaYQIIVPxw08Si+VxT7XPP6HYEWVQUbu3Jspqeh6c5y6jNzP/nMoMxbLMHQk0Izwud1QfdYN9U
rNYPN3WVWnGoevvT/axqdDu38qIUGKxyN5wbxwdN6wl30Lg4SdHdooaI3OVgnozh+WDBdkL0BJD0
PnZb4lVeTa8wrNZlt3b5RDi6u4rpX1Zp6ggUzBIJGMsax8bhT2n2qniqVEga+PTqk7F56qSRwZSF
uzefPbWWr3Hr/7b9j31eaGapAsAhRNwike+LPa4aRfr2y11Y4YehlM8QRy67hiYIs5DX8QJxNy4v
gfyTYnZOfShuw13g29PSqi2SdTUMa7U9/nhM5PcupMQBrizpYwxe3w0WsqEmZnlmUMWvPIswlwEY
5oB4jYeRXffCLbD5IoB4szW02c5N3DxXkqCo9SY8qZG2eK9D5dFyHnpx9AA7k9kulwmdwP0uiaHP
bgUkDi56rpCfqWxgJlNZ+Zvp6J4rnzgih+PRfms3/pzgcSc0RcS7A8B2ZOzFmNZWwK535HEYmx9c
Xv5bo+mRM+Dbqtbv2z1/XnSSayx6L7Md30o+0xKayQX4hVbBPIq84oOqzzGH8d5pVu68FMezJdze
gf0v9/KR33Bf1OdXI/h0Z1YVGRr8QlliwLoyE9TsPxLinZr/9RXPQZQNH1MFrHbdPsi2EEs2hlCH
k2J/LZXZMxI433wZMd47tevBwdlHVQ0YQLrE6XCr4o2Gf355DstIILYcvRmjoCEMy6dojl8htKpT
tFD+YNsMFbYAOUQtGQiqy2gOplmZQ1HXoG8OV1A6k3bUSIy0KciClrx29XbjOCfF1hud1BGYsYpm
wcpMUhXGfckIOk+XZyXzWN6ykGzwmQ2Ripme58t7z83EvrdFTY5sA+NfTEF8ZH4zJ7OSOjP8+veg
MDyMnkTQRZkgw0TQphL1I+wq1KP2IcDqpJmxedkgC32KYE1PNg+BdeDJXXRhcwlYbLNGhk3q6dvb
bVjO2yqyOR/fUPuYlX8GMStZ0yO0LMwCD0GRlUPoZWzuIFzj7im9VtM7TI62aSWO7Au5+m2KSekG
P9dCMeLBpzELn7fipMVrrSfMM8ehdML/ChgHnoZwyFpFlVYgQxeIO0+IvuA01vBCagvxHn4XwR/z
dNkJPqBAbrefBXyEbKY1PMDvSBU48NSQDX5q0909n8gujqZsnp3sXuu7JbPshToxUnvw0vlLlcZH
rTTnMYzYtTc12kE+5jh1R3NXk5WjKI4vo1+cT5/4Vdx3rTJop6zb3Kw1Mhewa2YVsKkyWRixhxbs
lDZdEerVCbqETm9AjGBd34mGTO0DX1pmSaXO1lUyZ/UJ+BR+vXpdspVOsjv5ST77yytrTScAB38f
FmTvcDRBilrLxmSM6RNEcVzwH0M+amiarYBWNi6ZgMifO+kKZ4c+/v/KCUCo8DNNwrNpY2xCOGVd
y7pGpSe33dHDFD1e0j5+3gtEC8lUV7vGP/JoEHv/l6CtgyQfXd+5++x302p7u/CKsTNdwl5rhxV4
fSkXVtsIvPdIN75kzsq7vwTJ60NOO5eFEclMABx5+Q5dFB5oDvQGf/XwywPAMx9I8DRX4PD3/q2P
GlOeApF4lG44x2fTX13IWIStasrzrUvdiqvYnVnNwIEonp8lCt4dzkq7pWwbjMbL2OGtYR1ZNAd+
WfsCFmXBxkE9rigTA0eGOZhssE9sWcR3i0LR9yn9FT96DoJnKPN3VbwNS+OQDIHJdw7edHeaUa5v
pVyKXnK/MaonC/Z54GCrD6YHWLpQiJMBfRuOCadoXO4xqrhb3VbaDOKkRGragioryYqbFxNS0IiC
f9wvHdgGI4SVHpQfgVd1LRhygttWnNcXq5Cs9MDbBHQoRIHZWG1BvtZrPOUJQJZLEr114BiLXM3M
8pqwC0sYSAv4mO74ELLLjRA+bidzJhRw4Bv1JoVMFfCnj+SKspTsiZvlwU4kYp+qBMjHlZNvm728
q51wlFa8shXRetoA/gpnkdyMV8Fg66a1duZ9UPoI7LO2PFr1PDjubAUKLRcVMMvUJpnwg7WPp5oe
UKj+V+zcuzor0780tAFz7sn0DO2FFb68myP4SIQrESr3DqmEFQjzfzZBMyF7PeLrULe6E7YUG8qZ
kpguwoy9FSB2mDVxPEOImcIHVRHaHwROyUl+DajEabspj7OUQDJGTJ6aqeWC0wW9NdcnxB2Uxcvz
o339zZOOPEM9ENqtr8a5+Ct+l9EabgXUtXZj8dvobI7cmS7p72Z+6RJ51/rcWGOw83HX3Id0zwvD
JzqQKSNKLzC2C6kOfWY8F0yQDZ/ezAmNa+q56tKLELCvKau99EHEc4o8bdZA5Oxd0JxB0GQO8zhA
Iq/lMUceqYwqQoP5COMc+7VXdS0+ovCp0Q8/6qCqBnN/StVOWQrZ7HHrQlb0kEdIeIjgfsrL//MD
x1bfp/uo7lrQNFkCOWzf00jDeqgEkaJbl1mU22n9CiTu96OJ+iTouB0Z08TXf8rF2PYndiCs1NAC
NG/nVYCjhd7yforv9LWSI35YBG50PllzTUbEL4htBpvZMNW+HXlb2JviTMllS+qizS/yObhpgQr/
uKOu5Snip34+crokxXM31iRH9Fle1RGzSjye43D/AFcxCNAW/LMfk5yyB+idXxEjQ5UKMPBdxug5
/vbKvn3DCmP0wtK2wtO6Z+i30PgD1emj9Urqt8bvLZGsL0Wo4DkQxAzZFwKbiBBpeoF5oOfr/0C9
eN+HwuTJda8MYM1FxIIw2GoT9SVbUXfU6qW3omq0fMUStMoyW3nnEgL1pQ3sK7LjLZF9C6vNcOi0
Wp7UtfwrKusIBfZJjFAlvymkUXEJAcXmcotNHa3zM6V/KR/GcmVBlaJ4fWdHH3mwodPUvsADmQWP
ZMnMZtjNUKW2ncaqFGttnWeupdAw42qsW6CpbSVFoJ8pO8SF6cuYWh+bEeZcrB6aRF/Zx81MWQDm
8sV/G/E52BLOjDfHPXlpidOPWYXwWjNqkmtfoGn2bCIDIcabp4MpI4VoxI3wR/fwvIKr6Nqgk6xN
b3Hd1PJLKDAO27XD9iMrq/6Yt2MAt+Jimo1GVyLK9JAYia6wMjaw7YGsfC7oSBm7T9ubT65csCrm
vASzCJZ9jqdFC+8vhtMwybgblhwLUNGggxbRJkaVFxKW1kSa4qO0P76kZz5ffrP3icolJYEQMW9X
6YJuxzMwziOBXt45TSAOUJjebFfHm0wreM+5ggmR0PlRBAi9I2RbvLl4jmVtLXHW8ELsEmrXMIEp
5bE2DakD3HWnsDmztrROwqvCTlPmGERR6jmd4no36d7Frv7kZYK2pHA8BdLjM/7OerTn82Y6sq9h
1pYf/hCcRS1CGKW8cOSETc7++AAbzgQ2omEJlGthLIx0sv9ik4f73L7gRrM7ei1ZErPDU5h48y7A
hD4nSDI5lUZvcrnTkBhQo/F/QtoTUiJo0YwT628rxEzo8rF1fFIfgoUzdotjcbw/g3c0zAXwjphI
wiCw1xDzp0frSeBVCoq0tqYcued04rpQAEM73QNxxxiOGm80sBKMejgykcobTkXzFJQnbgkQFBL7
cSB9t8bAVSux+j6Ecp8f8NVEuKOPgfugNEJw3sYTJVBZaGvVxE+eJZ5n51lBD5iymeUMOgItq/pv
FyQxAR4OCI5RU1gHhy+DfDyGStZ0AMSr8V6aC6LuMemEy+Py+PIO69MtG2m5X7Ms5yGqyfXcoXCw
YVPy9Etpmaxl49tX8bdI/bSpmQ60PXFhczsoFlPc1k0AQC7s2G75eU5QJavDi28FnlCPYjsJcTsK
BAnvwlE/74+poNGHBF8vJAKSTMh6xfZYTvFqm+h6Pa7aUziDv9xWR4s6WLNw5NKrPDnkjDi2jY0s
2ZmxIfDvTfz8TS0G/Tpt/6PO08ekXQkrAL6KMFyiuzIRpZ/FG1l5XHchoqiTy5OFYhbVVmhRQfTn
aM2r7Dgh6TSF0FhQDzsem2obsxvjtglS01iJbqAzzgT78PN/1IhHxXB2wmKAUTOljVvjF84sAKFW
njp1STFI1qceJogpsbdFugSrJfcAaTD3s/B/A+DQy77J+paQUC62aug7IUpB1JgzwjbqIZbgESki
AoOPW+daNs7Tw+gx+S4T/DwWbbgz8HmJ7OKz7v6v15K4UhQjZlUXOYObfMEfYWgI9lhsUDEx7DfV
D81TOVrMBH13jE4oEjKmrwKcVWluMN0uB7MihiJF/y9Zkp0jM0+RTsLRzDs5oU1d+gJpBHZxmsdO
1DsSB9U+63Oo1WGwA7TAJAicX71Rw4mES5uktfnkD7Dr/WUD3e+mbUQQMfQGNwGxQdUKaH8Bwv6n
V//vrywhO7xE4a21T6TRWINJxt0fo+R/na7c3d77sX7vz1SFinqF5jpMJkWlkktw0ZBDfllCOrXd
HautiHnbowyI08KSIDz46ZDNGCu5fyzphn8f5yqRlS/uKYg960rWvUoaI9FMi+0aYn/5UsEK3igI
mDqL2yV3zTWyuZ+SR7PXvSc8/Inm6sbXl9Yo2ht2pV4sL+xsva/gh77uIWkfG3nyD+nM8cBFCwci
/TJPuYpKQIKvRwuPb85NDQwZSmBSogIl6fk/FFLc92qYkiDYG03zSVvDnHJFuDKkclZTjEzcAZ8P
C/NUU2bB4aAvd2tR622+q6hT9vJAdvm+XoiI92wy25o9nL61B94yPTL80x4zUtK//q7QOfgVjrNd
E6iYOiSii+actxiPjMbpsy0674esF7yc9qDPswIj2swYyr5IUiRNPKKXQhlD4Y8XRD6+nkgpKFzt
5jhh5pBSEhEOz/mQ0+ZrDO3XOG6dzghlm1ukX62BJF4FiwQ32kIShZu9B4ut3e3XZgXsTGe4BW4p
CtNijaJmAlr8eYhcehudWxXq2NiC0C49Vo7x9sOU1sSGOzptaj/i0mG7EsTr8OOhZUG5ThX6I29G
fB1R9KdRiO+FcEn4RkLNyp3vj9G56nrPOpdjycRY17feVHCBwvpaxMtXbe8/LWp2omH4yj4N6WFI
D25wn80uNdxbLxB/yV/yM5iXHs/COEWLQwKRt+6ey745WBf2OkQDa92zgHP0XuAz8X0FFuUMFakr
Vyl3DnFukEJp2UPpeAcCP3Og4M1iAF+MEpdQ3NBL/j2IGNNWlPlPjRj9FOhPJFk0M9kWr5XDzA6R
KCRMQSgMntuY7JtkPnGJegHxRzRyCAdSagOnzig5P48V1Cy+BkR4IwFg8o+B2dFr06Fw0mq5ozuh
H3cko1RZi7kMtJpbh3S8rcP2256/hlwIYMaKqEonpRa6Fg2Wuz22/HaQ6L48G3fi7yi0YHU+b19D
N5bL7fvgnEZSWzH0Pg0+1cKm/bn4Xr78zi2OVSn1H4uJ1tOkfeign6pVE8eHVN/rGYoEKNyB4aFw
w2pkq+yfrzoExgT3glh2bni6metLFSBUcGoFUhfRg/keSPyKbbdLggtrN0DqGcvRIrt8KcGXIJAJ
p56W+uBPDDzTfykyA4nWTKLad4az8pQvN1cWmrd2U/kCRZkVC66UYT3/rIXyIYNpCmOaWmrnj3eK
zMdnyHWNnxQS0mdCCuSHo6aRiqX8wUtSXAvGWMAVKfJNo3IL2ufjoGS3mI0Q64+MQtmvKarWunuL
BEkMgYh5B+mo4Oz8Pil559M76+k7iABhvPNOQgQgBqxsaBmxlLJy30HKCk/M3l/l+zFHL7KuwsSq
iRTIqeQNczF8p4onInTJZ4xuY8aTSXEw6skrUq3ftlfdpsYE5RWyMUucUZyV3v18b5JIlExYbbFb
6C+Iv+Iqhf9jtEcbJqVd/C+KrhCXRzyF1eFpq15VgArhTLiZJwYTHVw4Q4QrgEwG3qO6Ug2Rc1c0
9MAavKIocLl/FUjfKwdtRw+B148fC8/KNY54zZ6T6Fx8RYOCPIYGpKQJdK7dUsYp1UeM0MqXv2Sz
3oXvS5CXk54RZ2v+faQHel18ntCoLYsy3jQgrajou3pALhHnv1zNz4l+XRHFO2UEvvUKss2ImfY1
TWBY2AZU/pzjdBhTY/S0EkaYmjqH+1VaJ4CXAF7iwwtWZSFebhvWMfAW27AHTOL6tUHAD3jtx/TZ
Q8LtvNzBZWcWAndgf2RiyD8iF14Tr3XVRvGxGdv/6qa0oOifYCNZfHoetWPrD3pVNqSSnJAqH4TN
Z5volO32BM18IwSOFO9PoYdjNGFRQExIEi147QqnmS7pk4xtel2PwPoOPLuPXz6iPbuaKwnEVANB
mI0XjskkvwHQiB7bcHjJo8uIP+XW+wqbJIHNonKp5g39qKLzRqI5isU/XWDY2IKF7bEeqORvKJdF
4YGiytcrmFmEnNeoUd5sYCew96XwpHYqLplnSyGZ8t5i1nCF8oTKnNwmKHT3OWXI33a/IRtjxFXW
EL7qPDJFOgc87qiQ3f1VEDOf/wUFf++8JIEatbQlMZbWn3BOXP/AXafKIykrvtBgNV2FS0Os2guf
xwbwOwbrDH0zoTEtZtLt5glm4etHKBBlKsB8ct+dOewcFwthprR4O5B9+HQkzjcBs6y5uQ0x+p8z
GTmmfMP0MZqHhFy6cx+T6dkzdxrl/X5A2/yY6YtAMoQ+vvAQ1LjqRij+yYOfarEfI/X7/gTGPcvP
iglxyjVeEH/aRXtvoBhNh7vs2aPnaz16cjhqfK/10MIrS3LylaDxm75cUdIhAHSzZKOmB8arDXK9
3Sa6dwbm3ixE0lzDU0OSAv3pmj/qh7UmbAyBMDtv2hP6r+BNHDkcJ6JYImnU2XWKZacutYaloLUu
jKKGO+s52XxxVm6TCasHrPI2BGyC4TSg+cq4Wj3LEyuhUtU830iM2BdD4hbbywi6JGxlNYWC9h8Y
4+1pLZjHhoJIyXyO3BQ5sr7I665Q2l5fVUcCcS4pB20Bi4ENc+eWF7FvgPpflG0sLOe5IDxQgZn/
rydzfi3+oITixqww9qJTeDydfnT4XD2BZbN/OYKaD8eT/xxTRa7JMiTlCDFiUBTwWs5b2u0xatnr
poEIoyY86lWYSaq3bvU3INtdCYoqbUmJg8eb0/c6R5hghmk8hURdb66k+iDFtM50FL4s2I/S6Mh6
i4MDRNWniyZTiAvpRqy76Z3dCPKReQzB9d+ZkfgnZSzDeCJLmjR5t8e/yEiLE40JQVmgTVd2//za
Tb1XXSEJ404HhZ55Hh2NXO4NQmtU6Mnsy/iRI8qRMNeZimeV+HXYKDzAwi25fdlm84bZjukOGWdN
PRn7t/+a41UNl9wczFvEOlaXbetY2sJoWa8q+KgjwBkhJx7Lo7M/YtFaDpBeKLHyxVJhQG7KNEjR
KcsGb1VMH0W/C6tBEO6aTFeFf7RXn9ed/7G+cylyKDoYaoyz9KqrJX5o0IsXu5jGJ4oDjQREgKkN
BfEJE8ZnglbE28656u0UvvQUQTj5ZCfM0Bu1IJVjaG3EXe6G1GIfl/2M7qzxsBs9RYeoe9d8jiOU
AUjBN2HvLF1HWGXiZdAfuNzuh496f/2Cy9oU4pChw1KvPnEIGTlEQ1VqN1T6upd5SX72vBEanHgm
ElVBl8slQKtr46yaVmGx3XGkQT12LQENHElxLJ77VIEX75AQ/43sOWesRnRNuzqQv2bZLXqy5aor
6rtCNrtxhMVy3Z+bebAwqvI6lDn+zRqVQ8SiKI40wQR+mD9W4kR6Ce6sao93HFUWqmTFUTai2F5/
VCPyHFLlqfpwdg6wF+tLNJ6lZI0Kkd7kO4LRw8FZUugB91O3XYRsD2o9J4SAegA99LRQDOLOhYPz
r0Ea/4GHx5qwdeP14oNN2CqBzmrT8by1YjZZOS4i/nPgnSE3UC+ghRCNm1Pqbo0GcpJMFYRhAzaF
vQ0sDLUJykws2NsWFDZn+ohzARd81Of10ncoNxVF9p9DdC3qAzuYUK4WtzO73sqAAPY74A4+0NgQ
C+XVXWklyqzwV9VfLDDDHijDmxQ/V6zHkr9KmwX+Mh/7gQkVeK66RtjakCotPt9pw2BF97H2OVeI
BMeaGoUgsNo6133ZPL8unho3hYxz74XrgpVk19+Pp8InLjTCuo2hVDpQBGCzk37WcP0mnaDaqQ/o
+wfyhJbyhxuNtxZc3sMKoQpXxLWsMGvE7EE4wYysfCcWkvHuqT2x79ZhI/HWH9Ib2riSy1rncr8W
i1LB5XjzDWX9Gzv55kYpRgtozSH3ARijiKgc5z1sPwoRTgudrxMBbtMC/RAAAMoVZqtyt6GB43xb
MmBArkTvGMnxrJMCE+HwwBGqlPuwbQY5W7bZTUatJgNyfG2wk2FQ/kvTG3yKjxt+nuQLw2uHTCSK
ooO6c7B6+x0Vj/2SpblGO4YimfCktn2pPLnYKi7wJpX/5CLDTofjdcVfNyi2vB+XSg+F3MRw+R5F
W1u2z18ZfOiP1AczE46SWry9czWLxIwE2M2Ma7YhT2ZKmfSYNS/de59CJQ+25PjDqgI3PF/lyp3s
jSJP6rgIT13EB+2CL3eg4UPVokSFEGGwb34RmNfle72OJS1BYstieiCxoG9Zw2uUaZj92Q0ySsu+
PSGzquJYNB1YC+57Z7cp01Ttkq7woXLHZZtcfFp9OufEsW1Z8qlQ34Mg6R3lbsgKECTuLPiJUJIu
snjGgxQ0unY/z+gl5qv7Te9OW+TSn2SLziJAPWhGML9prlQqvnSv1dQ+j8wqZb2n06aXHdNsU+uV
koBZ66HmsvjnE2VCHyTF6xDq9Z1vUfvSbOOFRnmRKeph6JL7R9md3//s1emiMK/BpnwSb+lOKvUx
6/GtN+Bk8mCf9ox7meXcs4DLpcBhHfhINWI2jWT9EYoh0rRWSb2QktKXi/L23x0qbXKErcst5bNO
B5nRd7LxPa64u7pf+ikm0liGkToXBypoZvfyUisWPqXMhjdbRPbSbv5AwJMXzTms5CDqrixHNNkL
yuYzauTlMksivrxPFeo0u9zXrsYBIZqDWI6evH16gdNNoclhMPqiFeXQzIz56AUwElH4HErm1dbE
0nmr45vyg+t4q164+ZsGQGW7hiGxXDs/tSVlrz137vHYr4QKSnBKzl77WgmOZ/a0pE40f+JP+EwE
Fl8trJsSGPfdCix/S9eBx/pm4NItY2E4LTPR0R9rFmk4JWdsYRkkcCQRsZmsncKlJKsUeLfqfUfJ
PkdlB971AJczUkfWIg/0pd8qmSljNvIvgEiQ6FqqloyY93QkxVk8FxXjRDndxnA3RSi55zE5Ll/T
thn8kl8zv/5EcdEHbwv4qXmgtIYHYUGsYsIUyt6feVSdn+yGhbNus+/FCBd8WlquIR9ykNm3nmn0
bHvrxx4eOXrzK0DBEW0DlBT9IV8/52ViSiuQbJ106JiAkc3nz/hBNVeaPC3Jr5EeeGbRPJuUJ1eQ
RryXeu64tK+ue56Pxxvib+1mUV3bSv1zez4+ihBeWYCr67tFFlY1Qh0jcVMNYPR4V6WSVBfG+cSC
tIS6j8vUJJYD123fOamb6edFyfWDCDw56Hrr/Etufzn/ZFLQmbJothL2d7lFCgQqVagvO3whpPgk
THOr4Wmd0L5l8N6yUhhc2Bk9Jy4Bj20uxrZTPIlpARV+SJbzSSsHgN23ZJdWaYFNzFX3oH0leAga
rqzaLt6YzR7lKOA/NEd9sqWMVIYQCSZ7FMplHuxmowVZjZhyFEmcT+hRAJ0qF69Af54lsVhWn+Cy
qGk076CkkOnMaIupznAHG/xpT/NRTE5dB7pZLYzrluKiZC4CFuNTy7gY+GiYtN9JPzCmKX3Y5sfr
ie9WlD96qpvcFppiUpg4FMA5eZWjERTdGdwCDkcb/7pgdX4FZP0O2YnRkJmDyMt2thLxkOFpdsRj
wHHxAV6B0Qw1455dD6SEHPCbFSB+Ht/rfXV4wuq3EdtyWS9FG6PBHGs5hTIp7iazrHG6PbV6dthO
41nRGP7L90CXix4EiG3bM07pjg8zfLTWdDOAYhBw+eaiouLZupoVSpWssFb4h2PU1pq+YZllvRHq
923PEeDxJOKcsrWYS2Rq5F9LPyPPv9R+nwoLzsbfPoi0A7kDo0w8bKE9V6bOmMYxs2P/hPR2lFRP
ekgNi63VoGatj2KWdS+oRGXDhU7YYuS05lVj1CVcaizWPAO+2zM766MHhyj5TTKTmuzB2yYHjhA7
6qh0aQPTsn98zgW6ofB/QQP2oeD+D88a3m+tLh4QFEBXTu1ogVcCricCc2RTaTmgLrmrRr3xAKV+
7H9Yl7KG211YPggHGqxcij20MpT00OqOgDhSa7sixYUlMq2pipewHtIMWPP7hGT0eZT2Hrcjs9X5
S0PESKnhNoOa3ntaIDdhHwaGjkJ8SGjnq3IoGLomSVFipNcuE2H/Mqli7I1v9f4s4JgdfBIWUV9l
zN8bLpyBWg8tXvJLFFl17uO0C+66D5ZvIeL4uey84nW4iXvX9ktvGNEEsH4Ekl+6KPO+PCV+gWes
usBuEJA/8Fao+ncU/3N/Hm25gwFG5kQ+Cy7O8ZhNnkPmronrTykycwsGHDaDnhp28GPIeXJPSveA
7DPja6E0sBBV+OyxbCFviatm7vlwCnyz9zX6lNMVA2ZbJWS8S3yurSlqlRw3zdX2Jveh/y7uGwST
fUOPhyb4aIyRewT88fJ7+tHymJswFbO2D5Aenf0khOItr30ETQpURb0o2EkXY5iVLPnF6jcygkNq
s/XieOvqD6jwVECIAPyVVucXbxAOL0Iai00ktW5im4jeIYiRBD/5DBYmwoW4IukGyyYwxejXnvZB
EJRBDpPxyHIRH0hdAZY3YMeA50zXRPgDia5VNcnHRLynC/UDvJsn/9XJRhpAXQVcxFqYpjZl9Ywv
a8DvBUCf4mfwJgCImXSNm30LyzUrAgrktcoSeQ2u6dMq3NwDaVJIVcTeZshBMbP0wQ+Np3SDjbev
uS0/uj9XlAObYNP5yFy1JqfUEbbos0jqRVrAilitUd2NZNQzMU1XLfaDrvky515r/1vpqAfjzbAc
I3W1b1ZcCHNdSlKLLRo9MEA5cOWgwwD2f5Sg1MUVsK+Zn1cvJwfoLeFQL8j241VTgBTunsMxs1Hn
VsyVckN1eowYQHs4W5NCdlIGYhDvWZhZJ4Y1d5ar40EcihkLsCSBHTr9xPYdthpLGjrry7o+Q4bj
oHMBww6PvJ0Av6cRdOR2nd4vcgxorNN0ie+YlzHrsv5Kx5NbLxg9j71NsVSQmabUuFaOZAqQFoE6
qkEGfYU2nAz6dTUSg06+DbYGJBnQGQezDlSDyxy2fBMVACegvG8jJSxabW6Mi1zRYpV0g5R0xnjF
vug7w1wWaW2eTQxkDYJ1dm21It6kj8zzDS2kPQXeVJkySfHInkICv5+aph6tMCZhjjYHZMkmuMqq
EpVW7x4TdTz/MMJI7b2FBocZ101WzElS8SWqOuFkN/mA+7FQsE3N+GwgndtmHtnmxNnaulrUu2Fp
c1PglfWNwUgCFGvhW1GiyRByPj9/gTrAD/Wjv8mAAutm4ogbNOara1En29zfcu7HBN3rQ07O8dZF
Gf32kld7sAXA3fL6hl8zkIXHBn6RXLg0jbcPu3yKfbQ3s2NV+KRF8mMrPLF/bDPQeCsNKNg2gU9l
Fg5JdaeraTBUNAnyNCOWkaAB4wJYpEw23SuW4o4/2JMR6o3RWS9yc/llmKk7qL7ZiGkYbILZriHT
lcSCYLsGWntBDls8zrB0Mb7ZfiWB1mJzS/h4UorBQSQpuzhV/S5QbBZgdZFgwPAIC+TgiOOjYYhQ
m/n4oCWNQVM6hhgT3P1yYxhTRL5lHC3h+tVmGI2/ETTR4uW8qztE8k+zMMz3an3+5fJQlrnTd3Ap
Ea0dAs/LkAZUFM5gzM9wvMl+fGpJLXbdf300QnkufLngT1NAAetIJaX6369qwAES92n1CqBMwRCy
Ks+3X/8GBP4Ox6JgNWBHQiZ+qFJh+3hkMMfjZcStyLx8mNfc8rBsq01OI6mrwfjp5EusyM3jSHpJ
DAnq9Sfqrns/qEdR4i8Q5Of87Al6xU9mj5L1ne2+bZKMKk0trNmkT5cd+a0uyEXn+96EeTnpZ7vX
Gdo9Z+spGHXTAPwvLb8f4gKl0Ow6sIUuI0imzNjJGL++jlIJsQ6MB10vhI30Vis0njsyK1PwU/Cb
bNhAnyIbWPNLRpWayECV1NDdDFj8q+X3ts1Pn0pB/yIQny8HfNBWAaYXsWvNnDI8+2TU3QZilT6Y
+UZlu/dvP/+FvfS/aX0TeMdnD7zDQS0z+6z8HSY943UWhdGyhAP1kZve/oRN4VegS+ZDXEd35Vmy
jB7ap4qA0kzAUV2/iu8fwOAr3G628g+aw0Ik4sSnTtjX9uz1mGfdjRYPWggTuQkxbgFhEAqL0z68
S6/3mIbFnVpgrwFDXQYowuWwxMecMfisy5i/TW47jzVBJ6o3JoK4PxzzEQ2cqLByRjgef2H1ET3d
mOUrDCtT7c1J+qFUDepyjHcm1Iv0zz6/XWfzxxrqfiH2O0dCEUYr9ucfr5nmzwWRWTOzAIh23cVz
Zb3k+fytYD9mfkQM78Su8o99BSfRS6Tz19av5LOZY5oduAwc4bPzWcNDXaUKQzDxxfchkJ7R0Ns9
lDPBfUDcJJoETVhkl/RbIl3ER164z+4yrEYmw6XRRzvOwXY812/eaxi+aIiHROSNAeNr+w16iq9+
7zitoJe+aMpEHAQWMXUvVrSUMcbRACf5Vx+fz/Nz6p2qkFpEp2V+J67eWiDZPZYRYdZcjOneRBuh
My1D6KduU9Y+mDyM88gbsATvbnsAfHMdKLxVhdogtP/8ADf7v29tTXO6B719t7kaNTWXSDhs7OL7
zKInNjscqoyhOBx0CknCp2pBsu06XUw6tKTu7hJ962OL22k0VHzc77fJlBnZ/cxx7zM42SlePtQe
4T+f5HIoE6qEPeXy60EbiD1BOgDX6F/nIvvl6UfQ3j+dSIKF2pBH2YXntt2GbQ4+c2rNeZSAKBo4
v8gytMraLWQ5Oc0IsS4369KlI967lJg5U6sDVJMD9IzI6BrAPi5VJuXDKANuEdoH4iyqw6KZG7JG
+daMPpwQcI7nVZBdbUJQ3qHu/GRxY6ZeT4HAAgglMb1Idb91NkiGNezKEDoCD0ZEA1JjApDPbW3h
EJmfFA6PSOZ5sBuPl1AOy04Is8mpqxFOviqMzgj1p02ubrJF3ChPsKt5vcblNSzEO7p2DIoGNOPE
oJuTAXnBnHMp3BJqvfqervGuTNumVCYZfUetBy8gCWHE9VexkY4N7gxYk4LDu73grprANR8yms2u
lDQpN2SZBI6G8QkP8KNUC5vi6CXkYoHdI08P222CnHpf9w4ZtVLx3ZfirxY1WKrvE/XVyHBQe8+p
ncOJxV3/3f0jOsRPHjY5QBdwtggUZUihb/+lgx3b9qAsWxam//1yk2zcgzpX+9Qlws0tq1WpamNf
2Ix8jueWNR0ZKmQ7AURmBADZaz5XZS0lVUIwjxopYn9muqYglzWYwcb84kLM0GxpSPoPzjLUMR4E
X1qdXcyFHUa0b94+Pg7haS+ZQ3Or2rrLMLu8te5A4iEJUBYoc8AwtsefqVh9L9ySqqhC6ZvRhSEy
AWX1qQgEgZ32+CID9Uwae1bsvA1Q0bsb2pvNhD2T+pfZa/ZJQha33OCksT6f0ies82LGDrKNSvoo
krbN6NdvPJnphgSnCLgHVXmx0FbXwwtX1F7HLuD4LHUW3VDas9Xru5l3RzLugWcGBWY5v7a3jvsK
+wh9bHbGtGP31vVYNRpeZ2dU9jZOQDWLX3p6pxcNEx+TVOoTqX7HYVgEYM0WsmkEBsc2Nl/S0mPN
qCqFshKkFn0GZeVPEcj1Yuf29BK9RyJglmJPT9K0ig0Ko0BLNt8ha3fukuqyenODnskYZdCgEQSP
AoNzIdsoYduUmkwrgSYYyThbRwn4CRkB+dC1fNCiNZKzHOJhOnNAcu/r9WFjWTWVm7Ms6cE5eAKs
OplvQPg3XbF1OaGqf2p5lPS/agiu6CmGjriKs/bYIH+NXjbal6oHtd13o2gs+ptRLUDkuGppS2FE
8uxfNPWhUsk3TtmWHf3GKL+Q3cV+DMiG/AHc0pZ85pIYOTiEFA1JWwjDNC0CSxwKJDCsBxzIb0lw
mLUdyCNzI23a6zp7fxOvKpCRv7MH494OtndocgWZZ63QNfftx4IoqYETgARojaHYrT6OVIMy8pO7
khU9/L81zmC1IhOaCS8jChILgBygycTeMblY6+eK1U/V1juyZOmQ8g7i41R8UZ8PX5DbGcv+AyJ+
Bsig8tpHXY5PkPuFeXdwv9Ub5A/JoOOtDqZDaOz3UCbc1HkxwBGS+XH7ZsrDTIMLtfDbzlj6qDFd
iQxHWDms2Mxh5SIAZe8q5qwjDRDTCsE65Lybsrdo2mbB9vGvDF/+KLLey7oKEnc4kwumIWKzCcXm
Dc332TuQe2LzbAbDeMLorZ2EPcH9nI393xf/d9FjkkLa7tH7nr6+zNa0OBOUH8ZiT+F7NxXF5ZUx
oQ6yzXOpqcI4D7MsvNeDlQJapcz5yCafs4x3MADzTP+XyO22oKfh8KXBobGD2mSt8OQ0m9tYGPl6
Mm8jfBB+qQe5gytaRwk/lO6os1gHQYnell6MZtrNGY93P10Al5Hl7IZJne5y5TcmZNvhO05tYsZ5
fS4PDsXLXYvlomWyk0KWvYZiDQycz41kP5lk4s8QtD/D3FfCmr3S2p9e0EGmt8P2MYNkqraw8cq8
YEtjTfmp5zWYziqNisSa9dxA9OStLu2A2htIHJgi7oKDouiEZVKjfcxVfVRPMyKcqdaUh2rFhW2+
fcExnAyYW/CLVka7++XFFLQoq32eLlWUvP1qmqGZbZEZve/tlKbZpPmKAr7TyJSyGwcGIBZvhZy8
K2UelOHnBHMsqtybLuY/z1kEcjtl829aGQ2TtMnL1ya6GiEGkVBbbF/pnMsGuCHtGe7fm7uzpqiP
etP4JmJ0E5clMudUcrXIJ8rNKXIczmW5lChIoUZtXl50Y1ZLuWgxjC0OeR5dYQGsKB27S74XeIYy
rKZF5qfAjv/TdWmFLLUqRXkJvkwSxTO1Z9dx+k7eiRS1O3q8aogWyTYHgrgvKJl3+Z0QmspUDJga
LDpTci8KwKg81SoM87jTlDvyy1ajqeHJMwmbaLg9mOqdFyUEgNqizx6gnBdp7L6SGbDi0btWKMeg
5dG1qZTi/PPIfbAj4H+qiFs6zB4NUZVpN7nUphhGr0W8aPWat4aurM6sBEOIgGeR04Pz2eoVCkAq
wlRUFUsavFyi7Fzq0kSYFyHeIZu7leIBPdAz5YErbeMNa0yVMKws6bLjbGNSFITsxdx37p8kFa08
9WoRtq6XZcKGdIA00vpFvbaxhGVvSw/3GUAG/cMpXCRZ0jKBoHf/CK9Z2F0AbASIRHfTHuR242sy
4z5aDD3XYqc5DoOQL7V5HWKX/L8gdp5GCR9McTqlqOOxeBL/sqaqYK0rUw+em239doh5oLkcP+yI
r0dVTmI5Jibq3nRWRQVs4auK9BE2MShq1REb9tCr2qBsDpmcr0LZGu61gRUaRgykMwfxEQ99EhG5
DE4AVHd+0YmlRqiURWRNN8wYmfS0jBvm9dd1IG83jkOFrZLOY77pdb47SgY3epVnYA+/aVZ9O9KT
ydn1g0n/s9b55HsDqR7HoE0s9y+PJm4zYdOIDW5JRYRiz8s9MKjbXv3F/SY6niYre5ksujKcScrW
69Vuq8EyaGRp2GwrlXMw6sUmHY02ht1TmAum+JD4oqloE2Um6Wzwq71sT4VAd2PQtR2/KyAHPEQQ
v1Byt5bApXpi4Qc483IbZYU94dCEnS7AeF71CRGRrhGijaKraIBwoIP8S1lzrDUJV+Xg3E3xopYb
G5eivu5TtuJ3P+EzDj9J8A5hdYuZz2cJD09H79r5LKgVe7vxHHYnw5SJ9DxvZ/nv354kwCBWHs3j
KUFnjq2MEA929SR/vLjni8PvXiqutEQg1ffskcnpbgQwqfk89LwVWrZ7rn0buD6TIUsN+ho+131N
0NCr3flEcVKYHYm8Zzth6uGEZF9c/g2JkXQDuPF2bnp57LEzj0Xuai37D5cnv2uU8bEK5RkA4XpO
6jnsmZlqrYHzLj+W+yRcVsGgjIX88UIH+nE7ZtVBlJcnf9elDuz3rp+cFCxLiBXIK0nbNImlgTQb
24pZs/KDW7dS03nEkzE7BuRBmjcYWna3Um8YvIdFoJD7/CpboEBmhZ27WWgEIpYETmhKFcA0zeY2
MpbdJnpMYEkjzVJXtQJMBhMccepOS8iL48Z9I3of2NS81QcefPq/yD77XOF+LE7it/WBhq4fSx/8
JI+FGhSNOHV63iRHpdnf8bDONN8XtejKmXCNzsK7lhaWTN/u/ncd+0wx3IOcl7jsYpQzc4P+HBcF
r7o5aGPDIxAnMiS85Gatr27n/NFuRrgKakG0CCJ+HV1FWa3hJAvStwaGWVYn4erQzBVuZAX2TcuM
XtJrEHrJ/CLUKbYbCCXAeInAn6NbNHujLzYwnfM6FmAh1fo4L19oCenoLYlOPh3XeecL/C63iRsb
pyvJqvhjwMbbK6U4Im9DTk3lcYSN8a0jrD/4fSulGcnSiuFD+yF/JAbe7XDoDuAS+MqzlR99yv3c
4EjpHp5SH/mOIUMPeLK6t47Z7ef9ii8PJYIxqrOqiH1qKqB15fDKHdc0ssoD2WtHBcVg1o28J2QN
NioQKve6+srqXX9p5xH3Md2bFBE5aGP2FtU7tH3RiqMknllq/WwuD5BdcrYJibn7iFN108/H8WCO
ZpETpZNdXEkJ6LVX7WRILPnLznEFhttIlCFbXUEfgcPNpZ943IKP8FqPUTFNIXcUU0PpG5ULAjor
1QGXtbBCWS1z2UnEOAXGxqXd27RopCaOzkKWBabUtDp7YdvGB4EdFPlOOFwPJJ5Z+JpKIhxxNszQ
lxp1gNkubUOJP7kMUB5ghguJBJl6/guBy7Xy2baWGS9xWD2mlCOjBOz1a6TYuhXGVmme3WpexVfP
ET01qbYPUw75XFd2M+ycDfyKDx4xG2bVMyfP2FMFvqg37Ys3l/WhkNN4qIedNr/6qb7DQPOgH51s
p0abD9rfqMTRwyOrqZoYHZEjxoYWnsK6QLhxl1oKi3Wc/UZg3FrNBethPps/e8QEpriacaY/nH1m
3/pv9xJktU2Kphvvo4jIUYSTaW/fzA7s3VqgNSHadsNQhHDtI6jUmBe+xluBwLpkFM8IgyminmPj
2vRhlb7VrgK5jqK+zFbOtMdjnvKXwRtCNf2kZLkAvEALN5GCna0rPP4jm9j+B04Dr4fZJM9Zcdg3
rlMKZ3wGP058WsmpWRR60hi294TVI7VnxFgbElTnowx3VuVwOK+I6RzD2f1Vk1wnYypzmNA6C/Cc
8SdQCdq04t2jX7LJEiBYG7j/BvTqilhYNPfFHgAs1k46knPtib//WtUP1fCUNgyXkUnGP/WcFCuW
qNc+bjH2tlzg8F5cXGJ6vli3NdVubEETSAMjxO029z0XC3WuATW5myEWGhTi5gIyokROdD3Scxvr
cIjtvFHJSDK7zeX6xv69fQuhJuNOoAoH2IYIWSVULpAVzx6ORSVYo66lHsVGqZwsxHQL6AdCHI6c
u7cifLH4Oe4SLiYU0JG/0JPyjf7H1AqRCjlSKTFkndYS9zQK4GqRDPIRqs6pFbBXSOPD4ya9MZgc
k2YkT1clTJFHBokYmXzquSKABTgZOBBE9sGYpmy0U9bMre0Z5Zu8Xa7vdY5kZ9sBiZrLu8Jcr1P6
rKb01xojilvn4mrY00tzT00kv+fmsFHdypseUmfBI8HxLNYILYaacdtMiiTyJ5Trn98D4eRyNia9
vOIVXiF8Q5PpCeO5ZJl2DMztynwehQYMMNe+i8EW7aSQzAsk+fsoJ3obsH2u7eBzUPifeNRcxSUj
Ww3XzJoeXBbZnqC0q6YtALGxJAi42YFNOgKBFCPzIdOBwQS6cwTh1ST93SldcB691z22vyVgfq43
6QOxPEXOFccWznbDuCOx4efAp2IK01VXRigkDg5Z8Z7buIjIYd7+xFG1MU96ZPimu8XP2KEqT5rB
v4TBULl6BWjIyixCW0Ns/fxj0LCl2qm44Xh3+iH2/dGA1elIQddA42sWL2uPIhGN0CKKYOPmeqEu
sYM5ZSu89V0Dug48zypGz/+DcMyt1GYKPnuIgdciJr5VbAc+rZTZVwfFkmQvTkrMEVlgQ+aaXB1J
tVWljQtNJDgIcf9YUICkCU06PKclMRB9+nXLYxkL9BQjWgwBPFLRcEROFSzElms5TMEIc9BrK49h
fc8CtxI19o+fWDtC7QqNSZIOYbL9dWGLsX7s6imyKlZXs9CCfsFXovAfgAvsuflUT2eIPmd4wTP/
5CHUYkmQqpVLU2dNgMt6p0++azZsyHKwtVveUqrKkPlGFhEbC/Y203svwfO7nXWaV3UXZP5srlM3
/1dBd5zIYdpF2hqjH//rMH5IYk5y0dTWB1EayXaGTfdGrfHDYJiPWTrT7oP2zjp2hiIyf4KRDSM6
04QtRoE0xDwwacJwcdbjBCWmkfAOqzp2ho1MC3n3f7Hz+v3s4j6TH2cICsYGe/rwHRXxvRVK1mLA
eTGVDaurxAJLB+H1Qt/qIPWo8CLtpCSfRogOUWeVfRas0WgEvN6fRGKa5fnfq9ptETSNJzFpCpM7
a4X+gg9gwf86eB9ZcQwNhCccAMzH0CECxZAG+KPds7IW8qg4QXTVmPUxsYagZWjztjxlWPo+RGAr
IK+TQzw81IQjcioGcykvXwj2D372Tk11ToBGPUFuwvYncKMCt7AmjhMjHOLIlWtq2zGbxzBjPwga
9k+LJDiDl+R5KV7BIFPASDzexCN/6PXEwy7r/RJaB1dxqBDmAxzLXvFvsNRt+fjHNbzlEh5kyS3r
o38xmIXR/o/e1WkDOINiUmfey5O701eXLP/a4QdzDXn8xmeHKntl1JDwq/Lfs4bvCnl3D5IjL7iY
fdizGt+1RlQNiDosaq7ZxZyR4H8+dBonILzNnHo8JmVpvoeaK/bQV+Wgc6Y+sisBkEggdAT0vpxm
7PWwv98VRLt3RnqgsLn6+yrdk0I/wQKSrqIj7O1AeAgCqKqFRwnVaad2f4vSXsa2nGKi8KSiysJA
qIfqnxwGoR2WWKXOFc1puX+aSOvFKML8obGWXfQuAqYWHWBvycR8aYcZgOky4TcES/3dZdxyFDPy
QZcwIKa2ey7EihKfGBwytzauhAl8GsiPfVC9d5d/5JwcgZQuEPU7yZaNdZ3mr2mYyoNljULm56p6
A4xU9y9yhnCRNccrsjLzOdV1q+kN9iZHiul4O88+Hlm453/0puwtrB7gNN1gBMSrLy++aWwh7zVd
arPnc6q9wURWIeoLigbfjFILImQsT1g2yRY2YydStsMCt8HWCC2eN+M8i7DwExYae+xypvxBxgiq
cr6sQw4peF1fwTtKAHPbIUUq4gUVVpuwFrRH3qUEOaZeKmxnEorcjvhhCJ8XDCWfZ3JSM47x5seq
QuheIDX8RN7I/Gtow2lAOrgHWW+VioXhqKzjkB2MSVvTI7sgtGFyXGiBBsNG+25Whtuvl6QQeY8c
tVDp+a7/cNbGzxbWcdCh4a30XezrnxF6XVYCj/tpqRjuYsmSKBrDl273y3Gd2vrZkZORq9I2P2ql
3eNB8bzlexvn6R8brmcteuVHtG5UXGdKyKUafVsA4dfG688qTRLdOwPmzX2793lWBlh5OR9QvD+F
LlynGTooscQaCxBsXQzaAohKApfGAkDIKrDVQ7G/+bQYS/lhtA7e32E/sgsgFt11lrVn/nOyeB8R
21+7uIQ9ymr0CWZlziLLSMCSNS2CtRV4AHckPfCCLW0ZbYGtF80CFnKVfHTGWk4I48BKfJ+KjQfw
VAl3DQM7gLdnhmoVR5sP4VCUYf4yXQw6WDW7ZiQRgsxZVTaiP+AkWoWHYKyhu860j2pcL8EzOe8t
dNZS9WBDOfDMQNM5M9MBe7EUjN8SPGs7DnGEz6bz1jySowaQ4PxOUGUi1lzlZ/esQnu/xhu3a0GI
jPzhZzJP+Y6LnVVVs0hIaE7g5lsR5HKkcVeX9jpVOGVmdUJBiEYzDyE/cFGOeZsrQJBWDMC5Xgno
jn41IZue1XU1Z43yYB9jegDz5ecfGZqkJYWpqPwBY0pdnYKCsbEYtBTe0l7aKJmVFAp4qUxBacSl
o8wAeUAo8RmkcklQj/CAjXSAJ1wIC6blU40bZzZSdfjCV7z/EZsw/jVBmSvepelpf3mHdQUDBGRA
i4UFoywUodK7XXG0HFYMGYRcY9CkGV11In2fF5ZDf2TqvngyVo2FSvHZZIEwRKUf6P8WovyrDnJM
8jOBWcLQMBBQi2KubqSuEwusBLcmmDwkIRLtGhNn6m0RcXFpF2NLVK4/rGG15eiH6nH96mjqx5Vo
6WOFoaQxx47I4fc3POG9VNAWi6++B0zi7cfo9WEsid8D8rivso8fa5Hjyj62sD/EFiASPbOGeus3
nekC8ZV/OLAsddVgXWM/1mc/yMGk/dz3LVCCS7yrB/wTguMkOy94Zc5p6eIjiZfNAO5xC1iK+D+C
fESqPhkO3BJqkF5c2/ClF6pRmiqqJI65yuqlssdafXLCIHJ346de9a5UAFZ4/54O1xYeAZHbHwLy
rQomzgml669exGj3FNOl/ThUZNN9CmrxiPZCpW2lIbtOaCgJF1TnXLza4DhJfk9+jy6t1byGogDt
l95Zq2kjBZ+sCloK7kI6sr0N7q3kwAf0cCb3ldRas3pt/cEIYPtztOjT2CaDgnS5e1GYMZ1B6dRz
fs0DBwOYQTCWhXuesRQkAYyOK2MaT/brYt6qQT+7wChE38NtYitPDNwFvGGYqfScpsTxpDhmNadD
/W1YYRAjv/frTLtVxLC9z1cHxxAjnDz4nCxHXSogt1S+IDA9yUTwjS30Tnamcw3/NbKsf6qXoTs8
KWptDgaUhR3MXmYXfJ+Pnvy67XGwyhOwrIz9L40bwUwu9+MaIEWOOR/KsNGILXqk71O2PgiBTNmM
Y15HwHXR6WC2bj8b69W6GouaDhck/rN1IqZtu19IYDHeN+74glKNjYIxqiGZ/697gk4RfoEDc0Mf
kGVRBpM3o9COa/kir5sNqaO5iwrk174GaPoznkVZ0+SBkzBJsYIjcQ5CBX8mA3lctwWQOGz952ch
i7AiNFnL9/xVpAgW3QSBCUa6pBoBcyp3ME2y/JnxD6XD9/8wjWSO4ePR6Eh99tEgV+RFG53+Lp52
yWUixB1RVwGsA0vupBEtC70c7z8ZB39EdZb4e6NUfX8syXzzEjWDU5cVpop86aj+d8k2YQvpmATB
rOh5JDHi1Pk+a46fjucMIvMK/jaWX3253IB2CS0yld9aB1FHy461xQPtQ/4I7EAAobCs3jVyXzvs
nCbDP14rIDVeeE1gO105L+LdBeReY4d/W0ivIdgdA1qX73zYF38zJo84wABS7WLBQriYnNDBkluv
Ski5GJ2Lhb26emLLx+o2k64aOlyNPdAxfCdjq+SFu56jN2uzs7M5EuFQUuKdGBn+v2ZsVn7dL8fr
cuNy3FVR5EvFho4i+zsus4U9BPNwpIxzMXgagyLLws2jlG2PIcSnD+DE+amNi/wVDweWEyTKTPfO
lzx2BBYdygKgNatHFUeSlfTIviL5t4wZ8A/+tEv+3yLxLftUs+GB3xwjCvsfU2uCO7Is/HFBSH36
0d70CxMe0FLZggrhrHCDRLkbfOveMwaeWa+ihRKeFpuRuO6goGESbSxTxJQGXOF73FubJx3v49Ol
epGIHbXOmgBcAM3F28gPlK06u0yTpkh+i5xhKwLu22O1ntgXaa96YKqH49HJI3CVQnxouBbWCTnZ
Tsy9u9HIN9J2s6hzPmZx+fSRRhmD7lwEjKlejVAoPwnrRsg3XL5JfsG8neHfbQU4MRmsa1cO7g/e
1GlQzrg27UATpoZnzHKtewCUDlbFT3GKwkrqX8xoQfJ0jpsZ4OCaeen1hxa9RxhjFAA2EEwr7iCy
+X3LcQboBIqVI2R5v2pzxZ41D/Cpb3D4jQKhAJ5BZzwfHS22btZqlCAkB6NBLxY7Sx4leopHs/TZ
mWIrrydNt4QNP/WkpAs+Obm0N7fTbIjGRMdSclnglnpK+wMaCr3G25bLrMzwyKoyWQH5YUkyTRbE
SajLp911ceZqR4FPmlqCBWKXJwFG/tLKODB6mGj0+enUkvwyADMH159AYk9DK7hiiN4x7kghYTkS
KLhHx6QgwLdjZCjG8Ly/7cGk92zIqQk3qBfjZsR9HENnKvIFyRUi3BAESZueIvCy4GuwFu3EXaHC
A4IwYYDZ5uUK02S9rJf8O5iUde5TAxB2V9kUQi6S2YF8Ql1uK7ouP0uCm6MZsOPv8VQhhTveIwvz
3iCl1538sr2oSVSvuWfWYpNfGXmDFrNXjdRbIUqivyRjFSGEkYxvAv1D4k8YxyL8P34Ef98s64jv
spHGsdHj6GxiAhJeLU6BnACkcyG53Caoy01hBVOZ8wNX2XPRrk+KUlW3ZA915MAbwMg794VejtBU
uxR4VxCpOpxz0ghF8jiFyBOSwoukFSzimeQmbva3OG40uHUrtLpxLWhKy5yCfIHqZziSBD4k94OB
Yl1zhL7XtU98EoGvdydopGCDnUcHXA8aHOginaCxtFh8tEuxj5t+Deve2dnePZ8dZa1hhbtnaGn+
BB+QxiR+1qlB7RJkEXTm2jB2PaoHXqapF9ThKViZBG/pJC/aJavi1kaI/d4sTihfCLK/whNKhlbr
Bh2YqoqF70BJ3Gjd0zf4dHUbDPf2r5M8Xf4wtWQMeN8qY9wS7Xym9HRpa5NnIQJQ9+CDT/sm3Img
1Khgmey7S/NeiWv74O6RJZu6GtzRy0/fhc1+GRYkPtcKeMQ4nkCrJZvGLMhLyDtUHuY4Lj+zzV72
p2MGKFjfPW04aVej/fiGaiWfuSG6e/mvqPVKFfdyHaTxOIf7fvOHED5Izta8otUZW1yD9bEd0xMd
4ycdyy/g47TACUYos1lRow58HqxPhZLIH3lBp6phK8yQ0Vdc0/Vv+5uWRW81gkNshfRwUFaG5aYd
ajibGSGmOK5O9+NtkOawywCEAEdVxCxML6BeMFXcNTpXO562NajVyDQxEV10WjE8prCU666pRAtZ
yg9GsguuXMYq3pKnArgkqZZlOcg8fhC/d/dB/7jTVbe5Pdv29d0yXVfoO1e6l/PSx9ntJ2Q06STH
eRkicYp+j1fnZ0ATsvs22nDuST07jSEFjCPTPqi6I/GZrvGcNu6heIMUKP9vIZnjtW00mdhBezqu
33hxK+ZdJFv24LZAeIMHxWHJCoH+LgMn9r9VLppQ8v6P1k4ULeCOWfrp91dBzhqeCaPwjE3d/ohU
IA+QH6NkIZADkld9FJmy3PSlZVEomGoTnQkncyh1tVmLDeTLQbx08mpXBqaqQLyH9GWBuUjcvqXr
AiShHG3bhZ8hqFpsKy0UyW4UdMCn6ZXTC3KyTlG7x+w3/4pCxhaLpaMwnsgIKlLQaisTnFFsyjav
SP1PguB6a0w3BCAy3Z0uIsxOIg2pjmLxf62oA/IVJR4R1Bv0TbcxNgR56uRsTg1MssjYCNFAWQC6
gdoj6enJR3hE5xC/ueZpNRZhO9iaBxaZmUuuxC+U5z0sUMJ+ECTPa000owaHuXeuyzo9JPwg4+1M
KcVJ5Ix9s2Y4hhMFEyvFIKmo2K0sQaSPvl0iI4N8FXSaqj1mK0jQVaS78lARxqbkv15DbIjd8wDv
dps3k6DfcKGvZDp1LVni+JeTRg0Q7u1Va1+tB7zOl32GumGoaMxASKt35ECxkRjTklCqWi8mI0An
3xLHduEXDmTRapgwzzt7ubSNsiHiIKKkOw2+GLCwyIUXg2II87Pl4htNBRE3WsHdnd8nKDojbzXV
vYBQqOx8SjbNip9TEpBdbqhOWw4jy/XeLRjOzlpBk5z/mVCoXAir5BV0tIATcXPFWG7xwVGzeWig
bhv3KJcuBIcI7AE9QDu/Nr1+KoTb/I+wOzL2zKTpa+7KKBWVti9AJU3pNvYtXGiYVLYvNlOePgjF
tC92WlCxatbVosyxhLsKzQwlQPPrfvXa8cRqKU+LarNk2Tkzf1VNYs14ZZe66xzopuIAZHhZkgAa
NobLsSM8xw8HHMLoUMbTr3Nb9nEX0wkrAH3zuya+gh+SxOauG6SwWsE0bxEyt/JcF++5ovaskByY
lQssvN89F6t0FbtSuJhmj/P+q8Cs1bmieYd1U/VKHpDK/d9lAuX+eNgMzDKQM9SEdI/4tamTM8eA
3CL3SFWatK0kpXdOmTiYeTshoJ4+8oYOiQ2vKqgPpEYGzF618Gj+A7hvvQ8ZnRBgHqXFyJSUaj64
wGNCpJ7Elouog9wPL5wl85kugSyHBsNBUi0AxisSNx9lYcI1+4s0bbcU0SssWZVZ7EQd6y+HrhLj
SqN95XLTb2pRRv4bWh2kQAQlZ0jdHK3tiUkuNxOxmt4Kdo1J3CP1E1Dm89GVuBtn7DneUnGyZJoX
5m7QJV6bIgVfx0euGBtYKUCSArsvUCGsuN9qUFdruHWB6JwPE23Z4pCTfw3OAw54hQl8zlSdEONx
2f6Gewlk35K1BszWrxnDlhKgur4TNX56OYTF8M81GM2WOlLXIlxiQKRuW3lh2oO1MqGiJWJb18A3
SK97uoWEieLA29KJrnjrNnNPRxQtblGNnH7m0anM6C61RFZEQB60kydryOpsA1yMfX0ahtm4PRRJ
D3bnDHsfxd+I/BnHxA7w1w6lh2berQfFaxsfu4rxsWxzAHe6Npx6cw7ztnhIMJNS4xI4T0IF5l1/
tiSJvGlMztaZTR/uNlsEJti37RT4qzUPLLSbEyU3sxZY6g7vYya16z0O5k/BhhRbVH6Y7W/HW0Db
hoNNVpCpVd8jfmMQbNQ71gTC0LL1y565Ef2HU2P3B9g640ehpbkqob+l7p4FFujNXINYr1RKrfzs
Wj5jVzntmJD3p480LeDythwuIcBw1krpyLo6lc4zMTGkOfI7d+ZFqFpBhQOXWhr+8dT58NdJoLEi
v0T2VK9jYA27V9h4MjkYpud37oq7Aq+osPsOqFZHo0iy2XjjcVvaqyJv0l5NVFCGOf4PTZAMCTBE
BxAKbSzjkP6VKsiZtE/VIa0WTsNhJ8lXnFavPgfCn9TocGT4F3C4c7fum6MORLfdFJ/6hxxPHAOb
eNRvZcFULkANCEWVzvJvdqrJJt0atWEaXK6iMfBc5jT16LhiAEw40E7IhqDyJGX6i6p1a6Bf2JPt
3fFNWHAmmp4m/gqsGyg4AOS+BGAO7BwsphNknipz7H4SCWPopu995vvkrXg80FL9G1e75xuFZ0NF
F/itaLbUSaqu2hVBp+PmByuOezioNtdZ9penRvD2JGsbj7sI3hIgotRxYnxFimXBmgM9aVHWztNd
E/Or3DV1Oax/3/3gLcLF4upPeXGKQFTb5saEm7UclvV3akbUxQ5yd0rlx1tqJXYaLND9gJwoZ5E/
vbylmt7/0PZN/u8iDJxxxPtyhEoEyCGobKuoGK8OYM/zQ8PHJsDqurtjytBZENhoMq0N1ry52a5L
KgZWpjPop6zcF6kIuXRkYJCPfOkFWKy3G24LDKsO6aLw5gnDoTztomS/MORAjp73NVpzqmL3lFh5
pRgvvUt0dBBohlsO6D9XEvn9rCm5iq0J8Nxml3mUp2w/cszNyoqC14lnf2AeH8AJdHnIS5zBf68b
wpxWSgHKei1KcXx0eWKe28OzyOaOTzv7GLedyKv/syGygDLWlOHENfBhyKdEXvFwGqGMI2TCbW9n
VUSlZPbWjUwC5xs+TC6IHHitN5ipZcGvjcQM9DX9WTL1YA00t6NrKPfcOIUMWKM8PmMOh2yCUVoz
afbd9wmsoACzHUWzQTTQiIblE0FYM57khoC3At0cEffWADag9xtj0EwD/5xMW/zeG9YNUWkQ9Dyw
u0ge8MDoPjIeibKmJr9q8N/3ytmGd3La+2vscSzwnrO6XO+mYOQjT/Cw7AS6u09ij3ZgCzIfyIuv
I41ZUTXlQCrsLxMZGuDvnmZEsC5GwmKDM/EmcVSLwV5/QOHaYHr/3fGT5nARI09ZZJdbD2RCDWsH
mNZq1xjV7cdTkKQGbV/d5N/iT6az6qnciuOm+MBUVZsSiOUir9mLhIFAUR+W+inkne9V+bx6T6Yg
epLQrxpSr0geIKVDQgwFpKrcpUSCzxpF66Nf013q7AXwIcYMFFjW5wAU9yEfzpzdLxHyKOxnmrj1
Tc02yxf9m2LXJZLxeiQ/8bWm3wW5SL9s/LvqVhKc/e3Qn24FrP6xWhJegwpLuIvCwkBtmR24X2pG
DTBKqX0szEoe5ilBOnw3TN6z2g2ho2l07NhyXNL+ybzs52pco4iGb9prMlH0rl4Ux3edBK6MHoLF
RlOkOcmU+Az+5QghVbNKFOeT0uB6pobJ7oMy14RMTDbFtnBCcEUj+uIP7aFXH3hxHcsAQkignKy4
sb6mbDZWUdPP05NiTDDULT0Y8Dggpnh/GFR0IqxR+PRxYAW8wNfU9EPPaymsqc11lbuEbFDstoWT
4JHfn8Hd0Xdy4elwiE818J0xHQ2Vc8x5Tbfd5CMEr+UTMj/4wKcE//QczinFOhMt66VQzPA5gdEa
yrdx/dDwiIewWTZsYwpusEK0VOgB2MONJv2b61Vg1B88enJ3Xr6qqvoY/S3FOHBQ3YINYOq0zoVV
kZTb1gb7+5JJhUhu4jTg/pml1hLCaD7DebQ4lpucy5Mz0xVGqD40h9h5xJU4+QuFRFMiLNR6W6rb
S3NnHrddHmmJQWvzu8pa5sn8dlWhxXAy4kdnDfZTnawkfsbAbfKtNZFzPPSbdYwKkwcAphRR6lHx
H1kLoYte6IvMTSYeTVhgK6Uv8xXKC32/i0MQFFxiib1+wtJotrqIf2aYpnHYwvf6uGuIfx/XLmIf
zIlk2ZtLeXK71pAthU5IObKQMllv9Ikz5gQ+/pM4kzlCE1noIcg0nHoBhVjzR3zft/1XoXM8w4jN
w3zsvxWuqXfWJpR7zqUEI6tKSZPwLJnqS3mZk7YXdH7JX0IhjAvWRKN0C/Ty0DJbNGHGd0xKQhz+
z+LQgka1rrEMYKChuCxSjy951PfbUizC/R3KsfduPbwI0G83gxFX2SfbxSbYYl3JCqq+ta42D5dy
gth1T4gfSJGSt8+sOnKYIozsDuTAHP5ajvadpB975fKqdQbPhl2jT4OzDsOw/r0Zov1CfNp6cuuE
95Q/yQb1Bec9MuE3xYmUNZZdeQsdznQyf4ZDS6efrK3WTVV+NoJFcr0529sQa+nXBD7F/NIRRNFZ
I6AYpWfHvOLvmVJCw41/loUQL9FSwSCBS5Wh0w5vVfaBLxoVjk0H52SmH9edMzgYEi/lFIBjl50K
/lwHUFzcC2qOV2n+sdatd7u6exbbp9ufOQeZnLqJUCwg99+PcFa1oL5IRHJXvKz0uqFDWM7/+4Yz
MRwjoerDJp8pEB8jl75WI2QSm6LoAcCfzHtmOOTZ0Kh7foOT7X9tPyeHjkQXULeRPJLTK4PJLWXZ
tuYj5RXqHbmw0Cqfc1A0Dx3lv3EeE6JV3DOyAjY5rC/S2J6SXkVMDF/XQIia5wLaNJYYGMSjHs6M
6bjgyP4vzLueYk6LGEjYl8qT76zpzWZCryaTGXPYVbkTZhy6kmF5dLYu4PjikXak5XMsHy4KJhmQ
na6wWKI7WSiH7p8dmttMf5Dsm7YxJoLkv6+wfnt5f5y05g8Cyiy30Z4Bsapv+jxhOGN0z8hdD8Dp
CFWsWFE4DnBzZSc6GhxAtgthohBS/6MqdB9hQ1uMEAHzgyPRa0bs08+PWiRFy9SnFalEKMdFOURy
s9LeJu43x1cK+AgNalR+YL1AcWA1qCy64DkrpEba4m8aUekpDVbjuNZmpKoTH2fVwFENV6LwzzCd
FtDqDuG0aRkQHQWZOAC8EnhdT4tca5RRn7kUJXBh04SIy6W5GxoaknN5/Nx67E66Jw6N8Zl6+QDg
sUNtrfkh3UZgQOG15wRIvssx1coNPUKpJlZPPsJQN+rVQTeM3TgjbYCieFTA4LRouQEVeMm/lZID
iadGeQq2v5mEV/OsBmwB+CywgWIKnePwi3Z+MNZb5icE8u2jc1nPWfoLGBXOy7eKiNPXIlgfLlUc
sx7MeIf1ZINZoN/4wm/PGcMsNCupLMSNtooqjAgwfEQMBvD2aUc43CCLPSFuhE1cl0tYcSNScQrX
CyNcSe6efxu+m1NUA/EqbdHzFGbg7oevAu5gBe11iDsQ0NqaU1BKZvnou0wf4w0nGd4HuwR8Gdd/
pWoiYKsYTydEeQlNFwqJk6BDT6W0Gaqoq03kMc46m3RuD1xaMJPPE5QrUI2Glu2cF5H7X3BRH0nl
HAHN2VL0+tlQV1cjBlXiArkx3564H7Qte9XIh6XF+PvZzTH0O85QiX1IWZP34u5OAaiEnTMxglYT
c2mMHiDg7Ahocqb7+YQc/o+FLUTkhxB0CgwP/N1nqne2I/IOwQRk6C1bJqK/lZhV6NzzYU+neF5a
+FYtOPWUw2z6RsD58OXAroOaOzaW1Ipwxi1Kc1hKKjmuKkedBiCEoR52ywxMVmZGO2vsItWHTGIO
kRSRLmKsnDIriCLKZKzR8x6+5AfcyW7VLpocptqUI7pWY9DJZ0ApcHZCtAZ/lvAqfT/Z2I96BSjR
jFV+eMJCGKyk35Z9z5MLf4hFyIyLu8rpvNHjebr74JWMc/8t/6rTA/OcH3KqBbA+lER8EY1GE0Uj
/Cs62ObwEnCRXwDQd7UfBn0MfUG4oYYOGa6MH025UE2Ghbfjkc521PuTsN5PLNN6YE5U8sE/Y2U1
fcqAywEohZMB+QEF/30FXR4itz59MnJKC0chMJzDi12HWN2/rgEe/lFghWvRdfCePPZYcJWDOFHG
KM2cZDo/H/WHPIdwVmnSMvGJWNo7gVg26TmSXINAzWSpl6jElo+Wl8e4GXQAseXFgLwCEUHPPoCg
Y8khJVC6lMt0Wm0HfNVu9jE3LpMo/I6HUHagX3CE17/CoaU5aAXwj+15fV1At+Dgoi0WNzX5ifAR
esnuA2kqAdll0Emclkez9s2ySo3NCPSJ1FD/obC045wHXZRKOiA7rW/fjO30oXDLyYvxvj3o4ZBL
7zdhBKnYt+GIpdza1FHKLJW+dHm/jjiix6OxXSZCMcbiqbrBawDnDAxXwIZk++vWncCT2dwE8wlg
oYIVI2ZGyPBowz4WZ1H0CnRlpxy5s7WQnrWBAvYRf71Aa3ppFsb2EiCnRZHIZvYfVPSknHbCNzSd
Vj0ZPa9ptzHDgyLcIp9b85WmIk3izItsqgImclMYIB4byxN4DxJ9uPuSNrNCKKlGwgVm4CapaL1x
/+7FUGkpEXWf8DxnQJFjCKiKsjXYC3if8Zb0kZNj0M1y3gOfbzmvszj5PZCSmedVLvrJH1Qn0j42
zTqnnthWukESS2HafC9nCkhNAdQgYF5OwSDBXf70TljC9+VBhxqwbbozr+lm6K7lGtfWcotd0+aA
VE7wPKNww5qJC5SGA45Ns65hMCAbUnGAkmGVjNH9rz1PQ5KSYuJFo1YvX9nA02vYpHpHBNU9MfaK
UiCfEubMul8Mjnr9npTHp59w4jvyHRQsPGCeo1B1MI+cNq2O2QX/5MRSzu+esoCqrHL/Eivvb87j
HeG2SKwkXHgBKzArRO1EBbskA32s3cHEVjchd7RBB72Kyy1Hcb+XAamy8VuPxOA3nGYA/vlXYOkn
y522uo0DLG+B2oyBmttRfgQOUtZSELCgptQqVS09HV4X+falY6/+yTdCApVXEOfpm1iiqqTM/yLP
L6MPqR7eHGQaBmzrOCn3fCI8T6fsAwy2aS2gUTSN9Uz+pqlsnAI+Bxv6vDs/vEqajdaYi13AxreF
Cy9I2wCsensOEimhtkwR2OBGupT/Xh1KZG+3frCjvPFkewaKE4ghS1C3w5+xE3gL3LQv+/ctMMPI
9XZE5F3L3YfYRb33ys+CGs1Abf+YqNdTUny/yq3ZuUcFDW6habi5dCzZNWwFibg60I+O/Es+i0QY
q5030tcKzAkoW0u0WbEWHczJZDJEgxq3VYtacB5t+JHTWz0kIzNK1nRhzH9iRzMRkVaxeym5yocV
0VrMWndCUIWHauuI/uGSiXgP/gZepBkiKc62SJsEQwh/EsudzYsda2dcWgjkUMvUc5mLOP/F7rjC
vXAL7fgJ1ugXG5pUnG0L77YsnSLbYbqhRK77GfxA1CTrn1DwKB/JUrVB+IZM8yqYh9RetM5VyBko
3WADNxorcAE2pkqUH8I4geQVYWTRt4wUBIHGVrKXQ4qD08c3ncD/y8c7zZJlK1QKPuKqfVPrFQMn
TmYfhLVXiIlkihlNujRtFMV/n0fWjqLU+bsC8HfmB2Plq7gCrIjBMuiyxNtZBwC7tFs2Ca+c+wEB
+bPcDskJAzM8pHEv2JamB3b/73wPcD3udPLH04bt0yJ/AmAoq+6IpNxQ2H/lBAbJe2WYSVQ6N3cZ
RkQwSwrIdT6pvxqmu9OHte9JkpmZSndWalisKx8frkl1ga2adx3ZRVE6YNteosop8euCTn5j92nm
0WDn06pqra3mxHzgATncOyoba8lNRqSA2tOD/0UBZ9jDNqAiIQ6AYsioSev5lOXqusdS5AsghbrF
1FwV4mkaY4eEMlq6fh16KXUNZQrhf1fBtCXB4kB1YmY0VXrLe3WgZhFj/HqKb+QTHFP3ayYiVn05
5lOWQgdoT5G6lfIxrugsWwL5MuIe1Yqx+deCkLM7GSciGz6gGIjjFj6jcP90zwAUy/ATx1UVoSes
Tw5VhBYPwBozuAd4Zv5+8ky89Ab4gye4TRwYoQyEzDkMsRRWOiUxoAo+bqyzyiRGTLkN/I+SwMqF
4YwUdMLt/0eM1xJzygFlm2Jlda3tA9VjnyiyktEBKgdwy8PumE17oqlqoAKBP25WLyzJ5qkeX0f/
q12/oLogjk3idiuuYPst1V+h9bH/BtdQsA04mDRRggHz40Id0wIOZdHkuVjxQGAiA9/xeCMgXcjT
phYu9H+NnSXXC+xnwFPArGf3h8A6oXIVeTujx+KFfnN+ZssaWrqyc+x2qv4LNZFCbcsgGFYM6QCt
NX0Sax91NtJ86UOxZ6nqeXdqkErIbGO+E0gobHRlloG6a9IggslNDnatf2CVhF+DlYZuktkUtnfv
ato8WEBysAEZfS6m/Tayc5JHyF2Uw/pO/rh6GLdOcKSyvA7R08Z+VHCnEfAZwOWJMVcQ/7hE4xyQ
I9NAwhf/sZeze0dhhUJyDeWuJDtHQzgSkx5pJiuRceg7naal3DUv3Zs/3IPU1as5aQVrU2AJBNTu
+6r1FKkvs0oNS90Xg6XcqxJ5baHt+yksHdoiqqIfofmOkd5QH4NUORLxkM7xmlrXpB3wDMfD3FOU
A7Z4//45QXEZKFu0yq+zcLlRQrCDCTrxpPgul+B48mS6WFSy1B5vZ0VhKNye9pHPnPHd1PI8UaOz
JI7BcTEuCSh3ewVzsAos2ccJzxH17czB+26o8+TY6QM5oMLNauEITASvGw/hl8K/7uQYQCvS6Qw0
pU5T0q5zXBsivAe33kqW0j35YShnUVEXNL2HB1V6x0HqJ0BBEQcpLIHywOQLzJAt9PQJETzIIqB1
JUPm57fKfHo+D4cx9g4Dtmh+kNSbfF/Q876Qri2iGcGF9qNqZvs2y4K+mRUA3Gt/YSMJVNGqwDJL
/ACESdwouTf5ZbLpFawcgZHy9NTX2ExreDRiQ9JScPeWsIncNnLuBMc531HPSIh47+R5HPskeAxn
pPIUZc15JCKZyatTjvwAC48ipt1jWuNrg5uNtwmJKRnjv3WGhbW9NaCiH+RJunqK00glRYTEZ6dE
hZH+UPzbfPhdd07HzQvQjeB6q6LxVqZ/9RutCCppFw6/Eq+NYOu4LxYuRtvnIjGOssKRBQaXlgoZ
mjiVUpBDdwCeb+URbjDG3rWcHRbyhh0abtWdzjvnIh0OgZcyZAxMbMVIXUpHb77VR5gXYXHbRZ1m
JKQtp7Ztj4SYH3FOjN1X4KaAtSQJ8IA/5HfQvrR3ZbtwBDoIP0L4YujZFCsJi6lKmnltpU2ond8d
eJ72oG0C6GJ6iGD8aMDPBKFxcJNQoJN1EVFp9xeUtHSFOWQtXDONXqesiPcDBNr37Rw+Glkj0uZL
Rpo23jhDsj7/lt0gnGburFFhgN69vx3n87iB0MtgPH4QO22g9hrdTehEmVls5uESoGG9brsEMWIl
kXOTgvhX7mBzl/CI4SLO0XeyfFcECmH0mHW5Jo8lKS9pcUBad3lHfomWJAf4EYfy8sx/eHbap2t/
3MQQr+T5eg/BJxrpbsEEGsUkuu1V17GWI4YG4ABpOIbaPakSlwu3UOr6qYEtCzYdLuNSGpg1Nfvj
TDMxgt81bHtL+gfhC/e5i6qIVByuDdBg5Ced5rYPPmZOFYAnEpxmowge7oKkt6hpljgZ7EQaIOVe
XoYEShSM2EizgFCYVH7fvgZ4nzA5ek6YglPr9b0Xia0xbV/+f+svT8TgxBE8bry9/x0hmetqbBxd
OcFqAUnNBOq4euKzkiRTIKxg/vp7WigeGA9mJEAPDtee0YqPnosxqIEf2BRJJuav4GzJunFU3cNT
5E65Llki3aPR9RAWgxhB6Y+VE3T8j87giPYMJTiAxp2Pgy6Ccchvi73UOWn516NtN36DzMP9MUsA
XF3VpwKulGiJbMLbY/M06PLGSPJ740YVjY/8Nxqkl5JygxTILHuZ+dOR+UMNys94Wxm7Kb1OvNOg
zrfV5qus6Q+hih1CM2RYhjevWF7DKRbVuBzztUwm30Taw5rxtEMIsYf2cqbwzMp/OGW7iTsbeL5Y
PywXQNxjhuBOXYpKGRsF5UlqA1qhlo8rUfCk0kIeiVZbdp+fNMxYhDBkS6MLBycuqKWz6sC4JVNd
lF7Z0ID3/ke0R2buVzALE+N3gwObmYZU4AOJZgVkthT9qeIuy1lYGB8gawtgmMOp+RHGCT+SKoG+
3DhfGfPnsIHWF8UEiPa4bo18MwoiCGjgTZbtl5ULRpa9yTKW4AhTIMZ+5BX4YCn24noBOQtQcBvC
+fkYSd2LTAxOx6jERvyDxBQ8biz5BW1JaQeClN+XHxxBSXYL5cSm/tPFsmJbvLp8Khijd5YeWt5J
S49yeJdUPEFLuAFoVM+wZGG2zh7QW+c0D6t9dCpUpJRniqIvhWZ2s8lfkCwLffJeNTamLYzMu7sX
tT5mFO4XFbYkigOWt+ZiPn0x/Uma0r2BsQYUocqcco921R1zEkjjVLsbv/FTACxXtU8MNUTaUfg8
B8c+m7zmcromTx/LbHj8pckryIan2whl80hHfafMhMKG+THpOZQeVBLeViapqRrSDuKpyJN2xj6K
ZddV6VzMk9GPvQ/YpnOeCNxb6Rw0cEonLE3HYnyrj4NVYPr76pCtxtLY2BdIGo9TTjBeHW0Nphnf
m2yP1qMbaZFwjBeioxKJzQJy7thSuDy1OYDbR98COHXwpe+YwEAtskkQeEUW/fDbnqV/ip57qoiS
rJOwvIAe/exWY574wMEWYufVG3ujoI6PZ0yVrIwMh9QLmCSajaUxM8P6V30JKyndakJt2tMPncRW
IUxepGiJZEQ4p+6N4hUdHmKnCPNIqeFXzJkfyx0dsrH1J0NXg8swxOu0KeIdYijwbA630m9XSXE3
E9mP22AKnj1sAYJnVU7XKf2kQAMvce6CLNw/jpOcDFBcrrl3+t7P0fV9nCvdG4UBy/BVPhIIXmWp
pDEKDxxWEsvUkUeN+BTBbTqyuMRJhQqK6nrb4mR2KBdXcX96RzFDFrAsEnSolp40a04rxUscPyBq
g3xmCcRnkVYAYv36LZu262gTIxtwA2kPA3PFf+3jUBQgHcQackbjnjxsUD24FiBIj1zN6/lhTkFc
WQms02ShCFQ1L+SaYcajJGDAzkLuKWM12EUC43Hei0EqeJrV14mXFYRqoOPriEsa0U4atIXf0NlK
hmkWM9reroeGQhRoK0WW1PuE7b+h1AP9EM1WXGCWOvrMrNj2JWsGfeqOk0NAWYZTDqfVkTNcuTu8
OFy8tYNae7stD5Dzn9Oj6FMll5JrDcbvb2V3XInAU9rGIO9zM4JGZ/UhhNskBtrHCUrVFvtqqkoF
cAOk1aKZL0x0WyLYMlE9mCYk83+4PynT6gkE7tWo/qWGeKdRUG4JaGg955BFoBh5KUwOmv4d0ONk
2EpEqQAr442OwLPXxcRG16RcApEmVv4EHSoeEc1v1mG4KGDkmU2X2d9kLFit5VO8g91v5I9qiG5j
sZItsS7TEwdn8rPmrfbeO5ngqf3S0tSmlOz8O6m2uKwNZFamDrfO++aWyrWgMcNc3JvXskGVrz62
dxPIcfH53ftII7jZZz+70MKRl4hCXZ9K2GGxFAeNScaLMSsRJ2dyhsckFunuspXU7DaPZbbbVNjU
pS3IJgmEoInLcBUB4Fm6Z2eBIpOQ9HmPjLb24nHZIi9YnAsDmhXaHahyXk8NgQ5cPGvmpbTP7h6e
sSxvczlpdXBSQuCBW75/hVrUu8U86Y57+QbhQt9jnr06FW40sqyLkh5UG/6acTSutriY+lKnw/wn
4JQPRFD9l+O/wuA6Vo/aZ8yk/QN/uETEd8GOQz5eBHDfsuMBjt0RyaQRp8xfR3+1jKRcrcEWc5l7
VRSIRSxJZ9QFHmSN3k6kNPdtZMZ94l3R3vQvUSaDIC4SymY4T4qB57vB3f4Nxihr2cf+lgja/xnr
K1o5OEWNLXgTKDy1d23M8+P0Sp9kVdnWWl/+XdZ14TKkAISOkAXXgNteVeGDykZjdwIXlz16k/X/
A9XPlqbMveuMhmHjWW4m/KL/iM231jThPB+MVmaeoncJ/6iCaU6lAto9C/kgTTYVxK27bYyiDCmt
5n1cId+pTWk818OQ1t8dOGAsG6v5F4Jj/b0bBD+/kmT7C/uHRNSJSj77PKoFQQLuUIIgUyU4jUu2
XYEkpJelatnq48RzqZOJ0b9wR1EEpf/FByuk1N1P1RhU8mLaXakFBsgtxxX3rMfiJmct6xLRjpMq
/NXeqrwc/3cPGaOb8VIWt63fKl3Cllh6P/BU9XTDkZD2JBnaZPsfzDjHHb9Zq8LxW3m4pXljZg2R
flq/fjr7g7+daNt+C5Z1PTBFW2KVD/41lhC542tRIaOp5Ml0gb9yAsd7osMlU4B107CRw9qyj3xg
meBWNAvwhRkhHa5bm6neBo1sofYKCqM7gQ2qX0Rh+eq9L7wR0WjFckJt93l1IyUow1Xr1nnfr+Bq
rfQDdhFnZCz9kKXbwymCsS3L4ZNoxwgf5SsHl5bh8Dzukr437llk2YpX17UISepl1j3lCYjkTRI+
oAtsVIdlQKn/sIbvkYICUVbBWQaQWoSJ0Ax7niu8KwyVF0m/gyywBwsYXIL6U97zLgiTDNqkifxr
KVvnd6LOA2tbod/kphg10EPd1wp9mOckUP6k4RN1ng2v4LvJ1MXC8znddBrcXWUQ0VJmWozIRPDs
oKn3Ny3lNQ1rftsDKgxL2B4Uz1JFa3a9BGN1WybjifULSd/zsXX2n7H3CidfINZUcOoA3c4XD2Rv
RbCv4qWPe3XvhJW1F95TVxSs4JjA87n4h4acwMbM/0Ep93o8OCZT3cE62Qj1TlxDPSgZN7HU9c4X
pEgS7lqDv9Zui7UzH22d3WbawlD5oOgs61ZFyO63cZEoySI0JqDfIvtwVA6R0X/sKE7j19luvxo7
XMKsydf+piwjQ5Uo7MkCp19BFgA2Qz5nuUIwUn2pN4CtWVDyu2vlWOtud4t2VkHTT1YKPuH1NQtv
JHxAqlHz9v0WDl13hy5asGWc+7OnJgz15n3Y/++5Ttu58aCYaAe1io1DJ/l8sXBJSLzOx2rTbsa8
IP4C3tIUQO3alTj9haynn4L0aKA1z8EXa+YnX/+XZneST7GAMK1JkPEnDD8H4Vk/7jwS+ZeR8/JJ
BMfNfF+4a+qZRD0KG2ef2NtpJ7Mqunt3Z0kZiCllyzG/VR9nM7T1dy/tqVhi+9wxAYvTbU+yEjG3
/srMWSgZj7PXTtKI9yhnPvm+Lwc2tUIFC8y1i5OxACZZnq0wAV2qt3fsfBmTjvE2mhBjVUWBhC0o
Qnfw6LTiaehp/aQGrN4Wg6eJYbHrce40eXvJHkO+j17TfWt4iS0x+JTO5VEG3PnT1FPm9yEqwZPQ
kOGfrPCLy5C2dGBZ1q20gK0vLr1cEjOo7c8kyG5RRjMSyk9gGCUuYWvMEghMQ8zZJVVe6ic2Slrp
OxSF86QfvunlLGvSMOyggFVOKG+/NsOHjKy8QHnmWqITk9gLn8vP5a38LjZqtjCJClQqXHW6m6JU
UBZUnrJ0o3VuR+pCS/1bKrHxuIz6x/L6kQxkCMhWDe2CmOWppZojfyrRx2Egu3X3Ivd8cxyTd8Pr
vHv9KNS3Y/1mj60h2ND8xdM7NBtbBrdTCaGiRA2hy7zyhRmDlFr7e1CxRB8MGq1Sqvcb3UYYsJUb
M/1MQFPTRQ6Y6mLjTZxSgtjyXrYt0bEZcVJBEWpBmEDjAWwaT2ZV1jH6DNpQhxFoCmpBYaPO/HHA
Jv41pgbFt8crEAKTif5KbVx/aDyiSdJXnKfJQRKuaQ04nIqlqXGY8hnT48hMpe0xtBmvblCKMcDm
Vt+AwdT7s5Zv7mCKgGoi4c/UKjavw3biT3iPrQejnfKtNgLcMe3sQIBM3rMPrnfkHAl1Yt28AdF2
FXoF0aO7DuVIOyFhbc3VkvxUoYPy3eJtHnSCYe9RYeGuxeZWDpXsE4D+0JW9uhIcpxifPlsJO/CT
6aH275PmNsR8Q7cOoDn9ZO4Fu5w975iXnT0QTfV1BkVJnvFVCdl5RnGcnZIEHkVuxBuqj7bwxb1C
RBnFdVvZX4rGqPAYFJv0XxOWUdgkpjjGYh+qBJE7Kwz13/dglNXY6IKG2P3eJy1Vd0EujleYwJCv
PSOHa2OjQse4KDwdyjvSGlJQ6whuxz6Sw95Q6cseX3Z9ftyLWlUfcm7KlNMuMxgDINtQ7FTgQkVW
mY/YCn8+VgHVQaFrOtkEbDO7JCTp/laRPH28waVObFEauwd6UsyhfGjm6oS6bYZvjsU1wGbU9h4X
TuD773llDkObbMS58hZ5m3+4ELU1QiQ7cYUq7LDh9UY64syfPj+28RcNfBrf0b0woElueJLyFVuz
ShCy5GMjzBVSkVvxu4FG8B5uRNh9VykfiqtQCJgXnopW8lkJE5rB8buIaBYYSysRJGaXniHaNEf3
A9Jppm3KhaywNbqpAauim5ijapULVgouA7luOOOzqEhjGj7p2EQQOsv29JSayp4xlrDveq8Nseez
0euBIAp2hG9itgoSSqChvK1kBgFw/LXWATgX/9SJIHa6oX+ea3TQ6Y1+CtHEuV51u/TlV0O1zPa0
NqHQRz5XlI7RQmKL8xsFc4+WaY11h7TcAwAFO1WAUF4XZvHc+tRD3VGKrukbKJhtNPz8XEaF41jc
sMnVpippALC0lsfLdT3vIYKjhQTqLnqWYe/NLdJxRq57pGvlzjFUB2p6VoK7ojTdlq9lb5eKThjA
WuUigSMkzFoLuCULec67R3T6SGeItGM5hwHDQzBUMZ6zg0hNb6YZiAnrfopwJ72yi5BvuXOm01pm
keNxikU+zLcetwWyN1toGofQBzFy2UGLvTj1gQLfcSIFzuEFVeUJvbe6gw3FOcuygou5r4CI+0fC
7fP5cOkzgDZOVNeqLWJYC483HOHKc84E7TOPbZUtOw2EgAAiYZKlbZXNNMtfM4Goto/cLSJkQpEw
R/i/udZTDImn0xxjayk6xBsCKeQXhYFfX98sYtlTZHvVaKBCVpDKSd60+90dMGtLwidlehYLPW4a
LXzyguAL8QCa5zulKDliQ52AxjeDd0tbnwGEI19U0R+GWu1KZtnYPTMbX89Lp2RWqEaKMQWe/cHF
JXZvhWKPDcsmRzHpdt32AIFzxQeEYn7QXwQ/I9NAfsUN4sk+Mb+MtL7gmHn/6R3KdMtC8IGUa/My
jzYzanGUg2MSbUh9GqYkc6aWYL/M+dTkv82poY16yjShkXtfzdmMsoq5yzpU9A6m5WMJ76e7FQRm
lF+pGNvCYMx2dHA31objgMmygBJGm7quUGxIuC8GR5RswldOJj54YFClSmJTNPCI96hUrfc7ii34
gWa2EFti6w+tAagxqN2eL/1CRPNZP54TpRK2uoSJbLtcWbzqAMr4L8IIbowxpXDhjVAfVOxefSXg
mG5tfTxkH4N7ZnWUN7nYL+mcAJyrfkrZXpuMBs2HqzllKu4iuvhO3G3ybjXxBB8FIvVrmhcqKJXD
fo/S5F03T1TnHvD8mB45OTIaVMEcQV2HHGnkA91iF7NkUw24kgo4XoDrju45Sn3sy1cUkeqt4gw0
Akh6EHTkHsdLmBseKdX6qqACpR5eAiVVnSkuKuXS9q8pY3xOZKzRuAY9ZLWH+3AaFJkPnwf1YcFp
LZFWiZ8Ii9CgIqzJep07X8veNOVah1vo0EM+7OqAc9aLE2O22LyyPYACu5mmkJdSmEm8PoQXSDCH
u+dQJYJqpp9SothmeCNjIVrr3usVMyzbnkFmpllK5ReY41to+e5IDoStE8cb6RZIDBNg9d2Eekwl
GnFGvJ6QsZia3tUiYiIAh1jF+vexWg60ETdDDSFhZSrE78zq3roOWNCaxCVkTJTJgGHhNbkgTiXV
RsmPq1AlFJDjFb1Rox9dHGWL8BIqGLMjoLbBri2DOzEAAscydAyW4Q8zvBck8BHWa5IuEiDIX96c
pssd5b29QL7051e1rSv7YLI44I544w+X1vzSlR1e40kC57SFda8VEGcn6ZJasOiZvLpTYQ+l6vcd
/TVYg4aupAA1kvN4u+ZqkZfM2HZcZnzoeWDjCipSscytVNIiSUTCJYvtz2eA6gmsm/9QOSMphRyT
p1YdwzY8GHbRHDHNcId56HpIDS6kq3rvVtYI2Ql7VHsDewcTKxHePXLmb+gwY8CXlcMevrH0QVtF
Is9oP81ybAqoFbYCkE3MiUCSK4seSwpJkLzVqr9mKjCqT7YI8oPSX6XM5OjlyEZLpJtJha6g9+Og
Sdfi8N51bkn9lLmuwan52RSePU8WUVHZiFhyDkSjMhjugntrtJddGWgCiU29N3uG1znNNSHWbIQj
fQkpEUpUSCNoHGYpo+MYUjYdo/a4osvMn3pb2+QGuJ/cj/m6spP26tU3/LiNcQiFbyf2U9FW8peZ
FI8yti6c8x+UmncTjxQdeGr8DeqiUHb8PYsy9BEVKsMyzwCIjonBiCQiBotaBXTDCOY1cwwtZD7R
hjUQaT9OTUaw3hi7n/t2Ly+ZZennqm9FaBHGt8VDV+xxMZQlwVIOEJbBBnZEZceJMb9t19eevBEj
moJBkfCCXiJNgdwjLdQkS4H0kR3xlqgIsf6Q99l/unaQRVhBwnacEB/kCXJgVC9MjVIBFRUa64p2
h7eUxspdXxq+cYCFViZQRuBcsPXWkuNxGEF36GMUfbnUOOR/d1h3x0Nmb0EIcN4k37wsCHEdlpqo
96U7zF7QPNW8gMZ3oz6YHc63fs2Ow3Sunw8HqY4ZQeBRARq8oEFjKI+SqTZXp1wyPHBtiUF3TPPY
YR6zpvo8IpKx/KE+p3CWc0wxed++kKa2R1MecJQgIcaPv/6zrgXK58V0UKCxLPU1F4tPVYuHM9y4
E5L4phwpOvLD8nkzZY7QxBDSFTBEqe6WNlf+8gaTNuNjphEBbo2Py82hUUjGWnIf0XqamvmOK7bL
54aIu+rJEksZYJhl9Grg2X59qO4aQj4vIvwKdipOrRjLPJgbEi4dYD8hJnMx/s70+Vu/zIItwOLU
BYxIMLw/S3/+DyHSMVQlnuqlqc/pDaQD/EGR6ERXQaFAMqD5QYGT7yUiBKIn7xV9GaarLBocexmA
f2rOXyZLZSX4xCHYqVeUpHhLAx3sxIs9z+4Sd/Q9rjHLrUmhuU7McZ6/fVPWQC5HZVf+6vteR2hM
DrV0cyBSkwGKM8FQtd0HfM/3upwZh0J74n6Fxt7wdeYTiISzHJ5QgDVAzimsM2AMSKnMQ+xWb97a
CjDxUDJZnikJ7iCzEFdEMD2tV4m1izV6QUX1jZpwUgq9m/eEr4kPV+6Zj8wISM9x4xvTBqASBINK
AOKbfbU9W4UtDKTQ0v3zEiz28+gpVK6m2CIhW2eAusfiCK2zl+/u0UH9EuW9UAhV70qcsBfmJKOa
/iu7U/IR6WJF/fQfGAFGLQ2nUvg5liMywuQuapqw8orVUnzl5TBOJLfxap13QdOaKwItbsV3nTWF
yMwxwStLAAcqw43gnzt+nN9+oPXrHezQuVtWKYufVjn+3JZ1HhmEhJwCbzuNlRTriuaEhg0o4ozi
VyoLYlWqoqDySdLfq11CE3e38PDnTo7VzLJ4MbJYVGmoOtGx+/tVdIAfjGhCOlLeWFlUyeKcFfGB
oYkYZyLJX3oWyZmTKXX8xOs3xBbDMH+GpnRDJcODmTrrsuDM20Bq7m0fpxW35Na7CbLm7naRNFz2
Z+aFcg6NlUBo164fTrAwcw8PhJTfUB7+UjZkbtL0dNbqbdQmgrSGp/XWvhSJlsRjtfTvVpa+GQTb
/iX3pVEP32FZjw2Yu+ClI9p3lPcftoXGPSOGxhqQLcGY+S50ZUN109WVS35YMEBiRP977NEV9zXf
6VM8qSW/TKn/7XZhaO899QsG0psOJGDEExQNeOqdu9O9kAkQjJJGt27FZj9OG7rs4cpaFa1iAoYV
2ymfY/KYKxhrzFlAyK7DVSMWhFI4ApNErjsRBT2+gAYGfQEmE+896lR/WrganbvtDh1SEwpMw8V1
tvXHfF9F5UKM5Ut+Ah8llIXnA+kLaQUnQCNKuC8UgmriewNRn5erbiyFYsEEJCBCB4R6PV/wjWiK
2sJR89D5alIV7Jmo6KzQzVj/e2RYt3QNX2+UxIKghBYNVMxPAU68Kzp4NVAImdDG5uUg4bLTsdU4
Efd1dOU7rS4OjGqJqyBlx1qabDssupoh52sTWDcgNO4SJwGiWBp2IDZeJ5PxN0W5KyV1cTraPIPn
542Q/vW1XD5UdfoMjsOtZTorNhJVDT1l8pByUL2cHhdwSbSvMaGnVJg738ie2nJThMurIOrpKPe7
QiUGZto6g8ZB7RnIBu8jrYPkispUWIrmi+m2GYZ5scSGDFX5RJ7Ur1NbVe6pcjopPyi4hRDi2FuP
EFN4RW05uDP+24GuJTXGfLNpzAdKT5WXxMHopke37vzDb3cE8bocQmbRXagEg3ZIGEmRV4CefP2B
XCrb/6tJSWwIvZYUeukt6Iyci3Z1+zVPIAem2yI8fgRzF7NvZqmwwPSWcS+glwhdz/WfP23bhGCT
lSGCgpw7AQ4hPIDjut7t33NtOCKXYb8/SU9lDSabUcZttZpy7Phk+57zakkJZp9zoUWeY7GQg6Fz
Hmn4ayTE/mM6A/JzrGXkeI916TvSEHzhcco3pX2fUhJ1inwZ/KDdbHBUvY5ryAxCTnPIM3gQ+y2h
vg+hCRvEJh3El4bMdZVy45fPj/bfnrW/T3YvnRIn41KS98R7eLW6XO8AOrXgEnqxtvpWDuh7mvWu
kzP3vqsSo2oz9xxF32Y0wC052zNDLjzq0p5ampzJvauDM811n3WZDd4jrmgo4ftrXsRFfNZJypZQ
z+VYBJj8ofticILhRbJEeZF8fXzgxWMuxoa5lyT3I7PV1b0qaYbKINFHpZatWPR7SYt2OQhOU07s
ncIt8G9Sj+2oFPhMgV3r53mGZplElkcrGnQBXw2tGpR9oV6kSASVYdLafsJ7tuKnjFH8FXH07Qd9
JDuPPJOAYlll11n3TAtx73LM1JIMTeHNIsgu0mxhvR2gQRrCqVOWB+Xa8goJWtC4SAERsrdugigD
2TA6cx7/pHO3h6bnRvd/U9+CP6vAExs61pjjMDfygkiylHKodYRokjH5lXyjn/vW49/b+3jV4ez3
SUHCZD28vZCKsP9NT2Z+OvckcnEzVYqAtsnkgMDj03wMOnGCzggjSIdFGQ1hmqdeHg0+SV9Tjwjy
2TBbT/kKEMIqPDiupsbX6gTOiJ6ciQKhwwpsZ1OAbjWxbxfQeQAKcsaEtQn8FjIoscvFTqo67tKl
jXfEH0jzqeeXNjqgg3sloRtoCttY5XEZCgoIyUQSoS22tgkFx7Jgu6AxMPIunQiBvjjv35xgKfXl
UlI3Md/M2Uq9Q+jllNysc9YJe9j5n8JOu+N+Zn+qiV9yLTLUExkKni9tWrE1RbuQ/EqjuXdev+jH
an71Kobx3aFbynORUdKuEe25JLZUv2IKi3+YMiCsu6LM2t74GXzdv41Bn8uYXdKzmyalC8ImI3p9
4+hVcWBLjCaXkb6P04EskBBSMlYugg7XWKmCL5gaIGcmMS6puo2k365la9rfCjqr6QAYOj+sGy9y
VO5C4HPgwZ4MnSgO9M7HjH+aUJPSa8oW1yMtF+RVneJ/2kBo+tzr75Vglf0gq4i9l0M5/KsValI/
jnnL42tNdYXkL09y1JBW3pjSKdCwPAvcw5cjBO5dFBPc3X6VA2vf2IuSmwqvwjiV4E70DkLDrqLN
CCXnUUTKW0jIaapuwC3pW1shyr9heEvLOilUwM5HtJckPsNJQvFagMqz5d3jdKITKiFi/TVyMEp7
4mMxGv7uX7+68r74ZoeeDRikztivrcx6rNNb9pdPEdtv0Dxzjhxq9vsunbS9elC7WwY7zokgG7xV
ENFP0wtbwX6CwhQ8JT6+Ri9mGYfc/H96Nj6jLGfEOPnAYbE/SCLUHRIQ97Hubgjwphr9RS6ppSgI
kkYmukLUjq4/4WaEREXlKGfhrHYBMLIC6zyyMz2WSQ4Szt4l6TYitUCHPATQRGGSgDzidj2kr+9y
97FiGFj7Ph8J4q8MH5s8dwYZoKVDGLDpT7ZbVnmsAzdQBTKi42nJV5rrySdxqQ1rjl7YoBGNb7fE
VzmWqqWiESKad5vbOmzIDOD6npQ7aaeR/8BNrVsJu4vxT4MEXo/eBcczIo29VBSlzAUiGCIfaf+a
PnVcQDBoeK4VZ0O90ahiwci3OvrrknANbtmRjVXsUVVx6AalN5GBFjgGInC52b1YClWb53G0RzDi
Z+irnM5GWqg9ddSTmj0CfP6CdUeSO23Ted3i1uNnitC6Cm9cRQGnPkG+uC9B9laP6Av04GLDtDC9
qenq7n9EaPXjLievypEjmgSgon1w5jq5NV/yNBLvfXxnat1QF6mOUqOoxANKhDfXWc2QHPjV7mGg
4W0PTPsSdH096Cip88bP95sydSaFiL7IC+RFqz5MOLqfKa9FTpRyW244kd86/BHYF7SCY10FWzQx
tpdOkNgz7E66JT5KpzccDe+kAhg3hpDi7BTbJVWZhjiQBosRytIb38aluVjqAe9GlXgCPhYzpA2z
93bfxcZCBzDIN6Iwg4hdMJvNr77gz/+ua7vyhHovKEp4N29crYRGYudXql1S7LtmvrbCDj2nMx9n
zg9ErNRFlEfI5zPpdRUIDAlZW9LOIAjHutBHV3keDZlEAu5iXXLowLgUmxnGlBXCF1Dmv/0qlcqX
7YvAVksp34NstEeWL3fGJIe0T3LW9jIsJoaPAYzlMu+osX8j312U+OQZiM939W2HcTS+MtnZCs6j
o60BXSj9o+1IK4lXMg+z2CTBUB/uvEuBw1RPb4Cd6bJcRWtplFSx7a3DSy9Mtj8g75K8anmHYUR9
vyw7Xnim2lH4Mecg89yg1M8ClFE4BQrjC4voxyEsn//OFn7wZhCoGNuZrguJUvbCRm9eH6NzVgln
IxpBvoT6Z5SKwJsjA7Mxb+2vdMZ5gQe10ovA8OxtiWNwcPdKmEIipSr6hjWcWw0VPeCW/e/qaZIA
daKm9/nTj6JXWPbNoDcVL8tcR54oXdOIPez5Bm7infg0b9uF9es2Sfe3Z7GaVk5inxUM/9XQuwjj
aFk0KpbLXWWeVqcw6s21LamY6SQdk/StJfBYXYOKE4EFnenrALypG0P5uRU0JZFj0KiXVsDXfJgN
ux4IFPD1crlxNfIsLR86MCiOnR9HEcSjqg/Toypk9xrjIn598vhYi/+HHYqgfLUU6MDJiSbHpwsG
gNCAZ4Oh/5AnAT5uct60DHbUUU2940D8ZLAuvHHKlQrL6j5eO2f9UsbO8dG18p7xR8AsxX1eAGOG
k6fgRHqLhMeaF0h4BPzFhaC1M5pdYMss4b5JkN2TybGevoxmWmNy4GgZFXbetQpKKj8MN7ME/DeY
J4QfjbcI8xoZN6fcBhPkR1F9kzf4vFvqydZHre+NBO1ec3UqS+naUfjxuYhX6JnMITaoaGjKdCrx
eG0vLoTJfo1BPF5nKxfSTDSJAq8tX3kGPPChQzPvspR+upyog7QkWCoDMp1hLyME31pf5RW1uXKo
2OSTv7g07BuzVf1809nl653UGdT9wxfNxAIzquLN3kq620kIJiTwAoIEg9HMXOCCJhmhMW5MOCoP
e8yNHIoVSreFpKu3Y3H5QN9YYqgeQuSgyVYSSZO19Nbyi65Dj6DBPf1OnIRUf05QPi0iXfcJJ4cf
6NXPoNsiEXAn0jLlvOAwNpS0ILbfLQ1TgivwBIJnAIaETJsP4UX4B8C0rh3dLzzmifEVQ2VCKGYc
QcLrfsz1niO/K2L5SZjGzxVaJTZi3zLugjpXkrZx4RjAIF9sTueb48ToDrc9t4h0B56irBvN5ohZ
bz7vjr0wz/rTM0qLRg2HZ81F8fzIfrU7hgci4oiCvJqR/lrjYdBpfyN7XHedpW3AzZvl3q/zA6gE
AKH7btaCqbFoaRBMuo8ryEhaD3sbMa1gsjka4M2/7G2dWu3ELhd/azxFcSGUHuV/CA/CASa3D/FS
XEynXpTj0+EJGZNDMBLXx6V21S3EbntK4Q3XtSI4Kp08tqO9zHduFfv3L4srBsakjoxXTzxzoXuR
+Vq0uf9p8XZDupNWW9upn4Gke6wHvSzpEXtFObrN6hvM7yATFem/MEveLDrVnbORG3ZPgwLmD0ET
BSrzvm9mpgU3hcVmGinMayQOEhKjdEUGtIzycztuMkjqAO8sZGdDrxVMmnBeVoweGmS9yFaaFKYC
CKU31G9a2OjSOJCEDuJkpLK4RjUgIJrGsa0fIPLJTupxlW9eLkl/wFEO3iKtgoFsg5985g0Id9PZ
+pqtu8TbiltqNQYUBvgdsVyy7mWcYX6qPkSKZtWzOo7H/AHYtHtLowumTUxw1ec77oI06qkvlVtq
JTrx6qmLoGuxdccH7fG4GL2RU1/g/nBNXTLJNQqnBd75HeAW0S4Jpuu+51qRNKMhWypQD3sThaod
OLyRJwL9hBGol5gAOylHIM1sLZ3jblAXKO+spc9nCUbFUq+GSWPBaAcMH07ZfBHdQ0Gw9yXBaWLb
8TrrIFDB3w5wNs0tc40c4CXukgJyd8mR7k5VT2qgnjwU9o/0Ul0M2FAQoy9yRsznoy8orAaYkGk3
EaDviAkySzOvZobxkh47vJmuKL8GLUP3QlpF8EwP25G8zT9OwTxRzta5G151GLl7BNx99lSc6FWH
2nPabBUMNdaO6Qfnr+zBKFoirvGQ8f/Gy4iTHIvIHEChJqT5sXcx7cLvJH+Kw2SH0hDzWieByLZp
Heqmx4kt0CCxRnecRSL/HQQuzw3X2em8cE3dBMiWyiqQec+/hl2sYNorv+l7S28rRZK+bWXi3T+u
zgKlI3iq+ydieC9E0tbpZQire3YfEKMnhnxp9fasbiGWeb7H/aLe7go+HZKSUqA2IdGU9MqpYOXn
woco30lxywIRn3Vh91yBqUeSFDU4wThNiHlXWjs+s5sOXNvgeGFxIK3LPnt0QTEJ7XRqQ9HOvPwv
EEwUanjHVv+p5cyYiyV6O3rVT836ZQKvnzBoA3taiWkjpBmwHKjzgjtN84wep+TvktwOjoYV1zjt
7oDziW5ohWskEINAQhgkroxHwZIf7vx6zEZTW8XCp+/lgY6rnSyyAOOsLO2GX+muJm2zvXX0lWuI
FUO3JjzawSkX1Jg3O8gM+vl847Jygi5fTJ0igOOYnA5ABQXNuFKtq5swXj8HqRZlxN11fCd28t/+
kjKcpmXDlqVfKCYGJ51PJpSR1YNwJTU6shclmPR0Yd35z1fXlv8oDQP8UG0KFzgYyhDCJidjOeme
E+rz09KYAXpE835jYivzmy8aar24WMTuA5zEHfSr69ex8CkmXV8qWrx+x3pfkJP50uGVOSCGcW4F
KddQMmDQBObEWAqJHmAd76YVmH5M+NryhVDiQRN2q6N5QhnW9pKlFEKt4XCpetD0LuzDDfG1Saxt
3/I9kn9gT414m82VTFO45fm2idpz866pnmIC70gJ2f0PIlDYxSqTiuT8s+kE+8Sc7E6vJt1LMhXX
OFjnRgjVJODB5ZKhqyH5hTTqL/0UxhrLDzjSGz1iQXrs0CdIDWifGS42qZ5RDBTxDqw4/N9wAWkq
LhzmHXpCJXVDfEOJ6Mus5m7e3gdVbgEdSvKOTOaDOKUBFHKHO+TN28X3o5NT4cemXp+s99iUdbQ2
IW/ukn3rHYna8LfA7t/efBfZKLRBZX09zAJc/baamYUeRBBMIBw/yhEomtDDTN8lP1S0zGhmhuMr
scc22bOt9ntz2Q9hvu6HxA0T6lOU5gRZwRfiuNFi5p02oH3tvgb/9EmLkd+bbtmlPvs23Oy8PUT9
epEwh+2v3xR3Xxuq0V59S7nqAWmiCvY59/5FoBAzkQ3wxHyjObIjCCmGZDdNeSg0/c5GnceXSpcC
+xpZz/Us3W6aJR83F/VYUyxRSUY1Edc19dOAS/4GV7fs/GDhCF65AawehghiGkXCqanYPxVoH2xX
2ZKOqMfRkxFK/ufB3n0amPek4KN7r52a/xNX0/+YgU3tr+psUPGPJYAh45gcqr4nxD4QWORaJPiB
YUtMhMU3dqMqzOwV2Di655y1aiAaqZOJknsQPOfj+t9sywO4rRMr+ONWgvfKuYkeD0c1IkAuaTqK
8D05wJjMJ2zeucCWzeHs4yewshyj2zglz3k/gkGPlgWj2WXbNnlxzZ+Pd6rqaGjmEJF+oVy/fRB1
anItEb7ZHjk4VLNFuGAVVl6s06AWEQD6xp7ohCscAkw0CEcHQhPyCEiKKx2Wtmaqyc0+NUKnbbde
9jwtpXhRGFOOQTgV2xxhFu6KWel2Z4n8Mxxdj7S4P3WJinfC6I8LtcMJkHBxym4q1EYDPLmTG819
89k95niVKmWqj78oZGItRPLxZBAfJH7F8hVnvA5vU04MoK30BeCl7zkancarPBI5fnNE8ynVfGdi
7nBhTLaa3iQA4pa/7YKBLi3s9x4oRTZhuVei3y4JYXnmjsMhlpT0Yi3X+CDeuBSg0kjiSnx0hhO+
5R/hy+wZ4QrZwPz4WIrHC7Q9pX+es8aKlO3hLri7aKkVJgVXQ61qUKac/UuoDCmfOXa8Ivsp415R
/FSURyblm8sktNqcIkGs8u15GhKJonNvTm/Nv2qaZA8P4mjIQya4MyZEzrC9kVavapYzbZMF0zle
DNm6We8dg3sTpILdE37iIrX3VaUVKSWsU5goRMyOB/wgV2ip+CLwqiDdSDScNVlTCISJIccibEpO
+7TeDmYD222u7+W2IDCKOWHUYb/GhXn+GGncOdp9rg/jablowKAcIdXDbSNWvcU7JNwwVxHfBc17
VlJwenwuwKgfiwodAPA4S1joHiFLU0W7iGkPDdCkW5aXD/dRr+9Fgfs34oEsJBlvobDw0uXMaT9E
fo1N5KYKIAJFVUvpT6pJMJ3335M3ddb1ax3utDL6G4v7pAuiQmnrw1oLkW+lsMAm8Mx96O4Rc/gX
k7eFrOyDduu+hV4D73p6IGePNqx1s45uIa2I8VxUFsD6OzMJrM/P0NHo74mN6URxRl6jtiRMMR+A
MYLqEsvbtLahidxpVW4jbL9waWqqh9wnleOuiO8wNmbJqG41DDkCUzPwICzxtqtxLYUhxov9OIo/
z6HPzeA4PkSftplkS8fbnQLpKAtWf9qG/8tLvCqK+GBLgQR6iwlgDyHX+apZ8xhbDgPuYjUBWt4Q
XlobYUu9NHTDLN1+wAJvOteq9WPZe47fFdtISaCV9ATLZE3NwI07zlOlqOcXdOEYaU/V134SS3/t
0ewn8i3NHhV3yK2vgdRpWUhQgQRZv4lgZr5DiJCnpqgK1Z59i+J4BkR5dMmCHZa09Xy5VlCAxeYw
8M5t3aBbIAoEI0Nijah7rcFlVVYHicSG9SqiWASGjV1tXTCtz+6wnylkRXpOee7btjsB4uQt3s5z
kw08tVCmbtlLQ9J3Hlms+EjCKNr22iq5OzrJI4lw+mOnt5WqShxZEsHclhwQSsbVcJgQTMMvMPCi
iBlRjs3kL/bMsGF/nP3fxihLe2S5NsfT95nVPIYUaCnX7Dwvua85RDfvKydxW12oPpEIChQFvXBa
ICeF0n94XkKJ869Tb00+V0IBRmAjQE1eJF9cK4EqF411kc1ilRfdm5Kwg1dhYuZ5iCPRx2efiTs+
ddxhFGwfXc5nMiUeGhawWqLjrL5Df8zp4xbBejRVOnQrjmWni+1j84jycuU7g70U+VZb9WTha3P+
tS+goA1LHdo+zQJutn+iFh0CFbQxlS1o2ODP/A96L1cyuJCfAVx7OM+5GdYA/Jf/fAEPItbDCnh/
QdqT01QowL+ZzXzNdEaZEk/lSSjCFhXYus4sciWjVDwYAL0GMUt3eK1hE+R+KuGk4WOmWsfdrwge
nj0oX8aHrZDWZL8EgDsCH73gcZhPg4aInjtWglSZ7YFxo8juvJSHSdKTOKoSIhZTIPeaoDqg6or2
oPnNx5cC+rVWI2q5UB6X9ixIpo374/apmaDZP7ZAo9em2ohpagumSj7c0HBLs4oi7pPUtF4yu2eX
uOd/fFsO66NxzZYIBi2QnYRECjPVmhpDmDkMahjCE9PYJ0mr4SlB/mzXocNe96GSNJ46SoBCfSri
zR9ZatL//IYjRIlDPvCPNGDdFcAJeGBQ3s/r2GSeS8EExjQcvlpgrMQmvP+n5P85hAsCVCT34F6v
hc31rgPHLc6XIBmb463Gj7bLmwCoTG1vBbNO12X+EHidG2VRhBq03iJbcNbRDA1ABC5fOhSAF00I
MSnjejK1G5/UV5XQvzuwpNxxY2Hrxzs1SIRHF7lbtIFeGzUeJHDOXV25YJB/sB98PYG2ZgC6//o1
hZduZpySO9Z00fAAskZH7WUt/x7NFeDQR/UeQOxE/gk0TjPt/BfVedDrF+k1BIwsmGY3e7G6i/RH
Rm4ZeMUSO4XH12dZaElzmiBhJz46wYH3ZTHbMXQ6kZlkTrbTHuQdhumyy7fCgMySETq0ZhQJawl8
d4Xs+0tFiAdzYfIV8Ito0jAb6Ez8jEdL64422vSvIvcWtonGd3V++eyPLKlD1uFjgY0tfdSVQ768
2PDp5wL5nBbnF3ErjY+UsiEbbYrK+NcJtBbp2SXl7TJxkaoWu38Ec4/Jt5q5omDxe1S5eNR6UGVh
ItxdjkUr/LOzRdczlVYQCw1JlmZIq3qiwtBBHKMbw/FX9eVw2E5yQRf7DAqMByP9LXYMSp/Lq9l3
2ZBu96L4qzbh8KyNwFUYO5ciCob5riJ2fJBzjHcAA5MYbduib9Pk2Bk06v5RyWC/tBuldlR4TXne
AukKHjbKdpuow3LRhIKhRUnRrbK86MNJfD0GKUAWON6xp5aRWi39KOOgS1d2uTAAvCTBJv8jMllM
a+SJwDzCSC7bwuh5F/VPwrswL0ozlaI5qZLkerwJKp6T+ifqxVCelSAgx0G2mgrRAQWvHxWwHhvT
hv8j/riogQT36GA8tcyDEiGJchWnz1QOJ/g/Et1THDd+GNFxE4FnZlgSQ6tiONviuwIlqQ6Tb+vO
X/DIBJJEH6t5eFi3JxaYqXh8FOWDwV0NJq3jsCxlGSYnLrJgoutzml7SZqdNjdzDifiwCrPcEWG1
h0TUnxEv+p5w+NAzrjGM4KtHL0ApPlnkQaoEc1x8BU9EExsQUN6rjBAzSLjbpu8+N2megOeTVaKw
Zcla6QEeqadUoxK2Dy2UJmGbrFZi6e3OQfPjLGBHruZzIdscDBGotfy2mfX9uREsm/lsUoV/G6DP
D8MvrTsPDLtQGATH9Vf72QFiD2OzCLDXZvsjY42YNilcJYO1n/1T00uP9Tq09Qu3LhhhXEldcScw
lQSbuaHVbUnWxMf4Rqs6LrjoImpg3iE+yDY+njtOqyOv4xVuQm3NMx19q4+Posr9LlktxKaUzOkF
iiIbt/rgUzabi+HMPqWEdPtvQPlmENotwU4xYPqb2oKtq3ofOh2MsF3LxloGmk6II9JU4oI5YkfY
VKO4w8OdnEtY/Tm7oQpQtbheDUvbAcVbI28mk4pUalGIgkQwmT4y7peun90d+217vlPJjscSuqs9
hWfd98GdkeiBuPFjWpHUf9YBAn0tHtsfktC49bpc21Tpbc6fKgHXjCp6KKtUNXPLOyOoGW05h/sX
O5eelXM7ZokUh2EEViiM/9XsuyE9uNraGe7fGSJyZjCmtLp6Nh4rIuoTJPIfyKmXFrL+QekgT75S
id/6uneSZjd1Mer9P6LehX1XN3Clur0kGhCYY1LKDRwvsvltAd4tWpbiE6PsWmH2ITbQP7GiEBg+
TfE536iL3Zw4g8yIIWCrwNqjZ5NWEqXwfmXvSpoynfqUQEVW5NBioEbANgxqO91Afwm6VJZNwCMN
K4uUaqcWEj6D66bPlNni3AAKLdaZhb794GzLJoqRdfKdhBb+eZlj5l1LXgU+SuThR81ruSVVhiOx
b2tGYcuvKQy8U5FhU6sE9PvycxdXvJvuW6peLnIIeKm4a3CC8BPsC81xpES3JN69NXnGCRnI/Whj
cnmE2czFKzQGNg6kYNAm9714zGtV3Awoa8uMFTrO2i6fMVk7AUTEefSUGYUdYvQI6JAfYQ4oo02x
pk1o6Y567iywv8DJbpWkbl3YNd7AUl0+9ziUZtQhRSaM4D0B6ZuSvlcGuBgwUw7XL4YxnZTc0p09
x+xe4VjgM8FPBrEWJhhIBBeSkcuFMrOvjLgL/KF/S7340NglUk99nacthzgZNQfwV0VHCZJhjDDL
P2cBiMVl4hSRIzKSEOC8bmrqDULoksXwYWapjPJuQ7XfCwh7FKLaKPzUlApNXLY29Z5wQS9maazy
71zeFrLMtEgp+yDBt9e6n1EJhhvYGJG+KTr7ByOZV7Qqs7yCttkDTSZbl3VkocPUhcDdt7nOIZAl
irY8F2d5a9lmGp7SFyisVH7IPuCrRA84Xu7ls7u/8pBgSbIlbRgMCvdJnbmElmaUgRnnFgvITvq1
Hl/Q0vJnl2kjNPH19avRO5X4KNcqqRy8i0MhVHHyYtGT2+B84kcqg4vQWCLQQXnlWfc3XYugZ02c
B2kyPC4Nji3iP3/92cBvWgLauwfZE2G0NH/lg0TNraxgdvFNo29KQfVwv6B3BFLnldpgJSgZ21c6
Z7Zv23s+wT0YV7ljO2O95bU8fEV7xYFU2yRQhY7BoH1XJNTdlY6yPIMMUkzpGdL59c+z6jQ2Xhi/
O/XGcXrQpL+lW3e49MnFTiXyC4ZgKGn3KVJBRORl32wDDXrxpngpYC42NkDZOZ+uxXDA88CADnYn
DSeRSc+E1y3vjuc+WVGhvL0oT1e0CCuJ47MS4ZTscGRSzAvg92TDNZ6g4hfY5r6SVNUNtAZS5u1d
Ezgj5fnahMpPyqNrXtNIbVm+gqUior2GWcKIruGVH/SkA867LIHcP+UwbDrG8pM0a3dnF5ZxhROL
eGtfH7em5nhM0fNIE+eac978/jYCzclVTY9WId5EYq6uAOSSCS2sX/4qc8ryKzb1d+gBO8fCPwNq
QsYCM70yP/m0EM/310W6i2E9GQG3tLZxlH5ads96WEgPFKMzi/ScGTz6/364NQTHx9fPGfVV/2/4
b+p+kTBoBnv8m1pBhAtFhARbyLw/oOv0WCRZuavh9ymNFn2+vr6pNHjF6/aYA7Uk2DK2HXmWiV1w
IFntX+PXMHd07A2tCcpiesEwgKyOXcS4lGguW5B61Wlvsk42gN7Sp3PprU2K3w2BXmZzpdncg/4T
ejHeOHJjiUqOOCEQlLjDsWqAze+JLS41Yz9RgFKOA7VWiOSEwnWa/S9uYoqzdb+Sns4M6hR+RjQB
xzT3OqF4p6vMh4jMaqu1DGohvHIwJcxuC6rZKrSjMt37NLGspjuNEhD7TzEL6M+e9KFL3268v2H7
rA2hJ5y40Z0CHDfRavSvb3sa4z3l5C5uNL28benp1dxeO/MXoeD9Mudu5YrtSw2j0R/2e1lk4NGx
MbJbr1nMHPIsfcozd68W7Ufp2H3ghBogbDyJXLoY6B1gmcaz4mQdCXnu25kHaOzSNwc6JXib5FXv
3OQn0h5Cb9bqoMoQMXtOFkKt9A68+PVraCaVuyi4hMolB5hFdmGaVhOBCNk+jdf9rESLNxcWNDLz
pucBlL9Vzc7+VSJHie5vgITNlEhXpLguvfdp6Sk9y4JFZmxUk6IdajlojalZnxL+fj0JIvxCpAeY
DIFZPHw0hOiL49bjP3dP72yfStiCDbHe4PEHJzs6E3piVsbqOMJZKeaGSESAaN8UWu7vXDJEvzvG
mzsXi6IxACMXXQ59/UByIbwE+o/Cxf5sEU2FBCSCwPKcySrcN1aDdU8eAuOKJvQmM1/rxRkmEAI4
eoKbYAxuTKMyKLxJHoJcfxteJpdRnu45QV9yasrjDMRw21KKD3UNL2l9YU/cJPMi76eRBGYSdQ28
VgAcbFrtHNO0TaKEu+bdIoXYFTqHNQjm1rRI+Zn/w79I5L0UwquvuU+xO6P9xd4H8lACF2NDbMCb
zLR5bJ1T9osvsELBKQsbouKNRBZRpwbZbha24sttkJnijcJWPR6YPfZZhDVwcsHHlldRIIw5oHcH
Qe5vvccpa73euFFgywmVP0hzQx8LYweC6bp7ecxF7CzNHxKihqjr+RcU4aIwmLdy7hOEqeBbTE9Y
pxzSNACj3cl9Q4AvWqBkj/ZFpcnnWMSxPIaO8PTf/oLqgCRnkINUPEOTJoBfraHrE4aJYErYZXDr
ANKEUELo+FrHRAOtqgj1mFudw6yEEVa2v4sq8BIEHdQHBRPrg8LrknR684+VvoiRv3d8aAjsl1os
RoUe/vTZy4uAwvNiMXPa6NTIbWcJiXBWFftfjdzM9YzMxhkmexwas3L3X2gzOkR6V7/o94P6wRhC
ypv4cKgMEwlqyyVaS9O2NDc24hhBR8vVbh8Odie354ItYVe4NC+1Fy4qHpjx18RC20TmmfXQYtkU
Tx81/wVQQL3+ohiird+VLNskwtga95+vHQ5T+s4AKwkzTQWMZYvXRKpG0/du9JrBoNHr/uPI9SVt
pY/6vAfltrLCEBH098y+70sYluADbkQEGCVUyRAesqZKHa4PAVzGCz1+LarbEtxk9HFlH1+YRL7E
3XwwOfRlUoFElaWPjGufyr1fWvDWuNp8NGW4+qDx7RmKuPJjc0IFBGA+Z5nl6hE0OiZ7p4KXo9pr
kwYFS44qWYpCBy61f3pEM1mJVThaCMObXfUB5ZlCshITmVzSX5znTpsZ1RD7D6Qz2xwjvMs8B6gR
FThf/xlfRxcsp7ueA16w3Rb2n+GZGt7hMnzMs7v3HBe0Rv3kJxCITcnkZmQU6DDzEvKc/LdZxh8C
TFH5Zp1Z1R/Rzf++y9/snnLZMAL7OdHEZ8CRA+fvU4ODH30DucD4f5wRzhuTBg1lW0KeU4bW8ohP
Jh62AV5m0jEWgy1v4FtWBDDvVDFyEnd9r0npc1Vn/Jai2p9/2k7Cer1BKsGjNBC1KVCnSKpPlCZB
5gtM2I9uU9crmigJn/ipAEy70AGGIGgN8MUhvY6dSZJkr4WEiATY1CQ4X2yDHeeHUSeNcOYIxDYD
18mKEd8DnRwalmdt1faExtF24i03PSpJqPhMc+ymsu4jl/1W0lvaB6y8JjuKtZSUXXyJgKJ2YKJ5
NvyTihznUlePrBOdX2aBYePmhFBcAue632llvBRGxNA3tUyUmA8pIJCTeOC/7ic00oQ/zPWMtzSj
5/GHrkfBjxCeAVs0qbFUgtI5OEYpYI5tryAs07os5Qe79aHQkxGSrr3rchQeQbyjmpS1ADCXT07q
bekzisIZHvX9cFtc8ecspAXYBygldmOKpLdjWdGHuJfRZVHQfleMLNTDuM0TdFKpb4Oq8a4zu2wY
O+PtuAZYSNl3fnPnn6in2LgNZv3Z76U/jfcjVyCZETl39McbM/J9AZPZ5/d2NK5ewP8CM1Wz9jwC
01kPItARfe/SlUvZSCsfEAr/2DARB5VT/g08ApFpmHUwQm4IcAmklq84TkjBHXxDXyFd/G7pAVTW
mz95M/3LkOXn5j157ORhrITE+MZqDxSIgSx2JKeUyp3TyEg68jVVP5hWrdSFuLOIxxYg5sA7K5Sb
t+pwqpww2JpLqE+3hdnPAyslnGX8DpJrcxZG+65C3gNh7U3mF9AvpervPO2cC3XNnq9sy2as4sNV
2kLMFAsUfReG5IV9z1FDMJKoC5vfSablN+0AzKMpW/kIghC35P+w+cSl/ERfD9S0pseXVGxt5H+N
aWbjxtvKZv5zwqbCpDAvJ2VE2VYAdq2kO6lkqF+nLmLDOc+MOOfFpVQ5anzlpAe2G2rHMAsXahBV
dd8FQzHeIFd+vRfbU7TV+40ZWSpSlfefBHibRSqG8r50rwDDpOLaEVQ6nJ80oTphx8XsEXllp7Go
HxHE7kq2V0FsYwc47KxY9IefVQhSaOQH/CDGHR7tCtBSKvdUInWUxN7yuUa0zz48M+L50X+sxWrW
84IhYsOl5hvkNgujH1DBEzYS+LIr0zJ4I+ku4d1gB2y1W5oOZQy6FD3ZldvcR2lwaY8ZviTpYfuu
qdOMC1SiatiJdOJiXi6JuScGlJ46OVjEUlQoqB/i7dWVDu1lCESyA74dMHnXEHzetqoqFKlvJ/l+
b84iCNUCDFh9EaOoVYrtRUuxaU9wpAalhXSnWed9/520jocqNTKKVbzz30e3rlw8n24K/VUhi2hF
UlHWt9lcYYC64Loj/JPNTjoDuiBZJDDWGEYLg9DUSRpwNVP2trz4cvfNeslHuZURhmiME4falieE
VIddrQGgQx3P9/ScoEk/KMYkxEy/0krkwOJjnQYLsgCdeYvl3rLds7wXcmyXmfYd2wUKZGtjbQKE
ARGswVPycp+YqzF8GCefAPO9c+ttu5jYF6ID7zDs2zdVtuVzdo+5ss0F4vdaxxvUGTCYZW7BFe9z
36IsgybgeLiz7RZ1BgH7tvmQ8TPfVMPmn9wEHf8rxMJ2pg2+h55DsH3wSX+4vws2OOgPeKiup6QL
6HPZpfqv43WgcXAFuNaA24moisl4Jyepq5LFJt+synmt5oCy/zjxijnXA0THQBcZF6/IR7i04v9T
55B5w7z0ItI+qFkGnILXZF5+R3GiQ1riuY5zSAGLt+2OdeY43GhKIvzKCtdEoCWuzYvdQko1xcoS
yOrkiIBegDqkWmFRuWnC3e1rkKf+ge04XwS+Ren1O4uK6JN/nAtEdZxreSiFZIu4766G46GSgZPj
dABahYutsDEQyabdgc2Xbjrt8r6fK1LXGbMfrqUJ1LdNJ6rqDBIIT06Cv+56Hzaep7FhDMpRym91
wm39XyXhh26phIKl7Q4UCBX74uJ0t9FtEja3PFD2rfiopu7q+mXVFJeYpFJJFdfMKm5H7Vh9MI+G
35A5/RCeBIyZYsoPM3dDwySVtWD2UaFPqQ63Fi3B5oifyFwBNgNjE/0Jgwm1BWo6d9DX0LXlj1ho
8PUeTCm+OOY8Sjupqa0Pnva4hNCMdqXBfjBEUDCXvj2+oe+y1ci5SPGXz+loXSi+iyYLiE9tMp3P
RPCPyMQjCI2zAy5vIebmo4hab/GsRM0lRr0kwbS/HHr8jOLLFSgBGGZqQMbyZiwPEeW6KmVbWTa4
2riky5/Kag5pqgvTfd6vI9ALXTF63LW3no2oWe9mpmKwhlT/Cjmydt42w8NDENH+wQc8B2p+9KfW
20pTKRSHUabtxd5hoNkqr4D9X1uj+lgLtQTT+H+nvwB4QxcozLKFqAGlloVLd12ss79OeFyibmOF
xs36k7SMa+QLeXV7DlCfrnZ3LAs66Yl8uTVKFcE0eHRu4/qkCICQOj4OUQ5A9O00r6iSZtPO3MPK
kw9AAPo4mM9y/dfxdDjWgxe7c83mCdJRVFx0I1h2K3kHlKvlAvE+ZIfmYMsKbtJG7zBI1Ajlgr1i
Ke3asrUNWm8gvelj+N9SN20s42YrWE9WKLSlsS8ZLfX2kQ/mSsQk8Mae2jqdZm3Wpq8drb9IcHEe
6I08Nv2hsHh4SFnhz1P32aoBf+UwgW6Dk+24E7lZAmvBQzwjcDMbP4GW5OAs6niTMBDGO/d2ipd2
kSd43HST2DySxGZv7gtLe6gEL/Wt/7vshfGvXQLdlTRPUHf/b8VUoX1f2e07gU1hmO7jnhihBWs4
jylCp1dTpglvzj7I9MkM0nkkVP0ItdNJXlVejJGF/e/TFJ2Icw3hJqmcR4Mz2tpe2N2ld5/LhIsn
JjHM6ZG9p7meFirDKDQv+HBdeyqFJWRxZTkwdMNx9h/cseC6XfQ1MgDVw3TkKxrwpjjBcDrxoVvc
GNARQg6AoGCFFhc4hQGvt11CAsK7sraWAYSHIcac0kY6N0hK7TyoBPn78nAQDr/l+VsvxT/vw9hE
BEQiaOkXW/Cc3+OfiiN9NrzdumG6q5tsus+AzjCuCN2lBFGyeGN35HsgkGThdFWDs4KL6x0it3GE
NSvrYf6TC21ztXcySj2v9uatjeFon7idwXKGdJTgMtn+XxnnnYOaPalOEmVcvBVjjvNjXNomQ+g+
2DN0+Cag4DV48sQQ5EMlKEXdI8GbwmVs/Nike0Pac67gxxQI0A+8hnTbipOu8aEL4cTpJB8zAIkk
ITpEqGreSH2/Fu7zmU5bwxOnFbN5gxcty/s02HTModFk177T3ePFiCyUx9pJ5YUpQfh7kgC+bk7I
dR5apTOizaY1WE4nJ+AHNdViMu8Op4pb9olkhDZVikzbhF6gSeWszTLZFil7nYBXYIxVPWWAO1G8
+PYohCmox3TR8EIuedshoR8Qa1VqWiU8CCALVzpPCmTTIzp1YpOKInMk4lxVcBd1J0Au6aycTUPY
b47nBJqJJO+Wi0A5hw7om50SFTPZZLKWYycDSiZX+uTfOa0PAW9fFYEsV4l/qv1IprxGdibucE6j
LmRakW5S6HWkaIbc0DQuhZEF9wuh4W+LA9fKfaz4cpYrWb0psjpvxd8mj2RDEsSXldOq9rUqu851
MUA4VV7eBFs6sQlWDBUaOlI1CuR9Lshbho0/EQEQ6lhaCZxcBQfW24kKzRViy1EtEIVRrxK8uU3g
YpubNjTMHFprsNR3rV00vMzjp/48ug6lR/KAxSExpxv8M7/ssnrIhW2J6/KYwlIcznutYdaP50rc
GpBE6vP/aclgwopzuqKMCVDIV5hGralkNyL0mlWEpBs9woN+XGVI3cJLUzZtvSAjmf1FBrcliMiP
N0pHvRQavghUu0mgKlyd95eoJtsRKlrKgBD1S1A5vALPQ6EqXWZpWVvSf6qWJw8jeIQZBOlPiqV8
wa80QFIS/0re9IqSZ0unddcqB3Av5dY4B09oXdqgirFAA0lICOReKgVpTK0S/sbLcf4KbO+bRhHS
9jgA6MmN7JyUVjL6lL6pkEE8BWj1RoSXKBNt7dyYdXxkOjjNmxTzhkzE6U9Gow+UnYRXEZ5N8P5C
biJFfEQruGaj7Ocz1rtOzN78r595UQfKxMQsUHjdJzCaIXZvzIHGgNUf4lV00iTYf9RZ9ATsNYmX
hKRZZyPAMLZBb1kA08SlUNOHKSCwkeyIwlm6CF1pM1qcaywf6mlSa6H9R/BefvS8gUZlQn1s+ytF
4UF5ls35TZ+RcF9Wy1RTC8926Xm9QMPNa/5N854IuGD96FlceogpUEKXQdVAqbKbRhcaEAEmtF5V
+JlbQ4Ui8+Uf48ZFJb38w3QmuMscyxLBdrxQ4nf0xGBKvsrxaaMN0CFWImNdu92bhkKA47m1qpL+
6//E+TS3dyKnONuOY3ZrPK3Iyv8YnTxYK9XT1GU/V49WHxBvx7O4e0S5HT23Y8l6q2iE34G3lAK3
jtydWRCa9MJQ4msrqJ8yLxi/A8u17XIBLEFe6XbkKJPRmkkYucBQ/Qwjcbve+GNaVS9y2vt9rLA1
3OEdJDBnu2/gP/ZucaeHh2063zPzWX9qtE+Aq4KrZXyp7pg63/c9IyM5bRrD9zi/qFuqHDL4w+xk
qZBXBOnwmIPwXL4E1huu+i6T43DzwSZNKduFQoGHxPXK+RLQgJYShUy7RGMXWDYauwcsO3nqmUrF
4+i+ZmpNqJxwdwscKdTTyY9EzSV+oAsw9uRv3aL7k+2B6fPHOT9fq7MO/TDWZdvpUyO+HjSk2A6h
UiwSuwMNyz++80K5x4vFUfUnnsxHfK5M54scPdPFw+t4Noc9rbHmU0shWpai1ijbNkEgn+VmL1Hd
+zPZaB4d0+yGoq6rSv83yccyBgGH51RyNBHYkOnNmw9yZ3GdWL0pvIasEM5HewjGwGdfDUmsgxSt
MCJYmUdvMFkq8Qrl99YSpWkv/LPxrXu7CZNNAhNdsyFF+wwA0T5IiuCg8AvUhiec+gBIMRGsK45O
SRgzaBDIwdV2Fu17yyBshHAMeODJqNB7clq5wTvzRLGy4FPg71m6Xmi6XENhmgZb5FD4IfFYHNL8
g6Fjkd93GOdigUEgZuQvSa3exVsjRZOjv3hisQemDn0gcQDXVdMp77ES8OBwissJJPYEHKR30IGP
VoktoQDc1Qo7jBAP/lGNH/qUdZYWDsyoKWndX08CDMol1vLC57cl2Vq1vbITN/65ajdbc46YyrDA
FL2+taZZd82CPcmR20DVZUFOHNQkHdjaTh/mzrzLOyMPERVfzNxSkij+r2JUqDJL+GkSNndPutEz
vmqYWZLULRJvtBTy/exVOdZ0wY0BhvAhnFZYbJhgUESite312YSSY46fPMNa0Ts95C+pdfYPqGB4
vesnBMvQCsG9mF6zEJV9TIwQvLBmfx+VeZgfvQuHFWqk2rqnR09spvxpeFuy5DjUiNtI4Qaoa6o2
dZ4JSIO9cj0P3mjo2kx2BFCZI5WMy9kMrgGO2HvqEFITNPB7/M2f3J9fIg3srQQtmTi7LNTyeCIf
vbiBcdSmytZ8k4bt7Q0iCQOZRG4JR0j250OFa+XmCkGtQKoR21O90NqN+tl5nlkrn/siRAFnTLEU
LrFNBWq9Pq2Bot2LsZqpfluN0c60oIz9RQVqj3H/Ykxl58Bd7RyBE1IderyLG3OyQvHrN2EsqJbv
JJtHfqUhmU8kkwRG6vb9LVMLgtFXm2N163f3SP6nla6EWT80I0jLXAfpVVVI49d98RsmWNZ66tY5
qgBRJ3he2zQ58al/ZRv3IzoBt1d3c8cLI2BwLnjFmfZ6WP0y2503m+VU1Nehf2bUeC1iVq+g0SuV
aYIqcqNNjk2VLEqMMeEkVQ3lfAQRUMM9fb1e0KCH+EPeK7Npg+13qLJXYnAwyIagkWo2dK60ACbU
rj387b1XxjfNZ5bj3PSjDaBxy4md+xRb3L1OPAiyjEiNTMne0f8f76wt6iI73JYxeutv8+1Vmvf5
NCwgfLUzKtb0UhrTt5CtHrOKzlishvxIzi9qUil+j2okFbpFS/KI9fUWPpLkKyGnvSdIdaMCxs4h
mnnVjoQHxH9vI5EuZ81kw9bKmyLNT2t2kWiSpplHLO92QCKGhiSxgb3q6jLtEKKtM+jcFpJ0aKB2
Zl+sMOA1TANbJhFpgyM8SbAhzYr/J8hF0PNG4nJ7KyOxz6vAizFBQmjg3XAE55jf3KlKAxjciUji
zMkpl/f1HgnMVpyKzvRBSFvgicO8zDeDsOWTFeEu1knufsjAz84itl2fdkoPaW2z1lQnyAyx22Ui
Lp213QMt/pRISauqie6KqzuXgvXfaXzlCRqOfJjcoIXnNyc2F1eK2HQEuWQiljzygTMyoitnX1SP
wVYN6FlUS1EoyvJU1yMXJEJSWywIp//xNdbnR1WfpPT2q5Oqm2c3dQeAb8IklCnOjNYCDJZ349f5
xbJjc4GYcz9zSQR4fNyXHSCA2r6ZOPitTiGTIFMbVVW8vmKTrtXea/TpJn7OTVbAU2CwmK/eQ/yL
Q861qTn6/kHzyIK2JZEsoJabwU7Y68ff2X1KlOrcepbjj96J9wqrwDnneSXFoDvD1/Jd7gAOWk2u
6SkWwW3mj6LJoEPaGxQP8943PPfLrk+XHMYiqWOxGxyqu2IzPgJ5B4C3LlGi0IYIQYFuPih7Rtd2
H7MnUxoF6YjUYURVuKxPdya6/qF+SBWTgaRf8BEV3J2oywZO4WAeSb9AqfvuFV1IXWxKB5JsNsAw
l+haNosHh9aOm0D86Oe//sRCxydmOFTQuGPAiQbPNpr1Ysxf1azYMjs8QEbnqNsPzLrUiYZim4Ge
f5t9E941DXyl6ZVmveTRFPzqPxW0/8QKGv6BZjlx9PpYde9N5e9RbxO50USyCxC2zUz2OiiYIDH0
PMosNQbX5mkBVj6jxsjAglPelBSSkAp3gnoJDHj2vUNFq+ODw0/lHJZQfL2SfbwBEMRhJHbLJRyt
mlzL9dGSWdxd/vYa+GWcK36zAESJIqVF7ERTKDoWuXb73imIpPqRR4EoemnFHX3fSIpA9ppKhRjm
I0hm/FTkGX83Pxt+In+AQ09WMC6z5Ypw2wNVsg9KjDxkq7ILNGPjuJNHAlzB1v4QG+k3RrcDDlK8
ZMFHH7SRVxYgttClhvfIuLkE2eqI9TGuZ7jbYwLO2Z3FAUt+Lwmgidadecby+DYcYHNinsuwFbRS
iRP7ZDbG3b8V0RQAvldhoilDSTHs8eIkC+TXwk9iOOeEflrH4jLBYN73A4auquknB+E47wlKTH6b
T3ctwT5ktOcIEpZsS5qKjRnugFtuF3iBaoETeYeksmufm6oinAiNrBsvMmwlXE0WjHkzlAR6ZaE0
4zvPFHwaydnJ+UQJtIVDwUgTbai2y8aakvgg5M6+XC63gLmEW6RYLAVEJO5Io24v7KjIww+PWInT
Z7fcQ/ngheSJsASvzrYo6IkTDA3Ns8U5xtQ2SPbLU8Lways7YxbNsSFZ1x0FNO4+Uk6DCKDTvYNB
DabITjY2flJFHCI4Ybe8d46rjrAtfcm5kboIsgFvAiwu/P7Cq3R55qgLwqKjbQZ3Q3xsRKg5YirQ
/qgQjkYnoBhJzOF8NZxupAPml8Bp1n91mdaIA1++SpOzfWPswuDuhbsV7YHyDyM6rgZOYoPmVQzi
Pwq2QhNenbfb1eQPYywE7012xqearj9fVhEo+JsLW0LT341J4OtapwD29wzt/zzPSaTadTtvhkdj
fDd5y143bx6nFWFWsueU9JvshZY/R5Wfs4HElS9FJTLRMfVepIXTiKTDrFvDljMaHGMCKmc8ec5v
5W8gYdgBD6SEmiOQdtluConiOYtbQmZTOSrkd+whxxZcT/1ZKVTpqmWM4pgVyN+On2eLu7LEcxwR
3jm4LnVG9TawXvKVtU2XwVk5tzvqxO2ONfobavn/SgmQX9Gtu5zZUyLzx3RNhO1539IyhBVmpEN+
KY9WOWPErqGyVCMDshV2gWiyBrvyFtR6zZ6sra67cuiUHjLOMij+X1atQKzXPHVaDOe40CXRFBB+
LAbiLGaiz06piZTI6etWMtQLgvx+gdwL7ic2PblTUCPTweV8YzHwyoMtdQ7yZy0OulEa4hARaLUK
grywyJQIaUgmL0knGgzIEevyItLAPLmpDDjMXjKmF9FWAGbtnHDa+itflOSUhlk7Ay8n9w1d5ALh
q54UhUxwsadC9Z9pq6s2SgxOk2F/mCta196xgjL9sD2sUQaVSWLTTF5yvsVHtw5qK2QSg562K9Iw
Rl7JLaKpyiXWYwsNHX1pwqOacl1z62Rn1JFeSlkV5I5XCuEiiHy37sE3aEsSoVMMKFBfabc8doVq
+chnXgQOszrbMzuJS/2/K7P2/BZghYgldeNk0C6oJAGlxa+KjjhCBkrkfKRgGf8PuPSBXm15tA2p
2tAhSGb/Np0kmqiUOlI82RBLZ0BijLdWLbRoJYgn3LX1m7hsx5AJ4z+BRwc6L1zN9eb3/qH949IY
+j2R45Cx/iy/s6cF59oGyXUoVQwF/dQk2Drg1m+V4AzJuZePBXd2hhCi38ubL9A3VgEUQdtHO/4d
TXXSPHEy/Ng9g7RsBL4a3tphVNjFqBwNTUicg7b0mCsnV4fi2OBF48MTwhcQ3Qti5nmqDVVbM13l
PscC6fz3eD6c7MEK+6oeBxaoRTF4ZxouwGI0KoLf8faQOdi9HgZDAsrzTF3P7t1LJ6wUHFc4RU+u
6ww+502ONby7X42GFLhDrRDsCQZZmGixhcR5n4F5F+sJYkTnCZzskFtrJ8BbSGzVnCq49lazPfx8
cUEsDPIBotDm+KODmIgczw5tB2gXSk4LY6zi513gmdNlVnYZFvhcBunl5IuW2FY7teicenD+2dGe
jV3isuhZN5tib5dOTAhPZMrtRKhO+EHrFt9VpBEENucDk50TfGnd9ZRVXGytiw5s3C14h20RPBoN
twJZS9G/TBB8lajlRDaYySGgdjjtttqFdYxwl7hLje6uHCswnXxKvKEzwEC2nI51uh5LjQfyscE9
5n5RXuIMstwYFuxSRM985L+VBC1xUSKVhhdYOmB7ANf+ogPXPg2UJa/R2z+/waXzHrX6eYtoOHVL
l2nWvi8xHOinA9u9ca2H3kRm6ayWorHWEpkf63uXnMzpUpjE27l8PrS92l84Y1Ng0rywoqDX38Qw
o8eE8eTcrNo0a2l4QSOWzW36VFSGRZg6nAyBrhR1Y+Z1UXX7ZUUVadJV5FzcjZ6MP0SEYAS2hNr1
5jAZxyZH6R0aS6HqsNVfX3zoHSUSGd+5ws6Y2786cLNvlbfopOneNIKsMxKI0Qfwm5YxFVH2nTfH
dqSdM14t1Hvg7mZkrM5PktNXVFptOtSZf7S+D2A6b3+sqTli3SOpScKzh8nvQn+8bQqmcsQilA/m
iwBo45Z5be2IYKL46Dzen9bqjKlYEY7dWGe/lkQlhK2pfjCqWe+i5wj99MwEkHo3XPif7DUeukCZ
HpKhBNSm1/ZNW7Ox8vDfKjxWUcjSOZBMekDc7yrMeixz2KUrYQAvWL8L4UlLCOEEds63aWHSc6eV
QnFcUXorGtmDniW/+IrGwxKE+bXP/UTtFLpQ7nRTnuEexKjznSjMMQZky2W+TqSKiBmSsgDqNlbG
Hrt0GsrcH2U6gmSjf3/WUWIkEny5Q+fMRrs46QPOv0Fro+/cxuDvwjUZk9qI96+hb6kIJ79Crube
+vgaqUeo6tW1j0FoiWcIZxEMZcksQ4hS76mjX+HAz3VDmm9n893FTtZXyQfUXfDqdMh1YAznn+oj
Zk5aI7cE2h4c5HSenud+7eAMGiotUaFoFicWhdH1y/kcwn/kXxRiR/6/2JlW7HR32mlNGdYs91do
3jM/fR5aPzIa8Cx5UHJ3pjngPsPjtvVrmGnWDU/7/61XPfVfhOL1v0Td3lt3T9RebgPae4aniB8s
4rdmC2a8utQ5/0EnByPscYD9e2bhBqjlyHNEuDGmBysPf6BY+hz2vfP1hNkQGq5TjAP5MW57lmTz
eZgbbgl6CGfyV98C3gM9AoZzbYvZh4+PFnaMyfscyS7gyvMnqjVMq+pOICiXzBpoyr4IrTHYAxQq
EwvAB6O54sCONOdrZF+liVZRuJhrKURo0ATRxAUDLhUi7jneZHXVo48onFn3xsxig9Lo1cEV8gGb
uKjoGhPzb0SYpo4RtbfYew8CrTI6KnTu0Yvfkt6/NRSIBSTzrm9sPtWLNKDslo2ix4nNeYSRIyBx
puuCH3PWtK3PeyUqpm7hVC3lvImfQmvFsoUXAM2EGvdQpVIfwiIEYl5WDfn6ixUnrvRoj5s/L8hp
hnnAze2smYK9rmvZOU4tn/C7WStMGhMAmFqbHzCsXlQ7fc9FOXjaFkOdx2aoXLFf0dlgFpFz2kAH
nu8vnMLnG9TK6UF3McyVDFhCbyzs7r6AYGg5kAQN87RxY5iqxpoF63XuaYvUnstCw7sbtTRr/fPb
wWhcfgUxmK+RNaIo4tFmun9BOOjYQ3g4lj5BN+UHHHDyMCu7pQHhQnzySmYrayexklBO8vKN8kbL
ZH6izByhzx/KujQ2N20WYFrorTU4eqAfMDmQQmgq5zQbdgITmB4sZK0aA8Sl+fm06hY9AC3yp8Yu
kso5SazU7q0KYoWTxEFZkhx6tOAat2Ypkha6w/t7fpH6V1oxkO4fSttk/7C+6VQM4bQcwwqy8mlM
NDCP2nl68xbPeYRNfsNFQJAFiwcf8P2n2T5NxGu7iL96SfyytuZSfIbkkTJhxTEG0AmuYvx1y4Ab
OoVHi9TXrqSft/KZ5WQKuALmA5/kO7oolJR3qRqeAZAVJs5BF94di/eRQjCShOgIb9vfkV2Ciu94
DpvNig5uEEqe+61EO/N4FAaxdt2e+YX1pNqyO0SaoMH4FNF1KIA0n/+2C44apLI9ia7ac3QSyYtu
Ymh3V6KezLvGnKAxX96Q4DFY+JReqn9rj8k8misNCi6gT3q7IQsatq7AmXAySg//mma+49sVmimL
wyI4e4ToMKGIdrFuVYyB4Ou99dw1J5i9RpzF45iGIGdJgsqU/hygkGgMlH/LZKBHgk2lpg8k0IR8
AC/+rnwjYV5CViFOOj35BC0dnXqkw8XUbhR5qRqeqOIyGhHfVuQXAkSC6o/N0Tzs4IdXi1gKCZU0
EzYWZiMwj5ZRBw2SlW6R4HmkMEET2jAlP93JG/2vBjXFXsBHoPtXqPlrjD3s5ofSdd5z0gC0U37i
qpWqvwgF7NCMHkZMbHONzT8n162F01LXBot6Mjhk1QbHs7n9IkWa+vbO4HBuN316XiF7Aiq/Xktc
MhFJrooBXS+JjuOCKL+5KXFBcUHyHeXzkrDVkNHofjXnpm8ZKNi7ZF3D8qIUZvzHvtgxvBYlUDOi
6moKsc2aTVIGANCrKe18VKwa++jrPYRgr/8vAZGqMM4ZThy/P9+r5nKZF4ncIQwFJmqhp0B09Lv+
md/qA+fM3/ZAuPnetU+XQMxXnnCt6mm+wlLLAlzLrF04Es1kmnp0MKoJea314p4TQ9Kt3hGyupB5
/ltIjHyVQLP0AXnwMPPasnnDGDQMot8dedtbKqC4cbp4wje/IiYBDOv5pdCe9jaCwSn2y3clcrW0
pYLJehe3KZR3NhF2QGOhH9p4Zk5cesKoQyzTJahOefHZU61QKdJCTDtC2FZC4PvYv3OiWUED9aKJ
4wQNBkGgJzXbOlYrLo0PbQethb9ewBNFTz84DwcEUt1d7cgnTOtoGps9dyrVMDsbasmN/G4PmM+h
+Kj2MU7FT/XIosbEsmwjAc+gxwb5F13udCpJTfA4QagNhtpOMIwY+zQpXRqpEY+cyV8pPsMFYZAg
uVfq+TbHYruiKcbUKd6xKliS+yGnkru8xNt6aYZUPQyy2ONYR0WVKaSK8C/vR+Onn4dJJNvymaLX
9OduPWzRtesjg5FrUeIQ4Amiq+9AnB3ANknPkHVQBY0wq1EhzAojJPd+F9LgIQXuluLGGRQ7Qvkt
5ZNYeAo7njFKtaIEDtaGc8iJN2LJrUHTZvP1R3dSfWuaMNZo7O4jwzrkRfe4WE5iGruAjRVEJZvu
bEkJvyV4dmu5d990POKLx828D6KZUVLOk9BbxX3T5jC/24samdvUptkpdvuw54fZs0ItJhMnCfT3
1Yh0QUhp4ZQ2uO9Ej+MJoPufGuDua1Idgt7d2Br1dhOCyHq1s+g2z9HrgtGus9NZUeIjdE2fEO3H
dVJU40xEkAfbGstkFDXv4zKg729WrlPsKccB930XF5KPUlLSTrppLqepLd/1QLnIPhZvB7fcZJx3
u/ubFCb4XfH0mJG6Zmy+mg+YWpa0Kx/KdS7aSdMzEUA/zODPFxMGFCacpJVYySZ3+zXR4KOftceh
uMbj/ugzptJo79hfzkd5/g+y5owjk2qRWADlo9Tms0PosS/28i/PzG8CwoAGP+ua3h+FWME8FVOK
KDyb0E7horC27rFwUD9R+lctfE7fd00XCsMbiNZdEDjaVKMksyaUm9LTq89aJLY8j8yyH8W7mPkn
kf1BlHMSHuH/9rRnliGOPnsTiKjBJsCMtb2RR3Qls0WY7tLxdabKeOqmn2Jbi9NFe1t0TJg/MLm2
RxXGLnzJatScEOBTFTrue/Rq38u+2PgY3bjn75yJXMqInbRZ4q8gmZv8XOCXFc2WNaUC/fUOib/v
a9NsydCqCxqFlPScQ/oSTr7L7kM2OmlbbsW0Iw4UO++xwCXVfuImckIsWfDMsAlloXnNPYH1onsi
/6yH75gcRLlzrltTPPv07WTgWZ47hx3L3xkqUe7aapUzpqdm6PKhY3ixqtuluObq4+W1QnGEpJd9
YSutu45zAnqr2hvpVq00qM3l223pxAZ9G25abO3A6TXpWbxZWmFziK4lQT5PFITk3ixVhCNOqu8k
R2uvjHbGTjyd29vEU+7dXxFMR8z9AHfbGK/EFEpKavb2DUN4K0t2xa/uY1MTcCJkBK+sK/b/fx1R
WrTNdBOFoi629xAa2me2sV8dZTh6C8x0Y4JJPLK47Z2T93d3nw0QGQrr3Lvqyx8ISCPu0CHyuvHd
P23QW3tZdEPcDQ2pQAak8BVbo7dJt7LLtxk8iMAcLDSZHiZyhfs43PkbxhtpiiwSARe9WGWcQprY
ahs7byoODXaTU1/IpheYO0SQvIt6Yd2RuTaH9Sf/0NoFqM7xvjmYvi/HXRRMu3YCZc5DwcrUCtcd
4BLlfRU4UnLawbGTe0t8h5Ds+2ZHR07IrkdRr6cEGhUvhP7kmCGVZoac0ae/g9QwZQGnTmTfxyXC
fqiV9V+sRx515BGaf6jKdVX1ki6pCowu/vqptMC9OCaKxvwkxOysngKppbl211K/ZgNN45U6Fgkc
lfInfcuQ2Qu1+7zU/WmyrG0SJXub1ayupcBX8uedT0yeFm54qHSkMnyD+UN1Lx8TOBJ6D6jlfs0c
X05qSCqAsrfg37/UK1ugshpi9nYGbVs5igsbPq99iz+lbxGWncQh41PKO1nORfCT5QiVVLvT5FuC
C3Cyw4kO39YAPtVKEQ2fxRP2O8iMBpIhoYgSKX2u8mMX73/PdBqUKaueXtIRAG4ZQYOltnkf09gU
Oi1nBuMyRrVAHMnfDjzclB5UXpb61l0PQxqePY51fWIXY70v7S/vdydkdjhYDKCIdDbH0HxI1BCr
M8NPgmIFY9C3u8v3JRo7VYZNBt9iHFRZxYXiMWPA1xKHWFOTTa+ZqcQl2N87RVeyxnJzOqdYfNcS
+yU3T1lk23Kcsg3rJ2YxODFtOw23SgwSKPTinheyTEF19rP/2kaqLm47vvwAqtjJUdwzz3/w51eA
3R/AFvZgncameHNw6kySJuse7devJNfblFawLT/cXDA39y0i4//2VOfdnFdIB50rf2Dh5rD9WinM
iUqJh3Kopl6les/lk/+D1vQl7+C5AL6ztV+MZ2gMS2sKkatqEXQ4VTZ5IPEcwTlaQ3nq1u0tJc6Q
JUHED2poyWB29rq6MwlxFU44v65M89Fy4gHsgEEgNXhJeZp4eD0QPfjSWQwsKGPryVgz+oY4044T
k6TC1C6IhgnJW+AGDLqjIA10+VzxxW9qq9cSdKdFFVVtITyhoSM3lIbq+K07nRaS6JeQW52it27i
iFjSCu18flHJZ9jw/nZtu4vsMuAU9TOIic2orPT8DAcVZrNyZklv3MduNvRGYVL8BFpMrgxnyTAM
oayMY545VDiz1oryQ9dVSjG5drByEtgSMQQ1UMWGkD1uI3V2JLEP+1GasAAw3IS81VtftnqOuxb5
TpG0+ig3ylgBZvAaRwwEr3GIns3V+DjQFkR67jWJA5VHzHoytMiFOhVs+Kxwv/MMwjM+StYC6WaB
cwqTiUEps4ZfirDer5gFgWcFF9e/YJ7/eGlMH+vBy8RP6ThvATK8OtDgjhQ0zxNPurpUhf0hWe6G
+ifq39LgdyXnNbz3/9eV/9JHIa1iQhCcfeQ+6lLCdMgxDdRdQr13R9y6jUvjQ641PHWG+QvJM1yb
saemvXIDWLNvt8xEjAiZPrZ4n4KzE0znSWquC2knTVcvJSFph/L8mp3qpBcCe0Nb4vVsSxqcBzmN
aBA5UdP0eV/h4QBijNqrjZnUUIasBQmXeraxuBO34hAPcRsOdArNpEYl1oDe+Vo5+uSNcgxDnmwy
n07tFA0sqaiZWyTqutP4h8GJS7x8Mqfg73HjFNHPQ2xDb3x+492vStuHqeHDcnhIeMvPBhuOxndr
VGSlCp7BHIorXWYfgMOKz3X4lNgCm2DROJL3xl90aDwynuX2LMk2lLREmu10liB007sM8AM55gwy
VkxhXH0Qe4WmWVJ4KUJkghlrYWtct/ComSlxk1DSX7oYrTW5m1RQuNBSGhEoRAh6OGompnPGLR68
ysQk6nmJvSSgi/YLUNOBsgXAwbkVOTEhw1jAVRtJ74j3tSEiJwC/H9nTmXJUqhUYkm1+fGYLIWo5
pejJlTccl4NBe5JPSou+lL1nbIk7GfLxDYvMiQIWY04pkz5+e/IU6cl+Nn3CNBGiFvODUZ2WJZ4y
BmICBd1qdia97lRuca/11ovCF60DgVrPuLKgwWF8A3vbrGbC9xjFOJMLJGlz3e2VYPTJGT1lMLr/
N3idhJQZo2Re3DuApoO4FMvaco/jhRcuQXpXpLJawuM/Tys/QeJAZf/LkdHXdDJut6OSUWFFqqYj
omJ2cGH3bok+kW26T4fg+YAMGm2O6RSOh+SjhdBCbEEGrHKYOyQpYRd4/wG2sGTfyrvRH86z14iL
oPSQKIrIUQUaMDKjSt0txeEhN7eB7013y5ob2AIeBI2Y+/u7EyKBOZUhQjckSNTtZHnUR0zxIZWl
jwo4y2uTVAMWxH7O3tIOpP56nVb9LBRQjnQ3Vl3jQp/XX+qWlSzzohND/whdFIrk7qk8qGzWtNqx
C31WDLWnEcTYNwRJ30329+CkbFCVw9tBGAMdrZVJdWbJo11JvSHyIOCjja2U27LYvQQLtfXp8hO5
ArAXMJMO7LlgbkgO+JMfrdj65hZsc6Dst642TP2dQ6m9tyHI+xxC4o5s4a7MoH6UgaCC5Uxe7ca8
dVe7SjukMrTZGEeweBoNyExmIM3tve0NT3U2XQXZa56mbDSbpRX03+0ACAIOanY06P3SXaB5qB5b
LWR+Zv5cMpIlG8+O6Pxo2ZtQECdtvyIhI2NFTytZ4ewzRKinATyXbDnsT5FAPv1xd+iw1DiHeIZh
PBRfrjDoEHdaRlA4RMq6nrg8dhvozXnLgyIskeDHU0lI6NjXRcnHT9GXtVpycrKZFtcw1P3yoeyg
GJy+NbwUwZQeULiGPPO5DR+w+Vh2ZHmdJT2KC++tJPwBeZ77wH8MT07TBXoXI14r/Iht2WCR6HNg
UXx6M2qVQV1jeKx5pVEkASZi99N1LH0o/XufzdC3ztwT3ZQ6AL8sJ+h/TeXm4/dHqGt/ozdqQUJx
AUQPXwKr/ykpbmQ75N/D4gv6mNUbD6kwHoLLA23rWy2ihPWaQxXSEmRD/HasIhT+M5mj8QvPf/aI
7mkgqN4iHeBhykYpe9X0V0UmPTCrEItFQYjqyzy3CvV9dGapGfxz8aosWl1Br0yhlj03CEmUiLA/
vcgqpuz8Iq0Ud7X6OIfGXLfUwtrfCYRHgg39fqpd3tKCi0kv2/E7ifN2I1ueQou1f/iDFZAj28FW
50fEB4L2GFaGluam2DE+Z2dLuy8scFaKnCTE9ajPq7eoBFIdgVYAkMJA32rkCUkFV/oCMlARRTYE
JRX4JwYKLm8CyPvPQZT+UxqaEknHoO3niydW+najqA3HmWSws2huiZWLNeNmorQBdDxBqyosBYV+
/QLt+ChyRPkoZyi2qz4rPFDb7TDCi36DzDaRQAWWNCL0/gJPd20UQuU2jEBqZUgseLGieDsH8btJ
0sYKyeWrdiFgZCp4j6nnY2EtGhKh3kdKzXkqCoZaU3aF7t8RL3jlP6cibyIbspB+pmsmR4PXDULu
m7RWhvdSZgSKkPWNl9DSlIHp2EzLWQ8IBc/c5SkK0YBXtHvU1xdXVFRQ9MoZWpSH7DLu3kBCvFUi
eIVjdlijeFgqgpIZ7ij/WQhvvaSgqfzvoxZYN48cMp183CFw799z5j5aC9LgUqL5ieRA5mXrjiDE
kbWDssivNi9Ifd6YhxMnIMDVMuzNSDN33LfTYPcR1nw3bVMD9hiavC9p4ey5IhVxrrYf2A2UVO29
v9bT6K/0U36KbuYX/fx3pIZtLym0iX7XNCMDs7lwW6ZhjIgUrkGOxAHNU2vP98BTsSo0gHAxGABd
Zh34s21FRy+qQPpYqp9kbWVxae/09L91MUp11atmbr8fvw+W5YR2i47E7hsz+pfp0zgP92ubYxrW
Md+gAnDh1/TdxKdvyctQDhOVODMGpakYXjmcyhKVMqhF9PdOTFoMOp6ltUxqL7HHqCKO7HsBGTuJ
Z6lpn03V4b+NJYM81+ls0DsxSEooLJHCWjYjcOBdNQl0ROPxBllCfr+ki/3qVxyAYwh73PDlW24w
iijXB01kv/m2fum+M90OvCAnOMA0xrHl0S6Uf/IFLVfogwBTKOK6MMvMRKSgE/fNi7Xc6cgm/tco
uVsYommDTlqR0qUFYCdO12TDA6BSZu7xOBA3NUO3QBy1d2NAbxVuaiXZ8dQ5A4e/K9ATgz7v1bwU
R9Q7qCmL66AfrC65BewRKuM8GxMvzsygHlCEPBWYgTsgY1Tw1im7YMSkEAnOFYkSYjD1JS00NJcb
Tyyx5hWt8jCfPhza8t/Utc5eNw7GvdqxIldbvPCPy7Joi3nop+KYkZbk5SxUxXzFxcNa5vL+Fco1
+AOTyv5IlhkndxEoNON7WXa1E3VfgigN69xvc8TaF4IRYasX9AsLWyZpt3RYhs+KGgftiQjSOUhX
pErpm+Oip28+qp++Jfb9WhiC0Pj8O+4mr0Vn8YPgdRdT+c4HHivAYFKQ3/DjSXdjVsoviHqUJ8OL
40wglHKupHE/XoDitx+lwDJHmrsjGlh5KHnTYnpLPqR5kakjr6pPjRnWWdMs4u5ukcjUua/p+mF2
oxT990jRP5HeWo5TE5eg1FDffpCZnp1pImqqKm39LNM8TJzsuth5wpCSgICE8Jo/ksUMpqLLI1ho
duywJIgKwt+yORIiOj4PekMzCcEwFU8neTTIPHUu8TolLOtx53GL3mxYsmF2BEGRVHaxZ9RPiplu
GAcdIaIrooMa68uI+GT31F4O0ya9cDG3SeCI/arCYbPSSweDCh2UsQYs76h8F3Mym/+wF3zepBts
U3YDApf2qdGkGcpFeHFsoJZjkRJ/rl4DItXwbodqQvLSeVYJ+noCiJKlk9THNdwXFlJhbqGpzSBb
RpDzCDVHkEqG0GT3SPyktMeN9PQjO5ditcuevhIHd07BBm4HirwZ22fWy8aw16qF11vHo8uRzawC
58/I3ouYDIYr/KG36hoQB1fwbtD/15g0I+A2mR9bA9Ibowhc7apaGlDOLPcJYJmlGGeiwvV1vXZA
fv+7HHonr78C+vWuCUAIb0RVH4jP49C5WXpQY4qa/gD67dLDl/+suQLYWBrolb5ad1qjXblLB2+r
KOmTmU/NyVcip4/c6A4QtLr/ntHeBRy5xE0plfb404uCH3RtMt32paM7PfE4EEIXcHkDXgl8wGCh
84rhF+A8KHHdqu77rJU/SU3DlRki1vL5PxXzTZ07qrK2yTpiUPpCi4HVRuHaVll9PIYT+FO+k9Si
RntOm42JgM4KHBy+CegsAA10lwFIiZ//Gz0jaYh9IWwEOuf/VfRI9Q0JWOIL6DV41XtyaGG6khF+
pK9A74AwfiLCaVtBYLAGMrSfxN0y4s98QvatJOG0ZQutzJKfDbdZ+QFvrUDmPprbDuh8o4VGllzc
iJcQKEEEupj1U/5s8gXksTfC5EygxUzhP/IU18GSF/DJhUJMEtLlt24XT6GLPDMgkSDOMk9YPeHC
69xKnfSL8yitCm9isK+t1XgnW+92b7orsfWp6nJmIHQClTrMJbiOQA4iB0f+si2rS+KjXAe5PGyG
4riX0XbHTG6Pxu1eqwiRhAV/LkJkdiDxUgUtLCo9c8y+08tDhan9jnjTToyMpjXjGt7k3XR/wi4S
j9F/46xD2M+LtrLU/IsuU9xoc65VcaWsxjloZaMScYME7ArcA2eUzxA50OhYk2zXvidvigU02UAp
CZdyOlbnYrYi2s5N3N8gOKk6CSQtenbD6tP5t47BqdSeaUmgC2BvPSVInSFKVDEFFE0MBDOMvDqI
Qg/elP5YmO9tvCoTfAlWM35QZaG4vdwekZiZIH9DKFQ6I2quTnyst6eqPP9YGR99jMWAZttwnB3v
74JXniCWmZc5PIMxVLORzPZZgd29cAx48WNde4fhWgUBktOtkk6crJqB8wqQKsuh97ruwNpeHEyB
jD8LHwPSNAVFHMWPJUYxiwgHBsC3y593XHtvHrtG014K3DI3R+CWdpWRs01+tNfkxncIos/W+cUI
HEJhVYEaiZku3TnSNmYk01g6kONc3QCdi1TxYzCmNTDg8ApQOHmp031IFSga/BYefkT0DEEuZsfa
2XCb9Xi0MyRAGhkQe/MscDRUSL7II9pTb0hMkHLb1yL5GRvt8S4TyBroOcEO/U0PLq1f61v+XcPU
/oTSOf0Y4ivxWV1FbZIK/5prX4MhaonkDDjvwOCiKYnGsQDvRPSeRyPgTHoZbfWlgg//bJhoZUzF
29Wt4KoqEvS62Z6zQtepkHJ1rfir5XbwKwjVJF2Rd15W6AKBPR2daEsQd63JA/8pYZBZOrZ1DqPj
N2VKGn0+2w9lPH00yBZxycloA0LhuBF9BeCqh9SWydIPrvJPmYYoZtnadXT55bXUSSTWmH/vg8bU
FvSH2tKb3WMWdRe0ALtoeJWSvRrWGuqsfUq4LQ7gMXO9AacSkEUPSvOqjYD+3LeeiqpMtBbuHLyC
IA3xj8RzMAKAuwpn4+M1MfaSdPfOgEs/M/RLS5lbOFF6QWPmo6040hY01RxPzchdA2RKgGYAVjxz
24L5YK7adYy1Aj9q2587TQNJVuo8aYH5kCLF4inWhSISsn+kddrAngl6rttWS4Hn1Vcbdl5RCri3
5gKQlBvRD7fNccwnHE8wQm8gpvFlqb5tThrtNW4bLOS4Vo8WpFjV/6lEwoZu2FaOKaVfwyDpoAqN
9HzNu/owYjQnPG5FKA18gX0CijSAaQtKGZYxmmdRObj63XlofzkpGNsXYYbteh16Jdmy7JE1s882
Sd8n2Pc1aNNuryngdnTLKmmW4VRimGSnaTf9Uo6cnXf+kgSJ184SOwZ3p6AIe3HUCEoPl7H5qU37
8+es4CKhidMa7IQ+uFHuP9X5ooa/J1yOZWEzlQXaQ/NaEOazBY9o0j5NvjGSKu2eLDtH/jHCQ2XZ
U8pOzQRtjC0EnoNiUM0FGt3oqCzHcZZmMVZIKLVIankn4C4li10S1UaGxdhjRWBsCizeuF1OB6kr
Dp0gk6LYeiKT/98iZO7d+VrM7TDaubw3HdHd/mO+7+WslYxvfcM5+okSdgmFPDu6yLrIrpbBPk+1
X9l60/MIo35gR6RopcHL0sTSZpohe9gHaRsDeK1y7dgkSLIEG5VlEgnP6FwK6mggiSthJ1OALUAI
b38je4gYQEGzMG3xzv+tmurHRKPVDMiffd0Uupgi+rRmJHAkxR/lr10JVupojrL4UgpWeKmUNqJe
VTngpnChZRKBPxtrLUSj/1t9QRZfsb0a8MND4u5p4VRlxS7MeD/926zq4/NrWnnflhreVNeg3FXi
zUvBU+O/CHTiuQ56ikScjk6BndUCsw+d6QM5hIfWbUgryxBiOoKIguoZHX1rAqbBfL4TarIz15ny
6SGzu7VxIqTFDRNdq00gEq7ksbAdue3nCyaszxwGaubaT6aBeJA+IC4nr4v46kaLkPr//9FXlgUv
+DiYr/GLdpqwIGzaPxx1eS4N31vc/4c3W0l0N3tg0h4M1iNBF4qadN1Es3YIgK4oMxST7gBMPQ7h
V73q+qvO670LlQupZ2j8zanASlApCsBLx1bjHE0IBtGJhCxNDgdkmKlGVFmAiVmHo2l3dW6o2s+d
ktyqpabcc8W/S0D+2Sdx+sY/KR+6veeNEeOz+kGjDIhRcH/xchA2KzhGjwOixge5CyyPwGjhNPql
XqVqFYOIO+cjYD4EEAH0N5EXGz74FowWhRG9Y7Dw7dU7Apf1CPwWthG73X6tfPxQnw2HCbmGSwPw
akVxYjg5lSIGRb7F0RiIc4EI2KKn1734A5xC1oRUpYIo1LaPLRG+KS8YleSVSoiPSD5h/BOMxhAl
cr72UCokiq17EoImLq4MDAVuhxQALp7uSp10Q3T7q7mxzQGl+Fss9Bqj+3JAq5fMWkLdhG+MvFWD
5J8KREdSq4dxCohj7+iLfoGHRQjVcv0Mmc8gWu4rK9f8o5UC7qWNpOFLmUTdrOf90+xeKdeegKE6
R4g/+6HRYmCz9vpWX+gzy9SUIfeDhpQggYUea2vvyNxVhjvdDECyFRn+I8b7KHrUdVQQDkCxcWs7
dL9DE6jbG6y6RFU4ACqvUTDRHDps52UnXoJgbP63Zym0jFgt9wRTZZHKC+Wq7skXDezyAAFOgjRv
MPaqFa82ekCL/v1ip+x4bJc7gmXwrtk2rjgG8DEgJhYtUITfwgwGvuYqawgUX/uOo8lOhkH80sRl
oFQ2AE4xBcqpUU47uluNn2nirnPgk0E+0Yz/j/5KYQh4R8TpWP0o+xGDq/fQ0EDhoFUbBLoVNCXv
AoCHVgjCZzADNuJp2/xiFOLiLmTdLW0Wmd6I58HnzWtA4KntvlbRww/bVVZoAnMfPc+wA8zaiz6F
gVJLbgi+NS8Focbx6LDUjd9rUMQDDLQuxDizRTY82dZP015aOjVVR5XHE9L0aO/VTAMsRshhkX98
zJufqDbLmU1L10SFI4M9gOmO1VdPa15JPK4kJ5qX1qCjlVE6tKq/aEk+raVhjW1wFYD1oWFwFp+0
I8exAZPwx3U5yE5AGix95QLW1xCeQb/0A0MqWE3ZDnEgHgiwewwpIVsmVOiCCBlAWyAYCRUgX9Tt
Bbq8IBOMeNfVcfrBB48jJJCKUqEdUUW37wM66uc28zV/rMqAcQNwj7x70F7WQgtUYxFF7R2PMmfc
oP4nxJtBLeo85rq65b+lPnPBCIodLj2t3eh7VR/wccn2oXofn0tRzjNpgOpBUeUR9Nt8oxjZUGvm
NKauFLOgejDfDbXeWFNV69olhp3dxKQLDyfnw52/fkLl5Ts6cczM901HK98cyjYodp+Thw+1DG6m
3Rd8HfsQ9B9/08s7AzpNavUAhIWqglHjTINrgtMRbHnJbq1xSV/avYHOEXT35gW70m4sCNvl2YBT
IOPE20nJX0x8lK8ZBpsORMUSPKidHJo0YDfq/aYWtuBrxW4rOlk1BqrXJca5YYzeOJhTaEzdo7Eo
+cK7MSVRyqzm5zM8R0weeq+Vjt2+5Wd+vvEM9E8Oehk5GkBUtqpNt4POEygjqzIRbQ+bqVDeEQ3n
BC8M6NNUjBtt+enAI65Ttt5XOuVio0PVuQz8/6wQ/+5DDDwx3GCYz5Z0C/iHO2OaONhx5EQMTdwi
XvvkfaXL9aqccn7sz0O8sECwfQWInXxFU48R00iDaRMxk4t+v9cwTAhMiduKhWpNfNql4JVaVsYb
ajdcjeUA031K2mnKaCyOlL5eaG4UqjLmdD7ybcpepF56xGdsVWGO3Koj0kFeWKRz/LN9tEsVzjLC
qtDI8pjolqURM2loZA/lCmGOL70H2hpAVbKhluBe8KeWy7Vl5c4dFL21+Cnh2+eli7mBQevlQg90
vaxgtBwRYS2H1NwZfdLgt9KLeezguBTq6jNIRzynB44NfRgAEGNJxu6WUkOiNBkFpKoftMtybtXk
k/1sG0X0L+X50Bu9bUxCXLlUvzOVkiGikqOQ3NPZMYnR4qf+wusHlw727zO4cscP42hwxjKdsIWF
0rp59WC5R7pOt8Xx3u4Plr9Jn96IQJ2C6Btti3HJZ+askWjtGQePOAnKfB7nGY/1aMNOZWXN77IM
5E1LxZlwxPkDQgWfWPklTXnfp3HfFG0qiKDHtnVE9cQhuuwL4uCkXo2VXL+48ARzImSrgMp8Z8DE
xtj8zHWTCItFUIvKsuRUiRe7ClTP+HaDEaB2MUnjRqD+wTmIl9SHsA9fBE1rbawQVIHdUSWRNe/0
gC/RRnJ3hPt/JpNHyWd2HfhzeUMX5rxxs/Sg0IEL2AHtU22RYFIBJO0hv5GTUxafccN/EaDgj5Go
WCaMOENU06DxglSzz8qe4fIGXaNTwTJH8lG0UvpyDGvHua/2mk0sT9NJNmppXcuCxahXmLLlckoi
LsO6wq5sY296JI1scLvF7yTarY8SHQIfnHpHnBD4OSJqPjA0Caw0Anof3dZalrWsf7Z+YpiQmGxl
0ZvMba0UlQDzqhCfCYs/oRfyHHcZSxl0tnhcBvNjQsJ/tXTGeA3ykkqvDQ5Funfff2BBNP+h3nLr
s/Flpfrw71vvBEHlYzSLqJmallUttqjZz8x4ojcWmWCgt1+GcIzESUi3kVI7fV7lq+TTsIgNmqSd
2Id++4o8Lxi6gAkQLzw4OVBd+yI4dADbWsj9kkJNjP1fnKsNOxpegdOtoNsFi8uMQt6ujdE8OKK0
8e0dy1sQ2aylreaU/DuMcxOs2v+pnRXPbeWVWF786EJMrE8BQ/gydgAMUQ1EhERSp5AgXbCJyIzM
7ywumFw/ar0OypBjeWMwHFl2/XS1U5Jc7hlfoHvphEog54gWacUPspRqZWqisE5MpUKdGL1edTBb
at4AYW7yjKNKcjL1lzcfC3eXp5nsArcAccngNC5sYED2JSih2YJhUj4w6FPKqRqy1juMO4QOwK9t
iDqMxSB95dc1MSX6XMkCiaqVhCMPmQN/W5XDgFLlb3oSFf7erWgA8GK7hqFcC25G5x+y0qA5Ca6r
1GOVbjUcuALjWgxtYdpumyFqVeD0XGLsD2J3wkASmEzIW8XKsgyR9HS3W9E01aua+UsU3keVvCM6
jGMlj+nJR3V1Qe9OzQ53ZG8arrGWB1rdLrdpb6c0zz+k1Gyv4BWmjqYDVp/rXR6sqe7YSvTU8UFg
VXlUPrpH0Kd2pXyoBQhO7Ew2B62TZdVpJDMbNEzz5mWBUelf3ygaHso1S870pwaYjjDGR4aVyWUU
rzgFxOUrs5zpvzBqCZx2UvPtQNqOaT2doNy057VjJ74aYorUtLoZMHZh+8bCdM0yDTcP1ece4kVI
X63mxssd6xb94abFeKoIU+4PEcJWjE2ATfwPQx5ix67bzM+fKR0A4JfuG/qO9Zd04NHnHEDFjqPk
QJyH+EkuVWqye/PRSYKiDwgCaONXA9n6RlvDCgDA/9yhG0bVGA3/oiaeRt9eK1AaaRFARDtA4SSm
DVAk+Z4GQkrZSorRLIsBCDLJYQF9ikcYHJMg11OYkbfAzXXjJ18efGLfwq2akI4htp7XsfebNd8e
SBu1SoHqPdZB6rNiHHJpofY3rAYXuZQofVU/zX4P+vZOrW50QEZTIo146wdT6THVnN1ehUNo39T9
Y4em+6RUNIoTeumQ4rzNuTmE+fVfv5r/9+Zg+71MSvPrYKPazzvMYBWZlS7qxNz2GdEexLwIdE8U
NwFqfSXYSNuVPURLzMqCdt0agtkH/csLA0jiqx2LYrVUITknrGmr60n9aloNBfepnoVC2s3jfvGM
2lrQNjeoOApVrK86BKOolyB92vc9oKv6Yn9n165ifX43TnMrQVHlEqkF0T02X445z2Pf7qR9dbsh
fPc7pJ1NfZaLlmBHSLRiJ1W0G3Bo/BtGlx95e59Um6c3ow//U/f3oWBrVSZ0QC4TMB2k0ddqWfRA
vohVP4jWxjTbaTB7viIMEI2neuHpOABLmPlYauFQWrlEa0pcSYKTlbx5mtixLuYhwRO/O+DjwMNA
8K8xQbe3nbwSsmk5lJWmZhdWMYnepAXQMh+ecEQ2guLvQb58RreZdAiNNsz+Nc+4Wr6GBQYosDc+
xzKggPj418DrDkHX4yziocMlS9D7D/9ZpOMlhfa4HtLpcD4LxUMTya/+uYcm5+zmIDitii7u6/vw
MM3QaTmbAGEd9hpdcTr/RT3h7+YkYF5V0WzDIdpRlwL/vCRVKbVIvBBoZgBNb0myVpA6A6ADr0yu
G+vMhT5fhgSOi5VhBzJNekD3EtOUOXSdocIabQi+B+h0kpvXlHB9PuUVM1+VEUjloZSriT639mm9
9Q/pTqRIEEnTdoSSsTY39bh6R6u9PqbUJFbZ3h3jKtWFOiJSyfghKo/uNQ+Ov+CGPvu4dU0Iz6zG
wc3jZu+xSAkc3ojQoezQ8q/dFFF2NCpg5VmF/kGXENje7fTfxvH40mdWmgQL9m+0WUyfWr7cZW3t
AOD5lZjPlRVZ3F1thpvYtuNkLQkUQgbWUqIRv3kZu1eddmzg8Xz9NLrW8mDPca816P4JJDijYNfg
DoKzT6G7R0vC9zmOtYoMeOpUno9IWINzDOAJ4LgRhuRoLEJsk5hldEB1yRibjAEJ/HJQAgZsPS11
QJeavgyb0lGVzTaaeD1MrRVxzdE0llhVUdaA04ykPzCj2p2bAHjGNCpCOyuPBvUd0rl6w1oXhTlL
PZR2F6sQ0Zn4lRj3+1LOZcaULSFaTctXx9WBpCJwW9NmXFPiDK9TwF/bD1U8IE0KshXfocHDfHrd
xQVMWRH+3rrrgtapE/QJ0oZQELp6fPnryxoq1sZ/CWQe6XQGb4BHqHm5p6g90MW4M2WZJHjYppk8
Di0MGHWFwEGi/5h3n1piIqV/ArXTyIFpTIYmVm1r6SP2AdAesVRMGxz3m+fKMpmVd1qF5Lbn4+uW
EJ5kXsBQoDHNegqzEXKrdFGDyDUzpvLuwZR455dQuKooE+sYojar/cVMuMAshgFRP7fHi9jg4BzI
jbzTZ0VYxJkYJeoQh+rlpyrOpy+A9iGmrYaXhhR54g8UFsMmabxCxA3RJM7jS1ULuiudZK02ahdI
WkbCzEGenUGLn+0i3WVxKGOjlX6zkA5KcmUkkMUABqt0tuRiefPRMJAPm1LTfY5xViSqtNIG1MXq
qavQNRKm6ARSyXZ4a0JMd7tSr8lihHLiTm/5DPoeTbsTFrLRxM6SWIq19RiMjrgSqIGvsjqedhlx
B56xqXv+vCpvD633D0xl5WgwPWr7MkAljaTPGj7P9prbF0vnXZEQlnAzWKtdrs26tEQBmjRodYkP
bGZ62vOXI3dnsD1vezWd3saAUp7OjKXBL/L5EKQgrG2B9l33+N+UvOa5Olr0Ffk90g/a1c1QFVKK
48IyYb/+qQLReT5Scy9GHIuA7R1dbmek+Qn5B8GXo27fxKWK1sM8HTiD8RvmE91ATWW/2UOut3k9
X4jpLRoja3Lp795mRvyJ0DRJkW6pl5GsA5LtUlLc6IpHiO3ouf9HNw0hh4lUME3JxH991U12MYL0
HTn8fgnz4EZwmGYzEtMtd2Du8Zmk/tN9ucBHEQyqAWcm0PHzIm4oGcNz4fV3PBkFkE0qyERNOgdS
wencDqVvxFtSY6t/sbUMMenV5STq5wLnMv+ENPReBPvRcX8mFEaLbzC5kR3W8HxB2sHU5bAuRNDc
D6Mntscc4NF7Stsx/9wUxU+bo+m1EztwbfZtvfaZeRG1KMuNMOnmvQn1QqzuFZiCG65ihHUqrEPU
7/XrjDyP+ZHVbcRrIrfQCe9YB8cd/s+GkUYafuU3ce4BjnwyGFqig3erW86bSIcziZ2UVPppZ35+
i9b5UlhzSuvWZDitJlLB8AwXw47S5bVY8knAzmaZo0gSOhlIK7BnRMrYdGTpmJyiJ/IlUXaiebvj
Q16e4/MLm2i5Edj/VVeFAP3nsGCuhlBGzNTCclR3kafifLrSk0ujnmnIjRjVXTJS0eFuXeKq2iWI
7SGxLmqLByRerpMD1SJbdQ4D1Ug23Ao1Km7zktfKVpZ4IgidxCTrWu7GIZhpZiwVn6GZ/Xs9sdij
2U2wAqYx46qqhMU6NCjVb8lK1dDHJ3BjPoQ9Lj5WshGrWNDx5zMk+8amncwaNrvniiTEENEflaGT
zZIQY5h8fC8FCjwc8hpLYtaMGWYN1jcXiclco1r9Nbr0rOztXUgcPaXBMuRL+gK4MwUr7QwhHtNI
NbHH2oVj7IEwuKAhVOLuyu4bagIIZ91BKUr6XaMHVAKkxiHEnHJSYAYbYoBLNzInM+Cokys/qYk2
COBE9sPez7ViX5hiGvg/Nzn+kcAmKxFmOp47yaxuCpAV6C3HkYFjymgDdo3d+olggrzjoZVJG+8q
99CdyqcXVszT+VcCy5chRnm0ZWZPLQ0o49XXgGBZYXJafmsmPLFshjgCy00sSS2+xnB5EkfmGyAi
uBzsy56UBAJNkmHa0gYuny3FbQHl5pU7BytQN6CSSV7SP/AHGeczyfye/WEYgLzx1ueC/cK448oa
LGuKnK4h7KzeYkDlRDAop4O+YsvME/SpMnI+X75rXrPP6J+IaO2kdoK0VxPn0k8UeN2NWvEFuDqH
a+vcs+r8vbdBRNPDHWJ6X81S+mB3Y/XCyZbmsA4z1weo40ajP1I+MnVwDn/xLdhaq3h3QFQkyaOK
L/9ujZOzCf/YQt52hOzL+3SJBI0pFc4l7+jCuMJi3NaAy3AG3WIWBpczkHCSl4cWjbxpWTbJPfLh
eh4SxfrWUYDs/KOD5C5TWGJXIxGgb487hIkw9DxT/JZ9rbGMmJw3ZfuPqZP6x7EwN7MQ9/ccH5tO
aJ+s6Bai7E4VU3mEpdKOjsSygk3bsnmDPSzQ2M1oNNmOLDPwwEIqGp8g5hL1D59UA5tDaRRxLEwQ
o9l7H+XIeIzw5FdxPz/1nKN2EBWl5hkAq4uz9KCpA/oWmzCESgdG7lMbAd74ORa05DwUIeJdeqtd
ehDOzVfwdiirr3TSSI4c0c/wLRFTdjIs0aDfBk8mxvrBiehIiPQUsezpEz8llXqATfT8E1SvWm2B
LgebvFrf1bDPEeK280OTBiLR7VTdPiY7qgGHIFLhjgrGPuuoaKnpqLBeiXRcP96qowA62lSn52Sh
nsz9cC/Ru9xLgExIxgon5gPP89okrfA+tlkG+XAKX7ppT9+sOed6T8xdkF9jZYgWO3dlyGfv4KAD
5ZrqAUJSWX5UNuMO4UaP+8Vi680DuGdNQK36HFNOI2FePQNFoRaNuVGGe0s/l13OJQrfHZoYkvy/
3sR+mTU8e9GKk33AC58aiiNKMFka02Uc9fhUGAb0261/iuXXkyhpoOuafOyg5BxV2uCggdY3rP9M
zJuf+XgIdaBGG095mx6h6UzpyZpAlu2wXZus0RiltE0KukAgdqC1ySZFnKnNEe59azFqY8QUqslz
b7Y6YPQ/Z+rgGXff27wVSCvwTurMTZ9EFIbnqWkf3kHvzEjXsz8KnJWd71hWNoUYHV2LRdJRbKh7
bFzgDtaOVLWvc0RXRNGAHnKIozd8iH1fAGcmW8Asav4Ll79LZzb8HAWIbT3Pz4fgXzftriqZO5NV
VFO8FoX5E5BTG9Co5PHMi0hTNlvWc3uwVZn9nlwd9S29rYys0sbJ9jzJaX1jfPGhrZCJwvNy8Dz5
eyfFoTeEHeZrlEb5zsGehcyj6Ug2tFEuv0VBnASDjj7uT/S2UgMDsSAHpO5WxjADoL771VBTkxwj
SaZ6GeUHKzqKZ0+k59fBlH66xuris6WwqjBxG7JXceDfurVjf0t6oRdUHgsRlJK2JakfGxBs/35A
4s2fNLv9X1aFcAL1T1qdYHmD2riETIkZuGACAlhm/2hxqgRdCb341mkltptNyLtWDpdOXjfCeE2x
2e0cRivWVEB/S1YZ+lR9CA1dpGDRJHU6T11uYaQ53ZMGyvuYvovytpbcWFduML9s5nRtmpBvBSiY
1ASI+C3LhG8qTHWNt96llRCb82tc7sQW7PXpOTfM7qc50LMnnuMoyB2nhcxXkHA/qlK/iXesFJcF
qH9TG4uYv2YxMY2e7Mn0//F+/pDyrFUH4wQivA23N/NtFZAZnNPCpnWIIrO+QiOfIV2hprUoQbVu
8guwua8vf9ZROAoN78imVXIVq5uBWogJEHmrCTkD5ZxLlwgXWBQQUYYt9rTbD3Cf8Ll7pMbluoHE
mH3bFYO0pHTOgt848ffXzA+AjAFIkHvMKdj9uz99E8xyWGNc2mByskn6J4XbHOL5HJqSA/csgk9x
fuQGBRmS8zC+LsoqpuTYts50MaVOF9/jhJ6OzRNQ3tEBqFVYd4CAuLi6n12UJxOZ6lFwd4yfHNn/
k/x5+G47wZAwyCBFvQJZRbdAsPJVc1byRLIC6XUgd7BXCoWlT8W/aoIqzFnRlkhs66EARHnURi59
2aIwNDeFefhPIrbSeDrezlA8HPGQOHDXWZcDwOJJlY9i4dtby0eot3jDMjM/9L5nseQfiqFbF5kM
2LHvKE6x3BSXVwptV+hgmyVYjCcfe59wiZrBF+wE+cWXcUzIJsSAq7WG3rL9IvxXa0aHQYSLm0C+
VVZr3cInAqfNpZR9NtmMy/ykn7P6ihgwHn+h1pTzClU+zKY4BrXIrJ+K43Zvw7hFWJx9VsJQxeC1
P4NHiqJWnw+Ef/PLbpVuL49VSD6o3W8MHyHntbmbbZ8pyAKgzUSlH5WHSDqIrlMZ1wws3avYgubi
RPyzTmQk6j9whfInMYOF9LW2x45gQ+gu7HWT1kB0/4DHHmzyRnWxM0KTqd8fYM+CdoZWykJwXC95
DzcXrEmCyeGzAIiRmuEEYlsMTWT8523agGLUNaBW+qCRvOQ4B1KpTmLs11WHDrWy1cTzpTeFZvQI
9pz039Fl1PBX+CAbjO0xb28Aj/oQePNK3o3xbiHAdOR9XsTlhWPCAEXuQDZZsgqv4qPihPx/JM4W
vxbGl++WvUl3FW6aidFZk0qeks8huqSf/RxtgYtqb8airbmCPXa2no1oMdDvDG1NJhQa1mQT04m/
YYHnbt6vuH/UdLWVwFABb4ckfUPv2dsJgfxQUQc6Z2MDT0xoIj4b7dYGg58rn2MqIIFunVKDhswi
BOrZVtZbdPS+ttOhA4Um+60HUcBUCaeFP4Y5T9n44EgTZutP9s+Pu6neH1vWMcbpS5dR7ohjiVv7
7LdMqiyzyxG6Lj8X2HUAXea/u1GZBX2sLE49noYluiETj5XshOMUNVgIntUk9Y0frzqOx1BT6Xuy
RU8AR5np8NY8Zcuoy77gcgEilAv5Tguy3VMIyUgQ1F3Z9NQaWeDUEaq+znopz+XWXxfn9xjvWq6n
JHZHWn/CJlNQt9lJQI0TTR2DoadWh1HAMLex1yluRCn2BNY1/20IubFiBbxJsb+v9mdpCSlwcSzz
XsagvxzUKzDqKzH0tzKvPkDEQXRVDF8OD3m6ZcwZBxFqdaO3colHENR94yceTYE38svGa4vKvv4A
j7dLG7SYBvtWK9mnGSNaOXRFcEL7vauWsnNPapBdkWnPmSg7f7h+YNsNDLlY4f7IgODsczJrer3B
27jZsnGMRoQnebIoBZQVfeIfgbkCS6pvLBYT66xIVa9DESwBXgr/CjLAkBJ3KBx6PxNcHGFhmQdp
vREF7bUIRZtyRRgtGfm705lzDVL48aMCQtYXFVaMZgItLWBO1zegCrMp7MOdE+RyzC4Vym5nI8Bh
aFBPP6EIJxisFJJ+QJ/KfsvyzORMnv38M9AizcE9wsHfbGC0X0ZMV9ElM2ID+6Z1SvxKXI6XA7tC
qPHy5s5/xtqOHSLzC4uQg0WjbqhcpYVkdPuedPprhYZPTUeSsatQSLgig+bmb37widmI+3bR6flp
g4dlqyEtb18Y5e12aeHrzwlZdAyvqRvmsEr96SPubzHCaWyUU9h/hbcXlsUU1aPfH3x0f8dn6KG4
rGWWa51zSJA/fDc2nDh3tmgbugs9qOj9jteaZCvrHvZPAc/kzXeSyASPUI/HbA8kSpARQ6TG1clB
keZQSwYmp5PLwrouqMv/5PYk0+hALThQWsz2hxTunSq0O98OslRvX8SZjgg1PQW4pYBap+JMUcw7
QFh5OSOWM7708FWWLVXhFR/iidWJLObxYUopKR5LnSrWYXviAkiam/TYbFcGPbQfrJCSLLc5q594
IjWSwvLEd7EuNcO3fxbROoowsP4iR+r9z+HqD6/BJVSu1o24XK1wEdhmsGVBd1yngtbZ5iAG8cwV
u84gzifouREpMMLQ88Leiaxj8YfjV+DHw8kXV6NXR5CCdvV9SoJ3qg4SVOM6rzHIMPtcLA/dG04h
9obN8kfkwqsgqx1cRvKf6+MOnLyLa3FUddg4ztmuOKMQUF5Q9ux2bnJ1Ycd3Dy1rlPiMOE4/WI8B
W4AqGaMSMp12MDm1lkwlRyK3XHlhsxZgLS3Zgqg/+BD/S+DqOxSc1rm7KXP8NgRsqvGWtTj0s+zc
+IAxGOJMeMd8cQC0C3FruzNZNqxryT1mSMlQ2vjp84xTfp+CF5U2pwJLFKSs03StgORgbqGR8ew8
+AppvefyWJtxKWF+4YxCfnz2VCXiVM+Q1Qq+QxDpF2oov5KVD9405qtfw+Uza0xo470CMTWOYHpL
VpOPXXQrZAtyooicshO1nEcAeLmt+OT7ppb1hwKIfgEJQgdDOxTeUwDuN6G71ffuwFBX7Bmv2EZT
D8MSUFsOAFLQq01ff6SUnv0apprZg8mmSvUCgVlu/peELQHVh/lhTS2MFH5Ed/JPcV2ngavtevLk
9xnDh0uqo//t2zXoZEq2C9W+1/fqxfqSGRUELpqSoUcIXxOTGMk+RXnG3K3NHlZjVXXsQg1jRS4p
DJ9hrAMrkcq3w+5PjlILBqmz1rcdiuWtvkTCTujrVjoHkJ1alZhsbbylq31nmEZBWpCoftb0xTnb
PsSIPZOFfIKCx/h/d2La3jhGlzc7s4QpB3W/HQfb2Zc2MCbXuwAoYfS9/3fLsRnFBEA9YMbtfpb0
ovcOwQ6X8wcqEvYzMfFGJXSuI45nwGtWArp7XK/C+al5wWKGH8dpG6wZAxfPTT6b0CkpkCEE7L7v
p4AF0CEfl6KP917FAUHW0jhqsLvQmgwlqazY3LOIKEP2OiIPy45beHUGcQ9XifLe4tx78f0c5Od1
H3jcD2obNdj4JK5mc/fK20InnnYBdBoVvv4ZfkwWIl5ePbiqccg855Xveaa1PjkP/VoSinj2HAmJ
bsTLlVJu631iWLoXh5frX32OyV6xXBtRHa65PeehbvB1TC9wCtO+a9FkSR9ayv53vcdvp1wzJssI
kj1uawDOXLufWigfHQSzyQvclkpkKejasEW3BIxug4DUwVvRf/f9Ie6/yE3/ApfahDELs2ESeEOq
FSwZ+V5bGIwmY+ZU0T1LGziHox4H+U1fBMikrnJsckI3Ok2d2+sTXYOijeVKF9t5VchbvZBjn9Ys
Rzr2ngo50A76KD9AKUGY5e996kWnAPs0/CUznlezbmYDWyGwe1x+CKqnM10bRLz284je6lKKfg9I
BWAGkCw+xkRqUzGHXZuj4iNnmiWnM1w91Eata641xkN7CQke62oKvLGZmjalSAGHkGqB98buj0fV
YYFrVZ0KnFsIXr4vg5HOrVif26rJ9ag4zldiN4hggX/T9z76mdEeX0/pezwrUPSuR09+AY0uQ57k
1knRbzb4nhuC7rQedhClRicgNmorgU/cAvH5SBaH/ilJ14waa+fQUtp9l6hH/cbwY3W5++UccNfW
l/NYhs+UOMBdnkmDn2DDJOF2CPwk+pFRTHBFLSsS8dKskuVD8S3WBtN9gFCPWTte68x/q4b03ey6
CqgsKe91WCcxfQKjiU6MjukkfbWuLhCpZR+zXxpo+wFTO8SjkLH9xBbRDv3XR0Yt43PvGe4QUzQq
q1/q5AQUZ4JRzaGiZ7dcomTxwH+ZJoosMJEPWA0lec1eJ7d1QJlg9mz2sqJpdYhhrSfZmM2uRg4A
r8djnPwWcV19YQyJHER5YU76pQE2LzwlW0rqdUQvL2uiIYV6i0uvzqSrwW2SF/7FHxHOb2DpHP1y
ClYO7zzWfoYqflgccxnWsoQzHPPaBj6gMOss5vdo8s7N48dl4uv3VQ1pTg6RvaLwI8nWyBXmepVz
Ae9ngNz7cNAw1HTizCV9KGibYFtxcapO+0Qzp2rIpTpUXIEz0jT96XtNhpDddZNnSncH+dGlTW5W
zAXFPKBHjNcWxz6q005ZcTsLEHun/xavWCY3j/mLtkule9AuTue02ShvBS51+1iPXPEZrv4N1dwF
/ipNCPK2T8A8eMXQlJq/epsW5DwGvJXhntugy7vT/Av34owDlH8IRxBExkE9dQ612EboX4zPwHr9
/hweVbeZoB5wIr2CEvJuCChOVbGELyPTHNjVBVCURVK4ukYkdsJMwFdVAcmZuDAUa61iEhCbsBFs
/imdHVaSvxsvkiMrzgnAirLigZqQfmh7GG2haQPoxSb8HgiN0V0ut9BKtEpeMmTgrUV0kd7f09Sc
BnPkTf/xcO+k5ET4HyCLZlqQMm/Tx5T9a1Sd9zasPky9Er1ZS2BirqmTDYqtRnVXO6yRWySYpnc5
eUUlpLCdtgG0G1IwLQU7O6udBRBDD85OAd+sFs6FWdxpkCTXznfsDIuJkgdZBnDhSraeMElVybvy
JU1+OrSwBPtxwfmq456XLh1+Pr021Cy+Nr6Zz9o5QlqhdxdbogLx9SJUjL8mkVXnv2IqW0LJyk1G
WqDXbztHIEI5TfzZ+6XyREHecW4FyFWwHLEWLiXmg9inwAlUaGZBvTRTgnXZz9SjjZ3u0sAa15eq
eLSXxHoSLMCNR/M7OZi6f+0e7ifZ6/XJLHSzWYUZ/tyuTQFcPc6/pKZt5mZgwIybQT4WIFr+bgre
OtoNEc8Q2qB91PP5TP4SoS55X3Ymh9cboyu0qMfd1DPF5MyXAJxniViCaHDns79Bq0C7/IoTDN4O
PkVy79f6Joznd8k7JyiO+w0uDKJ0I24qAYVRJ5x43pEPUOQfk1JoJ/nPgsUGar4qeNM/5A5t21Bl
KGaqe5YBVlAxzSic0BHcR7cDK3n7KIfAC+ns8vHNfJ8Hj+JvDfC8sJKdGCw2pOhm1aD31O2kKnyQ
UDbDpAML8Kn+IWCFIaNuDtGA25X5YBySgEK4hPCpuWAI+Pvn4Y3nqjcDNDinQPY+hVYFJIcLPOSb
uUf2PHyw2/St3u5f77tZmbsx9ysLwq5VYfmx2lO+xN/06mqL0aEY+YEG7uoLLnhK/uMyT64ctDtV
MwOran9cXjO3inPA7FMKoc0SCbdooJiwZvPTG+KP5dZnGOOet7sMQrcMf+nfUKoV+HhQuZ/YL0zM
Iaadh9/f2o4oWLeIswj+N+z12de2XdgXvfvv6iORGKpVB9pptBj4XiPvJQ/z5dPWE1RQW7g8uek6
9ljcaUqiytJlqHL3JtOWb+3wyNlPT0MfT8CVt4f8864YTEHBJ/8f1gPwFwzlP4sD5aWDDEn8Ppo7
LYKuZ0+LZT5Rh/WVyodPZnXh3z5hmyx8OP1ICE/0b48bfoKhba3Lzsm09zwTbf6iqqAsMM1twk9a
kNtb3VbfXp13J7V2PFRkVtOtKbdBXqySEST5hBst47pYjgL0fDB6Oss554U+MJqAksdkz74VNuRB
wiAZpey3FjILEyfbuoSLKFt+gvnDGM+q7iS//vrCScVhB4JMukORVmSpyMSaeAh473aQij8zJ0gM
hl5WGM2VgMXQf8ykTuFbgwyGBp5/j55Ahm6ZPjProsfBoQwLyn/axLfu9hLv2jXI7kjNtbobhs+g
j2mNeNte/+MRkANGkuAbFNTaysyIXU3qx/p3GrCpEhjxQIhzpwmxuDTd/+PJgrMlzPg8iy4IrDBZ
DWYyHx/pHOiJTHcbdjPIcI6Rf1ke+mpz2hRmr8giSoIOGG2ZpuSXpgs04jQoPSHG7nHu7cCR/JUK
PcbG7WZ8IaayFPbJF+qMiRW5sh+IHbPZ77HfJnYvyV13MRuGMXi4YvtMHBrnB4W3Z9rllsOUnoQY
Ass+WNNLDhzhq6W8rKl5cA7IC/5UMDsSkljQ8IsVimrFAw3ISz9eU5eWtFlbrNxP/hJwbn/j7TGa
pfs0HHCf6cWsryDAtu41mb+hQWcfpwXtKM8JAXF2ToLlcZq85Vg0y1vjMLzXyAKkkFnMTG7M5XQU
tPzm4Jj5NmhNmkq+WMqXvWtu9EUBdk7JotLe4mkOH691Xf1p8QjWbEHEAk9gH0r+GSJsJG7MJLXf
MacvsG31R79/Om6japetcjh1WocQsJaBA1+DnBh3R+YozpGkN4FqlYHr5YTz88ZhHRxPrn9xPGqv
ntkp17zefYgPRwqKhlLEuT779f92nGTn5wh9cWLcBvW8sgS6AmRfyAQOyykvs5CChPPXx/I5wH8U
QMoNb4O4tk60b8QbF/NRgIrC5f2ebIOFmneZ9y0SXOHD1Iqqnc+3aZFnaSCgAVPidzJkFiT6ik09
8c95NGqkz2ovf/9Tn+ZJKOsSC+k+l5bIgxzPoqkGryxVTLmlz2Ihbhj1jE+Gle5F67wHH0ltiCx/
Ew+fkt5406LTczkSCWlB4LcFtYcFzvtOqyfXuiFyO9sdQbIxmdZoPKdHOJD3mfFFIZGs/tA9bzNU
CrIRNLXKY1Qudl9po2WpMb+2qtqWAuGfX4vf6KcAJakzXde+sdwutqx9LXg96QGEnG7l92YYoDkz
ZFNK/9/j3azeVwzLd8ew04bd61xqzlxcneLCVhOkbSh820Jyb66MOuGHlqajQ7yRewaw019L8uLJ
2NUo9arx9ypwlOZrHMaUYG0NucpVpuWoX7zmOAv7jrKBUvzGEkB3y3JP5XGG0qU8RXqIMoMU+j58
ASDkNDhZA1+PCKsMe7u7UOrWP7CpNwQqKLBLeBuZ3OsA4gghcYS9Z82xx49DjdfOypYGt0wSjs/b
EOQPOtxd09pfG4dK0OaUzj7G1C3YpTRcC279hGCtj4XTK5tvcikDuTpTomVlIhlJJKAIY9jvTwq0
SVcPlw/iFK5daCSj7aGJjkTQQttuH8UVgs0TYN4VH0Q2fIUId3o5zYeLu5JMRx6XBHCcmwzTtALk
cDwEySkd7PiS2f3/B6b9dx9jn1a32AE28J9oJl7UOQ6j90hfBGuyEYqqN/yVKtNCfVs33Tl3oQN6
KhtrcfajwhjceR1whnp7b+4IsDtkdY0C15FgX9amwWRSykkPd/1HosTxeYSXK4yJzE/SCUAU1/AP
mVTKKwQXtp/u2CW0CJgEtJ6k6EmglL/YCgLupfgmx2nv8h3XVJAfX0sVW09ieQLo8It333csMWsq
5kICQJp/1sFfQcjK3O6fdkTP6U5Xfib9DfyiWAPURJzcRdpHnke62603iMwxjJySBIZyruDqpFZd
f7gdVu3x2isv6IrII2hmGfzgL0YvKiL3OzcWBLw2Fgau2jOUTxwqpcvHs7OlkEUlHVhDBqAN8vuI
MXdGfIufEEPyHkokaWQo/iIU1i+n/qZqQJSpfDEAi35NkYY2kOz6P3ZBvZKm4UIY2QcOwnM2PYIO
EwVStv0APYaN+lHRp9+6F1sv6Kop7wELTHyiR6wVV6BIYjh197ytxZ6SYvT/f6GTbjJ3mvvn052s
XsU4sj4VOjp0TAoIBEU+J/tnBKsWFJRdxD8cnNZLozUNmnurgWS1s8zb6S6/thv91IuGR+nznUb6
dfoB45qsFNxWCobqvJyjqWF2p73yonos5fW1Mp1JjDfFlXJQkO4INltEQcsa5GjenhoPmUCIJBhW
t424k5W8Sm1eLlHxT4vMy60B2pANbuYpzIi8SaBJdPIaxCQzW23F+awhUPJBE6nvqMci6IeHp63b
AZAOkE+anHPFbXm4PdqVSqCBCk0YGnZDsJUqF7h7AT5yRp9yvBXiHmEnhd2uVsb1o94XXYD3CVRx
a4EPqLlH7ndec/zdBGnsS2UILgPjIZu+ZQrAZhfHMTdrVIP73g+RSmFJj4Ya8m/Fy6mbImzo1ROi
aOwPXE1QixSY5msXIel/o+gUevySfQlB98WPE5kJTx+AHDvQjugEfWL52mM7D3V/U3CPWT9BS5p9
OwYZVF64vpBDO0On2wIUWAxo5NDFn0Nf9JFqV9b+RawooU0Pn59ZZqCv5g5RFessRkMG5BN/vWF0
njGcFsfuoUTnXM9GtBSCzncZNPt9oGnaorRR2t3KSqijzIPZR1gHpFMaG5Zncge3YbZ4wIWERJhu
qKC3xYvVhJmW+kWS5NHM4UfAHYrHWls0RH01esRm//Klpyq4lB4unEHSzJnJb29nzsYiv66nIfLQ
g+RJI+koIwYzCJE423wR0dp3kXk2I0rouHQ9FoEKWQFEstckGE5FUGEOduJg8a+U2H5t9s+PE8TQ
NFg/5Jfg/LkYMzhxDwofNEiU/Jm3aULU1lTprr+NZYumjnGYTwRfzdoERW074NerAFM/6VxiCHSV
7nOF2Vz/kCclJ/vML4+2XmiDJx424VgjH0NdZpGQLIVRa2qPiAbv2bXQ2PiTyTpcoeKL/mh+XTzh
/bxi+phgY0GLAMxaJOtgEAKXlxxqG2Qq3rFdaGWC2JR0Jvw1swM88/0+biLI19SLWMf+rnk5vEpQ
37noU0Jz3tVGAWy9Zn4+wOQHlk8Iy+EbkOB/zPK7RfmsXE2KeqamQsA/pCVvudlpBDb5jFNQV3X3
C2KHTy303Deakm9bIVxdimhOGtVB/oz0Yhkkp4uo+i3tkFCnPi63IODWjObkHqSHRarZFWMK5pQN
smzMBUWRibfffObcGKNv1P1hB47KzhzVPR6jP9OmIevwMgYyLD6RlG9or/hoMlmgyBuYRC/Sgp6B
ha7IO5PiFCA3KudHEUAmcOraTF9iMGXDSycv/LEI+Zt0+h9tb4TAJL9HDyKFKkayDN9JuuyRObiz
6rqk3bDZASeTbbH/el9UBna6hmWXrAR0LwhO383YjHKjzQlBy7uXxx6iQevogmnskKhA3dqtXhrN
qXQQLIZBCYx4iHglVRTAVzYTGXolcP3Acq/95h3igQ4guFEacYuVHoX7hEcTv6/axZvfk1d7Cd3g
GqDuEFitJiKY+J1Y/lleF0U+gwdr+n4YCo22ajj3p5fDCZMtQBazbe6K/2mh7VJyEaSsCC/4fr4y
yS+UXmvEB3S1t8XJP/7z1OcycoHjzMXDnNn5+e7VIwkGhJ1zjbDa7uTTW8nFrPTp95dCKN1c8arg
h7TKeIHsb6CJ2f+03R8EY4Q0jDPf0ATWDGPJBVlf4IzvhqPBmP5rOPWWo2Om8rucXd0ZWd1fFcGp
U+OQ/eNtMFJQ6+he/kAv81qGFH4uSAVKN3iWgknqRdNol4P8GMIiipms6eLWK9r2XrPMdVRYUESQ
Q8DQKOhU4xPK1Tq2dPXaYPZ9wxSjqMVDL2Go49HUOQ5WnoYGPI3cdXegQd7vBtXqTV5MyRUxpCVJ
cr/hJHSkZkM23YTqdYWGWtige0n+k0aJrWht1kapXTsdCbqhmq1yZehktxfvX2x4CZIVA5SjSORH
tArJVZv3EaAdzla3YjOc3C63vlXJ/AaH5aUodfNe3QxMdVX5Yfhtn7ETSOayiORPsXcvXRFzREq3
lOex71Qt1SdebpU2NV8nfYMhFJ2yiBATAIJ+CsLtIsMAmunKlIgcc3Li9GYWtHo3wVOnGUSd1gk/
ZMNWV3kd87WiGH8NBhqah/tmbZBWe/40IpSi06c9c/pqBMO+gNg9BjpgwUFsSh8DfJT19mCqGElL
U1HUIZ52nnRnvtOBoOrBgAwdlKAAEAfJgt6Tl/wdzmHJg8w9IjqRZBhNSPntX5pJMhGJ31IRQ4Nd
GwJIFFx26b1IYmu7exJpPTThPrnAvwItjnQq6rmkR8MLKrEWEzZjDeMFZoJR0vEABkowmYlmb7Zd
eEcMrmw4PCBkgOGzctkNyXX2pSMswalORCzRKDmMBRAqOFDky6Tmuzpik7A39XKPasDEVdXbilX+
2Ob3Ekt6BrE3v/ftHcs9KRvoVygtrbfbHX/OSzTd6F6n24JyIohgdMlPwyi7IYpHBJOl3Tb+iZkl
HfBYuQXmqBgoIsoN89leTuMSlrGg+LIKaRScnik6nnygdeEyNHZUNlzsG9i/woCAda0jV3dKG6Dn
UJFqB3p0jGdC9QyvsrZlcCHQg5Ea++F/E9sYOecOhXKpBXjXOMpNHmGOYeQUvQFSqqEMfmmPTW+U
mGSG92sSF0QUaZAminhCMwBGTyV1xzRcaMuhwd8TeUNyzidK1w0B4JIQyu+RA04ehYPyhlhivFJ+
FTXduj1QViMrpp0tD2NFsRIMGqIX0HnwPujS0HFm1ID33VAj/ajPksO5rji/LPrF/ZOcEjpEfXi2
k9CZf0i9oEjveVMsC1ZpfMTNswuVcYE7uuWfuJoZTw2Jx3FBdMdrKOiTd/1WeN0R+pd0T44Ha2ct
CKdACmyytoAc30EqI/0OxM2duTVTek3cG2Ng/h7WZOcBfgqXW5/O5F98Y7FGbPTQ7UxsVPOVP+CD
1R6P8g39TcDSch7ap6aMoOzngZw4V5l591UjmlyNQ9sq7lggjq4K2XMevEcXd/RlD7RSdldCcfex
l7PDt9KJB5ZZoBVwL1YdzYCVLLXNc9rdqk6BO0/uiBgKJRLftUmsJm6nRR2MoG1zzytdikwuK7x7
iqHGH6/vvhLHbHgaol4YIRHiLirVXRfZg2l3N/zZ1fVCAiKDKHU1X9420GEyPqEhTuMWlDZFNBbj
5Lm6g0F4XIjb+LmDpSV4zHWVvPRaOzDbdIG/2nlhSIP7aovqx+L4/bzSzkszD8oqBtEclFpR9Vwt
i5rKBojj4o7YAgCx2UajZhLVVwRmEAXS8QA//mTj25Ey9sGsZPtj9ZilqfDmzhjAwImmE4t6+wxR
HcIwBZg5C28tV8sCtbIOMgd3Yoia/x/XayGRdsXCmQVMdhReNF3xLLLUGIPU6uulpCJQfR296JHd
8aP5CThm0sF6SktrbLv3TBg/8BZBgp0CUAswWA6yRHCDEw1lstIpkAjazTqarT6cktiEZGbq24Aq
AcvjbnTIaIQ0Ww/MJi0TI3dHx9KKXRy2E4kacsNX8GzhXWZU/Ei7/LMIy79mU2fnWNVazoS2lGnj
POwVK2bj3cuK/ehRdEpAAo4i2IwyYrIFI17mZGFsUY6QlnJQWj3WYxKqhSOjt4B6QkliX5TAwP9D
/GCd51VArpEEVY9oY2QcUO18R1kyG0E0WS+VarKFyqjleoUXGjSRIsH42UXbJVFIdgJ2s2Ss7rpk
sJeDsEzRImI2yH6JcZlu1qhJZ+eVcRQCrICRNCMqgij9NbDSCEz5VPYIQG2fhuPTvk/O8VqvYm6G
NqBCqQIW3rbHE1ZsS2glTQoYN36rBYKRjKKj206vYs1hQYBxb/cLJC6E2I9r3NboI7Abxl1CewZE
acinxxFV+Snta86hPgZjY6uogBmIjz7zl5p9+xIwq88lInYURndsBNnjGPqNHC5cE0tehlkLFgv8
AKZH6cjdyxZSbPWcTTI+1xL2NS77MZcxd9eSYZEi5lAUw7bp+7u4RAUSuZmFynsswByxu6j42kvB
dAiKHHI33a37WEnVoJ2CoRyqXquLuoaN81SStRQu+7Rz929+06M6zwedrR0frbTocZQ9rukbJGDP
v7swkqhn4HA6zv8dOxXqun6NNoWUlS1wfvtfeKtSAuBf3x6vHH4pyItivDhG0hINpCurfqySlAOF
TQKX1v1S+01X7bLyISbGlKRItmlbbsJQNq56d+V0rcwB+Wi43JIVUs77uFeWfJmsLOPplvowl0Lx
rMTst4wgOklGwKfizkf5OUrJmGCpa8AhcH5Dw8/0tPgwTPsoqMbEP1Tgyp2hZb91ZLepapGfC/Dr
9nWzizZovNXqBF+lM4CFyqeOd+lXQElmU4xJV7vQzAMhHLvPh9ViQUEYYmIwvxMss+tCtB9f2Bnj
y5crHEmBorvWayT0J7eWNyB/Y3h9x0HnbMbhPjvTcA/8O5FLbeFi6hKK6OIIRJRbxPtVi3PYVVjN
xID63p1+MhLjmmBmXwCzWQ63X8M5pEzP6ktuQwCez0LGNDiIJh+lhNUFT4WjjcJo7N0BVV1JOOXq
v4KM4ZOvZPrHGjcrT8CqWa9GlHYA1grBeee0TFjn8zW37fxmo7DJLm7BFsIWUipCeMBgB9iJElgO
0jQUESe66qe4bSzbHvR8XD+ySlWRcpNPlb7NbbGYPdWMQXenAiIXGH1vZS7jGgNoD1buOvsFb/vD
kF83eF1ksGoyBdUlgNrv1HBW4e4bb3D+voyImLEadJWehc6wPS+4OckeybPRqem9RfuAjZq7zNEZ
5qHM3L+Cd6bUyb0EUN6VJYR75CqSOslpRWgiqkj7Bbo72yZpPz4aUklFwK6Ftj79p7/h7Uia6wBC
ji9D1ymhmy20ZXt4JF6Flj2T/gxSe0nbNj99CiD3kKAqEBek/LvEj/BbUg1jPlv37P/++5BW2Xm1
I6DcwCnq5Kd4KvgmgC0Grly0h9E7XKrhrTpAHBjWB0H+YM/WZINbMBX0OUSTWdCYJVVDTCbbHVz5
ZuQmaHkR7D/FEfZ0VAaf0vtZVcun+4VyXm3apj7rR016VJD+ZElZTXHppaKt8nbM1KTSUpiljpsi
j3P5Vit9Ru7naFNIK+fOoJjpoIpfV7GU806CmqzJ3LaKBPTu2KB7DWZyHuaVZ3XNE2/i9TZE140D
mtYfeh1SpMLbSl54Ft+Fz/OgfbW+anT1ksOEAw3K3drFZobz06Wakdi9GTcv0VEckxG8oLRr9nHk
OrLeEDCbYpsK5+HyBNjfDp4GAfM1o4O4yn3T8MeliDmKH2QVVYLP1mpm8gsf0sRLPbrMtU0+YhQl
yUu6J7RV4spXmmSQtcVFWJV3NxmQCpCL19q/mvguVtZgpPQI8HmB3XAFRADcZMFIwmIWO74nfpiC
50Zo8871fpAgO1GUbOlys6DWi8cX33eNDDqIDfvQVV+rlqk8NhXGCThmVoeZgbi1ATtjw8aHtiZ3
6iBGH5mAGz2F6ioE0KrNg0Or0QDqjIvI3/IrJByd+ISMOG8867uhBeXcv93zcvZZTFqxbuGaoWEW
v2Eo6p1pvBJJwxohQOEv6v/ULo/bgVK6Ejkuoxfd3rbhehjvbToHeuGdg88j2agEQ8fturWtKYsn
fbVJHaSZzzyD8K29sNfFaA63GfHIPM43DSJYbUotyzEBL1B2TW5s6MOFCr2owakI1mjCJl06DDeL
O5dRvnAg2MVqXB0RNH7UzVmdvfz5/fz/8NqN7+S1O+ElHGSRh+A8elEG1weHbBi6VQ1SZkr64cS8
lS7BWKh98c1mvIOYtW371aj89l1AyKAalZxHI1nK4cxJi//Z/V/xb0Qu/59ric6Xuz+JL6HqPR5j
eYLm2jpOVyPJVgb7W0xgzRYKszukkg+vt3wmmsaQbE61wM2+3qwbPoA4dCpqs6Js6LPVHdlXio1w
yHWvl/AqAWS50zufUWr2YKSQ8ns6P7L9zz3N+KpvXnptnUw66aTUmZXBjVnpfgW4t2m78CDjrTHi
iRrvKzSKpii7M5eC4gRqTbtB3fk3nwWkLG00WGfQ5yjYfMXjHS1lnQm36gNvxY1Ps07UgCN6gFO5
GGmGE1ZYnYxf6/Jt0F5xxhMxQEYYilA509lLudUWrc2WxAa+Vt9n6xxxMt2Q/ySZMNNITl0KEKSz
nE1YApr5HHVwlx9bLBDvZ0M/iKmSI8liHsYpLlGFbcgizsRaxgiU2nG4u8DdAJMNyeDbhBfXPgCD
qp3eLCl2JlIJUqdPLSlJiiOFbz8G2+Tc+/y1D9O0hbXLXYqMeIiVT8cblCT8Jo0ChCXlriEEgcqC
RI6TJCA1D4mGkjJ1sb5RyzKQ6140lhSZSV7+R5QU6rVrdD8HFs/8GeFn9mbFT1RsEe30v4DzThKF
C5FOM9P2MPfWXc09ANmvH8BObQhgdmrBnhYpMbOtCC3FVySXYvX0zd0POebLr0rkAtWn1vtx1yji
gTJPfP41hWekOZibh5enVqWIRgo1YTYgnC5kV0z/b40Nqt7lEga/ENK71d+++2G0C433NYQHTyid
4WYQPGLDHFefZeHrOsaZJzuxd+uyxFF+jsd3W596rrWUOvK/CLm5mEYnmyypt1wQOF1X8d2J6PLU
2lFevh2ShFrPf9h7ZiTiOq3i27VtyvEM7c3mg7lovoXcQPPXgLL1CLqzUHP8787R0NecAsH9dYcE
Eec1/2zAi0MdSlglo5K0FTqr8c7gXYsTwHJB5edP21F1dtbNwxBQO4p36NzKqX3IiPIhZ2uAFxrb
y6WcF00vtPeNiFVLyZlHjMa95OuswjZyO/hEYTu+pqNYUUD0vBr+Ps78WgGU7VvUuM52oQmkRliO
YgmRoT8/Qsfud2AkydfX/uyfDLkuhoCPW6sNAS+RXULsFY4143uJ3hnk3rrTlRBNyCUOJ/izwx55
5UqVQVHE3yrsXJD2RaMoiZD6/zYMyJnxM5C/ihpO9TZR/d4P3WQmEcB+E/VN6RYtFL8cKF+n/KK7
Z6pE+hGwbw/gyO23MdiqWPQXzmpLaHbJLmyiUO2S1DHGkPU4UAmI27It22ELWURWpBHLgZyWevKx
mlJGwJuBWWNzAmCqJxCI4lIRxL8sy0+cbLD85wuAexKlzcj8nvCuRc1ILU7fesUBaCdvr1LnaEJL
uO99f4ZniEGpalZss0vkAbfo539MZsqP8FDqs+LLRcJP7m1idSjcxAIo3RM+/v/ETsyxBnQrwf0R
RgwI7iIagF5UYtMmmJMSKkty+jBjE2E+WfeCIesd8RhzXka8qZVUZGerEn1mCztTSWIQr2odHlZk
8DQAJPvZ33inm7g7wfx4S/dBz6i89+NI/ZVzBKtLrmm5j5CF0bNXlnssh4ZbmxDqIJvbdOKjv7gC
6LDkgEVUwXqeUKQDaco8c57/519aDNXVj6Rdi3rnamPSsa+IeFi74IcL3Te7v5PKEfKxUEUA/3gU
LPETg7T44DATzm5NN4hCpCiXQgOtrAUZ5i7kk5nkNCCw+MuKufU5Ni7IFok/WFl75TASsoUlDkhe
zA8O4k3qh4UQhFk2UbEmOQB1p+eHZRQWW33RizxbLwM1umeBU25FOXXG/7oZQ+JTlg8W37PYIRY9
7q4RRAhZ+zBQQeCHdQbGhb819MEalFO1d/OgE7VtorB0+RMWL7nkxz6n49uSjK6/qzjRkHbOolKi
65xl8gXjVzOExN3fj1g0fgAo0/sHU8HtcSXhjdm2o0dQK44T97JGHlf2mS8nUUht8F0yoS3u7TP0
nVyXUxj99qoUWvrSIdeLxObAPNqx9pOKGrlZT6IBjgBYcu5RkfkgPz0Rv+aVdQZd/dejthw6nKko
wdetj+OyUpWUJJjLUPaS3igME7uDMZ6gx/IKjbBQIpLwVR2Jd3B+08HROxKC2Z/3l/IBUJavIyru
dajVb6m50DWtkK9Y0AKvMKA6tCaDEGSAnTM/DlZrt3QQnYs+VD9/awohscp4cFjuwMQ3FbtWLoVX
COqivGtiQjmiKXWXhQ1zUKCm8me7i4zM+M4yavX1y+W6r1veS/D1XVR/jVyp/mrdsciBY7TsDk0e
Q+ifCVxZ74haEMw1CCeh9+fc4yOkfMqHKLddljH+2Yx4dOK3eaU/1iPCc/1mQ+dl4ZSkNX5Kp6oD
8aaSrT/34JqeDEr8dbVdV7aG13ziiGEwIlo1xzlZwUxmAtDdblFSnP7Nm7rOuKR8Nfu8MhtR57Ji
DrtllYJt7Hrn6zkgLRL8KIQ/dBAXZ9wy3hR2PhGayTG5cLexeBYaghg9ZxCf1ZR5/Jg0YODKBmLg
kbMQWDouO67F5xBaWWJskA1emCVttFtdW/0pKHTh59V5bBTOUngSLNwGKXyKVlOqT7mzsrCvD5LQ
86hdIOGY8fBYfkwodgFCfzI5v+tC6scgwmdYofs5IpdeV5to4tQO1t+guB31AsZID9cgBIaF3Ntx
TRqcTCUx3s5LIcBdcWXRvhlBnrTCwVppP8ndDGe8aTjrSdy0FOO0aOS/XZAkLaNfJJQ91UcI+Qf+
KppfUQk6LKrtX5L04ypkr6ZUSdzuUj76yBL0izcWmQIe8ne532JDYbVH1mEPSYhjl/q6dWoMZBej
j+/bxIX0oAeEfh9z3rby7HOJguCSrUFm91N2Kj7zOcGg6BXeQu/DG9NJfeBiB3tXCr+LdhuHsy8s
BgX+7iOqnBB29Gc6kcOJ09W7AdeXvlp0DniBsIKKAOJS0jEexxpw4WzoeTopKraqODIduQ6INkMh
xGOeLheBgeUxBCGVQAlcygmi4sXYrQzPXdTNEQG52zNm2/kAk6iNLLTrZExZf2OcHRlWOR4d5+pu
AhRldR0xxeWSvVhHLNQDTc7QDk/q88/9nliitVTgk4zEtQKdmuGQy9/j1Q9ldGZ2c/Jnv4j6VCEb
UcB8Oe3sUql1+2KGsxjUnG6+UUjwA3F2tK5zf3XQQr5haBfhCLBt4FhX5OKaXHDhqndjZLYa6uZu
N6O2aBNP4JUUL2894fn8VIujLQcH/79m/vUK6Hf/ZcnJYEZkwMkBfkShnIYwU5dzkesm9+oAmBTl
yxBm78gAXq81XUZQ1XtyGmfPhvyrQb4STVolvyWGrbiu1YVMhLpjGbZoL0GDBnXAs7ARZ9+s1Qvt
BwLU0+Rt9NE33QTwwTeb4MEBo7pepwRDkSpl43HM0lHv/q4PD4Hz3C7EZXOQ1eGg8Ae5gVVBp36I
oZ/qyuhwrjdzB743ASdsAW1lpEzWyd3EaBYtJ+G/7sDyibXLtb5KdMrZRBz111qfqp+1qWokJDCf
KasVNa3x8Vuba7Z/WC7TmLtCbIQrBz+pAIsyQt36jJsp5+tV3iTvPcdvlhgb8JjQMlB6266CbwLW
KrK7IlP+TBAFQhmJpeMD7DA/vTGacYBKLuYTkvU/XFMYg6vtJG4TGCVwK7qfUVeG0Qw1OGoAkRz6
qzToaYELUPw0MhfmhTw/voS9dKg4xENHtTm24XCc05TE5nkofCmsoWccmeWg0v7LqXVeMv7WUNHH
sCAeO34aCA4qdoSeb0kxpyFsKF6swQ/DzLZMdnGFXmhQYySQZZ2XjV/0eEZtmgbnMaGwaLMoOzu8
rDcNez3Bv+Gayy1Z0cC2YEWjsadmexiLqfyIhYqzVb2NdgmyaTRpp5XudzzSNP3TFQ3q9zsKJspi
JgY8UIVnnIgH5DxnrJW04ZdJQfwr2Vb9plhIi0Grt0KiY8f3ebeP5DQGbZssolkk7riXirHgysqn
7WPoLu/ucjLAbBGeuIxu8UF7R2l29//bjhoXamHZ/ECjiHcXHFj0u9+Ctyh4J2ZqiOk9Nk59VMUn
YN26N0p0sJuV3eo8rFu/YALrWZS2rC9fVT2iu9538y8LfFwZnCzGwsue4tTvl4qyPQYSgv7ILyyl
RVL2rwOxEQ/SPczD/64mGWgzgeiwT0oY2aaByHvMp04Q2Jeq4wMkjBfdjMWfZnEnB62W0YoWjVDi
72LP6TuDM57hdGAY0pIfUVvV7jKGfTvEIwi0IkKaT1fDshJLs+g+7b07WdYo052U6rJREBt8yBxa
ZSa2tddg3CvnQxv4sGAEi9r4pA+uOhNxTpW0BK01LQlM589QQkcI8M9kJivN7b+1pq0DRe7X6esv
PubkfmDWtEYHEFkniVFlF2o98uUAY+NkdAfV+lxoyoNzUY9C8gWBKcU3kZ25KrtMaJAseYgoRvbb
5U3dr2FDOZi2QqtE0e0+cGlbk9TOZ1h1mct9LErPMpYuFOEjk3wNWSXCqCwf0fS1RmSxly+IYO//
nPTJCouz8cpqHha1OAXbdt3T55nk3q4pwLIgvnRWGf8guiIYontxsLR7L0zrkGLlDQKQIMQMtUDG
hsjFQjz83roEBehcrwzUpe+pix1UcdZCZYrs747GzaYdjzbuKwh/HCBpeMkuWBkrzxXKgFoTw4LW
q2BGlCTlkIMYLVYcO4ARW1HNRQoaD3zn6hXGP/1Hro/PTWIygrjzs9s2vNDacfVX0GzLOH8R/FdU
GzkJ2Dx6JW/ujYrPIJa//v/Tx8NcKFXGGLH/kmKeXSq1j+9oVaresyT5kEvOTl3uoINDFaHJaxAF
LSJBYi0yQutlMFELkr7eiVEfb7eWDo6wWgVVcxtuLF43NKdzumu3yAU7IidOFmgJab20Rgd1LZc1
zhPGXiuLlH8tbwNGxSIrK+fw1Wxfax+3cgvLlOdsMLn5ifCWHZqvUiCSzcejQt6905dtTgWjj9NY
7lMLiMYKbMoHDfNrsU3QzxiN2hgEtYaVtIvbUWHummqW19bqdxAi2HjeGSYHN+0xPsJD/FDl1yev
Qxc6LTZWs0PH2+bC04o8vTpXOXdPj/Jn0LgFExVvbobOf1np4RYAJx6qox1l2hF/a2EA3Mhy5yL7
8RKal2FReiGYZW+RV0Jlc51RfjZVhQ+0ysQ4vtjI9g6r73wW0AsqFRm9sMirZeVdTOCYQAHcKTvg
3zJ6jkmiSn5itxIvXz2DwEq6+YvU0oBK/d8BJ+g34kTBfLjz3GXzdyUV0k2Wcc7DD0IB1A2Gb6Wk
SU3KmwBRAgR5hRyMQ/ngco9SYECTxJGK2EBS63l73DzKQPuTu6D5qaFsLIDdfT77Mk+5Bz/677T2
eXUi4hlgvzYUVMuN5gjyqFTBDW9RsfbafsVV3GVgZmeUOK0fsvSaopVYtNVKXTjO0ldwHTOap4E0
E2eR1NDproSkpYitFMqKoWrd/1Vqgq5FjRqVvyw6QfrIb1i6+sQIiRdbcLQXeGkU/puH8tBOyT12
PycsUvyKUoxPsqeAC6hKx2aZ7TD5XeE+niAbfJIguz4GxZsxai1DlLcueEO44sMilssdJkHmh4EN
+7e1IueMhPv7KSxAxxVL9YGBu9RWd5+Eh3Ce59hmKOhjENZCTMMOlJPbsTAX4OA1+Z2UtYeE08xA
uAWErF/75+N9Too/h6OgpAkdU/x/xhrIAryLbcCxSCAFtBGOwN54fqBPiEkuTZnU6DEUVC6fP+Lv
0R0i5LFLgdj3LCiUdl1vDCq0Sv0I4A5BixAkyCEv69EtMr8p8gMFzavPzbmckVEqAOYOt3949XRo
Ao9pcjnIDE1itFrYFYgkamTgddQPnTBlvZvoidomHc1LgsH19FYwpDeW1TLPeRz4dqTgsBwpCzg+
WqVw3e0SDSTYI+5vmQwPukk6pK+5qPLMV/drSR6v3+dYVQ992i6bmLQRDfRMF3xMhGAlUCXTnEaX
ugH1ahzCb0rZ09SlY6lTmQimJ/68SB1bHnHAwezmnDI84rlpEEzY+eapfO8Gg5zkZEYl/ohNk4zq
2bBiGLMJykXHvpKCqK3bNRsIMCPhVEOhNeUcLAwyr8jySVmyOTtOW++f2A+QnH6KWIfj+jaqNNAD
DLH3mg85oatGEK7aQyDy+ywwBmegNsDIZmmx1yejCh44QKKsiMmNXQMIByIj+8pp7udi6mVfWEo3
CYJUhvSY8bZjgadUUtXzSIvWZ76mYIstT/MFxpNNquyRaHYf2MsK3nbd43a6mgaVkeqbbliEWZEQ
nwPUsh6hNv0pLGEZJJbKhMefUTheYiykchxq1c2HYW0GCKhpAyW75o9HtXpXJSj6HP0Ms/zxocB4
QeV5srtZ0P2OezfcTvbgA7Gvox/OrURTStZSsT22RXz2KZZP53OLczv8eyIJDT4M/ZNeP08fHfTt
Y7ZODx/L/vIZCi7oo9odsLxHqCvQtMr3v/zgXdW5pUBM+3l/D/o4SzxeG/e8iWJ2k3NT5NWQZ9N8
ZI1odLlW+lNuoeBVxz9nz/PTDrLRtc5oxgot+n7QJ7Cv2+tR2VmJL9D1RLTCZ6eZrI7zPwsLl/sI
uqr2fiRO8t0uA0RshzYbtY5Gpi/1GnxbIAT1vZ1fv8KRWl7cBKbYxYygDMyparlZrUWwiSRMrhQl
V4iD2b8IHKZdIJxuP/lriQAkPxHpXzskPu+GMKYFz1UPjo2S/Cdyg4GwuEspQVFqWmTfrE3pNICw
nqAWS9vE5cDzVTXQYQZw7MWluAz/MnZx/gnZs9WB7HL4kFLs0O3Eznqg/vIlMth2r8SXW4AJPVzA
AywIEvvWo9kxTbiZrJR4gl97zwuAQLWFwomfdq4XP9rgf1C5cN2qXjVumWOtMcmvu7RgJwVXPLcp
Szx/LBuv8ZHoqpmE6rpplYjTg0OniFHY1pWEOXkiHAFJMQl24vmfmblM2LnJzjddACgHduBL/W1M
AIBPMwkMeaRdFj3bM30osKgaay4ey8SM2xOLwr9oNbKEbmpYlBFjFtG9rRr/FxelD/rg0yiB0xs6
C/KzUfMZtW1TkhVfBpfkRDDjOHgYI6b+h7RbrpgQV8Yl+W07LS7XPphO7EwMehqgGnGh5jEEilju
454FUYxGm0l2d9OoxeCcU60okZYMUkPMHy+GvlJT/pD8IpB/0MAp/FsqKhsEvNeaoyTM1OV8oFmu
eHjAyKq+LA47wvGs3tXsb2OoiUT1z6kEzvr+5p9cK8Tr6D+uYzQ37UayYlIyVBsLbh5gd6hkXk95
xahORxvBvFap7w3wwzJiUoTaEWLA7xhsuwG2B9FtjcbweyWAPnINb+HC4O/t68bLxDwzGI9+ol25
kHEhwUIdiUwOztjwH1JrXmR6TA7Oc25sOBn67vEccjHdFWj17Mic8w8V7vq4UH0arA9f6fiJgtfF
wGtbOFhg4YarawzhZmbunL/ClxpTs1QRpvWZMRvTVHMUkKM+GHPm1uXivFk4Ia0Fb3Q8K++Qhw74
CUZlU2Z6sJ5x1VvjI9Mb1Jj5p6kfM2nm9yzwfpJxg9M5XfOllcs/w2lowXWSROd6OcDt0qpUxGuX
GN2vMP+igkaFE08iTleLd3gwvUE2PXqp/lsbXjWlpuwkNmbyPCSSbvYEZqhgbRnU9BgJBA35ht0X
sDKL19bgNhm5mcYEZ/ESN/QLO8rudd6jhiFD0bWkp4JP9Ep3HEcUdcfhRUSFccvmIgbn5m+20XYV
sGy1KePKhfnAoKCrBiN8UMg/aZbzrViKnxTGJ59I9ppg+5nLgol1xOvNp9ux0dfQqeiQx4BngEDC
/pfu0QnETnaRbA2C3moptPyxroPWI+HDiQDwF9rczFgMrVXL7czbs6dybjD59qpK9q9jbH64G/xq
SuO73/zg0dQHkiIOxpSeWYepUNljxuXCMlgXddb8Ndm2UYJd5/Ypk0t3IakOSDTioUfPROaCa1mb
47nbUriCcPeUmzagwWco0tIxse1iCrvtJSltri09dOY0SoFKDhM6Dc5X7vCExK43E5biQEhzG9Ti
8XEIhXphtwPxQAkqLj7feJk1QQHASgyLwu20AwrshSBPUoXKOdfWaM9MZu0yOrDmiXbtAamYPuT3
KaXwdP7wpSB2vwro3zIo7uAoQq4DB4wKhWVqF/GuRvohm7OpXCJaeVpI3y08gDtXoIzA+4RP1vZC
ipqN7mRCyYura5FNiLXXyCCAYrJ0cpQ5dqnvMwq+P6IGyQ4CG5Y+oTkKHpDV7DIqxLSP5RMsGvPk
jK5DmN13yI/erMVJUOgLJXNktOyjHJ59FPeLCsYl5yAfV9HYIL4jfxuYmUqAW1pLV9vAbU4WviW+
j5lzIhWzUfmjo1aHWZVEsNvjZDLTOF6tKLzS+MQ6X1d8prWtrMkDMg6Hsdc2mKUT0oikt4Hw+I0W
OIubJHSJInzHfxpAz+kDYO/Witezl9q2Ip7/h4vRpDwrQ2mVlFZ9hq4mO2OqBX/W3QN8EYDBN5u6
lBcfEH2hAwLNGPEhw2GUSf8g/uIwzg3PhiZfpCv7thIoz+vk0yx8Xtcq/WODKdhLRELDTUwYGHZt
Ncp+bqtbxSNKtM0mTLqL6Bt+0+1mC7r89OZSrCJabzONyzCoWFF9xEOi/G/u3vA58o6DiIHCRF2J
5oZf9+edWdRYp4JxTAL8vcLFUYY6U7Ic9VxyekUxPrkvABY6zJezG9XIv/iuJxtHG+YnXWW5eJJh
qmoBTnjV31H7qlZltPylKuNdTsTP7AgS0VNLGq4SEUEoReVtJFWXBNnhExiaKjtdDavkvh2gTk9g
MRXbpobd2mbTnXczlQsOBo7SbEaM6EFI8sXX+3Qd5aCeEqfTy1/KBp5EW9csGo3hCWvNwHUhhgW/
iE0kfL0crEf+YauN/VmqECe3U6EvvHzs4GGfd9eAVma7OcQDPwqIUUvlPGChg5w3ZNBwl2rydy7Z
oGe1peB+65dAD6Q+IOXuQnS4lG4mTEO3lUf4n3Qz/zBb4cbGHNlecHgHFSjdZ22ZG5X1aUE5itmV
qK0IMVxYVIJgSpkDBKMecmaeWczT/PqSbBveaFRH7kU35/lLuVVKB0Y9UC8Wc0zK/kHzM1DmG7Vd
R8/Ag5iL8Iwr5lEvIhFZFCunrs8po1bpfEnvCV5eM4RyuFNy39qJLvwO9Nrd1u3dBWZhIAFclEBr
sLSKWZql0C72ewnYwLx5iQ/on+thpcl8H+TBKDkRy5fOqDzPcPkm73m7ttQ0JptLmBmjqrgjtkhh
wwrQhRpFFL7eC1oCebssNVMrCwFAzyu2Ed0p73gLP/M8RD/cT1hpg7xtlTCgivtSUHdEqPyo3sr5
TVgmFf7iSYo98zAYy8CFEQY4Kz7L9e481Rxm1D3iWHuue4qH06kfkLh9T3SJRmEVnqpU55BLRa90
/ReHLBEDaHAlMsDOfvFB5ANGkWTgtp8QMbg+j3aNdRJZh9AG/oqXnB8Osxjt7f/6Nzu2JvrWgAVg
XhEYhQQOvARDQTltAbZffeQA4RkD+C7GFRxrbsnFWsNQpVp2xXvqMMpYVfisow+nprg0eCmu6yVO
riAIzZhS8iGhyNxd1xDO78FSi2RCbiqYD2WyE6uxZU/5jWksPsdAiZr1ukxNagA9xSqlUNfOl84V
Adp9e81Tt+Iti1h2DpMmyyWL5hZQZqs2OdHjQ9mXXMtVM80lzKMFXtnABy5dgdmKMrc6TBEpzvpl
d7EqnJ04I/rj9uby6L/CwXXg2a3Wy/6IJdayUj6LsTmnu697Vrx2TQg6NYGKOYE9zv598V5O82vO
gWrUjAJgJM++jV9NXAZWR3jwyD3HDUVbSsiB3iqOYv4naQzDY75TVAhZ0NBz52u+R0edts032YZl
TgPr6/hg3BbPANa43UzSGgjHibdymd2q1gLEKGzEvUW4uLhLEYN+a8YWKDqutMuJK2QAJ1IOBhva
SmG+pQ0WdDDaprxS7hZNBSDsbaChzmeR9yJZFI+GShpU+GLxYaugGCXYBXY8wrWKHufPRK7FxB+1
HBib6oRsKK0MYlS/z5tWV4WQK3tLV10555/XpfakLFaJHYMY6E8sttkuRy8wRWFl+hX4ffL3uNsY
S1ISdSVeXFoEYO3RNrpK/auDDgnvyjsdNpizd2lJCAUTrYYbRzhC96s0iy7EzSv5+3HRm94ir/VL
4cCUCBTcRY50vjMJMgCXhMszGMpR9M51+OneQCwuDn3QVZzO1aZE3nDHvTMaJmylFbrfa3pfQ/RO
JRH8rg/7FxzVwXB2zGwz2/Lm+V+ctvAf/pBqAjBMIo9iAEBkeHduWxOeCOg2A9BG+V5xe4uwbdkL
wbE9JoOO1Dx0OKGkYlLqac451gNSwR94hQOR8/xWNb1zQ9WFjVbgic6A2Ughq9hVR/j8oIYWKOlm
RqpbsZN8XKqyX5iPC4reiEipaEnzuzUlUtV3SR4701l0gKjBUC8jeUzMQB/ITxKEdfbA5vEKm2Ax
JYf/dRk6bTDWzz+zUHbgKIM5LYDRBGJe6UyacyqtZCmHRmK0pyAYQX2V92bvwAumMP544X8alrRv
2kyEbPRC5U0c2mwMnOoConXFetZBDpdJXQwZsLaaa/YvrW3/51uVx7/lVrua6aAdiI98ZJsEx6ta
vE/tsljP20NnCBNMjmNEbcmLvsBnYJch5admAVmFAUgL+AjkOqOICcZnWojoY/0MttK+MezkyBoZ
/09wM0xUFutV+oyoPney6r80izASDg6WkLglNPAwHzoi6LkQ7sRnZn0HFtyF4VA6aNBlG3BKeuNe
f7eLUWHlugX52qey4mjpw4NpUKzA6TDA/ZXbXrVvXWKGhHvb2Op5mw3DxvI9B0TlHk7zejf6+x6I
71myo5rXJ3AeREfdx3J5gxFra03XlNqYV9tY5speni0pNYZyTk64ZJyyCBHKyqS5w2Qsrw37jrq2
eReqJA5W5BeJDMLGgmSqqy6nvLnxxqNA2TopqXpS8ZLMnXf2vzGAuOw4BDeAPcg0gdg/5vGWTPtZ
ABLol+paUJlKbXe53FWJW/H69T/cYvOoLBXjzOx4Z78gQVZD3R7nOShZjdVkBLkyLOUZmc4dHYFx
4OHqenrCpVYTUojI2/2u08tm3Vdp5Qn94SK4IIuD8MzN5oMPnCzLQhmLNPZ9d+cJyn2vppWjfuwr
lcHlbMryCxxY0drkbSYXHb231G2+AXJF/mniveDOvHvpCjT9Tb4q7ngHNL0DbSkhWTUUVAY2UqKA
fDrwgvaPmivMtgQUkgedb5n4YEkb2aNCrujHP2xxBoF1WomFxGplOgm5tpSlOtqwbHgv3wrkBsbN
JL4d9gONLJI8BgDt23fBboVtEv8jLptxKL5uaE/1K6BY6Q8ednsMk9E5J0FrpBXt0IaqZao6NGFn
KQ1hSfa0jcqtQq/vYIib+Uj7Aimj+q+Njc6UuO6OtIeaVkrg60IJbW/cOQfsIT4x0ydNiebD840Z
V1/gj97+CX7MMB84U0Tl68fRHqgD8Jb+JB86qqd4qGVSpIPsyZ5J+bSEi1WbtZ18HN+x6MP+KmDI
AIFZIPekoagftSYGCspqrW7hswkR16zHEiYJJZ1ghPkLcrfmdLikl2SGU+Cs68PEn807n42f+uJv
G8l+ZeK8p+0ZmvPhQlJlUqAAJD9LfQQua+LhHE3AmGzGVmPQE+MLcVTzGKJA5MbgqdpbOmBLCGkm
Fw45vza/1kwdxuLxUjN3l6FOWp1LfgjtZdbdtYzTtpQUDaqGSiaxVV1NTY876GC92HU4AhnkZHEC
+332ub+SZL/WYFKj85s4T5NTBv7rwm71wyfPM7s3RUDCt0n+7WEzJ7ADlmXD1GCFIwbPbLEHELBY
iPVFWZW/dCk4nskBgQFBIvKRmF3Vfnb1vG7vquZTX9myu1zLMpulC01GMzbng9zhxgjBhCsmTw8q
1C4koWGd547RvGjUxxHOpQqgLcUy6Rwn5dUX2hlJhxPzmSncp5S4fROjO4llFltSkVCkQXDlbdAM
SzCnX4+sdr5GNyK444g3Xg21uhsRWvYPdnKkAmMMaZA9RbH0lP7DsGzD/TvwR41GhxMtJ/+sjabP
bVpRvF7WtMGgoF3Cu3WXF4+Wt0CBxylMCOspRTNGP33WS7fVprtRbj/2Mn63lbiKlbEcJJCPkfjt
NM9JGbBPOAYuijntbhLwIdr4bqQrbwtJKNNKvxY1y8LAikKPeTQDK1gIzPlEgUl53gQPMWH0iSG7
uIdbU2E7XQ4OiBsJ84BewDusMW5uxG8wj9IIGCDk60eCu2+vPNyQFz6U9SBVacnNS9UI9lY1/d99
gsiVgtec9E9Z2cy0S7zgU6VbgmiRLiDEnSv1EsMEG/oEoxm7gODRTMxmcrBDHucwWm7FuDnpy7Sk
zmBjS+EnNMgl0zdKNrErxlFZoCVwDyEjUwfoe/feYQgtUMtwZqDUrQfET9312TC/1mmFJXNPUCU1
6pzvrI5F1mZBVXq1YyKN8F8sINIUX6prwwduJl59Y4ielActxnyiVE/i01KjAXB8/ooyTz8+WdZh
vx0rcdJVe07DXkaXCwPEQVKWoGtuhCWPWEsWYEvp+d8pmf/BcxanG1hKVGCWd/iV531c0anMKraf
3VDuoJOigDE8aavzjxjqECw15iL0e2GZN7+6kcHF0ajSPuYTAbeLZqT1c/l2SoGdEJ89QDIFj6jJ
hegqTto2cNyl+4Wk9/5rVf9Fbp/3D80S/vEjPoBiHGUD5zap4bjpCgm1bX9lmgVu3KYWbJPG3xbF
e/7BD3mdz2D4W4izCw7seO4da7Kw2fbYHTenlTVpEEXJw8ZHQCPmEaXlAZabW20U5VIdOj2iemyo
6Wj5xB1HpGjNjmuelYBA9HeK4vggM6XnzzUhphfzBujCoCcAVQuXJu41Gllvg14ha6PCOTuhHcTf
sOaDQeGCxdbkE7eujogy0hhLm7JpuJmfpH8JrNWaRsEcVXw+RXl3u268cq0HgWC3Z3BRb9V6hQpv
+6CNT/vqwSVnyjj/aAgQ4k0pi+xpt6DFwO/3TKO6mYaCcs4gZD0uVLwM8lngsbhRVqUwZO+q94rj
g9r0j+yGR59L1BXSY9VSkchNP7oapoAXDScOplnKgHi4id4J4ov8tVrIVqtLzqNpx3wkHMwM32ja
hf1D+/+y/p4RIsdl0Av8dPS+CeVn9UnDH585YutxcEpYRWHYiELykiHnSFpJK7me0N54k3syd70I
Vl7hJllGprxpIkBNZ76i6HLIuqMDQ/yy0h07rR/C6wpAAg0x0Y7l3xbOSwZ4bOPoClPaAD4CLp2j
KF/74ChUbTzRdInbxcSCpFRa/5cTlhZczA2Gexw8ODGyK6jg43mlvsoQ/lifS49GlfG52WsfDVWi
2L6QCD7Rrc86hCZvkqkf8Wtx9z+F8tm0NvpdV8m7QJCN1f28/zGfp1IFSUMhK1Gw3FEQBGSEc1Ar
5FpwQYPTfaJXhHn0Gl1vHn41lPIq1ESFuBKz7Lfz62UhsbyWI3suacv6GLGgG8DwYolA9n/l+6GF
sxGaiXRxpemnKc7PzMpWi63nJWY4oKjo3CIctcuZ3otjIa2bYlkVYvenNWsvNVZiVe5r3D/j8pUp
EvQWQFJj9FvKR/VBqZLzEvDvPMvJO6kHvE/F8a2wj/KII1ylsFVr5ipCp7zBVKFaEif7a2CBwt7U
zLf7UoZZ1JenK+he0rALZF3ohPi5IGF8Co0sLjQT+vnkdvb3PlmFxNwa46LHWiJ7v8MBaU0kP+sF
rK6RugIXSEI5KC3yDbeDb0aHT68m+8ROnqvCPHlqEH9j/hyB30FFbzwdfbWrvKLfVT8lL3+6NVXb
pKr+ShjEnZvpBRR3ELSEJE2qiCFxx6dzY+cq2jMzQ0XY0ja3PVpuNCDUWpRkGZ2j1FRgYQsYV8vb
iIsjdcEvliTpqneF7OQxbta7wFdnF83P+Onv3qJOsMoep6u/XISmqozOQmIZJBKDvca/ICA0eoo6
37AiMsDu5t0/rXeI8h78l0EI2b8CShJ5eDm2/FZe1R4+/j/eSmh46cDrSEmJgsIdqMTGbAm9f/uZ
RAd2OrMJarAf/ky5/d7a0oXLCLx5xzQZzmWmKodeTSjWjX1fDXZi1Q2PvphjCwNeNAHBZc0UWhrW
goJ0w2082rB4fLT+Pt4k9pDIxOTN7+a7l+XpdTLL/kCyfiBlisNGMzU7+kSCEWr1/6wpaLJtgPlV
eoxZChETzQy6kXawy+TEfhvQ/07uWlprXRjnrTXiitSZR3D2qHnHz7chZrsIBzHckWFwupudOCSZ
YktejRuycndvHJu5LQuMk7CJ7qNXMSBlspzbe6dV+c8d/WNtKw4bKLHdSHXunc0fXKTGkt1l1Val
uTvjfpdC4Zx80c/8qLrJqgOep4A1Ycou4AwIKEXo+Los14xZ8hrB93KJE6026F6vRbAb6ziJB+Lc
2iyXiyca4YNauH362SIAxy8hbx2aFrVDejRmCjTr2ZZNmKBAYpwPFxojBd9aE2dxA8sbtaLLVNoZ
GnnA0v4/ls0CspMnBXFHNTXvJhSPtVvJhW0N0ESrhfyKmJoKXQAXMbGu5WrSEX76bmF7Od7CAH/M
/AtjP5SiBj4oavbGRv9PnHeGHSJj3uuZkXgETxuqMLdFqJ2ebVpPQQXqUFtjEHvGQbE+Aw0YS9SE
ENeBe5Bun/pS02+OyyIIj0D6UuiPhiEaVZvAYTim8rP064YajOpE4nujQgUY6n+glnxwre8W98Tq
y5RrUF7LJEzsrOYw/4aYcYLmEjkZxRlLNQnAzn7BVmtjnIEHGjvfRTIR783isJJxLxBv3wQON1Sp
ttlz0dccftP79U3fvIt1qJEv4AkSSZ1zOB37v3zhgOlqHP32Q9kT72i+FYXi9xEq27tum221xfup
uVZJMb8JUpgp9NkngLAJnAYMJiDQTdQp9MP9aY4J5cTCMQ8VN5MgfqNRzIIzJ0xjlsfJBbwG5km+
yci5g0GS8uRCZtNroq0FYbQEOVHIVzLslbJlfqIZvpDKy8mqHtGoRcL5Jw8MiBjD5EPHWabwp1zA
J1AmxpR9/vk+lFP5EcTsPEt9keJcPAd0UQTrv+I3gnm1o3zhbD7lPlDZxuZvxuSdfma7aI3Q32lw
oZzrlSNV/gRTSALVRupIRWnOZkFPOWon6XJfoL97H8VY844kIEfzaTlNi9fsPsYMsFagvTgtfKYC
DKqTiEe5kqJlVFSCIby2GnBqFl0AAd2aLvh2qKPrSyqFGcEUN1S8J3xxrBe0u77ArSJuK4OtZ04E
c7NF/ZGKs2APq426bFPVV6RfArFHMhJ7YfAkaIceX7JXE6pPL67sV1nb32AO548s6sXkwd7zK1NJ
cGY3LmsKRqLuN7mu789x8qC79Omqj5/KUK16Twh9OXBr5q7wQ/YTNx31sdBw7heaFeIZ5WVVCAoF
omrnIFi/DPY/a/Gw4aqsq4Ywl+6CSUnO+ka3JcgKRbDfWe1wOVbdTA5iDFF3eXMvetTlsVZNbAeu
EPZzw7QTuN/ESz3OsnopJmfMpV03nSzWlQ1gXYY0TujwHRmxdCcw3IhS/IK85auanR1HCcpoifiw
P7h0jp2CUIxrw3jKzO4WwDZ5ghDW45y6MeoAJ42IZ4er6XizEqZFtsIgp37LUpWZREQ/l1lPkAQn
Vybxq5mBItS6uSxicZf3uaoOJctmf7CMsdXTcg4U31luLtWgsoTcAtPOIkU6bpkCRBoqZhLtpknI
kJTcuOvSyPSz5Lcn9kwMDsXXYFPirGIuyQQhb2Ok5ERltwxCfRuznKUmyjvVOeBPUcldETJFSGts
oxH9TCSVw5enDfAmx7rAlfRA7LFcikfUi3jpkSKcBxDaqJU97TS+C5C88+muWzFWOPucqSpk6+EJ
OV1NnipeMCY3feX47cytpnqBpY3CX0wy2B3oE/rt8Uw4oVpGttYTozVrjfJFMVwiYXO4vNnypfa+
oSwUAJiD8W107M4DJVK97ZOXh7muAj6YwzcbfCN2B48O0oIT5IFgxhjmNR5f8DhY4U+lStGTSHYl
XClui346VdTUb7zL2T28p4mwrMSXVIP8kDLKpbh4GVx8A4WJebGED2QOMaa3SZ6iHyA+2BGjHXep
Az7UNkMbGnKA6OBD35TNu7AooWXTO8dOfZloyyahnqVB1J0xj+NTCY81jebBb2eAlv63z4VGaqwx
QI4y7iDMjBf1nQuYaZBa+Qr6OJifDIPEE0IVPl3rwR6raWz1OSBM0sMWD4eeuA5H6BK57YsZso3d
0gDtZi3GptRScEsNc8v9WfYen4/lGE0O1a9IhuiThpDBpWre0schLVx7VslRSsvsy+CDqHNsfdJ3
EIUHsZzLhBOXAj4EDEeR9L/n6hLZM2TBvy8PiQcOyY0mDIHKCFzbbAAAXwQPilo9LQOcwSox3W86
ShJCd4YlWXDZuMoDV7gCv3gnCCM0c6JcC+VHM6FuHDoxYPrDfp7NWlyeaDp2FiSqEnJbY6ZpGQZY
AfkKB5cL0dbXyv8lof3LAQDsVMpvPlRsBI1gpzHxIGW3924Q6i+7c8jAr60DsKfl/HYvZHQwATpk
9b7l4DXAOasxbQbALdgYJvOa34fT9LqCgOAX+XjMP+WhBTDOQ2E7oftiJWLcYQW8OYq8Lv1VFZla
2YoJU5sE3PnmWu+7kixHYWV01gsavV+/dMaxbby9BfocJlYVE72B517sv1HSaLsfy/xZlpws22ny
8NYd9B9gyx3Ww1yVX7sToW1kwxBVFTn8SrlXaa4Dh6NoIDgp3dE81dptwOGSnmiwGtIVIGmG1lm6
+Gt0zT0b+GhWp7kqHAczaaW6JkDGBAvC0H92ElDBNXhEpIZo4g+rpRsfn5Pghoj5X3OmNcQrbC6M
I6Dp1YBl+PxqoCurtaTNtrUGAjGdj9ViKYLPrTgde/dvjtYelBJcNI2QjVPtQtVu4sopxo5UlhJH
iqHtuaCumThn+/ZTKcToTLNm272VdtzDUjA6T7VzvtXRCUs8DQFjeqBJQLhffJlwNxsnE0/NdHUD
21BoZGcl0e9M2ve73CamUAxdgldcaqw7e7toeFdTwh4FCj4J6X+l220tnkhlr7Cmmes7USQ6A842
GBM0lhNZheOozKfoIGK74EEyncoYBU8HysdZi1pcnUPY7yKbItaGhbusx7Je51RtmxNcUOLe+Coq
HaP2ejJfavJ69DKBIcgdGFK3uJfnaLND0oQPyN/2A/R40KY6WOikVNSma/9TKH3Ixxm+h2F0KzZB
Q02x9oxMkwWx7vwJ0AVkxybMxAYmLbqOfQZTsNd7T89cvzA05OzV9UepN6XnQavyEiwo+SIAjfy3
kLOZJHtDS3XXgmTLCIYr3VtbXtIgI+VoDZub2S0dfE7dhoiPZ8gwGa/TDUKUi6tx+Sh3qGtlwJBC
6X8m5K6rgKRhenCyqIRkau7+HiZigUfbpaJMFfqXqKAmRkDrb1VCGSOIyQGDlLwMd0sJLPJuNJYX
7X4qN+/vENlnQcWjq3SaekKTfSWEaW/zKlMj/03k0BFCMDU+TtOLoVmqwm1FngA6z8susYycjTpk
OiaetlzD1X4Td/i7iH3svhNi/sW5lUFmuvfnPzcSKHrJ/rnbRrcP8Z9Gu2L4dHX9FANW4kvP65b/
/22jnkm4pskvMmcZ1ec6tPJ7w8QteCawHGai4qbp8/rkPQIuToefTv0z3eTNvxu0sicERPV/O1kN
l3QuDrZ9MwT0JP+LGQjCncpl24XBsSLrhMspCEc3JqdNzXUF4i9Ipptoek1N4Fn1dhEK9TB81c1O
Mqr5WSjGlUn8Fp5mJwIILTONOxBW2rYuEAdE2YTD+YG+3iNShSmswd0n+/ROMZaKbv/C7DfxJgf6
byepfHCcJphSgr8Hu2LaecE/hXOJYpG1+5nK1DiOudxA4daQOUcnzmyR6cDEYh9IVyGQrxckCeG5
tn8Jyjf69mRBZlzv2BjF32Druk1kI0BRg+G0qUvTqWZcMqcAOSdfuo3tACk7/8qYR5wPWTJ6hWcG
Tl+TBE57vs9bYdgRiOyFFIodM11aAKF9Qo08JlsdqbZEM+/wNnYtGVAN8khBKEOLJImapG1Mp4Bf
9rf45g+9APshTcmiub7PSoFfxc6WwhhGPQCAcyquNtIJiilc9HWxJzACF/uqzrUEFXUaXtfJ31TQ
Y4wCVZGPXH6Rai+GEBfdagfw5w1mgZI27rkLlCZflr/0TVKuKzBW5OKXtWzGegpdsDi/gQNN91LB
jeEQ3wanF2JodzWBCo7EO1s4LwcsGYT6HWNPrbVBsTHeKeFOTRJxqCMk6Qes3uxTK2ekd+RKx3V2
vg2dch5tq5KtLd0txCK3t462LGAmJHaTBKRNEHBkCycTjtVVZJf70i79Z2MKNPiATEnMJ2BxTMvG
TFcUx6Iyh+MLFwkkEJrYZs1ehYMFbDKDI20h2Jdv5937x9r3BZdI4qCkGYbPRvcKbH7PFuoDH1TE
2J/yVEH59mtiRiiVNmK5M0toWsRjj8+Xb3Z6csbcpffcIZiBCNSTDVSzaTBQiXoS85trUOefcg2I
Q8nVK0bVN+bOk9ncYCTJrk+y3Kl+lTIkIGS4AVUb1PRk/TT1XeNbc7RldpVHYXPnM+d1DZwBnksF
CPxhMV3MqaGw376TuFWFkt0n4SK3HLXlSpiqCSt/I0DK7mReh7OqXG3bU3dpRa1z5w2ildEhprCp
4DCtHeFHYziHfnNVRjnxHVclxOoD0D3IhD1WhjeVWH+GAS8IO9yZf3BdBHh5Kf13fxl2sn4IbUk3
Yqe0xRUTtNVEGXcerlUwq2J2SDc1gvnZWkzVgm4m9YjsyPVqgMux4UFOF95ELSAFHE0nX0IcNpnY
Wun4uCQiw3bH9Pu/eLqw0QWGxCjSfciH84+We3ogNwnn6iRztN6Z/3RWYgaaueRDKtmkQL3wxxY6
6szDDx7TSdV5Ghb2s3vpSgwTUuWxGYg4LH28gMKxwvEbMupmhk0qcpOhDfqlmmI2aEYRzsv3HiaA
f8P9bwqUBAggQp795I7RYt3/a5Tr8pFaCLHLBrj94EoTA7jFt5Wiq70tZ5HXZWFKVfbSrXX2NFxY
MTdrzKsURe1e62YN5V1IF5sSQHmIs9GbKngiRIEJHKqsiOw93O12midttJLR6v1RnLaDBMsl827S
8/upHf1gDfMSDP8DDwxmeK3cKvTRVW2fa/zQnpxWhbnRI/jVveFrmvRqbSyUOCJY/fjme7ee0jFl
lETLCNY6+roJbdmKhxRtt8ScEZS3iuCAvxuw9gIfPkHpB+0tJ3hAB9VHS8AZxFYiLzoQdMu6S8f2
Eq2r6Vkue42hph9mzHigxUzGMr+oab2Ue9kYAofZ+N3vL/l/LnFLaSlvDrsfMh02M35Zuk6PZrZO
3sS1EkXWlw4YHmIMzY8M8jTGJQUTsLKGqeMWTmXezn49R98EZdJazotHjRCBX4ueuBV2M/0eqd12
pbzgwPNHR0mDZq78HgBIGJYgU1KZFBMLf1vBdX50nrbdkbMaqCpCl7H5JQ3207mDO7wL0ReWGZlR
s23J79j0IDU2L139YwDbr5FA/I1Fn8Btu9w6Kptawh7LqZQcRgfR2aBFhFaepyFFwtGqJ9mCqfx1
i5gYA1vemzcJkMLQwIusuyrTUgVXj4K40YBIVD/UcvZEYxwUc89G9J23RDghUGCo0YT+HQeKtSB3
/DObtnFc3DSJ9B8SyK/dR6MyLQBEohpxpqYTEcSYPXArkSVom8WU1Mf+HGFtrbzrQ7edBCD640dA
h9r5mqA6cxfHehRm8Vc5IM2JtieM6UIRP6ItDleDfRPQ9gTsZ8/8r3NI+13meox4iFKyp65MJbhT
fa+o4rQ3/IDmWCS75h7lmNDaurP3tMpyz30emb2rE3rtZf2y98Qt6S/4nWy4gllHMpgEsHvKNMxB
hGGeP2dW1njcVUT8qL/JiU49za2C4vnEM3V26nqbwhgckGKpLzpiY15+2zBhqbiDwiH0GGkeNKcR
q1fF8Kwqob6cfi5x3gcWEYmOuj4L5gQJ3w+i10w05rWRddl52iv9FoomiSIfCv3/B2r3g3X3P8+w
2xNLX2dmJ4bCpHTsXuo8kGOassiXyRgfv1pVK4yi4q9spcgBsofzzBTC5FN+KXoVN9fUAnPmdN1v
41urY1OKABJIdWYBvYna+1JWNp2fu6xrmTHh73NHFLdQtacYvqgSq9xmb8jUsSPZDK4suMFckSwW
kDengw27cB/TCa1J1tqMm0gkIHFqVJZbman6c1B4FfgZjOtUg/4BTbJqzJwsBvP+cY58DWKzFEGW
BehDKv7oIAC+WMXpz5fEfrto3ITLyUkEHA2Iz0BYwIeJ387XR1oVgWklTqta+/uWMUi8UO1wY1B4
WhsB7Dx6RbZEZfYIAzMu45MrTHmQ5omzutZLnEGlquIBh9NUYRTFbSo74py1dwR9V4pq1FsHMyDa
c5Uad4aXlYVWGyw5Qk3RCp74WrYaVSXZfSPYmlR3ufUs/5VUTrKtb1KH5o9hgXZmt2xxfKyQfjEf
qhLRdUtTmzaPjvokP0f6CJ71WH+pqAqJlr8Gbpzt6/aXEWrKp+sIxYPqV4dxpOUdHSOmuYc7qv3y
8+ZiaqSP5h0IdZTQJydy//fAz9J47mBGXhp925bvQmKhvlczIRbk4WQ/fzaha+p3Q6cMiRTCY6nZ
998p7GRFno8CzJW54EmwpHfkDWJkNVG47YHxK7jukrUgp2HTWQIyHQpY8bdWS1bU8J56YyAFtlCD
lprlbQyYfO4D/9DLjKsSu7smntDe1bZQ5bGe+iyYpNdBLkK/ItHuXZ4CKGBjTDyBeEqYi9Id0Xsj
BIGLWIshNd6m5f6duKj2Ok//b+06kMwbJUOHPJgJQMm+6bikfOSQpU3pw3b18XE5k1c5UGumyVes
Y30TjxwRng2UYt2+x//Ns5Qy1fySpGACJu889ev7yUKG1DzM4NOYiliKpQVZixEx9LGRR5LLdgCO
CVfEOXW6wksgUus6TvFJR+gRh34OeV6R32i9Lb20OoIFWNqHj3vB0nObUfMxD2TiZ2SKHGaegTa0
DZEPN10Iy667K4dLDehq/aPWMn2vp7WNSNKOvRL1Px/f1ggl+8Hsa4jBEJ0/YTC5224VT2IMKBu6
oMYv8ugBU9Taz0ZNeNINtEBFPejsmfiP8I7edOXEsgVcEpswQtf7caa9mvGZjPjKrJefOtO+NiSl
e2A/CQ34bhwN4OIFh68RWYOZ17YugpwvQSFxZn5SznHx38N6MPQ8dA7y93pKHfPtm4h3Ocw9E3Co
6i/oIVmdGYXNO3JhNZiGA8xmwNAuMT+g2pVZ2WdFXVy1Jocy7T97AfVoBc7x6iFalGbkOJHXZhX8
xM6o3oUScKDjzKKVHbbYmg7R333VDqPKqRMVpwNOjUX6oM+FXgWIXCm3Bi+ebc8Mtow6mgpul6pE
cuL6VffnsDxaOnB9tWgu1ihgYxeRofrNdtKFhDlSlM+P8LhNXaRIelYhg9IqKznLeea2dwI2C6Sz
47O5wxyeoR8jmxSps8o8uUQ/m5ywQKzuNHAxYLHmMBZXnUKsEdLVW7zSTG/oU2h1UOpJGPFwDaPv
1suHHC2foZD6IosQ6u4AKmXHF1ZFdB7LuCnNA+1yV3jwSW4ZrJVwxXtm0etDyn07G5QT8oxeF2n7
g3cga5HUrDzqrbWzmwFZchaAc6iSFuW/8TSh6Np22Rz6BuDwqY5zv6m3C/WGBCT1yY7GMWNb5y0f
01Gtw2bvGzfn6dxPbaJ03DmRnCGzFZn9iDm1I2y3LHpEnB442l+f2AJVFazv0spDw42txklU1r4T
NQNiXk/kvW02IQi5AvVUk9XUc6VIv3IgVBk1ehSEYEi/8XPATttCHnuby9aaa0bXjBd9zu+q1Pyf
SG2I5sB9AsfWQBuM5MkHHTgqOURhFq2A2FaC+O3C6wmpJXXjaufBg6x5XLoKhOF7Izhj4XlmJNmg
CeUCKReZ8vt5FGsfQBLsc3aFPfu+6kl0uY5r7J857Sc9+oWZdr5x4V9hZKhdjjYxPCjBfINTgkSK
EIoggJzVrcQSFmnlNdOKxjFvZf9xnyySe+J/6sNXQ/tPR1+t/aI4YWpXlUSfO+4ZvGuebuGRS5bC
h7x/yPSR21QLu8NvQnYjwQZtWqv5BR6j3UbJdbAKWetb/go8AnvAwpcoOc91DC8ak8ug3x5ZZUNs
Ze6wjjEtgAo3Kdd4A5iE4LksczidUjRGxc09ldBb2PRkgZRsM6aUcYW7CR3rJXCqNByMZ9mCt4vB
KOlKIIyD6bjOc550amTJ63JnHrmnZMO6K+Obz/LsxRCXsKFNlnp/V/7gqEw/YEZmfwQPGlNWRDHW
uE4qJRdqeT2MIIqX/Ns8WC6IRgVzoytlmR8RAuNjAbNVdalpnTObz7OqaoS8BY//mp6z9Ol38TEm
bZdPxuU3sEOQ3NVTxfGJOmL+Mti0mIxvYYYX3QyN1aivVo2H7S52T2lgHo6klM+tvnx0D1X7AS9M
kZuUTzLkVDKzF2KTV9BtTFJ8eE84MZOVnd0zDw0cpIHj1smQ8/kLKGfDHSl0Mn4JpPGofIju4cs+
gnZfFq3W3OKkFpJMTP+4P5LxXN+SSvZPepwdK70lwBmGuL9DoEDW8u+ekMxmlTCO5gHHtz5Ddi8m
7MbqLMZJwfpb/BnbEXdJLjPGZMFpNpAl86Pr+P+WRai2A3L5j0r20OyYCUDeQrQ+8oPpJV1XKjSV
LztHOrhgxvV5jVV/AC4VgvT2Efw8wHPW/WCJWsKaZ8nMbvpTNjshoBYwfV+iwEEkeelUPOecI1l/
ZHjq+MNxvXMx9QBzA7sgJTKYvyPdIFwbAkQiJ2SaEn1Vrm6sSyFpG6boKr6ml4cOVs4J/tvPWwm/
kTc7GsAbnYZH+QjzhM/jw6hE+wNU28t0fSHKPlW8D0txuObi1ihC+6oivQ8RERPs3Ex+UGGRvdeO
sQ//3zV3GbYT5L4u+UOTuXfJAtGYtjNAHChHHLtHsCPu44qWhiCfw0XdpDJAHO2rHIwYqLmHsWLX
loK+O2yoad+/bZcX64Ykqqi2dEcKCpwftW2CmqqglnBvgS9Nh8ggSdWwGp4Ehr+nCAjhskrll8T5
VJv13ciLt+JoIOi/VElTFt9zwLRasWIWxae2yrrI/bYyXEqmaXvoQQGhj9SL3ag1gId6qN6W09NM
XNjCbeflwLZliU0kIole2NhkT/g3gO0UJO1S9pJrSbs9uSqi+baJetaP2Vt4AJQcWd0pZ1DSElST
e+a2YSp1A4f6O/n+RMx6a4dTaE8gWIdPqMW/DvXL+Lv49fhv3jPcNJOSHZ39T9pi2sJdR1nIiOHI
plwEPJrHFgoAc9qV2q2AlcTuwHU9nf06VIA7W92HXjV3RM2p2olc+HWelS6bdhAWI0yJXP3s4C8K
RBmt0HnAtTnXfPOwUu7Thd0iuZbRTfJJwXm6eyGjkhFmYFfeCn80h5rc6U3ZMMOA4AgOfFD+TTav
haJpLuaWf9St27k2cMTC64Fhy55SGAO85WJ5ij9KnYmc3LpviEGiRD9D8zDhvzxEfFXBFsUttLpY
ZBjycnbsPJX0dqD+KKCMUY5ResykE9LuaKxDyxmXL47C3NX80kx43Qg/mnpTYg8uS5qhHuc1Ykp1
4RwmO7pGEcGtUH8QeE8IgHvLPTsuihxK2PDKv/5DuHxsyTJ2oJ2Vvt5YZy4m8YW4Uu+n5K3vHWav
J09wA53XYJyoXv+L6h6VwljCuXjkbmHj6Fhro4nRiApmFz/PY4j48rsphTOAfakBf7ogKCfoaDF/
3PWsgj2o9Za5zRxtvA0lHVIKZCx28jA6BlGWrfm36Pw1r0Fg9cLVCO8fdeSUOxgkPhaZt6TMJWv3
ve0ATp+iKVOALNBIbdsgy4Fz1+axKZnFFqxHbP6tsKEfhwHRzdskQoBhSqcq+FwYs8ZcQEHFh4AS
/8wp/PxH5VzcfDf2keCC8ZSvqiLMDxxSGBBbxhduF0A7rdROQWcDDwd+C44UUQn0qiauVu5igdPB
eGAeeJnLXZ4NOCKBROSbQCD646WMOHWAP3rAvXL/TMv/cWA9HIRNH8zUNLbo7Rq69hYjnW98ykDJ
nanS5nFJLXCy7Zsbj7Q7hdTzAzRXKLcOrZ8cKg+SzTJ2X7cTtV36ceqRdVa7wxpNU03d3oQqgqDR
7ojwHp4TfYHirQkpw0CD7Fuzt1PPLG0rn0ad8OJVuAR4XssnNBPPv+E4rW4rHeUoeUHfomP7mwMC
P4uXKV78jpqumyBGteI2fEnimDvXC7lAvoNBdUZy5Fs1MFyXKrsSPbRouZ/qu5kfBj7oQ0MZiTOq
u73Y9nsxWztkYfV0d3Pom47GOHXP3TAsTB2duXbZPunrreDfFH4JfCM7bh0A2msQntU7L26zuYui
OJpxKhxQYc2GIu8GgY6AUyv4K7lkT8DfjwvGqLCgvrOU9Yi4vNSY9+G5iG/dgu3X97hOopkVtc+F
T9mcVagUL7qysLAk487bCPY+cp8CVt58uvRr4nwd4B0Zu2UI3hzlXe1Lb2gaTT+meZUyi1tcm8ji
beMdtra05FqpHuZM8l8eDx1Ajbh/jAOUHxhTIyJN/XiI4ix5JSKzWP+t/oSIfQPtnYhGfk5G28r0
U/PeYKQ8d9+WjbHMaJ3KA7whIXKQIqCdAPOQOhzwp3abNHSuWWBH0epzbMcKdiGcxuHEHmHoD/hy
nW3P5WuywIJz0otsHJcllK2pArfuwo4hdSa9L2c0YEgVpT71fqCYSceLOpOtee95y5fiYLmKtdUY
yiXeFOuU0DOcwj+isD9FB6WOW6t96EbZWXmsEnhUz6eSk8ZNWKZvJm7HfDDIlhcrZnpStmsHRaN/
K2lGMQX7L7MqbDeyKlalQyG1qBqG4rbG6z9QEUGPGWwnfb/h2jiKoVBwLRYexGRaPnpQe9wie63O
IPqgntYH2PVZX3U+E64JE8i8olaxhpYOyiIWHV1PGVxlgqMUndhhCP0adzOxZq2V6Ujt/TBzDjuH
cAkoTOM27uU8+LcsMamF2n9FN37PYqviZbDvLM5p546KVJ32i2QwDjGHHIYxziwNIVvPvW1GcMG8
4dqzA5R4EQ9NvG2HBiD0O5cjBKTO5OTuYvO2eILixLSccO1HRSmftV2r2VCg90aNLNUkY30uiVyM
KW+bMMKMcycT3cHw4f0Dkwjq3Vh+uvGBNmb5fTz9UjYDPzs5eergX2J7F5ph7Ba+Gnp3NUExYXIy
gAWN0svmuFpE44U8RzV/MJURJBJifBIXlDNRvJ1l/TOU2XqR6iZZ8cEIBKPEQtnUve3Z0L6e03GF
fcUFpsqiWiIejcBt4nvHL3wy/28dOc4osWaujOmEPRRAzXOYqbElek1637OQVRP8jtct6DPZyBwf
xkoTojSMEc594RorP8aJgiRoNV2W1HJ0h8sWnOCRkaDILYD6hlKKn+dCCWXLmCQsPLY59ZRs64L5
7hbU3IIqdkUMaETlI+0giga+c7VujBbg9X1DZHtIrSUVGWJzmoodS33y8Lg5+aSLVzSZZkK+THx2
q203dxVeXpiL2i+b+0/piUntLARdYVrFla4UiZeJflSHwlPu1bhdMOIZkia5WFMKT06qb1gwnFv4
cCQXL32lvdLvjOENotcbed0mrV9ecb6iCkVrrV8Mr3WRm5NBI0XSwDO9TaL6Y/XYzq1cdlmQ9l9I
CF57kOgao68E9HTYaa34fdE2wcZkdE1L6f3DtDHZxq2Scv9cE57fPtpR8rAX1v6hvLZa/PrdwlNq
fsPcgVKn2GjlDKeuDAWnzdcxm7/qREN3C+LZw9lmM61doeWcSUK7ph9ccY++0W0yPbDEssHtkSKt
kAep2FzOJaanBmWNOHuBBbFla65X1YvehFeQceKzzhfnvTsY+CWnU5sQv3j03HSqFAMr4nmijyZZ
3lfE34sSMig+QEGTB10N5SgkVuVQCKQWbgnRUZckrbnn4eRMvBAFVZJow7CQ/2xYx6GXlhhjN0qD
fjOE3AlMuJpyHf3VeBdR8+PgPjBEugpAIf8gjSW3Bk45FxfhMMFj+I2wfnSEy/cSI8KCJxgKSrqf
rwmk7kN887S7npF08V3mNLc0olzBVJuBLe1azTRooX8FHY30rAzA+rNFLxDnJmWQ2U94RJa+Mc6J
deap4QqJ5k3o5nHRU4Sy3O3OoSwHkdcwEuZYdP+o9TXhyMUd/biLD7C6BXfFPHiv0cWxLj3sVbc/
Cdvvo4M9UeAp4CC8HE3fUQNDKlTAZ4ql3zW46evazkOhwsNxNSypHO3Y4ZcBLnm6CVOm5UMusRN+
fOhkydK8CKg3XGxX2C3VFg64vwfF//C2D/QbpRjhWnrQyyJBDP3bLeNNn5GpC+JyCZOAj/LBfzG4
9w+TDAzo8agGdHLkFxqCqT7hUoknd4g5u+1KIO9UI5Qu2FbVVa2F/vUOa1W6YO9qCq5H77I6brt8
hRi8ZPOWJ0PVRlA/QIk9yBJbL96OxhbLzyFUduKptOfh8s/radETvCjb1uhU3J3QLffU5UzNUSHL
Tb3L7DAnpmAHuByTF+HzKdX/hyKzEfcYEwI3bAWuIB4sQP2C/0ta7bM/T6zNlwKiLX84cOVoL304
rUkN7As1C6gxShqkXhp/kCZru4o6xtOZv+vf5MPYkRaQaDLL7c7e7WZRf7h2YqKtK8hz2KINVPMR
yiOHO6TGk7b8hkm3HvTVWQSR3eMAbuhYdDvL7ANINOjYpwk0IWO/X4fLdjSIOg8P4HxT3oCU1KPz
R/nC5hTjPuMdKP9EPoYpGVWr1Kvs8YzzlxPBJn09fBqvbFcE9dSsoGPYw58SGUy7vv+uSno/24gH
67KA/mca8jHo2yruCPMd7Cg6EGKBDxxjJhyd/DHa9Zgp2ltkcvI7Q3NyAZ1A2ACv6j6T36C486A3
1/6eg+L2pR61U7SM22dM2bt7Pb0YYf7c4qRs8q2NyDBo8Kwsuy4idNKoq/LtEe6r0nVZv6IhDRhr
M3B3k4S/o6RN8xKY64FaDiR3Zrx0NqZX6IIHZKXT+0/3U2TBVwqAZNkuxHycyLp4dnhyYLqOO5eV
0m5CrG4dkAK0WLq5N1XPkdNqZE0dfq4sAPtHeaNRwRcBi8I08ZpmFEppYXeYc3SUoaUt6/+q7x4v
fkPDOJ/c+ONWGEN38y00Ui+3qp1J6ckvawcg8T95wJOe35Y7+eBc6w5IO3aTWei7AGjGgWVdH3aO
WsYw3qwAk1izt3K3oY6MqmDUEbyHO+xkFG3DFNrGj9XlsuJ1pzbQ6jCr9SpTxiWKdBVtu3dCbFSw
3+Ju2DXUJCViQTZdRtBvFoi2sqLkObG7zFPKYC39CvdHe0j8V5uqF7g74vUthTNbgqxylZZeepub
mRt/rYMyYwfZTzDmiZCjCbJrhR6TlT7gywVe8s0WrkGxZIDa647tBcKgLW4YPNMv/FmJds7l52+X
JDDNMWhK94Qby0oM+W8mt1Ms5DjfyThoxdurivaKSU4dIR6JO7cGeT/7TAvQtClp1ltnUHaetBO5
R21XjSkHsOcPZ6xpd42xQv35klDU+NHt5/uI6MYgsugpFQR0yOOYXzWeP9ghu9ORUb671XMeUwWs
MH1Chp2e1LhHqY/ZeVeLuiJlztc5OqVMBoFGfpPbqyhIJqd6/miiJlGWbGYFHTfI4912gufgRgWr
M13/urPZOr9vIhcB7DUzdXPbgzIjTT28VI9hrzeJ12zvqwWo83S/rOwz6AaJuuT8uvcvK65aiUa4
uo7tcQ8Pi3nt8WTzF+gploV87d8h2pkBVxoAWemQwSsmsGvZUGvQUZDWOY4DWZaXybM5RQCjB5oq
91TV1lMAhHklHr9EPQ658GF4G/ME1Lwt5mtkm7tr64THe7SvFHsEB/H6YM/G/oAzpsG3Yew3feRs
t+gaiHd3/jk1xlvbh47bBruGm2UJFF9XxI2Os/+R0UhSMnSF6O7YUjoz2pP7qLQaz5VmKfdrDeIK
naLbHh7yY22J/po+Dy9KDFriKp8MyYENY9EiNssVQennv/tqZwp0B3fSEqhF8OD9mEhUZoA5p+pP
ekMHi3ddkGIhanUanoGho/exWPrZ7LrE8wf4R8+IWghHewDXbFkCksNkEFW5bTvVT1Te8MPfjVrS
1TlA2wJ4JIfJsqGrWWASBw2QXFRtNbpGopPRHqfcMOPULV89FqU6qSTAh5Ckaz+soOeV+Vrv9NAo
ZEjZGauuREwv+rWsdDwLnwadb57KdiIguI53RNuJWFY58VIfv5bHxpCO0oqXWkkDHvXxFN+Z90kT
ku2iP7FUEst7INkeuC3d6YLJNMVY38dW3px2PggeHbFtiXMBOk2ZHIUe1Wfq8JX3fCkm9TwzEigj
b/r8gMSnVUSmmPtQkZWyuSiJfTtG1zq8takBLcBiOJlBVppx/+udjGUshXwAfjtbq/clxJSR61vr
7WA67czqDmC5hsoXvFjmmHhj4wcCokSFYa4NlpLD8uiohqtPuKpsvAM9dwSEj9jSU0iZ29scbj26
qRqVvhMtZNFCQEndX8GG5XVuuL8Us2EDkN+Iq+MHQqsy7HDj5H1v/rKZc3G+g20p5b5Xrm9C0l7a
BFjwEBksL8+vyVZeW9lTRW5zr3pJ0XgBVKsjG2RKbS/7FMJNawNvtrASyYUNH8HeZt+i6jFMHYoH
pPk/v7Px5wyc+IpgoBFLHUm7PixqWY8RGsa+gij8qQTP7+6sfzyV0CKsnXlmolLv/ZuWSyoSroGX
0RGkx9dkXxf5Q7nLzzmVlcO3uluLpwm0/vexPiZP/1paL7+YPV022bLzZGRToXItCoogBjrwYVoJ
4E9BRX6jlgVgYk2TnCrB+qoDCQ+Yencp4t0LdA653dkKi2fLnEsH2SYIudAFLKzGJHX99sTDS6D1
39Pps0E00ix4fex1IZbYLnUD/Zr4BUL0UOw8j1XZ5A6kwBaTpVFB9kV6aI3HhtW1sZ8mSsB+WoAJ
s2a6F7vNHgxlYQnv6yJnbPkIfIk8zFH0UkEv/sBfpg81UWXkriUCrrAI4d/BcOmNDRMqFZpwbwAp
YHUeEmzo3HV795Oa4JiOPNH7uf+HkPZqf134pyl0eu9IqTBUHqlGowuDDrbuLncSKm0YehgX3j1u
zqNBRc9Sv3US1AeF3zTocoSQVm3BvsDOBQzUNRa0eN2Sx5vAJWImfXrHBuvp9ErfET4SJ7UDkpWT
g0wmBw+iGMKYJt43VNEJ30qpb+euU8ystEM2Rc5+UOvMeAa4NXX+iCHUyB1SHwQmgZHNvu8p2ZCC
+ZSIRuDREuWeLYjuhVH5mtPAwtwDuVnkcK3JL1es0Ur/7SK6obBtjejskYJ4eyECvrrh0Yz95Xhe
z7xy6KtKm4QpT1XT/UbfFhGZIFIrW/bYPW33Q6ZQhXJirQ948q19E7tkg18yCob7Byxoy5uBtjHg
2Hbf0HKvXpraGMiBX+5Nwy+YUgY2zP0AkEaOTkSsCBIOOm66Bcr7t2UfTaq6Akh8ChWhfnKxm6Qh
7gNtLmlOLj/neUjDmkPW86sfRkYqq93EZ9WYhCJUP3NwKALzMc0zkr602q+55Lnv6m+ev80b6ncr
i6UQIVO7mm/4jPHnYayYVc5Kio65xHRN1RKnXStcUivGlKHOXon4Oif9TlhyWJACsNH4rVXqQxy1
EOxGbnb0/fbF12zNbd9wE3G+5hg9ALNuSZ/nkh2VDyRzLiz9I5iqyDNTLCKMsmKZgndsG5w5d2UC
GQqcGgUa6AYvWQA0EmMVPm8C6qzXOSxkWxF1PEQ65A5rqgcYGfFGl1St2koBtlcrMCn+2OwvMsWN
Dgs4vOyykNR+irXxKiqevSZTos0t++Mp+/8aMztAATu+p+oxcasZNqRH0YCpas6fpVkD4f/CFvJn
rdsjCSEamdLJLtnzaBI8XmUDRIjudOH0DTJxH9N3MFlwYkQl4JrUx39cuaA31+GydPSfe+pyYT8A
VnDBWEJKSb8+HOqtBIr/GNvkq7yaIwkJiMBrcXtFOtogflDqXzlDz3M8RvXKkvSqMakkZ6LzVl1I
nyvHOb4ZKK5rg3Yl+8KKI0o514tC7x28a/izDI6NY+t5xOiZUDkOc1FkS/voLD7GmVu+B7BlRqDb
anWfioyltXQNu9zcnu7b31rkrIMF9K+w1bxsFFVHt6uv1BHLuW9xqC0gKoBO/xy4b7BTuH0r97yg
kQXysKE7ptLz3EnsrzwUkGgack+SgBJ7u2gUqHdggxRQlnQk4qwcaEAG7iXeHyuosgD8en2laRfM
pXasiFCAjTAZTE/8Pw2Ya1aJJWn7aYv56T419d6crZi2LJH2yj9F9Vspk/bn4c3y8HGDhxRfgbX3
/LQIu/ryd84v/z9GKGC2ZY4510P7gbkom2aldrRmcwdRtPM/PxIJBNoaGewyzJ4JUt6Dih5+FbvY
JNuavcTBkrfLmFRcQjDfnCwDEe7Xh2TE9tQoAQpwqUkMZVHpfK3niTM1QhxK7LjcvuRxA5RHx8r+
pRbzMLTUfuOk3dB1A7zttslM6D5ktvqZzVxgABzbqQEbvUZfGRg2pXef5fmuTzDLzHMUy+hyXZ/F
GkIPxOJuPYSYAibWFnVIwAaK7hDq/hUfBXW2OyLVecxxypKCWBd+usxAiStTbJxj6ASMzSMNG3B4
aZqTpX3tJngUXpZ+9reO9COq7FpDUrLreAg3t8bRdAhnH5duLlBX36PRwzrlV0XEqAITzKVQR95p
mAPHjNJO5ZPwmkdpDx/gBo46K8WsJAz6BNXavDxKTxByXNmI3g+ngtuySfnHY+11tuzQ8s4uMU6q
pM+mWcM/b9UkLMSUVeQS/x5rCDHZgvTp5I6zriQt0/aDoFIwUTFRjsx5dtWDs+wlHW6mTrE9LE5s
yUeOzmnX1xk6Ro36s6DlIQXBYjRUfMd7DFwV7eoeMz+IlS37h4+bFBpdCyoXpOXo1azCIeyidOK5
SxEB6Hq0MQ6589ee0E3iM3L7NP4xyHRBuHrs0J94Zgta5lEHoKDAqS9eU99LgaQCdXCp6XadaMhC
w32Ic77svAz+W69SAszY8EYT3VivdCTuOOGZgUDdVug2Bg8Lfvh7/54VSZGHLUH+4B+n9Tv7Zs4l
yYBpY7crdBF1p8jnJJB60QbllN8aFUXVrG1FoD5SmgNBqbM2ewH49Ix1oPJIpPjeANecx16UX569
vdIec2haBIMF8bZYixo50qgsH1gL/aVuK01LiNvutRVwTqluE+CTz+RUwEZAEmflqihzi7TI+5zv
12rh5wipMTxHExve8kr/iv553ohYs/Mr/3E4TIxZpFup5KSazkyliFq508d7sgXuBfjqI+Bje88S
Iv/pj9uzoKHoDSPcjnJX97N6BRVhHBiNNReDms5JTNQkKvLwqRajdx2VaLm432+wD29bWEzAYwLA
lDY0mBgzjVOET0nYvLm/o1IgOcGn1n3yxdRnUqIiim0bQq+j3iUafnd8fGbadlMp7Pf2ft/y0xWY
GzqfFZ8gbeodVU97Hv4v24NzZlJjqIoGDRvhaQ2QAYuBO/p9A/x4cJ8w2MVRCY4DT6hlRtQDGZsV
6XYCI0MZAVseyrCnE+3ewtQGBlFhWxBJm6qyZAatzEC2pdCTyW3dRScnf01nRTl+HnJKFitZJMM1
fj+l0+EMkJI6nYkYY3aw+9lvs/NuJpSwW0KWQsZSrYUpVBNBMtJCXz720FGLeVg5q0bARh8FO+vw
ngMBA2ZMa4egb9HJ5htnehvGbYE/GC0fd16zvVKOnVYpQ6i2NfUAgaY/3aFmGVyyz1XCVc7NdFSv
9fGlMj3+jCMEtI0x3bkLVYSdvt+moln2yW/h4eFCO5I4Eo4UDKac2x9UQk/3Z0C0DAza53j60m4O
W+vdpdLyR3yGdn5XxjfKcz6F3plyWNbj3ckmO8+NzoUdIteeI0ZQdVYYIxW4IwDQyoM5f9304JlL
VM8HcEjntxuNITrQfC5jA72SomXM867GrL+LRo1ZJjYuqT3jk6D2XQtwFzUSEl31LVoiMUiJy+U9
vGxpUnhFn5vCO0Y58jJGH0/qBXAcaFycBChc3i2CR6jmj82EFVq5gE/iHQd9RynrTWvE/flhXncg
HrP5zytkJJFdwaoTHasC+Z49zNt0AG6Ri5e4fnmjtZQyhEBYl+gfNfPO+blP39B3oMzi320poun3
uBGarn7IpzGRDRSE9gkkb0aQJimi6vxsrRmDx654bN0/ug7iGTnifkvq7rYRlkqfHcDJVCVbfel1
UEp23LiQUNvVcbB+JsO3ZdNOigJWZG8UJlkos7zLbGReEPN0iWPffyyr4+T6KIC2MmJeZ0C4R+Ba
XYBFQVkPXdr0pi3rO4UaRqh1a93ncY3hkCmsqmNezoj8aDADuuezmTnhg6L2HywYyLXg4JjQZ7gT
zyCI5XRbOjtuhYVn9x+a3DF4SSCyZ6zvgZYm2vZ8YTUU+uAR8qBH+xyua1u1iAaB6W1d8eTrzx8h
b6Su7f0ZXhJJQ8iOWQ32M1l1FjQC/blWJeaydqdy5qenSseMtQtW/GKIMRURJWp9OqHk6SxI1wEg
kJrcFMS7rILI+WNpiZWi0bQZpRZbJIh2ez2b6r8qygd57fJbjB7ti5xwXeE7fs5pVVDUDflsTDJh
cz1xOdPSsrzednTADCkSceGSJFEWv/y7TR092KMSYE5M0aOe1PE6MEXE0DsFLehCZhsjqiVKz8zc
z5djJMK+7sOykX72b7eNwFEvstYl8yL/SoIbEY7DwdZUdFy938IflzVcGXXKS52e9vG1wJABBa/0
GHADqyahWyW25/L4CI2KCz0XnQISNJcnMWeWIhD10imVBd4JZmnJQpq1sISPS1+CNoaQNu8fpajw
dHI64/d661E4eu8VYNBWineFuQ5E50llUMT3OoNSe6r2/v3D8/DjjaH9vUxTnvTpmgWPrGH8YC8Y
EnVNoUzFQGvPxEFBQfC15bqZqP71oaat4IgU1y+QXvVCG/V1DIId8ygt5Z1et9mt/ETGqZOfYWrY
zLneTw2UBPHDdgkBXxGbm6A1303O0iscyHZIXjLkh7zS4gl0GfwzZ+4U8aHcIiObqC0gmAPmoKR6
k/MmGeJiZMn1OVdtYOcyi8zywwWhMsf4uaBXfLNOUb2t/ZTLnOTjsjZnezKqn42WkpWNOBlZJbCR
RTar9Aexn78Ku+hiG6euMVozpze+9HB+uUYrliSQxdbnS1KO2ffQpX/mPgWEXzwK4nU5tBpo6aVN
Yg055v/wFJ5M4zZHXC+YPa8+P14XCDr1hHHFzBh8iGQ66LqkNWlOiq6hEwXbzcYzR00DXJTkfuvu
BNdaiHABqlV1QKqhGONj/n161gD7SY8puukLya+A/JEOKRU1i2AcdSB8K/su7EarMs/vJqw3AAXb
O0nbJ24+FcR4jc7D876OysrvZ7ZuMbbe9Rg1Bd8sq6kTwe8KvQKO+gx+vTLi7s/8D/925Kh8RCJp
gno8ifuY5CdyhJ1KWSFgX3eg/1Q972zJygXMBAqbK5sC02/3PY3kjLaqIDnE7nD+o4HPGwAnEHN5
CTTt52Ckfv4BECYwlTtuzHdsjNDgX+ESoF5ZH9VsI5/5jBTj2+iBxTJS8b2ifAEplN23Dr8gc+RJ
B4ypZUQ/dulD68+sTbj/Q/SQwyn9QgFBB9T9I118vHDPP4L9iNDZ1g57GTzXagX8nn1ZFWCmPH7l
OWfVzmDFp9+Knoz//dqrFlYMH5JFCe4dEr/2ZhfXiE/v7aUibFjNi1odwM8ZHdE42TyA3K62LyPh
FGztK1c80JxvBP4q+FmPCOIRFK19KtD1Ze9+pHqd2B1txvBkogIfmtxGjmqd/oxsssuj6OaWp0n2
bhfWAVaNALcki5Z9Y8qp150RBcCnE7WCjBQBecRO2O4FdJv7Fk8fRz7QcSOXC+Dtb0T6W6aAtDlQ
ezflekCu/ZQtw8JtnnMYnh33+T+CrFbdTwRSwZ/jqHzjSB/TYJjgM69l31NF5c+d7nKE9LaEG+88
2ycuUe6c4xrhCKIy9uvc7iYZQY9q7a/JPkMyd6QqWR0SeFJBs2ZpBSCZdg8QUBDrBD9isbgZjWhg
NGFMVCFvSrzTd99VdBcpSFwsGFipQbDUbOD0Vphc0Grn3ekCKxs6a3CwRheYm42LHCKKejzEQHCF
loO3oip90mplTOIdQjSe4LEOxOk3Vcf0KYZ683J1HNFzIypLEnR2h73aKTt5KKDcmpY9XajePC1S
GtH7w/6VXSLXQT6imkpFrri4b99EZRNQ2Y42JCAYpDU04QKIW0JskWpsAfxTcPKRiJHmmPRJbgM5
msMp9I9kj0fee/agsoPJMrtkurEyXvJgymEOqOxDDYB99ysY0myjCqDz2Xcs2mtiAUb1sVsFo1J8
tICqp4aY5ITFn6FNJ556KtDftSkfViaCb76D4TqQLnIk8ohKjPDVlJeJBxadtxVsrNi707GNGnDn
p0qP7UwnQKEX2HC6ntb8z5ycv/JOoRK9DAuQJnQQNAL0N6elXEi6+nrzHdcoWQ/CjOsIjXHzEoVY
RWCeF52TR9W7biUYS0g9pVT5tM79GrBdKlMgtWC/2Nc9DalG7rVPrd04QW5YiCn+6PGXDy9AZnXy
0dxAD4W6i652tM+r1gXU6WOrT4HdWh7TWgsN9Iwfedg91iywfN4CLA3J6HBtFhUMlMV//VPT6C6b
pRcZWfLx/kClJGO3ViHEOh+zu01RB0ja8q+OZO01+GNVmNUvdLwGTwL3mXZXz0VlbxphLYmuW7lz
khUAYjB6CO45zGR/2IsNput89MklifjP5u2HsLwDAEJhpKAFuzH6H+kA7rAZTL0flBVui1fQGtcN
1tHfmtWikTo6Z0x56SstTUrCXYK1G2dYYgD/bEy28ouGtVnTEMilOJaXGXkJkMLzmhMXymTchEXd
37MDFLe25tdo+oALBvxxNwxdWkoooHXd3R5kTsQFx4kyCmjGgDjt+VB5rhvbhzykGCnuz+EAth9z
t0ZJrhxOZSktceKr+ZtjLTbvzKRp8kwnA7VSoxv+wFSIXd8oRzDd5tjVMxs6txbHSUmz9ulG2JSr
LrerAQf+Z3SxIrgK2DiLuHmi3rAQxpBI5MBWD1IdiiA0U2h3rDI8VirnLl92QhAG/B3CV1bBNoNl
M6kW1hVlb7tIofbdLaUlp2ZPtZQX6D1n/QkMCoKQ90fKv+YtpyE8vOX32V60bq3PvGJjpxjKPLQd
rJm3gW15wjVirUfy2KJwzXrGLNcx2gj3ktp24KgbXUiaRY6m8QuohqO7I7coUtUwfmFDbxyiwJyQ
Cdn6E10mlAxiXQDchaV9dzpoSAk5n/H0PrWAiOQvZZ4v518Sg8aOy/z98lAh3BGGkPEIaE2T/jRM
diUOnpDHBavjg2Kb9kU3wu1Y6pUWfIG5ZWqWyAbv+tWmXCm+czwl+KKNHG/mg5AXQ8Q56qcE2Mdd
KcZAACzy2GymIDTm7AClvyn2q1hbm4TB5iA+bV9ET0Y9IdduDm6L23K8vXAwYqdHmDpGIhg9PW3T
jRd4jp5xbcnd7aANrL08IRNFH670uBgIMgDdcUTAakV358jv4miSNPALy6rZ+lOvf88k7rWCbXzu
thtvbDByg2rn/hIVDUYWLsHdZ4xa1n3yTWYG32S1J9wZ3hoaObo6oXkrcIrWkB0r9ybbtCiFgFUf
ZNJWqtqZaTjhG/FZ+U1biC+s2NujxaoYjAT2b4zapJ6xzdC7Flb8Yekfpboy6uyCA9Lak9X9VP6l
BBuRKBOhGsmnlbUNMeSf2yk4oyYYzVirqry6CCKzETiynVT9w4/FxSriPKVfUJjC9+e1Wxjq2NQz
ZRHybtVWpzr0kEZLeSh//6FZ+hOJKiKovqv6OFZISpHYsXS34T0WlM3Z2mzvodoMcAlfbhMtIPsw
qd+D/703Q+pYWM8dtWq03SWTONkVPgeotTEQBMs5RtdPjExiCK/wbpNC7eHZeoG6c9BTSLojqWGj
Od9U0RZG7Q2l5ZSfECgrz+7aiuo5E8VGm3m7519wl5YyAbL/RPMa53dXO4X1/y6T4iPQcC5n21JG
QSioYxSnrSLwBIlaU3ePPtIbBGeDpaI2B+EqUSL30OK0WUa/RUnbGjmZNLzdxRd9sL+NhrZjQoM3
3J3OVvGDiIlR2ssqoZTtvYQVtRKLjjsroSvnIbyelumRagmZl43K08AwxR5a2nIEIEpSlVE2W5C3
ZSjMntDmEADhrIiF2zuUxsi7ULCj8skAmRNEVrEpjQtTgCaxT70qL92EaVHmaki1HufiAjUfjfv9
ksudinCoTBkS2Kzaz1qwYF0h3Cjt5yHJYpMuGJvE86cxuzZiytH6+U3RD7h5FV10xIGlOM0NhiYJ
wCFEAs0iHuE7OUTpf3GblFSuIxY84FoBJYw1RP4uElyiLY2ijv0gslxbKbHMAQbkDlQspdZ8t0QH
uAZooNSjfEflTK9SKFeHBcVFAiJHZuxjFk4l/JJVqpEPVDc5eWqOpsfimsB0S3W0f3NN4bw6wyg4
zchqBtbWwWL115/nVzXE00MunOif/ye+TH9sq8AvvAPG3yeNkhhNfI5vz0AmzW6TKAFdRoJ1iydE
7ffMHmD8b92bqOPcdCeRsZsmKAdfFCInQyr971JS0dsgYRqc1d528hOsom57xI3BqHEbaogXlQmA
+cgYd5f1D+BM/d1HUlWyD9VwhMjxgswGyzcHtvZu6HdqRVW87bS19lDwFUpcYR0tjxgngptP/s9s
h+aciURNqb0wt9G7TGc+/NUC6rIQLAERZVw0KunQe9G/5Cb1mJK1h5v/M1V83LCk1BWiiFo/tg2T
l8AtF/qsPFFR3I095w/dMPgLdZtxB9inLY6ps9IFymkTjxKe+MEBruUnI/zhBBOFy0TpFBNgFdGR
2y33o5fsEl45alUpuTzy0LKJN6l3ihkbTL2ZKRlHuNi3MLfieiNPkAs/lmcaDD890dhnYOib2PHp
oQQupc+3AfwOJW6ZXC0wpEJF11dOYYzV8OsZuK/j2AdVWLxc5OgZwm483vZhG4jRMnOq7pv5/4da
hU2qYis5+aeJj+r0HN+vwcys/rlek6BZv1QHxCXJduDkehOg1fOpd1UZPlUS4aqniXEZC8MvAtTz
zGj7RacmxqBnjTcB4apuESDjijvtfGdW+Hu/V3v0fOYiPJ04THDeTuxXw7QeziQLZeKdVI3c6I6Q
U0l0eaPUxUFdEMfW5OhijqARfasxQllEB9+sqvCGMkUpkJ+bxgUomvQrFcT0c/TI9iDQItTwjV/j
t47tO6fYFDlmlmPn9sBc7WC2VnJ7N/q25+8EHqKcY6qap7e9EWGiYM/bAmPpWNQGiEvSEi42fk24
48ASgePiGZKuIEtb2I5X4LuF1GJg+qWsw2hgrhrZIw9W3e+uFnyTZctiSc4tawuI3dtzlMBESgw8
qYw8GzEybJMh4x/hh3S/clBj+yeG2xjBSnaxJOLj8TFE5OgY9wQC8w5BKfoqtAoLVMMCL+bbKi8m
+lKZw3cj0EBLs4REzzuh5tPWtKFsESxOKZD2P20wgOyXWyJGe1Dr5T2hU7hIxT/MWAbOoG2iYBEn
lONtWQifKKSk+TNSEY2VukNMl1wtBiUhSS23DG3MH29HcJUl9vkjeT4wbvo3qZ9Hayfqz/y8aFwt
Ot4V6DE1gR5CDOpmZFYb9N03WRtx126xAO7CTlU9JHzp7FmmjEl55c/kxtk6Ly/R0knkNcKpQV0t
irJkANNZ1ypO3fjjgFVtamnw6M8d3x4KqySWKEds57Xen2C60J2EN+xshoGmqOlocBEb2yTBlu4x
OWoZkCTCDUFhgxl3I0mkfiwqWgeM84AtSaVVRBKdVVjc6th6bPE3XslhxCBMjVZy3/YrA+dS4pAd
MR2e/vf7nhWGbcmN6bOBto+NCxVk3+0exjHeNw5WBmZYZLrCdpucVo8piKc4o0YTrBbY+ouZv2ps
RHEmamj0yVi20th1QjYgDpV1pms/KvgQhdPBi8Bir8NO/I4tnM+ELtL2McN2pPoRjQ4IZphETRFf
4r+J4JmwTPUKd6a7X0RYwtogocjPlbGmxf7j9W2yjK1YLvd5lzGmNsu5nwpjC0sqdO8MAtfG2RZS
X3YWrGr64s7AuQ2ZD1r4va7OH5O2aKFc3C0M5IRD5Er3Eqy3EGwxiRiocnydkRX3amssXbR7k1sY
bAlreZsHAq6c99vqJ1RzPEv1mZJ/+ty06YKer/MDNvkBslGQ1qkFgfCqVxduNKoG2dSoQmG9pQRP
LC84s5p3/lpowL2ApRzgs10xEivP0Ud87IZIeZjpR//65wEwA08QZRN/nkqEVGfEU6rcV4D7Dw+G
oFFWd/lo9E7KCrT0jsjxcj5YRU9MQXr4pdQIvt1AzD0BFKmaH+QiLhmgyscX1HE/CPvpNh9X2AZy
jpvfFc7OgSkaGb98uhYXTRGwDAz/2sBc3izUWQI6h5LKg509uJQ44/jte301hSqKnw9wYeFrYSzb
WGD/oryEctXGMWjloWd8fqbJadm78muVGZtOzWjHyrs8XJ6NzXrEmz1oPGKeZbXMvQEo7MCXpgTI
QsMvQlCR+gK2oedHaXQ4IxM6S0a/zAIEHID2UbNN+ikOu6CUdzzNwE0avG0tBeQHys11Nq6+ebGb
VTbdJBpPgbKrCC5VEG4t7mykxSZo3UCkLAgPRKmjVvDnQD87afGt7lh8ZGh/EbziIfcNuh9vN3+n
kHrmVwIKaqJ92cwedKgochLXuZUpqdxiY8fdE0qFn7K1FrhMOYROrgf8UCrQot0dKrr7YQ2NO5cP
/ArtnKNw1Gg21n9QQEW8Go78D7z1D60dUoE5kFuksghQjlusuSJx3TUCfYYNC+qIOXPdYgGjSEZA
1jFJuFcMYTrMDlZVwX/9dh2G4U2lvMJ/N7snwjoOCuBkDQmTFRx13rju1zeNfI4Vk/hYDqFjZ5Ri
6OLQeE8vLKoI4dGAz8gebBYHNLqfhsqUFvq3zHxHtGDXQHI4HHTexZFvAmjIMS+XWPtrwohVj9Cb
r0o9yiWC1MD+8cezkdr2lwNAKrCu+VI8pUQSX9e2fjYIEozO2sbyzzMxRBv6KIUj8J3rWn7DWv8r
myWasu7RIznRgJ65+uO8ANmpFFbXoZOWjMCjrVT9swHW18CAEhFoTp4e4eTMJElii0vPLpZF6Pfn
Y1SW1O+Ml0Mk/PXJLckpUB70LeztYhKyXvS1eFxlhK6R22LQk3NdKA9nL9bbRXFAW6z8AuL1/Q/D
ZYCrSa2S4/z4I6q25kSHJ8q4gYy0SS8FfsOPJMS6DpY8e2YEwsAH5sPgPItDWEQmnKX4XEuTGjjD
vhe9e0+pC2cPOMOkC9eeXB5ERIFk0PL6JKRt5yUeGXFqLK7jxKDs2j9qIscuuBfPtOXd44N0onSU
DHxWhak313GuCyG3sSNSGrrO3Ikxh5jgzozT/MQprgWpUTkukJvP7zbvrS6vgbRPGhSAS/Abd6tR
EhW9v2tiqnOLz628TOoMJAWsMVva/9f0V/RGX6qe5tryUBpjggl7laP8490n5co/XMTh/0PewoxO
JP3D9IzmKGB6qU9kWCq+2sLhvGdhqKBeIpMpzOtexKwbJJG1swmjI1xAwa2rbPlfCtSDsBvAdjxV
Wf2qQRVd47lZCtJ0mZcoRON3mkl9SRA0S8EdLdbHNU2qu7vR+n9rZS4LYVKhgSyVnVc8YlVigj7s
bCi8G1O4HdG4HnX8iWTIWxEq3C8e0i4Kaz5o+nJO7YNdF1Qu2xbYdX6sK3Rae6UXXVcgs2WaHTd7
DRpnhHdflHWb7K+qeH5raGQUYGyMqpRw+dqoKCmjWRHgUh+DLYhXpKeiDumUD75AS7yFRLjk7Uj/
7tEnHLsT+4GoQ5sOK9E80o36QT8vIqjh5pqsLWX0Vipf2w3RU0dMDX3yNWWzqjX/CDgzbrZPZZS3
myfauUWFkxxKwbAyXyIz9VXAFGiUuTWtAkOEiHhs1kvThBqu/ShfLDK/jpnbO8Et+djqxbu9PjwP
PXadBE8RWVuSiYrat0syr4zGuJVVbPv9/RfNZkijVtTP/f73zXu1gqyZlrdal7humiuewBqdG7ip
ZhL8t1cb+xc/TfBtKjYMRp3zYpC+JCfc8ToryZ1PvEO99ZdTyaoVn9gpmYJMH67mMW46dtItwrQX
VJR9HoT3jQGnNaKGxuJA4hJ0/FEZuwmRkosfj9/39eRATw1dXcW+EukZQZZ5Up9xt9p6FTF8+5Ap
9iED6NLa0ijWb5mtIQ+bFZb0Js9IVB/fm9aIlygN6v81i0kXNq/xqkYrMSCYhj2IrldVQzUcR2qa
Syq3NJ4S7uRL0IT5f+MTW4ulNmqAir3VzthinTKA4SmNhnwOjP3d3vERyr4TzNPGBr7YCWJxDpnt
LClhR1jG77oUnmilxwC7XHLS7dJJhR3EFFo+l2IyfLrqrrQFKsoFhqXEEHPe5ql9WEPjahgT8Egi
r5DenQhHFIScuxNO064lSXYWwqAfKK2DMoQwU2F3XFxBHk5xCgYkN/MVIVSvv74c9up9OretJH7s
ncMgg7nzQWWilfkhLLMa5DGCDcDOgZjOdEzYrzXeKobgQxDDE8iB3mXNVEDuD8EqmL2sl8ex2bKo
xOiZQD++mxtJ91fyhmFtKBEzY3PZbMI+sLSOI7rKGAXCCOJa6pNsDDgAIgsO6w7AVHmPQrEnkj0u
sn+AyifGGEwm8/l48UNCNk5dBGdg0FzP+T0rSUfsDHC0NmcRzrpjqIMaJuD7PoXh9r21CJJZvdVa
+28LdGo2yLdNgIJiIkC9F9aMFbqi6MFDUvb3zi0rwEVYfkL/JcRjp6uxEeExXgG2IPPNquzp6XXv
2UnOizFtqX+blRTrZRHges27/yZ5+7+USzTy2XRLBnhu24nTQjK1E2tCiRd3sG582Tz5jQo4yE2f
dGKwYYLwUbAt9bX+eUPMTykVcW6XG2hV8iIkSyx3PNcwaFey/VndQV2Jg2rAq8hKX/uJFyOMw4Zm
JKPMLcHuWLROtpAnU5/7367LHLHXwVfbDpwoO4L4Xb5YauM4oETmmWv79BeFZE/UfptILMTcxc+x
4pGuN27mmUm9n05Xdx6QAyujbvs9jygVi4Xbofg7uOKnxtDoB5cfI7N20IL+Qbx5eU2FsNO0gcHl
X/6Po7ezlDow763YNR5rlKBXoKYBMgYF9sIKpuG/WJYiMcMC2TBUEkrfSlTPBfLJINrex/TIokc3
b/dGoHA+XV+LGKvULSDD8+f27okM9qSEmMQlxt6BgONR/IjO9hFZKP9zvXwPmbXu5Nakz5ZjMYMV
Arqj95fDqprGFPbqGeHUlGLauHtrzfTLUsc+R2trwsgjeMbJ0DUmMDIckGOhj/VeddbQFiELkFj7
CFKSZeNQgdAZLSawFu0RUPIYkKOuTJJB04s5VuuP5PuTkPoDNd6ZukUHFqBa9I8rmbAmXuPsy/gM
z+HkfUF0XrQRDqJK7loQSrgoYabw8ssZ0D3PF3ibS+ce9urGaNn6DCK4ZFH3Ta5VaFta3a7E7gLt
9RYv4t3wuhvljk1uxUIK2/Mqpzf0CXK99+q8amZYONApJYttqny2qNx7Ip56IshrHYv8+8PM7Z8q
3NBDURZTGKDucuEclFIaHIhOF0KmxMmq3lgheDBgEi7SzurIu0LM1/n2/Jorc+8n8pxf7jX7UGaX
o4/lAXLfIRye9ll4jQ0mLbOLzKLjmEvwxZwBAG7hNU5ojF/w+Yvio2jf92W3DkCbO0sT/QaBgwfR
uVF7fHsQ9sZP/bfNTuak3geMKbY/euCc6rmTEibSWTwyX85upQh/JznTse3mHhW9LSAZsMeo3ID6
G5orsYWmwwzykqEZlnCjv+mLwUHT3jJzEkIKgu3NsDKBiwc+XpURkp3z4Q31pvWeeNePxfrj/j9O
jx7769eix7O7dCaG6yAaX3II1UX6DRB0liQI+sh6vbkaH2FnjoaGCTF1F561HOUmdAUQe8pAPBuy
7wuAAhN7mV7TfmX5juU+HrVd9rFIOa1zWH/lnSb7YLy8FVw0CV0FFOSkFvwiat1KhX3bZ5NFLTSv
zdGeQnHp8lc/I9RKsH7IfFaWD5gXvwUGCcX6A/Ir3Zjyrzq4mRqMd1dMwJHMQe8AkkNlPNxrEZ2z
nrk7uuJRWTlWMB2R76f9avSMVaIYEWIJZ9Lm7+VD+S3s/UZOahWvBvn52ATzCGEgIBEozFy6J9G3
RWMnJ9ozeVNH2KXQI+WE9BqDYQl61FzR/pQW8ejrCDV2VtgqqXalApPnxlp3/92SQ0Z6CPN+X2TX
wifmvrXcY4Yi7oh+DhITAD8xGUpAoZxwSlSYR02EmsY3U2s0is9pEiTE6tZUzO/AlR4OalsW3uOu
1s3ZYKDY/Btzwwfd2lPyVgXoLN6vAhKPUDVU8JEKVPfMZAzcuDlrEPyHXWuWpxJhf6n4UNV2vYzH
6hrZUxslJDydZnksGHRN7YkYAUP/rHvkQ2e/fHaOOQe/pNfzEzbW6Xn5UePHD1PBRXtbTTv17c0p
Rk3GlO4I2sGbxotODxaF+XhQfU//tSywxPmKtwOM/kIDuapG3RpUkn85Hr8dNQ541lZe8pxdMp5o
il1Jx1CEHp5j1pZRU5Bhv0tIhS6cuhlDoaykuwoJ2g2eiBUzZoRbZxM0WRpRLScBx3+zDz9pbuIT
Q8gbZawS2b8JhdEcKG+NRDLTNmBZuuLds8syh42PO0GiZYvPSVLfprLzigFYg+EUKSnVN03CvFlR
vbxt/622zc2mQgIMgaB9I1VNTmDOGSCBFRKqxWoKsWFBoPFCmejgjgXPCj4G/xz5rikPubZ0MAPe
GgiSn3xXXZT7h7klHE3wSusnPRkUzkfVZOnr/aEuJVVKJVT9U9w5dGcPvznPPiLZ+wMbGGA8vAIU
mRwx73ob3R9vaINYq2iKVDubkZSJJaJ92fKuAp/PTpjkCqnZRBkDGd2n7jC1A0U4BtSs2sI1+CL/
txY579LL82+ks9TQO9mU4F/OisXm1zkUYgYOzINwAkQlBf1lD3z9ASfa/u7GlEtv8NNVClSKTKPL
NXxUtF0UU+GNFPEVyQ5x5FiwqMX6PjBDfbbJiep0AWnrlMN8/kpVa80ucig70mCcfz1Kj1n6OPpV
9G2R1OULDaA193FMQICXHH2HcHPag+VVmWKOA3igKPdCuCtbKWhJxW42v2hMkp+vLluB5YdBY4Pd
J3Q2hBFRRKWBNqiRScp7c+Vv1+AtsBc0Z+PhXbucfZ3cMhRHV7haxk8RRd2DmzAI1fHNptvraNVb
ES1C1aMtpa4ZNqzoM5gh6UHlh7kLgU0C2HCG77k7sL3p4a8awgAVhtETdb0V9NO1HTFpt0XBngaK
9Vs/0DEwVkti2mGUcgHhRqEFaWpg83vDjZnjgWDZNbIeP8iQYs6+I9HMFqMpzSb+ojG2jr9Tqmgn
nttfMEj4BVzincrrZaQ+Mf0pDeh0RHv2cMucXWbamYJe98oU9dJCI7/Ogy8As+C7cEmZ5+g4LcM1
UpOszT/AU0XeOd1TGJQ3LD8Rfm91pKr8XlYB6MEkm81ZqVFeIlBwbF5q4f+QRS9+ScQ1AD/9zSuJ
Z+paU3tW/OKp3vjJk26OGBdfsVNgfyg0pOxDKCsxQ8rBPYkmRPJ/ATKfaB2KwCtEW5myBd3MyZ4a
dci06QdjPPFqVDckmpWOkCG807BxAG2ankn4zogiqmMM2S3jxgLiFHdkntYW6SlSJYlN34OT2TRv
KAbSwfN8r03epKIFbjcyMovpe6YtVMPPwUEnWcHI9JwOyone5nF/tcWi9pKIsIPOARrulPYnPzaG
gYUbS5/Ji5WuCoW9h6zH+MxqBNBsnTQ1sM95OhgScwK0snRD/o112UbKS/evJEQ3QSkRei+5CmdF
zZ7LI6hmaXmbY+mouL8npVe7BqerAFlACl6NjJh4yzbDpu9xDimBxe9TWQaY/VR5M123Xj7X/Q7v
og19ECCx9C0CNJf+6z+3BQz1J7qohaJGVUDQ7hNvOHdS5Z3UDtQi+6qN17eshUypLRYHOVhraJXw
pLRZL96oE7jBl0A9xfdBJ8LOgVTFnMx6+qXnWVD3IZr5IOKWpFhCoZgBBAqxXYscIk/vqHbZrubQ
MvtdURurzCJTU2DpPZB5waPfWNs3iMxOVRkPmOB40H6dfFljsKVYWmfzLuDBmUk6OhgxjzCrcaTx
gKEeXNcVXJBuQtiX9Wbq1N4hPGWAPV7SzY6Qzh7lw2UgAbDg45yLT7mLm6+RIX/MPd567KhRJBd/
cn3TmfYJ1KSMKRMzbQEv8NIyMecZ3pBqMkxP6deQXsKtH8OcQ3xxBU/hwhCB9C2uE7u/gqOOQf+c
lW1hOu0uHmasekYcjmAl/aqBLGBUWawr2XUqy/wgwpmqc2S+PkBB7OflCJEKk63OJF9lhM5CXyeI
m4o7so4GHMXvMN502QHikn/4y6HFReRfZmQ1F7sG6VVtvWxUnLCRripNtTcHWQoMOe4Dw5I3NAdE
FrF4FZvUa5E53ANZNgZqhwKU8i92rFfsn0fJ/2BvzK71ioOIZqdd3TpRbdvv8CHQxK4V6WqoaQnq
duZHuXl5guiSoe9mTCHLSki5UCojUk363dXJU2eYu91K7V6BwtSNPjySMtJcE75DfIRxGkyAyak8
dwCrki1wk5kZCprDPQ9r3+EZsGWdw3dWOm5f1NCC7c1qMqQAGQdIbTj5HtWSxwqr8PG0G76SN02b
9738eozaeByT+++zAa4kriX5AO1EuTrIm0W/VzrmRFTZmluDf6ZejJe3YfYieuYepL+T/RwA1+VH
O4Yw0bBzuCPg63+yuYRoj9CVzbz6B6K8ObZca9tZaXRb5IixsBjmBsSlGTAtS5zdQCvx6hgFOLlA
FomoHyXsBQJSWLPzO9l77FsSxSyHAL5PewCbIk3yDnDgDljI5nlD7W1/B1jynJp2Mh1GerMvgEAG
I6oLGWokwhxl0rLgs72gaXljiIYdKiuAFoqDTCAadflOLguySBYY4WjrryQx+RfZJ214daQ4WkyA
dqvt3yzwmP2Xay8v1J2jLQc120bGZYthjJ/lQR5X/qMo0EO0Ud98S889XAM38eRKFKvYUiNyL2kk
4aZHqjw07G8zl9MaMK++f4v9JnhJaKsmdL/FGCJhCUmvQlJ9s/tCYlzHl2JBtIAZF0qIsGrv/1zh
stsuTTENXS0JleGrS1kTcC7djCsKkkr7ZdDs916H8EGHwKro3GlvA5ZrlH6o30pJvd2AufkvTz0g
o6FBD/5Ptz2OyyIoWxFVA0Zy5vjnDD89owN1rZlhruYgADD23nSz9Xd67TNE0zAMzdq2v/Toq9WX
rpqAzb8m40c/6mgMdi8qjmGh18amIHcrph+Ej2A1M9hourec3aOKSNyZjocdCOTQJmv6Mp3v+SLA
FZvKNkOTXVEcC/Swes2eGh87TMJy4jQdxbl+omzrGq4BU4GjBbZ/OUWD6CBqfWnNtzxufWFMTZY7
xaTOBtPLxvjTFqh10v5CyNS6yDusv97l7jOWWedcH7cWYBcppohEJRHp+lpnaWfrH35um6+OOWm/
rsnZDuFBpiYxjo/TOEbCaLM2Q45reKsVygCtdZbIgJsaUiHtf5rp61gXuZrfFQIIDqrJvyLywS8r
tTKBv63Od6BP1onQuXNREEQMEXq78OWNAyyqEsmXBLjBkK+o1rsDN0/0eyMWGwTdxxYaQaQvCSVC
dP13u6ktFDHjO9KkVGyb9Bc9d/EAl2OQ8RSPJDv/obgfj4NyYju9mZAsZJaXZi+MwqO4pn++Odwu
DZv+5/a1RE1WhYU7s+8/pnapjuyRjWbq3OTkicfOy5cXNC8ix2iHwBC6K43JGZGUyVwvDf37sVya
AJPWe7XT4LPJCMbIcUUdYKDRIi8NUkSiKxAeuadqSCYiGfYtSIoZ9Amd6U9DuUdtPlJ8RrjIO7Fc
quywbMhO5fMLnA+1gmewhO9YCyrG9LvMuAQsxbMq5FJr+E52knBDP7tYzMS26c4rhYbQBJ8nBZTp
1J12VP/76p25YBG1ovjT5zlGfXTQeGIoFa2OWq0dSET9y6LWhB2UFkCv9dySlh7mGU8E1uNmMMcg
Re13lZ9mVcAM6dk013ytU93SUIQQGjuO6srX1bAoQZ4JeLrtkj2pYrJrWkVeWtI7ZSYaJoQUHPPo
DPg0uirCDokfkzmoXJE0QeDPUxdddDFnMTRMaVgcw+poZ0sFWecO1dXkIN6quQJW53nVJvjJjhJx
rMDYk6FQyjYa+Yor78KPi8CYiDnsKXDk+oL+5fCQyz8Sr5jEv0L5bbZuZlQsK8W4qVr+42Bc7qnr
FUN4UScC6bWX7IWZVYJHF4Mj16Zz6FRthihY4qCIK7vyzAAOcXfuAUmRcAKM1Gnm0RvflqNAjEKq
6DKcdwTz60G9veuIyzJj6xu2nBUJ6puVHWCkrQVuLoN6xH22pPHMxPqn6e3/+SRauT38mnfBlX1a
Sx4J5/2t18W6vSe+A25BHPXgbQh4plLPyRlADHv/wBTtWVjJTXLj9S2V8RmvvlRam4xVWfgMv2R/
u4JZ0TC7gGkCeND4r4d5QOabUVYNytbeChsVtotxE4GbxB6Doi/8cDeHL/klJpHX1cEAcKB4fds4
omI66ikbDfvbwu0+ofChN6mMSapTfd9uJc0DAuULTR5QPNEoDoDoUWuad5TNjIzqhG6HvxK1oBpm
rSHeBaK1ntJPi4kBMDc8OD/kxy2YBNis0eTy53og+727UkXjW4NAxtdv73UG7t85OKxnryu+hQrG
DhhlVoewujfYzkOyDe3UMDhgICrk6DXB3mlvn/aNkWioPWvZ6Ay58Y4puMB2hgFisV5+YN3sqPna
pA4WSO43Lzf/7Ct33F1f3cVH5hXLILtmE5krrKd1Oxmd8QjyxrTwESVTXmVtlmQodqskCOMdD9lA
MBOhde+rSNY3Vt8ryPrYeSXVJK5VYcZj4+EL7og12YU4GGmkgB8lGm63EKt6ecYwmxck/1envX/0
4mbJPoGahwm4IWMKaHHKm5+2jus8HU1f4cxBcVmZeRu9aux8Q1OnlyPgnKv7050p5LAXSBj3+xGc
YP3cAVMa0BeoXmnj1ogDj77VR528yo55nLHef5cdkqMb/PAlEsYsYxB+MaZCVkEhp/mmZcgGe/2Y
VH1q7hEeUdEkXb+zZqeb4AN5tWtYU6vqBGTOOzOMElrIPJH4R1XG77us/vp4uaNljP7bIGp81Irt
4rI738iCzzLIBqzi0zB2plDqgFleajoOhdXTBGB9l/KSaRQ1E8chL2g9WQ6gASCeoFORXDlt+mfK
vKwh98ooPkGs7Lo2OLmvIiZjEZCALYjCdOLa9hcpHxLkGFDoETSrzc7rRMUVf1ygBAEwVuuXjvpn
wwxwja4C/PY2yAxjSkXXHTzlZiIkHfybg7ab5PFaf65Pis/qa4huKrUZ4L1aYQ2vG0/qhdrGx8W5
U4LL8QAGdvWIhb0TmIZOTNDCtS0mBrzYaFYjmluP5k7ENC3rDb68oZiMnk53ddfV0f6MzHbRifX7
GJd1cKN2haxlqFyZwseHyTmgb7ctuC1qi3Toy28UvCABwEmV8Q44pHvuhPRxKBpkF6OJTSHfXRqS
NWSGuhagoPyWq69X6jFCphQ6HK6SeM7WK58PtLiGBTzAXsUHItnvXuTHuClD0WHQy/qBh0aQQYBU
K1cmE8Vsr49LcjfvedXzXPSxIirvQCRlkXK+fJR5Zhk0mTI6OrIckdq1Q1i1D35AoEqMMToRbdO0
NliPsR/jUgdJvIweQTLtA0jadIu0A4UCa9j1YChkvW5PkpDDFeKUIlthIk5H/mxUamZbMRWCrGjh
CV7lO8zvB7dRs1DwDInggtoCKJuiY8AeS0hh20zoUk6ArHYOsUsyksS5thOBXse8muMzqpwNiwY4
oWhNs2vgR99Mjwn/RsLfv0/2ksZ/AuaAaysGWl+NIRmRBlzQIn3F8/ZQz8zKQb2dNNsiCarvI57P
KbayMC9eKOl4mkBpVkSBwe+gta/1ghx/OXMpkvPJWBm68cnCwjTmGCIawcMdhQ2UqQrqVi6YklIO
Rn6/VoHvbIxCGNEC+kqGnW5BNR+wZb9UeSQas5e6SexYGyoLQgtC7CMApQEQCaIewAA+yuLS+pQk
kriIazcNSDtlfbWgE8WAnA52XH92Pg07Dq/dBu0yozbRsfZUL7R1Tnk1hGSSBz2ZRjHwYp7s8Xg+
khHZ8Rqwvdb84+ErEcBHlL6wGIXvOsw9U3z5Ll+sC7cYLD9W1+tmXIXzxaOm065E+Dr6sNnhmc4u
H9Aq26pAK+h5oG3DkDttgljohZoQleLetENZ5LILxB7L+7RdFYsjS8dDQXwu0rtzGbKuPDlBSBwx
hLaiL1+oRhqvDDAjelSPbT77yXGDi3aC18uaS7BtcPhdaEzJEHavBKwIK3aVoe/19hgDZJZ5ER2D
Ys/qpNvOsxGpGsW+HxQ970f1jKO7t5aUkDu21DtetIi4sTdm5znr8ywDHmfB+0Vo7nwBlP3V4rJR
Wc/hnJ5qQnLwOGEFX8EOxVhrivzC4TbfMIX6Yf+CBTdIvs97QSnXl/X1+3OAujPpI7R/UknkBK2y
F6BQ4C4zSSzZXAPVI1TDuwUd2nJ2n1loe5HsdVy3lgP2PQ6iHkms9DmfsTXn5CNHSsyXM2587dt7
C7AAA04okX8dlYM1G0Ka8G7ykyNKSZlK0dNaMF5ZiFCPbxN/O+kxJCBdTvRbRce6HVXT4sc4qf0M
KIN9mffkMRETFCH65GlildMLdRhyHZCI7DbRfnXFRz8ujCd7aslSGuNEta4W9oIfsO32SNQ0s+0s
QBj/y3TZo3btkTD2edej0OTgNltaK4oPVsotWsKyjS5XiZGaSQak3sqUdyRaXiNRhlIyTjZa05v7
blfqh2PTPHcSa1QKOpfdbrnX3ZHfz4Pgf1pFllvWirPlUo4LXwECNhm++703evXGcIvT4MFsVfcU
tyawAfbTosFX01tsLPXfauiAd0wdSaC7PtNMu++wLKHVocPvLTqsSP1NDWjhJkOdHusf8NN6Lvme
FEErzKDSPDf82REYv72h17YbOGfIwdBnLGmIFe6U7Mr5FiJy51DbQz+eYQEA6acyYqniLUpIGgMY
OdYteOCW5RiPub/TOX8N8Qs3l3z9wAd+yKh3Tky+1ZcJ2KdWyuQjqInAuIdZDT0/BxLVlwgHysxC
pjOHNhmhW2xhE+u8ROEoy2QhGmwamTSN/m7YOwmkFHrnRasIrpZc+e5q/yn0Rb5Y9zg8s52a5ir+
kH7Oa189ubg3eRdWN1dWv6ecG6+oVdnmUHTPzzxwjmHOll7QDP0RkwhUSouvZaBeJ63QbE/2qbfX
Od3KM808nSZw4ystAp/uSy/qe+2h1WIHA5ni8d5SlNlSqv7jOgzIO4Avgm7okWdqoaNMChP9Msft
Adc10C9RQlMjB7NHtKKP7+f2T9qGK8qwbg9c8ACe0H3AzaBpKFDWwTqHcWjsyyls4El5rJTn+/VW
fUCk/9yRfidRDy1eeYBl3Dah81R0EtKUL2xEeuxCsNysr+6gliivTXm6QppGU4vuBbdkRMKmASaR
AifVfnfGO6w7LywUZSPhU0tXbtu2vMCdPLTtL2PveKcFRBN+4u7EbE3UMC5tiqmgd8vxGw5g+ahq
jxonziILPvD3958cFcb2WQSU+X6wiqg+2lOHlKBptO3WU3SS4gRNJe8wXEFkDUtm/tHeLX226Vb6
jDEEuT7c27QbU2oOikTrm/6SKobzJtIVvSO3nY3W+SVWsAj+NAWXawq8u4+cYiR7iZSKS1hR/hXN
goEmm79CzFDOj9YlIEZ1KI5AwlH48YljA824NfG4v9Xqdu7YbMlp5o/pN/d0piqUQH5A4//E/rYO
Fm4QwpNAKIy8r81MVlAcQJVptVbt8A2wLu1xG5V3+wYXS5WIcTWwfGAoG6anUDEX4FRVqWocV3cc
8f8NQnqpRG3Y6o28CKz91CqQBso5ek/KbSQAdIT9rfhy5hZDhl1KsRGHCR0wQTQz8u/LdpZ2j1ZM
VqvwkksyrrDwp6i6CdAD9IZtVLjWM2PQu0SLEt0exyPZY02tQ+LXXwwWzwF2/rbkitjqjLrvG9qj
ZeJpciHmrdDtejdoOPDx5RCUEo6FndmNMyLIRevk3FnqtdjuAJM2DKwhAH6i+sesFvsBTNLNVNSF
F5pu0WEk74WtZTPMJZmRkueo9mvZyM67pGMF4L2bhmUW2c9GoIJZraVuFwNBIef4Zg2Lsr68eJxR
+4EBwbJEShk7n11wdV9gdqtJzCSnH0Yw4JcLi5/OspJKvssQ3a1Xz2545nQj0UrDoBLyC7W04drO
cil+EJeu4s8frXSrukGbvqZNu2zFjd3RlR0U4l4GaKM0ThUEmnitglO/9baSJCI7++BAGOMbdL0c
APr9ZfYddCZEFS3I21hGnCYioJGpT6ndvNGpvslfYpVq4mRyJc0nEq0vXz0mjo2fEWLZ6F6qbOkU
7a0fbfgUxr9X5XC3OaCTvlZvdNubw284c4lbHvxMO28YTQhZpYrtGnsL6RfmHaPlSBr9Y503yV/S
c6/rfqlqevKwPjLsBXL30Uhn53buJ0VPsEqxF8Ov5qXhu+3GfN8b8pU9/78a4CpqXaReDy4rxYdD
3XmwDEvrFMJcs1m5GLNPTVKS/73kFII7EWcxpt37bzE9348I/P6jeTWIDfm8CYNqfmtBj1qwS9kb
+y6PEw9Pm5L7SMbLlVHIgZzjgdQozdCUFP86g0GDLWxQNjZpZ8n8RoeF2amkhWg3hKS0JUW/dnbq
K18OpESu7aB4P7zWFeUM371P9R05T+vRmP6+xpn+9972BLTnw6VItqwQYotM+Psv1kzlwjzjaWM1
XvkeOFeqqzKPzzpvW+TJaToOyCRBoCb+V1hG6p6SPXNXiVMreIZduJ9Hl2QGc4Ex4Fy1z7gzZgeM
U4Pwj0vQJqrB7f5YpGdj5/0H3MKsFuyNehQl3BRbfonSB5RRFS873L3jvYam683Fb3jVVsCgUTyF
GCcF6QE1/Ig1Vkgg/EdBci/zvciJGTMuOQFsBB5rmlNlVun4p2MecIg4gI6Us4ngK4S5zWPT55f1
SIbhK6V5KC7g/QKDJVZwQ9ygHQMVWgIv7bEjivyH2rUps9WL603BCznJic9b+/txHI5vbXfqNn0U
uY8Y93ZHMgmt6y3kahHfFrqE6sGDX9FGyoYeeMYsUg4T2oIT331huP/GxYek94oUY03LG+LBwQdn
EJ6mv/x1SRDhJtNWZbrhd5FNNc3G3NcNkyE6cMaQaG8TR6Lyps2Jss6c1o1xbsMU1WMifQMUmD2f
qFf1xF4yUbasrcw5U7AI8VaojCqJjMXji/rB07Q6dSr168EA8zb+x8TPvPZRZhDM5Fx6INpihs1J
xZOqD6ygwSQ3RJgFOBHldbTRZ2aclbgYVdob7Vb+gdR5GEfSEaIwlWWL0x0THg0Ynk21z7p5gdnh
IZQfeRsalnG/XOLLJipIX2HFYh4JeYh/dPpMEBweQZKquYL1m0b0fGPl0heRSFjHfwBkk+jFDBFM
9woACnesbNTqwbXCFsGmooydsEO+211lg/fKMN2WsUen1lTJ9GBATuQxNfJmJ2oLjaCXkO1cr68P
24BkKnYWeCyk9VM01dnuD7cooJMuXKtmpW3h9lXolXJMZD+e9n2mHf4jsjQXVlDUOe7usdVERtXF
aPP6XgVr7zs4uXeEYa9HPnEIMkIDcy4nKWBu37W48/1Mtn3dHYxfWPCk6yJ6sHwaPFRHS5CV/jKK
QfDgwouuugVrTrWF9kPymWAytyQZXQJkwh6cR5vogD0BKfqjFUHx7itpgw0arqJVI7f4DfzUVIHW
X3alzMJOXB/eWe7EfH8UkxO9dSXIwkNBnmzSN3NUyCARHtRETKixMuouy0r/8bmmRrcF4y0x3fCq
Wthip4wde1H/2Itnk9lEssqrq1fePtEqrw5RfCqluPI9OzVgn3b158mavV+Aqi7wUCsRkrs9Jmzd
iUAj7tKSPQXes+A/LpTGSlWFMPkl6gC3iO3AyqO+SpIRizu52w64gWa/zwA0cswwRmlLqn9cAUsv
tiEtYylXYUvyJ83EjHPEYg2HLG7V/OssrP3RAFCKkEMPZmwwgQPUKyR7eH/jISpzFvK01cAjBU7i
mwy7yk62Z2LjQVpTwnEZ1qvi040dxEx46nM8vR9puyS+RZgrn5AOG/+pIxzTa/YoAFDFbEHsebNS
f3sbGa+LrQxjHSPHZYLai99jNUuadzfvWcIl3B0kZ1dy/DYQOq/yZNOecIYvC4XycTFQl2L9Cb/B
sOJQrweHNM9pov6LL8aLmCe7GUUgnlYrqBS2Buvk65ANQz3Oq8BOmDZv7Su1KxKJyV8t+VZkA9SW
uDSXB3/bnW8R0CMJU7blSs8T7dlMl1Wp53e95bmcA8Qnp3lPAanC17s2hsiy3cso9nsigl4XXf08
5cuzIqwTjG5M8Tz2QRxaFaUcnOXOBZLCrtbeF4e7S2C0gWH0dvtNdJ6vN5KBD6NGyhjWoE231T+W
CP0Gq4YVKvn8lDLffVEiK28nkyOl+NapmFLUgMghuIo8HnWooQWxMDrlgo2gmjjKzf0xVLnGyOPt
7VO4a4pAQbaAGQAKerDmRoAAtHdN0y5o0/tybDe2aFo19No7oE22KDrEQ4fcWZhsG9qXwFVsW1Qp
DC50sIUK2zjoaW7XVDrK7tHx/mxBVZVEA5j+6negbxi+9nHBR01BoF+0U0Bn+TrfwWa/NAR6+Is2
BiUlgqF1/xOpGd844jsYeS8gxYX9/Gd/sRS4zDeiUxiKgqlLYEEGtQ+WE6mZOQlQQzOH+Mi3j3NK
7ONLfGiilmVB5bBXXiVMHX84KnJwbQfEqnaYMkkf/eE5kXUKKMTXN7cA0DKyd6wQGrT9qXS41/E6
su6ArhxN4l+PbvVD0Yu/ikmghHpIT6zRJbWXeRkB7EA0vcnxLh6QuuFfJ1Sq6G9tuMBn1sMPmaXd
L/YWFHver+rKTV2kqw3lAM0MYDEMrxiN9TzsxInBrNqgiY5t+eugurr5it+zKbZvKYNYvP78rjpl
kqxSk5IeJGgTqF4pZujHETrtGy4H+weYYZDm+LfqiiGXfZie7hHImtKN6yDTJ26p1Xmg12Y++lbH
vu+tAlyyUrNH7+Ly93mYfLM1KyHHZt+YqRMkJewT6xGTpwNu2eIbASH3qczfsdrq4Z0IYcey8vdy
FBB3MdQRJCrKZ5+rvGj4C4+dqNntORqPe7p0B6BXCCxnOnR7wY8j+UkAYBTxcd4oj53Ndyu7JgtQ
Mkc7kBN1fzBHHdGWh8CW5JQqiUDncqdaQ5dKrXsrxxsj7/4r6AGpHPD0Rf2c54H/sZDe2CLzhv98
Fl0lYu/A/TCSr+teWerkyvESikiFwYm9ZK0MjYHhvxlQ5paxPPdufMetkEE8pERzScdP4Oq4bZfk
4MQ5JOsXdf+PJQsJtAUbpLSeKRJqG9/gtpcfS2K0ff3armcPyFiFvGZr3zBOvB8Sct+B1Nc7usX+
BiyQPO+QrMk3SmffVKiiLVKHaesBT3OHT8riumUxymaTkjETobz/EWEvzpvLiPbn2TAM1SvLD7AX
H5VwWaSmW7RGF0f4jrNWbaZXGFsxodrCjeIJwEACrL5HOpSWIDYZDlg+1lyBuGBohGVWgXOXKSX0
yecqczathoKAGA7QKPVzE0/SVoJiIRHbegf2LRoHsK3g6xH/G5C06fWzueA6juNhESS4SPyBRP9R
Qo3T2ZT338T8j7Q0kMZXH+Zz1mwcJEP5bKu+9devkIck9rHZ0G25k3eMhrixqQhKSEuiAaetzoM5
YTNjduZ7GZwmPQtGWBrvMNyB5xPkm/JtNSoqL9RnjupdGB0TDgLozi2CoL8vn2xgzSjzSXujwcj+
DxtRyv8EljIkzzyeidBgZnJKXjfBGTFpCRYCfb957D+SM4CAhHDgbLslFLA89/+nF0Sk2zvPhY2P
FMweKNb5QFCZJGmMc9aepjWTExk4l8UWuTniI3n5xfWAcOUEjIF4zr9TzZF6Svg1ShKfDByjG7HR
MUK7/fr73ND4oMdcCO1w0Yzy+OlYMWp3hS1reOgDzQG+c9d9AaAydOzxqiBsDGTsQ8HxlGAQw7An
h/e9luUDFuuPhzZzwsbMNtOKQwooPKYgkcI2sU6uoOYXLgvMtj632ZoAirm7kj+eUsX1/uPJLgUK
WfGY0avOLvt5TK6zjY/gDqpAfurntGkMMkBbSS9aCn7/xbCmFv8dwrjwInVCXdvaUbxy3DZwFuGl
TZvuHdqWQpYgm6wu0B5OUFwm6foajU4aQDbDdnZksePby6Nsl7PWJKNjS3d5iNpHYij85JrRK01H
FMrbd99a9HfEOAjfyhitK/Uz8FlwQEds8kgOWRgQ2MbM6VlCAUboN/Ean5C2KnuPkXeUl7gr1DJQ
JA9xa4ZWA/v4NyxdmLA5lOhxJxZgsWlCG+haL2YugyT+9w4123jigDoKH3PG9svxUXF35l7IcoSN
n0LGDo6qn6VUH8vLhckqXrrum0LHNfe4nlDG3JkANnie1BnsH/JT28nT9AOVozoB21Ap6V69Y8/r
M2Zm0RTEvhGemZn87RAroIdP5ntbRN9xPWUe5jEpbQWwbC7h35J4jGxJkMrWX/2kU30rkzZGG8Kl
HKZFZvZRhSTcUmAVnkJ/yd/LeRq7bx+OvegcWpNqTeE24KIxHxCpKuU5mIQFlS/bEpmlyg5KDljL
7fYJUZTxskZe/DPbuLGydYExwJOKvpVBcwlesl8w8ZfWxZZv+JQgnPBWFOXVN5dmEsr9xSBLewY/
oh7ZsXBAguSH/4tr6CQX9dz3mF/BHG9JZXpl1ui3tDMGDHJCnBSnxp8+hVWCSIVVqQf0nMPmrMCL
9NqUrC9OZQoZRwI6t+Il9b0+hEtp5tCimprf+f/jLvodP+xWDilPyhFo3gvcFTbrJlmbI2L7kRGX
ewxRMeE9rpKS13IHFBorO5At2RHSJQX1H1t6DN0ndnFen46H6YKE7GgMyKdpvgsSn4IM68ZXp4Wb
xym8ns3z+hNN+kmrlXWTyK9hsQK0KHLzhBFduBSh08wOrntmTn+TXcAGmg80NSfnJtVdqkAbrfbj
APHJbkglCL7/v0wgzBV1bPSEPhKn9zAu7LYMo8NzJKkXZgO42CYctMOQIC5Z9jG3scWM36F0fky7
yClCIaNbctfQnkc48oSyQdaPrBYMc0BNGopinq50BsFhhoY/SGsYSaxpTyCWLKMZVICt+uyg/u3i
kCHBK/yRzLYtKA8AtSH962wWG3KHicsDChgJkl4v2hIHtcH4eyDunM/v/UPvz8V9I64pSPMEt+fe
Ok53oexY4jG57+nT6Z4xGF9pPrHRQCM3U1orefAxkfQ6Rdor2p2hYcpb9sQlU0SLqvFkkm9enGcL
TH8Q20MZG/m2P1B+YRifY3FRvSxOcnepNZLZpZGIOzX3qSUxtXE/36M90sHYbdi9hVMTv8TmMNDU
Q7sUqPsXqJ9EtTT9JQzzDOxlLqFRI2RRqFZ07zbTy1N7l3yZBJI2qpy9CevA3IUOkqSu1QhMUgxD
fMyFCbOYKXDIXqzsUt8FpW/HILsdPnAn6VVsycVhDDMpFzd7jKfBFfwKQkvph1dZc/eP2jStChlc
vBBnVY/aTyfpquD9SBKpfAazh7dHmH7KKDxn9sLszeoKqOdmkdZ1Vekp+l6rpKIVxG4U0bSJHi8H
bwbdSrU5MA//mpCOMmMcSA+lCwXZuXZ94hboTP249v8rvFfQE1ykXlXuLd6S5kyJF65kEIddZTsY
WS3Sq64ShY4IbcHyltPV/RMJ8Rwg3Q+lxh5OTk2Ucs8UcuPxYLMsGvH1SqMWZg5VYVrQjItKdZZd
BT3PY+4XpqSqT41Ptg16PKd6qj6f4IDrioECx8IxwV+/p5xxGNgANEv232wTuJnPU4jq671IJPxG
k5DI/04R9KLyiWTWkR3IoK2wlsnJWneCjMnLhgcagJkrK6SpuAb2eg4QSwbWKb6kY0Zd+4hKPn3Y
Trz+qBGSPhj0KqYxV7w8f15s9OcffTqPwQ8gPlxB38Yf+2HIVbJRo+bGjQygnC4PioeXW2C0KPxZ
sVimiU/Tm1941GICCRZb25uL06grEvyqRY8z8ynf9cLo5ksehhi9HBf0IRWAxaomdW+Ici34ERjk
NtNDxKmyp9PO7FncY6oqZMB1iLicBmN4ZvEPQ7lLYdaHSz8EWogYfkYLRU4as8R53UC4YliFEc8a
lsvi+YYXz15A4CyAXHNHuZO9A27AxJluGse7ys5XdYX+spKsKkxR6JEoF3I4/5EgonLfjypm8BBP
ppM+WhoxXprKnbAcZZoYv9LMWedCqeRNEeoWPuQwwasOnO4eswmXs21gaoXYOs9cM7f5IAFjMItv
tH5g943/nk5W5vUjdIVgdkmHOZTB444upAGTctg4Z5bobCePeWFoFdPwgF0cuJ+SYiPR9D88bK/y
nnh0NEeGXYFfUTwpWUvPnnanUxXg+7fjbONo2Hdwn59GHR3QJ1Lxp4yzgrH0HrT2evPGut55VouE
SuVHr7pUT7QV6CPru6qymnkrI9MgeMvJnalwNmMzRKP+8EPn3shDvQdttZq4lK9/mWtoAdLGb082
j24to/xi33fe0nGv9LhHC2ru9EsnECr5wYZhsA/u78rEKt8CnQliBG/sCIrlfQ43EhX8BJVO8Ldf
0Xv4LQRzRdAi6fIp3ipqvxFEoVTbiHuSLL1JyHF1gTZ9C51W22Zk2m7OXvlRaI/g7jtzK2opodaO
KdszDm0ZOFL1OU3soyoFulyT1Tef/dL3Me61sNRn/CXe+5V2nkLNNKAdfVLDGJkEQVUV77Znvnjd
21wqZdiDuu7EplJo7kGcRQGcBDklndRTzL4cFWrKsy5uM+a+0vJimIzFGHwaolLL9w6N0VWOdguP
AgOnIdQ6hyYrt5y5uCC5ZVX/a8YDomkR2ZOQoXnF/qWNNht1IRAGilToYo0vyXKkLjaRIfol1o0F
QL14biBglf3O9bglRU5xw1kZHR0S8+ApfzFSxk3ShTpU+xNkWgFl6b9mNlqSQKjC+hQpANKyeAIk
939NeB2UFdKSwKvHphfwg+BqlYUIfsfJwSU0ueOrZFuNuX/d18Rwf9azCg59lfKWREQ9YS2QNWN2
kdpQPrs/21Rb79fnwT/6++zDJKs7FwzZrvLJqa7C6Q5LA+SNnqKiTln4re/IxVKFIgz1qitbBr0w
xCDZf4E6s+s7/KBcyYVjYrlHA4GibiFs8ssYJiNDJcdvCV/AyBLh9QYhqLneK3K9GMBd3TNNCQ5Y
ovsBF6EaGkwX3m/kmKhiwSirr9xAblYz3ImkWhYHeFip27A8bCkNKuSH19nckQ6YCZyAoJKecfd5
y22A8IEeLfWPUTn7ouC2oHtis95i2Dn+x9DRaM2gydB9t6d80GXxllA2isq0JHH+mUX79+qal8qe
z+/MH5KdJrTBvdIA+grVDAl0JHVuXli7zqYZuDdP62UCyY7sqMzE5eSbXbL7B9IAC2W/OoOqTdI9
xZPBYebCTLUFKBKrHAVEITabUiXppfPuvgnuiN/o3S19Mv0o6NUJtjpjIVbXaKr8EHYGX4I621d9
CLPsIz36fFgQ8XfxmeeCAvHMDdV2gpXsAZs7ROZFaiWsRXoJJreYr+y1xg9IJcRyvErCJc/ScDN/
EuwI0rlYfj80C8K4UfBDbm54PPe19dElH0Tcm1rStZ9ngQpEUUCh6Vlrsz2Q8WnKDREy6rPAgKul
fJrEvUOo65eDQcz19KQ6lT+Sl4A8RnphNsNYiePV9jYNv3wrvSVxtKIZL5UZyRXzc8VIocAOaipn
NrJTi2P8e9zjm13k5j9IGoPFOpD+t247bELrUWt/2btWAjy4pzuXipB3J9C9Pn2ZqrMxBIW60Hon
K9Fu7okI2IkePLhUKGFDNGXwIsj61WwB4bF/HwJIxCjVghcPfDxVqrcyRK2+K9M2AfCfl8lw62Gt
83YAvUIN1m4Y4eSOthZoUx34brqZd6/vb/VrJ8AHNAG0t/akEX74QfG6/C+f4r83cU0KiUFzPDR9
iRjVRsNpUw9tYjSP+dlYxUU+tI/6E7XTR4jqW4rLoz25YgaXaA3FkmwiexDkNHuAF4qxhBWCFMWS
hv0HS2cjJK9qyAKTS3sg26xaBlNquUc43XaFGluSGgSTVTtOgr2Wd0f1efaJqqOoMWZVoHWA18zr
KmpzpoqfqyqD3dsEhdshgiQZvkLL2CRTroJ8JBVDUHxM1iTQV8b7KiZXV+D3StLfzcjJMoYchwSk
Qt+zvqkrm8XmO+6QYx0yCW64w4B5CgStqH7FJ5EXOa4zqHfmXNqE3ed8skwiO/f8lQwVcB66hL5F
MrqgHZumN+FXWP1U4UR55LTxBtp26S9GcjKvpNuIIoFTVqHz6QeKQXwTR74S4nbcILIaRUuM8J4j
zeybXNbvaCBCLoajBT8qFGEW8rJPrMUASIFhdZBn3ZRSYoLC/G0PdyfcQP6vFybIX22ZdBdPg3Nv
ikrTtXvL1xfkOmvESChb4AIZnK+mnNQPtYtYZv9EUEVFO8mZM0lZ1xvpNN3yqbdjNRMdcjpHUk1A
Oh7AWatEB9tv6qO9qbNqdDopmdx2CZU1SSTjapRNhJ0Jf01BYUvbuUQV2o95bUWbjjVXatJfOt3O
E9x5e1DU+hpHwicNhb7Wfadq5Al04Mf6cQbC2TM1ejlgeRSD057KULzQ47pK4AEsQCvp+1+E9YYd
o5Gh9oA1vutyF8g3YIOcnsCs3ryXyuTt7m8asb7UPUuXcfcxu9O3kKNS4VvKHzcFMGd/AmUybb6h
eurSp/AWS9WjGiALWB1E/Km77d4CjQtSvf7eV0jB8LVVqPl06khH+PiCB/jluSsRAznHh0zyENPc
wsOPZnqjRyOlTe4iOU3wS3xIGRWt9hrCbdn9KDEWAWT8KonLinmbaIVvd7pCkVfUfNIqacYHv5Nf
EI4sQcBvK1GcQJU4oLt5432jnUBuqv/Im3vRgrYBKvS3ZoPMXl4s4ntPXxg9Hl15aZ7PKottu5MT
FXJklTGD8B0wSfqx01nOK0Cjub2anrwza8Pj0hIirr77EcIhcQlv90M+gxFuJ1p0cS+wkBIsFPg2
Y6TbTIWnrLv6ryd0iOdgEC/qHrINUOiJatvlB3n6kRKJR+wS5gxzYochFmNly4UwfpujvpMzSTxs
nlOD3GKn7wTOsUXUrmbfNbhHouoVIObIMtaMfPLxSe3aDU6JCtzG+LGQz0umhmT2D/oqU+0vy9K2
JEooOMS35nr5seFp9MAQM7TF9pWEFD3AdTPbQcgtrqGr80CiygiI9Tq2lrESqxf1S5HhCLxeYhqe
G1hMTXcf5zkk2TVSO3htk3pLVrhBTC5RwwBtGTLHdi3l7zheiaWDCJ98GBXfwE0sV4K3Y3zHjibm
Xj87Eme7EPo7kWsp9NYh2nHKwFXS6iHY+ValOnPneVRjtWcnivBgUSXqg7i3cPwCGHzzHuqVrBXK
0giGlKkAs54UFGykKAhEyqxwRBhIsZXZPB9hibGuxgTMULpMue1lLZ+IKZkW1QwKYUE5j4gY58rI
Fkoywk3laFofAWdF4wVGB6ym8X0kQz6UuMdMTqys/kpXhFzVgBJ/j7Xee8cMN0cLV58ie7FJE/9+
u6Fd6d6j5U4nkSFbSZ9S6drW0DXPKv2KfkrWz/cKAoUF3PdS1dn1v/d5pYab+VVtY9O1cOHbb1Vh
5Taz0IPVWVAD4hei1/LpwxlFGjmG3wtbRarjuYAoPeXY243XR15W+3ppm2H+/ce3UZ8cFXA2PjIT
9xiby3UYB2nid4XYrd/+apfFPBlZ4ROCRizeeazPjFtGYqTgMLK301OhS2eqNGIDZeGVkoxwrJOg
uHiI6Zw5s25wmht+/07f5qqGEJAuYveoohsrWjRIl7huFG5h7lYbA0fq8z4uLtIWwXyK3OpfEwwW
1zeI3cYzFVQr5xCweOhyWJc9SQliYrPjbqmPw1OURAVVAxUAK4BlkzyZjCmYYGBqat+0+/CDW8/U
GzL68++cMJ/qObDRvPHPuQbw4qkWczquJ6FJg6mI3BI7zb0NkiHFfQcFcB9VjJSjwRldC8lhOJbZ
RDV0nauhIgBIDwjimL7RoRCCr+T7aHqoSVbAaUfelqbcli7TMZw7/y9tIN2BYeqB0SB5Z9VzTNwq
/7WZraOWNy9mu3/3TjvpNyIJn/cZKsCoOHQREJImFaFh5XV7HrrIPjeJbNdvWA6ljR3JpZDhtOhp
GPi8xJltOLRjMc959yRHM8KRM8ICDO4wlXPEK8rnjudUup7766XxwiXtcOSvhqIN3MvE3ng3JXkd
0PFp+J+6ZlEtmfhH8pbrAdaiIAjMbovEvy5JaCX16cCG06L6u0A5wHI0UqeeFdM0any+PdbMEbZ2
agePE3C2KVR1N3OEQqzf5etOSfiVvX/bJcjJdNxpu+qYBIMZyu05n+yf5mnnzyV0Bl7E9VdXJam/
0WrFQpWOJzDm37MSHxLUwa0hEkKLKRoTbBJV2MqYi2O6tdZu3tGz3Lbm4h0BonPkgCjUWSj7bvAR
TOSeLsZSWjvHDLoX7MUgQndoopW9u6uji9kmMH+01KB0jzL8oSScePWQ67to2Jx1ymdghFzdPd3g
Ji5bPpiRvyoTJ0cqlFbQhRFwU7XVpxiWzCpokOqS4zMKA0CNKegXcrCWUi9As9kd5l8OeOSdQHlk
ScwziSebI19jruzVK5QHS4FlT6vjcjbBRA765rnb5s2vt96DZ3IStCGe3IavwYJY3yImiPaXaOxP
8ZNy6SsqZt4ZtrWUSWdeMS3efjTZu+S7YxOEHKd8EW8aNvexkzZ0OwkKkNPlxp/jVMIUrD1ATGgs
MJ/ZYwlAmSRlu0TFCNPUlYcAQI8shOwjRlxwhyggHWe40PX8JVBrLfbXsCP01mpw9N8rLlVgSyTq
FVM3JerlvQXGyRGm/9vDEEqXVd3YNfs3Ozop7SSmt0L73LbICo+ZP56nTNtOhJig743mPOSLPEhm
bRALN4YqB4PEUtsffJR86QNWlMmgNV/ouWIhcbhdcXc0JA+JLGp+xJ6vMDuAsZ2sw9yoKhcyNtlM
lNwhx7eT/Lsk0erFl9g/aKxLSKYGmdukhJSRrPWHZHu793qsQEcLWaFtjegU95fZaPAWupAw7QNL
A6adSGRoAFdE4B4Xa/4l/ho5ZAVW9QaR4Ol4aMwUCmtQaM1Iq32I3GNa1GLoDZXj3VHQjr5Q0p00
eo75qnfH2sOLyg7g2J5cQo1+4g3Cg+LkOxm8+pRF4wVIEYhvHc3Mtgjm3uA7lVaPtv/HJvuS+z5h
7BLmfSDcv/VDQdNl6yLwfex3jGKYmcC4+SYsd4R3o4b4pO2nboAOvUNyv73wp/DEvhYNCxDVR48J
fC9Ef4uAGoznF11WIhqZpn/37NrdDmzfd3bKxyXlGbs0qWDVor1vKGAho7jkSt/RwYpX+cN92Cl8
ctONUPR9qA2c4wnU/9Hht46Y+LemfmhzgCrVnyfks9xcJZG/Q86olrcC6PVMBtXvVQjNGBxZfeqp
3RGPsWreHINP8xltorxi9xl1R3oOBQ3OmWN6LMqPvVvTeFMbO0g+i01+C5nO43qXNCVCbR+QptIo
Imhm7Vqebwh8oqssdzGkRZBFfaAM++pPJYV79DD/Z8Ali795ZRXcvA5ATIEmFZ/xu5IByWJy33rJ
ug2Qi3rfbcinilLd/Uaj1vXk4WPvFc+FrMqDIDbhMMbVC2TytP5g4hFjfAKUOcjvl6gzBsM9Y2xX
XVp/3Gj4hUvF/D7jKK0+HquuPFgHdv92Ro7aHVu0p5kYQmTWlYWqhua1tUlGSTCF3HyUjDS0ouKe
os0gPn7G9Lws3zWWkrCPHKGlcTVTkyXSpn1OG0Q9OVnU3LOd42Q9wqfzj/YA94W2kSzkeKCzatHH
K6sqDmljApqSMELjQzpD0KR7MvG7wNebUeVrLowldZTn8XZLDJwCeKoXUY3LyxcDvcH+uq/Tp9bB
NYbWkyXCOcVvB2aQugNWBrpL6MLMjvnowfRpWomKKsMgRuU1GnHbeTi/SzWrHUzgKBVDs+6bD4FN
JfkHX9rtelPDa01c/v+HJyan/r7iQm0AbbFW3+FHE5BH6eC1yLYW40BuTyLckNSlYJnsRRK4y7JI
Ic8roUGvFP2N3ABJcUsVYNDVtAZXiQKuTJBfgnucUpT5B94GprH1ggvzYVfJWe2Pe5huHCbjq4Pw
KQSv46/4QmmNK0ujpy/s0Ddvk1LTcTybomTF1mXLcXgw56YCqEK22RrilAWpgUdikTC/8m7olW1c
jNGohGHlUigtVwAUwfU6zNyvKC8kLqodW8/gyXTP0lXDz1qfz5wD+uflc+xJBaSt+dZhueSR1866
6+7QvlJTxDbQidVB/skpPmuNewRDqMp9fNaXJKMaDMGTb8lRk/wI8GSeUZ97ngLIFC+wi8PoBcQR
JSj4ZiqCtgjKEvXW8fiVggsKILPuziIqN1oUwd5yo9+deq/LDxnM2PVEj4/dM4Edblf6293mumUi
cQ7QLKXC33UEnjznU0NIB36alJwfOl2l54GfKKK9RLQKEx5bRFEysfViSb+4avi+5zCWsSnd6Okb
5v0LfMbOxNa6inLFaRmZaZ9yXOqrVQXXPqu5OxXJLqdrPS7mreAUyw3fXk4tmtOp8qSQTzSkiHCD
CEEpFk2ajo1tmtT3UC72L4yHXTLNRRJd33N450EAATh3rTDCEFEu4Z4VsODo6QnXiZqR7ZCCeHII
zDUOzBGdGFRernyppyR0ervEMZImp8VFDYEiLjjt14ZJjIJqS+Dq3eHt78WFXBfv44fcUYX4lVTl
VgBMVQm7XXuPxMXw24tfv6giajqN639yVA9beKj7BwVq2WP4DtHivs3aNbHEp1tBGuuhrgNmOma3
IW4yHAnsDYfXioHONfHXf4h8S1AswSBUEhoDxZgEiJmCldNA/2hfnl9S6TYvfv1yBeetKF9gGAuB
sA0a6/YteHg5eXL9HDWP0AxSbN/hKmJCKHwPbQex1xMOQ8CLlDm82VHIkYi1uOb3t7jCFpovr/GY
wDqXQBY3yFAG0Drzdew+xW7LqppvqUXhhjMhffRKWRO9hshOFzODlLWI7LrECFgrsATmDW7yyFty
TOqpZo4YbvbX5TrhbaPyD69lxNm0TMXAVhqYjcP23kOyl+RQTd6fAZ1ttNXCHwHa40VNokWapw2s
gjBnseMQPMU/ZUUNIgS+pTE82cyLv90cO8HqXHuKNDy+kHVc5YIG6hSV0RhsLJspDUpjGrok82aT
uOv91rg/KDSvx0s78jLFF+g2ip86ZB6bVDuCPeB39TQwtn0LTysKuRMZmPM7XXVj2Zd9IxofO+dL
Eu0LCOaAlA1rD+Sor0RfaE39V7zxu2VuB841k5p7xUAzdXLj/keAIvT0WFPJXLrc3eIivuDKLQlK
OyzK62GV2InwMJYZu1JqrVbz3sklIS037BjVvzb36vxvR0iBE7TRQnHtuVLhA8A+rjVFMtl8me+4
bB2FXM9P/uQi8JUUItLTfuixAf7VtUyEXLgD5lx1nQNlgtECg8SNXdfphen8vkLDGZnwzRWFmcjU
3Mptjf4qMifE11oooFjjx61YBO132yEizKJHBgXyOQ1TQcxtir8eXauR4QjE/Ji6EpYNjHNneBgX
9NMYywd5H1njYC5HAs5bW6OX3Y3pxVMw2nmTop4S6oRCI+tS14j5D44jEYvCgG3AxOsXnmfgBTKc
Q3s0Y3pODjbr1mv6e5XuQRCIBIrLD6PSYQhJZ3IpSbcXSTm8xH8Jdcg3gL3V9HgsO5Wjx9Wa7kGL
4TTft2X1inHXs1xORfIw88JcouU9LajpHK08ohz5dUpjVg4TlZ9Tlah5S+Z+hjS5ZmG4H9VkvG0J
R3WphqQSCBUwXz7F7feWuHJlPsRxGve+HylktyMv2pirKe3gN6J0S9bNJsOkB9EPAqzPRueZOWwE
ND0M0+DIMwGHo5lWd5cKGw3dQqguzbnzmCMrTCVjUh1tMT1VqaOo7UZoYKK8moRFqQy4EjQJqCtq
lhOExHTwppXR7oxFy4YBe4DjsK9WqXpkEcegoMlcSLAaLQuLoaEo+p282Wc9kHeQiRErbXbPWyHi
0LzWl6VXfpIB5NGVrpPoqnq4+qmGmrfnRAv1+/aly4haeuDapj2y7zQdJkX3GTf8T4Jbrfu1daoA
rClOu7rTho2qqvEAd0vxhM3Uk9LXOm98HSK4yEJpdQe2URQwX+DwJaMHT1/AErMLjOd+S3yoIrYN
HgbReCx4kvzi47ZGimf99TTEJ1ua07i9BhnsiBDI1W7AllbP+fcvkyOIXLiQVFj/21EE7JJ1p1Ab
SylocAN5rzK3BAo1fYQ/S9nAeb6jFF+xyumWczKP9TQ9oZOnHCBIL/9hi0TZ5svCDfexF1yf3H4S
fSw2q1cmiYWLrZclw8PI7x4NTGgZZEwOnROIxQ0mJWRa68L4zof1BToUuoBB4X38qeHD/Yemjnqp
x9pKMM6Wc0FojZtQamBg0CtU1XTqZo7GOrAIiukOXoOSK/fo/OcNBPHCssrBC9NYJUwq1dAfrsvk
48VYXqHFymmRnWUGvYfQRCk9IzEgHZYgXGwDYs+DasPunXrwb3j8EhkAtSI0F9wOyPqrDP7nt4hw
sePIdWMyW89Wpjm6XENnzNNMaofrxGFABuhdSf3CfaZef6SzbeDC7IPgqHcZ/J0fjYA710smUGyx
x4roFjwdlFy2IyxhaSlTgW5UN431RBfn0q4gE6SaavK24Mew2Fsxkpj479tQ9rSk3WF+wICSletc
OnGXHJ9gP31XYHCsLzy1SaFJhvFOdILUiJbUqxzHTK+P7j2BBCIw8ReSeA3ibRmRkXPjZLt0n/bH
2FUt/APZ6MXfjMK1gxkjNJbXuR6CLpQ6HGNYf1SdBPx6OK9JBnZ5ObE6sQtGOxKOkUtWAZzWbB8n
aniEAfSSfSZU6qOSTIHV66JScBuWQSlZeZ/YJJ5rRufN+qUsb6L3l0+HM5HnA+EXfuBwPlMneGmK
3Y96QNucfWjeQYSs3XvGdf2s+WiOxXkzpBwZWNpGsg+yI7derjZrVCFuVT0zgOmJCG+Qc8kzH0Jc
Pxf0SAbIr5Z895DLQAoxaODrAEZF7KJalkBl6GPqDZ2JGqqPu+AEfxbGX39VgwRmOmPxlqIGZl/T
i9UNCSbplHza28jdW1P8hsvKkOzEJZYUa2ZS82uCLBjkT1cNBe706iCIQV94l977eYrhAU/G0Bu9
/Sio3aLRhB1amQ5+ZnKU6kRHIesxOgyRJepij3zI2SXyVFSuEopokwmXrZLAk510k2D2oxImZ+Gd
3hBkM25NwLaUvj/u3YiCThcyk4gcqoRDo348DSiy/mE/MxjOFkN17rVnKARwyfWzgWawjrXJGcax
HL+jqpDVKmqpy5b3pMil9Ayn3ZZPhSIBWRVkNvN6sCwFcx/gQXlMqgwFphEAk07zh1Id39RNlAXQ
KWLYe2Gvpbdiv+gEjXnIGzW10jove7oMGbmokrRofmloKMU/5oHoHvaztTMNJxP9jfEl7dHFLOpi
+HR1ZfWfR7LBG0mgXlRg758eb7fdIhpWVkJS0wjV4sTOXSKHWHmTju5A19w2bKd54cC7Cx6fG7Jv
914teNq9kcmssl7B+SmKQXvTMYP+7Ra/RNwm58pXbOemwZ+KmLXrWt0/uLaopM6+Hm2x9dclOxlF
IM9JpyInpwQBAC/VcDt+75QOCBTDfqu5NZMKX9avIHUDviXvgRBAjUb+T1xDxpccQq89RttZaF27
Wezqm/ipdu6WdMCQt9A6QKOOddk1Igzx7Etvp1bPzkcHJ2M45/5zqqgTuwLpJ0DaoqPLk1MfsAg2
QQZH9LOX4h+4uVUoWS9epz12PprXJQeGB6/l9s/u1ODZS4ydZ+yerhbm2Ke+Qt3LwwSOKxHGXmWP
XZ9yHDKPuSGZ0hmmk8uw838lqCa5f4iwFhG1XErMlKv4y8baDOn4aMMoAUG2zRoVEhk+UcU559T/
pWI8zZdxFeAkhGgjQY8WSOPmvSmGHJwAfbsI3DprgqW6VkD/m0M/tPiMYhS4lljTXa9T7rggtsyS
6R1Q254zfHfWlxxtIAX/zWN3RkcBO7FFEFVmOgAJExaIpoMJ8XLN3lMuDjheUesWuaatEIxcGdxY
/sFocHzFdF7W95wTYuadql8Cdp3qPbEFJJqPIQ3wMToFMgBJv9NruUEnNquljPZ2waqloKdKGQfg
PkSsrIgVTuS0cslsIZzh6J1UrYiDUyehit+zQGZRrqZ65X1Ndaf1veGFiwkf8DAyeydSqMO29qH4
gFu95kA1oreYFR7zufpY0K7BEJG+5Ff4vce0XTcOZr3WZNwGp/BQHpQ0Nwv+9LHo03bG65voxudA
gb1XFzr06lvcud1choL3fRyyMl3Smuhu5bwv8R4uvHx9pB/EosTNEpSh/s34K9JjtMKEyUmfNOeF
Eh2cf4psSESEee7geAWGrXJmkbLPh+/rgB8jZbzXm2pfOT2eyT5Lgkrh9GC7C9FBirc0zoQjULya
tE+Nyt56MgQMHJ1nszxC4eXj6ouPHOiRu/RAuJP0bDGTMm2lT7QIvvpVQkOD/s+vu3q2+Lh8DOna
xy3RZQ3BMBQhP7QcKQClTiafZeY74d1jIbfyC7vWMeJF7HVLiTMLHALfJU4IXaN0o1fLqntEz/+i
oTckNhsxP/w8kMWeoNfohGKDqetV4Er9VELyH6UZ5lYiS/LSYLoSckzYzlVzv83CWMzJDe8UAoUR
wZN3eB17BOqi/rxNIR2amPjDj2fbUaBQzZqHANOIfkvSfJGJTiiwgCZuqcm0+IYXzdNjlrFWbmZ8
mUMMf5+qCj0oDwZo8VVRirVo1VehsTDzrooVdyPPJ4dX/J4Lb8SDMkWNkQHyzmiZ2Thot3GiqocO
u0valK6KbFKr9YlucWjnfpCrC4dhC0MNXBDAjJYXpNQx0+wPOhDgEMDuSy+WTLadf0nQdNLUH4Om
oMgqT9e+O2SapraVvl9rHLPDFa0l5+ZIU8/cRe9DnUCtP9Q+xWcpTkrF3vsRyE1Qff0jQvV7qZ7F
YU/27GYqcUE1P+aoWyyRpP0JioiwK1WWblklT4+OzvY40o2Rrj3cFHmvzH5JMs9cUDq5Ya4xByq7
OOJulwzC7rft7BWhxiHQ+duK3804V7iS2X3/ubop90fUBILfzBl2OJs/PFegnowynnAJ59PBUK6Q
MeQeNuZfOnkxQSvGcMgKHsE1clXccCwxBnUPqXXFWxN5iPikLtwlYuvss0L3pSFYovpbru3B0ypP
QfkSZjw94zMLQ9wVmW5iZylluI+uCJD4tgDMY+JQ6Ygmz0O46rhuGVMIdLWbs+uIg3QO9EYTOTW3
FSmQbsgdL0PbIJTvaToxLWt5DO9guAm9WJ8fYgwCQhs9y60ncEVIocJBsUl95x8aT7w0/Yq8YtLZ
+GRLphlX+MFco26Q6jXZHQoX8kwnRUhYb2aiH+eb3xVu9O6nRyX8K0N7YOJ8gldMdq53E49PSWst
4bggjVzg4bUbA2TewNSNF4gv3NrGNzrhvOv1Rjccv8SXO5CPw1Lv3Y4pXBEBwvuPbJ85b8vv93y+
UtgWHmIS7DKmGbz0ryuvrhjk6hXzksmbCoxxIs8CT0r4WPMET1L4v9ZJ1hc27QkdNQs0nF0gdeOT
JHN6BJ/U6fD6AscsXeYIxblR3R+JHdITdC1CCQ2g/L3MwQrufMPMFGGAFiNASucLdyYgI7JeZGLw
QWBeH55r+XzfjhjKWnjpomx6giy2hE9lc+dZoVvbqkqi8Kfb27o5EiN7O3qIhyT4Lo7i22p86BLk
OgcYgZak97phxdpS16++syESUX9/ECYbDx91J8MjyPtvTJWyhdlAVQojvINoQOUSL7zrx0cchuQD
qUR1O6ao0LTh6f76XHhkhap63aw4tWWsfc7A8shavXObxo5QraNHYjsUOuDevX+oL0sQ2rmyMAD1
GSv1g9QhfFKokAC1xDoWwvFBkfeXFOWnyTlLIg2JpVEZbNvUEqvVThrC83SHwS7ghEkcC0fUrlRP
pXWAAKGENBA67uEkvdgADXPvRynPSY4t1xLpSNbvwse18+GDAfEGUEIGOeTssD+O6iowHh2M4KdQ
GsQH9e+53gvznYpt7wFsBKrvz3COMCEa1uQtt/WUtnGSfs4RQa741F4WTE2eZ5jEfLGknEpSi0wA
uQUCmqbT11ti9k43uIDSE3IIOlGs3vtsEisordnW+IRlyd4a8HLeCSuQm49wgs2KyFzHHk+R1tN3
zTCVAPNZxCzHeNwWHYp3Iz3054OKFAP7AFaa12KuXhs0d+tiGYLvmaphbO4PxSZ9JgUhPyRtGF1k
yRz+nNk3hBXVe+9SLsGztj8xsa792OZ/hucDEC3d+D5dUKjtkTtwqpdDRPWFpezcs7Txo7ambULa
Kvw20VdhUiX0mXggw/EwYQf6Jifpv+4yQcUhBZm94Iuyvr3Nchm6Pn2nZbQZZAisin6fZqZNewAd
1d1JcYbG4otP5VBiQoV0MTCNhqwNF2s57+UXiFvVs8U4ozPQSMS1qwKs210oQBOSk0ztPTdjYDZ0
1FBjI+VtQ4Bg3YTj1E3m2gAhUDSblJSBaA7KOfLsm3kjYLqi+LN4qYO/+COisofEUNwVb7dubE+Y
P/EtTz8KarxLPLENrnfWjE7XZVjDuzgKoN3KSgWACCq8uE/hPz+unK8bQ2a4hpts78es8PGBLGqE
QWvWmF3O9+068hSQvhtz+W66cpuF+ISC9OtwsgNgHckkYYq1eUKKlgfKdi1wJlKX4EftVUyNaMKH
aT89FJT8Iexakh/jmskOJUanJNNimDil3ftLLcq2HaodfgBHMVaWVc11CbK13byq6YMwbEUQw9FQ
BIg+/7Xfq0zj321leYbOiLFnjjg7fM8ZSPXR5qkRIujkKHGQc7uJ4hRCIwY3LfcpM6IRFLolDT+k
aoQrAsOIuWGBuAGGn183MPitSXFrmQHyelvQLIzP7+NfiIT+pUujUa1rdCX253p2uYbwlYmHoWiv
iFkYG8ZP55YL0esK2EvrNmBbwBvOXGFTN0PMhNd9UQnj4/gVnsAWf3nbIFte4y5lLObTdCp8nCbi
B6+u+q2ITcJkAG0tIVILRE8fycN6WBmj1bdVglYt7OD36enUVuyvaAUHw4wuAxf5OFbbuazPcOVA
lEvPbmGyt/YKMTiKhiPLiXdQsmgWwdwQRdqCtXmaFuFdptaQjL1HUXUm4vLIsGCSLMhfvwVsyu30
/vRxGLD65AeU0qtkaPJlqvtBWEEa6Y5y/GAEMKGrLiPFHsl7uyMYZT4NFIJei7wb1TCtY3XAwI0i
H23HE+bzWD9e82U5X1akm8/LDsv3bTnplNI/sza2/xdXadw3OfdHXbmuCeCRoajwrEoPixyR7gL9
9zeTvRaBB+2d7L0LLZnSodr9hHBIWw9re/696GtYjrrZ88lEx1kpP4M/B3hRx6LHbuaz4PoQSw4n
F8YRzxXOprMM4Kxb1Y/w+OK5vbDR7UPJpUQaf0oqQeuUe2QhF0sxUvtqjRJgYXeucktgw/AL9E7V
PD0DAQrF2NJlcOvUjaRMBPEajm2wzz0SoD2xHLepdW7J7yn8KOAoU7zSTvgDf0I0dGf+FVRDHJmU
5VUjGkWuOOi5C2P6qJPmul7UZSYQklxCjnOWyTc6g8w5rtiX/u/xp7O+kcdWnBVY2ImbGPjma/p3
bJF6dGad0llWkV/GCk0w6qRTsBjCiEBZReHLetdeiOYIMmimazlCYPt4YdVdbnbd/hHOvNM4aZ0/
3sUYXRm95u2/H1gbGS3XCE6izVtzvi3Wemfbd5lpLR2HEBKTR8X46gWT7bmLnjDcl/oE1FO1VRRd
huQ7rzr4zj2kHejDPWlf5iL/YY9lyvPkvYBsffyfbHPyckT5f+bQRP5PYc3puM1Q5pmwFgx1Bnol
hLOx3TjWrKYxUyvNjvdjBisTgDG9dUz2mst7JX0asu/n3HTNRESd0OzsbQ6/7wgN8lWoR9u1m2MC
g+Bc9I3gbKdAPUP7opl3AiSBkdWssaXzcfFmyG5lW7ia2H7zwY4kgV32fUCJrZ4W3+F7+pm3KSGz
hf7kWfW77S5avxTmy4g5dPoI+RYdnLRmfQtbG6Fiawk4TFgPjXbjLEgHB4gMLuaygHKRgHktC7C5
9+24kejL2fxVtKqUITpfF7UHgjohhC3LYdUmtT2m5UPKJo4Y++dCJjC22H0nSg6OcaDNbs79pLwX
BLLIYNzQPkupyoE0SU5vdnwnEbF0yT/GPLqk8Wnuq9Rn/Vz+81ajyGhJET+zbqN+iDh+OBS2SHd4
ZUpo3OHM7LT3pxZGkL5OLav/3F8YiLvtJZ3gS77cu5PQUjeSO0hw+QRBnj8KATkja3wWurIZVhdz
qnxZX2g+c/DzqYqAtPblFhDZGXGz97ZbKKES+qkiuD9q4OrxrXtq+cIux6BClviNyQ9Biq+f05gH
dvizfBgzyqRSStXkE7o7vMXGjtoYrG57V0FZchp7AhATShg/LLLm/IYZvcKpM+YC42GTFdmjYEzI
bHoAXhdloGCYyr+0VqrB8dPCeTwzDFxOMgNHlEeWpYy2dbOT+FatQssHwDlf4DZ7dYcbm3P0Nj1V
lGfS4ZF/aH6ehjLUwh2+dwKUMjqPaSy+fhuqjiNcCR4ozX2CP4LdRZDABAnK/q9QnMO1YE3IGLSM
ekbAdcRnL6K0SxPx24dCQ2hJyi6BOwmPwpG/ZPyi3sHymKo+dmauxmkCyEJcEGM/7/kflVK4Zm06
9v6e/I4mkFSplFN7h0OwlJHNK7mkcqHK4tHHyRMBA6T4OAKiAUA5q5KLkqMZzZhVuV0IpIhak8DU
ITyJzlvpUZlfe/J3TvuRATgNnX4Zuplo3jgfDJ6hmpRa/edmGm47jkML1Hj1F5HjzCouYzsWko1f
emXlHER8Uf45/F85teZ4pxMWZhQlJwJvSFTaXFB4qHa1Tw/KcO3H3/Ye0WzKUUHP2nBkV+lhkpuG
eJGa/Z0aZXt/0C2E7CZ4oidckLHxzIMyknjJ7kCup5h7181Dt32sx82itRYE+6j/vKvoZV4V9mna
yQCDXXFiwjWBoDHoCwTjtcpiFQgYeEVtDJdiPloc1HJPpvkDP7Sou1OsNvCZqv4d6BJaqkZN7TjU
BtJ2zKISvBmGw4xgZ2rIuEoT1qQIQSSVfXRPE8/X0g/R1df4Dja58aMeDkC9jIndUQfM3hOZPhSf
416QK9VoCw5wJSYzoCNtRGptaeQ98MhF2mULXhm8tDXPO35SMwDC/115BwFnoQAklsk2GCXxmAor
yj5oWdZVGuqSvugwsztUQgs9DWky1TBUQjExCTGLLEIhwZvdj6DyXvbtMd93WKFj6xHKQvdhlVAZ
qw7Thvky5cQN9a+QGu+hZFV5h+UY/3wJxjTATYDqrx/3xDuQmvtAngS5aifqLesx2y734OPBWK5z
iroVmQWuiMLtDNJjwPEAW6Dts5igDftbIuQ9+4DIDmHwJ0f9veGmHyl79heMK2MLzOpG9H9QACZi
y5iWFNL9vIasfAIjva7Ah8tldIB1OtDhHWBbyYnrynnoa22T8RNOf0ozQvRfxlCAh+wrABxVwsmJ
ozrE7ymgzU0dr4IChAcg4ca5/0OJ6ii7lQvCBye3eWluyhYfJGXZOrWUkSudAI/BXVKbncnmSq4u
kY9OxTchUUuxk12RM0Hi2uoOIXk9vL4KfUGdqX+2GMhm4b2unHiw/WgIvhtoxLDx7bmxuShT7IF2
UQ//t15khema4xv/VCB1pIApuTDuysidi0X4YV92ll36RJXALiGU9AZX9k+LuaR2pazsuZ8KOIdq
Yl4qxrisjDiRTYuUKi0NoSJsC3BtqcAOU/5EJqFpGbObxOjGak0n8QiUVRaNrcjF0mHESb95qep7
ft7+KEgi7tsbCEwRSlKbVIsYx3Nh9AXqHfZmmjL57H3tXkc7ubuHg/WSaD+zGjzck7yOUq22pOVc
H3fgrToHnukIY/ToS94muJu1wWgzQo2ooBpRbnoP6A9uiAzxfHt45cmIiFaBDganrbMqZ8w6Y/kJ
DNfC+4lWVJTGuGHBjJjUt5L6wbm8XjucrK7aw7Re5vNLzh+3W5b86itlxYRadaxewhPXQ/evhlAY
4/rYMUfHHey6OIKOh6RBrtoH+6x0bboPrcHQmcf65UPIDdImMzjXFcbpILGilgZfCzHEXDsljOc6
GIyGebB+uHRtSotDC3lRyIkxswuYc8pW0qm22cF5ddd40N5hpYgChjVuJz4W/VtEka3ohHQ0Ko5G
RJfN/04qH3R19rIuu7fG55RlJ9mJl018CRui2QvWcRp3mDDfvGJ33fg6jimflzgx1OI8Jp31peV9
1wl/KCYGf3QSUAIK1QnVYftQJlgkV5+EhMR1L5XehcCL1HsWwQjm4glPhHFGB7DHsV9Ey7fhBJ0x
khsRppC1P7f26V0fMWbKy2/E38aOVCjx+TR14bmAKvA2kas0UmcZn3vOGr2abxYvzgb/MI/6jRwD
dPgAaDOt2oYJiWp+wG+2uwqDAsxlw1SpXyJgyYme+OBXX2+E4gKVr8X/l8yJqRWNEuTGH07eCofP
42TbkUV5hEF9WeiCGA0NWihv2Q61Ddn/7nDmFnN9QSvJR5Emre9bqVt6UHGFw9ruZ1LhgUV8UnLC
AdG/vMynfpOj7/WDH9ER8y93URIvgFNHgGSjeuNHAMdY/P/NIArcQu5kmD8MVTS2PVkGxbIL6sQx
50m4W+0VU+g+b8ToH+O3IYtY+U7M1IbrdjavR8lO0wPqtsAvCYw43+ZUunY68SbdVOZFIx+SfZ2B
0ZxDqfNgcp4thhwVhB76PTSW3YnBXxfVGPFYvL4ksd02C56oz9Tul8bkBnGKRcudrHpEXgcvkADF
0DBbJY1XkIypgoc0KRPZ6Br5nJ+c7YUoeLXm1qhx0OBkRN/HW0XjeovVg07PsQXRsoP96uqzqqU0
hyienKRRlaO5vUQW+bRXzaK8ioEWB7hyfExFv5Fw4/K62WxzVVLiBTjpnjilwH+L2F00GKE5amx4
pAUtYhruDPVTHAX46AwHIbZ/M9X5bBhUygkab/affLkd1ynI6UsigVfkDuulxSD6jM54z9k1iS3N
MdECm64R69yvHQL2ukdjHX4qMPn7ixbmMZ5jBBLg4j2QvooTsrhIeeBJ6ztRUsAP2g2TGuobIgLW
9jOw7TL2tJLbayGRpyv48iOR0JD1f+/xlSyqccG5Ld9vVjvFDsA27NPgPHENxFdRG/lj9BYtySsQ
JSytreJXSZUS3i7WCP+1ECVCZnSLmW6AG2ejsqeCplCLcL+7Ys3aDN3sJAtZvA00iLLDa186Gz8l
If7AnPu3C5r6tPaYqI0/QEQxCiVupketWhw6eh3XHcWew7m/Js409a777liaJdHmozBkkbtAqEln
CvE5cqYw9sZdcWQ+01BCler0fP+paJf4Q33Tyz4HiN22utgj4x/ArzPuIMHaC2+LFb+wib2Jx1yn
HvZ6stEGnCf6SW4GIbFcgZTChmqN+J74shcX36VB7p1paeQxf3MGnKmret+tIfxhQ1VDrKSBFrnU
h/JBPysZT1zvk23In+ysnraoSXIqlQXYAoGQHWywvEDgsObx2smtFR6hInWuDq0jCB1wzvvdOzoi
XknGdZsDLZf1SB3lUaBw0unvimMMMzxNB3u3O6MzaTItexlRRhhy/QtJLVl2prSSw6g+X1X136hT
QYsOr0Lp8LUQ2C+JdXZtfORalqX/HfNHZf6mlYnTFq+/NMBkgS9+gIhopj21cJjCwQkJLL2Zq2w+
o5iiouEGp2IEtJMllbT75kk6aLhdPaXZQqsHFy7NiSB18AuB7OpW4E8GFB+zPTqqBxj/s927Um6m
xwgy/91TgR3IlFmwVNOSOqcLLiPnCIgN7hZvm4s5zg3aqZRkBlOk9tQueQjTqyCE3+6Q45XIrp5j
J913H0fMM7DxUkOuA8bh0xnaU8O7ZgKIYhIze3XI6HBi8v2pZX7C5J8j2r4OekZVp1kwBs+uu1zZ
8yMh3wJpaYe10FMJ5d7TuRHscKzxM+BsIPdyxHt8nRj4MpXERICRUEfw8Rnn9Onf1tITreVCK3f8
F8LhYnC+Qp/HxK2KioSxgd45oaBDmRz5xn4bakEPwXeD534dZ8xtwEYAfx+al76TvbrMBlxDm3iu
FtIqm71EVnO3nqEA/WM4ALjOMYnuC0Ubqck2B0iPsd0CqFalF1sCN4WJTTa02x8TpbEjPMLc8HSr
tQ6tuhp83JPEBOxM3dHt1IjXYTfsrXZoXi2I6viSg2iWUqJKdHF+w4U9URMCThrXu5AxQzjq4hlO
Dpm3KrKoE/B0l3WQawOQkquPTsyGkWaGxAgm2sFI2lkn4t5Jp5tqVg0fI6hDcrMIvFOG7XgKte65
UKBm7UEPo3dWcg9LZbdhVVZyc6sAQ0vtWVinxZc5yUeMYPKqFjEeJoylTWbr8RGjl3gT96mS0uSZ
hh8h2ZoWojRsSE1F+qvrpHVTBZNL7MtJgvvACM2O7vwuMh44mmaOWZZf/excFkTOYU7LXU+kljul
m/uY43ZQbErZH5P7mRD5cznciZ6AK9nMrQiRGGVhLOAhss90DqRgClO0coY2zQr2uFmZcMEIbClF
0rAqg72leegvBaVnC3L2hkhyjs0g29bEFb1P4BqzpwS+2NpC9A58s0BeHczWF8PemJRTzkoTaaMd
ZN6wEcnEgE7Ln58Tv/4nlCwHurQNoXAwjFCSvP0LACmu+Qb1wOfUcAEI+6HoDPbCExXLaFPGCLOR
zCzZcRErJamgn7Jcn8n7tR6s3aufZhMTQmKCZu7B5pnZwsPU9NmMxsbAp9D2aASV+c+0uY7MrJ3f
MfIhVFswcUFqRQEdAEhGhdYrc+Pyw7LzdExWyzBcG9r7E5zGS+vQKe55I+Dka9d2KmRZFW/fF+0q
5ZcKI+B+m8raW1yqI+4B8XrOzja/2ixu4qwqu0zDqfawzx+XgJ0bSkbaJRuveGcNaXNfIj4WnSV8
JqaEUA+zRK9uqhcljYgFIU9PuRJIMLvbSlNEnhjvAEPeEq4qwLCQUwqnqiQqhfloAPWMI91PUm4b
/VIK3Oa/gN5KmFpKiYoinTTFQrAYCsb8z7t3Fie0e/v3xkfS/C1m4Z+tvPycCfnwc18TViFClNAW
8UFJ9H3GntPxAJHmpWEpLLwvIa5n0Dk+cbK9A0uXbjopDEM5PSPh1T8WswLZzAjPAhF+4FAJJx8i
+5cCvVhGazoXomM9SsFLPObimN/I9y8WY3Caj6PE4nix1W7jv4Dh69liVnmy0pwpdQUkDUk1u+Mh
BXCkwAwUksVe39o2ExF9rt9mu29ctSqd3LO/1Wp2Qvyr3q9RMhbTUtY/8pVp7Bim94bNOGJ+Ic64
wY42tnbiJdOhP0EiswooBUiuVcfHyYIIx5Kwy6x0xSMTjKNL+1Wb4/MC4eUtFU0ZbcYLeu0pOvBd
kXmERyZEe8MrECaucCTCFanhDmXA338rPor2oa932KpetowCkk6kZPY80uNnVYUFrxmDSjGi6erH
7+a4inkUgCyKIFL2kRE034sScT2f3XgswW9qtgYEwk9t76Ls5WO53fD22U3xuBMF2SmsEjpsEjOf
rwv7D9IZiu+67jRdl4eT5dkRfA9NvQAR215oACPOGTsRrLO/NitaCqfqldaWH0XV459R0z6nMcm/
XJyubZoCOVInDkeNwAitHLhicGUbvikMgAexuQpuGUnaGPGBsStmFyXBaOV8Ai7wov40xngMwY4j
E+/ESpq1OVgm4n+wjEY3xLP19614ul1YjWSVxsOPPnciQwqe46+L1nltwh5zHoBRMmTv8SppUIuf
TctoEpPirzzErpSJNx2AcFe94Fp35vtdUUnl3z+RJZyiOkWrfeK32yo2/Ggo3GeR8NbzT5yGs37k
/VUT7YzjlOXoI5UE+D5YBuMx2VmNr6dZfYsNgZ35PreMkmfBmOCxEgLc5G4Vv7pPaNyyqsr2RXrD
Mzu6/hyfAZSBkJnYxBijaamZGrNf05Gfdl+YbK5jBUhiW9kEC10Z9TUkeMHowgvjeDW12kgbOOgB
XYdqZ/ufMK/xFhAEHFsKPml2n0nEmdBBr+FYr3K9xTZaVHdorkqOofezx6bmF12dFxfZY2eUd2ZF
if8qaPPUToV4XZEolbolpGjp6CrVqtISbKqGZmGYRcgNoU4i1yB7/kg4+CablQ61N1vvpUxggB50
k22wG0M2Dqg0kcA0LJArd6zijokmOWcSICTEU4JsXH3rYytgzGz6wPCnsM7tPG08jVM0/0RvtpNQ
VCGX5u4c+u27LXVRvEcCjlATU2GZCf0uap4BbrjVqfZ6wyJa0VyDl6zo4Yfx4ABALAR9w/prIrLC
H0f4MQhBlgOu6XkcX8FlCTtUsUwifq6YIUpv992jelQ4ibtXKgbPoGxnJnuxNccdYpazfHyYIm8J
fSpM/OhAJeiBX4f/4qpNogJ7RVmQun1nUp2vBR1ajlnBgynJWueuRISN5dmaGkrehAqJiYJicBoJ
8Lww8BbLSS8NytIXrjuQvW9cVQKz0G3mVnAf5XKzIpCzKzM6NJ59TjCUjxpM0voC/h+OpNQM3S1y
TBZ1q5AjGRtCdJszu4oiZmNAwpsbY3k3aijt6ep/CdOtW0QzORIru/mTB4g413gkTzPSUWBDLrEy
7bFs9BJQFkNAwvbOGNTTDvR9RbA7rXWg82b16H3U5gYIGF5icnLGcz0LVUei3G3U+LlH+A5gLuii
a1EWoDGaq03RAFsmLEJImwe1HZchBzYokOBZmlAbUXMwriMylcRIeFYSNqwaWopFyRRi1gNIG8bx
Ejoewq2CIB9e/yViiYXF/aWfO2mcXt2yinWci3OgW+E7XxGO1y1V9t9mK+j6abbzSqRLUKkLno+V
B4CCskNTAz0bMlvzQx5BeNILfrdtvi9iGLqLpmfccNxzbs3p2vcP3rmCBtH0j5d0rm4c4x4cE4c0
ELj06lw/B8s/7a5fuCrCYJSlqogwuHcEvgSmPQVhirLmsRWXkFQxYfYfmNNR09kyFxLoGf+PhsE9
qUW65d/iAIkUH6MGGMOhMsFCcPvFLtHM319h9wnFsJI50upjlGh5Zxq0Q8/1srJYZSCNVGXv5QE/
TU4CZyZU6Gq8JTVCGvXhrznL0tQfYo9C5FTwyo4iBeMCgkPb4Cs54VW4LvpRlEyUsWKUAVENcYT7
7OgDySrvwWt/xiFfCSXmjDx5AED0BNdOIyTMTTATzx3v9YClIYjZ1VqR2pKdgpF4moNd8D/k20Ne
4L4MSbgsePxz6NJSE8urouenhZqI5RP2juBtsHCD6sWmyp27s+5PsFACutCfEQFLjgTCW5n39uSi
YGEZWRhWL4cKxx2omlui5NKwbTPfIAYLS/5kmqPNYgNDBpDkNcl3vQXNWbnSXZg4f4Zc9zZseBlw
EhFeRqKJssMK+H4CllgNj+a+GHxZOvUcMyk0eyMV7VXHHLuRXqbMTjShaxJF1wHE+6HxzwY+CLHb
o8Yo/LabFX4BzT0rHIF8GH0tw0R2tcH+KTqesnJv+6lA68cGfgVn0sjoM9OFTv4NxnJcdfUVXc/x
ZfvYNVASw84kqwSNHZ9dk4M6eHTW/xc1dSavQURXZ6TMyw3bk/vgADCVxB5NuHf3OJ9l/XbRf0JC
Hk2HqZDDG3wRxa+Z32cDCsIZWy6KCHfwjsys6IhTfFDeNBZFFWESwYppUFBWX69+maWGr++QaGc/
GtVVXk40OsSXlp1asRWRFjJiATHc9Q380FbNwZJln7xLSYbSV9okHPnUq8fzBzLB3pFJ1ymvaIov
BRfHEkNll301R9nd52XEUCzLURD1AT5eIY2fXNl2vvWhM15Pgv7aAGpkrDTK0rOeiv5kQHNMYX15
ao0+J+127qBcNOdUXrJsXo5CQC3X2sWF+Yu8+nEN2e1BY8BulvYILZgrDXbHU/ykxgxHbtJqqdVP
w6qAcS++Ta1yzALIyD1+ukhOUy0MsiogT5pJEqyUaLGisB3/tSI9hlrkttJBp+VwECs7HKZcbyKV
ydpMQOAUk0qxR78M8CtWje9L95vM1Flr/aq00GaROzSK7lSlicvIIA1Dm/FCTg+LHXnU6dN1pzUG
i2LA4lxN6ztjO8N0h8qE0R48eU5SCWLrqQKiPtEHUhhIT/LDevKIkNrkhTl8PyuGzeNfeWrTBgc/
YugcZxAQqTKonQXluNb+zRIrpPyDhZKpAomhMg55aawat/H0fTB3AQ8UvHLQlelXzwLkG6AW4uoU
57cd0nRhM+4ybubTFboAa+QOQnBsHNdNZaO8aBE1vsUnbx2IKjYlZFCRZABDcro1KYiTzlFyI50S
B71t0PDsn5OtgtW30QvPpHZrU9Krcrzc0P6af3Hay1FTI3LWMr8eAuOvPlcv3xoXscEybN/QTCyw
egVrd90SlTubvr2U/z/Uojn7y3WCXNsOJmYlrbbLtAzqSZl1H//HqYS8hFLDvlULV7N24WA31lRJ
Kh7rxgwOoiFfYVrJLHrPEw4NICE1YgRGAIiFdb9smRIkBX10TRKO7IepRU74Ew6KfjH9KCXDTXOl
i0125hem8zqKMEfmcNJITTLtQk68l0hBPWkSdcGO0kzN3H7YLtOmR3WXDx5ryn5pHsnzI4dbm5ZR
jj6PpfdJIi/Fd4gbK7JhmZ0v+f8+Y7/ZUAaFn6EHn0G7grNlFhYqnWRGbg7UAEr3Wal/ymZN9er7
5bbkQZZStM9pRotQyNGKXrGuO2/Ul53DYDgBPjIdOynj9mimLZycxSXiqmaHsVx7exyKIMe6knAo
jbpHZX9Y5IQASIdXbc+87TRjWWoqFdkYxNAPE5RlgzfjL9YHBTOi77WV1FWzAC4YKHioXKbVrI2N
xFDKYWCqeMA4UFXc/qFqbXOWV/EZBCdqMws/FqnFrYDTJc81kA0PQwcZS15bgSaf3+Dlkjfhb2p8
qbTrWiKnqxewhnh1wu2XGXVAkz2o07kfp3CCOkDCFTYW1xRmltUByn0k83iscOtNIXoJACRqo6mU
S7r243aybVTX4UioXPA19/vPcYSdXuMnrTHC5ZsCzKOeZDOymVFcMYjMqybQOpMBrpocS1sSJVOG
IQE0wqeafUcNLfuzJmUwKife+2pFwozXl5IvPFPxtFcUDTGL2rABT47bu6ftb/4lUJlg7ZDUV5Va
VUWBtFfSIz9D8yF4UUv0sqe6gwNXDcanjBdUP9ZrGt573NX4pRREyM99TTMqUu8bOipplyGmmN4I
z545BS8fC7Fvp+Q6ERRw6Hl27TXHN+UXw941/x/riCIBIVoUwPZakQns59fBWGcUYmc4AOuPlbwn
nSatglB8XmlxtH3NLzWKYnfKtnTMlR+QnPFl7K9Dw8AvY+rWZV2FXUOygt+p4s/NLx/cOgUHPDh1
SOm8TQojQh8aWvuODpFhAUbo9vDHXZomHkNJ+aLFMepktHpI5WnITIGj1MKCafUujX0TfrOnlwS2
JDA/M3Rj2Oq1slZt6yDEJo72HLk5Kgzpxoa+5Zd6P10XseVTiXDiqpdnMWY5JKbZhkT1Bc6gkklC
u+MivVS//MvuKIojY6h48ACl0NU5qqiRGxlz5r7JET6PcdWxY9vIlFtL+I95IAJhCQQjfdDBiqEO
9qXbPptCKn/+h3pr3V5qWn/hL114h+LcsbCnxWZNKxPaAI5bZDwTUV68scXAeKWvf/uEUfLGWdhM
Juo8menW2o4SWRYodHKYuoqC4Jx6IckFEZ0leTcLPO4OZCE4LPATiLzycwD4nzk259GNrkVrIMrb
EIM2/anFHdV6gnsNT9A1SoGPog1+B54nYa7aSd7q7TkK1Da/tzxLgEDpHhQqwpH9aIFDSGIAiYao
gGj7WzGK81VkoQQXntQ0u1hr06Cmnr71AdFZAZw1bP55J88QTUBXHsf/Tv5iUj5keEAF+y29xWOC
hajAWE9hlRXn/TgXt4JyZiBPwuRiscfgTFI6GFqXucrmln+Av7LT7waamNHRPe5MxLkDpu41lygs
3F6XZPI7PwqgmqSu5s7/CY882ShPAuzkn3NdxlH0j3ypgBybJJXczafhnD0ASDALbxDE+VtuY0to
UcaCt1NSDoXrwAWdzZJpOYqMD6GLLqjbFz3UrLU9C5+5bvBBS5pkXu1617lX6bgG/1HP7it13Oc+
dbqtdB3Y56IRhTcSjTgPNgrHjlAvt1QhRldNfddas/pHIofrZAJS/BcjXeRMnbZZ4C7Qj1P3V5+u
Lv5Ydzl1YRN6zUeFyTh6r6CiaiCQf9foFqVFo5T4H/3U5m3GCNu6l1R17QfrzliC9bvQ5SSk8Z21
RIfKiJGGKijWdBZj7NbCIfpmG5wIboc00mQtgjsU+WVI3KrfjjpQeq+BBaKDnROwUEIGGadXKyU8
8oBy1rK0ERi3RBzIQrOAkNvMPpWTobw17/sCgJviCVOuKD4bLPaMqlFlYPEQ0xn0TX/YZCUR8XrP
bVwWPh/xAl11jIH7SZwmPQQF5f4lo7q012msCeeGWZiWXg8K0LYu4ArsXM5jkIIjTCY8FHBaG1Ml
jlJ5d+MIYb6xRKCNyK/dq9AcAuEzY+sq606VezbPrbTFfBk4V/b34fyfZeF1C+xnsYfnfDx1FBIO
DHfLN6gRaNC1asoAH5aDgV+pgbdUdr6eggVknXW8oiuruZ6iq1W++Q3V7eLfNVl+ERsdOEympjBg
OeHUIleMvkRnyUsl4qmw8UO5y5r5HN2E1foxfo9tlSu8SYuW+czTUgwWNdvB8UrgtYYO2S5axnRr
bqZDT67OJ+BjbbcASiPcRfpanfUez2v7jdF17U+JFxMl6Bko4o0zFmHWouJao0lDdbSvQJS3JDeX
AkN24L73sylCina44P9qgWR9itUX+l9rtqCVfJO61ZgGW44Z43ZaaeX9rHI443F0I6KNRIbuMxpn
i6C03Xg7GKEmY29wS7fRbZ2L09gn91RASSqypR4Sk6UGuY0BQ67Xg2w5hGgB5kgPXorj0uMARQGo
PqKOJYeU3pfYPKUhTjpctlWyTgo7ThvcTb0LxlXE0A4j9v2LwqZRktLYg6fte/T07im8+FkIBPnh
2FNIKBu4jnoH6KlpKUftRKna9392dhCQYH9ZZ4XN9Yx+VfX1ByMcC87aWBcbkmegAqv6hZuphv9H
cQArwZEeEHmHf6G4VSjuMGB3RxmO+HBuJbVcbrRpTSwVMKGrl/iFZt3yXck4ZMNwUM2UOCv3VNzm
6mLmX0JUtoDeCdhSLEfuCmAGpYqhjA/iMRRV+p5Z5/Xy+kOtMHuW+N8pYewVsi4gTxtVdbSRx4v8
dNsAOGHy9irwdA8qVztUEoS8ayQEOwBAjFSZbzyhQmRoY4jl2bjNzUsN+AVqoHl1W8RYxzF4z8HR
FxjhLL1Ur+hjtab8uVT1ArV2MkmYMyu2J/Hqc1ZPH4emlf10ZZMVn+H4nQpIKFyiaF80XKSdVWlO
oFSY9VcGqhqnShRmftO3Q1yOM/bw/Dfgugz1z8VPAlUUh/IgN2Bo6LS1s6GO/HxN8bskky0eTSMv
ZM0tH6l9ROIbSb5E1Di1KCwFBhBkvWcOJ6USjTKaaiqElIndIzc/QH77sUEeMx3LDmArwdLrekU+
L7VSRlVIpzLKKLxcHMQj7h2MwSO9MkTS65ZwSBdafWuyMuMCXdWFEIfZBwY30OWJNX1Xc5Al5PLk
QQG1N0xFPij/mUOjLv7//B3OMKbrb0/k1KO5w9HZuDjHkwtqClFyXX22fC42zu5/ozhepo7pQBKU
GSgYn48mLzdMcyszjqJin4L87DU7AnKsjqqC8lF/Dnmcs8EgA6ErmzIN78fa90wMd1kyewjc5q3K
f6FKR1AxV8DAQrc9O8AAjTUz3Tt7/XKhqiRtvgtS1ZYz6Q9WAe0RJQpGOWoJ3QLy8xUW2Aoa/Ev1
PVjT5vKL/rOkBIVAUmzZ5cIUvVCO4Cagm95nczajpwNjdcaWTtrirDQJrGj6TjKUq4/k7Ufb5+gg
3Y6lAdng2BJMnO22ZbbuoqzXnJiQUba4LjgqGVWH5yDymKq/lBfinfkRmyv9+wNILmv4Xksjmug+
G5HZnhbBE1z42jKnKNrwyTJ8pFsmSpOfxXAbIxe7bslMOd+j5g8wc831MmkenQE187P+2awfQXub
33gikSbxP/v2OhZgK/QQEhqV1dXJQkIGoODZIO55UtfvSN3h/2z47CW/bBaqp5B1UEavG/YteZnw
FfoHQLu2CFSIxHkePfrIrRL1rJvI3G0Mmbr0Y3nniTHpOHNRc6feUOXeNZsoYF8MVEeyHAX0t25D
9epnBEL85BtBnnCgpKTcTN1g4xF7CGfMnpaOeFHcuC6lTkbWUK4747M/Mje/HmCgdtfmTCA62Vnz
Ry+/k2MZIo9/UvhtosIQ4gf9AlSDLiunwBsn1OJs0WWPvmxdJEKNXHNQzu7W/bn7BcfXNuWNwTxs
/nWYhyr1QzPlZ1aD/IVN+0ccr3To+9HpteijjmscXeXxsbkqmpCTtS605dHUgQchKwKj78upjiog
pYrGXWODv6LvNBpjWiT4k9t7QQjXDxw00S6kDRvYN1qsNwKVrSgS7LjSmpknkZXhJedgSSZKqGhw
I1CByY3DAnCFrgjI3yjQfdDBZfGZDbNmLgR7FID1vdalAKDEB9ywqGtUQsfCg0SmaREcZ0FTeOO9
ZWfST90Y640O31a1SwxYuhMIsLrsxGXCzJQUqMTMNtc39NLg6XZ7kQTOVPlWoSIhkOaRLXrQRDsq
rZygpQ2STI1cjVr6+Pg4UheM0Tg1WOpR1qXMpoJzB+wZsZt8jpWkZ/pPmWFB+ozymzQwDFh7gi4W
p2RCpJYH7ADNGuXsR3HECYXZTI1oX2epL6mu5kDkFnneRufWVOhxABrbnMxpNHcaM1mJ1aS9xFmL
MTGiPCpP/7Nvips6urpMOrwvoRcQ4Ks+UMD7epZQh74Np2FjsbHNfaJc1DqmqByN9+q8nGt63PXn
Zy8r/9YXygzEr5TpSGMPuU33UJqNwBRWDn4W3ZYSeU2D6MseUPZgk6fThbyOCZziICTOilw8XhqS
uN6qkKPJFverrSWutS09quUOHDT9TgN5nbpVv37w8qV66AfTxrSurufzwFU9ERVwo4eP4i62PTyD
eM833IZeQfkvTb6vrI1WfZ42HMdS2AIUdiloJ+HeIe3lkST9SPqA3ngwe0VVkrLGJiRSwSHXGJA9
Tft5PzjWCKVaSDy6wZOgxlwfL4JBUWTSEufr/krJOYKdzssHyIS4v3mGqVAkIrISBRmwP78rE8hI
KhrQk7ihG7HSJGjVg0gq1KLFRgRNltVCsQiluyMb+nF1WbblW1dN4srDK/E9+bd1cxcfvyYS/xNp
3Ux6odDTDKAD+ytXZ+d7jU0az0s9SYFC8ZuhfNw2yrucVSvWB++E4kG4dX9tq4WB66cVPcGldH0Q
2jbz73O1m+LwngGSBOP1MjGDOZMtXuiPt6T1+u4K1cFztA6eR8si9xmw1uAdZTedm7GvO/yQVIu/
Ku171/gvnafryj/f2bxbXxEJqVdOmQ8o9Ds0jxDMGiS7qggWDgdUpHFL26B4kGqp4epQxgsB3iBF
Th6KBLi8L1p7m+1qJpDqvBGG70IFYYSsxNFNhmwDAJ+TzDl9ncjO/f2KZEncl4JP6cu1NV8reeMS
IWwWOuRnysZOOda/WcQtMTQ9u6ktcprzaJ9hZr7MYYcnAlkP8244RPULdvwf8ugu642pgglStg+1
6i+LPl2vyXdEmQQM9cCSU6iomZryrMlUXv558g7cOctXGe/G+hf8BGSJufnDHrnD1nE6oN4W4yKS
xswFsdd6tjXj8jflcMw2UbgMcIzBzC8aDaW+dbtcAV/faO33+4+aDzbjeZQ2czdaJUYZsYGldkSn
KVSBBMnOd+db/XotjB9Oh2Hml/hqQ9tUnJ4kEnIpgA63jVr3jEIHw6izLzSzoQKzvxbPGEF/iDdg
FyrcFuPNZvp76CI/a0WaxITVdQt5vyAiPxs7yg8xWMk4UAvgQUgls4LQTS5hVfBMgwcJhaAaOwJg
yh4KSfRJ10Y1RlJvfx5lT7+LLd06xFfS+q7WjsldgIQSOMhfFmJjiewdHP3yGBQlsWOvMVF5cJE0
MaXQBkbxuLhKzQGhqdsmJE4IG9CYUdPf4YXV87y2jXy4eG9f6M4Wv5RdX4YcHisDy8xVDnM7EgTJ
jmeCvBes4PWJgB38DIBgYBUZzov3Ys31I45F6FiWptQzISROqO4mQcl2yyk2nTJOUSqSfenFQ4fg
PGf2YsQv/Q3Ch8f+MTMfn6nAs5GQJIVg4HEugjZ0Gzt/zAUbKN28X8CzK5mCaO88KOV1DtT/Z8zX
1L0KcpmQgVDYNyFgREDI7x0z8eWDM4ROjaasVr7TDpmjmkUlCuqJNp7Ugj86isYgAcuy1jxpiMqX
8HIeDKvX9LE5hIgLoNdHACeciJa7oQ4IYzTFHiIgwQjSSI4uxGsXPtAg+p/suf4XzNBhkzlMa3/4
IVaenyVcE/mjGZ8WZYr1I/11dBwzmAsaq5h1gKFVYWQxhrcfsTWVXTJP/Atz08qUBU1TSC3DTgbw
RvKGX8qiYy7wjBeqt1Ow4+r96f97G6CL/GIjD9mK/pdJv6uG3Fg1BO8LCFRs91TkID+X/zuN33H3
BIhCz5QEcTz9Nnk4nX0j3H2v4r3RLg6sybrv9K5JFMFSje4kgRk/q4IEU4Cg5zMe2dSlnUX8Eko2
C0BkAEOrftxhtcS2pnE9vFFMHKcVnNNg2s1fESMtl2sgWd2/trD181jbac8/ayBkh6K24sqLz6o5
G6t7yCch+GTB+X+6z21yUC9fT7+aZBwLhJrJyS6Btw9Wv2VLbzzQTN408qZ7gPNhCKFHkWXczbr1
B1/oeOzCLqMz1u9cB4H49N78ftEJ+f0b0RH+LIktI0rs1QLEre0qvvQSIcDhAC/R77ypRdyuz2+F
cLE1Prb4KSSOwTHxk2gFsh91oioU+VEvtJDDhrBGRFTki0gWDrRLTck6+/gP8hxKV+cmGzT5TYso
jl8/JNHL2h+WCoukDJhXNMaFB61BQVd9KVPHMRxccLz2MKYtcws7xLPHsdbPNEeqt3rC08RWSr9U
4OBesq2WJh/PEBEEetHh1NFyJftDFdzliJydZNEUP7wAWc2zNGwtpBM4ujp/j8Rc/tsw0XHSnXwM
7Gl661h5Hi4AzBOwCWQavU9mNuygAm4Kf3oMyfMYKJq5lBDKFb5PwDg4hv8mwiue8FXbPMRa/HGu
MuF0b68lLH8Mwb6+YUwOJgYjF9Y8kFW8hKYFwdsqzxdC2s8E0WuiTAybopPZ48iYJ/drHf2UYqGC
Hm/g9owpMnG7BvLmOxPJdP871oW5vAA/Lnozkh7jOjy9OvY/OsGE+6w2jyqwboGVcy5C9vF/xyGs
BHkFG2lH8/bztfsrazD7IlRhUIXRAgSPv5xciQucj7L9gRZPSyLthclzaUbyIwTx6RDSx5sY7tou
XAP8Px93R3W2Fr3cRPLQ/4WsDcU6S8dlv979oF/mKE2GJBo1bz5VqSIhIm52Ix13MF8dnjLtzqZV
uWS7z2kjAjUc6xSec+1tx8jzqPd2yQD36E45n7l7o7VXuvmj2Zubv4Y3q6c2/ItvkBxb49yC/LLf
NXzI7KZHVPZnYCCRJ+4MVYq9C3TR91IAJ97SUuHhPQevz5K6IcVCYpUZRn9WQ0+GoyYCHpjl/UZb
tn1q3Q24UwcScfoGxXkdr426Fu/p4WaLk7rR0h9AsigriQJtjd1RXFX1CqbiFgzIDWABS484wCII
Xj3u8PmJ88k4i6YpIlnJCRcKr+CDlvNNXCiHe3G/dE1m5xx4Dzqz3F/0TUELNPBFJlHrgd8D2Li7
xS3Hc6EKEDEGGbs6ghEJylKIzbiXcAZBunVvDmr/6oAyC++OMWkqi421nC81c/OeyP5TZOigWtb3
0rvC16CYumZqrYizyYdhF1GUrmj1P3Mzy5Zk+eQMA1Q598eULyphrhL45MvVEtWjFybhf+HG0C1W
oPlh7QAvD+PPDD07dL8s1pDgZT6whJuqIh+cZWBJPyW8owxCtTXlp4B+QRRLu0Hp52+xlwCqIre5
v7qPqA6lbz4F97Y+aUYK2S+yLCdak4BjYF8TKL58zwC/cQ9NO1RLi7M/oZG5nkdDZv/pkTXGT3cV
hEP/yKaWrTjy5iRiDBaKtgaL7EIyRpeGNDt7wvlTIoQmZjTsVvkKnULV6ag9uaBbaY3TmZJSd8hI
K3WvECjbUURKeRRBBEHNOsci9jkGhshuIJr2FwPgZh91VcDSCJ58/+CyxLcNLHma98K3iKPbvRk4
wswUid+VHmIqTrY3EMVejeOVDfpoluKgpRigm51qhPgRNsK3a5OKenHsx+RFeCbi0V6YPppzxjlE
jpSqbXkq35dQvFdieb0ieHtOmZjnyrn7amOVWcQMFKiQxUOqMHWpdCR0zp/2gIVw8hX6BA+Ewt9d
K0YjZl6sSbrSK2UVx7XfankYKXNRvLgcvNad/iWcazwY7zAGmyOwyTgHBQ47uGEdxvCFiHP03EaE
oQGTW4xh+Ux3gTieMqBB32/WBZQnyV8UqhIYxyswW+do1wccujWntduCAqfBnw65iTIkpK5gkBKt
4TH8YIZlhaz7iPcz3V7dDXSNCEGBGuZuIFqG8Xd4GONZmRHRMzeb51j+Wkcl+fuZjYGzL/AjLoo/
3OEvCE8AuvsfDLF9yOx+ippIP/4tio17jmvyi2PHb6fSoqkp8gv7iwOz0A/uEPBmN8YErWS239dT
YmIb1QXxWX4qkUl/gnhJUDdbHK1CYw2MklmoBAn9zZEvd2pCIwFBFUaG7uBczNIi2N+Oc7ITKG3k
4iiJcRwLiRdT+Y3p1cV3hVNrrRU4MThEjNkiUUqCgHan5zzQu8vK6BT2EGtsysnYJTlCoOEacRuD
a2bB+6+R06pPUChCZQcPoF9UwJa1DbThWYZnEWazlnoH5w7ZQLhMiBFP0ewVo48IeIlQcQSl0Fh4
NPJyHmo54byBrAFTJAXpbquHk+msOSP7x+PYPGysFppO7aw7K5vfvu5GAm0h/GFfjkC2WeySg395
+oZf/tyaVq+kT1Em9KPmL+OUV3XLDWupE1iVYB61Wd1bn8lWDocuNH9M7XYUNKDndq/SGOlpXHn1
5G7P9TDMSTQtSifEKPPjeda3r/yQxRDB8KR9wOCpEVp1/VZmUnT9JDv3tc4NZH5eXdD2tixUa+ME
tsTGxgDg7hJ+f0/1AJVkbnPIb6+h5llarvmrNjbuTTum+xPaSOoj7tlQfcu+1pAfY2jkDJpXJXZf
L5hL5u1P72kOogyyZRjgaYG2rM5JR0cFRZ+LeMWsqMONzRaS2gdQROkSkQI/vaWQLbI1WFzG5l8G
Nr/bFMZdr45d987dqc8JVPssghy630qEuLvsNHYz0q3lddtco6wyuwibwURRRZ256gPaFlxm+zTG
LLhPeNDUQibjrtpFjQlS5LyOYtDZ8GJNttAikKp9ZlpFhuPnHCoUnkaXzO2GEwGZ7Ju21oxLWCqx
eawoTlu9xXt2DtMZa94PKMZM6/pMZwg+zqPuEgK64dl9IMpMgcV72l42CszULqpnEI4VcgpkIiss
j5k/75IhMyeXVzHnoPcJxMVbw9hVlzLD1aK6zpG0QVCYP7E2t8Np5Twd7L4ON/rmKl+U0qWDXirM
5vqRkijt5URKyGahIXxf756ywRasiF9im2JvAOwmECpTto0Zq3KGZjK0GIPmjw/ZLOnAikoiIPNP
4xWztkZvYK2P6LCTsqRhl5WTaaO/nLXIA1MwfDJIJCZ9oh+graBcgdw+YCjofzV1nc4Rfh+j+a8/
/6ICrDpxSkcsIXOJK9T9cVJfIxZzZw1+WZNALszNZf8TFO7ojSjoKV/QQyDAr2y598W5kU670G2p
BWy+JA99XemCx1RMgXe8vOQLiYUmJJA6xp/uSwKpl5mojFdDgiGrwjZLo/GDOjyXImKFk+iIZox7
pH7hOsyBZN1jUcX7ATxHTUoE20ExBz1MPZPF1zRDJMSBcX+xwmEbdtYhccE7NrZdRviyufK1ViZi
5VXVfBFUCLDuZh2kYhVMOlt0RHf6+FDSjBk8AVyCEigbxmqOhIgyfFpFVKB2uZUntMs/WM+3hWVO
nNrokCs35yEvaYM1JYKft1EHOyw7KZRYw1AqoDIYhu/FAFXbEMYzxrJr4gy7LedzZvntKS0LF6P6
DSIhhkBk44YgI673tuIsnXQTgmZKywBABPJKGzGALSBJpefvQ5hNumKu0d7tdimVFZc7wcI0KP0A
WwszpwQgVhBj2O/KpVNeMNviQXfPn2YNio5UpXV8rlF0Lc1jGrqkIaumUKAssjrLJtg6fR7LCMEa
+UY4qpQLSuIrx22TYdCxypG9SjD/p5ZoncVyAokqsnfEb6YiWAycV8DW2JIltNEhfrU3W4+1kfYc
0jDjytw66mFzOeYZPr57Z9qqTeruqoyj5vtkUafZLAVC+L5yKBh1Kc6QJwB0iwNGRvv6fAtaQzP1
s6MV8PIXQksAh8tNUi4rT+HbgWp6yT7G2zYLWl0rbI2uKkgzmeIgtLxj6PzYf7LzbZVM+e9byDfI
LCh4bgjsHwKK07n5R2b2I1fxsvB2mqZTsby2rLDs2aNrPP8uHm54DPMMs5hVNl1kcN09ly8TGl12
q9Fp+e1qzOxOw/O57zztFKcQYnkzNe03umlcM0K9LUgmUklD2ddO++OV9qHv9k4Y2w2FpfGJYyyu
dVxhQO9hsWv74IKcNLrof506kr40/zRdVWbz6OJtTeO24+t3CKqLolv5auF3Y3Pbjh3jzEZzR87v
0xctXEH9KzYiiRjDt9A9Vku0tc2flYmnS13iXp25gkok35pqKTENjMFGOoN0itjK1FbdQIK6kK/j
xEqW1pmlo+Edk34coYJ1drqVH8Jg/+qfD2PmwzWifmxvndC0/j/Fur59Ns1YKTpMM4iOwk/Q+9eO
xnSm09IQoZaW/m0pJGCrhT2gfhnHbONwncXHInYmO5iVH14C/xLeSaH7FWvCH/AX163djn+Wqder
tsgx3AIiYaalGsQlPwizRkGsHuzknu2rkkK4F+5w6LX0CKZPMOKh4gEXD/2zhOC7uDPZ9ae4VCxG
CD+3LXxHwNw2Afip0VEeXY9J5Khe8b14RcrKBKq8CuwXpvFloVDiwwD9lRlrKVaHhvFn6zoE+vdM
J59NJLr4uPFj7gjzSkexL3Fmx7Vdn6+i82LhJzW3hvZAiOxRiE466CU/3moyludsNEUOEto47LkH
63duKZlXWeIvKS9KOCyA1hexJdUgrOcuEEk8TbrrExOC74esoGJ/vfYkIeBncxTFUlyvJEEWawIZ
19F+0/aQKialtP/IIo2aZepGtPdEDWwSACuaa15wCOFHWjaXQvHx/OW6nd25tvY0p1r/gu2JIxjB
JBzoDdLRkXdxGLncfBTi/HjU3g1akZGmo2Azy5KEdunmqHmbnReaUNrw/z+usZsm9YgkVHq8i61H
JRLLzp4bVv5TCKIwsDNcN0z79h7Itqm6GTo3qLLHR/WPaVbcq9Mni6NjSU7jLn3Oq3nOwWDZRKQH
FRZvVy68OsuBcPlacI/cx8mk3he8DQnLSCCOz5lztGxiNynY4WF/4jNMlzifE11uXpJ02Aex+AAC
xeoYP9jNNu+8WN/3PzAFKoQ8uuY88LS/Z8lD24D07Pvf8gjPLxt5V7GHnLe0QhVVmx2fs4tbgZh/
UTayC0UkQ6xbyKj/Er/jkTklaNtLB7RhaKes1HlvLc50j6cM6ZwF80++DhWzP1+ii69VXxo0G/9c
HJdYcajSfPPi7KufUy+BRxYCs8Xt/HbCFAQAdT4VU+Z4a+8t5clLkZH/m3ZtqXNpLqET0vWrD80p
VtdtbHERMoO0GOOz+OcMYqrUDUIRJlUSQMuzKW/F30KcAFIzhcvPhkoHUJnblQ2mYfepYtw2KhhI
oeBHRBTRcE2E+Pw34+PiaOeAO7c4KgLI2L4Gl6FNaeT3KUQZWDNCNvZbAf4H7qVgPT0uXt1gwIRx
IhOUYAFOQQv9oY2Cz3CP5UfTkINIf4vthF7zgGvQ3nTsaX4MXkZEHAXTBbYZN0FTcCuQT20F9Nai
+vUeB74FVq4avZtqEEqGLEj+rqNiIgnoh4uceCIpFQB9/OOM+F67F/6nReabb+BYjA7YuKZWvSfH
3DBFXuqw/sVRox530mkOtG473WssPjUDrlEK+pALw5VjdJl82VZOoyNpWBSXg5EN5KGaEvGvi243
hvJtu8zw7RCIKrDTixDcvhDATlnh+1kS76G7pWJHlkbua4kVp/2YACZbq0eURJPHB1g2YhdCy/1A
cxXhCQS89MuzauU88Hvk5bRgCFbHf1bqZJ6Ae+ZMmg97lvjvGSfI5EXUG5d5qxsENQ1ZDZexMCwS
BdmIXUBXHdcp9ROrWZtjSq6HK9K5RHTSR4nlWlHGK0f9+Nwj9gPTIFk4C1vq+im9qKlJDB4nRedu
mzaaNzkhS/Z/iWeY5hGy0FDYONJ/ckmz+80wjudtda3hBbcJtMpJGC3aU+KEUa16wa/UKC0Th1vJ
O5zMjOtAgtRTEQVfCbWUj9dXJS0yo7/yPvgKlmOJ2NJOHfKTgHLTC0I7rWtOKMCDv3MM0oBvFl6c
JNTloPyJEaCGDHg5EWEu1xavUSUTyC73dfPgCR3wwc69D7kIWs33irJC0T28qlj7CFOXUqTqBRNl
zznKRUhqWEr4SAIhdk+F39abjPsyrjS70Jd+gJai2PLq3dQWFPEiNEpr61Vkq9crohkHiEFwUymF
T9M5nB9OIVg8yoPOR4tjzIGid2hDsxXAPBhc0Hjg9Otg37vHuenD+INd7FhE0LvWfqow8kR/1FiG
lDQ2LexyKeyhHdq3D+Lu1/AXxwDvuNoDmNzmHJVg4XVF7O7GG1xmE7xpf3We7AL/COpB0JjkCerp
9otegkUb6nC6YF/JshjW58gojvX5lcebdzlnRaw3DnTgewc9ZG28J8se0RTqpVOZnYcuZimQII86
UIuluD50it0RYzjujj//yb8CJjBknhlVxJd+zh+wmSW985Y/0+MVhDQZlHeymgIE39ZWFancKgva
1VZg+DX0IYziJyLsB3kTyCGCfHsleJx8RZLapWjEAmnIVFXDbQp4zQcU8HXdiL/eNktlRae6yGmV
+E/0yNgOlgyVC5Fq4mNQCkmL5WX02pg/eaGOBBt8/wfM1qUICNBHZYOh6VVY9rUPlEbFSILLwVTg
BVbRgYp5mgoMa3MYNJO3EhsdbvFkw68WbO2Bp0gx74sso107ugLsA2wZxbT5nG9pVYSqRBGcEizr
7y3ZPG8T4buvASE59ejeXNtB32cBSxItIy/RzB/gM2NZVhEd27l4o690ESK2BUJOg8jaHQ3jJvd/
62aZkMNDU6FED4Bm559Hzc4uLXBcO6KldGfB2eUjlevv4zFrC6EkYxTMxBZPgBlkUSL2gRRcuhd9
3XGlc8+aZ5iz8/NExDCJxCJOiX+KVHu3RUQH//50qGE4wZ7tumqvIDXtv/xlFQ1VaoXQw/gayfU4
TedP8mgGwpX7CqnU5ZQ7Gb1ZwX1rcYkascjQ58vlp7YOKqgH0kgbrF4xUhfejIxUux8nqD3PlBev
pilj9jj30a0NolAt6p22ssqaf/1Ru7snzs4AlmmPwTku94DUeIZeAHauUKW8Hrbgzg7EwnuJf9yO
JgbpacIm2rXaQ7+Q+SK9I8FiDiknvaggPoscZ2Nkw2YQ0qtUmKp+ka5bIegZm7dIiNFG5qoYtEuz
9e9HSALh3bbqGnjo6oyE7l93W3rhriEa+T4+Ff4lXauxi9q9WJDGu7VhkJKOoNgaoE2TYwU9O6W8
bA9zA+Tewub4OkCcr32fy+88KZ8AJaPi5/GWy0h8ApcWpqqVDFXxFoOp9Wjezm6Wa+1JLSJSqNWz
vRR4jcN+PDun1c0J0A5UWWDCxJNBd6Dh+6TGFPWBWQUzJsyhyHGKf+ePw0Rw9TyVQjcTeQVTRDjv
92IzxAaCXvIw/6mnJWT7xVWaPYYcyuyy1YsSn+i2HQDO2pM/3JRkjYhyAKEYzlawFt1LNIDVNje+
svvUEwss4hsIAWRuZRVq2JLybfeZln6iWXpxV3icJYnNY1Vxg30muEoDMFlqtauDlQW8lab6VN+w
hfdXJy7ZXi9ro7uQN66KasKAW9Y2/UVz+kKjyh3iSam+rMWNu+BwDSAIHvLAIBjyGIf5xDYN2CVP
SXMlZBK3YeOHOotCtGiXA9a18jnLxhwZF7U+AY0LPJbyT8oNy0j1SvonhE2174c398PDoGPtgCVm
3K/7xmW8PKSQu+A+/C7NOjOWeCbgAqz9W5V/zH43bvxHK0m0iPZC2igtgHgPb8uotyeJa7Lh/aRj
SNvsNWcjlPbjKqNFeuw0JyZZqtOZnmxUfDH94gGt8CWwA6tTIjkaghuT7KK42rlMCoqEQTWz20+1
6YiFt0rSmlPGP97ajUdBj0E69o5LfIdm1G06ogUxcHO3kGIrJd6onETpiCbSiB9ZlLfOPlJVJiXU
7hS7SfeOQlCf1W+CiQH1E5SK7LcjEYnlBLQR4H7zJ/E1PCYBYeiviSM05w9IauidyS198viqfgDm
z0TJT4/YKxsGZl4V1CxnfhR1Tp4lZCCMELxS4dkHMteLnFREp09pAmVYfC5SYAuIsUra5mVdNODs
yDbEEHVY6vA5Td3Z7+tnGXYxC/T2cBz2LlZDBGFebDnV3eTE3hFaHxZKt2J1a0FHVGUch5D20/6K
INMDT5WXivhmvbKSG6GIFZBGEVVS5AtMmbDoM/oR94X/MJ/NnJcly9mdCVCu8/WDRIMdoU2vbiOO
MmQJen8cMIsGBoiN1RrKC6zg+tDy022MBJIdb5DqYpoNvlf6XtB9BZQSloT9fsZs1tgIEMrVmD2d
agco1QNLPMIAx6Ig/3hGpNhdP7CMAT1Go8NlRYmM4c0gN/Va+akKj/gDB+uyAiXWHVn+5pWhMHOd
HeGSMQimQXTTeJYLo/nmMFa57GjmJZUyNXDvyA7eKOeZ0cPzmDcVbmgEvzo5SDzw1cddP/XSk7Fo
d6Zu9fUxOIGhax47CEeZZsyVxomILxAcnjd+xT6ZhKHDjc9BXQ47+CfHCuiRTYcwyXhw1YCgxiDY
+t3jTvWZzA/N+B6kP7K8mB9gEgJcWaFg0AIamdK0/ZrOypu1WNA7663UOERLeLvoH2huxpCUb9G5
V2Eg3DFjsSdMIeCHJDCLg6Y0uAqhB6evmrHqHwB9y7Qh8BDjy/Wk8zfnbqkr7Oh1+HjTQ11XLD7K
VMac2ZP1Cv/2LgQnG+191RPI5NB9dZwO4OAEm6+jsvaYCzUi35vgxprLM4jKic0mvg4yc8jFKCVw
TEFT9JxQX2flGvdzcrm+SL25pyk0NJmRs2cj1kBePJ+jPZMRqOgD+408N9Chv9T6xUeIya1pxqoi
mUljqL8y/bboCZNOF4SE/nLVO2espVK+QK1DK3UOeIzRyiDL+Ve6CPacAtbHysqNyoo6Pjzis0vr
lwGouw5t51II/Yja6ot7L3DsRlp7KrOYSeMym+asdJnQDF3XLMHL7J3TU21lVYvMMML+AMBN2eM8
92XVSj69cWG2kULnWzUekRHUOKx3ebIId0ckyDkWwSBZ/Y7hoZyAjgWuAuT+jWjqyUqIVEPj+Z+C
NTm/6iOw00UnaUK45AFRiISTTSNwLZwr2nrrLLMCJTZOfs7KKljMG7NaweeC/x/uWw+hGqoVENau
N7BxADBkFzIWDEnipwPfUCwni01PeldFiYsBgmwDfWcNyvTNY2RFVgimO1UAZIdQvBk/9SFdQgb2
Bd4Dl8eigwJGi9AWo6m8CMmbV6MaO9lyPKJD4/kcJRXjb0Zxf41hB40cvgVt+gVF096YGGNrQeYh
+Oo1NPMd2Quh1VHYmwdiNekgLAIRcdtx13ei+72d3XCgpt2UnUTYBRoQXyeY4KwmuYRpEkvDNCzQ
LuKSo4qjfehfYhMBkI3UPBQw4KgZR5P5LGk/ozbCRVeqxkT0BjS1sXo5O9FsZJanvYtOCKVdH7nm
aH1kq9AIyNHMddoh356YBss6BY9t514gghHXO8k5/juWSK/lsmx9LKk6kBe64AqUOmKnLOWRCSzO
Qc40HTog4jJlACK1ULP4Y+O+7RqzpE9cDjjNOuJXFWpzypO5BAVQ8HK95CobesRXezSq5RsUJN37
/MksZH53+tJb/h1/RrfhKlfzc7HvDV9LaFhvM2RpFu82C00y50P4WJ584L9CWx+jzGPbeW6Llt34
sUG+mv6tTTpiSxiPchBl0XW3VvSgep7DEVTj9YG5DNicnp/Ixq29vj4HOdHUx/7tD2FRzWJU7OLy
jNMJhSpsmUo6DyolXIL/4dVnabea7dcDAhUxGAAoMS84GHwhS9P7ZiSuVvieHskh1CRY1mVB0C/4
dZgfJWPxAIqz//A3ywk3n0AMnLbbDHr+BLHVDou0tJsHez7+vzidRS5rpcOaxV04k2SNGSuw091/
CEcsTdrYwjUB8cAA286jpIb2R2+amCy33RYylJv/av4rYMzIgOSZFCyCQMO5Bq3CZUNr4sxU3HtQ
Wev9J2uO9VgqhX7Ezvf1Ia3zjVmxOFkttS+zF2ywwccDH37B9WcB02bzCam+lPSU5gsYs+jyKuVa
HDlIcbEirB1EAisHJhaZA9FopdFEZzF43Ly2M//DAjK0mIB5gNtcNEWyOsdcSGyiGPCaOqnRiC7b
yDsh5zEi4ilFzU6IuA2J5fvdlMyY+Q2pDL/YdSuaEwmopUs26rWCdm/gGERN+tEsg2DCewLLOlNb
Oqj9GeCs8gttsjyAmc92D0Y6JvT/2qOPBf3hDbLw6TTJiiXYeW0/EvZ9rt0cmi1PQj4sFhKni9CK
ZhGiA7c9y6NfEZK54UkB51hUM+DvLpXt2R0S4lgYHIWZl/8ss5iM9YjY+i5dgMVWhflmN5dMDkZq
yPlcpv+yN60IAZxT8tMJWxuZFJqqa/1naaYz3OFDyqoT5/wzXEpbgHiKe1h1nLrTnb8as4heCiRL
cJN3GSaggYDT0eKwBoKNyxRYZMtdlniRJwk1LPxkEa/FXAAMswxREQJqMuO2rI8V/4fXM1YQ/aq5
MhAvDaJzf24UTTVPdMYfhqpo3SatTLF4fsNk/9iJ14bjEmO8lYI7xG3KRgwIS1L0E1NAZNn/tkqy
yWZbdtCNETS023jST07YsIQEXuCxtASBCeL2/TAGWimiBQyIWj8Ru9zc9Than95usjoKUvo6FGQb
qn3n/PBL54iKVJaA+h/BXhFr0Br/5FV3e8+l/bipSxCu35/HcqQ5tIHbF8tQ1G8NbpT5Qp2ZNKYh
C4vno6ZstcICsQPN8NKPARof9OjiZPuag/r5LVc4KjKBA8aYWbO9PdKZGJzTaMFPIddQea3dsUr8
reiA67WALLtgk458jyvUyMK7CLCKQtwXRkRNKz8FVUJjUQjtuPjuPRTARaV8Gm3cSWTJSCd40fml
FDMbe/S3Dfzy5DDei5J3jJKdkRafV24fIDBBLO5YQeD7y2QpFg+2+ld0RqGLzYRtpEy6wDXbjXLA
/62pMRj047xL3oCVcHj3rTomZpNWvKftV5mLFZ9QxGMWh2U1BMQGB0GW46V+Ql5Z+OkFc3pN8kyp
lfiBINbavB/JuoNd5jaKZw+ztmnQYaZmW3u2mmOTAvRY7CtDEXJBh/RtvjUWSYeUruUc1NnmGRRF
9L3smWAvzC1MMo1CIV7Lb0KGGsYRzolDzEIi2HpUt9hvpGcLFbhRV+lRSOTyoItFZnM2crNQXxq7
ZGrx1nwdb6MlAdIXctjBGx6ea6YcqnlnPL1bx94vwcKUvTHOvcFzjapRDd35HM96IWMd3aWlII+g
ywUxr31ttm9G7TgRzPLAzQrDWSzFmM/Pb3Ef1nkSK5yQ6neabJNCpaL1pCihfggfzVRyhRww06ii
NyTNwpV5MCxF0BWfEroDLKGxZHSISshEdBlsitzIpibfayOWdjhWggjIcWl3eLBlrrpTl9Kj20t3
tS/SY9UGLd8Jk1dxgxwVseJSeX0p5bMbgc3kA5FbAaynLpMOfnuC18pZl8R8L4/LokpdCGItag1t
oBcUVSAgXqX1E/yroFrnvkvbqwLKroi6mCcjagywwIzf4/E6y4IptG+3Pblvkp1aQuHXPXa2Bqj2
22Ns/ovq2Fxv6wHT6ooEYwP+Po6I55Ta4Eyb8DUszlLBLB2cvn+fPsM+Z/1n4uENWSBSQdfUTL1X
y2V9Wt4fPYQPDVy/TLPgicxXDMab0WYRym2U51xRpNjiQtmvrj2D2QAS4Yez6FBl5nEbOFQw09kZ
sOjYcYyKuhsQ0oTuTW4oCqodbt4Pi51zvVlUnEV5raiCAIdgl1T09eM5/H7TgDN7jHXMQ6IVEEeW
Rc+uAqfkB0U/PxNpwW3PGrwVe6qHWqqvodcB0eQBgpZTUXe7O2c8ofaSs3q53OGaYEPjVycvS/cg
10TMg3lpx4ekXRwc206Da2aDJq7LVZ5FierpImqZuZX7MX7mkJUC/XigFgDMthWUn3Yd/0DhGCwP
gUi3LeyXX+FcmredvhK2luluOUcAgGIfkRmSQA2pxIDzQa1EP/yoGSpEDIlE4HCIpF6Nai2SebLw
jJTESwREARmLLCMuE+fZL9cySecodemqGFk6lmmYa/qO+NG5JtB0Na5/UfFp8VTNO0gz+6MDEMzp
Uf82ePaA4HGDbx6GR2Y45u+x/ZbNmyFbk/mpS+yYiygDWC9Apte0Zx8jQh5ziEP83Wy/8LucqE5b
UOiK/tfvIKDIHX+9jk+Rsu7pBmfi3oycGF0FZ+0BEak8GMV1VGGFqRen53wJ5CjC9Qy/Hl41qqfi
zgQyFgqZqe+9R6YEzwNSP0uQWqviOa09a8yaBsioq8sQ9/oHhW4wcqpOtuw4J7gt3ApZEgwb+5hd
TWd2wWoh6lymvuyZgiEN3qq2ZDqV5pL3uHGgae4qz28T3GKDHwYwa8PLOqp7wfZE3dWJnj9/0zWI
o3M4Do8ecDU8WtjDh3TOEq+jYZ9aGsDruoWBmAJi/SofrpMm6aP0kCjD/aXzlE2t7XuIJrhUP5Ds
UHXc6Wo5MNMqx9YtoZ5U3jgk15+WhmlbQiYhiy/MwH71N1PIJAoJUdbizQhFoiI0eoceqALYtI26
ujINvO8Aw9CgbGnfDW3nB7gxAVCjrf3xzN8D9bdrzLrKeP06rz5fLmdXgtmiOahXmldAUHZmDSwj
+x5hH06R9cQg1wo1TUPfb1lnm7fp22uL8QhTniZiqhxf2vKL3Z+sxK73QTOFLg07ZyR87N/j4ur4
P5JiVirHv+wVHYKXTH5SZy099Jl0mL3nb4jycYnNs6xYP60gCREZeMVqmWAV/GmO+mQirnSJFqSh
yiZUTYuikD7mq97yNjbJFLNIA4VRygM4Wmzd65qePe2nt1vEuKGaaCgZayC2yRiEU/x3TQi0OCuX
Dn96LoHTXILnCaGJVwZ9lb5vgRkmvMFEaAyVscB/bZEoK1J4K+C6CIEFxWfBpGIifvTzZaV5gGKS
tAm3B/7xg33M5JaMmWvufkup5fKnaEuBX0ukMJLdQXUOTHudmf4ueMamax+zKx8UO2hk0McSj9AK
aewAEopYgvEtYsibffaaao/52joTlku9Zv1eeNU7xjQ/hIIMlxs4ySOiRp2sFIJXTulbehOG1DmU
/jwuF08pJVrt+uxvwHERiZTrXZqTvy6JSKkXHqzCnQv9k0xTzhllAJFgsdx3FYvaaY4rNFeUyE38
kFlaxv9eEG9+6JunCgiJKgi9n6UJqeJHgzgpLrk2olsfIKXKhLigFSNrpdW014Z5yEPVruHKthX7
zPRoeeIHZrZbKPLfallijs8l6PYbzYlvq3+TQlwv6lF9CqB319TS5pbaGNom52r4vT/pcUbB+KXL
FrT+qD80iO/v3MSBLq2skJVLXIuoZX4Y9dfSxYDsiS1ckPnh0mZuCS2Gk/HBY9QdfpmEvbPgRfN0
2WixV2NIvXHUWxDenT889ePRuqGIO8vKCa9aYR6eY2AlMe7BAr0xi54RchRxCMTbO7K57vulCN+Z
VM1zAzc+3XxpA5ko/LeURZJHU0x0qqLGI1hz0W0N7LdpMTFRzg9SJgNk2MwaO01WaEIft5lEzy/h
YhMiRqcI2ypm9jSpF66TyVsRJi+wn3FQZ67cwp2A6Q6rZg8N58uaV+vQB1zH1IL0XHH4lpyD2JsW
0Y0erYNbI0I2XNcboMTr8ezMjpA6RhSyZQAbAjEgo4eoKCyasGYhV0L5dB//wloog4lvsgy3xxYI
X2GtpDdi7eMqQy9lNP85QYnX8WFwXF9N00LjO8acJp5+4qSwiujO2ng/UBOFIBWs4+5vBqrBqxUP
4fFGhY3ae/zMmYA8hhQY/T6+bSGWqVJOm8s5YRgejEKcuDStknycJXHG/JgrN+8sy7/oukOzKbP2
xK0QIzpz13QPHMhcukHrNq19Cw5QMvb0uBafI95QyOh615enFCcKPIEf5jv3opUTnMDZgtOhN5dJ
pZzUzZnHnEQ/Dr/HBZOje1MuOUlhPPTj9NvxxEYPlUrt7wECo9sybCblwxlbaQ4/SeMO7tmzd1SY
3vwtIWVtUynSIi1fcMNe8xwpp81fnqRrdxYsT/SAA3FO7Yd8EA3KmrlAYU8gs7xt10CtFtK47nEB
4s3WioaA762watRgrXl4rqwDWWXCGBTpsh3eGtItagcUE2I6qWb4pV2mINPeeHhVRz4Kzp11etI1
QK1atBKGv7U7GBtUw7OfDJjZg0zqCBehqZ0Iw4ceYAVNMZdGgj32s7XvF+2qEyu5VwkNNt2YNf3e
wbfQfiisjE7TZNqXAZD4ymGGNUC81ip5vFaLr1wO5ZN0/gxkYfHXukQZ9vnjTwjyWI6t80BrbKcO
k2T7e2Te8U5Yx2O37vF4exIdsNyo03PmX8Xq/iVYYFrGhclDtTQnpWQeeICpJlA2jnm1CXHAYwes
cbbz1h2jVW01v9NjHHq+4VnyoeRUsFM8dxN6fl9fwC61UbZT4DZ8mnczyVLyEfwu+lyVtyd+qdDV
9eSTJxnhAJp32/chjmHXqm8k2Lw+QXjrkDrStLF+qMRSAfA/jYv4LscGeN1lQaiO8Oh6MubImQ4x
G0pEru2pFbowPzB1E8SeeI9sfpEkjSxL/bMaG+J7nZ98+FuTh2OYJjnV5DtdHdMiCY0t960NpESO
A6aurBj1v2wncxFYUc7xB/Wegii9MEkYv6qgOs/gyoY/rHvxy9BGOGC1DjJReJQoO1EhOXPwtH5d
/fifeR4oG8cgdiLIRw4R+MMYcPp3cp+IhLN4Qpo2gxZYFrBZ0SzxZN9iRF6LnRI4vAweAQSkooUP
P6AUx//e9O3FVNhNDKhmD5qz4YGQzwUp3Ma4yl/kLeIkBCjrQ9uTqGtmdQr8TdykbKtbvIyiJt2X
AGcC4q+CRtWtFBSJuk7182TWXwot92AWxcUeStCvAsVsSmvI5ks93mJjdSFxxol6EEGwjwrslykF
414qick4pbKlWNMks1ueEhGWnTfYpuznKanjL4lsAqEuxD5lFc1iETruexoMtcs6/3yogAMvBiGD
tjSbSNScu5542av2VGAnpP4GRKNNsCc/QfcHlACvQx//jhMiBGi5CZ97QguV1NDRkHNGbHOSHC7i
+nI/v82Thef1nt8+4u4vQnGh8LsTL1gBGUU0IceQ2RPVxAyLxZkG6zwVtmoxBzXwQYrAw4xU9Cj/
+SGq6OhQ21IB+o2CbvA+YVcUvA9zJBz8dK3vAmuDGZw9VKj313lYhyTlbodEcPAKfWLqX5dAZdmq
aVCJYb1ImiwP+jmz2jx+xP3phAJAzjWd+4lgH727TbcodsSdRIuP3JGaxuVvZOyxJgoyLVmQIsN5
gwl265RETvDcWtETbMX1lgbv+VStdJ4LrEcSNt+HIcU2M8n9VFaHAelVQNMTek/yEBo/iP9yj03s
00dKsCQzqtrNFtAfISR0Fw232fMtbMPBanjrgWmdIDDSGm+H4c4jtn//zKDbSHY/VgvGouTsO9cA
HCxbCxIpaSklSdwM4WANtMTufxEUP2ogCmFmy1V1YeEHIFU4I6DnLu5M1TXN+DJFGFXkJw6jPdxn
e6I54+DbqvTtDHm2O7UY13T0gAfyfIbKU0PsMkwTh3Lxk18nWKeTAugmyeG6BrNMQRZlv2wUYX2I
1lMQKuWFiQ6/Phrg8m/smKZppQGvcydtcsmETviUqtxTQCJbGRjv1/v4CfWsUPGBHFfKicN48NwJ
qluGJlRHHpemPtF4m5zB2il2oEy3zQQAJAB4y81i/NBi4fVUzaNTjqMDmKSWvdILooCgZm2tml8y
0MTGf/2t7IiXWX9m/sZTTTAilrB4fBsqSbaXdWdWCSUZmGHm8POdZR+I3hOlv3EJZ6PevDZk6qTS
Q/bD4dIh/NYcjr8f+ZHgE7HEYxzKGZP8PekIRJndxEcZT9duvh2zO9XFCp+05IVF3NS6Pf64byGY
8VCC03fbVf6CzDb/2DAcKFGbTKshLM5PpKAGg5wMDpGpM2owvlxW3y3CB0oArxKGEqD4gIZBSEPg
SQ7iyl2feKoVC+4eHQRu1BR9S4VF2cKUMw309iWDoYbtCqXJ/sSyQqgWIGmjJuFOebAC1QzwB7Is
fLx/BZ2sJHAsBGkaDxvqBhs2OW4N9a80HMvNFR5/ks7aWvFtCveU933FenooOqf/2mR2es1IycPe
45bt+9EyLk+MHwHHkgRZqGPEGCN+BMFqidb53zV9U0gmlPAMB1rPT8dWlZsez/6kkgHXZKeLFUOh
vvDv3oT847aawqKnyTh3R8crywGKCPTXOREfeIZ2U+QK3JU943zBOwSohC4YxFrxtYrIr9romPS4
2d5Hc40KPL+cD7kcACbK97851JXls295qh4M6wsnPWjkrtFhrQoOUhP/Syr6yMIMX8c2jSEllw4Y
Zv86lT0DPmGn8aBb4AzaStKluDTifqa3KmsDvUDbc7bM5/WqkbwmgSYd8MTMrr3Hn0R0hH+ouOoT
3TwHyCHvTk5BYO4EVkV21PVnLHf45qqVOs50Nmn4f3asDSNGkIB3SfzQu3xfgj7fhaIkIO92pZBa
wnggWeQAD9w6NcCtnD7woC7Jqjabw8DYlGMxND4xtzhBD9CRAmTfsDH6OUaZdWdSH/Q+LacdOEB7
wR9o1SK9YGxCowwqof6MjU36HgRoy0TUomvklX1f95A/DdBSWz/E4dLIUXiTpA7pCZSTjmvzCRQt
gTik+fFR/LOA+n98YpFZXC2M8C/zKw6bHHz4dGIJ/pbB2Uaq2c3lTqkyVyrV5qD/onuHBhCkJdsc
Xt1hZUxNAHmg1MF+TgH2osJ3+i51JXDeZVrHzY2/G+0xskRKwbwKFH/ifHOtF6e4W4BGoFZexspx
oI/lFXjzt061i2Uf9jWc4FFH2sxi+EbozqaIlyffn7NW8gU8JmTL3W/8PZe2sR4h3kMkjxZVMs7d
Bkdcrci98AUF6SQzij+S9zP8p0m7SotODlSRqiA2hlFjV3Wm6J8xeXi/ilW2jY+Yp09Qe70ZEaZ6
9Sv4uOWdhE14I1DoVb+ofvyYyiej8nmI87oluVlsIRz+kQDv7dX2J628RWDUWJZSY7fBKAwFcjXr
y/bq/bIcH4PPAaCManweRYDPK/taUQ4A9MkoOjUPKDUlyhdsVVzIet4JA1wjdQVFSvGJNPmUv2Gk
F30McTBu5H4cZbV385cGfFH55Xr06bkuuIpNvxHkV1X/Bz29l9+La1LrA4Z4mK2+r1lsV6vEqm+H
4xAMtZRmp0NYep7hDx5sOYUBpjGrY8TBg87KUck0z+2+InE2pQ5owc5UoJhRb2d9zIsYZTVkDT9J
DpUqC+sh8bqop3g+XSODNZ0QJi6gM1O/ciTYTHElP+crtSbyWwHiPWCSYIvsoj09mHeuyV5zoU/4
CX8brNGk/nfYz/hjIOCt947HriPEetjmeXA8qT/WKp7Ut3WG2JJyLnl7ynLYLI+wptvXZd0jrlv0
Q3C8Hnve0+VLC6ySScI896HppTvnUEOCaei1x3dIVYOwb4RzgPTUk7PtI1Hhpj4aC5tsvl09fS2w
kufh3XCh0ZEtaIcS9xrF5AETI/g2ZRdaL7Pvd6JY1XJDDTNo0X4wMHXMhjGmCwMzbVvHlBibbQpD
2VrU7e098d1Sd+GWky2P5OWdaqEE/GoWNnNj1t0iz1S6sZFWWcpvhMVpJAOEVGgYK5Ed51WdoWSV
EDijchcn+dEl54TBLmAld0DYRX9yHEy4t2cnUHKEesEHczeX8DpW/gK6NTxRtN7omb5SBcVZNZ5P
5aDU3ME0SbiNa0109w0u3KUmDWyi7R19t86mSPnc2zeCYb7oRIq642remj2RXCvGukbQBYejOOuY
77xua1Plkp1mQUliFAPPDMuqKhT3Q3Xij6W9MIVe2kNDTDFGKVVGv9eOQ0WimSaR6mtzc3HW5Ih0
/aO1UEN8bHI3V2zmOQ9Apqn5x8+MpxBMRn3c53cqKNh13Tf6aEDf/P4egULsAq4Xe5KfQMGSuz4B
SEj4j6CCZcPEEdhy0G+/FEEvIp7i4X2HSDIFZkT7+T2QYmmUyy8xoLwrARrWLdzkakgrdWou6VzL
4tlU373Whf2glb/5P+opH+OgIl0TI3GMOiNQep74px5X8n+xxySyz4fBccvavCXAZhJVWXCX7zsb
1dVre5mPIxfyasplwl8rCmKGM42g1X21dl41jvJ+yoeMfe7f3d+kd8+NPhFFzM7vGkjLDtGBqbMn
XOZmmgRQMP0pSrObBcw5BGvHuNAFDEjCBb6UrMm6SwidjNl7gEL5/GzZxhv3CSGdWhbp3YVOk/qo
sA1MDuoMgIMboOqNHDzn02xPK0AlBPipTRTJKzsgB/iBhllgK4qAmDwZM6XHIBB3CsIK9OtClckE
AxvHtdcLdgRZt8sKGVbHy8zOR7u9bKXA+6DFRRvJkPKfGtyHL98VgqdEbo+GAsoH3xo27GmER3XT
fBqhZTKZpJ0WfJEIIwH14rjyJsVTdgzklcfHNVc7MSCh5uADzwVy5O8ZoX6Pw9zS60LJh6iut5WC
XI+sjU2c1awNC7KuskqEJYyPv4ZwwtmNBQpasWMdi9Ienj/v/A98rFe8YyjTosViSfyd69St7axz
u1dYfjMln9K6EQkyFYgAvwm1LdB2ZYAXQg7Uxx5Hns0sx+bIN6kK+Yiew1Ld3Y9d8TuWEpAxkU1i
njkS6zLOPK+E/KFFWIXPgGbFLPpVDLHZ3IqmO3H74DV7hnLlAuf97wFyL7nEqj4yQX/7Gga/CE80
/wehvny+DYcPeqVfmehTvn7lc5mwTJdrMGgt3PHkp5vnP8GMK+zmabkB/XgT5zVV/68Wj86CeQEc
aHSzxzfG935unF8u3glCVGlq+MI7VMIg+NVsalm8DpEQdMjn1k2Z8mXCh4l0z6ydAYjCOkqNYSwo
G3BapM8PQQW6XQGP4sd0lW35ZvEK72BjKFiT9yoTrErgbum0V7SYHgjvEJ5MXyDOpB5bCjkwRez0
uJuW8rxQHfuYi5mweOjzcyjXvulh0FJOmGXg6qQBR30Hwid+/xWkDSFUcvT0NX4VB+GNaWT3Lnf2
t3LM14giyk4kp2ECllR7IqJ/EPNqIH4fEWto0cDo8k2CYkhWOvjc1MXBYk9Gti9jvs93CavqKHy8
sutIdThzk6lYVWpmnuQLj6Xj3A/zFNs9KrI4mIyHEpvU9s03Jy/95UefhCdSA9xD224mILrNyuC3
895NLy8NcUJGi6W+gnAFGJdPMZy3Y3TP9Kp2TCpqzKT/UiAFoAiGidktp5/nFqHDeLY7JNx8RDhT
NmTNnsu+kQohlFbgkL+TB5AifC7jg825AuIKsXMaW/upaOSrKXRzw1HfuKvdOfq9I0MVEhlkW9w/
zyviJMREvV+RvDao+smmUfSmS1Yh8ePNU3Dp3rR9lIUBc+5TjxiMQaFKxmHvohuQ/zACmDb/d4Km
99bpOccd5u8GI66hhQ+u74i3biiy0nsNCf4G+VFZiWt/l0aUTSDVZHq4dbIVkKQZSzpSNy0ylVs3
A8+yOS6GfQscfAu4ueRyHKebT0Rbvw4cL2B2d8B6GGvIpNNjZmI+/q7jwO6TTwBROXR0cJtpGQQY
8iSAXYdBmWWS2ThsOjgS0PbMtEKzD4ymrZNl+vxQfcsLVV4dfxmZjtdyQIhnJYrNA/+xoCi7tzKW
WpgFB6vChQZHhiCAjPJnmiNaQ3zq8sNTBU0zIiV8Q1V9/aSoGcx+Rxg7sCLwsSN1EyNJ+3kKsvaB
Z3xmeewPU/acNtswyj9YVHS6J/YvlKw7qdix5V3obVSk97HUy217CCJ4mFNXQ3mAbPzv8jxyAWfb
WamTOYCUNqK2tW8vTPKduBm+zSpySvzrO5majfsi5miYolfV4Fr37Atx3YLGkerJggEHBox1Ri07
pIQqYAhqTO9zSopVXBTZY5Y2H3TRVdqwaucNZq5gD2Z2mcC5/dDSz4pdwp+AaJik7Co24Cw15Y8B
nSZ7m8lWj5X17hxnTtSrq5ffhZuaRFI5tYwRz3VK4bBTaA/DTZheS8IM2vQcfV5DxZE/mAG56G3I
nRExwZIpXitdsORQTqM9fC95ikQkHcNyTTObv1X5U8K8g240ndo4BB50GvHZramfZXjx7wODu4H7
+lDXuym8PBw0S25NUi2If80nBg8VScWahIdep/tZxyZYtdaUo4uKPIUW961RN/TpqxJ5DX0ysPb7
0+dYJoe2gbFGiylmMeeLdXSWQUDJ6BkP9en0nHtkBabAjtSy+H0PzIW2QfDs0suE7yw6QBF9t/Xw
JJWfSecZDRa+zh30Puk7N1AFHhwZ0Gr2naHCQnaT8RA0RhsqksMhyD0VzLIiAfoAS/vDCpDt1JF5
OuZtjSJI3zjTrWEWd4UfN60DKABEomrkjaeGsFrbUwc01vH00PUOylu4NmVT66wlVfIGehoE8m35
DDVByUpGuKKpRi8Osq6GAbXZQeaHk/4XEcg8eRwkArMuZOAypwA0X+m5TZXF0jjX5/thwj/VRZdB
oVdgU1YVlINRnQIgI18g7pYTA2ej0C1BXbNvDzbKc+76Aa6gBnD4mrdFxDJ6wRIHlcq6GGfuN7tR
GgfzGz2v/wMdkW0sIvA7o/8W+md5IrxBtiMsNpkPzSs8ixFudtzbxxH7gFWAPd3JYW7E/qSwvuq0
7/Z45W6ZpjNErplk5ayG9JifG0ihNUoDzcFR0eRB7nQHEkY7vZ2WAZPdEANRtSb6pJHxSFUxdEU9
CTlPUD9NZ6wlEsZAZ7gD/3Z3kdI1iSmYLfj9dqMA3RhnDFHUkTLAU+7gawA0Z6KV+wWM401g9dQx
mM29484G0OfJ0I7RWHJ0KjzesGGNYVxssR1U3T3q8gqoEyo1sZA6EJkSc1qMWvEDtzhjwhgDdTgt
UKXUTW++49RelOO0PWX5/1WHfVPh+6a0L2HMoMu4efw7KB0eFuoNH0+60zxR96zJLPo5icThjcf3
R42sSha+1KwAmNurYQqN+VPYL38uWSqx5kVDa3if3xh44oMw3oHmRuJwO+80P7iq3MnSWRxtPxl3
4qdvzzbITJS8i6U9wr4w05CMN037tz5Nt3WpNYDJ8ZgEWsLD32jj6YYJh2wGy4aWID9LhM14tmIg
j9jYGQcErSVCXOG0pUFOMvLndKJX1CiUG2weJ/PRIz2s5VeEcnktfUZpDdWhCWd/Bsn7t+NFqQpY
en7z6Rq2uwGVk4PjajYlwSC4jM6eVafmZfURhnf7Ezd2y80IpXV3CwWh7yUvxs4HODDgpsCPkDk2
fpPrElvj2o4YN904ZjtV0Ts1smgZCtGs5TS6KxIb4C+gug62Ce6UGZB6ZkFVwHCSw+TL1QQ6n4aR
EWMFifZDQ6iiDI12j9eIcG7GsD13m6PCQvrjHsC1pQoW89j467PTvhfuHKnT91t8WR5bdc1NPs6p
jBMh6c7kWje6Ewv2bKmyRnqJuGeStusfAxTN/Nzrp6Yg/+3eeVhlCwDU7BnmMy32SYJNCgyKcz05
LiR/rnbAOtqkiER9ABbK+/+pVqNE8/BMuPAy4UBt2eBAxvGDh4ILGq7SeilPTz+jYCO98s+wdZgp
1WcX3lW7rS7Ed5mYv/yFbMKrp/9GuIxQsREIxuZcHhLdGBTixt2a2vrSU6VayAVy4a+KOgJYbYNH
C8HG+zMwizwOuBldZyrXk/Sm6qIbYDkyUIPwUGlpRTFAi8rIqlD89ep1F54f7zaGwev2RBO+U3wz
rn0gV3QbfwopEPAeCM5m/EjPKxUnpjUHWJqnwDLbCc/9E96vEv/kx6ATvFVdcdso458rIN97vtrn
UVfrE+HDa4Yb1n/RYXVOHz2aBFxKLBHdm7jJEIi9+VBP1BtVV7r+jxhKjyLdW8B9iIjdc9+c0NEy
tKExn/0LrcqD/glNCUxO6TiliiK7rqNx1P8qdNkll5Cr9Mx9hkohqO1QkitwH+ttixmUsa3IP7qu
DXav7gLR6Ko0isZb4PKNHE05Uz/xE4SNGuOLX5clT+/oKWD5gnJgBJi8MXScJAoX0LmAQum7nOho
c/hdDXjoPCfYJsiMhDHoP1sAw5mAtXHSKylNKby0qmFHz5egSMA6hPDdrDYiLNwjUYombamd+zJu
kzLzU8wEBmSsgrsBqNdBFrajGZWJKTdkf13oWYoX1es7MOdltWRM8HvwjVl0Np5YQdTi7d19PkiX
+KQubXgM98ewgq14nmkmcucsExTwaPmRWzos06qfO3Q09XWLmFxchgWN0L60EMWZPlBTSwJ4ndsW
UZdYq5bHUJsTyFN17r3qO28RPlxllLSgv6LQVDi9OPRqqT29qsl5kee3NvBHUgIB0zETOrpvotZ3
Uh5mM7aQmUfs1kIRno2S4t+uNiRpdDUbNcl9+UPSmBTk0kFzqLRCKQ8zvntT4e1kyinNAYovK6mO
nKAg3oYxMWEru1JYRZJCr8cw58e18SgXnyFjhAgZZ80xdWacY92dl/s8JmC1x5ME12nfIKba9Ve4
raQHLniPU2TVCgkr91UgBzXN/R1Ew+SUzTFiVa+Q9jEcVahEMB2fq1C3VhkgRROeNUiHCf4ZjT9K
UIy4EeG4DPpsBshpzi7WjL5wPY4SoYyOXtQ2KJWlpjpIWJzvRxyp5JiCEwlB/uWAY0MexmvG0baB
bMM0AGgOYxNy65ZU9oQRYXcSOblKvA1gNFlrMgP+T7Owu+G2vqIZmujkdTsgqqMsg8B+iYR7leke
CusW2F5w+VPMO7YJ2A8Bmhik+UEoYixoAChmxOkvtpHve3PcjCuBlCYZ77GIvc3UOYcKR2jbD38g
YU1VCycQSD06pC/u1Vq5zu3YSKT9ypsK0UOiWDRP/KxAqTV753c1tC8P5I9THSxIRPkUR+S3b1Qd
yZly9MowUEsf4/4emlcbIDrCPxgE0JLIVZwodt5MlylcCbMC/rRSh0TOdc6Bd6EolUQW9sNV8g8x
8+uDbjOspS7WBviEdQSGU8EKoP/pgkteh0DEKjuQe+A3K15DkyUTjEKYTRmb/htHnsRR8odPNiY4
l4assD9i9HnwtKwCmepYLO0N7RBJ+HGW5R8K8214ZBMBeT3bZmvyGY/S4Hv8MTc8KhdJpkY29izz
0hNVXrPOeT8y0bAwNOSUHKvdDV685GOocsUx3+OSdDnHrnt1PVh8zWgyffm9ZMIFB1wOubFdhlos
QI/ZfJU5ui71ezTPd9z2xP5Sy2+fG+gu0K0mLS8q+UURyENZh4pFFzCzHjfEC9CczHH5iE62caiv
ZFdOGnxdUku6UtBrp+DqaI3Ky+ee2Mh+4Ez43dnGQdzqDmUiXHTFNw7FDtRWkpK+rwJqC0UA2/OV
ru1LUYhch7S3Aoo6YFpYpaaqPmzdsoM+SkC/QgR99tPGkCHmZiymTBn15/0XN2sbeoL8IlbME1WG
HqeQBuEtRTTL1mvLwmO8XOT4N1tV+WovDlyhq73ZyskpPyyjgEDpmk33UXpAaf/H4sSR9U5l8VLc
z7bC51c8E+E+EYN2bcp+xa6Ev5gjI1bIMIlqsjcNmYdl5QY/tkz9kv7VV8ch3KzJiy9ruGnNmh51
rUEGwQb/add7+1mZ5Gm65cXuWsxp/g4/bPOtLSARye4awh7eM5IBev286uGYd7co7DgOkDZeJrJS
6uQEzkQHVkGS12Zfeo7pqMZjTpCBv6pM6JNrZJ8uYomJr3I2ieTFVt1y2lavqgXaP12IbHB7ksWZ
ndf0w1ygHz/+1TxuCRrVmKmjQU4fCySNKScLQZWUOnKz9BWtM9mXbZwheKytBU/Aslky0Kpf0Z7c
xmyGkpYcUIxR1LLgplvGVLTzMmZvlt6nKVVfLoJkV8YJ4wgO+ZDSmkPA4uTMMO3b1vdwnJQM+Dij
wCETp82K9y0rH/ns3OdoEvhxF5DQRUd+2yFvMAGKvEfq/5NZfnOucIi7n53/SP4vZMUyJKmhm6Wk
CcbKfPmxBEgINYsxtWS2eRkLcLurdEfJzq5EowpGqbeQmfXuvRnNYV+pSxmvHwcW1ILFEdbpYP32
2wbS6Q9io8zuwqUSFAxBtdb/+tcLtMJVJU4RGz3nza6YmMEhabFFNXaF/iTbjtyhvdrVA95HKXT/
AL0Avg6U3HLfx73moOq7dLKJ66HPUPDoizu8crrPVo+/C+EXHrc0GMW96L5LnWr8SAYqI+x+k3Bk
O6OflIbrjd2M30wPjw5TnSRibikpjSm08t/rNfQN+jFz6obrixBrp5xUpr+67XCExavq6FikUwwz
p5zMe6pBV94NHZCZTCnWSBQecQ4BJVcduwyGbb/S9+fphLzwG69uKu1vCbhUYmrUGgOA7QN+LSUq
wyOa/FSTE2QE5Jk/VCgk5yWc9SMYm9oisB6awnG21B4mdVkXyuyEQ8rmdY918g6GKjZtHBX43Iu3
m2KQP9yFvR2qwOl2/dK6k9OvJTkxfdX3ASUyiVzJ6NtcaZ4MHEDml8DP0ZBY5ppksLw87gRt+1ox
tTPshOG2D2/sYxUg3LrlwjRgrZJPyLb/O4Wvz98w7hUHn7VfGY92/2sygee+SNI7wiOFXpeRMC0s
Juv2MZFidW91ijR9Fjv6cvo1wmUvKaHB2n3ON4vTe1EkmqUTovjukaTFALt0XxT3rWKKyshJX8/s
rSKL1yrYem80GUGddPeu7kLrEU4lU5ZbtQxaMwBq2QVHkoUW+NeASoZmqn9Mv0Th++SpLYBT3Aar
P8QxnxGgwZepIN7t0n5W1bOgiiDzE2lbNdGN5WkJ+dwzLUF/PJSLGOUyd4GSKr8y3Pire7AvXIfs
yxXYOR3Gz6HmQGfLik1DLs1sLDkQ3Os7lLaW4+b5aHrqaQwIA/C9kX426j854Bxst4OMcuz9NV1N
a4K+K7Gy2kAN+Nipr/Q+FT+N29nFyFcoLcteYqU1GnlCAePWaw8YXY1aqZA50b2Epe8W1Z0xQicC
1mZOzxEIxx/nbqSdnF96DV9o07Bu7xRosWrcZ4hZlfvtf99nSdvbKvG5NXZCwpeoOKrW4IwIbGvj
/Bo5c6236EuQp6OJIN+kCdGqFVuBVQywIBsQd13rkP4eeE9bTZxPhnetfFUTXdzJD3RGcHyX9sHD
MoxkrcRW70AhiC+bvxT6PW/qVQ73kca+U0Aj/4W9VCZeagHgSwZWGH8dWWn1ZkTQMFJfCJ8aBnph
N9LGMynblmUrKUfk8nR8LMPBpDOYFgOWHIzQZK2At2BXjrfCC3cH3rFSOFbEEBT8V8UXD7B/K3NM
2cLcIn2m1Yb69hmyiEUUEukKnqf9g2KbwJTuvbEUsxKze6eRyAntkE8xbuJJZSX39mHDlBRTtipW
yR1QAQbV7jmNvRuu21DyUF2z+uNUPpjJTsNd04M78tj/Ew6cteJhv+glmB/S65Vzydz4S+oy9gfi
1B6aDNfvmyRjbP63EdFoQqzc8ENILunG/0b/+Vhd1VmSioek6NemCW2EgmowxlYHZyMum4lEuEFA
/HzO8FZZVwU/MgYH6oa1VFaBAeFzgxvo0O/tLgzpo2/vndE5mLfcopBkqnWulj+IcZRKhNpJUEE7
1txO5gE55kTYdEu7ddyOla91U7FocnJ+EisGA2w6tvMjCqpf/HtoKEX9AcqAnpMcnsYyZCLWuFxg
bSQhBmUs4ZFmifpLPFNbqvarZgRh/3zONt8Vu1jIsoO+wiyBQ5mQ/ZDOXh/+DkmaRyYKvAbaJ2/9
+S3E4x+1hQ9O5ix2hJ7G0DnlrCS/MKojCgDguIMJnEqmzDlGN4BVlbSTABtMUpBwqEKX/yFPl93z
bpr/FxKu23MQ8ntL9JumgNrM7OjPTE+IAX3JEXY+nPNRydIw6QVkndTBFmRr37Vdr6FPJ4uSgAvU
50RjHKo/R3ZZUMXVlArS6i+nvaTIdx/abDE1mdQ/2pAuRJmcuMBlkg+fGACYPbw/SFbK3giWzQYQ
BtLNv9/tF1L+/w9z4I7QsxqxgRtFnMBLj+xK0wQJ6ij/F2fp+7xwGBesdJZ1lqQ6iXMIh8nhwpLf
1AcyTlkJ9ypdOWvRJz9smTCkMvH9u+Gt0E1nhTCmJ74B2Oh3ezBhv7gqU3YsfXkJjJLnadk3YTFU
7FvRmJxp4GtAU3Ys7gJKHozvBHngfIae9+ZrFPsLfxtnk8MJFmLcUhmN6qMu9eVRCqB5WTerIOrE
fQKoUJ9Zz4oPFbq409CIkaRKITbEx16BFiBqwwz6FY3Lj2QbrwkS5P4ZBdnrUESV6eaSdVKVwRlK
KqemsPSPfcLMlsAsWswA3lUyCzSK2H6iETewZ52aP47rPoQ860uAQrwt418N/3/Byc2xh+9yF/jU
qtpJr3KhomuM8T/R6yYeAfitJDP/bT9OpeG0cKG5AHVwf+nFRDw7uqvQ1VioB/aralE/NA82sJ6Q
w4o0IJfEWP/TlzVPTfr4NkJ7jaw53uTW7TGwyoizQwxZGUKjsPCKARP5fWL1aDQHSCvJ9VUTbVJU
c6MU8zsVEFCVvtiuC5yOurB7T6LGJb0zwnAp2lqu+HX0vQZ5fC1ua9TdZ9G/ThBqCttEif0UPIze
doVCxZQzPARdjDacJ4f1qfhEPuY31BBQY7QPfqzZnINlPvAK0TdfkRxtchPPfQ8AF/x+9IJQ/TAw
wDDZoNnX8J6AyNXe4H6Nc+CLPq6s9ntC9Pz6XSp8+qoSXoXfJyV9U/KzDm1gbB0pa7HJZMDKFjvK
9R7C4irnpbD8A5zp0nuW61DIBC04t4RnU5Gy+IefBg+MNr+869naD/ZUdcs0kp6pSRFbIFtcCg/Y
uWXHqOAK+mjuFXTHRfORsEgKZNCDFkUs823hnezSsSOA/JIeoCoMuyXP0U8Tnz2JwhI+9gewHWGY
qDTn8zoQ+vT4zAVgAIy/7rq3KeqkuqkC660kLdtFnbxGXrnZ2CvSHNUrQiqsEwAd7OJQkDLcnPu4
jWZCjBVjmSPG3VgTHUQnSdJfivcyn4YbhgcR879ynnFjmYxTYrEbwQTWZEHdXvvIOk5OrRHgVStw
7UXig8w4H5BN89X/ZJcWC35tUsFOtCd+CfQY48/+mdmVeHXMAHVF9D9Vs/sW6lE/1F+OkoH9Ur0p
3J0pISUIh778BRVlLkrVkOvsqMLgukk+OvHJSsjhRqe+/BeLKxiSOLdd8PA3Of5jXN1XQ2aZO8no
PGqKMgQoj7xeJD68fqRY+4X1qo9DVIZv065qz6cvS5QytK+GH/7doRb1Yc/qVTKE5E2It83mAqNZ
ELiPl9zcpmzvKoJIjdXgCn7hZh3Xh14KiYh5dIfCp7HC23hKq8OcvWGFK05XrsL4LTE9xuSYOxhy
vi2Hopl7A9cEmpshbxV4PJfaxv9oxOGb6QWgtrF1AqrVejkEJQaZjZigmzHsWRkt0vj3ijz6UvnS
lD8mTNbfAwY9LuGjKg+RaD6Yf6hI9ZQWBHE2DkjDo3MRImeQCcVmjFDuVzUcJe2Nnr/Um224XKI7
GgQ1cKn4Vuf6dsg7wVpTv+q4/vgs8SaRkB4Jwr5ftfe1w5xqa5fqwiwehiHU/6/eAYhLb+/UYhdx
n/nQYxnrvrN8ROYlgCiJokhpKJGtGnmajzT0es5ON0Quj6r+0MRdy8o618le6ZIT9t1fSCgKIOno
bOu/JM4okW555DDvEFKXA+WpmQqSvFg+OJwWC+6Lhe0w2jc6F2ggchzSCmPcF2GakvIFPOW40OlH
E7e0IR1tmN0x+1ap0v3ztV3HlgfqHV+4q/CBk3+cfI7lRURkKzGFoMOYTwiicpLLp/Nnp81CNAqD
hXolV5nLYMOe6pymo5XEAdgCe40Fy59nwcwVhiobw1AqCoqjsrcIIDLU3Gxw5uG0xcelpnyVFWZb
ikPiYyIHTnPD/K/h17/DS7GaCS849MLSTQIu3eZmzjQetnO8iJZKbkBA0r5x+q+xXwmPmvfGDvUF
T8eWSNTdQe8W3jHYsRW6jbB7fn1A1Fw8cV4iQYDZOb0GGgIXhlWwtYQQME3NlUaSszK9j4P1eEj5
oOcyAC/F2/+o4DAVuNQTDTDlncnG2Dd0n84nnhzOvCmc3rai+phsey60qHKi5UD96Du3RNkp2/MT
6VJ4XT1M7uBekjxr4pC2u4Epwnxvl3o9owX43h5KWh1MhBV0ca+KNfsMOTpT8FMMO8FqFWTyi/F4
QFotzpjsw1hpN80MDpGo2g1wTxBpi+/S0mWZolnH3FUz9dzowwyqRviEMgWl+SlmV78xc589zYvx
3HCMo2SEYyXKyVyq+E0WbyXKUayAsO0Z7+2QYZiUYC0KwO7rAZA7AOJZlJsaCzhYEPZFX/BMz+VO
VsGPQARXLyWLJ6ewIOzu+0JXhYAcWTStOr2fQptqoJMHJRaT36Heu4Mfm1wK65/UmzEkgk2GcRxQ
e6TRsUjFpN0Yh8zkJ/F+NMUsgY85bmoEVGx5OCKv61de5P76wUVQrJMgkZC/8Pb+SIFSy64MC0jY
E7vC18SD3iULqUg+3IuEZ2ou8bign4Bjc7oAWOupnL0efE6vSDO74SMACn80/G0hP8GTfJhxsQo7
EJpL96jW0TDf8IN3WFA8DNdoEl/cifEpVlmBpi9fp7vZvOa4u/h5VqofcfosCo4FaI7uAYK+/6MY
O0M3nFMpMvuSA2ECZwWPSZBA67dvRHnkz2Y5TDir+K5cKgPGm1vSm320uFJ9QVHTJopmVNWyGTaQ
IS8jp13mM/XyFhf7rFGWZcO+Ew8U0azCn3yT0SGw/cEQEseYnPEqwut3TArQ2d7WZpLAOdr8Pvsl
HN5Jfw3n4iCXGt7EH0elrTZlFLtLcqz3bVxTrq2Dmnax1WfQQvGBhoGkwKSEz5himHI6P11gvoll
MqAjGryo9fni85hOdI/Lf1Y54Mob+3RLoorSCFjjQYOBzGW/nwlZe3n1+5LaOnsNwo9V2KoSBbnZ
XlUdK6mHS575Qxro/KTioDj+v7oXakT4wtSsxQISM7JjQ/QVc19TDnKVwDi/laihIqMC+OaHeDmm
sMpoGe5NDClJMwgglxtTZ+JjgDNM+eddz1OWPiGlwE3jGYI3PH7BcZ2a9kuEy6SCAvA2BS1quL4H
r8u7s/VhZf7/DuN2fcuZ4nfqOvBcRM0rV3gpOkP8DeH+bEP3AYII4IchS33w5nitxAg7GPcZ1ugf
fVZfed+xzrY7dCDo6OT3embE/suSQMpQkFg7FiMXjfkrgYjqsKK3jRuH8hRpWGaReiVEZ9/4hP/m
Moaujy4gfrdga+0clIba4Wr8tSK1Pc6+h/QRDKK2KL52ALTTkK+ITq1Xwi8cDIGp9i0bUNwiTB8n
eatywFsGyqPCJX3hSc3OA/lFkeJSD/RO/SPZ9Wv4/t2SA4zsLXQpWD+CyOSxa6Wqbj0jYyYI/8kZ
v1KkBrdcxyw1FfKntcsYci7VgYeh1YSou0u3HZME3AIU4pQ1t8cH/zhKPA09F2Mxtkz7G8FEf76Y
s6P5fWoDJq84PGLPkHqYpTnVWx1GjW2+m3f6A3KIooyELcLbdh+sZxtKKpE6y4cu7jwqEU9FuUnu
6COxY/3UDHczvNqMA+hId07al0EnpCLgjX8neAuw2fQiPe8x8bcd6F91zjctC8PnxMEfmGGuZc9T
T8OsBQq2SQqUUgH4q5lSx+0u/vErpHBUxD9WWpUWhrX3ATpv0KjmLCG1QrbGCweOIsxCoZdj9e2B
wROxjSf1obzygE0o7Rc/x1Sh7U5vv1JXcGx95qqpx1hOgnsNCEXbWCi0tk7kMiTB89ljORwQfRYx
ZxGfuuMSKr2KiX96WrRGI93u3qZQyjmYjwaACBoskjbvHetcSpny48jk4sORs8VId6yJGoo6B3QX
Hh+x3R0r8/iiIt6R3HDKnovNdAiCsXnBwBgwDDjfdDMNdnFqMcukeImMllT9kxMq8asFxDbWEgKO
wB2PvTWFrEgkt3GPp9MPLibKKaHtuJtM+R/X2OneoUR+IYT9xRT68Vd9vmGAV2MIxcccCb78ObeB
hYRde+Y+pcV2BOAOpvPMKVyDtohxA6wwmkU5RjhhUgEQ6Qe2fYCyCVpCiP2K03zuz/0x8lcfAvzm
dIh0OcaHO4e3kORXHi0fyUsV1yp4jtek7KV01T84AWCpA5Jp1P5dzhfl3HMAGEUdCHWmJW82gbl4
BI5Z/SxamFjjduuNfdfyksYsB1BK4y9gCkpGyZljTVbEMrvgka+MAkrRT8E/gjjGFm35w+r3kX0/
kx5Qh/FyBAVRwebib18FoBJA3DZMKSLnzBpLoffeIxALOTJEmp6vrFggvh86bH2RiMMBPVznKeoh
PiRMpskIcIgmOFcL89px18J4aSgpXieR2JbmHF63O81Kpa3stsBZJRQt+7ZvnQo9EjnYISRzORhQ
j1inKTPu9adyqoHJUOJHalK/sYf5i/9mIxpy3Yi20X1IjmqVsrQk37nTiVWhLLUJnR+TjhPyJbXz
jvl2Ee3BX/R18tFAwBzHxD18FBpUmSIv+lTKVH4OVsHPUEr0e4qK4paOHT7kuDxl+jml1s805Qqr
pE7dcn9c4Ur3e7dzMOnNaWeK8lbvYNrXvLpKUANqEo42aDQ03ccD0hMmOCJ7TB+Elm/pKNsdCvyB
IwOxZ96jrML4gFRyBTKbaulqyYcEcBmFoD8vUtUw1bnrYlSDMJOfsWV7zjZ7mSpY2gDJqIfqCayv
3al7j+aj97yWWa+yj2mS93QME13IOG2er7yRrMFgM2QqButnjnhzneHoL4IRd0l02yck/R7tvysH
G4NcB0wZtbskg9RKP+GGKh8mXNfEAbrZBydQNs6TWil5KZAeaK5t4Ylm+dROlizl7tK5TCPYt38W
qW1OD0HC5sLpw85PY6wh2nnIM06nFLZ9gUxwknTEsk2rgGRviMu6Qcn8gY1UyC/g+vdG0uZk31tm
M8lKu57zWOPSytDrsBMSgcH6Nde+kwXAz3AANOEEy2LYKdRqFUhD02cTUt+30r+xlFJE/Px3uWF+
vS2+1c+7VMCZ8NNeBxQckHQRCxz/9+tjBNOZKx8ZZnXI6h0v9pJxFhTTJGCEBHdDScG13JhSm/+L
sNnb3Aez0NS3EHWxxlkpg8mvW4dZj78rl+irEXulWTiLHZvMZrEUfN1YqtQF4ly6IbZ/6gdXcOTh
LFV0GWaaqPCj+rS1nFnw0PE61lzK+dWmZa1BgM93zeguV/qm0HuZxh7Z76lCLglToPLm7N1ing60
TymenQQaL+grjiIVTmoAa3P9a8SxnZkSLI3Cn0ryBOX02YrUbuzdvtMf36qjNs+RVnbLMhzzP9v6
+fk43GMLhZHKxlUbks6dIm4xPFKdSessnvNIseQqw1vdCeNSTiczDbm4otaDvo3oQVnEu5K5fuYb
E3YaZ2kvFkSE7PzUEjjhG4v6U/Jnovj5n5kkAIMVAiQ8LuHjXTQh/0VzsvNpvgyUWGtJYlczdbrp
XyevcZY7XADYF3du2r0n0C5FWRmyr5McjwuCbWEx30cHcIyrujKMslUTKFRW19zg5OH4ljwu/low
hyNiZGnfe/YZN0zZJfZX+w+jziBTqEOPi3Cu+rvhzBxAMiNFA6xM/dgvDplM6vaFhJ7smIRDrHxK
qTNmnJomPkwUKsBfqjJm9mcYLtFQYfycrShiXbJckqJLwx/ZGaPzL/tlGyhgmbA1qiZL2Ts9iGjv
Ueu+CMhE5o1HzZ38Qhe2NGRd4exbikl0sYVQny+Q0aojdu5WkFps8keEMAt4ZW+PFOG1G32LwsV8
WMGZF28rtUHQxGVoWWHtpD78yAojl/IHGkQyeyVBsbT6ZKEXCef5XQM/Xjre/mYvpfZMRdDpzYyH
sHTEE1SAvvNK4nNfz8wRA7Ztut6xvrpJ6dsNaTxKVHFbkv8tZjPi1VQpobu8WfXqlw3HnmIlTtr1
xcyeYy7zUPR7lnQxWUqoG5QS5GLwnJ0eu3eG9vyb11t/6VuLd+2S4E5I0MUTDx74LQlU9YdBCuzF
9moWIJsAD+8sOwUUkJcY6Zcp/DJrJm0rogkh9hc/jNTUEG0mZ4+PX+vjgeviUtq/38Su2saEUeBp
eCsCwE477OA2e5nQzt59SsKrM00HxK7qaBmgB4edsiSlnjyB9CMbiwJu93ZO/1H9YsJ//gODPp9u
Yv2WenKY9j3TERL56sur5yWilixyjU6kK2IGo4j93AtFAImcCzz/DZDpC8XVj3SKyprMnQo4nV+/
A+UPB5shsvIYt1e8DwB8ORdHkAT8kn1L9DY47H+t3OLIcYCCo7uTOjefdHtcnlcfO9+3sknXbTaH
mDi7ZT9+m5AnVnhna/MTS/aWu1Gp+73072r3L/5kmHKRMLsm+hvP6YcIpXMtJ/KsX7+CxjMxZF3A
h1Ap2Tdl+oNN7nzye+XKJBXPvh+pHn1wQ/WnvLP9ag4XZ+LaZbAeNeo8YbiV748J69tDTIqtB76H
4pYpRi/yIA4hW2PQCjs3FQYbY53s6xeODInkKiV5p3KEiJ3iGPcylPUW94ydzxJ4XUX7ROM0pgm0
n4Wo7xSVt6GVN0vW2QVVbPnSdrAbC/jx72Tw+NnXHSVve+LlfgaIS9/DDzaqCooIuRVLO9wZhsLm
GJcxRXNLcKfsVtYBfugURNxJRhmOcYyZzVg+EiXFNK1djK5NkLKTMH8Tt6PrTWBMVsnO7oFMYMo6
XjW6UxP0AktvZFKvyWHkefWYO0ZPW5j/ylKibj8yoGkcbHxuKASZpMa77wxIORMeP9J5agtqJFp2
YKSKnHD+ZyGynPeEcAwFLGKclrZiRuCm9RjCCIxTmn7Ejggvl6gd3RkQRJCSRUbqPxpelKkDha/1
ZclUf5kFNoEP74upPkFBWV5qnY5d2yryqhWqyN0h+AjbNSBG40PoLTNx50wmUQrVqFZufM65JIUZ
OEkYBMxJ8TWksxgHTfNXir7ws7MbNFrprrtNJWsQtTCiXVys3+F35FJxEjVgPlQAhifJgThcUaLQ
/fDOONeM3B3C97HR5iWNO8HW1+dKvCJMHHRUdZrtjCD1JFal6tCAIgpQbuize573CUFuwtRp5iHI
jsnaX8j8GQoHNrHZIaSRJwI0Z5m6F3ugC42rdPrL5gnSkTsdv+giNbDbDZwDc0OZX024zJyNcORv
9Dbk4dq6+DiiHn+NAQprnR12oe7lxdwDola2nZG8LlcxWwQJ2ccBp19VX8pDATrY+IOVmPi5x4eH
RHksJWckRbt8LKGVwmM36gsUxQVJ7b7YJNF2ONGIuHMYZ7caaidzeThqOFwjXOhD6hyfbozS+yxj
yVTDdLIUvitO/N69EDjxkvma4ewLvrPEoQgpw2jGReNvrd3tvXyCcFkaSBsxclmcYchWjXL7qiBN
2xhx4moJqzKbI01XMPdKHpQ5sEGojkQ65awZMjrEDHnN1Wr260uXw2UdcklHyQRjL/mHFZtXcdfj
6IDE0U7UfAF9svJsgOxYkUdNY7xg98FlJsD8DSc/1+rE61NU7suaniD9RbuYwpfbux/cS3lmPHy9
tHqWKMKqehXsfd5idJAgWnotTO9yR2Ocq6+w2Et2Sgc0/qsgtEKlm0ZrK5ZHFtdwUBIL5TB2IGcN
WXHhlCvPSw5Ack64xUeQYboqYJo9orCJ3ODuprl5l4kI1cXnOOaEdLzWYTR69Qi36e2mOgpX+0Qm
mUFuc4+L7XHDQQURah6iBBBGJ3mJ6ACMxisOO/PWZ4fvCttKnPliA14UR3MlJslGjZoDLnLQl3G1
VDFT3By465SHEtJDw52MWrgopjR8cCqimwBdp1S7sjxe4gka0/DQVU7QQ8NRzxW75BGxNmES/G6C
XFyu6tpzBhhl+RaOWyQXk/cQ7GhSXqPFouMEodkPfiXG0AARb2Z9y56etfIu3JAtLN20Kn4Np0PN
n7wXD1ErYQgHmQjg6jlV694nXT8paGBa33TKfEietfNB9djHniC8tlgJ6zYR5yNmpxQONv6QIaVi
1UQZcngI7mB/Ithx7D4FLfi6kAaR4ckYHWKscJ1s3BZqdZb1ls0NnfiNigairP6+358X09eYy4ti
30q60jwRPm8aLPf4kt1FMLOKkwOi0NL+CkK5MJ67CxPMa8ytq4sZELYspwRblBAlBwKbfslEpcJO
gLbPeUZTvG+SWTW2z1FKJsXedFdLBzI3Gvf25amu2YWciIJ0jqIvt7qBunYU0rZ278ZOESikeO1L
teOQ0QWJzvmC6mcNhTdo/1l41fCT/JerJZKt5D7VZCJkPeyBCkO72Ht7UOYnL63viUJdwvYzY4gi
/zKCf251fi5IQwJSBmEPrj+Pkq567LWmqSOtHQNrl0TrlsKU4W/zdgeahonEDTYg/stC+hJ6n8uq
NmXDNldVp9V7/zWzoY8InR69aCqBNqhp8N32WG5XsFkrgYAz5c36AHWTV758iXkHyLg6Y1Oqxp4A
Tjt6DxBWcv9DwB6LYWkOHHLnnj3QzMeRMwoPXcKjjq5oXqh89+Jzqs0v0guvMZn3k33vIq96ixFR
uaaatk/SnXu+/kREUH+a+0cHytpslmrgVM825I8C9uo8/c7uy34Hi+o9tP9m5zVGOw9r9w0WG3ZC
Wv7wUCex9RQQMcCR359TCGa5OH4Kn6amCUy2On62YYaJSMOF4eZieS8Atd4zsaeFUdKgdp13BocW
GI6keqFvcXri3L7hFi+ifp4pLs4lllrQbjfa+NFtOIScWUH7uNDtFbLTBH9hIKA/viZdlyQLaD3F
MrWGEkSxGTuqnzAuXOatT3iGf2JClHnbYPXZaaTsCwBtlAUoc9UDQejLTvdDVPuNe7skxy0JMyNr
L+aLV3+EcP63PH2l3LDZuePzLjQAVuOlxmZsryI7eWJmIQQIA83ewOuRuh93e6XXU55s/aWAcZbT
PKNA3vZWCi7TPE1ojX0VvKIhJKbb0zjW7csyVp3ujywAkggVhYE7v4y/SO4Nbh/Mr+XkyAWxn8LO
GSZun5/2b33+T72qgJou10l0lJP9KGzSsL8KzagTL775b+U8o0tPRlTAx6RCgQf6SkmCN+sU1qqh
FrQY6Y+YsddrwO4psMdCw+OpE3b5BRmGVXvz99xxWqVqRywP3Kluet4DppIm9wz/gFPBOF70lRyT
mfxBiiFEhemNqXOccV5Gg9dsjX192xPmzYIzNhPm9qo9fo4zJ4ufTrShx9F4pMgpvypHoMGu6m54
OjCei82z5cg9ipipRzxYKYZDDXJ1MP8DHGWxI1i6Sgli4j5wRGDhwllw3RFs+BFun9QuD6T9/8nF
u2d0Yga/xX4lNwAY6fETUB6tivsYrulM+0+LZnd5T+2+FFDCONAutTKEflperUn3fLKwn21joeM4
lhwizYQ/SIfBHQ/zk2w+w6RfbMiW+tcQk7Wt7JzX/rgTg8Ro+SZHekC7QkqgKpfYFVvbrRGODp2C
fBYHdxWYRihhMnfP3khfsmWUFwcuduLpdPPrxtucCrPuqYPnzcqw1Jp2Zxwj38Ieg9XXIh/RuAeI
vWcESJhEhjvQo3HedvFhjfd/cDBLnxAb5Dc/uy91oFaDs04Fas4LkI+QMv+jTsFL87b35F4syeiu
8xem5BtNmwVgwFlMaHQdwC8txtGUDHB3VEPzP05k2B5pVquSH/PfnxCaKtm7mzfiAHbI0mOcYxjD
lb+rEqoG9BE2S5PlQjrvVpO3BUtjRKSOeLB+L7RibNx2szIGa6q87BXUsm1x5ogxDCnGgEH0eFOr
2OTrLT4d2O4NdhrLDznxHCfUdSpbmZog9LJqKchzcpI6bWSqLaw8Po5kIC/lwk2TT5jXHrVrG/jw
bi7hvmHOlNhGBnuJvhdOOvox72Tba+tfpC0qPlgonodHcUmage/jb4wfH/aIzclb8jPjdeyrPqfy
ts5REXcNukYLpzWO80M6fQr5Y2KsP2zh7bTPmvSJVOCid2kDFQ76n2Vw1exWScgTCD0Y99Ejb3MG
47HLRwKQ/6h+c8ptqYKfkrPd+P6rDLhMqG1+GGxfoBSwCkb/eEVWCZVBWkbMAYjChGU3QpM3XGXt
WiyF0ZvyRN0tIcHuRt5HRbibdz8/DKTN3ACb1Incn4GkH8Rtn1cGu3ECfdM8NLsoTKTgGhD4pf+Y
2MyvzC0lFA4ltV9nBlg4Gep9OCkzDDCxFWtebv6J6RrnzNb0I26YNoHNGN/7ZRtFJzMpq3C8s0ET
j0PCapdCUYElDoVtBv1JLYHxsdBk7s91O/6FKsAA2GPZMvndj6IQEA3jgwrw//oeUGxWWuUSgGEM
+pVatKNf86dmBioxFpU39jGWTBgLo3PeOWuMFKQjvN/aXudwdCEW4Nf+OziwSb12tBVF7gXcsLN1
nmxGzm8BK3tb+SVOQp+8tcegor/qmUApjred5P7YylaXXeA1ELvP56Q5zdJ63jy0dhJ40FUddTEx
Bz/uB0Di/5/ADwgZ+4hvhuDpJWeZTJYP9w6rMuScZbw6CktXGhxOOy3BduKOW4Gts1Ljwev+1aEq
IokvCFJZR14B9Wa/L6DcnT4GEF7NGnKh+zZZH/VPWcnkOpdQ2p15k8AZDLoOE341J97r6BJqwMer
bclRuZZxHFH4XgFwvjMJG5fP6KGsrz/ivH5RQ6cJqt3M4AvGF10CfDim+zDcTv77Kh+nFw39kyQW
NWwJIYzlM8/B50F38wc3ZZWCMWw+pGnWhJrBuGUpij71kC/eNT9rZbos/8e8tlBpL9faSFfIXyEw
Q/HH+gvPqZvphI7h7+EJwlSFQl5bhYz86TJFxdIlHlolmPC75MJiiYGbvVW5IMtqsrkX+oIJkJWz
RfqLaXsLvL1j/4nH3Z70A5hcaEmkXrbU0NRSxDQjyRA50SAAKP7c11n3kZR28WbKWJ6oLgOnXOi6
lCETxcZgnpK3APJzSOJNAm5BWvpdxtBTBlhkyWv6VZ5j1cAOrRWOflO8DF9BfePA8zaVduGvoGXe
KPo9eXnvf6TVAifCc9/fIHDenW0V++bU/m223BQySLCodo0TqTbP6PovmdNtV5iO8e8U1/vE/WtQ
RXpc4T1xNsXyLsnTtVN8OoqxQqyuDlE14P90LlCPW6qERYH3UosMQe9hTc+Wt4YaEPKuvZUicNK9
GSuiXwiAWz3zfg7TJLSetwRJ1SWPnuQpYkpw60/nVP6rDy05z5rI2HY6FQyVQLVG9mZjuV69OeXT
UjRYfjqqgEjdbBl7Ndo1+o0oOcYLJR7wWB0LnSWuOHwomkptziZPijVD5M2aEpT9tqPEuB7vXWb0
7Oo6oSznihT8ar2Y/ehCtfw6unU2Dj6Imj5NLUg0wJ5oFM1kBhh2ca6grSJU1APF7nmPJX8A/62y
PROukmY2TSE7Ez3ewo7e9VZ96WO0VSMh+BeMtA7Gk9tRnXtr2XolUdESSSgRnCUI4n0ibAli6B+E
lHojx3Br4g9c+e3i/j8bp/BblgMRvdMIGmBvzqSlZmTwF0qUFKuzklE6tVWf4tIwwcutISlEg8Sn
BeJVkI5mPwXF8FAT5brbNf5Q4rV24U2iSeK4NlwfQTZczAN5zt0G23MkDpm4w6e52Z+kIwhrikqp
ar7NDJH5bHwE1MotqKn57yI3fTQhKgu0Tzv35kyP53kvtGdWXcuTlTtQBsRjkJ9x2jJrcMdMCk9/
HYTSAS601ow53cZfUPK5k7MuOMOZiG6763rxbgi0OkvzK//rneKETd5HTg2ucK79A711i/DJQj+m
RVv96KgtDFUylgzH4t0prxwSun7tKtxSl3N8Sw1Srkl8nkNp3/PAY02SbnIrok/ZBgEfx3taozx1
f1qqSSxrbHPtrFo0qrR1dgebrEGowYJQ+Yo8/O+pttfnBOFb3WSl6q69kEQ6/pvv75Z+RUhvxo8o
yYc2Cn1zK93oYJx1ID4gmIhOa2gY/BMZM1c64BW9qWGCUe56hOvo4STOGKfCjHw/AXFuNG1KGIR6
/k5GwkeKZVF7dW9kQDwWe0P+R+pB6UAggZDaxv8eoP5Me8Gf9lC1klKWr05psx1nfdrmaMUAE9u+
7i3gMc/wKOvcXTjYRTUOULb0m0tiM43GFWbEztHNan63yDJTr4Dv21aEq0S0xrTq9Vd5aN68Wwe4
Q0gbw3aZYrDt9g4gy1RtaUWh0HpvAjm9mYG5rcziXf8AqlRgWyyt30RQjK4o+M+5VFH3OccfuZcV
bWtpRX2Wk/yFqjj75SsUvyciTszyW7Ol6UpgXl3nPnVdxCjzb8k/MZC/i/cKd/ZUuk2sMFdpmfqP
zM28A6u9IDLdWe4RMaacL4nBdlQoQaLY5CJyVRspVxuYYVVWdSxPVpBx/vQwflslzFeBVk9zYjrA
qZsT6OS+2au/pM/1LeoMQyHLUXef3jrcpaKr87P2kfK/qzMDMl0X4NmF8u3hHBVHfk95wSxoICa6
tjdpMBd4r36mZaDynOwhrDeZSg0Z5WKJOC9KMdtPn36didRykphcktNM/ysKwQrOGOnU7J66nt/E
XH/iTEuUDDbiuHDj3BLnUWMrrC+7N4vUxO4iMolSrui76zgWYrLwzpy7xnzfv1mqxKdF2vFY6dCH
rSNx7lEYSoCUwC7nZwOps8uH4NNqeo3G/KZkBo0R+/Vd5BVDsD2O5qKr/dEf3OlIfOkYf9DxcsMJ
xDcoZ8QijpnxF9qUS60pxcl3jS8pLlKJ/g04b0Qic7ownyGXRKOLgJn7UDDejkMf6q37LlMIjYav
9EOGVUM39XdX79lM7yA/cePg8+swV9yD9An+WyQLxseiNFGe0JlaoaLK8S+ov5BIOcgwEXzHdP50
PZ540ecT1pmWnVoikw6b6C990L3creIjDMspzKkchkRZ29YmJSjW2k3IMJ7YeeZIvZms0OPgm6S0
/LYoCzHul1bCstMdi22ZEFOVpEf8jHEoImF6tG0iof19RkmBDtpQldfB5mo4LeklPJcUFBeVvscD
JVa8qw4dYtRcZdoKdQIZLD//sW8vCP7t2I4NXn+VBDStotRU4A7yHaDsP+PSaNnVJoitNRqDziHU
CZmyp4DChjLrlqCqqmMkX2N/hhNlynUNrxKa32+t6s0mI2xxIECHq0xOJzafGs1efEVDg98zE/CV
eUDERioxeqa+vfvOWFOS8gYhAsjLAc4k7pVO94u9ODmqSLifgc2nIzxxyt3TzggHM2E7LhZ7jJ9i
RY212ev2Ui8eL+7vDKWifuoCmKaFDJAESRj87Rof6wzdn9id4aw2K2dXZpecw36b1mwKleCdT9Zj
5+jnbcE5Lm7YNqjMV3Ox0I5a4Kw9Zah98BHhfluhmZBKP60OfyzUr/BZh3m/QXsY4fO9Zvi+snoL
k1lLu7GVvQA14bzd69Wdvp8zkeMvzWpv3IowyUp371bViB0NxtwDHRbA8NbwwCa6mJkXsbf2PEA/
Hr0WwD/k1a/522KLu0dGecO/o3CLC6bgz3mmRQ47uQHJvJv8j/V6DJ4nVmNnzZYDWDoitNnRdxbW
EboQJAtdGhxCr3m6yUcvLVKQMtEUaexU8uZqgRcfaDQ+xzF7BsLyX+ZVhrIq5j8kJbqdcIx/YBEI
du9YSxzriQ5tjKqN9ehleqYHvjCtXMpCoUvp/ZfA3EK1s98c5QkwuMwl0CHEIVL2JpjXfvLCfKcm
1vXlW0rB3vmLkPuoMO0AB0fMAlGi33LzBwYKyaCdXzJivM2DMEW1Lofav+HR62khR+RZIdLk+mgM
m5KDHezoneJrFPX2QyPO0T6oEjS0Tqf9ONW8sRSG3UUCUbPKff+T6Fig8+vHrjPU006whBVchpWh
WoOGVpJAgypVB4BH9oK3uz9aiFKYvDrbgzJkshEFmoorDINnqSXiretnmenvNudmDD5vGlZuFJBD
qBr9OeUmd82jjNiCDmXx58cLRYjsmHHXDNy5WVknQ8ikcPg262+qvwRxNAmLYDTDsro9/tWKW8Xc
kSxnY6RP2oRLtQ1P1NXx5XZ8W+Z03CTvjtw6O0CjMn5GeJm/qG72emkK2knHUb+W9yMxWwgg6gRy
OFsxu1r1IazNdplPxNPNN63GEeKlcK9y2C2XoNdm5ORCwMePAvFjw1VLG1kwgfGH3AecPyOYlp9u
rLvWztpkt4a+a/6tKkskeIImvqEfX9QrmodY2kVGubPbIgFIqJa8aW7G9c0DRNy+j8KlIYMcpcRA
m15Eyin8ALUYstroK/h+eKkn3J3KUm7tkkdKDiNVInQ4wMj1iZUJQAx0i8xliQVAV3F0KewuwIrW
0uJNtZeJ8P/dw5s1hN5OsGwXMJz+avwfVC43eVNuT1LRmFNfrIkV22rk1K1Q5FN37xqL3lUz19yr
xCCHivEw4CANhgcHjz/w3Ra5upgYtfOnAhuXAOQ4dR2fxYcKv9orPkBr6FkctTD7SwgoJuDCHTZm
FcA2iesJHy8x5gVx3tKvBehA9xW9ZelORmtS/U38pnOW7Ax0DJTwGy5fO6NcUdrCbOLga2a3PxSc
PYo+c/JQtLaNj7WU+6floBPib7CdOtHiVvVYkzvlT9QEWXbGJco1jY239Fj6zNczP3BohasICT9+
n+HrrsxExa9Hzj0EkeA+Z8qal10PJ6zrUyYbGTIUvRmrQwHo+CvYxKiDsT4BUC8WYtcHho3M+8HE
M+D2dcIRyOZhOvN/EOGemOFpc+77S9GBITW3WBcEKSVUy/HQ0dY01bnWcqW6Cqe4Ih+o1NagnkmH
2mB7iplYxfL9oQ/X8lyHCdyA1GUDCvo3408Dk6QT0Hg6XkVOlt6aY0QFtbmM0imL/gDLXjDMS6ZW
BFVEweyWk21KF28E4qMn9enVPHqXsaZ58BJcY7W4Q51Jd6oIj2YFnZDEpKAGTkxLo/jMUMEfrlgf
cZt+2+68FVA+d5WLP1mDJw8SNDNmWW8qubGky3rmfj+7pSB6ub4jStGu8lmfbQ3ga0jnxaqUgJ3m
8LlOwpL+n6xROKcK0V6D4Bdncy2mnMMqZbtjnVm4hJiWw+phF56BzQFk+XmybhJaNn0QJ4GTcJih
79sqBcj11+8EsBWwKQkadef+rZDdyCNbcehah57IHJtjabYBcWJGJCWjm8mG19y0ceFKf7O7XAJG
rRYhOwbKtxV6ET/LxDyLyb/81s98rshJCqX+WCDM2i+YKyAMYnm1mlqE/flDdcOIMIgxVOrCuJku
3oLiyL79vdBiMoUVTZc23Svg64qqGlhg0R2zpu3tIfTZtBUAG8X/ztnHOcbERSwS2+mYxDsqabQD
9RNrT3/CxKRi4uJUWSF608Tiw75cbBFZwMACg3Z5t4r+0oQrsSAnoaC2EjJtr55juTmFojGgfJPG
0WaMAnQ4zA5sRp+DJD17kFHb6uZVesE9QsSPVanXDRi/E0HuIFvmbaT3jXpoXdEJ5ZuJ54VoSy+c
3lFcP0aRNaAWhI8ThknWZS4k7caBSJ+HUbqBfi4XZjInyFtb3VbxFMjo2r4B1Y4UU33g3iv1xnDP
Qbt45W4iOyzbXcQfktucm+kW624WzfNOpnGDbqj9IUckG+gtc7IV7CmcMZhGzL53KjnD3E7Nhdby
G2LbMJuRTItYQuZD4JfpwcBvbsT45XiNo4v6wOz1mWB8QEwN+ABRbyLtKMnW9bQrhapaKStAyss4
TeV6bFKCykx1Cgf+SV7UkIhAsd3wOZjcr/Pkt5fNsyVEbFy/r18yD+kImWS3nbttaeudt8chrB8Z
UFxu7zDCLc/cmqAin7pxNKBPUO0hrOUuk1Xq4sAL9UOjWoNZk4ICxMRX2kxNk0qa6P21JNMdxjll
QJkwoc0sboWk3j+OgZ3Z84ugmfJZ55Ux/dhMsxVkfDTBAZPEloulf1r4RG6HA4xo9pTUw7ygeE13
MaD0iQY/iqwGQTRj4GjOXtftDt6ANYEzfHvX1bWnR+lQ/jUh8hP+MTOrHgowiYvbxltVH1EhYIQi
mTe7u0Z8qBR2GYzza0gOm0dWoSDzLcLG3NxrWGpdNqtSnYpnNQJHg7CZHRUarUDn81ON+9ku/67e
OpBs+ZOjX3c5mbHvVgz1v8AzvUru6lvvG4yI42mdl48kEjz5AK5VfLLwOb3M79smm0sth8847GvW
XmdRjnOjM7WkzLfOhbI9oBsjgcjHyzoOoEmZANDmRGdal4BlJWnsaZL7F6JNnNvTM3lKENO+fBrJ
7FRiOjhfDGs1W0KmArVU6Z2ji1FT+L8Y7yv1kAxTgRNTZpud0WGSrZvwmpyeXAPCWCryaQ1qvvq+
z3T8GGvNiLh2ZDJwdEEvqWy+5pICeVIgm/34lErkQsNYuw/dGcPFOuQZ4Y7DQ8H5GSvLF1rbjfew
/HIUYJT4JObl4jGU4rehwENhSRb0wYG0TIctMF4W49eOQACDVWi7R3JfxxsTqbGYdwxk8+Qm5MNm
RpCgURtjOGP9DMlLiBiLfAA3DG3fBt4W2KNhcpFPmwzaK/58nZOW9Jb1rmGUJ7jJ3wdr3P2Ss4VO
Bge5YbL6CLQlzLhe7yR/qBPgF5uwW5ReSBcybx0wnOOGNzpWD1/1CJbW0Pf/gSVQHv3Ejl1nCqJD
j7DAdIi9FXPLBU5vLxL7m/lOnVGjbupHa2YTIEmQ+5BQcRJqxeKJ+TUNAwQyhJvaKSA937BzgPwL
fHA/8TngvG6tbF9Kf8iuP6zLGw11uuzScn9BBf+Q2bGLNxqIrt6nIElD5SA8c4THsWqSkCV9QdBt
yUoeMAM1CkA55AAAMt7it3htLc8zcN7d5fG9Ctu/D+myR6Hf2RNIl3jM+FYmUIb5dGvs0Cj7+cht
ten1aKyABv4jr3V2M7r/n0zqjmz/6So53HSLkQRS6crncguZRTfUjbMwleiqoQMFqHogVxuaw2na
H4N1+vH02V6/hudFNQ2UK181/mC9tqzgjvlGEQz7cZXebYsMXiRBiAjCGAssuAWr8uviC+D+yjKo
TTVGkmDTmm0gbVdCAoWkQ63nYaf5EY6BjrMzE118j6+C4yMybMMwXCqsjVja6BJbAtSoXfofL8tI
FNZXtqpNhkc8W20ZkfaefxlR+f/+QItPz0JuqT+9m3lq0sWWfMKQDQyBDNkAGcHBp7P/a6qYk/dR
1csFU/LAMaxpxeDjDlDVruM+T+5UcmdsElkw2zeWPsgRivqSEo+U7A2+CQIXHDvldcioApsP5RrF
EamD8lRWO0PHeWF3mcv8Er0tQ/ScD9j6AL6ElU9/afpQJGLfnHfNjT0wpowWd6730HKC6U7IMlLc
QPdpAf28v1cGDhlexOxo87745ymoso1hxmm2A/W0l5tomMvYRoD0CzPp2Z0IXE8D8I+t/RvAVBLt
+yIvlowxQh8HWQ4dp/lD89deltqeuCq63RGZmC83LBJW1XqOXyhcn2K//xA2MKhxP0VeMfLk+Mwv
wgMWPtzK4P6hi9sbO8TtoNywlZLHdcmt7kBetShxNZVuwJWKkgPlm+IjYrZDZs95QEe0qVClHSkq
+7bXvQ0ZlOFeO5q9KXZgLi55bD2FxxP+gfyQAmel/O3zcww9E73tF7BOhYqy1qa82G2PiDlof332
jRF/6Lq+/9M5T9VSvsacR3ezddb9f7xWyy8vH4jDsFgqCxnAMJrPGq/CbvG9KWZX+Ltk3pw7nF1p
7iMKwI04nfzeCz35wulkhMMFJP0tg+GZ/Sbzjt2Do2A+nM5zcgw5WUPgplsjAOoaQfoo4XBnVzkI
puIs0WXOCQ1Nd/5UE2zjFMAUsv1dtzDqSKBOv6oIboNuwod4B/1hjDItB4P6eW938C363gOTyLyc
cTQRVFLguq/+K+/dYvcEZEDxK1YRuBDHYZmdKR2LjnGwO4xRsA0VT3ADa/uOVYMi90I/ohD71sre
weHp9PcXFvWlTjAYKIAzQ0ImjrH5aQSAIAj/roLFb06dY3/GdcsW5L8FKy9M3k+RmdepZFyHSL0Y
Qos6/UgRsS73zPDG3H8aZ//gO29ixiQlXdtJfVPN/s33Q0hvntzyoghJOPNQ3QcOiX1cfHE4oKYM
ql4V+ig25C/16Ox4D0mYM3Qz8sRZu1wyuizYRlAmuhFJ/5str7FkPCKgMZaOA0qqMtwXY5zJdRdu
sxzT1/dlo+2fHR9nvGDGuLe0Z+wRQLIdCh8eBTamsINWefrcTr7Jf6Bs912qA7PBZHhZ/8im77oG
H2/NZWPIJKDgFKeWX9ZgCTK0L3BTML/3L0y3GCXlciFYJbVFmTewYRL7ky9q9VyAzXP0SAEBAnKC
0lG5LnzqH7KpsOmTvdqd7dHFDsUiGFRf42kmnI6bdWiWBvrjJiLHn62YIATxBPdfXL3z/KLpemAa
Az4n0r76jQO0WM9s/jjPOGFTGyy/ntecHCCW4Fdgh4yc8C34gUs10d62biKP3anFSv5nguaKNyHp
ZVSHxbesBFmXcy88ZXg1iU250oeoz3ZGNebFWKlA3s/J4fMrm1m/IgKk/SYJYxm9FDGxNVr6+L9M
nmh9ygqTPIo4z5hWHvUSnr4j0DJ/+RqzdaPxzHcwFwEwXMAl+5OyCW7IB52f8L/9i1NsGWP8nIlJ
vbk2AqAcSjkh7hilP+Ti0qLBfbGYzSCJtKx9VrtYhriRdJDeZLNNQBwF/hzjfr2EuhtD9sdhJvxP
9y15rZKkHFzgkVVLd3uxrYeOJrQ+eEOxHSpjxeCXGCUcUjgrk0QO3B8PWq5hBx/i84dTWjD2M8sP
6TFI1c2jRrHbOZp1dghvAwwwTIuCg8rNgDLNlV0qNMnZIVUbNgbSrSVlJhnr5BhZ82PQwhNuz3QG
gqzEGP8KYZ35JW6z8YQS1noU/2mD6PBexSKSqn8dN995cwqblVqX1JDHZuQW6ZTOyul30Og/VsIH
tTJshPLAHzofYj76iy8ADp/l+1TGBAE+QhMgXJU6Dgicz/3TWkJ1fOCEV6HeaIbguoUrQnWwBGlc
FH5GUhTG7CnOqXq7NkN9LnmqJBNYR9kobA3OECPMhCgMyQN+rmyku1x2OHXa7YDPfsaC1puK01DE
wS7Ap2cwrBoRebiRxtd//5z4zJWU9fAYkiY00AD/5GyLu0y/2fL8/8hekTGndRmRyMfW40GgwDII
kOmp9/nepsTuQRPDCXCPNxfd3BkR2cMZOLH/ZH4t6Lltcj4SJMAmgl3r35YMjZvFSx9VXzBlnjQo
mKEIubO9GV45kNfd/LFqkFjzRa8xFD7iIjPVs00K4GHFOXOCgMk7Lme7WTT8oNx23kcB0mG++Nxd
8blhCW1g9q+z8cRbm6qk/IoVGRIzWg4lWf2tZhTwgDls0SWhxa7XPodtqS8TCxeUYAw4BQbWkm4x
lRbLXdaZZxYBLFJ5hj/Q1AhuF1GlbZ84ut2EgKcZrKOjINVHy0/FgZDY750ANN+r4bP6dv+r0DVD
a9Zj6GVtJSOUo9FOtZspZEwPlYGKk1QnnN9uLRjhnmaWeD9Ed9foQbv7Dou9Ll6awutndqgofPvX
4OAOn+dJ62y0l62C+Snt5SEIoCTXmN6qtOffwm39BTKnn4AzAOEh5c59xQvJP0vlTf8tz6p57IfC
UfjOGQte21N7onTi0hcqXmTw75dePbFNCHkMW0MhJ/7zJewVZT7VCt3xIYyytnZbOaOuADmb28i6
Toc6S5n9dDq5nekCy3I3Lbcmg9iJGF1Tp+1LXw056O2AfwNWTisVQ8WfE5fnOM66qBFIM/H7P64x
3iuFQyxrJH+j0cSW02ccz5IX9ZJMegFYsB6nHry+t8YgfcfeWO1LWIKIDsg4FHP/hrfOKl+JTf5o
nc+/C1eLmzOMbm3RBoDNr+UmQGIQ3w/IEUrSqDImGvFnE+LP2kTMESjxR2omE0u8iDbkJsGEuikk
hNPPTERjGTACRXM3+5+1MVjKGlENGGkN5bfP0k0FpywJujXuAxE58YYXf4m3+T9kg6zVVsvMstJh
kyptrplhJaDPu/48sQGKfeQBPR/Z5scU2j7/HtAO9vdY5gsvpO9kwRPl4K7PL3tMOedLm9XM7xH8
4yJzbds8pW61N17zZa1U/MmvL8GGyRNQr7mgY9H1TCQIcy0wXA75e2yO+PH651r8r3vfUNYHPyox
uDvxrkUxrW8Pb5D06E46BWIUd0rEe1EdOPaE5Je6drlswSSNhh3Qt+E78dEVIQh9wjZ/Q1G/nCrs
fW+pmbf1Wh6IuUp8ChnnBQTPPiB4otJkJLR/rIqrLbbgBIVe+W1MGSqp1Ib6sbVZHWJXV4+685r5
9S/Nu6Z0dzP9FhhJm2PTTs2aJ94fKhbatNfde22UHsM4wsYmPFE5Y35tmwvP5qssc38VaTzxi2cp
MfLwxO43YQv9lVd+j3Qrw4/OBZ0Gn7u+W2Wl0a7ju3e+uv98oWzg1VOZWajXrUxfix9suxFIlnZ5
rsLsMxrxJCZR8/9R4s6Qt+DkuvPtQ45aVCwoY1NEQcKnEd5vQllwlcPaI8tAoChChQY6lKEdwCer
Ew4XlQNZ+nXewdNC3vvWRk2JN4dCkQTJSTqA6U69CteWfbtF4/mq7KKGkccqthyJpII9kg3nAsSS
eItrk87qTslRWFRgL6qNYvM/JEt+jwY0s0NbfjHJY/MkD83h/cc1bRHROeL18UvMFkUQBl00bOo5
sJBXh1Ke6foPIiSCH3KTZ0gmrtjlABn2Grm4kC1bI/dX7GK1jnhwgR7bPQDUXgVC0sL3rza1E1CR
d0wrqwxQoVPxzplJN55aXZ4pc3cTUwDr0SnoDOdJWvxPJeU25+/df5sGuUXOZ0Va2qi0ZcHNoyOk
5n0EUizzhuNQUg0HjIH0tBgIJ4s3Dx9zbZS9Wofkglbijlu9uXdsKZqC3C8jfQavfhE8GTLXpC2U
9XQFAtHYC5mOczGZjRmmIcolc7bW4KFQKP1J8oGuxd03rhzbxhEOV3mwVsVQA31gxi9elg3VA+a/
AuxKQvk+7sInlq4LsfDWAE6iVOKcayB9wrWcaZv6CECrnOncop3BmtU2Qg9nmT+V8e8dlwTiRxUd
hAZK1D30o+gGqdvFC3ItEq0oCWd/DKNH1pARGT3bHMSxHLiKwlWH5BjBuYgaYD2T9s4vb4UVd4XG
nR+UMVeQ5xiR3RPtSy+3C+DOHE+O1YZVDIe8aBfF6ssJCQS2ROZh8sJkRX404JlnJdYZD33hzohQ
kNvXUz6ORdTvBZdokoaHifndeA5IgTUb1FU8EfO20ugnxLcS+CO4/VlelNnNRa9D86XKBtG8DNVj
2IuoYnXycpCRqF8x/sVVHMduXDDlKHTTLb027f0SIBupxS0ypAyYG6anuWeLjvlsQROgEBPZUl4g
XRrLmzMnDJSRDFgNR95wpc+OUqIKwW8kFy4ebTByFfqY5w9/LesXpzAwQwBSKK3JZ1BYNfI/OfQu
uMKN7KJMsdE43S9uo4npDhcCoKjOVU4QU7A6IpkpJs51atNe21swj0e7XbiJqORhKpHR1ShNN0+8
rURL5HERN40F3JCHg0gun74f/ZyRa86kfqmWnpLYkQT/4XNnTPoFWECfxe/KeRZ6SQK67kwWkdwF
NYRNdwkInQUjKTLirRs4+ZK5svkV3fB1fa00Y7hAGR1f4AoBtpISGglirKwF2V2aETcz3OWqCLx5
HZc1d5T0tzE1k+Bi+RHYYBEAJy3/ZFRa76QS9jF35KlOzH/BD93+Z1R0Y6uUrkrD2hGdJvzLg/sE
/Mb8/BhneHCJ1qTRfCXobsF9stAf/VmK+yGmXFGC3ZDG2HhnK1+j9avvYOKuarMZWp8SzTjxzqxR
GAjoIJBUqz7mrCRokyQ/X0iK8XXeMhYUnypxrLwFsg0HPEZPNj5iHHzuIWWRO5gGvnA44iI8vJIF
yg/o3OeGCLiyiAqyJ4+wh1GYvzZw+S+64ku6g47zyPZZtM6BW9Fd4IelFiIifHI8QvBzApGg4tKo
LEmTAvcUVgDwgyUTr6lGMkR8HGD3oR/54f9EgAP+L7NurJ3GhqWAIgEMSwU586ABbJ3U4sQY05d/
tbTYhyeMcZHmeITWzMetNL4Ns/QdxZsGRgzViGICpJpjc7DQIbTY22zpzrUHORjXvCWLSEkRVGtN
sRHgNEyhznvt44y8DTBmqUjNww7lgG0bFoHk3RMl+cfKg+HMwXQ3VsVBr5hZMRwD6kCeE3rQasCF
pWVAB3A+FAjj4bSD0r/Z23tkLJh8d8avOFJCHhqTj0otcsdhj4wWg2sfrsn6ICm+vYGaGZxKEwB3
bJ29s6fwYUh3ZA4r8YkmZuJS6TFB3kI6ze4zSMNlOX63ZAAtY8rj1P1xZGy01lR02mqGteeqN9os
oGplN7mK7DLx8O95ge57XEkJkDIZQmrZGONni12JRBsspRf6Flw8Zs5+CDtyZLrqm/K+sDJvOWT8
QElWfyNfxBpAejsPwt4hSneETjRfxUUH6iVhsZ/4/Nuhgjbw/PIgWMRufOe3lBvWYvTpntsLW8VH
4EUvaO3+UqnBalXew8NOXPseqAZHVx4q+nTrl96o5kapFxCb5NrOQkeZ4vilab315Ez0Jzgf/SUj
N/fNPXKbCM6so/lKcvU1nbut5liBG/bb2sFGZT4pMikr6zsC0NaSDaMhjRdYV4SAfgSOOLtJIiit
ExYjqYAL5d7EcJsVJAyIKuP7KHDie+eEvIaoU5BlC9yjF/VQ83V0MN306VrvEw5i1SM6YZPk+JAA
xPEviZ3P90zQFDbm4g7LOJhTNEmA9Xa28dR/4+v9FBzDt43ZNluZ0oLz4KYGH7q7ehwxIzVkqJYa
QrL6dnV5nZhI8QIxTudgzF13b5SZFmQHseZMpQuK1WUlibeIbe8NWC0v7ZFi0+pLY8geWnnT3mNO
4sIMCL3HNuhb3icxgMiysMupLVh28ou7N/7TVHPaTrpEckV7wk5Dm/yvdSX55wl6k20s64bw+PyE
JHaMqiBYdByVjIoDi+bbHCPXkekScje4sgrXKe+iWZEShT05h1E3PMcGkaxTP++4MFsbbeV1sDYw
NW18m9eK7r5gYBVJ+qJb5NFvNQZeqRrssOOWpa956WLheEt+VoP2blEeKpzYSxGuXmkBXXqFw4gB
ggYxapHdgve5GSellToZ5mEZxhZ1WfPyN/2odHBRyz7u7KYN5JrXR8qgSz5Hl/kI1UgA62vwsJPD
kPEJz6zlKQcNhREs6i0hB4s6072+Uavha2DuAMTkzTFamZa7l6Q6gT0olPGRo1p7HEMNkZrAXqdl
5pG4TJcLuNj5OhynnMrxgS9URL1fAQweOX2eVjXy/lTxBPViSg22h3ulHROXNrEg8eplY2AncCcI
N+t4evaDWOgi9fRZfu0SAZss2y8YO2YqkDG0c1RyuiZxM6bKiH3hTnPs7JvR7y5DLHZEl78gq6n+
MP/Bxq2Q6PM2lNBCVOq/sW942JtxkfJgafot3aAIQvOJET4cFbhvXL69FGJQR7Yp7BZdeFGI+xe7
ygWIttcMp+sGjzEIyZbK9glvlQ0u7vV+YP6aKndAeHQoeIFeO+k0puQyLFn32iF7i06XH5vWxvyC
ZWH6zJhdvenjXBchEGNymF+dko18u/BysaHI97fGfg/w+4FUZipEZOAjnHCWwvwoe8m3jyvdJbnq
NcOky074fOm6myiaRL/l6cTkNIRNxayxjrRaDbgFo5YibPC3JgiXRxJcJY4XanT2wVqf9u5iRTeF
gZJJZN3HwTEaug+MJo5A42DDBvBL+pcMnbDkWrCtZHybpXTq1lCtB3xPpeqvOIu+ES1A8kDXF/n9
93kPFEWs35+jhXadGlWUWbunDto421YDpCLze0m7Z3c/BbC4s5scurbDjgJ88XZZwnErNsdiynQ/
dG6vDVyXWBsGssuM419xxjnlaz+DfqsyBZtGbdB3jy37I0YpeyAqxqz/R05lh3Ewizfr5o+ow+Rh
Uq3jhxaDapxkwSBcGhNYS2wn6NHPVsWHOJkT9js3lys68gJQs6CJBG/aTeB7dH7Kws92qXKxu/IB
SY5R+kHKssxKDnXRz4gC6Wt5BpUADwAaclR4I8Q66O2+B+J2CJupgJXjUN0Rqu1pwtvev2V0mwHH
a5VIK6GeDAHD61dB5BzX+6VKGZxNc3xQOD1nrUT0mOtqzl8nVt6pQJI2U/QTSdrUHtE1lKTpgT7c
tddERnRTceSEL+4w2y6mkEsHTHn0V+tjiW6rshxIPq6J2qbx2Ie2TyJpV63/LXvf6y5IvNpqz249
1CftKPQcPVg7J/GRsTjn19iPW8kDK7yWfjhyYHFlJ84FEmIwImAh6Ney0GKVNxRFkrKkfh5uGpQ1
+YffsFXl/3HgVjJTVUyy5OyY0W4o2tYX0RcVMiBk5V9fosWdwCnqx24UfPmBT9IWUpcjYbl08Fh0
pzClmdG+LjOuHpZd0dqBre5l8HNyyaRz/JpxpXVzAh6PUPfMQmEW3+gGggqLpVpbsSa7WVE6rGYy
RvluY+bbc+iy0toJOx0Hph/31RXJfxJZztsj9z760GvndONfKy5bziXBNRQL0gOAGaV9fBrukN1e
vJeQWuLvbVmynvwvggfU7IWQT8whKysvvyoELgM7Q8E76SroimNteJUpWgKw6huAC8vPEHgL2wpQ
z8+yoENr7XnqIJJuvg0soBPXDKcB7X5rw9AQavpytXAXgRC93rH1/rbJr5iarC4fgFHJdYcncox9
XZzn6KhwdsSWIXiZcricGzUe7oOW80+3Hp+F/AQq0lNKDE2ofHGMLsYohAoon+PTIYN3na+SVqFb
cTYYBxSkjFHYvkZsALBMDibapRQQNIU/UpH3ub9crF+KIZ6MitQGapu8iC9vlhPZsys5WH0XcK9g
8zIjfb5fbBea7Q6ZlDMtaf9p4cOxfIjDBPu4hGX+ObY+5XNal4H4GhE0dL2rc72qUVRTXCAL5AD3
ix3q5cGDrz8sa965TbjpVYNyV733BJquSW6/r1rtNTQl0CjasPNRrv+UQ1iZ8nqQgnwGAbmd7DJC
qepe2w/wx8BmSYmLs1/olsJnprxESto3RQYAvTfJdh3QPodXbiLjc1mSIXPhfyTq4pSs4Jb1JWe8
GoYe7WLGWDSY37xVqUkxTTvfoxF9zCNCr79Uo4/S1lE7mqDLHtUPPKjCrtYFNZRSTLxCG1i2gRtS
tXFPgpAzmZfZzvYJJW0o2WKhHWWeoi2NG4NbNe8sO1frgHPnxQKwSlKsp+uEW3jYHPTm8p96AnZ2
7c0zXCwsn8N9x9JlCNLf5ynPP2ToUE18FPr38goh5I8c9+1yVhQdNbEakzXLYoZKtGJQyAxy3V8l
dSRLeTPNj6Zc+mMA2dx95uM47IyK2L9CEJloUYF/kbpni/kyi/oJJSN3fxLHhq6c7IYXJflC09+B
ZPpGLrr69WadsnpNLGBw7zePzntenPYwes4YW6rA1ImLwspOGJOBk6okbcaXgR/1LhUcgvvheTSV
Lr37flj88U4VDKgXxcc4SrccCpEY77DUhWQ8bhZRJpuE7TRCrHcZ96Wsl9CbubNadg3ZNf5NVlhU
flWu4iQq5+XlpjmBZzpADbBsA/M8an/ByRQIYpmxhR7KOJ4jY81/bpScJxQnloGoqpk6NrZidvf6
1ezKFQbUVooD12UKshsvGfEh9i1fvNskMu+/QSNhsa1cqUyPD1Vija8GdmK5QlUCun5EFfg3L6d+
720j2ozg0LcAdKwwM5xQP9G7axot6/HROnr1kLkDAk/sak+q6cvqv9ncT4Z/2Sys69cOqZYQv1K0
tCVdLQXa0QyD+tkerOCWWPgXoqlUvfwAWXZHcTifvoA73z9c8CDU93QFwVFi3lcyodlB3pMHMykX
Yz9iz8womv0eFg03UjIZaMtXH0ISqJPEjGLIrigugBqxO6ayKff/DUqKrkJdy62Md5vIRv8bZ3ym
9e4fvtxXPWLqw0ERSoShoyD3WR4Klm+kmxTE0fujgerS+Ox3hfZ0yUZqAtw8bR3sEUq0HDKt5OzN
YVmud5Di4qDWsVoUeZje5P5RqfAhNsLLPwZK2Ck9Q8dC2v1OCRE+Zy+Xes4d/UH4Sf8o+mZq8an9
FNd9Q7vy3ry+LETwgEgxh3Q6QWDIbwVLUldNLdPL8aCUt/pXYp591x77rfSeF5s2z3XXpeznJ2qa
hKfalABgeQ3bv/idzjmQMVnZDhWDC8tE9o96xvUnVSwjhQdbio8YTHpplj4pZp7M2+vHg5M8oKn0
i96wstWhDeC62pBp4ojS6M22Akr8Oj6x3adL1cx13IyhImkeZ1sxhGV1tWNSPB81lyWA4q7Gsf/Q
DVYctqql4dmYcDKJkLGJx34EAifufU9ndxqsjfa14T4gnrgw8M60Xhk3keglKtNs/vWbMu2LD2kZ
CN2kkxjUCKMwbLmiKE83HA9GxiLdRroismWYuDANoCHm4CquSvFlsoLmk496xNHSVn+3w7Oq+Sy6
hxTe0zEY28wwY5U0ZFeSNJjoybhUpK7qiEn9RFvQUgq2Mz4jZaAMQHqEOtZVb3c8sk8vxkLp1W90
G6/NhoxEqY+GZhFTwUN2Za5JE11w0Yf1WfjSNRvqnREQDNn5wI2n/+AVJaI/gCmGADBp9MBFKAlV
evF5kKpanXoQwTn01oWW6DOR3ofAAFeZDhaw1DyGVQDCJfN0fbAdmmQ7/oDFp4lvEktyNB2N9kRc
VafLQwz0CcGSp8DNBQFBpwQZoVBZYcjXiYCWSB3B7aHZtghEhCKVhPn4lnNyfyCxufTBlp87G4WB
NXGKSrP7kOtQe2oU3TYNd76FPQRN0zhiUFHYspjLbQ6W6AfYURMBt6k0s1ejq1x51BEKxpwOeSWf
KG5+6VF+o5Af4otFfWWolOY19G0X2BlcRAcXl2m51L+bLhEQc+hdc42E0S7fVkMvTfvNPjHQvUr7
0M+D2CxlzdQ6e2k2RGw7aB0sft8/3eDud+K0mwzcUC9ejwklZmQXas+v+/q8P4xwBW/FjsPjX6vt
8Gwn7iaP83WlkILpWVFWWzGKdvsJKrgLFYHfNWTs9dO+AbXBkguiA53Xu1cpEbF4VVENkp9Tij+Q
VMrEei5u4a1K5T3yeLDKe9wze76S+jY08wzdM2ACaI7pP+RHx8ZH4+pa356YE9fVlQloHy80xOWq
BFFT64MklCHAG+7ibOLJ3RLnN8WAKHgDbAL5EJ9uUYiaH+JOfoV98eWpUZ4gNpLjZtmwHUbfCWUH
a1pwpdNkRkeAcfNxGdcxsf6xtSfBDROkhOvv5i0o3xj45XgOfPB61+2lyOH2877Smn2GdSzZkxCU
1ZLcx6op2AcEJbTLlQSyLEw0Gf/DMeDHAO9B/R294a1M4aR77lmW2lSVboANV1B5jPDkbVldckCF
bmr/C3ifL2Z18WNiE57eiWofeecJBQB5NFDO7LJUA7FbVYLBJFGnNj6II2jmMInKQS7T14D5/zjx
xW7FmUvMECrBozUtMU7g6epobpombsX9HIweBZ6Alnm7U8n5s86VaarQkQy5a0qdTfoF6pyg5MdC
/bQ9Kc//CEEDtkpaYdsLzfyRxhZ0g9c94uedNg1Ly0rKEzAaRVkZ3ZfmdAvIB2EQOLqbkMm12gcv
eXL/ryTAwDlD1QHMy1SIWOtCBQFI9HkL/wb9u1/dTAO9cg/ncN1rFppU6SF3kJT8jd6pjoS1yWSt
FUAmFS1j/HrkarOWYaW7pc41aA2t2n3+5PrhsOPPMaazYYqrp0GnATCRz+9BNPtMwVnKZMD4MCEd
RwoKDnMDsjSVwviuit8qeQPw7LQCeWv+7EmKeL7rzsssB8advcoJ6sZIoyIh7t7d+fZHD8Ok6sIX
bc8dlc4CkU46ClsCqHuv9GCBrjEv+UCXfV02hZecEGwXSiLT/m2GU6onl10tKNqzBrl93PUN0/Ux
1EubdyQiV9QzbOauJud8B3YaJZ+w6xtg7wp9h2DwOwJUTvbxPpDXAWDtG1+jpvuCyyMPSmQo1lf5
qy6NZdbclJKxYPwWYyIjmXkuTHh/dvw7fRsgiabTX1bfQRzWSwNOxYGJoGrb9WL+Ca3D03tPgFIO
IRdJaSxDq4v22l0+0014J3I7nyqiJ3JsERUwbX7pr+5QFBvE4f1yj1jMt9lNjzvM7FyIZpERHYT+
gTFOdcLhB/MvOH6WvhCYZ/p+eaXF5bHRGewCBPinYjqulrIcgdHLvEagzysTK1dNTf10CulPHQWn
AtmjWblpTD06JEYYcfEeCaKsnTw8exziu6Kwwy5Zj62ljAUtSaPaeg6AtXvUjgTsiIINoaw50/iV
56pA7kxxKRS7A9MW8RuI3rMkcfXuLvVbAFZna0Iq7vkuW6brSIYgpOWnHT2EVcP+nXXQvm40hfAV
lax38SX6yRPuyLCtz4q+eIy/Mq8gEgr/BM8HxLRwCkupUiOu7SeGCv7Y6n7Vkaqh87S4NhXgYqIf
rvfF/Jpz6R/Z1w1GC07m61kyvXlBMzKVvcDyVNZOCm+l9PjsuCKTEpNxLyS3AsqO0A3xmyAuXfn3
jWJ8GQ1kpNBYjt/WtvG1/OQRzq1DQ3xjjJsw5PtZutID3uXVJdQccWQrWGnNmUOocGyShkDCEH87
sf529EepuS8sJCqZdQHOL7ggxvGgdqOnJS/DR2J5K1t0DaJrFOg6tUMA/sVxHM7F6mkScnuejotM
Irn/pWAhT9WOCoAczmggwDMY4omGa/Gl5qlIXncIlmpWrJLU8sRUZfseYr+4QT5t8XjiG5XRppVB
61HBV/VxAFn2F89DmGLbSjwH1mrCF1UBCT9O7uBAtmubUFLH3zMa0lGJJcbi95UbviW3s6g5XJsh
ru+i1w0Z4533fhgIYD3CyyGINOUuCOQo9uP1VmQlaMAgIc9WcvO2Bv72zKLmVq+gH1BcOvUTzNW3
J/eOJhC/xRspFtrNbZW3Fhi0kYSc6AARr1dhvtVWn0akt5SYJb25gw4ibfIUFmZXKaroX6YTi6qH
oZbkRKRpYW1EuyiR/tuVGR62jnrs3Zpw0H1JVWepn5X527s0n7QO8opLG7i0O1DaDgiUJc3RlUeN
G3pSLwWYqdJ+9Z2+Paei7ajuu5YzM+SafYQ2xtncj92Z13EK3qw8mFRutWjCUYJ1iA0PYTyilK+j
r3pzj+v6ZzojdkT/WaSd+oRwPMN2bxfxS6JYidrF12LcUqeIFLilFyCCmTBD50IPP5M8MhQTtcX6
gHqezR0kv9e00KzPuQ0fVJXpOsxG+9PBm+8Ii9tiH89UQDojXm1NnBN0U/Un2k+5QMLwIBU7FZex
vO5HGt98byhjHrv1aXKbp8jlP2W3LswXv6J3qMZj5b1fkhO5NjxlCrr767TE0KsakaeTZeeaQDgr
A4L4HyMOjguoDEkkFVVeUz3GVCgSQk9dRq8zXwjK/TyzrI32rgXjFQwM04V76vTV/EhzM2virLS0
SA0kIg1XzAwqSC5uPG7cPEfdejCJiGgCrSB3EqnrmctQqw8COU40N+IVLK1ScejQE/HTnGOqtQuj
9yYk1Yu9+myJT4FWIWfpSiDpRHg5s1elG0ZvUO+scr0tRdMBPk4n7mIQJNTvZorAtz61ltv4OFVX
Xem2NBKLAVRVQ6VwYhFD9AtnVyfgpiwJThCufiqz+dnvLOQnpTf1bhf1EP9cE7W49ChV/mnhfOqT
dHs3QOw8UkqlchMOdBf4GQ7nVzewUrJ7OyRB7fevM/r6lemUqb9FFLZCghseUgwaa1tqYFcQQYdr
UihsP5lRx4W1n2QiWsOd+6OGc+tpYfTVd7427xb8+a6mKhFfij2MOidVRnJNTawWjwF6cEgFR/pr
udwjJS0ZB6VWGwunygriVWQidkNsrlNS6QQ9v6v0uuOtY44UFduiCEtOcmSvo7dOJT7szWlFXYad
iqLLL37pkOy5TMb/FZJ/cp8JPZjsTzCQGrySp1gbHUa+DibRnZiaiHXHTLSMVmQdurDWNluCN9If
egE9D+eypsBCCkQ1HWHcdBNWcdPA/ujSRzY1NpNaUM6b5Ikd6mvUcRH2v6mJzW8a9+Ei1nG9ROB/
kGUXwUI8HHwFOnK9oG4rEoXWt9JXuAur7ZhBbZplQHvFVQtvkRGGTlczauO3DjRU8uq6XjEN4hdi
irQg7T9e4KlpT4mYRPcEbdB0NXpgMhcfycN1FYZnXKf2YCKYH3t+Zl52NEUsjUvgSSXh1HQQsiu7
PuE0grxBQ3MyHJwXYk+Eqv49XXFGEEMEWLppS3wAnGUAM5T2xpsjhZ5zvQ/4RSCoxKB0hcj5p7f+
j/RlJJxTJGN1wvK09qF0jFOZq+jnWtxaKvY6WSTQVhX9wf/Z0AqnPbKscuoTu0qKPiVctj8KsN9y
qxLlER+hjyEsCMhxVStYBeFE/amXNnofgfLQIFPzfvr0oQxkV7bD8A92VPRf2bOqCONXmres1Oxg
jMCeJeUggG11/kjCUs5YDm6LbhYg7UqK2nT9efM39zuuhnK2ASUj8LJqzd29tnuR2tIe+FGdHnJx
5dvtrto8/S0EPXW2jfOA5j1Kw9WINHKkrrFp6FGDSeK9lRTyCJaNKc7RF7pCRuX79bMAb5Vx3uHw
ng+wy6kDLtjxMd0HKwc3xsiiySczzbecunoig4rxzCfIMnK62C2YXjSj92dMMZkCcofwWfK1Yk6G
bo0xOTVOYFvyXGvVDZrWIi3IbCHaPWESmf8N2KffZY5xOauefBYMjry9XX6ZG5tO2UibYRdamqkh
brpvlRv8yZDYSYWuWzpDvXJVZIZUoa77meQNQI6PezqQSaJF6Mb97N0xzuyn7OeM4+cLnqy6+MWy
3VRuUsp9FGG6UyHMCZ3Q+kh+MWfTO3I3gFt2ZNCbRTnJ7/dvPpqwDUSbiB2QY8nS/mreJuM7w8gQ
qbgJrc/KU8wId4ePvpgJoLCNy8VhS8DYiRomTBiNDv605O3vD1yoXG6iz2tu3lJn65oge0E4hN/P
5taxgSc9a686AZ6soOresSuTrWvt6oF7uTwY7wNFDdyv2jWRYkjB1AXWT4/BfPIlnGLd+wGZ6e+5
oAR1SJxCbISZDjZZhw5n/IxpO7ZOTk9+H49+kNsMZOoFVg9SyadoKqlH8sf/lfo4kZ/mPJqzBW8v
MejY8TZRb22lQy5uFE321K9YU5FTeOtD92fPIMQfEyji8jsVUCg8iVcNo8pB99vt4VFZF9p1ST1q
NSpwm9wMj2G8M7d1PshJzE8dEKg0PgI42BuntBSosg1P9f6aXwHZyBMAZ28wj2SGxf3nxg8N4cWG
NAx0pLThCmjIVlDEaKQz5bYNMsszVsUYnyW3D1xTSCRsjfpYpxn7gXLY2zmcKVEjH3P+Sa9s11P/
aaGiWp6n/S0cDpFzQHcyU1b1uq5wjzQh2GjYzdW68GiIjBOfEqK3Vf6liXyj6A9XEzsuLLdxBpry
XPhBxNJfVm61FWfFoRnA72DYtXZA1WiLrh63EtQ1ECLnO40m2ed/fLX2j6NSsdoeoDMTcz1EkLUF
G4UT6hQdFu8glGX72p1erBl32gujtBuUBhk9SaDEfgJ96xL6hnuB1XaMc8xEk5HkkUGe3cmQ8DhJ
GdRfs0DCnPlDmPvma2xFT+0LxFjBBMchpNeMd4jfGyKvgtkEWYJ9FSAqrfJkgO0M/f7hO/ozBKAL
0x00QhkcExyyuRH98k8Gf9AT8ANwaf1l/0o8FDql/cJosQ4afWtdVPlXqazqxoobwG1EForpsZhn
HJ+/4AMGybY8ha27f7APBlovmMMgWFWhGtdKVYGy82JZSeA4CBqbqT0CRNNyEYBw5MoZtfkp6xZm
OmzfC7omDc+TzR1vVTX0w8Pt3Zbv3kjXR2UFHIXVntxoRiVvTjwVHZW0nmGug4HIutwm2o1ZDYdd
OpjYOks4DSeUXK6XdsURRrWHbporP2qQpO8IVQEev4SJJySU2Ept0HqkeXdtV51lDe765t5ArzoY
YARwZEHAwwUm6auznxzCanbH7PvR1pp0vy0ws7n9+qosWFQjZwQovVb84pS9H2s/te+WDNCk/hpp
H7Jn704nIWrprk4AW33DpzQ+drliXBKhYsMKYUzxf+FvLLhYoxUVkUb/foeiYgkC9lDFxstDDaUS
BlMWWIYJFrxvK/niwVzK3U/qYgkxQfVDof42Ni6CjKy70hBIrWY88+BZL3TppOk/leeWLHMeD11y
Z1Eko4R7AlPQzJFYnViz45THc+UbZF1wMkVM+UosI6V3czTsYc8nZuWp2tChybF4r7IXmO0x4FFd
b3Nk9QcN9j7l4NxF3ZdpaKAzKRfPWK6oQi8F2kTtxhzWZBJIhzZzxw7pGPVegegxoEDN6mGUmDKh
xc2PIFvcVvzM/oKrY32StgZEWqXdciabDmBrxxR89fBMJUN4CQXec3ade3gycIcGwM3aQ63aai95
b3GEpBs4CSR6yMnrqBYCC5OosQuS6zYmXp1kgxQ7zgEsduIyl0py1+6cP6KBuaVNWgUT2VM+gDo9
XjgnaUUKyTsNSm7Z/N4szX95hp1xeVLgxKnZFxsz/fq0z28Q8Yh5EOsAsXztr0XB00Hm9nYUkAws
GjAMTMmjAcBrjIFDbzI/BQxU12rj3vod9wceCR+SLxKYwqCy5/XLd/VkcM5g0DxN+W63T3YMGrLG
Z2hfo810TeKRkWaCCJTnmf7XsRbD+/jpypGTsHX0EPSFyEdL/87WMqXjm36jr3g5AQPn56svse1h
GncITM9mVZm7sVHk8w/WNuFVGfaKsnaL2eBBQjn+zBjmW48LUENsoCNY+0hiLvEQXM56vMh4MPT4
pwXeD0cLrW96IEXkY7A9br3FJKk8LJ3rYZCEf+Bu6te+7XECwfYvyLinm08gLIZ5VSpTYsrQPxvS
lfWPMslw1k+5KkX6vecp/21v0KqkztoEqTL7zHqpHfkU1KRmz88amK50RznxAeUJFMe8dlCSsv56
k04uIxlX/o4+yM/PKQ6EA3HHFAfw0PmjyTLkq5iphAepHtaUEx7OMsAxYjcjk5TXaYFQ3KVgdOeh
aWNBf3wRjODBOubypWE5Uf6fr/Pg3FhAZ1YR5dZmdRfCFtGhQR4YWcLPo1rtDuM94S9FDo1+I9lg
83rrufC/OgMKa2/T8fKUZTGwllx+v8pzfVjR8SsEsSJarJmIhe389UPTM5B9gatvR5bZGcbAoBKx
9FvivfCYvshAniVk5KNH/ROo3rqmtU8mSpnrbJAQJU5LSwrZoNg5BlzxIvyQwr+TUOyQ6uY75Cv/
PAXZOgiqn1Y+PTdg8/dQirHCQ/pLPlkRIKu3oYYAznfSuehw0Cz2WE/N8gvtBy6jJPHXnIUaxzPs
S6MpYez2/N+YM9nHCa17nkQv366vppDgjqXPrseU4vOTSYDZVgo03YbXIDFHYnP8CDvpnvDQv1W7
bWTzLLw4dxTpJ5SAp1W7cAzc34PQu99fXJ0Ake9ULCmVlOGgrc42GwtXjPYRzalrdDH9tPZlO16l
JlaVj0PuwVFtIUNjE7tt5r1pQj5AHhHmHhPX2gIShY2D1K74wssj0Fm64otXaupAMi0X99X8KZKI
AKbF/4I/N1N5Cb0Es5ja9IREc2JBYgo7BeKlxK6d8OfxgTN4mu3v4SM3YD3PJEcGgCw/KHCD0VkY
6Oa89+bXINfywSPyloNhhUSSYU+tE0QYg7QT9poU7lkj8iF+R03zyMH46OHzMgS+SF9tZQ5G7rMV
EcmITQy7hmrTAPQrk0GhsXrWZwUj0xDc+5kaHS/ybQPV1z3c0OeHq6ULZAZoyC78bAueoT+YEwn/
Gs4fOfc0iJqoSW72b669op0wFkcAp+I6jxMg55tRtBXzCT0riIHn4GvnhdozvzN19zJ7mCc1aCaP
2L4xyT+NRpNzNIAaboiKG91oO48sW7QWe0sIhaEcI66GsNMvcOrViKzHGQDoftud4PmJ2ctPoyXt
kUZlKPyoJiP47zFtf/17OgCsH/LpEu27oUL8wMOqjHL0HQf3buiYNBsWP9X5Qx9kbNTvdaNg1Sdh
pGhBHo3MgV0XqZoy+s5+Gy2BynoM7/iXotndv1ptqPC0LbnigU5wEFTYdHvwzGMQjHH8wSkLKR6J
yu088gb9IvGfuH0ZFahgVaqcFpZ1ADk8bUfSwvKgBM9IN9Rko6E0AzAoFNT63gR+0H3QDgI8VskC
a79w63mzr/Pj5n6DL09ehWTKyq1n8xAtYy9JgobUAs0m1usGvQ51wEknunRkXHAMDr+bhjvoXD1X
xe1OOIqVybr/HvgPOe4hNrReV1tpcBn0TYT2l4gAA/xgRwjzA7z+THe6r2iy5QDWVmbaplaz5RK8
nF2Y+4DjQhMgAl6y94ubDvun44RuyF4xkTMm5PAxli0R4uoz+MenCcayqmyt6GQqyny66RSt1AVw
Kzi+8Ee13gzwPr6soxFTCVKu8s0zqlUDw2zW25ch5gtzSyGSplDCViMbaSOIBOp7MUr13s5NkN+q
UrWGa2YwRugw0PMB+wioJ3lbyhYBskni46AG3oy3PQNmOyJ2oWqSOtqfdUjbzzQGNL5QERIPLswi
z5KuIMjAsdIFYXje3mbf6sgxWCnGeEjuVBoLIpGBh0ErqVKOqBTy7UiawgnQ1Z6umvuCMCYN5F+E
d5x+2KJqZzVySjSy0NFgbyz+Mix4bew19D41B5KhZslsIRfkhhSpuFkZOLykHxGKRNw6xcxAiNs+
IvMtQm+wlL22xINZn9plSs/U/HObuPoOA1VdLpBRiDPGq0C3A0LzP8sPfTmqGRyZEvd9OTHqYtZ6
FZsEuKyepU/8JrTuHA65IsW8O9fpk1QvSI+sAJCZubUzB4DiDfhf4kcloMI2slPoaxWY8YX8vc/p
O4OP4P3+YPSTkbp9q1K4cF7lpEkmYJEtvGYNeZYn21SgTatwFN2hzWUgnX9EQ51m8bhHrq774XBP
FDyOOwFz6eixf0b9aLj6v9eAR7kciyzDeoSA5eKDnbitekkP8Zqdpo8r3CRW3aUN06qnB/Ql/QHp
G5YCd4RGf+iXbssqrPSQRa+rA18LxlHVEzcfvN9yYlLtRqjdSGeq7BbhOwriteqcLyCymEqfraZB
SunZfBWgTzeSlvmqK/DdS0uYGs5KwFNb8gQ1z+YqhvT4sf0k+4lAlz+Ewu77eIy701RAVdO5Vqut
cZRiSqXieRpn/Hg3kFR1IZb7jSTrzgsDDehO/JkyFLof5nYGIhskPkye2IpnvuKLRum09POvLSMx
s3f6h6vGQVQBVLGKyYwK5uGfwKSB1cDrw1FrhIaI5/UUm3WIYjqtRW2ErcGxFWrUTzrieg/1JD0f
IniaQhG+8tB1As94RA4EDVK60q3U4HJ0y88NT4zdRdSOiBBVvwaXrB1u09/hmVKKotxJaEY155Xc
epT5H7PWhvo2kuvulPtwovCu8gH/YCyxkRksUR4plXI0cA4Ex2RIEBRwgxY8wOCgq/PTCypB925C
50nKoZjX9QiqCqmPbCEs7LAJjin6iG+SE+9tzQv5X3SuW9lwNYSToSDBk7QTNiqmjTKZaDAei4rV
MCECOEmRj5CwFPrRI3fTTPBEL4WQCPOdR+ZTmBn8fZKrQBP51lfLrRDoolMTDfSJ7Snc047ppq2n
NaZ1unJGSFsbVLErjqkGxJcg8Ezr9s+lpkuqRpPIMl6JOqQ+iFoX8O5GPmuGMVia+R93h4M4NXOM
XdZwRxQjlZlkZFC04lsrokNjtkIRBMRU5QB6MeNPUagGKrmsDewn4yPpr7C5dtVUfV9n5/cWm12D
M0Ta4Sy3b7nlPo0Qm1FlktDgJyMH+7F5QtGrLgxYBFtdguLgd0wTAVYk8iNUTOKqrhI8JGzm61fZ
om6kqmWkhHFbR8vGmr4O1D7uamUui/cE7Fq3fSLZji79gceTU0hk9pvPehnKoOCOuf1bvqbGmzVe
UCtzhbn5kZn+5/d9jS+vt9oTQJYomo4oSB2Y46/uoUcVxHVTjigAQhARRFuWRSM+r82tnV/0Qtco
XshECAh1s4MKbjVimbyYklRVQzWvcudEowHJDwuliTZccBcGInoRaBrE/aK/6yHPQclw600//xod
7mVOJYLcmnHd+goocO+vJVoV5owBSqjjCsZ3UX6ES9YEQ/WOTqiRKkigwnPMuk0d7fdlOUxsqrsc
obkK5Fsa7ibJ9Uh+ta1WAkpgVyHEz580IrBetAB5fXSIuBeDBhXVHMlK0ko4X3VLabevfOPzz3eV
ITQM/r/gBrvd5XMniaiWfH1HuocMJJWGkUOMw1m6K52SBpXVhwRofAhXb/k8RqWOouv/CNGAXqaI
OJ3lhqOC3O5AmpXPN0g/aAUWBua0yZMbrxe+XZTnJLSOCduzCDq9guOdXEcoKA43d8YH9+a58Gwg
FicheoV8AbGtJZxcGABvir+mhje+tlGatX+fSLaNiMMEcwA/ExZ1f7BTY8VVT5jeSVmid0oIKgJk
eoR+alTLdsdoy9KKqhXOOP6y5lIzXg8XuaZ7wtmAC/SNKwPyILK1N8yOLuu2GTxz7Wu0m7TDCSsN
fYNLhJ+FqS/4BMa2w1zhJcVHB/JFGwhmYvQs3RTmGA4YmV/T+JQkYigLL3HDYmPFVV93lerfV1qb
TouTP1V4WRhztd+D03d+ICIkzqBa4qsPX0McGyifgKTaQz6D7oiy6i+iZJiBhFXghzo4CYaIeDQY
hlsECMkqCvhG9oZTmzXnDmmjDmJUJ99M+6pDYtTEkLO+sBqBs+A5OYCfwqGZ/MOFo+U4aqdBqnTi
583JhTxzgXrb+vHm7GaXwHigxPDMirD4XnHMYLu7T+DIFCJAhc8fp/N7qb82N3gC9yK3AuPvOhOg
+v/Mblo65eGg6CkglI6b5tn0EASbTytsGqs8nXA7NxilfUZZYyH/qupIdeYucmFbjobxR1d/Y9Z9
o+19/kJkLBrOSGyIn5g2lgQFBgAwFQcQCM5Gp2SeQaisoWb4i/20yRt9AYDID/XKYoN35/eZx55Z
b+EzR6o+leHYRA6dxH0f/tTa3YhkNd+jy1ycCaI0wJc6CZHabk4t2jwSQviTPHZANZS5yqDT0L9O
+sDdpntRVs0bY4RI7isnXOcXmdHeTZPl3Cxq6wUJBpAq4sBA2jTyv5ouqYAz8+QlnejSfFID9INw
SHjiN2/hziU+3Q+DBlXP6Fnkbn+W7PmNyBe0V2GZ2HvwReSa3MjGIR99EHYvd1GTr517xljA9SLG
Y99Az2vpU+qsj+20upRWI4uAhgV3F0R+5SqzAZKO1pT6bpYGnMlsxT+U2xipqa5FDdTN8zP42rrl
6YWnKOgs9d/VAl/ONXMFxaGP2Kl+1DDf8UT/D1w0Hug1H2iAkQXHWybMSM4LtKMMClZN2uwVhYJQ
ceyUjSxWBylHe3UkI83LShz+qFYv7gvWA3xrBR9QhT4jUAozrIb0zO03S7hN8Y2OyeraD99/oUay
CIhQwllgoGIs5PRTDmB6aa4eKRnqQhF8RhbF/pqJevdPsmH0gvaV9rIgauhEVHyESQ38o1PlOu0o
dZB6O6acZ1hNblz++9lqORpyHbCYryvU7ubRze92OqVi8Z2JuoVmnXW2RQn/owZKdBZTdLvg57a2
MGcxTvdPM3/aZYCHlgQauMBiHHfpQ+9bhnXXjh0q65wCMAAHN7qwKv3If53DA+J0zcQywD0/fprV
/gWvnXRc6QJKCdg8Gf28leGNZAJVN8utEX+i3CKdRinKNRlYG/n7a6rYUMMHcqHfmnVWEnYGF+wx
zvYKlRbNdhGHUUzussbc5c5UoEzCyzwSKNLpEOFGKC7G2k/9UJ3WC4rNHvSmhQ8ZJndJnOABqIK5
TZDASxH9TCeZOx1JyijBV7TpxFIbHiLRl61FwDcjGp/BaUiQOVFaSOlnJ9doii8GeLviGfsdbiwk
ek0TXFso+b3KsW4Ptk2PLE8xS5bJY6HERNi/bC+VigwclCsL0OPjxJyQWGPFrzyG/3Fni8zIWUn7
o/twgZ+CQ1+/kC9A3KQruTtD2/0ZUVE8yf9X2nTSItWns2uXbv0fRNuOhtM8lYis4McfWbdMfAZJ
kWf+PLDGM90Bvkn18xKP/TZ8CD2ojfqMpnv5HBQgVYg8QVQzzmhDDo6uFoSp8xWb8RB05XYKYURI
BTn/Mg3j/XrQ4cJYZEKaeQH26cvZ8zjCicVN2o3eD/AF7TSgWbZ84GR7zVLdS89nfAphumfHkaeR
h1cFeOqrk3UX1EMw1/px8m7MEQiCbaD+e4QnsJyT9Cu7zhEvbkrpmPT3hErYMiXJhM424Oi8UomT
GCRsfHQXbyAJJOC/c2lzeQVewT8bSlyMjt0/g/XF9EV02MfCEr2wzRy2U+MUy5enARijAdNdF+74
MUCoZh6DNjoNCCWcLmt2RnGvAP57OPVZcUEOgIFZ0lo9jM37kavGW8YpIj88hN9vOWaWyfp/muv3
QQTAINKoTlrlpgb73Sbx5JnNu08/y+d7SbX6i+Kys9nYGQ8Rr6BnfjXILXNIjq964/gHJI9K6sK+
806NWM4Z5Ft7af/P1CjPqkUfGJfegdqTwDsU6PXz1/wa9N1x3zRsd9pFmYS6k6PVAO4cVP/5rHI5
gdWRb89nrnonpfRJTA7H03cqdh8xy9BO8oEnugzLAwcrIODMyRQ9vR7ipob45nbHbgjPABH1Ma7i
qckHOq4auR/ik+LVaZwVt2YsQbyqeuUplNVV9vMi8LdI1PPO3crrYVBLNbajRNyRAnGympdWvL2k
i0XkXoiCdL5rh5uBLAIcF7X0QBHTzOSDACQ8vvV46ZyK0QWpCoLGqRyvWaNX6iMDI1/2iaAgbGcy
GSe70E9/7qqv9A6SuRJUX3utRUDQI0N9+GSmX+Ua1vgXXhYNI/J8xQcE08gLrrAYEOa9116K4LFr
bQGd4VgUO3gpjq0YhH25MKUOa+qbaRVj1KPpYsgVpmsvuhLXWm4wdt1p+59nuM8+5ydb0Ft5lqOH
FjeJHAcu8clVYXpJUjvy9mvEctj+8O3tmTRsoyAXKYvSAwKUy+LaQqXdGG8VCxp4iCaEoRUtKU1M
3roME+3GnZA6L+NS1PMWzlBMEJmrXIcaEPW1S/6ZBi1s5TFzWMQkEgRr11BT41Aqyzs/1Es2gxhJ
Daw0pasnzfOPRWFX8rwrwIA1Fvz9UpzcaLiJIZlyutS4POtiHUP45Gkct6g62CtiC/wOQD6XkAqZ
wKun0G7XBhSuyBkeMjYrlCeG6qXk8IoyTWT6TIZR7gqTv5DN7gcOH2TXu0+0wmEVedNt2gsENZRi
hztSErCV5NyNtH2faUpF0Ee4qIY+JYgqda8xMLbdGQxeLJRPZI5h5N82ItYVuhEtW7zPRFMde/jd
cYq1bV9k+53yCRbTM/1uNJmZNV8A4W4qFWC0B7W3//Y/FUziLq5QmKcjPE476/6LGOCbIwz2Sw8j
d3lL9I+73GFdGpikICf1XvuB6SnYK56zlU8blDHbIrq4ofzzXswpmVwGFpT9PnE638ccEDmnxKtg
sPiUdXuomk65Id38H/qeNwxxXOQqUIYyqMSrD/+gXQa2pdUBhLMRUJqDYvUIlGiftBB4V3ya39xO
AzLMr8OUn/mHXpHxVzTSDIDFHNTHF5iYzQpw56DgzcyPO6OZxl1YKWTe6gRGjdkxAq3LULTbeixz
LYIZU5LR/ADEV6syit++EaIPif2OAl3KmzSUwztYGC/LBWhFYs+vJj0jk2vRJ1BpR5x4E9U3exqU
5qJKXlgctvs1cv7RWeopDXDsTUsefj7MV1XT61fLocK+AOYgePkItMKUEeFIbeUuGKAb6GSZlvki
LddgVkw+AwjDQItyA4VDX75+ogoTWfsraXSSBB2O2Nxe6CGPptsrSQgCNXh0sfORPlOACWuY0uCy
yfXxLuifUD/4V7qcCsK4Wq3nWUdwu9GuY/G8bbLaBAIj5fWZINPPNhsCZavyf01USRsvzghEinUu
IjP6ssH/75OX10EhyCiMH2UNy4tuCkG22+Nzdd/j6RFDrVOqNn869/kdKPPeAxCgt/ddDKpGoXq9
t2yHIDgejLbgsxU3kVQmwpXP+CQnFQjnwJ7YFnZhzrl53WqVkHVFVq0oxbsI/XNnXZbx/2QFc5E0
jyqO28OFx54U2GQcopl4MwshHLWHkF9qQtDwVZtZIsqvJOoXF7c/G8/35s7Az4N7DVrArS0lNaqb
n0vXVgExfmpYY0EAfJ0+K8WFsQx/Fi74N9EL0XUOiEXxets2zbE3Hmro/dt87dMJMyKfp9mMjVS2
EjOnYdSiUyYP4hKjWeB7K70LBljiQDgdDXa9jSXkfj0LO9vechqtSEj9i0ALJY4fIG7gDRmx4gCh
9toyb8rrHOq9Un9l7MkP4/6PPVTZhsCjDJUSPgs91Y4MY25sWSEiPNR5+ocQsi/15wDiD0ahvvKT
G1EI11hPhb0jpEaTHVU+jo2T++I+rCWqMPGNK1TNwmnJib7tTvSi9jhZZZ9ol+GMq7dHIuK2szw2
45mr2YlkE5VginmEWF+RLYq3S3WeZoyovURUDlh4qiElo9g4XHenI8SjOkAT0opiokx2zO8W3BeZ
4tGPFbMENM8f5w+e9iZTHSJBmuwlEcsa/pPgUeT4bui04TisDyt7ALnoSoXK/Aja/VXO4k3uLTRw
Au91R7DQg7p8mDVILivGPG37WCVK/OMpJd0A01k8L1fDFBD6mKEomh9XQ4kRHAbpVYkUIncIq0Yn
xNEgOuBn/JYsSiSNeB4Y5ED+MCiek6Ana2JDrW1laPsD3nsCJxHoqPITRcJ461YlZCHzwpqiZdtK
3gqPOuimWiXSO+rQxHFh+0hdVr80l/hT/4kKN+hnx8ndSaOEEasNyhnoRsU7IgC+nylE3PHH9Rjb
4kgSj4qgabwCIAcrG5O0a5ol4hLtX9CzAB7fDdGXdb+MIO5/f+3iu7tK9cBcpU6kHN/hBybNc1sK
fs0j3EMEjCW7uF0LNVrj9p8p/3MXe63oMHHR5XaAnTQf9y4a7ER5gL38tyAIS2eL1uaxolwxA8xO
U1fmsE4PmU4XYW6JozbE0z2YmjewLMZBlk+RB9OR3fcHrpFXYlgIig9MZXOGbOHSWqOdxnrS1wD+
H/lcGWFl59WSN2mW+wdh4IZuTB2PnzXMQSWNyQ24qLlEurVWtFNCHvCy91ejccc35ANNDozoQNyY
zvKGUNWIlhyv30doby777xae/NCnzrw8ivYQQJ0l+tNohbaYdhOu55pMn4x+lvAancjuPffndXMl
crhuwrG0aWC0mjTGct/cPyiCX12Cy2Qbh0LY9U/kCRwDAJUEYqRABq4tCFlCDpUkaJ/Mkc49xfSq
Xe8QjM5YDDUiS55j05CV+kONdc3gdIEr+BTKX6MeUMHEIA4nIYdqJqQCvEf1WhyT78IgZqhcWw9c
x6qGi1WWIjVJTUcxaof2oVKOabWJifKbbRN4KfopxyEBCc5wAa/DBIzf3/lyhdqnxVidvEKUKCXt
pkiDDz6+9KuZMAVoINMV8SdaCW1sq4GYU6XGhnB3nqHR/WfmyzfOpeEQYvYfnq9fiuwp4TWo6cl/
z2ZSn1R7f7Py+oYPiEPS8/815bugfv+uqvTrLNhfKTBDTrjQEsPqXJqA9HRyCby2yaaAHFqOetIl
sew/UMDk5IvWZ8nCDm9l+6NGvtMXtL2cC6yEi2qkLGpyfvvLuUPWhFN2m6qSQyy5ldsEqMGIkhkc
6rATa/uhn0rTWMPwJcy8sCDj5moYZB+n9fye0ER2TE3NwT9Uf1WJ5pqoyMR5tG7KuWTOaz4LyR/y
piV/3TOfOqbo5QDofxCwGn5kuu/O5WnJcd27EAgj9S+E63g9VzNrknDE44zrFKwoVXK/XDi2SRnl
k/LAQDsOkMAoJTEQzQfGWuRUYvBbsa1hGmt5IjHlUj2V/FWIka7ZK/fS2EWvoMlOR6i8LJlqnnAE
kwW7pOM490fiiFFHN/tKi5y5nNUzA+MeNQcw09CLJ2Y70LnC+L3LBJstXvCfY9/Yx7Xs4Gwb4uFk
Z7jTAfjQnVSo76NCLuU8ou1gaEwt0evYkrwVsLsMSmYTunXGD7n5ZuMFKUj27JULDdy0UfZmeSw7
YoiqspXuZTB2rb0ElzgPzOt50Ou3ewmG4kqoeFizCpdPiLAiraActnz4wT2Py2x4Qleea8U+Abyl
gnWNTq0lUaI7WILlByDRtduI8wLbkEJJeX4Rmphhr6x1GsJBdok6MjaqI94vyYEBGcQ23FFd0UcE
5ehBkeY8oXnYh1YDNMzaoY0tnmzcWAiZQ7iJ2CoggAuVBpe5PvTEI3vnKZn8bBtQhvxxdG6eomfw
99CH65+6zAzCVhQoRDcBVwNjGThQVuBynCz0Exp0Ky/dhxxNPnQ4XI1g3R2gkfR0zSGOxCtM6Rbp
8ZW8f7woRR+b0l8LK3UwbBglGB/+2u31Y2GqT6wVshQqQR7Nv/2Y5N8Ei1KeM7LfScNQAt+6wVRz
PD2zROggGa1JJ7WiJmn9JmJdpek/RzG9/xwa0Y3uTPs+27MZRnkP4Mao+AWdHIKi/aoF8UulCyNL
8OERbaRiVA9qXqSZRDp82jyOJoK/lnHOZziMaNEnR5Ycvl9ZzBXrBXeX+Fin8IxN8LXsyUs1R5UG
RvfnGAGr2hHQMVpareis6wWMqEssNJotvv0nvNHISF5Qln82He4bUFFdx6cwZ6FxHUlia4ITlJhL
AqBEP372Uvb9+wrK2LrPqBaGT2NsIQR4Xf7FGdGISCnovs9fDKd4dKjJ2IReIGo3lTOLegr1EQ4q
TNiELBqMUtO9JVH2m+uMjAudPpQks5l34khOLnC5d7oWL1Oo8Gwds9bwk+YdQh1zQxT1DNC8bCLb
+GLv2ITztO+0b95pJm70meYyM9Obbxs0hYZ+Ip8cmICmBntda1ClSYgKmiTmZ7wDtSCF9SjE5dOD
/5SkBNV6kCUNuaXjwvWR76DNFiYaEcqxleHpnTOjcoAVU+kKs55Y6zQgq0kZyb6c/BfkHPGQj8qG
28WmtTiRGh7NicSskUFmEYtNZ8PXTf4gosjXx3KM8bOZDN4auhl74ObwPtJIrn44L8zgL2Pqq7Jd
4psItUDmBGqT/TNXch3MmLJlcd8Ktk8qAoZtD3KvdBlfXwmNBU4Gda1mWrIdu8ehKoUpAd6M7MeD
nJ0xX1QIQpJ9eu0O0qLeNbqp696js5ZA43+8GB+1FblU+Td4m/tAiw+G4GAs/bgc1qh5uuNCSisv
u4KwZ6SNfhSMJ162TUElZKLMxam4p9lYnOgU6CK6GvxhzzLbqTLZuAf6to1a42lcL/9I2qFN/6FB
ABkfu2jZwuuoYwtHCTNNPnO9rmePAl8Eo6KSJn/iZMqhcmZcK09z0gG6SS4XYtaeBv6jr5pmpC9P
TLoaHVp/AIZiZdm8qyrQxZ85xsy0BLKRx1sRqlaS9l3QN+qxD7/0dnkah3FsW2ut1zEyj5Gyng42
3z85hWdlKD/GmLxyqmA0tuwe7g0J2uIAejVmcNMOqNw2nXFEwQrv4wvPwQHqFjK2B3PwL6NTjYNY
zYzUThxhM92ugGJW4EQmNmFBa+7aUni5iLq8mMBPkZ9gHR6KqKnac503A5zZF6HyUf6HLJfq6kp/
Nfsz8CS8nJJ7DyC1uwJcDVViSwjYQ/EG7Hq1HM5WWYasmFws+EumtfSzF9TtMPDNXKLGUf01VqLL
XYhulmvN4dNeRr+epz9fpdFLYf3lZVrIscRWAV0kFrmYMly5GpjxEv3mSbjmF6z69N7X01hP7M6Q
67aL+2HkMGAZcWdzKZYX0OyoeVpWdJwNJ+G6Ks8deB5+zotmvciAKjTVXNRs8mVQA2AhHYSbGrYM
0B8BwkPo8eBTyA1EQCqYSUtlAjdwy1NqmTM1QpdtLylJOKuxiX7gP/4yVPBF5OgT1iRCwIA5U4/G
dV/W60ukeZKfu+hyeCssd+T8tcMnDLWjI59v0+VjRWxi4aAB491Zp8KFtaB3TBtw0ItOGXNRuuR8
hxDDzviTQWSEGXBTep5/RUG+3JFXYrBVGxl1cck3ckZK0viqbCGlkhmTY2EZYixthLW+EOxFrl/M
PvuKiN85RYcSZg9sxIZQxwcC5KHP3w6HNrrrj8wIajSJcNVEfvoIxxwaAVv/8W8WpBBJuGfl+bZb
Cfhn2OX0rfiTHjGrNecbBJV69IwZH9BZCtEUi2qjCdnDMgcQ0YT9ezNOpTplb4EMo0Rie9lmFHDn
A54zcX/qDi8z73LReh7a2vhSfgNNH2AczVoK/ZM5RDeZF8lRLMv3R9CyCuiKqUze17tiHB+asgMI
LcR09lLpiYoaaJVBgqNlW1hAH1NwLf4afKtNvA2+isClxs8WGN+JAPX1UT0tN40FDxlG++mIQzg3
00aYYCflmTz+IMTRkb0JDTCBJtGxh9P3MFyw6+GAAowccFK51kixWrkmBdZLMUzFPOKQqatyBN+V
hTxEkyXEAsQI1CxfcrhANigSgNtaZqNIdlbCN4ModEaKYOth3Q0CJX0QCFxQVBmTwtIMJ4VKNfok
soCTGuKFXA3kzja5DrB3tTL10AAMSAo61QrnTlhUX3uJ3kw9IO2ntdZVsxViFLGKUhHVYMkwu3g3
8g62qZMjbBbl3wbOMB97T3oJ6UBA6Kmqepn1dndBjAAH9X/Qto7KhAkEyZSpWmScq1k0DKs9AjLB
6VZnyq81+ZD4hStIalJMEt3Ugh9TZxjcU5h7zQfqqrcva5pQumNrYhDWNaKOkBjCd4IS9yemkNsL
cfaDFKBD+xfyeFfbLs/9RpM5q8mbQZRlMlkd5So60HC0W/Rg+az3ca2kr4nYY8IUqpuHe8D7hEQx
RYXUN/t/cpp7L5laFE3+cJxr1hWnPCq4wINjb/pUqn6HrdnHEMqyDRgGXfiQpbwWqCLcUNZcb3LE
9k2MhVveaJ7iixk8gpOUZQ5NHuhbr4CUrCCaZikT1jzoMCb8ff5siUL4CgLzb2UhXgVRIRqSWcI/
2vRpCaF7iWX9kB4O8QU5GfItRAj7MagLc0EMB7KH0GTjXHjOqLsXFGZpfYznqSd5Ba2ZHlWMF82E
TDVVSa/4EoenZ5vZlcWTKLO7B4RPCmsJe3w3ONd57MLadMVp8HouvvzNIhFJ9AaWTL6eDfnHnpTP
PQZ/EHpwTeFblFnRzvAUMJTcGjDRXH5kGc3LPsJ96o7YFKCPi/KrNCOHIkZpN0q4xyZmr5fdGW0N
yvOUEITN+cgFJkD2/lxqMi63gZtGeNo0tQOmX/rQAN5DSH2PU14niloh7wMR1QIpo6BS5zCMwmta
6+foXW4z3LaGMo9uGPsiOYrKRzDDDZ6Zyth/Ikt7jWmvz04GJvPagRu+f69GohX5CgCqbK935ngx
kCfgnitRzPE9OahH0RxJapLM6gVgwuIHo/yAf8zYZWbgQadZAZ6xMsJnayZGTxXj9+05D2iSTstX
ya8BNhLFh2kL460g3uHy/oH+RAUq/0uqGJ6Kkr5ZNo/pUhgBAlj2Y9eXdIJ5KD2nGiMhorXKkHRc
o/+HJT22Dx4RJkLEo1fdMjVdcmlvtwxnZ8QPCWFbZjhg8IBIB//XSUREfP2G47VOuZ5L6jI0msWT
fcVd9iqV+fXK66H47ZqdpMAbkOUqz/V2OCV46BGR1LJY6mFTZl3I3hb86MWBiZOI9akwwYo1pbIx
mOejytg7n1kpMsWMUd3k58LpyNasxuKjQwDJ2YgERjP41c6MHUomIwaoIk4AnH6/g/uwg3B7yxOS
YhLw85uHKUkKBYkdmukunyqk8g2dR3RpJCLQ9i3td1nNuNpXy7DtRdch5ip5Q/vkpvieSPGDSgOL
CUb6eTqMk8WlLyxEb8sDPouwpZUFyFaiISq0eV/jl249eai3PGyIgiqpKLzR0sTnLCZBi4vArWgb
NyMfDm9nzLBuatlcVhv+ZgfmxDOaVpFgX6+WFLRjJcR5G+Gl1gvyhHDobmwzg6g/ZAJRZCWmUA8F
6wkwvv5+oofH9kOh4n90t2sDGy28Jp6ZB0Ki8F0jao9M+Yid9TvVxn0VcCb/SnRROv6gLXq7/opz
yxVAX737OAoR1kYuCRzJhQN8HLj1naig3EG7cDuNI9m/f0+x4t/pSXZSKxbnitHunQNPd8hMS3DR
XXqigZi2RWMR6BaTvez8sm2/WeP3qE2YvBVU2Tn5Ds1Y4sYalOUJhNR45TeWtj+qUoWjYDHk0vYT
+nz+uoARie3+e2rkXtl5+RhJ0IRLe+msBR9umkhv6Jn5N2bnrJACVmJZlw+QYkIU5SvBNijLvXLM
YiUTqJMscVjuzLIYMJtCckfWRCUn7xL8nAh0acmvfxieRGa7yvFT6IGQ7ML70uJHDZ409jl1XvuE
8shx5RnXTaKkGkAcgeFmtdBdfNs9W6GaxewEKfGtYF82VlBGcFmAngh5u22SOGMj7Q3wLo3RwRwO
8fei5A7NgH5jPtBuL87X3BczG6M2QC6RoiqeCGNcqJdVuBTiZ9m4t7lCYoUTausBs8Y1Guh4VlyA
GWbM6FonmG1G2nDDohwENh/9z4jGeJ0yVkObjw2JSfi3uHvRlglgtdNRH2Jscn0RYGnaZ9BvO8oM
3+20lILjs4Svhm+H0+RvvYgockPW2n4fB2sSFNYlZSYme0hoBC6pOZucSXoDzbC2Es2UQi7hS0HY
nachrdmdVjG7xQEUxeDcrtVRP6wevp3cktwtHbjoSjADTJtEf1WGUwmCTARNHABxaHrClXSq9mE/
3WcG+2JRg139nuop9TN9JcX33MkAUuDnfH8uGj8BbtAgzIImTqj5B7/kO9Q/t85fFGAwHBG0uuR2
4IuCP/TUojCqn8QFKml2qW3ypiNwLQ1q+zdJeBT5HDHuE5EEtB121DW4WUGjHY8lpL1UOqvBqodt
VtcKSn/SHZiQnq49PTIakDyZGp/JvpNEn+nfkBXOpK36OQUWbQ1dPj784RXuRSvEsmhbyj5c8Re7
t75McORBkRA0YQZRNOfprM/4GyT/LcaszydxwMqo6Ejf4JRLoLb3ReBybfcT3tUGOvZFzgoiRuW4
Ew6mPArsiwyfk8k/VORHZz185y1+KAVdaiVS2/UwY+9147jcX3L3TIYyoCy4nQdfN5Ae+ngJ2qZ+
hlC4aDp1MLtIFOiG5/5vw70amKJ7HCrR6L4WtP+8UnpLoomddiYsfpailcswNKOCG77ccr6cOF0F
EmFzRTN769/SRTjgq10MnHdZzXLRtrmwOMFc8oscKeCidMsFY3ltJJu6hpxvr0Blr21RSylemZq5
zTT0RMJrcjqJWoDOd+DzKHxYZdkEys3G/GikHZzR5IEAMUqO66Tb3dUeXAYdRZFqFvLKtXO+hnyn
lZQ9YIVxgLc4RI0Z8WAePn5JZeTybX38QXo/oekmTMOFPEz+QLxiH3dCHjQNcYKRvKoi0FoF22rp
Fx3Ih6h79XAc7EN5XYWBKEUPaaIB9FLEfnZIRAn/WqgI8gnR/908vhievVUWGt/UFxyoWFzlH37I
u+6eeDswTwUf45cARWyM/uwgTN/iSI0WTXjU/mbS/QCVolmfXLrSr4ZKy0fHDWPsF23uw32jnEoX
8jpY3bvqg7tzFVGmfJfxTXW6qLb6H7qhLOFBNdDr94uyUoqalATV5KojMkAHhGBGzxjzG42tQXkS
agouJnzhgPdNYUm/gPH3D5HWbZMZ/n9NkQh+a4LDFnTWXSGMmHjYsUnXwlOPjNgcn/Oj+kru1a0I
nhHIy0w2p1QGWBfdWvUZBb9AelBnSa4kdM6uz0zDH8zIZEOYeCTudlrTYxjSmqMBIRPV5KkpTQnZ
IAnqMkKQJ3S19x7yrJDPaiiDQ7KPWe09j1ncCnZhYi/+++OSsRvizbtZ73lc/i/Mkrd0hHPkyqhW
thLLipPbUQZZIo3MWV+kn+UKKwMkrDPl/GcbQZRX17PMFishK/+7pbVjLFnupilutXnYMvxobl9K
zHsX2rVA0UvgU3y/rT5arVNXH/BhSOaGlTpkcPt2S6theQjvUoqjKcriliq1ub99ozj6PAM0DqXQ
oziaMxLAgvlsW0FeNAYNy2vBbo97tOSbi4yzWY68usLHrKG1im/SkYBj9l+zMYXW2PqLC1WvA+bc
gOVk2ibFOi/5Au51LhqKJVa/hitxptSzHHkb2ee+ghI2Eh5AsJF52AIjtw7Q3tXjtP6C+pS+uAJX
pe7d7q/co2xxjffiPkRL2W8iP4r05gaPmcHy59Pe8Juhpnr4T16tJqQ3IHQ3ckPO0OkJSiiB7AM6
mN1YWHlQ9TvkbMz1n5BCGQ6FdQNoGWpsxTc5pLG4G5zBTgPpDURfJ1fDGDBOc4xUXk9vgQ4I3hMM
rSvGgWryF+rmzbXpqK7vPUGB335KOLDzLBhLEw6GXKiSyCXe/PYjBpeX4t3gKLADiqnIGkSMkVWX
cSK7GyUN+W7RTQbT4KPZS/SrBR/A0UN/GoO9IJl86Gvw+93y5jVnfo5K84mx42qDe7YnN/0l/M1y
uM4H2X99S92+dK6/q7mDM7c5URS0YX5a/orAQZEFyQh9lCzcXtpMdtNXDWDFfVX4HpTgTzGBnGOx
uSLfkvZHdC4luc7EWlRAZgZeVMs9RKAKxJ0Dg4PdwlDIAk3j1j5M9bXdRnDXoYIkBvAQJS7pEvUs
VTAFl13Tou55noZaRRd2DzuZ5D5jx/lCz/5tHZJFEQD73hWs80WuIthvzmVJovdjaff586w3IGTY
cHu7aQzu+l/j8LsNuZadW3v+kjoXT95L2eMBa0nwY1OEYlMX7pkrkImNe1QUCvVCRrdzih8shZUg
xwqqPRzvZNEKl8JR8HW3SGYxtSs/eDcNXJhb0JFGQbQttp3IQ7xXBNJxWYmMx2ygyEOvgnpNPj3Z
6nqxv30Skwl2QtypSrySVA6QQfjIMlXnykP2kczCO499V0t/s8aHyr7tLXK4LoXx6IKfxsNvk5wf
xopKA9hPvGw/yRJb5laaT5ZMIEgDD8rd7eLQCvO4+8mbG51aVEbYD0Pzw4WCKkA+8NDUFyoyaxEz
Y825aVU5CFhsfpmxuJFgRNSO1cEHvYr+BbFhuUznvCvqeUy+1w0yukPWR+dQkwtB3VYJgEbTjW72
NeRZWZLk9qHZkLEEOOzIWpLsBLtwDgJWzSt5FG0bjspm0UytWYW6MTve67DgdpyiTFqUsZ5847Uh
22UJZrBfr5GK3tQyTcL72EgHE/U5O/TivMpzDD8ZI95EwHJqPR48mFnH2GTDzbDuU9IXPVTyhH1a
PrtLNJ1yZn5OhyQ1pDosWqytwlIScw1lnhU3R3k/p+xOteW0YQEGIRXBaFq2JBRTgYZKOnOpd25H
YZ4vN7WITJG9uExjmX5cbGJbVWQhpQGTokdr1CTP4uUMrGpzcgEdAbtvdPbyolAWdyQpj8YP5C3m
1mw3Iu7moIzG5G+dYQtWAM+v1U21zaKNRDwn9Opi/Jvp1qz1+7+buUWY7Z4iFRai9DtICQ2mS11/
Ba3YKEFvpx4ShUHpiBJEHFKI3Jngl/beZcLjEs5CUKr2sr1yrK0fq7K1zBy/Sfx56vjSl8C2lWvb
85Fgm58siifupVXwx2Fsw2FmJXIc9tMPMwxwNWh8xhK3jrhinUuHOPWMrsnR3LuKpA8ipBHZ0b42
PcvRWggsMO4/pJ+qTlFLXYOkIfZ+tqY3ac+R07c2Nibn+e0uu9alSkOATatHSh+aS+NT+n1AARba
oVaRwY9FonYZlWnoGdL6/Yxq5coXd6QD8aU+yB5qr5KS1Jm4yjNuJ2+wdySd8XgysS10R4p/FL9t
CHlCqk9pkHXDMEVGv2Msn5qsia3PFOyq79Sv7La1ITkXUFaG8T8G6MVKibU4q42lAG3UCeE5A4cn
Cr8xjgIQUmnVyZYM5ru9CYw6crkCXrTSxdv/qO1mBVE8YA2i3KTIhKFe/cnexj+drq4H4LjkPw8M
pfwYmK/T4JksiYpjFnIl0+JNoYLn18rZKJ+B4cwgI+d+R7fpV1V4jBQTqzUVX1+5t+QIrz+mM71X
As8MpaOJ4TgoZpmbsofyIYPXpYYBKC0+vr4GJzczXxbUarwEnTGVvpVJQ6lDqHbursCL9QoyXahG
5cvVfaMNxZMkD7w94NLGG/qJuP3iWgT52YXrL/5Yadu/cDWrXsEDDH6SX0ljj+J8OuARrqJ9+H8g
NF1X9f5jq+ZlodGESWp9/VYCfNpqucdR+3ohak64+jnOtzXrWPTHCgh9xTE8iSNTcDRX3Wees6xV
eOEzGu1j+VCsyqzzCPs2YTpjix9y8Ea2juoWIYyyrKl6TqVnpccJ52mnDMbGo9lJ7EQtJ3O5wfy+
PMU/JW6THDwAAjAMdfzfFJmz/7JTrzdCiuDkhl5dmhvNWKiWUDP0pVvo0WAjYSME1+JpkA4Uw4Hn
syez7Mw6NojvqsxfxtbJyvzwx5u1QOkhHx37MmH5WixYQoztzEp2GiUW11I5mS9K2tfvG8AcHePL
uPgx1FH1uA9HA/5MDk8xi0inKbDjRGp5vLw+Sq++e3m3mYEvhhsNAa6LYKklTyDLD5i5xpKyv0Zr
5xMdVrmKgdd1f995fAHPmuFtZQeaxsQTOK8rRwT4GEgAbiaj37kOoJ6L55bGmhe4KCDETdoZzk75
68jCZv8pAlcgR3vbjMchgT/LSGLOvGHjvwcoDunQhc7u+gTuYxOOUpq8rlWP8sF1sBsCvZhJy23B
Wt++1iDUmdIGILHxcdzzulOCwMu5DjPHpe9Dbr7nrnUj5vm4AANiWfT69TgwIAWEQnsANY9vdRju
RSssloFIrXqGFe6CnUHWENtAgwJ0ET9SI41N/xv4NmXpeYxen6k8Sn9C7GsKWGckGRMWMiJupksc
XLGFIXi7Awry+gJB0dtNM3lkySMVyPiDvaWUQdX3w6T/hi/MXTJ8V+maI74ByBP+tK/EmPGVF4yV
XERbUQLUH9i7eJx++rxY5ohIMq1CWjQCZu486JwCFFNv9BzdV0yoBeflqD+rmhFweauJZ6wYcM1n
oHO5AOgORAnXI3y6vtG0BJXOzPjZj2QOFLijqby4jPluNqVg+VppVaYeCLiLR8OkqO/BRXZSpG27
2CaMm8ld5o1caCQXVQTGulJM3njtjKYsv3LbnILbvaWNo6CGBSOkdDmeUXbqkY5g6U+YSP4bWq2i
TP4WHAz1bn/eYFa507f8mHMGmk+8Uqi9L5g5lczx3e7r2veQxMqgE/bQbdcxnECPFOCLG+nSz+pm
fSbchVp5tDZhBJ6oDXPtjodirr9VwN7Rz0v3TrEDtqlLIDYldr3xAaDXS0M+kqgQrr7IOqBexub5
CH6WDymGQiNRJWlF/r85amL7CRrsEOk0L+FKbm2zPmf1+F7GA8RNg1Kjn5haiWMn1e+DBIFtsXpn
Eyx9faYitnJjmcqc6GIbP4QB7JH6LPA9YiUWpjobHF1Oi4AsWwfi911F7gZ2E4ECBnOE2jiiwQLt
qMJ92YKP9/QQGM1moA6QVkw0PKvJEmaAU1eRuEs7UkTPmWOBgz9qVXvXVCEMjjwo06gKVRspBcUG
f6qgeTp2XqSUM17C2YGZ13sYWKWeGiGuhUXUUaZuCXnKIEJEXt2DtTNrTSj5SJtfK9y1NnKJRT1k
vMLjbfNYEAg1IoLMTv63evSjqRKXYhmVCP9tCyxYVTPbnyHohahdxBF9AkJrdFbuoGwsQJ2kNBzV
l0OOg6b1WlEXabLdN/HYjInAV3pkA9EETw2uQKwCaKjmtDMdVXKNkEz5Hl2aw3AUn4CPSO71XvqK
D/D+CRMJuE+qf+ssRV6VCR/y1AGfJJUeK8NTP6gaylJQIflMojTOtiPnXGh0Ar76TJehqRmi7UPy
BGzA4bU069YEjFNBwK2NWPdXU5rxERVzHWgeGi+YJNMC3lZX/KEX3sWX5lAl4bSakjBiIkO2+fcj
cwH0WUn2RKcG73+cVxrL4ZUGLSvrGnzYWgmDwmMsF7pmXmnEUMVun1sjrcuo0TUllH0L5a3oo+ov
6l6QGAhNdCDSwBFP5JCo0KpZMjdVW6UIrGvVqc89com7xzVYMBWpqvwlTYawNVbLsRqbRqhcmW1n
sbNORSvEEsPbhkCIGnWgU2sfUXXj66bLEda1mSKhSkhhmC3KaH9iscTE7w5774/0A997F2CYar2D
5e4LyLUmMJ5ZasJ/t5glGH6N9YlT/Y3IInun0mIyfiJe94xYABwKUlAdaUQBZxDedQ9MWSF/qK3t
1DilDC7bNXb6R6cw5/nC26sX983saI2zzqtWlV7Zfslg+S2NZHaN+csoAQlFuLyWDZNWepIi7WzW
qgsw1bixIZrKQEXwMN1yvucYxmUtL5bDq9owBqH+79FNNNiw6IZSZfT7AgaPzD7z9ruSLTctCce+
n2B10W+1CltrN0w2Ouw6yARqf1wMNX2XBLOfN2XYq18MEQYWIX1imawiulEV9JRLzC0BeIC5qnwk
5oQO0T0goxm27Qp1BCWeqXTYWXmkxpxPPceToqwaemz79cVhWxw3Cy1l/cT8Wz9yPy39hp5c+zJr
iHhBEdPAN40MhEg4ZFWHGPBMBinMQ7egZ+39BvxM1K+jJPshPtLF4awDgJmxHzuRMRJnXf6dYj3S
tqz0Ip2I4i2YOVd9TX9Xc8fPbwjrW5+aypnZSnK4w6Y79bvykOvVkICzPaJqkH2gzbv1i5gXZ4uf
vwe07L9wCD+4DS6/k+Jz5c6wrk3lZSXdhKnzAQFaKCzVGodIiVScTpyn7l4nX204dv+7ZHJ30M3O
1sqKzA9nTvRxNja3jA44J1ClANsgPTCj2oeot3cEtzGBBkoM91xtPJTweAVNbc4XCR1L4yGzw0d9
wIgPv9YnSJ1Paj8lofwKwNPd9jls2mhpZx2+2tOJ/SqeMd4tH3l+HxK/dx0ELhRLk60K6NnYfcIT
PD8YHBN+AjKS2KFhaBrrnrEVkgLxpPalZ41Om2agJgDrsL/1LpL6iLYTX7UBCmKl0irEwS3olGyQ
UnDQ+CVJQLUtwPFIjbByJEjh26tPEwu38KJ0fPZ85m9JRszuv6V2ijdCDn+BhS6Zw5frEEPXHMyq
sFG4n2izXeOLA7kCOPmfZKZhZi+fAbjRGCTJE1H1abjLdQram3bbRZ6wXm1YM+X96nmIkoLBQAqQ
8zsvhER436QQJX9FCpeviXoTEjr6TdPnkO32HU4gfHVdI/1NaMriylQJSjuva60ba+WJ0tRhVevE
fq25wuIYrX2V8zvmyTXqnsCvqdJYku4x1ZsziL97UVxiQkK5lDDE3v2KwH87q2RSRwX5UKSXhCk+
he7Vbc3f+ou29O8wjnoyvS13x9wLi594hmnn0xQjqU+WcNuw62v3NR1RlGH91sq1m44f9AmfY6Bu
4Yq1KA+3AV+JXsOXpWKtzu1VYg6bR/KU4oIMT/VdZ7NszwIkqz8qeSksN1QS5hWwk35mye3mke6U
mOPDeg1Z79s0N3LqYwgVCwUXBf7JqO7/w6ZC1rwOF38v7yVLuzjpsJ5z9ORCEOajjx6bgLveBigF
WaLRWpEipKIYY/24xX3GqfdVkntj9qgtnq8q+oQ2R+T7VFkJE2KHlYTRBrU8tz0bpjgDN4wLWlHI
58CMuXa/X4Y8+Xa3H5BNLav3jktP1wwV16diAE00rJ4E5lzJsZi6Urv2/Meaw3os+cnMmK2cTrkL
6erc3u55XFRMN3Jucs5bpSk0Cw/AJgrz105SQjXmlHQ02ZyvYzmltOhmlvVKooEnITiRdSKNwiVc
l8twZHzXY5lv8nMuICRqQ+/thpWek54OIzmYuEckOj5X3+HdEDTGRzFGYUoU3A5KUIww65oJk79I
lyeetrgrkDnmkiyR0zXo+DySvRNXqAuRuxo9/AUGLgIGyzF7faEN24yYq5/MO8dyHMWNfFX7exJ0
febNFYiVGBuJWz6VEq/HZvV+TX8G0Zod//TN7sAw5H9MCQmuJJxE9SK0qQubuEIw9tJ+CEsAK8f5
Q+XZ0H9d63krchWh4FhOEU7DrJLzt79v/eIwH5IvdXXqx7LsFYEA+qydQ8aStu8LrZGjfMRquWyS
zzFhANxRvv//TPPjUqWeBLv9BYYSVyRH4IXqb39ACFqZzCmfPoMYvzsHvZOcjammVySOYRZmmw7j
tJY+1YDog2Of71q2XJ5w1QWyQEO3jHgILT2LTs5GGLxm93KovoXbO02jfMyC1UQUYSvlocF5SM2F
oi8Fbc6XmNh0y5oH82KlEzSZISp8ncb59plNxkGyKGV3PxQks+gUZFNWecXCrTlYeXZ+W39u2ox8
eqlr91npVTpcnvsqm5Wct4N1Hxql+x8cxNi7+Gaa3B7Prtenydqu+EzRQu93/3mgrZz7NDC25FFk
MW/X5u4rVxN6pFKku060DN7fKqsdBNE2YWPbV+8ax+kS3h4wzfXp1qAUR1E44aOOTK9/+rLOwyoK
DvjWsLH5ogrrtBMos/dI5VEwd7Fz766flnzVD2apnmU/DLzh3bGqMMvbT8CugJ4HqOFEdOudmWqn
ng/xuvFtt29fE/pVXZcil/fgchmleeWsmwkj67rdPyV/pQ5pwdSnuVTAmGa/TkeD5uo7CERfl2CA
+Zuj9bM1XDiXwnPFFPNFJa1QIwyV4NmPWwpk4p2P2WW5un1QhhzKIaDKFSBjsi/8LzYhVndEF+s0
eS3bA18iGl3HCIaZxHpSlwwZ54txcUq8+H+nhBgZoEpx1HFw312bIWKl6kzbCLnkovMDwET/scKn
O+QdRHNN5T6eAsmvamKenGss7bKzTp79+zA06mPhKTsFx+uK9Rwxi1HTxdkXqnxeW/Kq8z0MkDsn
Lc748pwouemdyANBaRzNIcycbL83lGvwjhEorLv/dFqQgNLAhonx6g4YfNBF3ytgFG4NzFCFkfWe
TyCu6ysE087CGuSkIXJaGAphhROAC/Rii3uT0mUbvcEPXvf4Ju1ZSfpI89sg7SykNTIX452GLzxZ
hS60Vze1DO5FnB9v/JHPu0sbHAq45mdFQjU+YMgFCyKnyLQdlH5ewgMdaNH2VgrsHCO8zTPXbnzc
xE+hYwuqOdCjFymWsYQDB/zZG3PtA/C7PId68nPfpwUy2Q3W+9fEDY/P7aHzTESfPHGqIs3+Lmrv
mBO1TsAEwSMa/qn7vqMupSswsITvn8bRGsOSK0/UyRiUPSc4lR3/4qk5/1eKoABo7lXsNEQY6pVl
JWsi0UXytLB9yoPdY8YYz6LXCVhZ2EnksntwqY5xsU1k9wJgyePx2CP0hEjU/QH2F1aTH65wgGLa
MQ3pOuHB47odJTOcdiItrzxh6jyIFgIIvmXAV8+tCxCv0hNu2NpfrDruqVoH+Zgt2E7uSK0lgziw
WD06nq2l9NKhUIEuL/N50UcDKa0a0dJ767jQsixT9umvpctVcbUXnWSlq2FWKQOL2CjeBBspGpts
hqNtuXQfbYRIY1GjniLtMfcz0Hatb7t1wPtxTIKXplL4N8k233B6LGGkaoE3esVEBdN6WNmr/ktV
Apz6M80oEUhz8YZQAfhiigbgagylbotBlcaS7dqviQJlA1BayX6TXg6fwdgUbDeVX/1YY3cP7UmY
hJoUZUeZ+jvhvVejicm4RKrvknzOn2LWP2W7SpUKLg+R5wEnkHGOB7m14wzsjcQwSbmegnd9QxVD
hX+x1E3pN4D+3P5uFrV1npbvFd+32EU1N+k7RUTon1Vvv0NUk8qBszUEYh6B0xWX/GbRXpGlvGyf
tmEKbsxaIFM3Ek5YlFRtM/rOr20KQET1w3W3pBaWuKJVA94D/w1/bfun2RGY12CgQSvOQHo+fZiI
iPa4wqsgOtxc2NAn0m1XW3WihzjcKjWke2u4ogAwuXyYQBOWJl7qxmO6CVasuTHZrORU3HSOVadi
v1dXI9lffKNOlntzFzr1XadliWlVfyII1+JqnXaGoFbcV1yS+K6YcO3DFBbCsZuB0BdDeEl9s3Oq
UJ4HswELvin3Zcr6OXTsqBpK207FcfZgLtaNVZjPa8U6yFzox4KvWRmfr6fGUTn3ZMX7Agf8Qa1Q
tP4ePtdcemJl2QX6n5x4qR22PNLKwLGTEWLyGwx/qwgka3anjvpoFOf1TDlyISIA9rKqbryZ1+Wh
8ZdoglGqmeS/unTRwb6bG2+M+lROgoba0dFwPMmmoQBCLUKgPBvd7HQS72R3uERf33q3Irm1dHDa
WH0PpF8975J05hsgHDFiaoAHcWWTBw9A2s/SGFOzvdrdDR5kIt1HCePLHEfZPY7WU0yFFjrOEIB3
i6WbbGD3Ypa2URTfblZHLYWkGWJKX6nu43LjrlKPuFBFYzYSJXFv/WqZm5otjjLsfQ0qoYeIgVS7
ze89JHndDSRR+ByzE2Yo//ETBIRQHivBZUr/MPs7aR5+aGxSMOCG9Gg8Tmc1lMYw9CBWMufUp9hF
RwimpAgcjCLuFMe4jujKFXRImSBkJpxwiPQv1IBcBF2J6/Fp/B/E0cQI1aecwPJ14gRltPDSE9vb
rV60TSC2Lu1q9svPkbKAPFUUCaHrg0YmhRO8T6TKPgHKfXSrjJKnWkHflHzcgugJFOKhuTQ8e/+K
4xj3pwCOsI5uUqWSAscsbU+Jc9NMRTDdeIrUqd6UFQjfevXlQwKiKsH8Az+KDSnuuom7qd9dF3XF
HX2SsXXmKA4hFYJPJ1YDt3LUS0m2Eyp0oZWsjDu50zzBVbhMK+mB2W+lPNgfTblz6dgZbQWAXW8P
JadFO4DiycQ60iz7UhgzwEH9A96wE41HfLVtl/95eEeC/TOZGjRdMfLAI0QAtgyFgN5U84xNJtET
Tck6tEa4Uw0HHsGcrbILgI4rpR8pgmzweOznbhgs5mTQ6ENzReWS768Qqm4K0hYYfZVzuUmykF03
+83SrC4dSgWQypCJkFBe3y0NqjImBtxYHNp2y4lsZEFBfZH78hLAPlfRn03sNTdCixDmLPr93lIc
/CawJKVs+rg8UC5XAeJ+0/TCLZlIJ51QINgGHXR2a9ibvgordArPyuUBuIvfEYM4CuIygLryIVEL
1Yro/XNfFQvL5H/Hlgo2TTK+0SXF/uLgGXuNOyM1HOiX34tuB5BowTesaqLiqi9jhgzt4dTMWk/t
kFyuU5nz0XuKlbV+ckFLLrYb0fDXbdKvk0rEdb/PoEPamYuHpivcjlky/nusz10b7L8PyCELetD9
BdzE/Zzq4aIUZNH4znsAYFv1uwxKjiPkJR/4ii3OnR6CbfTbXDgMiWxt9YzL86YEHm/jnQdscinE
VvztbXhb4EoHjrkt9UhQ/vSuwziwLv4Gl/TKWYzlmfVADVn5juhKikmgvOwiIKgUaJfKEAEa4DIh
/DJvEiGd0ogkk/rnKJR9Kckg91NiNAdfAZvG8aC76Ix69G+UnhCPlAiO3L1gLn4mbv3r1ieAHc6i
68XaJaiubI4tCka5WDMfgQlEgOmUNFmSJfknEi7nmneUGDLLTZB3p3auUvh+WGbFmP0mnV7GeUFR
o7yBR104vq0aO1/qyfhW78XIUEsu1DDTC0YfyekkKdmPsN7KwsDEcaIgxlR5/AfrZHJ1tktMb75j
11bpREsWk0sDxkWY0Dc+pOtqGa7pHx9objPsftVgj9xB2/1rQywkRyUtccK5KGBZGXhotTu1spAe
2n2J/c7jurzoFYInCK7M9QC7K05LFCXhBhIXEU3C9+dOLIPPE11Y4fMTKbtRKqmxRE+HRX5fuabj
ZmTInWs+SL21vrJrFji9jQ8lxZuErzuOK6As2GPogF3Y4K78bARc7egLn2TkN5ex3MU2uGjufTAQ
XKNK5dSoQ8YgRW3EW1GWljl9G0wwBrYQaTnfBd4jt7mJ0JHnRFr+WssV/49YSke8SPt+77o7QKQr
n8HuzuBWvrjNj6QxeZsXwEes1jhc9unIJu/55ANbHg7G3jhoLsIp0yxYw/ZWT13F2DN7khkv5vs6
ESCQY7P/Xa84PCiEH0EVNOiVigtYDPwtTFMeJ6dlHlxTn2kTAZdVQtMbqxDyaYCeDYXJ+THQz8wY
58uIvxhXgHtKP+gBQnT9C6m2geC5ZMDt4Nw2A5TY0atkUE9+uBsoQm+KQxkON90JhMTOiCcDSx2b
ADQjRNoH6Awakq4wrtrXsdT9JY11UqRRz2w7Ik0DNTKJ7/L+3jZo8XdNJDAOi3rcw2Fl35OXTBKJ
yZlMnBVaRGu0WfLWGxQUeLul63JFJ6CW3xlkvLLEyTabqOSb6cxnaNx35zK98+7QKuvY5ri+1I8f
vKY184KPtTsshbfAMx+3/RyuUnyWgfjWLu0fZl0J8rjnEkKXLdUD7Mlale+d0rKXm+pkyoz8k4wK
Shjf3g3vd0CWhuDa+Tt/GrvunhSWtuOTuBCubv2aO74dBHDDF5vqFdrQooq9wQ4PpjjmzbUnXZhh
I61qm3gpm0/03o2X3crQuJZCVQZrLRnCOSvK3hylP9GMkGrfDr695stm4/XegsTnqGTfPMWRmXEi
4XZKBeUmsL66WH7oBpfmBuXAejIYuSoKIZ8Bc5WIa5WdGcfNpFW9f/u7yzP/6g1A8lZmWkjU1uRs
LdoENtGCemQHGta8FkQ6R1l4ZceYVkdQOnG9J/2YGXKYaSs6UakKbNsAN5k7ErWMf/JHjGLS2flH
3OrpcXrDC8hX0IMpPvYDxnzbd6m0jxwyLs/rbpsVdZga3sRgCb5kG0pC9bc0xEl0StuK3+pTV8Id
x9PX+4R3alH7Pr9aLIiC9rZqQ0T6LeUQpCIiLQ9IDIrkJ4I+tS521JehxyWgx0iKI57eD4dNSZ0I
gJ+E2TQfBelPxGbuLolhQ7xwwOg8LPd7l1oLYy9T8km+6m+WrnDHZahDz80JkT7MtJcKZ1D9HuIo
CsKTlTFleQaedTlJvT7d1f2jLnUyF2TZDAnpGobKcwMTrg0QgzGqThg0wFYCffvVrfSjaGJiwaf/
FYvGgg9mSXOTTo+jZoPuyc0G9JExU2GzVSmkt/HWM7V8CKsYR7Wz9sETY+2cDVSj6/TcJfBLlDTB
35k1j9bZ6PmPHk2RL0jm91UcLpwgN16A+kjvgwAmH3OHn5tAxE/coWP8RJr0kEb1RaSWsHmytA3I
tM3m7UzRHuS+zWe61P36XTjruzJX5PzFClgJZUXBOQ+/YD+O0sFBNopsWrx+7mzm9LuTeZnmhpJ2
GXKbszmOQ8soTDYNw41rZFW9sXsjraq4osLq8kZTT5otA2VbA2sOaBGle7x4ZThqBPxBvyWaJFON
TcANdTAf6LdXKoYdFNZiEFWaYbhbLScIe9QD013yeGci11cmQWN/KTXJ8wxXM9aTDoOAyo+8bykX
54N7LrkUG2dIlcL+O+E1OLiLpKrzn0LL/URPU6qV7a7m9Kfdngdc+47bRJ+TwHvlburHoA8F4bsR
PjBCsjrnZWCTeTo3di0rKb1jBo/FARih/NNqCaGaB+SEnDfqzty+3Dxse6G7z7gWLsA9HEbk98Kh
oPaVTCnUTtBeSr3T9L1XyF9DMjpRAtQigsDdNRtGrLhcz54hhVaA77HWOnBmxlAelY0HbvvTyPew
quK/P8jbFbx/IZNgjx9ivMKAN5h1adtdcc3mv7hn7cpjx4bR7H+b7T40DFtvzKFNFAu74sfE3LkJ
l0HaIe6JOZGTUnwqU+g4o45fTVQxXgc85zITCstyDeCos2HxE+3NiAGTXFw2AVm1Wqo/HqSt10gp
iZv8F/ZZT2xQx4FuymKrbEfFET7glmtkRhTjnBe7qvz2H1dwQMMG0bdgORvW6halbN+mjneae8np
/euBpYJ6TJDG2V/OMr2neMQ7FWrt89KPuz5CRaJ+MtQe2taIrarSOBAr4eTiASQgFCX8HNl4mTuE
VN/cGSblPjayVr00lCqTlO6FGjRmUQAO4FTOzEAibGd4nX498SV7VJ+d3iN5MIkD+l3I6ActVKOW
csAhFuOT/flLK0s1dnh60X0xj3l+6K7w0uzT4GjATg6sUI/MCdugNO9XW4nIL6sM5Amm4JvXuiVG
Ue0qz73SaW9wN1mr8XBqGq0gN3JU6qG5ZrJwA32SSmzU/IEJS6HpKVnGUSwXnm1H4Lr8wjn6zaWm
bt3HCxdoK+BqrP+V7duQOfOus4ia2P4qOEUbjZVSFD35LsKP7HXgP63+0CITKgqvpxUxSHTWsD1X
VHdvj/pheygABPrne5HqD4pbOYDO5HHWreYfaeVoFs9juTERRafxkBpfUiSTpWawmw6gnCoJPoMz
lkYZgMK+5hvmiingR6cnp3TmZdDPaR/7KFnVTp0wOQmWYnFWJdFbZ+Z7pXpZwuNFDNWTzWeZn28M
6XuOYxNbIH1Wl0kKD53lyJMZ+/rV72wJjwO2+y02XgKYjhvbeDr3CMvNz6cCRc3zYhjvd/H7fLFN
M+gdvlK8A/Efw3gmyYVwvz/GDpbHwA6dzhCdsPRybysVTMuGENqQSORN3Mgiy4elJkzN2vECktnQ
iXrMWKShGGCKyflunL1IerrA2veluUxcwdgkmbGIRQVEdhJifK2RcduNVcD7aFsortE6bYMUIY9T
RxBTXMrlG2NNqs/igCd7HW1f9EydeE5zzDZmcqmSCcJXlmNi+RtKnqvRdQWLn5LpEsUfXeHkAXkH
wze1CoPqnE14FouqIo0zhhCNI52RBSLNuPB5+oYqIF5zL7/+Pc0v40HzK0W2G3/h6h+sK/9KHAYf
B9SMt+sB1efxGpAR2BgBA2o88ZfibyUPtr4Ga8BBBKsHnkqq8JFKMSVFIIQJDrFDyiukM23CAB1X
Hm+7YouPrBnivE3Dph68VRWP+14LDO60yPl13Fmkc7pi28rRXPfHeSsP6JUUShCieuIC9yeW1vKZ
Cm563qEx9rM0WDgHM2CA2FNzJ52DBhcRZaO9bILyYl5YwOWB30Y6TTZEL6kvclMEJdMG6VP96Mc4
SHXRWcdWxDM/MUelNstynz182LCm5VD0iD/hP49zhy0LBIGRr3ePfFFSkclQd/7Z14wpkPmosdzD
xt8X5sS4Gc5tM35bugD6F1Sz7fELHEC+qj0a4wKRtbAD+Lx6r53xsdXKkTU0N2Ygzs7bA6oIl4/z
laNZs0CCiZKhIVx/m8T0lTsQ+fgFdfubdX5meXjdSCvjvwJ24Q6n/Bn7Y7VjCiJHSkdKR/5N8Cok
U5d8+DuyTL+e483qliRCTPcoyNVQxRs1sJl7MD8ddFHS8FQhnbmzzMcXlU/CbqAUrycbOQWJyWxt
AIK/I9vcFl/HN9SRt6lVqtBEFTw299E+b0te+E7tcQ7fI7rfWNeKbTvS3P94LserbP/8WopGCDud
KJd/WaZMvxqXF3/kp3Rx+EeEYoB2/ykGTZ919RbUDie3ACzzLUbRmc1nqypNG/++MdbDCG1rwbvc
dpGDiyp49P93ilj6UgcrQZ0/W0Mwq+yUjgmL7IpaRlZOUj5Eu6Hyycv/OfU08l7iJkUYfnR2MAYp
YE3uZ1vu/aKfpRqDRLAkJHsSZwpFiGvsAvkO9OSG8QGMC+NxPJuBI2eseBsPKyM1VQQOws5OFJD0
1c0mrTAX+Kxdd65M1+0mbOoWgWGzECsRdZWdVptKiA6WRFnvSWLCVykzZmnZAHDWoQcjzFSWcGqK
i+RNsUqj0XGHdCIbYoJL4jPyNNoddCql9KaRjA4kByGUTk6Lgg98aJxY+WLLR1ZHEs6mTNTXoS3z
57eOM7ZJXtPOXfl086hyUzl7y+F7MS9hT7POYiUsKWzafkE4uO9MZbitzp3lDrtJVbQZdYx/WcZx
EnWuLqqxTo6z0qirqxmNIFYegF/Y/QVtuZMMqWXwSZjtc62ptuVmRRWasGBsGu39WGt8aDoWeokJ
MNpHUSlI4L5rTWljOTcD/dpRBbP5ogxBuZx3AYPH9l+kRAn4Qj1HGKshvPcmoaerMmdBAhC7Jx/a
VLgHEI4veimLziSBes4Zx9LG22VvBA6OaARB/l0NkXramV6JLeJH2SVCnMIXHcl/wFF98lLOan9p
u+EcQ/YtkcvG+x32vEIK6bRcISSErZMJ3liuAsY6DGe8glcGky45lf5EERS04pFds+ZoNgp/de1v
Y7N+mzoRCDEnTHNDZxCIGMroqR6Vj3QlgQp+USsbpUPaVcbvQg5ykpEK2oSTmxT8IR07DYuPk9PK
zxJkWKT3wIcXvV8ByCB8K0VQVWUpJSweScCWDvVdSns4k1O1H1eneZ+KOV7sTusEhMvxfS7W4FPe
fJfafEwIUWT9+KekyLsxEmu3x0XnfFC73KIG+PfsPsuIvY+Fvggft5DO4L/CkkEPYEUBnknV3NHR
5gE7dSMvEINWvr/NbQRP1BdMVYDJLiGJyxsX+IonJjwiPVd2Res/PJNzQCxLbHdNmPRGbIcbUuVK
BWB+UUu0WxaAa39uLd9cOVa96exhyA7uceUaya33yFLfYLNUrRXVIZa6+rAdfBTLMh4ZDzZFtpnw
D//q52oV3u7/1CFgJiftH0V4BmNiE8MRXW/BPjMwGoJiOVoZ8Z3/Fk+k20Mf3URdlUXGiDuvMFr9
Id/0wWWCgDhdT5YLclQSNkZp5jVFjhawIVk0k0MGSCyxv7rorY3GwbrMcGPbG8FVNTOH2HBwaj0A
Mv4GB/lxkHe7ZAH4vJ61C+NuW8EOUuMXTyOeS5M3ojDlwwpQLNvhn3+aU0o3bLNmSjsWk17Nr4RS
RI9zfc/X3YMzlgBNMOtofscMdCMiOmWEMxlTlPlqR/S6cdwaj88ynM2Ku/5FO4H/mVmpkG53VHZb
UX0yzg4d3y3YkwVOJ5z8VQFX7uzBWYYOJK51IjwKvg+7aG9UHGhE0JiSQAdHVRI13OHGbkv4GwT+
RCjIzJ6rF3z5xt0MmmDWGoTn1EmxlCZYOGqTAsLgX6bFXK1lxS9B6HvPtHBQZ6xS+8hDnzIHv6Kj
9LMh23/59E37B6L9u1/D41deiuU9PqqIpi0632fnDqN1ziz8eWV876DOn38Xtti4Xft9A9tDExqm
WpiSK8cSgbRgoTgv3hnzLxjxLSkz2xA7hp4vvZTqb1iFmmG1BhRL/DPTcIlYffK3XiqUs22wVDE/
plClYZ5FZeqKVB8wJW03CSGkyOSBB39wmdfb9Kqau6Vfu3IEm2bsDwvD98MG4euX7k3miPfdjq+X
CabgA0JMsSG9MWRHBvbgPgydmRAl6galkhS3EUijg5mLFOHyZ/yCJgdaFEZQJvzoxGhSyh6EhFwo
Ipn4h1AZH2UaLyIOSIt+1BafPrQ3eKT+Mrt5Z+syFE2FJd9vBPZl5BAdNq1lAb17+wj9z+ks4YvE
rRW+DxqyCYBGJINGjzMslJz0ri6+IA79DaEJnKCadQv/81945okoP+pmiCW3Nqi4lyPrLdyWz7Fk
0abGeyGc4iBPGmtyrPNcAh504RG4BZfJWsv+3bSJKHP1OrWzHdkwSZEcHhlvAHp2zcp6myJUElhj
7sR2Z8V07m+UL4HYSR18gGOBjWDLYfvC038B5qEhIQZUTaoAs+1d9khd+CAQkRaKpLsnId/w+7xX
2vBhhutV1jiDBJjDhdRgA/1j3r9F0+MMIGnLiw7LWPvCQ9Z+VE4vWHSKcXYPMpIO/9lR1GorzDDH
I63XCxlMKp17TVMn9nJMgJz7EwumQuQBb6GSw1KiE4/KONsZ//JAmmOy9j2f306zgiteex6Of2HG
bXmtId8VRl8iV5vTi5f3VFzNjp1lI/H2Onh5UzDuomwChF15TVvDWyiO9FbfJz5OoQB1oMJayUj4
VwwM3mN9xqzVISVRmTWhfsF2m/3eurut5b9dBO8nX+mSoDWWdN+IOhhgqKKpFEPAUp1VfMJM9hzy
RkLQK5T5/PNpgqQRP7hO8J86cjmxYDzUcTAe8A3/3pgAcpJEZgCiQvYdG7UfNXxLQ97t0w76PcQB
Sl+srYK8kOqpmokI+MzSINe4FBhOsmH8IXk3YBtjBzrnejTzmNJFLZviEd0L0Bb6B6RaB3DWYNnN
JXcZ7wCzcnWnmQ7wXxxvK4gkuDTac7nGFeM+DGreWVEnh4OIAL/0+6KUKV/iEyturIXiu9ioYHP8
BNgSQEQ3f226P4sNB4Jb72VnLzUAkXraqlxPGxpyrBf9A8Jj+FwajDYxXeehcvWTmhvzyUW8xfSS
E9GE7nWmznZ+2qjm/GV48c2cUcJI3QI0V/ecgPySvebBK108c9GUA9lNW04YBPipA4mGZCe4G+Z2
JA0099cjshEjf9QYLlHKXRam8VEMnkDXBZPlIAQo9Q2LfzjKkxbEGC8gMhYK5K4U0ZhcuXm0sNqb
5t1w+JLaYM+x5q+Zu9W3Or1Jgp399nx/wz6owtAStbi3kLwkr0DMkTx5D4edRM3Bsv5cT/2pVPON
FYFST33q0o5YtTJvUoXn9dWHWzs+UUmy+FSa2uN4A3hcxknuVjjQLFW5GIw/HyUs8P+EhbE9jsSc
wZ6Nn8L3NjeU0AJMagbOjUx1meK5eCZFLKJN5NnKg8Yn6UHWsdPaEJYzDfF6Gagi4qSJmWs07c4K
t9HBwulBjMlSugj/TtxRIDDWtPhC1oP32QCkw/YX/Rbh5NubHacBGGDhA1RzMZ5NVJZU/uiI6d/Z
Np2MmH+awM1B+M0hjN9wSeg/L3LxGbM6nPko/gEQL7G9Ufpw1ROcG6Fk/kBFRozmMGXy2TMiJZaf
+FDg4jMgRJIG3+OZ1P2/2eB/dakaKRDu3iPPJuEsvcqM/zm3gSW7YNDSjucuMB6U7ocZ2jSZs+ny
r0sLIEdwT62pY0Vo+cqk/ed26g28yk1vlNIrqmKLbDIPKu2fXCjXEMykuDPWghqijVzTntFLfmI0
HDfyDJEy6AIz0J2f6XHrYK/yg13onWIgfE3gzx56Ru051iSLxymyEcFwPne9inSXzslm58u47vLH
NQNekbY9KnJnU+PIZExIVdsY6gxxH8rEx3e+WCtTTkUR/czT7I3hBvEMZabttyrF00emFj6zkA6G
2UKnYSEpBR3uiCEnwWKDcIxnJRBG9SdejoGVA1uLN1bhiBpt4bINlHw+MJkXlGIoL2SvPqxf4mkZ
m1lPrF/TKY5pqRHNw/jvdvOMqLntbKL3vdIUloop3lwR7VFjhBdHE4ES3cEXUSnrdQmm7b8ETDh6
2WJjkGPxqJKsy310i2BoAd6c311mldReeTUjeUIwSYDZrbh8Wu15nH2UemwYj9ypouzjwve6pYib
LzGW1Nh9lLcAkRmiAhcVHlOs0FUO6tK8l2zk0m5rP8nqTBdNFBLpNAwmLtkObLpgW1ahndU+561C
C4mkYM9wtF3LsaoFM4+ouSUSUsIo0IaL6YmfbrlBuKc6dM4oBGLJguRAfCrEs5xiPBKxGSiLtLpz
ta4zIb6DIJD7eN1EKMrJekF9pENWsA0r2ldSiuVlZRQY7E1RiMcJ+TThPHHZjbuYKBb+fIp5J2yc
L1Dd9mZM3IAUwsHOS6KRv900esExFLjTAacmQ9TMdskhGZWhoGMC/eE0uSCE5HlzyOgMdIviT4og
tyz8IW5bsd5JfaRLMibKK0KRqYPsxXYdaR/O1LO3Mv1REHNsjlNY3uRp7z79VnE05CcE6pt8Uurz
YbUQs+qKiRjOUZvFNEVM1aV8Vb+Wosa7b479V5RAjwMbTMXM9iFhTH4ID0dblIzsuWIl4oFsMA8I
pJm/0X/UA7AhAS3KmCLR0+EgXemWru7E2yoti4ut8Q8YU+0PeiN4Yr6ZunvX8+aHUv+Ngk6E8XzA
gRQai6U+Qd3hCvetc1hha4mcez5Op61NaIAV9IV1RfztCLcyKeqgC5y72I4KSfIfLKsm/RamByub
rGn6VW3G5iO7UrieeBYHfhB8ySU0qIzl94FDn3uMyN0J26eMX3sneQnb5k/AfYwxNRLYqzdUILyB
gVhGyBck28G1gDycw4e8p3Nsi29EDgIA71o+SMvjv4z23ufd7vcOBCwUK9IFY6jo4o0iN2pWEWRh
XpqqGWimZBaWI1KkmF9cIznBHBMLoSipfwJLTC94NQwxhHKzYIGZKcVYUKBokBtwVPn8e6R1tJq+
CvwrFbq4rGzfnss2dCau7au6ZoprXnGNmY2/alAdEnKOYFHwlN7psxsPhKTyRXC/rhhb/nPjZAv6
HTd/0puyyjGVk0m0Ju5cZ//FjXzMZ1kX0JV/3KxJz/y+gkuE99oE3WtZY84PgzWahKr5bPbtC774
iGuJnc33CQdJHGCKLh+Fu9jNy09DJnmONZMcvm1PICChA5bIYLAjFNIBFAwuaF5ZsAxeZt8082ol
cTgNVLe4IQMwSB/tHamjD//QF3L9eYbHd8u8dDZoCcctEpW/AVmosaAWeEsDaC+YbUgiGRglX+Ae
mhuNSjFBBz8nGI/o80Fn7wXqyqLg+K9YyYJ0qCBTH7PWQ+ZHWuuw86Ko9BMlNhb1ArucjkcuBDm3
MJNx1s6Yie8x3GGsemAW+jtyO/T6aOFpNqekKljzqYMYBVGVLOB0H8tsb/lLMv0tuYXm0LCMHdtB
73YZsCLXoZREs+zMmdc6+Nrn7sXX4mvcxIr6SGDydWZxhsW5GWvUmAD9U3W/9rdVztfu1eTDULhl
31zRWP2ioKbYGDTt1NrvX7uSZg1attDUWSOk/jhAq7zlxoDqiz7nq6ASwlgfZHZ6MB9zu6R59/tW
xvoFpDcSLHWUD9rp9VLx4iSreDOy031pgPGu4ID15UrglUXl3imNwTiVvGDEAZHMWtYtX9iQ6dSU
OST8JZHlJfCgsMJuUAJUOixN/nqARzszLX83HbXPAmDoyXMjakKFNsUs88afGVh6lNQIzjyc2Npr
nYWziVOpHIq8SFb7ErO05RdsGS+IsouzDifbhjHnzgzcbQ2LYU8PlPXW/fqBZrfYvYn7/uBhA4j3
WkWmog/N9pPIYGG08QUs5zMkyGGg6Goh6GDENqEOUNIRKinZLg+oHYWoI8waCW487cbn2URPYjfA
aPM535FnYATizsjDcxRcIoj1tLuWJUUAiXmKK8648Wkq1djStae5Ke7ZekdmwZbScLQaJo9DnIyv
8Hpm09op5DGzEU30b7jDxLiu1RfjytBkG7gyPO4Lvp3+GytpWVOtJ3NuZJ2lwN0qudcPp4Jt3aF4
730jssmdFtg3nUbzvtBI1JRFaMhqoXM7J+/GZritG0/3FxH1KFPTyBy0BTX4ZBPih/ghyHvUNEFF
DCmYqtw0T3dGSCyVoPkshlB546GJ1d4OLFVQnRJaaDe88UN/qTPfj4DiL8TXNMhFmI/P/LegQwLC
eEhETctwfTZ8YO3RCtsOxd5R71JML4nvN39Fi1RP/oer8bo2d/rSIQTXobm3tPhNHw+trp+UpYY4
gwOtjehexdM85+8V62tdtcEC8IPPM55NpoM3jkDdfxpIQuipWCPue0arsYU/N7iE9wPie7zNOMKu
lY1ZXpkIXfGJenE0c1gj+uQo0ybSl6Co2/GcM/BJo2wDU+xWMHnPZ9st2Xb8+XRU6GA0W0ioEmtA
NJy8YB9orTV1e4qUhVGeAHePBy0ZvYodZxdHkznSOlfjQTstMGolwRZHaUimaaJO/fRcJ3xkGnT9
L6pwwzNVt9lHUYNKK28V7T7qNvDu6hACSa1yTjwz3AL2p1HDwuN+bHUOCYgS8soM/v+RFaVyUoTq
9I+K+RC8aSqCE+5Lzz/Gr1SjsGJ1dv5x/YZdY18Oa1ygviZrfjmsXTsUE1uxFNILVH6VMrApHSB8
oTlYGkNT9UYNUKBuO045riXRmBXX0ftv5fv70/5q9hra/ppcxeF7V7gNbIoComf9ZBRDazrgUrkd
A5UjMSkYpz6sVEHXRGbOVc21BEopFH0L8GZGjnCmmP7+ItThW5OmPweTVioPE2Tg9vHWrc6P1jyB
nJiOqu8JIjnkRiWuxE9VX5lyM/kMPu2HPiNiNPPuvXPLoCgAgmi6Pd1lL0KIw63EsPeCZwy7Avsc
r1LcoziRueUnkglsXHQxXMAoPMGXubFczhVYLk2b0BxC2+EO7UeWBcS1LDlzDNOcO8rTRHnTnyL3
3WsYwsy08ppC0qJgDxIsdEsinng3WWTM1m82mxEqnadG8QqBp/k5u4fB9WEqk1BPN7SmTPgP+WBX
3IYqIPgvQW+6DBfJv8HeZjiwe9Y83IZz64nlSXxk47rYFGCQemfi/2skmvmDBKNkoZFwwVfiyrS6
BnjEH9VO4BfKXvGe05OGHE0mzI07+0Ibi6hmdm0ouDmgpCUy7YRRVzjESlLcE7JDwtlZjeZRZaHf
pv2fs5fiGwrn1NdXXGXLoVi0L+PVTvwOKOy9ejoTanp+b1Y+W6iJwKVp12crUpi8EPgQADM8UgCv
saaJSa0bUwleIdO9kuk0XOWKzk9MSR60YlR0Q9sTlW9sjvnL0Ivh3eQrUL2UZg4qIknipNFIFFYt
Jeq4rtaiaVq+hl+tgLU1qm2WFLRJzhJatsaAimXS++953zsuRr4H3owTP0Xa01xBN7lZ/8Z6ijCt
a3LR3EZ4p5EDchCrYk2N8k/x1qiHHjUtncVLR93TGzb26c5XRIPAM/Q4GZKdrK+Sm7JU19QjLt4/
M7eWJ8fEcuMhTMnqayZKZJZrxzDbbF/jACwa8qBXZzQGebKOTU/VvDxZi5jwzn3eiL0nPuegiag4
CO++8p38rjDVEN/V3hGvaG11giTlu9DsfCjCAPxlNYlUMvywWUxvXxFCZfjnh8mSmhal9p4miTvP
w5itXo8qrqgfjeTCkllAhXVbqhp4rdMMIUDHJ2ttOD46c7FoAOJ533u2StpBOXW/NQsn3QHI+7+6
sLsVMbKx+8fySJk1PWBpPjgF/ApxMA/v4Pj5bj2Isxo2OHC0jKwxKvRNbp/C2hORopCBrgphEvhO
oc3qxhCgZyot9tabXR9xZVlvFZppLK1yrKl++SEcaB59A3nbjbY3g48yVDp0y0+MrmabucT98bw3
q2S0fBSyf+ipIvehUw6F1t9ca8p+u9I13YxYCxmvGubAT1otMyWWcToyQbG2rFJCRJkoBUKVSiEe
dEpZe2sh9/SoU43hJc4I8we5MXi1cdv2QeWiNeNfpkLqrH/zrrdNDl5MHXcY0wnUQyaFIekBE4cp
hDP1EyQEmj430p/L1aEAIrIu4n4ACWaWpTRkOA5Y0Hqblrn01KmP4KcHgOBtKh6fWX/p/XqePeaC
f7CIztGLiYsnz05i6kmt5qsDYAdXy/b2yOZ+py0yKcmKziFrkpljHyo9GDPmeRTkuG6txZU4byK4
Ch84UcuCaPtmn0Bwh62iV3nrxQ1T4IJALSVe0JrDZdEzCDCpghqEeHWUl4+Xsa2JXfJY8/sff/gx
UtjYlpJWe3iub80Iinq6DHS5VEAC5xwrE4DXtt9ZFQ6ZTW8kfxXop+SfhhjspLoDCu8gyGKvPLUS
mKbhGhQgJuJN482NpAj+41iK2YPJFvqoNrI++S165Ft1bL7xzp3FS7ap0QEd4Icq6GN48moNqGb5
AYAL5gtiedYDlf6RllQCOdy0yqOH/1SShNlvoiamuUxqQLsbGyoiOjcLpb5QcfyiaX8pnmJjkPwB
GJEEDw7sO3uigvg0t5eb4kMxfE/THP5U/XDcd20O/U//PEnsHh//QGKw+aDygpF4XbbFgQ+Zo17P
dnsLauP8J3i8kOMLSEoqslJ/AkpScEQXdloK5D6gt0bPooE9XQrrd7gAfrdx2Zh2WL97j0SOiqYU
iCQ25fEdjSr+lewvNfztYQSSBgX302sKR+f85/HULHe4ecmgfKQjVZqMOpVAbTgwVs33vU98efL8
itmtAhb8D7S78nL5uYLZRzKPEw1It3sO1ENTjDiNfxaq0Baq9cR1ypAZl9nzPcI6cTv6Ec3k5JST
uJEsJKT3EQVW7KHucLBMuEtzF2boQXb5ScdVQXFbuQNanKOxGAv3SkjwcSdAYKv3s0zJUI7/yfFV
/N3czZ1l+tBkU+PxfyRYTE9w8zktPfjqeIBVc4DYD6GSLzlRCZrk8ZWyjkkFClv74IW19ANujRj0
amQE069yP8xdIlYnQ1b9jDt0gR/uwH6x+VD/JMfRnL9i8ERjrLmKhAeOzINwhvPM0vvfgIBAQQIc
UlCJ3+7+tb9XCbcZgYTVzXnF8GBptSQ+dVdUWS2EixMlqLCtokTko4UJz2+QlpJwsV6SpwOVRBn5
Lo7N8bM0NOKYr9bJZ0ngdf0EcLg+F0w8M1AFjAX3uFrpOR2eua8VVDj2Me+KtKA1P9Ncwpp7QE6p
pa9jrXqwmljMUQkUSVkgZOUWJHJjibIHRUUfrBKibT1GIQU4AfUGGK5pFDB+QfFPrRPVc4lonNro
HU23eBBaJMfY0j1REDzmqQoZDwkV8TJUpBs1KGHwWGqtsN2lM2CUCdsJXviBXxdI8HLscKoolDi9
gEfvtnmZR9JV1zn+AQMfcgson/FHvbx5muOIlg3XrlcCuZtLjfRNrMtkvfBxC4aQFALVNlpqU7NW
0SfZ3todbETdo+eESpNgaluqSpXA49OIaDml9X43KQmjaKHYlEDQpHJJxeRC87DVDtqqPG6mPGlU
76+xhkfM55w0BQzh53r1VNSRj9qMfsXCwsR1EYGZFpyoyUl0bCKJZguVngc1PMuA2TjqySJXikbK
2DCIl3744Iv0/q3sltj/FUennXaS//wGEkmQ5nAvcOQPK8qGe2+qArCRjLn/wWbizNYWECc+hAjI
9IK9IpGb7+7zcjPhC3mVsUhJUzFscquhdSXsxcqmjvZ6aUMt3/NCUoWB1j9lqrPq7TfH9bxJUW8j
Jj65NrIeSkRwEN99v2iDDeu/BhuvDrDxEWANrB072Rj4GeNEjWiS/CNdAvzjDaUx8LZnzJvvT8Db
NzU7d2CcEQIo8bvU+BPvNQqCKNHqnDV2MT83JD4uI+OHnrzDFC7fku7DCy0rArlzqzt+KysGFXZo
uM+AVm9T99Ok+6S2PlbQRsGoWsblo3ppwvP33xiLbfzi2vfpoNxwAgE13xWpSWR3DHpWqGsqBrNk
8B5Xi7Z/GS0MbPJV0mGqiuemWbbz0msqx8W3RMY3XMVCfLpGtgTb8uWX9wumJRSH2dub8H/RZK90
/a2RleDhV7s5EPN9Q8mDlypiY260ULGMr46Ke4p4WbMPrXE+1NTDOSzUIG/SMxD6sbOaFV4yNQcw
ycslFx0SUiI4DMRfArcm0OalmH51Bmgl6HLBbvcVrloNKHxuVFdOLzdzbBX7T/WmZ62rt8+7r/Nb
WqaVWgjmd+Z429jQREwg9q8xgGXT8qZMb16m3sET1fonR1KOmkzzgH48xLHFoliiOImamfAoF7Ft
k1SF68bDGBmUlpP8yFDnPQg8EWFXHQ8n3mLICbj6iFF+8VLa9odQuuX75pan7lL3i8O0DB1nu/nM
uDgBx9XMWnQ5FwIaOqnKBusdcGw33DwObbmjwNDaEtIFZDbuzZuCQrlhc9F1Zow+Wyl8eX/LPDb3
jI8mgh4OTMs5EfgLc8N8xkvQ/R5M0CUK5xPkOQ2DBqK8LCq/uucSwZzNlkTg8qcC3QRZY9QWdjum
V4B58augeSy+7Zg2VR4SdUTwSAuQXNOz67JYt946Wdj0s05fFAWSy4TbBgzt9C0czBbjvEo/12US
Iz5MDFzRaKxS6sBwzH+uXUeRYq3k4dfvydiNj8sOnMH0EVg7h2efB5TWmlVUZAZP1bQJBzr72JfH
otD5FZjzlglzVSvvr2ojmfODW1w/0vREdYDrK544NNs5Xqas8VGxAvX+A1LJ0eF+V34hhweO+z7T
UmtUmD3kck+YZw/R5srY5JDKTOW90pk9BM070Xi4wxYaFmyVxT4QVkJwoMooHm+HlFnqHjWYYf4V
La/7/0kJlyBII1L00LzE6azwfoZ+xKY/9UY6ExOXtv+iUwalqxEjiTYNL4AlxAGDLhGgDkSRkGFL
9aAQr38CyZYmmVMJ2I8+R8i4frfaexUS6dh5+qyytjmQbgZpn6Ez6pNCvv3aRkLxpxLcPizwDAnU
4PW8M/X5NK5govXrSFKlv1Wl7ZPBALDU8pIrbEUj7/qpHYQ8CUdU7u1Wno+DVGDRzw3U9wl674sl
fIYPpCEBubSdz7XgqoQZyEHu+olJTHLAaTdh5wZsZXwQlKNsEoMhlhWEOu9Ngv7G5WGdHPt9bkYy
QjAQMs0Yi5epDzTtNx5uvE1/flCwYnbrXypzCZC4vUUC6kWOTVc+kn4O0CWRD8LPfuLT+6nJ+2CS
kaRHcHnJ+PZ3UzkCvl+OYRPcN2WjujmFUNXKXQ1hiIyt9cJnk4GW9Oax3LDEVbcGt2FH+jNh3Den
xcerNyKyVXxDISvWaWILAAGB+cW7gFpWIqFpUw0RdjMTUAPCGNfrJrKZSJODxJIE1Vxl7pJAu3m0
B0K0HzlvgFwLpZsdo6afg9IhbSWpa3a7uj3ZSWCArLaKEkp6dR/Qg3ZYlQZ7aofKKe25oZ0qmfSV
QHsANPK8LaaSHSffVIPRZw56paTSxGk7IwZaIyg2KRDNYKBkVARDXL7L7YXTODL5NTO2tz4/ridl
SwQBbEKwyU+6rg0J4PxqAaUOiFCWAWQLy0mankwqSAZHY7XALZCG3wuDbHzM9BON51oFegyawbu0
hKpZ0VFO3UBA8rL5Mq2nL7SbhU+cDqrxMSOTKzSaUD8XpEXMSRmOyHYDDJ2LdAhOtE5/npj3KMI1
EfaczV7DQSQrMzm8f9IhZlMqat4xGs4Ytepgl7Vvbd0kQTLjBn73npAmP7GAusxNgLyyh5kank3U
x95nwX/UM/dNABNj/YN/Z+3SYBfzDZEc9BXV/BqrSWkqYCpmY2WZlUdja3NukYn6vQsLnhlBShDa
Bu3w/IDHjxnY4STBIk3L3nEx2gCeSIDag85JfwEj386tLI+QJ613msw6ns27jOkRWG8sPtU5TIIL
YaAzolrBfclk+vzU/7bLFEFxPUX8BVLhHDHLHDSXYQFb2qzfWNEu7C9FMOblhX6a2qvKedBYd4zf
2sFHDwLgz04LqZbC8AFa2p81NOPTkXTyES1zyxFLLtA0Kj0FprDI052CkhYDnW3d3vDIG1EGhMqo
GMWg6qBZBT6yqOLGzSYLtUwOiqGxB+05IfljPdx3fSBNsJBCwFGS10WRJQiaNqXexwYg+MX9Mcny
4ZE26MteFdRZCZ+cAzOGD4S6LU3aYKuN4LhnPdZAtWbHxVy6aD9FBNDd94DXvsQ1sj1XpWJ40Z4L
pM/488aX7MRwn5GZZxs7gIicKhwq+N++U1ymCdNg+ESAID4GlBvcPZN1umVYxE1Eq8B/ploGGRzN
npHhy+TYXNE7nweUmt3T5w9qkjONrwi0Z4iiFZU1FF5rEJ9kBCAj2j4CjNE4qcvvTch9TGh83LxB
iJTKMdWmPSmhKZvIHYH63106KFFVMk0jYF89dL6gY0F+njIJXwn4l8EoPNi6oXhlD1mSTZsIFqRs
ntrS3e+v2FP9zYV+3LGikvy6GYw1UYIx1C74hOAzXoD3v7PNYuLwjl69yOtG3VOZ+myzgxNrlykN
IuWVAxLWKswtZ/pFRDflajKtDuOEqdMJYZOZAcTDbuhKcx9//ito9FbD8NPkiaI2q88GlL/Mi72w
y/ZrkGLIS/8jY/8UWGltZNL0+EyBbKWstA8s6zNvFMlyaVYocvikWGXpq4wJ04X41/dR7xSOc5po
c8N/D71GU1BNP4/eAUgyxfyIv74zYR02EtMIoLW3cHBfLEAN/KPE/ECVGrEScl/KNZu649E1b4MI
3bZUY/mb/sghheOw6r62y0al1azavL2ZJRMSzXYq6LngdOHtvTcJ9nRY+qWEFW/btFIoreeEbspl
DTtne1rCbluJU7jlXyNIfxq94tJgQFxbWMrzdTvvypqQ4guz9wYlTwt8Cu1FfceBN17LBp3UxoPT
rJhqDZ3wOgNX4Ket8OaXOO0+9AXPDUpdMZQz9I5fVxN29Cw/zfqTogR2xL60zOJmb72fi8Mxv/Bj
dLqLKWSBDJYZVdq5GzsWWTyjJhT7lKvzUxyOLBK9F15X/U9NrQxI/wq5VLs7SDpnN+F2RuojFVlL
JdQU1n4XaL9X2QaH6H8yBkgJ08IJBpVyP8fwA/spBBxPpb7VYSH0kRBbOIDrwBnist7xWVKaDsFX
tB291PB6fR031zOXg6ldM7vdRdfEL4zKVIupamRKshZF+oZY4Unew+qCLG0XXnOO+VqWkcgd27FW
x3mcyEa/AFnW2XTTyU1KXYHkw+JsPSohHLXJEk5CGSrTgHm3kwqyH3ZVH+QbOWnvH+6wnkwuiis6
TgA7rjMcxb7XF7YG7VSyqFGleZaQa4T1US8rQDAXgta8X58iUC6kPwQ7PFer1tFh0K2Ah/inWTkc
gdK2Q3W7DJLdLI/pUd3vFwbjLTo9HJ9shfRyeQs/jC+V6KrwUb552nyoYPTBIBoD7RmnfTmcIVQg
BtNbq1svtqG5BoNspqe+2272Lp+PIUauVHc/zITqLvGKrfaNNjtIgkn7gNkq/F7YTo7jmhrr3Ap4
yEbD7PLXIAJkdK8CHO5fXMhIPkx866R7ZTZV51EF0U3gI3oYB2iY+cLRF/xYAazyKv2sB03yTPMQ
ul6CVAl3MTUTFRrUji6pl2vZ1UIURKgapxNqpBiITmdudFeiM1NcACQk10/OUjg0R7Zt4LD/k7er
OHn6mvRO1hTokHwYkXPTJlrsSIQ6ks1dIkGyz4l9IB2V2k73vHEsZXCha0T2U4daIWr56Jjzh0RX
qQAKzmdjX7Nt7Vrc0tdWKNBPXIzFfcF2T9eVS2rqGBOAxUmvuP1ieptkecr9Z6IKzd4hS+endVOb
Am3jtGtZnHhfu7coJ7dpKyEXLIYGDA+KGLd3UlM7DUw8F2FZAHlD7Q97t11Mys0V2L72b0kfzfu1
3AKMaJIPXO+UgBZJqWk7sDPsEJ/ZjYwUzHlh9yAjWFQ8BsLWP1BcAetX8td81gfP9vojn6GOtkdl
Ze6fwsmdyMNx34T+eIiWUCS4g1FM3kGQF4bFNaspcrdeI0fxR7CvHp5cAjWLv8NN5sOHA2a1ohFg
stQQBqN5Hh32nVlecTZPe8aIhxkfcZUviIiKFheDBZVK+X+EKTUflO2d58UKwY46O4bxVsU9KB+R
0GU204iSaazyfAOoc3U4mijVOzURQMJTfoAE8jz3/i1Bi5HEAIQLeKZZZHyyotJN0i8XNlMUdcVn
3UsTJeezAeAiTz9UfDvtvM5mHEJr+nmvTN0fDPz/Iz/h+ArACFzzxVQuofUYuiNdADzth5LTMq7O
r/vI3m1mg/xJSBVf1PaTm0Lv+9H4misClDWVQl916geqRqDUY5Mxx13reQsbWpZZl/lhWF7eVR6n
rRRHFu7T4ivXSHj8wYt0xLWJH5GZF+tIbwxcQ06tt8qHZUmF6Z/aT2OB9ijqgAngOEq/u+Vyv6oc
J74hEx0wC4ahHde33CSDbjrGnjBnF57vpcBqMB7eJuXcCmdCNLzTFRVtniIZkGMj0IQuW+TmIoEC
Y+z4CqqzmVZzPANq/Jxvx5LUKpHrFp/KGL2YPJT9eIrfvmus6WN7EofH0xNhYxleKB3gf1tQsY43
KV3gGyPuHMdRQkXACpAJ05ro2N2MLuolz672QaDwijVhh7aKFHg1BqhLN2Q11ubtta33GpIP0TfC
h99HsdjCWvHgTv23f9InUMY9w30CbRbFnSSYpZM/k2fx88ThXiIe7h16PNjg/x9LzYM2mhK2GsHL
D3y6zuAhyRngGUIqjgfbnbqxXeVaBk56CmKYjvs0ip0KZLz3Mfijhl1OWWCVDh0tJPZASFR4xoqm
cZt3mz1z2qz9yxlaMvNuhV0LYx0qIB29BkIdl2vl5tfxHfWcPCLc1XnPAgoB6763mperBYN4xANT
GFBDlZyk4HN7sLhRJnh5R8WkP8hGQZaCb+h7rjl/bwuM0WOlDJVuIwnNKHgJxNdGnL5onv/BKQf4
LpI8twYIHoE0/nYR05yNAen0EHaIV2y1FgyGKhBgCVHXlzovGjDU5N5hAI6Z76oK3lCOUhWoP3A7
ovQnmJcmSv7582JqhNOnVv0mzsYFr01KypDT2b4LWMO8K1y++pTdfUWtzwZw9YCpa8Xy1kvbmcSf
lZsFVFBWhicjUSZP5LDm/5+lGDe2StiI6F0zGnz461Oj0k/LpnMa+QlNZ8MdBIWi4KJnIO9C7+NG
MJR0ulL4/OLE/HhuPIjto5s8rPpO2ejsn35bHtHkOMUnIxuAnw2YbelyADTEELLW4hUV3K6cCG/N
wicmi5RnbBiF/QMdDy0zDzObordGFQlvPqdaaXULTCXKcxOy+6Tm4MOM4dYrMSNnl+iBaYQTQ6Rc
44m7ApJTRdTp+2l4FZ3Lfj2ho+ju9u8EmtFd49CyRnq8rrUvunWZLYVJvyQuI2HZa+Z3IMfxEXke
RXmK4NUbNHMRTDBzmbPq8cvNzcIrLIxpBiILitqmWVUtPo5gXPTFqtH+jVnxX9X9/EOMrJNcXyHs
lPhxvBzSXg3asWOC7+vhN+OkAfN1CF8jqZO4UHL2EZi0/ACbr0aX7jzLYZ6pO36RtOYWI59497Gd
VwszD40iJevWT1tcqDMYf8UWmYcNgR56jKdwwmPscIec4bFbCXi9bOCgA+7gdwxBfJf2xzxSin2Y
vnYqoxUjDle3/Z1LQE7Yn720TrZ5xqo1FC8MwgYX4rHnvM5AzTWQwqKngkKHSXMcNpkxFZO+0mLU
gAG8M2fSK5faIPQUkLqfZQyWV2XDcKRP6mDEFQv0dmJe5UDEI1SvGGwHbt8W/CVcnlklGK0Q8IQl
47y1jcixWa3PAU3mrWp/oNLjG+sFSZrow+d9XK2fmwCoMYo5fb16QB3KM+5TKa4D8x6iX0KT26NV
zvvQUEtiDyb4Jms3F87NKp9IslIufPr3vNmFOx3nVn32uEBUAl0p9Z16OKLtp6OzdpzdLRzN0N71
LjuqNRPt4JsMylg5dX/gdoPd78S8Rrk9mTmtTDn+x8Miw8HHDwVBIo/VzdQnSk2k0iyJQBmLcUcQ
Ei5oEC3VkMCeqr1qGkXSGQn3CMa7f58aAQ81djIaD5vyRaI9VsO32h4S/mLaDlubg1m0yPc5SZqd
YOc9+pveb+D9v1FHATDtu8C93USvs8SZfEsBZDhFg9J/amyyPk0EbZ7RNdYl1a44yT8ZwVWg/Qe6
Uv9wwhK4+YSh7iNANPH88w8zbDaaWm31whmpknk2OHdy0HeYKXQ7QZ4kz60Dm5U6uJNaEYTe8Cz7
B8S6IGOiB/m0EV++42vQ8rTOLodHuHopoIOBE0J0Kitk9wrecUdTaY+wGg71fZwOwG62FN3LerFY
J4XZOdvWmY0Nqkt5oyniTkfSIZxeDm+ZJ4r7bgGwAHFcsMBXLoRdapqKqVWgr6hkE0kuv9OTsnTD
9IQZ8kfnv9QYxoK0o8pAgnDl6M9brlGZ4IOSZFZMjw7HTfZRICAIMac+S9Or5ysGZ83WenFxVNaH
VNnTfkNXA4dPNf+5vArxAhPXiq1oBJOuLzU4lgg7YdAntoZmYkW3rpTTmnTbP4TeJxfGJwhbeJmn
+ZFrS24HkLAaYRzGGpv07ro9tr+/wMnFp+lqjXOQBwbw+nq4layoNh2W3454eKyyKq5eW9JGzkxI
E8CtDa91yERJkrGuxJQEnLbWM0coS4oi3IW5Sp7Iihemk9c2PcPBOIUA4mobQwnpEUb7LWSa0N3V
OT9o34WRjtjUF0Q8q/wjp2s7ku34Jh2fCyoe85duo0xxH21nS3r5Q2cNa1MjT9krjtYH1CBg8kr2
6RmCIz7tihVm4k1cSp0/tCzn4JDYnjghtfpPaJ6MvAyZ0iMc33uwy3aw+edQuTdmrhxu0PaRpFnB
f1iE0zbqECGPRHg7URAq3aXW/CntaSArcQDxw4tK23nppqolqBZO3ltNYvE1ZiJokHTxPmun1UDW
sOZQtLQZFenYwY3oc/ov/qxsfvVLTDzseVAQ9r7ECX8bCLJf8DUb7AkRvsTD5YTHKVjfAd367j6O
7iTKGVUd6mjum9+Wjwn5iVqKTL+XcTwA9UbM8CnuvhldHYWKq/FGqraM6kVSeR/iCR1xjFCp+5MZ
8Eup3OYCOyFFwG+WOC8T4zq1ADcJDqhXGvxMxQBpHdbKA/SaIC2X5QyRlEuOQkUuFjc0BOKtxxPO
IQ30855LF58NBHTkicqnhMTG4yB39MBLWTfvI19kUWjW5r1aXgstBjTToGW0bY/rXRMWME3mWrcR
aJZKh74wIfbldoPPmIb3+DjATlCIYVzYcOP70dPf8pTnvAvCgOBkLvoMrj7WoDOAeCtxx+W9Opqr
pZO+YEdbW6A8tgMBCntwch6yrrcu2btcJa/cwpbEs5ilJSLD7vvWdewRhvb0pHVyL6VsrprseEJC
DUvfbyebNDbENcxwyddgO7pMbGowqkZsnkOCGVNpYbvejIHIKCcl6IjwhDVF8lBizjwLo/AdE316
j2lg39Z0/T9tb+vYTQLPF1R/qOp/7GqocVA3vyY52vOYAeZ0nj0CA+V1tlJ2+zJOsBQ3NXtvkLEa
z0RhxLFlkQNlsiyuXl4OmEX2J57qwRGXUbhfZa/l9xaVtnV7mwR5EqKMjyehQagyx3ryEtUI2nn4
W/C4w+HSAtIFSa3rXps7Byb4beKWChRT0Y+xev4ACvp1/LUM6yxLa/J6a5GZE4NU3vc+XDIeIhQ+
Vq9ACGfkncSH/Sm00W3KVmcwzRp2nkXeeNeNe68S6oC0xqrphtciclsDelEVhufs0Y+2tt8ytZer
c7EEUTW5WNv74Jp2V9GMsX0zPPFR+Q7HUrghXSXHkl+nKPFnGXLy6viIY21bdct/oJayeyMW8i2B
bqv02gNlNANRMSl9XAO0yMmSql1THsB/A3Tf/CmpI+q4yAnaHLoYlP9cxSeY4LzY+C1pq7cunAe0
TrT2AQJngImR5C23U8PA26L+aQWg+lP6Vw7dUoi7z4SgBmx8U0zhw6ffw9P3sW3AjWTDsN9I3hqu
H55NONU72wY3MjTK1HNbBxZ91RtsF7WRerRKxBUL58/tZxFf2KtBuoh7iJKezjlvt+QQowWP5gqJ
gP+e3AkF1jwFR5kUCencrwuxIBxDkEBk5PZYnfJ9GiyH15YWwFz1hBJ8E4JrWFlhyYcr/ARmJGaU
O8vab3a6wxcLPSFt8u7DqQ4Y2yMBqlg/jfzMHO3G8gpaRxsVxNh4vA4PwEnJgLj1NCrFxHzYq8eI
IWAbG+C1wOXrZJuVDOFQdLHOBzs1Cs48zZtSVCVAu5uUt6jPoV2qKY3PISt65KSqr0a+aDdZYKOM
ZWoWEBeqXQIaQKHlpTid728vA1APYAmuND21TOiM/Ynpf1NQqfysYrP+F6bl0dgUq1M8k1nLyvq6
KCbtUsaG7Anx+uH8fPMRDVWg64mdvxDyStbEKmGZmlzHHYfpbHRikwYDN+GN7tvm//s57kBHVMuP
CxWveW8u1FQENhXG5vsAu7+ffK6a/ZYjcF+Ftjm+e3AsYYS5ZmFj70P+srwIVc3s+3lA3FxcXIOO
E06mMmoFL7zzkElqLqi2zmQyPwSPyy5N8EFyyVPzEPr1gRHkxFjzMtE1rE2tqiFql3T9GTNnklSZ
WJLFwXmzosrQYMXwalSCT7RaZkqbzMRFbGmmXKfroh0B6ceY5hx2FzQabxHSSUeOhW8qT0jlazI+
7FkObW8vXZLRE00l5AcbQsS3szDju/G+6+LggLstBM15VWnZ1OeFNyRv9TtUUPVmG2cdbb4Z5S1p
SEix61tS8asjtxJcTkDWd0n83u2v1LSH3yj/9poXDVpAamFwIsrfnKKkrp/XZYD9oiBwRpth/vrI
mZsKbVrjvJsEXtw17pFQXDmq4HDL/7VYYkXU+3OUWeLdEmg5GxTJaOnboOGXrS+o4N6yDR4JteNq
2U6S444NCh+PoGEDjHJLm9c0C/n3rU3SLMKO/IVd2Qv3lBdTOysyCbLf87auEdvTwlqZU0mwElao
ltLr5RmTKeUYoGbQwzVlmJ2HjPALVNFNnTgHgicWgy5HP0w/7dGzV5LqAS7a+5KutLUZ9TbY84xC
wC5UO7gKA8jI7TLAxX/5WkF/OUhyfKPlxyqqoou06sv1DUpD4sIeI3JKAz9mIhdmdrP1hRM7/byn
nLl98953tlOCWdZJpBEbviRNK9V5MKVLFu08QPRTEIVRZB6U2i3SVmGk9WL8hO1yat+KvH0QD12Z
n8wS1OYQnyY2SuTLiFehmOXAqKJaJU1USsMmZ3ZOZRf/KAAMtN0psGQvE7X+BEXnfvuA6THGv50h
aAn9OTKm5tOWwqr+1vTVuLm+lhYUtQILzCjoov9BDxqmzadEiyYrl11xKkVRDb+T+03rt8ZWMIkq
BVIlwnJ42OxNa4GGritL+bjUdb1oyn8/2fKdKhsnFhGhIo6nJ8xLBugMHZ0rBrCTLy06CN2cSv7v
qPx+IXQaH8mo2NZWB8VomA8dxfnPS/oU4qC0MFZz7BfxN58trQvpHhuqeOP2AZdCJcX8JVQkNKS6
YONc9zR3Fk/AoTbl5w0IIQdoKfBQpkuDWFwAVJ6VFwBE8o5kHl9zKNBFRIW1YSj6hKumbIxQnM4m
sXkAYFWjiczcFk8NgzJBA+zMYIR85hIJ/GjTg9MeRgFUiJbSvRG7IkrLG5G9Ol3v6QINIz0BHoso
7COz41+4NBVkyDzEfJg5ogXqvKnjAaXN67iFDWMkBGlwf+5AA6a/GCUMAjrcYrzQqNLmZ+9flVrM
shPNOhY2Stq2NNi8iYaMaeeJrXoZLgtL+yo4cYXNGOwVmQlsEiKggBjjr0cm1otCV0staM+smT83
dGlvHkOOOKGz3FCm6Dq7k2huHxB5pg+QGuv+k9FlZFDsDJRMdc9e2QgJJ7XvRaVYfGugSnMUDBsw
lq2y3HXVqVkzESqSKD8IcyXAhYn66+0hq+4SryeFa2x3CEV7KcRtM2Q19u7nP1O52M3N7vAO/atC
iAHYBnrNqSqwta3sXmgYyRJg6UrDqODkUKAcpjdOlI+XNNQqLrY1ylrqq56tqHqGHGGJJRuoGPNo
em4lrv2CK+YkSbmO7GP2yBuCkcqrNn2S0FfSAFUsZHkZkmHBkhGAaSYjwlKe+JSzrgnSjpfa/+2t
qf1VveDCOCxDpbHte4wNHan+V/XIMoOCoEh2RbPBHkaP4tdtFReF4WNTH/K4BNmgQhIMVYXN5tYA
u+/Y1nJBB6F0XxeC68KSHGTucBGeKO7dcduHAOtvUY5D4meb/ukNIJl1+kbjAKIheY+LklNwZi8C
j5jiaVamRXB/lqjVXOe053i32gC8N9v/zfjwh0pyx3tlD32VNsJ1QqqN7UBgkKKtZcmMzMqlo1Lk
2+Ewf1YFRPi4pzCc933fZgrCWF505A10mbvvGRLf+QLInQRUO2Uf7nm8Qq5skWi4/0F9bzBGJBzM
zlIApoqZW5DT0tlsvfZQLQelK+9IeMcACDOU0zDf+It33UMaa9Td1Kwj6AYWliGjodvhE8BE9Mvt
P8rwJsEj1VJOTjyFD/2zV5fI/sozXmIoH7ZtBMRMHz4z+A6oRaFgq9yxTHzJM9R2NpIGOTGp8G2w
YEhXmN0UCfnVK3jmcYJiB/sGQCY7tXgSuUDJWa4xj6rSDlUoleofqdEpVl77+NpIWsUdHL40lHZW
fbfU+8KllPKv0Xqv9t2U++WBGATgwI71p1BTv5Di+M9rptQ+h01AbJrxf+iZEjO+V5YLYB6yn3rG
gWCILPJ4N/F78kB2iYz+RUmJot54H6fLTyXlgwE8N5Ye+JPQ0oIx6rWITpoOtAlrN13baSNitH4L
GE/IgCusn+YdybHIzrYB/A4w/MZcHo2faDN1k1hibzFCWbGoG5hBUTb3So3sSkxjTYbPNogziwf+
3bzw3CL2XMckOg0MGKusFgc4deY7/jRwxmpHoT5d0ou2Z3Tl7nAw8DMs4tUXkQtaj2uaIOr1qQrM
hXN2JcHDs5UdtwQt0l+w2SU2kKxOJUQqVjga0JwvKWgf19s9HIIBTj1MWtj5vgyWyK02kPU2AC04
WTvE0kLqBqMWlTD8d5Xo2TbYLclWbPkNpgNJFChhmX+AFvH5tDRKnGCf99+vUSbxf4ZMuJrVRReN
/Bu6FdglciozEimsgLQa3Pm1CdxQn68+xuXLSMbuB5K6E35kGW8X2oXFAe20wXDwp4sRei+trEbT
tuSnM5C4YxiSAqVV8XjwaEvZLsJOmMWdcMzMCUbw17ZQLNQPy0e1Fx3H8nTevYBUIulN4QWMOs4b
myfI+Iq0gFskCz2kBiJIQ/pj0jkEXAbVkI6kx26SxPxkFOGF6D+Qw1wpB7uZkJ3G8nWwdnDShumV
IEKVm4O7qEkc2cdinDq1u+qCHcOoOmsaw+67Xtxojn+qJw8Je/FBQvbZOVk+pjRrtzaLmJRaRcQ9
egdmbXCWvUBwegcP+ILJvSdkwO0tB72cjYwQmdx3gXRmLlV5u4xojBt1kpaUG+wwD3pIAnF29gqF
NFGKEd06RWGTH695f179YPNCSGAFxcfWRMwPybMJz89mGFBmGvI+CKM1GPKS97KQE6pBFpJD9spm
yvRHwkr/mfFlS/SG658Lu+IZTD9I6FZhmu55s5y2j00OQyAWCsx7XFsGDK2oOJS0Y8F/eqFzcVZ+
626+OH9+a2u3KVnltz4PrIs5A1gUZvsZ1VZEHEcMF2zRuQvK13NKPwiRGI0qfXviloNs/xNYAMwF
l1Ly2zUhX9VdCDcbvJF7LtcVcEHGpsce7UbV2pPhwTONayfJG6sfxFIQYo8kIY9yyg+WBRhp7Dt6
3HEREDo1y3vmxgh908JuxpFL62c4BbsBJtjrNOla3QDRNSV8gcCyWep5WoyOVa4VFr7c1pWrMY74
cncSIym1iuRU69+T6mb85DZMaDsGRmk6XioUMC9J5+aGAlXPq6eLw9fF+LSaE4B1UHqjdk/7jW/W
JMqwkF0U63toC7k1kKXp4Tenw1pzKBy8H1DQWWv3og40j7lHGhVKPHe6e8rWfUWWXk2N/OzQ5/ra
vF+v65DE43FeqZ+F/AgApHdTpgLrzVftZDp64nT8t+5eV4alcbj7jGSyRy6XoOf9ktGVXmZLgngT
enSUMH5RZiDCnIQwEgGMDATd7bnLGRcBA6x1BX3Ww7DrHU0Jb1WZAH4LQoAczw1e/5BTUVQv/bog
qeURmMtv4D8SouMKQd/MHd8dtniXoT2LFl/YLPC8PI3cQ8gMPnqfY6LOsmRejthrLzskLg7l/J8W
mcz0eSCgLKI6NMl80cdjUWeWd/yADNeRvSsviTTostVaHLAy3oNUwWaLZdEoQgv7OsW4fOxP3+Im
/NMHeWuIyrv4uRgKswJh8yvCjobOkAxgecek9gDFIuv7vDnYygVQ7Hy1oTFm8V1Zw1CKoP7GsmlO
tEj17QveIWokjSk21XYrAHgENxqj+7UrvGso/+Yt+MtwPzqYuvsAsXVbFmhCAyC+256airSGpjzT
Rq+Unslli6nW2B1MzMCS0RWc/WVBe1rif9GpWd9r/m7wFVQuz4a9CKyuSTJKUHWTJReoO8WUDLWW
yZn2H21PFbALc6dtthrXYoxFlhsfVNO90up/ZDn226nQrktfkXKIRmutcVnu9NzYNbkt/YJJDLQo
tFE1ie14z/xezU6A7hVYVYZnMLEBvRvIMqlDDV3afYlr4vqW/Iug17zD2MRsuhN/LAZxOTqkywmv
D79T64qupOjCiSQRmHJUAv9pkPCAL+LHeGxGe2cjbaKScJ1OccyVgP1+5THCRToPORYle4repMR7
jUVUjRhCXHsge6PEzuNQkmGP0dA9dHFsHSlg7i1vKZ1sp0Q1e4TbzjCogUnq+g/nx6sFOL/zb9iQ
z3WgJ6cOvgYUFF9jmbDMK1EAWociNWShtgzPyMffi3/+StgS169u0ovSBmn+kRUjqP388xVMPQ7U
3MgQArJrDoNzTFYe2TXKuh6Rr18rwicm9njheOTsxYb5ovnl2nlUh3J3fRiIKrcwUIlEpLs1nKlc
LamAmGow9Pjvdj9wH+lMnLgL2Fk2WWK/To84dVokw2SEEhXXO4JZtjveyEtT3mPPwKvNglTuRwRI
gLfNul60qpyFBqFo+aLka4sGF6zWAMllFicfg56qELXEHnD2ujziuKpmWZmU47jyr+j/qY0CCWAZ
8u916bfub88TfnyqMWg20zh2d7+HvqX1WELQs+OjEKFmOlG7dj2kMt/HQ2e7olEN90FnHdnK03oe
7xL9nU5fJTH7tJm9fIUDfPL+6Px+4L9MUnZXCX6Q48PgLHVhIWUS0Ca3A0aHTydXKEUwkqI4Ped9
rT6xvg3i68szONKZ8YOxMWf7WsaD//+jyBqCFYxQDGyLEci8B8WKdA03/9NQIK+co8l8RhNOYNTJ
iqIOMkcl1jWJ/wOW2r5Rto9XdyHC6OQgMWKvmqCGXKYs6UOZZxSe1fI2EIpYddqqYK7TNcpieX56
VkA7UUGxSbfuqDZQGcjjwYlNjvSMInlGcPCutenSsGnvZwvSpEe0dk+da6C73cRBC4Tz952uMMrE
zhEvxcoAhIOgJnGKPV4QFPu0QfBl8E+CrCcGMadhem0PYaY282J5k7AvsxeDVNPF/viSaEcWg5WR
517c9UHA7nEfHpBKwD4DPORHktwOKG2tdq9KBONXSDbRiiYjsQUoJxRDE8GHuk+cErrxJ1YSWAn8
6Lzuil0cY0Fu0dCo0xSuiEF8X0x88PhAyQ39RoE6nZotsqIQffivxkK+zas/XsYbM2GT9sIdgEEl
uTbo3k220uqvUdnTjmLreUgv7+v+9x7zkou+RDuzL59KYaOrJLmFpl5MlIbcu66ExrT0ofYVAvMd
/p3uHuvQnz11Ri7I+MH/Ypu7viVBJWO2dhX+P0tBTS47TDyDA74j4rPklYHD0YWMyNPW4nRw79MS
GciUwG9GxbExc/5me1zX+LZLoqcruwqp6cMVjb1DCKutAAraczJXJJY7KfvZgAiCK1wUqyvAIOqU
XFLlXDgZXnVEbJbV3enh9s7xxzSTKr16L33+VIpGJ+qy8z9MbRMj6qNv2WFbegDQCD/Skp0nlEDM
WEmPB0apFdjpaOROFnNmv6yz3CxBhbitIu1C7jrI2JagBn8IupvO+5xmET7bK7w73hdMr+A8Mjsu
ajTr8oK2/31AlPSSvtn9btWXz8CxmvWtIVqSzl1X2G2gSiQzVQ1qf3wipeGYngRRp0F0e0E8yPDT
L06JJxfoRcYa9R+tcm9EdD1zpW5H8nfqbxMbmOHYCdJmA0WKE251JvacbMS0DnKvjo8Leyt4Xelv
+Ea+jLBQTIN9Oy+ZOpvt00VbhH29wrFfTMdXbiFaJvv8gMctuZxlJt+8T7T6gVcgrC27dVfOjX8E
6/VJtSyeYf9PX00NWOSUGdKtWrFq7M+2K+d9HnIb8/gJ2kWhiJ1t1h8r9ajNdUsiYFcP6AwLgrjO
Ibv6Q5yikghmsxYhwFeoYf0y5eDAlJsN5KQw3W/M3mEo51wqoYvwg4vH2eDmi5dpSx2ZWa5D5LtV
OeIzDPZ1K2gat+Q499X/H1Eq/KfKsKLmynHGPTwyJ23hgMEtnRI2cpxAgGTl2LBO8cpGVqFgyKly
4F6cCrYt5o9K5nSIFt8q1JrOuQvFNTl+mBpR3fITAgdu0Ggp+GlH8CpCGLxhZ7a3awMAxBwv3FTn
SflQh9qd+dPgBXlETrGlU4zTJLk+cDrcnNPsde+1P+yCE8mAP6WYcb4SagXx5kKBzeco+lbnFl1D
2oIcHWBNEFkflG7pNYmZyyiPn9zKMU1QqzkBeyq4nyaYW4rvMxpf9DEicEkWckdSPGH3YE+6t/g2
52Lm6uEBaSpDQsQ3wAbkqO4CZVdsCQWNaQFefUV8J2AhCCB3Da7x7KSgojjl5S8+qnWbNam71tP1
2Jay9N/ruzZClhzM5luq2PSZv8pimIBxuSd+qwpGvQulqEYYu53cqO/P1c/z5v3LTl7V4mvYD49l
xV2E/bodUijfdKoRwfc0V7Uvuf3k04fqGoO+XFtcN9RX76AkaGwYMkE7zsxoeNkaYD2OzZuXpf6q
Va1N0kOMnMogsgoXEIXyRU7u7hVbBGpbxYDm4tBMsf8jzJT7/7WV9FEmhuG7/6BHmlqQElzu8zwY
H9c4BJapOTlX2rwAc/Cpw18TWykZdF1sfeqfycorwUtOwur0sBkrQa9d7/IktbYHkq9pZpFcok17
Tfy77+1ZVtdyG968QhzzEEzZjs2wSACkYRPoVZkMv5EDiI8eRseZHACp9v/u+kwuXR7uNWxGzMq5
1EP4seP2G8A6GLrVLXmW3rSUny+ff46/b0EPQNYKbyreis4okFRceTlD5URpFb19VpNYOyHnmdbR
l28Kc3poyvLpo+EsO5WnAp0lzCp+b1oogSaokr2eU9c4w8iQMxx5B54U2OwoeBF4WCmB2YwzTAh5
oiyxxBmGbC8bATbK8FyqeqXOtUSGpvsCwC43JsCBIZ+NQ+gm+BpLihflohybqUDfpAtTGIS5Oa05
LF6aGoaJNhwmUbZKW8fAO54w+4BLLfTdPUqZOMbhKdZ2JfeyhiG/k6YracSsOID9OE9eBkQIVi4U
IORSuRheZuXTsObN+Z1pERt42S/Cg92eejlyqUQEEWoKtVmmNFpvIHwHk7sbWeGLyyQV7KttS4Dj
4lVggfIWyJWIyiLZCY9Z6YR8OdFwnP+4//7fJWepAfSVDlW0XJKH7vd/HnX9oOmNSpJoRIqoZ7pl
iRNJ3UGigwtsngnJQkKs9zMU304XfgjgoeRuEq5RfsBIQiaVGprdIsAQ9YGQf1Nf599rvoGtMray
hNYJH9TKArNwHEOshCVIr5Kpl+qVPGgQ2ZYU4/XpB5YqguUzxgSMTSFtJ32CKxD/uBHmmNguAvHv
BxA5ALTWGfHctHgv84srKBWOgy37tKnQRM/3PrXFK2chllL/DBe0dbM/2wGaYwOsrTk6FjlJYW9P
Of0VZgxeyY5Hk52eUTh20Q659Y91iowYbr5DawHegiB1BGNqHo2alPYQQxLacqkP/7//nrz+kfWQ
j57sgDjIHAiMm7azebTiH24W50l5XDfM4bfJf5Kr1aUQopsdPbUVj8kN3PoBQFV1Vog+JKWqJ0vE
aOqiDIxl7dob+r4Mf4sKR+nCNkSV9ay2sls2bvE/45W/LmNjSuCK8rpdzsX338omXcR29amYpsFo
9lmwGv9TO2Z8gLp0aTjisjOlZ1u98SIal3+ZKshzMd9li/RkEZ+FKNhe7rA7Y3ZypCpnRvM7suJw
vHSI81Ag7q3s3DnRC2UVTeqDtJr4MB4ZCSvRW/D/rq15AshPxGmyppjUbc76PcFkLraL1L8UOgU4
iDJNzRZo0mRT1cdmGt7tTFphKgJzBsjOD65ZLn5ojGCljfpnCaLqA2SXJx3EarUqBJfF3vPdvXOR
JW4994UuqJkqRxBpis137S2d73EAZseXQ/mBYq6WWDohEDl98MophD2G/m63TnY3ifuBspn1I4dX
ODweKG6RIMAAIzNACZYzWy33BZKGpK/2RxaKRtKFB7j4o/zHUA3KkYpOqDmh9ngoDAkqn89RwO8S
MoRfKz343djetnvLwNNZoqWzM9cH9HwIbMUdMdvvWednwzZpbHWptb2/DNpDtppU5Zh5lw544FO3
UemP9JvQ/Cmv6SPLzxF2sme35jczClewPHRFC72pata/vThu8vaPkB+8znCmJiUI5cAPy2EvgCFz
bpQ/LSk2fCTVZS84AHm1f6uGbq455weAXC0TkKUAClqWm6sy2KKGEPtmezFA80suNBO2dKJAVvjK
Q5VdGO1PpyJvvs+c/ltl6dlvaEdCe8Yj1hxmSTlw2V6+cZV/wgjQyv9aaHVweoCy9BAkLhXSIjnj
G5MYcTMIKIR/XazcytLTGusENH/dols5g0Qr8Y4M2DuC5Wb7HccgY2up3qKglVM7CBtl2stkQaIv
jIFHFhWLwudk2u34WKSOfIXNf9n+gS4BHSt6mrK3PRrp9bOvBv+ZsWAXDJilBrow55sxYYvZU9An
5Li4MXTD2j9d94NVuU3uLEcq64KBHUVee6pbKY/VQF+wUmyOMGZarTjDsvOA9UYOSpwz7gN61oSg
7yETtjAgbn1g62AnFR+H4ZhWb71ag2QSPzqP4g/4gdf8hUYDR+8sWRnVmuIONX/Zi0wThBN8EjIb
jOPtCTpjwSMVNeUKf/nmcbJovJKmlCgyC/aGHrhxzVASxaEJjYiMSZ3hjTyUIYQtAFIomKFG6rzf
TkocMVAL5ZyWLlITBRRjmTSxaTOsX4GJf3m56W1HwdCQ0zO47TS+mV/FON1s3Nxx0S3lhiOCLzCu
ek0u3fgh6kGRfEzk86bEwhsj+4Z34R1UbrD8VdBv8QhfLuQEQwzDdgmgn16XM6tP4CHTD7cD6x7F
/2Cw0LOvYoMIwuvr/MrVTQxmy98j0VfF4WYmU1oLtOymJeawQU4i90yLjQQUsxydT5glcZ3mCqUg
Ds34UzqHG1xbo2bidRfFOsp8mRkfG5S91BEfGQfD1cKu0sYW1lzvPmUOvSmrnIPykxeeuHvy9Rm1
MrUA/j1MLDmlLgKv9vYwHnt0It1NDEm0HQ2XSJgnTclTT3zDVqMXuXqQy1vhTNF5t+7d24vIMIC9
WoGtHC3ErhW/ozHoW+BXaAEzlagNAEqMuwHZ9iYH47kADGfBNn5v/USwA6bqFQYQ7g2kDBgoSjGo
ZVFcvp0RnYl/BpsojInskdDJO1iehcVlIy1D6QedBqmL7YoYsqB+MZpANuI7HWb+1rXoOkqTMpGZ
4/iR4pBiTvGj8ImlS6TNuvat3SJgC6Hl1ybLSKr4K4Ldwyzp4PZEGZyr/xTwrthqlZ31SzlP7wdB
/LwEk2f2SeVNM583oUraTdxu10nFC7/xDgHNb5cFKqv0HJyF56qDKdvqUiejcbFMfbG2c5/cbRxW
GRk1eOz6TWoLBKfk4Crng0vL0T73sp2m50OOrUCzQzgaUneA19NWfQ0aVrRHb0vnqAQhCl9RRARI
sHw6OoepL0HE1Nrc7l7vjGWN3HeLcUxFTpa6o7ikZOU9aG8SwbPOuGG8QsLkn91RSZVNWRZUO35g
M1tHu8A6KLN2RV2HMH+YJOOvY7FZRq7q2Ys+yt6drbGBjpNXaKmcwjfRgvf+TaKHhXvLxknpeFE4
n76bvBAOPLDbUGojh46mDDdAIXRXF7Op1oouoQnKJzX3x/BgEn0ejffFAIX7M5aSv8M9IPxSjMkc
wKmI390JvOq90+/TE1LOgNloeyw6qQgWtouOo8w6qWpxbiqumoQzKa+d++QxBNHFt9WKefmGGCjj
5CgztjIGLOOnvg+zfP0OzrfT1wbM0ttXHHpGdSPeAHCpkjuJChsR1cRquyMKoWPcRDw6+1S3Ksmu
8CQaDwVxXqAMA+iia28K0BZlSNq49gMPoBT0DFDOc9lRuMltIAmgM5QgOTVsxYh8cRytqdSYMqNF
rjvoYGqnJqfH325zdwCYGPMn/1uygrLJv1KfevWbUJc5MLrj4B35hVsbJHz8LX2v1dbl4Z4MlEkw
Gioj349X/p8wDBEotGDHeQW6gQLNtog1kOiIzq2gqdszPWCpq6B6yNRIuVEMZWLccYJ1j7uP/4QU
Ai7xFQk/nHcW3nVg9Q0gGbqW85hYJrgW//D3glgP81f0o5HFlt3dlVlGyp6udG9lnwpeax3RJNpa
g3UHOSD9M3WMF/SYQkpfA3Rlh+07HjxoyxymwToABc1CjOEr6lZu+POXbfGMWOksKlDIZDGnmEZK
44Bges36aYfybJRXPwWfP6x1t5dAEDZc6zNBMsJ0eAfFNtUneY7ftrftn+fQd8zXrHHJM0pGadVj
AhDQluSLBh5fsS/ibNRMoANUQBrfePrN2r2859/Yrm6+xRLDS+PBuXOB/NmCnEKXhdR0bpAiZwSf
cy2z0NA7DuX7YBnPzpduyf1dxa/cfD0DhEVfyVyeBXWp41RSXMzZ+pL8yb78RzeRcTcNA3rPbgGt
qbJy/lwG7Di4HAJJrxaKKTzgn3o8pctSh4ufmCsHBUUfIzkJBeZ3n2234r7qtD8ZcFIUCP5/Z3Bi
OqBLB2G6OnA03jTaAy90e651jFoK6IDJIAbv8pd/p8tB2W8R/sQ/gaAxCs/EAorGgnfYim9/1qLw
SvGYv+aB+V5c8EWPa/gaSxWq6yLKq9u30R6MvIXvdCiovmJYDJItXV21sUTN6q7aCauogQHQ9DA/
gBezZo1aXHRVzc26xkCzH7cwcoEXZorkj0TFuif7cXMrq8PnUXRbtDoZPsMXiz3QdsCWghCCGFhC
X47dhygMH6Pcl+yMbP8KAtg+ts/98WC7Huo1aRZNxUmlGmzSMk4GXRhBg6tasMqWVAXjnGg1G3dE
hiOZNQZmcAeMDNT0AUw+lFolAFSyGmJ/CAb5elx+EwLj2QWhUO+vu1hKd/9LGzuMQB19ZAkktGrG
cmmBlJ1hMzo/Wi84VfFiEIlEEikvBvtIWCZ8pMErEo9ZpuEfKm0SCWfrbbj7UWxpzy6DSRB8lyc+
TOpVIGPWkUSDa26WtMdH8FJP94xrlaXVD4s0+tLwLGw9Ve8v/dISdMPtVl3de26uQ8b7zaOcCwYC
EkZWVaxOo9bCMRMnv87wncWBxOqQwYMj60RgbOY9Jzrd2Vw0swoaZa/ft9ZthdQzCplR8uBU1Sfs
0nuWdjRIfSQhiqtGZRmFy9EgvWIAfXiu3knfOG1LWqIyp3FSj0vzwDL+MAxy0+bTIq2vvDwGzbLu
FjY+/XRj7WJPcZdch2Xz8bgZJx+DVL0Y6HZ1uUBmQWZ6GrK1MJSndrs7H+Q5mkA0YwJmQSX1Bhe7
Y1dlbeb3vVa5VPy2PYGEVXtnr/Vm1vu1hKB16bR4u7i0YLGvd9IzdzCHu9LvQOtyxDDCg5cGC5UO
rHCUDaDsKIT/dpqQajGFDdHcJfEmeX+uyu8xrdg+lMaK7GMp/d8gcVO3zNNii5VNznkFrUyhX3Y9
OqCTc5VTWU4Tjcfj44DK2lJWXgCC1KMTqC5/eqGq7ILp6c0HtWqoUi3HQyrW+QKHiKsaDJ7EL3v7
nGWNgSUNMEwlkjkbarzPl+b3fimRibtcTKGhKdtWVBsQYaDMJJhxRDVqbkF2Zma9lijb3Ob7x/1q
woAamdNY/MKoP9ruhQx2Gi/bBBgyg4IoXjCgOm8pDtuooGbko8KkHWA/m5e4gkj75SUz7wIaKfXH
Q83InLG4Xt/PC2OtM494dhixv5cZdw1Rq8LS3XFidlCb4xa7DxcYR5z/VfskGKh6nNPIbZu9MKSP
M0jRPQM1XkxAXy4b1h5OoeckDVMJOfCcGLs6epfN7OXP6x4jyn7MH2mVMwknJUI1bG3e0Mr0ret3
4lnpM9R47cIgZ1GyBr2qRqN5IL7DlURT1Jr/5qKHC6GrdG8nMVaHQZX2qXyPeEw9XT6RuweuzZWa
V89/0P1SiXry4XkO5lzl2TIz06Jpern/q+dpo7NOxh8meM5tGZ7HDcw+5W4gAUA5JHYzIzp9MLRJ
tNmtuqzNCJ1KlIto9YVaXcYmPYxm9AQVnrkX7H1NepsW4CapRSCaGVgh14m6JJwv52UvSTGC4G69
EzgiRYlkoiL7vg+hSth/R8Bwmpx2u1nZJoMGbbuauV5mX1uQSeiuJLYVOFYQMqUUb/PG11GZYdte
3rLOSPwpzZ6xcAiv9RB3hWOLrNpQdRxPLh5e+E4KFdhNtI2PAqa3ZwMefMOUjusEXtv5IDKyx2EL
STOxXbwj9Kuf9AnFvRgrDFyYysDV5jpMT51T2ELkWd7m9mpV17f4gYUiGySNwqmB269dz5m16QYf
z37Z766t//DuXwWa3j9QFZ5P5FTOgEYW3pylO70lk2pIxj1/R/9jZcpjKGdyLDUzMuDuSGQfOk6O
hEX/WOyzsrOF4kEG8CCLAIgs7WNMbTYyJqzXcwaxMKu3PZwohDnBFssqHCY/izGM12f2cCkchl2B
o24oPbzvUZ0dzkyaJUijvFNPLH1W2OpbUA38YrkE3J8P8VOgPhlGk32X/eJMqCYCS8HoIv9JLBkX
YQ5ymzsZgkQ7o7jmcn4GDOuGwFbf8iKW+sYMNMf2MRTaO/AOfsJuMEXvbY3yZdqWT/35+YaL13XD
Om/pTkMJ9pLCZjZwZfoGjCT1s63UbFMUraLcG+xRZAPIEwxp/8omSR98FcWBF6QUlBFcs8AVuEcN
Foa3UDtp1IU1QOdYQrBvL4xPUtnny5gkp3usk4O0BPViad+V7jV8xNUk9bIRrfwigt4PSRsYAyHl
Kh7lczGgI2a5CoPJtJXThGHnbwwi8DkTqbkLADI353Bxmsif6nkj6njycFQx1j5+sMoFK8UVdrcS
e9sdbAeCMUdFN88fWl32J9Z5KQ0m5QF0+vb7MYPurCcmQIe8dDJWlXxHIuloY/Vmqv+VJSWqZmnP
55V79CB93uKj5vod5ahHOcTYNzItdPQveaE4vvimkBrXMSYlaGIFg7DH2fVhvkIYidUyaqQzKjK6
/9WZb24W2Ivj8cxgub1ZbyqQm98ET2sO81pxmfVRl4NHVW6ihSseWUwdIDLSALhgxhskGC7DCOrn
TMMZ1ILGHGFFPT3wTXDWgIcRhg5EaR0CAflfYJ2NlBz9XQiCkOadcxCDYQSBgzs6guvXRUoSvKDp
vs6XXQIU4PNRRzRtsVo7NsGonHaAkI8MvOPLyqVSH8SLqJqVpzcMCguJSx+ji7zYKXmzSRoAOWG4
W/Q6bBJOnj22WnOfwYiLQeZ+WqjtvMe2WPvH9q92xAlzNWa0PpHKwPyeuOXHQG5Vht7/ViMebZkV
1ZUl4xn2AW8PTXaK9XbdqAGUmylPvHRh+NzR6pup1Io1ckrg6mpL8AMYT0sOslMiv2KxIaj49NL5
EWeNyMHatOI55Bf21DEcA2NBOcvp0nvMLraqnxtGYHVSiCefzvXO8rxqikaS/+bAex8zby5fqakJ
qqGiyxAocNNPyevVzmpRn3YnWmwF0lD6WoICo2PSPeHWM5qrQohtkhgPBXSbo1CAQoyMk3gLBRw7
Rq1PJMMq/1++nyftM+NC2Y59bF+nkC1YLPFG4/EK+EQ45liLTMAeKqHGopW5llOeAL4WpN0ZHAnr
yoTc8DPqYOH8B5oB1Co1YgFpWOoq3s6+Rse0fo5L0UCqkey9O9RfhH/2g+1SCN+tqGMA5i09eygn
4IoUIPM+dwPYBVbOZn+e2A4ev8H0F9tY1pxOzjsMfrTsd8+/rMM4erUQY/KAx9UEPso8HnTLujI2
j3NIV+uA5ob8Rmhv0w5/mvWUs4x6igIsyO9bODQKibT/BHPH7+t7T7U9yNMQrBPJvmdNDv4nDUxi
Vo4Lh+yZQwZwj53vItC+EWOZHDB03RIZko1cb9G/AqSPoNkJ8IdNNlJYO5V7gPPhTNorGTYPsEtt
3BjMBjerrBtZxhjC2F1vSLmEKGJhj/+4DemX8FiudfwG6pW7UjJZfdEFN5mFIITc8v+s9x+w4Old
rPiVq6CnghE2NVS7wDEf5HOQMid3XCVs0dOzk4klx+YvxVMXtn0ecy3JDQ6Oy49alZjxf2W6y/zT
TauOBCVui16Nj7nyCvwV+vsNDND0loRFYEQiHioasdSaH+XMO7ZQi8uhAuNsS2AAHcQpDIayPk+W
sKIHkEu/qof1GGu0nTXnIMhJkO+hl2F5qteG6zXr+lspZxKzd7DKtVLSfzONIoFenAUd473yR3CM
amWHIB3xPNvG22AP1GfrHvIUhmbhOO2PnfIJj7ouml2vBIrjhazFp7rftdd6Bt8NaVPd17Jca3yv
yIirPrh5NxQ3QFWkHyiAk4ChFo+Dh3SzB0ijrSMVDa7siI9qvqk7eviSrWUes8z3rIZVGacDemsy
UnGveY8aIdnPbAAU5IAePdHR3i2/uFa+GnP9cbxhkU5MdhrpMx3JMpIo4jH/A+A19gSkapZ0iHFN
H7UTzHW2O0L0U7XxbjFiu7bd5wSgTBKnIMlVAKCgLgH6GFzXLgSXul9e59Pqyq4zWFpSy0IhK4wH
LZU/BrFwxYbdxm3t2MUef/y0rzlMq1ouGJLUf/X9ul5ZKPQuq+mvbdpMoOfP/DPUdZHp+FcWR7sl
BKIf39BOkxw+gDVHSGlKNwxqfjHVtozXS9iPo26xfag2KikHypqXa1qrS4deP99UvFyqwD2XrUeU
9pBFtCJ+Y/inXM+vf7cu2FOlWYdlYHBLMQXGA2rc84uJPlMsdYfI/IVsh8aa4oI/O1L0kaoO4HU3
jcHbHCWyFMANbyNPFws3UdVHfdEG5dqkz5g0mFtuCXbyi6g43yowQEbJrbX+5ibqfThMDACeQYBz
m0+OZbKR92g9lCEVVfTUmfk4+NfFFmquLwJGhpzqDZa1Gmek/cR6XdeSSCbYNSbB6l6aP0LlcVyQ
UPxSKLIYUYhmswRqmfXgvEJyUHO7xTmIOOyUap4IEzRWwbFcOIpCIY+rak9wI7ZYhroxWHjjEKKp
hkoW1WVBrkoQwTiGVfoqr3MZguM3P8WvEQb4KWqqxAM3fqfVBqFfyOaxBpta+BE9EIVsQf+J3vCH
sZTRTj551jcwaaCK+peJEXCpOTq9kwtn6jHnK+akujAuAmPSeeL25a9XdXZU7txqznriLCvrJnlZ
v3xwj2ihDrWr1ChzA1RRdfvkm69RoxcFd9/OyMTk85RdKcE4/LbIZcGE4VY0rs3IZJEKzt/TFzq0
rkIGz++s2Pb/rkXRa8JY87n8+uUDuUblRoHhw4HaAp9kQ2Fh1StzDWKpFsNEtfQvUh5B53dAs1Ia
/eSh3CW+bVwWv+rsp8EQk8Te40qnBndeCB+nrOmxsc5Opwo9bgIMkdWeoyqCkJ76wEmhmjs69Tdc
WVOnJwf2xcdLyAsbv7k8Gvv5HPs60YxXPLhsB5Z+t19J/dKq+8jrhPHEBEaG5tZQeXCojVGg8uFF
JKY2+OvS9B9MQlLvjil1SdKlydNjlCgRg2fbL/mMmIwCvO+O7C3i6JqPJuykKC9Hpm4ox4aYQCrt
cSc/8LchLwxtwXXJiN6mvWOJjF+cmuACpsBuitbx4nnUut9w+7GAt3jk13yPUQLDriNuIgxwpcb/
NiXFl/UwslLMHM63wQbhiOwaMy/XgCz3YB5asN8FEon53Og0HletgYdUHWjpAYpGQAkQJzUFYxIS
BeI2rVQ/oNiG9WzdcYW9hB6UW6/ww7CVMBtd/+RpNbRsubj1lJHFXSFeWOHQCnvtunFTSzv806X0
navDqlyKAIy+4FKDgJCmvWway4lEtI8h1H2ufHSn86n1kgtCppc75RjL5aamgHmtagiYAWJldXiL
OTIcXkMiMwYSnmSdsfVZmqBBXV+GxwzMm5UZtD/52FZzWmIu/L/dLPplvXU0T99MlOUBbF83xZn5
9w1pZr0z44gZXdgzPcUtAvGp3FDCLMq9YwkxFXhKFLQt+pMsHjBHROBDCVQ25e3X7vU65qlLMPjQ
dh1ic0eISsuY+WLTMrYVRy+rI9HQTi2k0qyd1zpDqUfkIFNImQqLYAUI9D44ck91PIaSe6IkyHc0
Qk2uyl3N7W0zJFOgwQhRskD6Y8KROmfaIkn0UnDOS4k0Sb+k9DqDwp7X6+uCsHENIxey27X6wGYi
C+38RyImy+11aWkinZZ7nz+z9La9IXz53ND5ylk48MvEuOD05rchbkYHq8o/AjN4ZmhAOTa2l1Pj
zZsHsChWxDoDEnfMwp4xRxeEOXOxOMl/bhwTeFLeehVmlNisJPEqG6v6e3htTzBvkjjNEKFYx+oH
z/4Gffl6SrpC1JReNJu4gWKJ9HmjAQfOijdRpPwNCui7BhVX8zWp1EmY/RvnOvo4SP+uHojA7mbg
zneZ6UOot3j8RoCCzNb9XrsXmbgGWpSjQWsNzZyMM7DrtQQC+Ol3ycxLnA+9pMxONipRGXW1x3Yi
RmwashiMry36leUNlPrfC0mqaFqwJPj/pLvbDA7r4iv8vZvDdCTFA5BPtmWVvs4ecZTMgQ1wQFCI
sjHbTuvNWsO88xAmkUK0aEv0LoQ8neMtH9JoI3rX+STMzXuQN+UExFLWuhtGYxuVwvzzRJqeriGM
7j2cx8ix0CNzMNkd1LDFOUHj7yLiShR0pPkDdyzAJ8qp3ursF+bqAT5yEUofIkChf8TybzaBvGjB
9adMT56lvaPR+fGkFyVweHLJmXOI4kMO7OS+XUvHYeZChvv5JY4mobmYKMWwNIB+J5sOSwVTqKzX
ip+lOhB+jP65tP26ajZnjBWF/DRPcetss/0SpwLWx3TZomDLTLWIXsxH5UmumZuVtRrYK8InOVy9
5D7Y9p2Gz0L1b1Wff0GnfI1Su1UvHfCWO8MRN0oy17WTFZnMyyfJWkj7kIiocxGNLaVpCVqBScpL
F3FGrUM4L34xSIWNLatkKVwav3sMedHuPNYIEpgIHv8N5ocHbxyRAQRYKM5SfNqI0vzCCglB0Kd2
TBYMWabQaskWg90+YNw68xHmzeCavksTvmKJn4U0FZcRAayJ5Tty4Mr/MBqTI1VYourSbo8uKuOM
cU9cJjeQGFFiREBRGSE9eFsziYGV8O7/vj8cAVUFLUbJWOaakWF4Rm9+Rlsf/1nj6QSlhetpjs/J
fDRnnYlhhol8UPe5xxoTmKTJ2UdS1EY5BZ4ps+zyShigfFEv0BiG7rfaOm+Ec6CNKv+Uf84fV48b
rZEhoKUnsiWJq55LC741UMEddSzwLrx428OArThiiYXL9SYleTKW+2yVzmn9aXrxJJPL+faKog0a
fKFnNMltrl0koXVMVdhV/HyIYHDOoXTeePhRLcAFftYabid9r2H92H6s7DHSPk1/1Xj9hBJ4OUZD
yOmWuHc7N+yQd5Sq0T+OrGxGU34ojfs8j7kr+GY3c0Nx1LYvWo52eANC27uHeiLDToHIbpduiyp9
GODAn2SM2rnk1PS2RgU1Zi7Q1eHCTC86VRKuSFzJvsM1k9P73WQ/bMvx++boz6IeLBnjCYW6HWAV
cATPRIyz5Jl7eCpR3CsC2QOwnpKZ3dcSNDdWyoV7/r8IxVa3BxWJS1dy46+P4smA0bcMYy9RP+rd
CrxBAWeqI43I7xgaaPFpZnFBCnKSZhS61wJJy8Z04oJMz6Q2OdRYo1PJ99rb6KicQ0/oQpKHDXYI
rBeQdhvx8D378NiQ5xFR+N8/KSskkVKKKoDbVHhIPW3BP5jCkjrBIg2yrkJaH76qElGzu5b/9f0G
lM1lq7Fi99vybb9/hp8z1d7F9dGWBxTs7CyT7lHHlOK1XSRqKLlToAALULx1z8Gnsp5nMNxMgH7m
dWhinwXvnWLmIN2+56heWflq+HudIZZXvfTronxOFaMAy55uy4wkeis0tsxUurfd3heQaK06ld0I
MfVwLcJzryk7lP6XPGTDZpYoizUeQugWdRpMyMVZJAYc6nu7mvqqaIkqSiZiDd11Q1up78kZST9A
Eix75LauignYi0zDp7eLXsfpn8t+lQxZvNbjnETvGoKu0myL4rvFWD9jjWUTn3RViEhLEPq7NwuK
S78oK2j8Ara9pwfmedVoatTFabQnMu4jGqyHnZKnw0yC7r/z7BJT45UJkSOf2zxX0WzsAUE0h9dV
RzjoFbcvJKR04FXpcUT6pQwozInKJ4YEFUqDTSig8q2PrSl6/Lf2nhAvYX7D0H0sr7dHfmUhcWtc
pCWEn9q27MWT2saKbm05ZuXLx7pWXP/vbGZ0jeQnT1HMhH13CqG8qIC54IgA2A/6o0jBfq+BzyvL
oV/b4LIC4jp/P/jTQBFecUdZpEPKYCDrfmr4xFwJi25xV6KLJE3MbIJWkH1pTzmygU4DkISfZSAC
N96wGeixAfj2gh9SE+rrIs2XifVZKs3D1m3y1R5+pEFBrPh/Z+qqdldUfxQHFinpcufvfMaoJAaq
pEEJOZ0MYjVl/hw8WdGEvVyiOQvFU6vtcH1HzVYzhBNY8Asq1uCA7eNhP/+9LwNLpCQdOy2tdU6K
dEK2Umb5MXn0L8is0g14D0k20rIAUFlf9zbPxYk6ZAhSCNeb9F0i0zzHHfbRP+Ru6imu2VD9G6hx
iuxnuqAfIeF6daYniQiXXcttLi6QAVyi+FF7cHrPBpYLDdz+SzydvfKj25vpoVYKLlniXSEVnM79
Ef/DbxucJDhd9T/3DK68hNSdVBDMYGj1+oBkNTPybUAd+jBv4nTQslmkh/zaXa82h/vM7Jdv279M
jG2Elm9R5Z+byVw92UjrBdhkiZOq2PC7FDen0NAZk5JjO/9+Kway7KSDo6HUqxpsug0J46Vu5cqp
v7NpwI0tG639KSxnjdhbB87xgfiXajVAipgdAsv2U3b9AhF4Q1ZDqf4lF055dCgNhBsFtEln1Fcn
6DHbAwpY7ZrzUz9VRBMiZvzF6lZtQHnzBciZRtVi0Eav1w0eq0rb3vIJrdscVntxLeCLYgm0TI2k
HgHmJHFQjGX1LB9gWwmxzJdDtINk0L51mPYyjlWvDBjVBBjlaXSeNbL38cfsBLej7VN0vAbJ2vxt
G4ComsQzZ1Sxyrwl71FH5i9BV+kybbtqWxeHZ3LXtkWqxDQNJYZiQq5pfaOkmhvmuU+73j57qiYk
R9t3/9gqiGLqgMi73bu1NJ1nrrcGC8HBfcN4vSyDokRZLorveJq0eshM+ThSc3LIEJuc5k4EPXLF
Oy2zjTxyH/h/CYMcAmlqycT/fJssCHtg+tOPq1zTy9tu0HhT9b7ddssZtx6D/j1804OC3+t4Hk/r
2Yi4hnY1zKRhpaAlpNQoa8D6m56YmiXYl/ULQR6H9Fat+shFsCJeyPqKyVEL5gTN6HNXuazxCiJA
KCO26hLwC85JY7rZLI8T6crCaRROW5U6ghYDA7ixWZkNKMuppj06GaNzru86o6/ny0ns+fqx4emf
5XZ4tMZky25TI/VUUn8/rBbBuwev44uY2A5abkjJqtJsVHMl8xDNW8VKfeXryPPBOgl7wnu5RjOj
v+aUKyLFF9R5NgUiq+oDVOfW/GsBA2lI3nis9ZcGPeLb2hBW7JvRblrr+GgS2UYO8czBuMe5bxEP
8bApStWnYc15XRx595flgOKE5Y4ulirTOHyQiaHbPa3RJUt1L3TtB+CXqwjCSwuBRBjROdRLg2jn
DackvzpH70KFSRY3zmQCdCXqZtfT9QZ20jrMLmSFcFOkD7vLtjto+wwxuDuxd0iokLVRRt92dqZ/
XUkOcU+3gM+D9z8Fnw5ygaS0kyacOmvyghGYnEEjgcG9lMh6ovVxmgaRa3bTj5W8O5GkCdpzQseF
nWujQvx66kxTK8d0vmnuiW875XL5pe0FNrue25xv3c3VWTbqbVAXU22iKpm7GDTBJ1x8plhVnApy
jNQ5pRV6HDpFL0SGDtFCfsiHdEj9gmqvO3HlFaCCDd6bItVmwreQBgr9FF9+C22NioZx2EVMWn/7
JbwGSyW9eUIHkBPgnT0CsYWmskGXBsUUdVZFelF3OrwCutbqQxFpfUWSYWkZ7kBt45XrqABJECEF
Pl5DVMRSW1q7Bd0ngOyEibQnGLHNIv8dbAlZXI57AytQ2JCc6ll84HpxLPErsrItfycp4fZm5KH9
jrqQgGWKMhwyHsl0EJvWTuoSwNF0eIVAXcvNvNWP4kxThhoEHKRMmwCFpR8IQl7jvzMiLzoBNbMA
KmJHm+rChF4088nygnFcpL+fU1oHHe+SuZmGEoQSYX5TEbpwOTVQUz+IO21lDhDE+iiD9DtssKtU
w0hrRjqPfdzMAm2U6daQ9SiiMuOYsAsXTUrcctnHRySm5nKbRRwPA/7aba0oToM3u8clLr34GMYJ
c+89yk7VVNUxjRt6QklZG/vJB70ssz9w4WCnHNdU/MOMqdl+yGh+Zx//EdZZr4HZ4jiH9peRj5Nv
XQYt5mS+vmvk+hLrRG1KQgv2MVvggzadHk9oFDl+0o7N7nRquWiOwLA7yq68DxLGF+z2p2DQDu/c
qVXE1RZorxeXBKzK8AZgN0Kixt5QfIlZLZKAOtdIwzSucfi0+ZaEwe7x3J9CqqmE+9Lg2Ip9KdUk
/E3ygsmySkxnaUUmdM/dlei7aYuJEtGnHmidSHGOyNBKy8dhFfUmhTJpHUSW+AQVptfZBuogz/08
BUV7d+137PSGWDr1xdbKKgolumFU+EIY+ItL4Iru7/vXkaMQUw4wu+PzOue9xthYX/oQoGLARuvh
8Zwrw1/MC4ghYbrK2prr1aUh2ROfv63CbarNjMN19hL4RT9Ie5BJyhcoffAD4prE6zSmZ3gcuK55
eH6frLaWokrgqSaLgoqg81JZzYgEZV/CiiAgWURWDCC1tAh6dd4RaEJTkr24NyA8NsQh0fG89uIl
fS7jz6iXNUr/tBfngY2bCnWcJn9Ez/z6ICeTFzW/hVHwKPXJRNC5HCjVaidLMEky8ghah1ZdUKEz
3qMzJuRG3egnm+Kn5z+mxyJ3G/CfT9g35s/DEpEUVwPOHC3Ih6uPwfFvUiVrA8hkNHMGQsffLnrR
gNKOCP9W4zcM25XRiNB2TFmYA0utZpyJPzogz18H3+XqyVnfMnqvS1RA2ZB0q2siwW4NJm9N/4Ss
bCar3KDxl//Gptc7TeFO83V85vmC/tkMWJyqN/DUXAHDt/u0zbSJxtbLqQPp1zDtDHu6/FSQWbXz
53+JLztO0phn23NYY+3lFm1/Pk0OzcjOZQpTwxWyYVdGvMaDzfGbu0renIOVEYTiCMvnrdcDYRYQ
fLGc2Jqs50ByAmcFBRLGCTMYEoZ4dXiK8Nbx4oojhFvR7uWUNmULncc6kwqtwwVj87lJ7BNcY0RG
uprPukVQiJY53Ir77tuPcjKSQB2muKzS2vO0V/53o4m47Y0lN5/J3+KibLAiT3g4DqXY7SrhsERi
RdjwjBt+DvnzF4NQSQzI/I97h5d1PjW9RUIXQtybUR3+R2Qiaca34hH1thRMIm+FHLeeFXV018/Y
qBHOWoQi6JvnP9FN74FcrPcoSoBGID/DHQ9nc0DT6tKcnnYWcG+51CntReknadrZOaiVvINuPzgl
sdVuFEkdfiPIGhr0OgjtI5cCITH4Nu5y9zyM4fVNalptYHx8SlscFTI6agZMd/+5an3ob1gzI82Z
Yot6DquKhnCPJ9t2/Vfkw8ywenjsSrp0kZ8P1mSKKzrK3+GuYVMk4NWqTAaJF06FZWTtKgCD7MMM
qNu/xcnzu+cEKFHZLhnbMQYKQ7GkUzTQ+J8bKuKrhtks7ECUy/5h6uRmeLb38Hb2yD4P595hpUje
4yRSGdcbPGNp9mwPSE5XWSRXYsdQG71B8NNXg152+NyHTs5Dq/qpN+LK5na/OOXQiSmhgun/UYNe
tY1HYTiJBRgfnWeeBip42AFmkmUPKElcGCDQhQ4NEVzJkvF3JgMqCVyWfP8dS3MFPdFeK+CzH87p
7z7LSEWzZu6y9VleWF7eB1Ut1vdXJFmjiDsIdBP+OJc8vWmyxNzViJypKl2c+fKawReIGge5jskl
O9pLmSAFcMjJWCCdrBv463LNKpafP3Q5hqadsC0IzyEPIstEBe2Om6MWBzHZ9A+KPdNNLZKFoE5e
4ijlUiF5vV6bsptxnPMsxrvUs5+TTRiL8J7hkmHhoJTmq4FjNH17bQ2I6S+AYA7zwgPPnCbosRDL
eBbRHAwpxFsKevwsZTamv5JPbFqrkUWkw4DPoZy5o31vzVNBAYxQ7rqlcphmpiqAz5u1EVRZRJOb
2ODOp5Tofdji4Cs7TeRYKYlDPKAQ/ktYa5UqFDCgOR7IrzLetKAsLOxCk7/v3CI/X/jUaDSvcg/f
uVH4M8+yD23IESxZ6YKk42JHPn8R0e5HwQMrKAj92iBQOXqZTWvouuO6DGcMp4r4dIJFpAvgUjEk
89OJoFogqnFN8jGdFiKwXLBF5W/RgxqkH0U9Zf1pKwugj+u2GWSFmjXSo+aaf8azixml59Ltib8e
O2GpPCQi9Zj+0fTFnaDHV5WJi6uhQDkHHNxLc1tiK5DMAOiPiz1yTF4CkiqWpz00TseIxjYEMMd6
D7C7ydb7iqLR5HQjqRfQ9BH6C3UAh+DlteQHVdlLgY+N/cLOaMgZNigYsO0yqGtzu6gSPuUst6Un
wNutgF1kpLdP1nB3KbJIxBjyTS0lcts+h89uTjNUKVG9yS8flTfBEcpbHZHNcETqqK7EXviYQvsy
5F0C1kDmevwkxh9d09V2b4u3lyuQgGofiHngxz+McUAVJpcGKIfsdCUv+D6nzAAyvTRJOUGPzwr0
+oS0AHf49F/nsHCrcdO7IuqFKy1qUHZBkOYWpBwlfMvERda6l9PrggRO11ct1LmxleOYr79PxJ2v
IPYez/j1rDi5VBVGS6KaXloB8oV8IUsuBNT9uK9uUmqaXq/mjfXln3mrQryU59NnGELV/DqbTI+q
ejbVRXuLvNop+ynZC0qSc8eK0BJe1Ld9OQ0CMaAYe1CZ/GhvDv6Zh8Fh7FPARlqPqeW5LEdDDIUU
U4My5kVOIZvRBiLEd3WhofEhQzezTMR98t7BrwIOcRwu95R/2p0OQ8GR5yv3EToqIBumroPdHNU2
YLg/tPzgAvClfqNEIVrsqksUpbTfeLuBvpWU9F18nd6/d/8ANCmgf4v2SFiBvHep2RAutp+iLFv9
AVN8WoSY55y0FE7LiqUjhFiC9C70k2rSADq8rCmlrV8pISFs7XSE9APOuLmCrcAbnPZ4opfRMBU1
lgzSVeUX41yKNcXMJMM/DvjNcn7wa3VepAdmnNoH7wxbGaTwNjOYdOE7RyYTC5aYNyETajh8NIh2
7Px2guZVEd1+CprfmF5BHsHgmwJIxr1yAmAeax2fmFLbq2Xnbrm9j5Wbf2fSFw9QI6F+2SPSJ1mP
nc3oxAduGIbyDjDGhJTQfB3HAHxyzCjvqOMRDLW41NoiyhiEK4nUkd44FYPbkdMOeb90ic2uwjU4
JgH4xoF7SnRl/RlWF2L8jk7LJCB/jXmComxfR4qZE5K742q5kG2dTPwd3SUTlX4drixDKdviRjup
lIFH9TlRwvV+6Z2HdtdBtmWqYgV7Z1Ja0ZMeWqpFAv+SlQl8xjSwTdhbTs2zhGemGvFo+BlymvQE
V3eEhl7Gr8w9bNLQhNB8znr14FbFl1Ves1fi5vp/AzqrzYRTgm6yCurd5xQ9r9GoXC/PdAWBpKUg
kuiZR5EV2+rTOXHiWuVR9efIKtV67z2gdZTsjVLloNR9eEj6t/iPUImzu96TnJf+mkKF8uXfnQ8X
nXm6/edK0QGxTtochpFkl+qQLglCvq+lgccNEDvt9hsfssUyXaa7G9GCifi7Ld8lG4MDLCTv+03l
1taLjX5YssiLWx8gVpShHXd5vxrCSNqYEfHlvGy8+Jhl0XjrXiWBALx5+i+DuZogTaBXpo/ECFFi
VyPLybIp7SnayePSEBED7Rdw/69ktoj+jwzfymC+gl7IKl4Mh/hM9JE6eUJrzOuUn4CVdLWPn0yW
OQHxulFeG9zkzRuxxtCZGEVUxN6ie6wFpCm9/HtCNO7yt0AiKZNGwJwNa1cabmHpStb3YAZSvhhw
LmVXTuVMKnBCpKBrppSIwDwI+IpY6QXUtN0TM1xaMgKPJaU/f+2yxbdbd1DYp6nkG+y+Hj9BIHSD
14xvt8vf+aqtu+YLKlQYK5IhQ+FZ2U0Rg2w1BxPo7Fl+41wrLh+en3qsegAKRbbYAEQp4i6+5igh
AhanYAXSu9wTcfZLzLYWHFT5QrBk5dtMD7G0qF+RYxCH4cDzBBBqpvQubM8E0HSR5+UZl72QzDRd
wXAXjrHtTpTZcTe0tCOGyJPcDYpASHCTm9HeG7aDf3YFCq4IJRW91QSbxULM1LR9XxQSvc705yyu
Dj/J533fDx9ka5lOukVSZENdN6dpOEqcuaAWSzKyQm44/215SSt63rLhtMOBHKFmrXhvDGGFatxA
DMzm1bgTQh+1JXgICkfj2HWW8G/CeYJCzy9bLqQ74QuZxFPRJi4PDsJedExp4Sdpc9PjJivgssjA
qJ7QSvoMPI9y5+cpMNEEU8rhhOku1wrrjzgMCBHtUOSAJAjkgEkaDSoVbF+kWzQzGg4eciDW54vZ
zyrDBO+NEmdCu0rHzPwdXT5+j+Y5EKoMxMf5bxTQXQyHfrtUk04f4Llr8m5WrpkpYmb2Nh1D4cyY
p8z/cVkDUSWYsk16NRJz09SKelfVNDt4MTrvh9U4piL6UOlWqeO8TNBLl2UkHh6L3uPoBPmxeqsb
tHMk6Ztu0qOosJek9aUq7in/w1yrYu9QYgEsqRVpPiE9J5X8QWIPrgjNhDKSYG7HXRpaF9lg0DjP
C3RdGagZmqAc2BmnZ18f5hNMSNUWy1HK3iNaoEVZlzU7IrANlPiRmHZl7saRpkYd41/jLRldgA0p
SNKB1ghjPrR34bKc69QhvlJBnK2oe2eHYXUXacL+D4/z7CplGVrFoM48/pVWujft7AvbUtYB9sbl
S2xyrOCuJHI1ae/7j2+qqyJyBh8TfuBxucnGv8/3nV5Ac2ESDRP/lOtcIKumw2IrN1KRdK3uu57b
ijeHAFpdJLHe2elBlX+2UcQTJAyv3jDrAFp48JzJJwLFP/Pf04qdoDmAVN/QkEc11ue3ZRPMoEAX
2fjHOVKuzWiACy/nG+At62aOL63eA7P19LHn4/CB8bDaWA6786N/0iCuTFVfZam1Flg+7orzd3lt
Pw8vIKM6TvV+jmyIGTmnN05yGe9VALIeQ0a8QQEbmh8R5bCvH4dg9mpc+OWQrvirXQEUoFORHFUt
Yz15OdxfOucDVO+32ESVY8uvh3XAtYSA3uUWgy5GPqtXJ6DsTLunDfma8ZrpCbZxTskEnsEkuOU9
9TT7Ex0b6L3VDkty8HpV2uZ2HwB4DkG7ZbkjKocBczyKNFKRdjFVOiMZM2xwVlRzR4dkVR6b3tWa
SROykRVFJVGV63q9d7ITj6M/Kee1J4BarExQdIW/Rp3goA5RFwQgf1wYH0au9STk/cFfnmQ885oQ
Rpop0jBr6OMTIc7GcN5DPjQWNeo4w+IKW4Hnu1PtHBeoGlGb+sVaxxXbEVRUSUV/CjY+5K80PnNk
8+xATJWjt5W95wnTZIYxa89ufSY0Gb6JCJUgyprNlWIeS1HPq9guTxSNWsbrWXZPVwtGEKID2wIF
cDYmvt1ECBtIe8GqLCaYMRB5f2O5HmLcxeEKxAJh1gmcNYca3Kcov4snb8Ija7PYa90VaXdH9bwS
xBr1w3cl9xvjfXYkWz8oBZqlyfQfbyCwgdKzPE1O/vY/eGncSQZschuk7JApN/cj83ctUJfC/AeL
RresTTOqZ9x+xYx2TrIyB9AtaKlZwazyyjfid1Y4vTWrBI5l98C7cTB0mw9KaviX/VPyXINQGtyb
Gw2sKsx3yDdmM5RItm48wcdcQqB6xJf20TO4mOGP0Ew6v8YTeXLOv8VbQDgranxc/wDht7ax9eG3
+1S021/0oiY3bCzIXptGu34Q7HR0uDK3hBhs4HGozkAlkwQey7NrTYSpDqvy/fXN4nEOpdr6oME2
MxFqLVpd33MCGWlAHMCDkNez9Hw/hhrUU3Iagveby1ZUucIcR+CXUJ+kq6lZ9vD+4yr3dI5o39d1
WQeOeeTjN1PQXCOyPMe6BlpThGWwiGpUOSHOd6falgTeppAWajNixBsQ3b17YrriyS9nHDLuq7R0
hR0HCP+RNN0JL07UoRpTb8sFxb/X+qLQUDQ+QUn53KMBvbwvH1rlwEhniFRlQ/Ba0o862ArA/bJ6
0bR3M0wQcR4X9TFV2N8hThpN3YbYY9ThUAi1OpZ68VuMgQyxGqvDIP2twrGAJvUh59Z/byG41OsG
nwL+ZA7OinQnnHfiLuU0WFZSTed+8Q3sNnRGP46xlu0klDbnpY+MKzx+X/45IwrutbgIbxVceDY9
RCEp+p9Uvlbfltl4LQEz6hwCsC7Ch+FFY91OKUW19y13dYIGCfkpxAFRewkGwCZq029RbkopzK9m
fDQwRhkj0RtzHr6OxeWTO7XAbDKNvwVm4DS3V0GH5yNIzUx7tiOGIlCaqbtjL2Lde93bVIBFfNUv
FBZ8MFaBgQ/V6XHSL2xYPZ1Lp3XUR2sXaTfwEnvlb1DNdRMYDaO8oxLu+6PpYpoa7VT6BUZarASV
P0lgVA42rsx9HZu9dkgV+b56d0hhHeUPFA95nH5oD8miIKpn3R+Q1GMP2ew8OKn0p8sCCDIu14rr
mKyXy40S0DJBlDtvW/374Gz/mfqedfmyKAgfRxcQBX+YUTBndcfiF8yirwNGil+uWL27/dmFXFZx
egEhucBFrWW0QumU4skAjI+5XJoDS+Q5f2ZOgT1mnVuELN4jMe3CZX0ERloCn+yS8lKo2i0Ed3bd
OMcrVuy8T9j/jXZXVeZFw17jiqr71k26XprtMZSSTnYT7VFFSqsqOudkRg0SoqbGKJA90ocRAjdP
N+l5+qx/1n3dIcfrLDIKRrhRjvcLghShS9oh16gKSYCpXKHTnjZAk1MmBeHWBXSITvNI2IYVbSId
oTD0VFzGY/PCPeuh2v0xMW1UzLhOqEYM3EvCcDqB297jST8aKqrHVNMcaKqRQZiJ2K5RfbFVuTJN
eZBspDXgBhUrY+uU8IkEr9n8/kgN97/z+IzucxusTPoLBVmR0sszVpHklXntDp9955wt1Z103zVu
YNfp8viNsJZ9BMomqrh85ncWKjYe3W/dm58LbOyFn2ERS1vp0gTmur6oBwT9hvj7e6bDSBxRibSC
r93lnLVUaiWhIo6e199SUy+l8GWbbmWNnDcItxYoGjEwPPKJ4F5p+4IBiUWzZgQYGnxdVcCNk0WH
F/KMzG5f5sWc+XyJyweDY0heuTH9BUE9T9GnWzcE+/Ale9l/LDt3i+p7ETKIRfvpcHz5bNDz1Jtk
cGin+2x664OlzeIS/52S8jd+pHfPcvBbjsCpw5T9dvUyveOzceQWDczOsaynZP0kPIZf55N7tHv8
UwSeXSKGRZlz4zgbKq0R7dE65JTJddTzVkao7ZC7NRVvdUygVdLin1MlYr5jZWpAGjVh4WEyA4C0
fF2cNdRtHXvsdSmQjWT6oJdtPaf5qH/DpbnBOZu1Y2+ga8gjYKsAcfk98oBeMAUNj1UMVi8S+2g2
Gio6mG3oEnPI3HAKs3HtI8YqbKff0VeHTBfxFt3lpd+ZIffjH7+B9NPPIPVk0nsZMKzVypFjzVnF
nmFpJwA2rE7Jp5hRGSGuihRl2ahbK4bS/xEIrMGnX584xGJeessadUbXAwPJnpqlUaZkMtaZ2eEO
QdFMUrFEg9MDy0qiW5YVnwS7Jkz42+N0ehi05XraeZsVIbcfg0ddCRJRfqtPd9b+ZFb02TLfFb91
HIK1V8ovE+dhtRG92ZswtyPZ94S+hd9flg8DpLUftdZi6vIJ6+ta7JSwsgsVE/O/HlIXLtbmji3G
Q+PiVJixbckNvi482Boo34U/t91jPU2qILtTTeYYrS47sJU0Afqc2io1vDxdFRtdDUlg9LSLIEuD
jT5Eu9Xnk3/Hi3Dsb4/YD7Gv4yqr5haNDPCv/V1AsEVkPuZZ67XQI0LcEYwrlL9SScJK0WeOu7RF
+q7gB+goyIB4HQQxRC4qy2Em5K1srZM4I+KpF5RMAvmtgn124owSVs7vzIR9qlA0XxU/qqY41sgE
JOD312/0m3EvC/9YvyS9b5Saexr7a2nZMxUIp78p1lR79hrx7wRK7TrjHDuXuFyhpQQ25FGIJ1We
5Net1pQn6GxBVaZKHLKCyTkMiZu4rJSVCUviaNqbGMdyC19pgeZ22v1KYjoQqrFBQgBJ2PnddqOV
ZvRq7gttD7ti3djdHeIN18dpFhyWMfClVowj1eydbTBBWOwKpYQQCBBrZrOGSRV0qok6RwCHGipb
chWs84SWmWZLan9AmHnvTSUAhTEFiu5G5M64XLghzmKF87194E+IJJojQva11Y3fov4Y0Uqw/uc+
A0e/7aaZMnVlNi5cR1lgCiYPRUtOiNyLpESw9rLeRLVS4YT6m/o1MrZG4A9RsP1aEP7yWOTsdWDv
oN2QyIESA/xZO5uOjDDHrmhH6K7L1Njb8aK6TyXCbl1W1XSVBm/SJzPpSvJ9SERmOJTuYbiZoxEl
g00TDSMWlvqpR8+ooyu6FA1+KnseQyyzHQLk9qXjaeAAnvJrOnnGmscS8x+Efpa3eJ1I4WZYaZQT
zXQKpb69oX2iDaN0yA3mC9bWQJTFdvzqWPWpoZE/Ck1B1VArMRHt1ntLRcmKsbqr7h1XR++IIU8f
hZhhFvv/xtK+rmAIVSCfgXC4xQZX4aF4I5DSHU8d0KJ/c0Wqk6sH3Q08LASsYuxbASxW+tKfasKz
S+h2Q/AjCBBBHKIilh7oq6tj3hvo8hOHnwf9jZr57NDL2UbVmv6fGUILBSLyF0L8cIHALganPxaY
Z24lkwhY+nvJqzhBZ5F3xMmepKcbQdeCrUXadxPijVo4jsdSUc2PKiUhujxt9HfgH+huwkn9j7du
du1Qce/2+TYgZJj82/M/YmFujDpn5p4fp+bctKxEzxkQsshtAGlq4SgAqhKaKOsqC5d9osBZ3Iuy
6ANBzW4zGlLWqpr7tf+l59aTvUxWOUzOWI031SZsXuPf0APbpTRYP/iS/v4jpcZZCu2xfnf2+FTM
mh6W8O5IHsq27PqM6kLQvwW2GEOzAz8bb2GCen2++7tuC1e+yn1fTdSFbCmn4EY5koQyjlvd3Evg
LDN8DC8O8LBZMRrxf+lADG1uYMHS5HRj/t7+uCnp6AUElPBf9PqEZd8OkUrrZoRBxJhJKvr+1anz
vArEAksqt8EMyBltX5/DHKlRL0VjPm8Q+OjxpbAC9zUQzmHsvRBbMCds8qmUgW/00pW26f5u8ITi
A0dJSVoqf6klGrG/xSSJjYL8cyEr9zVHGPrFFgj4gCps7OXIKgdjFC1fgjX3mvkc19jFjJKP5VMn
zbGSDgMwQzL0ptN1F8cVn8n7nbcXJyxNEs4jRD5rCKma68a518neECrPghcjTXGsZ+3YwcWYsSEk
A+7B2UFhiw+PhU48+z9O7wWvHZNTUEjqiAPI4Kg3dlVxTTJQQnwn6OuvErAmV3oOSNRXN0uxHeXn
N1HM7FfqxMhnhH3OFYHomRVzDA2NuVN3kI5gbtWcYx364WBIpprUAVKsIB5zP++xPXYnT4uEqkMO
iNrNclS0tgKebXCM1FyZPSsqClekFMCQZwwb1WcikgL4Zu/v10gfORnyyyU9oq1QslaFI7EJAinc
7pGdnOHGWDck/m4FuR/Exv0cuhb/dwDtWANblWqxv38VD5f0yf4ityzXLKgvujKyiAYji4O5hb8N
rBpMAWNIDy5VibtcEVEuJVy2AwpUhiU1Q5xGvnRtFrfTQ5iAaqwLWWGXE0ttI9mhfrvC74YsVJ1G
cG10Khus5IXsF2y9ThXR5ZksTEGmJtAII8j3W66AT9khh6em/ANcRF5c1iThBMdjC3mMfB/d5CU2
UBOwKm5fS/+1ntSOmHaUSlR914q1prE5v82HgjNCifDSBWgY5sfVLLwkfNn3Gj5hF5x3Oc27DTqW
52gXWu8HBzhB27bbQR2oHEK4FU97DBjlwlFQfukujwK9bzh9u2tdparkIQy4falgapWi2bUbahS3
eDssXfPDPo7suLVCKGhWm52LjZ5ReEu9JuXCLYXCH3w/F+aDOm/GSFnC4D2WZgxHxndUzjB35jKr
bCUVVOu1e+jAhX6KTQiyZcGZGaD0ysAjGCYdvlvlkBxwxKyRjsE5iuIBFRCCHixnz/logamzWMEq
c8tU5d5q5rkL8IixIzkv6jZbKa32UlTpaWsEnaytY7ClpQ76IuPdIZEqiYysHYQFdCFpgcdgrUJZ
OzkP/e2eAEKh6zSGkOgpL9OtxqlpIF7hhXf4dCVnNB81AWvG9v3sa/DNGjPvHoLgtSEJdqXkGNVE
lwPh+a9CdcaQD1AOt5hSWel9uHs1DChDymTurObsoZeRzcfx9aqSjKyiAqW3s4T5g+XfUx6wOJgX
CWNQC+z2pkaXo+LgVX/SSbfh/lC9Hp4dxtXoKUKUKk4ZCKOQBJd1G0l9+EglybqSgkTsEhRsUqW1
TekKTXgv4bwXoORpqRFe2ziRB2lxsz1AIkKVIcmABimr1/KwS5xf4NIv7uV6AixaQ1Z0ZF7P5iSu
54f7VfUwL7TJHb5LCFymXe3JI5Lk3v/zxdD06MAffo49MBFHauSDBcXm9InyEa5DW5cqX/pv0+Tr
J010MPUSNVN78Eojjpghs5N3RBAslnnKxD7FaG11Yv460jQQ8w0dY0TzJFJzgCTeJIooit3dwIhD
UarSiuL25wPHbFewvIJ20z5at0odQWayWOorRsP+Uu4TPWQhxJt9n4uJuR+r+BNtFuJNkIiGwUFB
vWDFiFel4LMpnlqxT9c1nxtJDrnxwIsOAazomOPoMW1aNqMjbwfCHFbkscFLdTkd55Of/SnzSp0t
jhdVK6xGpYFBu5+D0aQK/6hRyt1bITrcZ9KqBDZFaxYpFfZgkNsyjJjv9JxQNMR/P/IMpLCH/Y+x
hjs8fga5D4LMliB3QuWBf8a2nNYGpTeYYTpcgYdUsyAD6JYKIpVhzY8mzXt1XqRJ0qNaTHk1Pvd3
roj0RAV+Fex2L5bob7OFHn5zt3PIaP5JSXr8lnEsvwsSrnJ2ler/QBi3uoBdWXckC8p9XTj05flx
71VOzIk52s4GkX3jtTn/1xKh8imyvwKd1m1UMHN1PUjcIYJ9jui37J7OcjplVkxE9vK182AEPOxI
NoAeyNRLzIngMhQJzTxKkoyn0xjEJJ4BkWDRfwiofD1C1Q+DhMTW9EU5uFH0I6DCMKCAbvf0ueBC
vLSF7qlS62CZHqKAqhWhn3zsbWzow+vwyKIsVWZ8KTL/LY10DIgcmk6DR7Mt5CFe3PfUDR0ydsdK
MlXk0VDVK1GqgX6Frv1mWXg8it+y8lCLQgmODhUK4TK4spcxRZxLb4Vj/BZLy/LZ+Pn5AOzKu4t8
Y3fhuFzNhJ6Yggs+7Pt0A2M8YRuEZIGUycJfE1JjWe7zJ87VAuNLBJCPzC8n3OReC8f3WNb7tS80
sSXIvTgAGn2xg50kdhuuBAVlMxKMS40eb2ulC2VNr4w8Iazkysvi3uEKV/ZAKOZxZKTMvffIwih6
K1mnTYSSjEgO7EA0wHLX5GCNu43dKWeZ9zAPlSrMUJwdvBB+bw+pdbp6KGkA3HPrVSGp0zVnMWd+
37Z1ZLxkinOR7PSmxP9qVY1h8bT/l1lvMNuhiakDFV//VJ5qrsqc+ySQUlMBF3bWWzXmIw9Rq61e
oN4UhGhfG1DLTgOiqSwua7VtJQRfe/eBv/6qKgPWO8rmAvKuk18FCrgG5Cwiunar7ygr43QV9Bua
bkLUjSlno9/XcQRJIAYf0WOwSAxD6ILYMDyTj48+j0WCpZGRC54+zRIq7YZYvG1bYT2cj7fV8EmN
j82sZAS5Jijd39p3SAFq2k/m4OWbd/b9tecOaRnn4+eM0fUUAmdHk4l44DFgYvAJtKnL4u+bCVt4
GGWgZDz41GQJaE7ZshpIUWiN44c5qEkaxwd40UVwObG5frC51P9bCmck7A/qh7Cy6oQzWnLYrwDS
TX26r/8ptHZ6ZNE4ijOiSlaNqEr4yboqQjisOGu/Svmvjw0ELfy+76QtkCtZaJe8dHT1mZ89AAII
1acsw2h6fQVOC4WLnVmKzoEAag8WgHwJrnc5VsqOHGmY7znj2C83Z/ek1oBQ/921EYmmL5ZgVcCE
Iyycrtkt6+xrd301bpGXJ5UKfEPCT4tOgdCcrhjc4lGp2/G8ar+PI8SpEkifiiftfRzgCjierfaY
zsWi29cO3PimUGeTmaZNmJJhzdQxBTBd86DfWveKSttrw/8bsUpesg291ZRh2mLNe1pBbbjytqw+
GsMAJHs1oi/u3fQi2XEQe38d8Xo2WAWn51kUI6Jm4Pjrs2SC4gRe5fC2Qk9d20gD/QYxlBaVWrKi
hMHdEa5mmjdjX92d+YWkA2J0FmIyzr7A5v4geI0xhe7PTjNhil9YmVVmoSC/hg4w4OMzbopUp/j8
DYOoF29SJWpTyLcfBribldDzOZpgLV5UftII3RX4aOfJEiAMsEL2Lff904zRj7S84oFhWbo4dtZ5
/bSrlpkxTarvvpyuu1k5xttp+R6VWfJSzyfIQx54KhIdwR6F/kHn3ope0ezL37HOBxrZ+JhsRtuH
h7MdBsLUJBgovB+YDuRBZa6k4+TgyxUuG9boa+oq/QY9VLgSpBKe3Xd+q1BeGLyHcCKVxpSSZiCP
19TzJ13MAtL2mP2Mfk/bULfwklFLdus/zKcH3x9c4eKBh4M3SKAAWj44Mls3lUlNROcUSvCvXF28
U9raMSOzkSe9H5tx35FJjli89ySori700ni1Kvne1rtEtktSxGdOuhDwsLa4AEVIsW44MtPOQddt
M/DCyLCOKnseGbEmUJ0dHUMGvR/gaUIa/uqt+FOpi7RNnlK5IyIwQpzD5u2jdMm/NLlM0rznr8bq
XqIQOKTrKvT86ac1iLzpV9JW2E8RQOdtJNaAAeAqH0hLY+TF3/KkKQE+EntFLPd6rvLzaBPXWwjW
/wuwhW3dRYVw/nu4hWmhfYAvfcZZJxrH6i91DXpE4IWzYmHhBoY29iP3kl4CdgYSEsOscUmoPchg
aMCtlhRDHHKW0avJX2mvTp5vXI0CGbSFN64q8h3mkcrM8KLXKb/2kUhQjzErgiBrmsp2Hjij0n1J
6BZ24GQyVhx+9uIdbfqGYM3zxwCpMIE9tdTz0PhYQ2ORvQBde9kRNd06gtMhD290cDjdFu8N+KPJ
AVP/mq8XYdnUQ+v4AHP7Y5h3TCbtX7+X6fiFATHa0Fs9Le1lY9YVTt+Y0XTuMBzHnZaGMxLjC4AY
ebQb33bitOho/bFBWWFfVGinhOpP/k0bm9ZSYn+rVgo5+s9BlHzJjyj6DZcB7tIEvpQpy5LFkSK2
FTyA8MHMw8BYcOKW6Pq/uWERqPgH+fPqoUbdQaP4aN+5tzb8g9b2unuPwb8dEA0/+y7B0nx/pOx1
pMJidakMRZn6HfCrgtrAga5VdpXwIt5YVqJVyG5x/hRZvtUDj7szQhuP4o3dqlrCrj+WQBnO+clR
YfH1Zgie2P2dwEQkYRsBYdfnlELtehS6gmZqQ1yAd1s+EUXHKCvFsD1UAgwJ8APYoWK2f1zQ/czc
ZgxZwSooCyK+dNFjZHUhtwDK5g/VCpnjR7hKlHQOXgI1BFqfM5WpNGZK0J2DBr7bbFe/LzEq5BFh
0R/40I7l5HKDYym+p3m3c7qjams5DmX20AG1mqgNZlj4IoZmarkr/FGwNLKs//3wADHB/icLRHYC
/s1rGr6MDQ5EVMBJya3VH9ML6ucQfrFvDDTS4Q92pHDMVW3D7+m+0ft9wca4rJPSBa+l6Y0sR5yR
ZpvthcuFkPG4/3qikDVJFE1KoXkhQhpxm4BEL4kEc+kc6bEsPCpXvHGGRqsQ4ANbCFJ2+Vu247Q6
GJlnyfpq08NaNGkiiGYc/qg/1UxVJLTpPRBbzBJsv2FQaOKKALr9cF82lYHFdRT5DboMCodbdcuB
mqAIm4hTGo13f/5YinFWAIuZyy++1nNgpAgNtkswyIHAwyXosax7nyNAUZPjy8qfsEkpRh1p0MXn
WXC0GEjy0pDH9NuNeFnL96NQwmfMrgHPudf3/K6j/GRq8q4qp+XsBJnL9v8qHlZ3NuDeIBGovR8P
Gaf24MabZzSo7F4017cxeC1oiTrN9M8VrcLm1pN9BK3O8CxVq5Sl9+Go0g3HZP3Ckb76n45piY2j
P4MKdlqL+2pozKaxZFiFX2khq5rS4NnbFydzKkgxnVxd9VBp6u7PpNlYz/2fDRaCXtOrCY212HVZ
gO91lKQR/gh1gzr+oIc6id/hWOU/Cu6flBvaqqQpFAUVV0QXMcayUFzoL51nR0C7g0YmpWbTrTGh
7xEVudX4QH6yGn/SHFotrzZlNZikcYcJLcV7+UN6hDru9MPIxuzqpcfOs6HP0IFaAvP1RVzLQf0B
Jr/HkPDUEhJAiCaOZh/jGWBdxlx1SCqJkSod2Fxy1NW/W81Zdcx6BU/6fj3VpLsg0zIwjQJLT7ae
gg3Nyrr+2ujS/bc+dyIh/Ui5DvbSh5sE1AfN593nqz0SyIGxIUlg3XhPOKobGZTgXegR03B6wzeG
8ozQLYwXHI7nTJoX5Yc1QygnU+lo2g6EpNOA47yaoOEI0q0lrrHj7jwEQZ+ggeI5XvnybHDOu2JW
UEBb98JMhawfF7TPa45QQRFAOcUtQUrZlm9AAGssOKapfZfpK58zjD/xmELMOnjegHvM54E747Kx
eaN2iJ6soeEigktVsArLuaraEFts2rJWZaU8kEy1HUSTKuj82Oam0uHGio+hkSwYsm1UUc79J5mN
4DYeTq432OZ8C5L6VMVOsifqwgHqXQRyMDekWTKSB/5RNDmPPk5xJSY5Qr+GKz2lSkd/iLrpo5/o
7AxgYFHCC58jfTkVCCvNdd0lSFZkOiNg85QYYgSc6/5cf7iQJ/uPPasUN2gZMbn6pCYKx0HUZb3Y
11ynb28Z1TbvxNx1K3tzw0s+dhOu/OP2boVNDz/QhT3TL50B+fNLQChUK2Eljfonw7M2y3mqimKo
/rGaPnVmB4w91hhLkTiTio1ByiNqboQt1dJKNQIwQbHzsDTARiDAyuUtN6cUj1Zgy45LEuFbLvqY
/7idG/YpoWJNc6lqt5zEvG7CHuPSYzV7jwTk4XY8xO0fWeUthoIBDUTpr1jvL3MYoXYcd2+jDNB/
PFwlVuWZGqffSwl/U0nSQage3F0n2eyZOAkBfn9KKsODuRKmc482G4J0d551i12Qd+X5EJuOvYLA
UPXsQKU7u7cAFu8xcDlswm8xV4E3LBgsh7U/L58XHONRlebWxdJuy4NjnBGJ1OzkpgTkb/PDeFz/
SKB0u+RlFdwqiwbTIKv10TXcVHMMK3zmtMcrUWxqAVhyZdWJ2Z/XUe5UBrIm2HG1/PTi9MXC5nWn
uTAyN98aGvjmCa7nxSXLFPYl17sagwX4+NL8STe3a9BSgIZd8V6u7Sb1bwoVI92h/EvDy0puwiUH
qaF16r9w9HDbX7yBxYx5ImehBywsWCYVeDxKRvMAssZuFq8DLsKqMGAWkBPciM73VOtA0XIU/+AJ
MyuLex/wTU3HJ2UtP49W6I9IPtzfALb23/4Q2bD41AODhcvyIO7Go6E1NP3ls8tcX4D9yCnanLDg
BlNfy2Av1Lxzu4LhwPW8d61zjMd1Dnjt16EI1F3Lz7NoveFhiEWweB8WW9c7Od1cPfoYSFNrS+4p
ORqlrMiApY29qM8fNz7SLO8OiZsCkIVfNds6S0jddKn/BgSBsQItR3G4P2NUKZliFxD7imMgfM3j
Th1YTJxnO10FgqGcnga39qTW1bsf30SiPqpJ9eX+mk8hciUCBEplpZkPzjCa97csa4t56LGlagGB
ZyCdxszaCG2tW6wehigiB9KATkakkyYSJSsAUiLba0v0Gi9V/ZCnpLF5em1F0fsXtAWUC7GktSf6
iLR6inb3VyijJmi5A4dIa9PFy4/LAZxGY4w0zqeVe267/8tW9MuMWvHJg1tBf4NySU8VSWFuDq4Z
C6A3kog109s3M+4fch6MYMtpOsAG4Uqal1QWz0xtwW+c/feiuu1ARIww24vWM4wnN1CB+pIshSaK
7+z6tWtSuxOyyAotLtPOszwVYt0YKH28KEetckr1NNsozYjjCjeINuBY4lCNqKeru+q3bTRlYNEW
PjWzBb8hkAF0OdpU9HQivtrEUl0PqWcyPFa1zxa+g+7QXcr7bTTIaYleurDqv+8M2JZcjyhK5Gr4
/yoyFIQzM5U/60bUXkl63lEMnoiJK8a1K0Js1vdjmV+p3LLmXk4SO+Yx5WoD/VTIQ7ls9tX/O0pR
9hb87AC6L6P6REBJOVR3c1uSlWARcTdLqhPe2dBoE4PN+ubXOuHfaDbn3OaZwz12khATnvRi/rMs
6zqXWsTCr2D6f6/imisa7AMJfc/KYNJEwkcTcNIF0JbafE5nL43nemln07h6cL/lFHkX/H6gu5KN
Q8qlGymgdB2yA7bxYPS55O1nVMsHU/Brucd44S8hvxaw6I96kQ4WR3X27Q2qM6MDoK78/bNa6XPL
i4+HTVaDbAbyHSqZf5nWt9C2mjOIaPCMgskc9JrVVzIl5L0Cb6hiKWZPvAgsYdD9sN86T8CSNAIp
azcUDpGQIZ51mTduC1SWUN8cZl/PO334qZyjgyHICrFFrRS7AxZ2YVVcKXyivIoju3VEPgSOrUQ4
G/3WfnMuV1U8fgUwWCwJiIAJ1AegJollyt5ZArliZ5I4FGqbZdS9BTuMlgWJj3ReaWYepx8bB3nm
4U7gNA4xvv81NBpT+PDrMVVFdNIfJ8yv4QUQP9UX5oHHI883MiXgQUyCK9zOWHzsmrCi03fQ2Dx+
PDrfM+xKSaUuVjAnCy6zDSCeIIVHiLfWcyFM/2Yc1xNgUR7NbRKkxoJvulTn4ObZcLZO7ADbOSMD
nxvMFLw09S2MQgZKIaRwcJwV9r9A1x5p8wUaHZ69usviEIpnw9RlfNY9+jk+0koDjSXJMNRDP+YX
JEn96WIlaDC8fX5NimBm7w3U2GkI0QYhBsIzy77IF9LNKVw7eSqaeg7zLNrc9e4qLstLV8jv1frn
1w/l08Me8/KU/7U6GBP0yF6g/Q7RI54UKQthCyH0cLU0RXI0AAzdolcFw9rSAfpwgD+CfCVJNnon
SoV8qfeZlljfd3xXs7YyG9nqoUQi7SEdrmZ2SHHex6xS+Wt+pnJ8+UQYRcOr6uettWtaUhuAh3d4
pAvWpb6Ku1mYmFvo4xF4t7eAuBYbqhj0IufH355+jtSXjOjcnPLT1SHpNgVGfBFgVZ+26olRctlY
5cq/Ppc9xSarESzWECfgw28jSQ7AXWNP1y0VXyZxVmxTcnu8CUMtcFz6etmYbVZOQY62d+s2EfqP
PxkaKkm5zxN7mcgPDIN+cGH29jqO7KBvNSIcDZaxKHMaoOc6BcfON1w4LP6qDcqKx2BHK0se6FLd
PtRgBtICOCn5ONTCc4G4Hah5ossPzymDoGkZG7pq8EY/6homqCZpovaqMkt+LpUEG6Wp6blrqH4t
XcT3Llp6k5gp/ZKytWhLB99HL+l1ocq8nNqOazkZM2tUtMHx2ZY6IuB8wOKU9JNaPQHIt0QEY9VQ
jhANk2XaCdH7Cf2aa9KecfFWM1x7ym/803gc7ST+21tBGmR8Qe+msptXQF5AvKAuXKH/GNEidQAd
oB6yzOGWv3mcnly84K2yt0+JCSgye0HMBqwRF6u7FrSPIOVjY4+pcTsQlTB6e7Cp+846ImgGoNyI
NWmf9gHJjrh4sLkwCuVoU0SuQJO1ZnYmEW6gzDT9pD2fTGTCnl+4YVWmNu/NhCIY1QMChk7s7haS
jNYoni+HocfN5kKqQ+sRi6gq7VHpZ0M9bDypU/ZTUQFJiG6B5mtOr6rMGrD99erheLkZFi+K8FXz
t3HL6GeMxVXiCSUqPN1YOpciWPn88wnQx89AcyuDic2haDyl2jo85W4WTypJFqWY2GdF1P/+a2JQ
7PLx4RJtOan0e269jKYtIT6Qgw+9dCAbk+PaW4UyEZgSig2vhlXaUfuJQcj1yaMuSvXPfx8cGK82
Sp5EcwzMrHruT5q4Gb8KjkFfF3aZWJvJ4+B+s9Zt35hw8NWTIdp3jZ1vDymQfVWe5FhiB0nzs82H
ORbDPSsoXMTuG6puzfAica658DX5LulCx/bhBJf/AXfHXVuxtpIEFtVipvZah9eqWdiD6jWEVHdi
k4WDfQ5R2Qq2KqLYwtHfuGtcNcqqBFxQsoZzZmArX8MVAGfrQpIArEubM+F3mpTvRd+5zJNWymhl
L/vOS1fvQkhicB8xPUCx2g6DoLTNZUkqm7J5rAcwT8iOp7M7dJFO8JAtOLhlD6g1K0Og9coRDQ0X
3C/XzYMrwsow2HJ2XpWaIkTbU+W7B1G6k7O9X5Kx5l0AZA8e9l7YBRfOjrlBlGBkrdT8cQ/MVEW7
NG4gdXItASOLuH9k82OHxlDFIAXSNmD7p6UstOagXCxsuGqTdQmJZHyHtkYnLMQDLNw+cK6LbHzU
I7IoqNPw5khIrNTYSeJHoICPi09RS3OOJoHdwiu4ef+C6BngX2eaw94PPMRPDh1W34ymAPWXuCUs
1GvbdAvdg0kWipB0SNq71IlnRVkq0YC+sSwDwKlS2oNc/hwdSOlmDhJk13F+lr4pBuCxMuAzestl
AOJ7ClkgNpBz9yfNnOJHrlb+ySiWijvk0qpSotOFFWYTPc75U0mAvzPEXFlbIJMOW+Rns6p+2Vav
mY73MxT2fwTfh45d//OTeyHjWm87DX4yIgJDHSoukXJhb13kGIqV89TJ3LpvPfRKf0BQ/TuBFggd
iECwna8gQOEZ7xHWOCLbcjE6qv+vHMbamT4/R7r04zkmUT68iqcEP7Iaum8FU6OiJZKU1KinQzmb
ZwXszCxG9sOnvAxO245U2vwwjDURi/62Vlh0dVUqtCwfMaFHQCu0Dc6+F8c/3Hsl15dPifnvDiQZ
UgyJMcMIsJx/vBdQkYNNgeLU7onXPy5G1mTSZeRPxXq1a9UGqVNUUaaHbWFhggFMRNvWBHAEJg3Q
DEdOnngod+Y3vpSMs5mJOR5lY3j2ft7e5hF5bsOG3JtmsMy6YN+JbT4FYrPM95+bocDgFgsKpL0u
EpYGyQTwAwYiS4v3SKjuCBJyLfZTsJpk988d2pmYuCAgazSzE9szpir7/wlEjQDy+ecSY2GTv5ds
kX7C0XPZzxBNZxgK1GxvO+iCW4Ko1m9ndX6IYvVW+54HQU6C5K2WpaiLN0AtU/I9YXxVZ7qEjSTm
QXXduXOOK7SrAJ9kq423kpWC7I9YxmOT5p8ryYOJYae1cArllaZxYe6L6ycjKlniAZfFtRk0JxLh
FV2CfXoBXU7CqS8WQ3GAkHZjLWUCVjEtgj122yqFyhy131HvXMjBUTLEHxbIqe0qPU11rpNx2Kbu
c0H9ZJcIHLn+pQYbnGQLpb9XQaFDj+k4mskdKCk5ZBc7Sm4r9yTEL+rggHDOPtOyFUpAy0OrkiXL
LhrgBsWlSI1xQ+06iF4Nt6CWVRN+871Ngmnt68tRUxcuffXuK5mKFMXBjFagHl5cq0zYNgTPNGbu
oOqw3BHbKoCyU79xupSya2yY2+KCi2MzEJ6J0THqt3eq1/mAf1wsEEEMq5Nadbr4NHkhlkygiB8/
8RY1KekOHmYuLDOQH3e0VObSYSSHmYH0mROdmbcSHewbPkFzPjsfWEwPmUw9Fr8IWTG4Fd/NqL8t
rbHGzftSN3nTeBC3pdcge2leOv0WKNVE8++o6fa+1gB9MNM/PQHOPYb4jfTbEDq6G1Q9CwIWuPdt
i3MWTaCpk8oLeLkfrsk9a+3aCV9vLw5fbo8fYmQSFDPby5+NlUzxq8Kv56qPyT3xAizfvF8R9RAU
C/r4F9RZIPd8mmtlYoRFzAT/PBmzUP4DLjUex330SR5Ik8zoWUu9wzHKo2Yf/bgtFphwgC77H7/L
WT5josSxQRO9LY96IzlPhUGPlOC7oP0G6L/WfHeRTeJgN0+qmgNI/icI84Gd/6pQ2jJ0W+VeP0QI
ZzVc8DnHLOBqTBo3sNrH9aZjbf3bwFyjYdS4yST946tqdT9w3pGcEQJCvFV6+ZOz+5nfuJ1Kp4e/
9iOBQe8d2GowICNlzies1P8jlBboOS5adSLvdlWtkH+jQwQQ7tLmSwbCiYR8dd7IbbxADExmdh+X
7olSgby9hDPzGeY5uZpDEloJ5ZDXBUsPgJRcgyA96DhB3hjCwMr8TqNJABt2FzukM51pRDV+1eHt
Lmn1MgDIoYOVMnxZFZO2lo6EBVZibHZQ7+LiZ3BjN3pvZmJiB+7KK4KUWUOHHmootq2tnQI4iYf6
vvJmq4QpxuJe77YvUyJusOn1jyqKPZpPi2X334NrVj6MBCZ1ZNBEx7VkJmchblnxqinZpWOwNqYh
bTzh67SKvXFlXpXEr3/99lSaxhnItVOc4yOi2drVF2VTbco45ZcbFQd1CLDREVowma1bsdwst3Bi
wwPJROGB084hB0WQ78dDlQDnuWkM0YgWYgib5vq3V3wuLDmBv7JTYEdLhOsnWCGhQ30662yQzemg
FaUKSR5zw34fYngL+46E2KiBP0pjk1D4WmWRtjdlvEDvRldxYr0qu9nUh1sqjYgWT00/XAPF+KGr
EFfO8KBlsijBzAYIp+56YkfHh77H8chi4kG271qlxrcv/75NN5XQztVpP+y4eJJI0ROyzAAex03o
FBEUL4Rf2uuL8IYTTlul6MlhsxvJlsdgxj9ayDhkJEb+Q8xCKibcNtNZ3YVmR8/JWdozlx5WAUnK
VByAH94l0n5XgmsJJlttHoAh6HDsHvNvi70eqtw6qzKTIgrwBnmWBMQ66A1uEz426oBL/wbOh7PG
hziK/lk9iCxqAFKFaxFHicT22MLFedaNnY5O1/AydulqvfxN0doZVL9DlL9+ny3EB75OsjPV8fZM
RrT39TSjQ1nd+UexNZ1niJNX9SAUnQH7idMf34OcIqsKxqj0dN5VCJE5ZYjYRInHGVtnHnDxMSKq
NDh+C2v+ubswi//WJGm0r5Z7lbpIESjy/VdztY1yq0d27bHwwuIH5UV07DiW74Bc1bKevkimhsZY
NOH15kEeUl2qH7K7nCkqfbYh/WAByc8cMI5kLWWNxxeTqStS0EnA4gjHEpmpVD4qak7QT3JZyx1J
7be4SBAzUJUibjdSpjOGQCyqgmXw+w1QLUkohBUn2VB83Pa9fkMiwjtD7sAJ7+e1S4JeCYQsXo+Z
ib2uwutigO0AEw6Ki+ANvK0ksQedqlsPzCxVCJMWU5Ja8PbWczd3WUL0ZAY4H1vBIiF9/6tnBF5G
OiPTeW32cOOHKbqldKo/K9BTlfp5CIvZFErPTxrS2bjjjhJWQ+2eks2jdGtrIRMVh+QNNwj9VcXG
AmjFypXacMOX7hH6yf1Ge3cKDR6B1L2Xzw3SGfJEgkkflak2DfrJXl8QtSqFg/hUDfOEAvOt6p1z
s2nd1O+edYEOkQQOwnsldgliuUWPgewnnIxIp1Bt9q4zOIrqOpIcv36r8q23BSgEvG9cT9gSteQ8
aB9NzY+3Dlsou5yg3woCa7lC2hP7xs90i3Z3ui40FVClfO/llXJjJsUT5ifiFFx43RU6ZvHd6Z+5
MwgbPuYLMViL+xnRGBQLPs8zHH9QZymqmO5YVzgJAReCipbxCbpiBkptLqZPtsv3JIWdmd2KODQY
FWYkQfOxwGAkLq4nw3F3XSSA13kIZ9tzAvYszS964SFxFmDZILnyflRubVd7eXpBJhSy4lzD9waG
2HGjQFpKXLnE6F1RJMZN2lbtpOIlMr6xQ74pBiYB/rABDY/H7i3hLGGLU/Vbs8tlQpram0Nn4Zy1
FURR+pWZEmy3A6qKAOmVm+gvnmncVGuAbCH8BFKW/qll4ByD2rJcQvIE82sKYE2dpab8hKbjFfzW
PEONzOp0UgxIN3RP3/Tvd/jliCRXURjUltE2embNEzQSEQljlM43I+J2xW8iSj1yUjawDn8UOoZ+
UMvwUBYsnjiLvuD24OfaBhbgou3/ItOcDmT5g0WLQ9EE+rtc31+8X4F7TCckrjkVzqmkEp3uUIwW
PUi4xJjAKTrNbCpQNCjgePI/IGYSTHSvLhnqKl7lcCke35wAo6cWjQEtr0sxCAt0lM+n9Y14XFqa
aOP0taqYR4q+xtq5nLMbxlAW9prjJPIZdHorvAtwuKrr8C7rDMTQe48GIR6TQsfCW7T+uZA6kFF2
jqEt4so8I9pMo6AMieJ8bMvlDTH6j0BauoLiKpipBpfCH08y99moOHjsNlcma65N/fU9JxMSiZFF
iUq5ARHIUjFwjgMeHkF0X5imFdNTuGHqMAJy0CqGh18cigmb+OxX9nsyNi+cwasge7IvRMqRjAXB
vCDfkKG9IxjQi8z7M1XN02CzboX30Y6jMhMxQg3N/tlzW9wNKOhkoRkI3yltVzeX4EvrVX8lEc8s
D9VGZlBp+btadcvWt4N+cKHd32qFc7+o4LJeA6SV/jsKB04M8Rvl0KB8HcOpNnDhG8vBRzG5Qi/9
W6hnbG5GYftWSbAzouy9HQqZnPXm6LfXBrwGJ2ZcpbAcwVX+lc+6T8T4dei7aLmjvp4bzUqua0w8
fGsAFbNKieXWAg8jOn2Q2lTF0rqifV3XXyV2jut3NZUXVuT/LFOX8IMYHX3OcPOjLxZjXw6gz9D0
VmYVl1KRzuwJWCaGgty6tDTTQRhrtxwQD9HL6ufesE5213GI/AAplvyiE6l3eMN9qD7ZoUObk0KH
l5/W9mPB5t23t/xybYVKUx7Y1T7NuZbDdWVH3H6GooroMQN2PcYNe4s6Os45X0kIK87iBd2/ZzSc
NB8w6Y45T8qdnAHGVDK7r1BkWt6FTWzAPIItVOd3fflw8EXKciPscnJ60+Bqht5nqqSM1SLWjWX9
T37JQa+UaoYDX0ekwiJvdq+gD5euq8aIcR8fqdIyavUv6UOJcp1Es9NMOj03M13v3vRYFtT46SA4
opg2vHwnHT7BGG+XwpQ2Q92X3lGTBEH7o7bN6pUPdQDQubr4bKNp4k7Dvdk1MUZzKqDl1ozABtBF
v+nQRG59sQ7sBe5h2tjINco6Ha/1noOATOlrGjck/5YdQhxHplstsi5lgeOFx+ILdqGRWjfN2hgv
2dFaL0EQ9y8pwBDfkYXq07Uvo+tqGVMv65LxPM0Zd9eK+XPF2ykjb8nT8gXE1NkIuOX5NsiLSxRA
E4GgqLqiAOY7/vguIgI4uvNvNkS0XM6cHxHOV/DIwO4QN2cxTwt27t641qWEyObF7fediyZgQHmC
9rlKQMSkw85IBfhsvjRmHPTnTZDJ9R2KzBmdy9S3MkkyFnYCb2pkPdA4dS8cYtXnjKa2cvLnINvG
sVmG97nfCp6GE9WIdgs5lbTPTO0JCWZrx9ng48CHLQyqBbS0+KPgrYG0MtHCCQJBQ4pdTDMxPj/n
OE/lhHMOpoMYoB7hzjeU0HQRYKQpBGxdgz5RccnpHjrSHFoMjUP7xNeAJ1dZypM2WRfnzqZcimym
eQozykwmba9O3dnSpPxGrZFYeGgX0fa1l4vLF2uynkL7T6BeYshNO5vI2hdOPywOS/c3h+KVJ9e/
8EvzY9zbGSJMeIXHLOhI2iQn8w8NXlffENM2lNQn93a9J0dyH4qVbWTWLZId3ftXK9fwr+KBpADP
3FgPCilzDKqm15HAkwZBua9ciuxLYb6naXdXJbFAKb4JKK+9enKOXVOv7TFf5N0SvUzvgwCP+NpO
mWlawmHZxbZnpwPXAYKSF5slRBlQqkSys8r/NmTr3ah4VEmWD9btOc5zKsp6GMun/nkmASbDVONK
DE33pC0T0buqgjZsUflkjDXMQsnUu3kehUAblzQ2sci3u7nbGl6aIKtwukjkIml+coNJTWqxNSG5
HditMRAqkIJ64s/E8SnrAI80cmQ/9TwVA7TS4Hjr3nF6LZKwJ8j92BKFQzUaDsyWMXZYtPEAv7Io
HOYY9nRRSRBR01UOAYtaXNIaX2k59g61DJDbwTEH3rd2T8KaiwmA9rPBdBgTWfV1U6S7yV6Fl1iC
icZnIYYq0PVZP9EMbGB+d4ZRR84MJ5whYRIMQ6b4F8eVyZ/jpXEi/3WhKV8yDdQ9HBs67Dneblq9
q5pyqpV27JFJMDqnVjwnK9qxQ8aGhramBAYDPkfMaN8keHJ8VIGtIL5PNSS+eFwEAIiNncmlRXkn
ECrRWkUVuOKPhHb1spFPU1zJGBMh1WNKmhmFJq3tz6icg4wtywDknCmDdVR5IKYi/vLKP9Z/5FZS
OE+PDxkiv9iq0w6+zE1hLLNK2CUA7Dyn7Eyn6DHMRM9lSqPirLDnX2s54vk0rAOD14P3agDSLRhu
Qym9Z8qPUCzlIeOqMbbYWsIMHfjiuNG4lS0TYALWwBs7JKL21i/p9UfLiSP6E7z6U2XCAVLXM5BE
9O8B9EniIQwIPApc+ZWZXP+RJqKaycECPWppX5vxJwlMU75wU04oVdd9Rt3o7b8HJuuFcWr6Utis
NZFsLAulXG72ijKoLKXrz6Fi0I+MJxZnBnAgOH+JSW1wU4ePS4Ks5q1pQDp+G+ODTvXQCURxxYhK
PQwAtqiFL8twpcDarHucf9ZipGuIHln+COxUffR6SMMDS7YJV3b1haQHadFBnYqJ3h1rJJCF3NLA
oaB0MOa/vABJ9+lDeoS72zTIXYawOEDbXotiwBZQ/tOkH1Zh49LEsbHWOznAdt/byiozRlEVtR50
UliCPyLFp6wA+LGEGD+eTUrQ1JAXGr6b5+kikUcSz05Y4KNB2gQZAZE+F94yECY2Z9YhzvbOPd0R
jrydi5Ci3cV81qXG8bPegPTRGalMGCI3bbhMeH8t244aQYpiNHDFjWTB2ihAq/2dPMvztV+bGkl8
esEjTMw7IoWlYcl8uT+1bOKdHdAb8BdeJ95H1Q0gHGTIu1oCwvY/KAh+MzZUJSMmLXq1q7nEr4cO
x+N1gmzdbVZSAKBKFb1nFocDS8bF344kS2l5x+rHElrE+QlXSd/Fh6AcaJnVqjjjtzSDEkBmMfA0
T6lgzMRTzjKJB74gGyje0mCm9ucQqfqHMZE52jlgg6/92cUZYpVIJnEXak1oUan2TV7vGP3qZjys
SY1xZlR8kMeg01/Inj/q5ENUZevuS++D+mRkCo3oyuB+IoxDYh9aBsszzZf3GM/OicDeWxK6ZfRq
ZLW/vZ9pDJi0hgev7mcLcfVWn9nxlvviQeCLY1V3AnXYLfTGzC/apgopH7BTMKl9/eI5i11mv2u7
ptUG1hoF/SXVTwHRR6wR9bSbQjS3sd2l2cjkjpz9oExVBjTHH+ImsjBcYN0ZWREKaBE10sRja+/H
ktcBVtwkPTzPVoLq7qJLwQUHZOKFtibwviNNFzHJ2lq/B/PRHnJtuI4JrLxJugcw8jXerZgvMKig
yagt6lFOl40mIEXBycCNHG5D/PBqkKs2g+DbaYSYl6PiJQ3ZBT2/zlVHObR06Y/hBK96RauI9SGS
B8BcoBw/Z33RuGnhtmjxhCojz2/GY4MV6H/2145/Hjjb2Dd3r8dM54O9cN7AI7/9UmhxWP2grJ1R
nU2Nf4YYLsbSRtY90K4zIr86dNYjb3sPEescl6SutVmDoKq2SHZHedD2TAU8pXqi8GJVNEdv6avn
Sm6cZ/EVpHpFqOWpNR7hiBWJHpRiRdIQ2hQIg8n8hzvfCMx2U5z6fSLxXw7lEs9QZLZFZKZFUrXd
kupJ1TFp/KdO7/pcSWWfawo8GpT8XiACV2+In4z2JJBDBma73jMDIZ3uo7sZ6MiPir/PFwFwy5vI
1uvidcOgpb1CahD63twrU0lKX79Sg/7zLAXnh0GeECZyZUvnWdknKlKKxoTnarqGcXjsP5ZpO0/2
qOUJj4FMLYNVhXU+YzMZaVQD0h4AtF0jgGoHD4bYGoXX9ND9/1I4NIrr31jD3ljbod2hey7MpGwV
R9LM5BLMx/e7+mw/Epfgk24qrkIw22RZSCYVLApe2HMQKdvw440QiUSsrvO+hfEVmU29Kts2QSQZ
PwMqsMM6lkmZe6nZKTcQMPNFEFJOzStlFnaTebE1+Z9nDwQVB6ELHqHGx4Ye6/5cgqOvMXZnUaFf
msdXdmZUb9JhEcUOv5Y1mRQ08PCC90R7RJIleMrt7Iaa6arHnytTaYrp8fX18toJkXUtlFdyyAjL
jH+EYt3UlVDoec4AvZmO1wnj6+IzFibg0uP70thAvjeaHuNwikuKUkuMzvaPeDGyeK1Wbgfwym4t
LodAq+LebgbGHN8/JFHUTsUljBvVs6iDTKuB/AlY6wgSW+TpwcUgLVyGsBMKznpvn63FoLAiywyj
lc2tDs6cfQE/dBtVfLaq6T/tkrrvh4+rSlzdjH16vkHYvPpdnzBNKng18rPKLHr5CTaGWG1oi3YQ
JupSah1ShUZ6Yj8k8j2VWSlnQo+031EA57YLH+KkBA32EAp721U4m6144BojEZxfB3UZWmAn/mMB
ElBqmadaeGqN3rgjvwJu+6JFcoE4pxKMCvgppGPn3drenwXaad9xXveXVEmLOMFi+emdroZB/rQZ
6QeybyfgQBog+tngnm95Df+3aTXkviJ6cWnSqE+u6Z0BptABStEikuj3f2ScIbHHpZUgmWv48+J1
w23c7g/PG9rV2wFAwqh8Yyjb0UgcI9KLbSjps4HjVoBBV+3gOHG/M1htaWwdxEy9fgceyytO6HNl
5/h63f5pWSgaqZcRhgDgmBxTcBaDwuVckyOgDF7x7AP3zGd/1zJy4c1pikPf/kmZ29Ui2kH1Y26K
Nd2VVIjtAX63xIxAJk+D+mfvmMJanSIK3rAWGmEztN+l1dJK9hgpHrUwniRutGTFrAKdwYduxR7k
7JBnBcg5+pnV7S+BMbqhHAvI9qHpwjmB4o6rd0dMwSSXpYWiat60IZ3PPV94hxOTKEiuEGTWbiAo
l6IBFu4sJsz0zb1YtDwS5MBJ9nPhtu4Q34ZiHIa+CvKiAAJN7BcNgMAUD0mJ63ziDCOA/LSJWhSv
aKsezy6XDt2SRggr4J+78RTXthixzDheC96PG/d14EgF9G0Kfbb7DM1pT93Az8OW8rusl+xvH3KC
h7IbNt2Of3zzhJavs2c0+FsuaNZHoOsRWRbNCKkRjVxOxDKJNOn1bsmSCfgcCmcp+jH2eA0r6cCc
99MzygZg+fuaKQi1GNVr35TuIjOsx+r+XZEJpU7CbG2IwR4SsLb+DEyNhWCz5L01rfS7Vhdpgkin
bZOYEtJ9sw806wepeYBf9AXYqAqYm6GaKbHxE8Pv14Fh/Vml8pxVSviLObVWjp4lvmcPgZ2YzRbj
7GdFtt27sez+/bHfY80x9pOcst4exfKtwXQJqCd00L0+tiFLNATZna2lCrS7bw5Slp1b8EQp075C
HzSZOOLGxOpxoXRqKrY3SVxhgFqbmcTOScWkVHooUKk/d/XdsRgx4BdDBRK6g96qFq4i84R7UMSl
2zo4eY3Ralnzvk/ge9MVedd2Hla1r8mjxvrwbg4RJsMztqZAQvcZ08y7hmM/jG6Q2RTyHCKq/Iyn
iPbvKj3o3gERrKGgSQEWdAwlBJwwfL1J6oWdz/x4Ek0tN8VuQoAKyrS1oLLrieOKkEh14fLw6oVE
7/37jAu4n6hw6sp4YMC+lmBQSEuDquqxvmxfHt3E+zo2CwJTaH/1IKby0yt+MMOZg3Lfi1nfhitU
7D2dJWxUXm4HhqAZ3bEEnXakN1t9I5XZ9x54QC84LSGqnjUcqVrQ7pcshG/Ztf/ZVyMjElL4qy/x
JIh0b+wQelIvEjjQPtK6QV2PvLgyj1qDzylDxk2BnpUddztnG76u62SFkMOQ3fP2V/BabdUg7x+/
rGFroAJADNnjAq8q0qpqAlEOkelX6babZQ7Pg53zarindpeBBJR+ViMizzSl1qi90B/TXllq+RMu
vtufwR4eVdv6dT9HUhIMxkxVyeIQy33cOmsrmJOuOLGO2ZwW+T4z1r2fP7MbR1L88pdJJOaEnIo3
oz7TG70B7SfHpcHSynfFLK3+i6fxXXvfWskhxc6y4UfCf+9KwCSMZYbO1VAlDLmVZQorjOoaVNru
z2se0lbEym5wOEMgvXmvx9ijmmUTPTi9iSSaBX7HZahebv/r4u6pKkgvBQZPrYCABiM2r/o0oVT8
DliKlvy1WA29Kz3V1yilEz07fmH9Q1CW8A53quAiguSKdiY3np3aMtWAacF6EPbhhOoZ2PdyAn8i
8G8P4VFyHkRO/DhNizob9G/aJX4R2NbUpjrJ82420Z/qA2ygdQARxo5nDqqbQ5wPTMVns9Oj9P4T
8NLjlFdFimy2+UbdjWkKXM5iO6eN9uVAaQaaKcAMR6qIRrdOhvtfCYa1Xcp4zWtdiNWO82p3BltK
JV3VL6DuI7ueZi75Sd7v9vKz1cPkogHHKiFrpQcEavvR6Br209Xu3DCz1i68/WrUmLkqkmPwXmtf
ZdLt3YL+OfTLn1EddXld+mwpibYXUIHAcNV6lVlViLgZj+rpAzhoyQWQ41NBVas9Fm6KnSgktyiQ
g/Pa69m5TvYktdif6dZMRVG/o+D2uV4QdRPX28hJq4U2OAR0RXNSMqXnt/r23hhmb0mlQA8IEaFu
5VkDlqlB2rw4ZQiwvA4oUyIWhWzvKHDrANSBsVdygA3qS2uJZrdvU2VMsuFrWjp7DR1fQjMwqfSu
m8uxThmv1vV6l2H+uzCq2zrPaG3lUjSlt9rQYrYImSbUqGmRB9g/JeqxyGe5S1uw/QYJZsMLKA+p
OOgFLOEHUMz7MKZR//cU+FYiAdYraq3JHSKTsq8gdGrANLAUNB75UNXNM3M715981bR1dgyzyFrZ
MhhHsRnZfNDoTIJUvvW+pB0MJsluBeJR9XhzKILG5Am9c3XEFLwr88qR9RJYEp3jhB0gNjvVrLBh
wW3+hFsD2ekExK52dfzZlrBlZjLUDliNXx8crzLPDq4ZjJiLsNE98k4gXnY/JgkDrQnCl84QQ8gs
1WcKi0XVsQLUmPtvAiLEwUiLRWDPU5NYZfv0W7Z1PeTrCcpZL/ZZlteslM5pUrK/+qJjHtxSgDDQ
jMtMoa+8SbveMFiX+if7xiYBwAVBAOUsFIqeVn4HcI6z6KU7wz6s+eUnCD2jx4YAVSJFCLJloaTO
Byo6Fu62S+MMYv60x27cLiq0+Yp6g1bfTiptmaGG/8bL4XES2ItAvGB0d4qpBU4JaMJTsaltBy7V
p1xl0uenq7NR2IrnnpcaVj1PWShfrUo5bgn7+UEXzFyoJvAk4tCwn1WUbvbL2QOD1lAzjI4iytaj
72nWVi3kiwilWapv0V+3Na3YcozTOoYfPis6sDr9WLdXUKrO3tMhSRabZ0+iPE17hIIF0lwNvPwe
mbrHBlhXNeCWmAEZm3Ly2Y5wvJ+kClFvAawhuEL2gTq2baYKZ3nYu8PbBarlm7dwltpeb5IyQ5pl
SvfLKEII+N5QkRLNFvt4VNo+APEDFseb4S6okRMW1LMl6hX/4inPxlUXozat+Oa/MgJ8XtXoK/Gr
G2Q2a65Xtl2SIftJL9KbgkmjSpvi1UDRIhPFteDSoPuzfx3kobebvle6cTSiQwySa8LfZc59HjhZ
x8+6MIuFVQbWa44A7GEJGHBfkx5m0I5vDljjvu7XN+9e+6gyhKgJgHI45+f+zZudO4bpla0yGOqe
SeZgm/lHJblLdYX5ugEXKuNzXYC4RCU9obGQ0jNhNgMZv8WWBdvSvxLOtT8LgpMtFF9pJWd8XhP5
+J0aT9hRs2oi6661HxpnsLicsqOqj9BvMw7aWvelBqatigpryDdanKUEf9dhtSRIp/9PsyqruDKf
6dt+o4vCl2I9wvq+2UlhS6yIjIhW0XYOATSL3t5nf/XRb9El48BOxL5rCEXBSUD+64VVtzhvRrSg
jpCgLcR6MdvXnvBh4fO8xAlhSj7LHQay2so3lNj0RWkP3K0KZJkX6Qab9StXAQWUha5cZ+lVrYMW
6c8Z00iGfBVFn1/5SKsO0lE/mevd06WkAb7CJobUWLfFJZw/ud9btCpAlGlWhqKX2Nd5zmuoD+/7
cviper3a+OLHshblD8YGuOOnt/wCxCYkw28KMJ5dUloqfGz67tAv3K5PyaLz/HFVSqwhzwy1VUNV
wEMnArM11UZO10qXExc0XyYQMrttcEWVqiEpNYMshFPsCaVa8GfcBQX689JhZTct/dxgZ1TBtgsw
uyj9s3zH30iHcNccYsZHOM0WiltGSTm85n3iAwaIvNEcWGlOvjU+LSgC1FzWwblQuWC580xv8p2i
wokFMSS3aiVt3vqD1Ik5xrpixN9+ZOZ0d6mLUfDjm6U0F+xNPRwc13kqUGm+OySH/2nnH6jMIR5o
w0QL3CqUBj3aAvnGtsF16NtrC980nQVd2XvHAcHvRnTwWeuVL3SnY/fMFl3EfpUBzN7RN6m9WlbC
PxFWFwPfdacpZMZDd4Y/Yfh1mh+Y1GMpLW/RyiPadwytMuFKY2bhy2uVcNKaz/HnordKkQY7/+T2
SDy0qjbpvIQAzwzq9eAW0ZwtMq1ld9jZdwnXOc4qeaso9mVnhu7Z4BORY7RDQGyUvXjXREJRvVGx
AyhAgHQry+e+kC6QWS4R8iJn7A9E21i9IzvBtqyVkNU3jV0guZg4jRavdj5FvKu9CI8IUQ+nDegy
yBmHxXTGwEYxzizuTlR4XuaqRnABjXpfmezXest48lT8UsMP8U8gWSAK3gual9WtWYcXJVUNdLeH
1jXw0Mmm4+jkwDT5RbFakqUAeH+SInoHzo88i+G+cdy5H10/z+BU1XFyb5N3864XHSjl94eqLRON
BSopckrzEJAqBfLaJ0Q/HkhO0zps/QWNuuKcvG/T6V/Z0Uml1Glx1C1DIWIOmwdxsetu9Dr4cu4a
47JFQYqTRu6jtFBKCjW3THO3f6esL/RTAAPQW5DUR5EZiSd0sb3lbC25OGtxA26bJor3QkriOP10
myIvRtY74qbKmYkEFDEv8rHxoWlFegj+I4DaT/P0kkM9lERzUHfwnhZCK+0tae2Y3ccQY4sg8dmG
e/r2o4RRjc8ZHKRSnKQ4qQscxKKq6uf5bcLu9IN0GQxSRJ7xeUA6aMG5EoKX6588tWlkwjZ5m7jo
y0StkEjyec1QLgX6C+gjrwqpU/saBkKMPEOc6bk5NpwnPCe6+0sN+haaU/bqfkd2ZwjhS7Db99RO
sorNxDCG+yQD0RRxrK93czSmib1DI+DBaXXbMbvek3ON1AqrZ4cZZSR6gu8rNDHHIetXWjMn81Pq
x6PLzJjwHrwJsZaSmoaqEMZYpC2EyX9tq7ztqjfsm5irrDVUU7514QcQ7UZk9Qv2gTXL33UCwQ0o
u0PXZf/mn1DTd2es841TD+YgakdPF6vv7JRADjOpPssR2ccUHwRwuMzo8Gqd8RE3l8WE2oaM9JfW
gaFgtOr2OTyIz7y7O/lmjfEA+vGNZTE+CnaGDIK6zwc/oHgziRsHi9GAbdhoo3os6hIrCFDghbaB
Yr3c942S/0eySLtEpWjzulXBg2DgtP39NW4ZutQlvAl2odC6tGnb5E6GvCvzvdU0EKLxB178xLHI
gZ+XOoTXlrhp+WW4ZsvkYTVAJe3EDDtVOVVp/sFCvDQMtB6+5wehYV129bunb5emqsQ9H/wjx4fP
qKgoUI0CZwHGxzPSfDm3sJQOsaqJmUJr4YCouzVvb5AvZJ9cBRoPCx+9tQQqtPRsXDVsodIESF2f
JBZIORsrsC/TqTXmJ7W3Kj/bL05cPYpZWuEXsxUJWenGOTTLMP8mytWRVrWN6K11cZ/nlJ6ql7Dq
LB4CriA0+rNNOilh5Z4tIwV4BdQaeDXN1qUKl1uLLDRts32cZ6fFRjzzLMdyR8YNsKHLCXL6u+dX
VYOzTLpvx/WSK/yMj4HUW6vdX1xffvCLvcUE/F+iD65SGeWXUSPxQIWsj7VBY98K8VY+d8fxBQFp
1tUmpD/FtfBUMpJhiEAigPp9Gmkow1L2/IDc7l0pbfnfTIwu6kOdCL3bcVu+Z6Ib+BCEYwn4CToR
JtbDOG2OcmoyVTIXikxeH1+UhIOicI0E1WwYYU+/BBVa6EeEVNQrw/WAMwTZwl46TK3FLLaoD23j
ZMGR/9lP+1cVU2E5s8zHzqZxLTGqaq5hF7yxIPF4AGA5QgU6Fri0TXY6tgKy7DNcg7sihbfAYLQz
mxHKs7+AHFLzQp5D+SaxU5dJ9JrTypcJyoLx9rml/J4OF38vmXoQy9yBVmBeFKKyXTtqjoRhWGR+
YOSG6fd7/yFWCrrfzkPh6Q+GIyCgmtBQbRoS5941ZKMNOG1bhA3nBq3Wk5CaQDf8uIlAcwMykftu
88lR0fPUPeWKtdD+TYpZf3uSNy/xlTAhQfGuC+yOFOOA661StaVA5P1kG9VPbK0cKaSkSetPAuYf
6oN56xgYyvl1uR+vFf/Cq/dq77bcXVyu9GUQPj6lvoYEbVmBySOyOrboEyPBLCukNYomN4PKt/Ao
Fyz6vlpJqBBzzAw1AX1/XxGXWnS7s6WCf26ws23js33gcw34xZhznKKp5oT2p2YDSOoMMrdt3PWa
l+bvDv9S7dQZgRAN+/DB8llmWK8Sa1ASca3H8stcDaweVilF+aZxuRmff6Aj24rPzFDV7XUhnWFE
7qQ91qBqzIl2p77bkIDiZQjIMl+p8+kOMd6ybO2zzNF3Jq12+MuqRcvXRU9PbJPFBihAtqp9nuce
CL7Ca+dgr+eihKRFQdH4IVuyuOKceseObfJx12icSywvJFtcUhTPKQWKcwAOJl1EYcHfPsvDggfr
00aluaHZpEGW4BoII4Ow5X8LbyjotfxNykH8/tMM+lT0gdA7dP5VzBUnsSmUmxRC+Sw007csJNxq
ZSi/pfPFZwjAy/Ien59hzsv3hEO4M4k8DZRjR16BQd0Bm1ZH6ISrCJuJaS+wB//WLX9epbh8Q5QZ
mvJ/qzaHTXx79ROM0smCDciwKHEEjmpfFs+/hZEPJ0tbVmwGqTa5nxiNH538z1BS10RM3s5fuSyY
7q5B4URW897N/a9ItZG+xvttGsHKooCnflfEjHCwZSPjywOqAvttW7EwBVQRfssllQzWv5PrQDsw
wLVi/3CYjrgnUC5sOs90OZ+0c+jonYHjz2TBENC6E+rlKQGDmaIPFjy8237Jrh3sx9RHnU7x0txQ
VkTxdD8PoPs9EnuKDFR8Zbgp3N9Wz6YSK1NGVBjuGS9I808O6sutk5ExcFXfs9vMLWqgFdXoxDk3
bkLTEQNK3bOcQMNUMZqN+lp+P9kMlxRw4RsH5YBnIuGosasbZ2VdirQ2OcmRXwxvtZtRe3hpz64Q
ssEY/FEDyAEWdIfHP88qtF/jO0wxVveCkhP7K13si6ddJ0lH+C8bKJD+RnaOAdWxY9sP2CQKUBgO
xDizSZdB+5VQBYrhZyEBOacP5DUGfWVAzusxW+MrahetuRjbVj2KjBsC74KRZhTtrRpJCUzADfvr
bnV1oE3Lb8M+Qkr71H9WUmQHtymcffTcu0N4Cjo24gcTHXmbUEw5eTUfucE5nMBEuiooeyizSWk0
JQ+9On2DdER9FGQFc1dVV+st0BbriUUPbnDQcKFRCS2x5W6Cr8fLWSAgtTA87PYjv5lGSZ1SQiEy
+DdSnJqe3iLOFa4gpRITS3vplIbeeqPJGdjoX4h3YzUxjNtVqK00k3XVs09qPlFEdzPBoQJA16E8
0Kr8w+uJ7DYXtJcMwOo3sEwQhkJYiNFV7xhdf7zYLtMHD0iopOFTiQcarWvLmXdlZcZxkeHrQ65n
u6n8co0GUPUgIc94CJhMZFX/xsr//p9dK/1pTvZ//ldn55yHUV2wWe2GD8+d132R4ZTwzEgLZ4Jh
Ty4a7BHi9pq4ZNrxEaNyufRe8Y3upPbGzJCHKASs1w/QTkCFXa52HOlA+LaiC45Sy/9ZOjrysWTf
MBufQ9nHepCiqWiF+voqvXCUMEPfFyRazg1uTy8opADZqDyi7Wve6qvNPNHN+1kGLPvAhguWUoCY
E6yw+1GMON2NToDB6juvoTEvd6rQdiu7lXAnAZiITNl7dyIujuCkDHjtomhhp69HbxdvvxFZ2OZ+
4APU7TLTbL1qCbqsuW6+p+XdRUQulniCMurUpBtSC4ulBXZqZHkSrtsOAU/njG0f3cimuQfStxqR
HxZRSJiBFA5/JIDEG6YZimJ2d2srgclZMSid2a8Rw0gmOmGqQY+MKu3v/b/anL2udU6nyeaWp7hk
Cpn4JbP2qfp2H+sq1YgtNYdcDAFCtBGzDIRB7SCoJqgFuSEpZUzSxTgaGZdIJ1Q5sbwBb1xl26tH
RgaIM7ukZS01Y3iX2vUSfegbapxCyGcQtneea+A0aSmh1Nc/ICPN9poFL5yifFAbAy5DWNInlxTH
7JDL5yZ+0Q52BAzJwDaQGAM2lSMczr9rU0DFUyeHnuDdxVu714IrexnR72KeXAp5A1d0Y+SaM4P5
8GqNnxhy63eGqYEUb4S2cW8Zll8vcAe7sz7CafTXk9g7s0l6bv2XKk38L3g3jngjFSg7wy6a1vkU
Jyv4m2emC0y/eK3dvTabMC0S6yD1ipBNcipABw//pnrfXDkirFxVjGRonXSYjeseX+lzkC/2CILh
W7CrFLvl+TaVl67E/DMpkF76WhTQ5lZuaaRPryzXOBxpR7wTeJbO8CL9mYNVgoqrzWk9lthS0z8i
o9RGaED9CEeEBZR5hSplGNkXGPmjrA0xkbTlhxHO/Qqp/xXKKeUPYTjnPTpVY/t8cRVV6WgCy/SO
4om5AsKzGlj6PYYyCXwwdslQYCqxp6kHHNh8hVeSyOCQrUGwRrFatOgIvglKVa4I43rSlh5O55d4
Ty7ZlfxWYRWx/9+Hi/zZuzeFO+XjZb/ElB1gujtNhC9NNrWqccPVdWdzRxEGvchISDBKrO9QbMap
QDkNnXAj8MmFA70MJ4rlsSm795/8UBbZU63AgzKcy96MFfd5hzYOVO57Xl1bZKVabqd1l/2ySYIu
cEXJtFqmcv26prQVBuXHBATAvGg20bNaLLO8VDsbrhRjd+lXzATnJMFSoAMyZySfRkoYsSc3PWv0
JS0TY4jTgvR63797DzOOGiOMCtfg+OykyyP9mn6tXj6jnOKliFKIt4NvFuOgY4XlpOaQmvBydfHw
xFnMMIwWMkZ0FpXdoHzm46JNzA+0mg2vLU2SpNRM+LEE80vA6BKQLVrzIaoa4hr/O+oRGOEiGXWz
tJIGUkvD42Oqd+/v2Y04gWCTE/l2UrQ1C7gzS0qZwESA7o1SbLQQ7iA7Mlluk3n5U4UJ3ZgTpxlq
Ot3fjWejKT/v5+Qmkw+R4VCvvpEsHKueRfxi+dXY0rMKswqTeCVTk/2UbsDMr7Z/XwifAfRJiT4v
aRixFbTElr0bD0xIGys37f23tJBc4Oq7mff1olzeiphhMzAwNEm+EG+gbvubMl5Xg03uG4/oniv9
rIuW8TOeF2ojo0sVNw3cf+CkIck2RR6sZ3iEAHFBms8GSYdIFhHTWt3X9tPhSLkqJDzbv9EtjM/6
3vzZO9ZqbvbK2yHEBiXDR06UmF5Da4JyIJjHMTZpgtJ9Lo6d0jpVWyWO8MYElX59EDP87FXEzNzp
Na+tKEc3Ch2BHbuaH2nltusc+G5z74ahqaGxvgjZkKpAA6C99vvuT1+ceYdpSkjhepgjMnTCikCh
mOvUOHLRzz44WzlnMADnOQKt0ja4+I1SzGO1r5rX8fdTyNbHMWVti3nMieA3IpkgqvCwDP8kMZ77
z2XJclFPjKkGx3fhBd+DK4O7DZajr4qJ6lkUGFtH629TAQwzc1qU0wHhvJHuEi0n8FEPBLr+LXDK
k81DzIMM+99C/hcCQav0hazmUYbSj7nGeN+ypxLATMY77PBlnJSj9OvrdZKDYDtMSCUmAv7q+bDa
j9Ml2cpnvcjTdUm16L3/zVBUPjuZQTJW3Ip02PHY3DooZe8Yq3VVwbd28UmTLotz1lvNtR6QZThc
Jkjv7jM9hdFMwHZw2BXwI1qtoBywTWxFDTWWnfPzEJu0EwXTWy/vE+38Tex3/RqXicjR6omSPn2a
E95vcoFa2Joi3/XPUmETb8edXblefZE5vMuAKWnkzaZ0FiuUfaeoVfpuPfZQL0sGy6rDfFPa61zM
io6BOfiDd6XeoI+vgy/qdDsCi6IE5ADX4i1hFFVeJcyP5incnzic6w4V6jWtCg7xRn3s9AnsnZKS
0BATylV1zvy3+/qzyH//HdWlwVMdhpensb3iguuzvjVq7hNdGpWDAOlLzbMBoyTgADSVfcNuwozp
PYNXdSIA5Uf8XrpTj/TR8kI5VGwErxqZHsqN+pmNepkZTAwywKNIGQEn/H9QVZyH4fOYpLeaGZzF
3it06K9ZBJxFdvxppPiC1LCz2awn7Q2z10X99BIO28/rUuFI6nE3aES9nwlAWWO97l9fv/z60Scz
KgVmRhTqjdqyYEFbHS8uQ6NH9FUm1oVJbNF1QiO0TqTGTtXGfcD+KVDnOA9a36fZlOymVhtMKPft
KzC+wiqqBoURj6CjdVHQ5R9rLPyXH5V4hL4YsdrD9PheqgX9jNVZaJ3BSba91Ha6VTPTR7tCArIU
EEPps356fMgbYYTOuvYIATfLWtZ74R3aKtnXWCImQEqjK60sqAdYm4DPRQRbUk22RWgUrYSrzg0/
ETALJkO9SZ286lAXPAvRPeMz21iP3v5dbtjn+cbQ6LJ5sJDCsqjCfJbBHeVPaR/VNF2OPBoZObwh
nXvntjUT3QLowF9fb21EavfDLG01bP6ybVKGfEd+C86tiqg1Vemtxx2Fy34UIqOupMjlGsSP3jNo
1ZrBUuWLveszuVHita7KiE+FfpVntFPdmtuTXceniH++6Lq+cHJxoYQm9UkEVx3Jy9BXMnEZmo5q
fhKs4e78zY+TuBsLvHWy9thXDO8YUteQqasKVuCsy+UCA+/eQkDhvmDOcrNB3iC7j6zy2M5yDPJ2
W6PC+O9+ggaXTNbBAmhHI6FoyLfcJDEXClsm+GcB8sP4LkAlWeE7tRcr2wQ3jLBPane5/f193T+H
Gc/bo75cf3OrWT9nKFDE8QY/yMOkOR/m6kT3OBpSgNIYXBTVrN0yPqaJTy+94+icEMuQCPTVdyqH
AbhfLsp0AG+LojIKUAQBxy5kkskvWiiSmRVEb2zvomsS4L3u2+sPTYmJozuQ4KVRroFYE+McyclJ
NBqBnkx4BharVWRXiOxpODTm2mR3Ngtgo6M+TEyRp2dl1+uW/dydYaiEFkFWThfpxgLyoYScuXJ2
EJ9JfULRXEaKvgLWzCoQ/YCGeQnNfmDr3W0kVFXlO0ZFq87eHNlhe0peqL78YAQzrz4QsYd4H2MN
51RLHSFnun/RYBmgJvQ3lBOLBNF6B4KfRJ+h3ol4azcmAVpH0J1r5g6u9I9PYcUys6FXEuDpJyGE
FOKkaZvY8OeX2s4catMXwNa1gLNDwvbDT6ha26MN5yx3mvhtohk5q7DAvao4/nFk94nNo9LBdTot
Cy7ZGds5nOcB6ImKDn0jpb//KqrEx5pKUZsUQKRYD20i0ePgqqeSF40srLGNPBX1SSRNe0l596RG
qgoMm6N3ryL2PX1IiuqK1AdWFWB71IcPG9pVy2C2HpSb5iOXL06zk3WRFlgDQCkETt5pBFHulv5q
/Xzg8v7B8HXe2CWp8jUnzHkEYH5qz7skolmfJzkg8YlZu2wawGNVH+3OLqnH3w7U8A0kTMZDL+/X
MzkS7SLOmWZnd1HSYdRWVO9ojEY9m8Ox5islMkJfKCo5Lo3aIaF+OYuewOmZ0LyOGqRnR0uv1eFT
Vecnzzxuye7cthoNLQlgURR/ksQoCyJI0quI25whNP0W3gM3BSr8M2Jl4OJAW+C9iQ+Iax1IfLtT
MdbAzUusEpWAL3yzuxSUVElyEBAQXQigiu8/ln5XB2U++VCdA7uUFeaAJGdPwk16FeibAOv+MMEx
0yQxlJ2xn15DswDnYY0QwjhnWbjgMZ+4Kr8+K1jQeRaYrv8e0BSKwxD9eYkd8xTd7KKBzoT+N0sK
AfQFtpM8kcjA8k1KmJAvhNMpwaiLj4y+glMQNFoU7cgA5UBtjEx1FD6m40tTqU46nx+Ct2MIrLCp
ctkkE9tJihH7GCH69iquU6IE1ubfoU53NtfmcNxy3suFGU4TYGjAH7aJPGRC2Vx94HiydGiBSZwN
ulWsFcojUP3WlGruPdy3S7taXdayLIKsu51IDMNHdUNj6/omIA7DAK0iK38U5n/SUNtu8yg9/aHC
KizjcVRDcA6VnpRpe98I2Ukb4GrRDv3uoVHodSdetD+sV+it08CFCQQNIIDefPoHoWzvrUowVrhf
bUODXv3sLSGIWhUYlAS9U1y1pXiMAZAeabiwIC+CgwWTz5p9awS3Xr/jhZnfaVi65j061Cji/Z1I
RRQuSHEzJrNtGiHq3GbliuJwxNnvgxcx7s91iZfkWyET4At8s+WpMuYM0SjCmLk4o7bD/qm/MLc/
ibmy0LuS41EKpsgCAQ0YZMm0rtObQ2ULi0r7g2lsJMKeIjTCLLhax8TTdmecmmWOleYSw8WZ8+lK
UjQDbkF95b2CeF//bUQn4Q9KZjqiCDffjnpk/zf3lKe9UK6lqF9lBwoCOnz1XG7fXEpHn6KfcwSo
mbkAcdlnO/xK5MXwFXnM9j1XAYlls1J0igrf2xuMB9W++qksM8z5Rhs1pHfuyYFJ0Jp/4p5D8wuw
dH9Y5KY4NDiULlhdUU7DZ3FNhejNC03KV0o5lWgPuc0Fku9I+98Kws1aASKWT2YfEwr2mkUNrhJr
zaje7knbkxjnVuoKsgqrmCPwyclTXACvD9VyHAwigUwudlr+LK+ZeqXKven2NgFg/CM0Zq1dwmHT
EuWw5JR8a3vKmgmAFajE2yIHB2Zl4u5E6GV+A+r+cYrwF1HkIA6EmmSpLnGAo8b4L+FBcSRgTWrS
8dXCBPbI5u12WahhMCwFleoHFNnh0/sfm4J3Ox4iBchivq46Fzkn+A7ntiXjsDDp5NZhsXN9vn7K
7lhX4K6CjE3uHQoekF02FOADzchAOHAuNfKW5pPlByzwSSsRQxzmd/oeVxvmso/MV4r9+lgyiiKV
pAAKHHP5EB8hPJiNR9tPOYLCtXP2JjoypdaiCsFmyW5cirNF8418zQcwF2u33hr5JeJjtmStQiOY
RzVrTq6bxmxyJzlFHXcl2VxnWLHr4BW7BzXBl7DyIt3UjHKrArlG6uo5+/fc6ybYxdqAFHiqE/76
TJifT4naGunYXnR39zWAyF3y0KNTZbhfFWwnlS7P+jhJS6aBwzsXB860Y7wKFVKrs7pbQLFke6YW
CWieE2aozuOOR+U4kJ2duBEKcZJwAHFegO3X9SGsADd6E/Cn9w4UjWt5cjF5jqeZFiw7f4tMzow3
FuQr7se3y/ZZdguDDu6HlA8vhoAXaDWxPFHUjYYgBLw5p8m3wz01KnYB5HYN+IseuUYWe10VKHXs
exmRGi65vPCzfMtZG5dR6d4e+3VvyXEaw0MX+yMDGSisR4Ou/D119rGL7tIaGgdHUq5VmKZOcYqG
0QRl/GcdQcDwWC4ybDHiP2rTQOcXEHxxHckAAue4hXjEfDl4Ah9tejph+/nWgdW55BtYWa5DFIuU
DODELhOaSeb93nDPP7nTPAOiw/VuoC58e1CZswaIE2wh8SyjPDseiOvE/oV5WD/UzvXelQYQUul/
1RPJ6v6dc8kwqjvBxoK3slDwr5OtJupb7grmvLpTmmZhGZAli1wbxOhY7FqqUb/GGpuUSHXuHrGD
6disfARoG47V+HfXh+ypmApgqE7uN/nHvhP+VFekymZ1sV4Y5H9h2b1FS3KFYW95TzSgncn068uO
BHAkCogehaCjl7NoG3G6qcGHL3nunuyH3GAZPxB6/7Sh4tvnsyR1xsyevC/AQ0aAklnmK/qhLdb+
lmGYor8CmBj84piSOgc1lTlnRqvvZJYQE12MxtGLUXwBHUceM/RJnTtfqzp0N2OJQlCXB0jnHN97
7cE1o18M3KPYH08sfaPDV0JW3L00A4gaDLg/07srz9bZGPkpRDQOZKFYQ5JD/joiLuDqQ4Lmqo6Y
RvDuaPoav6yP9m84Kpu4CwgVhqdLGad8/MNJXzy+iz10w5TzF+1LY3+4DASge8ZWXwki4Boqqy/8
gtx/40F8RHoequ9E2CIAYP44EXsqj0cBJ/pVs+B4L/8p8OJ9n5ZvsJBMvWiWkUj/KDXlOay8VyuG
U/Fsvvl195y66krdIeFdmstWGdZ0l9z+cKGRjR66sl2Dw0stNctGAnBXayl6Buma2jNwrEnf1drq
Jr1iCu3a82TT6Kf8AXCQns7eQzVXjV/ocfQMgXG/D7LmdE94zciCCp5RIJKAIgBrBjo0QAjVo4Pv
NgLVwF2GX5QlJwu6Py8HPE+wOz5AEEhcBj5JGX/inxsn+nHOkhiJdK9sPBi6ve1xRcqOFX2oRbiY
1mXrp6oYJe4KjyJZbi8Nnf4LGtL6E3ECpwPjkPhNxnOZxG95T3GDepE56gaXBNsZ04XpQ07PPEC8
pAKBIURlvMXQH03iC28Bpm3uN0xefd935ScXRhJQA1HF2JSEUE/K2j+lJWmf5pcWzYL9j/w5R7GX
ouc+MA8WOaFKSZHLNZR31PIZUFJdcvFmVOh7WAkZezn3d2BFZog62L2VBCOKKn38vPj+Bh6xylOi
JqHqYbD2ehuFtQZox1MmqWLxABZ4fA7EoueC2VjJ6or9OMtn79TV1iwlVcvYNCiC34vPIXE4kKx8
27ijHlaZHjIwITfYLdwQDb9ATcHKUQsIC1DLslrl/Npk7tFMfxbyu2JFblPg/NNru4C+S0ao+B1s
ABAZNQqKyqxekziJ9Plotx5O2a4/ouFHEgiG1WbOwX3li40hFCOpYlGFcnrgWswRvG9iV24gb8N0
130VxFZxLoN0VectvKU4/eqH8ENqqsopEDY6DfQQXO7tQpA4R2JI8UnbBdmZNvIMuRiq7gOEO+8r
sj39ahMJ8EThJ8QYa0A/BXRvR3WTgpbMVI5m8lOHQAVJbPFmQ0Dz0qhhbCSPSOnazQ5jURd+Iwxh
0kHWkjk2O+4tF0EmuG71Y9xgW5ALqeOW4vW30Ijr/R4ZhrXEehg8NJlx9aZWSVb7rKnYSlPUMPV4
O0v4h2Bd1vKRqCQD8Qu7zSDSQZAuPKIB21ft/STCWKlUFFxGG+txIJH+tyO+vnNm+Z9F4xaB5LlE
x4qGrlezLNSEim/60aNVyrmPCIf4xRaUAiXmvfU6M8BAhSNgeBonOKSiAX7YsSuj+I8kMm3QnWob
0RJBHnFmpeD/8GIUn0djTuer4sFFRr6PtAjK+2U2hBRroq38qEnYEgjcSxCt0FzOI5oYUO1KK+SE
GHhrA2MqGYhIQWnn06yQ9GVTYyvKjQMOqpNCXrVun2tTdT9rGOaNF+D7aO+6VYyJjnCcNG5UP73R
7hYwiKQfcY8on5Jm8TwdjPN4IHU3m0I8fH3f0CEa4AWIVUzD9ISc2x7K0LNNasDzQ0kIeGL7dCEs
T+CR+jcqBucXsuPSTjNvLpomAXr3xPInCu2UhkhyoaCZFyyfaCyNofaZBTUpc/CV6qREyZ9+BBK3
ZYECajx50BOeKwPBOI9YVyTPyyNjkZKI9nlt+BxXjzf6Wfrm0KeYuUmGzKOD1v6ZKFcpifzpyB02
KaO1mynzPNlCtpEa4YE4gdJw46YMb6OwVFs5Hb7o8H5e4A/aqSFObzrlCRL7/axJUVEh/gSzJIgB
rQIdCJTmBFhL6/6wBzUxK+uNwIOtdMCqBaKAxijrruxlEicXJMgK7ZZtWzUvsQuwEpHutMxMem1j
wBfp25ja4nlDbdv7gSek9PYyS46IWf7ueNrZpIJF1D60Plse+Wl59mi5CLKJvFX557UjTsMrIwOH
X+9QbJuIbPAznCfakaeGmmaET/qPX1VXKaEKP48X7hik4+igqllbW9g8I/jsIRSSTCNxfmFhKOyn
g4ky5Tjo2elm1N4a94nxlvj5jt//jc+v7VgnZQUQ58aPVntbkqS7+UdwuRoEHKkxo1fRJYJdT2lH
vy4pvw1KF2dnNwBsshJnvf/8jTwx+1RsbJ0hV6xXn1zrkGZE2ujm4/puYfrBhBCECPqJC66WKhWq
dvhqWK8fVSaeRbkIXBgN3YTpf3nsyJdYTh2W8+ThqOoTAoBNzlWKpzfeKb42RfDAvS01Diuby4Db
RN1zN95FSjDImBCMxzIqiV68U+kzC1T7Tm4OFNS9q8by7ucwCrkt3EgZ7DuJeUtz5lBEJzb3bR5i
OZ9pvY25koXtkyccV6wSsO9oSwDaCjo+VIWklv/Vyu9QeKDpnnxzZB1S5O4zWdCbppd68a2IfjDF
TmBUFVOxkoJETehDYPXrTimSaeVa7ffEdkeqw1pdoqTX6mS/MbgNozt/YU1p8tiE0brOP9ZebO7h
lb4WcoRpzQTdGL5eaGNCP+Ej0+g8QMMjGQUN+vUhDOLcNKHzp5fbgjldJ/6NsdYCEE2+R1xd0DMi
W/vOyZXrMhaCPWHV0hEraiD1JDVoOg2HERhA2UGqLT6MrhgTc3ygku6iCOwDSI096J261sPRq4bH
dtyl4/GR/KPHvk/KNoRu/bMr2ty1RGSW6ZHLU6yy+if1k2X8YtHfRjQtt3CTrR0RAV58xq3ePg1C
mCiS7SZfs1sVGGtztWqhKqqjHJrJRRkfK1G28dAwCk4etoVqQkZi6xV4Jb21JCqjiZMI3WtV1qgb
Tml4so7rxMoCCwsWsvBKupaMRbH0i1JBGnFBBsmsscfw63WNqAZpezrPj4zh58p9a8GrIvt+3jvK
b90f2lUBoYdCnp1+cY02pPGgjzdgR5vcW3Ppykq6Fr+FvQBGxaXwWr0I6WxO8H8hECpf9upBWu2M
BZCpUGPBMYQXiGq8tFpKui7quqXmjvLRN8O8rl5YzXrRKzliLMBOPx6uIjTLGMdkjfEnUJFk6Yg+
QZ6A+bwAO767wErTM2GiRTqD3jnPSY0UnRdovnGz/unqDffUZZt2YnT9XOOTru7aWzl7M/wXArvG
EGTGhVFrVu73zMqhNZAMIM0QP8wyFn28vpbqg5Uiv2/LDhEKqp45IIlSE2weJDLdI0kl84lLxltC
7ObqKacsPMP18vaADyTvz0sT80kBh4y/k5l2xkSHcx/YrKplQNpisrMYsClnx8cFSK+msK2rcOiy
t4rRpG/Y65SVbFvhs20eNhXQAtcT/1353BJCOc2Gwm4T8vHP17t3Xyo2Y0aSBORu35VM3u26jpgT
kKXK2gp/iFKTrsd5mXPtR/anNlA6wA3SAd5q/TZzlDGDcVZbgc/vmDcnKb6C621Jdpx4bwT5oGM0
3U82hYmBmnPiZRMxvBUnVFYOgUFznRq0PQPtpMAlYGahVyIfKjvgpDcWjYYpPdkm9s+RAdQpHpVb
URElS+IvDjTw6tozvifccJq8kZNmf8yE76aZUZ0/q2vh8c2yWRfknvb4FXRvnqEP2cpo40+pkQqm
qzMES2/pmNu6PfrJixCLpNk12CsII1H4evQrGGQKFpM4CKa0frSkAXHEobaTxE87s0o8+FYPFO8K
02c7tViyJVYjqcIswBmM3zCkoPl3xUb9sFE13oA7DSmytSEAxDnB7jh5/G6GmKuQkkgb1OOTLLSZ
KZJAy3PuWcq5Xz/j+pbYTufwZIH8Gyq6yGXjXw0xug+I+aBYMZQZoVmSpBYVK1w0ZobKuWTqjY8y
hDtIbdIk+e7PMwxg5e1tIpu/kp/PIQkrVgiLcamxgGAyih43UJ8I3akxnw/IfYghfibggkdsMIbr
o+z1o/C2GH/ugoLsUf9N4CRbNSHJKP3cjxMbpz7rgfIf2ViAOA15rBXSof/ASDa/UOgvjqq2AlMw
bBsmkMH8EabgzJcem4IBzWtrpBPh18/gKRtf7fb5jNtGNcq25PdlTKJH5sMUZtrQlOya5hWO6go/
wASfyXCpxnqVx6uvrvQFe9LHZYpjbRTgRC8zdB/nqH6nFNcOQNUNOeW8vmjmYcOAdaC93iYjMahr
l6oY+4LdNxg/+h4lNJut6m97mfJ/XjwxzwMJZDEirjX6zs+++rT5OF9HQ3XAYK0960xBWzsOCsdI
Z66DuR+ohpSeJAgjugw9jRIc+2WvSFtiMp0g/Sc0sXn766phKIOtP3ocKgT1uPSyaSxt1I4sBB1T
m3ZF4VHzyYsBgr4B5tuYsE0T3GKzacxO6bouq6KuzfxnOwXKIaE08iCi+l1Gq985bvIR40uLmNHV
YFMmBo+1m/heX1m9wIxqTBhws6o/U5Ac1DLrKns7mtaJDaOzBB3MBqnKMFtOkT/hEbIzmF8ogt5+
qbAK0fxtUgoMvmdbc7Hgo6+VG/a54/6M9KX6cJcPQysz+iFlFFHeKAaSkl81+FfrCzNfe9oIok/m
d58gK/d9CSwc4bTA2tdRrL2Ia6qiIQ4kjK//NfkcQvta6qMD/Vfh5Icv3Ag9mjxrz7AQgQQWcGfF
RB2QEBsYP0bjWYcAcaTHoWXJb/5NRn7u3rofjT957A36EeQ3miXPecoxoJEyiwao9CjgW7Rbko1y
2XyxF0PLbXJmcy0xczy4vM7+wEndUtDNQNCdxm7slTgSqEoOnRYmWQzjTuGpSa/rIDlCtgBFR+iN
DUukMlGj9TPvHfu9bW83BVVXSWgkLfZdffM0ohpwIQSN6454xz9XzCn49edjyDpiJ1WGkXgICkA6
+ZZqlK32Wd0MJ8J5uikypPbktjqokIteLewlV50q4sVA0pEWzmG3xyMj/rbKwPVRJRnuQkwwWuCx
x5dGy4h3F0ZfwNAAcy32j562p/Ii9775a8SGLlotx2U2uSZpuEQ7/m2IdDTTSXVkFzMW++AMA0hs
3ejQIx0k8Aa3m/bEjgXlkr/3alJF7u6CrMJ3hHOx30mpUL/vC76TG3xe7XQlH8rwNvD7AffSgxbB
uejsv0+E+84V3DHlEkp4qQuI+nj3IlJGpvMukPz3k5jNUAK+sYhYcypXb6/OWkJoC6POPu3yZOme
Erd8lpSHY/TR7W5ays41nplBZ1xlsbs8wjcQV11mAOTpbLdjbBgJ4788q5iRvrD6qp5Va1swQ8bc
XktVX/5sbVARAG6Twtd/GYmT0+w2dzwK+rOvFpCKuGJQ8Q6Zf0WkSaatsC/BS+mWqnQ19gxdWmep
GVWN/bkXgYmY+Aj2ChucSqbiW/E04OYvTaeRya4R2k8SNZT2j2SYp2MaynOVLC/WS0EIvhz5/EA3
uTgu6LhTPpqXeXQHjxlo1W2iLkBQzMy0ZZ0AUs/VU2VfKe5j726tTbPVfbvqbRdAZH3c1vrqrVwE
h1a5mKqACsvqI0JVG2Ao8JIY4AmCuxfN6lCC9nX7MP6ftBmP1lRrBRoj0NZn22LI6P3TNfVpu2Ap
2zL+lgqubJEab0zh9+45LX+MKzllgaAISjiX+PdbrhC/NQcXADzWLH31gxcDb00vRwiiEQr0RN3X
7IrKMZhbLx/Hivn744ufBiQYUw+jyHnEggNTxl1a/knPwZ3oS6iwH9IWfvOqsQdIHlRdz9JMvPBf
ENNWWhW8lsSkKZvjE9QOcTC0bFPuW1zBzRJHGMR78iJP7a5y7mwkUE5JnFZ8tcGq024VqWx6S+M3
Ede65QOXniM0PVDOww0NRsgVhKwoUP/3t/LJWrXv+T6wdqK5APyBmZvToZQYQYKOUBkO8ObP4GjL
E6zzuoKY8agof5jyJTo1VzfFLaOG1kr8PgviaoQ9LlEBNoT3A9LsamZ33QzgxGHylIjuT7yJ/n0a
6dRTngeRrefDprq1StKjz7AsALR1g3R0xhvK0pzmHgT+Ix/ig0XTU7G5eJea4jjUdmTzu3SgMZsg
u3ZRrHs6ONzwg2Vca44rX6b/M5acCuyWzqmWC1DbskXF4Qx0I+SHddtwgzqFDhQOORClLuYvRT2L
UD3lbmWxl8ezS1GXAhflVqJK5Q8MIO9LIKqC24ij4NU0/81LSviClOwzcgzTZaN0hw+cofVsZU8n
ANEHpkTpfnWDxr1cDtVoa0g3vkYn6RZwzA0czMrEnkRNj3G9vewL5qO46ZLPiieGOA7V7KRBb/Yo
umJGKomB43zlNZo0IApB6DB6sat7AOoQjzYAew7iLCTvdkThhdQmy0YTVIdgM6aez6f0If8BK8y5
Sufjk+XyDD3z5+7YrIgd49s4XDbbOszVF7VE3ARK/cE6fP9gF340h7DkicYls/f4G+Tjr8q0zt6b
2gSxGl3VfV3HXocG+qR290gNAXv9l1ioprvBOPPImbtBax2rUxr1t55Ku1N+tJee2nmnD+FP77e8
IzcMDmTrqayx0W50ZAfhXSXd7n0C9FWFVWn8RyPv+fATT35LoWMCkOE5W+AzrryThLEEealL6rr8
rw74Y8AVmzgQ7AsJcnoctOfIgytdj8f94ZjwvIXFHcxZagDd+k+17zb1t/1SBcghmIv2rCEeRoxa
hS+vdT7tGKgaYxWKkTMRzvmQYeP4Whp3UWfAkRRg/YiqMT/MhXhsFc2ebtF+Oq1sKT7IRCOH9gt2
w6OgnFdkKTKsZ0iCAoX0Uc8atjNXidw+Un4IzYn1mKncOe5vC3aMlkk3z23NNtyttn+nzDqomTvZ
kpyFMFYfU9Mnp9ybFVrkafRsPWffbRd4925F0NUfsgOzFI66DXq3VBnVqASvYhoG1RKTTJ7hCmzr
lNKiUBG+P+hAx9UMNqMczIzxN76Nox33mfYznaWWd9wIqQPvzJjHTu7DngoRenHBr0/++6gdpTBY
D3u6wJLcMYB6Nm6Lfu/IOFjFtkT98ivromkCSCQQna2mqCoPwAmv+FJt+hQ/Km+8wiC+OB4147zh
rq8t/RWQAGWOizjFOJEidQqLXACeI3jZpoOpbVaSXr07BhbN3ohzl8fEq77aXfYzPv+Vm4STh5WE
e3HyA7wOGvjKD+vL9L6wKWXCeDHJ+6bVQSxs4OwasHB6kacPHy1RNWqJMakDCu42+PT2M1VtI7Ov
tJtnKkWt9c54HAl10iukfXlwGJ7d1A+9Vqh6z3U8MKo1rXvQlpG0+chbLljxcBKEYOum0u6FxHoH
w86EdLFiqIT5CLc6ium1gY6vb9WQq6tzSJ61ZMUxSG7LxyIr3iAH4HGWBu5qCUrWFKj7I8bM6esP
hPKN7+XrpK5sITGZeMBlPPf+HNX2+x5Xe1x0aWm4MzObFQ9mNQ6+I7XBj/yPsLdiK1oF+vrLp/f0
r9in9PKzy0S9aWdIboo8J54ur08iLm7B6gz2YoJKB0sJi/ITssq53T4uoW/yuKMK5bxP09894bPL
MKbhGQaoRKMYC8dA1suX/VYCZ3xogh/hhf618zlkTvEdALR2BpsvQiEosBqM97G3FObR3FRNhxvE
Jbo4lP3VP3hSpWR7EdGUbtvwiyOIjuLGpQ6qBX10wZMUgIIMvc2fF9HPcHRMIn8ENmzZ9ypVkuU5
VCXmyA+NRU0wSVYuKFTwVlfxWBkQXFkQbW25hdMVQ6LJ/axXLkoQ7T7VjWUAfJQMaudjW9f4FFQX
wi4CzXOvZVgQFahKNB8VlHSrpHE7XTSw+9mHeHTADMs2CfZd4SeV0fo85+dpsG0dnY1RjaMzkas9
8FhqLfC/jWCQTRNsxNW6SV6c+ZPA6GuqxaL2wWDdeVht026FyRJxmvbTu/Kz8SROnbwSEwmGSuUI
HN9thVk3XjvAXtkgoqt7xG+PYdrCbTCC0xvCJWQWDjdBGlBEbx1UDQ6gXf9dGSTJyq8mqGXQhyx/
URP670BBcNL/C3OfQjy/Nsm3E/le490fUY5Jk7VctNOlhsl98lPzomBFPBI7JkoP8TyDQ914AsyP
1wX/0sONBtz/oyn69itYu+SsPwdpmXe4YTBCo4T7J2nY/k1yuL0RVGpqoEZF/N2wbnJTGh0+EDu6
tu0UTElIRwktCoehB8d5d64zCRNvgc8OjlLDrVCKfBApFzP7Z2oXV8/kCknj8x9h8dIxKHrziTsy
3ELH2HaZkAUKk74Q0TGu1ckD6W19uehcBSjUyR0zUX2VWd7mzCG6eZuRWLsgVkQqlWtHWxEUwTVT
ZK5jW8IN8WexQguZF5IQ/EIHRkUzoUmxEDKv/hcegxvpsXRVuujSTgra+j3splYJuGN1Ybe8g3J8
Y/RszjSdc/tkpXl3Y1b2hY4oiqNqXuf54YldncQ1/UBhEzGzVOK9kzOuQA95IGaKUUAcojMOwM5R
UJgsk9++kbSU3v8weimD5cZyrEWbRDwsz/SfDkm3AFTKJu/L8khL4J4Sxy7a0uK5gaQCCR0EO+zp
Kbg+SKlBRDFOH0sGtwuk1V67ed/0xs27P2zLU0VaLj0kn8p+Ugqn7n+AlWp6Di9J7cG8zNpsU3QE
kRziFedy1UbeJn47XvN7J7q46Poinvq6KowRcGlpANSX1z8IC1sypRYKLT9p/AOjzgWcaY4yTAlp
2fzHOzWDB1N6CHKoESvY0KrpiX1zw/+SHj6PpJAoZz9sHn9cuQU6y0IjdOGQ6+k+v07wegFeJo/K
hLpKtb3OP6MoerI67B4Kl3s00JGxkQTUidoVAyhuOCWAE9psnP+5F0Lnu/G9680gk6BauVBlsRZw
oCbY+tTtAZnTRLc2e+ddpuJ+bxe1krvj8i0NQ/taHjxm2pH69FeOv4PlzljUrcQXPa28730QrdlD
2zWzoEM7YvEgP8QtjjuEHTnmvRKr2TkCaubaXfcdOQNXd9PHSQHVBjNl4dEmNpBaHUWNpyyURLOx
g7mX8O/VyBJKKckjShZYDscp+6lzeLMMpOUq/qWBD66/u9m9WtgMqyRzhctgSFrsMYZ9EyF3XQaT
xDpsN8brvYLj61I9DcXHsC+uuxO2lVkxuW4HRSk/ca0OeRPqatSaMhlcU5wBv7tXpa0re9lFEm1H
jW4kTspqGqdtJXxtBlqIwU5JQCIX5affpbet2Iv3DSuZne3mV59ITR0QY8odb8mOYMF5zQ7aDw1B
uik4mqhNE/r9O1mt6gJnqQYD9m7WqBiDlmmF/RDbgx4BTKeXzkOML6wf1NUM5kxhiFT7SfxIJtIw
3bgPCFfxK4r0R7e8Y5k8f0DXeSimky3y81LzsvV+rPaPqqfisSppW8AGg4gW1OPGkPtcIGxazXl7
FCqFFnA2FpqRXHf0+VjbD7OMVSkCeStHf7BnYyv9eHsZG8ZorksPlBj601OMjKGGtkEJ3mFg03Wv
ABwv847UH599TUghvkH6hC3K+YdAkj+AG8MQ56uPYat+o+Uw7UHAdjMzxBSbxLmrrmhe6HRD5lsG
one5/+2HPBMQyEOyLreAH2RWfbZOaxyxUo+S18D4cxuf/XEENJdSSjhVepdFCXIrhCrHSrBXSPzX
Pg8ZIJx/VwxC+NYUFbuIsDc/jfkl2NBFaAfPD9Ie7dErm0cyt56qs97x/EefVJVbOkAyFA/e5wCg
ygOzU9FjMbHBWrFfGX+Hb04oB/JgDid7hlx48sdTsNKmjLs96DYpt0XR2JKqMBE7iyPIJDhN7WjS
yj2h6IMXM84JAtasarZ+L/O5WBmOW03LUuArXOtPiPN6XYtUy4auVyxF1NYc45r5ymkZjnjxdQ/J
YmeqvhGZUlSYiXLr52L/lyo/RdiI92E0zp+bOgPuUpM2Xf+ru1Y2b2fBHTHWJ2OhaQCuz1tUNbUv
0qGEQJTZE/8F5pcHxANNOq9VPgVhbwL3hVKTlFaPJkg60wVv2jXMj46EGZndl/fuDYKLFwKbko9+
705KPL/HPd9OZOdz27OZjxWN63CilO/VgwfzoWVP7yxphVy7YOXFdpkY5JlZiRAUeVFbc2zZEglo
zED7aOyC5CJUk7yAFA9TqRc935LKvuwAB8K7uhsjCKVxU/XdSaYjCjP/HHMfphUZHt5GpixHfVPq
54BnJ3ieby6Nl4sgvXbSg2SYeK+Q0RA7r5Yum472czOn0at7qyRis/qni/8gxz5/6EdOHlUq+sAw
HZrXkpxOrWM/dzUXi3pGVFjNilZXohTIGkBELhVL9OGIQiFhJzs14G3I9YUi7jBPV2GKJTJ0MfnH
CdZYQx8h5XIpMn0YiVx+K/Rk+gsGeiBF70Weablq7IGsvE67CxSxxypwRwWE2zcm2fObcXnclJMm
j6LyIuSLttLfJellEEic9ZbT8iZCLCivbbXub1B3enV5/EZt7v3o7Pt7mhKqhdbBpzUupwkgl9wD
ZniuiaPBUhpuYauHivus1CsJbThMM5fjyVFzfsK+4xA3RAfibhJD9SHK8ond1UXOKhYIVHnlIAM0
SJ2vz1C0lj6+Z9YERHjEjiDgvXCAiRmiVR6G6VmnKtXHuu7Ca8KMAn6bCDeHjl+MD1NrLvL1oTCD
G1PNNsDNKOzQYMxFQuFJ7gA7gOadXwiemrVPR90V7J1YvQOcqKYwZRH+f8miREl1+GfnKstbIXW+
GmYoh7tELLSGF+kBTvpPNZvqOInBYTY9soCmNmN3SqFMph/C4te1wi3m4iqRzQ0Mr6CIh9EseUvM
ckfjeskvUcWvdT8CIARPpGjgXCxY/jTgGytIpc3QyWbOdT3t+YAyPj4PpYsWAbBsdWAdhAT2HusM
wj55/jYCSU+mEn8cl86DlzPi1oGK4KBXA1PE2HtFb9iUJR49wUWE1Fz7q9L4QmcNnURri15Zwgug
MAW/kwoVkluGjHyqoKuWK4eVM+xo6VM3ljwnkS01XcyOzTJ9HygGIPUmiJ28p7jmA8i734Ot4dXR
JMcL60FPEf1OJzZYOw1i3SaENV57AAk2BSH4vjbPG/emoVUIhxnttZROUL/mI/xevyV1FtsyozGj
yTOnW9vafIVJQmkZwt2kn0+v/cTIu1wceMa0reVzS1uQoRxzzc5cktkqz3cxc7LUqmJTABxdSRYz
/UOnchJc89XBSIEfoXo4fuCSlgFkjbUdLjPFV3L95/dy+4oCyTnpzgKaTA3ROpkzCe44TR3yfRzQ
q2adNtbY1yrV8S0TOrhEAW0U6OA46jl1Zg/Km59vC61DTUcrK72YL3HeOaue3X+0twq3HEqn9PXC
x5OgralG9T3vuUzPGSkiQW/gspRKKN2LwFitNTh28+bUsCodjQAwoCD03Q0Be2XTSfA6J049goDc
ATD4x4rZLLXCfwNy9Q6x68Hp9OM4DOFbWmdMHEbjjd3XvPiNUJumvWkDlzjfGFMznyUEywdX+otV
KwuuMtu22lXk1dGPuvT5abQGlMZswiyv1XBjjhg4jfCgIrYDg1wD5LiDSdKAm9sHX8zAY+a3eWC/
eXYl+J0PbohcCw2EDgpWmQjtd76x0x1YJPzlv4ye2JnqKAY07GAZaSLzqNbrshAdCR/ojONRGgr/
RSdOERUWpq9rE2ffra1/T3ek7WNh8yho1PHLTguAfajl5bgYqhErttxQMGROKoAfnAd2i7o8YHtE
GofY4KSTrTSTB/pEh7K/FdI1lGkpumfa/Kt1wN1/Js8yYLjPVEAbYt6ODscoZagdUCOa7Qzyr6Fw
3YrQWJZj7eY465F+r1iwOwgdwIWNXZ2/zW1srSlKKZrNFLh/bRFNU3w2ta9reRQqDsxWH829IznV
XS/lPxyZOWYwaVmL4YxJVzqHhjkblBkSoPYsWuuBRWjtsmXDVANReis0NHfQI4WxSKXsCCk5W/lo
glq54U01S6lLM8yvTt4H5qaqYCJgI5owlWxf6v3ReiGU3C7Zi2RUNNeinEWKIficJeBaGxRdYS3Q
xnwv1Pz0j2BOhDOnNAhvLG3p8KrluTCOLDJvXYD9xWOvPKb9CmXEDUfG6e1XYur784u/WSOmpg7x
jV40aHPzWxCZZYXLrAzNDYPYYvsooWNG1etv9kV/qNvFjtMlfg9uWJjNHYde3kXc8W9Y7Z1ZQFD8
kvgjr151OFvO3MXHsK2R5PMrcJplc6wFN0l8wEV5rYX/N1c+cRmz0HaiTGk/k1RsDqPDbykiDXUO
FHLKrsC1CudIKiUiPzkojCy33RHwhwJtOF7YNPuMpgTAC7rJtUdfqG0PPcs/le3w5SmxNqeOZZGL
+g6O9HDhu6DMvoSODBEt0plNNvAHcaB4xJH3XTPKQGEYntdNL4c93zryAwlul6fzeA7i6sXBuZ1X
nSCQwtBJwHgJr/tgOWZTAhgIjMI9f0A5FlthNJkcHv8NBEuCcqHzCZPM1A0BtBP/PHqmw1pxZan0
XaNKbJ+ieXLXjechxNFPU8qRXM1zxxQDJlGqf9IdmKR5GwSKdHwStV1a0uP1mRjqdRMQ6C5sfMRr
F+KRc0nGlcPClL3I5OlaJKIU1r02CEhtMvH/tqR8Xl8J2TFwFKeGv+HTumABsaUYmDdF03SqaHjd
3vsl5If7MCebo93PTB8of722leVaKPxU09So9oTDMf/GEJpQ8Zkf/gI7LXnKIKanNiTpc2vDLT0S
0J8zE9qrIt973+G8IUpuXzppaqAqr9BguMDYA7jCAt6ys+taQwpsPKor0ny2uoxXXD9wkgnTTgf+
HkwyTIZKowg1Y40cJDy8y0p+ruMQdNxTpWbZ89IFzJ6SedGlN3zxA89i9WPa7/1N7JbluRff2wxR
Jl6UfjeqSCVO3vrqHfQxNYZUMmkkt/3hsOVkaQanmXUJC+cPr5rf8vLE8nMyzBEZXG3ZTR5/GWrA
bv4XVixwtEi+PHHof4HRdDXKZWInuY+BIOTEsrVgRFfpC7UOQXMEVQ0/5dBvpRmHGEXVSHbl67HU
N5I30Ca4A6dCLK8w2snugOqGpwXwc1D1vDpOcTjOu0QQf2j84Qre6lEZmQB4toviA35CuoPCTI7F
3Oh8KKtn6Eg1NNk4pmz0f0BlrZQqualAlrChufhi3LkxpqZJAx1xfIVPg2kx1D6/4FVW8j0sj3ZU
rFvDhT8LidPTm5fN4aTsEScdoQCqn2ukzzV5WVpRWXm5D5KPwR4xgmKPCkoi0SqxgzNbPd7L1YF7
qd1pP7hLCOS1h+reJtJqSvBtsAbMqGDZaAcHH5byYDceSm2jgF3QVDz+78JAMigoUM5i8FPfc66G
L7CHqYLzYZ9zpe7g0J3DdymnSLiXscvDG3rEWM+HTLBeMzf6ZBHWINfdJfKigERnSPx6Pdyhq9mB
Dd4pALMT3xrVjHunHgB0u/0O33nK1a7926z7LEZAryymaudJ9Zrcj24DBPOwfoexW7XVDviKRlzC
D5JzLKJ2ZfrgA/MAvOHup5qb6F2EzRa9uP1TqJgGydfg3/g9XDA7F+f0lneovFJ51IPBkBifXpiy
RBmiqg8SFtlTHUofeeMttff8do0KFGC8AhyvcaGW1Xu04PO/CIx8c7H9Ux3H8bZpk9Yx61DwnQrH
5B/n9QIadVViLRBq0Wh38ibFRxwzL36IOBlgvghtdOn/BwfEFziu5AdgUL2hESdR81WGxGQOauXB
wJcynsArtEWJhHf0F9cyjwF+itxXJKBOUZfpCkI4lXpNsk/tzahXwFX8xkezQeUAYLrM+k0HjzKB
BbrzTIOHGSUo0RZkcW1dIldkH1jWEL95gvaOClE3JoqCY71o0s7sdzRchWlZEwwkWxDfZgPI3CjC
6VeET6yzAhZrFJb6o06+xVIECoBkLidQuDdRu/kq/AkX2b8pT/ntfUShlBhG9IHApa5e4cygPdWy
5fzlUn1ibDFmUvKT/m942VBZvevJmMPapA2TEjw0kZcu51bELTWOWg/Pqdz3ag9txwIIAfc5hDQb
NhnOpWGdL6T1vmWoXCZXl4R7Rr9uKSW7Y3a8gQL6VATqf1M4Lj0n0yzUMUdXweaL8eTp5XG4ow3o
mfQQ/Z39saZCv/stnIE36mMJM+hE7/MYtsnosMfNLvo/W78V4A7ZP9frlz7NgfRxm7/spa6CgFIT
/ma1MDdw/aWEK+I8JNO43PWsWf00zfeknaHkdzps4LYxaD36iTU9XF0OftrghI2NONNVpeqfEkPV
RQ2m8evEFXoQciGkWgzAcWfTVxYVD5Pd6mHt+CF1NLRWpcc82dUQ/LI2XMlAhnzNNs5Ibv2oFxT5
x4QyRUzR2TkSGzzemVk5NxBl12fq8aLdBhbYG+0NxbiPb3rrJlChfjztRzy6ZfexnZAxZEBDilTW
CnKbrkCXMgShEoxK9xUF3J9lZBU6q4hZcE3vt1WNAQvRwslNhd2nzBLetkXYTEZtAY2sEhcF1+Pj
XivUEDjiryP4fnhGU3K7pngGpNgq/H4UwWJZaPmOlT751ZGE96f4CuNuWlNKkWzWVgmnv+scbqOX
bjg+heKknjop4QYkDPx629mVm6fUSSzyU4K/hrpPQvIj0JGEumHRi52YgJB3cr3tEiaoQZEzzFS/
wkk21VyrXzlzO5u5UtQqorSt48NTVRWj7GFIvHPsUMfGDzIGeOV0C/hh1lCvr5F5mkdfmUTz+KJi
Cij8EAaUIiphxi8j1JGSJKb6MBerJLqViybFtP1lGrf7bW1tBYeuK/kES6mcfcvaSmFPjPz7dwDh
0z0aTqXuW/2H5J8OQ+qp37tr7gEm4Fu72DFyqYRS6bI/YJO8sJ24Ky0o2c3R0rvB6zyo/9fmDRKN
LpVH9bNVUsHNjH6twLOEi3ejcgQL0OJ9dZrEbtYNUfY+njuasA8/TmOZL+2TtAnCHeXc0UCkX/yN
GrF5WKXLEjqKlZZBLL8ztEsnu7boo9CR8yZ2jrxIn7z+UvRVS/LYBTPKCSDmTaPkc0ukJ0dAC70N
BZnKZl2K9b0hjQl1TTP/puk+TnKvqrZFc6rckZRu84QGvekTnnk12WP1oVAi5BG8z9Mb/VJR582s
DtDHPD5iy8AvaBm16A7yjmEUmRKXz145lil7rwbAO6BmytciZeIlxx5TPN6Luoxd1JjEIauc98PV
VVphxMsZgYtRC//QThshkcyHff5VaHZUWkNxxnAp74S1eBD57lUs1ESY0mBhz/VITbEgNCcmwhq5
1iJO/F9VNGYncMqG2vKgjSzmpbgeyzWFbh4WrxWYpBuqyRA6+lqOFKxlf3rr35Yf1A7eChYuqDLO
94OSFG8d1X6ScAPewS0nEN8RFxxY+6AGbQcR1G/LEoTmmtR7jYEhwi1zx8d6fwwSb8fVB7HbzIpV
gLhr+2buFhsf9hgglQG9OCINgWTt0TjG2IkkinhiCLUcRXTcKnqMbA5PDE6wN07HT+sqQI+kQvNN
jDH24WsuemwNU66327cleNADOwrE0jP2xeNPA9lkBhLaY8BJ1aivwYCn2NxkcTV1SSHFq1B02ySU
YVeI34IoAW0hZpWTIuGzZyUIrVS+EXfon3x1egBy8oQ/LqNeMSw8HAqb5/MFp95KuttL8Ppt1Xtn
YVntmnr0SI41nGbOriXpuTwR0957rYmPaWpqYlubQPpWK7ZKszjdukyul1T5VWPM0XP4ogounLs+
2mqFeJNtoqpFcyGSY8mzUf3PdcdVhEB8kxvXS1XA/w4GNb5UoQwMVLfvUezO6F7i7RZhYT/wD5m1
Lu8SO4T62gg5XetLGe6/n36R1njDwM3rYgsUKi4zrBzHrtANrDo1i36Jfns+Xa6O+vIa9qYPZqKx
tQ1HG5Xjo4s8s+YF7KwrL+ymZQ0GVmBh/yrFLHhSjalkL4ntfeI3MfOgGHHKbjMkBU2iJKbKdxPk
FhOpAcFz8B/JPlWP3F7oAORhoyRv24alH7CuCyY8LeZ5m3Rf2gHlRLMGfIZTJQlp1yAJrQy+FUe2
TziOu06j+0zOsz4Z2rTXSiiZbEqz0W9jm7Giyy5CwLdsoysUSRn089mJ8XjfqGcXlLEnnbFaRjaS
1ldwLgXaXG2VkS1xMX1NFb7Nk9z387xClwFJzwRNeEDrrpREBmnS3Ud5xa6Jrb6hZ1HVdvQCO8j1
3BR/Vvl4DIQLB/9nxNvo+QSIWM3IlIkscgJ3Zsfv7o7NoLwowJ30OkSBWfkl9iCviUdrRZ0tJ+Dh
ObQIvOj5Pk2TL+WEUEhxkXr5wKbjOQ8a7q5tcjtk+cr69QvjhnCY7MV6VWKL1OnDHk9HLjGZXBdw
GN0/yNPXqQrQaypXGWG7Cl+4t2t8PTWZWJsEXDKYiOA+Lo9H2DY+xbmBUUCtO4Z4pSIGh3ZfA2eX
vn0ZQYGSLaxYe93r+FfjOEt61AfNUDCS3k9uYSAzmQPA71EImIb6E7eNJchUWEr2ceF0au5eZHqe
fXUKigQpP5W3z1lOETIBrcC7rQkvyBRfJw7wgT/xo+zQSY7xKMVq0qs1Kg8hi/rnwf0mePOX3PiE
aqD6ASgeP/Ez2l0HrWkRcuKxAUV6BGK9xIkrE+gO8s627XKkKwAxFkM0BYfMqxvc+Yf2/N4SqEyw
avcPsa4HSxtk3/ZDX7dglVnCO6jg1X94gkeUGuF1DntBx+lyOHg+pk6d1YkuUnfIEANlP7iw1TtV
jqZd+JuAIiAMlstbS2aTyHzIhNnz1vN0x3w6V3KywqnSzvQLneIY+nUx235txww7p22fojBceGCG
RhJI/LBWKYhEMhqvX1iQmOU11L97lKtePCKXqHJaWs28IfO4Asq6BvUWOWFsrJTDufrhHdDuRutp
xg50CnXm6viK6DtWO5UG6VZao1F1ZwjI1nF1jiAx6okytwCQCeNz91bNoc5ZGHSMI8XHTY2ZDFN1
2/O0J9v1oW0sWZgkDu6z+/Q//I++XK2iqP1j/Qx38IRfagib0lnsHLxXlUGFzlr/Nr6BGHsyoHxy
weqkXyzmfClftoXROY1z1Bi10cg9ELytoWlPZVqoQHFHZakzGlZoBgJJ8BqC8xG/3M4YEiCy+Knh
f8J9fJUxnfdrTGiaiS3ot0plqkcSE760DjWJHheNn9J1GkbPVlGZODiJgMfsZiyNvTDzRNxaupcd
CtU2Gd+sZ1hrhtMyQS0SRdeFofY/rONxCdmif2LavusnfhduwsxYSSkKTUoG4cqA70EtuYw2F1xn
FQO86W6wtpKRCP64L2KOCJ1rM/gO0f7fNEG72Q1O0S5Kj5z6cKo/HyWRvs8WRu7H7RwQ1gIkm1O9
pt+3K6smUzsPdD0P+raCVrl34j/lwI7ZYZdbiQ18UfqjlFUkcrVzBn9Xr7363NOXeJOSLhiszpFa
a4czw2a4ua0ZO4jCR9RPNSS1Ya92uWZgJ0RJVa0nqvoSK+cWysE0vutvXAb7O/FDkG7P2EDTXXj9
gQpt86+QsLjxAC3Jxonek7dB3hJG0vSKvtWYge2wT6Fxhyl0cYps1IUgHlFs41C7nSNIYt+hVNhb
l+og6xLZhZ9lt7S+SHQbZYunzbgwbVoJ+YmZpeBvbMQDmJTptH8jhDGBpT1rDziTNYAnf3RSA5yq
sypQRJlplmVVNzzP+yiUGMEPj8wXKK+sgwym0Y1RX7z3n1zTVi0r1l7IYEss9qbEACODAfQAyQGy
9hgPGKTsearvk1UINen65385BRGZdr8y8w48NlBTKKhsZXOYu0fyd1KCNAlH/kjxJPkeX+qOi6a9
sp2bDfD0mLlivipG+MlNi6VVIs0+knC2ji75srF3IHLtB6gtE8gLJUwj8CXKGW+YEW7R7K6C1pQ4
2ItuScN4dR87Shldg1/BonB89YltVJF5pgxxOlvgmMIyBeSl2BGABew1/bR4QBhD7PfAK3C1bmkW
mYFIk+RpXbWKocRCnEmB8mIxOAR4YVViuOt6jDzNWIBqaYDcvkeUJKmD440WOXxihq5HIZVB7cx9
fBiLj04QSf916e9tTxWHN60dtU/dD54Wv/v3BBAnQ1oLRHJTOfX4/DWW3o+F9vmLzNoDqPREsMed
OpTHUZ0i3gpxEMJhrXekVi0Nu/3TwFUGllazG+/1VdnW7508smWIIEMEY3dWEymxKRcaLYZZ7Q3/
27CxAptJnygZbk2hTUYh5clQHOXMRxuwG+UYeImQxCatoV+TVRYzXFNCzdaHiaH1ba7RH/vTdkkq
6uj0j5BU7BjfU1VpRLELDoRVyX58B+/bBUdqDtIhX7J2Df4XqJaMqueBkxL3bXPQbBLctRIIgpP8
85bGdAJw+P1BjJNHwNRnZmK1g5ai7D9ND+bNhHm+jfoLReIEojsEZgRCtQDWYFrigaOwFkVeoBQr
GShtl7yok9UXaMmNxqzhb6+ku+HucpXgOcCf44BiMoe+x73uubuYx7VQ/udeqn/1x2zc6Rd6vwnr
noA3J1WfulHwvoVONMRKi7iBUfUzQl8SAXwh01AbpNGv0hTumplda0TWLQk3QF7YUedVAAqYFP+v
/SIFRZSVdGSHGNYF/IS4ScigaWBC5UyAmG9PN7CpSbCzQ+5HVQz5acu1yPF2XLOd55wRot5QnWpH
MPWxEFJEjEGzQQf4gwz4wyyziDTP+MiJ4/nLz3cKRRy31hw4gS9vXs/+WvjM3xOSMRlmN5nIByMc
BtASrwiWJGKYW1Yf5b0aT1PdEBZqyLbtIsq9QB6ibze9fa5/e/NBHZHRiz/QiAa7y5LuF1FV3juB
O4InfMEXBhDzOFIvmw3wUqM6bqj5o1MyVDNj50sEjgxjlFrVnSZNjDx6UPv3RwTqECdOM5m62MOp
9Zk4W8WqQB/zwqseja9oEJOFg3Ek9ChQw3m+QqDO70zqepP6ebkVtY8sanRdkNPbWvOjD9r7YKed
q4GgNqUFBAwGkWrthkYhkWqc+QRupR/8QPVfrEbrS7lmN6lpOzLKMqGCYY8QTHCMcj5ZJWvBbk1P
e3RA8T24v0hb5HtRniYc8yTr6Xg+HRaVcJqHnCHVw9/p8hUNp8PkzudZV+2yluSia7WMko4NrU3c
bbz3CdGaZkmLIUXNxCtUd5/dm0Tail7KLpXI+8AQP2Dc7gKNkwQu5ktL3FzrdwDKtVldolIHICMr
Rpi/xN2TEZq8MiBQvmYVRkG0giQwfWyNVFy6dHam+Licc85KSOFd62NwUfCTCbS1b5to1EibGmzd
iHofSxnV2GQ5kg0dtQH0UczkKsm5lH9fE2DFBQrtNC+7edsjUihHhFNBdwWBUtd3teZh1ApkFLkL
AKWAEFfaY9edpCB4IMKJnytiEJ70CBY7eqGk8J4793JN6wK9oPj6j/BWxL7WgsOoI3eUE7EUjuoQ
NrZv1nkD01CFRxpU/GeRS0Ujx9vx+fdrrXl95BgfSfNNc9F7Kvk0Ndwh6dNspLwqlauSNo2PiKeH
khbq9vdeawUyzTJqM8Mklzc3y3JjcPGycv6jbXiYgv/tZikXl8eIrepEU/NpDlxGfe3RNCApvY82
C7Ih8m5+sYGL8mgdDXe+URF9GmelywQBn/2B1bu1F/n0RaeiQZa0/XQRabd5Rli59vuKcN2YZJks
guya8dDx2LTdAAlUnDGS0YwoH2ak4k5vtjQNfDI/a3a9grNsCXRijKK0UDkooWpgcc4Yf1YWc99r
Lx7xqViqhaUpHDdeJwu3hlSE71PQ5pkckk1glmTAv2s1MbgUASmw0eaYZre3i3sVCI3D9d7pB8+B
CIJbTL9GAgrRTxV90HbBeAizY3HULLU449anqQ+/ZkLAjQdrX4V/y6SPjwRhnpFEJ46x6atfjQjy
yFYPksVLTO4LX3XWH2XHJB7u0swWJa69g83Akqnxi/IM1IBkY1U+0NtsJmW7r8pgv+toR/NfGrEJ
qQeezStX07QRVG+voPnhO/uQiLsWbf8hX7Xj9mCkUJ37noPhjdDjIjT9Kle/ATn5O8wu9+PgaP7S
CBIcTZsMn2gm0kk6qPUXoIoWTqhyejDkqgz+eV5NSmXAb2S3APjaLoy6bvYILBsKT8yHRzSd3KPE
2ZMjkEyOM0EYhDlLOkV7/qIE0zjyrtzVBrnjpyjjTEwT3OQMFjXJKlagEgM37096dK9bEGtstKBw
djucQMH+f8HdAECIcqicQdzCfhPI6CErdrqUfvQ2U5WtdtXVlRW0rgtbm1JimMAPUbEelE1f0hdL
NF/XrQjchsRk++TPyEcsmqOXMjJfB6O0T6dPajsm7Uxtcn5r3L/qVTRZlCf/NqvoPg7FWI0lWF9O
1OJTK35vr4f/kv3B/1KYeHU1X92j2GIbEuVu2gmCcJNn2obU9SczUwUtiMlGhIVuKWFpbL+g/soE
HXySy7UdUXDxYsfmaI4mZ3cXta3Tp7xbNWbMFfCm8FkDdkSv+xZ/TfBsj+2g36keQu/VcN6GW2U3
mdnrsGoZT9e0re6Eqd3l14mgiLsTaqj8Pw2tr3ExFSN4PRzxMrMYU4QdjexrcNO20ln9xLvfzMdx
0f9AX7Gp7atVXYxiDZIPtvRDm5FzzcEFT9MKd/VsIoabEqSTyXnDVaqVeJJ/mjyMb2I+hX0xzI9g
1j2fdzIlBcAQ7BbrXgsk0K+UWYWuSgeG4lI4jIzdk2pjo+hoXrfd8lvS412GInt/H8WX0wAuLYdY
yVm6hv6c+kuMYiiG7ZuIvlbvnMRL4N3Ac7l4NdUjLae4ox9ezc5YtnN2furB/JdSZfuGuwuVncxp
6NpkhFhWX1NoLGqzMQxq9xBxgh9GqRO4eGFa3cGtiuDV51Ps391pyyC/PMRlnOiyqUQy3dxBdKu6
DT1nVgRB4r+HNooZ1XmHvsUqhTswVsKr5ZbYrBf//at9DMn/8gXxCucHnNu6emIbu8XymZtU8ZPD
C+tuxAVMBAxbWH2ZMWBiyvL0eQp3fkYbZOnjaI80f2nzq3Zd0rO74D1dF7z7cNWQ3vjXYyxtAI2D
4xRi2NsDsqp6u6SXCmti9GhYBon0BHvl+XmhwnUSVvgttsiyhhibsdpDrCZP/ncFW9kp6vS1olW6
DTz4BCSMPIsMYGExBZ3nHXgBYxFLd96G5fatUq59bUP9h9UHLbTKVKZ62EWWPDaeKSVo5KbDwZVo
st0esJEDWSFeDbOcszAPPYy6/U2efvf1jXJ4CABmzTxC0/HHdhaDVJfzImmNeGqo+o0rqA4Qx5T3
K0+WSowmGfxoBVbee1+roFGqbDBtWg2IV8t5TVgqjSO3CSD1rMDB2zn4TyZOC9A4wq/z6p0qZ3Jy
uj+hD0kyMCGAytejwNv0t6NQ6dm4Mn8T5y9O62WbMPKtexDY1g9Fyzwm3o14wR2SLlaUdRmHV7ik
gjt1XkAEp/8gV0Zm2c4ZfRSt48swSCsjbZEuDPbhnPGZnnpIAimqiuWFndoqOljeMqXtVkaMSnVF
Ye4lTa53nML7GaEKeMvbVbrSTqRzjB8e63qUSvQWCP84OtFYEGfM4qNTsjy7UO4mHZU77wMeH8AB
Mqt531lOdCLYhIAnWXbwXlgpXKw0kPSeM9N1A66zHTq/Wcahb7a32cssGGINVJj4bZcZ+2pYaiS5
rM6tHu9wO1xk9IGF23gQte8I4HF8N6lVmov3vPDyTpm+oQ0MJSEX+nZGOvwkI6x8+TU6JgGnpOu2
2pzTsEbxMuN9PBGAMg6HXR/rkJH0XlMYwCKY7NNgFFQTTBtj8nBzJNEYDASRgu/fl82qu7V/d1GC
WDMyrQxUilBMaQYiMcdPSs2o7xo1KTh7mTQzyyj8bAwypzqiVKBDVJpC6uC8kN8qzpkCf1hJF9VB
ciKE8EkxhQrvY+I7CB5ukzc/7drPhI90IofVjzoidCqKw5bqDKNWu45i8uj02NvoD+O7YH0S9Wkj
PagxjORl9NeIWp+MmwPZpid7MH3mxzcuJGuEwERuSXXBTPyTAFSGj/4I1ftrfyuJqIu4Z6CIwInM
g9s+ZyqhAl3I7gWfAqr6vFA1QRlXrUrdRzLUW0X5ReE8EXOyLD32lpOSPWSqHqk9U+CbcUNzUd3w
qsPai0/bzY/69NXsaR31s7J9CxJgrHyfKbG8Exo8Ch3TeMxcSJHAaPprVab+qdBRM59tfz067tL3
mrVTCNxV0lL7p3ffCd44Wd+l2Y42qyo3dRDttIq0jN5HDlyExBkdmOcos+nXYU1Sz2ByQlKxpduN
szktJbvoP57JKEO6evDf6CqvJqMWVHyeGUbfCwiNfFT/TF97dxjexZYMJutMtxDv+QCaeGcsbCQA
bZr+7q5ic/zVpSNOBxwdq/FcNBlEVT0tfzufxKLR8bSC0wc9qKOqFrL19oZNCLUBZi55h/N54jTL
QK1/exmU9bGhYcERPDPwRKselECDIyO8VDyXPAGhdNbFI3FnjVcRlbzPSGyv+F6CjV4kLWdyzrD/
sYbsKtHw6yzz8X7n93pk1K4+Mh9gLGHA5F8O9D7wIZNCZDDERwrhoyX94TBBLKZ3FSmBrNEICWMP
koTCVJkRDyDj5WVviykkdtWLAuJsCWasKGsvmNxu6zAaNTcOnFi409gWa7bCuEYU6TFO67lbNVWp
kAmeqNYi9lWRx1KfMtSSKXyklk06koBSdkFpHHvfPvKM3oPPM+ssCzYIjQ4XGEcp9KqYAnbTx+dF
sOBSu4RUXxWzWrMYnJi7SVizZcOGpEGN4ZrPWhkCyEapHnllHwHZLRXSl/2FkGmbNClKsDrZkePE
WSyBjuq3ZYcRk8dAqS/4MhjkwLTCEZlBgcxBLwKcIV7LfGj+dt1GxWq9y0/K0LcvZ1gutDhgDrmo
l1TjRnX1IQ5VZ9hjOIYy4jJLW9Wu2jikTOa1t4nh9zq6kCY4uQ9cNITzKwVcYbKvu9W6shIpxVgH
piZhLrlHcR1zPCHZlQLwmC6LDQlLy80tOeSHtBTtL9+oV7WD1cMssFmMX+m6fbJIGYDml/0YNLYF
rsBI9q3rsv/xmR/rD+n7pN7hAa+8A5+bT5SVHx0hhfVqV7XYb3vUug3VpQhtK7k6b7cR4W/HnzG+
xB1ppLLiUfQw9DSg26bb7gwuom2lbcJDdxCsbiuQn0sxbVcJ8Y+YNaIJlJfBsh7RtcUZcRaBaVO7
n8wcHoTrRz0SHLJjrDQvUa7B0GeW1K7CgVJuQ5ErsOFg+DnIygeuO7LCMIQJwTpzquHMa/siqqOo
XtDsOcXJY8d1v7GBwwhhSRQir6blKT2NG7P7NPjUMGJdtnbrlJXQfOxoscPBE9U/kckZJUhe93I7
3OZh+yNpkhWbRUKOGPjQTEo4CWUWyjiaflJjXxnGGRJbsRflL132/X7NirLAkwW33vLP6jTduXa3
GaQRHKIct0XO6YVnouq0bgLvHtHU+w7sollhFOdFj3SsiNwpdsrb1gZ+wqThylPRcMW9JNoOr73W
YG/kHLWhB6iWuRdrws76K5YOG+RnXY2bm6E7UC+My2jaQxDH4F6Wsdmo6sArrR2CbPqmp3mKlf43
37kEo0CG0RPIEP0mEzvcYfkPWD85mclwvQ67/K05SBSaOuOxcmrBwkhdRhfG5GIxfWqVGbasr9G9
po8T3mqvMjudCHe2Sy34YJP3jEhavX9eTlK5Sh8XQu5GQieHv12YAhTfBddUIIpJgF1kPfePGl4v
dBdiM2XnW/rvG+hJl3y4BN0ERzeFNExRrSaVrwaBokL0HshQqSZfEbNFuk47BjbsXDMguMvU5r7q
eXiDC+sQaZlbx7rz9jNtIHz8jax6o5Z6MbN3nTz5jBFq3hzfz5oXyKokJdiF0f6UcZx6VYVhQIGk
QitA5Fundh6wH6zwDembjvrooMP+c2MJi3/xbZQCqOEJmJrS2Cr+bwAC+SkOe7MIvnP4WKIlYumf
30lRYMN9BwOfUZxysYAnuRCg/Y5J81ChQ1QGmN1lPTwBwdiHCfwMU6ah/flMjhZ6mQHgNpt6POQI
gQNxdjyS/Xd2RmN60zBpHZyQ53O7yiiykFwtgj3pUc0LvVPpr7P2u9zMv12jf8bLtT+NicM/Mly2
1/m9E3SWwcoI8YXHfTmwM1ApnJsxOAcwP8EXF3tdCVpcsubt9g5V/lIsVEmUB9FwH/XD93592QAa
I6CFPfTchh4S+GBGfd2FR+uDxi57HRprL/3DhDlVs9ev5kObnb/6wGeco7phyRfS5Rf8rp53JNzE
UHkxzHVyXy2vuiFOAtCEvc+4SJ42yKY6N7+x/CVI/Z2Is4kOYWFQh0ENdpnCi/jDILchMa/9oGcu
4LGDp0lWlVx80s7sjOwbD9raDpLq6ogbCCNpK0XhfyPh6s0OKfHjxrUQOE0vp/zsIFK34r6vy4YC
hb/IKotibxzvGcGBLXnJHTvxan7ivO20RXlVkwyHg1tdBdUhCk83YThBssy++5smbbAJlpvx9A8J
5c9lifHmusIbGkwkeAVBp/W8207wbgCUTOX2SCJiZJZSisJMFyEej2rmm20Hb7xKPXUfKhrfCjZT
0WcQjgKX2BnePZLMDpp8eTEKmXlLJAwbEwcRvp1F5fsdigoAK30E31wsW2VczzxltMEcdw1RhJB6
Az7ytOscdQl7nXeFmECjvPV4nekpaxPtsU/JVewaZ2XSi9ujA1LrUFHO4g4dz5iVH5lekmXH9UXl
zLxM0wD0Y2GqdWkyekN1Iq8sgW0Vxz5khZBt2XVAd4dr7IDuu7PvhJYWatDoEocIl1OKgkcSUSqF
Huawd62OsRrn13i2miMgUKgIWCbJTK7y5evbLOBr4RLKuI+SAnyUSAsoURO/My/CestPX60FI08V
WJY7bc8cAeoMKgddOVUxcIRoy/shRx1U9f3x6Ns2KCvxHQY+0a+8pfNAm1rkUqnEPiT/V/zFZl1A
CDOUsCbPfCR5wnDPfKKrbli7dwZhssk07smi4x3H63Ieto5pZBhEUBJ80EHmW6dX5voQsYkG5iCz
0upkoiOxgpDr9ZRbMhP/xWEfL4qkry7LAIlRA5E3oLap51ZMIb2+KGuYtef/QCHSuYvM+hXn9avR
DpQZo0CXatSkILav3CWdLe8j4p59L4oLtc7+MAb/XcploHWKDzJQjzA25p0JgsS/Pnw6Um7Tx3+4
06CNbJd9bDBNG+S56hQcq7opjFy2X+gMqGarcVR4yJfn+72fxOZJRN0vXCqQK1AFpr7NL25J3GRf
oxHMR9I3m6BXsozTFjT1wvqd4vDUAx6r/cmXgNPBhYfOsvcFiHlE3jBj0UFwCc9KRQF1sUik+RUO
6D1TkWVY7RTQj4MtZmmXyawlp2+BvjIoqoliM4/F/m4JmBEOa8T+xdqLmwFgonTLih5ALJK7txmx
ANN3pUzlyfzn+9q8WgH32JTHruYRTdXDTRQ7MefqBwQZ6Mbs0ZwPMZFv079Ebp0BIAlCwoH3vuOF
x8BtDMp+OLUaSuACyOMP1Na3b5LaRrocsCFVGukfx20kcDY4KmEHh/m5zRiarsFNrOb3+5/kxqiK
+2gAaYRMW7NElGbd/FXgM2pR8cc/6QcpeK0uIjsJfmslfn4oH+OMmLQvNxtyJ5oOSe57TJ7FeyNJ
F+xnX7615whg26k2W1S6ZHyj5lAp/JtG+gF8D+91UET36HgTnQHc4aGLxQJU9tU3/9+kFXnnX7pR
GnEvMSKP9+ZlOdg5HEFGU0bTv4leTJvXIXLsuUQMPI3OZwf6jZON6AfNN5zPPqfxbP5OJqnG5NNy
pkARlMeQgezlClr0RU1K2OcXC8nHKKFcHo5AYeag56xJav+zllnFWSJunr6LCPJbD8BN1NdRuWIn
XKPuQNorrjhKoYbUpvzvvUMLzkHo7FgXwyw4Iw1mXG1YOvtHsmzYgorZ96QtbsSemZKFqVuF88Kv
UR6cXLatFAkxeRBIbe0yHbZID52ITgiPYiXmQwJa+pGXE3sh5RhWNFIxaSSJ9I1un2XdYtfkZcrA
MnoePcngyjsfMhWrupyhMtn5XfxMQCHu5lfGcyiFb3XS9vTLP03FRooDJmfu7d9+YrWvbnMdPLn9
JpYxd07vH2iOwKsNchqPSiVnknoN7OyDGmrvanFhIBb7IH0M3kfuqmCMnwVhglB8EBeWqSy/ZkaA
zU5PSbQTBPYffSEaM9qSFDQz+SBCTw2re57pFEEZwUk4sobjJpYKyXn55s9H7QffF1wBxHTVKSGw
yy1AX5P60Tp9QglPR7JDB2OddLeqfuaD3y1T98NtwaybDO6ZaRObqgKdzsM4nZY7qFI0BkGUBbvj
po0BIzPIbh7iYAbodVyWK1VtYpMglBRo7yS7laCNnT8bm6CSph4A0obooDOfHT2OJB6SIBICXeJF
Zm1Fnp0Dq3o4varkPXfHrV2RFnPc1aKG15APToEeRU5OAu+CWeenkiZzsj6l5lelLYjEEKJ9Tt2w
cHVV49rj5tRYgXtuGyM/rzl2554az1MpbAov2CgGbh7eXp1x+shltmVzZf7qrGNDvPr1UKNaNpT6
kaJt2Zv80vuG5N/VIuZATKw2lyR+T6K3kRBZ5tjKONcZ/wPdc6LoIbCnqKCJOVC5dYLLVOWlMfBx
lje2ATYqQoMd37OjY47ZDUbd3d18VnRt43ncFzYBgWdmC6jZ+OJ6vztV5YZabdGo1JK2AcM3jFQ3
NaV4duDzPpiPi+vPxcMsEyWMvCw+JWKLndoxo2ZFrpx5v/I+xA3111XCdYPprTNwCQnhPpis68Hm
t5/xNLCPMn4tn4+N+WoMn5SMhgkW9ap9xeuloTVzYad3NhqsRvZ66+Ui+YqLeveubgEe30cNBk0h
Cyug+5nAYyoc/fcj/LPXp4usjyj9ip1d6/YjBu9h5VBcwdpO5SoUNrdUPCe+e74YMS8sdzKNRU4F
TgaOnhJtsH6KuY0rFB1a4MElknkeQVIBL2JvHmRU2UKviUkmCx8OJWrVzkqSIHBykzTQx1Kiwsfp
zNvJCVd/EoW2oBvXwVgkbuk1YABqRCBAWEq7eIaw3akF2qCuvqZWz6/2BMVzOAf7/4KsyKePRuiU
IoM4VCc4XMimKVH7puG4/Yd4Q2tGyfEjpTTjSpgiXA9ewPDb4M6Ne0yuYD+ROfkbxj0zDTEbH8XG
lTCkRsKhDZ4JnoXsatLbAotug7Cv5QlCuLdkLq3ojWSCNDmgeWnYpVnlUSlXOYlebcyT69xQAtRt
THs88GRhvvA+RV1jG9wcd9SEths77zx29DAl6itjjQrZ3M68MP6JpiMBY5YszDHfaXorhaHn8Hc7
wtI61hPYunbR+VXNYOK0p+ehK2k9iEAbeWJqL51IuJBAfdWXJ2dUCXjPBWzO7fSbxKj71+7YSmL2
7U0D6zpIjdS9G0DcJ51Gdh1GvaoguW40kQ6MebZhcMbMA0rRwJQMeOpww8X/IXfpaHLeiocRRrFD
ZozDVZhx7vXK0VH3X6wIYV1BbPiNwpGcDDDQAhKvVxhjYKvaV2CCiI961y5PMjJtEBfi5R28gXBn
ekTT87m4+XUOFwN8sc7yJYQoc3L5pVHftBJk04VLF74c/a14NT38zzM5IZcJ5fJ/iNAo7wn3+o9w
n17bh3jtMmbmekSqpWUCf8zY+nCobJdixqn9F5VT94Lx2aAiISJxctV1bmdjKfmWZKxR4K34w+Xs
UO8rzL4VJ7Ky36eYKczLJUmpSPmRq5bX5oi2x7lmOyMcJu0wlOo4L5X7PqQvdGfr3W5RG8w+IN2O
v9sIsAcmRpnqBYO7ZaxUGGUoybr/Sr1yujdRqHQAx/7mTYDg4/LIiPy448XHsd7GXCUgGzQGNYmq
CRzsP34zsIvpkBTLsljJj4Sp5DEQ1Hti/TWjOyffZ+DcsrolfIZd2VhxB/7Aej7S2wRFIPYV8kRk
0y8cNQvWP2WMHu5R8M9y+uP4L7uk5iiL2CY1YQxyGSwiv96jQCGY14EvL49Srz48dfUYwlGm+AQe
f4Raenv4lUIK7ajoP0WFvSE9pVnF8aYVqbJVokeGEREl+Nf3UoyJ9ahimdww46UNHIQ1QhB9JUth
pzclYRQbQiwxV8tSNTGBL4hzSNSV6ButjzKga+YEwBlroXEJ2tZiT3/TuhejXUp1bthtRgs8QhQW
vLdywNAIRYd5aohTN5xpaTi7no/jlv3l8rj92RWC0VIf7wq37zQ/l+pr/IVHnImf85etkltmv5F6
tYC4FoQyGF+ouJVx9w1373++kXi2+WTWCy9rNpeq3IJ3g5NZNRMNgrzF9seUVF1iYLfO++FH2mC6
pM0+90eNHLKH/PGXwrcYMVWsUU+Qv6L3rpGF1W8n5r7VD0lyZ8nLYfGX5myDWaW59TtUCQ8akNJp
gduyaAqQseioYtoefbG2+ghn+LYXXfB5k0jRo9N08C3PB/dNkk/ZTpQsABjaunukHvX8hV+W5JSl
3UJ1Cla3eLRX0VoMan0NFeZW5Xtzu4jge9xesp6bYm05pGtoewNNqDo8cCuxYI01BBE4uIB5XVUn
ec3R1mO0/zQeNDtixXnk8nxektz2Sla1NEwqNI4rQ8OiyytdECs+JrY3/Ee+vDhVjDApBwdMjJPD
8hMkp4HIiuPWx+6EGUdtVXNAxx4odTKqn3yPLm5WKtChxtv3I3ADjnuYVDMOhSEvIvStjLKsZpYy
AwzgftpR/WhSB2vGWJ94sn/tKfgDCi8gQRd6K6jNVQ8vB1qpeqHvucyE/u/UHPf6zHC6tomVIw/L
fRza6x+pyZ/+P1n+FQrWxYgCU2tlFY6RGoEFDN7PwS1KdwOtzVGgyAWZecZVDqblPbdOp/d0wcLv
1OABkcKvHS7Gx55rnUzIutPnqUWwh3uNrdE8t7A6WJE3jsadnVcd6GbHt+V0JRSjGltZkRcsWOsz
YTUaC6ppDEd1NMMerwy1gCdJuZ/DeBZ2xGWC7CfG7HRMr6obcRHkwxWQKfIYgNDazweq/c/HvZmB
6wjbNiwOeuVUQTnRhnzp9M+UTFft+M1tgyDEcm8QCCvy60Edj2Lye5c0oNQYUOgYO4NVWZwIG9j0
KSu646NwvP6hcZ03EjM7cp5ckUBvvM05bnEo+b+KfZSwXyrJrDptwBob1TUarVO48zP3CVkM5rSS
lXYnLIU8KwLqWqG5kCsTWi6PI5+Rg3nZ6flBUxey3W0iwiSvx5eWbhE5FuMrzgUsFIxyNsVE9qxA
GEWjgDY5SKZn1EHK1xGzs+X9YDImBrrw3C4h22K6H7Bi5ZMD62b00JzFVs7BJqJMvLO49nbrfwRn
d+YcHG1/jvPrUvlxUhOXqEHu8jNUwgkszeLpgqWrG53rcqRYv49mVsE5o0HsYayoOQqIf0aFaIF+
kHO/QwllVkl7I3cg4WoBA7iVOtmY28CHjCjzQ9x99Kv6HCmj/8RSn6F+c8xvwZvDNQ/wzy43/4wG
Q8dd5yVOU5eONj4/wxfZUXpyObEABcp2RejbYB+mNad9ZZWZMkkU1eH02ZvRcuAc8tgeIb1oXcuE
zNwJIs8xcTy38Hl2knFe8u/hZjNUyEVKIP7be3WFfBY2+R67ilyz1wCm963kVsbSv7tOXgSoXEaz
9hlEw3vUw1d9jixD9QcpYF4+vuQL+hU1mNFtiViPVysZp9v3SdDqoQRjOV+MAMNy4mIOj/BtHWX/
rjtvTo1ow2R/vQyPJU2dMDh144gw7dGYRPEiWKZsuIUavLAJKlz53avuIQ+/U4K0hR6Zw8PiunbP
dIIgv1yYrAzXfcEmbEjES/hDABx+h4mxSEzPi0MSQrbDPCfJXNS+X8EURy6hJqAoPm6UGnhj67b0
C/lTHInGXk0Zkyc7hAWuKgVk983zw4DlkoqdfCYn9dcPo4og9GZNHI9TlKsKbtibeX7z/tRkKPBq
qoUBxUco1nY/Re/qcvDwtbIZkGUvdauhDgASa8zSWskZhCtKfLGbwCHLJ1aWdgyrBjB3+isaympM
8UpvAMbCJ2Jj1npeaUaM4LFhsqM8Z7/ttogxCtV/5jBbTIHjOMa6PnSvhsE0wYcFUwM4YSPKyaZi
0nb2XF6XpOo3Hup4r0/aPw/PXZFUQ3xCirzqEpNhEDPUoUoiSoSF1+3GjMKEyv8Kco2rZ4drTDpk
OlYswuwkfYFOwTpC2VzRgQuudtqY/FD54a99YQ7/0i0Cd9+ida3qdWGj2PKR/8hey9/MNvp/WBXS
OWKXvMaah9nk/z57U0lNUlcvWqgoG8cXyQ0bzvhjd1/5hhdLYYnblohgCL+lsCzCfEgQc6YiZF0a
0XgaRM/tL/2L7VhjTADdvkxa72PBpJ8skmiHOaglAQDrauvZujVLRJw/cLaINfE1A0iFNftWuJWm
POVjd/rBpwqRVJQyAgKQhPA2aDb7+qdzzKzQQLSN/+BWcVUqPH4MLZN9nqIlp24zffchEpSp/A2W
p+mmThi/W9QFS6T1yy5aaqDlaXU22PtMhoW4t98fV7fnnlauDPknHbBwysF8QTUB9SoNGWp8L7ea
BzPNPMAWJOF2ALVk7L+A65inh7jAWHdJwBvDTWz4q3QBOpQla5ePngpCTzkDi08IBQWX3sFyDFPB
A0iw4qD5AgD8XCdPd6blSaQIuUFDvyrDMoZsjyjYQOHyvqiWzcQqonc84tL8cwVYB3tbnJ8ca31v
5XrWZzUu9wwnPx7kokUboxaFUJ/hizHyV/sNcnLavLik7BzgXlaW5s79kuPdbx33Cf3OWDTgBnIL
mdn7sDTlXCVOAu+yEoXZ1N7wmWidryMM3bcv4xJx5axDV1RfUEKlJLB8+nkxmgoXAgRx6qJ7Szlr
XwYn5RC56wG5KmSY93JZwOTrNO4yBPOe/6HWlkyUVROqqlrSp2SpSxoUyq6HZH12tVObhMEEQcEv
VAKAPet7UA25FfhVDACQDrUaedSHhNs8LWwtbRmXEImKWGfryl2ZpBCDq7/XkFkQlvmRQaQFlbrj
gnC1+z+7yUjKx0ZEIyZm6rTxuA7TkbMSWmYHUsKG7ypeBvkP75ik0wq5kY1+Drc1ZG1h9jpUje00
cB6byHkKpmwBJDkRiK+nG4VLijYdu1J08NLZx1keGgNzJSFMcl8P3Hxb534PZShrcM9YMuOUCil2
MdAmPwfcTSHfV3U4w+Nc1E6GNDxjrIwrJT9h9+D12D3fuA4hDYuhOwyWGCoDTx04mCJvAZybs7jl
Ipi5+IRVrDGUFrRTcO8so6bghSXBLSMFomiVjArm7ckFa+TV8Xa/ujnYRhZ560O1ZM6iGZtwY1SL
F1aH0NOysZYNrYPXtBgRd1c2Rl03OB00vVZ+LlRmFiIdIf8zuk7GYeU/InPv1LdpAD2olLn0WH1B
K8wTNJPOl6PIi0lq6WQjrhex/g0OOps2ifGaxACbLEQUCaBswwHkQqobu98ogZcbi8dHymuwiq8u
GIZ1RTN7aMf5nLSUJSsT9MYKU6lr1HyhBNtgkcqk7KTK3G/+P+bxnpK39m6yc2VF7H6lDQaPHYyy
1aahIRBsCFNV5gMPGTPxX6/rXRkBESjAflCCF/ZiH5bBJceLTW2y2+irNpa4wNNrK7MPN+mIvjCn
AVfSXjsZBG3Jeh9MTSs2CSsBtwEkJoZLhUnSsCvlD2Z6M1odzxM/NKZJejj699xcxiZBkgOG4QDu
hkDPx5zbFOuMoP03g+xT7psLMolPp+Nb7kAvSXmzWMN/rDgorLt6bBnfHwAk8TV5SZeAolW0jQXs
ZBGOAP9tAw3g9mg4a1Yk7mIa9qmKDo4mJX/RhCG0Vm+g5FviZoY0DojRr0n/kUt8ywyJriyZPKkV
QeEJ2cigQDy4qXRvzPAbDmm66xxHCUZbLbVP4HGuxIpl1mftZVen2vfRk6YeNh1O916JGnzkOfeS
tOGdAaj73stX9SHkUrBmCJodHqMMZAl0WYwYFqpuJMMHwG3u1jlPtq39SreRBax/rm7kQLsyk591
G5yGJ/ymdytynPCXAUPT7h9GWbngX3YV979wc+cryVb5/pZMzD6NPeVa8jTK/UsoEeBVJAyShCrg
B9R9LMdmQt3el6wKXlV9k/q+iC0vpu8A22yFLFCBuSxCIaBMRflwTy19tuMbuTPQTTyAzqT47gpX
0m+WSFxp1aBVMNWcJfzbTu9IdltZgam/5t5hPuTGyM05n1vXpCfq/oaCrWps+MJ8WmtVsSqOpKzN
eMST8MHQx/61H0Qgf2gq2VeQ2pzxt+HEbMjy947MMpjALeMZEFrtft4kvUqHMe39u/eOBX6ZSzDH
x+hLaE0lIH+79fTj8SsGVbp703dbtakiQOkCUEmPSkJZOLt8kU+D3V4mhUPRYOj6+8W+cIfy1cI5
IX3/9b3TE9XMj80TeqJLtFux0jHI3ndpSpXnzWBHDwcLtQdeARUCx5KuccStqcuZEan2W5sSCNsx
mVuZ2ycW+VaXHBxkttCpma/npXcn25ET1EPfv1TTUTTNDZutDAU7SaDj40wEsgGotu/N1KQFFd8I
5qFohPiYjmjgKrsDqfKMcsOc+hTuzmRjuXNVSi29GTpyPuCILCNRs4naXW5uu9icUqzUGeGLisT4
os+omuyTGe6FN9SUeUDyQ4SXtFQmtA9jN0MXkYrQaLxWtrd78u5DmsmgEMw7H3FNX1qM+8z0uU7H
eHvzFEYSwHuhi6pFuv9+7Rax5xWkGGBNyeNof0/PVx0H8zm8zrGxEmLZHgiBozFq4mpxrPoK0Bzl
Msy35xnJyOLwu0KJqnPqJBQpjiDo9BIEgw/MAPjVtYAZPuADufLBqSN8+SBANvfhVeZI5AnHZ1fv
n+b7iXxBUAnf2Va0PQXXOU0DPcJYcbNI186kLRgW9br4vLKheOiYCA/imgqvSoukLTG9Pbns7a5L
bhJ7D2bpsggKMVgGwsnP9fjxQ/sLyVN09qBDzcG3warbpogx4bIh+4cZhHITgVJ72JBLldtoDJtn
D/z/VcuR6oLq/HRFPkqZ4MrSX3lEt1xRW+IX4rQ9X9o91zoEmaMWZiiTID4cP81l1wDmplo/Or8q
wfQnBZ/aVVmAH6ZqelmMJbjs0lP3eOIxuM/dMTz3k8GANlPE9tovIdfzrQ9AjgUNESK6QOGLoY3q
/zOFVuSo5B4jeN0odWhyjnlGVCAia0kUo8hbPIVoxW7ReGc/zQ4PfV4lv8Qhq2VFxY5SrzDGY1UV
8OId+Wpir3VD5DnD3MIqnahTVOqlBRyBZcxyBNsnQssEsK0UayZm9BSIAI19TAZ3iIlal1/UkT+r
S5jCQ0f7KDdT9ic1ozgmBd50Vy9BQOpMIZJnWLNJb1K6J3dWCMlVbxuqc6ddM8nlDJ5/jzJTr3Cv
b16COtr3htQcbSppv/E7+7rMF+kHsRyxW2euhGyaqom+itFtNPDUOhCTpkBQq0kX3vsnUv2Fuk/Y
lzKjHUggnN+A7H8RnfdheHB4XjjvR4j0qsmTlkDlc7Q/kX00Edp9U6sZxQ1wGtvDiE1yHnIHWreW
zWXkDBUYpCkVfpzCktXYHUKfcozAXzKS5KI/H7kIcufFMkc3reodqKt4HQwPXxT+iTQvHmz8UFIe
ww3gE7tPenkGhf6cyaSW1JGvhimzprDb1gikdK94x3P5ScGUIFmYpfV6figRwt4MWMwPfetLKkg0
iqhmPLUuNTWXP08lfTc9IC5Ayqfwf8wK5+LWH+renkIunfFOHNiQv20LY63K3PmEw3ptqEbyk/4E
33TX0xD6Gb42Mm2biKfkf3KV+jkLw8iZBsVnRFX9Gl1ZJ1+qPg1sWYkhnZzw86zT39rrJbUN/nki
DESJHIGTfhFIhw48//ltAMtdLY87tjclDybh+ExqA8gmePNgLOC1DmJY1fb0cCheYoVEZhZ10pMW
BtaIcKX/iDFfBV/Kyhr1cAap8HFaTDVBd0tmkmDgUG1wL/IDmzyPVsCATqVEPCLBJKmp/Nwl486d
0nP5TNz7ZeNY2pQzfT5cx5vGaVZaflUUmSPj0Q1BMP+Uco5pFybqUuRq8RYolBC6Em03sgF18d7t
tJwVPExlHSd4VnMoTBaRUsiRfdxk+sEzY5EXPcwdHyB1ZtOBQ9gMX3UUOrS+dn7rRbtMg/JFZxsU
/KmJTWt7xUAH2pxMtVLDTvQr3mOY9pSDx5uQZuecvq7vXjKBN5K9AGjz/hM47hOlcsnYestDVsJG
HkcENO20XEeRwcGBJ7eOhkM1ORzT/WwQaGcgkIQT6RpXPSWb7NOGiiGNPlM0Z8VXdc1ApInC4ppB
wvnCfMgBSkKARPOiNrgVFSx7FwW/ffkCwCxfcdUW/ujxrZt1xWOGAU873lx50dRT2AROEIcDESfk
bb8ChswV/QdwJq9YGZQdF5942mK7JP9mTThurIA7f6WkpIl00b3N6b/8Eu2UzkPZqAc4YK2XIunw
BsnjbLrZjIiBKlcRhrk/yeTmKkhNSv97HlAUWUKosTNEsq9m6OwO81nuaQ1vZlPPMFUYE7f7IgBU
cPFx7iojv+8CJtogiuVOJfI3AJvKtpWOvlYuhx643qzNDtCokHBWVJlSLE5pReodJWP3anm6kxkG
V5QgE/QLtvXdKQJABHlEp31W8mjG74A/+Tvf+cX5o5TfFUJPu/49r4KCpQyt2SC39fSBhi/MB8OD
4LHfc3WVLcMnvbxVZ+1rHP3+ABfUPSN0inxoGJj5ht/7JUHZQTNcuGagqEJajmn3y4Y0A8V4UwWT
Po0LX7vPwBx39zz+OxKSCDm9oPv//+uelWI14YSe5VQ1g09ujvUgwN3QZhfSfsicJOWjObMM0B4s
lfCoat0Er4tDjzlDJjSzgV0SGxmYL8H4jgMjxLxdynWvqvSthXYqd/kDjFxxrKi7apm6lBenJxM0
DjJQ5acwi0el5OlJ7m/6qI6/gBuFVf4d6N1EeC97QvSwYpXixNl1aFjfsQs3eNJYCW39Yb2GQenY
u3+8aSPruU47Fvy41O9H7HmOQJqF3z/Lt++2BgGdpwBUOs/EfgGbZWG7HAj6OVR2tFpOUSao5zXt
zySAagDNKkGM45gXJMr+E99riRC7EpW83KCpgnVRfPW+DREu4lSD6JqJylx3yXjAmLgjFVkDEDl1
ZiwE4zhWIz6vVIbvX1WxR9AgmUm9OJNAbAqrXwJmKp+//XX7UnYHejnGqh4cCgAysUKUevgbN3Y/
W30dzoy2a4q+Tz/WIXlvIL3EuuDfFQytPCF86Tism8QJGPAZhnW+pIlImxvct5zN5oue7rZZsdI5
YipRVu87dPGYjbUL4fjRveDZOW/ypDTU4RSnA8X+kH6ENLIaNpbEnLWdQg7QWepyxxUqKAsQL7ur
m2VwSyF+HGO9WUmrr23tdL/xzbHrwnzj+nem6Mm2ttbmsALtqYAUu6sCjf2xIG5nnI3/q9kHBQvM
mqz9nySo+ukjqMJV2cMcwE5UqgaOqY9jufwODE4UkRYyoIR4bEjffSNEm6o52ZweLRBMTZI1bewk
osharqEadqc/2gz5kxZQftMmwGaD02KCzLgOpYKPGb2dYe9HmiZT6E0mlkpUiS5CgBO2v0jkQrc1
+IhDFgH0DNpzzcUvCb0ibdHDRhPgYfPzXdyblpLysEwuBWNE2qbz0F1Q3K/CznOp9cvILEYS9BNb
v+4DS+Z/etbLXYEEktM+Wnr/jEr6WE1vxd3lxeZ1x6Vzr3QMh2mZNqOUmWkYKrH2zgFeY7bDyITg
KJ4JNY+UVA8RfZhfAeeFPRS7aefSPAIGY8nKOfNhhbiD/Jgb2siGnBtCquWqC5x7pgJuWWUjBx/Q
SRan0ivIafP4Z1q7E/JVrI1I62FDTflMmfs2oQ6QpvZ3bS2JcsoRjZ3Ooa9ztUHl80Od7xOoxMnX
+bCi4Dt+n3BwjYvNyYuEaZ6wLEdS74rBucpr1g52pMYKLuWgZp+dzF47sRSWM0gnKZVcKKcXStew
+fpt+Gx0DMq0WGoz7RA+mzMscAqxb1X81LMJuX0si6f2W2kBiafOVJew33KCNmV0rNjG4xf79/MS
h2rbeHxNzo0KEtII4xEE0mKtCfEqqQujaUHktoZ9sIf4QkHENq3tSuLI8h6PEira4sfST3Kk/jyT
TjduatgL0LRFXTyMGlQyUIoDCyePsEG7F35oMDmEf0PzicGePttcVnN8SM3UeHz+fSO34N0dpkHA
oJHpkG2n+rSrO7yUlPEBK6/CrLBnXsXPlQ4m9TBuZzCpHwE4jcnCyQw8peLZGUdu16/hBbVDoBtv
Q4bEV8AMYoS9fh+CCKg0qC8uweJAlXN4r1zU/NvQ5izXqFZVqJ4idObLsQlHqnMuO1E6s7v3aI7c
axxeLWsSy39jeHg4Lpo/ehe526NVjMMcTYauoOp9fHPfhi+5gF7rm3+11jhRyky7itFGZ603tl7v
q/qjxm4sqt38iDoybbg8rQLIgXJ9q0EFYdlU4c4Kyq8USqQ1+CmgXxr+Xpf4XBJ1wix2ky/mkU1k
trkOcCzdU/uNGTRT7bRMVjJ0PF2TpLNnHQsrzSlMuX4MCxhKUtGTILJYPiNxZByceOmIVZ3kuuol
zm6j2TuhFKBBmppZ0L2b59CyK4gtYaABLrGB9gnVrYIWiJmHDZ/LR7YrW3fUtlt94E4ygi+I55s1
EpyxRhUnH8XosEPBFABk+OFL3Y0hnWDlh3k4xyl4rrjv+kEgMrCrFhAVKXGgMwdJEo5SoC34rtBS
njS3CoKOmQ50erHPfE8Qt6WCYguVdyGzNcPpsViclBwTiMjA0WbkGsROCt0raKk2V/OZKWxVGbsa
Hg2/mkam9zf9x6LTYQOunV6GlVoYt6cN8EdWQD/smlR2uMElmK9+dtA3QWFC5D4Dpy+QLfR/HXaS
9cFhEeE7NzFd7y2SzrYUm3ZYeS3l0q+r7uL5nr3bFuJhN+oF5zXDOSUeC0P5x/ctaopjv3gYjJxY
OukZvr9zq36HBejnzMXELcMdfhj2v8G8JxnSTvZff1dZtWZ8lxUwbg5kIGF4v0C7GDnMsyE8qwDb
XoqFYCHWJ9uVqTYqc0Rqf0/zNAHL2kAJjuk5vBQMpGbn0k48hM87w42FI4MS/I7AcQmFrc0Oo2Rh
Kq8ZH/P9z5b3ac4uLkpRusWB9JEHMvD6NpV+9mcrf8IwSn/PbHNZxu4XOU81JRWEa6zUXaYCi6h6
YDeMyiXVBzYai4CPzUsWot23upphM2uzaJA9jK8vMgu4LluNV5vKlNe4HS0DfNNL0P7slOfWd0Gd
YeEG74/95e44B0w6rUeXFk5MwdxKtmQ+hIiXgEAmjEOjL/KB5rdtLRQ0ApxjJfSpmNJ7dpOF33ge
7B98E96pIm8lQoaiKJkpZvhwTRHVA0wl1eOBc8cWCY2tRNVrrkkkyAutKekijENGH4qwCesgC8vD
uaPb8wJr85vIR2bZektfVvvN6xVtdpM3H26F84FK2uXzek/OfFQMElf1Pg2dCndZrGfveenbLTq/
BRNi08qsZhQbVK1KQK4IEUcYZ4i1I3ijSyhBINEwqA6iMYxK4+r7C+GTFHPruXfiMJQ9aV5uAkbl
zFqhZOy/GupdhlI2SsByHNrWeqn8v0uGSfgVqfM0DgAIp/FK5IRw7ssPlCnWRuTmpfJ5Tzd3l2lH
1Y3T+k6qiQ1aQ+cyT/Xa0MWKg+uHrciWUDs53xN9qVxIssKd+9L9BIBjR7hzyi3hyBPtGHpqgd1S
DPMJVcmFlfBXTSYNUY/zOipZL+lPDLZelv9TNyNmD2rUmz4XOrml5ue3fPjNhBBqErd+duQkyIR/
4D2kfDIXwQt8P7ouiMhQf8HRntFsmJXnWimBwdvJvEZZzFRWpJY18t0nQ7LzPuMghWMXiN5fDEHT
Ab8KHvfq9trhXS3dMaNQnnDPkmnsg2c7HKLCvmgz0lL8evK9yHVC+gkptnlctvBwfSZ5KwFdFrxb
ypOvlnhL1oEnu+whWoIfuZ/gxaNeeg7xccO7doJwemQBvsGgTfgfomgU/dB/PrP17Sw2y4+rFo3m
/LbL58iZhLNddEhIcSr94OB+qhvzxxuVmVAs5Webp38H887ZcVKLfw0CMOQGO3H34dtTBzNwllU7
a0gcYgCTQsV+vJCdUsXhNmAkh3ITDp2UibeBz+6iZ74Mm+pcXZ/ywneO6k0Yw17xteAvMfWCZ4iS
CBzJqsRu1fYJK9CfJV1QWbB05Vk5Ca+BBufi/aJQM8c5hCFzrQ5YrBXFYKjr+aKc1RFSYSZEqLEn
Wo2fAIaFgs8soaPgw1Z+8MGCUHbeppYBy7nfEG1EQTm6zvxobq520UYU/9iv1p88zA/roYd0lzuI
HTGYvdJWkCP/AQODS7qpl/FUr30FTIl8XS6//3Wq4mHJDHqe5eykV3Kb0GW8x6mkVivCBRMfrCcA
LwIyt7veAZWt4R214M7f2ypMep34UiHkvhuA2YWwQjBaxo5YsufP/gQoE76SAcNmxKacG1fY8d8k
orV1raXYeRUHqAnVrlGjA+Lg8QaMnFT2tKNJbtRaMdO5XIuNj5yk6Q6HwS9XSCL/+eAoDZNCZtT+
pMSdInsX2oxrugTcq95Sj72YiipBpaUjwMzQY/8GBnF9uCygx7nurSq1NeXvhaaDtLLGdxE6MpFw
Q6uJWxb3rCQJB5oYhyOHqLWFiwDeSWF6NFMvYzb/cPxjsnKJzDCYRrYu588666riaeGsopYHFDEU
2sJf97nWsny3v9e33n5Mphxb/ioOiE7vocyG8SLznTxffGKQK2zTiYJe9j0aZj9cewpzguddPO+Y
3UTpGJIemNtf23aXSxMsDSkSBIDEmRnQlHL51nuR+nD054S+m6OJUaEZw00xqSrCs1e204fnnNEM
xenb6wRdSJZT5rdGdo/xzep/+LLeiiQ/UwfDTFrbJSNPmz8MN8PcADuzj79bV4kFPXx2b70anu8h
BlkB/snRSK1xAJvHVSciIOL7s0J9FDj0ZnazY/baNxxP5ukzw9ImIeSLagDqyXMdAKOd6vhiRpGf
JrvdKzAhmltiwB/kBRfz191UnnvFrWYchbSNgW9dxgbY51HjtP3ESOVKuhcAU/dyxFv9MTABxjks
hysFya1oXJ4xHPtSoKaw2uhQsXPXrok3bBQgNRuJBuZZpyrZsN7q3xW7DRUsAhVvw9Fc6tVzssjE
MLUX4qc+v26xeD/x+mpVz8i95TDP3RBHskAeHsW3YBtqYf3SEjGZMkBuOdATP2SCZvKsV11Xutp0
03Qv4VgomwGH+TFkcdLuEBAp06aJtkQZGLBo2o0NR4fJc8FN0ccjM6+VvIDjMvF9RB6bnIpixoVJ
hc3npXX55lS2LmSOPU/fL2UsC73IHuMY2YaUZEshEvEjfUDTMrkw1mDOC1bPOWwuhjRZtsPxeChy
GeG2/AuJamkVqY2213DLfgtw0avY9ZGLH5xuwe58WDXlh8DA+7XxYoQZH34RR0nbACkEgT32K1aw
wtgzwq1kT31fa03gVlaMCd2aUKiYM7Wpg0dL/vw67SDcnudzuBNg33gHRtRtJ4b6Ga1WeFNQ4bX2
rRk51yN4UgKUbrxcTkCe8sMDhqR9sirDDSYFwRa0A1scvjwvt48+WBXujq+k5DiWqgvcuT3OjCwg
EW2Q0Mx0u6YKz4DvEfjQcLCl4Hczh8sJ5tNEdt1nG8tuepnqU+Fk/XbgcObDgCp207aRfZMXukUa
uwTiAteK3sn2qntOjsurbAsRYnRv4s3RjgUp3F3Z0yyYRxF8Xhzvuc80829+oSKEUbDce7gZy3zH
uxF5/qisEfcx4F3Y3vmzyJR7gsKMcSaONPfeYyzLLiv8okIz33nDSOoUaI2ay2fa4wVKCGb0Y4e5
oSWHFFTKf17azujUpb7ftNTRJyz4aXsTKoJywy3weHWcYL54QvTdtWG8Qty49mIZWIBpx/iLoHhN
m306a73s4WBnGL9iKQw9rxYWzuM5tSHsdPqIDS80xwAHZ6gaMyubPEwlg2wrnIDxHm7MRwgJ292O
Ty5UiZ6O+jL145POkEhoJdcFdBjFD50HG/CuMBqWG4rqD7XctLDvJuzfAAbp3MiHbcZhvve30zDT
Nc5xvfmfDD+teRBs2g+eTxr9EAP7vV/jABT/9APOGEeuGqvmg3ZtQB0NXgThiSw8UnJ/QQpdFX2E
6/eD9VpvEzz/STAtzajYaHxiflZugaE2RXeUpVkB46A3rgFh7T2C9myKUknY7b8RDbZjvsIR4QYY
5dFB60yJLpj4MRqSq3mxvFUrgKHIRu5okgU4OaT/7UPH4N0hAPJVr9qOM80oTfYtnpEL8/TdAiCH
UHR+3bTqZesPpmHwL4AS1Oo+rh7oI7KYSMJoL9cNZP9NSCJH9odYSN2R3DyVdELsFEae/g96zAMI
GTxYV2M4aCT1kw0ZhCmPEKDUVY8vsAXo7jPQ2hQijKs5YT0B8H4ghNfuAq8pxPnRWxNxvv0tsto1
BOgMguAPhdnSnDmK6/fOENk8aTl954QV4pTaGd21UNAdE4atnMB54EbmKlTWSu77NZGzYAshBmUm
IZJn7gue5WFxakat+IMeBwX89eEnkyl4TkEGET7KYP0aQ+zrX8/o1nUDwlNGt4raZqjxcedg9wA2
WNHj0ZXMi0dN8tMTscHA3StM+HaJADUa2Y4Vysz+Pop+0GXhSMW6LY4yOc6en/epCZlbTw9IvQ0s
prsmglo+WFuEmOcfpRFN/JqEAA2+L/4PwnxI8bUGWPkGf11fspQqk5ZocT+VisMtrbuNL1iAkeqY
4R0AA1T4FIPdc9WpvctuOxeHESGfkl1cqzoaD/blzUmdqK3L4Rxh3BMjc4v1XUsYBoX9Xxqmkung
T/X+8CLKwoM2U/SUcTCfiOoHHvBHfC3EXRuxBtCTRZJQkOG4karWNzN0l/6keU58JJvTtu3wHqc+
mAXm6BNB49ivk6oYyYw/2Gkmz/SAr1ikVEMziWBY0UxO1FM4zgy51CUbWbWCtBXHipd/1WHSdJoc
DjzQTsTl86inUqzwE+DLpnNerHlfO58IKRZmCoO4YANYOJyNxx0bJoxl0pXHxfiYjuUM4dYYtQlR
OV8O3aC/uukI8vfTGJlYoclFzYKLhACtNCW/5hYKE94GCnK9D+TlB6yJHatG+anh+G0R0f+UyvAi
zIP8+CDeORlrGCm61p7nAmk+p75w9K25N7xyzhTsi1ZEpKBB2yOU2JFo6Cf3kf6qUw0/5Ca/CXp9
lVKoVXU5zPnFPN6U19A3ZI0IRzRNeECYPc6uhzd0isJDj9PXHTduM8UsxkWmxhOQZv0XirJ7hptD
yPQCstNSGaPvlJDJz2RlrgWt2uFYW0S1saBGnyeQWqI51qn/PKcIkmd5ZBT2P/eXy/ngvlnJDoxL
CrJ94Uwl1OM4YevzJitAS9XInqJTLI9XmDZR/tYkgjnWJ4dnN/OiNNgZvy0/GbS2NZf1+ovTmUkl
4vkLp4g/Kafwm/KFBHZFjlzJfdVA61N+5emtNVldreJdS05Af2SEQaaFWNUcHrlg4WrD9iFLcjbl
sWKdC+HS8rsn5jcLj0ljUC/jfmDvg2eeX36AnEfirv2VCp/Pk0SylsPNHbXDtp9uIJaDBdmvvgI0
L5MZDUa/940zu5BXk9l4W35241kbx3JFLPfYTqowB7oJ09Xki8Y/ECAuxe9VoUTdDM4QLk0VCsUA
VnwAKJ2yWVe2K8ajeNlyWGVtQlAu1V0QzSm8AaPxloVLuZSeq2bYd9MxMdSBwS+QTcOKwpN9G5Zl
fApiyrZojP9whhq6Suc1Hq5BRl1eoqWE/SVZb3R/QgYtkkqVUx4aTe4KZ3vNarDr5D0olXO2PqTD
wnadM7F5GcKMy/6TZ956Gm//CyfgQ8/ia9cGQ+yAICJikFc3Dvvsk5PiDzeJDdtpFi6GbZhRTpXG
PeZFknnKgfvNCLGWK1U7XoBdgi7C1sktHkVDFuCkxoAZl/RWaHg3VApXklwsG8u+yIphl8Q2Z1aJ
nhEkQYTb9qx0dKLVkIuSCxmk/SsQK2IJ5ssgRg5pFA8S3PO+nUegxMsg1WQz+ZRI9aRBw3veFpZw
kzKAfGPhJffeFY9cacjCEv5+Y7LZICiJGhhDXQb9wWsbmpzspgKyZMnrnfGWhn6jUeXINI8Qv2Fl
/BYia9XqF+dQBIzbRQ0/1IWs13vfog0vqFXL8g0/S5O/wzCRJOcaCUzr8aQXFPKTlIkLNtnoMy06
/SG5ttfZOhOlgQqPzSqQAlP479Npp/zG0YAW7W6A/1xZ/16YNE4dU4N5d1gy6H9tXszSd/UObuEb
aSVjIzjmiBSirmigBumgYZn+IoWUIND/SOVAGNlh3h9ofUC9YgQqVoIVfT4u9MXG3CIXnLqmCCac
q6qjOg4spa4W/2KppD3Ti9CKcb6pJ6cTvdyUaPOHEF0xG2cIPkPpvtbaWAG6NHSoNz+KMcrNxHdV
R0fFcl867PSAyqooZWsPf3ddhQsy0zjldnBEKdx9BIq9742ZaUYdbG6xbiyot80QHFIotApliJK4
kPnREVlhllfdslTSjl0lHmalBQYMdT8KsiHU/QVfvFxGP68i8r4fr0X0wRBI2jrPbAN7HnXIblvX
8ygfe15/xEdjs6jjzEB9PfBhbllTPT6c5+l8TxC0Hbh87efmacJvS8K4YzfGkakIiPGUDybiWgYD
xniKBF+y/kw/A4VAaro4riluPxZFXubjzik7Sppqaq0BmdDwHCJs3mJ0Tnag70clkN/DzM8/UST5
XnLymm8x/9MRJSAskBp1ycUHzuFXckIHgwqIcjvxPkIaMxSU3qoACrkdjXem2qkjHE6zN98GSVl3
gjRUiioqtWqklIbIG+5P8CzJl3YycQA6LSR2BOipJQw8hi++MWXHEexKcHplG5H5nRwhP7G6FGOf
/TTY9X6NRnk7OW8BSy/bPnFomT51eh1yeLQ2M6Bj8STXyazSk9Px+n/bg/VmEsw1TsLkHe+8YIBz
qEa3UvBj6ygCbtyrr7B9KaPX/Z/cAlslwBbPQUAJe2X3njuaPGPRQmbywt7AgQrUHD8LMYfqRvjj
oLbVpXn5myfOAomDf8wXyFLNUnXW0+wgJ4bXsPIOQN999kTfBMQXR6Lni8z0igJ55M5YRiJNbXu4
iCRCjizlrOulxBrjR+bnv9dhLTJ46ktTEEcKqGU5T4yrU9reG1F+H5tG6cq8t7sAo6LysxZohOTu
GS4otn2LkvzmWn3wYQfAFbrhC0Ohck1AfeS1jvH61uFp/pErSBU5/Lh9tvE7VIe8OOenDHFeKlL5
wKL8dAE79cXSTC4SP24PNZ7v11YZRAeSqMdtmTX7z0DRteEAKkfSb0L7QMMKYgMPHI583TlGHxWB
gqAHlvdaRjKjpl9w8ryvaTJPlOdjjspwZaGceBN9+r7JiXOJ2zwy1KnAXtwooOIJfWtUS7FyrQwF
AfGWVft4yLAtt7RVrRjqF9E237ho2SIwzC8wKmsNjKjlGzKgWQ0YrcVp8sKQgs7YvW9Dnacy7OUz
ok+W3+62FmVbqugnsJYOy9AUD63ZG+AaVpWKJW6REZwqpx3dRomjF74JekiisB6RPWwHitaPjc/8
smDasxPmUWuc/2bK0dJleKG2/Oxvhw85x8RBcT1iae8giWVTeL8BSQdQsCuPspkGPwVP6w7rU907
JGq9Hq+ewVhqK0Lsb16bB8K7/3l6q1Md3bszStUvB1m5oW+jAD0w8zroK9kgAg69vi5euiSY1rb5
nD9uo4nVovBS8dSwxHR0O8Sbddt25J69lC3mdIoMG255wnjL+1qgd0pfcKGBtywJkz2YK10Q6KAQ
YF1cDED/YiDM/r5fjrukFtOwditp+5EUoxX/HxDMPLaEG8or8NZtim8ZYZCdrjT5C6vCOhBsQhKe
GEbkCWzjfpaJyLav2ycvZ3gZX5ia87PwFBmzfTSgoFGCvaUoH9w3c0trD3GLyAqbG9GJW0b8p0vs
lMlKuTsa0W1EpCwyxoo/rvXMjXbVq9XnEYtUrvV9KQ82B3cAp+ILLPK5aFKgUF/UUjQGEZmUkLUS
8cbhpHLXOsGAcWnTB05LhItRsfOrvXuG62TDrXYpyIzHDI1bHlaIdaiKH60Emcfg97AZhAX+kOS3
Mr15qy8FGLrBeCRmGEhTkSeAkTpyiH/sI2UMuf1xKhZQGEEbSQqz1tOiZyjmVV2O+eie3jDu3i8K
Ro0K/YE9fDp6aQC6/XIPVOTTHOSCHfsmoIhaaE46ulRP9imBHylcZ+paJW8X7Efpn2YYE0kEm8mc
uBkqGgtzvEMYZ+6AqjvqFzP+mLNP5iziT8hPsz4u0a9K9uY+3BD+zc+LzlRe6OfODHznRs3BT+sX
faos3SGYN8cbyv95eFdm0peqTxti/vbWB1RpbofWBQAtRHtBu6FBdwK6GD2HWii8qKb/ctv8dsPR
/SrAqzQZ5HB3UCy7BZyYKRNjRrV/r0oRZI9txlxAIlF1p7F9SB6eJenUz7u4/f+RLwSH8ceWLYoM
5tZENIB94Hhd+r/J3LeVByTT+lCbrgHWB+UJkIhvOz3wtsQLlA8OBrd0Z1coVpVUjnM+CbBV0VEA
WSYArIWVdrbFwx/kyuxizLLMs5OoNjgFN4bNjiDPT6WaPknnouKRDGvU1wi33zamqOCjMCCL2R/0
Js3XbzxGG5LyPii3MpCmrkot9x1nesGVEE2Oi3f2qBSi7O/RglPPdDiqQtJbKq8qFIjbkGBoKTbo
C+4vs9o6nYlez6D2T9P0ZeYx88yWBoYLgCplLbADpY96QdK/1fgMNC+rOaMK808zSYnNYJyjuX6b
OCHYU23YPO3kdSAqN+CPT3uYOQe60yO9kJhDuILuOnqzd2LsuRj/z51DNTuuzeeZ1vd6LVoA6ywM
jznY67Z5xEf6Dlq+K6eWhHh3qczo/NBYiyE0EZ5tsg4k2X6etbSt4sHrQxLw+7qavnQGL8ZfPyO+
Qa16BzJQOIoyA679IaeftuJEJsNphCGztweByMvLjeJo90KjdF7m/snn5moyZ0CsMDk/BUzCuBwP
W470dWpAj7JPKDdULaZ+nQo9nY9ag6pmgnzWu9ylgnhgAEjrIUbxZTifayBbszbdht4ANPLbZ7OE
ih4fD2VT+9LpH/sK8IRMVrm861Dj+6OKoxS36ckFuRxb73sKFbGaSo6M5fOw/LmsxsknbumkzyVa
r+USTBC4RJZ4g0Mbte+7jTVdnjIfVgaQ2stsQ+BBO4BH1W1ECEfTIo7hofOoZXYxps47yEUDJWle
C9nBAeI6hDugwHaUvC0obC2LaALSK3gp4xfMd8nedLKkAbiyHjjLAzeYjN80sFnr0Yp31ymt6aeZ
U8crMZ4QLg1NRQ/+PqeRIhlFHzeY/D+FwO30AK+UHlg+MltunM7GKi/ubLi5y3DLMWTb8laplGcS
3Ek5kcwdyNzmr9kUI3476/XUe0nhnae6eUjBgiFSuL0be+3UjPQxdncHkcnYyP4TXx3teCaayFni
W11jFlTqoAqYyFCwbshp0GlTMQNSDd5m6AbuqKs23xNU21gSKc/9cDmAIiAM+uNPxI/3udT0Aadh
j+nKxXp1yuFGW8clUqndTpZ2p9fLhQBI/xuNIJOu7k7qGNIj0i7UAMnDoYwZEVycad8dO/O32AeJ
B0smoVclhHwlz6QONMV92gsDIPJWA5m+ATAEVmz6QUoLPnOvwkaR+mGGV64h+aoK6sCH1Qn19pFx
HVrOOJGnGSAYEmXokfpMF6WUjd7lSRFlZK3He8bNDgtzejQ41hLEa5V5nnPZhufsUE4xGnYWo346
4AQX8YmNpvjdK3TQQLf9s12FTC5a0endoCIPg1tZFRc5QN/m0NoR9ZJ3F+C3GGa3oLTLXxLFhALK
HDcqaszzZ6o85ZRM2vCVsndTyURcSrw0gkpXCxj7mq8ec7kSgaOqhdNG6s5xwm9aRWxfMngQ0sb0
bKFLLWRy1GouTxbFybkUnK9XX1n9H0R68xBmMYdXNgOMguZ3LvJrxnQ2MhvBEuFY2GewIRU5t+8H
bJssJ0CSm86u48Vf5fBI6rr0uoK5YBKMfCE4BV4eKwIdhIvOup2XR9ajP5SEqg26rfkwP9K2P+dy
J1TnJ5TTeNuq5J8WZpF4OmkDZbA5UD5KjzUFpEKhGj1gnQ7gMKUXc8DQAA5gZz3lMhzadkyh/DIO
ftMydiRvhH4I143xiXSX1LpmnKgL4ydRZgZ89OiGsUQCzFIRH4e6ILR5l5OaHLaNS0Mb1/dPHFL2
O4iWUW+6lxak2ve9aZ86CLJ4PFj9jT97jGRbgYf3Pfco9jwOUOxBi1EAC8Ji/VIHspTudyUmnkr6
2anb8lqNj564k3bwUJFm8x2ShKJk2gbTGdBH7L1FFvhQYJh6rRgffnD/LA6ZDSDyCsjcUg3R5K0r
kTm9VlEhDX9Z8ndT1m7qSXVqnAltPB8iaxNKNNTAdTwINZ82lcPC1t5fT0Zgfb4bYum+5+tbpICG
BK+gpBmiTQekQaJkTcYHx3z1m2JXiYW167Np8LgmuGOHBJQE+cclYmoCzZSZh7iZRZZZvKTg1TML
j7HDReaoNcPllcicjefLcXxjW9tnjWrFDiolIAcsel/zVotzBZafMYC3eTWNh4xJn2PnT10ZkqxW
td3forlfJ7BOaxxjn9qW1lNEIVn2UgjgOkxD5/0w7WNgDQc0sBYX+44mzaQbvOHbNAXt8qQoPWyK
AoAtm0TdAn+PKkRUDJnelZUU30SUMWRekCntMp1/f8/CXg6mDxi+wFAplLFTAlU7wpZyq4DUmkWy
gzWyenIy3cWIIjjjlnRFEYHYzF9crUfMevHhsglOC8x7rsizNnnfpR8nVGElO3qHTGjc7vQ14uuQ
mFBePPLSinipdRMAikx3GszSqCh5KummQe4KMhJ+1bKvfyy4dkjs/YYHZz0wzNhg7s2OjXucAU0E
mPhESpkbTmiphFWaCHEtjaIFDNd7MaifNlYxndQf5TfJN88Mk5NXOVZzNwFqNpRFdLZEINUTO2J9
SnM5pdiyVJfdY9GQI5VhX2PPZaDLxPf0YUZzQfwhoQH58GVV6Am5NZFyF4fiNu9eJNzYMOveh746
mTT9Yhq6zdbNAqXMCy3alTc4HYYpmZMM+4h+BC4y8ZFOwy1+T2pN9SSaCjmQ0fcu5Vmy8ZuCsqvc
3F24QHZaBcQJHpQFRurtTlDyU3G8fysqtIx/V0KUJLE44yT39yuQdaGnzLd12Zh6a+wB6/a8K99V
uoH87D9CPwgG7qwlSvf0hLpsVP9WgMMuryTSYOo2PzCsCX4kidQ54i8c17ugw/b0AeOXA69b9koh
HMXaSS8OmWjUQ1xV7p3icLL5vyNUeoJC18AlQiLUOjD6hbnj46BWqKYZuk7VFHXMhZ2QXjCPRKI9
wGPpx0PWVtvfCf33rbbkvONK7lBeZ8IzoogjdHJnC4qjHbwaMz78qxDVajbSLEXsLPeCGX1TCRSi
tK8GorIA09eSr8tUF2RTEdo4WdptwgMjL00Wpx7/zy+Fr/c3q2tTjm7TfbdoX2SoajX1JlyxElLi
Hpk7D/xGwnzOG6OkTrYfaFa9wXYr/65INiSeAKm9gQCk0M3RCDP79u0HxkB48jxSqAilGZh62cHx
iUR/RqAbJQjWJhOru/poR2if8+hMuytRSbkkparhBdpYW6OPoHIaEefdFzTncMgNFc87CYdJnY8S
73BlG36sPtvhWK2sYO0DJV7ANMTsqo9RJ0RYo+Hej6sWbwkxI92lbPypEHej3fE6vuMWLYBGdGYM
iY891BLSgR73HM52AgzAC0Fp586NjdXaE7N0ChhroC8wTQKCJSG9FLE4MGpYAUcGmU20BRll+jrY
ou7WJOy5jrYZXExlXeQBks6W7PJmI38T0zZXKR2TrH5ZdPhF/FJVyxJn2dOBNX0gs+ER49aXnv/t
CdX4hW/Zxrbww1898eIAlfCCWJvcd65Pe9Kt8jvzPOXOn8TXqJ6KxLMOcXewv1Ubbb0GsP7RYQA8
je4IIuL+9+YRwLHBcp4PhQcpalYYLwRLG7WUBchfLUwaDtMWnHmNvnNG20/SmVEa4VGisb8l4gF1
3+g94uGGZLP/3EiNfB3sK6IFwsLeoFWn9VBRGtbxkkRarlSDeBiB4wMXmQlrHNdbwYSPppL+Kl91
WOajM6ntDhtxPV41UIAn1aojf8IYXPbfAVs1xBGAEe7rDXIZCDCLQXswtDLmoxS3lrR740PYALRu
MF+xl1bIodeGmOaw3Z0wbmYRiaqKDCE+tOZB3qXaiN7kcEYfajnOyAU/EsaB+p/GP+c2ninSHCrq
31XAr/z5Q2jhUh46LUoy9IIauBzV7qD1DyRm2pVIRS4xcY/s24L4tPQ057UD2eWPHl7/FRptEG5k
BcN0kE/TTJwprnlpf/66r7FtrYV6re2OM9Pv5HpSLyIkaxTGdieNN1evdvYXOxLGx44LPC+8Cec4
axD6iVUZ0NLZdJe1pU3rQILJHHreKQEHYiY9zsO3/4atO8a1hLmeiFzgPQGTlp6kzG8gphvwMmfL
GRzgp34uSzoBcYRaEE0HvHgYcoPhhWDVDifyMg303Ew7Mb1RMWUeIWPsIbGdOi/y6BLSi/vBZoIa
tD2Yvz5xegGf5zYH7lNknwm8e0J6NOXVO3k5TszQiQZpYHK2C6S5aSJfHxX0JGDeUlF99PRIVY/S
OiLAorajl9P+5cf/SMj0rIYT88Gk3ApPgI55hs5OtshIVF3Yd56+csoXLklxI7GVBZxoFa1rRgL+
Utlhj9bkAAtI/kA4JvmnJIoK9OdGzWV2lRNR8aryesTe/AdSlwTUNgrF6fXvFu7AfuCfF5relGtf
noorUF52+lhqc/gPL+lUMRywenOfGVpLxXh3g9iQeC/MZEklXS7JAHYEcoz3U5reK0dX6xJ9Vms/
KCi6K1ce17O54R0KkbXJnhuo490jy/zlz3NXuz4rUEi02l7BSyktLcXLX/zXAEf3Rtv3sQUhSQso
dV61rzONKytIXjQUrygsUg15MkxCc6stBfG5Yet/gYqNwLwC4BESW0Vyubr/QWOZCEazrJO796zY
dlByuAcUpRxjhFguTU4LJZ5YBMCxOKUT6YA+Qqx+kRlq5/P9KtzaSXfEKsa5bzE0GOF+ETErdC2z
eOvGzJ8VwiHPFRgJNrrj3hy8Ekhk/PCTHU06J7I/zyChmgU+AIL6Vf2XCrMHbdoTZfIS1MftlFzJ
7WFXOVBv2DCbAKm4HZzOA/0YmRn/eYbwwJ2RZFhWENr1jBx3I+NkMVvteBwa4CG66uZo0XTGTjOT
9V68MfQQXZ4djVW4mPPBeN7Ruf/YFOMJqUFgrU0lTXzwIaWKD37Czig1eEzzoDTLW7/F2nuylbkM
NPF6kgzFAvqSq3XP+z18mvD4JBc/4FxlIc2i2ioviSNFXp4HArvKaqp3bdOaXjBxnHrBRUNrfXT2
tXpNtxsGrxXKUpIDkhDp7hctrxHWNrb9bSuZqMhxGLqMZMsQ5rZa94bH8Ekthb7SfENcpzPFOfW2
wQ0NKEw2yL0eYk8cXWTaq7enX0iyymsQUeSFLjAsPaCHPnyVub5CrxVdlUi5I6ltAxkDV0X1x8//
FScYzARdnsXyTKQYy6jvvr6EXSFnF6cL8//mVqe85hEfEK9G68k1bmso5SOWJrIk+xsjB07GWhS4
cRG1+xO41gVVMBvz32D9g4i34RAep0FKd1rz7+1/vyRbd4tij5A5phg0xzJk65AG0QHRkwC7cMUI
a6/0gKIfC+MXyxws9kW5kQSFvHWM9aZI49nPYYjBVSTEanyKrga17TDgkgrBmS75RFGDNMbjy/jE
BAKutr7Mu9Fh7pCPNhzUmANlZDgBbaF2FDkVEygxVqYmCjCQKYmtKJr89tJlAcerK8cPZoeaGwZm
IUfA2dA5gDc25DHCZiKvxYToKMBBoEYDYfaBp++UQ8rwOj8aHyHEKRh0SnSQ/hUeGs1XF/biMfH6
cfX97cp7fmbZboI5nNTmve8yD0IB75XRXN8rKq75rtZ/lppPiBTIeWdiSsmoG9CezEnvhjjNTIou
El2iGZ6pnXqsEb9Iu/dYRzeTIEVt9jPXB2zTiBdoy5GO6+rBClCa4jOUp8ciahzFS0H1uh7KdmVZ
TDbSWLFjs2tHd9hVXRcaM0bOFG0kXxq6Tgi/tR0qkXQsy2INrsfj3IC6lMnL0MJ18Sairaai4mgm
EFKssfFyAwAiMmBD2b2foIjlaEaXGVMMHpBiqCqqKGPSPNGZyoOHjOm0cYE3RmW8mzud55EsAzON
UzXbVC88CLXZ05r3PR1esOXPt4e5bfX0a7aDJWEhv8mZivom6fCjrjbUVlFIji+a6Fw613f7u6SS
DsO+uBLURmw429/tmo83jIw1cgPxYBF080jrzE3vsX1J/cTn0vgJWiaF0E4xqWdhWmYwWJvbnZJt
qx47v90VROfdUF59CPcEJ6Y5JWtn/s71QPXqX0AyuiJQz9PYmDuPGtYpCDpvBTsb5Wrb1m19awha
+PuclF6dJcLtRb5/HZBvDiwK21GgL4sxwuNn51WstGpGDbzFVC7SIXXo2NSUeIojguRhSEmV+DHs
Dt/mG9l+phDgVuVTsd0X94t/0wkGDttUNKD8R7E5rkIC9T4Zf7He1cgH0j1Ll7ekn7v8W9QLPTPQ
Fl83Ajbuni7Bxa2FePICuv0ttKRBh00gmPKEzch3NgsmCwBK05SQ8ji8m6GKYOEM//sdEOh8ECP4
0Q5ytIyo6RKdB2dz6zOX7r7FCPw6YEALRkzNDyZ70tXANlM/kFHXglNOv3MyWywyMi96VVQAkUBP
JV/0JvNO0d7V+9UTwFJ/BDS9AEUk1xLcoEMvUgJm1WANU1QOjZrs2E3phM7ZuTCbizyVRS0D1yDb
OS3CIqYdq1muuXQLaWMsOrNvIaZCTb65DMnDqYRfCV/ZC9CjIqdx3jvk2XXWybK0/kxfWQbJabsc
TRqZEPxJODmwASJari/Ljs402YHb4D5wFWHOxVvBiS5fwmKZV4lPifCO846fRZhw6edwoIvyKbCJ
SvtlQUlEkD8tYMSMPfUhGiWvbRvBQ0TzU+o2yVLpmMO2yZuBL37fvsiZ9KfDl+frs0PJO6hlJCf/
V3INapo5Cr770eHOD0+Wvuje7rLqCJPXKW6gv6pe0NKN5jpPFzQ9zukB6adpNZXjwWIw/ahX+YhR
E4BRV68DqKxGp0yJdAtVNFhXb4rv9lQr+jMWwYba4fQ7SqWNIvafsvR1/RqDLHktQ4IZ0AtRJK/D
50zmSVc6vRKcH3+DlpFOtVADWv9AT6et/5ETcmEGN55eRfTC9ysvzJB2K/0IQiQGgyNNsMSfoCg/
zZnmg815QB5DI3HNzzEEduMtupTMhrC3KapqZzIyp63OkdXvUqO7AtWGm7iW6hcgz+L8wLlI2XXo
D+GESngLqyDC8Cz7bY3t+BfnLIbTtPbAuJUcPwIUyCEe0oQEfIs4uPt8pN5rNJO0Ymf6SnjGXDr7
yByG32sQwv5QB+UZ510Pk9tPiuOnS8vHb7ItleOI7AUfMey/1YEV7Dz1E3hR5UT1L4VTZEhsL+Ar
Wafogu0bNBjtU9IUnYVAQeTY4padBMDFyqrwDxgOh8DK7GBv40rptUhmO5T24fE7/cBPVjuOPed0
KzPQqmXe9ys/TF/tEBL+JCdwE6rwdO/Cs0C93wywzBrz3HAhtxzcrUjInH9/+3QwQOYKdAckiZsI
+W2GFmsbMpdMnZBmp1dbnH7GlWzxrgV/7+GUIwMzx2NE7fSfIabVBrpjgqIzLBvFv40970yMMBdC
CJ+VfaFaxTA7tlunhDufUktGN4i7XDsy3UonaKp2RLj9dNh3gJF6ff7ghKXq5IUxrNTIbGw3uDdG
eMG//RAv3EFFSWrSlSuEtcKUk/b9wix46Vh8xl4TYv3aPKDfZ4ra6Z8fUI6bWKlew1Ia4O0GCVPZ
n+HN8PgUEXZalfXW4llcpCdjS87Niuyfh5h1kspd/A03NFDm5hF6cVvnIeo4E/uIWjVXkzc1zXlP
BF5x01778Q0iGyOOcHQsBKF6+WbAcJWiu5nL2DZy2KXuIvKIJUVNCPXUtxGNJzASvsnPLyrqp6nU
Eh8jRdwG7ufChHnRjcP0MA0Z7b/A1+FMCupI6QxqgyE6KXAISydFv9REz3KbkcCtnbTB3KjDUj7/
dj7yQifRHpdZdXNULwNjqK8snnOjhuMDSYn8rPgjAeAwG6CUETih8Ue24T5UB3UC7R/jCPclM0YG
oKZwxwrOe/FhV6fG4B8JbzUvVRSJjiHuk7fCzrkCF+WlhUQXfAYCpgH30vUIAcWfmbP5KaCkPQ3w
zHU6oohT2n8OME4fV59vBRPkSS6xzUPDBclYQr9PcuB66u6Nb4hnM/2mNz8ZfT+LuwwbOa8p+/Je
y8ySK85OQfZdNupt8isbAL5HP+x7JCxNrQaaSfZLYFvJ7XuNuFFuM6YP9bR5rYUJO/gKOHmDQT2G
KPfeAnE8T0LTyyquWhFMKYx2nINwB/9nqbmHG4Q/L4MTFRdey5vd1/IbxfopOFvG2FhVb13/zxCJ
OjfuGWcImTo4GqUs2PthsDCKIvxmKV7tJEXGU3yQanYl1nZq9zO60EofU2zD+9QGqV7jq5PpY0A2
XFsmSeT0B5CLkVMSrogP0wCd43LSdyP6e5yRk0wg+1jURFvp06fTx+0uOn2atl8hAgLvSKqKvQ0r
3DL7XjYofA35boLKG5Utrq4PVAdxbVmEutr0XHhEZVBgv7I8hOEniQlhyCHhjO98XefJt5vbKiLb
CMJFXI4El4X7itcsyLiPb4H5U/2pCThiMBnUl83KH4HK+WjYfq1CZ9v+E67XM28LNZc0F9r8Vfhj
avkqcJysJ1lqeEBf2R8iRVqfQZsdlxYbFBGUcVC9ssvdVLSfJAtqt26hauQ4MKCczYPXUdHOCoFG
JjdPEVrJQ/D5qu4diJ5Z2iZyPvqr2ssGY1FohroU77iiwKFozd84f3+pQEfHw9foxUWPZtV6754B
ZELsVT8w0HvNhEVwRZcKWXYr2G3M5o+ykOI6mXpTyQ+7kGneHVE5UuDlTX9zDl0BVLzTLmR4p3HI
7N3szA38DXbfTesL2GEgM9I3/51/6DiAnxRZt8SmzF3vb/x3nBZffFWtwG2jsL8v8kna5G7lsnFX
6WJgmOTQJgXQRmUzPlMST2W1aMZwU6Ks6SQKftQHX1V0ETwHzUzhvFznsqQ41y3TvMTuwLgY+MIc
1q2bo7q6qPn2PS/e1+kjuYYQfznCoxceyjiKIdJyawHaqIjcDLda+iaJF4UnhK/uGr5bj0ASS56W
PgGkahExbQzIlLWY7JCKd9CJftE83rxFXhoawViagAVUuab1F3ywWYNods5roknCaLgCTnE0qQD7
PV19GG+d6Am+g7YkPikUdbO47uOCToi2X+QGziPZYNZAXmivUZRzAjtPbQ/w1cDO4ShuAKHYg/d/
rrErGSw+2Ant5eMhlcAuv5qHGgjsHd3LEAtaImrgp282vfWlZrRdYFs/bfjBe5SGeVy+HCib8/9T
dLhCPa266rMKYA6J/hjKz0jKW+183vbGcbbF2lMyBj5gmo0ug45b0WbBjw6ZfqsQFD42yYjF2kZX
pPCuBX68eMEBZl25tvo4gLi+6Yh3eKFmsTUqplc+ucVLK8wlgCokScNlEwvPhZWp2aPgdNcQXjKy
bpAEuNAGhZMWniGWrVUpU7EohoevwzYdIeTQSyxGXzb/HySb0XU/4GurRSz0tckhwzmaicpjdY5b
MuoUT98Bqu1fO29D/l5PoH7ZQ8xh2XKQ/p9Ir7u2chNIgNEVS9jZzLU/+eoQG/KGxpYTgHUPda3g
MYtcCbiW0VSpGxUxC4HWX+nKP0PuBuBrCtRNvZnzFiAFbf5cwoC6JDa6sqx1TJu8RfCVvyIuUd7w
JU3pfkAo0Guisdm1QimD5RBZxVCE/gnKq94Q4THIVM/9UguRKJ4zArUX3Pntkv2/0n6cT0daJVYb
wkgBjK5U1KNLt6GevI/6nLVXzde0AgTtivka7KoCV1xoPLcwQc+Iuydot65EzdJTlxXAeQjA0HHl
KcwjnBB6QjzGQmWXQiJRX5p9nA6yzldjuz7h9/PWi9A4Drxal3mGwp7K/jlyuTma7VVDiaA5erLo
s1S/f2qChvuM+sLK42Iztvpq2QcyVVOnOHHeI45m9hLczTuJKwruHh9tC1cMWGmVY5XH1pGElDeA
QjZhRfToiBIPnV+ZdpPs3skf8ktqF3X2HlY/d2D6txw3JrcrNmPqApNqR7cKG4cjQzmO2e3AuxB1
Z5Vabk5XkxEkAcKHOSpY6DpNOw/ZXuJmCVVdGkulrdq4WdreB1/oiWSj7PkeV3zmEJOybRYZ20JA
EN2RcKaJ7dqiuG9INQzS3IGNgxcTP0QzNdgDfYl8ISj/Nj4qWpqh91aSnqlNqSHKsw1OfecPRtXY
+M1so46bocqIpobexifftiC4K59Ivqa/6631CDQvHLh7HZ8235d7l4cIiSglvfM3+S+GsFiJVX0w
EsLBZxpw2/IUGPY3bDWpmDfIj3okM5g+6HRVVuKQW8VpwXXPic/KZXvCKGVpJ4gwW3tJZ1fHKaY/
OdAXZ3X5d37Sc1lsr2KvKH0ZhvPlI569qyWz80MJE+ABPw8V1EzOUUJX7jpRHwOLh89e9Xy5qLHl
ANSJolDcEiIdrfOcx5BY/pvElSWjqpP0ltMeG9ABx6M1BmkB/t9ACmMP+9IssyyP8he4iXatRC2c
UL7rkoUi2RQ+BGPp7JlJfHdPwXb4Jtnu5Tf7itnkTM2tMelBhPpztNzuT6oNMnXfp4PtcAk+Yyry
X9t7QQsGT+Xqg93sqB1RfiIeq2KTeIbue9RhAfrH23ZIsUvGjH2tUGdQf4OEt22vLzhp7xxdWs4J
JLjOI18PR9zu2BIvAfUoyJxMgsmu/sLwk/YZq3xypQhPyejNKSjKOs3O29WRYIGKg9TP0KXz9w37
M48vV73p8mJO2GPuPymP4KEQAa0/HcQJjWH+/yeSLupKYKIOTyddf4dOLL3l1m7RWsNMjQdad75F
ZU17Ek9X1xY8uGxMhnz5hndncU6c4ZRygDYFNbzG7ilE4XYNfchlpzUQO8O2XxiKXFNtzqsj5bnq
64OFqaF6lbepLg6qYu349WEeprzGe6bopadTMH5CIwIiPgKFJ2Ot8cAuuBg7o6jgowUacUOT0qEA
ja9xG83czxSbbC2jlOKGbdfQbxy37ToY01i2j8qPVQfxaqlNOhq0ESmTPx9aKOpx273IhoTc3XIu
m77GC9Tb11c23Z/q421x69RjFjeBZ+3dsKfHZEyH7MUt5ENVuDpYj/f+q6q94Vn02Yy/6VJ5N1x0
aGoAMGrQQEmzSIBgAyRMGMi+nRv2BoPLP3CFMOcgTWBfxq/SOFUXipzWDUUiHAEZqHG57NnLi5hx
VSOqM75TVBAwIndz7U6K9vu8V35XWIbPZ/SiA26ZU0t3k9tTj9xuc5IwJrACi8DbTRKavqxxPnGF
bWmk9QPAaNodrdxpb0kCR8FngIwfeP6osLpEdu/dlMaZZ3VFDYgtw1uVr2DsExZVL/m1oJD5kaS5
8NA868dtpWB+/YceY9ib7bseF6Md8ytWGhn0rKNddWimYIm8rdsBky4xkahS6l2rKJ4p0rhmc0CF
XxEqMLXRRTEuItpGLBW/pYQW+Z72LWCyBD6LJ8P5MFjOauKDTYQoiyyVo3pl8dArbV3VYyez8+XP
FBxUPgbab4+ime72nnaX2B6beLsZ98SvWe2lIXzC9xS1qbRcfab+R+Vx8qmUiomU0zJsweYw9Q1v
yOEC3QLRrs1PinWYWo+GMXtoGQ8IziJ7uAyLq/qViJO/tyB395mMVWNH4TWe3ArDTZI+KUlj882z
SLloowuPYAhngZNAv7BFtLpBuW4LaQvinm4N4E8fzTSFVUZBAHtWG1SCZX5gcnRWoedfTFraC49w
ZX08tT3RIplbsgPY75VYidUCprGtuyYH4xtzdSLONOqKcNcip57WwQHbZWNMvKZuULoVuJgzXHw+
UaEcWsZwN6/npd0qcN6FGjCEt0MDWJrYlbHEl/FfPjdM6WYKEhMqngkhpa9kg/95zM8fZJ6HaVc3
gQWu3yPFG0Qtmpaen+sCXx86DxzdDczydGrDcLKWiyM3KK6c+L5m2q/gswmDxs8y9c7wtS7tT8D4
z22e3Fl+hmUFgzAxhtsrHHOa4jcaPerIohThzHkIinY0XBJaTx/gjOBV4m6D9GeA876E0sTqMR7x
nwDb4l9b4Ua1jsJN06kQCVg3hvS1S55AKATj8yHPtw18+y2ZKdcfuQpDF4J1vOJ80dQH0xvvUJzB
R2npMQAWyEfzwMR+uMyaRx3JmpYlaAOyVVvxq5AlpoEpxRWFKCJ+uaDBjmXKG6lAKGj9oxYdl7+H
CFC1cZXgWBi01MwCNvCazvw4R3iBTL82KTmKaP6JJytaBweMcmZtRu0w5wn1dlnccT7sqZt96Ixb
NtPh0CZZ+V8A4CCotlpBYiFXLlieHv/C77guK3bG5xgG+pY8PqjEl1VdWGHZD1Ov6x6tBHqcz7we
P42X8gghvfZ/l2PT8i2escQFLyRwTeMDmeosWSdPaF1K5ZGFMXKs+IrMezXHZBtXaO7audQTGmaN
9BDmFgy+wMaiDqNOpuFxhfYS1XlFVEJiEAhxzO8YF9MM4mNOrCZh+9MwESNU650JIGZwnw6nJr1d
zKXdRN1J5p0os/6XWIuiblDWQtt+Fj9xMHTY+fqiJb3eJBcGIY56HD3xW7tQymGcztzAfmhCqz3U
RrIqYc25CmBqzB5EPQCKnNaK/QQ89L+a5HuO9zicj+kgOdhberfOGxrDNLoEa7h88Ic9TkS3/jO1
O3T9sbEchnNTLXnkYgR7AYOIwlWbNjCTBQchgvnHMhovJV4AxGmW/+btEoq6vHgND5g0Nu/mMgap
4uy/7aOoX/yl7a91fjIy8JpsKzQdC5veC1s38OyltrHpQrcLM/brjpMRXZ22vuRw/Y4ZKfPmILz4
yLw46YyIpXdAaytduDkfF7iHX+LMVwW95zrX2zxE20pibsmC8jmXSf1jc/tLORYAVWQ/HT6VyPzX
NPhkVn8KW0NwMeswNCBqait1cyP4IUstru359yoB2yoEkUGJHEy6pWoFOPkyw6ckmqXG8H/ogVQu
df8LBtafKr5HGbaVnP2ahumbqYoeInHJZfzUeVJPMWHdOKuBbbArD95yBZNoWJdVtpFHCFeFk2At
iSGalqkxX6PeFLps+0ENxYzn7X9Lh+vqu0SBBF3DmF4lo46VJR1G3+rSe1NwZveBHRdXpyC/YbzT
GutisTYXtdScdM83sYlO5jxv0xoRdBPVJj7Zc9tmuLr9euCJ/EywpCd7Mt28OViWhWB0HZHbOQEm
/N4TbpCEESxw0bvJqvoHyHGQzM6PiHZdYvdw8SeSxAl8pWUsnjIY8zkFZ0qy99IeGjbv6CmuXtG5
9M6dPWbys49hhYr7w4kM5w88jY/J/ZjSMmH1kAPt4eqTWWwwTPZfagvzaBCO+2mldP0ztL+GEmRE
c2fF6TRCPNRHJR9/l+tMZfMZcNphYcxZSXxrIjszV6VS5pbQPJ8Yia1YGFb49eaZwBEJOk7gz/hk
F0pRWOTNFRAMDnE0/1aV9vRLMfVMlAFxpRxW4kJc5tEI/5erhxR8pnZoOh2ZeP8CGphNCdcaYK55
Zgrl5DLMOCQBhqKF4K0F2J4z8FgU0Oqy3FivUg7+J+a1JmATls7MeBK16uvHbXtufhpybMohr4p9
rFRQ1L2abL8fHJsK0NwddvEpgnpIHKjk/Eb+7IVZBO+LxUScXmPpKb8UeheUDRabv/ruHaR3Pox2
RFtUyLiB1viRY8PA6n4MfTyVaZFoWFaqzN8JFNjk27SjxLgqYwjqsIp3BwSsOx4Myvrhp3Jx5e+z
D0NmObhWiDE3pP0KrW5hcCNq66945Al0RemiuH3+Eaa+X/9rAGxjk/nWa5ShhffMXv8Z8ZgcvrMa
xTOL02NzFyF1HvtSZdmzPlYExklG8/oIIPHWxiLgki2PIbUbQnKV+CgFdjpSPZ2ftc/qP9mSuCHe
dJyJbo9J+y8/VvI2dbsvLlqw5+0l3GC71JSLinhJNN2H3biE1kROxMnTsE7qNL1bwzD2A1VR2DWw
bIGFDppvMbf1hKHSYO8VcWIYqO8CMEA74WtEFdQGqfn8pqqKtDD0mbtr8uyFlr7pLF8KIc+Wv4Cl
1OJNN9vWZaxr7qZ7R4PgpHx1ZviJDqc9we3rLK8rgXYUwzSwcktJQvFqUAd2G0l9Ung2kBAJ4MC3
VN36rIEkjiehDIKsX8tAIzWdoGcQVQjS//yJRLjAuduVdTodyYs5Qe2skGflgUYOF5bY3mcV62vc
eRScbSEjEpzcg5qyMV7AssvnkSAoSV6n4k+XC0GRlq8wlqOxKNjfnC7mcgnb7tniR2pGiVn4AUAY
XRlbp6rUpS0D9sxrU2RR0LwCq1j4CeIN5KvsW/mRnNbU4KwMWy77AtxikV0lfIrx3MVFVOawecZJ
X03c2yryIcHBPDFPe+B1RSIAQmbhLmgQ57uroMtjUr2kUCA/mHnGaRs/dyWhyy6Vb13yc2CWhJRJ
zLSmFLtNqb8pdokRZJ4nQtwXMlvqH5MQDBzkZGWb3QUQTidnyzDMl+0SnQMBNP4Wydzo60ylJWay
M5EDkP0vAn5/B1LvxRuZCaYQ4aQe5dbFta1nXXBnvczrP62iSS/mO1Ct6Fjka4FXYrrw4LRhqsrr
B+X/gYZ2p9qM4T3PBHn57qwGtfdr/EBGnK9MuJ36VcAvqpDIxHiWbm4bHYADpOXjPGefpM8zPSdk
qna9NHF+wjkTy1UVh2DxnMF79COKOBfdv6hnycE4p350iIcwPzyAAgiG5k5RFl3eVXrO6St3lWSZ
ZyN9+YP1kGn1TfvmlxTkT3prH5PpXlKmAvAMqkzC85mZVvuUXf/qzMbFI5A8wmKdbIgGArULJ0N0
MGhAQ3ahNmQV22JUm8fMV6sGCVxfrjI3s/l+0o0IxhSrKpevBUzrZHQJzZPHUrXV5xvZ8wkEAKFq
U2Fmu3LIEXJWV+DyizxFS9KU/4kfzNZcwyqWNO08F/G2TQQKQAFiHEgLNoE95dFx8mDTHUC09M+r
1S9VQ/WWiYSmFYL1k9cAROQIX5mS7Vk4XPKuN02K2XsVOT7QNPN16oFnjeB1FuY/xYy5PZ/rdasX
Ibg0W2zK243JThP7jxFLhD7u2Nfj1COdkCBUpjQHmWWDPVx8eNUqCZVkKoTyXCjLvixKpXNry3WZ
p7c95A5wqNuRcdeEsDgoyJ8OYlR1BKcI4dpEJlnH7gFOJY/aXm9gGO0IDrTLGXv1IRUOB2zD4aga
Mo+bL56ZG0OhzYx2VHwmBwE9uFAPGmEzAuSCAtQWEYtTPKwioUl54MDGOcUrL3xOnjlC/5iDJ7rE
9BfU1uzwCk9s2WzzZmfMHz/63CRv/MrUCSx5x4sR5E0zoUjjU7PgGfk3Bzdl5zeLW2txPFTiYnbi
z4WbJ0kpCAcHMyIPsP9l4qIXjWRxDfnt1hbZ01wjIsMmU4effBfIhaYMd70DIEaaD9WXae8ZmhnC
zZFR8lMQ/D2TIQNhcNjuw7sO0atDpnwSz1Z6UD51pJtJmjXy93ECFbtDiCpN13BPDYvnjQtpGmDq
EbV5x8EJI/xiwcFoZyYa5afqzStULog8NO5PLS7k7V4fnF3jBmbPAS110CaXwnHYW8fhvga9mJgB
fwu080nVyfdlOw0D8j8H/w+o+YV1IBSUzYGPY/5xaSvTTJsVlj769uxwZZyP6mdEMSgGHImw66y5
0RrdCupX2nFomC/MBHGoueqVU+glZ3LFsutRs1PN1q7o7EFCCQBSoDZ6S7h++oKDOixdBvjs9/Ua
3tCA2I7hoyc+1B+Hc8Ttuh9vM7CuccA8mPzmtDIp4D0J7KlVOWaFs0jCxyC/90oZeKuIynoJ9KxD
FAg3xEd6YhQzoPhBJYO+bF61T/IAUkQlKhFSz9RgNrrPBRB8twhp6S497b9whDz5WBXhvGhnocIg
kHK4ynZE0YORD5CrpOjG9Wk8aQptbctG7y7/yF+gGLnQve29RltdOdFrpAnV9z/7e2eDHc1Alstz
IN7XWZ9m6sPkUXaGBA8uhXenv8Xqe39u1XEAY+F0CLpWp94fHgSxN6k+roj05wXuidVIIyhgMhOn
/F/FgZbaqaeTe+yZ2cD50FJ7gJvLXVvAUbxR93NuyyBnsevXh1+IcDFnZkDpDfWNRkbSnIV6QeCv
CY1FQ5G6YrWzpr+jNKr6s/W5KJcqDcLicllGbMMx0w24nBDwtWTnLzv61Lqt4WX9ALbi4+hTqKV3
Wkz7wMYtV9EAHTLZSjBnzxxbzE7OQK1x2mzgs2i6yKOOW1tTjA219/96H64Bm8WR7d2cHBXp6IyG
Df9JkX1zf7dBWH4F64oqpSN11i/LucF90fUZeezbI63zdGenaj2F7N+4hrhK+qJiEVJPM2Xmk2Br
rG8egVj/nddNJCjSDrgC0DzvG5fBUt/lqa3RCLd2WYGRs0K4wHzoh/NAFwYKO1CzL1mjyk1QdlGE
C2Wy+cjpGkv0iIX3flBmLRiYfRQ9QPpyIrDqFKWonerpjNzSVWUKfzsLtp+6lXhgAvlVtzxWiMKx
gjMMEhzMAYDVQi9CyUyuhJIZslT67Q8Tqk7OSbRL1YnpfbqYUr2TygBiK2FIaN5L6c2B6j+Ufn6s
SGFQ0kMItgFVjFhcqn6Zop6pV6ikwZH/oenR79kphSJ5J7Z/2H1bwe3pYTeGOnFCMMYhJf2qrY3Z
0doXWBjpoE0J1sBEyv9GQ0X2MYA8nVahC5/SJw1peRgtFgej2SBSxK+2k0KLaZtdlUPP53YRmBjl
vuAJYlcbQyu87ANV78ggGY3gSVePLKfwXnl/ZwDNJbacAv9/MNp8DX99fLV44CQ3lxrH9LEpD2ZA
jCsh+6q8UJ1S7+UGQ3ksN7kVG5CpcYjAoP1HACPqDRTUrO3LyZMmzo5pyZdohfUn7jeeycHt5G5F
NHCiQ56a9rmj9q2thgN3qEBBRcuUP9bNoXQ6se2XUAVPDT761mNQUp3P5+29urvIV1W4OC3hHdrL
KrzEKd6cPEHwRJ6OQ420kbnkKUp8AKWpQymqg+kofZOgDyamCV4F9v/78hTV2caZcdaNnpxf3bWl
r50QIhbvn1vFBfTgAoFjROEDoMKtsggGKCW1c9ed7x+PkS7y8TIBwNuW5f8qeLSk3IAgJOXvSv74
CDSGBbUK9h//SavEg6WHtZ+cbkhjaTIErr5d4px6dJkZ4RF8cDLUmK96hKgFNkdPhSbvWDFZdNCr
C4XYktEtkd63ZW/ePwuGGJIP+HukyuF0qHoEgAzXImurn9WlKV2f7qgAqjF4jx9hxwP+0T2W7QUG
/s3vmkSX3MJNLWq3gj7m/+JaNmNHa8fy9mTx2tZx5uMoJRl6wHMvTvSBv9UgtlyqRH5lgFb/+aOB
e+WLoFcLExBZD59vCc5MRoPIi3i9j789+Qu4Mes3nxuqX4vPRVOi46ff1ULTD/LY8K4vEpSrBeL/
0F8/vSQvnwIaZ69FbnU0glLedABVRuNAHLaIs08SBfIOZ++lQfxL/2yS27jlACt3fxlM7rqghhyX
d3OdLcLWQ25GzejefQ+VXbCoFpOfEk1Li1Vs4V24NIiTaPvetopUfPyDO+Hh+hHonnW5gFQI6hT8
1RWa7ijqpFR3yupnAd9C7DzDRy+iZj1JARbrOeDH0e5xzXuzPAylChjHbea9ng+hjY/b5W1np22L
plh4i6qCP2hBaKQB4gA7OOiLxLNbpPAdY+dZnEkKErOP885YyQ5uo8sRLcueVJf48TeJR/Pcvgrq
jMyuXRFPjNjkgmq3mByJW1WsffXj8066DeiypwMmiXmFTDfpP1ws0mOu7RrazqMwuubA4hnlrsiV
/XfI3K/Y3puTSARLLxNH/NiYTlGPuWcDxqz7ulDzaZzfRYrSkVZp9tPa8/q88yojjQXl5nWDFM7C
zjqGgIRxScvBR1wBz6oOI14tWBFWfnRt3A5F6A+raz5t6ueKEfuZHnCT8uN+Gq0ic123p+Q7fTPK
TzK/nJT+g/LYo89aRkWl2S0Pki7Kx9dibEbC2Jb6EWN2dlpKaEscme/yuGvhVdVTX/xjv26GxgPI
rcxdMObBn8K0NA9QDCS/khff3yios/wi71CMx0kRTt8gaYG4ccKUD/4aVimYcpX+8c3H/EJBQaQu
N5XqnAEgOnpxrD6cEBNFc8H8O8spXDgau3cdJ+zFZMWisGoyvQakYYmpt25IsHpi8k0oJopQrpPk
loB5oFWM2cKUyb6m/oYn0+mmpMTEPHXfmVHCyw1GBtp0dwT9S26PIJMBNk60K0qcLWAJw84nd3a0
saO/NQIJ4i0L8bWF4p38Uc0TaUXFWVqg6a3aV13Mk2prl7y8c9DZTEo8mNakNuEjgEHpOQkf+Tqw
gcj5cMslNFXDgHWgWV0odxymSwgN4cd+LIpVzUiX9UHfRSS93CRDe1QE/Q8U+3F9bcxd2lUVU/v/
io30AsQ1MYKBdW9gMI+NFGBnZe5hVY5Qraj+pIk10Y9UXhfSGDBMOB++SMhG7Zao8G5Hcw9NYAZ1
WsF6ighhsS2Qkq0ixgiEOj/l67cf6dzIsiK5hsjKseMh99hMLKPE78AV3JtZt5toEIM54HF1R9xj
7bijVvLJcErV14q/D8fD+FTTztrBE5ljtelStA3R1B7JeLxocvXoqOsjaNvwLzE7gio76NH0s8f5
XeUq58Jl+7XvMj2cQPkowWnBcmBNN0ouQQ/Jh2T0CdMlwi4r4mv5xsorAi3gOEsyY/hhp13WONEB
jYuKiAagx2i74UmawFmWvZt1WrZmsTRRrx8UJleqSGaoe92p0txfeB9lIobXCQu7Rq1UJ7e9rmxr
DfEh9lxP7Slia37rHk6qhYL4oYZAEE8vSckKyPHei4lag7qLYAwqNcR47RG1SX+b+8V20ZVLJ0oL
8RG2CE2dWYwrP0dcQkpK/2jQFjcuy/1suuKuF/rqQOZyC8d4xGbrz+x1Z4hZUpglYiyCIb78eZcD
SxeDgAQO/p47KqKMKByRjh5tacXjGjaO6gbYh+6DfJ7Y2nXLOghxGj/7Tu5DkAwxe4cNnY6GBZLL
4ZoDjTtyuBhaLKakaVQosdbcBYYLsFcFg8bR51hZ6Jbftnw7RMWvd2wbDi+Sv+3/dXUE2ynW8zu+
bW3GLBISOrDU51mvI5roSzOKpzRMc1I5TAIU6MDogy0iQVXWZI81z03uBT8tPCZAu2PZGeI0bifC
Cvei8l4pT79cUPP+xGHKlqNUn0Zy3fPkLhU1kMLpysHR0ImUesQjc4oPZe2Wjj5fV6Ums57DKaax
7MANtlNlhamLGcAQX94WIxoNaiztkPT0nO8ULRztnu6Q5tVwAya6UD+UfegObU3ER6SlqKK0/Hx0
tc3Vo/ol4VduxosCyICZWDe6WaKnhznpQmmJyjgiLLeLBjAu5d4I4FtpY4yWSRC1oCDjUbHt99wP
3dWKQnhOzIgwb2O1FXYokVVEpRkhefULNx/IALraAwXQAru+h30q7U+NPwQDjeraflFNvFQCRUJ7
oNlSpsVANAyKNjsm+PTeYg1EAHInTqwqdWTV5RThzfayz8GXlk3N0SXsRl4nisssgYrVu19r6Ay/
jQhfLfNiGvkU7XZlCgQZmpnXMsjvLocc7XTwWWW4yUfWhIWCHntrMahBprDQ0smN5lvLe4dR/WkD
fzf29nWeOHkptZGUlwcVKzwAi+d2HD7/0z5Mh993IkRDjFd9556qqIU15Lxy7tRNzj8bVfM4iJ9c
ejUy6ol3DqZurF4pQc4uVela2/hC70PnWE8zkz6MWAvHbKA03nENDCsuyJgJJFPSonYFm/1Lgktq
1/bpVVCCuiQ9lITdeXoPX/N7NERiE7HbN6wPxk+wLICNM5qdjA3KQdJX1Oobs5PA68lLET8svst9
e/T/F2OOoicBojW86KwxdEfGOj35PGSvxk6qCagpmf/shF3FgenzN/xIcMz2LJE89VdIWDuWgh8e
wC3Ed68hV92q3SRLQHlRHlpLaKKjjj2SqE2qWIYjqYpGWxnfWpXP1ouelqKe0zq0YISP3xpBkiqw
SepYl9FyZv5Zi0KnUWObTPCN3JiCOFY+MVw8MBugvQmfh1mnWHf/At/6lXirnR1gMsvaCMvdOttZ
IKjAZI6PqlTtAssTRMHj81nycoepWW+Qkw68mY5HO7yQu9CT38V2vxA7AQvkQ0UwKsaG8koQpiSb
+/6uwM3D+Gla/vAS6DjD6u3vYyKs/jonPHJ4m/roBzWvWkc9pdQn5+OCVQLdNj8iWjDckGsKhiBw
CRO5CS8fT4DYBMAuZ4S3cp0eTBsrV9wjW842Is4JKv947LO8RSOgB21il9oN99zSdPFxX5Doy1Ma
klRHhf1mjaQMaPzhjc5tUPnFRM2AsPjm6eGiidpMlqIZnPZznDBWgZlTA8fr+3pcwTY+zX03RnI9
doJ/mqvvNzMTlpWMHKgcCB/O9969sy1nl8D2K/hDBkJ+/jX0uqEjTK3TYO0sv72aofU6GfeCMQuV
qDsD9YmZLzHPrCLOTisBFpdZgxqRBZRvHCbpD9Fu0lCqHcezakqMo4G5sqczrPmrFg70HsBzZyHT
6w8TM28CWjlUr/7IgVg1muUPosDuw8RiwxDGQu4kN27AQVsGy9FWzn+BY04dpInKtzcInoam9DO7
naVH6PBTgQVnqxH5ZJX/IJjvRHkkZIfSeuY9+5d55ppNGdqH9jK4cMJXSefppUJqAr3IM58dq2Nh
ANB4/PvQ+yLC2um4WCKTg4vnJRHmvGnkngR/5fBEYrAOEa8H+LfY9eqkFdA4ZxFqJz0CuzK2tNxz
xAuUm+4qR+bRCuAcDY3+nrKijMs8tB5TehqCUZtCgFacIAklAYAB+25Qtn5bCnFLN8xOm4d0zGYy
xqRjs7xeA4hqehI5R9hti71Nw9h6wQ2cXifWIx6vVj36H1lNLPVvkemuOaiO/3zvjKjIRUhunQay
/k/sHX8KrgcfaYqJc4Zf9eiknt/b2obBvHNqlvGthzDKlOAhLaZVaQalzlNCZppX4oAK7/TJmiaF
ZzZbWTr2UPU2spoUF2AcPrxNdi2iNcXU+Ow9o5dCdSrbAJPhJ0F/DUncnXNfienl9BkiKzvOIDZ8
ct1f02NgPOn2ZfxH1MpDuYYI31W64nPfOz9NcP/uSkwy6/L+1lo/7nvDzh0D+Fo/JbczXBG0dlwI
hk/ZWTI8zSxp2m56KIWdYhIMCA3KG1afpIZHZ1Dv3ZJvDr1MJeijN87pMVmqQ0x8BW/d4cb73n6S
fF/MxdjWLvb+x03vo962zn7QRTR0Tt+ycNAZgVaocXLWq+EgwoAchXT+Rld+jvFxwc7kweWQCEAt
4xlBHOQJsilgf4koqP3WAv+V338rWZXWuo4hNAfs5lYoMfOHMMPDxwYe9/IrYZxaLA0SYdSUI6iS
ehDRjq6dsaLogCCPiLM87Il2X9ju5RRVi5c0sYzvqxs0jZhbuKYrPOI2UJv8xRhxwOzOZo7ezz//
D0ULfiyualxzlQr1XC88Rp0GBagzE8TXvckvJOBF4z++xV8GRQAepzcrVaqeFnPkuL3ayqwb8Z7d
WQEcbgCiL7y3whHIzZz31ypxEQbyTVi8n3bQKRouYBvVENd7sVxgJQZYP8GqDnn1LAy6WOk84kZd
/lFw5S+40ORkcqG2So4bactszYqZyGt7b5I5RyF87/GA3OWKhB1xdhHnfEYjx0Eagw+PnUapUysi
6BEiORmV0ZAHCAu1on4O1RjFgKP4Uy/xJCIZ+Q+zfF/JlJizi8K9fZ4RVSGz6vaUA6ausPG6CoZP
iDTUQpgEU/Jb+kITjY0QFrZ8jqxpa+vSPM87ZZ6iPulcu2Ry86Xvpzetrn4R4RX/PeFxTQiJf2VS
NTDYIKuw1fycj80zt6vCoDMA1z2uSZmAyVA6xCpO0NnS/sO2K8LbvExqFHt8/hHDaT7NJJhzqCgo
9YzK7E4KhJZRLulqmqRl9TKlZRnRqQwSqBPGisesZTr+rh+gsb7X802Px++KDpnOURjJD6jxzwvf
bAVhofsmZTdm6sTw7AoCK6JFyr51863/V3tZAc6yH3PHL269ZbsTX1Yro25tgvPy6K0eFhtcNUhp
R1Fm9X7EzTp+6sORkgFtILGiqBLVe+4uc2tWwS0y9IcRt2gyY6KkcOT9+PnsMS/E++yoMJPBVcll
pGqLpLIMWPX9D677GKI5UtFN8KmscukfBL6ZkDnGw7dnJcdypWRRPd1YNvhFd/J5jq1ztTr5DJiU
1y4r6Kn7ivUMPTxI5309pwvcd40Vsqff4fiRVJsk75CFfWrEGw8MeRHVHtNPo7XBOGSumGbaeJ01
u8wnC4hQcFhGwgPvc1WPcRASw9+kCwvyU8TfWVxpiai8mIrVq18WAivK4+8xIJbjCDNUW0rqPEp9
l0280+0Ar0euFyfPKdy5FFjPkPHMXkeQFDEWwgVKSUabcDDnZAFin0hw5Ub4KC+YrKK8kjfsRBUo
VprVndYigzLfG3xQg514vnywawHVFIVxy2ohu0wAqpLudCPm9QP0JVyk04HfXrZmR2jHd1rrFGsq
pFLMcX9UYOmdj6V281OlMDLf63H1NbvnKHjP37M5myZVmeYGYFgDSPtBNeX7zFpJ7J7gNNtp1USh
EBFkYNd8ow6HIXV5nbuViDUaD73l/pbXzKtnsBDEkUAEIP6czriy9K5r7qUAKa0rFNctMcheHpuI
N1Vcg8VV6U4PvhqGt+tHEMkZZbxYEBCWt2l0wSht+FAQj9Uaf+mEBvzEcyxZUPfnM3TZVKbUP9UM
gqWNnsmmzdlHQg/fuOKJsswXinDvmYK2AWNydiZa/F+Ed5LUNluwXVZbAcEdMRNoq206XMdJDNil
q+l9ogrBRf2jP4QwVwz6lVj1bLr1VQ5bCVz1BKsIvFBkF9Aa+C91lbEPHffgAHLza9+/cbwG5Gvk
wWA/6oqfdayiYtf8acpqdIkgZcQhMf+Sg/FyMkoLtgpwf+pe3AmdSdu2FUzoJc+ZvpOJqiK8WJQM
mEIXivbeuAgBSgbeEXaFoZimsBcz1FHqut6NaUKjVrBqcW4W20A5d/HbqQ2RTlw3Z81sjEXxxBgV
pVrwM+MFuhMU3Boo3A+l+toOVz+SQNw7LYpFQuzV0uhw58Fbugj1rOmpzBEmKdIH6ZOHEmEP9Vfc
n6FXl94f2mfGR9QfmpvFDr2GrZ/BgO5VaBM47J8LsJDDLgZ/1PI4L4rG4S6rIJCwR2kjroGNyjR2
gdUN/rPZM+bggDtyUmgUoq5dFJ+DQFkYIuJLjqAr6BF24fM+JW+g1UKHdB3BlBBiEaxYgdMbL3SK
TH2bkKJWkeVigt+D98bOJTbX3LNkNX1jpdVgByq2TX9r3OISjRwjOCz4Owcxfjf+HhvDCQG16iWM
qGAIicMNozZ1857iVXhDk06EUbeoxKkQJyC70SzgQyTfWGPEXE20ClXt9Z1cMF7bKZzFBEl9McC9
O78pS40k/bXtNhNp992av2tqG3HHAHamhLb7mIvVFHg3J2E1wfcoRw+DMfEp8Kmt/gjw7fFHN43G
eMIwrcYpozTaPs5RnTWh/aejUbel2syhGAQVn2HqIWAMjLCJmMqbqcr3Ev/lTW5AjeITWLyoUX58
ReFjfhQ64DsviiYUChNJ4r3jQjz0ZoPJTVfR8bHRWCKgTXdJFZLq75wlwd8otCRB50rfttfSN0FD
2T5goXHPSo3FeK1sWbSRbZHLDmc4ndYzmpeGb7k4AnMfpXp6lsWSRGed/7cwE4gjzeVKKlquwhtO
8DwnC9otC9PGjpdNNLIg0M4DhFkGJG6qvz6bMN8BSfraNk8pniOp2sENalh7o/hCUkdfNi/pn8it
7i7bNRch1AFWauvVAOVHsOOToOt3eiZmXLydB8VJuJoRqZgzcOKoz7FCnIxyh8/gtGd03HJmL2lO
YN2AhgWyXlMflrPsJaRJi4qpAvRHZD3+ipmO209AnbcoS7dTKkdasPVCGsTG5b6cW0WyuzHwP/SO
OuGKqi1lCRg0ZJO5RAvxWpiSuVXHSRPi8zgt3aNCROeHT1JvQf3d1+szP/U0gekpeFKrkAPuZoDk
ch6JBxuhxigOfLwwUn20mGOo7bRArT8ys16j444IY5XMAZlD+juqjj8YXsPjimMwau88zmuF50ha
jnZiD2W2k7NOHAJoyeahSZuwgD+NIcNGuG3p48Xv6KoesAVUSkERc4Q74xnE22wE6dVhyqsoGtPD
jzLfYkPbVMnwfTiVkXy1woaHtXajZJKuxOL2w6Gnh5UxubCEbmdUPZMCL9bcEkwQFEgbl2128z9C
4ax0udG7XZIqTpaSz/2hjRsjIn5nj5lP4KV+wVTBjLg0SX3lHIzJa+RlbbJPT7tXrfmz2/WYOqXz
Uy2gZg5XZzZCW2IWApOUkhoChJ/zgHSYE9oUF3a1du+SJWpLszrdS2iEgeRCJEE+YiDp6vdG2Gn7
SKyeZZT2JgGuAYx1sVWz9QheMivKo+3ErymIzOLHMAeCj0Jmk8KrIto5NTR3aTjnWI4nx/io8/0S
2PlWKvFuVhyhUVvuRhsFHEBh2NuTudtYy0aO5naihwB1u6LKHf0EoCuCggY4S258ZK1sARbfg5Ic
ke4l9rLWujNGaCF9N58SwaPSRSPYewtkJGpwqAgT/FF+cEHMi037jWM04w6fdQiLwiYXZ2iVV4Kj
Aj+lsRJPTMHLx6oyACwvQQ38o8fjf0dPQ0+fuEkv7SmsLbMs/GwQGlnyFmzmrRDPdMoalqVKdu8M
6Bll6pdxEjrzjDWaIIFgs9a4CIO28DqFmjd8SNh0Z3+iGorR5CMjCBcJ5gHXuorYDwObI/cazPfq
c8oNAxyivcqN5rSrW/OMKAF0OKiRHHfc5ItRRgNWzA090qqP4X2tWBlIt1IXyyhovXhmMz+bgRcu
cRgGoN+AqwB55bNn6Gxn+JvRqdgLufNZb0iGHyLNItlWXr4uxTpLU8CNKkBuItRQhV6IkjGr8lkN
T3laDG5G5FqQxfHCBx+hByIWlwbG0X2I8vVtAjgP4VV4dVVFV5IhorQ8yZ52C3t4kv3xVjjWNaUQ
bJQf9FMzLwy/7Ts/Y0NIuEx2NDMOnsjvaM1al00zXe31qRe/jr5gN2zwGuIiu+amdkQFR79SF/KB
2i6qEub6mIU7qJ8d/J+fozNGEKU7C2T9T2TElMEEa5ICdOYnSfEBr7UXLPopUokViHnoFlsOZwUV
bHN6+ypvuxufSx7pA4dvq+djGhhveC8tp7KdvMRLU0fSJD1YqCKQ4Uo38b0qWWaU2zBWGizZz9XX
HlwS15j2E/pCXHjiM4HAwkLkU82wq4Yk1qYshUzi1iNNa2UP+RMhouStMPAkFLg5G8E/IybtIVjg
A9OyibBRnbRX3ieveAbgX5hySPXLCtllwfzEOvqJwZ2LPVNfkRldAovnTw4PLAzmImCkkwRygiSB
6mNRuGJS7sonk1JLVnM+5unFvo+Wa5dkG3HkqGiGi2+ZpefvkMjjisfaqCjR9UEEEgLEJikAZPYQ
qOiPG2mh2SWKBYpAkRKOUA17swAFPqVPI4cPYHcadQC+NMpMeKHDHV1pJgzqnBX5gs4tGFfo6RR8
089Xm/GkdYJolf3ieAzCmnDtqZyaVcn4BIQ3+bbNjg6ka/e3aGJR7bD9eMYToqEL4bQena+XT64e
/D+xmSHbFZJ5yAamGlnTS2v3oVvX9o7ECZ7odeQWQLUzzKml4melYc0SR5tzLFnn/IAB5uQS3+Iy
sWOCSd8s1+zdmAnrWjw3szo/Kd9pdXdWIWSJk+495rZGATvV7LklbUs4Zx07naCiIC0oTnWzCvs5
lr+wOzylg2vkiuWLMtAN9QqbpS6Gl6rpu3VUjSpolFYVLJonW4ZBctSFn+pXFxcIumhCLw8FXwot
28Gi4NsFmQiiatXiFCnHtLXM26MqUH2zT9Peala3FecDE2rWQ+RDSXgFNO3bZ0Ae1GxUJ7UdZIKZ
ZfCKCnllaPqsqkFbkVcQqS7rGAQn8REcNezGXgCXN2uAuGrfhWOLCfmJVKwDY847Zv1MudKS4qgs
bJ75JA48oefT70RUpuCC74vXrHW+sreX4ZBnTaAfcTk9F04IbHw1JKlFlj9zG/zkNSQNCErB9KRw
evdofyowgCOtqHarCx2nDrYVDiKiGUJPorSktyLvbLgzF4rAvf+S/1/QUi2wl3SRjcpQJAKDuUSG
XJp2NrVshuGP3m12bMV3HPLRQE0h5d3IWwuqxPrA2YGee4Bra1FKXO1QWEeKJMmmerIxOoVjSqjT
wDPnrn34YNK1QMrpRKIgNZDC9FSf74pWtbY1zHoRD7T1hJAxLu+brbEuZOutk/DP0CIuYIRzLAEw
jn99tbAkf563l3aERzZp4UtHB4hGldan008NEXGzqKDNrMtNG7PDwamN2elFvHYbdAEc55c7a4gF
ioBv4Q5GdS43R0f8OeXYErKy3Ypt+Kcgr06A6bz+WLBI4q8ExcM+1uRotIXRFfBGN1zElQzL0YxS
B9X37LKo503hjZ3T2n4+q/tgmZGPuR5YFW5RP0bBgNnKlXF4NV+bzUePwDDpegvfQjHwwIGgU3fw
ulmPecDZuV3ujLF7PoAnM9dIf6I5mSi5mBOzCSC4A2jsbpfaDQC9h8BYZw8SVngidC+kcIoldx5c
spEV1/W4QPdqayn1I9/7f+Ikm7jzxgN7uYErpSkg28P9vB1eD6I5qtDgK1W9yU8Lp9sjBtppjefc
Y2R9iRx0FG3w6Lgspy/xYnLgM3KjYwDcX8q+PJyQfjbzFtJL0bkpIy0DY6SsezWjSvIKOwxdeMrU
VCNr1Oj0b3nOI2pqi6L4zgousrBf2uZ347YGnpi1a+Kzk0a+pQnEoxTc4OxrxDswyY/8By6mMYYC
7Co3JaSkd+CxeleiWaCi8gP96qYqiH5xM6Oz4UT292unVvokFmiLg2VilN4GmspHByX0bwB8mIdu
HuhOMUZgK90ZBSHT+LY2KaLc7xd5GBGdycFmQ0vIaM0TdqLV2s/J9132YfpcZRDdby5yVXjyMKf7
shsNwpKa8LBC0jgjw3Q16tyA1tv5bnD13SQ+P1ZdtW5sMJE5pVn0wG+ggWJXWXa2OmYjNdWPHzyn
Vr1Dy6wg1bXk2872hnWyxFYsA54maPYHICT67n31Jbb21+E1yXftLUM9IQyViwOIXQv1lib+YcWN
Gh18W6ViAGCXroEcRdZkGNJ+Cf/bgll8tMlOe6oTeB1is9xadGy76HeKJ3Do6CzGEd0dVH9Jc5NW
JtjcLEjXaOUMvwpweaNc6vPRBJ/lmm+wn32LKjRsHsOyrhjyMgbYJBvza0IejNtH5bLf3zIJE3oa
0RrMxrTVg6E4L2Rp7LK4Xuem+4DwSDcRWV9U+xPZPYEEOp3COfTaQmFNOLYxOtvlvKHQlaFEbioR
iRszqaA/vuimpVNFV+bfKXpsKZpxAlMkogagPfjbAiPsJcDi/JC4pKHPJL+6kqQfvcM/qTEUpjJo
lp9DLrL1cJO/8ifKhobXLgaWXixf0hHN8Nez+43gQBot08PP3jMCIOcEO69/kv4eP+jrbdKpczDD
bfRUK1/Di08XjUb7IZ7Gq8H/ezFGUNYK7Ku+NEcRNziX2tD3h+xErxZcqRqqMQOrPHdOi26Qlotv
Csydi35nbwYKipqPpxcnxNNEZLdhOcgfdvBQ2TnXNBOV65rPBn1Ac1Cs3bLBz4kAnqMwqFy7Yn4j
h8AXoSBms+0WoZnHsNevDfZmoeRNYBrioVllpVcO4gR/hjdDiuSGfJYwSaz9a0VjQjqnJcCgZ5FD
bm7KNLIVNHn3g/tA7/YOit9ogWtbEL2Jp2NJNtZGYvAfUxjF0Gj9lBAhm8rqRQqL0tGulVviZvxm
93eCDT8z7daLgaMtXsVVgnoFNXzfHUu6kpXQyE8+zOU+mP5ZCbnuoJRnKZjc1c9GHcbnex/iPBoT
0fymmlApGxx3xNcY8+MSpnEOkSWF8z//wRdbZJeFcV1P+uhzwuSuqsTPPG93cWU8/pIeM2J5SWQr
y0qD6dYb7kIBqiNAmkd746o/k2SaqY5FYLTDMafZ+GF7Mqpu/4SJbnMliwY3gdfGtcL2XU1W2lM1
K5f6J8CjYYJ3yTF7IiwaJyS58wnaqlzEFzUdnEEcgYdGPmZ4RiXu/ki8vgzSjXtZLPRK/PXdt58h
V3dCcCdIkMlc3Q4B6XFnKik/bzV98McooO7Fxnu5ShsIQUro0FKIQoiJ6YTKHXLMJAUgyf72MNBi
5pFYinL/SxbcyG5EkL13mQIdrNznasi4ho0k/v+sbHVv6JODJFaVOoK44qQXzks+l1MYNoe+1RHT
9L2mkaBX9pniMXsBS4YFHuzoDVyIpkpQx1B5mAhWl5f0b8Vhx+IQk+bIgtzGPxnVWtsyQ7OZNCKm
Hi4a08zLJW6yfhxcjfYi3Hb4cPO3YhYLZd/tkO1Dw6GC89Z5oLXaggYCpS904VVqIuYdokc5JCB5
vt7FG9Uwz6oSQm6lFeKWefEjyd0QyT7JD4OI4E19MjTKtFK1sSQN+Dx8bBc6N8GDtZ6x4Qd5DMlN
dv/UMglzwI5rfRXmOEGrjeepI2RHq/yLvjJKDGLs0J/puJBo0RsZReTBnzdyKAWxE1Iz+JGrW7BV
NA6kw5fvMSytY4RTi3of1xu1r1E9FTJqcBgpqmZSvUKMv8xtiMaC4A3jslPH1LzUFD1tbg2mr6/p
rMK1i9/muw8f+8sOgqZFN2Hq/HnpqK4sSPFodXdOqS2rb4oLB4igGf7/ZfMCYpEcfc5aLwpHnmwB
ZztlG77tAHn+9GZhuT6kW2FOw3a8QJzIEf0RjDndtK1O+naesPHBD64KDcm898XXeGh+ZjMMM43N
noJ3epi4/ILX2N2slquMje8m03JBnn9xZpp+uLMBigoEy4JLQn3jne1Eo9lpteXcn034EGZ0r5El
SQNW3KCi0BHrfcQvErGbzGQTAmXsXgnv06gHlMzH/2CmGbigsoMqH/n1xtwPgIzCx2nYeybToMJq
aq8+49TYpiRFvOMMMQ1hD43I4GNyR7MRzuLXA/C6Dzmq5caLbsbkysJgDannmlQVdDigzk/il7u9
kR0qnVpdWGbMTIDsBdo+QadLrYVEpXYrn6KdL3w/RkcETYvozCKU+LksBTIz7rWQCA450IXcjsCS
kLm9cOqXLyXCG0L/6RQkdz1D3mSz2s9oiwgk98uL+sIcT0AiSJ7cfnoU2+oAdy5FlBbbHOylhQAG
bfkZs8cS4KTvY3WoFXthfHKyl5dXI5hjNtIn7iZFmrQpVtkgYZlzBbGgeT6DgilqHwJ7JymyUJr7
XYVT0hd1TE2shFggXYUK9wfdfG+nwrHpU5eR5IhHyJWkhuAERi8g3w5DD7iuUX2p35CgzKZ+RpSc
XiU2PrEGl/uTRyweWsX/arcWaVtSwnu6ZytfIS4HGeOh/BPot1MIQc71CRmZVkgLlYHNkirUR+kJ
p+NhCDW2+JOpZ20Kue4frc3jTnNMhgil+AaQZ28B3l+LhqoxHgWY5rElh4srSkWsy1SEGsBgF5rb
JOom3xnxrlxeKc+Thh+2esq4fDNFr296VJH8skjn/ej+fj7oihJyfAD6YFuHOHijSZZKFXxyo7mt
Ti/CKyDwNrg9caQoL5fNlcMNANDXzOURqreUx7qqUuL/0DmlAfg/5EXu5+3mLBN15q6J6qarLdsT
xf9/U156iZIf/UaW2mWlqjJbGAMGjjHyR8W9lVX7JWE68Rl+rmPv7cWT48DJfx87RG3jrkSDe6mZ
s2IZBQADwZgynWqfoeYpMXO3JxuuBWGR2vkXGm5ColRcxyUSnSk/KNL1Dxke6jjeRE7eKC6OWihh
N/puL1oFGZdgVgy8I/Yrs0FjQR610YcvUJM0C+AtzSa/37hfhn3FCclfalbX0663+Dw3Q/JyotCn
UMkCxIFuKiQGt0XnOJDPiDBqus9sk/a4NEOmVrASGHfHLVH4X6/ush0eMlrn5K2d4bFR394dI0Q2
AH2rjQmT2V471qVpsY68memDbKelMzWCRmNVGfppsc9RNYslEi5Wm1CLtx8kr+hQFJAF67aJznX0
ndWZaiyegLW6Y9JJhONgBxh8KoSl0lYyeYdbrA8RI4ViX8dw8SjlpN6hADWSjBUlQvOQSqQLkLIs
1jdRCMXTk3gld/0yzIWAWNNtXzSDm9pPHUoUbkxX3CHvnhaH2vIqS7BHxAUMwzCoENORsuTPhoaZ
+DCITe22XNJ/0EjOlyVqPQ+Ujya2Im0Vw570iEtgZTTntPjIbh7pHTMOlzx42J/kpCp7OlQimCyj
g5U4ZJyf8DV+VEhnJ8CScx807zuQFUP2MmPj8KbjlcikhJX1YGxQ5xlKdQbHsr3M1VxUmnMphPCn
RhI2H2U8oVCNT5rGsciRFXKmsFYCQDehaJrqmbm4f+AO4y2SzC6mfsyQyIGj3e+FBSN3sfoQiWQK
90AZQPqQNW1GDjCbmkTHvHA4Jccl06UTfuBPDRJEZn5fP/eJbShXFNjYT2ilIo+G0lu3/bJJ7yZC
A+4MWhFb4gtLv70fIQswqpaOXPmezrOaoIbP9ClLFx5H9v18cIy5K3V5RpQDx5vLtW6sgdstMRHY
ZInolGjkTaEL/eT1kNOGmmvk869kN38PyjYCb5c2TX3kHq3Ussi+KG2ruhm2spv+DCh42R6BnwHs
Rzq55CGYOwpyAdyPmlfqfX9H5wbAA9EkcXZmbVa/zhvoh5OJFCX6X8LLX6K1jMuXZJm8hFW9z+H1
tukiDLhSoU8ieanInhXMn+jOmkrhC1J3fBaXJHdy7HlROvVkTRFVBeiOxPpAAXiAPtILNB1L33bd
pxHoORS4nOVr+iRZ571JNIQgJUbxuxLureooRpevFASUNJmGuH74qOXRsTuEOfUVF6xC9RW2myIL
YIqLWoFB9PyEfwm5ZEoj6hFZDBkfjeVWCERg35oK7SVFk05qVoOV2Bigp1KxU4uQiSvb4JdlRWep
NQCfRG4fx3C9zdjnkpcgsrUgtrCV1TeSU5irD+J2q5RcqE1dm5iyBH+TtUY9l7wHXeoqnRwucJFd
8IbhyxrP7uircyi4dZUW1FYLIt1e3N4DrMjpgFF18yB/GXHVwXymB456W4vaELwkHOpCoVeGsUj4
sll52bdzIslA2op9DR0bXm0siVmbuejwbHyK/zRtGyuRAVsErhkVOyU1M9EWcm6O7Eoha/+kllCD
GHiAoAEMGK/Z/Gbi7P5jgckB/4GDjwYPaeMouIRuZ0triahQL08cwMUTDaF2ZF7F6qEnEzD4v74a
jbrQ+YxopMmmBIyrfO66/ulj9/620+5uX2VTT3fFSJ+lhroaDzKq9T1tKOqNMKgfxHFo66Q0LrBv
BEg6IWK7XHw73JXeJDERwCVK8ZQSD+ePvFRMN7rZaReL9aLjhs9M7BFvXxYkgs04bHqP6rZYuHhD
Bdb9XLE5KM+kFGmdq8up+/1gRxeLyVoC8LM3PKSSZU85yp6oBW2kb93Fxmr71GWbgX299c+68dVN
z+1aP7qg4wM9C+HMsl/ekgTBKLKyMHLKtPUOxd+kBhaKOKJGUtoCwCQmU7F52Xuljqtw2N2RDDrp
YdiJEDd6LrH+B0YHW8Kn3JN/Vo2yUQuejT17XbV7UYpzkOJ+3aSRsdby2Eho+l8h4Kn3Js2cSYMM
OHfa9h9XYs26z7VZOV1UcJw9UQC61LzlTJV9jV5QojZOAvsVpMqOFGfTcjMVkKYiqtQ6CnnJUM1L
a98eajQEkcG7Fmz/f+tRbkpq8GaoDXh+DZIN403MBPlhZEtrazq/UK9L+zcIwHeCYpz2AJhWyYCP
msOR0BD8UfIM2AqTVC8JdIGrSMiJRGyp3mURFVBiyNW/Srz6bMF55mMv7c6RgKtyqXDPdWIGbYZZ
H/RFtj4LhYC8L7xHGRFVwkWr+G0a89xqucSbJNxLWDZiN19YEMJazjvYALiLb0/3YXO9v0CnPpfq
z4N8U9/2fHy2Ehg9HBm87zUutDiIjnoTj/8oEM2dG5vAOrqHRSc1OQ84MNip8LNKZQQOotzyprH2
qMCSpqyXPrUQZqn0SfYglp7fZWBFxyTAYP1eWr1CJTTKg/iXZYmr0L34XfEBXCR0bbx5tomd2zT4
QF6zLdQU1Fv09m5GeREvuL5pC+0USnK+e9j3mobl75zW/XQaKlOrUHE2uCFY+fm6fq+1bKcsgUwA
xgeuH/M2dP1a/2UXBNdxGvZkYmX+HjlSF4do7fm9YD6X+jNUmALAcM7u6ASM325iFiYaQumDBezm
VqEmVAMI6PuQ0vxu5Gc7JY5VdaD2Fr3cuPnbWqTChgxY1du04WIfc0BF+Zp5kyCxh2XqbtnpvNG+
VaxNYLRGKd0Cd9XfgegSuk29bjGwB0F98HcqE44QQkh9tzJyxEkm1LIZQ8jiydLJh5gisz7vz/HY
C9VHyf1O3u9HCyFKj2VUD0lHB+4JPql4e0rdTiIwRj1U15or3yteLnddPX8YIWgCc0AO6CKssMoA
ECI9MA1vl8SBTn0pfUYb8h+1uIapS4KEf6T69oqheiR7++nuiR5Lw4BlSkhWjBb5WsTJy7TY2KIk
qW5lZryd2Pm/w1z42I6gLY5zOtaRc3t2UplVXPFoEA20HKBI1s54kmf01ldvZOoOkrcWNDQkNNCH
Sey/KN2VwLtKpjcWElapDMOuqSCuNwOxBec8tINkrzrloeaMQ4m72pmieGiLc1QcD9EsOwuehw/v
fuHJXc9GBTKI5wbH2veSt5QhLwdWIrHLjJo/gfe48/ANpnCg7peUYf99qjAlUdLxZHc9o7HIrI85
2SjbxmdDeXhTTYUnpLnQNGD07RnrB9T0BzfWc0rwWa5gAWRT2GDOdMuw7XAJ0FrbAHE+BvzbG4h9
tBJvR97BfhosLQk1B66Bd9KM7CL+W/cC/WWqB0js1FocQU3hWisPPfawcn80egLLy2PHycyAqSjb
bYKM/nZR7WUC4ERHhHeVqVMHYfPA9NBxfZvJKaCA66vuoRN1HbLhcqAM1oHancEQG+bGzFdTL6wZ
T/VAkkALsoUja+3PcmxNODD5YnQDfL8wVzhpeWC0K/SOg+RfZoLt2Zxff3F61OFpqkzNzsU3Pgq7
CkX8/MdMfbkG01MNYQVGChywFzSrhkGSmMavrbXKiJ+p8GX7ejiuD4ZB4/kH1UTPlluvIvcStP08
KBh4RXeZ2ru8F4j2Kn0o5S4/uk5fvVqzPQ6pEBkGzqJHGV+N/2ED23nF3xaI4w6E7UUWzoJjlKql
tvICzktEnX/gStNUJSQuwGhDiQvz3Eme/nEFWcXIPbf0nCZ+1kw5S+QxNSlqkdbTXTScsx/YniEg
ri18rMQkuSI9NFBGdMs2GGMooto5EiO141JyMVQPkW8I+BJkBEPCt6zVJOvR/cy1pH4s93DRVeVz
T1p2TON9MzcewIzQfTijvZv7BwQXqO5GtviEhtBovl4O6ms4D06UzX0WiYRqj11qFjSrFqU0KHmC
qsbAKJauyD2K17thckry9NhzY0mbXa3PoFEA4WD9b/VM+Zl6MWIRcMjpZ0tIunLmqvord2+LDeN4
y3NXPF6MDEO2XP5hqDipQgNpA0BOkW4Jnunat7IKtlfCfWjyHlv9iuIaqliXWfqOfqrlV+YMht25
ZNhF9j9VyC6D3S29kblfD/aThAVHaVMc0YDkrO9pWx5ByqJ9w+8DJ0l9awIybHkfJA1vvi7FL63f
taAKFBtPhXlJPAMsYJ7cudzodO4Gcm+CSj5nM10xfFDyQXAZh3FKiKHrSKqiGGNjRB3Vy63sSgfw
fqiFH4LJjiAJ++O3x7Uh+zMaJ/igbYsiz9/ijCyFG6tSyrGEJttrdlUEFBfKvOfzHXoKHUq9Vyui
jWHHvB8lvy3jnY2hNi8cp+AW86bsoRlL/rKnw3+UWcojmvc5zbxPkUjmQvQHCAd+DkQMsB6DNcMw
N5V6hLq2otIwXYQ7Bn4qWf4bKBymF+h1+XxaltBjJHg5KfUpqGzuotgFNcWcNFp2gf1m0hEd4+7B
JHVtktS/nngRaXIslUlPExqxyJd5cwZXxVhZ1KfXEnXibUcNeE0vaV1xCoBfRLoZx5z+EXfxTJhA
64Px4EhTSOcb+Vm5BnO4/vgStX+xrAhRglEjRWBuJlzwVA05KURT+M73rmhTdtR3TNHavAEcPr/m
XoVziZFhujl68LM6JH+Ehc5OBXbcMol+LbF6RQGtsFq5kCLyFHl93ftDoRtnu+FgnbjtoX0d6npC
Ix7P0IfZ3xsHnupErmOtsB/lgY1NybC4mJKZNCx3Z5RG9EzDc9baK5HErryQR3mGQydLHjxMktsY
vDmxNAyuToqJTLf9YS3udLPmQNANfKbyTrrX8XyfhG1Z0pm7LlEaPqmMGsBaqhvLgLNsaEAb9NDc
cViinFnQ3SndORNkeshaMKrb5Fwjif3zA0WF+6XI122pUCxiWzqTTlaWJ1hTIFEqAg+2cFbiUCMs
qj/+AkoSgGKcZsNFlU3zsW4sJYW1n/u/xaKHGT4EKJgcPE/sOumRykT7Gf82r2vsX7jdJkALPBOQ
hq2NibWZwDv4oQuPP1mY9IXGDjU/pdn55xqPfVzOuRidjwtg7w1JjcvABtjNILahNq2WQbRRYDj1
isVU5C6Atx+obFZ8HPlPTnka3dqcD3qH5nq6IJeHuP7PSq2HPrG5KQLaSbCPPH+a9k3BAwyWjsCf
oWh/dqjmdL3AluSle/ea24WfoAHI+hVsBhmphF8j4xI7XhqTbaoqwVi4P3zA3/GafLTM6G4VVQ2J
53HbmaDueFprYp5KXXF8rRBFbnYHDaPLSKGknR23VVmeA2+JLnHiYUfwmNdEuMMAAgUnWa3Wh43q
4md4r2ufubuLaG/kiDGhTgQo+s286i3+dr3MkxiZpD8OlaCEpAl7JzGJTCE0lUMzgBbVre+YcVC+
coR2j7r2dZEjysrEo0u7eK3pqaIQoBiReItTg9x9GKGiU5yj+TEia3CXZU1xXjKm1FLiHRpUlv1R
b0hqHs+Kw/FyFnkieD+r8D9gjfITZ3X0RQ4KxpW243CdpYK5tq0Fa/YPQom4lNLZrhQOHG6KLuKm
4KseV8ihp+NcIEwe1nhJ4yxQCVgUnvCdlpYW6MWsZJgM0tzmxddFufigqLIarw2D4ySzJT2y4AGf
7rIcdX9Qrtha9+u3+psLVfS4PT3XD2k7E3Z/x+3cuZMt0TcA4JUiFCb7kgY0AUUgheFwhdMnH5Dq
g51jSIq3AL7uHPUxu039T+Tkp2xZ+gwrBSb8FcHLp4jqhviN++ETF6nN7hOrZ5mxNAcu+mpwM5tS
k1g7nP3Iu6baKGeCVjsLU7GrHelNkoGsnNgGOQgNiqm/2UoHgQH39AXxNNbutnCxQZoajQjurDWN
vvrw9M49D9FA1y5usDpsjmuqv/fV3D+QOJErvIVi7UATCzxS/a5g22AUMIkPzaaQZVxsdCbIogcM
PraU3bJ5nr9eJYvs6ip7juSTM5IFj/s27OFOdOdUd515Sux/kH0c015gYruEG2UwfhKNdoWbW/jM
1KNnzsHiEL/urWL1fTuf3/GBLnh2t3efPcADjC5b2QHgAArMdKJBYB6PFpu1V34QBXOJSqb5Ayu6
r11gfB3L6nLWcDeGQ25KL2ZnSJTjgRz7bt5heHL9L0+Oqaogr93DsIPkGAkhJsOsFhi8sF7P3f3Y
+CRTBGzqL1t4VuB8ZLWS6YtD8L3KYJurA4JqczqlQRN6K0cKOQTHmWc8li9JpYqQc7RRukPGE77a
vn5DhaRInbhi8WgTHy8WNe3PJfENdEbwZvQftwYEldXx4l1NEfBMyZYEXkBDcLkHWQ8LWjFvhU9C
DFdoYwFJKn4sSmvR/AyhIMeL6Ho5qKbLGmJ9Eve9iHW9s6PLz4dPLBv+cznFFF/yJEMC9jxtQmFL
IvJvUbJBh84TkMPS15Slu543rLEeE477d8CKRkhN2pitbHEJPFUmo9EW4H86//8123w6N+uP5jfe
g6g9xm9q5H4UjFTo5b+12W+UKcvt/wsC/6zAh73+ogmmanN9LKfb/i9YXR1S1Al+Ye7D0OXTexZg
b+YG6fRRwTMetE3XCG4LhtbDX+IJffRB6cxIq9ftR62X/lxAe4pKuZuoQkW573q4/MZddSQaIEio
wtaFP8x9oxhUh3gbTFK8PLqkTwMMXApW7CQRhZ/HFXTOQ8pSciuYrLCk576bHRN3fQP2CQfWmk8Q
f+hcRV9NSwgxL/xWNnC/+Gs+O2za1z3GgnBzlCHs2VZMRJDJmncW2mRxd4SWL3FNGYobpOMGjLz9
z39pFsuylZ2hQft35Xo+/aikHXEY7goD8ClYRm0IwK+tE3DpNvK2vFntF1iSvPY2GsQ+WMRb+J09
a9hgb8foFj8H5ysLIdmlKHORS9as/IJg6G2twV9xqiPAxO8yHkvmGdvePTV//UP8M+qFiZaVF/Gx
MeZzTSSZ7raVXHBz1quX72///ROqlls5JazNWo9O4/+oXTeYPcE++SIlypXZtmmotyLTrSKZ3vbD
EJpDYogeD7HDO/rT6r2osH92exDnzAnfmXPfMl2b3KHoA6WnA7Dlu+cYoY56c1ToMg0rWJnK8FwN
Jk1fHh1z4BPAejm5EauHiCGDE9p4R7oJ69csmtQpsqFNuIqtzZfAusHOXu2YOwy7fSpWsMNONJqU
n9rb00+nemvmFQ25OCVC6nm5OwCVo6/b28zNzLdYBGrcHDlqkpH+QSUVhCJqCjC8R2ZuNPZr4/9C
Ad+eAXaw3p9K3cJ1LAeyE0zyOzObutA7LdSTp0KStwtVe9eKphtLBRkQCPx29z78D6ho8+7k1ZWi
AR4l5SYuYAJRSjgHGopQbMWv80uUml3mBFH6G8Dtu/gK/qfmXYZQQ4C8b1NyPFMHvcBTccVetQTT
wKHHUnGQGpzRoi98ZKR9tHHxFENskZtZp/7oo0ojzYMZSE3lPX2tP0J3KnBwTxiref6iqwBYCig/
uBaIqRsmXRp3gqUUMS6NGv8XrYL849KHJBYYn8V+eCdnRz8SJ77EDNMh91H7yiVTrMNdAOXGIsN5
ssImJvQkVVHr5Ki84L36D8qncmNvBPtyQICd+sgD3eKpl5ifQ7tPGlNcCDYoHr/VGm6mJT2VMiCR
7rMG/9j5FUg2Wzbyfoox66XeYm1k5UGbrZ8A1YYFNNbBuzkqAPkUkPZZzYwzba4tykGNW6r39Tda
qkaL/p5JOjW8kBXoMotO9kLwaDCezFPfGXvnng6VV1rvKgaR8rke6a51YN7DtTchiMTsF+99pzpj
IHIby1q6+l4euzg8SQwQQY3AjGopJvlzOGWDkPiOCQD7/JMaONMDCmg3YcI+XEV+lvEvM0hJ3LnW
h9+AdTEAvbL9DSwQSZH/u61vLqqS0muvFEsbWQAYlJNzQSg4sCIGn7u0h75XSus5b8YmaaeHdr2r
1465gLk582nnQwXwjuc1MIbaIXx4m7/7LSS0H/6TWKJ20CnfgR4ZeggxkOrkJmXiyxGo3L6RdlWX
+hB7+liegDWF5i8UMkiVjvBb7yhmyCkSR0E0SXZTCAYt7y7LvgFkYncoumSMhbHgFR4EheLtUSji
helfsdKIWlAOunyHGr4ZspnNE4smUwIkYJo1EDtabbWO9CCkwTRIe+3N79T1qS4VRibDf4Xuh2gL
7QUg0LVIok9KK65i58vc+v7zl18s6KvpQyCgg14ub5WLmR8JhJzNOXZ0lJxduXWY94OolQmyRgeZ
5+C6HufZ8JyKmJgosvHY+3V7Ann55x6PK8UNY8eRUXki63yry0w43Dhc0utfw8CXt4bh0U7EYaDh
uloMOv876C+l49Lx85JphSaENg26X5KzxhYhOMaLkXAarSpruR6tZ8a83QEiWKvIkNfX3S79ialT
jx1e7TCRlJ8GYmZzzLgUcleH7r97b5s3WlyzHXiYxlx93kmb+i2P98NYJvnDtx1bx3ppPzcLlL+F
pQxgSvzmVAEWHJO6Hj5wH0KnNiX8DqnoPv6yQTjqJhj70tmr/gWioWHyS8eYeBUoT8lqdFmNbF7W
971ogVAypM/NRgD0nRR5j82yYHkqkU8fsb0VDHz0ASev50DXo0Z+84WUYKIpQvSkoWps58j9tW5v
ca2/Z63gQkVRYm0owwZ7RI3HeTFYF2EnPfpks74YFSAYbAvlCbPqVjwBbykaSRNMJYsLGrRhCYL+
6sxCGDOdzECt4rLRY9x/48eFIER53NHbFGVcrTcp323ljY7n0ydEuS00jHHAk2eQ4CywDn2JEH6O
veImyb/DgQCifYFtzUBPLUYk5MUwZk76BqJs1ecwoRN+XFfmxcNocSzS5oZhYxvTZ+wvtvBv2GPt
f4Knx/EVCuxYeu1DBAP3saFHjIfUtnAtYM/EodI9JncKalFwoplcuAJ1fJEfpXuL5wO7D0t3j4V1
w9JjLTTagwyePfWiD24zr0hAwrdgUch8PI3plU5tdjXZ8tO/MyKavGjk5oGp+vNIeAT4J9U0/uDM
esFMIrj2F4bM5QhnPxXMHYZCLX7Ms8qGAkFJtGW/rPx0u/UQeA+WdSBGr1u6ApPtugKVrfNOl5TD
QLsHyIq2QUa/Nt8r+OpEuaZOPlxsiWL/0dbbUm8+CveGO1Oc7cktw1ncbVS4infly6RtN6kTq87q
VLPW+Laip0c/+hcTI5CSPqaZBtavcCFgnJr0Pi4XPjZ0IsrVWck9Z2zUlE0M5x57QvZSBnP8K6rL
iVjP++EQwU0sOZr8uxFHDDLHqFszCs/Qw5lzPJAjy/O0o6SnCzl3dI3d9B1ggZtHiDg4r/UCs1G/
7DR2BGeBlcUqR+ZGKOBvrY7FbgbK0v9OzBCLoSXNp0L8l3Lz4/G31x1MncuYR/OX1XhrzIsFUQmd
XlpZevD7nva03HkDn2Bdvy9cBDwQuJgcb0jbqT+0Ym3cjHXRZOjQ2uhbFMFmEZhR4bCBo/5FVEEu
+NK30OggzuOixCrXAIVcjdWjfVkK+tq/OoA9iOpx+G2n44OCJ7KNyaODIZ4dO/ClGEajMH5oVF/g
0r1OTb8R+IuL1r0BxsxbcRBZWs4ikImLwXM5Danduw4sSjmzY5tgHMIvKC/MWk8l6ZyPkh5mQnQ4
0RUafJGxRw0yXtR5zmIvHYKmkpTVksfCxf5d7AWdv6JjvFTkZIz3ZP5Ly1rU0AAeh1CaIpzaoqFq
KFdY1hy/e5vBduYHvAvfLfUinE6SWlsGnbasFolYXUmrYuCzih+q68O45OzTbguTaJLhaVp/qAML
5mkhcD16MmqJ4WuVTyCq77umIgh8tG7g5V39nqFp/CwUMOfJaBLri4dbzQ5eZlb/4kPuCXuZHBdc
L+A5L157HWQuH6yPz501r+XpioDAYYrPPWuzMw5fyHx/vVxImhQctSM0eFmEoyTZehZX5epn5mKR
EOhtgJJH4k2Ql51siXrXJ647x2JFUozy+LVV8wMf71Inhj7ioTw1Ie93rV3x/ji6KJiKcH0fwH5v
YqBUIolJHOpGmZUcON0YYnvZmWNRHWS53DyHr+Ybq2JflJGVqjFDuuzMdVonjdqiecmxPMkNqJb/
2dCWxxt4V05hfiUEI1wOsA88bHVhrTgUfJ9fGgrNhTT4CJlj1PtoogBlhZxn/0ErmLOUr+DRHKWw
L29HoYsTltjkACK+NjOCk1zH5m3596KAKi260kBghUehWXmt3a6OIUVHeh+8hVDBP1rTJsD4bGMb
QJfsz8OR2DY7bCngE10XNy+Ad6Q7WukzP5kQUkFzLVsEKboRKMPDGPTTPqjNRZc03jiOgiT2KkVM
1MlAH/dPHQLWJkZkL3s63Q4OasTXHhf1BoO4CfwqDtiK6AQUKYv8lAKNgMB7OuOUbVI1mM0eEnkX
uizqfkv/LMm0z+Eof25cTp/NFhnY7fmx3pYo8i3P+14mx+efTfZy609WwORjYNFk5El6EfP+L1md
QVDlk2U8SMXm6fcGkTCvb6vGUGWNnbtkAxFcEbwWsnQjqX9hbCCzCCZMihfE+bkkE9ufWp/WIXY0
EMpiC33X3jgHJyY/030HZKaR8e+RCSNd2P0x27RBtOZESA3oTdj2mcBc+1dTxDiwCoMthTORVH3G
3A2I3ALjwhcMUQjVNI/lOWnn7YNuEacgOcsGQUuFDV0k4+6teq7zx+q4/enltGC2L9tOTUUeU5id
I3O+WvKnfB/kez6uD9+Kr5J+oMVmbrhjVAM4X4Ger1Ja7lbW4sc3ORTdQjeCXIsdF1CyQPyT0fdH
fnjxXiGK+DBmL83Q7IDD91yWpkGtkSlXMACHXdyz3cxfUAqZSExm2im/eU5EXdGx0NuopyNIMe+f
yljpfiX0hryq9rbCRWYyReF+F4Dxv1mzSWnqHWPlffPovibHSW6Yfqw3KyaRjxRQURunwflXYKGH
ElD2y0XMmoHo/iscWULe+xmGPbq4kmnAqb15bVDWs2vAnXRPJ4sMMTqD5EPxQrhTTXUG53IEPItW
mkKRZ4sTu/2O/4daB8N/NBx3xjrFyVYS2EC2RpBeg+YFPJ0aPX/P+H0p+Oup6m3dEKRJp1+lOD5z
4IZWEbb7oVex+Z1I7tflOMgIbJ+za+cyacez6QGCkf+TcdaGKy0PUcAFR+EHbm7TgPzJ9vpwSNOF
cglu+Z+gUmpfHJxfIPoppEZ+UlwfhGat1NfLW7PBtXWekzerGy++qJv5Gdffw6RvZyE4ddpS6CCZ
LnwiQpQ9/ywEhEPm6ngkOtUyOFNKmu4SYSTQcvwbs9rloVcKCM0O5jzgy8o55ZABlRCe4yojy0yo
/zqyysOzfEPsKa8vB7RpdYd4lZQw8vtmpXCm8mImpmUR6qvWcLqHK7J+BzaiiEJR9yp/yOnQBW/w
a+OYpKAuhDMINczB5CJCIt5hyYeIsQ8FQN/LtXs+eYBbgZs99YYJ6pshzgpUriFWSVSJyhyX22Qp
CIwY5CsO0nWgBx8VqZ6jR1qgmW8F6IxAQyA3NBm2JSyZ900jbDZ0q7s3c6Kicm8iIaqB4d/XmH6P
aGhuCcSiMbH2bTmF6omDxukEIQQo7cvllloH82N7beNJGS/8RUTfgmZuipQpPXd5qKoxf5hzCMEP
V3XnyDp3KyiOBEYWZZK3Fijxx9vlppUhmCo0EY1K7k49M+Fhz0yMqOJQ2m3jnjKiLblHw9SerrRp
Qw7bUP79gW4vF1AdifI8RJfG0Kl/1Fi/oWLGn76ZH3eNrNMI+RIip93pcXRW6LG9HWR4fFmpwCPT
PU3Ah4nW+uUH79ntTkyVTS0RV6syW67RtQ6mtJYDEatdaxDAJk9knNjP9S/IrWMv3TO6+ixGyLq+
WhrtHeMk3rGuR61BlKremESQY0Zm5VxJUK2+oSInXzsRWL4+UCdujY/yThVQHoq5Xn1+uQx//l/2
N5VADEsn0XXIAokdGgQtgxYtA6RgModXDUmTSjn2Uc4fDxB3CMnuSoV1gjVNDFVjzi7tWEs0/1WJ
IsIKbm67HmJJQyEpbMwk9VcA6wLuZtQnToc9E7WlpqPMAgZGD5ggrbUPZjpkqf/07PK8WDaioe/6
37Zen2QYhKaI3uhBiZodYReQ+ZPn/ne88dV1b9Lhx74feMprR4IAeunq4jH5UGWItVmKNLEFVL0v
jXhksRSuJ6MMpltmDmUqj36+vRygJ9Zxk4EIWnB5YtQKATBrgs2d0P7eHXXWJJh7Snl6qK+nzLUI
2yK122nGrhp9H7gwEDqzeFumuHVCsYUeVvjaMLyxToQjKjCQATmPbhWELf8fnyeJhxJ2sxsVO5RG
EdmBmWeLzsJiajDCfRJm5UxOhJVpLTmo+i5ZD5K8vkTvwCzEgm/zuDgdfOScCgDb3OHnPcv4vcq7
F5aiiCpwy5Y1Hx2F1+Y+KCIFX9LDpNI0a5+J03toXvl6TOJw99M8lOUAeX7LSdKNC0S3ld3Gr9LF
VRV5spCG7/EgjyigMy0HMs/12dulCVe/IcesOpc3DIYooR9URx9cI3/30Ncirb6PF81m9EhOutaX
5aucZGLG3bMphWQaD07cwZCCry8+sE9pYAVY8eL0IISo6t9tSu1tdtlxvN2iXSZ39DcSVjbS5g4Z
1E9vj75CRSekR1OtAdcqe/66XRgkGSMHieTGi1en/lNbKSh761J7/6ameB67DfZLSk1QR1Unzmby
Uws38Xqg934DhTxHMfMzUnbt2HfAEUt/btTwWjP5Xj3KWYnWrBymsC3PK5QSaoZcTDDVizQ5p5zh
tmSPotHTrwF0l43LsdwRZ/6Tyh0FxN0ufeTQp7RGArdt+7cnsV3SJtfStd3ytzZIzb23iiA0NANG
4TUjdkkxbi/aXoxCSr2lCpIJVvIqU+CxU0USMI76ZVsrmwud0lxi6hjrtr1Hr207AivR5THl00iE
QpBU3Sz2YgcYJHwtAqRGuPLl4qNRiu9SvwsFxJfXjhx736Zwmow4Jaq8GoNm1mj0TK7e+g5AFYJG
H/5Vk8Ahds+uBS2Ioo0DEsmeSBYOGVGUboPC2SHxsgKexDv7Xfz0T2RDozsMa0Pf4713/scgaZ25
sKpO31aE6JzeqZ7jFyM+aj1pidBMSX6tQ1PZO5PcVkXh6sQe6al9XgwussCMLeruR5bgVBaoC4O1
4MA86h/nZQ9YqBk3c+zOxXPQ1btl4sVYW22StHCiEYavqSYxpYDG2o0OYy+gSlLUONzGYRy04/95
7pd1p6vgqW5jFPFUVcTRSxZYK8XBKS3hPUk5IjzlC3bFbO/EQ71AZzwQHR27NetAkNIQoLMD3ogX
DLqKPCH0hPI4yII/iPsqOLrMH5AJRrWrNlxRARt6HnVhML3g/WT+dNPh6TVNKPfhDM9pVlHv0C47
AKEe7ikxaH8pyNihYyPHoJTCMcG3n0hF8/1SO9b37vxQaLDMkbYzW7bJ49L77OvofNDTAXdvjE1W
gTV0tOJ3wll8pJO8GZAOtD8duw6DNDMEZ7tI9rASLaAHW712csmUdwAWjcE6o+Fzug8TF7QOQja8
Mf4LmAuOos3nr62JlsqlLmetSsd+C2gZosGE8X1FaA/J+C4VpwsIbr+O0mPjYZmEaBFRU7qTF/mw
i+c+WXdzZFpJ+qu1SJy4vbNX7pqIGk8z1D8krwbUttIhmhWeUnk+D5aHDV10yglZGE5Yb7FSG/Fx
mA2XTJZIE9wD6lIyJbAeIyS9KPdun4UQxidio4t2p8eaCUCDaHkTg2bvyVlCxdKgq2X+Wd/PJow5
NSqxCTNwdVSR4R4k+8EA/rRo7xXkn69caEwOmP88EZ6oisn8giitsopHbyg8E9pi2wI6UjIkV1bc
+87u/B422TgX+kWq9c0jYXsjrEDMDc7ICIhlm3HeqAfzgexUhgKH3rUvrlV0MFC4TdsPScewA8C+
AjctPjAvuNgYIy8yAdxOjTtxVuUrwBiM0ieYu1BkV1VCzxESxbVQaz9lqcrx9C8pFaFFMeDoE/mj
kZJZzNiUQE8zlzGrCnVWLi1dwz8T9YHWZDcpaTWCQS3nG2kFYn5IeuY6h54m4yAg3WN1lB1bZ8Ej
NrprH+MQt7T/4welwq2WW+c29Tjzxryhn8/ntjSyntcGxitgePCD6ln6tKDwI1e9AqMV/Y+sECMn
2S5xbjILPIzXObJo2Ukfjk0DWWA5IW3OKgDU2RNCRUoi6m8anU6iP3Wh+gvDdh7+5QLlTNrOewww
+AokcDmNlu1kA4/OBxCTaCS/hRDymLc7o+OTpVpqFu3igM8YhuBgbn8I92oIm2EgToQnn4bhdK2F
1gyi+51BORVi+dzFettJhYedw+1vXiv9xzxeA4XGCKmeQ9QzOVZdv7ucHpn5COeQh0zh5nDxInKT
JGXpJamOTMmz/qo/NaNDNHo2oF0CvZ305/d3j77flF/H84o9VqLKb+9A3zkJeEyuG0H7SvBCqWKg
3viCdxrHktKP0flEiubUurki1c8p1LsTqPfbwBAXkY1PImiULWPzxJUd5ASz5E/xjtdNQyRh/US3
1qJaJEL6wZcCW8IzpNNQxAdwTZzH3MFdiIEzP8kD0GHPD2ftU9rPONq7r6qPMYKzNMFi/qFJRi49
JkIwwiIWBkfJObVcU8uc6hwvBI5vtr7L3eiPza6R1Yyyq1nrRtD6iB4R9pvERuCfWO/6PROB0iKD
yHEnmV1prEalIYvgYiGH1rIEmRn1G/TlJAbCGsvXjq1cis7O+7bCRgDDgk26yFPh4v+eNQGQQIlH
fJFewxj0wF4zMiXY3T3aXUroTXlTptnfVCbVV0v6bf2w88za9/gygqJfboHnwPI3yd1Xo9qfHyLP
Ac5v9I8KtqiKOx3hukQjDpFWAGJEcfTiVxRW6XpK+amiwHiqPG/jVCBOf2qvUpXMOrnfPdybhtvq
EVZrnpmODcspKaEo4D93bnbCoSubIboGM12PiAWsESbe65xto8na5X8pooh39TDg7V6kaFmQmLob
Uo7vpqjWizFi61PcnfFiSxihPUR5h2GDU+bJaKymBbzXXIVNN7A7U6EK4tyRWpQ6lNokbH/EK6e9
bSfkUzv0Amk0NjdiC2URtzx2gkCzpR9kz03kR2TO8xqpDD84KmDE2Po5KwaRJ8UQZ4sLlq31OOet
IjnowDswrhxgEAMwN+y5XTTKi1WnvIDjFaY3OEVgtcr0OPdlM/gnZOPBHw9/QxYZoAyG2M7A+jYs
45m7ovseTiRV95h3RPNBeeLcb/avnk8HUVb8kfe7qGI1Zkl8FGt9U0T5Jnq10lVs7NJXWTXtwrhC
Y2giNQwA0bvdxgxGdOFfAl2c/oe/wE6aANY2XHfWndZpImFs103IAVg0LkKrEvMkn/5zMZi+R+Qq
t+dEyshz/4n3QBQwwPBZ3NuAzJQb8w80iwVVxBQnHDIXGtkKH93MqTylDVWWzFldnSj/poID5j8C
7i4QCr0jB053pOBZOt4xSXaosEC5ne5ZsXwXSminkh+onVVO1NwCkwOCoBJrBIGken+YpLXp5MDF
8nzvIWoBZh6taIdgkc9Wq0ac1ZBehN8ME/HsLJTCD4fAuOxr6cMnccRGcUn/ch/YlaEn9ECxbZjx
7sNg1KK0PqMt9g6+G7So6k6i5fNVgGCbpI4bE8RI5ccOOyaOmsIvjXZZnCSicpB8FJ1ODbU6lCVG
mIsGuPKegACcQfqjaA7LRz9Qc1GxJHd4HwP+yHUXpsofLviSxBQDb592vwlvTgVTwC3AsudRh7yl
W5xYP0hAuGljQsWGQt3yz+BskKig4FBuNVZbeX9A4bZrROWZyVyUcRhRbDqA6V49cHSSYjM5IeVG
UEq8V9zGarJuCGZ7BWyQg70nWz8J2TEoSC8qFtxRLfG9/q5OFuPvmPTCETo7epr+PTL0qW18lYIu
9phhu8/5JuTrYAQj9nDi3ALlMsrRaDNMr4K1667di/1/lCrk98V1w6JodOpIixJM05zb0it7UoBE
hsGQF7ZSlX+D/wNEhnJxgzwZVJUUP05rSBf9b5NMnNlvc8vTu1AgdH4nuWmV7Ykp79n+LTaFmj4J
dLwkML4H1UKEZU11xGuHVKtwBDxad+ljFc/Tf1a8rmPD1oraNnKm5lUQmL3XcrmemURNahhWX4tU
Fb7vusQUOL+gTjcejECC7Uut0CraTPPScPcw6FUFn+/F+2UufzcppdnUOwGz9KB+1W+1rdGPdehO
j4aVFcbjkFisLcEG6OmdVsdiEgNZEOBSIoaWOZ0VUVjgtj6MtFnp4hRqx0Bstlf7UydhIBW/C6xX
HfQZcalOHnVaviEbMydAmS74wIa3XPUXoMYSkm4La5DYfVWD7Ozv8FRkqMesgiEMDbls8My1jQyl
sT6gunA67Vx/ob4exB9hZluAwZ1ohYIl3lxQJiZAU0QG8HMWJ+9QEEXICnPJOPUsJSLuUsLrI8hQ
XcvaQRfqkuYRQJOhuuHy+jGuo2b+XQE73fn4czSV9T/W81l68lW19KSF0YltcKlwbUD4yNZ99AXr
lP6HVaPCAaHMGNmjSzVgk39VA/PeP6CUcCgwy9ceui9nsVs/Xtd+Fev2cPQYQNNA2f7A1sjcs+L1
7ZeABFhLHM5nVTlo8y2bfBNEzlG873eU5uN+BYHsI5mLynd3OksnmMFM5+VOsfv+nTleVrToxYax
ySR+9Z/O5Rz7poc146IZJ+k0UVBJzCpxC0Lv8LpUMt+cGCTs2cP1P7K7MB82B4oiiy08Jq4PSZgj
T7oToYvmZ3/y64SdCekN5iOKz1z0jMjuG83eW54fcqC6cl1TRCelIVFj0efvE8eJE3iM5z7BrIew
hnr3LL3gQMsgv6aTMF/7VhmRlhI3cl3sf4A8rFnPJPsbmCwBvHiH1oIld+4O2tYP3tra4zulYGi8
mLM6NLq86mSSyin8ieU+KEfXo8lyNYi0hi2/+Jx4YesKPaj+MvSXazaPROrtyDhLbcB5uUkA8Bdh
PaPWhEh6G7G8rvlTnMhaVDLQanch2jkT7MQVHcBE1WCujMLMT/ehIFJXjWfbzRTGlsZgc2fhLEd3
vgsFIzqbybxozr8WAsY4dVQdssi8/7hhoFvEZcFnoawyNgDYWFn0MHP15gOIFFchLtXZq8+fk6MY
hntEtWk6eqha2IPAeseWePwdOmrBMSYQTLcWEmtxoTs27WUppWBGucD5OCVmX446a143ngz0YCwY
fqBToADapmpdmJd1ebQR8prhMJsfvwgguteH/aeE5N2Se49idtPJPlTVTRGwGaYUSuhvT6ap66mq
6BTwwpkP2N+leqVlgMcM1rGMMtr2ZHL7U6tT6mbU5N9dFk8tOQC81YjWzD+qEhFNjT10AIWAPvA6
Rt+YgQvBzq4tDfQJdiEUJLa0BfCQ5PbeUTBmZDgsosqbBR7m5dblBz6+fU4Jnna7uzvsvMGUUrK9
GGE+ZCA5RZQ06NNclaL9nF98Ogqko1iTPFwOsAbO0d4R9FYNvprHvlx1HsxJjru7SyVUuSrdO7lA
Iy9hdFE3aYGjKJWb/mif4V5zqTz29ccsJvfTt9TsWW/wTu1bOhEXnBEAA8BZsNIq/pNicMv7mQLg
nMT0LUMHu7JNXYsE7tEnc18BEkA4GS4FYXr7fcR36NKLV3dMbss882ySgDorw8/Izi1BMBEyu0CI
ueneGzk5l0dOyIOnLdcXCFjgpjPETckNCLp2Ma4jKbUxEnkyOakzfD6QZNpoVepnLIm692Lu3Ym1
mx8l8gQPoo5iYQD0zG/qmDSqwyCsiZRY/3Z0xdAjajK+chI1Jm+GA/DK5RBTw25DDl9upLI4qCfI
dmRBAl0ejNcuW96PAYlx4WGKzvBvCvJttAWGYTdFmTEk0KzyD8jz7v7s+vA5q9oCSvC4m5KF1fWm
Q+p/yOqjSJcwLlzMubGKU0CUljjxQf6CaKz2qqJ99YJ05kkpMQdDxGu/A29/JZHMMCWKg5QyQtPe
8sbaCQaJsGUjbqlQLaNnTwlEKSu4/dGexCtQvTdNfh/cLGs7PVzyEKc6Y+P8AiuodM8Y4t0lCByc
ooKlNn1+yK3Za0cS+Ox1193V2dLFbYJSxZO3khkwvy1dxyrN4/URkmGNKU3t04uYmJWgzvIk3lsF
E9acmndFGoTnJzPuXwbei+GdewFSj96bca0GhS4hefAATip2JpF/UptIq9DID1ttIiEwbMobj1YQ
3n0bUtMBxaOJa1nEKhZ+HOxlC3oJ3vKxf73u4/7nVfI+W57szkgMnXNYvdFXu9XDfiaRRhpvRjQm
ZSuct4GFUYD3QWtE6aw+4B6kDi8b0VjJTo6FEXdGmfjoCZeiixSXXIvWgrHF19qgwOFekuXdQeDN
kBBKIgk2PvocxnngBgBJHFk8K/RWWd/JQul4FdVwHyAlDvapOt3tpnrEnmEhxTwXDO5ZFib8MPCT
Nsww5xCJxzQaYxxfxNyAmq7lcqSI6NilE45TU0+uFFU3gM6EqbC9C6LPdEGT/M/pzzRYVrtBwyE+
2UU0j3RKEvvplrX9beR1W+UwGgFU+RLD/EHa66maqI7SRkjFBStF/hRNsLSWe8/2l/e1XIZZRad6
vKPZJeqc6Q4vnTg2vxNL1Al/JMBzGdYOZHM80FF6wvqKufaI4X4IYxzA/NFk+lB8gvOU03LU5ktZ
ZFrvM063WuV5lZMkWVvpOjQ07mmrlG8exH5femEGt0esPn2oRlj+U8tZl2Eioc0aClWZkHL2/6rn
YyXZLU61Ldl5su0uy+Jub56xJk1sKRgLqKf5n3DdD+E09OdaeCPcmZKQA3G3kxVh5iiYkNOru68v
Ml4jd6Wqz88Glq1MWKdq8GtsEvhTCrCmDXKP0g+BHtNauvm9WqlNoD53ZHYL56Iay7sd4mizsQP0
iSm6AeuRrZzkHrKl216ulHRj4SQn29BOiURFUVavbkm9FcKdbCuRVz5An9bxuygzfnoe08RpN3Qe
9gL6ZfdlwRRceh74nIpV6hz0VPUuGsQEOFtkDwd1bVygnsZKDisnSpnRAeDZtH7JQk5z0hiKYEwd
2Kww1WGwy+ykchy2hr8I2TxUJxqZHXOnUEHOugWKa9LF7EaiPHWdshLPC5KVbusFYt+gCJTVw/bJ
V0gmAlnQMa//2IvMitLx3dzeDqwg0oUz/0hbheLhhTqyrzNGV1fhsyeP4KDSdu3T+HnJKhGmpPTL
sHQqxmH28ToeKsnQ4ZAU3zYECZXkDnaAF5+IeaYDByTcNckgjVTSpd+h6vw8OpDnihi3V43ZoMfR
yw5r9o7asZsKWfeJXEJb0GTAMkI4mQtjS6iZBzRapFtJXobKVOZsjOSfdM8ll7DjIuDjteUnH6Df
zDu/yPs/U5csTiFjf93u8Jb9Ni9UyVnlBLYwCsR1oqRnkLHNck6VsuxbDdrhUG7YqQP6sKu+Eahj
e3bunak0Vh6xXxk88m3E68bE4kJtmmgq0b3uzPEsgiF0OtgqTBnWoF/AVyfhc5JInjYmJ9UHX14+
+8NAHG2m2gsNjBcnDGUpnyq+nWbrQC1o79rYXMjkfq9t892aEjrUgk8C3SJxaDuPfat/qRUb54Wq
HceGLGEu7Px976OUFiBA9Le16WF/FwMzQEP5pLdUYwb2bZIjiuox7iZndD8u89p+zZRoPzOYuZIl
/Cmb5yEMZ+Ue/w6ffQV5qbE1/dZ7fTC4PdPvZ0q0ciErm8N/Zvt0qYtFhjWNeqjYTkzI2tTRdDzb
laSNLy/zU+SQ1u98A96gYp+Yffx3cN1FIvFpf2KFiwCtg2wTY8/QXsB7igHwhkB7yb2mFqwISFI2
291XYLK3phnWFC3t8Eaqqd1NnScYvaApmYLqtxc/AKk28zXuSgRogFC/qMuh6Vewwx7eA2c0acT7
05TCQJQDiYUuhSuKLV4ioeVnu0zW5HAd+KpmzA9JpHrS1kKWs6SoqPYvki3VH6XKlsTpoync00az
Wv6C6/dzB4n79Q5rlsi72/INtaccb/WuM0miGCoTEo0iloE+nrBg18XAa69SM81Y7PTIbofXu0zA
rh//YYkg3LvySWcNk7oZcqvHsla6aQipkRxYc9/3k82PJzQUZaSlKDGUVUc6k+ioFynaogn9JrcZ
eBFs2SBq8FjGfNLsMp2pCA0L9xf3zoXFG5txfGZFg7CelZ5Wx7WHM7q7H5Ge5oALPRYqY9k3oV4r
+9t4ZrWTh7JM8llQKNnFlKqvygk4SZR+DC7es/orFkpb6/kO3m8K3u4RIZrpIvaSOIgMFMiNRRmn
6AfSxnPHt3AG6otrV7e3hhFAcuLS6q62/xy95eOCGxqlQkOrTlSIIr+hubJW+FhHCEoAsgDsCpZ+
uPEqbGd4QgfcGaBwi/jIlFrWT2u34aVvEykyA0VqswDPcx7XRFZtFIX3/pgfwcWvDvgxDCklNwSJ
4gRqh5tnulWZrFCilrFDJlqmLEp2kubbPTbcih4cqQ/Cke+618EEknJLg2WOtj0+MLXHaqLPRbsE
97xAni63wGiTbeHXWKujYoDDO01tny8xW4Y3Of1wCUtTVDt4Ok3t9JArMLKZxBpJp4XgbFAYkpJc
WQO3qxZ3A3YUEZrwxZxHq3Pz/ggG40UOvCSLq0sEZ97hnfUVxWRF4y1Ay46dP0sQL8CL3XZh95R8
kFkK7XKdzTEPr2F2Rr1cNPDnychwzYD6pWF1uWCRzUWDqep6TMq6PhmA/tQoYkGZv4Vbf6xxuZMf
WvYBi2HRvmVVrPBSOSi4Qzs6QSPjZ6z/Y1ITylnIr7aLKv4/kjVaD3NbX6oGqJpkYuXp/8Z8tLeF
gcitTELJ6O+GLhDVd3SA8d1gplXEj2z4lSYBz1IflLe/YQORgxg+wVpQvLBrPGvjpbAi19MERef4
jc7GMoSmIyQGxV/0UjawuTVaJQ+jhynm1H1e5n3YdtoFbwTcp4E1aJACtSJsZaccuGR9kDnwwqhJ
w4PZpeNKugAajUpEjGsGKpwkioVTuyh8UPWVa6qYZjklLq0Ulv+GTayIB6gYi3/XACCH/KalPi9H
oLz8pE1hyn5vJjLCaCztdhI4KHNGxVpaHJ8RS1XBX/+2cB/nsrBMCUwx1eJxcKWlDyCKWKFDcQ6n
fdyvwGhtUgdhuNnbOxMoFNlnSLzuwP9Dd6zORUNbRTkohfIjvQVOLkZ+sJ3vxTw+yiOpoYWcwbHm
dBDNv/Kf6qlDPfeWx4aY9BbJHprQz72vkPtZ21a8RrMRGgK4riNeuzDBNkqQaIlA2BFwx/n5vwxK
uvONMr1a7Fdfpg5cFWMcg4IFYS860pog1/SMVouojoFlrzmOamm8Jw/pBrcKY1z2prTAkz6dEj2x
Gr8UExdTEtVpjlS6VJq2U+3y1lLJa7/FwQ83jdSKJxKZ1SAx8yNm8h0o7gBkvrKfmY1TRDQiabSB
9WlnBZtrQSBYZstjef6xV+FbvZVThw0b5awarzqGzqRvrwvgaeI9RLMzTYu024Km4yT0sCaMSFP2
j3p8+WiEjD1yCkDnQ7SiXlPSnHLTlnLvtlN9IPoM2J/QZX+OilBcoEM3LpunJjWK7NSSsnt7Hcbg
QmLazzLjQZ2DKTqWZpi4EDcIJTfuJQ1FlpJu34i2nUJy3YLNsO+1463ogjpkRiS5AQ+ZIN8FKLh4
+4QGK8YgQRwt+HV30038/c9bySae+AthQxVIOz+yMsLAKihAXodxxfHp0kqi0c9ZLdbuvp4E7IEw
C1+r5wRi5mf8iBCSgH/IWe5rwGrDHXQEuojjUae6OvqlSF2e92dZxuUbpXwe6Fk4cIn6S44Puny9
xQqIJ4Em2isEoEhIJrFC5jLUslkxJWh7wu2S4a4r506eS2U88klZbYGM+UPjXyh9q//ZleXlDREL
adxkgsrawCl9Nvq0e8lEZbjfwujO0c9LWG/zPAQlG1TEUhJ6ybE/Klvkq7OC0oA0V5fnrdh/nhQa
Cl3JqjjQqo+CHV+LzYC19G7cv9VIn+OlB9ZDFb0da/yuA3uMvg4E3J3Tl/gpfg1WptzLBCi8Ubit
vJC8S5lAbBerIke3lF2QZAfMoUYbb0uXZUrqH6gX3D7xYomsl2jkHtOWq1Edf9HUkT2bI/xN2DBp
1kz8uZALXHaKxbHHPhkEo/bgXEooaLDKUSw5hY/guzyycXGns+O2Wo5qVL3h1s3sAPpI94qukzRN
70wfmOKRVa8b5/AZYdsv1xSY8o9sCZlQEXvwaZlOOJovI4bHlmFQbSm1QTw/X+8BiYU95AGEu4wJ
6RHhg0adHX7StrKZ9tSwXm2qLjm6urQm1Kt+5VN/jlGUM2iHN7AyTJ3PJJkblrjIUxRbJSyksqI/
b+I+sI4jEcKqWcGnY4Z/f3YkIO02nZZQazxdbtsaGLEfI1wCvUkfZ5FbSb6t9Uosd0/vpnLrQuoA
X/jz+8pH4QBV242dp0DyQrXHHptNl0Djbej53NqDubRC+Y9DntXpfL2qqaWSS+mBid1/Vh6tmQkq
JxPOQdadiAJKINCYQASa52rjG7IGItBebUI/00jMuhFE63gK/Ouop2oZ4VeY5d44SoogaN/DCLii
lf/fJIUNZD7ru+NPVcZQxqCkNbJLPccPyh38oUv0sXdtcJw5irkhEgQmATmal4MfZysRqw0Mf3nq
qt9KDqpJgmb5Nhv8yHx6/3Ax/31j4/RuUiMdx0sKk8h4ft/8oTTurbbMgy/Du3CRHBuYfzxhBlHy
DZYvwQ9wc8xacYpfkeVD/f9pQeYK09VAMM4ZCGLIjLpSPk8kW8zicOqVYplJZX+oG7cOqmGsDn9y
6qltYeaCv+DYXdOKlY0ovg8n1QdqsU2B+hpr4IE1vBcWI/b3sHVoF7Pbw8Jy5BcJV9fWrYiVjp+C
7kbGs0YY3zDkrWcQNWl7sHORra1TzDRg6rToUbXzdJSRLwIW6eHu1JQ7wRz6yRmyjtKDw/NlB/8Z
FfjN6z6h8b8x5iS6SGTwhRQzj59n5rmF89A6Cwhc7gGlreKKGIEA6yKZetcuUtfVCw0rOaVGGp2u
QiiYD+d/5qed6aSYi7btlJoIOH7HeU5zR5kv9MHgkjPWeSbgFJ3qR31ON5KXkIxOzHDb9tzWdAdw
hMvxqz2i/YE89Wcd5h2o+Y7vWahaMlgjX0Y5ySso/W6pXN3gZyyF5PE/0QJtZXCWzCF3drFvWhCN
iaWN4Rusz6Vyu1wR+wsSBb8ZsPDuP8yfpf17GMmS2PK3hDcb2qnZymF7XANGDmsrhwRA6XcVlCdl
VsQ06d30x8KKb8dyn2DJBQo8xUa645hdoueKhyU/v1PECZ/EGVVwY7aR2peO50uSy1civFZckUJM
Re1wlcEBUmYkXu2ge54M49Ts93oWG54x9BMjXU972T2li8YFyjShVcb7hUui9xtPvrcCu2nedOjW
3DaztiSAU6rgyBXHqhyUO6DLitqHj4TvL+xSwmwv1w0vUljL8/N0olr/9iGUZVde14MoB26xN0Kt
Kj5Kf31u08eVr15a2sFvsPHqOnAh7eNgPStm7hym5SJHb3p4yqipTpyXy7S1N3HnWQ9Obwnw9iJ+
NbiUgDCWxbmX6JgICXDZg+TQr323+AE38h1E2gtO+cQDPuugmveoWWT6urZCAR9fKyhV0BGRda/I
mEEaAwDOJMSkjdUL8I+xfQwkBiecYYPjvhecwHIu4Jb61NlurIIdivLWBfV3nhZWIjW4cvwZ3UUJ
gz3zuR5/69GjxRHa61gk3uklM4Y4jbOrxllAlo8O0v65wYUGITS+jLj4y/+W2ZbO3qR3m7wlcEMI
UK3WOdbMrK60X12m2LHdQ/E35lpbYcQQNB3BvPhbR4BS8T/aRFRpKy/+x4TgnHJfCgFTNbanxDVG
n4CPF79vhinvMm5caqGJ4Zu6mqFyCJbHhvdrVW+Otik5WENJxqE6ahSEDhGffgXWYLEyOgsXckWb
vs9XlEwBgbo42IKFI7O5LMQAjiror3JIw0+I88fsiBt+VZlikL06aWO4MrPf02c5iRq0uOZUKu/e
uVgHmIrO8e1Deucto5pFlbCMMsUYeC5gXCzpPuzpU0mkJ+Pz5K3nOjZ2UsY+1Mwg1ZlJCn6UaSVu
e3KbWGh0a3/VzqGLeH2tnkZZNHPtI9SZYTUgbhpDNQQSonRbg0R81GFEwUyb7mPWqofMj6YiHvqo
Md00kToErGNNm8vFNxoRpl2jvw3YC5070tsYWxMGb+BOW3qnkLCgXc0HuwnZE0eIrOCKWVPtriQy
MqjHU7bz1BorgcT5ZUTdmRNMPNSukwYcNqFp12WjesyLsr3ZZweQXR+K9jIVo4cc2JYTjSPJQaYL
7M8f1+LYT1vLk2GX7lHi06AYHWgW3Mr/SLUJKWZruX5m1hnCku++hyot08zw5cHvQHEt6ALyposd
H6mxlM+br/eqRWpHSJRezPceE2Iib3LFt9BKmhN5G9DlWsulJZ5FAM6U7o9BQmD7YG2QYgKfT8HM
KrnyHL+VQonRUMECLy5Gvi1TOFZLCyne6XyKptOt1GJo3NRwQ8Yx5pe0B7u42Ror7s7xoN/6vdkz
U1OtHuza3203K2GTojm3/ZE7z/ECRyK03TVazolGdvENWSfXmBBmrGfqUzrk4yM1vHJuBFo0C9Ou
eNkEJ3WdbFbcxMzoWwWQi23harHwNd7F8u4Cq0w0L/R6cIhOAYiKD1MB2B97KIOHRKUstSbn4MvF
gFlIVI+ViIy237Z8LffIZgg79+ynTFRoy+CYjWlrl0xY04UL/GZrzO5GfnU8WUc5QB3/GVqXbiEx
Ya9ZyCext1lTtoMhfs7Lj6scBBdalnV0/i/z0Hr9utS10B5gFoILbTIu8LkSiWNJSjCrAleOAw3G
6uHSbyI1zBBTfGt8/E2wX5AF4uZjCQab4XTzY/fPLgejN56Xsp64KixxYpaoYuHQXPQlCfmfa3Vy
007c9GHbCclgATcqkLNHeaO+uCKQpQpgb0buftCgtOGLx3SRs8T8rxrcn7TAIdYCvPD66M9+tUu1
7i/jJRYZT/vcRjUqdso6rsUh8ssjI2s1EQzcXlz+5GfWgwD4MY7tOlyVMjENT6z3CBDh/k35zvz0
EANfHDITnulsZzy/LRl8OraYXvNAyj0RVBGRjtiG6CrFm+nRJHbg3ZdIy7w8XKPYEC0uLKzZDiv0
T/EJKES1HF8Qq5LtCAw27YNSCMPShClSXCwvmPMmsAtR0T4My6mZAR4r0638ndcu3dOFkixERlUl
vz5QgL3clYAs6Dkpc7VcCLlw0emjHnFq/XMvEWAS+1wDbfKf0ozLzvu4Nh9OPnfFDObHAcN6yB9E
WHIF9lPdLA31t5J8QewlM7T0DZvAlMqEGACujrBpp8Utxygzi3jx478Zpc3moEXZgoPWV88m1aMZ
WykrgUc2QxxYNwa5Z1Q8BfX/00XJxfG+3mdo6HTNlu40K7KHapxICYFYOsYDKpHLDRCcfj7qnGwm
Qi+KncrV1/wHebiqKCN21xwYBK7Iy7WPH2ffvE3IrK45cSX54V/ab7dvGoWLfU5giU86I3PeIt18
psHV1ylIMZGEdNPrCTljQlizieTSh5UMe6f6KK1huSGNQSGkUtrmXw2zG9KeDKOVxrmQdGjSB1xm
PgMZV6TyhCar3A4krLPwGUqefXfaw7G/a1Xh3PgqDyQ98zbV+9bCkb2bD0tabl4oGaE8oAlHnBY3
9581UnukesPvq8QDjLBr07CNttM8YNPqOm9gdV75Gw6iZxohJVp6MS4/pqhi0ySliKeG2xU9FnK1
mA9f7uwf8UAji57UYm/33dRQseVnM1r0E3p+Sw6303NHhgCsVgIFoh8vjbPgMIr3shIsK6Y/RepU
ORTq9hG7AerpF5dwY9VX/LyVPnw48I1Po7+uNkVsyHsmQFaqTddCW7GIMAsAHxhPNeSebDpJyG7u
DTx1Bx8BB3j8btWMQpB2Q6sdQA6qNGMPZ3feOie7dtmXb9tixy6Ue6zBcygsJtrQJrV9zrbqu9mw
SGIakrvSxL83zSX+P64JggknRXxkt811aBHhymzpiiWFqMuyI+0oerI5ndimBtSOPu2Qv7sbqGnE
gRl23Be3FLA4lTBfzf5/IdSSCqskOrTbQN97OvAe78kIMTuow4R8n9UsZY2E3ObFFrQ13W3a+oE4
ETfC49zFvYkXi5tXdHPHczdtQt2Dgq3rjMQM/f1PfG7fvcmhOSpPwF2y1aydFBzKOQtiFRpsBFGU
TSfz4fnpTV9n8PHfnz/0HuVTEG73kveGr5Ho9WYRuEnz3Lze5AfquN/et3UFvpVkfzdFmHcz8k3u
DnbMKnbac4MLRiuPIPoqYTMpvWRgGHGQEggJmBv5nbHMR9iXb2p8xZZa4cf9XwhEdaddz4P0Ulqu
qM+a3eINbcTwhvGbhTI90smkZxQp+JTfQd1KN3L1PLtiDcjD0vjbV25eoCcJWVJukAe2U9QHIJuA
DICiUhUwEfRO6+6x6/egngYScaATUMZY3MeRjzKmPLu/P12lwyvNuygn4Q/BPidVvKWb1hABl1AJ
TpWI10TDBbWP+BdSk/gkRJDY92Hitl2tVmcdCk1fDLU/IusMtZL67bA9sp7tO32Mwdzs1Pa1I0LC
LbkpAPgNgT26gBG8+7jx0KGsG/psMNo1P4VzGCWviaPuuZsCp5/oJGaSChHraUS7yn0QwlW24W4J
wzG/w4gsYBbLl8fmH7hX0YwqETC54kUmjrPQ+D7hK+FgjMQ9DVeWxmgNOtcLGkwiKSpy3wPK8WI9
NL8b3UJVnbjeOVSpIFqyzV683mL8LxqRyLCex2XiR3tP8/WcmPIzev130LjQi12chpSb/1ZKQ0il
BijyGpRtHoD/XHpDHgBugF0MO+hSYOpY85OD/WT4CLQo48Ws2j0lk7M13nVAdBTb//pxGRHo9VnP
Kl/L/1pYkXMUtrVpOlv6CRGq7EIaHhQQLRWd0mzP+3TeamUqzICQVgcBY4frL7vsHC3+nbo1Tma5
JMao4NsYP/p/EjP6D3/A1oLYUM5LznmNOk0ZtrPlZJxRB/sKMii2qXPGXQwx90TR4xBnG2WJiet8
7Fn0A1bUZIeY7MZE00ycHvY8dOgtIAnX15kW1Ab8zgUNkzHDKPsqapDZj4g6XiWMti0z2+EVcJa0
SJJDGbQrrlEiX10riz3QixZhyDieDGXzl1T9xgph6Yx2ApVh9s1thyWY4ySMhXD2qMAfPsyrGC9g
EQefo2PRFaJnB5fbXfv1Phtq3X/mSTL2zTnrenFcmFh8jgoHlELmlwzX3hlHDvFSMNOV+/xZb3C/
RUpFgaUFMvfLxDzcRlQ/bTqhgNoYB+nCPmq9epkQS41jYrkHcTnMreujqee8EDxXqFTmqnnbth82
hpymIPE/kFYrND05Tj4RFPdnqvixL7PV0FWgyiWz5AdRDgSPv5BZTt3LvaEC/mN2GYkmw9nhJVTz
U5Zt6Lz6YEsLAymUYCFgGOHhGM2orUjzRksffmsVJrgA8NDfeXd/P1vcY0lQPPj/HiL1Wy2ixI/4
+17xTjDq93YXoHCiGT3SVilJWtBlAOZHLkYRrYF3EpeoG+AaSC504LDWGgW5Yqk4POEi49YbeIGz
kvnPzkuKRj1c2+0WaOpjXl0CFEv19sXX9OShWMDY6cxo2IR6csc2CnGBDR1FWDsNzdEY9fgFkw/k
VOV6X75G2hTfV9fym2aTRg6TQX5ipIcv+rtpXaByP1f3wyuWThNrOJXH9gH3/1aLzK4d1p3RwoB6
r1Lziya61mC8go1infjoR6GUiJXL3g+g0zjVGpQawGGraSA/AbkvT0Yb0Kh4eKA/m95wIQIn8fSj
1LfN4j2Xg8qKwEV2aufCmmuEC749fK4wZ19Yea05EUPKf7KtX8pb3fOPAnFPBHiPtFsgX/jaBzDK
TpEhupikR36mcB3EKqbE3/Ne2jXYD2wBYbf82XNOJ1NJSUeVyceGEkW8fBNEpcikGB2h2IrcmiiM
y9zsZcrvHATUGcmrnbWEaLVwXcrc4jQohuBUQL29u5YR2WIsF2BdtBmRKYBtu2W7LoCfQ/hAcg49
cTcpP3gPCYrmmFMCSwfQXuh5tM6pqF09b9pR0MY3+k+Ezd6ZVazY1CWeGP9Q1tBQME6vS/RnFbbe
DLiU0n5VTe1Ph1BH589fKWWzlYl7mcBvlcHEZ5COXzJTpwEP7OxfWigjRVi6sEL4jarkdBs/PwOk
yO2q4e73NUigUXd47dM7hABnGthF/To7KEyDRXELzDHY86GLBniZ7EkcR31DzTz2GEMA1s+uZJK8
Da0XI5TGlU+ZcybG+EEBwGSUSFuGUJfVK+Jvdk0fweqpNqtNsFhu/mI4lCi40hXYVVseNJk7rxMY
zODlFEjv42fODr9DfAjfnX+WM/+uD9t3XIaP7hE24Hbu14vN+cHplXFbkpBX2ExFO1wfEd6QGlHW
CX86VbwNOgkwITiJOmd1JHrvn/yjXOVNktFPUM/h9VFQkp1SgawJ7eCvew552TDysInqi93BjG6N
lKOWHCqjJBhhON2/RfsWlMH9TPnmNyADnIAY7/gQbjdqN0/vhHisgAwhkGD8cK+gUGUPRzmHBpq/
y8bbDy20SWv9sa3viNDmsP1KoM5wE3/lYHvhJOEMleQwJJXamgMLklINFCirQ9tN3XQMn15d713b
Mo2dyEk2x7aNq7yyNcl70u25LhtxUa9YKSYaexfE3A57fVlEISP/U/mKDoaEYSs2j/CV/uo5VvRF
gXl3HltGUiBTf6l8xyQXc7jpECeWbrDnxoCwPP9qmiQVBAHnmZFi7mIoDdxbW7W9RRfhg6G2M8Mq
SN6VhldTLSx96uRQoSXaZOF0RX6Scga+mmQnex1fw5Su1H9F5Hr26G1Znsei3maQQFmcKqUsY6+9
Rtsls2gZXlKGeXzHPiv04cJD2+xuRyifSMcH/Emgv3rGngVE3mvmm8WxpyLLyVPbXdH5CTWLBByM
CYnVpGR5ndc59rqyv6iJTQvEoKwiS+cQHt2fEi0n/gwvMd8uoqn7mfu/GCjt4zO2eYBjWPSAGNZS
9/AEXTnXQ699fQpVslE0TdW+gqIaZeHBYomGuXiDimKIww4Y5ZR6sZ5Xg8FQQjVmq9T1isBroNtm
WOVXRwBd8x9E1xRG3eJ0DLe0o/rHspjTeML9H79My1b1QJmSQy8IMpAWJ+CLbamB0av7r8iEsN84
vRv9ByPi7jPJLb+yWwbQv0otMGlHPzeUEvVUewQNYHsSwOpiO54eQ9yFLjV92pVNKeNP1A4ThkTo
Rrp41ikNXG5R7KfjvSBSRBvfioJ1aPdLaZSyo0bza+kXmcrnt/B0sfnoJz7dRVd2jKh82cT6bwfz
90vKwJmObfO580UjVKcxS7edQl2QGE3xK0mgVHZycGu5KMMxlet657CuZrCM/32sFL/l70EIFIvL
ODx84aDnqbiteuXORcY+HafvFf+hI6q8j0TiIgGY3wr0s3QDEoD5mN53pOT6lOvAm/d15xbWhhF+
hPLJj2ktYjCGOa+nJ4dsMrPd2ZOyZucWqHUh77Kv2Fxa8cWiFzoTvV7Urs6BOzzyjbLzg/t0E6Tb
9PHhB7NV9u/dtKve1i6GIJ1iAMLl/KOC7cEL6942hBxlVq1RtII8sMk0pQ2ak+lONMVsi7Nz/vvD
GtDCiCvRZA6rBU9TaE03Devbr0rMqr7Hp+vzQ2xrEsrLORk88EnYvxYGHrvWPG/pT+V+NEeS3uya
pKXfO24q+JEPoTySYigFBoGdcfKdG4siBzFIMbWDkPs8tt1MH/CvBrM1fPVMWspl+LcqoCnS7ORg
SxMePAJEyu/bzw0NKgV54q91erbbOrA0jypA8GWdyvWGawKE7LcuSoSmaPRXTKKDEpxIWTV8aLQO
EwnNHcFckonCOG32YmQegfzsSozy4YIudybdPohBRhyHK+GEhFYum4Z6cSZNK4x5ZFFn6Fi8df6r
5CZ1hO/80ycG/HLE5B3+sBfXRbgjH4iBnPIbd3cibG8nM62ku9nRzwxkzVen/1eaMZen3x0RHFh7
a0sYriXGJyUWWrdnkmYcIMuI63BvOz9Ug6ZV61opCymZttzFqoilt8RsCOgXNZWXKQ5Et0u07P3J
kNbZxKFpiZLfCBU6Dss5R5tGoRs6EFGfbXRKGRqA/yIrfMvrenEfNUlkFFWg5YFIHRCnskqVqeyI
R88O6bPAuK02gUdSNwmNBYsH/oSEtj8a92B3wz/C2fR1q+C88gbbHY+7pXist2TM9WVe4JwS5ur4
lPXgeIlyUqAY2u9Jv5DMBKeK4h92vOsoooXMGYkt7BNa5+5J5o7a7VP0RRK4nCbnYzokA+Q7HSVz
vIipTfnol3nvr1sscffQWd0NfSCV06ZHzXoWgXRmEA3QlKUZWKrC3txNEX6sWoM2BlHo66aKLYa1
0JH+6ryJPmyUaCkaCrfPKXq+V68gDsDUXet17CmfBYWJgTVsgosvRuhsw3kerNcQ8FP0jPHmzhRa
QifyT/aGA0t0Ur6m1wTSuARNyvSrghRtvftkfckuqu/gmVrdPVPACQZ4HjFoy/Qc9VLXiJIPZimy
IIHZdRAJIr/nR/HP1eBlzhEAmjoyAbd6CZRrn8hcpICu4Bw5b2Fa5rGImgpLZToR2hZ0CBxSJIEc
hHGutDWdAR4gfosoDERzG7nVCdkeUOjRjZ9QOtWuV1FeCF3kGKTLeFOskNSLaFfC3e/CNVam7DEp
AdLTmy/UBkrtdCXg2J9Qaq2DM6SEKNqFaJF8CncPAwQAVDCKJaD89IdhWM0WXS5uLnebh1125U+j
mMz/yZZrj2k/MsBHlAVFobTsMaCrBmP/3ktCFRKWMMdYuGP4EqFe+yFu7Bb6qbh+HUQgmkFDN1ie
pV3j8nvCWObbFl6dfa8Ae0S+DashW5my597VKFrwC1lKm6YUlAeCZ2aHLI8HZd1G6ZYyzZMlb+Uu
+uCoTi9sR5ymcHSdLM9/QQF4RnYYDQz02PxRSDBmbUSBfIGplEHG+6Q+m84VhoqS+4CuyyAAiByq
+Q8f1frg648qsCcGgKoftzVX9EuDXx4XaBJtC7+cDym69Sq7CXtHI+3MYX3hNYvkmeIFo79LVLzU
mO9NxcJEFSnA0c1C5IfErkEV42UglRI73xPi/OTbC3Wu1Ol6G+PdTydsVrf4X4dzHRHjx1ijOdoE
clI/4MSEQDjmW7EQYz3UFRI3gH0MzSlTdBRAV9chJfAEuknS1QjrgdJaRGPYVzhs5Xl4MgcTWMrP
8unYA4DzdX3WiN7dZtl8+HNdJK32Z4OmN0YS6bX6JLy5n65q7tj0JmiztpfXxfGi0At2a18UB39C
RESE9jZhJEPu2kTtA/wbfqDMe7FvXx9rzCJQU4eJ4QyDBcPpwkA7ZQ8sNdJdHdzUlLLGOz1upGJM
gwqHv0ZsmBTgWS6KgdKTHKOHWbxz6uylx0Hl3tRryGBeHbXodDacY/dn5931SBnMdggOWJuENvEq
cW6CweD73sX44Zr+tb+tDnNRRy7xCyxva1a8unUIJybBbkwYxR9WPe2KWFrvhhib2aXM1IAp9+hc
dL7Rea0O8MUV0V0wlW8qKQG6+KvS5ZUXZXtYmq2ym3F8zz4+lGYA0LD2dlCjuPuDyIx44sC7Z8fy
TMTeBjWAEowQX7wWL0MZMOIsp96mtvUW1G26T1QS3ByFDIalRf/MJs+x+UZwUxRgmvriEc8T3HPC
Fqlw0KApKFPAsCjkKS1gzvSEedZP3TCHnRE3UrM3FT6prvfKhfAaHXAW/oG3WdelKGha115nIPfa
j0U+eSQkQJmAjdGd7TD73pJCd34X8BLWl2Cb5Odasagyq+CToturaM8D6gjvw0eKcBJM4Pu8rh1f
/0KIyXEjnfGBSyT1pWMG51ozPpQ2DgeKn+fApOcDigJNdvAPsG+zoQwzVEZmGCaDHiqJ01nl33Ys
UM/Y5j9OL/8vwvfPyd+8wvlytHqaCzbC9XgqfRvFpbO/d+/mHtgnn2TUdxFrvawv9+N2Uw9dbjqR
tzQ1A7tqTLxT6uqWle3kI2xjRCEJnK7OtPuazQWwmZf7OMHZnqXB4H2seX1RV7svMAg+nNH5gW21
mX+TVQmxd/iCmxSb2ydCV05V0Um/J4sBo7txsdz9kygs7BLZr15y5L4tqtlQSjFO3Z3qsSZ5Vj77
L2GX5Dzzy/xaq0JiM4PLzBFu/ObFN7Rc+9+xFFZAVnD+Ty/friMfjlRvViQSe6ogsqhqzNe6h8XM
/BrWxmb6ZLm/FuMt9wMVTy/OEdN7TkpA6rCpJlhUynYBUbclhI4yhJz3lzhTW4A0eWNbXMVWr3lI
Yje/jw1DL+5S7zacLU76wFaJqMZsQmzhigXWiSlQgCrmgr5ztGppwxTDtidmpJ5PXeycZm3guwiG
Lnotao+nH/2vF+ECpZRQje8b7STCr90kOL+k2ZgB4yjBrRTiLL/wXHnA23AEjreF1rYhnbE7km6k
cG7T1w/JXNOXNC5R1fzdeOPeHS3eY1Fd/aqVGcwj+w2BVIdXmuNgXgAynJ4qRcNE54S6j4X6Te0u
yKBgcTZlB6Tc2RQTv29CILQEjwqQUCbIzWZWGxiFFRGcNEsWeBeBcrrOTvvZIZzTS2Snn5AKdgbn
ZM6JbBMP89lfvXtEEqg8svtc4L+zO/oRPV5O9nBD9bQJy+7bEOGV9HDtlvKiobBANr8Bk+/7B8Va
JQtO7/Ys/HSzkStcmFozRvTvg0kH+PkBhyPH/UiSjIi+rHKetH63cbvz2lTR8de0b8D6fGz2Hslc
1St0OkT59ONKVPg/aT01pZYa3cjedDAENqPNv6HhN7KSQFg+LZVQahC1TzOcHHone30Mu+arhujB
O1sjNReI9HcCkY5quruPAHEH9H2vdAaCgANbFsyJ+hVqOCYTL7r3FLl6kquvegd007gbfwc4107Q
Q1UKM2N/SBwR/vDuL9JaH3Cwmge9OBelmndQIVBU4MRouW7eaTvrFrCzbPTyz0mtwOrfsa0pblh9
zeTFSodGhymMUkiZpid4hN6S7xj5IUtjzOriU0BuscwJQh8qifuaxzsCpFJOE4H4ASYMyH+0xAes
DC0vxZ+gb7lbx4EEW3pnJwm4WmchAJfYzd5A9TLn31JATspclkSPY3WhKav6BmrkJyfJaHLKpmp0
6jTgvKVAHvRcl+xHT07bDCya0jvaj2MRfN8F7KMgRriuYcGCBepfALZfbpS8ZgVowQFXwTcuEBpv
pSfHzIWzFDGPlEzUsGAwYkwn0ef9g5XVJkVmemgA5WEduLADjpzAPpLq+hQRahlv6Rhlfo3K5r2s
OrGBV3XoJq3N5ZtagJjKrZhhXrJJqV89zU+C6sOWTef7/v2FyQkqXFSuG6ac3NCGKcmdslV3E9/5
scwWuWINZqS07m08Ar2nS4cOpS2Wc0RySyOQZ9TpNoNsBMqlFzDAExBndAd/MdLrMResi24nHkVm
CUa7M9F6wGDVegDL06jZoYh13tdJPCjszenXDD9wdP3AmLr6obR2arp8NKwoV/bD4oJd3nXj2aWV
AUjI/QOVoqkZKOe0tPR5gqgRS0XRbTd7z9qNK4IbT0H23KMcXWRqknpK9/8L1AzG8ZknYpMI0d4M
qHqTDGR8srwGcEPFGJOrTL7GM+gmnJrQaivinJGE2rgWMyA55dcKk+vUfxs9Fu+tlaESkv7Er+0I
Vts9shY2TsBbXKHXLhkwWeuYap8FZSz0dsZzBaM5AxoEokbx69SIKiEqM9Z4gqhrNvh0B2GtOgGi
axpl3XBaHpl6xayiS1c/kc3sG1m/f5aOKedQuiieNmg4Xx49XH7cXEzxnjmTl1cq3MJZi6Sr0fmS
mi78LPMpBxX58Gx0lp0nJpsSsrYBpdgL6oSBEri2b4eKIefxxMXA+b/jVaK+lRGQJKLrdIcDHzMd
5dcG9FpUdFcvPRkWaBCDjIKTD4NrBKlVGRdEEylQC2Mhf2CqLRallUSt7AW7ElLh3iDrd/TMZ5Ft
u1cFcffRI2jB0WojHd8zwEtna9AHSgUnijllXkhNnB+JV4ZUVF56lLmVJz7mI1FTQbFvG2RVVa+7
oRR671pPFlfAjlzUkYNJHnI0ClKTNaBzJFObLuqz5PgPEDU8Hl6OcWIcs9yrc/IxZBCORrLK2h4Q
H8rbZZwYO2pB8yT5ckQIIq5drFHOrK7N/Kamvkg1x1TfoL9FT3u3KU163mmoXPaeVGmrpXOcIplY
JvdutZnjkpeR483a0te6tWnZqABzJ6xgJmQwhl/PYgTlDX+YXDyZ5EByqDYBWdQMlk0OlBzc0x2v
1tVI1ZDXTZktrQX/3flb4vtTSt5fAD5uV32TVdSJKn7Nt9X8QFQOhdpyS4y75BYp1fEOPadml4CA
GnHHUjXzfh2Mv4j7DgYF1DjHn5N5vrA/45tN5uaRuDpmBW/M6spGnC/mvZpTcDFTa7hG6ASsILQw
gjWTdsI2g3d40faFnUyFqFRkuk/GutcfgvJ7KVV+x+Wfk+9etxCMQR9pfiYvam/asY+DGmeY8S8a
EioH239bMt3Y05Vy0/cO1Fu6K7VjyzuMMRdNr6sME7j2/6AhbuwW0QVC4FFbkKmEabUnl74+y2+Z
RFZMUHNdZyTjW+90R1Dar/hEP0YeX9x0P3bDiyrkO3AX07ziDJ28MvxelMXV0vpjaLKf+DSdVrW8
K5NaqzHEPMAtegX4189GdnmU3ks11Ic9sZZJs1Ridon0Tg5b5vQhSsX/z4S1qQ6fPn0s5T+Z+pVb
mCTMvTd6VDmBPPPkexlo04W22A0HCNdOkQLPTKluh8sJjwV3tkjV0l887v+ejIrZ23QMEYlwAVhN
/6bHuKtD17BZLeX9X2r53uiZPdauuwwxgF9UB9iu0ZUlvbpSFVNeBpospkQcs7OydKJdVUWs1DPd
X5hbocbie3Uosb8FjWmQqPwsrka98xYBveCKYHHCS9Rpma3oXcYnyNpQ7cuNtlagiq9OHd9xeUHB
fyNhrYMG4sRMVPiSWwDCm71H9zm7ynVZVSf6zFjXQkLbC3XWKqRQXep7AkAskUm6Ll0p3KKk5POr
0wEx0cGoYUWuXCcJTxVOcDXL15F7b2HDjtkRecFql0yDR6/FMeHnKhQbt8k/gW8YMvP60OdD/eMz
IdW3TdXORp4n1yoBXKJ4+VfX8hGAootYBnorzMHQ7GnHWsqNTyMByHye0bqjonpMJ7nBs2zSdxz/
TkBlts4KVYM4vLx204hT/ehZ5T8034niRrFVDzL39f77du63QjJqxrbKqXo7NwWO24ANfWZyZjhs
8+b5PV6opfrv9ej4I2YqRRGrTHaqp2kkVH5VwA9FXQpPixzqh860YIPh/AkSxN3CAJgmi8HlDUDg
YX89d91zuzrHPVc/XISCj+xxiQRpdWTbYNXgVmR+01abFprnJKERVTBNF8cMweYWK6M1mWhSm5/0
8uBrNUxb2Wdmtz4YHDq50RtdhJEC3DRw+b0M28rO9NrPP8X6PKMKai17OPZAr8hVV+YvV5yLaBtJ
VDqiQK27xoSL+Wl0XWFa2ybXRb3detr4QUNGez/sO7j/uqAo9rS/8rsKiv2vxW6nIW4f3ZpI4R5b
X67COeK9u/2PdqVuCjDjjmG9Iipu7JolRCRDDokBgCczAanVMspp3n+u9LKELgm4LjjkMoFy4Yf3
oj34S1nqVaQyodr2xG/9tNQqv1GNHeypm9P7kUAPHI3plDb9Hj+kFzbZ5CcmKMd/1PTrJ7f0Ozs+
WLDjJpj0b/OmYw75m/OlYOrSu92+qleqHzNAs1tHhZ+tvyEY3ZNxoMTjwHxrBlc2mXlv7uY6lvHx
Q6R5QDOU9+W1cJG3mPxbbBtzRfu4D21krgYysYZy6jZ9igEP7OF7WbUFJXviL02b/Nk8dtMKOixe
I4bEcpL7BfFzHY2cdUvdeEnPhZjPvatR7lABpi+QzCrzU2h/uWb/Mr/524pLaon8RIHhzAWq0Hvl
/h+7rK0ox88cRz1KsPC4v5+LKkutbvMOrRki8ZhBAuuUxSK/XeN6n6AlHIOPfDBZXBHlvM3TiLlL
OSSmpeBompMHy8LfJlepRqSLQAvm8SwMjSB/TwbxnEeZUitPGuSdNZZQfqUo/E8JOWgutxSi0ubC
na0eNVd79hGMeKqdT3v0w083yaquVbfv1GhZP2qebPePYvKh0ST+as5baxIn8qsPsH3MI2BUEhDt
Sadu81cSGD/JK4kHQh06XZ7mjPh+oUupnP657N6WuwCuzBTohhWJEuD18+rp6G7aVdCKZzr1ArnA
gQY5ih1v/HwAUvHhjXiTv9n0g8vwRtCSGfkZtcT07cuEs2SHC7Zt6TauHeK+Y0Ca/lI4pNfF6Rq8
Z7Rduwv8gltUcQRmi0oIFSDIj+5sN4aNIUy01w/zHab7TCCqOGFOFVd7cRP63VDAz729E9P4CKpX
B7p6ucHk8/e4+P/ks24laWw+BL+Vtwyxdko69xBfdw2O292QQMkAon6VMm8bL7hs0S6KgX4KG5RX
0Rsx42ZR/O2WsdPWp/DTFE3lS5DQ4DGaLvnSVJbwDPGO7tc5MHzdu9JkXloxCKqZBs/HXLH6aUOk
HTg4DJr2y0zlmghJvWeVZ1h+U/aglBSgDp+oZ3ZgQmmX6jYbAGbUJgsKTqxzDcc24193hlenGOJz
v+6aOj3exWCrTuNPzdF8KBlqcVopGyXLtBJrp0eGArSm5JWWcj/GSHidmfTeGx5enXR7ra0BlD63
L0GW7W0ncp5wuyz041SztaRBhFYIOx6XwcN9tTKgC0ij+mPWoJEQkZ58ydNg2nkMtLjPp4TnRze8
jJuKoujr8GPPIghZCb7DNv75txi8SsqrDTemZJUg3T2fhnBVc3+25XRkHkPS+9q1qts/MKZRodhx
0JX4j6yKPndmE1hUF9NXY+IDHOJxAqAHI3jVNF2al+5ezUPITeZZnznSGx+7ryaqklb2QQsc/Vvz
QtVQQDLwwXJo7tnE+Oa7fw2mu+VkPIbxKTEAHo5EuC6j7TkjQo4copxZYZa0PELapgCF/XKSXEH1
NNNw8EdlEOEGvw+K8qzO4btJ0SrVxDgUDUg4UD69s1YYFDGdHk4mRvSm7xAsXVZ9fRxTpGIuObTq
r7GUzWInp8gmjQzMZ+71ggSjVR/6WvncBkTvkUtBZIa1lSodkWRtpwAOJdsij56hs45OL8Go0bE+
Fhhz0LCNXqTC/PN/pz6jsKxFLufKHA1OKG4k8VqpdtGH8DGGmsx4eDv2Y6e4s0kCQ+5Nfwm6ytTn
wkcchH5BVUQYlqShh2wY9d/LWPYbX/vfEJWvmPPERfChryPSNqtiBQMh6dhVQozVCHV77koQdJC5
9ZF/90VFcSbZFlO5J0afHhSnQmbiZOBxfwS0E1aM3wjWNI2O07oQBfSaY0QMguoHTDmbByrT7m4T
kLfG4IUDbz9n6iwWUqkmUMP10b4Jqr5wtADs8EIk7HnwfbqmuU3hf92/JyEJCnpwgeCxPiQCF055
kOKIZhkkps4PjXo8DKJ/Qn9PDeD0L8poppj/eTnoUY+Rwy/xVlPMCEFxfRiqTDwundNmHGaLNu2P
x5mpdgSbyjNxBoNpifke3/wDf0NNjCIptj5ETdGWYJNNMReMdEgX4oMbg2LzLgEQGJ3/JGoZbKA9
vXdQANjUY/wV0RkVF4JujEgOlNQbl7E8WKsvxQ3JieTzWYVD8JmTCmeE/a2mpjHIGM8HnyMeLJhX
v0zpfrUxN/E7bd2pZ/3uBETcHoZ0oyFOpnP//oyxFlHuPgvBxE/sY3ZPSTBEvKl9hOaV7n7wG1fo
2FF9Ih/hJQ2VcP5ZG7s35N5jHeA9spIYDDFlMaFl6pCGgITGm9y09QbrLkeEYP20pEPCLRLS2WOc
VOA5M/NJMNGwuiNF5HFJ+bBqf6FUy4TUi9w+jPNDo6/NrW7X4Ib3uyukgyIuCXJknGDanzvz9IL/
zCJKDA8hHxkLvyocZiYp7TJ/mehmvNBGngPIIq4DeQoZE2GiSaMg04R9GcF0NuktRoHiZReFq7le
DVDKfDtrFztgN0RTI+gAf0p6xoBy/SToAGFRraMwXdNb2lZypIusla7tJvlFaHGUyojfdjiVbXRF
sfdOiV/V7mPAwxEWQZmXogRc7/bvCRBc7oiPSQRnwYCMNxd2T0xoovNMLk2TChWdGtAHWDPcjOJi
nn4QgKkOWVy2Tyht/oGSyp77ffgE7zb7lLkL+24JlXz/fS1GveXhhBy33iyoYT+/CQUHVspofag9
300Tx3F1HjfkKmtWzjsfiJVgkXJjQNJa9ejuPrvlgy8ekskbDiBIP8rjlJvMf0RmMAT9fZZ15lnn
e6mQiQdR/dqmLPOEOSGKRhllJKaRmn+lLrzymssJ9BtECjMvgUkvntm2IlVLSD5Ix4ebnCb3Toc6
4SJrMTXl9Zl2xSrFa/U5I4kUQTWbzbqFYJzkgd1EDUTbVgzhLqpM97wwM7N1T2LA0/b3oEFrNXw2
7RqmALppRHUB+SSjSPiHjAfhiOPZHkxvW80PxsVHVwHDiVdXRGBs47rMuuf/8KgzfsNJp2KjpWNK
TxlacZWthu0+NJqcNjrTo3ofN64j+ecclOc4I18tZ2vBTKN+72tDqIaQ9rXIK41yQB0+FDuBu9/I
JfBu9Bp7tIxuV9INgupYydO2Cn8vxrSp9lQAlgZ4rQNDTd7QDgjeFn0aVSiuhPoN6dxdWesUL+Cx
eiQMV+qM6Y9xUto2Px/uWk0jv8ObsCRNOnkDOvn8jKt+KFDlr+++UH0whbBHbhoEYnhhf/VNj6S+
r1SDHAkROsgoO4HcHpRpUOieuQskVLyc0xhmYvhvM/eQw1Fq7SQ+9+noxFpGlSGcRJO+FQJl2cw2
g1NenSJejFmndLKAu0Uz0i1sPCuF7M2c0xR5ymGAVdTSRgTq7e9vu+u2GW41Ws1teoCsTX7pSFvX
utBtYwmKMD2KK5iH/CRaudgGhEtJo7mu2/ll3LjBSobDJGBGrfbGEyzqEJINQduj7ZcyxCUWqCKf
9QNJJHrhGuXaJsPG/4dAgg0pLzn2hSe9omAY5QRhZRdGUJF54n7ot9vr0mntdz7y83kkqgI4QrS5
WmoLYA+sg3RnWnpuBg6tlsuWHVkFlFHmAMLS6r6BexO2gP+u2x3jIx3XzfjvCspEH5/9RwcA+B0g
9XBW9G+xRhCHl9i4xWcqFP/WTJMaN9ItD7VwwqNkqC9ibdIVU4dnBeykldxvp7tyqgN2DRa2Tofd
iOIYX6WjxKBgN/AqKT9VDftINdqS5MVZO4hUiWN3MrSE+FnWv1sL6cAuD/LfoSNkayDS2Sz0iG7m
65AVJML6STJZ1WQHMhHmjgf3+3f4zyaMikIoG2drb7sZSTNfLHT3ucTuLOLxeXD4BCycB4Mrn2T7
QCCfRPohX8DpMVDOhfX7QuAyoG4jHEO5ZRHfTFWugIw/k0tIqUuNWSDujI4lmnNuoD5BqEujh5Cd
fWs9/5dHZ7q3JTvGc1kR+wfhodkexbUcpXGcr7SYP4spLNlXPLFvJXWWCNZVVsROvaPt9Ar0xazE
i+kjbKHC1PxhEBjEZdfV1QLk98ZwkyRgfhUeUMgMUKMn1vKa9tdk/FeFxD9zpVwIZ2U9qNAqxbHz
2Fb434Kug2X4kkaS85MSRwgKBDI0hf+mdRU231Hu6srdk6PHU2mwE4OwIOBuQsoUUgiiPs2Tua7O
XrN+GiiHrFYTD+Msgkbyc/ajFrmAZzE0mO3gnXKKdRDHh92ldj2kk1h5LfBDgzcyJ+dpRwTW3kss
dtcTqgcEu5o/H4VfdkZrDklKGFfo1HaLx2fJZNPyWo/7B6W4d6loCPdpLDpAv4+LlVb5FawFe6ew
xV9YifGx0eTNFTsf7JbJCPHtG1kjeVIbsLy5EHv0QoSWfZLOmeVMe9Wnxr3Pt1Qjho1n9MgJQGb3
/lh5lP+VbUEBdTtUr9LaYJaRO0Cmpzss+uCIbAhe5BjgVM9zJm1kHq5QjFT369Qgn9LIBg+AABpI
KY7KOwm3Aeyqgh0auBZjWcANe0FF94rGfwGoVqwwCaP8Q4yGZssSUuGIwfcXsmQc0m8YQCLTL1J6
dvpp4JBpO4OrU+ol5xy+J6P23sovUaq4ajsgwcKOwaOS8ab+QSHRiO8bjvV/tt5Z8fi3gI0+aMtN
nFjyPVUy+uZYsqijppdti5ZlkevVjzy3hZWm0qEIHTc5IQ9FPrrT+890bd6ugDM2fSQRL4jFYm+V
kskEjv5CoOFbJdILRlYow8G5u1LPOLIRVDii976IDqVtCDVBo8oF04R0fQFL/ZoO+PB9fg4yBTDW
ltlvnm3gjXpZi59NbTQDA7A8qVhr8ra4NCkaEzVHvyORhAUH7E7lYYviIoqv+clILH2gRJoZh3Ok
ZuQ/DWV1/oRjH0TDAzxhn3Z4v41Ix/v5szNaISdbzL1x3sf1zpUTchckjhBkJrSs8LblGypQguow
tXQ4WZJLwLkz3HOMB/qrS4cZ8HpRJrsTeBzmvlLIIY1gjOh+meilM6jmzqzvxh6gs+8ArXfCEBg7
WxBdwcJeWrqVhgh1IOxvOUL5PHCIlvMddWk4l+qkzZ+tbuhl4KWvCJoYPGUqiwyFwg8reVKBDIum
kMu7T6s3H1OB9D/tiLdxj1rEW7MPvHhd61cqcTjptkvB2cvkzVmHdIMZkv3HozHfHn2qUkW8QTZ0
dnFgstH67It7M0TYtZP6e7GVN/C7BDBZqlR9oR3+lqdRJxW1GhTudmu4Xek2XldR9LmAUnPnSnQ/
rbCaBUt3rGZrVBp/ioekknAe/SkgNzERr6rd/WuNnwEaryfWredmv5EDZ8wiSa5ek4CsATTaC1et
rTV3uWezZFSAEQDO7yRutm7na2eog4tKrQ9l6fSmSv8YNSHSDf7cN56p8vxp17z92MIHpbSC9FQm
L4YU8A4+GLZ4LW9m3nSbN+u5OMnv+VEFeUyf+5xH1rOnX+2nWehdkXmPrfmiMIVHkg+6n64bm+eM
RMxUVyOdZH+6ACIrZfqGRr3N408j88XPciP4L4BIHdSZQ965HzJKHIEgv2PZKxEHcHUWngty4BtX
FpmrW2Git6BcL6zLNnp9v0ojSvA6GcR0ojo+sVtfG+sfO7FGUs1hoXU8/apoZ/uYKT+j2hOyWzYQ
+kTAT2YjbpMYzCRe5cFT1IdfNVM6DLL6ixB3Ew/fuuQAZFlLwQqGIGgK/hwMsd0rl1VLS0BHDN9i
zv6x7550NfoAFE3SKto7TLq6pBh9ozlMjqHG4rKN++oIDGMR6rjbj6OFFPAkcRDGuw8/h0H+s3EI
uuuprX/u8BlUZSoRwNn+fi6LJERV6rAkydC9krDAScGiIIuJ8E9RrVXJyPb62coZXmJxjMdWyQpX
1tATOKV5jg/yCkxAF/G4N0E3bykxkfoijE5f7nBIQJjvmFKobwsZrRq05CXXs32DayRs/zyPBtcx
G12xDWPE2JA8DelLJjO0L37xEUpOaxGOAFU4Ayky55Azw5TzXUIA0wnIKoVG9rWg2g3xG+/zPEhf
Mtx6Yktja74g2dBMi0PpsfuAjH5XaOecsetwpsaVA0KwSneaFzkwlgLv/5jMydjk5LiG/NrOzCfk
WP+sLlMDJoavpJUnYuZztW+ybYD6DPNIhc0ce0eJM21G93L7m/2mEjbJA3XWLrA4qcjh8CjL5wN+
CiwtJtoA9iH4Xa5GmodhapWHMC/wuYPAibWmuu08VapwemjKfGuTMEj4mzxtFNrncxp+Zqmk4iAU
0cCxBv2sBdXJ+UfyAM+CQAI2Q+d+Lq4vGbkrUseV/t05Mpct3w3N4ea4oD8QC2wQ4CZbqp35JfhV
YFNKAjrJhhsUAEqtVzZoaGKsODC77juQMfGiDDMtlWO1ZciceisI6m7ZrHeumLjUmrDwhKjdrsk1
uvabEDbXY4XwS1Q8cZ5PLsGpuymVoNd+qNbyD02W1Cv0YIIzygRxcrj322hVTJORomQ7WYeqO7uM
SMDf0ZJrRpxP35H4PYcf7rSore8w7CL5q4HVlEFJ8dL6jnMrOtzsUSA/KU57g9/SxZxFY5M7KZzn
FG3uFhtvzDE79e6l+VMnPXbYWdwmHPUEGcKypm0SUvwlRWvcaJ5vDPLTCa3WTneC8JOKcuT6AV8I
tDHVxVpKOCqIqZJOFLQg9CHIJ6ucZo4GbP3NuWw665wYduzJNF/+6m4ulPN2C3TH5EnTXJpdJpVd
IDVDbRfdOywROT7t/HwmxJxgek1cU0cNj0rkTh0Bf3tKjhdeCEVzEXOBFvVkTtoDdzpHrBMME6k7
zzRksnq2qaQteh2oeubG0e6DZko/8Fjg3b7XA0TOtUnf3n+odn80o19D9RozKjH1nCwj6m3PYDTt
P6Phiwj67UwtHrBw8Nk8UqS+knV8pMMx4yje8L+jIAlZldtYbBu4YtGL9Sn4nbXWQvdJaZ2iz2u4
cfOeBQ1D1PJ7xq2liNe74GAX4nNOhiFpgimVKBRXgWK2RA1jsgbtJbKvM/7lukuJjvzJEkbRJDX6
6ZR+Ic5YCOhASHonlZx/0xtYamlysEcjkBpd9NRZqy9mtiZyBnMEN3R0apeWhiMohS+HREnkCd9L
/5n//f1mj7I/o71T7jnoO2XQYmWvqkftqCGYsbcGmtnImfyrQyOHzvsTabxl2EPcH6lUTJ62V8ih
eyOcopIxGZrBa4nRH8n07WJRN+lyj/7NIvmsem64TGGIolFVmjDr5yHaw9wdJA/bOi1iPet+Lzt9
n+qjxExbz3fHetbQQv9THuGfT1aVI4HA7k8l97XDLjyBvGVdkaKfT4Au8+NPoN22DzdubAZ4T42/
yI7n1BpvmUjezasH6xXEAvH4fB/Kr4HjnphLgZsdfGshN+qSRYzCEckcfFkVvlKIN+haf/zlkpKY
37W9qgX4wxidDTrDBhHlYOzJADrYtPwp6O2Q8AEDOgq/h1qd51sMXaMku5FWDqG6p5dlj8CBDDMs
yUlc5+/RwNtbzvnxKWAdpUPP9IP5yY9fbzJrkVZXNbLnqCdygAtp4mXyF1rgNaqopqhU1yQICCY0
HhHPtvjUWS38d5Klc5tfMkPXvoXbdXGy0HbWoJDl7d1aZiV1Mg/sLw/oYgHmjsoGv8PAS8DbRVGn
NqNruq/WhCPJ+kCH6lna9Y7STWCyGgm7N+7ziJQ+T+A13inJShNxlWLRRb+d3/gh4TV9yA4Sylxt
c9S7U6B3Z9Am86kmgmI/JE18uFiYHsaNfWBWuG1/rSJsRYcUk7vCKAs1ZlzI1Thhtp3kmzqLRZOg
oImIi0r/4YHKAHS5kEwElAwGtx1St7ovaH8uhRRCsw6XfMKnN5QPDdy+ytDtfmWZyPmPueH3mgKY
4iws+4qPpnF0iJfHBWBZEHiHkjGJNeDrai2Mziu+N3Us+Vk3oe3wk6yr5Osxz+gH8Nl9KnjzzYg9
u0tzwIB80zLg8AGcHr6IZAOtjIht+MvdvfZ9xXQCjXb0ja3dsiLXz+bogrGyxVG3cr2L0EatietY
DuceCOEg+neffPUm5QFlV+2W0N96f1+L7Xt4QvdZDrxuyUtE0Lq6WoPcsBu2jRwdD4pb5avKG7Cf
+Am5IHTHnHM03fNwyx89LKxn3sWz8sAKzvgeekvK1AyYD+ovQHeThvyvKTJYVqEUzYydJFDMB9fo
FAhWiTla7wCjSltEVib1VHVEw7IwheZJuI5/3UoJJGKDEpai9mjp6yLkTnqRFAw1HTvz3yTw12eA
F/ryHcZ0hiisiqlMuZVWpQgFAC8LayAjHG0UIGrLJ/giTwQdRzuZeQvX7isWvNk2EFFfntyURXK/
BJbo096cPCZLSCTtg5dFm7AHeMqJna8oYyD3hDtaFoABysevJTcz4yqPlRf/F+xRr85J1I+KOFwV
+VMUyxIdIbkwfVSSA89ROc+tM50bS5QzFf7PT9Tcax3bpXNsN+AaOwsAerMENCVuB+rU4pf3/z0O
mMR6rwuMh42MZkxupbkVnN7qFpSa+lUND0dgzLAcvY+bGYsUuv1HiVbBn23NFDHYhRigg4Vcc+oy
mET2u96Z++zo4McuNeXGZopUsby9WJOpMDqKiN03PG/fAbSAG+G2oMEuo55KBfUWP8s+KhgANRE8
cVlzLy6zzhcDSVg8wfRbtnBMsLaJGtEZweE0LcvIDgQU+sHLKpUXSZ4Pi0i2Oh8Gh0EaflVUdVWR
dFriUvZSVR6+Ikyvq27sJlMrFQQ1GERFJjVHCtqDVkcLj7WwjBjrUgJFIEqGFxdbHVFivH0qG2s3
PSybe8P11x6I9iZ0TgrdRCrm+JwC6Nt4yDeNOwbmlfeiMURYYGcZE6aZXVJxa4Wepj2ctVHcJqAk
5s/pLZpihGHNJr7ylBYSHX05a1ZYXPntSwBRtJoaVxIpDKsVqGKTIf6+ks5u52sh4YQo+BncDJQY
gGlBmXjNkdmFNHZlC/eckgSLGTtQR8iSC456ldsmBeHzjcuj6A0lkeKJcqTTsZvoO0weWTtDm7LM
TRcQj/jr9eLhvm0/4ZrrWGH0duLtwutpBDt0UtX41V0sS9RAhIIXeGqfPj41U+rA7EES0AF2WXdX
z9Y9rI/UNU6N8cHsQvqd3vkJZrNFIrfiLISNa5X/4FkNrXeIuTHwSJv4a0UfKZKbsUG6WqVVYyf4
GZBx1assOXualyOi5FzB8yrO5ghwJ5YTwRhQMyzZ9jmIYltlsbpRixLvC4bWGKDjmVsR5wuxRN8T
qIGzvY/c4YVQAaq/ZMZVWMLIBPtsLwbsfi1BkNngJFlImZOboZkVgYd/IRK4z0O5MCgSbuu2KsG/
WY3GXLfZhKYNyufYYqkDLLfiCg1azp4+Uhh9ZAiYwQ5P6RF/Gm+aPpezTfHaV5px/ihP54kgSnhN
LfrAf4ugBLrcA+cRN/pge67V1nsu700gIiMpOXNXKpVRhiUUGZJfngUuVMo7xcZqvP73wqLMPXCJ
cQypFiA9qfvfoUtnmNOS/MO+HsjMStlUZZ3r6m0vPLwjHJNwXRl1REAzCjDQ2EpldquDCFah9tXg
RexF+t3RcPQ/2sysCYJtcpWIdCMKaT1Rp3LwBrBhaHxezJIU6mEQFwCYoNKlK17aodXXmENo+Blz
GAO3EnZT4K05E+VmlqefM1t7djpoMa33BsyZKr7fXe5uMQUZJifgHyhEJszHZmzFcYZoI2O8HvFA
B1Pq8jbRISpLbkVMbCrWGp1BiWLWwDiHvYohWa96+lxyDtYdDI3Wg8V4oLJ/G/BR0/caDmXWJ+5p
GagVq/jiMtDkOFav1OEuBiGxOb0wQ5gE6G8erdR0QNfMVk3L+FFyhNzu4Ufw+kXmCA9HowlW0mge
9aIFnkwFAQG51wOQ0p3dpF8Kv38nobYGmcaE92FAYdJD43BVmnkS8PycVBUovMTpDrd/jkRUI9xJ
/Yhc1cbu6SIP56/ueeU+KAi+rMizGg6z0mnfi3L5lY8UPvVdqYTFZJzFmBIRDefz/KO6KaUz7zK6
J57CMqAJcwL39xH7Mb/YX6lh7x23rNY8gfh0tG574NijJyyhyjWQ3TVXeZttRTMQ8EkVZleXG4P8
9Cln9/2k3TDje1sjh3cwxf54LOlr7XEQhqTv5J0oXe/Pa2JWradNXJakWCC3oZv4Y5wIQY/oigJB
YU52rboYWwGjtw7aQnH1lwrbTjq15uJZVY9dJviytoarjFFMs6K/cV8074J0zByx5U6ZzdsRj/Vv
7v3J97Ntp0snHPbSbVdrdLUXPohiXf9pyMa5n+RNlY7ign/cjSFCnP4r8aqyXb6+mlGFNYCEjsI4
XY3qfRA6H0N2D152V+tJI2Qa+/Qgv3HXK0XhMB6tFZPm4oImU6WVu0BmFGs2Ta38aWUQ6hxo/q3u
1Zg1lvYyLConAJ5jh1zjMIxqEI1Cm+G5aIgYeegM17gykOmppgTM1tGfSC44508QE0zwMFtatSBo
Hozer8aLXW56bt4dTjL6M3EbVsC6LtqU6OltrPVALWZlqkvxgki6U/3vOXgYuMHSHoJY4TfWHtds
6gD9H1iLDCaiRZYOGfvUDYWoZWiY8rgRh5uhjb7qYDPf2Dhd6bxKZrlc61V+z7AWV1OK08ZX3rVO
JcO00uQEbtMOcOdU5s29kq+ApAbvu2M/YS+QC2b0Ph+ApNbCBr4QHH0ZUcGqagUTxbPK1s+cFG6w
DxX+90YQflDmM1Xy0L/XqjGJwxbisgLGIo8wHazRImvYFHPtovsPnjQ7Vyhov3Xwms0serwnNOdz
XARinmNrJGe0MmNktHakZ/DKHBpCY55OEfiBQlx0wj2aTL7aALGDA64JpzhqdWIqJds4p20GDl9L
tBWMORbRrg7mqzNOs4+V3VhX7NbM69ehfdX6tdVRxTk0GZ5Kc/VTmr+o/s/v7owAL6YMv+gRZIBs
sqmyKfGWlzG5vZu+jnC182meYwYvikPjlsWzqfNVNs0g7voofbdWcLdFerugsh9KlW8N+bTdLnB3
myb1GfyilxXeRactCiwh3NuHC4A3E6NSMt/shNddxllAEoR4BRF6ulkDjl0W927oi14CL7LKw1Gr
uiKPDOhSQhy9PaDLr0Ff8/3PEQCiyPOzI1xclkzwc16BoMNhB2wU5S7eUARTFqWhikvHTwgUE+ci
rtkpD4vkvd9X02KTA98Swt/0kwQxpBFfzZTkBygOkoWHkglQdGVP40Y+zPgyHX64klvxcuA4HSL8
QiSgE6PpvzvPqoe3KRKAg1y5ino/abvoo6otYmbBMlPF2YRjuQuggB6G8Sg9oyV99DWqxfee5Bea
TrY/I5bxkHapl3f/dFxTzoyyNiUMKQFxjMrYI57q989Rc01j9b1jBfmSvwtD+wX0XgfVuIFNw+v7
ZMV46wTQH964pjElLRA3/Pz9fU/oF5eJYSNfJMuhfdfKGZdgZ2RiUbWNbI+9Rb/atghcEhni02YM
XL1bU66VCxqiH0VAjqDJfEuDgiktGTmrhK7zWD3E+kjnoeJ1AjcfCmkB5v/CPRBHUqvUXIdmhG8a
VGnFKZUiqnpQ918AXbeEWA1vqugrDzmGeXFJYQ8ZJ4CJVuTp1X6LxyfPdmXu5pAUdW1ajkR3Gzkq
mlt7xvaZDLaOGTwlW09UYU8TvttZUdiBMSL6T3DORvxP1Z7HfaBT6glmrnJ57WUBkuec6uB5SIrK
n9noOfYryqlH5Xblq1dXNDoUQEKJOF5at+KAHDNP7DdD2nMXrH2nl1e/r6Kfom4PjYiRj4k8HzyZ
YP3uBFJwpHnF8ebrGjpnFhbs0GvP3c9HtSNQS4qf9+nxxc7ZL7P9/G88qnv7f80uJR2/YlblHaNB
QewnJkzP7tB4BkX9u93w2Cqcv/mPDTADITVObBt18lpn8HdU0KRwxgkIKjjWDxhz2fvgmF9K4UsW
q3TkSiVkKV7cx7619UsQZIfxEq6W8n8qlKsvMavxP0FmhScW3h8yHbC5DUAA4QAA7FZ/JyCbZkV4
xgnnC14DWPmJgIm39itLHYsDUyetBbXvOQVAZwooUsX6Jkw8dO6pA5IILdqqwZvsahGz57c7FGmX
X4tkeba6wo8F8nGFZEVwvjJaZdDZO/Aw13kFFzFNstGwkyZORtn9kWRRRzvkw46S6tFCDe1zE+V8
VmnbcnZQcoEY5Ab/s3t/QFZfBRZ8jcilzIdcYL9awU4ScHXsE5iWIBH7zksToMnfW9rmxwoQxzRc
wv1/K9rAFQLABwyvRiynagdIC1uJOpK2rYWySz9EXexrT/Lo9mvmKToJHB9i8hY7v0/oaBTnReiP
KaL93oHKf5uUCZnuhkbLkI714bERtRS8VAmj+XMtnxQcbXiNhZOqjljCgPxfE3/qso6+aCaPcf9G
sc2lj2y68bgj6EB7tfaKo2wf0vhTF48SfNt/bldBkjYRE3pLpDIl8y+ODnchuHfH7tI9RuY7dCtj
5TnGLfVNvs3aWbEM5dTttL7QLapL/LeG3dB0UL+XCzdpfjH3gyvI64wnLfkOxaSNgW29OUPbc+iM
6knO9LtJbJZNAGGm+swwAvf2QpLAlgCGKy7B0TPXbUEXrBWZ38jNn9SBV9ql1DG5JfqiFRGFicD6
u6s+2DTyuf4di3qvAG5+fAwCD7hZQNGaFmURzyMAnoXHhx1TryIY7xQ9qEIFgkjUJJMyEzdM4Q/b
nMmkBesP12ZDuKfZB/hV1pvceXWj8XPpINFqSjPOqabRuXR8u3bB9bNdivkgngO3mXAjwRbOmxdJ
2PdyXqsagu/D2t73smQ/fDultqwNu38OfJgZ1osbhwy+biOz6QBoFjvr0+pI1S5kYeGLmjnWDUZb
r3y2+FunbXuRa8XE4XJf9G9e0hrg7CwSKgeMFK8Mi4/p88TBEs5gPbl78GlpojXNsdBa8LSinelb
BB4mBOEl0eNBIvK4Hk1ROTnJysaNfiIlb68IMgf+ydphNJJW6UvIl3RD2FDX15gyOJ9kitfgxl2n
Egy8SvBcQg8/pz3lMB77zPfIQ4G4xNpejZI/3Kgc4/AO6zRViwUSUsrQWHK0WKr5cavD6yP7mmRj
/ucF4XdBR4g9/3jqgyLGHeGkmrQ/LUjwbBlrD6bCWQdplqApd8nIbpD7b0Fllt7OUlLYo1Cjo6aZ
pW3G6MFGcmyfg2OMeUVT1RnF2/AlEokO/Jj4sp6n9UHyGukppLWoZT8jjL7LDeDbfGw8MuJxzyW5
0NYp67K3irN9/aQK0B8dPJB28oh8kITyhjLUdFjw/Fk6YvHLKgvGlzjp80V++2qd/e27NEJE9lxj
8b2sBBPgdofHzl0W6io8t1TzKChxA9HUMlgmaHoBKPniUK4kr0ueYGNrE6PkXty/1eia1pIWuFMN
LVXWn1djxD1SsNoT/UNFdrjeLA7Jq6n20sWXzkQ+objklB//qSD14OpAbqC/S0IRF+slMfNM4fkn
cc3q07WYWDsNm36+AzDsC7emPjwfu8dv8Xm+2CimPOmSpPJzfdLMKDPKL8DWdHeuTUI0mace7mlI
64KSf0+SdEXnpb17aHQirSsrHQmgJaY7icEeQF/P03L8hPkUMQ9TDNF8agKWnArlL22ou1IpEGZ6
pisJWThrjoU8DR011cbkJQ5JT6Ybj1dp2l35JPM4rmvQsojitxLPGPTJ3K+lK8sZx2uyHPFADeIj
US34EWjNvD1En46svXVfV0Myzk3FAwLyqx7zsI8eU2+e8cDcNwjGeFsYxkZqXBp0i77Ryo51Pt76
1ti7Bx8PaP7AffgczRcjNE/PrThcQGA+4VRIvLIjPNv0kp+vubbCpa+XUTY60KzZHtxldcIFtPqO
9UMx2Y1/9JV2q4iEEQ/G2ST9t+WatODvrytiZxEugnkIyRtm6KuYCbzHSzDQh5AOZ1FtyfecoywV
9Zv2c+iL2YjJRex40KA6gZr+zRASPqtGsCjeql1viq29f17m6Akl4WugpH0xlDVA0p/sxfPEIIgy
gb9aVOkzzHWgaZdqWcmM+aqQ1bqv3HZnn4P8w6Ogx18e8fKAtmA4EkPK6YjQM18tX1xLvIZeRU/Y
Qy84VBY+6eMQ+HSPvzxGF/eb1CezF7O4uPYLzWIzEPWdu2mRjs3yzf00+lzkrHMZrqZNtSebjEVB
aoC9orL4lN8KCb7cPFRhTcXgLR5IzoF5im9VXykshlBew5MEsCBfOpxN4rvOwueVFRQdlPGMp0js
DL2n9/NDazygl8EONnDvmCHuKwvgYYwuI8tbKb5UzbNeZAnH1E8nKMzEsO5eHHLEqHaxOGlqmxyS
l+I2TdWt9vDv2diCDGNNAPEvx5+WfPiGsoUvpShJl/QCKsBnoW/g+xnZ7H/72vt43PB/jr/GZYBT
lh2toyo/4C7juhIzQ2ZoIXdLccREF4eTlTnIrt4CZJoey0/ztcvac4eQKDWyqMIrs7I34gcfPVbp
tOZzhyhKKq3DkaPpDwD6DOS43p+9gNvBkqqUwUnXuEXlyZV5CHYMtH4+lT7emoFzOkqn2+lcOSZl
ixj79UU00AJOqrH1AQcv+dlh1YntMpDPgc9ldjqIbRg1PV/kJKv1HARwOmeDaK5Uebh61jpcqEpm
o2ohvtCnjKWMhYv2E4J+eH6PtXfeIIdOa3yWCKkAcOLFt55a6QWApcT7U1i/CyDef0Vy8Du5HSCM
xAyABaGBk6SRqS9Xgjxre7NBXo5GRroIyez19KEkgLHKM6rw7EnKdBmWa3AnVNTuEjtuw6Zx/DZE
W1faDes3ijvKimFqlnVjI7De5xVMwBhKOabqIZxY1knY7lbGn1BlSN7/IfA/qGAOavSkQeVFJ9Wb
lrD78ii+DLVJ/WJcIXAQHmDNmo34FAhFwtZyGBlNgWiaZP0o0RfK2eNF9qOeJ1sLljoGPWyEhkyH
IAfgNWUdf+9EnI4fXF5wDHLugA9j1XeTh+XsFK/hvFDBip0w2YqnESFuynfKgsBAR75sVAzmYnuB
dcIu+cjnBt+ZJzzDFVCG6t4P8zhP4or52tkeWRfH8Vp98lWOp1QkJZizMvSb/DxJpmO5ZyvjpD25
eb8EYc0RH3qDLeJuU+S6B8rWVcCmz4pVgUPUjxWHlprbJKRUEhuc3KbvZ0R2uV/a+uF2kqcEoRw6
XX1CPo1WAJL747JLwEpA0/7Se6yo8N/6UPD8Mv/992jbR65Y5a7Xmlsq+Vz9E5eeKLEfKAnTPDCO
IwDlpE7/mWCRXfLmAqqcXgjxhx5QkrudqZro4HsrWk30Jz5j90nUrMvQlCp1bcUAh3q4VF/e2IUL
3SZ1rv92zfRydd9ShmfuW3GVsZN6hk3kjOHc3aAzo4PO8sTBEErYt9m64qkfe0hTf7Evu5q0QH6Q
md/t3DMdF8vIIRKfUfTUUdUm/Kr6qimndyx8j6JPky2ibjZRuwC1HFLjUkWWmGzbeg+kl4xrj5aR
8zBhK2Ce39IMcqjUuNsvY6o1Nky4HrHIlhkn2FAOlirafh6tItPegmcJrMAmIWWN4EzoS7/DvXVc
rCqL5hauueEFCz7HA665nCcNXaMHj9gNHArf8KT/vRFJtQnEUCIQZxICD+FcNdk35IrluU1/pS1a
zdM89cADoOSkBye0AMvRSBVI3gC0McvcPVDyI3NoBTDZ+gpC0jsxkDwAi/0cX7NIl4HrtgoPR3uk
fTkMoSFskX8Zzw/QO8YfUPuhwsqIlknb1W6IP8Lkc6qrdoSOqDqoNYABAtuf+MaCpKqqPizRC2++
D2wyD/t2pWJSyt+G6glIuQql9g21gla6gbMYsWNuEOD5sYXIw+0JEcmFFh8WTixFpsggs3PGpbn4
uyHPLb12HB01RTltx9btvitxbAFCRthyj4V0Z7XULhDAECv7TsR+oRKizr4wzUN3twBuasRi8Zf0
gpF4L8YwNulRph11sbua6eRozUzZBex1hqXyWTZk2rVUweBNHuArLSaDFvUGwqutHAeggwetZMMH
8GuBDzsi+FUef1+lXxHxCeDuCgYpl0pP6lZDtKn+8yRh1hGpnWVDgGs29BFwg04PcL8+hdrjtNia
vDuMRf6/JHUhUYfy5HxZvmhJyZy83RIfvRmBuWRErbj/4ndWgt5BBwqXjaWbp7OzunpyelRG36Rs
Pc9NSfaSKinbBRvfSk6jw0DtbOpFXy4fB/HNqJ6cJXl3NiK+sfCowpFSR53cJWQIbvCsbjq4BMqj
78oEvS+UcH2y7OEULCyKT90m7kh9NqQzOFJlixgdl6Aevb6ZQGm6VjnJMZzlOP8nXIkGKA2ofC+Z
9QKjNvb9/J72y9UmblfS5xV1KQgt5pF7eW8SEGIryrbyxWIlY2rwb62k7L9xO1go2AbKPoL11+iQ
qhUm7jFebCixKtHAFEQrduHjNDTqqBSkwcjv4Ua4jNyDTOv4q28WOU5vdqScHmTF44y1cyi7FlAC
sPvtMZLFW9LQgFkATLsFJJNfGk4FrhfxqrhUK76oSMRrbZb8QkQVKjAhp3gqNFr4KCFYrmVyrW5M
PjpavCcHLeDFsUUiqld+al8OrcZ1irAOro8wWtqnKNaVGEK79nVEKtOvOEyFdk/8kLJJmJ+dzTP3
Hxk9yWzx0XVUE3eaKK7BT+oIYMqPttu0AXhuwfEqeTUpesVVnFCLorsiz4nJ3yTj5oLu4Q2XowLv
FEc2wPA0cTyd9/8DlGC1VrxBZnwFZNhjtDqce8o4fi9j2uEVRHLSSRb1zovurBQKzx+ZB3YBDFWG
HsGDMIGQfEA74qLkW+jwWMb3Km+iixD4Be+V0zj1YPwCldMfx0rB0ZQPRPop6pORtDEkyz7I3J3C
TLF8Ha58GLpDT14j5JANuP8OL5W0UjKIw6vqIJDvHP1SR3hGzFlBeKM4m7jMZcGIb/c9JXgVC5VI
W+5B8ZF9Fal7q+CwA7uQwoteUt202/vKzxRmABXs3vCtDcEnrDo3+V9SZLTA0Wu3TNLjx+hqJpNz
EoLZ2uP5D82TT5AyEWPnT6Vc0u7TUvTdBLJKa4hZgaaypL+jYiBEck61/HF7U6BxFcc3Lr7qudhF
wcyTzBYw3zqlEJX311zH4hAMaGVRRyFKr2Wx9imu5pzt1cvdyao9224UM+9+xidxGjBqvH+Nh1bt
fPdlMvEnDLtRzALfxJMheAlQbs4IG6pvPj4kbu1aoQXMfkOrJuFNUI0uaKPzqc5KC+JSbVx9TAzF
Zkmj8UVbG8ISWFho7jCr4J/MF3kS/xe8LWuEQiqEe7jSWvw9Wz9zbVJNWDsAa3E2v8/Q1FPNE1fA
JRSoZNDhGNoW/wyCnwKxUQ/HcS1rhJ0PQLf6yLHahZDZy2EXYeaTLdLsnM5p19YRp0Rmp8NtbQDb
P0t7SIiFkkTTHbZ4XQaKjYZX2DrcABTjULSJaGDd/b8zttcOck0x/TjrrNB7/ihphDftFZTTPKcP
Mr2v/rlPYAZ5pEtxaO7Ij/6E/55cnN0+3cTeCHuPGbZBhtnHZfN7q0uW4q8ocpO2AxX4zWz2fC8t
7xOo7YwSuMI3PVj9btybd3+a63tFyXCzRjZ5pxwonnFj8c8rGIF9/eTqWrPCAllit9+grfHch5xB
cQWuQPhaeY6UNxGn2QGuVJQYf2REDsVnQui5Lv25342O5/ur0+Nnb/p6booX4EpgTOlONssha6IU
63Y5lOKVVS/hoP5/uAiMpG4hl/v+i//e3kOPMdGh4MHyv5dghwPWgrFo2a64c6kbdndWdVjTgjtk
8q/CZePcet8ettN9SwoCC9i/9QK2fbKQbHcwSilJgbvYHYk0Sy3Yz3PwRQRnVzLjKJXCHQ5AJY5T
0Nhq4weybdCAqbW0BCANnbpbG7VWoSp8kZLURPd4jtOhOjeuAebq2/cxm2IspiWy7sb4W8NGanbu
u9074DPd8nE93tYRrjmkWwfLN7wA1tJGXBqF0ut9uU/Ej69C/53AvoXo77ZpQm3xb/gdXRS4R5Um
WjRNCenY84tQP/olgOMgwa96p25juEW190RTU8fLy6jn7MdjHr8qWGPhUeU5zeKVvPFDJT4KpqhA
Z4wk56shNdIhY7NeOPvrXfFeFtMuj2ntGfg3AWhgJQWEHJhYF0RQL3TovvtK3Z8BtxJDuCXzMiiS
1dWbYt7JGzPOg7VYq+aeknAfaPOItvIXqmcx04lQNkvcYRGkNsU7gCaeqxsfZB/1i7nn8bdBwJoQ
qOvwu305pcpHYhtUsHnHX2XW6enbIgiI7k1HmRy8BJ9xyxOHwPoAYor51lfLhKGJ0jzFoblKpnIM
14mJNgRUEGMkmJGJcYEC75chJ28XzcGOBakinYhVYcqH1hZ3bTCAgHT0WFz/c2dTGHj8ltJ/bb1I
lAMaEej8l050EJDcNXjezoplGlR4s0QWU6xUsP/iBs1mlOXrajFJ6/A1JY4BX70KRl+BXnH66weN
HW7YW5PDaxSWIv3Cbe3FGZennkfnP0SdHyiHRqErmL6cHGxr+Es6lSP8kGMhY2vbQ2oNweImq1jX
m6Poa6R7BrDPc1gxHCfEP/nfpqKlaMgSDCpLOMkd+EPHB8iltGcSS7kOB66n0dFFFJZzppt84QJX
IOHZcK2dxghVMW2m+tw9jOxOeHBtWs0PgBFcvw8NdYQkDHF59wrS/fAQjeCD7tnTsn4tOrpMs2IQ
T9WTe/5S0OGXmtn4KfJsG8CqKeCUVGwN3OdS21w5UspU3dIhLCIa7IqlyM3WBgCisixDhQCjMksh
6t1QhgprFVR1Tqk7TWeDs0CGTvVUUctWc9J74sISSCBj5T2enDeksgOZ6jzVb+gRsUwFksVDd32S
BcvVXexL81zs6al1Lakt5mzCb0nNX1Ki3RYxhvu7CKaUwmtlUXCUtNi2Z6ip21k/11hIJWmZVG7R
RPhIqTBAFFLpCNIFEcp5TWahPyeUSlJgWiZnnInLZz6IX89Olp23nEIZs7iwJmSO9nol5M4AOWjn
vw8hbzbob44IMc9TyNxY7bnrNCVaGm3ZzUzA8SoVPa0Eb9z8IfU8bp32rxlt8tptFCTZWohaG7NC
aSgjnSweI8NtYrIO1RAKiL5fK6vuokakLQeAfF04NCekaUTEMiVs3JNIcz/ksnmsUyydA8vEBZtp
C8J/c8q8l7IiHFKTeOgx0vfDME+kVfzZWYnppoUqiCv/EWoElkXWN+lN1xxf4fyoR5rG/N7xiDyM
ofFX8scO9WrmRv0cRW0dBGjYvCaapvEdftz8ebjvidMO6W19oROnWG0OvUmb3l/OxORP1yLAxCYz
SzhKsmqO0L74xTv5e9fd27mvpgbMdYYG469Ft8kpLhO8BOtncEfoQRUJcIVq8aRq4Ohvbfugkd+p
XW6IYDxnOr+b+knLUYkD1XN1JDX2pLXUQeVaGKPp1tF7Jjxk3MnT1IMND8vN5RRkd+XWmQv7zpaF
6ZUp6SoH/8J2tQQaB+H95fGksGC2Fzmku1y4zml3G0gd2qVECRfTk++amtykMYxXcQPj9Vutfmv9
dtr7/N9xxVqi9He0TaI9p0MHoqwgzqFejZer8s117L0vVzrTkltvEhUyKN9DegwUKsXUi2oB6tZq
URWEjEzjzHgDk00XigICBpaQSZYuiZxELxV2Et/ycT+p61XovOygo60m9qxf84byOrDU1E1RAuYV
eu9t2qH+p7Xm8BEtWOy9lu6Q3yaEGGqsAti7kkC0J9h+S5vt9NXIh2boQcu22fwDZNL8deV2tMBx
RpURsQ2RR1xX59N+t0c+k5iODTiPxsSPF0YWwxNbt1O2ZX1FyXIG3XbPG/AexieLJn3lBQ8bmCn7
eOlSZTUaGYSNhQfSA+SMVKBLHDtR6XiyoWYDqePY624bvmHY0WK9LDKl0AB8sSe5yEDjIEPdekRu
lEZJUUhRlNjjI1k4KUPuBxjdDSOZ+bm4e+tjpIC7CG8ZfbEcmNoYn2cv5Gy5E6eYI+oo/jfCkbtC
OMSi9+CQz3mPe7EI4hl0dd4iK7sgUXhE+uNvl/+Iv0SK3bUzZGVASRtU/CyJIY9Twrr8ZUhHU9uN
q9c2tWUpJ5gd2KM5TZZDK+tnH8ectzBZ2RIHoa6CTJpSfzY/xLsx6uv+yP918Rzchm6FrcbdV6s3
KBrTWjzV8BtRU2zFqtMCDjetk1i6vuRB6qJ94oQnnxBUErBvGY5QNuNMgrxucn4o00qszsqqZ/9v
Q9wkVhWSQpcVdYUo/oYVT2Z/kXCdzLq6tPyT9oEgeTa2Q0CeOZ1dsbqdM+bnd0SrtZ6ueY+t7P/q
i0SCHaewHcvMxNREoLyDGeXxQZPm9aEv3mdR54IMNd1NtuW7gRU2AQEX0OtpbX4JxetcoW2y+vZz
iMfVKlXDw49jDOZZwrQxfl7QNmMwElseax2xszKBRC5Dt6BoMfHCtDOoEKfydwwNFh/K5r8emx9T
2NOj8m7aPlt3Y4f2UbyuuaipPnwvsMSEIlzovahZoT38sW39fueYhaTwZ42CpONC7HsOL7+0iDz/
j9JdiwCF4jK+nRHVLZPXvcXKf09gp0Yzb1Yyz+TFf5x78J1ygLGlofyruWgY8HzXVoPh8T+pqaGF
9qnlJi0iJs/N7L7Pi/V3prl5MynazkULeVAMSh/7GHBpc0jZqBk5RnUOQnpxY+VFoiDYKpuN/n/f
m2tF4zqOSZodYZeFbZg6NP3Eq97RqHYA++IaPNNjkk6Vuk5/vCMDr7SYf8GremHonAd7XwySgsAn
dG68BD1RtihUgEgz93AdvxhECrznYBCzOR7hPmgZTzVv/egheKDB8ZUXx7Ns/J/dhZIJYs3p7xfV
A3lzl+vZ+rdeURLBZDzYrwnDtG6/60No1gEGzsG9MqUsyoMpjwGPvAw+2ALhJay82aXUG026iHNj
730lM+LVneq3V+RzgEB9Pe6jm7NVT9N38K8q/sF1715z5wpqCksPjf1HaQHYtwcKN3LHABTuJoru
N+5hPVhkqpwwG5HXl6vS6kjx77x9vvztRjzlV11Nl2DkThhGDtMl3gV+XZf4y3e2X8ZOaIqPItTa
RPPlPCTkn/RJgm92X6EpnQCYa2Ft4IVYui2jKqWdwk3gCCkzNw/eAZUPIONWnT+vTBctPnx90Chq
msZ+0gb+yIeWI6MyCG81Gwqpnn7c6qsX4SuQiSVecqg2o9rfcJDuibmI8JwD5+Bc2k+yY/JLfW7W
XN0ki9ccVQ69Vrx0BUVP0HjPbFQCd4qyqhx8Xx4Rs0FDSQ1TlOzOEr9sPZ+uYXQIN6UKWbhbnRMA
7vFuKXCz7Evsem3uUqX3Hl2YWtjldF4FVgDh4rCRJyhHmbJxBZkLDORjHv9tGairmS2sb0fqIgRh
9pVBLHE95Gb1A7LGXU0GbxKGQpccH06bQHhe6R7ZOHlniO89KCCG2Rka9OVKZFhJceBDHBMmWD9s
h8e74tgGI0Fi8TJM86iutQ8ZP5SnQFMxjz6BqMVmNSAlkTVGr7LSf3FmF9eOG9rk+ZSgMM+DE48i
SFac2V/8l+de6hY4vR3jJXvURdZCWjN62DDOF3thRehaHOAQWT4rAJOxk5BfSq4BUAI38wsVKfOe
h30F2GR7Irev5WHI6svFmNaL5UIhtAD2rS8cJ0CD9/BH+rZWEuhbs9aahmjUzMm5BgS2sOgOnmzS
flpbEXu5/NbAXtC0yCoGakWeUWSgSY4rh/AyauFn3hpjujbyqWYW6AgsbBDoE/8CeBt++dTMmOxB
O2aNhuVLtcxMLw6oRQ8k9KPC+fTTv6aJVYmS2+1p48bIvGWNu3p8aLCEjK3A8sWmr7Jm5xpDElc0
MJeC8mmgALQM7XDIU917ZWLxi7gV4q4AS4oe0o5x4HpHUW3AnPk089EPknBQwyLCKX3FButFB95f
v5Ge9/rwO0Y3gtLrclhXBwAOWSqIrSvBaidVx8Zf38pvvrOlo/4peirpAeSjZWmU7wYYp0QwOWI4
Qe4yMj17mhXngCqTX2ic8n942JGm5TCwFej0ip/TgnEfWlh4HlTuW3iDBCQF+j7xNyNPrEFd0QBh
1nxHbSwNWmLDBBCQDn00seUVrweM4bpc+KCB2Ptu6ekxbB4qAS+1qxf4iB6+myIzLSrsKwuKTusI
zFK8NtNzY4eByX2uSKRLpICtbA+CBil6E0Um9rxIPf2enPvq8KzLpTVBG96F1KArCzXY4qAYKDCq
ISvn49WG3snnr0OPEJr/tf/8HWblQ/E6CrpxBkQ88H/u8uW/3DOHX2mfL3WHLZs69JtQxmLtQcjN
+S4opFlxmY7dhHkbbbMMBnrPBumxquzQ6hJWgDFZtFIeRGEXhtqBTb2damv6gHUn2Y1e0UMF9zpO
VF3j0vRTZ6CE8ovbPgeTv+QLAAsPWzVq6zuLi8pgamThNh3nWWzDiHRcxN48jg4QuCAq5XzQGw5k
G8MafEkhtggS8Tcf+sDbtURg4N74gZKxoycUOT24EBuiJzsGdZoAXPPZWfRmRfugVAwwM1eU3iIK
DVl0NvcgIr7sdN1gTmLndL/ckLYpOkPveFgix4VZEbYUQJFlIwGbJO0sYf3gP3WxSlwlP7q3JRnL
e3siIJAEwb0xADMSD+mJ0dJeN3qS23z2pwO1V+P3m9sZDorQD/kNCwd5M7C2H83zzhGyAfxuE+eD
0sJ1xrq36CJETa1dznA0fvgP6Vboqns35Od7UARY1IkDK9tJyfCISYT/w7eTjGXLZFOGMGZhm5UB
o+EjkKIF3ocEp/OVftNYkkpRcuLjniXrLpmB/XSCH23wvufCFFEbWMJvV2ix8lZb8UkaCWcdN5Dm
HbtxgyLD2PBaLf6UmQyEORAi16eGnXwksXbvR3wVl6ymF8j7ZHFDdMTYrwaCOY4J/u/Rg1mqxr4w
T2RS0Qa48vzw/5PhQlV1Z6S5xCxTbjtFMNADVviKw+WvrscXUL1MCzShHcH8Q1+HQ/0n0zdCDcE6
R9HSfS6CJw6AnBRvGsKi6CfrxGdMvKrsVK6nH3RoOUhx8FvyMlobft97yfcw8dwbHKBdP1GbGYgx
DSImMRZ8VMtLKZpK3YhMTHxQIU7fW4J4Lr4Agg8O5h7fI19XiL08Sh53zy8rfIyBM/xnpY1Prz/l
OZ2hub/jPHRwm619jHRaQO+rRNcXPMNIEBmW6BBdC6YRM97vNIK/3qk9sp4uhS17XB/yFxUxqcfh
HboLx8xFxLAz+1WLKtJMVam0J2/A+fH2kwnFSgNVzgbhmRsmiU8ee+mrtARGeAtKAd5Wchwpyd+3
JMMR0jP01sU9sGhF1DIZ0IhDKWxBNb+f+KCL0AdDvy+7Tn1dluvzzzrEQMYM3OEwTpT7yPa3ot7Q
B5WgcWEZv5fjLFa8okl7d5kJ7tbO4M4ueD1eJ3/EyMxZYFMwCZsnQIIgg86Z9/HyTwzfxAPjuybR
LobX3rCJbs+jpX1u16oAKXHm0AM6UvErnxtn8W+XoahaI/V11/b1dGz9OEaxUeUAxkfZ+H/pu0fd
gpUmKcMtlhl1sv9pATqT5LuKD61Biek7suJ4cI8bCNa+ZH5mL52SNoIjDXpKYcaHUFPSLKYReV7y
HgSG9yrd1Zz5oq3UbnU8kRKs+3A/SgTS/lkku4xB1ASe7CX0bMrDl5ogo3ifrprcsTzwi8Kn7wpU
vxslFOlgTwKAmYa76aEGxRfYVyrfTRUx9j8RZXBq2qd8kACZ50a9CNoQFn+5a5XyPO0d5oRMjJOM
nKF4yyEvWKbMXJR7m/yRN9tvR3XU4/tUFHlZ/H5WEHaGbvJ0BaFTDlWxg68ssir/eVnnPJY4OByE
nlEpFueJ9Mnjcj4Ft87oS0VmGpcbmkK2z+323xuvf0eKGg24tXoIbckjtSBowAqoQynOi2bOnaQJ
8K9agsDJ8d8D5Col9f1pWxLIUQSsDp135ZFBNby8vOFd/CCwtx1R8W+rKwflXLb3HmR1ezVVLkYH
DeOBaLZCIPf9vHCzND7Jufe5UU2giqrZ69yjNnkM/7pvNJX4jIpqYCVshB4m7DbUIV1RTmA7QdF0
haKDaRy5zVrLeySxOCH8NXuU4pQHAcxQKUwz/7fFPTiKimBuqyzfabN+wn+TqqU1VMJyiBxdqUT6
9MsxK8n6XlKR480Iv46sQsPNXGmmqrSZnZ6FqXD58PRCb7n5yIkbqMV3nmRYcVrWIDSNg225EWDt
GCGLjji5peB+ewC5HoneH/RGDt7YY3IKWPf6KlLMyRhD49zGPw+2606BeysajkHv6JY5Gr3mj5VR
1pigfG39wNOxjjeDH+77SVjDEWTyhmJ8X7q2e61c/zhqC3naI3cbLV+g5h4MH/lzryYHgb0ehIH+
sczQelM2b70KEVWc3mf/naAaMxEqyfOY0Pqeb6Jhyyi5e1j4brYuWJc74/efHZ+NCVC4AWT6nhyR
I+IuW16sJ3x+BHwBJMZ81FHr15ftuypdLmMHYgHnRy8M4DpHdt0lkMAtBCf9qk86y/Lg5yUSsMWO
qpfC8WklhvvIE6AGPxyrA+P0Cx3lcg9ybveFVIXCn1eXSza/2L+IfD3Q/MUerZXd6r3Yy5obhj4Q
Oe2j0kB9lqAGg3SLI0SmQyrM+PMTXOrULLtAR8Z9B4PfrAnvYxhDDpzdcReIJL1RiVWDtJqvrzZE
/SZ9sw+SSlocLUSNW3bn9a73QgPfYU2Z/lJwATys5LwhvOFI9SZDE6HLmJcMVuJDUUKufAy4GHBh
3QlXyB4lsMd+PsVVfTKSqprygziuxtMeu5vUEPeqNFbHYP914O8LjWHvMBi9MrRATFiIEjw+V6kN
1EYlWDhcV/DTa1w3rsmcIJTrZATTOp8b9QCNyfbk93nVT+dshZz9Z/IuGbrBrTne7IGF0rg+9fXp
SEiA3+fH71MaFPz/m9o5KI6R3ilNxBBbYIulXI+Bdq63EI99LCSXAmorZ+BPok+0g/ON2w/hoBQQ
zh+JlTTS8PW17ZWZYbk1TiV89J+zzyDwch5RZcGOn+2F7ZgNsiY1lD0ZhM5jr2t0+WfG5cGekK+Z
Fr88LZGSJng6r5BZmEay/NpYNySDBvPZo/suRrcBaihduyiNxoQnF2xJmlmvTRiSc8aGoFk+f5Wv
yEBaEDt0ShktfwNeH3thsM3rzyUF/Nx4/Sc5EGGrIYN+UwNb0Tr3ngRSHtkp6kFqeZ6UoQhnR8sN
oSQ4rPvqRFtGcQLD3nj6BkiOm0yoVyIkJHVP7uprkCbN+rBqNauW4Dmd3W3LxBwpsc5nTVdq0X6Q
/eDSYE7iLHHYtORr7k+v6NroGC3OpZCZb0xLvhY01MZj9MSa6NzDV5CyKfPJISthUAHJYIuxrdA9
vyH6bTRUe0RlKPqrNAuLJRyMcGNB38tSXmUytfZXdlQX/DDQOhs/nsbNsbCy9IM24g2/jnmh80DO
o+5pdzyhDWowqZY1pLD1rF7mxAp5NcnhkHt2YTt6k4pGHP+M++P26PjEF2mJ+GkW9Xxxb2D+Yhh6
kTbiOrr2Kbh8MF6g4/xi6zaAtCVKMjwqEuzg99FFgNss00ZiSFk65BJ//615gLvDsPGuxdh6fkWz
JZGJH5q63D2VfT8ZSWh6fDEa0AiD6c1IQZOyAl6JX05dU0M5XwtMUnF7wQusG4HddhjOPussonL0
nLs1S1fbXA538W5VlxDmgElL3vlOJM5QsrM1f41mmL4+As5a7QeVmN4Bix+ItXiZud8VMBS85Dop
Ns5p7FSeVVDc7+FkklrCtaB6UrfSsXvFHpUyBSG2EZIjs9tC3Xt38ieywpxwsuov3kRnkM1Lk1vD
j6tOTM2tG/DXiH6ZINcXkVR3eBpvqMWG53TW6KdCu8xyWKrR18zuKujE06MKIYqsv9f0tPhcps9S
FQ2V0YvUCisNEP4F7Q/YkbBp0pLRhqpHSVJoB3f/i4bURpyCiH1+F/uTROqnPcs5hibVZ9xPL3qY
YvuYge/eVKaAuXVIlohD95laTc97BWNMWqyVxIUAuRxR7o+XfpyA6R/D/ch5w7pV1/QkxNJG7ZP1
P+acmTVCxpKGcpbgQuThPoV1mBsjbqLKlEMtiP8Tw80kwr003DlooD6kSw3naZUMsY6YASsdr66n
ES3cJAdGFWYqF2k6GeqWhysVBOscxviKV4CgDQYXFhK3wQey9+MDU1YWV208jDqSCFrnW/hHOjwH
P5u6GwWofazX+sWlms0H6/guePLbORGGpDV9JD5GCjcbvIneoT3ldEMXKX/L+IL4rid4yVK1yF8y
ZG+SHyVmKURRIsA3wzdFqTuPknr5C8CDDXG/t3KwWvGfH4cLnw5gLM8U7m0nrtR3q+/JX/3ENdYE
HBaZEDYMMYy7kdHsfwaYt4p5CmAVXjPWlh1wplvBZObZaF4uSmiIBs/irSVdRKhnxjqiiB7LI3Bd
WwSG/21LJXEL58K5KBhNkC43rTANDAIy5RpDpAznK7A12D+0xa09dxqK33qw33SzpqRI85DkJm2B
cSIyCopgBs3KZyI2OeqKal74AJCMT825SL9TSghNH564V0rXMGupuOR14E4rN0qCIFbjt4PebebW
J93nx73DSdKB+qmaieKF6z0ARHxqLkrOnutCACouW/HNQZ9SaDwwZLq7fxbRHa8/n+t/ym8B9qb2
ZBVVpJ7LGuoTvf/P2qnrCL16nJw3Voig9b5HOgO+ipRx1oke8VjbiY86LnLVMQ1+Mw05nW9yMeCP
9dPzan/BAODf9+8HPwnQT1PGWh77/fWuRY2lj4bFajK3H+P8pwezw8zI3ddLJw8gGeqIpvCqRIa3
l5YzNiEkRNNe4J+cUyGbiut4genbeOWzAFMoX09W4Dn5AH71bE4YmKJTaXOe7mBLnebyfvz9ajlS
x8cjJjwNo4CBGwraLZGsvQAP8ZTTE3FYpnLTzb78cFRELupn+HFfc5uuQFsUDeDLNqHdOnNjTMpQ
c5o+MfVaC9nB+Jv8uaW/1lMED1WWsOJvkTWAA4PxpIQLSo/ycnRlgu2Cd4KqdMphsNNT/nJ6GArh
oQrOESEkx8yISPECRWDRRVWsLqztBR2ZDS9C2QUJAn0InlQNtWQuJ8Ot/CSKC4NRTch0qMlFY2Ig
MQnRdSCfLDu4twPPa3y+/hHyxewHb/9ufp+PYl9u65oX+JQJ6XPUEmVQHWA+hIfsD5aTWtXyjrW4
eVlzuQZCXlKTtNXzEK02+OUjCgTOZuxjl0BMrUSfkQW3DgDf4CxxKTZLhAIjvi+bpxZGt1e0JeZD
MbH15zBfC5KINBvVtSM9F22qKSdOF340s/ku+o1Au/On0wEkXrORCjq64/I9WkGlAmtzcxhbJHCW
sM5ZdxtpPY/rio9wCf9pPuZSf26eW7sIt87pO7bm7wbSgRnrb3tm5eebU8WoMp6XyjeP+JBG0Uz7
2ENZ19Qi/x/dppjYvqbROV9tLEbnDH18Cw5iOr+6qyp1BvdS6FCuaYi5vjENvFu9JrPPUKG8Nxn/
4R+vjy/fz+JR2HUk5ZXAHsnzFcLT7b+a4D4CCyHEG4T6HL7r3X2EvurfKxvvcLwb0Qsz/uZ4jpiu
txHfm781lXV4Smw57z4Ugds01enassSLeP98bMb5IV9m5xG+8KQYscA9Dmr9WVbTjFmHIDQGddoV
pJiY23hEj3BwsWkQGRn/CYmtB50iNkVuirCRFC8+XRZBxlqXD/pxjA1CJEdIKeWDlIct/oI90+7k
6yc1CCWSuxGYnvnqzVnWpeYZXdaUrehb+NvskPZP+kZ4Qs1rD4Fi7bkQWwpM+DR0fZp7QLUI71Bb
whdjxySBnq4G4MqB5V7ssiKuIDgJUSQqc6Ov8crUlPT3uZKG/zVhSWJ0ajeqSeLjNvI3b1KCRpq5
9K/WUJ1VQCszlFWKuq5y/AreY1jAK5pJNgczEouzPClQeyV/83y43sA8lAtEZZ95THpVKOOeSeFt
GuF5XoL8s1fLf/o13YCpmRIDIUH8lH2VhHg/n7oXPsam5QFJUAA+D2TCirkHQoJH89ogo3w5R/15
DcB6KOI8QS/ag2EvfzB4z2h6dK6VWMVwJSSatYuhwmRx/A8lHBir18F4iyRFqXppDg2s4B5Y/el9
dHaL3fYZeNxVFyNnD1Uc5OqNW1B1bbCOR1Egz085wRwtB8LyxAyrSnHDcZxcwOTHrhSTzsJ2KaHH
2ol06FC85gnUJJYN4Zu9X2heEMj6awSE4HSIn6RAMHZiQJeEy1VGcnK0c8h63+PP3Xu4CcEnL6ZO
IUCRvwi8Epl4ZNiwfsfQyCJ8ef6qEbFDG7vJlVA37N93HWGPMvEdHZrbL9EVMO/cJ3AGSmcE4qBX
n/uAEVMT1occTb6c+4XqjBfvtD0NfTiOFswiWv/a6dXm2Chh6D+FsslUypsC1kV4KNYrpZZsbtCE
3t+RuZTCBqaiq39JQ/Ro+pmfGXFw4jyrZR1SPHbunxHOTXhvzUv0Qs1crg6+7ra0x4NOVi2vE6TU
lJMxR9lVEqnBobk96PgV4ocBjVl+zbDxK74J4GKPGiI13p5EIzGeJuaZiaEjCPNMSvFivz4/QocU
+CkmbRJ4k580kRHgGSjXLj/4UrlOgxAqk5sL/aEI2bcbBHQ60+z4UDNaB+jBB1hI7V2xndSdOncR
4YvuOvByyqjTG7Mie2hpu3swM61+hnHqaQMaXkJuMw5yNsrDbWZWeqUlgw3/KSndTbAXWlCBI8r0
dmWNI+uNXldaVH/sX3Aj02T0HB5isC8ktpaRnjJetwmyAGQL5NQoOY8rUjsGVFLgZCTtPeidBp7M
CLEGlaKK21mi64AsiEvJy/XQwoyBK5nBhRTuVAGjedNE5RPNI3DpIGwvpSVJr+7UGIdvmUPnmHQq
lHkvCwfd4FK6aZviZXZ9qHAJfXVcuZpN/8PFr2HOvmX83BE4SJNpMdcVnkox3c3bxl1iArA4li6k
MZcbzP5FgsFN4ap9kptsDsvcfA/PauPVhowrvG+DjmI4eCpWyeFC9mJ6Dj3qdYVZ+QVpPHZUCYUJ
JhWBTKB6WuQF2rnir/lIq+PLZbQVmMCuImA9H13zjcbN1joOVwkVApeXrvVFdKW0WevjPyG+iH0M
jlBrThzcByONCTC6NTGQ8U0m7dPfhQ1jv04bZFl1Qu48MPyZLtp0Q3oEskpVigPlAPgjys6WnXPX
y7ALjzNrDZkx1+dPRVMzUaWCIDVAfI2mDezHbNfzCaixeAd4QHULbb5HFHTsPjGA29Ql6CnmicUv
nCsX+BCFc2IKWRSKZyK6qdGvdy0IuDDJaJQaVI20it9UCOL6OpR/3/UctO6l3jOuZmdKs714yHkz
vBMO5rW+OmSAEoltxM4lWoZU06w2Znm1q3trr20g9iy3y4UvAu42CcBDL4eB3U150serWc4q2eI+
MjzPyBor44KVCG0uUzAUfUBCD2pbOYiQzwyFV9SZhg6zI8u3DYoTQW04XEXB9wAciAZ/AMnsgi/q
rUg/e+SoHGol99H99vvWTf1KhKpNAiV47foYBKutv5eA14jVZQUQVWNnNsD73sUYfClzKG/ZNQZw
49BEtGRZdZ/1C9JE+AJuXFNzWAVDw0EHA3cQcLFuwT/w1iADuj/b9fDb5WVKOG42Ncf7q8SOB2PZ
700a6IC22vriwgpckZ2UT/gTINEIUUFwo8EmRMtvMJevOJCP9ryDs5QXW1NCt8n7HJGpNNXONthu
S4Yy8BJf3T2FVXKIHO0DrCWeqL0Vwj0JGTqAoTKQX9sGTrfmblZHJqIULxrBAQBCkoKnonSyFupv
LNyU6BkZ4fY/gyAP/9rvh60XxkN/Dw6+5YXqAuO3kgrA4v595OeJS06MFwISSIJmGTKTU7FVm1LC
0PphubrbkBKir8lrMFDZjICrjMtc3IrNeMGfh7laP2gH0aXRdsBFqp8QZHo/3vOY+sb1KBC/dAdC
s2hhiEEKysn7/jEypVQT0DJfYVPkEWuoA6Q/cYPvI2k/6whBAfEOQi1jgREO+ufi45kg1LNvij1z
D4rvtNKvnQVs9mkQ5SaKBZL1JiJkLul2lCerctyCLgHSTtoiHEKKMX6F5xoyvi8U2TWwsxIgysxA
HQknd19OfYwKmys9vDmO1IY76IuDrrr5E8m2nEZTGtexD6TItwAO79atbPqOKZEzIFlvHPD1ghLL
7u2VhZUXMjRBw+sG78ZzUiewUQyjeLM2NPOiTWP+RIho5Tyv5F8MyGF7JNn1ka03sNNw6zQuV1+B
4+/s53/DhVfr+yMs89hHvQRQ8DiZRyPMGgdbjsBIw4AUXqQ93MAtTvRDnNmYcaSMc/3hhzELMO6+
WDNUqcwtqHnCbjOPCQ5o5Qwht0/XESRqfx66fZJFIn+ky2FBNGkBI98uqo1fkHgagONO0GnqXSUp
ZSDD1oBjO5qC/tEdgaXJDT8b1INEgBGNTTDAdzXQAIQ9IpsllFjaOI7LPUnlaI0oBvViXZa3C9Sz
nFjcYP+6GXn9zsBwciasDUAOvBxuuJgeZG5hiQ5ZrZyjYWIkraUN4aONORMEaA52bAR1NrgmEtV1
sELd/XvHNmNsdK1p7qGFGDcKSeqJL0vpBeU6uWOqhnQ6uyyFdM2HRj0Ld0uyA24SkwzRdp6BQ1l5
Rlc5JeOqBzDVKlg89ib9FjICDL0Ajyt/FHOLhhrCjtXHtRAp/ulYZXxLKUfkhrKKl03gNiJu0fnx
fDOMheNmQy5ALWqjfp+JMNt+F+oodRX4puciteJtnMZHFRJoY+nwZG86TN7FYzMRplSjIJ2CfhnG
SpZGh4+5CA2yE7jgjAPxg0JOpL+asBxhzotIliQXnQMII/QE0htbjsDRBkfPwOiZkl4mIVofk08i
syIMVHMDg8cNSGwUDmA2Tw8al5pdggjff2Wo9mxRnfs+E0AUC+vuRBhigdpGJKv3cAHXzE68tfEC
pJUb7ZdvUiNqJvdtdIwKzgPfw2DBR6HZNtO/6AysaPGYZ7FDLp0+JfUJOc/oyLI3R8ERVafdFw9U
2Kh2xXmGXxnpmbi9KxOIEDlwKQdt1xXxDGqbl4ho2f/RfErlpIduQDdAkGz7BQ5elqGqR7ZLz9BY
uxO4oy+XNzXyhqyYSf+F5/6YRiqAhWdK8/4U2WwknNnB6w6CVcnTeyAp5vUvc2HL8XWdeZ3QcjV4
WEsLWt22oUUXJY+asm3x1QT33b2A0OoQImDiQcgO1iQeqZbvmHbcrYxVV6f+kwrANStWRzYueaiQ
NglpJwPlLSSRodpbRieckt8cPeT25ptHtzG5ikC4pxwhT7gbv/Ze8Jtsx0BH7cHADuuLVhaPxDej
5RCJnEHUvX3tmoFaXRUiNp09CVluNxQ7QFz3JjIzIfIRHzqiQro30rRAnfkSc8r2TiSpEKsgy3N3
+Pmo7cPU+mryhHvf3S+lpDof+K/DDUqZYo+cpEAFJe94tiCCySLm62tsKF1WjAaGbG9lgvEsWTQX
u2pQRdjelwVKAtwEok6NC8dUW3bUPTripOb0+BlkoFgPSc7wvfyNwrobSwqV1ErIMHHd/XJDOBMA
CNXbz1NRYmK4kA2AD7qJMIGtWTviXjHIotAy7v5aC1v5588JMwoWw1UBib+B2PtzK/lsyTJJGki8
E2PgF9xOi8AjjyPmJ/451tc4W07hHMd0d6NfBDQ+nbOCuu6yMELn1XOsNxwi43Z2CFzVpd4ZWDO8
oEwp3jNow8BjhmU1S3IAxMNO1xNb9e3hkmfJcX1kf01qHkihMxkCiaIKBDJf0MSx/l593PCi/Hck
+ceKIIK2eG8JS5BvarI0Iu+3lIlEq8bH7z68q00pS4jQwFfoiY1sM7/dRGM+a0K+dsIdgqaMQdrC
xJEalrvyfX9dlRYx/cDazinBNpt416l0ppqMLjyPqFZE5CD0P6fQh0G6sguIrs4FPHRpuuehK3q9
goAEgYMofBjI4J+l2iJqvCE82Q9ZopWExrYIrQeS8BxgU1CrCYTUUd/8l8BkRc7AHPTqmqasSwOZ
zdj5Kp3BihaBYwNx4cnSW8zFp62npTtY5nsFCtWrcWRiblfcya6QequSQtrRVZ2c5v/LOcXcqW7J
oiU/O0CGs1Ci5JtcNYCte+OEQ6MkOsE6GmHX/JmFp/8Ib45ZlKhdwtWcRELGjloC6WVaJ+UIRUQh
Z7tWNo3IBeJtSURs8f9BmZQ3mjFrVVcu02nawhi+gvbJo0gp6ycwsW3dKYIwu/IxMKkUDj7y9Ary
Q3dqgbERm11f3kiNgYLGZYRUJWShYDy2kMwexfF171998wIJg92FXO7/javHvOTLLnWDieOtGhRH
hQ/EMDqjVnbmSwdVqVBMLXecd7YKYuNUJLW8pnqaFLro/a8ZtD/dC4u8WpEbSqILCRn2ezjvvwyK
cff9IYSPQq9IkOTdLwoXwh8KEkZ557NNE9kEwOjKLt43S8n4X4x18ZFkVdvM+eV8ArAf7SxG87SP
eYjPZrqlFZ5P0B4LTdcPAHkM7R312i6bYyud+tX/2X3N5Q/9JU5mnEZa3pFqWI9wH3ZQDmP4y8wt
+lo1+9YVsSugRTU+dm2xtwJ2xlWI1sDHiIuXzc73VhF5pnC0sytjehF3YK4WSUxhpWFwHUcG2Msi
+9HkjPmqUxUyE6IuUxE2xf6NPXJAgBUzPE/ta39ufRzxN04TyDS14kJdNX7qBbn+F/Z5iqE6pg4c
9cuaend/Uoch1kAzstoKgqUJEUQWtXDviu+YO/wnrcXkxUvw6/Rej81F9eVk2QuKSf1pAQnuVNIL
HX3+WZawk7UKKY68dBRb8urImxe2jLrNr7E3pg+Fdeelz8pYulzUt0Zi2togKqHPTtlYVV4wY2DA
OIMgwO/mHuub4yg/jq45IxXTYJQTCHyGGV6EXgxKqV+iEDCa2C+Ht9SD66a1LmfSL0aubQg1yMQn
EtAoyvFlkZc97pHSRZ30EPnVgrqC5N9hIEYrXCUtlUWTx4MuPC3C2enUR646LHyGWCWSPIl4zHUZ
3kH1N/1FC2zhvTOQTAbrmhGz3huapT0F9eCXheFFfrKFe2DVw96mfJbWaqRRocEfFccImlUEcKR1
dwPboLvJqh2GMwE+YrFbqTnENgRGDWtnDaKy6BTCu1OL0bZSg8cA1Dl4Dx5zT1/Ru2YJ9f1pwQWL
LegJo5TAPRfJtYcA6xIC2TYSHaP3EiSccoeY/o8OeUYTdNGEeM2JCW3u1Vk3M5qcPq3GyY7h12Nq
prc7iSEzuIAKkzumR2Gfq/VZThONp4NM2dAbe5lhOvuPEyyfvFSP1CKywkJ5R+eZiBBI7P2qfEtD
3ex2aUd+z49GXlzeCMcdwYcAPndLn6fWQABWQvRtUhK369+gX71bmK2IkEs4Jd1ULwLg7dXnptDu
+BB5ObLJ5myL2cRR1Id737xCjlEYMTTPbsfmoak2VASvOBMBU70HQTWRLegiNo3h5Pj+6ApNK2wT
22V0bfXipspw0JgqDG2bLAQZ+o673VhVYvfb4NQlsmTcsBj/DEbgKII7X3LNO2XNJ2gOOFF2nkM7
9r42qDlg34I/AsKST3/bODIvilbGU61iAaSn+qurDb6eI9+aQ+fQ9U04IJvi/XnRA+uUslvL2Al5
+EOBv1HBib6ux2N4PhkRBdtWT+Nxp3yeXLbS6EZcdNFb8bznXPnOZjMc/Z3xKA48+onI+p3hWFiB
rfQw0m/cM9j5Jpi3Z+VhjYEIBrIrWTHCnNq/Ewp5FlEQD6HJ+H9okBTfwtiAJF1l4Jwy45j1hcqi
NMlu4MrX348Jz2YrMcab2wdqTkzuo90RxVDEBWxzq1ZV5f3QN9gCq3QyBlIviznUg6K/6bu8V29T
VjkvxgKaytgTbbw8bgMM2TS5AJcR2m4vOCo40Padm4yWDMpCMU8NhqQ1pmOJY0YpEFVGNuBgnesc
n9TRWTBWicPov7lq1MXF4ohlk+vpSIy90qSLlMPYIMfqfK30ZQfUC0iyYqru9V/2eNch2t4MnnuW
5vXr0f4C7K5HErErqOmOV4gMD0W3N4HxEbAhzOhhpreWsW9ET93tsENKV2imzpC7eQhY7bdgzGcm
cKtg3XktNt32zy79eChCMAa4uhIeKsaJH2wUL++adX2epAiO5Xs/mG0Yx3QV4SvH6AxkQTnEWVo1
XHhIIAj8UIbd8XPVGOHho9usUXuKaVgQIk7unR0j6ckNiIJYrcyrRsR/N1/xwccAOhZbS5z7hRV1
6SJKVLfPcEu4DX+9aMkIw2dsbvwhztkM+Yc8p3OVH1uAhtRZecFWQuTNAJTzFd4zvcmdrQwT6Wve
7HYDg2ICPxuUUbYiJrps/NL3z4Y2uTYfesVF8mzxkKm1gY6P+zuJV/XU3vunBy1b4WLMncY4yZYx
ckKQLA+qvGjsb9hdY+C2u5MktGJJ8reqsp9NPMUuNLnso9DPxvxnQoT2IAg8Eiooxnpw39o67NPU
/DNGfIy25WjnG+yKbdQhEk3KehJXVSh+h7r6HDbo2VEXjnWsN5dR9CR7OIT4iJCExOld6bzF3Paa
QxF5yH/mvl4Rqj+WUZRFnAWVhPwOFadjifS8P7pK7Ij5d5UV62feDJf3wPDRAMIJQOtMsm0msvFv
4NG6vo8vSNOiTjFvNsGdlL1fq0JAEK1LEuMSADz7YokwCjTaLD4U3fN0pN54/MoVcQon0LaCrwDR
aZXr0PSplo9D0KrQAc8otPHNQtzNRGbwKqvtloPJSAlEb48eQJbiQySM4flGNUsiZTGsxvHgGr4W
EK3aiWiBKETTAylKkqKOO0jPn8UBasxJSaUxW8U8oknoiZ0sCIE2z71QQUnFmyBVBrRkNyhogDK9
iAMjLSHmX8CEr72toKz8l5qgNRlJZtkwdTSK2L5dfSHGKoF4Syu70eO/3i/bdWIo5Ph/kAUH5447
jo4KguI0dZVS03naRM1iPQ1tr4fwCFh4bXQx1RcaeA0MKR+5XOOuWTeaQ/IKfrbmFWkGZwp3UFKi
Xezs+RvJvuX5bboghlLfjSmMA2f2qtGf+YrBk/0+XoHaAICGRzSvwgnfbw9UBGoHiGh2//g9E6hk
E+4Bz8a11VpOBkd++HJmwDE6DvjR0bncA/KBrr7ml+3XLIeUkmjuONVxxMj5VbcgT6c+NIbzgH7p
8Vw6d6BKmirJd+RlVr3Mt+K+TaRU0uOHVy6eaz2T4Vs1or0DG/nvpTgMvLrA7VOfHBJ8Sszmiao0
FavVATvCFB2O2eG8nu0CBjZ/DvKrGAdCLpKJMcYSsCRbu0clh5Rk3h7ucR1+wer3pBrVO6X4TL91
+NQhgL5dfaHTsJrxUNu+JbiObFWQj5hJZJDWDPsE4vMKRJReZIwaxzJjnOoGcNDe3zNS/vBPywki
NC9ga7+899QT5pyUYzO9y8kM50Ps+7MGzszpF+egXbD6GwilgawxqdB0+eazv2d95HvUpVtghsKV
2l8OW2paqxwho1/TMJYW80jsW/QczKdkU5wrxwMWPh4kjUR7pYAtiwClQ6aPR8vmB9MMAZuoQTYx
WMXY3BZZTe22p1X/xeyH/dSYGh0XvGJkRbbbBON/67l8jCmbKVrGYpmzObYjXIDcPMkTqoyCntmQ
jXlqAFwUgmt50fIukUdsqEJSoSiMpMWLqP7n36z0IMeEJNtJ+YnbvrW3FwAUXjmeRTtdQHNKCLxt
v6UEeNLM7S7ceQjS36XEYo23DVMlpGrTfjje5ecBsiPo3XgjqmXPvrYznaJANZX6AtWQXhwG5G1m
sJdjfNLMPaG5gIrKzkE+E4g21g8fgANRl9WcIphnh3b+E5bzT8WoeOB5oXc2uyS+aW5F0jEip/KX
VNEDRi9uVRTXUj9JtezX+n1AjBdWqt9cLzFsL+6CfwmSKnOt1A4f17yQyP4/VStY+dLil3eEUedQ
h5fOdz6RZDyThX+RV1+dRDEjEmpLfz1nI3x7MTX2H7PtvuHogEfoaXkGF4JQku8TIo6p8PT2mP0w
7yeVJKM0TznD8HKJNyquHqxWTX7eSKnw2ccp3j+gk6eaH7xn1pRuNSd3iLpbrcN5UdNMAdr2gYGm
IP2FdEYxED2iZQThVSBfJMKDw2D+mb1rnpC06inrufy7hlJ8KyMxaXxz1LFQ6utmIPhZvhEZ7vt8
Yo20mFkXIQs6xQlZqtjO8O2WPDI7AfmPMzsQo1uRk3WrWN+3Xv4A4H9quikvR20hSdc/DrnOv2I6
X0YfcA78DZw3bKpMN9lSxcnzXvDl6rqBJT5xo90kNhkXDIMblFthtZ6vWyU1w4g/gdp5Zxg+mJB1
gOPikvC837vw775Bm3A9RK8u6c1nusd6pdO8CyDZ1kYRomikY1cMiuT7jdUMxZTyitFilX/rlSjl
jwCFp3k0nS8p+yq93eSK8u32Aw/z2akPZL3HzQiIFY0PwEIjKR/CmS7jxi1S/l4/dzYHK1g6/hzJ
ncdtYjSZxJaLrhEh1gFoXLICwW8jnywZxau8Y91X4O3bKBDrezqv5cLp6Op1tOfEWN8Uys3UIk02
gsHtEpniyA6nkrH6FPtixhwsrSlsEo9KqCF7Wc+zQ80bvpA3dh6L1cctUq+LHNCf/UrJpJ+IsD2N
Qw7AfS0itHmU1xzLGmu8X34cRM3nIu1qs/0Z5bZ/X8jEYbov3c3wS7v+/Ni6MCcJuuAls9ugUZKT
goLivcc8hdSnZuI2Yc8Shz84dYTcLWO2rCjGUo1RkNgwboRSRLfvvagZ1BnrfoqhBKCQhtlrEqgV
hZNnODKt+AvtDZS/B4Xx7i64tGuJUGW/vMTxMlSzXFxMHtk+w7BtK2V93crx5lQmYjN2f9jD10Nc
5XJgC5zIt/QodIlbYwDNe+Axi9N58uTF9B5Yha98vxTEmCrc0JHw7mXUzH/dV9GQ+nfTgRucBhR1
AiJZ0TmxUUdd1aUGA1TEt5BoDiJeISTDlYZ6UCP9k9V7fuae7+nauWqvGqJxCaLCK01T8vmsT1/d
8IY07A4tAiweensiYTn9fn9ASJuzF27Qzecn1FQGafGvvAQioyZ/wircC/xg4Yx/kh9jKf/8z7bh
obhSIBR2z9SEyR5KLi71p9am+jUE8Fi+6Ag1hf5q7FGPFJy0fg3jHvvrFcut5mYA0U/xmRAeZr9G
0LqdzK4wyIkmM//r8zDGkbW6t8SGoqvCKkRqZDdCilESh+5gFeztEJX4KzOqJ5v+WAxbGYyiCNjR
rC5hoxQskAnJRDMHZBJwUAbtpcx8m16bsB8WvgZdKtyTTWg+3qqXZb7JGldWSdirj1FYIsZeRqLo
xayDFIkxjLoJrKMCcOXirHA1z7IY0tCNu2NwLc+VMIj8+CrmR5XlyugOX0NrwDavZ1YFPF4sFkKZ
zlcYaO91Zoyzl9idtOfninB8JgLRY60iyyZm7gBOzUWV4K78b1sJg7Wa/G/IzELlA+9eQ8cGuSTs
z7wiR7TryDGsIl/8UHXVV2+P9o5GgnByfSmVRltIGO3HeGVRp7X5OemHBkCvIHLobAoDBjBkIHkC
Cudd5jNPgi5UzX4GsdR4J0iA3gIbCkhZnaOLHm4rUS7h1zNcLQyEXJUQU/RMwlmGInK9lCYzMrbX
JSsHx0JqNTUJ4sL+jL2x/uLm4aQpI/oQDhRYACJX/e+lF+yLNSYRSxsuFWJRQcLAlkywlV+932Ij
GZqUYqiaM2vJgXnov/Pre9WrpmBk/FpnzMud07Pg617OajrAkknlrpD8Z3r4b3LcJeWw1tI5RTI1
kQNPjDcQ3ovaN5aAZ9R/CRFIOcuVah0iO4Aw8RsHj6gHElUaXXkzz2lTRNKOVWwhMG6G7ursBMOu
rPe3P79pqzflYZzZ+ynSjPQasR0LW6YAbryJRl99Y4eSTN3gLMtgdK6EHw6ZOh3i1SZ2F2frUFER
ZIUzXnrt+hxV7uIm4LjMcEcHpEyZ4ijdjkWS3Hw9dtxEQvgYNR62D8kgmsal7r5YM5SHUC8GLN4G
5GpNqU3nTKK8R+ejiw6ojIqlulaVWVwd6/gX+cqb50VtKwTbadkYpSIJN3xERZFIW1XRCJGOkOrQ
nFDqeEVO3u8KqwRtwCDQrgYf5q9iR5Mz0HpjFPmfQSf5+yS6wj9WVqvyiYFCF4qDhO0Xl64Yrg/m
1db0wYSuQS8XNfnrkNK5E1iAkAK0KyBf/ups1nM4uWQL4KQb5Czn/wYE1dQEW9oai1ssnkUIuwgj
GGHTQIbXE8OqqcDGxSOFy0mW0dU6RgXgH6dpT2KWu3lPZ8pYyTerUYwQRFNnOIUfAdLqPciXCJpH
l0xXDBKNSok4zaFj2hLMWGk+BiBYISxqP3lry9LvZAcp4DrHETNChgwKnkLPWPinxFtUekkskmgr
mDWlz5HhhzAfbb7oXuDcUK15aKRBmsfoxT5AbxnSU6n8t6F7HwrAAjsM4vsC6qzJYUCRiri7Xn0v
bdWHvRHF2D79ZZkp2irfXsdehGeah8ionp1re8rRwrbvO+gGqy9r0FMWRe8XNT2LjF9mtbNQNJn6
PbvQSWyl1QvzU1kVU0vhDU05ob7vYmi6DqHTFtcKzdRpC3OuRPi6Vr1Zuts5swD/c4LNBpk6neby
Z5HKK44GWionpstgoUfBhV78E4mQQJsKRUB/nobt1UM7yi0WM7GVWVPor2TjYwUlSv+AnxR5A1VV
EutF6y3FvVm3tTjpEIDnKw/nfrWxVETQdx6gSrfG8j3qYet19wB3YxpVMEOYpBsIzoIQLhm3dk1L
kzP6AfcsxYorDdeh659zyHBuLcvhWe94cF436Euxo9MnpMVYySDVDqijgFLsgq4nXi8miaX8TCaV
TBAEVBZph8uG8TpEGWl280jzD+tlBAlkbfi9ou0JKkcPGTDV5kmu9TSKDsdURsb/Bpb3U5Q/z/3m
PuEHHpbekJpB3JTaeCQBfnVFNTRHf77EuIOucn3K4VMKjiAjeEG4Ajb//78HZERb9+KKBWklX2zf
Nq7ofXW8AJ0oEBWWBz5xQqk+lCfmn+mQofZ+aSsk5/r8sqtbMnfbODwRb2kFCHlpYKVazykCUtzX
0aA2P+9WhybuDI8hTpApMoOvEHLz+9ucDANJzkcG084LM6z92XouhG+7bexurEHSUICfj1praOq/
0UQjcixwOqUL/GW81dKLDye/Fa/bL/lk1haElBTXnTBX7kX5e4BVBXre0/ypufnxfBX8HL+oMXE5
OiuIcAXN2uknM6WpgV8vqTXc7zS8wGKkxKVMeBH1pVSDbduDwCmmZuTyqwB+1TlOZ4muscQo+ClZ
sYFW/fknisRXzCwFO39KZtjWm1sf9EDsZsMApwvKOV7a4UpvE04JdoT8tgPZ84y8SR66zXLykrW5
daPbaVv9mefOH0dEGdd1wkUluOlvmS8dE9hYVMUw4Zj/2SCL+mkTBbS28X/m/Wdl4eM9b6s4OS4V
u5NhklphGnkYf8xPbz3SRGvx0IvVFn98KGz0j+CmU0YcYlqlmV5DsFOy0K2JKzzQ7S21FSwtClsV
MPYXl5GmMlg4I/PdxlefMN5NRvmL74Si/SF1W7e/6eaJw1WMSbS0gyH2VPP6M90rOayEpYmysjZl
aUwwu0A0yQqfAanZS+8dZATAwO6GkNfhyApsXvqMbtb+n1e6AbuNPmc2LGK7Hd+99fYGaYXkprCo
4UsMfSna7rnS7GLkYjPdMj4J+6wq0PH02Tbj53qjyJY6IiE1eGYYoKDnGOlpal2FLpVGhzG6PenT
IcfYGio6Fha+0fE/LLOb6ZS0jnxO3Mc49ZbcgIlEJWbMyimt6aWI0WIc6w72eh+SqXfeLcIFPQIz
iqbY8ve2TzVJvkrsWne6iz/y8B3hLLIu4cXhuyphf9wgxjdeF7oLuZv0DYJzrLxYtySoSl598JMw
zw0uWsQZGmMBGis573DX12FbkOkKA+RtEkD3CcQ/EPCVc76psEWFjiUh5pQ3aUQ6ytSkECgIOoKG
NxOPFhe0v9g3T9q+dWAlRSxAdz9QUAEAfp7v3GpyF+/DdLhiiocA4DjqjJRzq61g2vf2vIoFaEAK
MP4djBPhsI4G6wtbtqVKPEAfzytL2hy4MjoxQb7KKgHIoNliZILSzTNh2PQkflkE8SJbZajBVfvA
DzqfLU31sWnzswYleAM2X87S98R/hvGNCRnKJYrIznxJwIt22Ej/G5J+FpsnodFW4f04BF80xTP8
/OowAPBD964apo0MjgCFL4R2nPXrnhAZ4Mw+O3MYJMpamSLOjBTYfCGKOWTO/8K6PkaRYyz67jkB
CVSTFRzuMdBp+Ei8B62ysxZ3lrUAG3IpRaG+zpaNf6k22Qa7EeXNoWY8ScmdyhKF0+pgLTh+TsyZ
ppm1FDyFtp3sO8h5qLhslHUE4oX8ivoIxx/gChQcG/3RjUHt3qlpoZJg7XsBKvDUYfwthSblhHkF
/qFWchpzx1kS1i10pe+ZOQ3D+XbmRPE5ksXmXtGmD7g5DNJWLYvDt1Q5ztn+YMFOCd3/83UwPjsp
ENdwneocEiKfHhrZIcKqitepv1/c/9JwnSV4dsqC8PuejLvNyM8z2hB8gi5rqdK/fMxvIPHnzsQS
bjv3GGGqy3e+99JgoyjQUX9BMAdfgbQUovuQO8dTTQxgrw3kKKGirVNYpWF6qkqwTYATfpFNL0Kc
P7sBK1QFhXu62jFdHHbWEsSPMca+HXB0+ZZ9aHl09FBYj54cgr8Aud+f410ovUiyxp5QiBWtM/Rx
z+xLVF3nLcSD0I4sGTOfWGv6PTFHV544meja0pSXKQaN2dDkd+mau+RN1hB9SSy3pVX/QhKEWSw5
VfN6T2Qr0WINH6JK3KeIW9sXr3As1Gm7Vq0qO1iODcHweb3lg/STVDh3yvTmzcPXWvc0QGTHl5l3
3WaWmHXQhWINvwCMqRM8arBIuO/4OpWNfLY0uXGOn8G2/CLTVi/YfDO/h6Mjv/c4C4ap44xtkIh7
KfGlY+OzHtYpZekrPB32WoBie8dYXAxu4V9EZ6/Rm5VEa/THR7R5a7Z5w3pJ0yCN6K6Q7jns5+Yk
6haM2frdbuulA2mVR5yAQIdsd4vCwAQvD3uzAgfdqiFuQ3CImZ5P0NsW9rzEnwhuFi2d+QeFxQ7Y
TXCX4rdVBEoZ8qXrnD5Eh8iJ2p4uOSSOW5v85Yg911kkkCF26HzHDi/j992ZpEC56TNmQnUfeK61
EQz4MTz58fxRexzowtQ1BpzOLVud61IRSYzUlxPjlLUSZwatORvHkbqsZnjwFdM2CERtdwpR/Y8X
CKC7eiBSKeE0S6V2g7n3SOwQH5UzbFiDwvBPPFsvpJ9Y7CSP666qJpK3m3janItI5dQb142FyAB9
3+364TReogr6vgqr6keWsgbG/qV4Mobk45w4vuEGevk4wN2u+YUAkU16xLapwSQA9ub+Z1lx7yI5
Ztz26tQKsCB5T489c93TWKkkJFi+xk9qJwx4BtcYPH9UextPrOfD5j9NcYTVXj3OBHzNn2q7gRmX
EreDtpMC2S+OHwMUTjY13Jh+L6rA4YRmFUcFck6T6BAsTdkIgKR6gJCdYPHrMmIq/xLEc3GP9g0J
HQx8IU+le0aSsTQxwFF9ZugTLEfmrgjOLkmehAJqUeNoUZv7tmAy0VT1GHvZMk6o9EaMzD7iaeeM
QCdGzCj6JVk4tWyLB+xK8ZphXz3J1iMKIj9xDjP+AOvkXqN54HY3aASjMwy/Py9Pau0LXQrUTaUm
5/q46OISP7Fy9hgE9MvnB3TGDw5Rq3Jv6mUu1V5s1A0t0cdxYKBo3rpJzMQtKnd9SIkuy2+VNn6D
/RVpFCCizdB2vQ9VrkexrfPlN0dHhm7x5HRtr4st9YomTyw07gGmpS7z2AuLzZ3tyeFEtxHM0MXC
Fme1AzmLt/EbTS9hDgUAPmGp/IBX8WmwwZ99jqltyZrRUC2pLQvtv0XTq6NOyUk1uiuBSoXTBo4M
XRkSicTFXaut4SI10fAJjz7ynCsMSUQ6/MLN1zd27p6Wd4KbjEaP/2SwRPy0OCXMwSR3TkWqBJPv
kUhvmT0HFvJJujt960MZ/XTpab+sD34F/PQTrX3ENy10uguzHW75dqwEFY36zOVNh1OonSvm0leg
N1gmzriiRKWMT1nMjGokI8g7ZjIsqfiZX3q1ZmuS1Zd/7JajHzp17nS09quK+MRoOLyL8aFUQN91
CGE7GN1SXbHnRJ/zaz1WtgMMebZXDR83enyZdvX8UsM1Ppi2zm1woix/tq74DWBkZgl+evtchAbc
SUXrYEV8zWmLfV+wXK7suNMJXpewfilzzopiW/rRyqUbQaNo8QaPRQ8TnoSIWCHssKjuSo8qSJax
QeouIRu5NZpSzfYpWDkAaxgGpFZPxYUYZIyabfPek4wpf6k4IE5cQWMFc5c4gcm5arukqH/yhoU5
v8i+CP2guaISVVG7bpngkLJ5GVpAJrJIKkzycnGmqo+Qc9Og/Wgw7p77Sw2xnMh4B2AWaAckyHYI
HKkFe/etV2HmIluE2xfxSz9OeELcVh1WqCZsZgr7dgGQAohNpAlcDDQ8BSFf1zbdlkDpJNmSLDOQ
skL0EpEbQ9nPewu4FdNzDL4DnRPegq8uoiv9D4wjJ/JAAIJeZ6AekEpwLT/TSt6eN4evRVEdXjL/
Bw+wL3nCBR/6D+RuUkZbiw8OUOztz9+uJnqyYJpNOGzm1UhTk6GKbMY5R1H58SoF4kPlbYBlxtDP
KzftWJfADgsx05Syf/MKZJzmCBFDkvRJ1mF7T2bnYty3BFQ8ko3IqWVrFEgAkY3n78BX6lWO90Z+
jwWjaKDrZKFlhwvtcSzhikuyHqp18L3bE1oXzTELKqnmqXYvReBI3qZvp4dlFQxxNJS1WHqFlWzS
7NWeNVWxsYw6fubmhgHvYR9qxejihlO2wKEHEOHCw6caQQiEwki7aR7UhNfjLiPlVo0imThdW4iA
AlBpuhtAQ0eZg3KjRJuh51nIqxbztDZ/arXNUTPyx2dUV3AAMrB6EgUuhwOgrs1uYsq+6onsJbE7
89nUpMWGhyRD7MaU73j2o7Gwt4bOodBkKpXPmk9e9v33QoTb5QShfAoqxTllYHICeAej+jhOK5Kd
bg7ZGQMK+NEPyMhMH6jK6AsX3B556+etQa5xjh6QmbRfp1gXL6njHgF94dErShmDwMfi2qvk4W8G
uG7YThOu25nbZOQ60wcn9SFpWUnBU8+46PVJi10VkyVUEWYcsm1GBsS0ILX5E+sK/WZarvxHGFFk
wVKYV7upbnpEIAbSVEbAJ6sM30w51WgB2H6eIcS5q+xfqnJNEvRm+yRa5voyijZ6oNM34I6T19xN
BJE8ztgJcaUFm/1I3FR3/tFvChYBcueBhORr29OyLwb1Kg5J3rSm+F+9EPtv2vMyTLCah39WcBWO
Tau2qxAhTrZD8vyLkKbUyBu4VfNOS2aYEaq3QZbz5bovbbAaTeZ2sXCfcmZ2Rp/jdlnIVlUuFyoC
jle5gk49HmSh2sOpmEr4SvjwSx79ZEdwKV02v2CudwFU43HXIT+UuIiMV8u1cZvI5TmM5Qy01plG
75XEnk+6I9UndBRJA8sCnKlVHZQpdY1wfEyGYU4g3KAC72mzD+FEh+4PMkXBp5pVU9CV4hML+25P
zLonlAEYCL6q8BZc4MX1pgs3jrJ3ZiNptlP5j24fa77O7uib7+Iz/cinIhVuQYv7GNldmuM99Bx8
cobF6aGqCj/EEDJlCvX6hEIhs0PpVnXpx4a4F0bgHk4rFELO7M2R3UGlr4JnMJOIjwApY9184b2v
YUcfpWn4Ah85rZvhQKQ1O7/CmU3mwJ6evcAu0u19o/OcG3WTTmwvAvx5YhjgQooLTWhWFuSpT9iX
88IpCY02gckPhBldJrwgUGVamRz/kj3sn8/XdMTN5pv41inXSywpkGmsSD3dVJ8Vk011acgauZCK
poOJP/eKybjMdqTttcWCarcZzvxxtg/8jviny5MEl2TrkwXggBiOiK30/qZpIoFARsgdzNcosULG
94AW/ZuqaY2VcDFMbmxsHUAClQkJUaOWdWnaqA8ig5k0qJi5v+xnNNfiW+coSYea9cpRrOPF5RAd
usOsQxI0jpYLBNVG9/ZmCCSq2A/yrsmoHipJzqo03vLza/Oj0fpuTwqIJFkn3x2Vpw8mtVuBPfIH
Vj4yRjE/IqJXDdbHfiOhZtJpg7/CeXMX/U075ist5ped7do8VKRsrWqbW7TM2GiOgbd+lXTL0zTR
aEvfWJZ0Og+EDZLMxjGOF9Jjyb4eZm4BPJXD4HMxoPCcUbXaQwLlVOzS81zJFIsrdOU5kG+bpm/G
wymh+YoY0ikiASr2j31bntw7DCQvhu3dfTNVEP8a8j8C1xgk95yyhR4w124hCQOag80sODJ71vXJ
ZaoQC/4S1tImJjeaBTc2d49m4inJRWcIQ4h17sour4xCj09G+Yf+Pc5uYMOInD0RJhMNlgAp99Ce
H0RzMhp+ihHxCMSYbcqos85QgwYm4/UNtRZo607aqzZunknkjloooUCDStNCKrPwumB8yavQH2Ma
sGtwasozjdC+9z15JBCuFrYBmGs/LuAbTY2XNmtnpi9vXul8dzqHozgqEcXXCLNZ5zYbZ7zKfgbU
eFsc9fpRlVLTnLiZBvWt5MoTUtcBqkM9kFNe052NpJXgxA+tHUHJ8V4cf/5cl+HepztjwH0pXrLi
nj+8PsgwpnHybAfymvTBbuMCDkqqoj5+75BUgUxzyNKH6Y5hN9OKuqkArPmNL5yCKaZojTXCf9XS
w8zatfH89isXcwbXpeKNlK7g1YEYRpjW5XvTqgL10c1gOvkNSKWL9diOoqcqPqlUIZv9ocDaw6ny
a07qjR4OzJJrm2gs31jjCEOxLYz4t25ctIM+oLtG5HJKE8F+wrjz9lUPEq8P54Jtqd3fS1qm52D0
PXtsCUf9VDk4HFYD31XdQ4DlP3ohnoQWG/22QvgfDqvj6KzU/NMPcdHeombSlQ49d9+mJoEFshj7
/0/zyLlTiviBCzBPdY3bH5CLobv9yjB9s6xghSzvooHhLE9cdigCPOi9Mutys9pg3YayJPSEDpVw
VKKXLwTMEsDAi600OyQKL15/Mlhy8fqWToMCNA7DfStDYOFkix6i1uLUzIkwWveo+AQODRWo9PsO
FTnS9wtE0KvoiClW0Ilh9gamgwS7itRLm93F5q+KzUnAwmLp90c7SgVc38H8LBu2s50C01MBP8mE
RqvHH+NytJNpfeOhvErVtbrlkZfiY4lnEJv6+TvH6MwdmUMb1ScLNtAFoIZL2VwInEs/UaxQzmrT
NijsYHjqo9736W/qGM6co3tBOsss4bGgI0XPE6abmOSjxhTcdsI/oY+rpX49FU6/E+wZwOuRASs8
mSlwhXM4NAxbCubxI99X0Yut+D2CzB8ceXJmf7uIE8fW5PGVgEAFW9bV9b4wsxuLR5JN/af4Z6x0
QqQYRNHHD6mjn2Ag/sLs/s167/pUfzkD5MD8eqEH7+mYMgBsrhDZZlQai8qdrAoDTGRtz18lPmfZ
kohNqvR5Znk28NroIpAckAUh+j87cL9fATKDC1ieuNyYIazLfTbPvzevWguZv/4gea3vvCRCRZqB
HbpjHFbhrmJeedFRbjDnionuB/lv50R07Vpf5rm7037Umg80JJw6tPz7ylTkPY26Uvp44rN9AFC2
470+G6UwZJx/WFv11tM5uy1j6BbSx5s7yKZ9a34mZrmNEhMYwLzRzcv/EducWaQv1o/YEIO61twt
1jKlGNckLgLVqzMJjAfXA6L700ATaiVDdrExoNZ/N5fxxo4Buc1667DzXUa9RtMwrFbCr8fQFuog
4m3XWIcOj8fbqsFEvND6ewNGakte3HjBk9dFeJ9A/+AqtNygDGAWoA9MWlIJ2Yv36XuoPZFMi3qV
Gs0PxMeGOf/WgrE5Ha8LzEw+4RXoqK1pOesQweIgP/IpsEI5CMc4uUKd6YqKLFiIB2BwF2mTjmHW
/Cn90v6AxWuf084bfv99fYuMj1W2dgtvi3ydyS/xwRliMu9l+eQh3xDbDf9WXmMuR+H2z8fc+AA+
Ds1icTWBPkLiocNXbLHuLChvTX6S0clIcVqqZCCXZcOV9WXJQIfYFXfSLG0fzOdqpuWZyvr1bqN5
APZTsrS8WdBA6O2z6aaqFusgkLYaq34agUFzYOAjYCkaFUpZW9VvpROAkodUbgXKUXTChSmL8ZJp
0ZEtUEJhHtUw4D1t8Us0/b8EA/zpSgLNMk9K0KrktjJTOd5xruHEoG+10rmLmVj/yjqbyzl+EcwJ
SQMfjGQxkLpGPHUQMLoc/RnNmYuXtJYZm31C5zj5VdxGk/Tt/rIjEXJiDvSyURt+8+h5c8UBVQAh
Y4fn2HVWX3ay2ZctP/Dey9ZqRmtHvEccJVvkv42W4jE1IBqH3zFod1jQvze6SXSyh8sXtug44pMI
P8OCgKTkmLsxsxUZH7/MM5eaTvQo/xCeh5vFmaNVNBI+cRWvGXuWUOEp7cOXc799r2XKNSw+r2+t
/DoM9SyFMXsy04LzZRl9e+IDyv/wLntiMaYBClQCYOqPKn9ZH6V2jblrdp2SCWGots3JBcmyFBqQ
QTsOmZBaGpnPpu5hABuXyhuggIndl7drYbetQGBy+6UptfnH7LEtxxK6cYyRKW+sZt/PXZj06LR/
/9RkfRL6t9+peoILCd9d0RmdkN/e1g997RsRGy+gRjdcUEqiyO8jos7erzD09Yd7pv+U4+yqroy4
cc7vqgtX1Vv3fkAkZg6X6Y2AQqEHeTVowhYOwGLZQDlPe2uryIRxh+PI9kZq+HjUDGZFbigbX8Mr
ub6h7U6nfkZe1zOsIzX/A0vxv/GFp1qoMZNEiWascjWsiVdGizEMHXc5j1GTglSKAAVxcf6n0JhA
/2uEj1QMHAFeCYDpvC8mNpI3I0ECtG0qzjRw8XpAyWcHbq5d/Bzv56yzlSP3Q0WsM/Iu0jv46g8x
feSMMpaqnEm9zLlAHTjd7lQK5H5VlePSH1R4rG+u8S6vWsbGQ3sDucPkrEbHmDXjtg+7VuV3iQE1
FCs7QTAADs6w5VqqhDawh7eJKPImrD10ZTrECO9StExd6Ny1hyHZblg2iN1YAXZCOdufnQxrbi6y
+TvmlrtjxXu1LFtO09aEU4Pt7qdoDyiUxnKRxuHYttAIHZqZU6X9qxuxbhGFZRPQ6SnO1edICxaw
uMfOAfwpop692IU5faaTnka8YTBhEBptjvtKbB2rRgFZKkOMDWSDs+aDJovYy7MKEIMu7l36yRbo
1H3A5zPVWO+EEsdb+cDANI257FNGVuFNrFpxITzfb82FZUTXrUZZ5wjmAbzRyvrne1zS2amKbJzK
AdEhsg57qquxw2FjbLnrXqMouVb0RPUTH/5wWxi+/z16brlPToz52KbQlHGga/zs9xTbsKaB6bSw
s7E+N9kzg71rrWr1YR4YHRhdVu4QWFK8tyU3xYSfg7ck8Z4mdOQ6TAHVpKMoytduh1MHGNdDcN9i
eD2kqI4oWt00Pi8Uyt8P49vUd7n+ZVzl9IpiROiJ2SXEuyIXdZ/1fT4gTyUTRbyn9B4O/CRfaNZR
eHUSKdk0q9Qz1JcbJQUbYb7DnIF5+bdEbDAIjwqhz85NBrxfLFgBsNRjGRNi50c1WQFR0Fg04iGs
oo8PM2ofn8hP7l3xUQFi1ZjDdOOQx059MitZLrvTNIjxEfDs5Xel1eEAO7D4SsLe4GEwygzyW1QI
BvQYv9MtDuQyRdiAxRdrnAM7I7kNXOtX7wlWW3p4vE6RcCjEFvK8DmL4veTCl1i+jaP8ZzXG3hT4
tYfUnqJ43QybRTCj9dLAUO+FDj37S2AX+IChOTIHWGu17TxOPQl4QzxqKFDlZdgrhCoRiYB1YXsz
oXIsTwXkVLlvZ4pzqT9eGUKb3sa4Orn25mygWojiXj0qJVGuli0pHUMCyNshZJ01KHcXjMFtb9T7
nJsJynzK7UiV7HIfR6YZ6BmPmyqq/JkaQakdsrV+wZWfKFetH4+PwQc/JmuS2JMoaE6+BNzOr81J
0lebbcb2sS5mI4UrwZzAg0jeAUaGKuwlEWDujImnWXiqolYzh+tpTubrdPhruIE9vTMUqyG3i69t
tos3r7uSBd0705upprVdDzjWv8DKUPPesQvek179UdPee+pAGB9WPAFnLlP7KHOe+GYDwezFcnex
xx8nFA9zf4iPLsFtwDmPpWz2t5E2D5aVxaWVdMAFeSX1X1SLtDLdlffflFAwZ9bLs8L43YFnTkW2
nqpVtCxqNmqxLMhgsfLMAnDmjV9yj1x2TKI/33XXm9bgK46bKCTFaj7ILkNOR93RI5sKbD78aDiC
WjMv5LQXheaQTV/vIazc/vaNXpVtrKEL1Up1aztO3Uqg57rJz7Zr9gn2XDGg48kVLWm37qy9C+pZ
sFG3MVyKMaqAGI4J2MYEatxdbr/WG5D6U9h3Wbo3CrQgLmagLhF0/hGI56Vx6TMqGP0ZhxvCt6jS
lxquvq9fgZ3FbS3SafPrkcmYAeU39hJO4d9Sb9rBcNUKFdGzv3lzQjcPxV+/falvz10bwJzt8lPl
CRCS6UthtWFnnMgB54qv86V+zWw17eeorUkx/rQuKbuB93Ml1LPDBXvH4nXwIJkWxLp6Le0RObMv
tV16hoTLv/tgYk8oXWp5beIbQMZqE6ZFFnnUzvUsPef8kIrEcCnnkuGIDDWfIKI0hBcJdSkX62yu
Du50hVPaZOhKofIrnnAzkyJoGcXRyhbkqBawmazxX65RVVuPwsgk/Kwk5N6haJy4VxABmK1tWBnZ
Wt0sk8CnkPBiTgkkQqyej1c2Urs2VAz88x8tUVwDbuakcL/M42d+DLt34JhmPtTYSNRMwCv25bY7
PnZtNe1n83IXyFgGyOEAPOrNIjSwSsj8CNhmIaXtBmtG/bpkmymOhncEjHbtGTKi0MR2Xd16ba1H
YOi8CvrGwBSS2q1qNMNfyFrVVT2La0ES0pa2VNO454xgFQ3+DvSbZTqmT/uE/kLRsLC6YWlFk0Qs
t5BLZqxzBKGvgOa04fXZVc5hqqUDJPhVO3AUlSKjR6KG+N3of3UiDpwnAtQP8ayCcWXVIjAmxi8W
vunzFGUj9nUShMVLtzfa2+mHypYYYJWY951JPxDcoMXtq0yT4oFeBMhDwrh9FYTknASX9j7jR6L+
TLkqT98+7p60px5quGe0hrCdIf6iSoulafnQL0eyDycl4DHFGTjCPaEvRW5v5+3f5O/jL3RTlLo3
IPZizNeZaVQd6S235Af1M0Fa0pVv4YO0cHKuYKheYkZTuKRsHhV1cqloVb6VArFkI00S3FdMbMou
28nWWRSbkt0yZDS4S6RF4HULgXZFEKnK9buluPKx/erQaYXYPj8KFY3hN6mnq9UzP031s9juaSNa
VFgPLyjMh7VQYcRE3PMRK+v8mTw3soQyd/r0b7D+RzP2tMVa6MIO9LKUl0FAF4jMYcnZEvQaRSU4
e5ULBT54xaMRldYkIr8ED3K7vVc+vfc0krfozIiJgLysjq/A9/i/g0KcAqYJhKK6gPjM0QnYIF8u
CEmuH9w2gBWirO2IE4t9vrp7vui09SaJV41KbeK2JKMrCwtc+6EWh95xY6ZIb2x1J3fALZHI2jvu
85/IqDzLhSKbHiCD4PS1hnlnatQe8jpIs5MbEpyb+Xzjssww8bK3T7ChxgvYwUEOBDwOCPPZIKrY
0fqHrUQefyrtFxOjvOLRcFbJ/QTGCSlUBkQECwSZEZOopLSZENbJewHtNLe6avPWxu8R4pwp+0Yc
BQNkJxrtARHYibEiwN2PzpTfmAC9DKR2WHoP6Le2ehKHjShgxR7nMyfm2Oc+Qm6pr2+UvN280QBO
lJ+vdHNKQsW+n9ZWxZOLoELeme5ZrDkOh8sLDZ71wuP6JNfE1TUVqEZFgUqU0PHW/pIqz/J+AsLO
aqVgLrXCMPSBUPi7WQ0zAuV4lsdeUnE+2RKZp1iv0T1wI+dSeMhaY6dWrtUtKG52CTJzW0o9pCYA
C3VsDpyFmO99196zNb2gxFFCSI6j6ZtIhGct05QN8uXY7bbsbtdIVVVauL+Ri9wuv77RExziEEtQ
n+Vtunv/PX1dXSum8TYn5cdzVlZtTzIV5OMrPzk5/KB4lvOINnuMN4SRJlBeYZAxcWpYqIA+MN/o
aGMZuTh1eIvOycKLOCf++WxpXBNMlrVu8F72c0enxSb4inCoc8srw8JxlqtTt4EVle3es4FMXl7S
8cWcpr1KEDvysz7YB7H9wob06L5HOa5j3U1qbEetlNYIQ9/Kxb0TC50iKF7K4QmW6iLObi+IQowt
aP24jJeH7bS5VDhP2jvDv0RbSW4VHtrilIZn5I2IJk8Qu7qd2JCUuqkkWjcAoqA9tkvPZxxJDJde
YS1wgqP2rADBtj2DnLw6c3LhE1YABOfDhLIXVz9lokAOTIHUqAt1aV2Z+6l5H2QGiyqUxyWo5VrI
KSQCwUGFS3M8OjaeQq6Ylgwy3iKFU/E6AJk4eV5ogf2bbQ8sh3eLK4Xaxr3eA2tDH08S07DcDS9e
aSyGkuJfhvvmBCKtpY3Jx7sxUDNDm5UZ2PX2AoSRMm2m/caeTUTGGcYYIpqUSquE61/0oy4z+cZ9
E+XiM31v3sEWQ9ETwZoj/IE06FEKPJRTX9P84kXjCLbJXfTAhyYpBe4X0W+PC3TF6oayv0CG1o4n
luOIpRKV5ZzH18fO/INrXFgCr/fCev35i35AUtNjJvysAx+hsZ60CVj0/xT81luS/0VgD+rGxExu
c69iupaVMWeiEGB5vQKU9+RTBdAkv0dfFhswfkb+BIj+Amb7KnTOa1BkNGj0+sNzHayLgjDjuPGf
tRJY6PbemLPKg05Yw4hTM5GjFikFeYGwTpY5jLFm4L8FOz96lrVs4Evqh8E9nFEILR316yqr6HgD
P+s6qtoYr0X7exPpGLOd+14SSkNvUl8K5Abqzw4o3j3RgbsWwgp3GykSTEzeYmR8qYJCkRDb4a9V
K0Rp6tnAXex2Ukd5hMmvrDDq+PHKs2GteSYtYSLxTGARvbuG3BElV4QdoqK4gMq7G9otFsPq6jTH
B11vULWR1xGcKDVfgBYNGjupotPg680KcJVOw8rH18T5f1EMRi8sqQBRm9VUXadJemEnC5S+URvR
btZayekXmFi5jGgNvxvaGxf34OsIEbHg8gum5Tf1i/tEvqnFASOSprgIo562Lny6Y27E/9dWSz6W
Jr5c+Bz6kP2KopUPV9P3HT9nmS1Jq/vgwG5Lga+s+I/NO0wj6H9TIBlzcVTFu7jKg74LSO3OEKk9
FrLNdxUEVqSzML1Ks63H/ZJxIsqdsBgzFvvFbpUnLpLstfd93jwFm/v3aKlguzfnbt7jjIdl66Ve
mnToU5M5RL4bE8YlMFbGqb6qi580MoQ3Nw9r1JuE5Q7DkbRWTAa4gfmr9d/mbHdkGtdKxUX/aUAI
j4m1kqE9yKuAT1qYFQnhSGJjqiGBvofY0S94pOoPUF/tG4OJZc1ycfaptorup78b+Kuk3paCYqWN
EtfW+4Bq45BHpal8mvIb2KuDkeRnXiHpjDeHQ65+/ThpyNkBeMlRem2ulSKbpTfx4IAMvp9TmgGW
Z9eIVxdi0fb0wH7uLiIaRsufIFdT30QqQvhBjYIMJwFzUKGufbIfI1AI24nYKL3beeMw6wgy63ui
0+WdrtURF5esALyB2by4QQji+dZExAhphrYYOHMSVgegh6zm/v66VXWPrDUPjoVNil9EdiWl8//x
5uiQihA3yiYgcyp2EwSXisLKi/T5Zhz0qyuSB7k635aMsvNuIU+OolKW08RD0r/s8kLw8Rp3r4dz
dz71be+JxhJe1ANJZLsorbIVPNS92EpeApk5YcFS4MuY3aqaV0xkKhsHKm+5Pp7/CGez/0s6Bgui
62XJJiYOJ1IZquLZGMGDJf1eKwc4wTKjLlC8BkhucZn1nVUL19Oz6KYj8/MRyj/QBcDPrQ/6HFoq
VLXDgkadXme2xV9E6KLUtfWfBnLU24jZBd1HKM6QmjjcVKPeHiaFiMe1BByGwI1/FI//m89wxi0v
T+YVWRZp1jFVrJDqAOaoMC5Jp4khq6gaqO4p+KpkWpI/9oHxpBuDgqiI4PYD8N81KrAk6RKr+jAC
FueTqS7GgGfW/ntvzdHlTw28uz/6tQzo17mbxY3Skp2fNVIZjPFniqeskq5fyAeq4h06lalJHZLM
FzTjTlnWB0VpjwxS3sRKroYoMJkN984h86+QEcV0RwxS3BTsCVOa5wG9TMqrexap4G6Bm2nMbLk+
qLsG903T/4o/1RaVc8XyicHsHU2Qmy788hn8ctXlgw7JFuoYhY7PtxKqfuu922nW92KBuU88tn1p
KtGA5BEN9j7RSzdSyp0WQ+5kvbvfbps+oqtR1FLtWzG8XTu9LytCxojp2FUPRF+oNFGRDPPZqN4P
iceqMU4eBYz5DrF5TnQW59N5WC2DhvsKzzJODopH7mj6xp6lxftoQdvwcD3S8Hgo9gT8HtuoN99a
o6NWtQqkXlG6qUrJbTk1oRXGiGZmXOHiMSrc+4UV9+8WVWOtArjEuUD7xDjvDRXV0DkFE502GqOd
Vs33rB6mo/ibMwDd7qfbP2A1xRdGaVBK97yJv2bNBWv1oABWWZ014Q2Q49kqyPhNqY3hZla7LR35
hlYPjAT7I/tBxDQsLkQ0wrve90yKhf9uExbQJRgQIVBl5pzGokcY/oFhEmuTi7L0eaXHAG26ku4C
PE2HA7E70a7n+KH8zXgHGYa8ZHlvMdOKEnFzAW1Q1HnJjL6G0sxOB4ZrU/6XffNz2M4ub93IVTLw
WcUKInTVD4VoDyEOO3MevASc9QbnSrnFJyXHpXA190Qw1yfAuzJydZz1oWb0y99FtkecGRK+Wumm
TWOoYwZnNeZ+AVNIOahxwIYUz1ygN4JGpHHHO3mG04CGpQe3YyfDqO32GvDr100rMI+QIaD4KP7t
WkO30XQhm4Fl7jiWmooFtaMUwMjGdiux6N/Hhz3qKs+sL3ufDAvPmeNqGh6ufzsHI0R9KqZubODB
3R1Lf38nAvqYVOavJwAMeKj3pKTsN1y6AnjBLODOOuT9Z3LumTuVSTdjQitThjp7p/LW78BmOaQ3
xp7QMH93ijlwk96oUfzyy6b45X9iyEPXiuW6hzNyCHLD6uZ9FfcNVzEnzqfaruhMhrud43J0vPBD
keMNGD3OVawSC0ItLxq9iYLe5lCIePJYgDBy4WBpewvrFEZ9axCVhC3JOHe4VR9jiuUgP0NK7oqk
KSdt9ry9hzOsrrjxm5mw3FUzofpEcpMyrxdifuE5VTDuujNMoOdqkcGTUW2ds9m9E0cgsVLbFo7L
2k1w31HHzeYCzvTmKBN52+ynsHhASfNRWRRT7lQOznOFxD5RR3ZwYx5HU56zZSNyTN5fBpNMyuU1
3w/eSoJbcQCAUMoV93M1OHgmk/e2yLUxmhn7YJq7I9+h1zVk4Jll6CARCcIBwg478KUEIQtpB7Ya
eWNLUfOQK1zG0eBHMzGYIN9V33+jVCTR41tyVDGJFQ6BG/SbLeA/PvuoMZJVdlKLaAQAmrwwnYZx
m1zveNCGAPFRxRvIyW9rQY5ZUH8Me8xuTZWnX/sMTybUINlA2DHTOrjFy0g9+zJCRK9EweiTNGr6
FIymT82kXRJAORrCIQq24FsdhVM0Gn92KmA5LB6yc0/I+kaHaUtVF/owuEN7wFTXwccxb37U6jut
2eMMkdlznTnd3Qu4XV1wmLPNQ23n34gpS5Id74LNHyhUA86OSN59hfmsUmVX42iXCbGQD8JLck/O
jlKWyB+YqXDQcybK1GlFYSQtLnYa5gpo8UFzB/IvjTfyFiMq9++xbihsYgqd79vu1pWHA14VTAN6
hxNoIk4Eap92nB1lc+JRPZnRff4NvkjuOIeo11YZrcX3sjC+ngkqpTDX8LzCIdrasTFpByAsNMcZ
abQKppn8Pr2eMKDBDhEfW3D0mZEnpA8AyWxmSNlmH8Ag2Q8adBWf3AcGRfKmRbzHKZRbS+U3fZJf
n6rokYiG+heRBAu+cRdo9zxqE3HR8hkrOALaFxrtGHKes+SuWrpK5vUczPi+9yH7jT/P/camt3+p
smcBihKIJ/dOPqEE9F5u2yvLzeY1Wk2hUyft5+bUESSbZXGB87lg8V4TFE042tVmtONE0S4vh18o
1oQpfw8OkqBQ6TSrSL0nMkjN0SC+Ngt0QZRVoBade4ozcBV2rpNdfU26gQo7c/6k1870Wzt0RFfJ
a7TNYF8GQXyNW+HmYdJNm8e0a2Psshw4Q1+KpKbO+SknkIGHk9KJg1GLf4G88d2cyFDI/7E7hZnQ
630NWNv2D9f2Li+AWcg86FzgajNymx63/YDWS7k3rWXK2klHJ8ZWC9l1VY9VG1b5ZX/WXPL34+Yv
39XXjhSLHjKIn8S52Zgkbw0SWzGNi028CHP2hT06HeMjJVujjVx6QJb7c4fjJho7Nu1CguoPvEk7
0KtXwgphFR//a4g5KIXY2Otg7SlVuFLywIzGWMBTd2/mm7hxFk5BMCDBDRZ+hP7NM/UgSAGJvQNK
YaKUIMU3k1hbuHxceGcQipuQPW7pLN2Ytl43WsqCWm0HQJA8zuEYsY69B7ni+RR0bc1fOYou4ld3
5IB7A1N5lrTOc9K0AWs3F4u9A8pPgRV2QBUsNIGbR58gaw82VIa1nXRz9ZuSbUSUNhe5o/GC7LlS
+B3TWUJNzhjZpbHELw3un9m9Z4RBc4CXedL4ewh775jjC7rUXeNNniMQ15f7YEhnqd6c+F2TvXLd
26hBPE8R6JKTb7zwEKFZphPEeMFXTzusSuh/8j8OljI4ugWNod3wLFNXvMyTXSX2a+fUS/mU4TE3
uQXrxY4OOcxkTDK1fRpOYRYAHWFmhLezGiptSJvmjMxMWrlOSoNRhlkUfaU++0s+YUZ++ZDEzIU+
Vlbm02qF1Baf6qQDJuonK9jyQ2qDTsercCnzqzpihIlvUrmwwk3o1Zdzcpk1rVCMzkpJeDOezrmf
oDQDero8LvJspX4S2x8H1PEwCiqgUKONcv0YoDfIskQ0QlJbH7IdKZvSwYlugwSQ5RNTYLYXXKse
o6WJvt0b/lMPiIei7IKBbPwKZLzxnV/shjSqQPbNjWgW8Uzqqq3ak1rkvlFPWilCdk90VVKOb9bH
HxX5xhKzLjxgkVcvT5s+5FXHqTul/ZUDkhg3AGErDbvtJrinmEG+cwi/Eko1Q61ITc90jP9JYyd6
p5Y89TOq5Oy+cTzzEH5nvpHaGOYKJ7lx+udu3UaLTT4lDdnmQi0Q1ZIIHwKdW5SFkrUpKSouvPQx
itl2jBh8OYvPYZJDGYz48xOGHQBDNw05xSAGfmevEELLTxOmerrZqIJ4qMSdpwmxX6XKxFV4IU0i
6eE9qcOWgsdUHDURrmcncGldKYj2s6lPdp0U8GQX3Jvp43xHFqLFGjPneFujgPZwDwHZUGiqcOvf
wlP2fFB+rELrpmOBy9Ilx1W75ULg4Xemb9tPPsWXQiBJAyorJWyLR5se32ORr+lHpPyHzU8+9b5x
3zp9gLQ5T/yNlElEhbO4dC8S5bUhC7iOfgEV0pkoXNX4xln1WVVgGnlskbhe1ZqUA9z+dMKGaO+s
ozegcvEsydcj3EG66QuwwmhSqI8KnyLMrCR0dHA4rfLfHKU//jPPKPMtCf14UkmuTOxNE33rQwOt
dUxEciyHZMSLssD/UBPWPyJe2kDQZPv1J03ie0Zlo1JevaYwJlZJvI8PgzJ/qqG5dXUFFPHB+FAR
iXdCA32gVmJ5aAowUjd6riO7Z4ZzVYI8TE26Vd0xfBaGlE8KQqh4GmiUiYX8IewUpmukmj1C+Ppp
4qkVr/5cti9uEIUwmxLwN4umKmG6xiwqTCpDW0dzxt7Bn64fInz9avslK23jgO1XxKepTpUCTElK
KdEWTizZnkqm+CD+y7H90AEFLQPs/jA6umvap+wo4bLjBPvUwZv1cKp7nntOy4T5ffZwP3+gyIwW
abW/e+0WtqJA3WtREPm3wJK8j1ZeOat0Re1db/SaPQCRMxftGbZdlINVjH+Cg4VDt8CcYErNi/2v
BmJ4y8ZM/kbHeSuleob15fG52B8h7nzOeDXGRJHNvXdDef+STi4yLvnN2KT8jZi/mi1FijAaMk03
W5eIeQICTotCV3CJagKxORaILnAxWMz8NEhT/3Z2dGWu5LIFZEl4kvPJtXprU6xFTZ1g2iiE+t+y
kzRpTKqTIv3/6F1G4e2BcRXE/ddpZ/H6KZ42SNc5P8oK//vcur3GtdHIJYdQBqQG4xOoQXfyj7r7
V9yLFF1eH1fi/iJc4v5wRtd58MxQYqxTpTSDVplk6J6KEs9NdsLWQg6jGCTHdnFIAPF7mGVLEDhl
Hdm5sP0a6qnHaaDtNKUexI138qrqaJvOuJ+bh5/LM9pBn7QuJToyx1Yc/nhOTaVxMsAArY92kZxq
jGjl+9pC4fBJ0JQ6GO6vAm4jwvwx6Ay3Gdd9q4GGN14Kmfp4D21wWhI1uwzHn7Syf2MTLWZl8lni
w3skrTgEsPkHLuiqt4CIqW7kSh+nGU6sbFNrn47YXkgv/H0DMdjJFEP6925dpA1f9iY7jVPdKhkV
L5VZ8ZiTZVGMe4/8H6LpqQ4iVY6DdMNRCi36k9SX9YdA3+ARntmrUv6AfCPoEhNJ25TorNVFxYNQ
zE9JPYxqag4Cc0mAv/9UFKqfDGHTGhMVJwQZfudUcoMa3Enr2J6wDrc3doi0FpOF1XRkx77MuFdQ
27sAh2A2JYBu1NVHAl5AunqCykeojwqJy8KzuumEXsG9nQvpEoIHuEj+fQ7fW28CH/jg4yy7sOD7
g0U7oQJwwZAKAx6on4ijXiI3xEtDqy6iMyqf0OTn3qTo5Qg/rlfyrbmbJmVa9fYbuC48tCy5zV4w
GLpVD7eIrhdoNatwfr9byjtw699U3a/OMcA4BHpiLvfjpzMvjphzyDw/cfRBjnQlEsQELme7075N
j7NBkYgyyIwgEJ8yLlVvvEz/as6gcFA7SE9uIFLPgsRo075Rfb9Gow742mNRw5iKecgQpshzjJsH
/xLHRZW+wYgFizC5kS9T1/3cja0pfKQXRZTX2DCdkRpwC6RBU08Mg2fKNYRVeVjmm3g1exSk+fPa
o6P9j6kqrnqATT0OGhpIUFy7MIop4GDitHZF9ejtHxa+8kw28cjL7Kex1skk662w2NVJPmO5S7iw
GVw+VzqgQ1mx04auIEltm1db2R3TsM3G+Z8r32LRBlbkqMmkt5Ui6uEkrgacPSeTrUKOEk8VV/7j
/e33Laru8SrD5MRr1Tje5r699zHpYPNZPJA0fJ3QMtZ928/IkeMMJyORSpMLUzSo6G02xS71ocbI
UMn/lrdJcqo09jIksZIHGNFhlFRxGN1bbtdgw2NAhjLR7bpDMcL82KBFYGA1tAlkgr7o1/yY91Mz
q/QE22oxeJ8p5uGGsMO1YHZNdMm5zfyh2k0MLtmUoUp/4VxIWNUpbS7MVJiJ2f9ty0X3HdLyCKON
5LJOXt3VvLBN/XUG2JwdHUSujmH4LrNoXMoKh9ngeeNg1YC0UvoJpXviB8QZulGkiKCPpPuAQ1+p
TF363ebEUhqZip1lYxcgYwASm187ZKGxH65dgZlETq7D4RZv6EifnaKTh6CM7iferQO6niQ0wQZm
cXUC8q5ZnsV4BJpDVfjIbK1dKKrcfVb8NvCjqsW/sO9ejFbzfOzgsd49SKt+PpXqeOPz/ne1e4Nh
9HPW5LwfnlJThOGLpI3hPFtSQXt5fm9oub5gDQvSvcPSa4TZyavWuuqSbNYNnxZV/CqpTKUUpeIH
Ts+cTR3FgD/gaLpCMOVYqB6uSyYB2/P5IQgd6Rz4kyqu2kiPHjtCwuwQU4d8T8BV9rr3LzwTLMFK
xRaJSalO2wcGjCq6n2IBK8f77qQRbbuJpFlb8XdSD+5IUC51xspJ8EiazMX4zR5yp0erxjKtH+UZ
426iL8TAgzWUId1jkw8gGjQ269dfl8sKVHASKGy7w8uA2P6PVPP49qNACnEY197Hbas0I7sUCwL6
9rem7qOMvIAmz7Hs6yL1vZS9RqyeGVPcVirxHS7R66wxG8wkbOutOpQRJ1LWBmm0VvqFTvUt5eUg
Bw+euJeYQVlz+grSMT5k3jU165v1qn7vl0kIBA7mceqIdj1uod9LV8hhfRYKrhke/4hay0AYuvN7
9OHuLuaJGNnPNjmLObkjKannZdgE1k0GSmjdor+HV+hzMFxWYb2ZYh61Qt6DHL+b27DhCvIwlUjD
I3xR//GE3pJnJ5oARhS4IB2o+VGX++StEczRdz8OJzgsTRUc4xhAR6QD8uRomvi5AANxghs1kY3k
TPine0TSlVG4qyM2lk5SVenH2sZhaREDKfqPguPmCyUQhzGBFKUaNhL+Y2VaPkH+XFI4oizNboj1
9x3CfhvYEyO6zLIly4JbD6PRzx988jRipcFP2Rp9m5tpzN2bXnCrd419RFLZWAPwaewGzEqs7ec3
QG8hKCFg5fryjBaS3RnUA3VvP/zo0ToNBbhNgAFR5H8Q7Pfs3BzttYKlaikExUNPQNeSNRfnGeaf
6PGx2YB5LIBKUegQIA7CxLtd1Pz3zc9/AbbW/vniwKC3IsHclVunlrE8MYVaY4et6WXEphV3Wb6k
q2G87K7/kCycqURte6YHBByvJjW7gdAP6tJGwKbQGAhyBRp2I0HRCHfGcj7MG74DW6LhKvFc0h3v
cpLdrR0S4NHfQOaFAqyQ/r9+XU4WeXvQBtTivqgw3s14aQ/lsKjKisSxJliuWdutrJN2hW7eP3rB
36hI8/uFrljvdXJNTkfx4FFbc/eGHm5264OayGhU2ZblGws4VeGwUQncHI0YYyzu9nqzSR34gLvt
IBfJy+qe6oMg0zBEX/aqZZ4zlgNGH4KNKOLHoSFTIKtwZ02AY00THxzFEtNOT4wrWLR+Uv+stJxa
0UydqllolKrCvW1aMffsSPdpF4siND+jQImSspFEWBjqbdsZXboeASbARlQIhKX48vVDrYqyA6nH
CJP1SNn4W2fVZHQCjYWrHBYqJ5lFGofq4zV8z33jZbMMT/Dbfe4FZwNBZscXUaMacsQito5e2axL
mgGNLwRbQFewcGINscJLGQ/7A7pnqxjV/loV6KbdhtRrRuUmjFzXAAEEBR/4yOFbkeJg9lxH8vHA
6rLA+8saJH9tqfw9+Ux+Mei9F+FutrwRBaVUUBDz+myZQv7aWsMpo+h5FAytDpitKfNd3R0ftiLR
yzV77ggPbSMZ/GQ1DTKUpasMZjAKXaoNjzHXGb+q/S7vFj5O5cRz3icmljxZja0i4/odb1SNuybb
e1xFFDhwZzekpX6Gmx9JP/EK2exzLyEUWTrESdaGlNymhfqi11QPMhrOBY4nSeZvdfFJOBIo83GH
gUx6d5ApyMktIPhKlvA37Rosj71I9AyiNCDSze+uBvHpvHFzlLy8Qvl7vuB29/1ZxxiBbvFGWifC
Qp0MWdFA9/bTSb8yIY70hqLqePHLeuqcMKmgAttaQ4K8IngJmRHwsQ1FxDZfJhO9Y6CTkV+nWzhM
5R23V4K66PSbX0HjoZATJFAx2ndht165IL+FHqCiXpEcxp/Hg96kNucS+lPnjp4gvBgHhPej/c+o
QZRdEFvcaUoVS3q0Sl4btMiW72JSIv8GRSwhbE0t9U79L2wE+d9tYSC8qvmomsC4z98IqLz5QN8v
cfW8lj+b6aWFCxCRyEiouMXCk/LYkhjVVr7l+jO1vl+1oVFRc3SphbY9J+wJFTzi5aRPHN4lk5WU
bRYW2l4zr8J6sbNvFRR2KBgkV++Z5oAU6kOTHfEMAW57csN45W23U1f5JJiV5nRk5wSdOQTsEmHQ
xREgMvLq643JAUdZwjmiSz0yL+zrQRMcRV0JZhEYyKdM5sVcbZAJv016Jmjr8wda0bAD2L+MO3n3
obRcei2sw8zlwIiY7SQxQ7ylkDT4QEjzdhAiz4ujHnnXFZr3vv5gTlZJmnHRYCaoB4wL5JrI7N0x
VvKOLFiIlfjzsrzkdYDXpYmNHmWPaRK1EjTjv5GSLQYnwvwdX+nTXjD7zXPhTQj9vtugNcaG8M+U
icM1BhQx3GemY7oaxfxkGQWTCCyjIYcbWHaWFmfC3KYA9wWqQP00bIPOWp8xmGaYM8Heb1axLkbJ
vit9ag0LLo+M7nMG2InH+JPHPXcEbUzwfcY5FMHWitnxnmq9yTTDaZVi0LpVYaeqKZHO2aWRy1np
KMARSminjGB6XQ/JuzZSJVnPicCMXZIZvSayi5CB1NEDI5hDFB5OLy3FHEHj/eee7y6WSRWfORej
M0KywdKw3aJfxXkI/wACt/wAeknW8F4Poe2q5saNQI0OlWg9N6Kz2IqdOI7vkWkBYFYNHJvZNntf
foj0QMGzRoaO2hbfEjXTJ26QDaES7BZmdwWDZeufgMtBhi7fgn1lfIMTYncBEmlpRJyaM+/BAfba
hDF4HIcGCOjMwk25sr6bPMFOG049TSEE7N+3fvNenxCHfbGEAxXAMCVS9c8IEPxs3hMto8j+l6FU
GCppIMLVwTCra+7IdMbjEl7NVmjxPvkLwfa04XkNVJuXapdf1ok89RjJEib3faRMlMLUu60Dei1m
92I4zi0zSfEAV3ix24iVDLfCUrI+jux2egO9i//GfCZS2pB2D50XIyy9f0gGvNirDXKcT/rmcazp
5vInbXyqa8ibc4BycGwgp+Xyt23LCVpk9NGEZ8rn1onJaaCd6KZJymguF/I4uL9I35xve75/+Zj2
fY0Ug4hmp/AWKVJn97pRnHwiZuARCXX/sUwuhXGUlrfjjphxRfggAp3XodGxD5ZgcYVUa2mlIltw
BWeqtDJZQD456oLoaDp+GmE7qbAS4XmHyMki3EqWFdYqbGv+W8d9058W4E+W8drW/S9tCvxZ4Mrg
3LkA2IQtPegLx5G/GxnwY48DrHpUoaGRdf8xD0WaH7PLcpLlgA5b1tttRXj6tKTZXRkz+H9Bayv9
B+9bQo+x/BpTNR85K2GnM3cZ+39HfIEIozNyyVGhimZPUMWiAvxUIFe6HBAmv7mVvOfH8P9HT2eR
8wXBl7GjoLrlD2Kzf4/v7xxqTKKXVD3PW6VGN/Snh0o/aIZaMiazOSyavwy+Tiwmg+1p5WZt1qvu
LtiIp38vctwpj8vSotLze8vj6Leh8hSW8qBSqj9Af+yltRh774XJM2uEA8a5CR4+pX83rYBNM8Kk
IWKQBFeUf/0gyJk1Z1LDm9dAqZE0NuNEHMcmayMAq3V+NU4LFLOxiJJ+N6bW4YS37rZN9Q890oBa
UM8TlKy6hGuvUdUjWaKU7cqsVme4ZDAST9jwNcE1XJG17d992Wpu277ND3vdVdo21DqkW1jH5lH1
4/+oHnpBoDhEEwglTV85HFsZVizMvnUp10W55x/XPclpPVllT8ZNLrJ5Prihg13xgl0VDKC/yv/f
qLiBAZ61FJeAQbZOIW7TiS6KbID23IL8Rn46Lxw+wxM03K54k1OYpqxjZ8y+CWmro9teihwWqW25
aqUiJXbWjSmTFsf7ksI+TaqEuICCAZTpJrjLBj/ImB6sVVC4/it8g7A1VMUT0lhkY+AcmQilJpBS
UlFqUvLPzkYQzsdEH/9e2bGstkigz2sc/bg1ZjFozK3Jo88rvAuoh9ydHZiYxpidk1T0hX+nUOKI
LwSsaiUwQ+oGzwfQoTycKrRTIK5QwQh6KeZH81QV/lYg+G2zrECXZIMaMyKK4tqp55vbxRa+XCp2
jW5ImOehG4/AeNvOWVXaYhYo3r5OwJiiWqd+MdfnzD0pt1P6hmZZC4odByIReOVMPRn6BpMDbEwB
XA/2Z56TnV542zRD+QWsmMTwnvPXS5O5sSdd8HL2F/UBVRl8BWKRQqeR72alJBEQKGvAHaB+tE+n
EtVDWGkpbedinMFayoHlknuRaZDq4ho3vDO2w5LaNGSO4d34YSmrz6IWXw0sg0bidhYwrJbYAdrM
KBgvQNzeIozPQzcr74eqn1xG0yzq0+bpn+9SWLatjkEW1lFs8qvdTqwcGgUBBX2Ca/L6JyH2yR40
q0gUNMxUKYC7FXzr9M2+6TDyMOG5UMeNm5gRfgbp4Fz/NM0JClnEEpAatg3Cg/u0ZyvTh5QxwVoL
dzq/1M2Uq6uqtevFW3vJgSMPx0PRjNqNdu0hDOQQ+vIWcRs8wXiP9v60DlWkv15B4TI6O0V6uENk
xp5PD7nlifvoN3TOor7YfKGZyJBEbG/QleBMtkeeC4j4Xr0XOQwGhgj4INFqNt3ceziuQdurE2Sz
ltSC6Z9UVJlW8xYFO5VuYR014d/U3GY3sL2Cin3JA79NM8pM25jziO/vOBDEHzZGcx+U91O/TNLx
v8PXrIIuU2UHxtwTNOXT5DB0f5fVQrsfyjo3ExlvFK36oGPzZOzqQYusIXMYb7P7Gkv/0H462fOY
7urCBMEy4bDJS8jFtiLa279sPSAN6q+oPjBBc6Ket0ci7tnJ6UdgjrB8tg0JiLIXOk4QkHZUyjY4
LS7L99Kvojqil7P4hDUaNmsW2+8kevVg7oRDPBc2T7QR/zb4qqQoqNlCQr9ViFhZa5frioiutQVT
X+yj8CTrzDhu18L6NBElrHDEaqgN7DZQZ4/I0Pz+aXgXnfSDj61K3OVQ9SPMeVUP8LQGFIY3w/4H
DB4lv1mVFt13WaSTYe8DWVk/49+FJ/JbnJRMeKWjhD7bns9dukEFLHa8oJgRphxC7nG3Y843wvel
jPI237VGYPwuTVlOZDTPf5DdTUBNdhnQhDMq6kGFheN+qDKo4AaAz3WOf6S4l/5nnyWhzR9Jl+ti
ABeJMOirCUCC2IcBiSTm7vVVjiYLbrU5aUUZ6hqxbNbcqoLFkIfj7SerdnaEn82Kjz7BwJUop/In
z7J2dlcU4McDXC42zLlSbn9iui68hnmnTXMgAM2Jm6TWLBbyEJKV/kUQXCgshlMQowTEEhKoULIr
wJMa+t/L2rpmIBPJP7te86TvwI74iamussjJ7VAPtNHL7o+DnqWr876oed8nz6CcC2LlDSCI9SD+
WNzOpHyqwXej73scyuyKqAmFvmVVW4kcs8fg7qOGxSAqpRbUWzUKbgRJDT2H2LE4na0s7RxdCxmL
fUvFK+vopiadVaAJJ/Irsu/W+ZUgBgkFiwgOlaDn5WaMYD880mbsufdf3ay5y1JLhwa7GSY8jogQ
4Gn8K/WyDPl8DnQ90NH26rT/MZbTRZs3ccgYAcT79RyNxTr6gQXGNjK50InL6yuIwfQTEtXiQhuf
XX1DLg20m1YfAaBYivE1q73yXX1Sv56nc+d14gW6N8DO1dS2iMswfHhIi/ytr9KIWhZzb2E/7ZXW
D7pEuTRGOa3NFdyAeqei2Gq611gaoqviznG4XVAp2+6nlcJSJbhnOfakzoozmwQSU3Ky51jHSvpA
rwumCi/vjH2mw1UzuXApcC9fAVWUJldEUAcNaeTBbwQXY5Ka5FHSd7/3xLUgqr4V9IZS5UH/7G/W
tOZWQ+TbkrVIog6138WoicJkyGWvoUWSnkVctnxzdjIqEsXtVydaWJbEoKQlqmHsRNaExsBeSynz
1/m4mlG4TOk/7yEk78oWoNaQviZCwEUHcTgdcEsqLcFSd6/qUBeX6nhteQv9cHmkvkkC+UHLPCW9
Gm3cWAyROBaYIQYl7fZehvFNkjD0FeFYr78zFFPk/m7DRGTsPWtvv8SVe9cOuKTWpMctPrn4EugH
QmoAWil7qH7WL5K7oV3Fo1FQtukrtywqUgpmu8500Lz9Bz6Nhi5U1FuvuiOgx3v8TX9YmTdTK8zm
w/5n9No9dGlN6vd8o/fZrlYd+Fn/x7vE+dwEkIrrpWW1lu/SdmsRWkoQE2TNrwXLEw/ejusyr2HJ
lpTtNABzXTzZvC+U2177VIa6z1acWZsyYbiuinXjwW98UimP+gIxUPJ+Kcm8BX1fpbkOeeZA773X
DZ9RssJ1ykc1+cD0XbVXWEd9BZqysm8NucFWPRVi3Yp3qGZC6DjLfLLddCJpg2aSHWz86gtnG/0q
3z+yGXxmQYtmttcZ7mHM/ebMfyLPYKoXvDU5bAI2K528MeHZ0sAcehn+MERLe32O62GHM7vf0Mdb
9X2GeH2sYE4Ma/wIyKaK/tHPdeuRI0nhB0xm9gjwmU95OZzNQiMVl7b8DhW/4WREAzCcLZFpi1BK
VFTnhtd9OlyrL+TTWPoUY5ZHPwkrEbjtLyUGwNc5KoCOVJ/t9R+GeqKnlHzvAT0XLVqySdKFYQ2R
2emvDMaiGxIm/ky1rYwoW86X56YDUuhQUzGBydolDkCDg6l6B53U0Sh44EuZjyG00mfWHR083kiG
r2qGgVtJued3UjjkCGaRhGJ+eDDvjMWc6UUgXlOkCx3ldSjTdsWu4XVdEhJt0Wsaqa3ubV2NKM+I
rrHx1S2M3dbWs3UvesFtyrSdYX0qrSwK047y3jM26TR45MI1pP+dNj7JnKMB9F43LfHvj1J8K0+H
W1tv2g9DG4IOjK4nLH2h+Um4W6/6sie/rhbJvghrActJE2IJ1T4KMCEQb/Lfw0obth6sYUped5gz
apbmZzbjXxhqqEYjwRA5Vd7IPLoo67075550dqID3HfuYYfWRWMqrPU3SyQM/exu2JhFDth+vjhI
VQ1HbriBD5EQlwwpm+kJRLUAO4NEtmAvA/19zeDNojvQ588rRiE77HGwV82d9QwzJyb22y6JvfdM
Ico//JDdIZCj9JUV7cUroYQrrtp0gGU0oH/ITKmwky2sxRD+UaJ1YTPGYIH4dc4QVWzbWxNvT5Ek
lLx2eiwByBXxP83FaF+Y0/Y07h+wbMMeRP/RUTSxVD3OiyxI0/QINpr8b1/EVwBiRnqprUpSLiWX
/8QEFRWibNpAmSx1QmUCZcHQS5WQRtVv2RPe5C/o8ovTAZFMIVbnKP/7sXRWLgKZVlpEWchpaGSe
wYG/Ob1VPe5sCBU4AmcRh3KKDIbT3zeV7DY2OdPtynGESekgCt8SVWx9oqE7TQuhhp6ghwMfU6iy
LMOv/UhWl55xEobHAnqoKUE8qGs4RZZT2MzRb7COO9mDHC55KPWqCgSmKu6qfX9HuAFs7ZFR/CLM
btTvgDwS0YsoD6yq3bzi5q8r51Ml3T6tDsr8Sk2G8iLMHOTUR9Ad+JHh86cBUtMmyxYy97d/KRhl
V5VpuO260BqlTO6e1OrzWf/KEXYYU+gPaNxPcBHFKYOwQPTy1lYT1UHQ8uh7cZnNJCT6bjOoOWas
m4gnrdM0GyZcgTXKpXjZsfwbrlZA4HfA4875WOAgFxi2fs+/r30y2Ay0ZdZWF3vomUBWFqs2RbuK
bGyVvK+r5P5NQyaq4uuZA8C+yjburQ/5MFvGonEI+zCdVMrXmgM21FhH61TwHvFMg1IFBfaccbGP
OgPYtU/JD8VxaGgHpz8Ki9ijgLdUYY6sXxw2CCeXDlgg8Xzkg+C499R0EAfI/+qgzritBaoTsfNz
STNvbMLbL09yARWaNDP7pyyzE8Fh++zDRgz66YDNeWjXTmvE6ARIra8jv7e9CTcDt9u1J/foM+zw
vrXROt8b/1wmliRzJuRkiLCMVA8Q7BM+bLOBJtBdhuvnr9sjtgrCZHWcQWFMHXMRjoEHrPuRHV1M
shSGY2BA/bNPkq/5i9nJ7bRrftLKHCNAcoREyuh6br+fa2X3yWifqRSqu97aIOSgrsTZysU5XFhe
OrIGpcoRD5zTSTotIfxCGnA6cUC8vnhwFpSa27+Jl9/9LqpZHHkncMP90soLiphqh4+l/j2hSBWN
7631LWDeGhshOc1k/Y9PQpJCaT57TZzBwH0qOfC4b51YBOZiLr/2xZf2K2urQn1t0wtXbpF41ndU
R/lGuw9J3NQTsMCeyvaal7BaKj9FNu6RF86tHXWStYLXA3UsY9cqeoPh/MZMBKIIY0j6B7wuHDr1
3z6t+KzQ5pFTQw5Z/8mhrL4Ll2rFx1F472q8EQmRWlQfLGK7wP10mmFaUhWafq75k7hjuiQO05wA
/mRTntmOi1qX5k1B4DC8EwZkCrUWoLtUNBKhN//fDhz9HVzv7D9dOyamCBjp0FPk2FXY6MDYtK31
Ry4m6VRMXX+u+CP4n3QoOIpoApitzO1YdToaQ/cm2vcGj4lKCtzqYJH49y8okpURrt068/kfC+N/
ZjFPnykUsG2Pm1EmNleRWjK4hGCNFo3c5TJhEKDGkrmBcolR7Yu1qzJuPBeYZrAgzS7pYG9MRyJm
vhp8+kUyCvTWCDrIavA97jw49ueDTAFFTVwadWDSjWbde0tHtgy4rGSzaENvYrjcHEAFO9I/13Pn
gd0mwmedlAuxMxLfThYlUXCtBSAKsNgvS7l5s6T6NIjoUklG4qxKMrrbAFE+jizEKOqWjJh9Wu6Y
H+UJHk6si4TRMbDPeRHTvywfFc5gYwb/g9nF4+5oS1x4tNrzEx5OX6YN0BVwSh1GJrB5ol9eVj9N
QzYKwt3NrzukqrIKUN3/yvtcYVOxEAivrTDdkAFCM1WMojlHq3IFZW5O7K4E2p4D7hEdjemhn9Ot
AILX+YABDVXahk8YMEzkOcCcbP7oSWLUfjSOg13CgyMEqFbqNrBASwiVCSa54AuiYGwnPeHiiqBx
tXXM1oKgRZ4I2pO3IRjp/iwKo7sXiKEYLaBdtN0Bk+CYbDmHt/VVTgz5jTDqeOW0JeLBPoUKhe3P
wncDEhXltB10Y5L0WbDIxf+nR9EGAWQ/Lr0WGjGVjvzb4mDoWqatSiGLbe/D9whi/S0pCvqQWcpv
MXJ5qb/qlOwPpNPwpyPLzWd6yHjdKrXdffqxQilU1jRqiLR06jj16ZbvSpCLqcg+xam8V/yViGxS
4TwYG2HeNlYABOLdkrqiSLugD9779kxgT5d+OwN63D37SjHWwE05Earw/OLJ0P9A+FRM6bVdoFK+
ujo96HMxkM1tgAvZZTEtlz7W+yitp9CM/T5yklvic3c7BiNAxUEwJv3OjgWYoB/RXBwt+fW+rgBS
UWyKxV9JJmiDiuvVCdNGhdaY8lqaAEPU/sKiyRynsZHFCYo7fBaLIxXkPIzf9A2TaEM/alANTAZe
H16gZaZUuJXEhRq0/5rSnlzNlX8RwJ848wccalEr9ZP82L5v+QgQUQyW+mtbyGbmelH4TTG7fhSC
GVF2xUUmjWAgdIoi2W2P74iTKVKWR2c6Etr5jHLI8HTsL38fdTg59EHnjCrEjgME/Rcu+GwF4Md1
B4HQc6YUPXK6l/04RW5lO7LgsyHIIZ7uTM+XlBXNlbJ62ZL8k1aVOcQZYEHR/7qgR9znl9IaJuaH
/KgAq1dKxn5PQU7UisShyY27RgsfAJuYkieHCZqaU4nCnhQRuE70GzTOnv/aOZd+4XuGbKAnVeRr
Ix6U5FD/PsgT9ybWz3tPxlfE0bbp4bWSNibd0d2cURqDBtsmljptV4rVgsB6Z5CH+mMJoTVulDg9
LgCYxacZPzZAF4MsMcQZuZdzzeDS2O4BllxveSLpqUq4wkKdTXQgDHNZabGI1UaLulvHRl7P4l6d
b0lI3e2xLjkb0x5zVVBc/arc2Bwotg1fNbecgLwipw/s0zLfQwnwtBdiJj/t64OBNtEzdxHciIeo
COFlDjSL8iPl+b1AElWJAnokNkKIYY9IDqS1pMamtBjVEwH08C8FvGsSrSkwutZyUSja8SebX3Yd
TOSSHZPHFaRWIE51JMB49/kv+rwPfVX1D1dT0tTm636SIjT/62qBMBRc30+SkQWlxRBfaEImVr/A
PcyLiwTDkEn0rtwVsJRdI5YDVbbxWXPeUWCY+mZABG5aFIpRQvRXjc+gGI0jmnuSa29R07K1g2YT
/o6+hnlGRQK7BukqC9eXdDP49ZzgSOk3vlWH6tTyleygezvAtsfS2uazr0L+uN367EBYQWYmwqaT
wZcRY4qAnS7KFjnE1yMiVNgOwwAg9EmhdBLnwv+jGOtMp4vlks0/I7aui2p8c0tlpsYuIH9mkqbV
uvnFTXbuytK9zkkxGhDU+K/35IsLOO1MdpY82xYH1Zz8nuIgIyfRTf9DpGKY3nlDovrnRbsKLUhV
w+tnrZDrmY2qM3Z6zeIIPvYSGTzC5LYDF1bDjQos2b2j4cpriNRQMP9wgQx5Ie67ITlp68d6Ei8O
3kntmZazFCco0+Qd/1RxDYAtHW8SEmlB+jmjvpAdoBX4Z3P0+tfcN8JZVFJxmjD7Xk0aqQeBKGV5
P1Jo/bayppk6Qg3+fQAnkDwSbnl4NT5W3BzJLS6sfGfZmwtNoLQZ4PsKmXWAfMN2VRP4618bL0s4
lDfnUKw2bB/0vgKlOBA/1JDFfBn5Sl4jTU/V98mi5JjLWDLQUrS89PagxzHX8pKJSKr8VCnvxt9H
doPDCEmFEiB88znlT0iPiPwgBMU+bAm+01moKnWxvxX4bfdgdeHpmMhGwGQyUhUrgNdnJBVLJjTj
9cTYQyyWtLeXSfMzJPLl6OR2ZwPmmDk6IPPGali2x38MnJ1Z6+JUWxy5xNBGV9AySqIv1NM5PcKu
27v4fHpvPci1jYK382N3H9CFTUnJAK5TqrfUij3heIyxoLFYqnNkjuFU3E9GbK/a/W1O2AR3Xh8w
zyF3y9cDxMvanCXhpkbK8gbe9SGYyto9S8oEj7mtBoGGdZKHnN9HXsuxiFM66vbwr6sJn5QZVn83
cGt5n4fXcQZHUbfq5cc37Dq5ZIqplGArgqT3LEs01o7yajWhSY7yMGzKYVQRnw7HM3sRivrfQbP5
C5WPN4g08KmveExRFMRr0lpmUSJt2kUqpVT1h3dAVDwH+ghgvoRYbp5QOhogR/Q0T9UGM6V+fsxI
9fJM5GSl/KtK2gGVr3M20/M0dQrs/3cJKR5g2bDUHQBvTAE8SP/snU7rOC4N/kGP4zel9S8vApq9
art8S5pVSnUR28dotS/EeoOwxfweaJt5N2kSFOoicKaRpw9fE/lhUqCLLhWimEVST5U1DQJn8ila
wS6e6j1/x/CXLXNiTtiucwRIUpLXHHb9TxOcG/nLK5Ljp/feDdlZ+QBdR/U8u7/1ssLEQLZljfBZ
phPM3iUjSVqmo80k9Tgu6iNCkiFKLUvX9A/N0380O8J/kzczzEO7eq/0Z7hi47gwkbmqD3gqfIRj
HAZ+17yUiHEXarMqtEn3O1EEe0hmp7h58KRuCszVtWPDyUjMbW0bW4IfAjBUwJM59JbgsUY3TSdC
XK/eVMGnJlmdWoSWI0T4oxgGgq2upqLxPAj9mKSsx5P83/3ddpvTsWsMwCx5t1WPP/PfUuXHcxkS
5hYwL+UnPF8QOwn1K+dLEEoDCzG3+9Q1eCKvhyJySfMANu4+Aorl3cQwf5BThywND+wFfYhJR78+
vRSc55yNsVqffYWheL5OQ1FE1OJLkfTEUaHCcHDNNT7FMsyIv65J0NMITbVBRk6k0MVh4nV6NFrj
uctvyA3k6GwwpIRJGrrB5DSyYU33XYkLnsQroLRTCHnQvvxMy4i2jb3pPjdNL7dXCRDJ8RcnDlZL
Qt2vhUG6/UtTW9UnGR08/XuPXdQWtSQi3JSvX7ysAj7ee6Yejc7WrL1YcclChGdmoU3Y08jpqbQZ
44X9Rp1KR/rxMvstmP9Ov1+Pve4I4dIIaunlw58wE70ojake4CsirHXI4C5BkZW2iIayLg7enuXy
+Q0TMdOK4DwxVtTHDkV2xZjC/TmGl825AFys7ABqFy6+F1Zz4qnIcGWhu/Ft57qG9d7zqTyKx6fx
IKLDC/cDa2WJkqqOlPtWi3WGGYE7Pb4gBTN2NBxIbxREh8owOPtimwI0/AwCOIPj64KNaatg61Ya
J6GpcNq2IUN09G9s99HBggL2OjOSxpX6bORzrrPWua5O7kWTa+Dkr9U/+xm5bFvtVpU9eRAA/qyO
pPX9pCmHDBAoKJKqofqlHyxUZ5YW4VcPdbUBTi9kjWDs9T09tg0KHLBzj5VmkB8V5lodGH/aEfIH
R0am3P249sbB1gJbwQSCfm8WSsPspmiaP4ANEqdJBErCvSXd+gtYUXij3JUnNVvLvxDdQtBTfc7j
qgfT7UWc3vQgFyg04ny9HVgg1G99gdVJGg//b3hLiCEO+6XMtTo9MFrxow/Na6WQE4LT+NcC5wGm
6k26WPKjwyUos7W+RGXBUJN5GWy6VU9EGe+IdfOb97nJVIuxs6HXOk2rNe1V2bCRCvWXm2tTctyi
ccAnpcmvrpX3mRV7AyBG7R83IfonOKNUSq3TQ7GSk3IFWNLWMDx/eUtj8KlksTNTdgIniw1KaUGq
HYl/Gjz6YMHnrxm6M9wBWfuMFXEAxzBO4qHhk7yfLlsnQpDG9455WuGx5NEyzZdJsEE+AwZDPlzo
Zf7WmIghBMZiKMSWoWpjUjmgfj4Vdzk+EFi1f0XC5hTHFztpuPTIknTbCZRt5Y9rGtbpL7E55n8h
EFDwOwCBIjxkf0MluGz+MKHku42VWGAVzejiQnBiwvOPKLV7V0gKv2uTkNSQevxNs9ucf2VID6eL
8AF0cYAMWQwq/EOrjY+v390fReIF4HEEyIlNuTiC+FBuNDOCoF9ginlvnzMdivX+X8QG2nfvtSpc
OQQvIViJHmmkp6RxKJrFU5CLrt4NQRoxW5Bw71Oa3fZgtqjZS/am3Nq8TtV7A9tYX4KCY7pb0koh
iHUPnrVHmMIl6fzsTo2v5lz2Gpfpxil6fVYhT+kc61zFZjRgC6SvA62X/3RrWQGYBxskX/JmSJFC
x9VRWLWYI+lLBGTFz7C04K/dDUiFe8SA1aPeis717fFKkGUmf03H4i1sK6s1aFaT3wyX+0LtNHBt
LpqHntrY6uX2FQR5SLOKdZG6MFaer9azpKdLDLUAP+yL+qbYqwJ41FnF4ElugimwNJjvtem3gRU8
M0+4NZJAcNrAKPu7PwDMOgG7fo199frbnXGWUjxVv33CzDCFF5E7F68RqPEf+wcMRMY83xJcB2qe
XIRp0EzOWmjV7xCWojpMjrR6Nk7bVyEDnhF7k8N2v7xgkO19QezQWIQCmpxD+g3kO2rIlRIvss1t
GXshK9G9IqbjXUyicITIK3kcefJ8wkE/sA33kz+yyJyN8EWfpZc5jWgvMgcjReS0/5DcLribhnJX
vrDy5QhO0T7peaQyVC5V9N+p7A3o62zs1LkgJ61pnNKWbcRMMyEBW4KopJUUgJ03Ov2gH584fj84
BFd79Ck78QzPQZfEOgYQwE3X0O+jdfvPVBik9Lo3SBaspIF56GUYIL3GVb6HEaq2bbN+xPdhEIZD
nzvQCQ1BmygxSSH8A9zFP9UNWWkhsDyRu/9C8NxGHPnpKsk8kB+cPM0XOyPSRqTsdLbbEZZLO8gn
gKQ1265B7dYOse4opVVYNaycUqFhOJRCx8BoVTnToRnK2Ze12SfApxDvoM5EYl7Fh9j/sDSYygCa
WUUqL778lak0k2rkqBnX8t9KeTstRc9c2YsXQ5N24a18oemtRm42EJ5Y+8y8moynwoNh1aPlHjqA
7Ivyh5tXSXB0RfW4FgLK0sYt8ot4tMierzwdLGbrBhgwhBd4iOnzsZ54O1g24TNjORE03iChls3N
cLp5vcZaOktOvc3462F+fspxdo06c/K7t/3OBRpLiMOFvWrs+ElsdYLRF8FzgWZ87DJFlthiT9Om
VDbQmE1pQ9h8aIBjZPg/qiIx8XMKDLy/T5bToPn/VVHP3NjdMWwAK/RsoP+ZaxV1NDHoGRGgEboh
XTrxsXmJoxonqVV5E1wgx4jmnVG9Edl285TXwq9w6EBOI8hRRH94FomCKWQVNIUD6WIi2kDRMUmT
37ueDkhERPDgKTlM2N9Rz7jCg8GcwLWB7YwKOp8lQR6Ae5WwV9TsywfhH9PaEfq4/l4ygEHoWVQl
xrCCb2U1nU4wT/LcjEkU/DwO20hYVRKv5ilXBBanaRtiAnrBBad3AN4oIFH37FrccDekH7rSFqLJ
/nMzvO49yCUil8NL7PjXxECgcGq8glr/hD0Bfay7KK8uCZVUy8+zjPl7qQuySwxdlHkw6utL5TwU
g5AdlkWGU0mEv6On9DLZBnqqHKjp7F98/S02BOIpc4o1jAdqIvhKAE9R4jkF6KZ0XJJG0SxZ5fEU
zwP7d6ZYPPs5IIxfK/k4d+YftfrYvNUP/WLUY2c0AYNevcqo1YH0iDAPQyCvdtoCtku/Bqp10CGv
cCk0fwftSrLmNCRLrcP9NwtgAigp7/aoRE+leQha50RsMj4Cvks56r2WmfHyHpMXaEnqYJSRfykm
IiOJAKmUj0VoMUBSTa5gQuk9u4/IQ5kQ1c0wGMQiUVt773q6KONTbtGpClcQRsSVHMlXNmtStCFZ
51MihtMXvRzf+DqIDjNzBZaid1Q+ygc917a2+EMYf0G4CHtKCKV2ye9KScuSBaguW2KfxnDC16hL
iyLPbv6oeH/jD/OB+qepQRLOy3RB5m/xQYM6ZU7PE9+6YK7NsU3Iu+FSFD9YE83jjhUj+/oQsrsS
L1NgdTIE3s2mAcYcnkrO7edit6clt6aYV1IsxfRXIR64c2B9joSfPzwECkp7fAp7zYfk1gGFFgAi
w5Vjw4dGUW8cSC9zHPdZocNRvc906R2C84IXWkMZgKld9Q9K6Fo1oSdYbmxOnyZ2jbuOFyzg4vxK
cgnwSyhu6iHfTVfbVyE/VZ2CAV3loExL+orlO9eT2hQtp0L+8f0QuyFrDcX+adk/AbD+rldeMkNP
evLqbx6QaoG8ZoozLlpE5pE7GEZk5YkSnkA2ycx6N2hpVgZORKraEfZWn2Jjr6Ud/L77VbDSfgDp
eLlrSBBFb7Vn5qDOahBXk1jxGb3GXGF4OZ0moJ5ZvqtRt4F50BsrUeBaHc6S23MuFiEhBgfw6ldI
9wLBni/9A/zxeXXIu5u/j6YpD4eqrkWW6oZqQOvf2qPy76O0Pvpj62RBH1U6q3i02XyWy5mMqB5q
Cp/wgLX+eha29LvljN1UT6tyGGo1dualmxYXrvE3w3VERunmtoAfRf126SdsfpOvaRjxepBJnDFU
akLVzdkxENHerPQ3hCEyDZm1zyBT+RaaPz3+8hEaW8liiGni8P0xR4PvU90cduYyT2PT9CeoX2rB
2kfDlGZU8+IV0i3RnHaHkfGS/rJ97LNH2i59SfDtOknOft0lGkmx7Z0zVi02529Tj3btMV6DYnaV
EAMT0J3zekfCZU7094M31yPbdQ/0qsts2SXbv18eqx1FVNrPxV6SKSVBszNkgbgKg03aPe3ShAG8
INFk4GFhRQ9kHuyhQM4j8ABtPF4jXzXRx8xzvghwC2zKWH75tJYS5Exaq/sPYtTgIelbeuR/du3E
8EoCHTWVewBWBCYrjX4TsLyFDTZb+j1qd5RRpjnjPTt+Uye0C+XZZ1f/8PS6AHjtNQEgu0d/M0qc
Zg9/qCiI+j5iFE1RQN8mE8ZcrjtganbW151WtrycgBQGUYQ4Xkcr69CiWZjjFmcxRh29HeAWClEe
+iUfEjCi/nas6uB8oIKIlzeeVnbiMO6/LoCMuijaeHu4orMy/O48pfOJ9ZCTCRhcZBPUsDbxHhQY
awGTWRoOZrKNwbT+G+HciSC2YsroQPPsJ8L442E10l/ilmYfXmN/XNJtf0RGDguSyKpbwdxWoWsT
NiSWr21dWw6+eYf7p2Kas88UCuzJRibBetFvqj0QisEjf9ynOzlgqypabI/HTYrpkS0HPoVngzuv
bctR5PumKRibSkFtXPBwvGR2A7QWO1X7EHsWX9vYVxnFVKwnRKeAa/DN6Fuo5Rogd8qCQ/w1vldd
U+mY+60ddWTJ29GZ4ZuNyEAoyCdv3XmVzYMYBPGVG7YiG6kUWRahGZqITDP8Fc75NR3+kItwriVd
dCfCjvg6ZiMgub2oLbXibmHUcaDPij3bMjLmTUgF1vzNWhpk/yzLZrtsbT8uI+/WA/ea86WMxYc6
LSarha0S+7GiIzyUbJGqHEwdskJ6IbXGPWN9yNHog74rQtBZkBviHsD4RuRWDVlgvHszRBM+YXHM
Nv+PsQ9esRAekEg2XIw3zV69crH/J+zY2s8zHrU7adkuo5hGCo4+aLEY7pJsbxPAarDQdgtWmoul
TiQhNOugAbVxU41lIATXIZvnqrfjZoUTdDSzFJirlfpQw4xxuqOCzO8uQ53S33V4H0ku2bDoPtsl
ZA4n3xYiSlsk82+tDGzFNc/1m8GbkyXET8zlBnRFYnVwzx+cJZ5O4wcBQgj4+Rtm9kZfgk+2UBSo
VY5u/acD5hh54BGBVOk6KG6w7Ws28dMuN6ysFeZzK2fkkNThTkj9tsNwhWAKYweHLhfz/KycPwUC
gq6b2Z2iemeLGRPIlPcsmwCeYwYUm7It9qMm7ZVjJJvFjPcjBaIOrzi2IZ/mTMysrgvKvL8lX3dD
KukRH+S9Q0RqD/BqwuSx53oq3VNwaKoaACd6P4kWzmGOajgaNBFDhG6aJwR78eFiIei+iJII4Mxg
R87i2IrWXUtHHVYgDeD4v0/0Bywxjd0mq/MtPQ/1CgKAtISucBRD6AfDgrj/uVk2HEnTrEYVl79S
xE1JUAkhwmO3zglTj4bdiTbesGcCB2Tf2FK66Sirb8XfWGdwfvbUeZSLvOo2vc/x70rJbjxeExlF
K5Uo/Q/n0TjAYUfJ5N8OQhWFRBp+9KcTRFGuFPK0oNv4sC9Z8wylADhnbrFyl8mAmGCmLzIK3GUd
LGEMO8xA7aQkNJHgH+xlNwhPsAMyDSUwB49R5S2dLNEotm2qusFjqWxqUyLDuaYHFPRZ0jnWLcI0
x+0lbOkFPZNc8kxKyLsOp3D9LTafLnNUqf/mjZnLege4qOMXVt/zuIU2bkgUMT+mM+xoLmHXTE60
s5n95auqrsPvJtinjSc2HL81F/NsqJTukkvKpyv/EKVcV0R6cZpPQegdV8Lxor1ZYu/u/yCon1eX
TlWptWNVsc/RMc/+e66mTFN/HObC7WDfTRmEbIPUPe4H4rVw+o1l2X6jbc9SaRxxvVisJM6RMXei
xlhmnUvIL6QYBebJxtEJJGbbARVRckpIClb3kN0u2ZLqTVII0I83AQJDLvyXkKW6fqzXjitYKjdg
W5Pv6ikuNfuR4AlST7iXkz7Cz3mR3xpjZrU1RzwiZpM6ASwZSYAsIC9S76l0r+QC6EI2Iz/NaqRD
GPxFeOhHbd0rk/NQZJTQkImQjBnCvw2W7MVS+6egxW0ktKxyHXJIHmjEUQcQZF+jBJ3L9H+Yw/xT
VKPoQgCEHxOxc0cUJb4DtQBXkOHD1iFEFerL0hquvThds0LEIHHe79CCrFSHHdl/4UKOU1Hgu7YG
gX99vk/a3oIwtRU6QRRLVl+3W5RT4F2JPCM5xXEdEdYhNfWQL/CjVgA2DYs7L2sNv5N0Y+J6bAzl
2ClbfPaRFdI7ddv4QOz4qekBcEu6JHBhMzsJfni3ZciCh/2ITtR1R5c7Ve/G5vM3+wXGcojGvxD7
aUgicWj8a+d4q1Br+Hv/ySblFyQ6tWaP8IbRA+nSHQqwBY6sm+LcuIamUkEdTCHpTc+zvn/9tdEi
D0DoydzKb977vDrMpMFBVpeofgrMIbzcEM2WmzGZ7YgTYLoUjjTlDF0+gE7ZjLqJDW5VPDALITh9
C58F8/1KPQTrus+ctxWAB7YEhUNngJcEOjiLqMIXy8pQqqRDMIpAAGe5zYARAh9qsxZRsQK1NcHI
5grzO8NjkRyHieZbQMXDOeyincx4VmlVGu/c6wimCvNlJ3Ctq3V/hprTzYeTRgEurGSnv8pQeM6g
G3bizFuHQlvcqlk7p4N4UW8+arBlUhrLiqeSYCMF667/Wno9A0aRMfl3e4TjySyUIDmCP2ztiMa3
8JdNP38r3DjZ4iQsJJJbIQ0BbjkLQBp+jrVDz2atvciKh5myV5uR4BswZqXEepzUX1vsjs9ZE8NP
1hSd8DZoIgiTehHNmN74Szwh2QsxzqvVfu9aeSEFxsyOf2q5nTDjvFinNOAHFv3WWJGeKM1uwP/d
wbU/KCgWF/JRT4jvYbR+92/qjxOKPjXI9cP4WzaTauv3BF5mbYrGSRgkSMSoWl8gIQRZAvUaGYF+
+DotQYnYm0MMCIod7J8Rf0qfZYUg8chWzoJzVbirSycSDQ33Ldu5S88doQXJ/Az82Rt2uCgHZUub
UeOaoQNgCTJhj0rCcfUOI+KoCprCO5UaK9cDRXJW1SEQ4Ax/dzOPJiHObPaOI6vC9JGwmNliVltF
StBiF4DwV+1FCsgHErwxRAT42Vcnwa7wxOwHF0+c2Fbs5LCNBLB0yWoY7jQfNl2i9VofDZ/ANrW7
8PuMz2nc/76uTYBXoGeehq0KLkUdhflsS2s2Oh2tY4Sukyusck7Qu0vSPNzPAvwI5PVotGSLIMyM
78JpjG4CMKVFM+1MDi31c3Sn4B/hm4MyPFFHHxftUM8Imvusnx2xEjszgRxlveR0Xhr5g+JDHJLv
SZY5L7+bM9D3hxBbJmqHEqKxmuwp/2IsMhEQhqh5o54DDuOeEGAngDoLB1kTAka8WqwF90WyqwAN
GTQ+AjNPmNLJwBJHtkai8aWgTG/m7TpgZSC7b1WdduYbOjlsMGMNTAoUrORfCxey5/bRv8XGYAd+
ydpaIGGSej0j0S3TYRb/kNWEXnVTL3frIFP2fC93W8TP04uUilV/AEgcZzjwmLr2uwCSRespGRxa
xBr34w/5nCIYLKrZ3ENSlxoSuNExz9wvdRO+5Vl611h0K00ZLLMPdOiLAbSAS4OxzCeAyPpuOWHo
5TS5P5fSPo2JUXIHvrER33YqsfeCxvk9JFZu7+H+oztYppqrm1tFpk0Su3GR/K8JM6dNNlhi5LvB
Uw9o5mOIw1HVPP5P9PsPWfTByQi+kw6a77ykgHxzqUiU3sTOYDaFkQWkonTFiw0dWZfugoQWHn5r
Nxicu9sTsvxbsRIS0oG/og5IRX9WW77/WWFnf9jXmNd8YZAmOPrr4/MSTmFNuS+2gZR/Pt592zHR
PWhUNuXKBZi+aWlKUYHTmjJPFhzHxKddk7P8isRqqD0/cwiqOp0kXxrKOZwDKj5odPWKMxOrvEKq
Su7jZ/yvXgYrvE4ofOAYQE/Vzq60LAT5Nm9QUpmsvhGQhdPoReY03HtClnn1FGxMlm8w6s/BaAp1
yudw7gI+66DLrbhKRSJVD5I/cKP3TIdeXGbPrt7gxQ5F96GmHyOJprdh9eVXu0pBY5LAVvRIl3bi
rOtGC3SEZmWCaGlp+OZzT5YUFR/RzvaK7bqo3vSWWTDKWcReXySSgNE6MXQs90iVmizNgvdpIWpp
y1wtLbvMKE5wAsxMDp6g6ceQWlyAaKtfj59HAJCjvuGtvAlnjhJFA2V3V8MK3duTIOmuJdUm97Es
Ncg+gtQS38dZufDESXt5byUohACW+1vhzBVg5kO2x55x9Ccvbvz9jTJioPAJZlHH+TsvzeKmVRA7
Z91oOcYrT1v+VKRsYQoMa66ZovchOWlQKJudlQ/nPmWvJ4hNjPsv7iEBKgTjfODTUoVsKRbfg0YP
MUI6o53eYVBK+jThsN9kOHcV/2PmZ261m8/7u/CO1HWvUiRn2x97/e9IKw0BAOdMddJ9mG9ZHkHU
SWrqcm9fuPKCLh8Djtk6CIS7+nHPaP95sOsXD9BFQbbQ2byOydzOuFLvlp5eaD6YxC8zZihaqG3X
3foIOmPtdMEMKFBAWN3CHIbO7TkY3VuviPt0RGL/6R+Atr2skmHXQZ+6bunT3VjNhZFAg2d6AVl7
kRClw6BSXsa38xET14mJ/ZWykdkRL+k9jj/++PpVcq8ckqmvQPf1CrK3entVgtO6AYI8fM/HxY1F
eNrq+FdKNf4e0qKZolr9UzHPntmX1FqEWiUa760AlvviA77Y/SjmnupZD3LcYQ79VH4YY7iCaBW2
gYVDpIoqkHkSzEIzLAaDS3t42nZbldJ+qgd5Z5uBFyKgux7ThOrITkhLAR+oeK/cAem4JjQ2YV87
s4/QcyUoJHdclh7kvMA5Z5r2oss/in07tkHgs2AJZ/ZnM3VQcZxBcmFIielkb8O6tE4HjC0ITUxJ
ZheUnO5l9whxtkWOAcm1DUhtBtD9yOoJnDPz+uM3qhEvboLmYtU8Nd+5utwV8fh60y69gYJJ0Dub
bcS5sZo+KtwYe5aqdvx73A9jn+cfMYSkhJngNt79NC715Y1N/Te7mzj+j+1UY764NznbKz33P7jN
CCI5qXElMBxEC9GH1iW7gRIC3C5BHCu0SCsZJK3lfHgrleTlCc6jiAGDdJOSbd0EvQk5htRpLQrO
EU4C+cjNIO4b5eSYteNus45BVCOMp+L1vpVhPpAHd595aQq3LGjhJxLGBhpnrFYu8I84lLnASqeS
zlXWQmukLNe96GtZlt3b/2SnLsvDlgC/jm4BR3kPkfkq6FRi76QgPS4GOPTFH2u9O6YerAX6zp/j
r9ahtAPmOORerQTlhLS2h8uEvtEBd8SxLM1YXn4MqcSZfAkgEr8yP73UVMrw1P4W3tQqdTGnDJyi
r4qtWS0ZQciF0ITedbgsOi6EA60+y2bZ2oNDwZD6MTEUX9/zbX+FGOwP5e2ZxvR1DdhY7Ik27mby
KalIIVX7KUnxAlTcdNBR0Dje40DIiPfqLve4J0ZqF2LQFwQNnw0wsITZYZrbokum6LxGolq3vSUM
zR+2Repc8DPKssAw6LAcUvgt+KJ0k4Eure/8F//jLJxMHPnHXeRKImiAaIkuMwKaOyiaCqFL4kZj
178FWl6okU7Meljw+gI4yDqvGoq6JmnE7ndklzGTbNEnEUcMRYnB79wRMXOZIsVJXgBKWB0fkLFQ
F6z8IntfWvPMnJZgmmDOO8AHs4Dx2qaYZeulHoWxm+scRJpclZiLTMm+Qx9eDr2A55IytIov1VHt
arpefngSrqPbH8i2jmfL2su8Vxzy7kvBaU7xZkns+LZXguM09dkPxj+FUAuNguyCHD8YU3DIY5NB
uhg5nB5QQ1EJ7kKnZjhXHTX9pNjMCXTAGXTjieRO1Z346UAtWmmmRGW5IY5SmEeee/utTYPc3n0I
7TrDsuu/Nr5gps4mOm8NCG7x8RjnRmROrGmD8VcXQq5WHLJzG5bvuipTsaKWRtDr0sFZLt75o4dk
hxjasgHp/zV3UxPkS/ln7nn/SgK43bDUt/ewi6ANBE5SXlgCASHLmiZwFj3nUInhOifhwqnb9EX6
MOb3DxMHuUE5/4jfwzrBa5YR5XxHHrIh1WbMvT89MKq4l8kNgv4S/Fhpl2QaZcz09gJiqcYf4gWY
B8QlcQPvsJY8FP1oVXI7zkqrPhClyCGPGPag1C7FcAvGb8bOk43H/IbbggtPKyncWlsfhjc2ZC6c
HK2sY9RpSdINV2g8crHMmcbVmjUbC547kHor+MkQTMdgFvU5JMggfSjL4SFKwrOmqRvekXWo64fa
q9kYq+dSRlBqtZdEt2y9ke/n+2i9lXd8FiKvtOs52xgaKSMsoVVU8MpGyrlT+POc4pJySZZ2zggM
DFslmkyHF2NMPWbFw5nCPH1DhBP4UJ5o6QYHDK3E9b7MpOV0HcHhWKk3jAFINUNtLMDra1PvhY9k
A3C8EeHr/LYhXFtKHwgpfH8ZWOgCkisJ6vYT4/Vm9GpYI78d6i0VC/udqJauHI1IjedvsMUOdJ4z
sM2W2knsNLCFrDmV4cok+w+e5DQxEdTXFGHxgMiXDUXEkj9Bgf1o791Okywve+8yMwatUiA1CxyK
fgOqUD8Bgzn7rOuqogrJ1jUa3J1pkK68dX/x3uuP0ZWsLkEQF9hkjg4sEKFaIe/LWPQy1LAExAI0
wrMZqzNDDpvY/PTOGBunpEDM226NCHgHqXxA3EEdW1rtuXkHrwbwMWO6PyFtCZyB3IBVMftX1Lft
QJuhTwyBokBTaI6zQXwljJwzPAK/0Ky+6aoyMVDTJBxp5f0ZQqEsYqnbHbQXGehIiJz81GRgsu3Q
rAcOPz+cCfEVvEPWGEWz5gLDQBRfUKjOvlDSdKu7x0IX8o+w3JZpQgDPvmwwDBshbp+Lf5fNSUWn
WSlU3r3m18TriojljRMFfnEv18ygpyPHAPrJAHKmugEEvuFNzlCHGTNXf/7gqhGob/BkjpzOw0va
oiCkE1vTzfPwlvQAuWNPltSNfY2RBJYNolrCIcIXow59jbI+3SYcGXdBrtHOtPIuusmiNceNg81L
1zyT3LAEM7pG9zXyvLLFsYvfl//NplqSKITE3+J2GDnuNcZZL14ZCrv5QuU959aQY/fOM3hhXaEU
evFzlWvFh6L2VqUIUOSeImTEjJzFXgBuWTHN3cSSeeqQORXVpUjb4H1cRHDRUPDsak3TE/V/8BNz
csOmPItuBhGSslm1jTlZnlTVd+jF7JPO5cV+VWL27wcR3CZ//VTRZQzeVJbHJJ+FvV2GB43Rjhh0
PBtVv014potaGpNeY6m8AypUaFH9qTJL6qyv1K55+VN1PfmiuvJWLBLkqz8wDwk2ZHfAhDa92KHH
wakA1QhPg0Xu+BrjFEzQeGeHdLUOjLWMpUJtaAxI06/zHpI65IZY8rerym05U4USbXVcBqZzIyPB
Gn00cbUoLJZFqcgJ0uYnq8zS9e8kzLZL4su/sN1C6CNrbwilwrmkC4U01k05dQMrwKME17qOii17
PokRpIGb40Xtu40m3J1TTFgz3L/zkHW3Gg4lT5Jxgx414j6U6JutSm2W0ExpC4+0Bgwv6F/kRN4b
yxWw1lO8S34rKVdlP1JHOSyzrGAeACg3DYoVvEltgq4XfcP4UGor+AFfJnUQVHTIj6qh0dKUwoPQ
LaL5wo4TqYkLrQDYKabHIK/gJ7giMsbh7QKyo0iYNXrHxjImjgOGUm/6vWdgeaHbTyv1jPXezqOU
kCeisqNdbGAdye6Zerc4AdMVSD3Dxgdv0RiyOn9D0ValzSc/85gA2Y7olTtzNw1d4rMh4CT6pvuI
Qd04NwBBbfc/+6A7f87xnQnttS5gXSJWslm4uidll7Vi+Z6kmuvCW/We9eZXk8YdujIIu78UJDup
EhUG7MhgiRFBirdcVJpS3kO6qyNNvfPF1aZo8Y03K7D/3Np4jvYU5K/gh5MgIkjjge6nQl4m6byz
V+rRmqKxPXmqDop7TlR82V8Y5BGo00H7TJOnE7QBrGHJPxy6UOOTetVpEFEaemrWJu3yhplmtFaQ
5saEIKpt6AM46Ss6QJ1Kza+rJllsRp/riHHB7N6H2fUNT+RtnNjaGfXFP3q6ZhXkiLMMhGmnfE6p
kCmSa9YhGx07vlwp8t5R7/y379lAvD6ZBf+Sj1BJuj43zhUNwc9O6vh8pUk2/YXt35AMloqDDhXD
4N+OE6Cqf9Vk52mvIX03FBn5qKqq3FpJlH4MK3jbiPcleZzmSgexq/Q7VMHd7kyu7jh2ZlfGRUvs
A3ZBu60kL474f1fjVcxlhWDPvBvc0FfdlcIIEWzfScpyuu35AwkBM+AR2CUBqE8IsnVZvfdQ6/YQ
nPxQ5pYXFZl2qnbgQNtFdovDjsGtXBmhan3USjH97r45MqYxD74O9hOweNosTXI8pjesY7f2UbOQ
OLl0f9O3l01B3k5LnH71EZyyfXcY68Gr+8Vxlrp/3ZZzdMPcIVj9lrpQm327ECh+FtSOBRRDhdnf
bPj7fS/avnj2r7giEHcdF9c0kym/rfUsKiPnU5rFzN5M0rOFDkhj5+abPvaeD0iinBQ6RgFgurra
Rx3PbBTU4Aiizhek9c1XVzakxX66G8+V5CtcZarq1w6I/9E1dB834UwVD8c9Q4QIJLY5MbmnfpSM
GrAX+DMMU+2zVGReJylc5Rjy0o2WSLuJ8VEsTYp5g1h3CIo4yiHSyw5+71hWCQgnYMLW5IAetwsp
4z2YlTo5EV0YWjmetLUM716g7pgfED4mMs+DLTTHT8lSPeAxbjBXsHeKTYdmAFUqlQoGcEP6K1ex
CiAH72UaxMqz6NKzawP5dKfrH2mO+JKa0Bv1nukuVOP06iwrD7njHn34TOePYNRoTg+fBS1Lo1Ng
fDPNBTmPjRVM4AMCPPw0njjpRLmyleECVAq3lfYe5Aooz9ck2BhHQp5W8HATmLwaLgk3iGQqHxam
5p1zBMKWBy5llB+UYdixeL9XDBTHOXt8OGTsv/ites+aJMeke9EcLzgHdMLggIvvMRpX1ZegHYyd
IJaNZ6usm9hRUjuDGo7LVto+XnzcdEjWAabBEqP4e7prUPQD8OrdhI5gWMGw0mgpSWUj0FZEDpVU
zTPgQmoyBkAIhWgfpxIsRNYSh0M3MWX57BJ3HtNw7AE4bPbQkDKWykiixBfBYg1MOns7TAM1Zx70
bWKB4i3L7ibSLa+YhLTMjDNYaNCgcu8g6vz8StzmJB/JIsFStPaXFO4ER5vIhfUrtM9PRbGTiAUc
n9ZO+eOhioJuzzGni5p1AQOGSA02Nd/XG6UBfLhMVCbm3RZ+3Mpqi+y679sLxJeRJXkoYZ/9AeZM
c9Wn5OgqN6o0Y7+pUtaxkSNCjDy93jwNhPEQCnkMEd0Vasj3YxOs8gNh52VmkloLcXOHVVBJ5CXI
fN5lRO/7gZl0NlONdia4iuKU1QK7fj7Rx4ql7EGa6ko39bOpyrDPqJULymXt7Fnmv8Cs+FIuY5k4
0RlyLZiSSTWwambmw1XW8lK6WnUEko9uhpHDKMUlI9LrsOfyi8WVQuA8DJNc3s8UeKHiAhqA20Av
PNfrO1FZvtAPtatPGFgV0Jd1SEjFTg0nJWrSPK3fEHYv1brnJKgev3+O6tY9gAAFrZeqvhGsh6St
De6HxcMCAgpapURc6/ftbi+6/NlLyAq9L2tP2hMz9IS1OZmldcmXWsg8PTXPLuW/qPVsX9r5GFHS
JDLpHqptPEGud08HlSD+cIbYXsLbzXxepkJ9tWc8KWxs7WjhalCEmpdvFLzrWTg4CwR7MfcvcoZU
r2NQuKWgEjOEFuhIb1uUjk8BdDBhQaML+aiCbjuqSFJ5Fx84DdrF6QxXb7dsnmzcVnfSxNyoMNCM
82umsN2jGnTWPKS2PhZ0S4hGJ8ekzMz3jXirJM5vHOSjDWSbB7xERxkmbjhjUxtjRRTC5/T4N+Qh
VOhqrfzsZIW66GkF50En45jIWMi8785ekpjILj7zhojupWWOb1WJCGJ5Kc44KtlvTat6A1pOudDs
3b+dVZDdsYXDkWvCM4TyKSSmDYoqL7pq9Ys/WH2ui1ZAA8LE9MYhyfOPL5mdJPf9Gk7C9rKsRVFl
ijYaFAXi7xjuFMDJhiB7DAEGpU01hCN0hKqbqqI2MGze431NEZoSCyohpCE/heqgENt0uRRhSVFV
4kLoKJcKkPt66wmkshEsJVxlQ9rAvNLYGvz1eLqvL5AIMiHqdM4BP/5emPt+/lONkDGNU+X+a6U3
JAS8+j6XmHGgDi12NTcWe7hH9xyDdDXsk3AwRYBD/cSVPJ+oy0rVrY4p3mBtqzdN07uLe8RHT2Lt
UK480H/krVk5t1BZh8HUVC8KSEJ6z5z8gcCky4JaAJHQEWGoZKifof75SyLhof/BnCKPrK9qiUFH
+KBtiUYqVparp7UZ7pHe2xhCjSF4mHD/4798SgaA2NGRDCEs15MsE+BUJOTr7eGKkPJvR2CtV71I
abIvt8EfcD8CjopttBWZoxdF3DHILINMIqu6XBQfZhZV5cVWHGFaHWxncDWld7k9j6FfejyKdKuo
j8Y48CAxg11U2kLWsq6fgio63lrRxdDdMOUI2Wh9gWgagillRMhefsG1vWYyoncdDNL8ptT+Tt89
gXR1u0VpavAWBrssTyQ0ntYQuKTxOEsyZfpW2+C34iehlQLBDrnTNf1N/NgsClN6QCTRev06115c
REI4dWxVYDIA7bypkyXC/ovmaMieol86vvifJNC667ATEhdWQlleqtQhekdd1fKdWpNyP2KLmqex
H5doxuIfq4lfGeaF+JRjZ1Jng4x1MU/3gBwHe1Cck5W0LvdsybDSL4d5wRbEJ2mf0hPwAGmcNe0g
D/QabvH7Y5Urbde+QJIzebT9w4fb79v+HdRtHS4FBMvwvudvTXg/9NaxWhytledv4z1UnJB+pF6w
ycGg+4L5T1fEeZfSEhFcTfDTw237Emui6KkEukjohpZuH4BnBz48rOjmjRWubhwzt8QIH+BdPaJA
z1rmcIdOH4sjLTUlvXKpkyxrZMkAaIECmeovM8bhla75xfHyiyVUgtrliXqvyeJbPeV1lg7KvudF
HkG6S9ZkXHdhvwfPeXwH9uTwKHXDnaxSGb5vSjH0uF1M3QMgvYWsLPp5/k1BP5/uUBYzMXMZbh3F
HuSD0k8kXr4Nhp8yi+SxAnuBbVz6MYTrU6sXI8opDAoYRFEfRUiT8KI7FbLVt+QecHfDl1ntElYB
JbHiAcLZDOwsrQgSp9iD0m1hv40vkPtbPiC4kIDZBqJPlbbLRRtD92eorXj1wHdrDztHKCdXxIuq
2IO8oHTuXLNxRoPSmsOjkzHcqZ1QTIP9691abu7cc9mv8SErldYE1y+KSPAXnjwUkmksZ0kiYY3k
gD2Kwp4ah2CABqCwEDAGBMw1XxR0mp9J8ZldNz6WSTvn75eGhgeYbYUndqsrsp3IO+2vPy6zkIZM
KvUWohcGHNtPk8mkYWEio12lzAfGu1DgmxiCabiosW0hNcPN3yGSDNSHRDLzUwCBZRCikrlvSOSB
83Q3bbgllm4e53x0WCiKg6ThDvHwRmKgp44Le991Us8b9Fm2qjbLHBvvgDRsFuRyomQYbzpSZmul
yT7Y7SpzewtBWbBMLjGLhnrZ0oVb2NogtO/D9efXSvwuY6ETAFoQ0E0Dka318c4jcDayT098FBSV
526EqmP/nbkXLUIYHsKqxiq9eeT6CkVriKKIkLzZS7NXa9REqNoimIgN63Ep/sgm2fjgnt+6q3Xl
iqyRFUJJHmOrTguOHeK4hBmSV+aKCo3/7n4XRL37Oonotnua/YAhDUDe7kQkgDjq5OBfwH9MsRSl
i6d/sJ41UOeu8bnEEPHZJtKBRRe0VgQ+vMfOUMDubFSFvhrEHTguBnFGCZBLaamU2GjaRtB0VFFs
gbyNBNxORciOK8Alfr+mJSZp3A5hSOQ3zRQZYXrcMCkFRzZ6x3cp7YmDwUbnae/XPDnE7jltq+WR
J5Qn+TIF2m34xx1mCQVAmf5PLawcFAXoBW+Ldrfb80fk4jenyAin2j64F09m2FIiHA+k58W+nTs8
Hr6TEzjxi0/Uj5i/tAC0IbnBJKe3u8+8hL0qKndRwwGOU7pdogRj5j8P2rrxMR+9kXcJLbbEJTP4
7owCsVpklB8UtmnrjZg44AQcHL/l47EHkz5TG2NSCYc974gs2t1TEkdaycYooC1sT+Sd28IrgsEO
DA3hgU8u63MMShZn3M+mcC4yQf4B8m+yw5bFqT29DwsLizUvCEZ28WQ0SEWC76bf+CqUw7ZUAJ8F
zU9LRcPXXVLq12jB6A1uPMkAIz6plPBpCDbV7yr0VbudUuRySFl1hqWod6cFmN4rWQ9e0uJWZpxx
5exq1oVf4xRGTlWY9Xk2ATdkADMijd6OMW36Vf7yynXUhlEtJz3lGK4il/00KSD1iASY2G9k6Ryn
P2LxhnIGP5g87ziB1yiJHfWWsbY+ttZKtvu/hIRccP96MbwjPB/+03Nwndwu0XjiGkHEtyqIONpv
/S+728CZH7S+/ZBlvc7GaQ7eD61yeyw8JaJKWHnReTHJc4iDdbYLPQPDGmwyYuCDymzuAwuVZ5UQ
YWM8WTlFTusqZuOHoLmt/lwQ/QGOLB9lWrLeYYgf/9cCWX6KbnJdlK1Ma9a9yn6KuF/KN9zyraDh
nkhObf/NylL3BrhHc0bvciponP5ww+Occ2ELd+2HCC8PEiiE0zJAd+Mpa1UiACRv97dZgWp1ORCn
TnUqrGzuRCbsD5MEnOD1EDGLRjlCgywJNboEtCf+FbDTV69yZkrtfpntpEEEJqE/NKhQ9ClAKqGN
R1TBSzheMntbmcZbvkh9dSK/njXtPdYhhkfAJLru4msKtP0VlMxpy9ELehRTdTkPjWcnScJH0Nd3
9yKAWcGYvscNrG1VkUG2N/bUEhhtR4E4I5g1zs33SBa6vlKff8fnfUb2iSHMslnPU5GpsTZinhCu
p3guP3POoBYcVDx8kSttKD8Fb5L1w677dU4ScSqc/6QdxA7m5yrSqJ5A4XbBT7SaYGJhi/wMJB8j
v8b1Wb9RPpvaPVrZjQC4qk8o2AnxAfe0WOVLUNhfeuwOqeWEMmuT7viOBCAHZ9zMkep2aDw19pGJ
lFWHUEBu7NIahEuN94poEszUuMeD0aoVhfCnU8H5X+yTo/jd6vFQNiTmIgRk2Pf1aW/DNO9isAaK
15pprHlNKT71rh5qihf9eamfIwWcZ1WIMn6OuazzWy2h6EvOLu+kHV5940ZJXLRLkLourIOApQ8N
e7NZTKsAscssxNBbdJgesUN4dCvJ+Wd8P1RC9SlAilSoA9zo1PBwyn4sSVejypFfg2kjozjxuSg0
SdRlkArFzOo9WUoN7GjvbR+RZDA/a1TJQ0N1/UdIJv0OkJULbWdxqy9hdm2BYj4lkwY1b9peKgfg
oJoK05IT8XetcZ0+NFic18Fyk916kSeakkcP5jznP39n1I2oEAAaIV9R8bGqvMcrnaYxXhPauFQs
RFtnT0P0F4OsHH/07GERa06JOcjl1Rj/W22bM9KRZ5hqDAOLlpnD+8rYTUb/RpQ2fWmAT87Q32de
QujYMaqpn6CgrXZRE83n1SI/wqIQv8U3yjovtAeAxSFQ7sTC3BPXfO3rlEcZhCZbD1zUPBHfcHN5
+/KbBoPJhDF1d4elHhE6Jviicb5I9O8ugIExey663vv9lovIAE0DuDswN/iUo3Cq9vyE+anJNhkd
6eVPIM8PXQ/V45ghT5YkHyAUlVOib8FUobRDGPy1T1WMQoqI+nLLMF6lEov9CMYcpuzKwO9TisBG
a8MNAUBk5VKBSIol3fcpKrgxrYH3mMnOPtMBfLMpnnKs6F8JIpr7vxbTs4CYC15Gs5tr2EsiK7Oo
yag1YIqaQXoQNLNo557UO6uoDY0257bMtF71La0ZOs+HPx9UAGaaIGPNwTvHPOXJhE6Y0GXFdVlx
ORkzwStSyP71BXsG9xnGtinxpS7DS3iseoElwSHGCvsun4O8kR5br2frkxCc9KtP6V3t9KIe0ITZ
eUjJzzhEnrHFJ8nVuZuCaogbnkh1YAiJHre4PsmVA1cR/d4E3kO4Uc6yRZZFGFfU8lCzA49LaNOD
kN6b/ZA7WLwDL4S6BvnAFInM1i+ww40aaMuV31ZvXkuXDDlMG/uRDSVvYtxuFrBjApXkxJm45j5y
XiwuSwUKAQ6s4UjEB9IFJkat8suXvPAj0IGxJiXmDSD5DQvCd/j1/bOJ0n+npJ61WqTK685sJenk
LGojh/5c0Bn73MrIptBpGsPg2VfU8TuV58Ax8VLqDIh0RtPwIY67i/uiA7ybxt3bdDOmLxthlpQd
dydxeH7vAPm3N8Ow+MO45eDhgl5uCQVWhKja2zt4b6vPKEnqoZ6dbIBA5LvxW+++Pv4yH2Vmc5Fl
eJNEujI+4rC1GMyUz+24pwQUcPcWF/sQuxgJUUrR4lC9ImpzCIx4/aqV6dojoqBszJxbFboz6Wnv
b5j/qqvZ5GjwIm37UT+HR3iCz8QLrcf8B/lLH5HJ+JGLSXtrJlUcRxOvTHennlgQPiQ5s+sb1q49
RtuidAICi+kdaucONKYKagAnH5bpllZvX9Ihi3SXbMseTCjh5K4efdLlLazu2taq7P+e4KS5y7f4
BguJFQZ9IJT7eRt33KftNsZuQRBiTnJSCVIkJOo6nRdVXurShId8dUCrlAtHWMFN66gT7xAFc1N3
Yh+OZtFZrOkb1e98OBrQmnwrzT+DDbiQTu/QBkF9DLu2uv2NP1If4G7FM9NOvpQoE9AUEsybgl7O
jdKSiuiDhJrQfXzuWiT0cpOGuJ73qBireG0o4PLlMZd+4UigQT8WlyoYhCcGCCuVPDB9PwtxF6jJ
Rd/K8WI+bNJmIW4WaL80eGndGH1x9GUT29WPDMncnXlrFJreWeXj2apMazlEbB+q14Fg9ewGkDVJ
s156IA+fzEMbnoeJuWkAKFKoYE5KUSbzV+GnJg9WaiMS4K5xbhCsJR6t3AwSyJMsoG+VmB6woxx/
t4U9bpjFz0OtKMytlz7UVEPfnQZoL/NJgpLjg/5YPJ9v0z7Y07qWCtXZkmcl+mB75Jc70F9FBPsn
J3VXNY8SNSzLWfva1d+EIthgcYIq5/MeYNqJk6R9Rq6B9guReEB9aHGLV82Xe/tJb3sMfUQzRhoZ
bUn9cR87EsOVN2BfoZJiBP0FbashEnfWv6nWOQ9wMacT8CM0TH8Q95yXf2aMkAYGNryGmCgOic4I
DJRhx+Yw0k45AsC+F4m3Eh668cdxzG72q0ZQItzJpsE9vJ0TyplANwZr/iYepgNOLpHQ8HbTLdIF
NAa1+DQJcdBcF2nFw35hSfJqw/nqkNSjl3LBvCGKNC8QHhtV1bIrmlmkWrq4k4yQ3LLdik2uD+Xh
l4l8EWM+jlMGVnwS1Bjsds3iRvvnCnBbWnYGo7jQ43RCcqb06WQLDSrboTnI4TGNNwfMeCc56nHM
4wsieTqE+551c6RMzNscVXlXMZrtlI1UJrWolctKzfJcpem0EjfVVo+yA9uDrUz3jeuaGgB9NQwg
p/sgcSJzWshlxVl1t2bzXJqDHn3W0PKyaRECZE/v3+kVAPFy910X6kcXtBduZSg7mBd7pOxYOhe3
uj3wwsxzghPYN1V5uPKm6b0pC6EItV7+sEdweFbm/Han6M09yopqN7JLBMA6fvT9S8ntw8+S92pb
BgqrKt2MVYPhKybq7T05SHdFSaBQTyC1hE6txGE2tlTafXL2/WlnyvgNkCw9/dxQlYy4qpG1VvUp
qB4DdO4z2y+C76YE7xcq0cgiMP/TQjx3FbmHkxc1w1zhY0Am4tkQJOwy8J7ek/DOLEU+5skMU25p
+s9tzFVrSe7VCLiR5aVrSK6W0BHJzET9WSlN7dSsgGiFpw5fP64utLmQMMFncwq6fHT9TLfxino7
ic9h/oDMFrvi7SXSkxpL0qACuBaMxCi7M9q93dOr9b1jSjsTGr6BJ412dBCHtLKIm29x9T8DgKIs
QC06Cf/79QQUaJ00j7HCw6g6oDB5CGo8yHXG7lsMN2uH9eQBrVNNV45YrzYvSZ6WUabxQVpXQJog
2BxqJcJ/iayaFHmyHhqOQZFEX6mJzsfRrnngo71bCbXdisPmNxdy6c3ZjnKk37nGbW3eC2dFUq11
6q+P2HIYMAKfnK0CLUz5T0a7cSf1r+M0yVNkVBh5T5iAUjQ5JDL/gy0Z5WAF8Vnh1GiYLqVwPRLN
0cx/1bwhn0c9eWkCrtJ/KULP+heiSK//rFDJO1CGvNC4yFvxE1YsGHAFA+AbZxsRrqfV8cChyrPD
wDK36sn7OnF+m7gGuuaWNknBo06mnaIEmumQZNc2lPSSB5SdOn0p7tE+WBa5c23cXeyb0QvY/VBN
IWnGv9EiymP0nqX6rt0PIVe5Oo1ONqLR45zdjGxEDGBBolEOWOQPinpZ8mPU8EdtDWUPciY+UAFM
uHstvqXD/Il4N5G6UIRUMSAFRK7Ds34jDKFe8svQyaK9pGjdbZZRz7nB71VNsNthMSuXCOffZkYx
PhLO+UQ+7owQbcQBmuJihX/9OjatmDQjbOjwXo6lhBXrv9DDSkGjVRA0v1xZBi9cqDgmpW5FAMPu
fwYmTYj2Cj4RnzhCzvukJzcx6g5S6LLQyuFO1CFeoLXm80bacxug8yciO9VQt+52nkNXqsOvWfVV
FvMlD3ABMdnCZ5xyf1uUFgandpp5stmwntuH5B6SlavXE1Usn2dgAXl/bVnNPGMN3lteRb3Bg544
I/v+dRgXgHHQo+t7rWkc7RmBlwRZlGce1Lx/Ccz9zx9o/4Eiu7+UOikv3h8wVFNHlAFGDP1oDIUK
/hNMYjFsetB2RfUBozUSo3t4jhH7MMwdXxqvEiB+tsA7jVwZIaBNi2KH7MbJqnI/ciMWoZoZrLQa
a6n7buiaIftn8ReC589TXelH/vEIzo7OXgjP3fQRyT/FhlF91PPKkSdfyW0Twyc1jwQkTDBglVZU
rr1crM0phSrnZpZuprDXvotyjCCGRhqI8Vo8q+L5kyLDNQMLyOGtmu6yhUy3z3wJyHGWxuX0aR1/
MXfILqJFPPha1fTP0cFhSB9mk53KnEouJQjdvZyKGertqWPS49p4wzGGE7eBMlj8u+pMFOQjVI48
9H/BZeqrPS094JinRc2AmVgDEhCz4Tdj0FtBN9FjxPBe9uOg+jJOt5m6z1RmgsVJAif5DfZsrW/E
r4Lh3shvywXtdxD63yUsrMhpB3andSBA858QtyMcfvNg/6VS/CQ9DibKSkBHqQUtk8ndQj9c2HQ2
XItMDzka0w/bjggvuo23dyrcJ45aVwIWqH/QXBA7lnozDXfrUUaiBhayOmu77BKdHwx6kpCExtv2
Cdvmzj5P2r0eIi1lnJlhJsJBI+BmYeXVlmCHjAu0lw90oWeXolsSGklal7of602LIePj4cZCkNN6
jO/nKSIftkPOnkvWGGAon1Jh0MCxGwQri/3LjBCIBlUQ5Wi7l+Hnu66DEqQlSwDkM3ABid/60g64
iaqSgRNL7XfrdYENpQXGEOw+rQ/LPmDbCOoTA+RhFXGnOLm5IaovBD6eahASI/yXdsS5+fLIh9zt
HbtAfdxFjAx+j/HstiMRwo1J2nri9ILmOdQcTOqubZDMss6cfaWHcIoLBTsvScTfaJhgGZxT+xEW
ZEkDQPLapG8wSqsMR7Wn5RxG5EsJgGwtEE8mkljcyjJNY9MUzTRG3EOBeHWtK3nGLq/B4JaoDV1W
sRVKJVzRmmkG0Zki4m80FbUwZJwdtd2Q/8mDPQaDRzmZCxlX10vUZDrp0mr2C1e7T2x3siVhnD8c
v2BmnbSpZSqc4ALaVuzzBm8DY7S4Uv9XPaL0909/mN35LT/fEBuH9pp3EWrO942FIVp+C4KClyeh
4wleZhr1ZkXfugupRSa3hJtGCkyuDlAdD0DJPI4/rO3aZwe9tl4+U0tT1jI86GO5Mo3wBPJPbKO+
haqWBV0ODMGnB6Ty4waG1/zoJ3x9eGMizhtPsoxIVkf3mkQtxdgBchet6g86Djg1PVSdqkDGHSTh
7h+UDDhhIM1ZSm33QS4zHV+tId3TGeV2qgOzO1t6HbO2XZnGs03/r+quUvH4Qta5FHieZrogrUQN
gv3bHbQ/UqFloxfQpQEzau6LAWrVzg5EZBbyLJrJrhQcqhIjswrkBpo2JThuo73cjHgds+6ft3/8
uZclKD/38s1ulzpXQEPbmfqTEAMHhfpGubzSXgwGXwm76xChLexk6Ni4KO0BW6sMu3a1WfwzZttQ
CY7W2hEL9tdvBXpKNtWEu+Sh+VL2rZziSfFXEGcWwN3ya2Frj3iD5Yk6irnjlimR43DjyJWwdNqc
ILRyoINMarbI2KhlduC3MWBrpucQZW2xp+3nqs+A192AQXDaOrNOG1dRfOrHtsnv1eORhglqR3u+
ZpHSP/vSYe/nybIlV0ea+IucJYGqe/wa4ufwNJOUL2FrcNrY/hZHfH4ZYkap6HyanuCD8zAXFKyB
uIn4lwaKYQ1CgKiovMsGzfgK7K9+1CUE/DekctBTdCPXeQs/gRvM+Cu5gT6+Md9VkdrKH8x5BzQ9
DPbXwIvmp/CdfH/b1rbwVsZpf+SzB5nhnZM/GjF2kMCuTo6gYnTiJAAzD1OW5vKwdh1SZ+NcqT4U
H8QCQkFGEFTKFCQAhSTloZNgGYunPrSjXzQiS4FKEiMNkSlbIbEYAPf3swFpnh9/xaORiU4d5c8y
iwXNVDNnYINLozd5aX2r61Qgu0uHWBIGwTU37GzRZ/aafaRT5l4uN5EaCqf8p4cELPwVrSkTOBve
XKU3MNAyiADrlEbnKDz6u73Hl/OH2UIUzTMBKH+RalGbvU2dQsRDObfa3MVti9HEn3m9vIjpBWml
eODFRKpcmX+4pGG9YAnbHZXk+ezrDpb5MTPST27yDh15DMqoK6KWYNFJrXFx55eHnWHp4kiie00O
GnMbpPUeUh7zn/++1nCNPB0mW+KLYK/p+NvB4tRFhtoiUZ9vDlZuoNptg2QmhCfmRXDE2jmTysbE
tk+Bk4yxMhmOu0dUOgiz++xEcCHOJKt2f28v6v7MnwiTdr2ChgO0nXGwkczl1ZbrjOygWLORoouH
bm7atH9aNW1JcUIzDu7U4vM0oob1jdtXWyEZQETZ9aFXI2bHL0rCfmG/nRS/EFRprjI+3GOBo68W
So8Z6PC3rAFi1q2S4ZB1aoj6C98J2fyQGdCZSuLmPJ94deN4p/afxwByNt1F3BiAh/2sOGou5Suj
8bWQQjyt8FayraYUlS9foytsjGhPf6n6ALm56thoe3kK05HuCQvi1io+cYYJPPNd634deBO3Nkdg
go6k2ZVienEwwAndzFwxrWgBxQquFcg1fxpgJOijtzOpk+/ks6362TicSCmqFhwI6t/PL0I32yBn
Z9jeF5NBGI0b6Y4nkjMoJezAt3KXZ5ZX2art4kS+DJcrkKALM+5qL8dNHXtxgJLUVRS9nLPzboNR
KHRHoQ2Xo9CyR2fqqMC88oMOPKYp+P90VMNSp44XPvHPcLnG+rSPkowhxPmwXw7jdX12XDYM7eFS
hWZ3t3lWUY7/PW9J+OQOL3WZh3gKC5y+1CaLtcM0Hfgz7jo7d7Tqw9+dr9NRJxkrHDhW+XhGEri4
l0WHqjU8me7CYEzVFxPV8Rjm+ZToiZ0S8JMrx0U2PGCEGcPu0jY7H+IuI+T+MI58Ou1K2s4Ew4ip
7okJBegKNrEvgRMg+ojwM0bf3ALVX7t7bEJwgkqKq52fb5ZwVlUju3vgeCYf2yKsY8Dr9PiEGLBm
cOA6446sSPISn8pxU5OShQ5/wUkjN4cg/G6WNv87QV9Ck93b8Ub3qf/9e7p2I61S5AwWTOuYktzf
8kcOSi6T8nfEyDEi6qkH39g9Iw+2OFyhQgJtk0af/oTir3ups6m5I+96VENPgWP8Z5z8LSq6880x
TZYIf6SPd8nx8MSaXz2a5EqOV2bdcuuJcBype2frfGSe3i/1c1Kkjeu7/bFpKkiB63oePmBEpzbq
0IAvnV3R0JOxtPyt+dLtkXKuRF35LHA1Gce1XE8Gm58knFMyRnwrsdlcW3/3veIYMmIeJYR+5SXU
lpzE7AMag64utw87N0xacEOjlAzRicj99IyAz2CLpejyf5wG11zPNj2doZ4BfxOW5aL0OejCl6NL
69qJIrQ/ThrvJNRWayV+mOJXBbH8jq/6pBYkRIVWgXKxaj7za79Z8wfi9j02R1MWQkk3rV8tQeUD
hRKU5AqwkuJaI+nM9LVMJn7SYm/F7BhLEE8Vi0I/NY0QqGcDegtDXggaZ/EQmuCPQXn+GanorOxm
OiWoFu/Ylfgv+LogWUnjrCD9863k/+6mcu3FXSpzdBkMzGkcrlG9IpdMLJtChZhWgR9WPsdWVD7d
XtHV3byin/6QDApt5CjycdJ+TU6190hK+DAsCW6pJ9/PVdpCOgkpz7VkjE1aKg7EDzcBtsYc+vLH
NPktSfItsEPTEgeVRIt57VDqzYlGvRQtbbH5ULz4DTeQrqwcfthv6aLj35PJHTrQUXzzbSWYyzTj
yZ+ptnfbYnm/CYfY+oDMszU2knMxWg0V21BiU3ec6cQkaQwNsuj+lMvOsp+Gl/SbqGhGWy4jDnA4
3dRAsg/la27bjvs9KNUrfWHBaiUK22FXprb07g/qtRq3Y1aMGU5UgkCEypaE8o2f/uNHNyYbhuKY
a7ysF5teRkQrq3qWS6HFK9buloqSdxus05mTuvQjxgs1qOAayE7H6mhW8Jsq+8E5ZRCGCDwk4YnO
Xy+Eey6sv7eMTIJLjTyXpZuO1e4mzhNE+KVhgLGVSWz5/Q0UGknBSPgt5VYWec+xFzALj0mjKz1D
3kWbS7Fqc7HdgFetjzoNYLKy/1ortXX3jmUnSaTbsSWQi3oR2j/j312sNuSYxCH4yehsjwOyym2a
soul5v1s67Glbs+aGaZvTqY0HgVybF+2yDC34o1FSbFO/7cPrh7ymBwpH5ywypB4QUvZJJjAtYgG
asUD8DCLVzWtRqvQ3kYedE4AkXEwqzywJOAUFYKPnqZp+1zDwNOp+C7aDvuArcqN8WyJ2M7LMZYA
MAFR4zvMV5e1r9lWT75+Va2jaAf2m4Oa/vrTSKSteOv01Sdi2eIo444AEeR/QcsGqAG5BcfAo0V8
SO9bZQYm2TDEOTGl4SBi+nev9Y6vzqs/DW44McQtb81Ksw55fayKQZwkxCwySDH52g8lohmN2Mer
R9vGcfm1wIOpsEfleW/aNS1vzOSK37260B4URyVWU0rSPCxbj77thvoOCkZOge4D+eMZE6vzRR68
c1mdAHEiqwqYhboWZ6XeIYQ0fK41qR0ymushw53NlNZJe8FKayirdVcrnhHGq1pwfSQVYPG9yh2y
uHfuKlw8dVzO2dKj5XZfe7IiX+cdLOmOO3jbQcZWeYrjzDs7fLGmxbmf2/FobZe8KyJj69FTVQF7
vBeuJWl0uOWq51kn8lN7Aehxlc7+Y0THgcskduzyMf6MEuwqR7nkWcuP6XIj6Dzi75dcHJCfe40h
WjzNclu3MEanz6vDCRy8JaAJjOm6cIy8LvVmFTCrUqmh3t4Ph1WHwuYtJLCZUu8vMfyTjc3VITwk
aoDkp5hVuJA6NesDkjOcPVmU1LEM3gQ1xqvLRIWqNRcrfKr9yZZCu2RNWRjzSl8IsPmreLHJePQi
7YRaycQwQvwOuv38CYQSSz7kFkkafmdHOidtcfNjNJ/roG48FEh0385Y18NOK3TCj3yY2tpgspYO
5toqEUqM5NijAUHIzpj0fUDbnVVV7nczPG30iGd1UyzcdLLOr8s/m+yDBpLqfkDps8WcY5+IKHHa
yz7laRAiq/SucAh5RCeflr6JoDgJKWLQhU8M5xNlPT93lwL5mBrZetvGWTS4sa9apeias6PPuRFz
40Eb3vsTOI2SAjDsL3MwuwcAXZWTmv5b5057sM7TD8LIK7CNK8AMhK4GnvteFc1vCmI5lstIA40v
mRhQZVkvkmgxUp3g+ZOAeuYjoaSp5TRfe9VrfQgOBS8KqBkvrhiUaRmTd3P9Vtw3fdbeoDxmRzs2
yNnGo0+Nq6SjF18o1L9ktVxXC0hq/5E8QFzO3fnLFUEqGA8rLZgQmlNM2Nq/97XX+DJZXeYp4/N8
rEIqehC+udwIeedsd3zboVlp3zLPkBwHcO4fmbMOIcoc1sXKZNZqTBvvu0c6FOEXMvB9I6LvPTij
pq1o7ZYqTUQdgSLu0Zv+mZAe0R60m5VpnAI+vmJ0oT31+NLBqYxthpnoaT8L54k4lMLUVlZ4Sio8
dgO4q/mjJjF7AgWoevLB+YQgUvtrg+y3YxdmrR330oZKp+7F4agiYUnTrCp1Y/VkJQmTY2EBQUWf
/ktGXZFPSPvwZ4ZF7DXrSGhqA8zCypjdhqgpp1M9jbDaC44tibcG3v872wFrL2LBiPzBskFK2VWR
rIEiXYzTuiXnIkdTs6TuHK0957WTM9gnWqiC+miC+wod+tkD3tcWEjLIXX1RPAEEp5L/i9s22rMX
HUP0m+cfSum2ifcLTirh+7opj+5GJ0Xz5NOXVUMhgBFtWE8AwtB62a3oJXGWpjcAMz5GJ5OaYKW/
N7EDdmHhZw8yRaVcF9PqgOAm8dBViefVHuxH9Y+je9usLEKHoKsAkwkaVsttia9MIUHXg+v5bkn2
ycHN9H+CSXm+hnmGkIoJD+dBRZU4wmldG+j2yPzILLFdj1ace7gyf9ydq4FeH+WapuX9oxrRQElt
694NLSqGdvZHr0Gdwg8hn7ozxQ0bVtxpBVcVCwTttwQj4eV1RBDusBpHIkQNuNMDmQvSgDSxlFi1
gEIqm6sN4QWuHGEdkh+9dqC9hOp0HkEyZcLA4w68eznc2q8lhZQ4oygUl3XtPKDKy8gYhOwH/4PV
5Ji2YX1JY7ZXeQFnjSK4Y8RHUqzaihgI9G60l9NZpBnJcSxh6RD2dJdHaTLrN5AXsnGGqpkCz1x+
T6D3HxQ3w0J+wNPU0AZAC9fJM9qA0DI2VVoS9U07g0GP0bmuWVGtQdhEoqkyH8bqN52cb0XBN3BC
lM+GwNzTGdwzfZO9bvOy65SWhoPOumoBuAW7qnw2y1x/apH35vgccdt9S+OrBu6UW9OJDkDdwjNX
5bpaHWefCiVh3EJaUN+BEUuI1CU99QGjaLrNxTVKL4gVQOJ4P8/zvZMY3wad6rNTYTxU6NWBO4iF
aY/VBG9F7mzvS6mGjGzTseeKJCVERtcJURgS9FF3DJeXsBKakeU1eQRiTiO8O6yeij6xuRJqAD29
IdOSXChBdwHni9jhRA5w97B3840amlLsg7eZI+8HQqcoEKo7QHCCS1VtmKmau6duyAGT2H5WgumX
mj99LEUzhnC0S483G/9U1gVoA0d0Xi1Pr8PRQI/lQA9RPgqgExcmfwgvRtcWGykL5EhgAAH4YVWc
baAVQoF4Ad2f/LdfjA71cqB87ZAuvk3XLuo9mBwdfYO8rcP9XCUL81Pu3HjbyRBA+BQK/8h2wh6D
W7cQvbQVQuH2AX9eFzxmVAtapeE9OZzRe1mKauGtQ+m3y7RYm0IXxyrOhe567nBCr6qAn9CkAkuD
drqZu6quIq+Mfh6LZ0sa9g43afBJAfyyOiyABX5lOA8aRGv11liouk8+w8IsaOGYyLf7N560/H9A
jMc75jzDU3my3TzsgUF6C4nsS/RXKQF1iXqyoRD6G4qgzcvMhnUGvjR6QxHqHP61N8CKlID4D1hj
ZRGyrxRWtVsQCoLALqtFlzA3v54zEylXVQRJgvNgl9piKDbsHA1jvyYbnVsK6XutY3qh5KEwupRN
V+jE8u+nFg6/lnM70qQRIPVhhHv710WRCdDe9ng17QXjaesIJ9MqRN3OTslSBYsJcjZ+TTHerMm+
ZjOorGyAquGd0XTr7Nt/Aq0rfTzq9DyJIMWHEfxev+MNAWTkONT8kyzpYbHTFPQJyux9lzs7OlIF
i6/itTwPYPnXGgZA5ET2JLBK/7pXjjtOwPrsIWQkAdaAm30sZJ05qr6gzHd72IocVjGbGD2FdNxX
IcbxzOO1Bxo18wafVQuc/NU0l3F3NfQ4cWMsBiEEXWh8ZDjznTsH5PQRNJ4RgkyoIhmBkRd8K4vk
bcxmHfm9numGltUpm1lb9LCyTcWKA00HZkbauqEFDpRWsFQp9rmV2Oq+qjGYLBztgS2HeAw1FoUW
m8xN56FgTDu8P9RL0X2jqWfsFdjKNNc5iIlr8VITrI88lkWE3Gf32/wjaz+LdwLylQGfgnLpTz0j
l2HVidJgvqO1XoYv9bZTmPoO/kA/kMrIhedZsloMQEUYwPcVhMvQxqUWsVjyPaRBZPIvsdg/UzIQ
DSI1WKx5XxSzK+TFeV9/Br2avg3vCx4LDA03vpbr4/jVfQRPnSFqfRnVS/cmfiSeteuxvTBdI9z+
fBqCnMNNQg+ZoOr0MYD1TrQ3ExAqVry9MqqSsvYj8PdUtC52EwzkCcYh2E2aBMLjOwpFi6QWollo
zLWf8EY6S9sAdoZHYnQfeHLCdebmHUlZonBBiq92esUvgth+hBZaFVbj4BcPqX1bH5n+rpJISZqv
XGQ0jXlq47BpmUp/5YWfdJag4E93U0k7I9zF6/gt10nX1+38Be02jWPRHoSq1o5PWC3TVeJP+mbB
plhpS4qhGCuHQjJDm6p0ghh+LsomEIYGmHshwOsqZLj/rlElFxfPd4ZKnyVvWIPxKC4NXYf89y4m
5N4pDQriGUtNh5af11XABGhJd5seGmb5A/H8MfgZFpb7orYv49IM51GFiFrFBg+N0dd03gypaj+H
ZdNkY6TU0kDojoNxRI0Y9sCAoEpF4swHJC1yx8Pi9mogKmoPCBGYqJGmBaKN69Lfz+YS5dNWfWO3
SG5S0i9tBj8ee3gvLjz9W/rSJjzhJelJ5G7V10GKrD1rTzXG4Vb1W2pVCb9FHOHfAnLTkfyGivGI
ofTIPEUhVWlT5UqPdKvFy5+3F2niu8MYS3RrUoiEBJUhxKuEVOdRxR+RbG5u4OaNEKNR/9Qcj2tB
WYcz2L2gm9BoiWqxFuG8304V1NjxeWoGNgn+uLWbs+nWdMIHXxqcE5H7y+AX4whEFczKmghJjXWp
o0bb12VQZiAiLh8xyYhD1oGuLXFnxt5AWORZvaxDOo+CIAqsYCRLCZ3iKQl50jI3U3cBA3Dmh3+E
7XkKvaP6wT89uqKrkkwwYMYOFXeMsv8fAZQf2J9cr1rhn4k3rE/9Kyn09NDru52jp1EetsQYc5NF
em8IjqCnGSjvfFy18/cCvDbbGNWlfB/Ds7Qu9RdP+vfTe3428vTOtMgdsw/09TqrwHVZzi32mogP
l2anS6VsX0CDCwEI+zA2tc5syVW+rsQxcsYfeYgyB68rkGnYo3JT8mJXGpw65LjS414bMGXvUs6l
CaD1ZW1FRYtm6xZ/XG0LoOw8NhUfkr6XvLXxLsWt8oImucvfN6+TEd6a0nfCClbhIzJwInBYC8iv
vf45+JIKswOPsRvffzE6HGgPIVcPARfU76Z/XbiumCFqr9M01KJce3zrHkLF16gM6ei4rLQKzqlK
z/dV5vNob4UULeuOAMK0mspmIABlwCbKwWCHfq8bqQwXAGQaBh3gSlJrMyRLmof02VSr3Jddwvt/
VuS/XBJSxBG+/EHA0ysrNaW2X+1i+nvqZCpKPaxBG1kp5cQp2RoMR9fnogUU1trjTul61naWoTgp
UL5qofKVHX21mBp3OIf+8iCt5nE+6T0zT9pRkqx1IxEazrwFqe1nybOhkYA6fR0dcVQCw+ABkzab
bhfi9sq7m+vIHhtF9/NjD1MwZ05XZBImRMvhFNHDyZPQqTIN3s1mZBT9w4K1nvcqU5mo/9C0b8ov
ZAlRlcl/QZvoozwqx3B49VXfwAq+Id5Ltsxg0Pgvc6hUHuTMJDhEz8exyoRySSHEnYLZukDJurNb
10KSr/Kqr8fPZr4okD8K5MKVtc9ThoxhBl4dX0JRSusb6z+vPlUKUg5C3eXNH8aA6v7Q2i7o2pkM
bOHoTbDqWNE2F6A+h3b5gIeA8mZHjzuzJ1/Alf2H5ajsmoUkO6tycEoc8uEzUMeLeMIMyHbfiD3i
DssrfJ+f7OzZlaeEztRTbqJu2L5Az8DOe47xkNuxd2oUuqehRG0LculTZhJM5wvuCSIUjmsrnX9H
WK7e5NnuW4diGwb2vjTxXo+C8LKehBTVwcavwD5i3UxW2CJWBxlm1K4OvJPNJcTZaw11uWvVGviu
vkKHP9lp4D54a2PU+m2Bobw6K2WTCgZ7abFB47KGZsA5RM4ATYiCzPyYNaMw1vmj5fBvJqL5W6ki
V+3xKTMh0wnbR4EpwdbgthpZ9pbA4Dw0g6jzh/+rGaZj2zrY7qXi5QiOS6kZkF3SjVYUCT+/SF4N
yTpxDW7bfD3P7UK0Gfrb1Nsug7KUOpHMhZHAVwjQrapPoqwRDeFa+4wdcjbu7FpZmYpqxQDEwoGV
m1tYEvAVkwNDqlWQCPVKg5vb+y+h2gv5zzQ98cXcp5yMUaST4aza6oEEwO5AgvEpzUzbtDXIxEv3
lhK4Fe/TvHBuJ5VT4ikPeSJ3J3WBgUaUUC5D3ToV2gyrA1BuGgHUXCGUtHZzVA51gLHlqzC3ywuR
e1eSrj6Z8FDjTfa4eHC1ER2So/UPFciBn1LiioO9+xU2/1s//1ic/ZV9nWBsm0i/10ELnuHFyEZV
QjKDYEyYt0nHFCfwUszMkrEi3xZ4WlJGWVWPRfZJnPwpcplkyst34priJqIBrBE12uAhAabHu6M5
eFGEA39FuhkE9hzhCCnYahfHB80OzxPN0FqyiRl+7qrUkr8YnZE8JthHDtP1nYQVXA7vOT7y9Wuu
YNqHagEkz/AF3Naz5kOcprh0Tym+BG1Y9r3ky+TgGrKzv6rW5kb0KSn+8h4lQbwUyBN4iQYyTc00
MOEbQDFwNUBpbpOvDOyfa8QJHygQSzfLaztLL2g19+pawSRYEGCT8t6+7pF5x1Ns4H/VeujWkT4J
ylf7IkFURoVQwbDVBuBCqXcGb5xQwhDnyiFxJXTUM8iXoF6qb+HOrCYjzdszt8JC8e3677tITExA
SGZ0QP1y75qJSUrjcUzH4wIYn1/KsxuRqD4WMJaJzSqCPRRKEwFgM2anIePVduB5yQnkpdcpMaUU
h3UvFIv2dYZtM5gP/04gCR/ckThH+0sIO2De42W9tKXZrPn8iwJ4/zxdkfI6ZXZ/EvJoatRduldW
RjwKazQfqeCs7tdPBOVklJM1K7YhC6nN2KthpnHcWF4QzcDqSHy+bKZLLNyWWt1cNfeq4YLd+DSK
de45SgINua37vuWmWKCtPj5JCGGdnf/Gmh5B8i5idbPvnGRmijMsWgI8cy386tfjj6tvkSb++qKG
aJbFBP1ZFfLPTy++BI2FU5PV6V8s2ay18MWvMzhlWHqSrn27u5qEMbrnu4L8y6Zfr38+wPYZ0OqL
Xx/HLsVHSW4T41iu2uOQ/JxtVCrpvsjxJb1xHmKcs/3/FA9UHOieQMMKyOaOjdcdjQ0ImvPAniXi
F4l+BIxHrFUq8/pNoJ3O6JVXfZFRfRcT63501glfkGIxXbkZuFoB1lMRS/tz9GCjmwaOISBDUiN/
JlEeDlejTM7pWeqL/pyJPGWnpTZDkNkU5HCcpWzTJ4Ksm+4Zt5BcHlMt6cNP+9mhszgDyP0r71Oa
EIKe82dl4x1Q3bhKoMVbiLeo7sWh1Sx9AguNQ1xjGth8sTVxc6fQFBC9ty9V1zLMnH4crRHKpaCT
ti5rTDv1KfyjlP+Fus5bQS795oVtGpNapmVmvd6gzuGAAX747HSxKNMVczybjMj1sEsI2AAIbezV
GNmTwglQIz20XHjyUaJJoj7Ka9eyZnHytbxUBBlF2D/c6HkViEUegVyMb1TI7UgxkkpQU5nayACj
PCmB12uOO/GWs0OCb9if6ExGCy6ydCD3YwGRifURQzJbDaWcMb3sNN/54ioVc640J5STQXPGpOh6
+6Kvvkjrucx9hNYHYyxq6HumC5TnWYHGicgYgANv1PG2wbyBI0I0V7XzhizdAmSjbA4PepM2o3yd
E+XVwCceVirQWpAxAMNLmzHegCPEI51op3qnmVfqwrzJImB4Imq7ClX2ALOrTPNR8Dz8fO/j7kgd
H4TqDfIKCbDqRwmtt6d4URL/rGH8Eas+AafCsm137kZuTt5/aMigCIjC03pZYIyXEmj2OaqLdSVg
Fc+orNPVuN5dnkm4U58lG6UxpNi8AyS8gtQ2bl7p6HkebDjj7/TBf2dezj+zgiQtr19NCRug41bX
wfrO8EUI+znuaBHeu2/1MWKMhK1f3aMTSTZPHt7CG4iU58Vsb+iA2157zc6Cac6FOG/HxqZaSiVN
fECt/+oL0ZFaLVCUEiq8zAICSuutX5EqRgR7OhJrZxGe6mB0wMsUzNAaJXhBH8ieIvqwSvLbvSWF
O/M1kbDeokkY4IqUxVcY889GEu+lkEmCDIbCoJvob2xtExUU7VZBLCspRsSI48D+Z/2ShhR76vTk
BuP9ucz/zPYAQMueoIRZe0JvNYzKJCXzwTGhCke0wK+Xdq66iPlmkQ9inMi9fNFVaZBylmf6eves
fmg67A6pKhUD3aDilzLU0JKrJfgwbMyTumL/qRmyRXEaCn6Lfjp1fsln96Y/FsHm0KQpqh+H88LQ
iRfEOYwXlnHJdstLeukv2xxQRKBWj0D5Wr4IrPQCRhSYGHGFYVcgcFEhAm1a3pFe+B8RV8yPs0AZ
0FWleYnCtKBh8fQAvGees5x/4f4lR51urSQrPF8ctl2zXjSIQHRXvJp0HaNFx5+p7kR81QaZS2qm
NN0IGlo29p1/M54siagSNS8ODLjKEI+R4H26VtzcO+RBkHsbQ6gwqDZ/zm2R5kQHeocXPrxIu17F
zz7CMILuzd6NgVcqWjwXsStXJg9w2GxB4XsvwP+eOEBulw+4WPBqMmqTxaX+9CspYROu0orySkuX
Eu2OiC7vNZ30yfZF4+FJxgzM4x+aVBh+0pUAkQ/d42MmtByka/kw3si7ioNiqlGXFn6W6vUgZLGZ
g6i/KZZs1L94MOQo/tVvl1j6zNfEvo6r0E+1AyvSvN/r8MFkNWF5dUxY4r1e3O4eSHdldyQXawJG
+NXdbu6cB6IK+dIkUNwprV/YfEISljafQu8QIxb1gpUh3ksVeK8uHse7nQkyOWgXH819/mgmCEwS
Pjp1LQs7aBd30/CtczMDk9feauyUGm8d57d7Oon4fq+UylJvn+vS8uwhpYon2zR44S6ZeIgcqsLl
AkbsThe5ErZ9A5u8nxjUvgkgB0OKX7+uBPOhOH8xXR+cwc4D/wkjMSyoBWZ27pgFiqO3ny95Irkd
UEZuNy/vwlopKs0IXml7VRgk1i3sEmFxfM56Lg1VYgzeW5RH3XgHVnmn9AD1zSUz4KK/wOYDNH3h
FqcexS1eAngZJG66rsm9XWO0naI2QRBaKpPNFPBbi7E6gzGE8geo927ZhWGuiEqCbUf9dIjdlPpA
1GJZyCj0YNttsJ9gKBMpWT1Qro2zwKGOgfMxUB69g0yck1WUQkE5f7om21F3LUBeokrgHvA5r/n4
5DxxlqvFV6zJi4K+JpCv7apd2QUJHZT1ctSZfrQbcpmBaAg7L8kxOiMlMvw+t9lHINjo0h5/rVtV
PpZOYGw1t/k5lerL7n47Q5S5mbANVppGzogYE+t9F8yl25Vut/JWnYyLn/ONncPOIcADjtizO+uT
56QZr2RBuqGy+JTsAKok2RSUNCNbJ0VCaWZXrMRR6HOBhTpLmhudaqUBwLsXtIwhHqP11I5LQOCv
G313ARi1me7xNrMlXuX+s69LmuBUXFaJ65GJXUZ4+9tNWaaXzTKHgH4yZid5V46WyTtec4DiH1Jf
vLZ9ebXxY0R8VGw8jlxwe0JbvEZ4jSYd67chGinycAV18aWM6sejieQ8j10A/4ggFovANST9lMkY
+FNqbQHuXxmHWyrE59RPrOyW44n2+lnbDpG/DDD3CNm7F5DaMdAWDvwl13/28GmqIvW86B57r8Cq
+fbmIqa3vI1cgeMO38vykU1EkLOhdYHmy+v1jypmJLEQSiPZmOu2g0euwuIKot+fiyQddYyLGAAx
MSW7GCmCccDlB+PrSdODZSEWMfVcWP0epswCLrScw7liWyB5qvgJNeZ1sN23VbVNBqCFCJ3OQ0//
mMfRp6bD3kjP6G+4ujxf3aFiwJgC9VaEbOJ4Ygl2uxx5u/scZwPVW4dC5WzuhloA3lao6PQIVJCZ
+91bvHGJZW9pC998Mp2vN+TqWdGHKtz+6AMLs7w1ffa2axSBJSxkQCerncg+vDyXai1dhhx1DMee
c+/QrloByBpGvnV+EGko+v45/N/6fFIRUOh+IQIsDcFdt3B9zp70zOJ3+F5UNeA0RHmT5INqdGic
sMrOIbqGvdh28ynFx36RiCWJHr+mxiMaah7baEoj50IPRF8194wrHI9l7UnezTbHySGBKRQOG8Rw
dNQpXocJ51ZtF9qiDUY+n1Cit/zXLCW6v1Pb8qSKxk9DQxKn3TRfiN448xwX7tYvxQh658V0NgX7
0+UXsK4Z2l7GK6JV6mkJ24uZIUQuCvvNz3luZnqnjSnYUd8Hxcx6+Ix0EJMCHl7CAvUsmDwduZAU
WLe0MQxU+YAOY6GMmvQ/H8X2m34q1hPGMAC7wMsB3FFVnwW7khdez6Xa+/cKxa1Lq1yt4cH0GcZR
6PFR5JAvPV3+tdcf83g2+9y4zPcfjddVvglz9HqvSf9U6Q7TaOCZ4UgJwqK5BJv7dXquZ6VM7pb0
l8xctBbfK5TzrJGhribr6zXhS5c3WQUKilFN/Dw8Pjpay7UFPgrp1kB2StnrwSdeAxjzLuwvupzR
gJGokB2HPcPlARv5VZeH7NoXuBxaYuF4LJkEVrugJzJhnNFoDF8C27+0bqH6C1hq1b2eGuheThK4
TNp4XL/1aEj3LXg1JdzyR3dYI001vRW0HIMEedCG3vjyzpKYEwSPxW7CxIZ30B1u64KXeG5vvuEn
7SpMBay79O/+L4CRfvWn0lQBFFnrKMwxedYP6Xz9NuHq9izAABQR1ap9x2cAzbJa/eJKx45KMYnz
Yez2YAKCCEXcKhl4k0OIK+VnsKswglvKuBNAFDOJizO9lWKe6T8R4+sH/APHSw6PkY5EYWUivOBA
6F9oEv9yKK23iq+OE232KhEA7bRSQYlR/2Tu2HHtUx28Dty6uXWN+xsyyI5qR+0WuzDF8zgtqEHs
vaTwNgz4yw2Of5r81R92Wc6KKtdsqpK5Cm67jHRkeOZ1MQRPo/E7Gq1sS/qpzZ8/62gIZgAy9E9D
oKViXuScZodmh1EzHRTmy8gcNy/xdHH95yMWUgV7cdChP3IfX3qoeZ8lAu3Kw8sQqR1zeI74AFpZ
3x7ieR0JZUbWVW4iywKv0pajpvDEtYqf19nuAFjscwSEWIYLHu6dVcvIlp37tMGTFf6Kca6xx/HA
qmSQ/duGcB1A1gpBdmlP5p5zAYDmcFZfsJF3Z4y/g5RrE2TDxhBsu/1oLpM2j/LxzTuHjK2jZhpw
wF6VgZExCxSqHEQXpWInNP5UdlUZUkLDhKqbsnN6c2IkEObKMwGb9gqMKDakzdoSSVXAiahmfzxH
r0Makx1CgQB5fGU6EEgJKGb/3zQTqKZSu9HNifO/cF2vYYv23cg/Jzyky5AsXHFPSsOfWGr6XLKZ
6r1Otj8n74Om5lLWDBYjfxYHC2o/DZhvo/7OWKZ1KKh+7Br5MHeu60krnkBws7N/wxcJ0Ei7lBLS
EBJ1pTuqUev8dn8j9PdX3eYERKBYUVMje/v5ryesK69YTJqnWg0QUSTbzlHmMdWrLgNZ0M7IXAmq
e2MdjGWpKCXkqVIz1R66eJuU+H2eHsu8kxt5qE/xLg97xCFH6CnWJN5FomQN3VDMY/0yoKOTeA16
+DRxi/0zHhV+lgLbMeE4SBhva/jguuHmFQvFSMUoovabxLTwDk8kLUBfv0rwz/gVw40hbOkXHNlj
V3xAqFAV8yEb72vfwlpjT+smmSECOcyUry+gnWLf2VjKZFp6VR6uiF+Ue7w1B416O2CIh7UoGDz1
KEVZK0NvZj0eKtx1cKZKKmfvldDgyTX0zOqJU/rHW0ZdgVYnXzIIZv9Tc6PGjzT/ncKXSj2uUxJD
aC1l2HuGBXN7Si+ZBw45FLmGw7TimPy66Zl5gHQsWfQ5UkUU5OAJMZrLjT4hERnadjIwOxi9rzQ1
r8RZ0EEo+bwjZBuycyk7yRV/K87lH0QcPLWarm4zDw9+/FVmKnrMxBqi8zFb8y7tnJ1QKSSDFKXA
yC3dSUq7m+n9KS2c5onXLMZ5o9Iv6UN2hhTPQC247NdUsCrkqbAcQW7eUGyHXrK4gd5LGlnUCYui
DPIMNumPz0URAAp71FQrTZ/0nTZOQXnQFDMTk7c07yQialuV386Zm4QRsjM+M+8jryjwGBxnfyTg
IGN3sDJOymdhFVUDdMV4ecBob7rFs7V5DpJ3jbWM2RAJEG90x9rkA5KP4z6YM08XZh6WaEnB5mOH
ZNzo61eBSdNumAB+mUQ+KGXv1vTXZEC6jinaD8j8t2DXWBiCfSe/ukDesntwCkcY2czRZjdMGKyj
9BLr7KVx50HpKEv3Ik9jTMC9kSPRPtIhJUqgNrfND5I0ep+yk5nFP7vxQvskAQBzsi7m8WRjJ8hd
udsHxFpcA8n41oam/5GrO5vLJL5kLDEk4fCOTRL67fkAcCMEdVyeIX07IIaIb98ydHiJkn5nbT4U
GA+cjdBaIWaVUqAZnsQQSpvWmcJDnjxPD1oUYqFtKSBsVSLPhTPxF8L/F6WHmOnsPawGHpZnkXPh
naoN1NMmMD2pvqw5pvhAfZgaG8vO5SnkSXuYxQQJPhMX48LtTgYs7+6d/kem95ChmY7L7CM3Si6L
SFqEKovnXPm4W9b8eeMMiMq/uJbKmxPVVYzQwp0ugOURXn2eVJ+vxF+0JNHIBEb8MTUwmr89Xxo5
wdv5cL1V1EwJOQJAkZ+TT7jS2HA2/CRxyRk7wmgr04pzajIwv89Dpz0IQnNAkAchm+zWUX8Ce9Ba
Agz5q1VIo+B8kMEpmDuvkCED0sHEyDIVgeJWyxWGCeHD8aMKnYr7eXsQgfZ/D5CpXMxHJQdXtaAj
+0FILt41fSQ6i5XrWNtMjNzh6ayUKurFrwFamvVy/jog51vwcyP1Hm60LI0j8GR2S+4JRXHo29/7
bfuW2Eft7WYT/p83KPGEpZUEWnlMfjft/wnuvZ9Pl9g4oZc572S0ru0aWrvxsmRPNBuYbdb7A6nl
Dmiek5aFhoCgoDFcxgLlhE6G3lQiFRzlRE7oC9cL7vYyzvqYqYKmzaqHEUjJDdCscPaFKCDtvOBQ
gxqSBqqypFpD2fsbFWKxWqXvbDERygdIKuDNtoWClcR4WyeCyMVTLEzl12YlfF18QpVDr6HqVlAo
SmgtSJt8qYTemV+KPsfzCpTQD7DiZMQFihuCZTZqiCLZ46dk/FuyYDwsvJT4z1V4xDNGfRaP51Vm
6qW7qw/X1C6+C7hKBcr5qrNSytU6IpEoXPOzBgjYIgZYtg9ETRjd/YCT3hes6llziriinye3rGCH
vsejSgiqdsCIBtSRVjNqRjHLMm8Y8IcviRgPbCmN7HKBWSarF/cObdEdSxNBhbab+NTuzMySTQZE
A8XJE2JcR0EJYKaAfzymVOmi69015yKRqsLaa6oxXIEkwnT+DQi7H29wd7/diDnDXUEdbX/bKRpB
H2IuZCeRItdIiT/aSic1FRNWntP0oFkOfjqIVU9QqRrTZhlI+79V2bUOHZ0nX+616Defcklu5kB+
1RlL1QmSt5wb0TaRUp5L3RB2h36wRnzhDF3pFIWa4lLlmTpYUpwM6YeHGY6CQdTxBxe0SivhHNIP
E0FQ8MkvHKgqowx7Mykf6XOIgD7ux56TWzV5JdV7no29AYKUIYpc9jKaV5PMRMGEdM8EY4Pn3Sy1
PmSzDnwRLci6ebornXPLWJtcarTGuyUK760ZAbi2Yghrytp4KalUpt95ogVclGCVx1KTNKtlQVQr
qbhlmP92DP48OkbZsXvMGtrHaNeShBLgo4cLVSOPD+w2LnuvYxuDciLWCANl7LljrFvVcbrIkofi
6mSIGaBCjOJrr/hSeiPC1pNJHAz+C4sEKTaij1R+NOkKxJHrm6YwlttIEgp7f6VC1nzFHRWkqB85
9s7Rg/Q67iZAEjyBlz2aHrimzyW5DhauggUy6ZtEfxxL9l1/AhlVaz6iwiI8xGsqe7dBxXIYQC+L
yw618U1gnsehsOwW6OtVNhS0jeCsW/wzwLU6xlM7nulBvIcBf8PwJQG/0yIvoGBG3VORd8XIVXgc
NmzI2bz5QjEOcfvL+6gzxBhQzkyl8aLKklvsBHnkR+vTSS4tPogFs38pau9W7VsJEptlbblcvzPe
+FtGWGfecAZsjle8NzuXJasU6ShEfZ8SVw1DV5NxQdN80SWSl6oznGg4dJs242s7IJ/7slmg5iVg
NnaEuCMpa+kC07YGdCOh2wDPIetFmUM/hLQ6NYiUEP+BycTt39RnflrzoJwFKDmqnmIxcTF2cNdE
EW4UF1WLDLPNapLSzkKlbNlzr8dLgOXjC2cv3QNY+P8dhL2V7Ppg+WPt8mPZsAPFZk83q2bzfr2j
5fW91Ygaz2No65mMkwwEm/N4zVW5OYE71DChU5q+pfXSKXxhPqm42K3vZ+9ZFRSCNu90vQLH3Pb4
9Ztkpurb49JX8D+4evv7aYb5Dzcy9u0vU7irYi3C6JCoVoRxfWWUsOJj3x07gdSfvtj6mr2JQoo5
6Wuwslxl6qG5OrTzUJu/9nBd1UdB7R5WmIOC8FMGDJKNxCOP1KoSXtbgh/8UDTcdaKQfTvM12MCa
j6Mi2DVhQr02ynADGloqpioZihPqa5mwN7xeQzscvT9z0yEFeM4RB0epliu+XPrm9jY3IYHuLg3d
hvmAVMChQxYe6NHSu8RjGspyWFbzRfR1kXB8AjVfMsDvA2U/Pzh2OyvVjyigc6sduglFyx5BxGW+
63K+Slc4Mw5bPbFkvMd28e+CBZc6NfC3lhgoaAWz4TwbLASFnaBfoVsKDRvCj9BIrDZNPu0XiX4h
3iYqe9OpViWNWegf4M7PQWV5uVuezVqYrt0Pr8icXa8YU25+LVK8Q4i38/0YcgYXC2xB5FS7EFvx
fgMlfM9tuDOcXGmW+DDF9UPOi3bSCcc+SUyzoxB2SGePqn3jJGmCHuVOPBLsVk4r2jF1NP/8Qr8J
8yiYZXKODQk7L5Eeis51nYDZ4G0s5wcDcDVns4E7hLGucjy5dg3v209xzdKsfwIbz3KrQCUSEQrR
vza+TgwoeIIZq44ECHOVuQzDPLbjSjoinKibBpz6dAxf+WXoViSwLQVDXwADluvf9hL4iER4Wgww
n2G3AUkfQXd5OPOO/b6ngpRLMUDekQztw2j4J8nM63GpHD6keGXuBe/vKG6gSNpBmptISzXOxLqU
tJiDrVeqdXUwFd8xHKTugW8ci4WOQu96MDr4dzs4+4QCoqq59CSVLYDfCtWt95oE1v+Ko6vSaquq
1/CztIWNZuBFZscxl9W55XE+XQHMVS0csfZ6v/TTAVKBU9g1upNYUIq5g9pQcn26mwfhaYfwOcds
4uDtmeTedqllwdvIZcDRkdEYuuSmHCXcUVlKgGbj7p8zIm5tjL+wXNb4Bz9p5b7C/fj9JrjJrKTQ
6YD8pjE9ynoMer91pn/jPS6RN0N5kcaG9cr2EsfrAWl/bDqYv8c1Ofp4wCwMOEdXHOzj/1QeoidP
XNYkmCsXsskHbvxnQVNtlYDL5sUIrpnUqc3LWZ354RIO4KeNflp+VNDY7RmmOLEYmuFK6Vwf/0OQ
5EiX58egGtUeSQ5I8xG0LfdQ4VntQEKN05PjASWaEeoyEgoFUJ4yDeIxDu/p5zlrE4DkIx3uGSEA
8XBlLB1SexpkX/PdubxDprGxTMDV944W0RIMIgoqletHeE6uwKM8G3AEQObdr2NnbHtx9HY2S8Qd
AnkWXZo0vCN4PJzcjAOQ4LL+fAV7JP+F1qSTwLMPpXi9UUvOgqJpahCXY6euSwXtbA5x/1huO+N5
AzJHCg+UTEe/6oqeqNP+fAbz/xCzwHd6s4vCDL3i6G8BU19eRyWR2BZ1KDM8283vBGUEjewt6QKJ
Purx6K5Qa1yoDnJ/xino81fcRc0FcQHbbe+UaP6zPrguKNIXB3ls7FyUhXOuNyiUeJkClryQXf1V
uOeG7bwoEiiIySTF054CKMHkR9enbENW7ZfJW7N3dtgEgP14u+THAquSzX/ajAzCspH73H+2Mrp5
jearvBFNeHVisZRfsJtCRuc3ivPth359pRAJsez3i/3iaYfZjN0dJbyRqQ2NZARAFBSeEG9o9Wuj
JNkB4cpThGooj0QRttgbMsg0gUaKp/mhgoeO7ahl/53b77PUSwFvitG2JJmO2I83g5o1BGJG/n9e
fZgSQgFS5WqjaoObIr9tbo5yxUzIoZF1xe5dcRncXrbhHak3pT6RQkzenw2KRkAVFf5eOJVmrCMb
vXblHk7RrtPtFSmGJ98mKQ37mq86rvL1A759Y+WOnE5nfvFn3+EFMWaAKALqE8wG0YLWYNZHWn04
74p44sdtasX+CB7pAKK0PqZA68nPbbfi07I2ANY8ZBSo3eNj6b3J9/jmecVDFGyhaSwKISmm+mn4
BKMtp3Itzw8ZrXhHYVxpw4uSjy4HkoIAGQQuxa4ycuuAI65h68Gs0kFy/fW0psiQInMADf8/kauN
exxLXjVQd+qxrqQVQ8SExO8l6SGMic2/09BgCRiwPrVDNi2AgO75SaC0wodtcKP7jLuyyhTkspQw
u0T8CiflXnEEZX4uhhs8c2i5H4ersNgES2YQPHwCX10Ao3Owah/Q8i+CNQ3pJSs3ad0tTQWFy51k
DhU2949SNI0WKYamnDBVAfi/W3sPKMCIMS5v3ZZFM5ACJghIQOxmzjfJVNxbGLCVH0cenL3vRArf
tZbhH7nPcO9pTU0J07sJN6gUf9N5gzAEM0qGmQZXyaElldIh5Ft5OhNOBat/YS19dx1wQSLgzorw
Xc0iFtsyDPnhkBIzxC17AiBeyFhNBGhU7CfbfkglXj89MMI4YRN4lkP8IAbcZl7JhPq49b4uDkUW
LzAkP8Dk1GmNewU3uWCCAoMlFRCXbBO02MXqpjBgV6aTgtLhtTGRlLbvdUe88KrPsBbKfkZeKEFG
ag7HYjCwyg87qE8H5RFSxY6Jy5SlF/EZMb34M3HsNspH6fgBfcSxLOwmzCIJJNJkARd0qaozDf9j
eZXT5ujWgU2ypYb1QhlWshPpGUARuzGRqJgFj1cstH8N7DeIyGu88+8p7Oif0srai+LOJ+JOkpiQ
1+LifPeWOzVFXoG+dAklwpTr9NfSc/pOU9cF8ema2hbm+2GGlmeuoydkgkMlow9IKCRlqG8WgUlV
9jtecYrIwieNSkQOYRdu+C9eezFtQSlaKBbszaAToVaeufROAeHKMLxiWLIl/WnthpCVbBv/Y6i1
5+MJcPr7ekElKqvByRbK9ZNrtCayoyQ4T0qcW0N3xLd+nUDOtBNK1DN/ndWszX7nnHKEIRrKdbEO
1ayRNPrfFqmqci44tO7yRyrGxs7aJMFk1mnBQGpa5BbUMUWN1XrWBUjTpRDlXFqJrIHzPNvcoPWN
8tzhlYsrTuoXr0oyBjYFOXtu/Tig4KvwwdzxRNkg0W0kjR855+I698Ywu9j323QZBFuchyRk6jYa
ABK2hdvsoOXSQCsoSe/+cD2rD+52Szy899Y6zRzrBMZqbLZG8rXT9LsIBExD9XmVphanDFZAIixi
hzlI21Tlba/rLZP51GBJ1oWnK6H4X9e6Ud3h1W+7W8yY0aiDjLP+uLqXoF6ySK8j5K7d++YWjLVf
RUlUtVfnzsdGMAKwdQyM23sOsK3ISzLPtp6FuYi2kkdiEPish3gmyp5t0Va6mnZi8gLgBF8jPoOG
cK85+Rx0vwJUZ7lJN2lNZvCEl3bIG0xhTVGa+bLzxDu7MFwS7vD2GIMK3CJGnvb2PR2N+0kEPiKr
66BLKYVw4Hx4EqKIYzMFZN7LMHx2JvgxurVqM94pSqG1VDivVavHrimG/KDLlnXXLh3RBLtUIk0O
J6IHgLyygSlgpxixrJAH5c17jKS1hFUdjM043NeqUGaleMzFs6TzgAF9tFpO09IDgoC4TqEY1ktN
ALcI8HxQPebVbLX7rVtocOxv3ihgWZjmyIAM6mC+oVOdJI4Fc2QAFd/Vv9aCbOkT+XmXTFDk5qtY
/ziK2NFy/pwzm0+W9V4sT+XjRTXJaQOcTTCgooKK36I3kFRfUodANkheIhN/Dg0FDos1xugtTYZd
LkPJAFwHCrKTzky3uzyc4RXaFpQmXAg7TQtPc4VJ7WjgIf76RVWKtMLpHP3P8mWTNrggqfWVEsKt
hZwdoh/Gwp0M0gtWaxXgfxjHQ6KktoiyEnMvHpesnwJ10oJOnBEWw19PncMuVcReJaUaBkGs/hWE
JsQb8wZDmlaE7Bd8cdRKmOokwtcLNuRsmCx6n4NUNQEeAfsm5xXLlRkVqFI1UNV8pOv9BdYBPPsY
UVbthw+dxsWBm4oDk20yy1qzs9qfKGHkVDc1zSeW5yPAVEd/HkKHaoj7YCBw0vi8ETpF2yGxB0UJ
umXeUgzYQisln0CF/z2aOXfW/3/d6epHTxkiuOV3ZKCOhoeCohFVm5xYsiL8HcHH0DibG5hYBIM5
FGeZIK6/X4eHsS4SS7WJY5iX+rn6pkidvnxcImfsF++r8qHafOMznSWocWOmLZxhaHFXfCfRap1H
bE8eMA4lFc5bf4XbJfN/qLKDemEYW2M2L3UxLQsQkpxggKcDyHozoiCorMisypD3e6CRiB9tjV+c
toV8ugGSC4H8ha1Va+bSL2NTnxWpkj5mmSvHCOxTB9x4/Ta5k4VpV0weNuaJHe2RlKcDBQiDY2C2
Pbtv0tsxUcJySka2TFFrvAVEQkEMD1RrirpBCpLyBoJYgSXhJ88X1RBBqhPlQYZRIYUXO8+t2qX3
2K/N+otyeqtPBVYbqDdctr4vwaqPWMY/eqgGXHN80segsJ7DXAlX6LFWMB2QHqndYyuI2cDBGZkN
cP2cgqNaN80hlBtANkJHIlF4U/QUy+2ad0308wtFwJvyzW1BkXoo04LYdeMljdqb/HLqjWV7HKiI
zE8B2Pbk3DVfAHi+/viqqlejyJ0swYomkj95edGwOJ+1gDG2/iy0BLs4Xawwznp2p74C8s0lle7f
FNhQT/h9wFaIE44tSaSeWvGyPMb39GnjNTiwsKuWBPZD669IsWFoBAdv9WrfSkYaAhOafpc8Bd5n
MFfpP3vXYXpsr1KjXLyyzOyt7YT56OWi/s7ff9v1rXtroA5XAqrof6Trli05QrOPdBnQG5lLp0Y4
ekSeasNiqIx/FW8LD1Hyxfqz94Dk5idBkGQbbgisyMC5HOVJGDaF6ICavTc7vR00Mbk7jnx5mXSA
2mdDk14EmeotcNwE4+4Q4Kr5fr1JRfQjffrI/KnbEg5nGtLVsHsssLNQ//49Drz91O0hyOb0cbKZ
0vp3l6YLbOfbE4t+7xPxm3/eS2N+eIk3Ekm4y8LK9XyfX+iklyBm8X/2iaIEzSjJb+hFDxZW2QHf
I5XEeaCFmaLXvBzy/cOkYXjH5QoGkU9t4PLtBggFpZIY9ngVVhjy+pZN8f9gD1HoKAWip1DPoAlE
pWjYc4ECDwVd93v13sj9SHsiFbvpqh3Z/ZGun+ss8/RyXk1Mxh9CUaJcEiZdu2DeRMC5tQEiOWK+
8lLp6UX4+3O0ZHLj+xcXicrXYxafTNUA6/SVGRPSGoZJzvG/wv7DxQRTqJAtgQfRjbJCYzIkYuD8
InCpWV8T45btP64UDBac/WOmoabUYZYWZz7s5Up5RXyw0V0cj9/3xNF4/WmhYMf/35AhjRTWS1nC
qTaNxilnKUoN35CkGjkKmcjYJumnyqYaz8ao/g1ZI+JueHhoSqfYSahGUIF/raeFFhqpQm8Ch0q+
iVjJtlPRJYCoShd1+65cyeZbhwiMeXLuzeQE79qFCjMQ6MEOYEy/QaQkxp+3MLdmj8mZiO60N019
sgtvCMFS4xyJGU9pqSHe7z9WhSkAGmgpF5fXVl8HNkXdI/bElk5OoO8wyVi59nxX3FAiZypWrtV0
okC3SnnArYYwZHvfiWLanKaj7Pg7H5t+bXUmJND+p3t0pSN0N90m9UkNsYOkpbEJuM/GCU2tpGsL
h3jVmJ809ATpuscj7DpRt9JL2TYbJRW4I8UioDogyB+/I7iWzAWwivu05+pd+EV2WTqCvcPmN3Fs
IumvxGpY1YDQ0Co1B3moDhmPgHcNViAWsLJpmjA1ueklRxoiCS4aHieuPc1YtFRaTD/UqO+jRqRI
0J0Ew6CIdYAseRek0fQKTnmFGmPdbVmT5aTUvtigl6GWgMmAjBdjEZNEvSiJBXr0d5HF1uJxa0Ph
j1rezvoOxKq1Vx8cQ4O7W6pgdylPyM/J9qYx2QyQFzBjbbKNcXnSNO3S31dFJfmwovw4HCs7RkRL
5nBIWw4HNblU5OG1VpOy69Kt8L5kE0FDoVSxGFEb/w+tti+N2sNh+NxMP1dTi+Y6smI/Q9OVpqTE
9FpTmNN2V3ofTJ6QjF/dKPRLqwP8+KIXy3NKndNVHZ75DuDPTrVlPJgacGFVvCjFQCPXKqB7SkcX
h8YeIOMnOpEGHCY1/HQOvCjZ++T7nm11kxd+cJ2GZpqvxQ5J0lb60hkIa1s9VEMMUZIRtGj0wHpo
0qnzSqZqvWMHeMxxf5lDXWqx82alIR/uaZPo9X8/btrD91Kl9BAOpi0hG4m5GvXqXSAaX8kxtg6i
HBf263p26HVKj3ru7ErPcwOw41ofTGwM0hlyakP9BABZWFDfgk2dGZUe2BThWFsr1F3+KSY/vR9M
l4J9cKhnMzI6Qry0S+eWoOMPp5nhucxKy/Z9en8bUydJZMOlWywvKswYy/Adx44VB83yhKLnMwru
6AT5DIEfR+dRk+bAMKSwQrtvvTJX9MUnNiQAEH+mcMIAQ6jPIaRfN3/A3skAYkpGwDktMYSQHA++
4ryllyKCOq9wrbr60atMCFd7d+9jObMRRHZfnoCM/0MSgV6FGFhL3t2GWYOS+ktcKXnk7Lkqxx6y
ArcYxAF8P9fFcz1auvZGmw6lmlu+tuymGaFmX23YAe3l4qhwHJgjo4UvwrtY2HtmHsZNVkAh9lWR
usW7WvNG927u/pltTDU24s8jhMuOHBFhq54j3RGZWxpf0/kCZpnUHVf30IkIxGKIuNS28bbqcZq3
XrwzSkaQkYaf2rJh/Zfq09kg4n0/YTHNARwwGLJZJmvF3diBAu5mJncp+jf4joK9Me3PdIqLRPKS
LXpLtQM5mA2fTxcPNl64iRrzLIX1WJ1gx7wRWNodjg3t7MBW33eVXeefzUkhRiDktWJxS58JM4Qv
n7WROyk6FW5KFKI5+TZwTLcmb/0G4ILkSe0OBV5clsrjfona0mUMN8rPEhfkXrgD9bnn1+QDqDbE
mJz8+cBdIpPVCIdkHlISVcB2rg59RMi7UE2p5H0T9buSMk6N7AQEZJrbvwqAK7A4+cy/HXVvk+UR
GG7RcR8pmymUw84cVdrujcv+rkbuY/vX85qUJczXAFpUQ9RvvYptL0MzBw9jj2yg//X/KA+zpZwh
tdDFBw1Y01n2hNPtOnpKvk3AitRLAVOkTpGPPFY+eAcJMsAX9SyaD8S0IrX7ZGp2F7s42gsELSls
3L8lNPv7px3XrDzWHP3EF0ZI3phLVpEjDhtdEGs9jekbOpV59FmYhN35UV6L9CDleqmq5YJGSfOy
RQXAoYBdHI62RJHqT09ix1v7XbtY4Wv3eVIylrrSAkkcxL9xKfiVecxWpoT5jGKOzuVW/MnDmyIP
aMj7qcBjnDl0sRhzRrvO/sfOP0MzxpOXuFidjUYt0TjsHePAqbRMBT9YMVXcRsKrSJ5tfi7wR8J+
kcQLd4phfmI5yTHnlotA6srbg4y35PdjVFE9nAG48ZIsXG9eq2kpYoiF/Vz6IyBQJlVvFrDiCsRN
M4/YDEh70l0s5aaD5WGd/QtBw37c90OoL40k3BcQ/bDkJPI1o5M/H/iwJAvC8QTGRepcpQxt1MBz
LfkWj8XvZQ56KzrjftlA8SycXcZzqVYTpYcJkLG+3QjEESzrB+y6JT09ooH/fpc9jfwQZsP53P7m
ieEUcNpndd3kn3HutEyTTGx5vTcrJ+U/ADesjf3YGQV1bw/GgTrjrKX3uzi4Fa5p14BYXGcUubyz
/8snaKHfUiuGjU2kFffmFw7jdkkvcTYHSj0T8VH0MLG79Uj2c8UGYtWU0k+8lNyaWI6zBO0NJRPn
EvEwNusVVS2NlFoYo9y9h705eRp9+waV8bTByEU59JQlqTUy+v4GaBkkMuLmVTYy7neDUymjBYWX
NqvR8SwYGk+8OWcHFY/6jH173HaDbrsqXL/axleHPX+UlpLE7SAdq5zNoMj1E68cdmSafxvn/Mfv
YJ6GhNrF/lASYy8VVG4tRrF+OIvalL0Yl3ZpOdhiOvutTtZBiOl0ChwcYbsV1tdUi1oVJSnEZ/UI
Gt8px5Co9YiJJ4WvWFo9iysirm3V6e8vHCVA0S2pq4pg9adpw+/0pQIubbwpEBRuYj/M5R2Xmadj
A6LlE6MI0UwZV1BCONd7dJ+yiR1I8z6SKpc020ltk/KLmHbGeXGKcdsFMr19LtMj367CDiYR3irP
moPUgrC6nEdIzdgsNsxdfDdLbgYGkaSuajfoqGQEN3I6Ae5bdLvDeBUFOvqZ4bYpLEIx7nEbxVa9
0NFISakeVe/yfPVOk7pAL/uspi0JdU9pvc6eAhzxk7lX9p/LHPiWgTGRf6tILC4yIa9978RjHyaQ
11b/yG66HY5aWwlv9MjgP1sKCy+rg+vDSrTXNky02zCOdYqt5nM/TVJ1GYa5O8EJRH9hGN36/ZgW
ASmD7Fsb6vo7ZNiJfVUyFdA7fRhj4PfLcDCdpyWrg7Ub5riszGwfjAhnCwPmN/4DRC2Qg+fh4SxV
VzD0w0/4sM62QwF7+jPO9PBx0QQ2HI5QGrhzD6JwyjKzhFV+oUx2afGdFBmOaoF8CxBIXYpiHS4/
UrOi2MLfrLdu9yJR5w02kbHwKnA6jvFREyIb3n/QH3iqkDcAW29stKQaHNyTfreSe+1tP5hXpIZ8
AYKGBMpGvqK+t4n3q77HIuN7vYqZRNXy7H7fO6yP9SbVft1TDv/0Ekhh/vp7lwrLxyuw4Ku3qrFN
9GPiLQ9k60+DLzlGCITwmn/9jUTwwyaJDt4Ys6rGkLHWdaL1ZhOn6nh3UYGDvZ8GCux+iEEWRdPF
0NirHU0PKTz9cQpta6fN7dQB7hNYUVcJlr0IbVHCSJbGk4d9CVGcAr3oEt80BnEpPCeTm4nEQucg
x0sVHc8BN4OCcO0ujoy6L0SfdLpg7LwQG5kCEh/CZGa9U09TeCEswTKyqCjMyu0hh/wtEeXuoG/a
gexYpdiloc8gdOsTPEnMQaPNhJSOwkdjVjiUF/VKtcNACqVBPhKyKdy4BMtG3u0lYCpVVDVp5YTZ
Y0UMc/PHLuOhxTMDlcHoC3KUuXo5hqGX9NeT3mgYeuyL75KBF8q6qqtR6T+DJrVeBw+oh0H83ZJX
5ucrLyniCtK37i6wwXWh6/whPWzYcg3owAqD58DiAM0hxy5x+ne76ZQG6MG0P70L4S1572DhZDoV
InNy01keDqumuxLagUjzinu2+8aw9eTU1CXMYjxYWJYN0Wby828FYw0RDfb1uArmT45rCVdeIQm8
B3O6zRYX44pq57TKKi749TDL/YpkCw7faFW8o4fBBwt2JxRECKV/NOAKsc4mO2gH+yGrBNQVhYct
v6wQ2zn4bxfifS4QjfE3HxpEG/LalrtFj4mBXRrMeM0afET1kvcYddn+QArR4CEzNTfZEakH3lmH
a1pfSjVbZQaVIZT0+Wwgdif0es8TJudWRTxi8p07g8jwzmPOdwbSi1EG+SkFGgjeRq1H96sw/FpQ
PERdw6j1vvn+aVle4At/Vrmf5f1n0eSd3sz8X13uFgd5ZCNn7jqio5wG0dqc85+vTczMvf8sCYvm
WgqQiXTOMLwm76zk8s6pOezqmzu/IIPRnVeDj4ELecXlSjki8+E4WhFMdoK0du5ymmx16LGoSN02
rPb/XhyH+JiSZXvUkT35x/BXLiSm7vzexPIfN7NUPil2K7pHF+rLc8M8f1l6BJiNYAsmMcKUiCYV
aplBoDZr0qSpzhDTQO1vwCrskGuUbfegkBkTSx7XDrerP6+IBlKTbFCWWKkiFnrP+OVJspr9YTgo
S88Zug1dBrK/JvcJZno6C6Ae3Np87QPXotCkbfbYmNuDM56swaQoqm7Pj71wnrKN9r1VaeFubsGn
0159ekS5pUhFiN7O/RqHIsI9wfRr25WOfG4hjnQbJK3r0EaTv4y/XBLDvGBOf4uBaeo84PGQi6f5
A8doLnr08XrNeyqIhK4qnFSmzGyY3+L03IkhtJ+qkCPQgUEQZ0pg89FD0AadFobuAdHiRM5tJ+ee
7vX12InomWU53hc67JI12o3C9LupPYUYS03QFRd5REAKY0HGAD0oes1Wo+HpV7bix2U4BrNfI/jz
Eca1JdNWLP9hUTBEZYQYmb//ieogaJz8MSBpiaf8bbPRjDSwv112ZFDE9i/JTqzfVZWeIsJIqYTA
Dqcf0lBiJgv78Ut/3hZWdTpIxGmcHHjhxVpOuwZm4VvtX9lZ3dVq/mB3qIwKfsXFEuzrLkF7iFab
W0jJv3lKQzRYO/RvQed69Pr9Sz9TBXTOxKmmlcs1nhx08+pd3Tyi8hiZMIvm+oQ7A6DnCCG4OaFi
0OLD3jA1DU5RcLI44ClHcGAQPBHYKqIRYr5AW5e6EePVMtPnGMZeDlLg7RBongc/4TosGR/4Kdww
2qhsUdw0J72ZrHjdhuj4SH9yzji615lWhT8SyO6INDd0wVEXbND6LIdEvgOO4LMTJR20e5TAnPFx
CjxNLCw/bAWZOISlu+XljKITraANlG0Ov5iu/ViafEISO/Zkt+6AN0UjZSh55DrT8o3jF3SFucsV
DI9RvgI7ScTGwlbV2SH4UOaj2CidlPXZgtRKtcobcm/qdrLTrYExMUP8XmnLxm8Ox7Ph6g37vvjk
8Mq8lLHugfK8t6Hdl0nV/tlmFxmQhcHM/z1sxmL8uhCtOqcRG428Ma+gxY4x5DGB6TbIiDs3iePd
lqt561y5kFLFenmKP2wESwhkGHWeZRf8CHYPzPO6dlaGxIa34htbPxxY4sMb8vyl/DcUQ8otyRfV
pL8Wpt3ZtR2xabi5/cjR3lty8kNzelauMNNEpVX8uL4sVzEgfaKAy11jyraGva22XBxwD2AmVaHP
4Ypu1AU5w71TPFR95z5wJFPRs0twO0EaSEFIMaBOk6oArZMFSpBB55iktc8Ddy8YXar2l0c7qJRS
hdGyr0KAh8JZMucqfiHBDpCSoPCw+y8MvoB04WaFkp5kbGK25yPPIMAVfpxJX/GzJ8jBO9pEmZZM
PJ2sCtG/09uhJJG4naopjnWSdSNs8e280NhjTh4j+sDvSz3Ji3f2sAerTSoon/xTHl4cdLSSczON
ZY5vPPYRUosLUA+PhSBHFKqC6iD2/QIXhDVs9X19J6mZi1G20y6mk9EsCr8ZlHCTOkWRu5SLRcnK
xIQ3fJHtIGhYbKg/K69HgvqJALQ2B2gQhzPVKYkFt5FXGceMEpI5ogsVY7OJr6IGZXzhlslqZq8a
OsGCtbyvjaUi3sGk/kpT8xgQ4fHlUHfn+rXQfwh16k6Au+Qp+p82SP8ddbrP+5bVIyijRCbqM5nh
6F6FTsmdwglJ2rmcIAa/zNpS+YzLrcEypBm+q6BSiOiVo+fi/mGog2ZSDSeSFw+LfUp8kRe6nmLx
sgDcfxtvwDEXAgxcHPDDtKrDW9QaCKvwxdpS37FY0Zsl3MTYBLupt9ETvN3pwDgpsPm/oWLlbDdn
HsrGUpqCakQEDt0fPRDYUAzSqOkWKyOKgY3hOp+u1/lv4+5qCoLCkke1ju2P7bLUNUu8TahoMRAA
dKieW9OqYYZULBWMiSn8x3vKX8kirBEe0tC4KUUIGO0XxQNgYOqvyXvX9E8FmFj27N4+iS47TKRs
cL0GnluPoyl/D8utBiU2VRa+WhTMTFXa6dMMeoAsGv5dDpKZihCubhxxB4X9gq0fn+md79iBYy7V
LIi0uqKTWSUHt8sAkZ/eHKpYBzC+bVqu7ydiOW5GMmxjIKABfQ7cBFO/b4zt5yauo80N8RnDIYdW
5mEVLR91qC0AyBA8Yj794tH/BC7wIJIwk21mrIkXJoQ0mzA2g4RzQ/yAutnuT8uWftnKhoL38sQj
nFLCsnK4K6XnI0hQPmY5V+N4I9Kqn7TtT+b8ubS23JE+6GKeJzoLn11tt8NiM4fsUO1ccoklNicH
s0GtA0vOJwXd8uounARjGhcqQzABcvrNZJyJ263iwS+wx87+a0VzXobIHlA17yOY4bU+OxPzbC/v
xgaXdTDtGeSS2+DW697fJ1xXvxwIbLo0tq+PC+Z1q8VyiShoK82Tula+KnGZxQ4Mwh9A4WD9dHmN
qspv87E9n8RlzoXKujWAZRw0ou+7OzdGTqeVgYVSFyYo8HeIUnmH2zmJh+Ajmm5HVE0SuCHdX34G
IqkO2ucTUto1shJMdcjRkyWawtqAtra7kvR9MbLmC+kCxxQ38IfPl8wJwP3OPewK7oQd2NjkJ5Yf
iwABed6PugfLhJ1oYtxLYj3Fcvchh+phE6Odd+D6T9jwIA4a14IR888eOqQ7Awai+XaIEKrjoJ7f
yjafMhj7DZQwDPnJPTWpz1KvbK9CBMFUEIvwm74lByEw18YmuAVTiJtyUWFMtjdkiYJPNqCnHbmH
wYFdB/jN37JmE47UJUMHdCFhIWYHQ/OC6+9L7t8yi/02QBxYo+R2SbT65TpjF9N0/OKxJ2lVtNV9
S6t2cT615XQFB2X1hL19p+evJxxVd7yPp9bCvB00+Q+xscnJiJdF0p2CEGSvMtadn6We5yw9g0U5
928gbu7CwCxoH9/V0b2x1mRqPTznCbytQ/fMitb7awFZ7F+ZbvMERKPbQzOTX2Yf4NJcKQPfKgUU
6Pw/voSwmS92BrotFcGRTgHRV2KQQ0FzRXY8oAlRnb8frIkS9EQVanm8OjVd8sRnkPC2nh6DEOrG
IuDoq0hiT3Ozg5xnHKqxZKGVijoegka59J3hfM+T4AMK5+xutFOFfOJuCVM6oENseeIpShY5aJot
/w/yEbiB4ULzu/tB3IXEfdXFliK5/DgDsAVMsUFP2Y5szG3Ya1vuU6gl+VyeC3FSbKbHZBJpNa+g
QpKPevHvFH2i1gzch9p+RR8gQtPPkoomRW+CGau7YMrQVfzosSXjGrd5swRO1vZu2tTDYj2Qtwat
H4bNCkJNIgACdhmP2RGR/XqHdjWAblHNmr7jPxQMwCHSZGFZnhD/YzYQbTgJ3TJ7mC2xHgjnl6Tl
ZaqSwKfi/mJShOyBwO+bi4g736Mr3p6zq2sVlUJHOYFKIJhleaRtsaiVDZ0TSXH6r6o9DCzaRxCf
x+N3CRKOfWqfsGa9DAMYdKZ4Abh/OOJ9k9VmlzJeKOxkKa1YpVDSOH1XgrfRnp+809Nsfmhv/ZjY
C2HihUPscAoWMmwJAxH3Gat5CQxlBC/3a3dkH7y1qqQepPOhh3QDB3bLmG5jdtFtCebMG+6jQj/L
Pv0IQov79MY6Wh/5DCR2J7pjtiVA8kIHZ6b/8pOSGs9Twix8mTDiJZ06TmTNNwCKYQK2anqKjCfN
Nn2PZl9oFVZhD2md7VOoTIFF/VDwUZZ6g8it4Odcf62+uZZ1r3g3wGePYaFl8S3SZda3GCS5g7om
Ukap5dtUoas7CV8g/tAx96v797PcSG5zcS46oklP36nfRN+L7TWt8ibnkqDhrmYaDu09e9BCW5dY
fESKz4LevDXfWlNsr1lvohoCkDknteOaRNQAwYVu8iBRfuNQrErLksvj/hDZFM67Mi7rFMk3ygNw
O2MvzlZF/1nDAgXGkvKlKV/Vj1B90d4cdCpkSowbw82ffNTa339FraQITiD4sJALZ+zeclqP6rbf
IsLpNbWdyJ7V2R/ObtnqNDnruCdfmpaKoFYk0OGyQ/6BYd+BLjE6aZKM56PxDQzgMbiSD1mk77hQ
uM/KNi4D6oz+PEdxb3Q72jgQ8rMclBvX33SfVWNfLjZU0aGP0V7hgIxiuqgbTGwhLncumvYP0DVj
c/D3ik4mwOSJXh1VG1H8ElKMVKFgOXGXXZFtyyXe9vyS6VxcS47Kfx+tq29TV/DeX9lhsxCHYg4u
lg9X6Nb/s2r1qHQ41wcWVBW/1U+URcPaXlqj/RiERA6+fLS+DTT0WIedeeOQ+12AaEzjKpodFeg4
jqVCYvWfB4xn90JiCB5MN/mPDE8b+cmk+GgLTgxa73EJg28RTXe+dkoXrUcUHDwTXKjub5OimZ31
RsYzUbYVdxGcgPrLFxVOK2KRrmS3yvue0x82XQKv5hRtZ7e4n3jSiFkw38VFlsBGu4yxnjbdY9LI
Itp1mNIu1JtkUrmytUcxayOnt5xUAWhpWi1bod65pQTYGXcuhW/3/JN+aohUhOGNsHA/BAgWBPQI
aC7V17eTfBdJOiJ0gDe7Y59QS14prwu/Z2CWC8PegG9GTtHG/zLc+Ml11ko7KxY5mbQcsNk/lRzm
7B2wprnS8pukDlKOPXcWBBwJq0FG0cEGwB9HXQl7op5lmTMz8irOSxEW5eMQc2Ueu7POTvLvh8yE
enak4JV4Ve3cslNFcEcyy8QMZjfJeB+HGr1Kyw6+VZfMBXD8o2K/y3cRgMOodjEmwu8NCJImaFhZ
eFT8SBvi2UHH9C68iqxIVk+5jOUADzoMtflrQceZBQOSXnaxqpw7LPk7rps5nMUcGNmoFkw/OyHM
3LMKXH3OIFpPhac2h8JVIN/KvvMZJE+Hw/KFyY8tCecVvVxK1XPX9X1bOe2fZcq+Oib7mUd6YI6O
D/oAbb3KKLKy1rv5QbAh3Bvpfw9mb4c5ERKnvyBp+Ji5OhrNb2JEfG+cCRqqVmbg9LYNoz1Tt/cL
VtnsbL72HxO38d0nzMvNzZECtRlY3LpAxm7Q+2LpqpzXRhbqKL0PPFS/Y8H3JJE9pMQ3kF1zeYyB
DMFE+S4Qo9vmnRu3HoJoMgQC+WwkYfx0WIclPMlGV0W5tgaOCffWeXfh0B66Ix4z+xfCrJUtGw/1
W6ZhVZmCLzOb92BuH68A7JkXcg2Xn3Pd926kxIWsh6brNe3P9UAJRkedjduesvppht3wNfYu9LT+
z4B6kkiOCXA2D7icKfBfTn1Z1uciVdptQZRAhZSH1TFZ5o5HQMfwFPju6OdsE7AkhFFjtauAVf3O
+izong2dM6ep3Aj+Fqoq6hlPdQVSmPtl/AJBERZu+d4+k1aNNWqJYNSC5VQkmSrP+rPuFZsJ78Ro
x65hxlUwNl3bsg/pV/DB3fs5buVxn0bwKtGpP896HHy8M1TpRIeIwRqShl8lXH2BYJ39Mw+viiG6
Eridy9arfRKLE81tDHjk9RQNMCC8Vz9RtEn9FE6ztFpI8B9uWcJCt+0wbSjGy7JBhAklLKXRJFhJ
JxSWISCc35sgZ68+IJEzXKId20tZm7bhdQ3C78MQMCVs9l909vKdteRA595k8Cjy5xgPXrLnwGTl
IhB6Pq1O8FLfxcLcYJhGN8cZqrStCledV7ljTlHymW1I2ZmyfAS/POiDY7gy1uS4v6x63HpQaj97
iDLWrWNnRYD4IM2gOY2l1o8eg9WxpozcUMFZ/fNdT0eaA6rWUi87h6p4HBLMYiod06yWvQ+xevE5
hnNE3s7/idGhKeV2YivDGsqgXhn67hd+6iOUNJbV00mrRMjaUzz2ey7yMvp2Qn7dOh+/8erp4Pia
uNrJHuaasZKo8InZ7Ufgj8j9e9Kz1GrcRq14biHi+kqd0tkoH8yDr7d01H/eesmzvfAQVSP6xkJ1
dcxaDqG1mEX38L9ey6FEeBYvlL9UWV+IvUhH8JoK/QsycfJ2NYqU2HivL7z/KHDZVA3XaXvPs+zR
ttKkuTXH5KH6zJcsahR5TvqbxmhKFJiPEaXAuno/ESnUzszuok9lzrZcjdpa9BtVwlv9T2Wvtp5W
BDX/PszMwn7+PU8VZkfLLYpCcuiRVX3gN969bWgdOOy6NT3+k1bkE75X3rnj+/GvjEACdje6y0xU
SUWv9/H+1WvpTrv/iZ9uJ7ChN6ufLGfGoDrcwueG3bYpKOSHNExlYWrP6MtL3g6B6cwr0llfqVTS
lE17nySUBRuFpoFaYWsJaBKMHiOUtCRCa3VhpfbVOw62eUsHPyE50ReyLcNgVtWZqmRWZmR6F/Mo
Hkio4l3wJCWLkQxtlMovFgJdsH8vDaI29qykL/Oa3bx3nLiUagF5vEE2oOLCM6wsMqGVUhFso97a
6LNgDu3b3Z3wwKzOZT5sMBb6XotSpGcaKjjkSjI8FLVD7Di0cE0xKm2ZH6Y6QNTT9HWBKsHXnqAr
k+yuksJNxAaa5unWstoADVjVB2kyAo9oTJd0Oc4EmNv6yUe9qlW8Oy4qbUv7gkohKpmJR7QeYYvH
emR7iAi/sMsGaW6K5lUJpakcoCv5168mUFQ1J2t+G9Zfj4Uc4zG0DT1giTm/QI0aIuHyoLWf1/tC
4NV63bhitsjF9nVqfzpQOvKaLWjEyvhywYiw0xbOdAn9gzN7Eneim5cCthBYcu9y3RLJ5EpBjW/W
LI3KiMDcYGZyqYsy5wolbBNOvrHuoe1tGTRc1v/w20UzwmDTF1oNHMNxAMijvpHVQhyhQ7nnPhrP
KmuEWIhB2dNkH5jtM8uZlZRSAl/AYxEI6wzohRYGDiYqiKyDrhNjcHXPPttvLjILEEyO6pzNDJnR
zWdcZM4t8DuThYG6fZKXeCJGb04ExYoT8RlonShZxHpWlhS8YDHpKDdJCZN1rZO4sIlFoMsitcgt
wunewYXdoAgxIYKQgHEy6zgVXaNp8EChyAOgHA2cLXcwWtqjFlTjZzNRhJsS5ZmPxXK5hONrQRJP
M/9Y/KTwSU2JPwIWWZeoW7CVp09196HzX8Sz5XJ2a+L/nwUUz1IdREC5sQyvcKZbJzBk+pKl2N7/
fOpFg6c7FThV9spOEaldeEBD83GCECC/9Nj5uEg0rKivYZSLQlVyT1wOeDib9euZ68sRN6gKaZH9
/ZRzL6ArKbhy0pRSom1Y6KP5o/8RpFoLFc3KQIiZjclWcx69cVsXyboLLVkA8ow2mdI9O6Xb1T4+
c+m+yCmpNcbzGNL86+lks6tjVx1pPEM9fhrUFw//55dJ+wjy1h7XOApXdwhYzQHTiVY3NtQLqXGk
+oTRElXA3tBdB3/GsC19tljnZkOGg6tPvAgWLAY8x+++qBvaiRMqGuUjRyQbbDxajhgSDAU96s6e
YU5lyvocLSdrgRoLuDtGih22bzybG6SQNFpRMVM2Aoar9rzLvsoxvVCAOdsh1hydbub9aPHspPq1
G2adW9rarJz7/gmj3gcJCAX8vtqhXSzEHBoJliUvz42bBGtpHyMUWwU/UatnrsqGt77aBb+j+O/c
RijWvT5cte27VaacoJbN97eY7q26hMNyKH05VYVAN/qX6Mw0WN6xW0czdK3s5VA+xl9uI6xWN2jy
xuqyy705d0EAgsjPvMq9DLrWZwDMwkSMA/qfauBo9OgmjQ9yPmXebUSAUNse7DR8xEVaS1xxLQMV
vSi52sdvWRbfX6GI9qbt3DSTr6FTcSSXQRLw+v5XKRXjxLF2pmVYrios/hKymKjmbVpOPN3c29ny
w/G84p34bQ1euvyvDc77xIriR+G6Ih1z/7+CFNwxHPRdsriyBQIN+4ldSB9cAxANo50lDo+hjAe7
q22Qy0fFQRsd763FD+L/xjn8mJ8t7i8nFE8ev8ZnFxAAMmUiqRp1yQasU1rMK4noF52qVo2mdCFB
6nngWLuGTes+QpAkuwL2/QpS+bXhuEHkfWsRGflrnLF9f/7u50rWk1zzjk8rNd/fvJUQW5Ezxs9n
PTrQsjdU8M+Dn5Kv02Xw3nCGoxKXm/d6aNDsGhiIcDDFsjQMWx4WqEkT9VT9Z/8peoFYFgfq+JG0
0stmUYuePR3to2WM5djXrLadcUOXuIj6S92dlJHijrxZ2L/bJ80ypRz0pCKq6gv2BU5rAYI7CNs6
kyf331KRZOx3QCEHqdCNSJu3Tb7vOVr+4q/g9q2LZDsouqF3cgvmqa8SF5+tblO6fj41qhjoxFCA
yw9UV4d3vJwuv8XMFSK5A30mNs01RmwBkeOBy1fir2/ToYuZCjV33EuCrP+Tdqbepg+ZuLyeOA0t
UELHQRpMDV7BjtZDK6CAt59fd4OVwDWyZU3DwaVfa8wUOH4wtLdC0sH0j1Wdz4Xrm5bzCDiYg+sP
GFP/bWzsMByP26+iPQwuADtg4BjpX7bM5MSNaZjf+wKu4ZLDLIRGK64FRrN/pSY5/H45TPOLrgsS
wx0L3H7AuwcBfag9BY+Di3+YOp1EUu/7M7gJTfXjyulhAImbBbrAhrlDKwYsHbGpe/aUKwVU91jC
QC8Wmrpg2UO0JGWRHAWij6plIo7Sk/4ptB1GVKaVyADtJBpVoYbz9V6/Oh5z3ndEjblwKNNQv1qP
LDKBVzedfpN0um1SiYSB7udEETEptbvYL+m2mMyvN8gx/nUyyuxJY5sXQZGiVE84t+iiigngwUDk
aWcLgbR/MZNltdat99tqbBjCd8NwZ3esCf13uwpYEl2LKt8bGzKkxlFZDWFWT5ERp5q9qvB6FZu2
07j2ZYpk6Ahpj74SSm411r1wejXWVG86Mufd6YN8dY0NBWYMwX+ookFsVkscmSqr7EP8NmDsjAcI
Ze5Eu7SK40JosY5apVQLDtFdR/6secNxz46gkTCvASVTfIwUs4pLWK7gjZvC/2/tupDJ93kNxUIc
PFHfZ9UWl1de812MoB9+uD5e/uWC79MznNcvma0Xp/CjLOx9RecV02sS6ZEQJbVa7sUFVeQ3h9iu
+1kctT6R3y0Tq2/lrQdVZJkiBl9H7pdqYl5cZWMlwXQDp37YYV2ZkA+y+PB9C9nBjC5wud4vsz6P
pfTy/8+JBJw5R6d6FLpU3Hgt4m+c2qdBtDpxH/iM3r7GPW56JPDLdDEjTfWOb4yGovkgRDMG6xf4
ItLz9HtjAYwHK+vWT3xpPLDMwiDquOrqXEXZCP+i46T2bBZNFwx9f1q6BIbwXRliA2yT1AC7JKsd
PxzDcpHpWz3Sdl4ymUWW+mV6gtHyWEPFaNzLrs/nDwbFHHK6eiKyw+IvYVoGGcJlxi91tcXnxGqr
Ko1f/kcDrGKBqaBVuU6I7l6Dpu+mqoT8MoBUPQMXMKVdpikFyf9AifU+Qh29zdMEEcuqsDPblf0n
OIBMAYJgj9jxKIzVt/Gyfpi814wo4KcL/CKn9GiMBdbIiKRi+lKrELC41MnAnPRaKAFnDBFUHiwY
GSJzTMGDyQCNW/Z35ZKxXxTwO+9r9RPpP0pAhxsaeBgfJmCsPzay/isvjFzf2WcEkF2MQ0GMKlfL
iM9Y80ExQN5vWLhZo5+AVQEjf7iZ9vnAM5eArnATbMluRddd9CR8/MUK07AfSC4XF1wM0iBcJYDk
4doCBctwKIaG2aluDr4qvs8GyJlOmezpbNf2YmXsY7Jn4766bhCE9bFjWgcwB0rkFl4ZMIiiorqv
TV3GEm9yaH9OVYDPvIUXETVO+Y1AUqsbRv2NYas6EiMZLvEIXXg5ikJcAEe6W+XAzTrETmIOPAIg
KCmFWwzTkXuWJcSAcxmwdSFJOqsRW+61kL+sL6dhVHgvlTq3NaX7VNq7+SJE4DAewwNImJs5sHN+
C8E/B8fQDFZ9DyU5qXmDKTEuaGTRQYCjadoEhLDpavcrNDNSUV3I9W/ky+v17+4ajBj70nR2Szwz
pNSTE7K59EmwbspzqllVsOBe8WMg1tCTUyFSGixHOdQy3yCjImIpYz/jNETehVGGOKpqCmEs2b+S
QfQl82wxJAdd98e6E8IjXBR0FhW7PnSamIV44Lg0LjYbXanQH3ojBELTZLuYQ6AdchIAie+i99Zs
IdNk8L1u6fNd2OpGNVMw7u3nNmoPQ5DZbAT38jdGHcDhHCoRmyCy3VtnLBXg7deceEUGhF4/pXeL
PVvNFxsOr7VBXPybcHxP4IJy5HjLprCcNlsMv1PTqjonJpdWfSZKuTihOYJCJTUreupgoQYDuwCL
ep8H6GgKvVdnkvJiBG2Kzwqsue/Gz4ADkRmJncKu6MWRS+KAflLpgkp5R2QaDHATv733ht7itJTL
VRNBc2BiQDtR81SwTDEU/m3hfMtMLcXeHXX0AJqWc2RXdzu5OI63kdc9xOwtxY6cIbvuGHzB/afn
Go6pTegIdnZx29GcC3OscU3teTdo18NTRZelFO9rriVYWm+CHM8qHZuiOeZbjVAN1TYIF6D4fVks
FTXspBXCywyfMrQRurcEjK1otKxCI3dXrYXrVPnmKEI4Qizv0TOjTrmBq+4pJnGsTpwS4tqM2cZM
0AJW9TrRiLjHK74bbeMp5NCySC052cySUywlAEb8U0yLrnNOyKqzZ5fwiv+J/iJZOcDCTVikFiCw
D7/jkn9881JfysB04UxuxMZJWwsEVkr0MX/OJR+BjOONYchEJ9VyOC9/2tiQbbWFNVJks2H3Mtbw
YAMRWIR26zx7tp/eF5R0PQUSD8CAj+LyuztGM+QCpmMykDmHqp0cGVbUVjFeF/0Y0K2V1CCFYM3a
PL06g7Yc/trTqzw+VGD5HcCsTsKnZKrvPAoSgEAPrlhp46Fv/ZqYIrsqw1lf1dYVm2fhH2QBbW8r
yfpL7sy9eaZQz035sfbY6U+XZ3V0FGAbVRXTRs4Ux9rk4CqXSRNhvgYBkf3C5Mce97JpP/WSuxIe
1td9GcL6hjqvxdFGONgkpU0LkhbOJ/aqsw1gJZDd/tHLOrVMCW8NWi60H+7PO51gTOaddE2O4v2J
VyoqMRlrlWBCtGjs0PP5ilScN0jQt75P4TnZXzVIexyoanH5FV+M6FFM/GWnFlvBbSt+R8X/u5i/
jf6MkAjBFCualYr/6dUWHQDQPMYieBMHQeCF07ZzQAtFJK9tb60TkweY6y8uQInuF3Z9a9y60rnz
Nve85KaJ6033qnEvnsBJlGnc3kpiC0wWO3k5n3+u2XDW+/lePoVlyslOLTS2GSGnFcgVOPv7cXSS
ecYpCcWWg+bHkN3D2B5vACFQG6AKcwY3KGoQUs6KH1LmTlX3rOVCsuMyVNBszg5xcr/K2LhhD2Gg
DXrarTP0+1pF9pO3kdt+wmlN4TkAm1d/GL756XCciV8J1n0ql3QXF8E6tjnScKx0nRBsli/SEEqv
Rga3GCaY2GznT7D4jy+6CjaDVGRBHYE7v2aWzVgrRT2RYHsfRt42LULP8shT0wpnE18zO335WwEN
Hl2dFrA8tUQKTIrW8mmp++IHLC8XqwC3uT8I7+xf6VaCmy9ne9PDrM4o2PUudikMNC0dxzPxlsxk
+zvQKn5FWU5gkWiuXdZ76R2ksScMmgTXdQRBYdFemMoooPR8ekrrAKW3nuG1lT9CQnvRdGI9P3EO
MnU4FMPCvYPWY2X2b8W8ZTSzYCReamnKLOFlJlWZRqsqJPy8Bx2h49o7NIR/s6twWkvCmbzejDfP
IX1TYqpOCUosNwia9aNfZZ+Ue+l0UcbJF5FEOV73AB9Ihwd8AJweBiO0tRcWwoa+CbNFYzM3xs/4
xK4Gsq0VT/xsZvicKWMPsy5DkiW1Tr/w+vhB4cuhe5Qd9o6xWhLXDnsFM2sFdw9yGXC2LsSBo+p2
A1DFn3VfjWbKQq6sMrSZgS3etIv+ZT/0OJ+jOrEAiTs0iqktn/8sZOHtuUMvdCq4XAukr2ht4+Hk
iSTxvcCxWxDyN7Wr+dYj+8GfJ7agkvXTudE2HSiBbak6YDtS4mLu0mVOCc1plKE+sB/Y9pGWbdcz
gERluu5dmUA2GUoBBaIetMU2Bw6thFDvRmSyhDC0k2FwWWQmFVb7Fnt8Il/zV05Ffa07rFFzvVsX
gTgmAg/fPr1HuVedUzvuBlu3fP1rjgbhmCOKVPULqmsWsGVXws3LeAEAZBJsfTrRHCZ/Iw0wBnxi
uwOtySrepquaC+n0fmrOG7jfK9W0a/07zryrSjkZzK706r684FABZTt1aPGD1f1sTP5+paV3gKzU
HY3kGKhgKK0KDlUHtY0IAIl9YOGYMqYbq3Jsk2B+Y7rRk/SeUkn2wH/m1vkLj1lo5QEM8Qauo6FN
h3cxyubONI359iitLfYvcRS+KrS2ZTQ+Zut+qbFT09AZCqQDWDeTMk9roLMGhiaCMfWDVCb+gv/F
mmW4sXixekaRZKpXNgTiK5SrY92YHEQW4iIZHAi0QErcTsNQC2ygQTLH/m7GCXyflljZBdvn+cmh
O/MTyjGr3P9HHUbMKKqkjmlQiMz6/eTXHzQDcvnSW8cED5ltK01FdKA07RPDle09sWc8Ci6ufTIN
3mTOrMzkxOxpLe76Wqf5+Kp7zstKQtpZhM1fqfvQb0qtuSc8zjB8qYF9F0t1LFuv6+wvxGjJlZBo
yAs5PokhXSOAoWM1yDanGSE6Knr3cUXeg1RyhmJHsipq6XEiQpADHl7otjUrKbbcF0tyECiz9vHe
Yu6HktBRoSlgG+sm3NeY9oThf2g9KpPyU45syttbugoabmr4ByRiq1WHxNtaYqtUP/5ZHAnHBy5D
H0Za2WPRuo0CmJ8xpy/P5uxwAdGpqsWTneDVn8i3U8n1j/TuTceHYAFJw3nudp/obM7YX90DPV3c
+5CsnEv9JHABPUY98CmahNcsAa0Vgr1z59newuOls/UJs6cuamMGRgqicdv/9GMMOGmukTgOw5Cz
82OyqBpyBgFy+GZDhw+WVZysggkDak2eOhK0tO/Zk0cKx3MdH9Plog1nRpIuFjA52evoI9Zwczbq
EtGeSpiPUX8/XZKuB+aYC014eLHBUhk5zyLzZVq10ioqSg3O1mRKE/z1yZknWzEhwPD7MjZ2u4Dk
47qFpUnZPiQSUJhTQq6SwhNlZBD8KJszd+ex/glu8uHJfA30waWgi1sXUcbsx9dy9OghSc0gpwrg
wba0/ECTdvJCs/zijNU1dhwHWqMppzfkH9Ci5Cd174U9sfSXC6WWxJeFODNePfmd8kKdI64i2CjF
thhMiWVF/NKSsPIcjonjlZlWjPh5TymIJn7LM5lxDawgkJ6TordaQwNsV6e0WAVRW8uAtykwnQ4x
qUOZ8m4TJ8jlrZn9GYkSMt1BXaXQlcqwnuHjaw5G6+heW+6xVpd4TEhB3PWNUFZOqQ8SOydBHQHF
BWWOf7+uifEE1OX7gEpy0xZ2GtTMHmaNUxc19iUEV2Yi/IU7EsNX9351TbSgGSYGMpUnmROaBmT6
lq/bxaxDiyBw6CfLrUohMlLx6AexjLQP2IXfcZmA8JedQDvf24lPad9NHFnlDS43tYUaJ+s59uLn
gi2nOFUvlptE5DNlFDLXoZQPpZmgc6dGp4+AGtOdNsKSJPHcHgYPKAHxEeJyowk7XWo28MmkSuz2
20rjJkBFv2PJ3ugPcdNw8nYUljzYRoGul15PGHWlRecwMbFvBo2XHg1eAwaPWSt2btJTZNQm613Q
QcBpyxP9xvWQ8Zf7tkMNywBar0RaZ2BNfpnXl1xugP3ELCyx68AFcqG6pp9+/kc04NQqjSrGPxTl
Q2IodETOJB9KJJli9XTqa6GGoxoEZBS9R7dQ0ulmsQlsETAl8Diw7d0mxTY65R6kl1JcPjALZPc+
XsymVDrUiIkvhvsnEvppvXXzIQLFK+5JArOA9HY5eCxbWWnqXOt27lndLcB/gGnpV9EzsFdf7ups
kQSQl2EjODJdzrj8+YCZhrJ80SUxE0GU51mtB5ueRevqJzPu8jT2pCfxsAWW97owt1gyEC6RgKLL
X0Q2LaLk6szbPW9a8Qhqjkf2w1lrZF4Y9Rg38zzSH2KLMEi6p8ejDIvGJw57laA6/m9HJCkyzZH1
Rb3OcIO24e16L+lL1czHsmveG48rOoRC70SfpqnrrhvHmtJotHR/GL+qsv5TJ7kFTOrUYkkp56CC
SNfp674aSJLqJqp5Nx5O4lvQicnOabrKGd1+kuiLQmjneJdntCJL+iRjszAjXOoVFxjg5fhpqO1F
Hfh+m6HawtUcXoA8xPpbecmJ+M1qrMIQhMaX5cC+AmqAJEREcxWFZNi1ZX1hovAizRBoAJFxXig+
K4p1dkAjYvsedimg4h3mqgPgX3NluELrEMjxHMSGC9kVnN/RE0FhWlqGCvTkOP9Ttnxu46mIp0cQ
FZhQaatlbKTqf3DvKC697ln4XzwrrNgMzqSdvQbnuPmO2mUZNuWuw9j8Y7fF7HhJ8sPGyl8koGak
0Wkw2eVAJNEtD8MH0kZANBO9GcheYIXNffS93RUiUDSEETZD9fgpBSr5ybsXFW2ioTGeLxNbGJ+z
7rlRPeDw9Ycc6DGsj1kr9UzXhmo7+ZkH4wRm2GBK5Czd1Of0NbRGdONlIEYTqT3DekJ2qIHYe2hB
bN6x8nHyiDF5Y5H0+fFZHpc+Hvkn4n1NT1xSy5WdVHPZt6p68Ps/WFEBE8Izw+kbS9DoIe2j4OzR
yrTAPkLuRg2HTPMBK4u59/AJTpWeI98xUoecGNFTbVchZUjB8NKTU51fw4GatXiWi2UJH4bB02hx
mUiMfpqit/f6FqYk8Tym9qcQjpHgBWDGmPfBPZ3WkbQj5Y3OMvPa/L7DKucSxJDtimjYcz+R8YnK
aNxyhJrcBVvGP6v7/GmwyxoKeckZDTY7WI0CbcVdA5MV2U6mhHEhdxrgc0+zR4z1rKcMTX6SwQcs
YWH7HX5cVGgNYNpD/pdD1u+A9MRvOJQjDTExb3Dwz2qF9UtIHPMdTakws2O0/RjvEJb++Tqe3mzs
S1mmFGyKZjE4C18u5T3uMrE82criIYcdC2mzj5z4++A/cDbEr8X4jnJzef2bzq98shQhTUQsRp76
cBdUKGZWmsB+W5yVjBHjf1UCa9+yz2k7vswM1/6tlqaInjOV64XmzBrLAGZA7QwS8D+97TOU72E7
zizT9AmblK+2vJckeTs0Ctowiq2Zd/DzfQGZ3hLONVLmUUj5xLzJWdSJ9yTTjPNXIIZ485EdpdCP
4fWAGtoxnF3NTbdMN0DRTzqbI0wn/qYW/I7wfUfm+Zdm4IwhZzb5ZVypOOBGJmK5NuUu5z7W4LLF
HFHbUSiFXjQhcasMG+ZIIofaKCH8N+VTVhJEvXOvJYcdMWyC29P6aPyzBdQFKbqJRihD5uWeUnwn
YrRmPnZnGjNj/qsdt3CJPQZuabuauWZzSKeR2OhDREKFuIlOh630TgScLcZTZ/KFLF4LEB+I3W5h
K0F7NgIL0EJgOZxfOuj2+tbxzdwY2PkMp2uGyQLTS+CojSU5W3qmKNQrGA8mv2xgCnq//+Nhgo3/
LPp4GlL0wF6EySNDqdQDDKhhU60daDjbOHVv/rKz45JdKlfhgPRX4K67wY1cXvqbbpkWPIP7nI5K
InVGHQF/bAb+XdgUtOpt8D1PNliGqU9co7LXTpLuvfrVF43Pl/0xTVQUrq0RuUwPEsHZWEeevxpK
up2amNMHKeB7Rw+pDE49SUISccsumj34u8d2PZpiGvAEmCYqW7BG4luS2e7/m3iQRL2zwbQO8aFt
GlY9rsqW3GGKlwJ4BZCsNnTSukfrM7Nl4RjKfB3naGQFDFrD37Gko06oE3YeKaYR1yVy3+jlCq17
SGhJTvDOj3zP4WlmP5niBIfkSraPKeNdJHvPgIUE+Sz09uqf+Kxd4J8qvkzLpnXXv+4xK3h+hevM
G5rwK6TYMzth/0E7+RQFBohlyiHopAg9d9ZuWQfyfRjwYExRzZtCSjuHQB/DLTodUPn7yPkRJ8YN
st5DmF2h11ec5lFl9duFBgzrm4kPsWvSFLwd1qoh+FomgLeC27ZRCLMC2JH+3tXIUuRSjcnjIDIP
CVhUIrZXC5tqkT+wSBcwQ9LLr9Gjn7/LULF+0cazGwkASfnjShNV2oe9c07/sEzLaH7IL2AX1i2s
bGBWyqE1Fs4DmIPz5NHQk2XYYQdohLnE8s15Clj/JIBghVlfL0s289u1tN3XJ6lUpw1bHgGn1JmO
3TS8ghbzvHhT3xqLVn5d7sXalfA6C2fejZ+hSVBPBaEdfznzL7rPuROc4XDgjAEUwBJDyXz7/aZ2
M0v+8/Uv4CadJObnGfohQbrATA9qlbPSDJ66IMzvf/fLSzSHX/GR7iw9gSmgoZiq96gd7cA54+1y
hPLkOsw2JBQR6Rcz760ZGiMb4ubX3Ah+9k2qNDGtSA2leBpzgRWIOq1ldB7xBVN0QYX4DZGh4Fux
Eqs24nVQSdXq2WzvRarPKARcS7SJVuBxhvfQoFmspm77uxOs5HHNwmHPEG5+CtIew4IpW0yME8QF
hE965VQ2wddCQM13W2JpR5ZoVdiDEz//0IsUF6CfCQ0C7FBF5i14GUp1zXQhS5G8oTGzZcwnqBTy
DNnhSc6t4iroE9WusFD443A+PCG5FRsbPVfEONjotwfHVjEEOfmhIhfYYO7z33wDC3YSZI4XJQ0l
HYco1/pyBi/KJ5EWds2ifTkt1CIPZGxXI3reCAzdV99caP5uQl57pKCMYGBOLlW2e6KEfSwNVmHT
E3yV+J+8ZobMFLRj2j7IMiXuXnRfnTZay36pYI/TEaSlSmGeQ69iANW2qc97FDxLmJS4LcPZuK4k
MbINMRrh2NmAFoeEtHUhmdhSPhACANDFF2DIYLMst7t9jD3brRHJgCKiXY/Oc4jz/3ESj6EUHCQL
O59McY7xvma/BZNaefaD1zol7JoZlT1Gtlost2uE9uOpKESh82LbeIO/wgLEEpkrrP9l3Knl79Ze
Sz/oZb6JH4+8mEbsB25M/FPMmtnqv2u8FzOjIv8H/mUIcOlcXXsmM/djC9vjdgGblUxs+qOXr0F7
YhdTpTldi80oblYOlAFW0iPKpxalZV0srKGPXzaMXXmdGYCCxl0lIqlsam1O8xE0JAxUjDup4fpz
wou5S2lc2WpI8NWCl3DPHb4i6xdWjKoZTdDDF8CX6/gJ8Jm4LeT3/1or48D3fqPAXduRVlMmC9Hf
kuL87AAO1oroF8aVdyDHMJhUm7N1fftNmnOwy5WfLhY9udvJh8N7l28RZs0XIiuikwNOFoRa9ZDT
yEcIm/6cGR+fPsbawx5sCiVhCNfCxf6M9BLwXxDfQvHmrY8a6v4+G6uyS8vdIVJrwaIzZ4qVhwc1
x237xguShJkwdkPg9nAsPbssPqoUVHHxWERwMPMHVvk0T5hzEProKi5XCbE1FeobXupURWUzB4By
DPoh3ECw5cV5mEJ/nXxZN3EofVJzhpVveAL5hJCA06b/eM/ZpX+eGpnfWyU+mIKPz01umZpEjhsh
kMbAlG2CZfxCd6JjOXDTHnLPf+7hD9V8o3AVASMmGbiNHBX10RXYNlglsJp2CdQM1AvQSitq8muN
dQ5K3qee07xEdfrN/i7ZlRa7zfmzWhERXpLcQnpeLqGs3iKO4Sbhl5YoxaAJVkVQ1CObH7dLZjQo
5Y87lUHzjHwPl/GJf+G6+d65PIwY7FoNCWP2UeX1ouxAYJ+evd2GmOIdS0J3REa8OAu0eMSZ3LnJ
nfw9uO+xZwZYz9AhuZMLzNU2dNoJsfaQpENMPWjSQiXlfGolznFy8dTTSlDrb1mZDYJYhKuHPFPg
ouo1TwHw0oC2zD0HQXdBLKaj/LEhlCxj4Gmk0pzA3hmuJ6TwWjZrx0cMSJai2eW3rLi+o9zbGHcg
SSZbedhEFJly86ijYEOvmVVvYU7VTaTa56//WtZvwwNnh7jTKsgIACQarSTVfd2ez96ItNieGNQx
qBZo1MJjtBB5Etidj2Zr4+vuOGFih4/GmnJvf5jZSw5vCR2A1qXLNSh32JnpICaR0rRrInmoByvH
w2jAxLjYS+UFBhqstlcG2TgvWX29UjfFhbCuQj/LJIerlIy6U5wB1fmmqcnEVf2omwc6Y1KNc2E+
X2qjuiIHE4bADZpZCdbzQjPlCQ5SJQEED4EdW0hzJn6QCFuA+MOQlC/zrPiypc3Ny6Ex7ILugO/1
lTS3kQKh98yYRL+E3NSd1UHAkDoZ4Die0vEwka69HINIR4+Vip9jS5b0VYz+QyvP3oMi5WjmSpKZ
s0LHKG9RbeVlMgiUnit1LeI+PJ3fqIbSThO/V0PBiUQSyLS05ogqxw0gI3ajoh0rri7evGvu+H+B
cZ9VTuvf5P9DqZ14+47DcVQGtK/gObC4kE/A0dPoaUwl3nobRObrpsBS2VsiDi48YiF07yg5f7xm
2WClk8nW7FYeKwwBPmqAPizuPX8WxFxer5MPENtX58Y4ZA8mPuZzq8pL6hhN3+c573YVekIAjEdF
4Xz4lp/sQDHj4F0AWkRipuNMRvJxyZYRXapXHyitQWD1zDgfopC5TclHdGwa4RMqjMHpnKTe4gAn
lLDwgIVPADltIdqbyHR8PJmAIfDyfrx28VJ+AbrXdGKzwd4dV2Ddgb73D4vcQzkN3Xdn4y+vBUoX
r15trPQmHKiPRZq+rg0yi5YupEgL8W5oJ2hfNcEB9ws3KVrs1TL3jLaRqotNRYNx95fwBEgnBPEk
Ps0lRQ4+Ifnc0U5lSZ5XoXGrpC2BqGFjESth3rX8VMr4VXAQZf8FBTxxYbcwRzxV2Tt22qGLzjUz
oEJU4mg1CsWPhgqj2yp80HTs1+KDG3F0IXpebZAH23eE8qJG1P/WV+c1H7auqgBJOfO8F2UFaiVA
IcUUNAhyUyXs8q5Kwho5Z6yfgZzJuDkbezrJTN8EvWtilS+DJut2zL7/+fIN6t0ckOnKsTkcdMCq
0RtPVt7+P6SEx2Yva6il+vyATuj2GBOSvlmyjedJ36jT6e4O/ARrW8BeJUm5wJ3AA5it4OiRaCC0
CF7NW9RCfY2g9YxeOpO9VJfSZNr+3onYAwFKWmZY+u1VR48z41nma4qovtLmoy8LnX2ZZzrNjt+w
Z5Y/CCvkXubzSHq+2YYLJvjE9jc5Gr17+nhE5FqZH8C6SochPYgpSbB/6z4hJaPy7iudehSaoVuc
1fAJoKaqfLVrgHiBM2VeKThtFvqADcn+lDAvpDCz2MqFxx97L05AomO7/Bvosp7ELd/r1Jpcw7Da
V1ot/rFpQR4aTyWCCTXXWAFzD3hPWAnn0npSA/yr+1ACyIB8Yj2n+aW3ZSQOEZBDoMBnDzJu3tEa
YLHJQBPN+Z3HAAZYIKAm3PGi6hZls26sNfkqo7adwXRDiNxuo1E60DqpICh3CH1bxkrqA9P+KURj
ZNSGdxhoa1fEtQ+B23qDdrgjkS/FKthAu/kYZSQ0qn9SIWFKIdZzSxb0e/b5CS8IdpfAy5ibCueY
ZGJXbx4VeRCgXQBT3ASbVxIGvDKDySSfxxz6R8Fw/Oe59govbeGQu3ff1mO8Eh++DDmXLfvVy4Q0
TLindYaRisfoJ8Z0qERsGbaPNvcxrebBVk1usVOPRHvGlIUdDJCSTEvJZb0fNI0QN5w4QUhWRObj
EyBWxs3+IREUct2ksKwVI4+AwP5iESk1ZppbqTY+68cw2HVnVudPmDRxvpfljieQOcXI6I1CfIRN
lnjtCYAPlzpY39XYEsaN39j1I7514wa1y4awKhOJCAw1c9lBdcZS0f3PsxhJb5V67wiMGgKhKfMq
EA/NtnoBWdiODAqnoWF8pknqMObldEbwmbowJe1yusmd/kyGJfYkipHi2iWjNLClbYEcL90Ez513
4JqStKbmEEkiXxXgnhNwFsZGf71hjD+CVztDZUo+WX9JGnLQYjYpsnMs2k845/uncf/ZwWqeuZfE
5IgC/oiBVS3pPI4tAUX/eM2ZPQTmxVxLkKOHi098od+eiMVwPU/tdPVaM+E/lDzUnHAXs6jsreOj
xFoOFDbQGkATpHtFX36owg/eszebAWO2Z93xwLxxyVoicVWH41iBP+t6piKkrPA07NfCGJHct09L
iSEIPPt9V+FO3bhD9av6udBGtdciICcs28VxrYI0Kr96hS1z9bzDWYzYijyReAjnrD8dCy60ZNDP
IR2uD1J3XVblrawvNo6rtDAg523xa5yCHd3uTN6dPO32rRMiQXbSpE6Wo5m75vBL11FXsW8GWbHf
FAt/oX+f1mfgUlXRaBi3QGy5kOAIqBNI0ULoBNpKBhgbEKV+fXV5DxtmnQy1ecYfmPy8TfOQRqe9
nStIriIghVaF41prSsIwmggPxIS/WCpcjN8BU0FdUDvyvGtyAonS/WbIlwKNfAHWxmy6d97lD2hh
pfW0u5nVH4S6n/+XhI+manXXNZkD/lybx71GP5IHQdT/05QRkyK6o8+fTjcoz60u/4ckG28Ra1D7
6PTfQihqgYdXbBuiKRuJpDRKzzTHXg5UjQxDNgdo8aBkTmZcCKk2G7BY4Qwjl/odIa91qnOYbY3P
Tk4L6alPjiUD/yEu/5D5/kDVNZa30ZB1WO8EOk90CXaVLdiOoy3j4kly3kZstkF0MDI+N8sjko9x
PHbJN7hoHg2TZ0s+tEX90hh59h+DqEDi8oD+k2GMcvRjQOpw2PhSEAbV9wc6YuGl6iDw0MPggZVa
VlZIGFhNQ+qMA2bWIybTHMUUogQ2t0CqsgbIzIzF8K8MdktnUg/0DBcwniZLv8jFogW0th1vLCju
6gAJujiyw6/Wf2x/sIVw3/dJ7QOnrvQLxLH1CXpLxR+nOTBLySE1muE5e9WBoVHXj1o+jxrujWpN
oz5TymGVONwaxbW8UnNr8mnI6FJCrC717vbWDGb5E1+xxOaB3B7DVbQNFjBVGZSSMkpKI4I91GpP
zYW2OCkSJFfCSopor+JbhPEER5LuzYHFa2F0RE6YocIVXngruLsvIGDfYI5XSCcnbJyXpVCMq46Q
8B5S6MYNjjvBb+q2irsexCBiQDg/pVHhR8ME8dnQOSVcEqvTEBQDO7w1zKW7Nb89qSBt8pgdTDdJ
giSH4h8HATVHrQ1bKByU3oJxrZYF2WVQZkdA4Rs+/F/ZiEgByGko6RFhy114ris5FJEsqwuOROlj
hu/nGvqICT/nRjaROChcFeKp3jb2lxoa6cfKUYwMVVTQ4lNnISwfFN6c9efLNCj5xUE8PxhKQQPy
HUpF0SAiJMq1i1eYvYDASkUfmQq3ZTnd7AyUbD1EhsbLnjQ61Y7RY8oBfQXAL/JnCi+Ss77Q5Toj
WnPEyg3QgmFhltLAXVKnT6D55BSIGCMnIIiFEjm3hRwla57hRw9z4WDtRF9fUeeSDJMt1qRebsGG
HQ9imp7uz/3DTCNRNIbeDjNi4bpLclu2m51F+azxk3tkJaTZDn0S2GKDHDBb3oXMulRoQukoH1a4
vhiW+0Rf4fZJP/AVaWT+uCoBssLzdpm+poow2oecw1eU2jiZ/WJnBhLIW9GV4l23Up7FFPsmQWWY
uruCbGgxprAwXVAKr0qeEMi7Us7TCgY/l9Ct58IzDPjI2zj0l5FMDS0mWPuITUZPzsri3tjRf3jP
geBlt/dNS+Yk0YN1ZI822QJBxcXQOeapZ8lg46vSoOk4jcVUldxBzbYcTrTg5dhc1kx+6OsoS4UB
sJ5GbVuDEduARem/1lhj+XTD4Oe3HZjw+Q2OEgiM3yIdC7Hj9aweXAokM4GYVHxYcWWnF/cqi+L2
0ZblTzw2+F9FC/8uhx0zqdEWtb26Gf0EUZ/t+MktRvVvuLwdY1Tc+QE1YdVP+sQJypcmjTrvHjU1
0MyLQtgqRGNafbtde04bWVDI0YJB/Eqsaj1np3nkNfVoF6wsxxk6fimH7QlAqEVbEAYzuwyAHxtb
aLT9jICSogJj34G5KA2V7nM1kE2WrsnGkq+O9jiINP2AGeRuZNY9qQcfkhRZyz90G7bLCnsWHhee
q1VnVehcFKLju9NRF7Dk2cpNK0S8tuK36KXXCpuc+oRsnWWAUL6RZTAXX3IqtTvkLJQirakyhrju
yFb74Vp/giU3ahseWmMFItUAjEidIkVMIdSvG37refcaFGlXZIGh4qfGgXEnsm0tng+yxvEl8BKN
c+4gPIMBMaQnwPb4S0vsTNLWJb0DIHgFMen5njPe+BGQmFUFwxqnObJbAGwb4shBiEX7JNcla08C
kXetvudIVBR/X49D7wMQC0fW1bm77btcHzG4FVwNyak2YhjcDZMyus05iMkkA0cgJnd+sRNMCOWP
pj9+5zTb/3vB8FeQW0cC8PHfl+VvnMKFe8BbVBAqkR3rqXVreN4sxK+VNneBE1xkEq0nZowlcYiO
iAUIY8XAybL39ydyETzAzuiL/V0SFn/rSJ3hQwPNrxOQcaAUezVXvHy3e6K/6A1DqLeN6cDAzaE9
aAJBrr6p3oCRU8ZQwPwqxJoISpAykwizITjPDma5FSS0OzoDqnUtL6y/CtFFhnnOXozoJx5CzTmg
v0RSiND0fNORUkXLlfd/eYxiZv8HH/eGN8CRM48gL90r5LS+4Ak1XkRhEW3jbBm8ZMZ2+7rXrNNf
ZMXABGMs53rs/q7FTqfNgfEWptFBybJi/2ryt7SOLP94+v7OXSNJOz2OL5FgcE7nMkUbh5pidRvB
i+7LGgBQFmLKZqNJvx7k2xlPE9mnudm14ZLrtJWgpMVQhlybetA0ew/6tBOUNBKYKzRfgpGBeD1g
L7gEj+MrLOLwGca4ROFAlsJTgMJz/+iw50G55/D4tfhS/lqLl4CHrwJ0rIyk3XHAJYK31blx8QtQ
WQ5UkeYix10T2aWZpQ5J7DlX+EAmLoQsQIP5oTKeg0vpRPqaR9xITYJCChmr53XQG+APaE1rCpKd
yHcQw1K5b92Tx7OXGvmqRU8qsAWh97+R9281/tDRK2xj8GrTMxmdwdi7KpdXLAvbye/1QCh4H5eb
cGLzBJcoBYlgzqKL7pDWnX4CqGz9qs5Yam5tb+cajfl0hgff9xieehbTd2JOESV3L4K3wRwja+KC
ta4Fa/Ta2d9wbml9L1d3hnn8fBm2+AwgEObemrNhKHP7RefO5JmSj4A4gKyZ87wRyTba+M9ZLLge
PljrZeNeosfqy5t+hLq2Zr8SM4y03NRWkIgZc8fmPqsRq4NOJg06kn0ZoyIOoTFAj9QXEx8a5DGh
wX+nc2AI8jt1ierygEVKUVgnTf0DplP+1Mv+OwFzlaab+rYEkKnEL5niIiecfZFQ5QBLEy3fkbhN
L3IdGwlNI69pTIhHkLYmlBtrvOocYzLTNaGwKN46+czHWoyFKGC97q+va2n3i9aRJUU53WrGAxg8
azORXgL4BuTzEWY+XZtcBC/jEVIGurm5eNDOqW15dbG4zdnpcEzr+T6OT24SE3rjggpgDHRImGSj
LY42/LKyCCD0ovUyMoSkIn32i98HvfDjIFw08Z14Lgv+gqAz5hOZG65MIlBXG1JyDaJ1m770lQB8
mQaQPTEBUZ2QKmPctFNUwCAMGD2O0Gp75ge+dZT9aP74V/XHuebUgN0a2qQ+O1a8xOHD/fAozdRW
wz6NhKxJ50VjI29hLiFNgFgpaZP9lBdjEdf0lLkNyneNYPrl7w7LysxfN/+kQGzNE0nBxsfgCqUu
k+ccIxSeVuKJdgsn6hu3shLMdK3kHPrQJFvWwlzjGtd9etJcpe6dTZgWW8n3z4548VLtCp4I5OSo
hksTL25XoGh/EzwwMgyZEn9nBx2mKTHfpuHbX+Tq6uMYyPS/UqkOGK1I8ioreh8YMKWF/+rVUa3t
sC9fi9i4UolIByIgVpODba6ZHznojz4q/2ncHWc6rrt9sU6I8qaEHyrtt4oWrFUK8MxvVBnXePJm
39HBdgtRYXSdeUDcJRedbERhgR4u9NCSrmVQ7i8WE28ddwkDUo9ndKYeexo5LcbClrQvGC9v7atu
jcXfNIz/IguCiGZzKdLNRT/Lx19HmapHp8vOE68D6zzTlST6qTWgeEW3WrlCp19ONPRdcAC+/9fT
mRgM6GSg/lzAmh6M58hAv9XgR6oh0K8VfrigdBRYgXyAYqtobBz3hYYtPDvYCfMfei1BFAfANd/w
Bw6EjeCTVISr6ei0cwpbpCNzQi9hFTCDvlj284Y/ahtkzIWR29FG+FMX+jd1iQnP3ZsD8XKEz2Kx
ny+qLhhypsolvN4JaV+vg05Oi93vuxQov2QZbre6OjVqPbP1CUjHffgKgfbAeS2drVvywmUDlMyL
D20rwEFnfpPbRo3vM4I5ZUKEj1fymdXnpkNiiwSTbVaG/fh8vH61A670w4NtArSEFghSu3+Rr+sK
SKEB9MD2lA9BYEirT2dmST0/mFrmR35Ym2RnUJIf+zYxMoKVAlUpnPW4MKQT9f8iltwybG3UgqON
EgMmbf/CxjVKrZEUGTCdrmWYt3xJFqlSsxXbFIGb9z/BdBZ4XnL9cvpbthCgGMqkkSIMZppSSxnB
nbwX/odmwbK6nutvR5D17lcGa8SE4Mv2a7VajjhZnNpaqmKNm3ShCYk2qFm2tjMfY1XqDB1HioTW
Q8xyYZQt+V5e4hpz7XVzI6D6lZ0rFteNTpuhN4+P4VVjTDSxlhKLMcvvHvjwYEPFiuOwm/9i72kW
dR3/bMK0c9RhkRuH/6sh765giQQMep19XPgRgLiAFQuP9tGvA4kExVtq2iwkJHicxFtffFlCsCMP
ImVIsdJ8fBwYeMcreYd8fjqsdFRE8jZnwyYVgbLxz+X4PtuDPr5pa13BXFU6Gc6RHwGeA6BFom/b
mVjcVDl1UN+AO0puAVUi3qktQFCUIvQquBz9qU0/NUtAnrXMCA/1zw002cnlvGkZ7LgbcIP6CoBf
LBK7KJmWRvHpEzYE+qnIIsapKcTGcxLsUlPtKhVQQrN2ZSw5HSo5AcmKHqSM3h6jbv7sOimIRh5U
DHbCOtUSGvbb86x7jnVxeWEa8aUvQcKkz5YcSD2nDvzSD3gRRbwMtYf4UbTigeCMLGRYfQAMU5hh
uBlQDuuUlUq9mHgkaqdalFXHPJ+sH1g0P1UF+hVSNIEwSE/Gkfqe7uCe9nvlt2bNLv9N4I7GRbAp
MKdPJxPDGpatOB2b8TTUEtErDXFPHUj30t18t87NS4oSefnhRg6WQce524wc/xGuqgHsyhP1E324
UxU04sqFv06hSOESqufr/GfSuBJap6ilxCz67hQBIVU/r8bURHuyXo/jigXq6v3JghNAXJTfUZWh
o1IS9LPpmrPBVLjOobbJvJ97Bk4N9TBFAahShMQgN6IVgEn4C4UlIDFG1H779Ykp+raD4CL+2S7D
Whvim5IXIFMMWaNzNUg4q7w/x1gpr2v/DEUFFMyqty5efK5m+BI8KYc7A1Fb8M17AQpReHWM3uIF
sVWXd8SCEpTLv5JIrNd3S4x36a/LfL5fFvUuyQKLBuI+tvCgr7qQgEbq8zSQlAFHNxr1Zpyo0qH3
mZffd4unbK0VKQJyO0XiNjZQBTwIl9h3EP4D9WgGcuw6YcGH6Kz2rq3vCNsmv5CNNEz3lR3qTpja
rAWztiqkp9NqGdwBoP+PDUVDykKKS/UKEQMzotzzKohIo4xScYRf5DufQmSWEce+clTD1+5eP9Ba
nP54uSm5prONALEo8BR0HSJIz+NcfZNo7obK1BprZtDYE2WcJDtwVFXsmb8kYqiEufw5E+nxGPmO
yuW435kQDYVRpsEVIdxBjYRz6jWmwbrMJvbyIoCqD6vS+Psda4p1Y6KYt42gceB+zWqbXMxEcpzy
0rZsa5m6Ew+ssLNLDvV9lfpF+A0L2m/jbqpA7acLwQQPHDbDH0dUQNqkoB8M1Yhi+/14IIpTq2ke
J+0fj9MEKc+8b9El93V6s32H0a/zTOoLIkdTUMcH5rpCJhEqkOLg85vpJ65MRbd4HE+W2MILerwG
qZtiN33ftB1INT+R1bnJ9y7MJPQ9IR5hjXhCzRGkuYgQJ4Z8DwyBZyw17jGbYH2rBNc9DuWOWMty
yoFUrJjsVpqKk1wef1CXSFoRzPk8dfBnMKHfdJoKCShgTK0nxLVbDH8STFgpEjA3B3tfreoHn8Fo
V9iN9oiTUmHV8CnRBDHQ0n4za5vjBBQfVEbP/wtX1OhDSrHngJObjpS7WMhGf/xl5muEhPMotXnl
WPQrKHVeqb69mt6kyyRsPEA7770lyAU81zk3ZLdpYp/hCwEACIHNI+VW0V74RYdVBfGl6ERMy/XF
jet5N23ujZxwzySwo2PWSF9P9kYmX4nXQQoaa18TT/+EcgdfZL3tjwrFxhHbW/32jV3sDp30MiJ5
Sl45hY4SyUoYwTh05opm4RnRDjPqizsuNJ8yJgdrWRz8unCNCWBa5CyD+ANmuy60gjTz/1YIaNJ7
ZBiiYAb+5EttPNmQuRcdSRwCwyyZGtJPWwdeUjzPzjJUz6rwHfZkhiRQQR0r1o36FsbtJWzVJBCE
n6qEp7IzR3joOyy9FPO7YEPZntfDkcyAd52M4Uyb67OX/tyZu4pZYCYIRrmoyTO8tOhXtqpCgHZJ
ec0fvjj2XdZg1x8+NfHjMyi9VD7C1u2BQuwC1HKeavlfwqpZjQ1bNWvE1hsbs/+75g2pHAxbiwEG
ML7Q842iQoRfJ39OrwzziLATrgcqLqbURiNnYOlhRo6OfBt+udmvrewXTeuJ41WtdN6Zsdszabgx
u1VyobTRihmG9m7Dbo4pLQLKBLXRaaLd8eSTFDxQi5mvhnKxWBiqXMIddG0jcCGB+d5CVbZYgqYX
+qY2wNLCCdy0e0JV4L6N/o65xd2jaOoo0tcymnypEG6gdOAoHN1Q+CI9zEFMOcsGU/plbrPCiPCC
0sbqqIQ6uZJDC9XSODFYBJMsmU9cgFlBGM5mXvHNXFFN9TjTaaaUGtIYX+oCrW7RyOBae+sjdQvf
BgydPrPgYkBymTWybyczadnQ2dSwyLhkbkn8YaCjYekBClUnqhjZ1EcvToaDQ4iO90cE/bcWoOJ2
EvfaLCNV+BN1TOhtqEiy8xiktRqBrdKAeqYsRK+k1fSmue56PiaM6KPdcHPFwCtXJiCdwvwdyVvX
OKYc3bY0LUPxqDyqXCTc/S5oaQ6V/iSqC7xCw4l8CnHrYchFKacwlxMQFIe19CIVQ/0/1VWfy48O
Z3PhoLmlVeN2V8Q7RWVCHtzyNFDglGTdd2nnPbo3NowxbgXgS1v1HUa5VF3tp2C/91wjt6X4xtH7
CzCjmgUg1Gf3TOB5cYxLVwSmUi0O4ZWlwL+M/uHb43gex6b102M/59MKrIilOJweW7RHRd7RtV8v
fnIu6F5vpTSdMUyaznZ+ekUrWLiZDRpcEBhrGzaHQqpJFmT/UVWz0kioRE5hemejPJ+Sj3i536mb
jMMUZz6N7TmaaL5938fiVzgrM5+GrxGf3HYboQvDgz8I4sI6Se5QPd8or3k1/SBuHdEz82sIYT17
WkoePj3+oLtn9bzmyDvzgejydCQV1Fk6nktCrDRjkZ41rup6gDbQWJr0rAyFyNhJA7zWxNCOQGq4
28fN4msky/dUgX4wdAMWolY+ERrrMz01bua5c/VyAytsG4KXjIvXaWjyoUPHaBRbC31n3IZz7rtG
yFkKKZOTgEomqp+tb6x2yN3aOHEUg7EoWmDgdeakKisvC7yty9AQGdrD5S4uhd1XHRDL8pq8D52m
KUDUCQF+WLlgkbGOQ40QNL5pE8rjxS3shZVB5uNjGW5eNvt7/StAkyleN652MQctYc7D9A9QSfNp
CAF7u03kzw40TvueXSy5nM9g2wZapOhD8HmtdRvSGfPm+BWla1rVAp/2hCawDw1sOzFPfzC42mYb
ZoQl7W2PtawrWEvbPeyC1E2GzHCiwA9+CrFvZCVe5W2rk67XR287yWrdXujejTLGDMVj3z0Aunzt
TGicCM4QakCfuN3A4ovbZYiTsyo8P+zfFMLjyMdohXaKxct9WJ9G/tQoWtNR+R6j5FfFT6n94w4L
3ZmSGqJ+QhjMu2KjRLaPmoSKhHcy1rkJm+kz417+zKhvbFbEnVKBiaudNpj+i6ZG+oirHCQF81Fo
z321EIiUdrRwW9uYNbXq1yEJ2lVWZECW/205hqK/EYfuOw6TYMurFTMDpuJbiya9+IyL/elV3lmi
L3Ix7m8VvKLYbJ8rouPhKN7795qvLuJLbLQJHg8h2kKMCbJM/RSkH0DdGYh/gzRZmC7VIX6jXvtc
4QqN4CEQ5Xq4r1vwLAZk2G3dJ+calPuThYd7aUxoHYDjxSOIKDtJO4ffiB9lIsuiXDbLjAGcD0xv
bC3LI5o52cbPWneX7iuBi49OPP1XbihpO4Yc2lGZ9c2AsNhNXuTUJP8PDCYhaXiHaPZJA3a57/0a
zr/peojgWeghLU+LpEaBxsNpXZ7ZaKFDG9GAcH5UM7MvUb6hCQ2wMNpc9wkc810UyW+ryTYUlkPl
y8fMLFip2OQDF1H+BTHPuk0VdFTMPJtUGl0l456kgI53fIXxTeHKe44wnBX4oIPyeW7kVm2lE57R
0CMefiwjgi6tim08/lqiKHNlFM+IVeHlK2rbAIW8CgWeBc6wglx68uweeLE2+QRg+cKhdFMfck/t
siMfep1OmURvfOeb2sqJwti/0K3pzUQDBaAp2M9rQ4a57eSfGZWMoV+8hYt9hEs7U1CBc3rTsOMl
Q/b0XElPfxEH/EBk1pu/tNVPjznsMEXBl+uu1mQaPrlv3RpUEKRUurkxW0N/F8Y3V4YBzQq5o9je
PQK3Y41NS+51i0knVQjgWYJ5ZPNQxa2jETyPRIGMylvjqWv/7Xtj81iTU2oZa20VE8SSKsfN6pQt
+zPjf2kZ+zS1DTdENdq5s5BAzGyKsXcVBKQegLLrjFXEgXqlz1NO/JF+Svj5WJrdaqZcLhmrsh+b
7gaL30ubWlY9a2j2y4KgeR/USafW24XvbTvPdcFb9U5TcycH19IQdlJXucy3v+8PV1pNkye874zI
cl9sKUNzDhxG1EkzEzoNzjRDfqqDIGgAHVuNetqqeAnhrfCl36ttX3htzqA7joaOS5wNr8VAVv29
Ks5KlRRiFT7UIIHNOtOijAcCpgzIbwbP803734S1Ab7BGfXyaJZdQ9fOW4unXDT7EEvjl6JzukX1
6WNAJDq0XtUHk17AWJq/JnsokfVRUtmxIPbriIVCW8VLTtHLB2pzbP/5rjXuhtrcLR7L81h+aH1x
RrFKAUW6qBj/p9ypB1AHhhDPTl3twWujUXJRPANKpIiJ7Sgnc11EkHnBErY2KBZKw66ZUyqwmvYr
S1/MFA2Qo0BF6CIagyo2eiLa5o84LXdEa5cIgaxGKSm1LLBTw5D9FTdg/oOeefr8OZBE1HH9W36T
8r7WisHO4syF0O6xHbtzjaaM8WHqapPRPLT28+KMbCEDHDf4USJdLJJRJL0zHY3S1ivUZ2hOYSq7
IGtT5mOFIkA/BW02gO6/KUbkrQ7qrz5sTA5smtgbQ4CHDP+agzn4Ppz0zRdvi4z+INfK04/tTX3I
erH10bsWdLLnXoJXqd1XvLsC9vMTeNdotLIWsxyc0c/O/JBx91RJ2/E6J+ijykN87xhTUycRCA4c
i5VMuf61SBPjkiujUKJyZbFxDXhk6GkC5GiZzVRG+wT74ahe63NEbiumtcxhv7c0So6tMF6+wPRE
l0RuxM2ZCvDll82T17uZonuLubWuT0kAC+HowTL4efH0Hx7BdCHKQ4KI/yRGOrfUNkBhIsFYUGz/
jwbVKGES2rsOvOMvYelm0RYZwZQtyl3WLBXomW3X6mPUXBJeMCCCISPFb9KI00NlZYt5fTbwGewM
FQkdVFIh1Tp18GyOvg8vw3/PmXLJ+iguqMmiMvjBUMzkOIERH6qxwOuKLS716Ughx90apbFK4CN2
eoF25FxXMWT++Re2PVpF88en/nRGy/gnR7FQpl6zpbsxk0RlyCS5kp5Apx+pPE/CD3rtua9liLfo
YztJkaq1dxGLKnXWh0GURdxybOzyb7m5ZHovsfv8QY27Ao5lJwXS1P6uJDqsh/e69DRn0An5Vk5X
nrvb4+X0K/aOvneJmALNUKD+nNJLYd0uerQta0KVWHeGc2LjQN4L2/UstpTQtrIRtxGABeI80I8a
MOdCJNV5k5pfCoA4JHiZ2aKA5kbFm6B1Aym6V81UniJTUmb74LT/rknv0GrsU/sZf0xYdiBihMKB
y6nzb8lvl0GgFqv5V+gKjyGFgjEe4803Yvb8NJNUFXfBLI69AjyUK2bmM+H2HLMQFoY9l3DJIR1d
i1Cta4aXmH0bgH2wfU6VG2buGPCYaWTMyOfj4oHpcEKVn4GdZ7AozWLi9Kp6Tmq3NbzdYlwjKsI9
u7uJL/iG6wJJJgUVfZlWPWHtledSQ8okdMjP8zLFJOfagl3q/kgO3mkrOLfNOJ/eSDpsvx6hkoVs
rrou0Ifx49SuLZiFf/4v2I7rJAu9dNHN7vxAlczRd8B4ay14N/hTIfKlbEeMpPoHYlI4cDX9Ojt1
cHop5K5sWgto624NxHJ1T72Rpm0B+IzTbNUmbt/RrrtoOZd7d3xfmsXYWPAtZwhiBOo9iTDokmdR
vYJXwuwrQ/PKIUaFgaQteuoEtr7kPlZk4KMznPfIuqiWAfpNgaMYHkqSsgjgXWHKr76Y2hxTItj/
F1pVQxUwRGaAVzjJ6szIuGm1BJ4+bnQ2HuxO4v9pYO3+c7e9ZILE+Ultc5Y6u0LwgieRM2XnLCsO
UGdjuLP/MLfE7KmueKqOBup4dMq4GEF/5yD5gi8fydagh5AkKsQi8xwkdR+sLz0rXxSFIV4b5JZj
3UfGNvLWkAkgg1RO2SKSIC8w0cHjepwTsPAr3bI43hQ2THlL1YIm4NZNjPWPGORs1pIYojnIqmMr
sMYyQZ6mZSytPoSv52h8CqkTJKP7xeUwKh6mj1VOda7R2r55DjEt+kzjigtB2yS8VYFFrJ78Y1US
VoA/Ws1mAEe2YhNZEPga1IO4tibK9kZ7xI97qwxjDvho3YDPfTy/a+WJoOHiXj7ie07Uo7CwILg+
529N++xHSn3aPBY4liyP7TE6cW1PXnvx1Gk2A5AHQ/YzCuCo9KJ2ZyALT/kwlZ8Bhb105jVgH4zO
XEORCt5DJ4Irt1ogoNXR+TJoVjdx3dQ8C87S27tH6CnFoMpOn4duzxnh1rYixIqVUFfToUC5UfOc
9dUlcCWsyV+MWvuDkMjSq620AuqZsdqiq19BJaJge3r4aDV+PIf3JyikPYKbzdzG/gfU62ksPS3o
a+krLe5dZB/Vt7ASe+bP12hgR4T9xoCqjbst+ohk+lBHI3x7CyGuYatV1lyS0rXTZbZ044ZXnr9q
aBC6F0ccTiUlAyjPzKirE8lu8724PLrtu4nHup9v9tcXjy9YNeFvV4MQY+/8pK2ESxyIGFxanWQX
9g8GputmfrIcf3NQSDoXavM9kI2048o8y5rZ4HwmuReIBdASDaNo0uO77bZH5lg0+6dfJVA/RsAm
NwjD3FhyhmRf3n9fZCi5Cvf0zPN5lDbfWYsbSMtJ/OQxUIn4joxQNQFlwENko/QIO/dmtHuBCVoI
4rtm4qY3kefJKOiW0e5lEjn2GjVmclZIpuZIUJh7flStrsv8yTq6SJDvKls2PKPyKSdcCuil4wo2
5pwOEF8oDXToH1coU2ykxPsa4R36LDexRgesryoX+YuG704R8tpcwWAE6Q8ZYm+RgkLGHVnXPDDs
cknIS8SJ5Z0g98J+uuYAqQcfoPdp2n0ts+X4NfagA6/IpQKCYN8mLsGLoJQ6CwCOGwmOoZWaHS7l
iWTILdXBH+aEABaGW+vjvtYnUVhwtHi9OTZdpPf06dumhIOpGShvmPge0zXmAqadp5PF3Hyja+6g
+I8yf75DAwNFPyV6yAZubNuUXpWf4s1DaOXov0kkqcEuiqCsj8Dk+5QPKKX9K3igWaCUrPG59UlT
QEcilttX8/RHVqyp0gMqDwQVBHXl/Lu0nk4zyZR2g9AKsTJ5x8G2zooSHdrV2jCz+16uVkGRp6NN
XCF0R7SSH7jRoyy5kH+FZ+nrGn21UxjygGKGeNUK/St0i8C9KgFE4w9xJamTzEVeEKWtC0uQalsl
y6H/0OOK6CiS5bDuueKgY0Ppqj58VkEbzABNRFvfzAyDKPacaYW1EBuqBWNr2M5wxrh0eVwuQbfx
BOWcxoJF1wfK2Zefb57Ip6K8CF89D+8tgUThyEMY5Yx7xxHXRPbNydV/TmKnQsddDfDVlVgjiDrc
czADtUuIZNtXAlsImJZ6vwVUXLaOMDYogMfbPiaJmvKKtF2OmzlEbyP4xUQ+NP+U0FpoWIbj4BOi
NM4YmWxsF87oQoaePMdUgp928mVDPrmygIDMmvRdx2/braHEMWMyBUuWc2FpbQvb39ChlOHkt2jI
TZ4P2sm651/CZWw/Q83QU19RsaYOoKxGiOhn1oFsEoKyo9xMjik5kgasoN78c7/Jbr2d9Kg4M1Ki
LYJtIhTj8vHEqdZkNGiIhUSv7mfP6wSC1Myr+XRSj5Ye8/YWavarLvdtNqYGmVqkXhdn1hAd2Cvl
iFUUOHPTlLcmpzu4lA1SXcYN+MBXEJ9/c83ouCqnJxPY18ac2I2L1VzmFUWamJJzeWv6mLj55zpK
O7A/UFNBDY2wS/kfs/wb1jntk7RKmtSDtCh4J+sQ2pAvLOj2tU3QsjCLAoXTTm+cmiQEjmzIyyuJ
jxGpAeB3sVos6oFbKWBDZxeEgbUqe1bqz6jdAvdj1HUMxdbI5OfKxu72Gh+jl4qaeFKRhOGJLZ+j
6vdFdXN9Fd5mFUgDNyZtv/VU3bSrG3Fz0zwRWLysflyL7eGov+FaQsba85NaDh8emr2KG9AxbC6x
CqxR9lwcHYmDVom1C56rxYUzdPpMEzXnOUUG599XXmwB2nC3ozPqtABIa0I3a8KfXHF4FKCGzxjy
4KZlLZzQBwAlIcpqsEFYzONXVH546AO6mAQTskrH30By62rTr8hWO+TIODolTVFcpVzKewi4w/GB
eDWoGnI/a/mXVBO1tuuVj7eQV9ULXezHv3so+v3b0+Qps79QGv1jknXAbaR89Bs0tRVIhI86Jrxy
U/qCdjeX7zEU7D0lJ82bikITWddV+estVK9bR7d/NHY+ckR3SJRFkB9QSTR5EyySXRAUW9xQe/QG
OadBEqP7zxxmadWOHwfmmCXnWRl48ZRORrI+DH3S2kS6l+4TxCpHdQ+379G45p4ox+4vgjOn/wyG
VlkoLGXLZp+uJSbcUj1lH9fmePLvnJ+AYdgyndrmUc6h7lv51ctFmodRw1DCmm5Ro3NT83nHi09f
NFhSeF3Lzu4tSZAgXwgNNTgQypfm6z5OTNwhSoWAYncPWvpR/Jkc49/ttTf3fxrcyO1oS5ICc8i2
eWnVtU/n6r7oy4ClqYcGxyGHZe2D9XL+/gMm/Kw0U+mOM/RPfCK7i5j6OYgLjMM0/gCUHXxVjGLE
sUA3UeT5sQndPeq5IdtBeUuTb43PTRbDSvlDFnc+4ymkIpv6Yf/y9vfsKjClYcI4lWg+8HFnbnX1
94w5LUa1npsmee1GOPLtGN5EV6isEXBCgwGpmTmDDXgq7ysI99HZg2o2mKEsVj3pPb+Vq2+acRTX
YAx946rXH+6wt3MoTAUJoC121CvMOM5S9LTuI9ZXkVyTZR6MY4wVA0IUxZwsxrC38xW3VPMF0btN
H1zbgjVN6rDkhyvNfRh5bcIANB0yrZyu1HEc9hPRDW2VEncegi8j5W88tgugfHX3w2wO2CnEm7+K
fjec7prkNVOHh/dky5+nClkW4RI73i9eVo2335vMVkY3tBCSIqqw3FLDXomX6avqNk67atGtJ9b0
7qn89Bp2AsvhvI2HkY0IMFQDEZCs/JHb7yUkVdA8dffUs/jo5qkLouw/iti1h200zCv6C0MDp63C
GAPOXdTMVhhCA/CPx3lPLfesbX95mMqsqa0yEHuNtqMn0Z99gH/vf4d41UrP8sg3xb+BXgCUW/nT
4WMdwVRWli2/muw2+vQ5GGQ5KNcy8lODoro+dC0PqlkvGaVdFgm98fhpIx5jxRhp9ANr0bGewHC9
x+ACvj7eFCz6uQ/jQov4ssQ/MOuk3e0NB3eAl/1VaHLJuk+NOK/uNy9sCeitUyx0LiMkltO6DN6C
A8ihBCqLmPlUTnns9s+0haU5UhsXFs+kdKfIKXszeCJ/4bX9rUlLhvwH4DT8SeD05gAX31Fp63lP
Rrv9g4Azl3l95xU4f5YItHBDIRWqvGARhvac8kbwXxun/+z7PaUAmxkn5Kpvt04Ba2UfLd9Fj73B
Pbcz2JzWUnF3uPVB/hNgVzZv60e/lPVzZB+hbox+krI4h7WXUwMSNUSqtTftR97iDWpC5sGnHaA7
blqdXg1DWrwmjIf4YA5muh7fAi5lwkuyQAi33Bl+7zUQ3muPO08cQJ2S3sEq1f54NOfM3qYf4ttl
AIKrRERLUigtloXWkstW4nSpmfOG5cWoKA/MCuakMltgMKmLovSh2MjhpXOV2Rw7eVAasOz3c+g1
Z8YgoYAh5QYaD9sgBpg8qvGcNzv6D9tilvR1dUnUkUCj40Fq/Jr3Oqvnv3OJn1LIZC+5Nogt52WP
KEBhALhoE6AQqEXgcSDoA6igBZQkH6oa7B3GgEiH+MTEhaCtMfMUXa3+GiWjTRV1RvOYimK3jGG7
ky9nO/035ViAmyYtgG0GrjmXyv5fzSzBsCmB8U8loYQO5cuIjph73It66bRqYpxi/4N3jXkdIod3
bDKz/MqUfwIgsrPs5T4S3K9NPMU0m3A2W72YKgkYlBCSZQ0/a7VFI0V8SPHeA4cri9MuSoYMLStN
N10jB0mdK3YtsaUNGipTcZo5gJVwXzo9j7RJe+eT3OFYqQMLpn5i4DE1a20I3G2UJuqEIqL+X8AY
eE1Uvyo3S8PMLHMWubILU26GaO36CXX6GgkdiaGbg6PrQYBNPACEZ5en8JWicS8KH8euQDJg13nM
nFMICEMtAAaHDW+1sAStje60g0YbNxu21EwSccj2QNGTHDa45k5rcWDq3BFHxBOD9TTUeGjRUgqr
Vhd59FsLEVLXKQLz7BASOwd3IJ54qKAlcLuWF6TPA1j2cbHuDVYRvxViKWRzZAduLIxTGO4RJxsA
NZnzVWWSR2a24EhrbeU4gAiqxZwaOv1dqgfUKSxlXWzpSr6LFctAq4qxjK4X93DwhdLQCYufxfn0
sz0lfnZOkEX8iMKrqP0eeBIh54GqrEUbGtF0jNUoiVvabTTjTNJEY4wNL3UZmGDPJLA24F0gYNNF
IgdSP3FBEwz3Tv4rjraaEt+tSFs6xdJRAxa1MabfjK0eI86neE6TpjpHwA76awV05aJ/zhSelR95
NnWuR+mmX5R/Jim0NAeQSzyu6w2C3gqtDW/SO4Fa7plnPRntr5ybVwQaNAAC8Rge50V+pGRUcO7F
NKAHI5IbjiBwL69bQKaVpxD/o8o1f3qXCsM4DnwZULkp33cPZuit5574YEj7BXeWrxXgHLRX+Oqi
Pu+Aq+nouzcwNEHmnivi8RGW7nJTVTfNUpk7AZgsZrQebjWstnZ9AURFJzuZ1CvgruntTjxviv9b
JWljIHtxCm/qxql+7RZJpzRWJzSyvPPWRQ9CCO3o7lNrzbcLUu8+DqMwAzbv7JELtrw1Q2eW2Tlo
wiSCRDk2+IJ+dB8NyCWjN2eOxrCfWDXFoBZntLscbmS6O6Uzr6hTmPhYgLY9g8Opv9PKMAy5TUbf
WUUFGk0EBoY0WJExeqFJpE+NjZzr+Q83w6C5zdA2rJsmmCClkO5RS0DkBBabg9ONJdZ2Drl3ME1+
s/IWU7SMEbEWXfEUnvWi0jHF7GIxWcecjBazwLSKK+6baX/MRDXIxj2egyCX6wtcxcj/7QBrDcFR
naJclMaUaG567/1hOtX168mFb0q7jI14b6qlh2ES8JBcc48yjo7vsq4DtVayklL7JT4HQw+m5vCI
Dros3ZviCo+pYbeopbvvlQsjylb0kh4BPB9n/Stfn5UXuWmbDQ9V2vaWcGUN4Z1YQ/lB0suVG1SH
YkYtJ4ye+dcQvI3J+m1x5u1F2tdpHGbPpjoHOXGBfy33uxPJp7wdcKL9qgTWQp4aicKKSrH/R1C4
ht9HmiNT3Wij5qAtaDx0aCsBOUl9kgnSWvWZqk08fDZRETANPuAfQAXlUPMw7GRCSFpTCK5+3HKZ
inXwKzwpcqGdePL95iQdPQWxHadLRWMobDc5/PeMpbC9zcYa0JMHYHNLhPsRwsEer8/6QRQM+JIx
OVBpdafRIlqDUarp4CXIjVRq8xfdSrv/vTSv4zzEoYIs2sowUB6/murcmez+YBN6mPJ/xniTYDuN
jB0PQVUBHvT54Gi2I4795ZlVDZqi+GMmwv5k1ruI65p+U64V6N6AmejAE3U0a3PKsmLUFzaIa3ky
KMGCSdJ4I6uaxZ2uVmvtMJVsRDPPA5mnXNa/hrxeFi0RuF/9TVZyYmyRqmeUwIcOYk9ZfezC7PJ2
HoRTN8DYk7l3ajx0z+soPdQjVbmd3JGAqhbthWIUVUqLjjk+xFbVco7MeDKF0KLQA7ag5cHnYcpJ
fyn5u5thgJx/I4njAtuH9VeZRuuSWIiv0p5M5/gUKCVgGIwYx6IXl3dGKpbfVV8Vrb8Sof3kjegB
y7W6kpaeM+JvWQSZKlCktYazBCMf7v6qHnaFtddVyNaRHF5/N82TPa/G5O0N5VAQ66yGABGVrBwp
5YnjNRbkKauWvmNnnNehi68qOkeusoDx67TLZhN1TRBVjv+R77GjwzuZRtYFFhJGuJLpVIQAUyor
x8QfNTMxUEEHHor/2r9pMFN8ju6ljMS2+lprimHfJlGzbGr1iMY2CBmfpUCwR4fsXUYt/wOshi23
Cvwx8WZwGPRwzR8gAQlxVB5A0XXiyxAB7SCKJQmzuOtozwF4kYzzhMN0mwv2yzOyyYMZa+ZhiDbw
ZhqUjnpE3H43qWCkPUaPDwIWqL+pYqQ8KQa/07U8SXirL5G3BpYFKHq1aDSnPZb6bT/l96wVvb2y
kuWld/Az60QygAj01ijPOeF3UPXWh4ePaMZWo1Mmm7HgMeWJ+Z7t1vIJv0PpwKubqC9QWU6b1eih
ZDq+M2DxtrfxrNwbdrrVgZOlEi2X6mmiikrB3KPjgAxJXthLlMqRUEQiEBZFGEmj3hYYs4nplg6a
eJbwjFTmPM71agyOBsY5dxb/T2SOLAS7a1nef037OYSx3lANeRjlSflDRXNnuCdCpNtWYHGEbLha
WyzB4DMZ1Kcq2Sdsj4NK17YUWxvWbQvlKHRgGWyZyBzG9YO1DNmKc0JVI2fgCWFyMtf9WhMuVxW4
jH5mKpIlgpvnTGAA6f4zsRJQlkkl6XhHty+YGtw5yO/s2hPgkcTEOVbisJH7e1LwFfUQ9vk0aEav
aJCVpl+o4vHpCwHNibs570/rraKAV0mP2RxfFLdCytuvBiOpeQBbDq7Y3KlYG8PNnnF9Fxt8ed+z
dex2zzVJOPXire68KhvyHi1yq10tek9dxNIsxIRT++Hjp0NNXbn5dWykME2GD5PnAWzv7wUmzVaq
Z+z6WJ6DdJOMXjO9c7wBOlnpp+TGfKMdClosRPq3xhYUkqbiwSpiam5mwsKMJ+g9l3d0/BZ1wRSq
j3oRLTe7WmH3lm3EuihXyNjxEv3AGQdxhD63WRRwB92kBClv3Qchj02/Z28IvSvjA1tCWqlTXcjf
jTgTby4JONiPXcF6u6QkjHBQ30e/5/TKJFRZiTzqX8KhM34hq0Uqkn9XbVDAJ8ve8Oo4dJqR4Y08
1SQM6a5G86CxigHqBdsj3kxCy2K3nRXjP3mxx9SIUbA/yQ9jxBnYqNsSsZAXmLERiJRxYfM3EHMJ
kfbRTnQag776NPnpFodHb2aS3tPvbjJ2xZUgIQ3Zxpyn7wlKzJvuUCZtJurJTDy1S8NXDHSA2zv5
+0dAFrc9FGB00uZcODUPV3ecOEuLNgtuYYZXfE//3aBJ07g+tSh0pttP9D7ScEC/UgL8O432MMCN
aRKwHlkqvp6DU6sOPr041D6EIGnW5ozfFEzaC1/oGvE4AMR83yQYtxKt/4bX1QmAshC+x6gF2JxP
g5le1k6r1cCSNQXAg+EHGEz2/RbN4yQrAowCjpCPdDSXQGqLfy7QFJgk4uUNxObmf63j5VxGShua
T1dBHpVxo6xNhShsCxPUKfdKaKviDbIzVmFBl7RLctR5sy72ufHl7c7GprbfE2Lakg/GrxRI2F35
DqTW6ru1gTuHM6UqU3h2kof8ok0IDYPMWgG3345GBs2UnDVHAYoew/TZvSGoFfscbUEZjqAmdBnQ
2Al5V2mZeFvYBElLGA7P0IrN0z+DXj4rp1IxhvRzAfARKT4rVBj1J4cSHhdVq9WvGsMMG2Wq5sHj
LnK0PoNcd5ZgnmfrwW3C3ViCzi7kgE+eCW2gCLfmEw4C18NowWxaGyM845mY6wWFxcbsskAE/ZDR
6P2SQ6gCRRbfR9YgD2agIMLaUZr38DYVR1KdQ9+DF7VRBmA6OzHw9BfNb1tfMeyf+nLmmEXlSR1C
Sh3+pgNV2kuBJGIMb3P4f6CPmZ3bYyHEiQg1wa1RDwrtrsg3LW1aXYv5QaPcW0UunmfBP/7LhUjH
NyKlrn6ooKexSBfT+eEF5vIMrsfQbTDLAJSl8f6PZX7vrHKCo+fi/0Xe5EPAqbShpGEEfysZPOS0
NmASvG3ro71qdzJyw51bpTcnhK1u4uZzR4Y01F8dHvK46eOeUwbWGtlGM4LEx8vWPQnEbh0HMbbC
3G7MPkHYZR88uxOrbk/rUfHNzMruZhJSAIv3fgBb1VPUT1a4UmbnYnrMD1aXv6wOLDMOa5Nukq/y
Bs/NagDelaiNAwH1AqJVMnBbzC0nHsAmMa6o5b0IoI6Jwgiqe6MU4Jw4HjCxSB3pIxCI6SKoSUFd
FyU8IK3z2s7JJnoOWJv8yMhDjY7YoFcDzsafh1wFaXXoRZL6wg6e4JqjjDuwsssJmxI6gbIWtN6F
sQYLdbs+wP15hEfl6Ci0fv7/IIs3MRqxzA/wYdIfSOAoLdO7z6NV95VH95D0deadGq9i8YrJEcyY
amYWe9GWbSfBa7gLVJlRyD82R6fcKkJa1oO4O92/oevMIb5o102YELhYLyoUQCitRadPzXyhd8GC
1oNTF9BTHhvJBo0ogoTko8D5EZVIpuugVb9LEf2aFcibgt8iw5xBCIEBUFb3Re5d3KNkpNK79SkX
4r2nrhkBCGvGmnXKYxto4loUAuN5o9slk3OjDwb6COKGM19bQL2lZQhQ8D3KbmtXW7uYnPXqvYp2
rIBXc+Y3V0awMrIDHvsGUT2k4gjJtzDzKcvzcfP5SvX6MnMrLjgfd/dDVT3VjJuW+sIS4mISMepv
6bttS34vIBtXOvAzio2ANGZ5d5E+d+AKQLs1/xF7Yjh4iOIz7/gBW1DLnMa0t224rwKa6K/+dnuM
ZgFx85g73HK7v6a8e1HxzVA8S9RPtyTZ6ubHIu6w9MQVadd6uZjzOPprHzwzssGb8Tcdq7z5Dg4P
n0xeUKxNVw0NzkXV0xYDY+b1jMY+FdIS966k5A5WFCJ5kbaE7rW0wr43dzYkGji6YCMcEG/rxd8G
ARkXV+G6VQ1inbpn3/zQpbr5o76jodv05e2LauT+87pw4JFVdV7wFuc8C3fqCujBejmsU6vEQsnG
y5KBSK+fULV9EZhnW/wjxSWORgAhDWutxeG2AVn9xKFulvkz3VEOBOGFdq+vIz/164rxHVkNIy22
hP9LcuEpqqg3E2UsIhyEbn4haQinR3ICnk4bp6xU6XEHFU+CMpvE+4o8dQncKRGkbYnvttxGl4mH
whZNN0ThaUd4pYbwNl/YDM0hjHeUd5tS1qLRJ0v1HzMSDgCeRX7DDAbMp5JrFawV09EtNzLByCK/
YXf9TiRudovUukIOXoTkSDoE8qrO66zcxJZDhzgmIDlWYzJVQ/wErV9lSc8GR/zm2eHxWcQew5zM
LC4CSHrTJ5tx06DSdeRLTmFEI9jN2ktCmfm5p7Kqs4GGKzlEY5f2P4AAPZHNlAjZTZ7vK8abGR2h
ZIej9VnvGTz6faaRDu1JTSQ7jm0QdDFicY8EFafRu7iHZyz2Jq5Q4P8BL3fGq7vr16GXZDrk8Owr
dKAgl7UYEHTnC7pTFEsFZn9ifqzwtcYu1UGzIWLNBhF9dIjjW+Yw0GnS5FvxriiSC6OlBBsAPjV0
j/wH/4fCbJNFXQufudrZlEQnMHwPEAaKOvcrqKDtdBjJ+wKQ/jLI23Ebdw3hTNJg2rkmE5m8oH6e
AHvxKS8P7Ej7ezSbN/QAtRBXWEhYPy82oaoWVnHHaKXXkhQVNW2u7ya9ZNzuO4XQgCcazvw9UqPZ
A4kGa7V23Ivjxf6lXL/GsiU4U6MbfGfq3A0Q7qyhhEQhnQp9rJgs4GCud6GPmdhT4JuL8PULvbu/
rmSclVnVJ1ckBS1EYNn4paFd0KigGlbY4CUCR7LRC8Icl6RoaqNfpxhK07BR5tMoNIMpq8CgRzoM
0cGfPHXSYGQi1dDQV/HBd8IS2jJt2BBIxFUUbsrErtJid2jinOqUIEMgGDr2d1xvjd9iWDjrMB0X
bILfcfTGfFf6uYI2aEzBCU70DxIXjzBR8gU+FiIcM31a9KfovWaFFPLgzIVdwGMmQcOUEpYmFSB4
0w9KMVpbHNQkQLF2m/mIH0ADh+kvyYXp7Yy4Pxkxwn11YpZUCndCqrtOph1KRFcW2II5NnBaDY2E
44c2z5UNLL1eaqjF7HacrPbqtglpaXB5W9gmMPrEUvM9T2N8rzGM/nEkHFJNoxg6pZFbXj03Mf2C
rL2iGCvKBLXuHkJm6C4aVs4Ng85zhVM+XCjq3h6IZsDhs0Q7C8BS15exWh5bs+Tvu8HpkOKv+W1h
GuprVlYKK8T5hQ187AbLx+rHJiumxhTESUhJOTsoIsfK5K9tNGhKO1gELK4/ldNumyv3Re9CXdXZ
BkFN81dp2oFWVOtxQEyPpJesDpB6YMLWCD4sUmDDeBe59HK0InvXMV8M47MK6zv5P247vaboaf/P
LNGTtNL0WAX3z24tbkos9bZ9OllGoMy6YeIGAJ6k5QyOOHjBowW2JeHg20HqdyuQeLVCBoDtcaFl
mzQKqO28VbdB4DcJ1qEh4zT2f4dD4nFh5S12AUyiK/Ex2qXpF+lnGW5mmCXHtJHetHs2C7aI4AvL
mDWvFS8LbriNS/hjNBgpmtu4yuABsWMf/9b6x/zI9+Nxh5IPY5rj6SDaZ/5BkkJQsBO/zWdnk2lX
up6Zh1bLlOQlASPH7/YS44xuIxH7aF0bxhIRTg9Dqk3lzDUydkkREzxD4u01oG1Y1U0AwcKftg4c
NMSdxteVnZBQ1oB1peq+Td+bCXTf7bkzMJv1gXzI2xTqMnP6NYc1yOmLEZ8i3+CtV9kCcO8+YX+y
BoD7u9lHMlz5r48uPqnjUDqbm1BsvJXfCRsSpLwlSzJ4XYmeosg7aWEUwtdw0l/1aQK86WSCocZA
b8FpWc+vICfC84Cxxd1pgn5I7YMvheZskWgxN/GFEBdAARJvik30YbN4vskV+lX4HBXqGgQ3l108
bTwqMGzo31IbdLyh/BhvmUO9xgzaDodiAdvFx5dNxLWsa8wun97GgjEwq44oZ+XqUn/JUQH86fbK
SUjo3z3XI3BVcDL6waJJ9NVc+DZ2JaKH+aQ4v2KyjJro8evGBBxg4Pd0whpdzjyrQiwrWP3jM9EH
nrRSBXjqngYclOR1R81Wwri9ya5V0YEqL22GI+1LWEPoCaZ82WAFzC8M8nEOXYdt3D6pIwcSMogu
Kjur9W2hAnGzpK4DOPuUa79D7aLXk3orDXa2mkUan8jXnakClAVcI2pZj+f+dGTpOio1qWy0Dnev
UCZR+uNnU71qwwddBBYZqhWx8RHaRB/eNnwbBtdnELnaC9EWbNTpIHHY0Mkd29h4G0OEq7GoB9ON
4A3ImyoV34vM9wnF8wColIgAEf/hZdd4O4FT7KRjpRsOTfJIwwrFSyWJgIcFOkImgQKzojcmK4Gh
PDz2gRNNhBdY5OXq3H70pYZZEyg+vepYGzxFFOopOY2dPVD7HhWPfwXP8GE6vhzWl2Lxcg2C24nN
dxKkS8NnDp7/BfZXweGUG0lGeSprKqk0qk8GEPH4biRsFVul/Nq+6dTk62O96SLurEKLN7ba+QVG
H1Gxo+wOLNGobAb09/MMmr4mfFeBwRNqcmzKuoa8Abf4r+bcxcDOFlnZw9LS5RRRyDS4H6hnLqt0
vbEe+gLUszdah16nZFaOl/bnv51FZIcRXBMly6+Mj7xAJEIpbSYBYKIO2eJMHzokDOe7WAgdlR6B
LB3qHdkcCx6o7cqURj+MtNpnSXyDcW7YQGVNVSqLQy4NDekMKNvlok25nwJmOOCGHMnog/plN+bF
hvQ5G6qUZXCX8KKkPESSISXv0CH2PQT7aFD5CyHZHPqL0aC9Q77E7bvS87Q0+CBEoYG1Rl2xsIJM
j05CZM5c0teptfMQIPzRmb793Vj6wb0J0VZLp1F1FFKPofSXmfcJHhwpco5xCCGfCnWnV4dv/pVJ
2GNOWZ75cECYbniBTYaDcADly/IoPF99FPq5biKl0x3guWKHLxSDvyRnKzBp0F8XV1Xk8lyb9oeJ
Zw6lfOo0JDk1B/5Nb3Wk/aUwgrAlq7sKobj5hr8+rqijQrWoYeNy/g1Bdr7/tL0AcuJ7moCuKcCY
k9kAy/xQiNDY6/JEX17cpmYsDy0/D+d/YdGAqdID37yBRsJAHapq3ToX9kyd5ahwpfIsxDm76YtU
MjxhfrBtVuFMl2m0u8PYvFtRUDOs1WmWq3md7HdznPF1rqne2yY1xPEj3kFNZDNM/puM2nJ1nakf
NUPKZHTbaMsol2tmMzX5MZgJWVnMwh7w6ot21v6YhWW+NWb3fTj8XLLcCN2K00Mpy2ao+WaOAC30
2xeKGhHUyA4PSGBEjP1SJEtChBCZtBt60fN6WW5cyAs/7Y/u3YNRzW+iCPIOB7xLGmLVX6XqDlhC
37Fpu2pn/vDYIavtR6TtZyOb4bTk4gdRnaJq3FfktPDylsoOWgMF7q+GRPzjr4j6BX0NleQb8kHG
3POuM1I2rNma2E48LMT5aNn9JmUS27qv+xSa5+0oxKVu2vqq9jzGYl0oa9HiLaYLvpQd9a0j02sT
AYmgEJgIAWPuY55EpnAFypCYUToyekp2VLm+rsHkMK76AiPPpxduk1stxDl7ehSDhmYTRapyvsrz
TiEYOLIoM9hFUsM6VAR7TddiUDEThM892AMn3UvwOZatgpQKkdRm8HS7Mqi/gwHIEeWTpmrRp+Hu
lYwYGtr/S28MIFiOXfLCxv0l9ilLaDw6CGp0bPex8DBFSPvcMf7lec82hEdkmJwb8j+KuGdcClpf
HkEQ2cWmZNE+CuGRJoebYRJomeYizMqllStbLv+Se11ntLEAavjqJLcro/4Gnmsqjt0lmco38ltM
EH5jDmKcgEEu70n0WGhj8EhyXwQDvIbgbIkuzrUFqAAD3LFMSntGaPapkXnol6UKCnWbqyBJdkTv
CR11LjVksOS98ksEU6OS38s7BKIeflhFfvGHBZgUmIm/dESdeHBwwm/R5feHgo7yAXLB3dgjhgyu
ZOPynnZ6+Aa9iJ1sTHK/kv1nf2E28ROFgXGfIciBliSPkR5EVikcp2XkGk9xEcWCWEiFaxVKpDQt
SifsYy1dqb4xYhHn2jBSFShD1q2pSxVX5R85ImGTDOcapn4v95DzZfHWbiTpGD6HJxQCnYPSODu8
F3Q4rFHF8ISTZgdYRvfT9F9I6UP8SH6rWV/FNR02D/cB2HKlZTVPnuxKZFWoHAoHYwQctprIpBfs
TiTNO5yQO4IeWHk7Twjj37j+bKZmJ6IbzKT+io9EdK2S+uwTfxLK7liytOuZa9OysMtwvNmbyKGu
mw3evywJ/45sAk7Y1zgnB+VyjE43cLChhvwl/dcTru8uJg6WzhJ15512CoQk3Xhs3A0PvprimxcM
1nOD1O/pR7WR9N04tSVXIQKsF8UTK3zo1cPa4JCj9kJfG6uJQrvWeHspn/9AaYqQVxAkqJRAXlzA
AMgrG9QdURCfFZbidSqJftjPtLvPBsomC5eZpX6Op7quYkikfbpwjc6Pag4XiB6/5oK1Rw+OYSgJ
lfZWgwoRzs/sruQAkxAVeTPoP7nb6qA0jtd8PKXw2icB2WI72oYNnzdmnml1+Ojj7Ntjcnk+yCHc
SkA9j5k0cKsc5WK/Ii5ijJ5jOV3LMbaB4swQLBLEq74AneIIxAWzIOHYgLWcbUBJKKenJptBp4d9
2gXHwjdCJLQhilQ5DFqUuVKJ9GRL6ZTjWr0ScIB8qZVGJoOnAERRXZARWAR1xjcmgi3BOR36JUKE
oj5cn41jAKH6/WMZTQKZ2/RBOH8fUkzISI8iwZvPS2q4xa6ptbzVGywMxhhlMRpJuGeIFf8uri6u
6WJv+xmZKxbJNuI6uv3KPb5fatgBaopst/schC8z1hrSa9relhIvEA02Rf2E6SzwsyC5EdQP40v0
lylVoHyzB6xD4YzcDeNhjSCnhnXo5LnrzJ/kK3Wqph3R49nGKIiPOLZtTxzpBCd2mNfdNzd5HjpG
wcVRbydn7s70bWcl91mQDdw9JyrE0NWcUr29b/K1phMez4U9UU+CIy2dtod4PySFlNnO9RyMVXZ7
V54FVCXrfZh3PpFSDKNdzQ67kBLRrIo+biXjROPb55F3J9VLJ3DF1OBvfpSrTZB2/jzYmZp3bGSG
3fnOytZhtXgMAYZZ++aD+Q6iRVoVU5fe6cOSlWcHfFWnNIJ3QVonRgQBJngPaitgjSVQbCWlnSvV
0OfbO8YtK9eC53y36htLlpD1VqzcIDnSVNJaKn3LxN7KFFQgkOIHYp2GDOBKOxAV3upyDKx4aqlO
V7H2Sl3ygC2EKVoFI5y1JwjZSYLmFyiOpStvwbYRY1+HpP4YwyGJsRgRLHs8CW6phgv4M5l6N+V7
+kl6cenv04kRht+hFsG5DgsWboYytHnfvYj2pr+xiEvBUV7eRdJCxOrrsGVJARIOxD0lrOfqZKqc
h//Dt8LiFxJvP/ZYC1hWP6Z7eotoa7tv1y+T7rQqPmStwMTzDJIeolV1TO0FwO6gAXBJ5p6chD5f
6TQIE8x5sunv9dQQghaDy8s74599tZi9pD6Wq0ulFkyPw5rVQYbI3Xuw99rtQK+1wMagij6fgGdt
JmkfEYR5pvmmYGFK718A+0VPZq10HZJxneviSLzxk3TnmwCZybmqwKhFoCCyi/M79Z+FJMmVxA1z
TY1xY0vFORhxK1aDrEYCx+najjw5nthnV6tojrJrBY91aLIcyKqoZ3qBZmD7Z5m9ThzXqtxkNZ3L
tX/KpSlb6gVc1/C43Me/GdeNfVhZNTMJ18SXIe91UcZEROu+fYFUM+MC+B4kCrLDpGrY6bW/z4A+
oPkQxix1Vu2+VjACFYr0MPnZHELNv+RuGyDOULj7j7Qn7b7QeYKewPiYjCpzTqpgb1HzT1Jr7DD6
3MtblP5fWBmaQK3SysAq6fLUJroqY8//WuVLqOIqlMjbJleXdkzIZKCc02uhTKmjnMDEVM3PD/pE
vt/7HveqefF97btgZtr1gTGmSYsnnYTawBlgpuG3C2HYiRiM9Uj4aKLJPGXUDKsllcc5iFY0/dkY
yU70ccy/r7fOn5+NuiGn5ahNCS8VSBBnLZD+AgM7cJ2dmEEVAmnaMFJEmeWZLQjDuPQ9+YD333X/
5z/GtwE2Y+6LJ13/eH/7dcCQ9E33yB1qaAxNnvNzgBqjbsXiO9lw7s8iiepnE4bzAV9LK6mAeTSu
KVjivb6s4MfbFgBxZPxiZ02N9cVVTJ+eSgsFvzp5uAbuCWy8TnRlEBSFxnZk6dVf8toJ4gMbXD3H
/Wn/c1cDd+9zM5wbnBNQhRjBEwCUrIZpKXwvU4fIWvVtbmXK8BVvGW0DqujuKDxMGBlWJqfNP2pr
Y5PrC6YbdraUMJ9lLKdH93qSBwPamuqL5AnDtZpo0IK6RakEc6QlCSupJKi0d/Ml2KoVJMOeYmTd
80TXruXpm8TWIRlFRRq7ylTAuLXMCh73HhiSfV9713eXzXy5h/UD4INvwmbsdyu4uCNVEsZPE0jD
vel2f2noaaddXmco4BBrLCi9ayc9h7A/Rc2i1Io0sfzeZI746m35XHs3TjEpv/RRvIa0EPtWOHG1
19ZDiLkI3IkSWSWxgd8PrUy/kgJEGheRX0LF/aNq+/3uM2qQYhWoPeZBytMee1FNM1C7EuP1S6mr
PgMa1Xlw0satrknz68kgnnwS6rkc7XWIktJkV+QtHr0iiW7EwsbUFDfxIHdREVmZu87j5gs6Rut0
pPnl1eDI3F3xshw3CBBl3uQ8lHBvoyofWZTZNGKeIKm8yT0CrSv99FItr7oInXV92dPdDlsDyHne
EZ1WCWvqbU3bG4QaaeagfgZg5lVArvnA+p5tYXqP3kDTFF9V8CaIxJo7Ow+4lxSErYobBtXO3NO3
Pzc13iHfzlGJ32iGw6yF6rAgxZTirzaU8ubB0ucvucBH1GrGiqj56hCga8Cz790sLXrqqfxwihVD
aehjSoMt4KapWThJzjNLYp0ylLGiy4U8u3y8femTh33rQwXj6ER/jIaQh6OJL3m5sjb1WT99QOhr
o9H9H3uQV/ra2oBq37w6+Iv/GO2Ip3dv6L1qFUPlKZZ8b7upBivJDu2TMtSgg2Nqm7LrHf+ucQBx
fWFH/2hrnTM0jed+V/Uewg2iuWOTJbpfkl1tgdYIzFbMXrf3/0Z/cQHs9pE2XPaVBsbPFPWTvWne
U4Xbfs0xHexzYvr+5yEJOPmP0V+OqJXxHaCVMkwHFvH2CmRfwjH3Olk1fJhs7lPFkXjVSbjjTyPT
NrQa+jqbG+s0gehl2QqDJveDWGyj7AxE8Qm8c9m5R190Xs/aEsOnpE+qtF8L1Zh68xrvDMlSc8Eq
zlebBaksy1+IFgbF9Dd5mLNP0ETZT0crTVJ66wK/bcPc06driSKKg+0ns8VdJInOsGEmXbcn7u1k
GKp0ydgH7pXShuZcsD5cpEqj6AFOfZAQVKcQrE017aPL2USrZyvULIBJYwK3x9Ax9lo75UwNVXOE
wXCfqLWU7LG3T6w3SFtGpV6bWOLFoLSClGt1eZghsop+xM98U5Kr+ErNedYHinHD5vDQq6mbzhtp
MZtR1CmG3LQt30QzHphlr0dVTDLR4nPurRYMvnEUYpxJOZwsy4NjXnyKgpTmzDCiHkJOPndRqioP
qKqd9CPB6Q4JhDiHQkyWcOcf2H1YDyBSzLA+jK6ulG/zJhgygfjY9CIZp70tfmD6K3ZX618o/jgX
KkBIIv1lNkrJ4K+XN6ZEUfxnjyMnXkVqEIX0FfACf98NxE0pT0yBgnYgUBTy6dYzdeeqh7hR8pNq
TEdYfhZiDwU9hFReFT0XUgeZrj0/bRivPrdLm/vqi4NW129N80O4vxTxfNgxACHwQ+oLjqrOi4PO
pLkUOC+NFAG+ms8g1qrHttkJ4Qfo3fwI3OY3f5LQKT3fuRa7dhmYQ9VZkrgxWRxK+AvpjBHIRqBp
3RqiGIzIZGrvVJsAJcHxjka4OYtS8N3NWc4p3Ay+w/qf116pwcmQTbjn1Nf3AtfCC2262FdA6heV
2OEOdSUp/6saX0uX8ksCo5sa/ce9ntsOOKcaAIIksKKp79+MCL6MmEIj2BwR+7c1hiSa7xkn24CA
9Dt8cS8VCppLZ6+Ygljo59SuB/E9x4+HvErPyBRbIpvDEbkfX8eZ9HBJwwRo1hR1dhtdx3bZIpKu
CPe0ypF/Z/tcfiqkK9ifUm61odM7PgC8KuUy4UWR7ggyM3UUkxaoGT/2MiJpTpyMLIzF02jz2ZU9
UcMD2IG6STjGEk8KRE1qURVOMm5olIqu3+MIYIAeEQWFvOTodnr73v6TeVgqBq0Hi8yy7cRdA0qG
NLfdZ4wTEUupaL2eCiYanYURzLmYQP4bhUB6z9vi7AORl5y7R7prsR3SAK4GoKLy8bcIzonLLItY
f4lDRP3mScmSDGwFWtMEHYzbwhd1RixZB4fu8i10b44Koqw1lYyQoG5f2ON7QSKeVCpiV62cHffo
tmIRyvjcDCaRxOloD3uxdaWi7np35wmAloptIQsPXDApoPGOtmz2MzGyqZf72+4usYB7PqBbGDcM
LKvriBiDcGsLjUadV9wMrIninI86CFC7JBDBLfuZOtyzEmoB5vz0nLpxSGeGHnbidmhrxobh6xFh
L37X1wnul49FylM2kUNbKbbI6pSpcYi5hAbkSodmhgkQwzVp66EeJvO7MPfZ+UswbYX0qzxKFgNd
qLQPujtbOtHpAN4ploIJq9ZcAunsDKYd8r0TpqC/xGoZzmDg5Au0W2q/JGJQ8fo8+zlEVri3xzYV
B/y21+oo8BvVCqXHNjpvDxjTkIjAYvS0D0qwhuELEVyqsAB25GO+E/VhvGUqGr80cClYGiUA471j
ANTVBE2jhhD1hD7QvQkaoik+cvWOFpmTKe47ektYrln09RSNlblGYUjXh16JLCqgq50lcG6vw/zJ
GCmmybcT1ixtREBY/YOl1l8b5Vto0TagH/ft8NP8gL+TpQlTBfHVl0c1A0AKOke+ev9ay1MVbq2N
qpnDCmMqegtGkCEc5LsU+9OhP1cpVJ+woYVJUUR/LVRKxdS5oxJdV7P61XAI2K7p0rc3V9tpVPWx
HSxE9UhZ8qmDNwgJPXguSdqUKoYk2/5JTu0oxfLjnFYRlLJdMn2+/ZWzZFI9Fc78Op6+5Fp2vWTd
hEIJ6MLX0M2rW94BJ1cTkbXmfKS+AjNE0xRMHHL+jP1Aba8vSh7DQc6Hqp3+xgoe3oFlIoQxCXaP
rHpXXz3Eb4tMxSk2KgE9h0x+sf0Md9DOwBVi5txSqEIn9yxevkcUfG3x/UUdi42+fW6CbSZzlrXT
kLmpsfEIeuOwxliZ5AaQ3pUTfZgX1/OuGnqd/CzW/9xY+OJ+Pv9GWZl84gK5FBfeNzPf/WkrXRTi
AqEgYSRq2/pW/1A8t+Ggaob4IHGx8yf4AyVmGEiQLO3fiYd4nSM6bY3FaB3tHgcd3VUKl6dv56PZ
aKP0+HmQvIqJfIgOnHD3k8HmVoMbc4wr6p5GVFCzSqnFLlXVjSW5i0ljSN1uApQqSgPW1KHWwKOU
xvgtMnp1BIMlVhlWCBRD+lBU9AfF2ibTPQB5URkCtK0MJYSDhx4GXC2DvcyRQVbzD/6LbhrzZa2a
IU7gnoL1VS78d+2FtFKc2zawD6TooL4Nv5qzhN2+u1E2Kd5tJjZ4wWyT9YKgtdH6j7NYwnyZU5uj
Es8fIut2CYNq84a+wzYppwyA9qNp2IRPqqiotEMGbLiBTkX5CgOYKdr0tULJubcZGmH/j16hAwup
dOFMHTFfc/d0ZgWdsPSLrOYRHK5tHLzulm/QSVz9gkzZU7dl7OAeMNJKYh9JGE9ABQMdtFjBsxsu
88QYDRbkgLIBaMwCgBjpHmV12iE8x823HzMFwXW3j6Dhf7C27FVeizHfQcAVWkJYp9L6/l7Dj59I
wR7LwyxQKferBJ+WIBGrTgF90XeWCGhkEihebruk1raNPbr2NaoVXAsEeKuta//np/9KzFgPymve
djqDsPJs1eB3NtBVzVwqc9HL0cNRXm7pPihFlGvza+FJgSIK4YS5Ru5Ke8c2r0CvIyVukOQKueY0
LBg5mfQrIdbIvAmxnE/wIDi/X0GuXP1cMtZlKJB5tdyqInK+QSn2fhfQrA8vJ/v7Xl+xcSDWgxXI
Pux+lXFtgbg1iG2Id1hkKeiEQMSB/YwM3IvuOBwEusd0hu1u9n14/X/HE0n/pjYvzzoV9GLTBnZF
d633+YFSCZ7NJErmtW1H7gGX/8j4Fel4YOfH0wzKd95v3gyD/lkqOC8LH37ps5z+68zTt/sd9Vzt
XJp1Y9HEtjIgkZqp6nDI5Gx7qT2ui22oHkDNvMiUGroJ1OS/21l3hHZPC7SX8sJdUk1YwwpQPTv+
2l9Zj2jfDzZgOHhrsBA0wNUNX/52m5OxHnPCJoOJ6i8lDKSwcVb1kd1aRrma5VCUA0BAiCYvvLSG
gjKITn3M26qXoFvVl3PoAyfOUb1quIbi+yUEp4tPRXOex1wb+E6IqXegu6xpfMRCnh8y9TFcT4qp
XZtFsynifMWP1M5BTOwfu5UirYm9tGnGAyOsSLTLbkcQiPnfGawA71vK2KH0iUEbnee/xB/6BIMA
tktnD0qYZkeEv+jRAMauEoO0Jy2J+9yoLLXw+Pm3TIpBPZtBQQ9KjafyifT/bUmx2JPresMGdQSh
0rV0IDMTIqcc2A+Jol9A+XiuihUxGglJ/FQRQT6FWZjffsh/VOf26oAbHJ/2TSIpHhE6RXr97md8
aXj1lVIMCthqIu71HlhLUkZjtBwzhmzl3Smankal2M0JSxNa1djQQ3AcpMAbqm9xgabJvQiAK/5S
+lNyd4lGjUwfWhsc3CLs+QSxsg15XX0ODxFCJ4fg+LnwrScDmYeltzABPL8eWjmGyfu3oJzXVT+W
OrnJ21j+TJJomWDTOWNWdLH5gAob6cpzd/E0YySfRCzWpfpBrNX+/JHzOpaRDA62lCu7ZwZ1ERmA
bZ/uG3GCY0qJyECJU9yGZJ79bw0cS4HBkcFn0kjW3HcJ3Sksx6D2J5hafmCmuP+v/OnIOLHVY7Zw
QzTHoxHWvSlETzXzGTlnSfc+HFnIIm2SjNI6tmEp7Gtrstdyut9rpOQYYgZJYzpIOhAs35E6O8Ro
P553irBKjEfcD64Ng1IuzGVPombBJZwZvtER8iMjKBmj3czUS3S1yjG3rqQy2NEMY1wcbzLXIFgp
6Q4RhepIIbmds3NvH8A+Obapixsc8wX3wvfXpFYROIfBcqfsnpbBqBm4b+KHIc+6CWjRYbUnkHkU
fPZJjpZBp4Uh0oBoyXL/vmJ37XwVTU+enUHC6BKlt8KCAgt95OfBk0tyrZLnG6YPCevdnVNe+DFj
4zBdMV8BIaGElF7z7urDBWas0q9keEU82wkg5AMqt+BkNRGxuqHfHpBMyQ/vnHnLAhbtMxtLIuRj
hFGW/prTeX52bfCBorU8nn7kYvCXe7XTa8s96R9FamxNjYX0f+UjDP4kIOfpazKPntFZ/o325Tuv
DCKpkspmSgx/MRl1WCfLisbn6wPs2Ql/h2JGj2tO4m494bQB6rmzkfrwy7HLv+QglQZ2djUh6W+G
fQ/ZA3JXP7G9x9ROWEKL9fM8kZDLDHC2j77MUQ8OzyHssOEO5L9oU4a7xRKxVXfshQ9TvjGv51Ph
bT4dYO1En+1TogLwSzLcbczVsvxc/5TuJkIGArL9Ucb7WcG7eePZ0pc/oLgeXckgp7vvxf2lCOEj
nM2MILXv0VzLW4swglMY9CfRZfoy/3ZsvSUWmyMdCKatB0dQz71CHFDgdJvrsigAuw+QFX2BCCS/
qKRrc0VVSagCtgGfOlQKBc94n1/3TYiV1We0oZ7gFcM0lSvpk47IjsKUygk/uTt0JIymcBphWQRd
U5Q+lB7+jsQTLr66Uj4dSn45Aj1KMiTZM3S47NcvMYRyuS7FSIpnMV1/7kQm6cRoIiNW222mb6Ct
sahQ5HxzY1Qa2nBo7DrH7Vl21ht+22e4p6Y7Cz1uXTxjcHTg/9FqMPRZSQ914NMHPdmPXW0Gt70z
l247oVmaonr4D0ID5FAvcPdzNCP8kN7eN/nrxJJIpMZLX6jEOFgE9iL6qN8dJh1UFvcE67tBDxzZ
qVkfbrjt/zY7mSSZbMW++wwnqbRIkkZdrVqTS/wKEWe6/8hbZ5AsXgkw5pOgLBFlZBZgtb4av4If
rvyOtpNVevsQbLTyp4NzuNZxL4RN8XsTn6XfkF69SvE4zf2rCsXjbHokKOnw/Lz/Pay1rhR4wGCO
N8VCVzKs3XFXcrrZIl8O484ieTnyGzNy4D8GTPN/3eDMIpXsL7tuqdN//bwDXq52MiBoKJ9M/usW
1TvhLHcOUVvRnsmZ3fYttsNuLSrfDoW5gfbtxkuq8ShCydLuti6vBNUbMpfBvJNPclg5IH/ntHjw
kC1j1xQpohBSpHcIeUBRZOeWx0R9u1e+iYGFPYys0BrE3TnvWJ1mcNVJ5dBGxYAM3PuIWACNjiFe
a4deO87txTQGM+evt2utVOpCdrGV+nEJ3JY7kC38X0ADLloWpfYbBxDX5PyLZq9NkNB88Fx+1Jrn
vptA/3GLEVF4lq76hyl2zXd8U5/UuMokdNEiTU/ODaE6OfzsIqAl0KztKPZBCQBnOgSB8GIkXQsS
U4U2oQc6gy34h83pgMv3UD/5K/QGBpYADRpYPE7JL5ZgI0nJclrmm414heviMquqWelPnb8VvtHO
467XDG6fSWb2d36G3c22CbU6s1wxNjIy9Yz5ySlfXHYdyMz3O0aoeQYPs6vm7GcxRR7jdX6obaPQ
a4UfbJhYkqHnc3h1F7p7EvTMfaPZx+tqcxzoNzQHEqmrLin4YX7dL1M6FngnrTV/e+nVL5xQSbfV
XdzC4ZmXCrG5KgXG8f7x1T5a542cdOn957Ra+MHyKqX7cNYbrzJOYUILugDhdZNBm1PEl741Gun1
EZtme4XMsKAkg3AYLaSO9j6sXk3lKfmb0FiP5nyKB119Bnus8j5oAnzU1i1Lraidt1IrshWo9G/c
0W9Do9gDRE0mp7iDJAKtPHzBmG3vPv6wcbPe58GuTMtHNOGPJaC3+QMx5kjYguDeAa+IJUv4G2Aw
2kkA4dQEXhaxcEITqVnf0EUUdXq3D3guoWwgcdk1zxK0o6FLiwgzk8jBC6TkyhYWvokn4EFCqm72
xKSwbfrXbUOhG0/zJnVbKi6Oc91MR/kQYwRjdEbI5fT5SEV1r7BmU2/ebswwBrmZLmFaQN/yiwpB
CfcNjguO7LdOhjMR2JAmAkpKeRe7lXVr3VklvOnsKzD1WjjixqOTnmHUgBOlewwNRbmzy+PHovZ+
7ksO/FNFUlyfrZE+xIjqbZyoC65K9L8qgfXWnaMkET97eGbydHNhwxm/hFWMDH0R47bKAWpwABCm
nZ7ypEzq6xSr2l/AJeEKWOupRlTbY1AZVqcf+tmF/aFHHPzfO7cSGDq/Rh3WTZG2S3RpS2zUsxe3
SvvUlpD1A0mJ9x2K2yKU1SixqdAUesm2PKHRbkQ2+/on4BKXoXOlcc86H3w0CY2y2rzw4qf2NiFR
6EyKWNnyLUBxdBB6nbNdThK/XzI6fnPloIIIwW1r9UzlBzCpfPdXpuQIxY82I5imNqfaipZGPWpE
/9f7j8Uzqowji+BYzOEMUKK+9XYHpo01s01XyeIWC0Ccq9xnm2wcT1rSNuJP5iGGkp0U7y8gRG0s
Ne5A0rL6s2DV71BXMTWV4IVif0TWuFlCeANyw3P1DFl4sZux9fN7taqotLpW7MmtyN1Ns7Ob6lCU
gDrbJTHwI4qfnaMsmE6IBwI6Aqf2oHT+u2tds417sa4UF0k1KwhEkItLHUFX5/LIq7Nf5m6Oe9WX
x0/E95AD8ygz8XcLpMXHqIa5CPDPA1Mr/N/M52CLl5sIGCIAhgncfd5bjhOXY481ItPbB9xsddq4
aHSKkllPfIo+FJUyFrt9n/7pmD+o7SAE6w7peA0HhMH+XPqrBKnXaCQ9JNsemXG4Spbt2elJcTv1
xpE0JdMh/zKriO4XRzQImFHmhjk92+ofgVRNx3yGGD55yd+A3PvqjZYL1ub0rPApRDrWJTaDVcEz
iKwbEjEXRQNVpVsDdjP9H3CqkAU/0n7LoFXxhJx7QWrwSoSfy1iaL6s6amOWnZKgpWdy/zwVbD+B
MfWvIQZe2C94RtllHL9fRgAieWKWu90ZvzJ0i/NgbxKD8HbzUMCipiU9ZdUWpOTcfFZpqXRtiF15
HK1zUHKnnEscMeGA5IlaKWkpxAaLETzF6kUAFD+Cs05733/O26JZguanpsVHgS6LrzLRLf7SD9ke
wvZNAHpbZUFKCrVDaxbZTtczvx8bC6dQK63nH8YiQrCElTR8wH7TS2qKz3SWcbcCAQo45CxSFc6r
ee/diISd3D9c4D4S5cbneoqmWuSZneTsHR1FaqsF1v6I4rQPWn0aeLV31MUqSflL+qXxp1LWSZVc
NqWYSb/1DFR2khp0B8MrTy7iL9Nw+cM9ufYk2LoedwE5vvlzzkqW4myLgX8C/LCMmmy0hRK5jG2Q
AfGEWjKL3+jrImnQY2V8k3pV3JcLPSf8X29+IQDy5PdQt8ZNd5V3yxNhi9FS/vj+GFWb48omP+pO
ZFAhT8sxPXBGaU07oyT5EBA/G0uHfP+0VbLI/jGJOGj4Vy8WgfOOKYdDV9rTPNga6cH01yIIK8SJ
VeT60jPLP/H+w/qZ369zVIaJDk6mfrC/sH3eaTvSfYuLS0cSB/HVGzNueIPZeCubm/IuaagK+nOR
gdlm1stN2cLtwFs9mCxaz8Xs0sue53LmYI6gnmYdp/WuLJHsIcHxnj/WYBeGdVho5MsfpvSNZV/T
OzYchmWzBn/Rm2oO451gr5MIVSb6ASS5a8gSs93vEh3gMKeCrILekIqo5AARC7pMRBRavt8ovE7E
Mz/6Np37afCjmwD8qR1n/Y/ywYbViYrDc3UoejM2LMxxlItCU78KuEANr4o+7Gf1tp531tNE3O4x
v1TtD/jV93kF7NmIWkl7n1bDrFXcxwxO3drlkElLJtVCNm4oo8Uz+9vCvEp+TA1UkvBOzj073yYi
gh1HToMTd/2/Aswc/8U3/d8OyqSTg80qOhPsO1Gu7hbAefKGZJLHLqFdpqN6dSv3bryi8UOp3Dlw
K3NmE4T4SeI2WUILESLIqRVRpFzEzh+z3cGg7LcuL+sazuVhm3hO53oqkATLjfPIMWfuD1RT8x4+
RUkzzOCpElToySc01q/lBpK9YwdP/xYHFn7SjOuDvkfKrJlXMcicZZ5R1RxtnvHXlxQJSOPRtEYr
8le/1qIf4FBzC6i6PKPkBaN0qUuA3fLgSMGjuG/c0KJuBaOLV4SndJCEY/DAV+WHBBZdOiIuBIXQ
dpB2L6HwnRPT+it9EsweUTpo43EHCO7gmNGuBFLZnlIpSFsWnozKk/5yJnl7rL26QcIbKIGDDJ2P
82LCsPY3hGLH+eQ+e06gZNrBZHEl5DI1WpLbkaPXZS2mcUylBEXsrJJhF8mA+1N29PN0sLvO/DkQ
ngBM/6NfMfafqNhIuHqxXLO5EXxBaOrA8G+zHjxYGbL2uHFbT8VLDRKGx8jAG/rUK22KwGJgCZH6
m7kPKvpEwPhMGjjq1v4gJi1yscUkbYoKJC/9sYN9zscvUB4v02MczaYmOGlnAgfNfiXJOKPBum64
YWMQua1ww4/K+efqMXJzTN++uaOq0kKmVF8RFFkNRHz0sNqEC1rc3J5Q1aJD8qrp+scG4SZ7Rbg+
WhQeyQ7YkLQMnc6zs/b2C9YacZKBZ5AY44ZUlOIpyMFlxLlt+vla7prHNmKRb+DHV1E3QEtFhJ9J
XvurLniCwTW6g7Sknw2uurmXf4rtckc6bnF0nUBa1z8zwEoJS7J+B/snFPub4BpJ0gedey4pvd8z
1PrjuNGGL3YgJ3wnEFtDh+sqO1YlA8kUzxGDILY2ugDvTJ4wJlkAT5VzaNQA8Qhce1jzKXDemo6t
FXuXRaLqxvQ1fu9ESzwJJpFtH6gZe8eUOorW5mXlb2JlVZhWwQDnnYCcHnrEtsApttIMar0He/Ah
X8QdDtMssVWGU4FvIP1YRn3cphmzVT75e53JkBFfmi6YaVA4pgJ1GDtODwTczHp2cuEG4F84gh2e
FTBKj7X5iz1GEWlQNuf16vrAbPXn8AJuKaaBb2IrWZMcOzHmbuZ/vSye45grW6HTngqE5q05BWlR
x1wYMjgsSR256DqzhiPgTRmqf825HBNKBv3C2xHctbeVzb6rupF8dNZ9TIa5C3aBrkXUlXLJyEL0
HmAjEt50uX6d1u/EXnnm0VyVQT/haXljsGMXFFKv5U0SZ44DqbJHW1NU/0uMuKIf9yR40i9IxU9i
Y/jXMHPjKNp1ChwI7kCAuKR4dGhxP6aaiu7yzLCbFb9gRfrIgSqstwKJ1OhaIKGEuWJSwe+hkD2p
r9HdBd++8mFFDGP1XKAILpBpJIcdg+4/a+Pj85TuYjlYVtGQRGVVc3DFbhfv0AXBcIWWYiTkje78
c2dE5ppeqOo1+QLLAv4LXZv9XmpLN7lAGULuwB4C6tfFFZNLRLblCByQSA8e/sr6WhLqAJtFurvX
hMSMhPAEKAZke/SjZz5kLIiqMjTQJF0WPYMydL4Rdr7Fjyp13jSiCmY8U7ZO6HbZKIWoi3iQrfNT
EhLkOiLAcZ/YoO+FG/p+msS0XsDTFNtR1plWnvS4cWlNsKqZaSGcQb7bV8lMKCrSf7arMlJ7u2dt
8MiqDlogz/ZXzGKwTrbpPfEHigA9LLnJJ5InrAXStMYR23hJVaBrYezaLeJgqQKKoaCA3ZAtedNQ
flTwI1khQHlQ7IMAGkxzOqKr3Nx5jmxscB2M648ZfU/eX+OyuEys1tkSUVjHpELiQrXWXgT6i5oz
h0dMqkHehzNbKz1+sv5nnk3g3nG3MDVSJs/cl/wWNV4v8LVkfvGL7qq0SRzrrCe1++2Sv+G6hsEg
QWN8JIL6ruYPQp1FsloDx9T9V2pxZHxBa0rPuBM5ASEJPqKUmr0pSxg6nrKcKwfqOtCtzps8Cihw
8bYvLGvBJfufTo3OIdlq6agsGZLDgeSF0AycOIKkVSlY41i1WIxkfxqHUQDWkFpyHBFReHhL4I+8
tLwjkGY+F1cu8SYYVV0agMKAjomlwh1HJWCPk0KpcKip27p6fpEx9j3rozUqUQnRHinFnhWCbE57
cGrcMuXmHQoxPG4EDL4pjJlVUcus25wJJlgUNNmczxHte+2gz6xELdtEHmd+30eNnt8OwBQRhD8q
JSKRtF9zpEFsjxoEQ44SfbpBaRv9nrSJRuxTromuVLP/177zDW8LIId5mQ+1edtZJf6i67MNOmPc
5DT4dBTdJiTnruwTlb8hI2KOYi6Cly1uGh+KCBt73x1P1ZCrGC46UC0TWApEyeP7fGpO1GMrbHPY
yYVD7q6XBuz9wn6dsvse3vW+m1JhQJynj32BYDGSBJWApKQOB4vq1vbFKu9YgSWJyUcoBIzZPIbB
AhIMn0NF/F/CB8tEv1Z5apyGfaFRGoNDDd2UCNlaw8eveke9eLw9+xzdFZdEzxX4JbIH96/2ds+m
cdrvHNP+lanHET3lriO2d9wbsKjZPn5+ng//u4myi94GfrDEesIqJkc+gTWzhpcHMXYTDZLvHL3m
K8G5oPtTVmWIwBJ0DiUTHCQPi1z8jFQ/+LnTm0MnQXkcyXIsrn29aCkbHMDx4EmOaO0F4Wq7Qej1
qdXgnpl5ISXUDqhYwHTdWMA4M9HWx+xj6m24TPHF0bdjkWBzgyrQYZEsfyfpZlDJh45NLdXGDUU5
+A7SEuPhnqPyJn6o02WiP6iCLR77FBIyIqihyrAjQy3kBCXANwy8b5l8fye9P2H7SO/QTYnFrf+R
xPwhSY5HB2EJhoJQlmfjj9QOMTDQ34Y+vTHQfXijJgidK2k6p4OaDmEsJtHLt9YRlWPnpNq0QCkm
akKluNR+Z279qGL7Ejq+nwucRPNBUAndhEOf/rjpC6YQsegbPpf6cW1020tgR5MndZ7zJNEZqtOT
Fm1OcGJEfG0Mcma/mRv067XAOorflveGi8P3TKjeDHHkq/dmSCqeDUFqJwbsFxxA18vVFo4ks8Q1
zyiM0rKW8maOqbPj/WjJZu8BnFDbyXzyVK06BxDRXoYUrLOFdmG+nv+HWRB6I8ZPNFtZgkGUjQZS
Is96xlgoKvo5nS0YisZjYouI3DA7hRK9eDTo0LlyRaGawFm4AzX8vPrQCyOf4GI9msXeM9OZkIoo
qsoUd5WVEj8/F6KqXQl/TmEF9FWPgLPk8iDrY/xqGi+B5vbqfNXglE1SK/iecM7Jn5oT/u8tWS2+
8kJ7dvKl5k5iGjJ4NxZmuJx1upyewvuabBhCluYprsfp3aKTAn4c35Oxxm5umjMwsdOyXY4D2qXH
7uPZnzkUf4SVaMet2hQ8hgknfdo82OvbFgvAA29D7huMdZ8udfV0XopJ2XPlRNXDASQWSWfyWBZE
ayyhpwYfIC2PqvzjNKsglaKg11iTFo4yhgFC63zobwQ1DfDVMPDtioxYIk+S2Khn42gPhzLV9rGY
NcTZfYhjTzcrhLt1z2rPZ0E2yx90ZCD/nBwylfSsZbDhBrycxV0nUfB1JzTJGJ7Q6kAoUGYdhPhm
SSJJuTNoaQNsvV+drRhxh1U5Xt3u0D3dU1hdwXjCAEmWA2J1UANf2RRUayFuMAmMxSUDVtdTPrzV
lAcxXzYAb0X6drAfu1UI2qNS8Tqc7NTspKV2cW4JOyByOKzkXBLn6/P2+wJU7RwS4krrykIWdjRM
ZRz9N8pRGaOxa+0LhCS+NtQMsPjTzWxn3tjlzw2BsITLP53BBAvOZ63jp9GmqFxnK1GzY1yb+ICz
gdTZbkKr0udXPjvT0aS11pugBWY/gtjJMtY0Y7vn5uxO0jf1PuNwBr13CQndfR2//PFpPvUJAg65
GixB+mzkn4s3w8KDbkFKORzLSfMcBnddFRDSixmlLvaxXlejsvc25Zyv1P9q0DJVIwnuNxK8Chtd
jClmscEYjpGReT1sXHjyIg4uvpQ6WjLUBr4HkSeAHVQYB48PCNI1T8RA0ir8JpOKCq3cNQb0xn1w
AdMUNfQ33Q1NEwMykWv8sxBvH3nlEQ2bZLK039K1QSf8Ug1PlIEvMY5cSypA6iLn437NLJt/TxiS
QWgNKqnQFwlR4RUape9VI/OMeAQDuSz8U+mEnnF4gtroGe1gY6nqGlI+eV43kmdj54ovVWoHtOO6
Q2KDUPCJhaYZg8E0c4RfXPJj7pmEGvvRCcErErDa48wZwjPl+xcWyIGcHzI4wkWcyVyctEu4cV0m
P3+RjODeJqA4iQTjJ0AdnxcTMsjZQgYPOnelXesZxbvG2WHE0kCf9tl6PrJCKb8DU3oQntCraHi7
s+BwaPR4PAtk4yVLOhtdJXtfl2z0lYKMFNxpfX2iDRYzGt4y5lU00RvPpK8bR5mds3vly25oNlwD
rz18TnqlUUzDlQ+8gfQEI4i4dhhjm9KoYU9DLdFnef2KXCUroxSznfGbW+U3CTcpaqVvh9Kxi8gY
ZZ+wHrCVSmMHfqZS4VLFG5WrQ8n65suKh8IpVD5N8QUosYK206HTvuI8lkiUsUmFG8GuwHQgzsqJ
cLt/WrTFiu6p/vsZ97mwb9jzADcxmmZ2mwH3LFZWx8Lv/2gljtG1byfSUJbSSviyAuRwbr9hPRw/
UFqI04zwhc8mJ8NLavVmt8Qu+jva9yp3/mjI9RqY9WVNYlCLsdRRVCTrBvDe3kS3nzua0Yoglvzb
U1I0h0sezX1+frcj9zMs33Zq1SnU2LCOzL/RpuVbAnITfn0LdwZTIp1RknolqhxMGbMBYyuhF1jH
ht1ru05ax2euOuqGLgkzf1MUGqO+3m3OJOoaCewBYB3PZLDmmzCFfL509F6QVi1yi4aB2sTcJ0rM
imw5W+lu9d2g1vcNrYeDKIT9EolZ5uYdIaqEf3bfC0zBs5ApyvF1+VJpytrutC8otDsYBQbX/ZfT
wR+4n4i1EqW3WQYK/7ceeHQNg6NFJOGzf3SBDQ85yXrw/mRkIubm7UGgdL/SMmMdvapNKmIzxwED
lMq4YkRc2HRICoGcmQ3xwKSz9Y9mNqm6juSeAAICjVCyKvZI63l8RJnMHHKgxxXrEaGtYQqFFQT+
am04ZVOYLrneWCw+hzjK3U0iyvoTgsyi1Y4TTYrgtNHsZ3oWGLTQFdGlsnSSevfD3aBjcguWInCg
lpMNt0EeIx0Ce8zseVjnqTkb8asKOWvr5D6MEIlG4GyPJcWlMQoV6xXGtY3fktQhAfE6imd7pAev
gIiGbv7H2uIWJpTb6SsR9AMep4lFJbL92FGEwtFG9Su8rdYFLi0D14DzSXZxkJdDcV3Xljv2d6dC
HIRiuGUT7q61cuI9JtB9x3/7KnGEn5/br0Bql54JuAnUPSGv9O0nD20+8n5Bo1aDy1zK+WuZRLyg
z/owaSVP1dFHboAw6EKXpKu16MtPDLsGV2JTGJtJCeS1tkCfMk/sL0aXubP5A7kBqjsvuflkAbgC
G8cPss6het9Eh/KDa0IWdc225p25IIrJN1VZBjOp6VWUi8Ei0MNyXjvEXINOYTiJN0HRP9qTK6p0
K0SHx16anlifdt6K+GxEhYOcBi8JqmqAw1sMu2JjMVJktRG4ZDJYMHcXr/XdRz1NtgrlLFCPCfd0
EEfelKk1pCmuCoR3Ra1GhaEXXaL6AoQtz2bIjqydG7aMeJ3lqYEJlCNp6xH9jjT51AfpkWtbp56k
Wtu6JIe37ShL5s9Tv6mngWnBKRD/uTLox+ymJXA17/GWW1MOK8nPODFm6z8gMOowosd1O4d3CguD
o8NSofjlRciWbdAMTRCXsZqCr7vArSLs/9ro7xsPyYJHJt3yYUfx/B6emoFxJTvQhT+9wNhIX5t2
l4Eir4A/R3uMh5OkMKDp/1xZofGNBngwJuK25o9P/C8T1h9J2L9HXJfG3Nt0Omi2eIYHbD+e5Mkk
VI+MD3TlxUqCHdFYVP4HS1I9edTz0GAxGV9QIwYwf1xrDwM1cwJCFjdBCMXo9gV1kdEtbkCnbjKt
5ZyTRozRFsp3ZOuwwjmGUXq98zGcdS+tXm+N3vxspulobrIItV/9ssEWglGwbHJvkS9LTCxAFWr8
qTWmIJ7VtxHDkbyOGa6SicMk812XTzYWI36POyua4UG21en1Z0MOxPwRk+tbZAiWjdIRCMrtwkcr
FhsXAJFETIYIie9ZR7Q1cyLkBzL981g33KIo1Vv7ihXo3mC00HvKAHwSo7Ld4TnJXkR1LBi5/ZDW
iNIEz6bdVZlXFJKEQndFOa7wBSeLtvcko9Annzg+2t24Bv7/xATN2A1M7iFbvHSShp5STRhzurli
SDFeg2B3y5tFr3ugGzO5NMxsOP5GYwPXsczCDY/pY/3USIg/tAwmTvbm+YTtGZkf8nQQ4iUnu6Fg
hnuysis3CkmTdb7AUQpErVN733ep8FIaBv8vmkbX/zwr4FcYSP0kz4dzqD2hYRHoAaYr/IkZ8vkI
xg+CnkXAMGrTxDKQYhkVAtLCwgrhqSQ8Pb+VJ/R/IGDMxu+Og/C7MtCyTxx1vHU1voNPX1wqUMic
VxDXFsLi63dmSQ0V2diT5T8rrbdIsUWDZbFifIW36yu8sP4/6++qGLWitnIWSKX2LaDE/SPurzCb
fCee6IsbHfJNrDf1onvUw1Fxj8xxT0a12qDnuCOjBWHkTfEJWwHP607sndUvhuJvP674z3TtdAZe
eDeVmsWf/JY7hL39KOmshJcVIwIuVD9QHvuzpmVL9cDnU5l74+8M87Jx00arj1nhLbiAD0x5n/qI
34KCGNZiNUWQXJ8ar7kPbeHbMheddiO602fJBSfHVmNfwqVCwEnia2cULokwO38Ia9qc2VfZhlT/
bwY+RXpXABd6pIbNvodXVjalSGYiU1KYMnsAFIbkLT+M2Vkq8m0bZuO0BEEKRv5vvLs9GmRtALZU
nykqwoKhWd0a3x5l0c7iDUTsA7gpva39IcYDV0cUs+45JhaQK6fI28UEFo+pxBzw5WGLONvKMuBf
wJrLATgfAVgMWdxp1vcnFQBrZTZ+NSJLcP6axeJtaiiNsDZx43YPq2pqJNZGsccb96eCUQKZhW6k
dVYg/FiUHMOboWOBPl2QL4viwEg+Wj578E6JHGvexIRxlqNOjIJt477zfnhS23hFEr3kJIERUItv
HP3WjaE8020/2T8Lqo1zzfm/vKLqb5PtYq3XKmOQ+ell6Y1vrkCbem9QoE0gcJBYDCPhdNEdoBUF
Kh4krmThGeZDdlXols2qocAXQCj/26kHK2HK2L6DKpfAqBWZSdH2iIRDuYjOUJETbfeTyuBZXeBn
X3onnKq+Tq/gQLmUuX4rcgP8vY0bGFUbw5HpAjMu95M49zMG0LdsSNhhF7gnSg2BKJzvZWg98hTR
CPpZ/1F2zEyiLfmTzAKwwju0CERcaXM9ElYNKxWWTLlq0jriMLqpicrVwWl1Z4QwIFWT0PjGPnIQ
CXEu+XM/siOJl7y5x3i0AwY5MMPTxk2K8UEA36UCtUyRjDc+3kW6BPGENzLqzlseUUxOB7moO86r
XvEJrSceFRnNciXRyS6CweO4ljBUlJKpQPTic2bkNl4QVnKFH/Ik2KJ+ptpvyyXWnck0lJS+CADV
ClkugxZUmUOo7GuH5+x4UsPmcKQTpGpaDeC0pw72DQuR478yIX2RPDt6BuL78o9bzN78AAVVnW7G
4uHiRCy0SxWS0NNaVsRVVUEFkP8j5QIDaUldYJuiu51NdzvpBxjXTyHLEP6LLFlKzE5PUlS5CAUV
48VyJjbkUcX2m+3iQhpURjdTJ1m3X2MSX+MvHZL+KLZ4LAFr5Tq4YHOiKtacJJx2Hw2ENRsCV1jR
1/PtHyInCPqzldWd6dyXz30ZezmMUUxtOXErFUeheyIbDmxs5yI7+jOX1njcxA9y05gS/tOX6bfJ
7naFLuK4a+/iTdj6Qnt19aLziLy6DBaqu2u6ptHMey9Z+k0AtP/ro1PwVma6xTDcnhL6uFs71EGV
an2+1aRUO0Z2kyOuJ3X7Y+ImyBP566QHw/wCSfGNmq8DjTvfjziXB/McIQa7IsgWQMMoBZcg0OgF
xlnwmpSeXRA/OswaT7FED3t+Ja+2SyHJMWeWpkG0FUzCnyCrR7JSZ30rJZrIBemXKVXdwlWVuM9J
3RaJLB991U5tRbcf4DSPk7dK+PjpbXNhyM3oXzbMz6VF75j6p1afJ3bFh8RchnSlY86wc+rDSJh2
JGXWjGtr/TuKP7B3bmP4439DKKg9uWxiUkrpAu6sCojuS4B+RPMfgFjvM/WRDoF1raKKWGFC5Zeq
ohgBqcaAmx3XcgmoT0q+/X55S/SHZcVUIYt0vEd7sUfXnJHkqpNGyNvMOzmI4X44+x2MV0ZdgB9P
6yY7wG3+a/wFcCJTwdVhSBWRMm4az/JVjjf3kTicWSdQ3Dk5fJpNBCHtF5EfBULJVd5/ZMBTB1VA
T58jOfE8BLPzynaWs+gqZ2c8SkIOHLS69WQSfwg7/7VxcvhHpqcl6gQiGwWMOGJv7i7IdLPuPcYK
TKonqYGGQuTedQFyzInOrmWAeAC4wISipIGsqgetfoI+nF51LyPwlrv0eIiq8wtdRXO0qog2pgQP
rw5SEWRVsMsKdC/jMZDY67anrrZjEfmd7pEjUafd8QX8kb9197BqQBwAE/v5X2F/3AFuu9UET/uM
NYMqDYSD8lisOfEij49sR1T8T6RAdawWF1qAz3sTtY3UCeZgOKl6DJuGGPlN7dWrK+GPNhTmLyM9
Vo67cZSSlUCMsrNZks01d9EXrQP+dKssg+OwexxwNz+P0FLXHHdxghJeYeKSNuKDVEk8WHaznG4q
xV70/vxtm03l6b4kiCiAKi1xXAJb3iA3aDjBDldl/PQB+Zw+F/uQUgLjwSvs1faFBbHEWDq9e+tc
Cc/py6O4klemVYt4FMJP6HNiAPUFJ1FnBLaG6JOq3vdOCLIeN1N9ubUU2MH0eZ7H993iYDcxic7E
ZXGIL2yVC7yIASaxg8ZozecQPEO5ih4h2HEeV8GrHUJq/2i8u4lEHBvDVSpTlITiWBDkp/oUBTnV
gPpyZqGSo5rKoqihgJUSKDXNxLm+kBXEeGWOe8uAT4wTKmBBCUuPyUQJOMFUcK7dz5fy97hjrILT
WCTQQVeMpkT6DlKGD0FaVVV5mLf0ejXnjtlTvQHAotwVogaUom4J7gEZATVJs+UtSdwE+G1IZQNO
PsAC8zmu/T9rE6XAMIVheTdyVKIu0b+p5z/MTNbT5F2wV7ai+mMXUHx5JkpF9aIvBCTv9aPGPLgq
cYcTMWb9MgSYvbGeIZsZNTTSQ2TVAvmFHJFPZFdqdy9iLdTvE7V8qcfft88izqt8D5JjSikGzNxW
x84ASqoBy8ig3OWi0fgSgJTyboF0ymacqAJJ9jftLfQ0XzkitCvOXI9xQy/z5hUsYIO7ziExdLW4
XU8Pf6gC02qiP5u7DlH3Nr1M9fElFGFgdiFaB76hLRfd8eMGxp4AmZo7hCdGIRuVNEMxbtUh5/6P
Cfo/an/p7YVoLp/0mwcTWqYCQMEa/TKhylD6+PBgxZxImGD4lbMxbINRn5bD8Ke9TTtK+T0NRDEY
HMxoiFDrsJO99ZjHYHW1/oD3VN1kCEMzNwOl8iPRtDm2R+/3SwsSn5dwYTQyNODqAGiEPicSMZhl
hV/4pfiedukA+MLgoh5kiBa3mUXjmLmrOX5Aroo1ODDXVXZzunbKJWHczlpMm732/lsyGEUl8QwQ
gQCns51ZSshv1653IBB33PH/rPSOsnjCUc/m5zmWq+Q+WMlTJiAjmD1N5xCYYj9i9JkSmG9QJEcI
h8jG4wkcUsEDDWnIfht/vvzLIgujX3uDSkQnb8ENM4X+NaEhv5olxqkVYukXtvJqDTdui3piBJDh
KdByfCJMT99pEcWPl/4UYgjnk70dtS5WEX4D1+4vTI83JWYxX8CxNBzCdBYnSe+u+OFeB2MA3ncd
TTuNluLxwfFvyzKYE8HM5gxK76w+R/36nxIcDyLpX7MM9jUvxFLyimtwRdd3GOg7HADTPUBUl4+b
2aNqwp5e3ZOfypzgayWfdmKgkdVsJwg0udlQ4wSpup0gkIDnUkJM4Bg0PEuKzUwCkwzdMXesbcRW
+HCCFaFJ8LxsOVFZFBaswzsvZz9/KQXBPKvv9rHtPc5tdvj5lSTNpry9az3AfrVYPrcCOJC+HxFe
gXlKworVQGB0ZqgfEPE8kd5Xalwd7hFjZ0k5r8Uny3KsbOR3wL4IkVPRrif7tSQgcAOZFQOBHyQ6
7sWamZAVvYmJ/dbNl1aF4nFdpiQANhke+sy6VES9NwayeJtov6+Dmr/jvAMnoXmu0IvTMk6GMW2G
t4Dks3IReBINfbewIUCLttKXJGsht5/Dlkw3EDwYaYkXU9pmIo2gLNlLBQWXPWx+ha38jn006ihR
n3C/83Y54S8ti2GRU+5jZ6cz7FDHpN/a0oV8vRC0WEIAqsvn72cquMPjvpLR5p33EMBW5mfxJ8x1
w691FXJR85cplFWNTbE2QQw7T/alvrvNEc3sVIbgqMcT5aj+NmymBrm90biuXhF77d2Z5cYlmv6a
RGNKq4y9MBOvTVjxP19P34H8+vbWYyixwP3Up/JS9aVPto/x4CQLKOUUtNt96gTxBim1aJ4pgtc9
8uWSw6LNUP9kpa2E8biS1hOhfopP0MqZjf7BIJh1mO1ukRKH7p/OqS4TQH8wKSDVLxHqfq+SkPLY
dxkAW3NHEh5F+Xv91epvIb4c14SSXgv/3arhlYGX5Pxl3kjLdF5yGGOngJeeNNY9G/RSUMygH9KF
na9/yKJb7+9NIJZ388Adum2aTy4ITEB3fOEbZf/6wwbpRv4m0GmwAiddVJ9+UscXVaTu1/GFjS2P
92J4CPmrXGYf7rbNT4OGOM6AMwRKDnO6/BC2UvIdKhU16be0M8qFjdIpi1EhJ03mrgXMvigR8wI2
en148VdwZ7apB3ryituDKAxWAda1k7QsOO/9DG6kPdRi/+xdBxN9VfdFkZj2gPf4Py2ZWbHR+RhR
VibUh82g9gUZQNE+3bJ00/Cey6/2JG0WgU2jxSaBVEHcIVoaeBviw1kIMXk6MATTd9DrdHIQxnL0
Ep5VkCxRDhCrpRG8p3BNEVzWUD4REk21+l+CcJXhhSX1HEGovzEvdOVPbq2Oq5XYjveKd8HLBn/t
U/mMHxOEHJQlRdzWKo4hjl5qpXQGl1loo1DzCzkNx3a1ak9jJzehu92aA8Ujf7AOrFmtwQqHNh9I
+ThxSM/E+9KSLiSyRvKbuGRCJELmwuEPCQbtvPDXQbPIShptq+7rZoJFOcHLZwrS08J0Rs2lIDVq
PiT0SROpKeRPGNphOzCLHtWh5HMPrfcai+1JIiKm31I/NU4RS2107UgjdRzb/5nig6JJzBCnTedW
YahMDExvuITmUtZVidGiPj+ylL5CbZYrPGPoSoREg81WQYZa22bogGQxiR8IQbJrxSTIbAT1f73h
ogNbiSDSysXHLPpErovKibeme5MJ9LGTUfOWgdFLMCd+PJtcEon6HXRIZDJe6q07PTwuRMcdS0wd
oKnGxnq4sIqEXq/7zg13/BtwwX3+LxhKFmvLwvXfc0iye6iJR/laA0KKtM/Zat/jc6wNJKCPQ784
mRU9J5Hnf6dOoFaTcpzc6ns91FCF6JVPjC+tPmDDBXwZOXZ8+FleufpuyIUWUc9PvGNLHnksaYeK
zNjCQbcXZLuzR1vmcAcVzBUaPT2FIGeCGJYZuzg6C5hBpnVbQLd+9qN+iOdvBMW5ewa5YKfG5F7+
DK6Cvkfy6M3E11ke5SKc03q/KYqaE+nGscVRnDjl69YGfFNJP83tIALKK4iS5FZhNF8y58oX9/hd
h/GUknQxrS+3Q35PJ6u0nX33ylDMHymArCJ7DDyVx2qtd6xduuNWhM9AlotJLJAE/j8jb8sc+NMK
dvPsrZLSQQw6kXhVXijUiBZw5JoZVT7suse1ictYYW8WQWvgbOe8UrAzXFCNoZO5QNPz7MHBeS8W
W+K/ldeDP1i/wBFLpkWOKkGUixceS/zsbDK8PO7+1/thGuqmljGUr1VTGaf4+/T7FK0pWUySduzk
eceD/WmtjD0+5gkqnAP8mCfhr8waQZatSAgzv49X8GV9YA+gvYoYuVccXjR0dGYz50+Qb9TsPobd
HzwEYV08hkKjHNisHgBPcnaofHIWbuTy8mOZW+TwAHgD+0c0TzbHhf70xWOcuGB70QatKElgmpkk
nPU9mmtKrCNeTTIrl7b8yEd+5+HVzOY3txouZTIvRDo/X6aWoZD0+7o4INHku9n8cVGLRbLYt5ec
paUXMgdPgU9RUDoPqJJvcE+ILb8k+M28tYx47XeaVZXZeykNgZGiV1hLG7QPePsaWcH2of7Mik8g
hdG2+oTFoj1wd9jD4YJrb4swjFBfumtcwd8b2TIEnRES8W3HSGG/n0ldtx+vIayRxIt0rYDATxvZ
ZJthyJFfgadUIjkYCoX/V7ByiExTgJxmNreBwzgzwCVpQENss6rTSzsK2c4YwpyZCjEZ4oLB3YJM
b5VsPr25MMbhbhE20o8Em0m1vmnYa/1wy1wHeWx0M1HvmUS7pZEVyMHdL7SYYHPH0bumjo16Tngu
nHZN1/q1QiKxNBXKbIfFNF4zSGUQZWD6dXdvAVGGiNwoPHmUebqa4WhMkW1Wt1LVZgK45+qUX7mO
PfDHLKK11e5D9JKV7UdtSDMQR7I/lZNRc4xC73XwfRmuYe4FeEn2BZOuXDDGM5UMzVoYcRepALKd
Gc/pxWGVMAxnHnNPpKxR4UECoD5p8OWd13wYt9fxNVjcukiTWNSQETz3sSyCmulC7kI6tQXq9dwi
1iNjUtuPr68+dt97/A77SDbVJ29bs7ZTjBru2F3R1dWMN12aGE8EZKDMz9SPqtjK97zHpgrZ4giO
JB9yhJ/x9zeaWio467oeqD57XqWrGAHDgafUfhanE1RtAD2EzS6nuVvO1xm0LhyG25IuYwwOxN3K
2lObMR12SQrR28B7Ih8GKNdv3E0egSPm/6vyEQwE9mk1XOSwf+KQebGH6lRs+TALpZXbFl8kcGKC
eg/adRZoc59V2QvLEl+oSTW1BsCR0MZydWhJr7vYsfmlZVrByUDRUxRMy3ItOiPxvgTtAPO83K6V
yxCqFtU6XzWg81NPh+YjXf6qDk/BmaKwPjJ5KD6i5r7Vax+3778rQ83CUcUiHMhOxV1fveC0zmbh
w6XEdx4Yewk6M5y4WsiWgYP6SFF9saoeEdPPjD4TrrH98daS1qLI3GSDFRgA5gSKt9v0S+u1kZp3
2kZCmFGT5kmcI9oWRDD5l6nN+cDa46FMVYo/nyYxgAAk089Z7L7HNjIqxo05fAVPKQvub9XFA+7U
HWSGD37s8tjaMmZvzW8vF6KklqrfSTx8J+YdEiA5HZjvQ4rElxbz0FqjJrFNpr5BSiUArviJ5q+X
i5H3BNlT63eF1RkBfTv4gpltfrt6udeaJjrJeZoIkQ7i2koKMca50wmEgKtWMGLItw/7rTx5gwsV
M7mcE7sxbkZhK+5ca0ISGaFEzxlmVBDD4uMDqvVykORL4CftS1O6+mMFDAaCuLHdj84RU8Kb3bYI
uQTDUOTTbEQqELus2jO5MR5rxBhTg3VmVseo99gURhc1M6KhKBSPsajZkLp3oEUc3JHnhfNkUVaK
GfRFTAXsgmVR3Rgvct96B7M4wo29E2OdwPDe0F5HERXKOepbqwaKAuxdV/Cbt1IqdZ1ySlMDkbkE
sNNMdM6lzU44xFaHkIaSRCGBn5BG8a7eMYVW4fAN/E5OqOPuA09ZOc6VSy4NGpHJgH2pPjjDM51H
PMyzwTcwmTaNLM7oucn9W2K5see34N2KXru+d6XJW0azixz4XE+ewPkul0AeCKx5m4tMgsSbRR/4
2tVhOVugyFP0125fFI4Iht93U3zzdf9qzio7JqulPfnzcv22ivBi+NiWJ9CVqSeHOE5b3YYP0CC+
pDijcTTTRRVZ1LZqrV+MY2VAgs4t8fCEK6Sh+8AZNmd2Jg+EOhvPTY7a8TVMCZDIGW4HA14fosYH
eEYtTcXLG0CIo7Xdkr7zDLUBUBpiOpmp2HV0Aeffx9zvSx140rtXT6uWiXXLDcIHLHrve4qXkAbB
MWQ2zTFgGo7AdQVkw/mQcLVfse7UXCBWAHPrit/4dN7V95/qD7HpE9LkDWTBQ7RQWHO5HpiybNP+
nhEfljZi3G2qZC9sKSaVof24f74UZQq1ZBMlmriNFPAyEHTPp01TOL89p9wmEnWGZeEJIvy4ZgND
PP4rTeQpv7K5au+fqGpqCXehSb0OocpxGmQp1ZBdXjSXIjahkWDjU/IL1oR6omlOhz1N/WFlKdUN
8MTQt+VPjoojj5A0Fh+z/pIrMYE4PV9Jugr5g6slMmLAZgtYHYxpQ8aa7IsyLk1+Tr3l18reZQ/u
c0QTAS3r3iIQuvRqjdpYy0J10VrT4gWm9mhQ8uPk6P2CrtK0uKVY51DMeozV7y2WBbcukAIf46fd
FklwZs9OSZ8m7QDmAOAy4Y41iWUipxSOmL9drluH5lV2mfdaUeGBn8ZAjzeMsr65bMfWp0WeyeFi
0Zg8p76wbnpgjfny16TduHq7o4sA88T3ssIMvl+XP256KDkUvfsBx943VO3XDoVvuGGYe8OLU1zS
lpDsTq0ErGVuYYGF0jse7H9ffBYzjgjtn3y1zLWEOEXMjrFCncskGaBIXS+vSQYtHbTtjFmbg3ch
MrJIbyjQYDIz7i7VZHRhBa9WafiV2N504ig5v6lB2Xa8B1O3uH5ZT/42zzImYbDsgQgLR3CGqZdY
S2WF5M6LDnCC16R+M7B4LKtJ3nopxAZa0ShnPfLAPDT3rtk0NDQ9Xwq/zAhVLPSN03ab6sN0djh5
xgHqZrYZa8960fjsEXzIaQ2eColq2utMoUf8m+lkW3gu5wyUQs7sX69ELT9Y2rIcNZytRvSjABbs
i0/gTH1/D53zGJMp8pnBFkrMO59RBlQhy3DPSUbH4dUU8JVdyQbD/kv7Z+lNct5lM+tT8oupoUp8
uY8+tBUdmC8w19BIsKqnahZETqryFuKlynA1X4xQvyC3Zl4BRgqpNJ5mq1sUozolqDGfsqO26AZm
0KFHI/7Yzrwz9SpK6KQHhkFe+25eXwRQybWeCWGPE+KDyks2QOIkZE2AKFzXEjTGBHcsNMeLeBFr
fz1Vl8QIX0Y7jq+3r4rK2WYOqzj94l5D+bXUaanlCdmJyIgzVXeEFtPgH88y1AYPTWkzAXXDF4Y5
Id5xwabcSM/a+pv8Ox9OwZfQpGosRxfdsuaTLMm6KnBT9EY3yj57unx4JjurwpcubCZLu5JF1/G4
v+geCQkGS5vk/oZ5GPwgh/IiwAOgGh8WHzQNRZskLnbMSDwQgxE9d9gvQy7ljh9kQ4MOrWlwGMon
cAzfmm4iggCGFKDTqrYl6IrHIK3z9nmzHaui2ABNZFrYFKwx1chwZzJQuNEOQNrJB2ug5a8VwFGA
UaiRo4B5Sn2BgMrhBYzdZuboBDSJU+0lt6p+59xRvKMllmFAE3TKzlMPeJ6qjwzaSxGJXtr8Fi/3
WQdTx+aTNzf07DDAd2D8cjYCowM4ulYi3w9nK7WTMOC9UAQWxV2BoXkZ44l/nSv8lWZEDRCJkkgL
bflRI0dK3bO2AruO5olTXHLFjbQfmftRqOydVyAPz5krDxlpu8cK1l9GHQcl1w7F0RQvCoFZy5FS
E5hFRgp8dg5RPyJUZt5PGOXM8Mru6fmcBdKhRFQ1WdhdPWbU/x+XPTDVUrpzvJOdVl4mT1SLkk81
8O+QHu7zfzW/6QSo/W05p1aFI5XEvhSEzsf9MbCriIIOvdFg+4xayKwd+CIB4ViRlSN3Tviolefh
kG6u+6pS7hRffYanq87gWM1U6rl/k8apzQRW7ybdElyGNTQbTYIYhaUybw4dpjJoshnACWadDSGY
UO3eWYOLPP2UJvHEK/abQATUEYnKtZZyGPUPPnO2ZOCzAVJ2KJx8s7uPm+UmRsOS2c+gIma+hFpU
DHQCJGvBDqbzizqi/4v464R4ZyFaW+1PRkvSwubUm+M77MhXA5Ne72EDzA5sKKRJrd0voFes3q7v
cC7lqt3O2RHUvlBpN9CucmW4utEEztrfeq7MNpJEhiwpW1MyPZC60iAlQ/oKmZfZDAz9/2hN8FcE
Czlc94n7iX8YGsuQuWJuI1Q6WQeZIutPWxM83L7RxITV1L/w9RZtWV+xGmofouP8fdImzlAVHPBe
aRNefZRBXY+clKYsgFXQjW2a/wV/uaXJB3W7fJJU1mTJUKNjZKuy5xo9DJ5DnVWE9D6nb4/pYy4e
GY6Edyk2jJlCrgel28DTlE6fLI7PgK/Us3tc9tw5sAKDguO05XL/MTVNWAxexLA4ARgHWz/pVU+Z
h8XSjkEVfIvUOGz8Ywf3uO92prFvpiRnnsZyEcDe4sl2gjiP1ObtGQW4hlx4BBAnT0gr792VVIR+
3mRLUBuiuj/BQvvy8qNTxABLsOQ0WFjHVUMgMpTY4rhlNkCUqrRrXemN8mzckE+dVPTjV9yvb0S2
3PKIBh4ipnzwB2gJ7f6qKevIx88Bwqsmvrlzu+umBdRq3sgErMfKT83ZDdZvYV7616RNcIei8zwW
SZZ5xvFGpahL9pMPjyOJ7eqKo1iijA0bYFcz2F9fIJdSTt3UwsxELBE4TnVMMYiDApvgM7mh8GRY
plAyj7GQlwZEhchZ9KBgAxstlATAh+ax9iVf/jEi9VuyngNx+f8BGpdoYvn2ADt2F9rdvnKux8ub
UglHhzXwxIbSO+5bx1tz+ohmLbhDi/KIn6lBti4UI5uZHwhjOZUdAgMOZEHtq1Kvp02J3URqBowg
Y5GhQ9iDsQCGUjnJK+xaVT/WQ4vazbWZFz+eAwk7iaa49BBc+h15+SxmmUl4OLl/Uhiz4NWYkBpc
GjNpiFd/27DzXldv52C6Nhqv9mlvL0ykwn/KpAWc0zLl5/4faWmCR0VyW6qMbhayenMt6X1j0ChL
DaUwcwTwy9V+7ZHP8YqTiIDLCuuQZDQMAxUvh+VZARDMddG3YnfTz2k2wwfDKmAU81nPrN+SLEVC
C+LKARAs3yom+3a824/IYON7xO3tabZbhe1ag3DlC1UM8j5Ome3x1u98svVorgXQFyfsd3L5CefN
VLLKDQbTW1JMlSRjulB9C5/MrOyNIs8hc+fK3sxFiXF0SuDb3LvNF7O+mruLR6KaEr6by0raL7SV
CouMgL0faBTBoS38pldB/TTrjiAYsyA8z5tzxF/UmBsOx22vTERUcuM8lPFrIiNHUgti1EfQ1Y0/
iJ+3KkkHpuE3SeJEwgBVzJ8+OGCglgthPX5qpomQwtvPLfGVQRul4XUW6CZ4R0l6P2dfO3f056ra
e1J4QMo4LhF3zcIdPK8feHZ0n/5N61cnwIOz0I30/uExwApCPD3gXRhXsl38eWH6zBL+edOOy6kw
g4ghOL4nwwnAF5ANGI5llBluGYe0+IwTt0nbcCk2Em89b212j+4ecoQWpHOobXpRpHVycgJXk0QP
Ko9mHKvG+kxL/B+VDTdgJlqd/NOgNXZSJQb+M9+emXhnjXoBLLqLuQdpLFW6lFXHtQUY45755R1o
8ayLvBit/7e5+cSZ150W9fBlS8h33Ysb7HCtL7XFyV5kWlDOE6P4HRtCKUdiEK+ObWbI3HPzOUk4
POrgc/7dxFIGpy8hAjG8XkSEg+dC9APh/CknsXhkcIE/o98iwL8wFmKZdAV4ZBOQml7G/jIVktS1
nwTmBOUA3gh4n07xKUn09+5WLKRzfE3oVdkVWf26/k7d8JRkTVZQy/Gbni5WTmzT1en5Tzb6kLkQ
eN3sFlGS+tIUix/rqKitCoa0fkr4wfG/AJJ7INIobvnrZBH9DK8+I3pXlw76VEMW/YYut2tz3GbF
gHfH5vgxxAwY75ZOlQogQfr7Y/Dw3gpG1NqfXyCqpceXE8p8q+KG0DFKlLzcVgBKX6cF2GvFyGgO
9UiGmQ+dKaJLmOseAViKWUE1zo6HuuOLW029wMjsICltffI2KG/vDozGa7dh8kjteWWcKPVlnmIg
ycS0cfpFrz+0QimgoEVCme8ZowQC9l8lix0tLabmhQdM+xi+LWZuOxVQLXWE3cBq0ssWSKEa2F9J
W+MWI2vA+mSAnkXsOD6ocWWgbBVv71aP3qBiZYTMBZbzpwQmJDpJ7ibg6pn9+IXiB240qEQM9edC
Gi5Anyxl2h+PSTPZp3Pphybke0HVDNeZMjHgQ7/fmPizWj1+xW+CJe7eq9NcR95qrElgh8BHdrJM
K30swFvoEsTSJH1FueQCjTb9HcexvSBEnFqvSnm/lGUvOIRYm9IJBpJljcAJZ8MBS6xELalkSjnq
rrvlI6YL7cKAvdKknr1DnSes8GSWeppWKV2XZ6mbudHVLXlMFHFRIAaGDQekm10fYVamDkf3ytzP
58sUYEjvS6gGWZ0QCj6+VfmyJ2QY0Zme65l0ElqfDTY1/1mQdvlB1x/w4pvgx7gLES2is4N4QHUT
9r7H6RhUvBT/2kHdngd43ZsvWvedBz1nvRLf36+xfhOSoo5idF1kaoloFSsmuAEFAbvEO6nkInVa
P25uuX+ohlaeMElKdixSYonztRv0ypE0FUZCMxKNCjYKbrwrBfib37Mx8y6rOjkE2frpi96gDy3l
OzmTPWNr9SHxqrhQQrKBtTzKtwOlzxOSDXRk5QHWr3VUaTu1GEBQyud2TTQYRjvJWVaTcdPMjSzg
2PiAk0RBZb5DMHLlku01ZQBX04wQ/JV0smO9ooFEJwr8EzKzXrg4UTsubeIhG5zEVhN5zgEq8Ag1
usPfVUwD6cLMv2pl+9QMQXgS3y3MyFrAmORp6ZQXLF54YgouL/wH1jsIx4oiGod5nkGzwaQFY4qJ
lgijtSTFrLKk/F9gnlmTu4IaD5se+NhAG64AEa70buWWfz/2YAa0BaVOm67XOnMeExfmaH6Jyn6l
JwZF30zCKqRGGPXnqGNePEZHJigJkbz/5AzkdJ6ZfkqrdvQ9bGAiH2SB8fqML8mdlOsCqETpF4Ep
8itNgjewJJPpSHsH12E4EL0F3xsGck/2CD9AvkT367hhIMr7BYoRGPzqRIdjupYPaBsCOd4TCjdk
114vJkq4xjrAnnJs9L2DiuljUUciBN1tc+qKc4/X8u23QsBk/n2PtBX4z90kdVzmA4sXOF6Ig9W+
L6jGDYvlZPm3WcwOyQA5G5+rWjKuwHHDnBUQ7RG6CSkNmFkH8/IV6Vgtd96KDUKh4xOBp9s+akDQ
6QBeEopJ2/RF1Le55p/7kKLBQ0T9spq4NKmNz737BHlMfpx7OH4WLyyKokrWlaEzIVKNr3npxmYN
DxgQDrwhNFpfCAT3S6nFrFrLUvOqteG4EeUba05iDJxOu7VUKM0VfHnKVfsWRPv9BemYZ2kuOlHg
8gc40jJ5lH0XtTxTbK6S0b/4ebOzf8tjGT47eyEKSFUj0qbJWSdzFz44IecynhqhuWdCdiy68MMu
VfDgUZJe+GytDZEB0bgBfKlS6zEzbo+Jq8VaHHkp9VWsvFWBPM7r55ucYN3ELkT3gLKEimCi82qb
vkeGwpyqrYZjiAqLqD0+qJhdCAT/cVrmdwn2IjWYaHLLcJ8HvtT46KRdiD6Ru5EoRS9usg3MCXNH
4YHCVK8ItfeakkMLYvwrplf26ue4py+26bhdaETmKP0MhFrvwTfCV7LNKfwj0jBU5mXZhvFEtgre
y007dQ36U5b0lg2xQSFoxbBHVVyovNETji0SDgabVlblaJ+UIaMbp3DxlNG0aLu0afZhCdNHji11
GWWr89qWHW3LPd3E+MJPuysn0gvKOM2GQ+z7cfNLSg1Nt8xLROzIstuweT9WhO6YCzJ2DJkkqaot
rMfmOIXJN/87TlyX6SZV4p5KLFeq9FXtatXJ0dOp/WN075dsVHYRx9u6sYsl4Ix2ighCRKRewmBB
YrpxCYy5rPaZnlx1JvpTutDjLBgtVIe6UPvkORWHWNVVDjLbYxroo0cYKnGZD1qFPL1bEZqkJB3c
QrFKLsX3Kkn4XFfNJ8CBiQUrjdu8tAQxg1Tq8lmMKSUbPGsN3R7i7hYmzdbCOFj3cIXNsR89ZqXu
y7QCp91uAj8FTjr6M/2635427UEhbeKFZdIxamStpR0SVbyMk1c1AWlS2fI/+wik9RkH9LU9Fvhs
wiBvS7i4P9GgLysriNJIqUHl302hCMUN1Vlypy8VLT+e2eBPyZV3Orpw2G482qTZ5PiKrZQULgEX
pNjZAGWea9ou7QZwBFm41fN5ziEvgoKbEPZCKJaOBayDFl/Ot6dZm29voP2BwybM87ff/MynMgU1
DHRN218vIsVhTZd+bOFD7SSgwUCdZ/FAtnDI/dQsFmw/g/ZXCb5oR9BMpPRBm/H+GeaExUwX49VF
i0qB/qtD+pszn2QcNMVP6MIo56pFpVYaCoSFF0H/Vj74pzqgqA3wK8eaQB/wSudQ9U4uSPcYYX8a
hCaBQlP9tPOFf6EzsjR17IBmZPgRBKvyGlgjUWZq0PXM3guIl+f9cotuq8kvifnCLAqMbEWrRkNn
jzJfbywKOMfzXZjwiFo6vqvj4vdiiOY667nA00UWAElz1kYK0GpHLpsjWPD7V7mObvlcZ4JcrEh/
/BSNtBgzA3EztEWK5oW8PMqI5AumwUncVu/VNLaseyozD8y9Xz/q9QHRA/Fwrq5xPey1Q8uN0XLr
uhByAKunteDAZ8pjkXpfe7KaTMhul8PFsl597Yf+UPkAKu52PfFsc0I2IpscPAhSWrc5miRxVSjv
JTmu2ulSR+qltYXKboeb6vKElaHL6VY/xGP33T/+0LNQmKbuFYZNaZZsks//z6WzmACQ8G/xD8uw
7+LYExgUhgXJ3LdeADoUfuoSE9OrLBzE2MmRzb6uo6drz7edWouNumMTuqcAev/D472P6D+jVYRU
DTWhT/SxKcs3pIAaqWFvK2O2M6YLMdqGu6hlON3JBpQ+IbM3zSXWyKqjaqj88tLBBDIkVTXwHs0k
vUvlnQLcLnGEKuBJAOqwaNlpG4Qnl7MGoRL0YEiljwBaHGJx4ukeCkwvspP90PX2FXoZpcquA/42
NrjlxfNdpW2rYdL+m+cmxUYFPebSdJe+4QcnnmHAp8i7Q3Ug6h42XZcLIYw6euAVuuU1fIMaDdjB
cw70z2/iTP2b8EdeLGhbbZcTnoTidUyUXN6GDkHQHDlWG1VcyNsvDTlA2sbflpy1UybgKK+a6Re4
txrJX+0hGl1SowMsM0ZaKJ1OVakTybr85vwS4I/IN8i+YMcYvyqTuEZxjIGZmxc/gZ5kohty8/f6
NMULtr7RojeKVjnvg/vQCl8hnjSBC85dD1gVUNlINRdzvYV2pcP6zikwWmt4YZSt72fZqQsygqZ8
11w29AGuUFqNxHCY5HYTHwj6IjXPxKvEhCPwdz6pmzLJVA4p7+a/Ylv7ZuwkqIqE4klG4oyVQ9Is
v+opLBtjdAQ5xUwjLQHXVF1AvLAbbAhBbnftGfGHsorgY5sKPTuF3L6MfXHmyLnmitDWlIGVm2jQ
q0zom865G+6uoORnRhysygs99yzAlNd2YlW7K/8+TOit0jCSB/Qwz3KDSGcp4Agh9KhfArBtUeyd
CZ69+IoCFY+maQI2Bw7TFrJkiGfeCupBmd//SfdUgPkehc4xhPrekVUeU7gR+iOpBrEFWL2BfUWu
oK5Ix9TZFEJabB507/NuTKvg7oty657P6ZFQ5Om7FZwPRcVlQtnulfXzr3Wy3BkLVyE/7EoN9er7
hTLG8BJ4SSs0jVHKI3jHlIIusya5aO1O24UxzQas4BYLK1GvlpUln/Ullm7xZkMIpNBD5IZ+6YdI
WkVeH7ICDdxLAvmYKoXyCMkgp1/dj6XIu6S3GMjogJOWFCU2YSUtkMJI8Ggi6weFVsNXg24KVczs
zQADmfmjruwz54JpkeDZ/95ECzfgTw+DIZjm+4++zokmygExnb1PHVg1YSqzYhH2SEjN8WGwLFcT
8DQpjTYQtlv6S1HqpVTXjpYZLvJC5kqz4kknxMCNJnEwWcNlblcoOGHsRwi+7VckCuWzNz1zbGOI
ZXtp1SVlZY6aFeyWhQOm57YJtFnYwKCqRRkUTNmas+Kkxx+W4Bqvayn6UY22VFAB6G66lCvdRbnZ
1KxljbWuXFjECOHWEL9mZZb/3YJBSdg6umqfcPqRtjlOtGcQSPcgI37uH++EeBCRKR9621lRrQ3F
t//lfi6Tz8uobDjZ+d6K9jqXhNvcBkN90W2CVAI4MCvNXijPEfaJ6J69Hn/r+HJVVik7GFvIknTz
CYa4hSiG54N8ahr7tSNIM9XvxMva8KDqyY2SgAjpY5vxqHuJz1LqHLiDTu+cdTKwgDDT33toOA3+
SzU3w+6qDrxaKEwzzyOU53e2p727lwcbtfjxPqxJnpIgN6ws1rHlcNnD8DVGsl/20YALyipv4AK4
6VGXafttr+AILHeJaPebt20trPORBHj1p4w7TGA0/rkjkDTVb+jc69sCEIcnyfYSXbtq7GTy122V
hwYxt2438ZOuTsgGtJaHJr/+YjbSn0NeR2ZMCaNs5nOeq8wf2i94Dxaw2egfMiZ+6tg0QamYNEeS
DNt4Y3SChWIelH3Bfa3FUdvYclhi3irwvHEpnFUTfRetcnHBvt1JESm4rED1gbaZ98+qhMY+QEMQ
blYCqYz/1QB1nGIBghWow8u+zILiNWKu8jjQLGl2W3nEibc5qtO35kQrjjxdEid09KvKzFP3imlj
7h5yOdFeRmNDio2rtLks+iBafYoyl//H1DwI5sNnNc1qvvChkAn+As5YwZQvTYFQdaD/sbzk/Cj8
MRCrcKGbuQwZkQHxoeHFhDC2J1TV5X/Tx0LsYtJTdJvOz7HtG2hjrNPXShya5qAAS01NTrKnWyyg
euFGkdC+n5ybpFSV9MYY3HBf/tEJy8xBVCVXCNWeRWncJVNYTBOXylU7JM+9GS2R9kKyE5P2p4OI
Ku52fHJT/Wc8RoTu/5hQYYnWgm2ZIEnYHrXecrxy4p2CPIT/Ka4nb8W4fLCeNDnRocqVxacsDmNH
juLaAhf8Lh0QyvoN0RicGltMgE/+mogpgzUxWgh7e+h+cciN49U5m1GgtdHPCRyfkixhiQPaEoxE
Z3/BUVKya/KL6nLXYCeJz/YKAZKq86Ecp4y4h0UliwKkkBHhg+XfplePp+lhVfTMp9fOMoYyrOsm
3C0Hhw+9t6h1ZB/aUbDXDTnJzooife1b71KzCYDxZpWV3NmmROslcRF4WnRV766k1hAbzp0khh3g
7nE8zFTI8jXIY4jkkQTlApRPzXGSMD+GO4i8DalWHFHei1Q7oPiPjn19CrXe9OGNA8CJOvmY5Lho
5SYwwyTscmx4LXQm51baCVhqFFVsRGhbl7Gy79e7qlX1HjRYAg4/XYYjOQEuZJlJVplotIDZZ9Yy
wBNHd2YlLPONAQOckQ9HtdrqAGjnj7Um/ZitROCIpAhP4LeawXlAwC96Vg/jal5tyBwe54REJWBX
FYJopA2RURQwAYivBjJJINTGMS0lHMIrZTU6OakeOdMXlYcWDdGUxD7qz6gTCq0/w8BKFuoY6ano
/62WvFdyNi+hU/aIcrzYISAzIlAc8tSqRSulrIK1XtSvwcJ4eMwF2ULOt3CN9PY1kx9I5sCSGezs
YHlDLQcrwNcFml11Q+Hgrrpjx7siwkcP1SCGNqfdSJlCUWphOilZi32UL/kE7sHq5mRgq2hrkflI
WP/ZIDWwTKjrubFFlqhakJAXZt5Th2CLZQkeXwz9/IAfHOU0MD5DY9PgmwESksMN0It7EmYwKQ6a
udeWDk6Fk6C7yWxWplI0NemwJNvX7f37EYG99Sv9/YsXOCZlIU8K/YrWaUTRifXC+GiZUzZ5gTas
DeCzudRBnaO/Qml4QGaZALt1B99/ZV0c7zH+kDbKC+3lpbm+cRuxQYneAc6flGmqhM9jPCqK1Rn1
MUw5LbSt0Sa8AGHrT0qlzAJHWeAFllycfSBfZWQsG3DedqCVwJGdnuX/jjq/Zbvos60d0YTSy+aK
jOhmnWncmktOuyxY7eVxmVwo5VJqKlItxNPxLIaiXwKATCWdXe2y3oWAk8Xm5dW2HlRX69/sG6rF
cLLbKpUXtLlubhORzg56UtAbHqSBBTGUSdmE4gVO3vdh6x/DSalOpD5F7pV68W6ad9T5odze9e2D
EvmffXCaINbZMcwGc7vO824m2VScijkas6QVYTjkO0kOKpHh3tGVUIGPO8I2pulzOCwjTdL4omaN
rUAzB9v696vXftXk+JDvdfcMPt3pb/hRTFMewDRxWqDGmJY2HIk5JcFwPGD5lWATjYxoIfq4nre0
KLO6Iv11t1jGEXWmeKDQ94v8AufM7Ljxu1loruQ6blIQmJB9EP28NWMRbOp7mcj/UgJJgMWRqE+Z
64t8S7olu0+Em07OYlFng2p2O3RLv80DpsIHr6l+UpqWuauxyRBCWATwLdE5vbKwAUR400r2YOb+
IWLB4L8pnWiaARIUtE13kO2fMPS3M/qAoW2gIHzx5uJTcg9hJ/thFvL186+2uNaFK/PLI78RwKVK
fhVJOngRV6Ukz9WkMDrbKUTcIaOZ3ZHh68GQX85x34B/5F1F2/PcwrKnICjsCFlF8i35X7Lf2KOr
/9mpZjcWn53iIodbPvmHegPyn6+pmdv84XjqIJKXZ+NjZnGF5l66FhjAU7ffQLmaVzp06LZ5UMlc
NAmQNwrCExr4OCFeTukSMtDc6w0GPkq0YhioK2Fgmr0BwyaqA9EutuUUpJj4LPkJoeun3zoyTDsn
QPlY1ThavOyI+TYS4uuuuvZWv0BuWFjjClBycMi1h0Or1B/DWd+PaRBlAo6aaZVFHbZBD41nVB5w
6N1TFy5ZtoQgyAzod9ze/uRTVX4pO4yleiD0XI9CuLGdyfjyrRtXe0fRabrtMOtBiKeeWOkN0HbY
E7qmNG04hJyskPmat1in/Gt3ufGevxWNznfoPUtbLoE8gosLrzFqieEuYwtGCUnki9MR1drvrFiv
FDSwAZF87yEBhRjO8UzLpQcNdjqfOD19iptKkcPy5Hp22U+KAZxyHgL38Y7j8IeIZCQm4MTPOqQc
LX7SgdZURTBTiaGTAYLOB9lC6QEepy/nlV+unZiefbiE8pW1awqRVC0R45LhjEG9GcJeK4MlAUjO
cun4z3Q2JLah0dh0+bAvZe287HqDNJRJPkSnXX19YunDQxDXwLvYhgH2yDTKawqCgUQAGNDmLX2u
1rbTIWirQfpsrk9Avlg+XZta/i/Z8+9Au4kix7tyvXKz/JQpO6tgsC6OQ7kdiO71/EJCNWfinynY
yzZFtabzQqxYL2w3j0omJSLUWrIwoQsrEV0Exr+em0CX9JGgedMYIA+8MfmPcr4NZD7MGDRVuHpl
CcU/XO4zMGJZSOqx+Y47vAOddyMMwRJxXzdFj8gKXxtlMGBVMPmUD/skhyDDyhpmb1nnLJ1goxwC
tATgLJqsT/DTgw0uEABDaAXDcYN5f7Px56J8znEErVCSZ5MLJJX9WnSppHbXrSr7Rev2+ni3W0DM
ScKm+TXklKmtWUl6VYeL5gRFY3q/FwRzo+jVm/SUnjbtsc1+mvCxBn32yaFQKsNqP9wj56aSOABP
if83q654j8lMl0yKdVAGY6OpuBElWiyIGNZtljZGeFVCh0j6ajpwqsocCItQWrP59rIK13GGlljr
Vl411FfIiwzExdONYQty9Mz3hj5niPAAbsTRPe2HaOSTf3gfUOOnvxhfmo721LIlu8sqSPmYr1wx
1LacYbyC6RLWtnjYNkh64Kh4IoSaySKwFIBPbQlJOWftL9ZJTamn8uZyyAxFpnXqzQC7eeZjrcMX
jVvhlvUeOHGME5j6bhM8DpEcfSZXKrbw2RDq0dOWWBdvx8iL0Hhj9t9V07zfhgwUP1CuDI1kcmSW
vZtbzyzvKprQBpzgtILHJX+bmAZi9tKqj2qWtUaRjPODrMNDuT06HANxZ7nGxLa7GsOl8MP6cbJn
MQw1+UCHjxcAsff4AjJ8TbopeFMLLM8E8/yXrCup/HXHwl8BfZsB71e5CeLD6JsBvWLMbPGalL62
AUa+wXEydcBuGYGapXGVxLkBwwCurkueMllAwmh32zcqkuugw6vQQrxqFUjzmJuLy0CEXV0jbrbF
nBovT4ONi+8dfJlDxhdSm02dnJuLxHOqbwNPB4FCloVjZo5wp6T8auIyM0SKikUHBZcKUSpXHjpx
DZchIDn/4xRtWT90MDcirdoTg1/1YVflmLI5lRI7yOFDN9rCbCZ4fNvCQzu5iT8+MANf7w/W1VrV
aQufKTkx3WZfR8YOKZTS3fqJw6sETIFBIj/a0LzjqzzYg/5IVRDy746CNPeRvWcTjcYbY1TN+SVU
OcxqnhxUNIIvc6rPee9uFfEC7BcA1JIr88SAFPPzVMAKrLl9heeucZ1kDwCua+u6e/i2cR6L6g+h
cSizhQ2arUOSSw+6EvvsqhUQnzACQZkRYWig4lXMVUy0CcbqSW3e06AwSe/YgyngoZM1kiwQsDNn
39N5jf0vfgwikB5psYXcSjzHhDOfyjXWdqL1tFLW4bMH5Xhf99plX6P/D4F+LIgu6goLBMzuHr+X
60daIbQOFC7JHkz7OBukLHTvL/u3Cxjs/MDX5Pu86Wot2Zv1hzfp/bmWLh/+0mvNG8rF/jSnSUxB
a+9/P7gr8MSb+9/yb0KU9Bvu96A3uBwYu650SUbJSDOXVMLLPyjgPffh/IZYmD7cBuLxrl/+rOdb
zgzvWWrXi9JAjm2wQr8EJb0t57e3Z6zUnEAb9mxXVQXxM7RJxKjcvAfhKmY6u5j3Y7TY7ftexx6C
pGyaYCGDI2Q995rBdwOVyDX4r/0s2NOV6IzhYldwg4TrBPOS806E62MSp1RSBS7n1o7ES4I+VvD9
vkWzUOWmoH1w3teblNtu4MS9i6wDM/H94qYg/wxflsvGddu9N2vcDztUBC5ReEy2PGdAaqW9OOre
TiPm6R6n4kraaQAl+AmnGWRxdnBjWKkQ6DIEyzEMWDDeMQMWH+5Gx3JZblWZoCapnIBgXATBxkIQ
axKD3XCI1JTq2Yqc0O13+lJFpOwdrzkJSM/9LKGmXBGgOb01D236pNXj0n0kz72zCgizQnTXEXhg
CoHBzPFh9Sy9WQEFek3hEIOLi6PCCjj8vaPhoOAaUDGH4VlqEXz56qq2VuIrdZo5fY3iF3xX/Njn
gRlpE4cjhN3g8XbV9MDi5VNUpdn1GfNtw3P18g3fiS1XAOkTcpKMoBrkEPttsYdIids2HGLIEzXe
v4+Xc4CHz9zBO+/IvyHbCyeeNQglT/ka5ptzb3/O9+G7PyUCGggPwfNLXgzLYCCMCNNNz/pDlv3s
32HGiYF8Cs2pGwpV9+m3NCQxZGPFXkP/2vkalr2Snn4vfpJCVLJB2lTcKTfylAqs+jzRIGZAGA+B
rRnU+xCgn7aKDjzcxH6RhicwhYmk+FeW7eFoMBO/8jRNv18Lf/f2JIvDAo/mFVwSvU36ZxcRX9/4
d6hiOlGw/7O/qdFjCCioHZQVehGqviOXWlfqSVhXUU822TOQ3ApdjN3b5xXTUJQJdGQyf7J7ikbj
rEgUWGmUYlDuHUrM6tepRGf5eTaTYao0HUOztsC6PvJIpkKGfNVMEb1bjY2dqyqN5v1t2EpXlnHI
g08r6sg096P8u3N2ExL73xjtMo0o3zl43vgsrITLchUu8OYBvOMDIefq0qTw2v39hX4/uMGklPJY
uYXl+3jtCu8spZt0AOkdjk7uA3vTMVGAR/buczfL9u+kPbNcsUdNd1QYYIxRHPj9AyJMBlz9Tfrr
PwzxgyXTjWUwfSsO+MSeiug2Lopy+cODRPn8x1Ae7Qska9npRqioquOlqqYuWdixVmbie7DuX0lg
L+vW3RQAGj97wC/h4nn8ensyOVh8WGMChEBizdVM7UbMr2WKOKOpuZzqCVHh9FRwpQNPCbmR9gQO
tblKRNbhBHlY6agq587MghAFaxuWxsYcB558/od4k/H0TJkwu8QjqMUKFlOH5h89lwg2TltqoOax
nqzHAQqUPARZMJcviAcAtNNGGxlXGlTATWjNteySeimI0yaW8rIxQl0v4X/SAUsZYfoZ8taYN4Ys
1/WTXi/1ndMxO7bs3Jp1owG354bUdhX2wQv7YzrgCN3FogEcLMLfB3hkmHCCiAWVlh4MEPR9CcWI
xFv96Nq7o90f2HLG+Ad/tMNwHbxvXoBQLxDo2HAEHQHTbt+zuNgTxiEvEDHj5UMVGJRHQjtRf6gV
NV3EcC/7eGgp6PsUlqtvr+HS2u/ULtS0Sl4+ykOEFa6LflhQU3NmS2+GnW/1Ze34wP0tGMSqEgD8
qOqDwqgEHS4Z5iUrpyYzolc140/GaD3qrnlwK1ybPei0lEYJCBxLKqZH98ZBnNtyzwbbZ/DP4N06
iA5TCLV8TAOdFfQDvPrpgx5+ThcpuYpPlouM6tgU+BJpqkk45HtBfHb/UQDEoR/XZCChRGvouaOF
dsz+GuKlH88gPmJF1aN/U+8pFI1IJaw7Sds2elRFpdC49L6f1IGqVhOxqJifDpEOe2ZWbkgRjCm8
oKdVMl3/fGhjGUhfpBmf4iRSMqYLL4AT6bpRSYXKBNI9oyDvj3D5JP4Ab11+9diBcrwo8VvwWWp+
W/VzRCzVRKA4BfIWIY6lniktnu0evWGJ14wp/ShqWNGENhzn6HK67rtwWFaMp1Aga1sjFGZ3hQMa
JjBjPw6recRIS0EtjCzpzGBqvj5q4UiduAWwOpzyxAXeAryZ+JGi3azKofCii+i0od4CrijsoMsj
HUI7SZxggd5QmygnizwZ6tVHay1VcD1ravcFfLSkYom/jiuWHAINkk9ph+SafsigqSooS3bH8yiV
ZEQ/F6Q6MHFqSis5PuLEIRJUJzhNxWvA5DpcQA/bpHAPrivitG7HE4O/wzGZETB8vTTKFo4tZWjw
UiuWvOquOq7QeiqpfOsjZ29wcQLHg3PhpgmOxtKcTYdtLC59SvtKv2BAnWbC/FmXyk0HdorMCE3f
I0kM+CT4TP4VsV5fEdOHtAOiaKNnvNZQhWZKJxUkKWBlhLYA+Rf896SfiXNPUZOaBbynXu6seT4X
FVh2FEb7xcUFzUxie1rdD+ni15hwb/+cCQ+hS/RV2f+tfY4pspWZav7XtmMfMrvuwyTIk1D3v7do
sFwQUlYWl697ugxmkll7fbw45um3FrSlFgc+YqZZ7J15RM8nf4HUASwOLAjN86+jSdX8A8Ffr2b+
DlZEvredLL51TjB54l8h+IhD+iZEI53Rh8/b6IDEEiFF+yY/IFA5LmZTCr6o+s5M7FnXlGf/BBoX
8s51bAmRqdffZsYytaRq4E/UqJeDvPwiA8Lzw4wPEqbvx592RV3A7qTz459IgiFV6n6x7uL6RGPq
aDNpjlexR32EQctlJ+CGK5IK1v4JiCu+vX0DqYrlnqb3SFzZdcCQ8seGqu19O30vv3Spy4kUkcul
dk8O7P/IVUrps8dGynVUbI3qaA7VjD/VrRGV/5aQqbCYs9N9Wt9fcVtD63vRo7dE8FsVT3TUNGQ+
6HgnnkH18fe53W7fbefNGeVWMq72UihcnOXOoWXO1YhY5gP2K5lR/WYcavg0Nw51kiKLH5CdcVNN
+gwUDOvqO5/1j0bu1+N4Oi08qg37biVQB3oK5xD9ctUp34VGSadvtuHVQd93QCpgV+/+pEodR5so
J72GL2DNGtl1PsGEg5vGVE8Ff0ZDYhtTMZJPqxgK0nfLmztHkNbu2633fEOjphcLEHtJ6KG0nJCc
P5ODQreHSvkK2UlkI+nOMZx4elMowfS/ZM18y5yJ71uyHWY/ZchT38tLNjM+NCTJ+Fgq5djIDhoH
LZQXKS6cvLA1i81I8pBmUeGNQMGIbswIGdgIB2Kw3wwrdkzC4j4xVim5lenc3WsAcNh4BmZuYEjB
Tprn0dQ2NcYwrhphBNwY1YPToYI5yBpPndVEQUveWnCbiaQZu3uZDtCH0ZGRkkR572QJaWCDrEAE
AtURdz83XxEH71StTnSwhH9ElqlZtqQYcPp5QYKC2nsNkhtHb3wHyZ0ErK4YecNpIx6WOQGIwpAi
R9q0YWbzpuIpxL4AiaJXRdWcMYBcJpU/IuPhs/IFA3+eakxbhFArRnvKh7MwK/sqcf/wh8/kELtO
S5MlMjzWdc3qkJiEQjJPzaPbNkHWKD4gJfsZDn6oNK927YFwLB7XnmG5vDXQqcdhBDk4c36xbvIC
umWaLNKfhGfvU5HIHl9kL1CWzyojQCAQDcuTZEnAuMdGHTVnOMEbLasxUtkZaoSDQS6vAv9/nb9C
0e3xnRQFZ5ap5E7hiTxhURMwcMxVjDaI0edqH66XmG3juF0bw+gtOm3p+ixmSWNROQz/KuTo62uc
xVNqrW1lHpFfFi5VNCDuPKEZU0+XoZtJUeLqDiLzLCLsnAW1zTV1iNd0i4hRJU43MjE5mx01WgxP
dYRl7grQhUbQ1aUdFG1h0HisNrZLVM3eFriwVfTIROsDX3Mst+FEbm6ub4ebwgbbFCU151DlaNDI
AWS1/7EfKOCuuPjgfl2lHzo+Rz0qOH0r8LvWVXXbU+oND/D7R4IxPP2K5Ir6UzJGSz3Kleuo3u9N
TzO68rBaYqZlT6KDS94ZbALFZpRwIOyU0LeIg5gypB2JNpD0+fak3Hiu3Ux3Pa3kgTqwKdKTpsZM
mCLazQHSzjOoDMiczDlxqTEBFgFOCHh4YxphfqrYX9OOy4xGiBJq4vCycME2D6bD3v2dn8I5WODx
h6Aujz8qtM1MilVqcVH9CalZ6j72qGoc7Eu1Gj5K2/hf+VxLa4mOcxTRHxzsIkz5ug046gEJ3siN
SpBbb3pr3FMpk4GKMo2GY60AGdKG9Dr5YgpJ9PUKIEC0aBjrm5qz69tu7JNAqobwLNl4XuKcm1Uh
Ug7f0GQM023Iv787mTnqT7Izj88xISm3WvpyQFbwn4O1YCgeBBBB+z2Wzu+Y3SC70mV9LeGmulKb
o/5vLNICzYKqupuBSsLaZOsNTQQUplL2dPS9RhRWSo2qke58r1GmxPa5HZkPhOdE3nmYjn47CA5D
BSAVmlvn4hFsXPp9g1lSHr49F9/BgFBBxO49gvadS2HRrs30M1EAIXFUCaDZxaTyaV8EIOS9V27w
eIdymVIen7ZlQ4reYMok4h15APWZ3cBnI9c3uvKXloH8MENWBe+MSXTHfUm2+7l0etR8f5k950wJ
gNE5NCYGH/yojKIxuxn9VSWU6AKt8f9C2WDO17UaCLPnFDy0G1faYDZ4C7kVJRNR+8szQ+2IwDe3
aXOuMpj16WAow5C0yKnzpGUXX8yU/9mZRrNKoBdAShgaCYbxPdC4UvAXzyuIBolis64nl6BVSOZg
rHpAord1iQJuSpBFSHfNGvKbczOWE+Yz5cU7uFYDBl7kOuSDPotb+zklaI5vfIRYujFfPZfhEp+9
rhfK9uqgZ2uC1eisBzQBJbl1dbC/igyHAZneqjXwvzgSDZCinNoXlHVeTW6uJAnpviJRVx2QOxIK
lP9atf3OCw5gKejxufGlnjbd+vLUZZfwtVowCAhrdRU7+b7s1TYzjoBTCWFffsfabEGbTsWuy5In
wX164MrLlRgSFTKJg9EzmKNrpvcKx1eddFntMyQ/ksYIDXbwDkU2rcfbHW8E70hQtbmfOqowzeWy
OoQz+UXpjweiecFahOdMm8x0sQBbkB2n0zDTT62XObuNTYV71JyYAkM3d0S9uzLhuuMRYy9bgAhK
ehRnGVlwcfzQbM8p1l9nzI3F1qowxLiqnLD+mIYi3bpyvoWcM9QQfROGz15AjiZ0jh4+t+tmLn5i
ohCMrUmbouNc2wMdt/Z0oPalkGj5G9rD7q0m8Q89k00/O/qCxXssW3heS1v4N3XSToTaf3l9Hyfg
Tty+b+wwjdYINnaFWTRNiBD22ilv5/0Vz/KERaJhZ3yu+0CtDE7gHQoRO4sUWomhNr+4PhRK5LT+
halzFm9LUiZ8BRA/IW3KmSMgZxilxscbzniL7IKftQHTf6ADF3/AbzXWRlzIvmKXoznODxPlojDB
P1ZPFz7aCMqdkQtVfMCSpMleSxOwmFZZ6H7wwUGu88TIVQBZeD5rJ0bQNQq8jtPUjUwydc+2oSJW
uhsyqH0k/PrM/e3KZLNOHgMlc4iAExEiiKWnG4iV5+FYT6QOLil9ajafUUWQ7GXAoN0Q+Z2AwtQG
kBkhnbGPqmAgd5DtqqB8/8adxP+cdipU1TdZqY34dnOKaHH5iIK3m+w6CWgX40wmBbgaWLRozXsC
2p3BU/pF7NRx5TU6VMsN/xYm/AE7PD8I51dM9X9SFZWZOHbcq9IX8Wzfk+EamDKzxKLKb7NW6043
tuD3/Yikxndanx0TpOGJlOAmJ731Qm7rHFH9Frq+wtVdjAgWU+fX8tyA6suHKhdSD+k1KslDxrJ9
5p8vmxzKRSVYj7dJVD9HjWQabXwMNLUGtxV3O0PgAQjDCRBUCaZ1UZRQWdyV8Bb3mNHCJdYiAqj6
YsZU4xnvwT5vb6DK3Jq2mCyUNiYRzYZXDRlylNDUQWV58jqzGyQFS4Q+bT0KvFZYmr0nOgIaIgQ+
wM2By1OMfl4AUKdvus6I8yAI0CHkUAb4tNgNEOdfEc8hKX1n6kAl2xJVP6VcVsBz4NLmtlfmwzRb
kT0SWBgat80TPeWffw/X/v5yYjTmw7NL6FFJtAPgIeufuW0bR6SwKyM7Xl1vjTqHGOhFtPUBe5Ua
Ubl5tbnHqAyt+WdRYdytSHJwlGluHX7+KSOf5Y3+oCSb4gg/wS6tmJFyi0YhPMaZswO+uASVQCGq
yNuj0UiLycG2x9Qa7VogD0+Fd/7+iGWxRos0K6YOLs1qPK6UT40ukNQXzjdbDuqHs72chX2wPOQR
FRlBW4UVIb/Vc3ZX9KeeeYD4RhyLqJMuLdPASe5YfbKmrmGqK+e15uszlh65tirF4Odskhc9KySP
xKEtiKpQaIcSMB9Lvb1uKfLUP6fs7205yfnWrQD3ZGO55U2u/lkLjLPyW/jxM/zzBy+nLkc9+4rH
Co4AuZbuzTDai5/mchKYB3PUY+75dsO6kfZkFKHY2FefQ1bIU+dKI1SLrpWp4oAhau0aq8i15gAu
xXPegmQmyPsomgzPquX+V/6p9jQyP8PnZgGsHMAj0Ypxnes5qPk3b7aSClCXvsa5veMoewU3Mv/9
3gg/bzHiK1TSc/IAQhfjTXdHTf8Tdql3GQbVSA1zfjI+3zaRDnwjcoA3wh5Lg3Z07q1JWWepoPyb
56RjfeV39kFrW+GV/8mgrugSTdtcD+J92dG7en1uEbvj1FF9lZTR/9AHj1f6a3jGoHmfkfESpwkt
uCIOM4LtP1811OOa/Y1AUgxeFMvC4F+Nu88y5XKsrERFIcFKPfmkHXiviNF7L/TlNnZrhOkyMqPt
SvCWzOfcWyp+UJm43jmFcZtImYCcZPWbD8aj7RzDyuSjM39EHr4BXIatqBbdNaIaC5pzc0jNeXxK
uRaiDXWgIcnDsM5F24irCspIhA9TMni3FKjlSqrmoQKL4k+BUxbYgNGm0pdNzq4jxpZ7pl6mdplc
NbWrHlK/9tQgBRdS5dX/xES0Iv7JDMM7WI4Mk7/efTRMkKFS1PzqYDU8H8xVpgECH0ix53vlhqAv
Wic7Zf/BqfC1GHMz2JT8i82AwcWJjhke8wwgCyBvJL3/PEay1FHXQKirWHquk+tF0j3sOCkC8IEM
dpTRomj3IHe3/iiEepemixP5bfV0IQNTdjNqsaSgRS45o4Ov57u1KQGtLudmt0dnbWYzCvcixT/U
n34+amk2XIXfUdwhbD6lFylfbkqwRRrl7GH/eniYPmn0VH6KdzC9SlV1QpGGuvVlxaai3xaw2ZRB
f30c9rZBD7tqKDA+9S2dgOlbxhJCux7O36W1+PfQILd/Fu4RG4CmriCGlEuKT+73NlpBeykT3Gwb
o2bM/ROKXkGYdlNYLkmoFoSZLhgRj+fvISLzz4GGOjAE78H9GwDffw9lztPA8xGISxk6/ywq61iK
svM3CPbpfEdm3gYwQsayHjJ9S+1F8AlhzceySJIXoUxhBzbPHfyNLEbzoprfzhL6UmdjaDqrJVhL
Iygh1O631rMiGahwrpGpjQYqa78OVUi97gIGZ21KnbgrBucNONrKwbzJy1VAur6xxqX+Rk3inPo9
X61cLlVhyWgCB6+NoNxjBI2QZbFvp78u+gk7c9eHCHJwmvJCuVkzk+BgB5dghAxULDDvfwCo5/lr
AGTYLis6IBPjNbChQRzCGUKQkbIrc3fgfBB36IfhO5nFBiOVk7kQpjFSTiyk4IKmlIhldW2Cil3M
z3qo+BA9w5mVD1ncWDd/g00A0fxGaFNpIyOa6kVTncdFVNO9eJ0bDQ6tnHu8+wuhzGFOFKWJSu7i
OMlMBV6vXErg3AvQ0m8dSvrRuZN+cl3VWQOIqGsb3qwUJf64Dtt9o2rk5OoBekdMhwU12ILh8rVo
6M4PzlheCj+hGszt7/iWNjYJtd4H/55RYuIqNlJuNgyTgjQ9XV8BskY4YFl2xmesN2c5mo9wGv0s
SaLY8eflSl/abWCEc1pfZS+S4h32Fu7iMhjmIcro0n27ST4cdid/yCLAktJCjIi77XF0cx/DiUHM
y3BnEOzsMp7oOseZXlNTd4M25WRRL5aasM4Kfj7mpMFJ3xN8wImaUYo7kkcWZ5qgn6lQnR0EYqQs
DxA1Kh4RivHblYUfdcwTqF3HHATOyTnDfzjQumhM3F7j6BpeIrObbri+0/bmoG9MhdHXWpj8mkWn
Pt7f8X0tnFuDCp2LNhcj9t0ldk4da6mD6zWJP5fwnrpdz5MpwLuTO8x/QWWeVe2PWOEfXX5GyGv/
GGxzwQJ8KLJTnxD5ekQj2Pp99incnMHzonnwwUgL5Btc9uzTVWs9l00UGtkwORY2e5qpWb25g+8L
EZnicuOOfOmT2uSHGdjP65tFqcQ4Qq0ZPbExhuH1gNuKTDNBf3uKGFScbNC13CxhwlJ8XtniBU10
Ab2Sg9u/8lp+sPyscJIO3CXm2wjo0hVjq0nWufSoWksnl/gFQ1U5t6eoMkPwG7Heh3Qtz0VS6lZ5
XJ8QVhj3T3wOTa7oXP1fmELU5H6BzzTSwctY28eJn9hjlcdAiVmyhPWSDNlcW+FLlznTwhYDafrC
Bf5Q8f6Z1Zil1Yz5CgGhJqM6lmBkNnh5QXQlw8PYKEHPVkhXyr/LULaydMBtc+1dacAfuodLSnCL
LsSrHoDZMReo2dBluyoGEmUq0R5H8hqXBCH3LPy+YwnXK50p/ZBfN8pSOKIsfnrBtLpSYlY5maEH
pfJ30q4CTH5WgC6S08WWscdaTiRSA9Sd0no5oVP4UGpbBZfHnf95+34zy8WWISzO0h2R+DjHVNcE
JNialx3SKlYBkGP4qV8+LkMyAa4fXrdKhPUzslyXWhK6vYxHl1VVw/EfMXlkAK1kfiBK7eA6WKO6
YuC7KM0Fy5Nr7k2rkfOeZSm1Wi07SuH0rqZSYDl7ZPqn8S+VlTursbSY4nmacdsM7vNbFTX6Fol6
KKZf6Mw6uuU+Gyvctt2AxHnxQmd7iQb+a9/FnpSRUcJAaxkos0M3WrbbPxApNV3q80C0Ah70KFA4
d7ItAjkMXKvQ9MnPDrT9zNEBkzsY9bfezhJwQiyB6YPdnNG7gxXLvnUApg1HXBJe5Zdnd0h/mN4W
WumbllgoIbDxpLegaC5YGJr/EifcqCF7j4w5K6AhX+sgBILq1HJ2h7uWjQ+4tJapGi2xi1olC9l6
YdpUOlDOT88lvemopcIm53Chz/IFPoPb7Y0V3vBoH3srRNvFtvk7dheVRC4FWSs2NiGkPxFbfS08
8ZWYVdA0rcZF9ybZvXwqHaWhEFgXCZZSCYUN+m7J6fytAnKm7bHPOsZZVbxyxJSzZ4aJvk6TAbza
tWYTQK29LX1s+wXbkU3d3ewFuUQ1rAp22YCID1azzka5zI9BavsilMsvYEojkQhkSaJC98mJ6Kow
Fhmqy6IuXU906kBzPJgLjKgR0PsLObZLdlkH+tI8cjJfHWSwG6NBLe0BPYXesW2p7AQ9D7dOtw81
FcmDQen97YvKQgG3v+ooRxrI39IuU6myI37auV/X73MUeigdR8tNdqojGLNF+ZIGmhYETR6mFWKl
pbjKVwVi0LpXizfR+Y5N4nSAFiPZh0DotryMcDpyGCOJa5HFfc4iMS95yvKkUI19FD9i7nF7RuU7
tEyVzJQJJv7qQUWwWTtSfW45ns5JD4X70zMv9cW2C6N2HYKdSJfg7NQ4NRuGkWlVMQJYpjD+goGl
HgRtRi+NLOjESpB/2HQZT5ZtMZEVWng9g5cV3nLy+Bpze8b95hD9PG8QQESnbXVLFj2vfSBPH773
avXsnD0ZhmzpRaqTItdVeaTyNXe2nZJqRfruESReUPZaA6lQidG3dH0B6g85H+LVb+xfVdGRnydL
7Y1nBR6BkixPooCSyrFJaWHJxML7JX4J6iF8M9BE+He+gC83Eb2xej1WpW/wb7KS6rvCaf+vFXJ1
dEpohYv7WoEHwI4Ma5sYyOo9MPAEC91R4uypdh+xrpT3w2egjm/HHfAnV8Ixh4uhpF26QfRDufvO
gcyXpdPV5gm6fKOJotB2DX4RlTbju30pvlVM06TXMtZnnaMtfeLuLnpJ2lBOZWqGkNJGCaKECfyy
JgdXJnb6vHUA4Og8hnSnEhusLyffFdkog9W+qlKhZox4IEPvqfYmRA6K94FXrsXM7rmccPcnxoDq
rrFSuFjWBK6cNNueNcaUVr0PO1PpW3M/8hHlPB7ZdZvrRaFEI69vrkqe4WMC/CCJbPfdJteDWO4h
nQWwOZ4odaRqPfRS78aYlKRsT0wvM1VUeNLhFAwo38h+QsFlTX1ONJoFzMZlCLRlrCS9hacCjKUX
QCI2fJ1i17k7LLhZBoZybLdOdpBG8dnowQGAc5k1Jw98dsWvCZrjj4D2a9pCKAr+ayAsdYzwLPkl
t7JvrEmsGV+org53Xd4GKTXP/16BBA6QtCOHK+0W/8kr0rv4Bux/dIkOU87HUNGPotm3UWwkucqU
NjwduUm8MJ8kB6NJHRJeBpE8ZWaVWLaXoO9vYRV2F6CZLrrzk5NgqKip8KnlmX1y3GaEKW5M90zP
gpVypjuLESdLBWJu4uBHoU5yPFk30zupCAxbOlFOq0yY6bJeuOZC8WjjIvx0gSzM13+utLfY+TfX
UB2W3dbxHh7VZ8GvLUH4DjU8t13NfXX8BNnpo9+7Mx5H0pqaWwiDh5wWJuGBPfSRzjIaxkjqqhI+
5yk/xFL0OuzIwz9Y3sq+qG0w2BR7TmcsNaC5hOIN9GilMUjy/9vUToaUPPBElHTTluZPY9JZGBQM
1newjuR9Ix/GtmXg0y2vAvoHS75VYjpbEswD6Sl5v0+iBWBHiEJ1BaPlEESWLCWUmO9PzPnS3rLb
X25RVaDUDK+SGfMBTDEBvfOyKmRA8TUq3LtCkAGmGD+sex8cQuxIZY/lMqZcn3qfRgvTzW1/523K
qYD/R+Sprlmzyj0385xny82EpfscwzFMgTBDZeI/Oc8nj05jRLJpDAZLyz6p5SqW6VamQmnf6his
GRGab0nW0YSzc6T55Sb0st/ZDLbOweFQIIusYesSTdWiyd/R1Vd4IlHggDcpm+0c+gecBmjPQCQ2
GitLPab1+uvpeAwrKe0sJngr0YVT53lzgh8QaFsFD679NP45Xms+cbsQLnm2iGSU1Uw5vly04kjm
KuIfOd/q4/+qQXFY9nnRm3+t9fUsWLWa2eT3RYgRPFPKOxulCcCKPw7So/hcWlhqCs62/mAEKOJ6
b6wqqskfjakDs3S+cqm9v2UyU/RAmRUt0oaK8F+7GSxL4ETcpoqGs+D238+dzSTuQFy6Uot+FhEd
1DnG38VCtw/U0GtJI9HkGuTjNvFq9WFqROuks0+e7oEDneQfUwYctDFDMBbGGDI3bIun2Up+J1fm
JWYxXgxC7NqwAj+ikznhINZiSPxRZfZG26FsCg/JcL5gTVSR1Rhb8rOhQxfkcLMqWbLXqk0hs1S7
yZyVn5RHgPjZM6HRnWeCtpS0CQ+LJrrJK4K+e2ZlR2nHYhhnT+tQX8XouKpSg3EV4UMgH5pR2CaO
u0QruMJgTCvX6aaGOX2YOICy39R7qKMnzF+7fIu7GV//J1J6twkXjC5Yfb182TRqsqX8x+++YcJE
secdww2tGTaUxjf3qHSEYsMkl+Fix+qmW/TMtfYRjaspWZpmm3lTxyssSyCJ0xFDxf5VJqKCn+0L
tP3H3zh8tuMGx3m2/rUmymqklMu2KX0Do9UiXAvbUUXAbL0RYDONraGU3EG/l9onZjwPYi0ByNeh
2X5Iev7VdOIUhe6QP8qANgSiORero43hglaGqr/lUaqIQ+wa6XhkYGCICkdpCmXY550U9hZsWGUT
x0jBhg+6Xhro6dhvK/C7tBrfSgivQgQecwWfNJ/5ctv9Fk2SyesnPQ0wgDuglVEtLPuLL50Mzajh
09SOuTyKxzrFBoVRByMXF2pkbBSYBYbLW5kyEtVgDRyXtamEcvGsSJWd3V2eSQtMAw3NFfxNpfT8
6ydXGVSaXProq/kPjg3ruux1py3L/yxgxvs5HVuyRYVlmtj4Ts16/DXwnAnktsAmlFyJf4t6ZGFF
yulYOFiiYqNmpvnAbZTeGDHdcv2Mb+q/CFErEWaZXh8aa100qEqlBY72v9sh5yH/TjR7Fxvdjyyy
I/E/H3viImi6mi8QPh+vPE5Wr9GFkrf12fyRl80oHPPzmNmQ+CqrNXmNn7yEbXkB0flkVxG+gNXJ
NuiQqHvmGpxBlygT1B+nU8zbSP+X8pW8cW4bVKuorqw3//l0KqCbvKrmF2KHffcwtt5DMA9fen4H
YbiBNtsXBKMTHsv8bnrdHQOacL/66BC5QS7QC1zdRgKaczkSpZw+0LyLVPvhWoQ/Zt4FkOqRITfn
TvriYHEMCWOJb4W/h4rwrE/V0DtkwPCOHpuPXfarTy7hyOW+FAYqrwxGpY3nJ2rcllt9ZV+XnJxn
rdIuCznubS5/0Y0hZ8GpxiEeGfTBaIYtqobmYjEb5zzuwCtS3uGsEfMd1a8OdVilXVDkcpTs2WNc
EH5481tmIoabs1M7ZYWWR6AUR84PPnyoBQpUj2k9zwGbbBWUs5m8o7VHQFhupQzagCQVId+YXy93
uh9kaTnDFxF5awFoRV6qa0VkUSzRNNphqwXcGSGpey3P3RwC1yNlds9wiH7l1Nsle0O95lIPIMQo
v/2ytnjmGVpG22r+yPGKIyMFrbxNEQMNW4j3aYiz2ZbFoJD9GnIStuDKcxExHgIEdTHd8EsRGL4n
mfK9Xi4uL/ph3CczsW449rv1pu+YaZIGKwGbPxuMaMa9YHkKUF+iDIP3PetuH1hxb0NKHtbhhxLf
2ULWx6v5KA/Ua4/Ds9WqAEPEAyJB3Dt0EktV0OP7tM4Tr41hd04K7lOQJeoUslwJL5GfzVBJ2OCV
lHMacK0hMYdDkjh+yoMo1tgccyTyChnvllG6+ogWcE4RGTpx6W0hFt+kUu86Xe4p/5ePPgOJ1kw4
jeZNC7ieDbQc9OrjQRjNcq8kyLy2qGj+Rv4yRkwNEaRU77M3hQ5z5iLOqmlDb3rQehpJp6Qz0IX/
XsyLdYTaOruC6176WQHK+sK6Pe6gaVy3Ndr/6r2wPXGNDEY9DIcCm1Dos92KizkAF4wr80sjOeAc
VcvCA7W91ec7aPDXxgED758sBEqRkXM+OuMOuV45dOXqS9fpg0fe70/yHw+t9YKt9442PD2Ip3Fa
GmGO/KJovihpFErKABv3Qi7YQIkuP5Xoh6WJulGbZs/k/PUBfjQWdnZsR2Sn3+uI4DwUGKUFIbYo
1BMXFQCmyXnJhIyxKvQvF/5PO5IunrZVQMbxPvdDDxEsZuV9qJ2DL0kiu1fS6JBenL5Vrf88k/JA
kQTFZ40p8xf7PSAkfK47J35Fg0YtG8z/+6uL3ClcvNqLttu4fOEGd8CP9rxSSBCGrdWDwLEQ2GK2
jUz0a2Ng8n+Ev5uFOIehXLQk+vuozd+5i/468v9NIz42oozfMl9G9tsozNxINpRdpkIxmzC3xMzV
5sbVt0cRGcEBkK3ErgDFd1kvLNLod0ysOdAEvuhz33BD/WF0ZTQk7+UfG9Xym1D/Wcl0Ofazf83s
51Sbzu2yLUWCA0vHBlquqrLIB3kW+kIUYjsoWjZ0s2aqP2lHRxa+BRdfDQK/7ejp2cvXiWBJEOPq
keLGr9RNXkxXp8tVui1R/Q+Earh6TylcRROwhpjyzV9bt7XWj3XEVB/+IfO/WYw5jnjpvXKPZr5h
yuBI6GM1d9m3KmFVQApaLObpEinXHzPRI+rR+q+E9wRrEK1liPR4tHneldnNEYI7Tbyqsoi13kWl
R52xkj0iYu9VVd1cceSvREPDLb7+yxTzBqqrnNUMH0B+ygqtNY5twUFx6dQVmMYxoMIW8OQKIa1p
7QVbbA/nKTWNWUrVG312N+CaAE0Kr0XQgVIJFNuK0YEC+96Xn38+/VQ2EA/Ck/iI0FPK94Hc4Rlv
+mnVVcqNepgRUcUQDRwRtPQYZcRY/IKWVJIdkzfgk57IQWlAzqyVuWgwlVZG/l6OOR51dJpw1EL7
9wIun+inGdMbsWOF77er53SUgreh39ApUE0wQuppWwvS5ZXgh5j3hNnW21CWh48c0EWtGRWQyAht
kUpcKmz0N5ad/WV7TNwAm0HzSMI9td4D3soHWI9YRHJ2Umd+zHEaSVEfXsRSlIucagQmWlP35nGM
gIprbCRqq7cvMPuoyg5+plj6SesjF2eUhvc3xp8uD7G4WH5bnjD/PLcE4SvLubv8n/wV9Ck1zsgE
mIjRnTC+lSwMK1zaz1XUzxfv8bMhoq7E5KUc7XRqZGEcKmSdHJ3q/70UHeM52Uk8y3b/3muf5Qso
uITKTysRT/TUqImg68PhabFHwRuMaMjS/lHBR94MS15JyRl8YxvBNTiPHu6cmqSDml1wkScMu5+A
GK2+oW9o9j4qLXd/q3j+o3lzclrS93SJBcP9TxzZPyJYIavoMCS/qjO/vKowiL08NeALHiKLXkPa
GIPJyM+dbsf8rkArXnJ8DAjiflPMYVshz0GnNu+aMdw3Uyohw4S9joF3Rtnv35GtbpfLLA8i5KcD
GriH8Hw6l6lss9ssNkRcwjXXdyRjWotsoX1ONBZ+30aW3S/So3JdtSH86YY4nxb0+uJyPF+AdC0N
lUyl6KrSXb9s4KTr/uRj4/n9lTboFtu7j3NVNYU3RwfwQGTtP8BjnC9PwAEo2UeB7lqr5ZVytXYE
blMrPvGQZuqD/y0YBEbWpCXmcq7PIJOAPgXpsDGBJKDoMCcv9n9gW8zBk5P2j2b9k5SngdCjj1K7
WJivkna8v8V5XQ6FG+TqBB4pRT5VV8WU+7qQCHUJ3OIwZpaQHaUSP4bQEANiyT3ueo2aqQzpNmwA
WTHqBsQCUyRYXd9m9gOoc+qMmC4ldJRmOp45nlibJccms4Itf+hMyhmSYTRjdPytzX2t40TflJRz
bXHeB4doUo6NhlFuz3FR93qhcRfrHJMYZR1TJOVVmhGDFTI03NUtoWKmwph5TTcTgx+Sbb2JIlb2
ArOcmEGCpJnKNn5VwwfM2JWyHRutxj56EsUTL6qr1H1eBsuCWoDve50awHu+AhQHujNJyuyvT848
yuHgJ4TLfvEtX+xobPLjeA31Zl0EAIkbR3/ex0E7NRwy5LKiVEJvhm0Op9F4UqGvHqC+x620+2Kx
vL0Qc2OZc9x0xyBqCGag5R0leStVolE0lUGrI75rCC8I8jXdJQCyGnL0dLyRDCNP7AEGL1MsAAfn
/geWd9tqxyNLTY4PhlU3BI/XAIBsY9jVfRSs73ZPZTNKlOb6Lz0s0UaHiAymNYKapTtTqJ908mhC
FnLzuPY6MXnI289+WHstpjE6i/+eB48NZKti+WkCqL0WA9LoHYwyT58M/IR220qe69cLuQGOHv/l
H8k31ReUTCLqv+aeeYHnlXXy19gjlXe5AskXJyRiUakAFQuCYezVYZ53El9UEZOfY3V0VF5ZP0vb
SdTmsvrBE9wYPvDzwZGAnetyzGwPjQH+zLSUlpXZJqLr39yUo/XXf7Kyn9IgpMx3dIgD1FtiQDE3
tNPShQpydBeGc78qPrb3Q5TLvS7O2pLwyp0MKhuq9JTP4mdNpU4d+HKuNVhxnw+PJEAmEVgW1OCN
B+b+oPik6VedTbOO77WvPg3nSQyGErFFQtRB7C3Dp8klE1eKGzqRe7ES0Rj1+jSbSnxHaU/Fiv2d
gSevDoks1+UTujIxHxAjyFEq7RLZBYs1LZP4KMCn8+1tBech/cvCvz3noEQmMmS9DMIjJifqE8fg
Ft4zNbrF9/KUt4MFk8UhM0eEvLsJn8e1YT6aEAdKzEmyXNpiIalgoMIpY9/0jXZcg6gXS+P6OetN
7lzlPumLWId1ZdeZF/cz4IxgluRx1QLpayfu4hA8t8D2JRCoUGAtBCKFbSw00Je/lM6bp2CNlnxM
vWmdIiKQXwn5GUl9gKMULUZN+84w4Z/B6Ci+R8sGsTsa9J5bSjeToQ0Vjd/hDVAMz1NVFyNxuN+v
wwegRgDkDwxb0MfT9iJqokhZ2XMRmEfdbbjZke/L7zsDcd2jKA7U6A/5Shqrk3wYl4b7+agUF/4P
Cte+NxqWDBem9q41XjNt6aTOq4irNnn1U2BSAjzJs3z2zAeR1tTcd26XxZj2YLt/cE7za1l6BLG6
PIdde4XUtRutdahHtzwWAIhYUMqUXDe78ftUEvVcXrrmWLEVekzJFih++REjCosLq75LsNSCS6TS
t09lBG8pqUZXxRuWeNXjxDWEVDKUzqHoVHtQstQTb+CjZanXXcee/RCjGBAHsBpKyhCeXluES18u
0Q0X7V1YIrsdVbRDzizom46eI6aoErro6ZvadKJFYuzi1YGCOt2XGh+HiP7soP5lm7Izr7y1xuo4
SAFJ4D4/OTMXEG678/sVBOrXyiRha9RBsiaVJsYyhPV+AkbelMSXuq+XEQK9I/LvUgb66t8aMk7e
BnG0fzLSzf1Y80m2i1+R68VulCtTQjpK061ZgNq01ondX9So1tEtoeim71TQSumsOeH3LSNdy5y7
hH24JTc4n3C0gH42Jsewv4SA/ouEF1i6qcy2/fx//Q3A0B1NO2p/tUy+c5Gx9kv9HRKp4fq+ICZy
W/3uGUJqmtscZPB2HcVjgmQ8tvfmq5+uqHvny39V5xdk8SpTkbvx4+03c3B14h53qWCytFtgALwO
B3JHrjXOqieDqIXRidYMtuKb3wftp79OGgcm0We0GA/CLhzQMP0y7YqASS1FHUGOPpZrm+Y+b63V
+cVBhUwthtXLjSI+27srFW19lXzYOYqwOuJcH/xgiFfVu2mQN+syzhKOPr3Yt6bfqpwLrevgUTiQ
p6p1dJ7+2AxXATWQRR2kpq0edoh8PBjJ2N8Z4nsYRgIumaKWEtz0YGdsUhXV+FY5hEAaE3oAONBC
uk9pVWM54YCvCop8DS1lt+qtPo110O99z6qxVmD76lq8DW0xro/z/u869nG1LuMItDMVzkM0kcfN
EbTr4rf+PL3vVLH/FjFFU46MIp/WDDXK9z7jSOxI7PBRBAVQqJK8VDuY8BwC6COw7Nv7ENQo7ock
jpM2kWjXXEcwm21XKlh622S7p2yWvM9Nzg4arhcuw4UM2shEqTOgk51s38cUv56AFlOo3ERtJU3y
NXsTNTSAhYbzQp4fyAqhB0ansQtcf9YRXmn1aoei9cN7PmSMSupdTlXeU5jdeNyIpo4EBLcAbKY/
VqoBMDUUSf6l5u7OveWXJX3/6STAuo35L/xIZltbjrnvooBhGms0BhlMouruGqYjclaS5eFxS15F
jO+Bv3fXxWO4790KUc8aztFdP5L0ye+b+2C9SxNJKE/MrAWruyykhw92SWigvc/Z4VfZ2FMeVOQU
sNB18WTPxwvHv2XLQl6havoGkxuhjgSISLtujnBnXG08Wa87EL/aEH52qmcdcIr9ToTx7rgDJuAu
kaNsgBOz8o2XXn4s3zuB5b4jSrSHunFzmfj752T80eH7sKyrQ4yZPju1SqjKcvBwEevKb32tKbAM
zZ14mgJ1P4WrW69f9XxCFsPkEovlYemxcSfS2weD4vqONu0FXwErxuiNTPFGLzKCRC1tod2y2VGQ
sGEI/EKraNUt39KZFSAjWlnuzLLaeUsTD+hJMe8QxHGUy5EvnaqTxkT6XHAKJLs59bJToYJIMljo
EKfKP3cIdEJbtUr+t+8+A/wzhSMuMK8sMGJ+VJlBPSn0jg5Jj0Soa2XjRtjg9Of3aRn26nRFdA7F
YRG0oVHtSIeXX0q5NhP7q2VO/kNMqZopOCgPjTuzjsAJ7+W+Ptz/6bRhI3FlWqG8vlHfY0gojKJ1
FpxW5MH3ncBabe6fO83QmeOycniyrKuTEjRrbCMs9FBaKNXjXwjfO4AHNB+bqKwkUF3iA9hY6FMj
LCTBfqjbLEkPbfNFkq+I7YA76eZj1uzzeiJ9plKqHrGJ3s8daBAnVEsg1flZh4h43AAb/UI4uwN/
mv4cM3GGfS5nzOJG4mLtCA0P0s/SFyXtGzc86RR8OgmMwQeBrm7HRKBnIAOGaQ2zIDmzNcx2aG0c
I+yUti7LZiC2lsK5/VXN8g6/x6XMgNKjGFLLLWCQXpIXK1h2niI+7yZrn0Pdz+Ds+ibaF/KhizHP
4qNw6iywDWhxbcHISOzUQA3WyK3uh8Nq2APaToUROJ6FzlwF0f1Yat2Ba39fKhrhBXZtXyRnHgIg
QElxMNSnnEC3Rxv2dm9tQgxt68WMCWUUdp/rBb6F3HVuqYIiyEjnAgwZ1ZWTKlx8wbhfn0r58BUY
DyWmLQdajvVOxebhiXT+wM99KiL1DQlm7bvDa1MKb/Nkws4F8eBgq6VNNBuJxN/96X/MNArfDPag
2ZsaI4MqEh9olzw8EDZiBY7LWC6hp5QE+oXlSL/Ki40ZA7PMxNgeOnyfs/flX8qsHfUp7br3hWz8
55t8ppA2pBDW1TUvnbKX5giSOHrjpRVa2vKlw+sKSRW6HRcW+HdenSklKug9GBwzvs2mHPFpYUgl
amHUBS8PNl5yHJ7C9cTXQK9Qb9lxKmE8tjLHAuduXf9FzChVp6/VBilYHKuTX6Ug1kV/rlX1WuNW
N2zjIpY1ImtNR7x5VcSolbRbZqiypn/jCJz7l8KNQGOJ7dxCcEcW04Pk4M6nsxNZeedjA+oR2s7k
y6ArSgzfcf6h+ZPH24aqimfOkrarya5WkjCuz2vPNBLEmkKLEzCRYL4ui0+iAVyMtVssonf3M8MK
Ny2wPxfQYJJCZbA/jnffORSnMNAtE3yszyFbxq7bthewn/N/rUaXmQSOpihL/+u0Ww+KDE5C4Lvs
K5Tn+CBSHtiP0IKSn/P7lBJki4VCuNCEFX0xpjA72Fce5guPXOhIjqkpX22/WWmLPuAy3c6TrGzV
zuJAQljP5dCNCLunRh+hjyU5dYBIV6slkEwRPUIIiik6vlYrmpN3IXvHoak+Fp8oIFFvKtmaSdEm
Bad5SYxHMsLn1Kbc5cTe5CMzRbOonsjxiL8IEEa3wudOGzl3XJ4Y9ZJafU5mYsvk7z3i3xO9iMkw
qeb4UwHBLjWNMT8rnFKiJHlyhdd05sSDv8srVa/n3a88WSUZul3+MJHyTjWhSu2ZaxR/TJL/YiZJ
fcxwhMqvd1B7PIPlLp64IZ77xFieHqtX9wAPIMo9bBv7oPHwd+UTSRO/hyqSC81JR2krnQMF65z7
Egy1jyVy+BOfTZbUd6Qnf9D3/oZLyFxavZDaHSTu4JkbaOQAeaJ8JCpdaKjsY5iAA7/993+koSwZ
UDDNPSndyb51OW6t9J4pOCVlLwVIbvysjpKrObdRepIP2Ho8SYNZxE95cTPzLcQIjCtsaktstjBI
X8Wt+5UtJGDlvnd11lG+cc25smWigZ1nadWLx5dGTtQoamZGZwUODocee+kErfzME/OmJ7AYg1Ff
jI0I0+HqTGpeSDxdHShJEzD0IoeSm+VczB5MTTkDV1zNmNOGdZ+GwATYO6e/W1XGU3nRfxAikfuo
qa6ZvNPWWYdTDRsQ4qCMvXkxYZ63uK1tTzfqed4bnVeMg4IJ8vE9vUpxGZdrDd/Kmjbpj8RXY/9z
girsVCTux/D6FlfFSu/yIKMl7J5FhFmYjtVSVWDntPCfZEozN4zYdF0yj4p7W+VgRf7k1inqFnxz
Y2PHVvg3SO9Ilh/mSKPu5ITg1ixPb7a9F3yKsOVJFPvz4td4SGLMHpOCmPRIbzAUqrg/lMYnDrjH
2HB0u5Y4wsLVuc63l1FLQA/5xIHTk2dj1T7Cac31sXuPh8YJTamoldAmajv5Awbxc8Bp5UoRA+aA
22nNJaQUICo5z+TjZQ3Zjv1RoJoVktJRLZu0O4DThmvKSHLYKuERgVpCnd/rBuwuCdm49iL1jLOh
JA5DQ4qUejU8yhD2noI58vq2e6XtvkufKCcwlOI2Ve705hznDla6SxkVmyzaXQqus+eaYj1ORFdf
fbCKu0gtDtRrxgw3E6vNfnilD3T4aU/ly70PYy6saGcVuPNGOcRfS9UEwHfKyF38fshuzs5W1uXp
KfcYr/BD5s7L3B+BJtViMzBRpSevn0r4QE70jTz6LL0wWtu5wgUg4Qcb/9PZD6S88Ox1GmgyNf4m
qKqrSi5pCjC3hhEUV3Dp/MUTfr1/feIXUSZHpJa0NCzHJ4gjV/cnOFjVSM41+UH0NeC3Lh+bybq4
E3CmE92GJCKp8GeqVVVkBvIdLbB4Bee2i/Dn4QDG+9rUtL+gmsEqk4qLo6yF9pjMe9Jz+RO5xFIr
D7vjVcr0qNNFiVGnZ1Kpt3NfGiNt5sKjrAX9Ya9vRcaPqn4Hi5eq2ddg9O1/a6ugrjZNRj3ejBXO
tK1JXOLDTmB+pRW/ftqGYJsl2tVtRwnVNjCIAtDWDI7G7Hlt+7+j8f5JRu4pjOUky2hFO+0dQjM4
vY+q5NpNAZ3XAWAXDv1O2E0H3D7mohIZiNz1cS+cBxSK7Y1MOtyNvDf/AHH8ZUzEimsRKEdGzZOi
cPMIciHQ7NpZnrXgwQGE3EdnNdCJXZ+PlhBVS6/ur4F4mfkoTf0dGpVXNMIf5O/v43Jq7p4mxN3z
qO0UArWIlrZlz0l6nJQoBMMgJP3EZvWI9JbZaVlQeGt1QXfD+k30y4yChycyScwMNSPM/Bu1OIx4
BjomlFMpesWHMM6bpdu77v/gshS/wSS9vBVhKRMLdy7YxdvXCMIjjvkwhDmLaKHTeu1FDbTWpdD/
NEQMUltuOiRWZlzBDqkQ+AGp8EdJnCoGpZeh5ZMKjMp4AgwCNU5TjBobjUjFI206Uve1Dn3LYLSj
E3BpjizVU63srsFAXoY+OdVmnB8qhanlQENj4OBnPkyERjYuu27irNkY6UbyivZe+zhx3zxzfAAY
YdtuAZBEU3OFaxjq4ggCROhdSV/3zdplblP9+w04ipl9Opecun0KbvU4IHk9jUjHjBoM5vyOz+Bc
SHYnVQXVP4f4Tlj3enDsA9CB1h+wq0AyLK31rOrMFUFhiS49JqkXFzYcoXsBJ03Dh/T5lndMkMNe
d3IUTD0drmq09hgoWidx/P2kwfkNjXsoNBBovSClmq6ZXPAl+38uSxmw500iQNiax80R2pMB2uqG
UiQ5d24OchPIRIVnKPOiRZsagxEj5JQBlbiNkMChFVh8yidUwsCepadvp0qZk3QFwH6iSpNINxTV
PahyxG/fGIuQJ6+DRAI6kySHRoQ0B7hcMQepTb/NXdtLKM17zExBgp8UVCelqUVBh5s5nFfhwNxz
vd3uWcXcZQEGC7a7eXayGWqcweOGysAF1j3F/bPPf156/3R3remCCrHdX6HLCsu3fYCV+rUOEkpi
wggERintSxsWPg6rmvDQJmyIXdYrA2eE4wyUdx6V+5252+z83INd0TP8tJRQa+H7Hy51GvyKiycK
b5mAMpLokUYmSBDAkFdVU61VlRnOHz0bKllye7WDlo7AovAwfGNA2BgQ2gufdrIHnRzNaWkTQpYZ
uIN+pv5d0Ba0PLW0LuNYVZbfETYh3hMM9LmhAQxUzwBJt78K5yNkIrk2npzgI37e9VGxPDhZjPtQ
IJNHxDQMcSvL6VnWQNmMBDc/15FaT6gXPejkI8Y2fKrrygavt9ysThaPOTT1tB7bgwlqsXkdOU8V
GpXFnGqEyNtkWxzvmXI7xjvUMNYFEVl/uwhGYmYzw9vr8xqEQHcl76oU0gbd9kaWnw1FPqhszAYz
CQobisZrifZEth+3+7StMIJKtAENlanhAf8tMXU7xmF1JtWmAgN9p58/2QSSn1h/absZl3tfc69O
RddIIvlmQz9sTkT3Ci/fT+3x0QLW6DxmRffBN5BZCVEZgSbr8GFtWdI7dp9mNkLaWWbwnHax06Gg
X3nERS12GWvzE/G+HUdUQc+mqRqbonDJA4bG6+i4xgD2TGb705lPF0ZEYZC4PCGMYQ0FkQ01Shbg
iT0XfcFydhe3u9wBtAvN5mMyAKU3H72p8c5+4XRYJI1LHy934vaeBbDl+0oU6Q4959JJZaP4DaSI
BOVmV63onFtxMWpNBtPueumB3DrzCbEqwUgLf33XdLtJKljHx8g/XUnvzJ2VWBo43aPhiHejPCjW
xaDq28CZjdarC2UI9cNIphVLC1Dt89H22Yzuc9WISyrCBDL6Ut9+vkeqCAAJn0jDGqud267q2RSV
sPPtjf6Dgk+WHCoRdzxBO1l63NGE/ZB74xq1C/tS1fp02GYpr5O3Bt9CnGEVhA5wxtuf4tnwrZND
okiksdlhLTs5NauvWlLWnFmCM/jHuCxGWyJuoW4snT/kvqRfq9O2yilpjwB0iKL44BJuRbluXakx
BfTF4tVH3TLgV28w6UmPRIb6C4GiFzk7PTgOCKH27H4HOukZqXoQgG9QIsc4UYucWdeDY36iFVRo
9ICVmjKBdDW2gGgZKMiUz/1WYzz3g3IQbCV+pL3Qz2KEr9Cz8x3J8J9FujVLD9Fv0kaAGOyEbsan
ClU10c2t9wGUbZPxB5y1kIfP2TU6UlQ/oL/1Ml1zkhgDvQy4+guG8shsv5/RlfF/920W8FwERYIS
0c2jcFEJOO0yacSuwfGtguPd2iCBsLDGEqa95tdkEwLb9YACnaZyNY75Byo/Ed3HIm0Wu6eFd8DL
yZUAe5Ryg4AVGr8/TC3Jrjaad2TYT+yQVyW9VySR63TYmWjEJVC5Z6JSrnYaWX4IvT6qQ3tAGRvP
USo8zzumJ3uj0AX+oiYoQtpjpk2h5BVmpm7bwTPUJIEhN9MNTtALotuerAg6CsOjbiSNzGUX4RkH
gFbzgRYCGZMtzRwUiksxZ9qwFNuXwn0YxR4sr5yEcWnC1VVBzc9b3f1alqTOSldfzByT0UwOhRKY
Oy/yR0Aq4Qv9Qx62A9m7KITFE4wu6/Dm7J/w67ZXm86l1exkDsXqMFMEHJv3CjYtQ/Cpguk5WEkW
fIPmb2H1OX63V3khyPhLvCPgRxSGGtcDhwsDskSuZuCwP9HDMWGjSLZLMnqbgejYiPKZ8GQ03C/+
a1fzHcRY2QnnqN55TCsc8nnzpEYJ8rPJ18W5X5yAhjKLzFLH9T/iUF0RhOhAz5+rq/jLcU3V3H5C
fpVsNoSbYQw9j6r4NAPTQK5TCVomfRzUy7l/09q0bXamrWQRj1Y2dFe7M9rJATbWq/Og7bvLIBbi
cWJaRQ+yIxcP1stWAatJGlMog1ZkPz9iJyN3xwkHOtxPDhpNc7FqY+IjbsAC+hcKZdPAs/PNW3ab
dwPpAO9qE8amHSxoDuY3Gxetx0Le7MLVWZjFdAzD9k1IPc4ROurupqbwq1l9gsuyAfAcI2wTMhe6
4r4LBlucG/Dzzpt3H67mGs9vxXd6pSAhEL/IoS28rvnrT0jsq+1IjOceA7eUv1FlZyv39dtfJveR
DtKIp/x92e6hTQ8wv0WKBugJtUSWvNgQwb/TJjdu79/mk8HFeCRk2sjQ2laRk7kSzF1FPKHKFx5Z
85zo+YJp1zMNR4x9hhFVQT3ufJWUR6SHWbApXTJ7LDkFjGud3Ap86ljCK72Ei6Stn7t8EcJHRR6d
YKndgvdms03N5cDb7/x6jE7IeRNpjFuid4boFT4NVlkvFq2Sdjfh8nEAvWERtva5dwljzHhHJmqf
FI9rfowH29j6NgrHU6xYKe6kNUGY50RtYYLvU9zdSiwiR3jUzFm3e7p1xJ+2GXvRlOyyMu2nUSwE
u2xWoeE9dTyFoixGI0kS6SAipYqESF3E8hbIEz2mdnh273GuxDBzmcBpyP+UaNuXMgrklm9OXfDY
RMDuSag6+HMYwSVoSciy3iUzHkcbOo2Lg7O25TFdzopKdLdRbPmTRUH9DhqdjuQhl7brW6xRMrmm
bWQmqFzC3lsh1Ej2Y7bN7vKE2Nsl+7uKuufYDX2hh/Ut57BWQzmPVXsS7OZ1d5Ueg4z9V+DVmTwd
EYxH/W+IMqu/KQ8UgQ4D8a5UJ4mB7GfMbGngwJiD8vjIoCoSkiOpEXGFd96/A0bXNTmgjirFmKKs
abr88GNYHxEJLFcqcC5cMVtiW6Bu/BPmm4ZZWeZOcl88PP6jBNJmgIGn1kKhaHUI4WFs0968KRZ+
YIbEt/KfnDUWXzbFLPxoBeRkd0ae5BNw1JCWzduAjqcTPcIZXR4h5rdpK3dX4gTEvRlo9pBMoSkl
Ls8GVsUBK9lREFEJBGLF9+I4nP8R94nOJsoGrkJ7vz4x7xD3mHvKvEgxPpKUqB8pPLjJBCfYES5O
fQy8VMcYfrM5nz1xhY55/ahvu4PzTW5VDw1rtXME9VZpGC1oTlaY9R8FYsy1WSPVU8qg8iBXeph0
hLgw7o9HSZpHOrsRftmdm61KR1JYL4aB/buM7upjamDygG+2nXzyd+avgrMgPM4u1ufasHVRpENl
dbRa7YQwtHlZZuWQNbcsA5nOSqY+w1x5tDNYA/cPVpK5CnA1hoYIj/X8WZcpNF/D+da1+huRFP3l
9lIVvHdqsqwi20iuV4OyFViVxFWmpeLrkCCJpRR4TY2cG0l/af3Zvc2r/ul0TI7JC7hQ9JondLc7
HH7FsyIlsSfC7oA57wgiiEKh7DHjW2M0Da6mCmVY9qzsKBiRUWIboMiVTAln2Lr5xoj1DwPERlCV
odFyZ1f8cqLfjFZoO8NMC/NfY2xBW7pygkepoFlaW7s6dE/oXcfZmfx1LuFM68k+RXKItB0cnGrb
TOgbHFa/qLSCp/sIjf1zuei533I/JrLmzt4b//ax0EvF9FX1xhmJC+Smu48N+smnG+vCRQpgxAtV
yrLWnTycRdqDyEW4hORgRDRvuCHXWDFeFBUQhZM4nm9vskILmD+NiQCDqZTft71AtC+F924hysLk
ZVC8AyB4UCK040HlLPWJx3hM4W6KpNfjYucMSp4Gv01WLdhDFXPE2Q1W7eL8yhM/A13Zi+v+Ftxg
O/ntapkw/zctahpqBhH0/1Ic3tFCpWbTGOUFPVhz1ySwFnVLNsI8pHrSvBR+jWWH73lELFRmMh0m
E6vu6MXZC2VN6kGKLRjBHkIUrmNzWf8AwlaStC2Kim5nm442ZS7NfDzJKoZ2TCbeDDf8CIwHjJ72
h0ZxCU9MBnBMPwhFrUwWO0Gh9Vz9+bndyCB9IaiKu55vaFzRJfX1N2wkVZBRf+b+AH9kaHARZzMP
MKmaWZZJv5c2G814C9N7hbP1bPSQrQxElgUUL+D78dlfx0kugdh2vM1WCSoGUMfsJMXpI+NiKeQR
Tb4FNApKOaBgQZWVe8rEhX3+jGTF45ijtYirCaknB9Tk+ISZSNLXNSi3uLx4Z/84imOgpUXsLHEk
FDsL8kY02LPP/G6hSRCJCIaYbAh5ztXt7lCIWMBDnpnNQjjrshwyk92cWuA75QCUk1dYSO6gDkJF
8r4f699tXx063Z97t3WkYYMEmgY1+a0Me9rHtBYP0lwp/YUHrDYLzz9bFoTHBmLTT6X/lJz2hmFc
8r1JdwsVn5yW42AtQaIOWUjt1YDOBxNntkOJBKldx1HNv63icoNFjoLR0r1v5CwyyqEf969P/n0A
v8lkaeU/1VJutkvYk3FSQ/pOPotyX4IrfHRpEJAL3m+uoNSjASwqpfDLj0plxNVk4oRRddsbUw9g
+JDfzcW+uuG4862on8LGEKwg9cxRKKuvo2YKAD3hLlgDpK+es78QARwUSfa1EvJ/gmK+q/MuGzL6
O6nWTqy92esSFH5mBYIkOVcekJUpWE/ts18xPgG2dfpK9aWAoSSSRVwS8x6NfnkWeIwh8AlUlRTa
WjH26rGfT5omogUF0rfmX8C/LxfZcf/tzksCbVFBMKeFcbqtkLGDGVbHruTZJplgJrk1Mkv14cO8
nQKdR35ofRM8T+hsN70vn/CHS/V8V2+MMKsQcrsxomEzVzB3d5ts8ojr6+6RuaJMIjFsA1VXdllT
F30xLPDdijkXphqkena2LIzJ+2Ab4Qcdbfy5IZTITmG4LhVxs3GHJ7O5a5ZRRkWDvjGZf8Gd6xDF
nUdmE+sBIo217KGGMKLMLux21RCZ0Dt2Dj0lDw2V4qLJMPskBiRbAY2L9ngoA1jMjaY+OgIPlE4k
r8+lxeZ8uDH2FcEwd9mfqcdS0kzIznIM24Q88AEk035sbUMF07uU5B3jt2xm4plSiDMCG5Aw2NB8
6gQ8emjOnO8u/pcnxymqvm0a96ixmJl4ZXRAr+K2XTgVQFhH4BfhQrA7PCf+S6J3KpgUiCj1ezsH
/Wn/1GRhWtLjypOww/ldsKAa1fdnSXw/UvvRkVoA/a7iSfggdXuuR2vHlR47hSFMxioWpDCcp0yp
xSFV7Pib21LGpDPhcPyAGTorfnOjACZzP/I5RcpU9QZzJWEzYVapSxtFiL684K6Bs+hoCE+CJIZD
hBr0snDNxIiBFxOsvN4zl+LeBMD7UxMDbJSxVWRGRBc3USkbHAy09KZUJZwQp+fs+/Yw87HSdgHc
3vABuAQmaW/1DIWsZaE2hEdVvhd/yG4ildcGhZYWr2xMT1zJlBOmRpM//vWZ9LJpzWaukuvV4ZZM
vzneTiqjwfnEn6iz+Jk9ohQYw3Hu4nXxwLnGQwUgRp21zGvktILraS/4KKE27BMCQqkck4Mqbzix
h56sm/Eaq7hOP1cF2ZIh+dhmyyBYu5u6ws5WClWjdblJIgR/T1sowW2/f0DrzKGqV7IiTHpg4TxJ
sMXKsEQXOkKZb5eWu8ntWNptCyVuWNLf9hDo3OgDrH6+7gSGmxvBBX5CEFpE2Y2mOqdO5spZzm7U
UrXNh+t5m5vHsvpb1nnh/NxWJYwkFMGKJDjWHFZ5uR/BpSn3dFPdmezsVo2TzrXtBMpcHNfcA803
L9ul4iBemv4Gccut+qOe/VtBRt4itDfotFSgvVS1Xlc2q0VKeJVijUQ0U7hUe0a48UUsgR9DjarY
8Q4R/hNrEG5HayPJmSVCppF4MhbwqCwjzHqrYdblZaqI5cnK1YP/+BEsULyM9gaYpbBPYpqo6ZRZ
A6Is3IdL98dyJI5ir/8xl9++c70Wogc0N6Owm50HbNccUpYyxwpB23eCqXKpI4IoQgVsXmanN57w
rt8DLtLuQ6T89LT1NQnrdkRwrT2FhwWv5VjdhzfKLKX+AUrTs+MgiVMb+AlreRFvHrztTXIRoNmG
qA3jQQs4g7l3GRzWQksktZ/nROfDgj1kDFu4dSPl7qz6t8Hg5mPRPZzhGuyI0t48L1g2pfnw9SjD
hmiuxVDU9ziQmOTN8k6bw2mJF/zd1MWTDS5FjppVV7j3mBZ6YTHFCfNHDZWMKBir9v6Z3scvK1TA
FDveOaVeqM/E8uFsyV0wgysiaesdHe2qEk3sZXPnM7q1eEIv7VkPYPoH31LBrqICNZCO7Qg4RFk1
HJ2nz5ewGlhAvw0+fDfo/CFXO6ps/5XNumi9beycwCpd6PPGRGxf/TJSp8d0QNnpU3/Ma2440bki
0B9pzd7vF8i49bBIeytHvwb81MzSV36RUOhLTfqu69LIatHqE4cEP1IIlE3Sy8vjK+Pu3qqclEko
DSIRPKxGvVOJz8t1n/W9fJZtckrhxPM+nBvByLbi9Zdd6C3fSbmdW0ZkL82J8G/vNaFFrikR7MHT
XbVfA52zuCO/qIPEC4kDL/gC2+t+MCoAafvIyDxuwEDU7uT0XmFWR5r5VJqUo8v1inktq0nfnth/
XiZtSvJd1TrHnUxbkQyfkjB/wU3uyb92QATyWa5nuQauzV/Uv91FVp2Kfk9hRU/idWBD0G3XgWMq
/qUJyDcXDteNaGYioS2KmHdhbD1KYbaFqyd2Kcv/fLKMWygKwAILulM6ZXfxTGiGx9e4/giTlsXd
cLs5GOn+/L9jGKWfuFCwDjKSXwCTclw6ek9PSUqr2WTjDz7hyOK0BAAKBodw0iwXaNuxu4mMDWpo
8RqJhx/I1FPYVZX7vlnOkvLqPn0Or5MftwaInrCkUZIIaee3PS9H2Iam2NuS8IDH8peOuZx7oZLE
6nS3X4A9ImnVLH/58LtOjhcYjNOeSQjTKKyLzMvutobmufCUs4vQBBF6zMo9PRWecaTExj9n5/BN
xbAjRXlyNY5AEz3I6OEwHD3iaRyKMo6FGqAzlTwH/i4MkdzzNbPrULjMyqMyxn94f3+rcOiYDQ0y
O3oRuHTC3+fkYomDkgBx3v0qg5pE5BDqhSKIjSq6Dm2U4hpYMDTYYCv+hU002e6fLjmMNT/Is0rJ
5xrsyQRCT0LnssJyG6utwxB6wf8VLr54TWHU+SS4HE3LSFi7gFKhEQUBTxR9VeegmhNpF0M5jFz3
DQIhBDSrKmjO7IH9dl9ukeZIg3nFiC1mzfg9hA7Tv5M5ThO1TgewjmNWsRSn83tbclbZaUcrT+U0
zvrYFTx8RU3+4U2gcz5HVVPy0J+n40qOoObixyIl2LSE7JnrZ3sZfMvxhqb3pCMGaUr1AXxKfm+A
/mfDUXmgSAEBM5pkQtgqjkHx3lT5w3uceoKhu9iQhECuUzgiC1All+FqUDr71QSxV2wln21fslRE
emjpfMDau9u85NMnMTym26ujk1ArlD1z3XAYssRsfqdg9QZ8zKLR8ny5aTTiyhkobb9wGMci3/Hr
irWSqH/+MVexb6i1MA5wnI3Miov7scyx7VAKW5Zk2UIsLSrxG0rFgEfDAId6x2GzIs94zeB31f4n
C0WKYW6QnG7Q548UM6z+FfcK1pCOwMbIT14JimdoajsrpEbSOSZOjaj+x3lisTXpDe++cOKSACtX
2hzrE6cNc4DRLOZx+XjPsr2EoSXs7kFyUK+oLUwZkuHmK/OaEAoOD4XupAachPo5lk3oIgHyPt2j
QIntdTFBp02Ua7C8hQv5Pbf+SIw4SccMrCxzkc7kOyps0QrzzdynAIFuvKtHKwnXB5r+HnyuPFcY
DkaTXgXSbvtQ4mWGWqWoaBNv7YzFcmvAYIsk9xmzSOATGyK+pd6XyoDIs6fip828qziuZTnKK7sW
sbtlJU1akEdF+XMn+KIvws77IZiSB7XCTbD1DCIuwwk+soBrMMVdnEfZjpDOlnq4WZu4g7vfTqJv
W6qJ/bmuzGEdTTc+hwd0mMP3ceUNiOYzGowCYlRuELXReNVDGSJpbQSmOCX4vs/mR9pYtBe7Eso8
O37w1OKT9mmqk0AoxOtF8MdFRZyEQOt9/5izCH+KDRfzXdG5G5DCuTHa3005eITqcF9NIrVxBpw+
IJSQ3gEjDEp7SonfzAWmnWtGiNejEB5VnNP5CDtnIQFndkQJ+SMLgWBHx/89m7ogvU9mszc1D8He
T4oj+vwuOw5JY+F9pWh/YBEflbD6BcfAPlxtqLCDhrt6Ift+GXrIKWEX1yoaqmT4foWBlKFVNLVd
Dc8ioOGOB6wXTZMDXNOO1KcLxl22zQeAXISV6TszWOPOFBAgyW4VJl887if6TPL0nP/W5xKY/ULD
jegbsPjjCkhe5nOuBj41etjDfcoJ9Z+Hb73EMXklQijhZZpDd8h+UbntmWieSmtvdRZ5f4MBcrCi
+AqWlplYhurGYHa8tCO3p1QNrX0ZFCb6rCXoRbgO3ueW+S4YHxobVP6Nw5PJqzk5jwzKmXl38WE3
fLsZB89ZC5fn2s4Sl1AmJPAES/jJ6mDSGPrc7AdkMOAV1FcNQo+x5thlPx/jtZztgLRq5g65xk0K
4NkysD+15cw1TBCoJh4z/gkv7RNm/jYrR5e09O4Nisnnq8mpt4PEnPTKR/merfnsmwKZZXGQZ6S+
Bu/RRfyPKi45dyto+ZVljo8mnxJTOVC2tmDMLcGIGWUrA0Zspudaz8YzkHkYPcAdcO+DLJ2LGC08
fBTCtbKWuOr9F1R5iDVyXfgNMwRnZn4OjzEkzYZe7qSUGJ8YlR6ilQcjS7eyfd07KuMLW7pmzF/U
e+PthwovMoptQPIEexOfVRiSRu6JsOgosjz84Ss2rbVTYuMrlPpWaUPkSz9P+xh9ltfTzUy4w88+
os3K3CCGW4WII6Y91KY6tduRTjRBB7fjyqgNpwR6tBMXhzNI6rUnReKFjhUZr1ye3JldSPB30/Xx
HQlFr8Ob2p9o8g+0e7MrzEwhbyQsmUL9CbftvPrrDRSBm2ndDtJpvmZoJe3vJ4UfXf5JUsptWdR0
rnezJ8NJHkbX31vq5MGt+I+iWZ0djhRicmo43U0FCVvSs78HtNT5ET1BdSv1f9711eNOD5n4jOpT
i6pnLWHnlS3KO1PJFaVwBKJJfaIsHkkpg8NWCIedjcOfL6qLqhkXDUdF3Nh3V2e129hEAAn5koqS
HsGBPVmJ87OfWw+T/fMnviYI43I72P63+0BDkC6rpA6+qRC1wdYdHiI2qCKPVhZB3vZ+R5gF39P4
6kdc6P2h+ttldr7jy6UfE2+AXvbKD3FplH3eFPuar8meklqDaT5f+ZLTRvRN9N2EYSYnFSDOChDW
N2fkCnUtLRJdXvC911Vmn3CpVBf4PE8MegxNESQlDk2XCZEIwSqyG3u16OkLOoNJPP68Tb2b4ftd
rHONQXoWh3M4CvP2GLem43aIOwC6DoN4qO55xElaKDwK1Tgu21h+4dXsXuofDWQZbse182QDBBP0
B4i2Gu0iMdlHHpm4hZ+o+1qUIFRaKdia7Z/sLRneaBvKUiCBeHT+d+l3RZdyZaKuNpx3lqbHvrhT
EFyw6NGyb4ucgB+RoOjonk92LsSV5lHs7Mnu+R/rlTH5ui2OaQjJ//1NmjoKn65mNegtwWB539dk
guykUHsObM+QwLIa64vF+K1hdwciGayyPnO7BetFnC0SSUeG7XW8/ylU60FphxyKRp9qlcAByuKl
r8T7T+952dJ0NqcUIAcntnO+VEErg1dTXZI9gvaN1hX5y6aabWrXvNd2FGBt7VxXYr/7ZDcz9ust
Fy3efsxEmjUKjU4RP7l60ELWVG0T0/u5mkPgBj73/IJCy4PW5WVjpqTkdVMTB/5Rk3CaKwbGxgnl
vgA0dVuPOcGJuCBWzYoPHK42ICLISXvbfs0qWJf2YQHQN2GPucmRDs6Fbpoup+zQ9v8Pe5RV0LZX
IKRNXyV9x5uC9TgTMfh7sgRXl79WL1acTk7Oqn2t4hJZceBlK2WrC/xyGQakUuslqsmQUW2xwn36
lyUIXeKV60GhQBPOfU2PxJRff4G1dAjhu6Uba8IEd2dZnfLLjONL+Bcgstn+iFOE5nNlshEpapcm
4MLFLQG+HxNDihfVuYsBitE+KF0XaGk+HY21dsFZSyV+WAiwrJduL8oD0fE8XLSK484yy/Xj8DX9
zP7T0XGxewxBW1LULG1JBjKHEuLifg1VeHsyAjEeiJuRJkoeDP72nwNB1CHwDpMV/NtmxaXLG+s2
+QcP0vuvYEYhbyxQQcqQzXkz4kOSvRXGZCY6S5++yyFGAFhihX9geuXDjVWPuuEK8TOzPvT0GUiM
9q6QD+iQwLaeI1Mg6A0fHAVKd1e9mnE7h6f6PfmOWeSo+aIEtMrdD2Skl0pg03+Ql4f7MW9V0yiq
FewWd+YySafY0We59Frzvvwj9C8mct20nKmhk9LR7LCpah1WwqDDlaFq/m3YPG9oZ6EVZFWbr4hl
T0BZe983YTvmACErFzc6Wpau//wPrtxcgdVRd03H4XOJwnDH19uchWQwhzibVWhqigUuxMH/gm3A
ccv5iAqUuxoJ3QRJJRKKfxIDYIxBCG20ZcazIElOsGOjLJlPfRysJxR5jqkg4QHjQ1msJkHx+7T6
fhXWX93x+AKB2hutqfJQunsg8tEhfN7ePBqlF4XbyQL0wgxSdK4Kqx9+Ax1N2WN48X7ye6PRqlmw
fjHxsZM88Ee6a8CJUfLUbRYGoVCjx9yePk3SXjPozavxNzRAi8IdXaMEhwGzTb8ebIp/dWijPjFG
GSSH5nvxLyZUqk5bqE1TYq4ADjCljtI/sRk7QyCcOnbgYElykJbYy8QjjEdXegL1Mai1qIxRkRZM
hypspue/rkGnqWOar1doeu4INZQV7gv8aX3Jjx0muxX772yAHvXSptlQsfm1TFAtRaNY27XLiqOn
cr8zTtJSr+5S3wh0p4anuFKmVj0WYUVXpW2yGea/qfjFvftuoP7mEpWQ+VD9jHitZ6m66tOERWpZ
5Vn2WSZz83e2HJBvQlgQ1hUxKM2mno/CdRV7qP40EVDPGtRs/ssw+LgPbpaQyVJKO6qxdIpmkvqb
JvaMrAZMcYS1b41HJaIEdlFi3TpTSoz/eCTTM7UbLT+s8AOxnkDdSX8fV9FSV7IDzLxcAT/GHqsa
xnVgjhJvCSyLq1esMm/eHBy1PvVHnvSZX86vs5jV059QrZ8pCs56nWNshk1jj+vAZ8hMpE6DJ5px
Jw3xgFSHqysa2LR5gtuu9WJmfnXtMbK1HRva3LjkfdaqSF8WvGpmBB2ZocwupGIhrUjerIdRYki6
63Qdgin9L510DdQfygJssisXkjssKEmkt1EudBv6WwL8asbtRq4cQZYl38oBzc3nicCXVmcFMFG9
glzY31mMAawr8Q7HdCs7Mecp06KK9i7HtCQqFyJzmTL9nNiIfRa143gIBUZRK0L//X2PI089M3nT
a3RxAasFyxR7CIpk4GMQrPeH3hhCGWVHIqZuGG01cbhJPtDX92QnMeuNO4afsW07ARtkyMivgZ91
X/CufHktZ94K7nvbUJHMBfjNT76W74ePEMu3KRO0c9AbNnp8JfnkT5dvMXefEFfyvM0KCCLl2e4I
KkDOhz4t1FCeUs8Vt4uEtPvIMGgGWd5TOW+pzBAFsMyt7sp5tvz0CdfRVAIhbvPK/ni3Sv5OORTO
5LSUNfw51dIXG2nw3Ig7zy1AZ+WtAT+Oih/oyZ1o8vU1ek57dC1dX0BPyHsaySmLrZBcBX4sdS1z
oiB/l0CLjBl+e/sSy/JCb8EC0L+cb+542ZrhpbVVctq1vgNlFvRrJ1JmOHb6s1ez50WNfDuqLsAh
5qo1gGPRiIvynVXcUXOqs5mDHN3ZuHcA6yoTW/yz0AtDujDtwVw3DMqDAirtL1pew1Zwe1HOMA+3
pMKDj9+6Zv6wqWdS5RVUe39xVZzNPWS0ZnmdkNdEaUzjdVbunu9nXKd4mKNqRkGw8lZ7F1oXZNBa
qzwO23AmBThr0UK843yCuZPBXfKlV/jsQ3BSCODU30mllaPktmDC8CHAD0j/gvBGqmtQRdcNpwyh
5/ks8wfG6mgxkFLi5qBvwLa7GOyCzoCyThzbNj/7iWnQt+IgAno+fxaWR8UbO3g/F6D0iA1vP5hR
o5HFbNi60cDslS0diqj7l3pFSw44+Rgyqtf1m0u0PRWxypjKVL8XRpQJ+zpnVTkOBdAXb7c/Qnr6
my3c3Jsk/fcGcY7tLPXty6XLsFj7FSnS8JAWzp4J+vHDX69Fj9ceRH/HnSlSD86avLtjdmnNmI48
PW6YcERJpIICK5qWN2eBQIWCGx0lq+jFwayGaIKn4WV7B2X2Z2UWirM2r/MJd/Srm8Hm+BjsqmYg
ViHZX+XLvsXsFmzGb2vRtdxOqX8bJ4699CDTIG9JVmmOqvuSumlnRazblDe/b2NSMVbcKFFwwKdu
/WF/RL0d6c9ZTS5pe0Rh3VOct6HY147Kf9qWsIzAUeS2G74GA9iulODEi1Fgom7ZW5m4ILbwp4KE
0q9fF/VHbvhZwjfmwy1sj/7/HJMZp4kbF3A+psl5xzLfOh+pytDCJuA6Ht8IHZxtq+YMHfIFZ/M4
yhjB+oDTBm1Urgu5HCoIG/yOhvWUnV/rMGj9X4zu32GDOTttFUEB/kk3GL9xQLJNKp3S04GDDI2R
mpdjk7w55EDitOFdeKcna0Mnbe3I3/nKik9MoCnWfTsxyhcf9Dka83OdmF3viy13k9p82YEN8Y1N
NqDZC1szlS4a75B7psHbDvq0BNs2ueJWSY1uAvcKW7bYiQ1L7Va31j4zdcJyfPUX9EjZC+WPduP6
qpmc8VAbfNjN5uTP/Epa55D35HiqjrH6vujaHt39o0rg7UcLy4mY4RdEJ9rRXcFSQodctWmHDzll
EHfKlG2xjC6YdFHvnaklgaKyfYwdHX+FUl+iWXeyXbQrpMOJpYxm2BxHduKfFWap1q0xpdRgctJa
/VngMb+jienZuW6+e4OkJMZQLBlY78DbOJZdwiP1HH9PSjJGVjOv/JZh+p07cJFcXNCA4zjTMlxw
4cWjXLLmKMgQ1zvEdXigrns2CjK7W1cg0RzTP5vsHSaMyggtYMR+3dN+j8RTqnToVCUu1IGV3acB
8U7o49tU79jKF9fbfIG9ZQQMyF26aIe2D77uDGT7rsd6glfcpKCqt3REwSAP+6SsiGxXlTwCJqlD
6813XP5Fc9xie1Vdkkscp3eqTTTl+P3AqOvwVraevhIf5bk/UGGr+O508tNObrnBYb8+Lw7C3h1+
iZBQNxDQHciC2e3lUgkqm5KogGmeu+G0MNR54Ei2qvqfJqkD1YH8rGMPV3yimrIDQhWLdvjCjcv9
Sl1OkumrAAUlB0kiHSgNh9NFfJYWDzM0uASFCoJ7hfU0ERDU005ibmsf2HP/NZosbrRG1EwNx+Ek
Qtz//wG1ganZcKyafjhtnrAS506gIjKG3N/viok51Owd3U95PQd4ZytEqZlIthnBBcgfNlCk3ZTf
CAHVxZB255iHZhQ/4X3VykGPjnTjme1XMjx2UflO8cV3y1UNk1+133ihJw3//MvSy4DMwFuQeHfW
9UaR6jWkpHZUOTYeeTtBYyJtQjnXvTOR+5IPkhHt68h40HlJv/X6bHYcJYSpWWAO0y8v0C+zErB5
aXAE6O4hhgDtHm7pM4vKK9SKSs0uJq96cLcKWQpxON7Y45fdq4Mq7mS3QKFqSS5EK4MnzVuD9jkO
6UQdR/YI/F0jm9vbE+7muMNSxe57/jM8joPL/HDnVakEa6NFZuETSVjlN+nKkFeurc7Dd8GXB6dL
eCShotxYWNMYZzEFKGKeL3clJX3RlbtDi39zlmdprhngOqJ0+CLiCs8he9+DHmTFY9r40HJa5z9w
5R+LmcWu+UX176M9UmDkrRr7kLCV18GC92MoNXUYXiBBRNyIMCEa9u+cHThst9WFfjcMMgQwIXx2
NxQS0doUf35oEuycOpvKZln92A+W1TKu2N87TnxAqZzY/iGaeicuBihosDwTj7VEjk7zZFiwz6pV
hk6Guy7Fh/0a8VIAZL/LizK4JuG+3gtyY+hJki/EO6zw97pBPeAUpSo6LXjnpdze54WSYvvrmDlW
SmDCbiA8Tk4fEwG8J6vEj2f0S8/G0dSWprQ2xHKu0C3aJo9denpqmM3hs8H1Q341gR7u4M06Eby6
XitQfyeRxMk4yKxJmx3At6Jft1kieJYGH5qGiCQ3q8A+H1YMDCFZO/yxL9yT6DNR1nDnU/+t/M73
yqm8wdKVleyyOIwBQRmdPtKRg/D0d+mWU2JO7fTPVjgiU1UYD06gN8wCSCnK0L+xwmf4CScl8t//
7OV9Ug5KYRLDbyVBh3OC+RcIr9lsLpzj4QgpY7c8E6U6XHf4hULmCmF4GOeOib3ReMP/4D+B67dZ
Sv8ZLFZx+UXewScXIOnp3KlT8n3pMVCn6dkcJGxwig6pHMUdmbKj+E7P6mrsitI7crJMLxedNSRl
s5ntrmz0zY/MKK9Z2JQEc8NnagHc599tzD3Dg6y2a8OOrOXO8iOZbZmWR/dNTIdX/AApCTsLi2ez
jlsOyuwMNlSzVGIuQ+2PzDlKY9Y/CAKV/gW9PP5CZ8V/jtAIzxOGOkAq5snjORVnrnqiYNiF7hVw
mAElBT4wo/EuTFhb+28PfnvQzN6RzQmSQAV0NsJsoR/cmNM5OCRm7u2pYqUn7p5vTNk2sbz2LtYq
SOcE4mWGneCvhsFcMxWofMRx6XQaP0LqpdB5at9vMaAtmKSPRg7LdgVY3ZfZ5AuuGgBCi1JD7Kf9
qVg0HwhmawlcifdXVuzxz6Rs/CBE28XnBmpKLLHxCLHHP15RHKlht3I2HR5YuaG9oNnIg2iZHOvF
ABR0EqzPmMc24kdrcVnZgAVYvbepCRqO1SjkcHfedHbgYhDG10YAz5GCuQGW3BOJLHxoLTT4THlQ
p+z6gwnMJHGOkzUr6bwvS53QGyO4y+1oEJRD6fsxumDAXfQ48Bf55/4MOrSV7bNC3rfW6RZxlt/l
MjhUYHBswIFjoUjsA2s8xELRFCvJnJFoOJLfksFk8H9ETXdkflCOSKx3HQLp+g/NakbOvd7vv/O3
JXbE65+tp+42GIaUS80QrEcZgq3cE2FgqQcqgHNQXIuGM/TDMwBgzhUhRmSAs+u3ZEpqojNBO76n
hiE4DcUViIEZ+AQHDedWZSjEImD22cb4ugEUvURoRD70GqySJ8gHwDn3DeK9VcrlT9lWFR1nEhfL
mYV95YzePcDuZpKkDutofF5w2t8SpjUs+VyxYJIOq20Azll3WLx6yVw8IDX752kVOuOwFC3R8iAs
tzeNLBWkH4d3eVuYX+C7w2WIDaaz6FtmJ/YArPZA2UJOxZ/AEGT1EEy4tSHYy8v+ZMN2YPqQbO/I
oO8T7knLO0g6B+jgKjGAuZ4OY3pNJuVppACHPTa06/evp6fFFWrLtT6+U01xk5bfhWnMMPjoynSX
xEo+ABGTRGcP33QXja+ijSsghfCEq2gUyS1rSZskQRSKoTkpB4L8XF/csQFvtQKy2iuKAk4c7eGp
ybbYAeQpuUB72l5vVkrqbNxMqP4/y0mK4wLzaVV+PBuCyZ/qcC2GQpYk88LxYQEYKN7MPc39mz5+
eVo32crPQJq8jVu99xCdTcS0efBRTQlzyppHm528EwxhUO5tRDYykEWbLJtZwX/AKxW1ghtDjpEF
Dao9S/79VjrbXSgt02HmnrG9iUiwOswykBmZfBnLnTOCzGJo+0fPZtpZorERIlTlgAA3ZCmXEbX7
axFXOsGw20Q4d6KqLHRKPDKbH84b0WyIIwQKAUDM7BOjtgrwl3d34eDrjQxjdGBaxMh3qfW/J8jj
YyBH8voMrLyR4rBvWG6f9S4N9LG9WcMDG6PARTLe6UaQ0N7HjeYF+iZEtGwEv1zaqUTrib+sBvFk
GHS3oRa3NvD+G3CSRNxE4baBfL9z45+J1KkFzqxKLtDwTCqS5GVgtnx/BU9zTCBeMLp6/7H+f7hy
SR76cuh34ZWaaVvRseHg5OOO90OKvGkDlpVNE2hTYEIEmPF1eWR6cSvCSj9V8naWxYs6F5A0Ybx1
YXl2PpOKAc2w/E6z77z8NzYrXZMtyb8dikGUAfmfjonlArotGxzAAXPFj7lHsT7fhZnLf/a3H2Az
IE6w+kgr9C8LCFKNBkDhGRPV5sGry/cRWG6991av98NvOOJGph0Ynly1S3fXB7j0atlJhw6mSUYE
6zwIDcpvEoaUTZCglENrDLCp5S8WttXeHzcpWg52ZceO/8XkT4XBeZZWOjbA9u+nw/rgjixSz+CM
WqF1zLU4H1Kcgg5jgstGXNqx2PrZMTZ42Ox8Sx54Zr84LMoA4IB0b+0p+bffuWZd6cr0Su4mghoN
xehvklgj8FhK6LnBQ9v9FdDf17FInF1AJ7tnXmp6k3Lk2H0rMMDMQHSfLSp1vAI6LWYVeB/CWvg3
izJr3UY7lhn/zU4eSbFHeglKIwvwMuXCAY0Y9pIoTID+8Hy49aPtD1Ua/XD/DzgrlJzcG90xKVTD
t6JVVQ0TlKZWm9pCpuQhBly6xN3SvZKPgq1rNe0DcCm8yBfWUVV1T3RkOaX8G4QP/SEMQvLS/Bwg
CASdTcref6ex+BXt4+J4a6cQTb/wb90pUeADgMtS54Y8Rindq3OKdXyjGkj7UXzYdL37HYF8bA9n
1Z52J+jheJe2oZV9AOtDVFDkAVmMmsnLZPToQLK5YKRDnZXiNt30yoSgOijzfbUkaXXAF148s7+a
qtCxmfYVxVjJZUyq6BRy0cklCcncC47z0Ih5OlT3zPnsDMfJIPiTXFzZKj+tri2cA3Z+8IwclU7E
JehH/jfrZIvFCP6UIDEf7ZcEj2s19jEKqMDGsazA2dskTHlGd7nEz3DUgrv1li0Fwzivg/J1+q7C
YuFM8pokeAxCM5kcY4c2p1H/yjzvuUbwr0xO8OKNQXCndd9O0BDXG20WcUF3mm76rAXsZoh1dZMb
k3vSJDIm5aOv3fuSkyiFr+j0qI8VogGIwyQX47IB0At9ZY7sW03dADLcjxpwMzo3eojiCx3Sqs3D
ptMooYG0yHEtNMFUuHdlfphtV0RUces0HWUgOcb9t1FBwuymOMI3Pw8Jwn8SLixhd/zmQ5VOLrrl
BtlI0emNWKV3puTfQetoJle/ohi5d1g7n1+oSj7pN/+8gYSMEb2MVGZ5j+hhiT2xXu2apPftsIhT
FQQHgEyYkp7yUWKxSBECgpqmcVMrnveEWxCGOIRz2am714uLw4FkWX/xBo3yOCaH4QC/cb8xro0e
HWbgA4p4h6dxrYff05bNIvJ5m9Pdy2qdNsP+drzctUi5cdLgyEbo9DQTOQg4queGWF8+pK8scWcx
x2pwqNw2framYh6Z5PEMpfImnBnian6//Y/PQKykVP2isKpym0u8MzjuCm7Ebz0XZgE4Vki4yDgK
mS6Oc+qcXn7emXQI98J3lSIATXRJ/zCv9HgBEP7yhcQTycQJ9KMSk/ZgzH6l8e7NxnBQccjHF/cT
CoBnTvuFHEBfMTbzRn7vAO3X2xuFYxtb5PgttNln7OK//BCVGKoVVZ+Febp9QiEtggAdwrVR05HI
FTRw/PGYT3WGni1/eJz4D8dSZ61D8OVseGkL1FJgz87ERoxxKeDr17e39p5xVMJi5AYWbHkEwBQT
3+zyxFdo5WBTcRynP87IRR0aneCNAIjhHaJEvARSjsLNNq4ozxdG84zWXpCb5kwmPQHgaNlkZ2oG
O7swU1Vupd5MsuV7kFY7ge068o14zcyFeXtfNH//Et6eyaBCZUyF9KPf35YBvwWIHRPJJbkYO2XZ
1lMeohYe3qaTlASTFgRWchPK+kCrmGEmgcEv1SGANliy/u1zpVaxCqZAL8sYLSbhAcKVJJ1ojnqh
0VE7WNYKDAh0ksAZsBPn0jmVBJjnPzGdl3Kpf7bJBZ7PNTQvLi+oVpoUqy3Ed0bicWCSu91qr/J1
TWkKtp41BYXtRUDcOvqTGF8vrApDTq3Yj7fj5HBuSBOY9NXLiL61726NxQfhEcRKuiIDQOfZvwi4
uaxOmHNX1CGOb9ZlaIsqDYNNWFbKYm5lRYME/wIr8P+tcGEX7TfZNHBAfegtbLOvBkL9XdWDmcVy
E2VQC6z+HAJUbB+Kow0CsG4tMz+wfBf1lEJfDyiUJL3G3FlpQbmVwEMPphmTecoNt65/lJfF80Qy
l7MK9t/eF9jj/odjK928IJk5v/08m4PnVU54wTUdb0xjs+Ch/espINU5KZmGf+AdhUhnL41xAqjE
mqMlqTvwNpnbF6LHZ0lbInI+GX7x1ghoERgcUCoNYrFzq1Ea89rbfoakA69GQM/WXUMzTQLsnMgI
14wCfLiAAH+/4AvQFtTHL/oUptgkNxrcIm9KQOP/yO74XdHnsaCagRb4HR0FH2RWomOX+1MJxL9b
XhD+QoNCnl2AHQE+GO5cVVVSI4i/jI/ouCzlmZqE0xjFhEwX+OsLh5/HMKYk3VM7whbeWs8UgARB
JvA9ii4kkpPy0b6bt65oTHyqu39SPk1lndK/jWAF5z8TK3Sp2hFP5C3dvPvQ0oR0FfUJlmm5Nqfh
ooaV1ekPSvWMvXf4CyFLo6NPnimy3XhxSa9xiuR3dWovWAvAanc16xcyJP5TfTeUrUKDkc2LRILt
wLlD9CR2qpyNFQPBp5BlVZ4OYTAUS8LZTb6OKJhSXNQUlpaujeBbS1l79Th+cJ79G2IytnVedCf6
b9vqgXJGLgXwTWdcdKnmlaAdAkoG/KUzd559x8zFlFVIyLxxyC7fNUejrPgrv1EAeUCdOalTL2uk
nN+DmACsgiaRvnwyHn3lNaroJpKVcvEaN6GMZ8jgvB8fzdVdAYbBn8zuhhvMHWfhHr9WuSCPG3N5
fUDYA2bdlabfQGIbKzZcSsB9AyWhlxU1Pr9UBJY4OaGZNrD5C8WXfzL3j/9OCso9a/f/PSVCIQ8z
orWCOHdrxaMwmnULfySD4TBO6i/Jeyaz758KFvCmt9FBOLdpcsmwSqtxzuGa8XmQFPOeZR87RuYl
MFz8iP9Gm9ZwII8w3WHh2J7pR6ZyLkqji521ffUBCJifuCyfr72RsRMZao9lwYbR+SZPt4ImDXao
JetGRXN+odeMjXD5qvLdStkRD+HAbV33UnD1rretakbVejhI+sF18aX7zngFeNoD9VIZOmG5v8cJ
usiZ16XWXUm3GSZ4zlfLexGBBtBt17mnRCPfgYquGEXnK7VFudgEeuqj9PX6iCgGDmbIbGRAilzD
VWIu5T47nY+yskGdU9BMhSzwtFgAjQ3VxIPbHUha+Rp775LXSsygmsfM/kFek1tuezagVGtS6om7
oyJmHOs2/m5UFOnbPD+K2d1jYARAdQ8mLC4tWkG5zMowsAku2Sn9W1GuoMkLjhnuhEXRHgNLYYGb
lCXt9aMvUtqZxXoh7rd7SNIF4LN1lAI653e2uYpKGJundQJzT4TrkA7bm7xRCImKYIUi/ZcKogjv
D1zyRomRSqTAcecIB5rL0Z2eCWr3FMhRVJAYvJ0X+fCchsUfpE6J/ytN0RVlD6cUw3+r85yJ2A/+
04XZHP6tw152EJ5QogGZI7tzxzNlOU4LndudmdtWMvKlbMOJGnPnKvt9PMXUXHUBmH6phZkOvFxN
Fe0hvNLEJ7VQOg6o+NopbXAGqpbxO8rBl4PuuwpJTcGVD244BpoubgRg0aC2H/N1w6FhzL90Gvu+
2/Vtt4X61fKtYTS0CpQ6YgASDbv2tXyK+xz8Ct2bsMX6aZTPgTacAEwzKBZn2mZ5v4B569z1VyZa
RwH30F3uGsfHr4fZ/rwdP0z2J/6+SQ7LGQUyT/2tf2eC+/MqB4O+68IzEZ+eihUOqj8/Sg3z+m6g
vGV+uaDzFxToVa9dtdpe6IbjfIiFEyoeidRYrblKfN5d8EgPEG7VN5VA+DwEEhR379QXndAN8BXJ
fAEEDn8rNOvJpIIteShDgmuePpDqRO5VpLqeSOOuTSLHQkl7sj0hT82Vc0haw/78mjxn/ZOb+xoP
MFHrJQqxooqfk7ClpuaYwEF6Ad6uEN898SlXIh03YoZ40kSkGbh1IILUs+FRGavobQ2njuwR6cBX
Ch9Vq/d3u1ejKKa5CuQV6MU6HJ0ov4sBZqyaKkd7fr0qmyTK+xC+hHp9Uzmvd6XUrAHvQ5m8W0QC
e/7x/cVzA800WMuljz2mqM3adu8OKQyxRKyGH+oJT0WwZip8upjgareU7HFOYEq/FlGX/UCaQceB
yAgakuVLJEBqNcYLb8ayvci9c8j1PQ1TvS+mGaBAZjYRdw0wsZrfEoRMCiMLh3Hvu9ncPT1td34f
5hdcjGZjyTDaIlBRBwhzlR6feHqxBKQCO0hX0k/NOW5AvO1suwN+Ysh4jaNqpbJMra69DHm6gYxT
9yTx+YKBrwh2SkFNe+avpFk9Fjskh2r8vZ3HgoH9ks1y0gDjlPTcpESdCciMXLNdmbfPuAvt0wkD
rJ6/IxSkf9oIInfp6B8A6AexpZ06lCdLqQzMqT81UPYI3whaeA75WkS9jRc8361jGICvrwhZtzbm
x0I4iLVupts/D/35vjXVj9/tZmjgIdD5o7+Isuev21WKQdZZR1h52IcCFHBV+WvEwIkPEPOLj8f7
pxVVY+FYUSrxkzB//WnjQAScJcgmnXiTkS+PK1js8JvHh/sa6xul0DXTjHaL0DDV4jGmZNBpfcmM
asKMoKpkIKaoVdXeqJJFFEENXg7en8yADaOeMnM2NAomm6R8DY+cLiRRxxgyJBQZwsXbeWyWHyS8
9Ahz5YjKYsW2qbnXPPDOpyCLVn1tZ43hpvCock2V9sjCtkFj1O8kM10kOkdYt5N4VpwYU5wNrZ4v
gLaT6Rd9ggrmWTPlGO5UDA2ifX49A0dZER/d3pyXTfljysQki2B503N502MvY0orTpiTFNm8DyvB
TP36ZCqs8aoOjYxjYz1ivuhAGmsJvErHeAhsMXxPUqcDdhgR93ERd5B1bDwH12K8qXLv1vAZfku6
dnJs0JDbZSAEGnPMRLslG8dgTOurLL/sq3ijATLc2iu2e7KthzYS15P9dNjycdf4H83RbLqqAwfB
1+MSIGJs72n+U18LV3wJ3cgqLj8Xeyjj1SuMWwVCANIMKO+0YNpxuFQr7eOXID2xb/QhEQ7RtZrK
+P2vBu21iXE+hXO2ihV4gYfHD9kngpUjO9g3X4hImczHg1u9yKbmhpsGq7qOAq85V6KqnKdZQ+zi
0IpphGfBNUoodCAjJAGf70TPP3y+YXK4g2bNDPUWqzC5HmoG4j+p9Ik/IctZra3krovqkGJvASZU
GREzScwwEDb2CGj+9gyZ5pXyxuaHz9LzzQFDG8oLuCeFED1tvfHqO2o1sc6xYLWakvDRoD1K+lbn
EDOal6jXILJmosZ/ikpLaNexvLabgJ4VbDMrkeQinArQbEZE/kn2zG5pLetEE29MHMTzip6QqkzX
pzd2GSdVn9z4Azdm2WkAQu/HtFWZeogarXiqom0r+tYrDpjKSXkV2JgOf7BMZskEKj6O7pXKLNTi
xxjliM4OBCckYvz1axktxAde2ECE52YYgpgqUDhkZIoJj/1KWnviVlV0Ej9XSWuFgFnmQqVPbLMS
NcSnr669WWZBwzqOlnJtM27KvGFm1re2hhS5yqxQ6IdBHOdi5VW11jMlhSgARsVUWldpPW+mvDdt
CISeKKkFK2wBnHUX63op/Lvfek2UHW9UWpt5MB13ibupHOMvsPij1qDQiphI8a9C8ODWBYWN9Ahh
KEl2h/L+kROuwfPShRL+YrWM2AB6Yf0P8OnwmlEJO5ozhqsiVv5MXS37667BDCwIsqmTWSjmIwW6
xWqCyFC4c6tjBsSh9ZaWl/LOOiUafZ3FWErpI2Or0EI2aZH1Ub+3vM+/w0l/owSaD1hnBCfUI1R/
2sKaduU9pNaQ6k7GUdcqUK2jN2ro/BlSfIlIxPm631ASlzfStcPTH08nV8PmbHSZXTfxSVnvzqeA
QTLkWSJIFcKGysRqiAwCAdF+k3ClNei9FYuRJyRECl1mbQTMXUmhSEFeXuqKxy8zTPfWg3Vv8Cmd
K/4iNzJRFJvkDiqLiZCScUzflfO6rfO3mOGWnQmtsNZQKyKMdtggHt4FGAA9CIx/DCiHi4qiNz0L
qrHFx6Gf0n5p+tacy0J3o6E+hb7NXVyuh3zj4S62NNstQgrfY71bHOtpeH+ykpGOwV7fsil1urzy
rF4frz8DqFCzXcnsuZnvRT88tArVKkxra8msRrVV7gnNDmQu7GL+N8TW/QEXrk1IGoqe56BeYbQl
WrZ5K3NOezWD8PN3MaTo1eMA4QL3yunuP/QQNx61jJOd9yihtLFPUsTQUON1xjOYjnS+EkNcbRll
xpAK6q4X+xVmBj6eHSorTmqKjjvGrBeOZfCeYrAVGaHbbgktF4KMC8rfCegJp0O+Viog3GFEwCX5
UVDZUYZpg+SLzrucDKbgbqyAKsIGdp+IboeZqFMy7IzDT1BX5B17ziyy+wbMu4P2j76/luVNV3I3
YXmvv7s+SmKRCAo4+cjfAiYW1NoxjDpCD1KeyvrEg1VxZ42gyVBx97Y5cJuanhCngcJIOqcrxZt8
m/dI9QnnqGAdogCEQyokn2NmWFmaJmDxydfF99P2oNCEDxg0SmYr1oJgSn5Enl9YKgZVNyX2ZVy3
pZQW5NczAB9Jy8hyf0TysNLJ+R6ja4XC6SQht7xZ8dimnYwUX+St3EdhlVQWFy2gFhdaEoccoqSf
cjgR7I/PcWY6lLk9yZE07q7vEpK+ao/tcrBiwJfqDSPMma/CLPyhUu5FSxYCQe004RhTGKnxMce5
jrPCssAyS2Mbas20j3R+pSBH83ICz5UyOeSu2l1d8/QfL7365hWH1SQb1qvqfSUpEeyK9j/6gjmj
nGlhwdk2AxKq/6ntbDG0gDtvKE2LUDLVROQqIXlbejoNBDUWgWXjMGYmrZ1MJV92DV3zmarKBX+N
KCR9Y/K2wE0wCsGfpbdg03rs9HqaV4s9d+kxZ6kl3TxizP+XOqApGsqqJEiWwE2vOpIE6NCgGb14
56XvA4rzFx3VxOo0woINioUqIgsIkrsi7R2zub/EghEyDcuv20GWDjooPPW6DErfKp02w+NSeg3y
CpuoPrTK4LuT4Y3OA0qeGFauprsVcQj21FB/Yh/rKMA7WjqdoOUW3aiGMuMPNH8qpk6e8rtThBGt
RXC7nbwdIftHmkPSImOcWn6yb7b2etEW+V+JBN53YHoag2FqQ4/Gq7MBMzA6paX8/lRtukCEMMKN
hjH56yGAJQ51PiX1lDW1TgyptjXTuh0OwZm452jQlsyBJCRw9li0txC1l2ZmksHPn7zQ3x8aFeMR
0P40/ZF1lgrviQpgpG3Ro8TOZ46YsoHBj2Lu/m4s4Z0Kr/wTU1CaKXoLB6nLGNFtMkT0ereKi7Yd
0yUx5Hdbpta1YPJOYXQDcILmO8UlHANKDjA4JwrE4sUueUFPqBHUYC09vgYYs1ALMIrdSGrNLzoI
K6f4uCEJoULnL5jAcG4yy0J3V8GJYwcoSFie444rsASFdWeudDp7WBl+2TRxRBuKBjT1rBylzNYO
xnuirZ40FMfMhp5GbCEbaSItPUJsppd1KanTU4cnkaMlb5b2Umjgs6H17B9WbYUGOYQkE0Xm10fd
NOMfyzf+LtuqxxPdALM+RGsLtZ6fI6/oUaokNeZybjYtBtCijQOG3Wz9D55k3uElSVlLgDfamqhn
Pf4NQDfmtWBKttvKQtKPLSI2HDPO5xeDxHxnsIrLSjQ+BAg//GZIAUY62rAlbitmh44RjCEJmt0x
JPKjA4GSC2+q5j0VQSHRW52ncKPVDcoVd6qsF3IUvSVyjN68Xh3Iw8aBYZ5bfCCyxxcPNGYIQLHQ
SeySvp7h+tPHluGCzZGfNW/t4dgD7UY87PGByus8Ow3JQ3A2fnz/ZNRGrYMgJcrA5GsFuv+TGP5x
SmTMB6EYqfOBJWKoAOwIawA4Dny6hxqPWxo/QHe4Eof9aCD8g8eIeJkP875mJ1Oai6y2wR+S9ECP
yzwjgNeVkyAM2YHv4CLhjoI+szRLOiOFgP38HZnDPJdOkG9X7EY/VYnUYEDb9iwHuhGbetWG64Ya
8dnBtPdp7NoAmPuDJUc0hxmY831qmynanHMiUj44u4wgugWlvvUrVibYl2R11cZlSONyVc+1odMy
P7vH9wJgU8UFaEC6chOftFXW30YUOM/AY20GkiH3hkljoOYphFqZJSrt5qBphqf0ifrS73Z7nV4N
Ex+vHLEN/AO0QXz8ES0Y+k3Ns59ZWwUxmUWO82+s9IfcOWBfjfhOwKjxMbQeeAKi+2u0IcR/XUxk
bH+Cy565xHjlx86h83p3S1bM4TMPEFMHRhsSFeZX8iS1fIhnuovvRLOYFm/QF9cE9OtOxWlVHHIC
L9RMs+9pshmz5fqy9ZR17zdqT5Uc0VQCaSYLqGKmiG1t7oHPslKf4POwTs1rl9/ejiKc+ftOSRWl
HERkbHei5Yj/N0G8Momm0bP78NmbJeW+zWMe6fyfL+oDZ724SVzWNVmCCCiEGq3XsI3g9+lPWl0d
WyHFKR+rbYFg6dzYpzP0wkJ03OKMwDh2i65vusUymnNy9/9VMIk9zxbu5jHyNHhwxojkXFYqOqBP
X4wHNs2dPymP0/owvPuFzsm0lttvROlmG9aAo2LTtLPST6me+UucQ7cz/LAsAj954BO8YOkT0WjH
M2mz6QBKhvTI4nqCrhLz4LKqPqzc8gQj/JbVLZzBBIJ1m7osXPSBpDFXdGrCTfuoSeVBpggbJV1P
2TVVcLyExLwkkSrW5ePxVQ64QpfqT8ovUk/Gmnbgiu9zECObaN0SWHZmKEwCr6iU9jOX3Z/vN8C8
4AFOYvgtl0N70xOFUhGIDKaSclGXNXe3FAtbgC/xNkC1QGVIwdhIsuKpYvSEHS7XSRk71Q6LoZln
+vZteuBJ/PsB9d+H9CcVa9AWwEb3cBQ4k7EMFATuHcryl8orTs929FcUiLu6JFGBfvrYctvLixSa
vg8gJn3wPdAtLrtMTtqn48yXkcuBbqQLn/AheiNqnd0yJFRsqrdJNRViAKxwnuAEXbqHV3/SmjMa
KBqr5dsCXUeMx0dycjaewr1pSuvaw6mzYPouLpOba+LFiZIcDSn01GQ3jiz4mbQkD94/vc1jE1GB
JueJ1NIUsz3zuEgV/h2jdpyAoDDPPCxvte47wFOPJ/Uc4hzwRIN50mrMITBIzm14EJZac58nUFxt
zrL8pLImAcY2QWa3hbO0l1oFrEqEF6ReCi0mBrYzah1N3lkxcPlt9Al5yiqCf08Nf3phDSpjGk2g
x6HYXj4GCRYJNIEQvnXWutpKG5hG2ny6VQqNh+fMYkp3uYkKq9Q4eElRf3kXopzSwyiLV4Fr65xN
mBb6UmvEIKwFE++PJ8q55lGrNwjU34nUVoJEvIMftLnS6TCWKv7NFj8WOCEVWGnm0JZVzgvsWpPv
2/o3vJW0s+xhVEMNSyydV/twLb+u2svPco96C0Uq3TuABCbZYU7qefI3onzLEZMmyc9RsFdgbMIl
9bAeWbpHeAYqjP/pZJAwe2U7kb9zOj4hudKOX0/oLfgOaPpNiMRO5Mc49uae+Pj8m+Z+ARddkCvF
Z9DeDsHtsvN2v5zEJ2K1p6TQCedEixNJkQj0XK2ASQwNqazvJb/8vYF39uxbvmO7XeyLs3ccEUej
T7UnZ7wHnkjPX/RaU5JMg6kWlLaldFdodpJo/hTjPSxTOXX+w9gKOkhCNjkLw1hnhLpWC2D9OEu9
1+zSnd9dzLIB8Ws8johufeFL1ekUmq3/7ePkBcp73qvK931qnXbYqaaPOuq64hB01utcI8Fm+biB
8fJsXJ/rKK3cIR1Uf8MrbfCtMeUyWux7B0rffSRmfVoB75cT8XSJ5LAMPyQkW+X0F/LuQPJ4BE2q
TeSmWLFqV6SaLPJm93XPOe7ApjgyOEsLO1fw0v39Ja+jQl+1Eh7a2bZYLfqs121Wj6PIKwS7RLbz
ni5mwoxGJ+ulTV0spbCWTcBMIdEpjjnhcXqb4f3KCtRvumnK9z9oyUJJuLrjh53/nlyWeOMoP4lT
4XfqcUMtdPAjtUOhHKU6Ehafz/VThzKyzOtFBzWLYFBRV+sMtfT+TkCGP+vjUpo8BKyloYnf7qwP
0vApI1FUUXTutYbr4GeKPQDGvd6LGYvqZh9/QM5JvkbE8kyLlC2pppIFbpWk4oCWw8EfC3v4Z1vL
FC4Qr0lgRntIBNruxVhZXzr3yKH6/cUffsChJnUhZCRzaKJHaJfAaexm4Bhrz87g8GGBIoIt7l9N
QtulOSxE6WOw+fB4l9QslxRhSssCMSkvEv+eIIWDjou+w+BfEyhIQMVqpHG4hPBrg/zKb3HPo7HB
i/+uknVO9MKX//1H/R2YUUz0EzoYrWUA2dU0Xk5GK0jNmMOPNqelCbrPCocVpyTBvPwp466wxF8z
7SA5E6zlW2NFCTVmbNUYHjgjf9OULswCSHPMQ+2w3GNVpHwpUY0nB7UhIbqmOEMOlyotvZUwjwBJ
uJbRQrdA6hCWT2gVMm2YmrGxIy6ZcbSNi+PsXc0OnWwukWXb4IqUB8098sOLA+9Ldi2KMCFSYXXN
3CHBFz0IiCWadUUyLl1LxZUDQRgXxw7SkObhF4c/FNEeDJMsRQ2/kctMhj2j7K1dV+8TBxYXmyPm
StTksiEN2UtXWWtYXWQ+zCX4MJskGcW8onAOjlcpry9YpwX6/EAekmXo2HVKEjLsVDj2XKxiHfae
Xmy1T1F/syyC4udsi2fNs73YaJIXUTLhqiEHg7JdqbmERxz221YekW73TLiJV0vxxZuCKDpn9io9
dL8wwSSeViZbzzFsmnnRFdwTyPDO4ZOK9i3RnbDKBkZAvM6ajBekmMTB5RXnQXIgxGqDzsRdGEDm
dAnzqPFtln0jRxIL0uEKj58ug82LYjJ8+YMpnazh57lKxk8kmrTyUwdmXdDWkIjLjujV8YK7kVjh
JromyYaGbijBjJhUlVB/1E1tXf15ePES6v7x9Hz3fRobUJvTfOtImXsdMQ6aUYOJZAO0P7r7arPs
ZDkt5yZJNIbTgsU2zjGHhCeexoqu4HnexrhvqXPAzuByukeiDtCzDdp0XlT0sgVi4kk8gWSWxZ2Z
nj5S/o2rDQydENTQnjBKXuWSDDlSSE+Xb4xKBv/QW3PLZAoQbfM98Oj4Sxx8zB6fp2tfR7Tu3Aa2
rnIA+LmYP/ofFnPkVL4HUkPLnGaYv5s/qIlvh25roVA19m5DckDrxORRmR/TTLmHDXlxDn2b9bYm
Yg7+8m+26TvxKnBObi6PPVuz+WCTSDaqt7HAmt1SyAlIH0EyEEz2rh3Rbsk37aEK7PN03jmLNpi6
03KIslZDgw1VsnBH7iuENm2HSJCT9bZf2LiUaGAgXO7rzTU2K7hpoN/PwWYjO0Dx3IMpqptkdXu0
ADSP0QLjcTT+G0h/iwnYY8K/u8unFiIPUfYcWX/vUPVSHcP3ca9hewXIy9NBaU0gVvH31+WTvuZR
1F81vNxc5ySLCqKSwMrxD3Y73jQh6RlF1UheG/VxZcihJSqjtu3AgpwoC6DkaV09tomuG/0awXvp
UuR4OalhTrgaldptvP2tK1Fw3yKo/B31CLzzGIdrBqq1Us/lDPlOuYuyh1+i90cNPKu96l3Bz0d7
ykppcX6bicGxbzsPdTGj8cUJxbnk/Y86GRZXX+rmjeMT8rwKEscPVf+I5vZ4eqftB5KWxxS7gkTW
r6b5y/aE/wHVk27S39CQQ6IvZ+kwLAA0GJWGk2c2UttPHdSjCn3tr2QDMpspr/OCzXkO3kj/dwBz
4WvB5JMJdcxbfBnK3FLf8MZOpjISDhvy80YpztNas9Wk5BFEemuYuWVczzUtRZr2rT2fGWGv+OHb
4vCsaEqnW91K0o+CWX+P33rGoZWxUHz/GrqMBhDbG7vit+HnchidDUz/fNrRtZ9OFicUZJHLuE5L
Sx5aqTuCokBLoTfCTx+KJfb2EmrvTdWnHSX2QjhATZxQhg5NPwNR1YALlRem/Fwpg2idT6ukOscm
pw7/7kt5fUwpQ/MgKPJL4Lz7Xw68uPzg/YVKNYPjhhfi6zikANvx39YaQQ8yIOdQYG76+FZ5kXni
QQNaHpC1L+EJwGi0zxz+a5WMTaZuoJr7podR8n79fC3qhed5p42xDbesHP7xNL5AY07pbZUnwEl2
rfIml/+eDbGhxQ4a7xkkOu+s9nkMx4fFZW7K9qwACaEsMyqg21wmW8klM17ghEBnC9u7yvQUPIDt
YW7iUbBFoykR3liE3iiPAMati2GHUiHa04QCylG4dK7nyGQSRWuZGl5yypmt9jWz+ttM6rhxBG7W
8kD8vnX8pSsVs1TFkUj6MyYY8yO4hR3FsZyKHDOEnX5GTCKBc7K1+BxLprm6gDYNFys0QPGLSucx
oZTo4IqY/dpK+7QnQ+CMsAcJ0NdlNSdmdGoorI5rE2uz+LxLUqOH+qrtrXobeDdeAjLFzykHdKnS
fDpkEB3iT52+tbKWopjPcKwoPUrPJxrQW35JslAL0abL9W+qqK3xGJTbI02Bh0ht2/OZTQae7rgR
3iwKhi9DAJxwcWyObI9N38ECXLzC+l2Lt8FSEFMsNNSToVud60vzCisJkEyUZZBRzRP+8YJNMUOX
W17pdr5IbSC2OL2GzhUMOGOYe3nj/M82mNnsH0gXl3dTKeBFKFCvuLnnvcNtPlqBpDOdc0apJ3DR
eZpG/1S7g4qgawV+azePhjDOt4P2nlqo4dM/LZUXcc8yw2Qp08gPvGzxVza1IzUiA4zKwe5QsZIp
U/Xh9QeR+LANuSMQeSvt/RjPHSO5CX/9fj1Tf8mHVegljatsOw+W5I68qjAMKfFSBneKp/Hj+xoJ
gut08zYgw9U+CexCS305lfAIY18c2yZo3aCJZmjxXHMZJu+l0dNdonM/5EMFaK2i2KmU8CH887Sx
940uoDlpl2qiCJn2cjnL2fKPFA7/dRX1UAahig12qg+At/qFTOnpYPNZjjJTjPzk8EuvS+3eWkH2
POnscv+5gqoxorvRZbQ1Gh3635j9mNbyxscARZA4HdaGmNXC69lGGJZildshjpbIc8cc0ymFSbjt
6oUQggWQDDQcR7V+5s2kWp3vX/67aQOTNE4sUognlTIAtM1pHPlX73TCROt0qUtLIVrC/zm+/qzl
UM/1obzSBDx6/RsM2SCRVCXjioez51eJPJr1yCJP6E2sI25vK3RXIStOmqJRiDdry61KBlkLgynx
0O3rwcUxbH+ajVU1c2OO9R+uwIBa0I9T7pF8AYqfjWVVRp99YyLJd5JAS8pQetK4FTfEZ8T+lpBl
DLqFHix4rZmg8iFWO/AcXZA9zUtWXEXZ6aPBgU5uvxTWVIL+MbeJbXH/86o9OiqeHaKT0ziZZ4GZ
lNjlpj8BckIDFlY6SYAZ1LCbRGuA486MZ1vIhCfez0x952uo++gK8x+TfbdhD4e9neOrvp1XT74A
sCp/9AuifBw54MNePy68H7hIwgd28/BtNqju9iNu3+ZrlMLpzml6UfxVE32XENxkoTK3dSL3npH1
OLAovKTnurlJzC/04dUbZpfXWStU9+PUtf3nRbxCMAOzy1MAYGbysSDQ22GOo78gDmkzXQ9nW1Jj
gKw1LrhoyyDjqwxARZhXjEsmhcjWeWyZgtZXwwx8kyXnhSc1wHxrnnjyU5sigh9QMIvXLlNlip/D
xixi/tzmkG9gFyYmNXU/MC5jGTvjvlBXp3RZRksLwRwxeQwvHwXQrRrA4lJ1CZpPum5p5ICH2p+r
ufqiarRYe5kehq3PNghwKY/q1FS4OS9uC7IfikLGm49jL0ahAG9ymER1fei37zFVgLYIyrx+xJqi
aG1u25vy5ETxobCbHUjyNL8HzhgbbT3nVmatCUXON7ajD9cmoJG5+gP8V+FRJgePOeQqTvo410cP
e0EkNm5mhGtWGjC8is2l3yj+7sq9VoxqczsHSkeDhwHpAYbklY94aOW7AbfW/pthyUsKsq0hwAmX
PQWfIX35i/G8bR+GjueYc+8Lk48V23cLsxhQjom0vzqi4MtYzQEb7ANxqO+N9BvNczWXtRbI3tMl
y7i5KvgUnc/X/FfdKRTRUtuMtMVf6PghgtI11x5ltdZnsPDl3YPCZ/JKqrd2boyhZQzv4X7QXAeX
lA59ARlcypVhJQJk4GePrDat5/z7cmptUKRt4FD8cwTL1obslOXGdvRoNlAQPxPq13O1zoMTIg6V
iyEY7LKlhN1GiOKCwamvVWHw6P3E5kcoG8IEyxzg84B/k4/7eyscuUJDUK6M3KsV+Mjit/Dn4e/g
ErV2wtfKKztgK4H0+2jSH9cxZQ3zKMLRdzbSDMD30ZykXi+uPixbj1WTVyocdPDwS2zZh88NcoMf
fupDOawJnWX2kd4Q/IcHm2gHAlrzsOo7ApfTrTobNFfRG4WVKoLuUq7f/YWZY+qFx5vpY+DHhB8K
dZmkQPKyeyuDc7vHhjdQTc5mvi3NvdVXQA4bU2Q26DEpve8XrPQnLYdz/cH7EtYw9aMC7mRb4j5E
i4hvfUizrgP2krtKRXRnz3xIo7nlbpgSpxCaVfALfvxLngBW5hWflIDnIDU9gGLOZ6SoidOAhgkz
n9GhCvOiKP7cTipCF35vHrWfym+tPm2QtJfr5E4QMeOObUk/3RMy+zgqP+z6rdhICGP03jh68bQD
N6AbAwsubsum3mnSAA39vFGbGI2hakRSzryQdnlAyjav+/Qz3DAzz2gaKcmhLoEVyOUEN52RuIAW
1+Asrwjks5mj0mWEqCVALB71xkFrMpA3MgPk2GpkCTvXmhX259k1NaHkYyFT9OAYXzo803THQvYn
IGEJuK1QoRabWK2kKtgx+UvEYeKv2GpyLIZ+EOyOEsGvqsXSO0SNxj7JMhJ1WwWW6wUiNlAslFy2
lP2RqzuKS5/XiXTe9Y+Xtm7be4Aih8pX3joGk/SyRPKubTVWeOA//xuFm3POjtOvw4RZbApN5I5I
a8Gu2Ceo5iP4iFemm+jRZWuaauVPCnftkSTgenSC4tVgvlYVtEkS2mB5yY7boHGX7eGcFiFRwXeL
3DxWy8T+1Pd8qB7xd74WYkqq6dN8VAl9q+h8FxjL9+uKi+mIRM81p1Su6qwSpW/1gQTQ/z7M8rRf
4RHhi2s0DKt5zOc6cca3hyw1269pql17p80Wgk5dc8m1/b+5KGle6Cz9tR+2jDFyc/VgeWZwFZX7
rUHskgixKKU4YBPPiKf1Q2u2wrMQBNdvsMz6QGkLIW2R7XZ0unE19HfTwj/Lp82jHIQCQTFcA4jH
s1YyWzx5r3mjH4LDqGq13CgTcM+CuRdCJh6xIUf/SI5U1DqtBCPF1jHGcHYqFcE01j5DGc2on5aJ
WgJQlWO4ySJw7/w6VXJtGzOCMCFomLszAjpQ8zBflyIzci69h+3dY86cCTq+jBSCqDhE70eIUUmi
19i5WXw+YSLFTyvAnFmwn+WVDARwD1O7DZT1bKJaogOwbfHdiHSlifK0vrueT5oz+I42tg3xac0T
G/VzJVXIPVFR7R739okz1jNiX7mT341bTAc02IDSmcvm/eCZ7eoUPJtM30ZeAKjbbigGWAXuwbaU
fF9OaNxbP7y7niZyBhfZME4AvF3nIYKJxZ3y//8kB7pB3MIfo7alEW4T+Iju7wMq0E0nFUqM4nw4
QLmzwvHvokdSbOkmmR+PqcYxh+nmfqXhVh3tIaGn1xJ/2fV09DpAZUnfAuXYpWLkuPjcBDNjmFoa
WCt7eFHycGsN0g21wsZOsu2UNAOFhcMpTJL2lsfrlNk8kp19ra5DtadpfFXQEfgbTDyM0IFxJxQ0
g6JOLbDi2PUjobphle9WdEdsn530JRpuGprL3uNYKd8ii6KczmGqBugjxj4sh8AVzxwGmfp+lewS
jswp49Dui8fFicmCbjS60CXE2IVLOizdvllILLseTZ8ff1d/fJWNFzZjDm9h1cPAK4+7gwoIEyra
BBGtfw7Zg8I349k8lpvNFJ3IDxBnIpArE3bHQB+7TunXzbTsCxAuiBCTIUX13oO+jvBFUlg+VFvZ
5l2RbsSXsse8kO+iJN6cHhCjriNZMrAl/WolUlWU2bKAgDXlSHeAb566rr2Gfc0/fzX9WYMt5GUa
K++yHhuHopIGzIeWdPv4N4L9MqwihGMQ/1UWrB1SoyhmmuG1H3wflhX+syZDZSOW3ptTIEWkEILR
pzrZZOx8CFA8gwhK8BnlpSV+Ty3vpOFNCvsRGQqUCNSRLUhPkKWgLhmw1IwcOHTLerBGnk/QJSrd
EH2UhrvD+MkkmFngJvv7gWhpxipPDPMw0LtfamcPPqzlyy9ZGjHGPj5KTUdgg0XrYPOIxx1VSXgw
jjqmip6rOQydEc8n2hbTWoxTGz6V2OnpUy0Z8xDKA35uHSipaqWzsaum4//27gKAkzbE3L7giii8
yCyC+uCPAmUxhJQFVVir/AcY+3eK6T0sne8r8V41VkgV7bk0nxMEkJhpEBjycW5pqQBHWDi+fLmL
Sh2TtHdGeZm1pVKP6ijRf4JSTPaLPjeApl3MNLnXRDoPDpJnyhSH9MhIaBj4xdtiLtP4lczi952n
MInA6ErrH95dmOOGyB4nVy3XGcG5ykLu0MLxQ/5wzskAg4M5QyaEOcIEFaK9iaNhO2kBPR7/OmrO
0wDOv/vSbO+VpdVqAwMoERPFbUNkP0gMqv+YfYtCkUkLLbNKRgvYfo1d3PxdGPGk+8t2pyLInNDZ
vmU22nmFrgGeag9/qfWAsrXVHFm5kGvgic+njSvtiMxX0Jh1iqd/Mpn4/Rfj2Na0yMbjKJtHExw+
tCiBvnut5aYQSRT6KfjEu7FHG+q0fzM8AuhLviJea3fJirQB+nEhM3+ey+Y7r5Qg/OrNQnzmIZC+
/RZ/I8Ih8z4DF8el4gP2Jajzda3bpgulAWdhYfirAYMichwNEkIjGEm32Fke4YEJGHG80+onOjXj
E3NCgf34DchVQy+v902YS8qRBr9XJCJPbmTMdgfBB8ZEscy73+SO4jKchS19K8t4ked7H2j9Z3H3
ClxfjHYt9/OezLOlQPqKTqiYbQEfiq/TThhnU1EBF9szjPXi2f0Avl9QlFjuuU3YJZnse+WdNPJ2
CH69Qd5dOrOx+oKc4izXJf5JzZVw27+8wsdby9Wye2Bf6P3RcD4B1i/5hIsCVL/RuBqSSdJD2IAD
momy5AMjt6awmz8w9d577mkmzeBHtUsCuI759GH/z5BWoNLiUrRz8AOIkT8Hiw1EP+TN0kWFTJP9
x6nHIqPfN4nXroXRftmwOK3Q0+HXs/pLz9f5mej6HnTRULNMkRFAqD5qaRPOBBTpobQjB2wrlTxl
wy5XW0SfnnGln9grNE3rDEge2L594pOVOa3SyBf5TL6BFI1Vy5JZ2uEphUU50f8GOjqfU6qJe6nT
fTkJUd6Yom8yaDNHPclKa1HaUPTVT4ft4p3nJl/fI7FZwkhWGILTUiVyQHz6VkfvtrmNTltz+WPd
9KhQn4A/LMQWVR7WKR5OXjFts/ysf53fTVDNOSE1qeKExTQJnoe5NaLNpm0cHtGk4/z5Of6fpT+0
Yf7wColcXT61OmlLIqgapLQIOoyynN2EljcAD8DsO7GRmh4gCn3IXMDdwymxajw1CJDVbIEJXCEV
R/fC7ji4huIGks7XFIEWWtLbPyTw2Q6aue0pI3+ISnsFK/ZhTO1C6UvpkgLcN4o73V4lh1W5l++h
teBNpmBFWjWL+MbBzguDRrUEmDqTQBXs6HxjaVEkq+Ho1QQgk8vTU18N9i61H1GJa+cRTFu+/V/X
p7VS30+Coip42I/mYq4MtMlUFJh6U7u99K4su8OSIQ6GoJxw67ZL1lNv8lA5wRuZt1uWeZe9hPP5
58pt8QJxu7ObYtzOwrDqOd6PVPlwUVPuhVGzWWQdieHTkbxkrfZJOfXjdh8mkZ+qbvtsxv7ET3V2
SNhlrezga+8Ur27K4WeNTymYLA4DdB2C2sW9STwfQU/Ck3duLW7nMBVYO8Cj44/qQcYNCCq3i9Dr
rPoe0+0L7aTLounuR1GNwQU2EnGvCqUQAbFnlWESsQNHHgVyLJ360iFAYeFv0x56+neN2Gf0IMbV
+FJZJUfZkEBbib1ZWIILjg4ehCShrIPVsVV9s632Yy/+5KkYud8kViFv8AnamKgxR0yA+1FEt4pK
sY2kXKkYHxn0bqzLTq2EaG3nvAtDbLWKWDaBvgUFZLOiXXlaDffv81whp6tDRCfOL9fi11cKaQaq
rST37hyNE5SKaGVI5ZSS+3MulDEYg6OmnrsD/gCCVWqxowbu4M7ya44PrHqqAivPi7zOKCRdYwsA
L5z4QvG9KPyKmWuUJffWLViC+m/STPFgiGTow1mVRhGtX2/WAxWklfDRgBVnCRu/Pn59mA5NMl7b
Is3cw+aNjDkRltyN4YlCEeqgRs9QwXhY7w1EkqWbdjP6DCCb1le8bEC7YZ0UpxKl2hWZB/Z06FPN
SdcK66Tt14jxKRy7OzdnqPBCoaeSaURTwSJ6EakWYz8QehvBBQYFidBlB04aJjYNLZqFNzWw4SUt
49II+0CEyWfKa9Unxt6glRK+2EsmplMkqLDGaqaDjwgDL0rI6DfYRHlJbNJ+hb4dPebtfk5NAbPV
/4tpe+YdaA/R5G01g3EAnrqvG9yS8kdvCN5+9pC8xA1lxvmLbZqN+WFZboxh1nDtg3x62BqoEdTY
V/wm9fAyOvS+q8lJWRaHdgJJASNlLlSB30DIzGFqKAm8AceXh6/u7CdCEgYzunjxtZDwe99SNsp1
LdUE6em32SlY562n3BPRgRwUa2JfWMXqYOJnYUVMFEVUwZf5dB6/AZtblS0rncvC/fx9l2TaIL+Q
kXxqb1i6PiC3irbbprDn7z6rJMawrYXsnRb70K5XYUTcYg0ouWtP4pSLbBIV7n4hTqZj4RvLWT+n
SIi9hITFLiKwqtjyetsVgG6ZEqczpG3GLXIoTzM6WGUgWgvBTz7YuesjSgWRZnXyt9Dg7TOIbYnE
p3tiDOSjaDskZD1HVbwsR4QLkj+3Au78VmA38AVMNzxAetgG5vP1/KWhY/CyQuXYxMzhzBLOdtKy
80lHYtotgWdistdHTE2ciEL019tIpETgUqstVZYruU7lLeF2CGhmjdIM10YItOZs0BxF3CD2yZhH
g7w5kRH3p28yiT1d8p7lNO6JX2mgYVNz7fgEp3d8nQc+79twgxCbA4L1MQjbfLRosXb22S57MKcz
+GmGfnxmt426twwidmGPsq/Ya1wzmFdTl5gLG4dZc26FXYSOleRUhcNyLAdXR7i6//HZbqk+S2Pt
aW0Qr8JT9iq2yrYouVGpc8SBpkl1yLRepVxNU/E2km3V6ylbw/Cxx4y93Gi29nXrfzdQVmMK+yLB
otgLExjdnc3yMxHJr5JOxYoZz+T37EmOzR+KpITIlW1x5WLXYXjSA49q/d4C9J2ko1awPBJrc0+B
Ru5pEXOk5efgM0Avh+w0uyffwKjrzsBzP2zxwyvJ9n70OFvhuVgooo9+m4qgC+IqTJ2K2rL3XVhe
J1m17ICONNSOoSw/JZGDOZtLe7BzVPWESktxzrsAaOFoIqxxFnFZSQ+8MsRO9I1UOi7Ne8J5AjZq
hMZ0tg8//r6V6EU5dRJRl+gao+PplWuNZh4ZtJgGJuUimt7vIRN3IBwqp9oNFcIUb3BvIRYpkW6l
7eFGbk4FDOIL8EVfm32TQZ977vTlqDxbwo0X5EjWI+AsZtZgEjE6qGKLjHuVbNZyteb9lALPSK4T
+7gIgHQAh5+LgUh60agRJhamy3RKB4psZZgmP/v25sBEhmOuDGqL4s40k5NriWN5hvT7Mb+lBleu
joNjwyLp6ONHtlfjN6svPlqco7UnHnbITc3dqyQ0T54AfS11VgbWh2D1yLtg8uE/4oyDhRSzFaua
xKAk66Ow7Xm5Trj9hoGVrEkpiQc0l45kFwWyj0mH6gEBCUS59c6fEv1N/5yGjsRITYdkB/W02pyP
ZGb/Y9HCa6xEyPLh/s9xBvjPIMJ1SFb+mT0UVPsuxgYRgwQVCH7yzFBNGt215nRRnm7lVH8Yn5dF
Pdk4RASl/cF/mFhQdARkVP6zn7uN9ZAV4MBZLX1qSBl1X992S4GZwk/B+jjZ6NW7tITlsSQXg69/
xPxqtQAkSC0ggVdOau+5/KO6NhFC09JegIUIh/vP/VDqrU0g6zu1Zy6Hili6n9LS0FHIRfn/siI3
IVmlqs/qXEP29/w1IdL7Wr+zqopa0NkSU8lpxROzHfjM8UFK1YdycSoA8BFVX1SegoXmLFxLgY+R
ZQDn0pv4/6gqXtNccTMxkFzy93ugiSi9xVRijnAPIySJyvrDhw6yGoYkl+5CmrvAZhTa4G7vTRQz
lz93zGLcaIbdHrucPDxGVU4ZLgKnu+1p6kpyYwlqdZKDG0YZv/eXdKk6OljFVpi0HHb3RO4la/JM
AXyoGi/jKyCN9ntIlGPurb6bDCaIiiwewdcQLOoUhHvWbpcwFxWoUY5FIH2A//LwkUusUtQlny2n
gtNC2BanGc+NHCWIUe8/wGCvTwjp7I6D3Bm19qgd27QSMkxRa+l14cN+jF7OTb6+aOciEm+rnayX
u46X4tujhAD6wXeYdClc/RrvkAQaB6hcgfWOVGUuIoDg6Yqn+OS7PmO3dl2zhhV567aB82dIonb1
M2OelKPeph5ssEYEqELnumIyuUKmad+XaF2uK2hpWFzxvrPcHMnpnAAlL/CW37lDO/2KCGoSv474
ihRmoU5UJAypMcC0PLJ252/h+laKaHpUh2Sf+WtGRlMH1FhAtiqiCaGlePfIXr8vtWfyk07INntK
1ukCjrfDWCF/jGeqiZkOXHlk5yzBFek/RibTnqXllFdBCO+PglXUT9EbNdgrnWpX1ofSA8a7mjAr
oCr8YRwZDsDNQIfuzFcQCGVTcvhjOeRmcxgWFGiU27j9foJ8wDVvHuBWN2u9D0erSx/mo70lDmGa
o+0PuTWy71d/0mRAQWiVGUOVrNBI5TYstFv6RCWeMed8Ry9m8RfYKxUqd1jAwYRnd33Sj0Mzzg3R
SyCLiEQxIttXZlrI1db3v2HV7XdZbrz/LChwEDR5th62aOTNS2gtaZSDNm8N2aHks9CQTPf+OsPc
H9qeYLDyNJHkJPtank0epnNM/DfohnbBJLw+rPvDUX+X/VJziHCTu+46FqkLbfR5i2rzNwFB1ah9
yAigSkI+IHR/GThIpwPbZT/3nC7M8qs1nNgeDfSS0mIJsV1VmGjrSjjBv+jgzUjl8PG9OF/L6zg2
iCsssDtTW01whvtHufmk6VitkVVfShxbZu8FF3E8x45OOr9F+Oe2fTePcoz0V8CwO+GrEhcry0BV
xqVFvETcsj8KbiAGHi0CSYwQkP+D4RGew4dv7/2AqFnYlIXbhAAB198DJxkrwzDcdfX6+HdeBgiO
8XN50Wd9jX0h/3xG4EiI8OyzXrnhfTu5nJkOnMcwct88/DXSmPBa0eu34qTXSe8/f2+TEWqiiupd
1bmrTT0TTLWg4w5I37X69kLgIrrtXi+nlvu2SWD4She3eUiR6P6y1ZXur438jOmJz4wkjTebu1s4
5TFSaPbkX5/Opy4yZtKYiLwkFX/binkGd6FzpnTErKGLjZ2TbSE+2B+VrSwITIKIuxvXcKBGQj7y
JcQ6M3VBuS9H2bC2y0fvfhKnubF1taLvx1aSZsV8EHWp/L87EJMPrunafY8nJzksMxTqrnczC6zG
G/re1PFAoaN6vC2sA8e7hfzoTI2xwzWNDzeGK0uuBtyE/tTuy8lemIkAEjYEqQyoFw+DkisQdQEf
BLxWoEZLkGEgoj8k02eoS5Sa4pVa7oj3gay4U71yhzXIVeHoOjkmtzr2UIWBTXnb7HXi6RGn6UA5
OcYz2x1nza4jwM3MyFdCGEozAqsmZ6CEVmh1fQ99rF9icZx/sRXTUkIGQEoWT0rpc1NdyxtixtwF
GAzXVnM6Jk5/2HjAZq+RexciQd2dmb6U+rmWAI/w3Xfr1fnuLSYWy3geHpSkJxqXShYL37cJxAC5
0s5Whzului4ixk5EhYt9uJCZeYYeqtGR5/NiIFIYhN3LMrlR35/GeUfEAptdA7fiF1BQL17rMISq
cyE9HvvJkqDw1xqk0HSACIylAVQ8+zg9/Z4rYCAkOiJsrDPyi1IQVqxp8YqI7ac5fy8FfsqjoWSW
L7RDJf7v79K76fm0Jv3e7EaiwV+3Rce5VE/jHVvLWh42MjZJjq7b6LGAIVPnKUU8BlENbf/796P0
0uciMGDH1PIr3rmG1tB97BNsIuwK4+vWFw5b7Q5Jm9oU4TkFU4UmRlfKSDHt71K+fBRblR8eJeN8
7bj9OAM4t1gGVDMhxkacbGeBoV+lpeyuj+SY98VSWbaRmN/8EmqBl8nYYQIDadmgqNySauA=
`protect end_protected
