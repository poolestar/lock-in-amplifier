`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ms/kGAvt+G3oDCnERO1eycJ2b90ZudbNptdHH38L+Y4GQelWq/dBA5+w8lehdDT6+wilefUiETrd
yzOT1V0X6g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Ma50tP+5k6PHGNbYhVzuZHTHAlUzrRrURKkQAn10mVQ+0FA+BJrnWXMKGgYaN5PW5jLKRkqwH6f4
+OPU50BZRC9O/gxpvVVAFHL58/d2/vu5JIbeAxandLPAFA00Gkku2vG3jj5JLesjKHuD6dx6X7kt
ltc1Xgv5gMIosw2XoI8=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
V/moDxOKcJZbPbLpE3UFgrzhtYX6V25CwXFIfGfgEujL4kSJhdHeqUaG+J680LW90EXDUJN4mV2Z
+5/J6wwTqHzq82YXHEiFHyVn+UKfS4SgLyuITAeVkbGJ7gYIetF30b5cEhtrK947V6NfEdKEiDzv
+finYCL7sk04MMrJamE=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZeR2RtoxAcS+eEvdoEOH6KignhKIkusNMpfM3K8fkH+CyRP8yJGwkrYREoL7pglF8bT4NyO/nnN7
e94uwKTGyQV4b75DhIrvlVZdzQb64e9V7E0Hkp58aVMVrlHLaDoDEzLv2NcufFLAROTHeG70dTuA
psS/MdUEKT4EIWY4kNfxRbIrPwe1NVBMyZm9ANTNsqFv8RztSt8Y9DmcsjQgPXvdjXH7RgOe4UCH
EyqxbXFWetb4BHORSIwRDO/rHW5zc5FMALVjZ5Pb3ST9gzQpNKfcg1d2CmubDXPFLQVhqQllXR4c
DtZJQRQxunJoURUONXMIbEV4nVEEVddf4EkOEA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ta6p2ELMVjppL7BP1tvafGWa96MSBCL/Efwc0X2wpgefM9qftoAke5Hr9CQjRrujaAeRDnx389Xq
ZCNCqwMVw+BU+QtNG7TcRy6KVED2eSkQogAl48DeT4eRRkdOT4/PKwFOYOf26ioPpeJX0KCHBA28
MrYyWDTrtKSlglqzB5lGEQh7MTfAMHZtKzsIZ3dH5/XmiHxWuKotsFMIW7+4vyUqG8iiz1QgQZKa
rKhkzZh66Tw4SaWTtmiFhOWUmAVGaA2ycli9svcdoW4uoRHZmubacxWVrupNeIdSUUZNUKhIUymz
OYtEXLYMKXFPFuJSg6Lf7HSKNTzWZ6gkp8Zgmg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ftAN96inAf8l6/mVEBs0oGDx+TLuDZe/J9VNNs9WygRsayoieIiCpDcxcofMYgCYPhQjxmAueFDa
tr7WJHxy1AtHMXRriEVgahexvtSLFeUKVltgt3NwoM5v9xZdgz9vtzruyMokKiLwg/J7x3DVEPxx
zZGnmoyRfDY+Jz2HpbpFFKridenliFuNkbwh2gGNv82CNMIIVMDFt5la3+s+RmGMgAMPBHhciUp2
iR7N3Uy6PAo0WHs0CynuNPk213K9X0hgntcRbDiFysBjCKRspfRUIa8vLasutwFQ7KbuiaeV7qrG
6GU4yaAXmnAqkTUo49a7KmR7cx1OMdkAGRLlNw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22944)
`protect data_block
DIWu/ooX7TAF6q2+XfGjIUT2sdZdtmKzbksvsOyNupeGnDC3woyApoczRRK9eiOJ/GfG8iz0iX5l
JGtqVIAGSwst+cZZUXPpe+z2G9XV92N9ogb22y2xHqlBvb2szFf51/un2OjPUNScnBXsyRS8trY1
kpe6aaDXbpJvbNCIM32O06GeJz2OMQAJageVIrc0BfP6DrUaBOv90cEwe4jLl4du1thbfvv/DPhA
QhH2iEWjIkifVRRxrMfy7vpwqTCdID5LO+ipHv8j6KUP6BRJUmupd4n4j6bdxIyEuc39pxn1Go/5
/kipwYh20YX1AqvCqh0wMyO5PmPJppR1MDWKRCNDIuvWnAr7Gdd746ipMC4SnCpCb5oKIkR8YPen
g7Vqdazveq20Bz4p24nUF0NtgeFpe3TvRrrEbgwZpSJ53WiZeko1aSyyHU7u7XWOJhkmCuCVm1+v
SJPX3/vc9a9wpwmPWbI6nu6USfmT9UvJ+oPbHJs2nQyzUzCzC4AzbRv33SVD374DxDy4B1LRBYiW
er0XVh4TGdUHg0/gVcFOeEISNuA88h3vJeFv4Pb5DuvWKi9vAXjSio/So/CyKt734ynSEnfPmfo1
sLIiqE4eWR9p1yVX/GGObsgyjJmGkciVqQWu5hrc2rrv+P+PUsS/Yk15oiX60Y+zmauj/p5RxuXW
i1XVS2/f04olLzoW+DLGoJa7DtFEDbweY6yu5+3LrPISkntMoxdPv4GqCu8bUz3w3/R5FNeYSezZ
foD1OSQyDY3M3y4qljThuia1ynxVQxfoM/jTC7NK6y/9YUHRIeMHQRjCxUFsZl5OmdciGge63aEZ
wJAylHTA/rlZdhU9FdFN3oYN31iiVZg1By3QdHV8EWdeUSEN2zRR71gawOy/u7LZYzQjvMeeE5p1
IWWFKw/7mQ8tyR+qf431yERc5ZsVlZOmvFYDLuQMvDFj7/5AZp0HJsKs2iSuKvq3twvm1bgb03y4
W3h0lvTDLDuqPEeMJjP7ZlEOSaxzb8/iPREm2EoubeVACniwgcEAuW0uMSFCOxWmg1hu0NIv+mca
OVquemlWA6/fDLLXN4NXPDhkrs/v6YfBlm8+CTgq2KyBCMqNtTnb2GkP4IoDBloiohwS+kJRAb7y
Zdowfa14hVF0pm7FighOmFIuYcg69dsPaH8wnnC3KujFrB5yXvRHDcu9aHEV5dqVMSq4ye0RkEkD
eB4x73EcU4qE9qdu7RTfOad0a8DFp8meWH+h1iFl5NYTWmyHNb5O/JUAvk78ieyCm/hRFW4WhXB5
lvtYdhX7zeTL5UXE1vWi5NE1VLwWCk7Thl/6azv/DSUD+JTzLkBxy4N8s4BTb47NM86vo04zSvuL
/MeHNptZDjSzEzWopJ4wenb2a8B3pRLm6qq07aDOPjJsa+5h9c0PVyidFG4VIpPQVEbXaOomeR/E
NflaO5a8HQzCo4QP4ovOoKXmUwfCZmgOhget/E+XWtEKSXAFPssVKaZAxC8+x9eugT2K3Rs7K/fz
4cEPGkdPnbWUFin3EwmQ7E/ML0UwYx4usBZ8VLH2nKQl+IcUO8Kbqfc0li1shkdaMxyYgd8Z5jzg
WCWQl0Ttspt3e5aLnW+KtA1zVy5FniVQVieM/Vmw1XBk6A58ArIace4o9PCgGLHhkUdVkYBwhkGU
dxahiaRe+vGSwBlQtRy9luAEVY2ORV5SMwzQtzhMCe18ekxESGGaLiLun7aLBVJLXOVTUFZsmUqY
5uc0NoDODuh0X4n0y3n2SCKkknwIYHwgAkH66zT5wVzKKYVAS2wSe2UyuIkPhxB06gAOLAuzPw7N
pC0F9oqU/LWO5JyZglPIvDUHjQL1F6g8pQrL4NQz4ZcttleBjX1dFtiC4uYFHCrUGDljIPrHiQiZ
7fYq+dHcrlG1fUhfuPRasNkpvnGPlK4ide/SA9Hg3DuJRtssCfYXHb0MxO/v8iRLgH2/3tNqAgP6
I7lqBBLrJTpMGQ++0iCzzKDNfXYsaZ/ZKMOfeXa9oGvnvedE4ZRmf8cH73P6ZSjVmwGtQ2pz3y+X
unYJs/iE4JeNTZqF/EVoXZmREp5SrPCvNwTf6u+LhPluJMj1mZ9teGi6Qatm6Ui7k4IPuNCNM+Ol
Tf6+hLRmb6dIPc5lPKfeGp/t5f+hEPwu3pviPeUokgvTDxLhRMEZq1EYzIA7DTCDN5EViPF79o0i
DYOvUeQGQLinzhMwSvoDv6S2m5p8JxbVcZo7xX1UlDhkMPcFdoNGK2mEIUbqBNbN3M5jbBb9bojs
XnTuRA2mDtPP86tWvJ6TnJ+6j6Aglw8cvlt8p85dD+F4GQSWejXzkH83k48ljCxWJpfwpBw5YqF2
xz7NWgsNNxwFfnnuo3B2IWq4w2FFdnaMlMbku57T1yoL08adqJ9xFkDZjeFI3yl5cANS20rcmYPm
gbYgKjiBFyhQCaZ2JBtZI3JXdVMtpUuTvcWdtVbfQ1Q6H3VbW7vl7Ow7kEFTMPx/x+UGwwxablpy
+IwVn3kc8C55uhsJKrbZ7HpoDZctsn9eYvPTplNX1rP91G6dTc4YhhN48GHXJTqgyPyF0JEJde1P
vBw+dGuzTrEd+Qkm5aDz1Ymt65k45bTC3oWLWOOZbjXjz5ME9pmAGOv3Aa7tDd8kr9zh7vnllnTX
czyb5zwshJaAXmlVJbDjCoKoeZNLOvCmmUgUqK1B8hTX/meQPT5MFY/RuAsJzOuG8TlMFtW14f3x
0zHcqHo3KyXZSRPDgWBBPOs6BHvN3ROs9uXD3zofCZo5n1sXAfwrI0hcbiogfw8nQhvhaNv1Rtmx
RW95Nm32ZsZJBsiX8iATIQoToyfukC4/Px5LVZe2bVewCIVMH1jLfIyAl2MZiXp0AfPVcpolGGHJ
Liqk/MHrI3FSzutKl8b1EpqPtOGdNAde4uASLCc+YD/Qyly+F0VK+PKraM9qeCrMRmRzg6W4kh5a
b+0E2UxXIRw5z7uRSNYtyheZGoV6cRs6In+669F+Q3fqzirG7VIfYvTeuO7FlubotmewImH6Krb+
xRLNahpnlujmN6YSPgR1twyv5z8nlbMKlm+N8RCndx6vaJW3LUb0i/w0g1DUyHDjRSDjcDc04vMm
8pUW2pFE51eluyl6sugoOG6X4tlJ8DHYJ8u4bkJP03jSN74ceTq2jJURAYvD0aKPsd8v43IrCHIG
8WHOGJp4KRuAZfTWkMSrMIlnIlPXrbqXxFzZUd37mmxy5ABoixO8v5WBKFFrNhuVmtMjg8m67bY+
+EQHiJ6t1DS8OuhEMGV4hfR1+XmT0BG2MZuQIPfSvnS/FKNUXRRFyIQkzx+nK34/nEwFuiTyjt7v
EKUTWDIIkve96j2UbQSOVeNGkg1OVvActWZFCoY0vFFCVU0RCm2AXzpuNmOUX0kcgECpFkYtJesQ
a3oglMN9B5KsuDe6q7j21JIrVex7S4LuaPzGxxxEsr8LMYmRiS+WMiAjVASGnseyDewcfFfRqMw/
He1P3K54Syn9Q/jKFw2AytoxEv1s52mhx/vwsyw3BCizy+lkcMmgAwceB1KlRZ4fKx7RzDDu2wV9
mJbQg4DDxdw7gV8P5hTLKET8kN6M36EJ7s9DVvhlTICp4pTGOyT3m9zg1icEqfhh5kfNpPkZxO7a
D92cBr6Gkzn7yDwI/T5F/y4gb/8MIhnsdMy0MIgBsyaeiZ9T6fMTKqc1XyHMJyvCLfkbskz2WqPy
imxsTXYFweEBqQEKFkp3Dg2uNJ6lRW7IdG/+pP0be4HsOYk4+Rh2c6EY3+9YkJwruCgmzwkWW3k5
wuOLtNpCu2dGH4pjJBLSMkVtPwGhQQBznX2NmivdUghlYdsXILb99K+p5SfJJ7C+fXylE7HZYZpF
P/xA3s1TEpgQy5konARcyqbnxAKFb2bLBNpMO4MbxhJG7XlT21JNuyn1sVCMwQLWw83Cj4VSm6GD
gi8tjU2g7767O79lKOPmpcF8KFyQ+/Pi1S0S8gAKL5HB3m0LwuOvS5gRUnDEgt6KePtvf1Yg66IA
iys0sIuwYhDzjONFnrQhDyW+6YP7rda20irykHOCL9qFmXP1LhA527AuHfMYJprCLozj7qKid5Ug
nm886IhtD+JYhcWBthw2XpnFTPZRnf9P7acoWAlBag2xXyELYYWRu5cJRpCsWxYMzuy8XbufvS6s
fjuZ09HZgA2ofw4re1VGcRENpMbwjtQLSvPgbt/tHqR0L0tljY+QkNS03+woljPYRLegP3QJe6df
AtuVTvBTsY9nTkQowv1tyRF/+rnatPReo2zSBDgW8dRwcLFnuNCNXmvJiAbzcJtBiOb8osbDypNf
/jp13VGW4rB8hpMi8aiHYIaQWFqK8M7AgkceXX2FuaI4QwqVLb98XqJVNc6qmkSWmKmUl8mSKvHe
Jgri7wm5uckwGACF55WZo0wKJZujGEJ4BlDs0SCqBbaCKVKptHmiB17Yx9/iDH35Obn8rPp0iQc1
R0vmgXGmPtqG/MMNdGePxEf+xtNas+RT3iXpwzpYgJvYmoAhXd7PQHoPJQ4fWgz8LNE1FvvznkzZ
1Qyil7H8HPSV8nJL43mX2WH6m32CFmqI7FYmMq5WkOf68xoBI6DKDeZyNT4URxGH39oGFGluZHNQ
rRK/RmKfiRiaCZWqMo2yyhyfl2/W3VVQKvoIAKbKahddpq0ER+lkqZ3ral1KbFYC2ARj7VNML9OA
/oXqJybH5vcVyh6GMPEPtH16TE6SaA/ux7fH1HSkaXASIAkckmGMTYh98/9f+D4c9QWurO7oTpbZ
skMOetXLwC8+uihr2XjGK2f8ixqVk5W3VRFTZ9YqmrLxRGNRTwrK6KxePEF3/tPw7Hc8JE1ZMTS0
pxDaZJNfMTdmKEHp1KhQXtWhl8pi3K3QoX7jCS2klpZxtxFJsJdYMZ7SsrJTmGU5U9BSAHu3jKt2
G+BsbcFTekZp6sLWxqVITYKXPfDdNNlU1XCEbOzYsWCPlGniLZbdNhRTFdNj+QjUMc36qrDvZQ4F
4UnUxr1U3WdEHhb+P4iKikOubln/FJTQoFFZepjPBu58SgjV38etIwlE1kAdAe8FI8q3gW9ztf0c
u6wfdAAHcL4wjowTOUUbqM49MqkGtzEPigsuBsKSBnwdAVY8bP9S8nl4+WrIquNn6whjnlswGI6n
EhlQ0W3MSsVGYrnRn6IZOnw+JnZLeLXHYrgwNVITz4Q5g/jnvYibFB0790GIJdddYfEkWcXN0G2P
lLoVidB4xWUQt5OWWaxxV0WM6nBXJOCaNZuigWceRDDQM4dexBZIgzG6bA6YIYMNTlA8rFods1lw
MmvKvzPrN9ju3rdvROS+9RVh+/YJ9VHvcWSfT4092N2m8vFhPNE2u6NhMhmfZu+G7N6C8TiM3xFa
KrYdPr2PaxArChjObSF4UBNPcXhidkjRPiSl+SJSb+9B8YZvbhRzAnnvcDdo8DpMDWLg1TZu8uUT
THgrZFc6taDZ0bJW7pcWSCJlcu9ZtpvdoQ5VmktK5RmbeTDHSsBXJR8WQLuEQnMcYkqSyQL8Wv3J
P5XlBnuCOnLfYaXVHc/yUNoSu1+wRPTraZscAa67Y3cgP/l5EY3yhd6C0Ys0m+XC3NrmZ/JCr2wR
cnvwSyJpRUajmko8Tkar0h4pez7W7p1/gHniE7lmInGr2+NrzaiFxGXxIcqPIHlUZfevt6yv9uya
eEqm39W7KrDpFw/WNyihbQCF5ppoIPJmtqPMVVjLfQnG1bBbEJTjgiVgpxLG3HEEhYO/Dsk+SVdl
Gb2CFoToRJQ3qUy7V54byJ9vgLFvz1OEioP32XFH9vaYAUkrQA6X9mHeWsjdfk29sjAPczajCNpt
X+n8gFOS46+Zioa31C6QwUDpJ1sQyy5hYjtuofaA6CYHyXqlgS2danNNNSQTAK2QxvTost28P5S3
nzEBO7MAjelU8f7nD24mQNZc2oO5NWansb0tahwtmMsVG09EgnS/dNH3XpGSbsFDD7hP9ZDB7fO8
pAZkPdPB4hwlmUELkZDpj87CFZ+ZpMAYbDT3sZ1efQqhJSEk5Tz3yYTk2ZFn+9LiA1lUkANA7sds
wjeDtF9RFhUJXVdGJT9ISW0AlDxvwSpYszID03+1xTMBsj+6Ie8v/kdJaFc4Kp2dFOiFDOeDliKW
jQSSlE+GrnyDT4yv+DVFSgOttcle39i4u6hVtHaOn9diOJ9bq87XHzEUAfG9AjjaGLuYZGsNVfF3
9JWYIk2xQbjDxAdNeQiZS56xNb5SSunuI6uVFDaTUdHh+PJMIOG35uF7QOOHJ3Pbvmdgsv6fQanB
hl0Je3DRmvYSBsA/DFSMO4D2vZ+ore4ps+3MeDwn7PJ6OORI5PqiI1O65L64f344aN/qV9TM/Jx8
w+QD6KkBZYXHkl7WnZRMVGRpOoOl51x/BBd6qovkhRoLTkCZe09RbGwk3SzRUJ+Uem/by6SmvaqS
HkCtPWLAdZENJyFUTPVmpLrbh+DqKXaSFTnmjoBkSR/n1WAaR96wdsWW2b5U4D39L78QmgjJKfzR
fbyQU1yUxf8aEe8rlskBosaGk2bf3uRHOWnWFP99ZdLayes7xobPYAjxzchicsAle3mha6BieIm6
NwBPy4tBygWz2kQovFLsztVACmvsvTR6GEaMXFxW29f4x4OJI7YhQ1JvGNe/LoIkVgJakcf6Wkaz
L90CH+34NPLsIPasGyHgX6DPq0NRRtNJrieLbaK7fizcv357bzUqAGQlBa8uq2wAv+OwxboiwbTU
f8ezpvsLwEFfA/N0xmSnjrmMJe4q2H9boJ4GKt/1ClZOjGlqPUMFBTjHsYt4ERk5sUHiwGRi+DOB
ppgcrINodTgHE1cUKXNlSEy1om4CQTcFobxFb59s2bBllUWaCKKC2UnSo6P5xltWEA94phaq/k5/
uQ5uGLupkykowEV4DTs073ulKii7WKUpaGNuuFtBcIeCO7DhJNk0QW5v/LVgxEkZBKz9R7eyL24D
vskejyxAAE17HHkDQq+0NZHbpVeCLucn7veHANZXp7Oe33zdaNkCIE/2XS4rU4MPlMPauJz6uf32
OLi5Ex+ZexYIp89nydbQjRL9CNT0K5YsOrK6uCfDomPwfCM5W5mKsU+zeNSgOMhRwwAaYibUirKf
pVPzG7WlZrQ5xGeuTwqg10ud4wnsAc+5666wciDabwTdWBFJ16dlF1Dapn7DrsdH3m5d+0IdUZ6D
9VfdBJvDN+YVhLa7z5/C20SS/Cvm2MRuKyhyJ8SWk6OdlyNLbZVAu/KqRAqO+aCQttAPShVls7ZA
l86uiHsNY6txp3kwkUL+L3zfrh1ZuLRQ+ZoXAv4vR8L03et8lIQe+sZXvrt9FvhlLzYPcq9YaBPG
ZaMSgwC4qUGatVfhlwrKrcffUbH5QXvP52wmNSCeYRKF21m2jEB+5fzzZrWxqptMW59q63qG8xFH
5Ub6MslmFn28aZIANRB2MTlDiBq0aRPF5MWqIwQpmWgDaQ2fXto7MgRD8dl+GTzk0Zx1saTTMEmN
oX562nxIBb5qUcEDnXtfOowtrUNzMdArZjKSp/8XevdvNMU/VejsuB8onn9tDVQYBxeEPKZm+JhY
w8x6Yk7jnVUVcaoaKgY5udpgZMDTjvS2zbPKlgjsD6HaO9EKbc7pDwC1vB2Kw4pHSsWCOY44Gtgl
G1IoO4EQzW5PLG3M7KxEXY5fMJ+BjFwNGrOhcjFUgA/uTuXuqWxSqcI8MhXyi3Q88tvjjoh+Cx4Q
a29G7yTC95FAIM1tRgiXZmOEsJr0kbMCzXcsC9vR2XIgUgVsxepIkA8G7IdKNo6fVBsw2jxMVrJE
0dQKmAygSZ+azGr8ad7I77ZoFz9eu900edwlQ6SKcJlB+u9VW/kcOHe3scNrFksSVML5ARlcE2o5
hnx8RKtOIcvHlAM17ouCqyEGsZekMif78Nwq1W3/zNJRHU0yuNOnagbBjtzQ6TGhwJ5bon5fqqmF
mpj+BGtTy7YiV8eqJZxdNSK8hjDIE2SURU2vOUsaCLJ4bL3k5fXlRboXoeWbjpiyLNX/ndGS0Bx7
q9LIBUC00UR///qBuVgQAEV6E6Zgi62PlIJm2PPx8Lt0xOIA6vM/b7nP7JZ97t0upf75v2xPITc2
JYDqC/IZmGoCUceGQtuGhjSNzQTK5FSk9Z/ihDfTm0BQYqMhmrkdM6AJQQSxjXU2frjyFkJlmt0o
OM3wrBnZMhjbU1bHcTSWx1f+qSSrqNYBBfE7oPg7bxDMK2km/thvnueJlyznghmwkxxez20+exoI
HwfUfgZxdfz67mFepeSHCCO0rplSRS+4ux1UjDjzksIjg4riDdrmtf2tAXJp+JJ5AwXS9W31tqiT
gjcEW2Ihq6QXr2t/M+uP9vcNyDR/FksRM0HbZk5uz5HZLJHWCbIgAwL8QPsGAz5zzx4CVkXiWao9
THAsCHtb9fKXlyRRq9VF6lKN9ckPcHUDABmTfa6blbNS5wVu8Bz2CWMFge9E/ekQVtaKWiMuxzB0
deo61n8u1nYsFGZ+Qy79Ol4zo+6uo8zmeeDydYNPsyjrhPJJjat6c+Jld408h46ZhjH9i+eGlJGs
5ff3FrF8cuJS5cv1+jbFOR5DBcLB1+L9NCcDYHZawhytGJTivPojX7gqxxhEoc6QRsqXt8JpQWJS
LgFI66269RXBR29vQ1xK47/oZERadQ1YxpefK0MQs2xdWc+LH5WWzsZ769HVV454jp7xa3vSQImh
a+aSgfNA9Egzt/QwGm41W0CMWORPJ5WU3rdxOovs2tEbRbpQMKu8liNeUkkLxJ99r4kXI/fqeL6x
ZzqRDFsZyuT9J97s5+gS/qIVIfe6yNG72gIgeURr+W/OtVPZquesXevz6HobjtEITzjaEcmvP4MM
fQPMa8QS71ciYniy9mFjYyKYTGIuStvgSmUG8vXLqp50ZCsH6ox4hv79Lt3ZPn24/FPaBF7nZerD
5qHhQbbgt2ZALeTtxKRIAKGab4a4+IZlhUqM40fxBfQugh/FfrQqtpE8ip2cGp9OvslfZD7dnRxA
A11Qy2fntwWmIwdkUMQeMO58E9OO+cT8SYx8+fj8MAItpVjwUCE7mWRFkZ4lWs0808SORWuxfW4Y
Eh81lRgWVNmPXL6hbpTSFPhtqpkiPfS8l92ESRLCHYSkCiA1PF04hAdI0fa05NWtbWEb/iYBJTG7
nPYLNSZ5tbrW3x+Zpm+hlVs+VZG81b1goWWmgBIbS8uJrY8McpXOOLB4KYCAnlCiF0FGUpCCfgcc
hIVpDHESpECBfh+q0QL2GiitnFPZY8QY/qR43h2XYqsWZJOIMi0brr0b1e4IKjsSpu/ftWGfYPz/
a8BivM5LG2XRc3jWWm67/TGf/D3VHLTywk9V1ku+gBtuzxIc5pO+SK5T8TgO1s+9ErN4ilqYSpjS
L7R1OOkDn9gBzqBcMl1eAttUhEFJr9FDxWtSEn8KrxMW90u7G6Cqm2+K7362SqjAhvUYWJQB7e1c
C1aAa+JrQ21txKroMz57SgDnQvnYbuWXdNFbWGDcvCgThXYRswCh6QSnrtZ/5eNN5wV6ECUrcS8a
/XQudk1GOFlvEAmFrIsALFPNwsz3l4oLU98Lgi6w8t3XlplkFBUiC9O61beq7zwCZv5Bg+pxSkIA
IK3laUDxzwhwcKbY42TY57yA5HREAfstpps+MCSQuBVfKMSmz34YLKLWynlfShfSo1i6lRTLWULe
iO2ukBYKKHXsNc4g3+CenMMe8vjgj9ekodMhx/R/0VlTfC2TxosqDxu28owx7wihJnIo3QcCX71H
ixrgQ1qg/5Vw9eWxxeJf+1nW4B7tjNIfE2/yX21dPXFFrue02pASd7p/MzR/CrtLEdSs4iOAcUC+
aCNmHl6dhNHB9PL0UDTgNawyMxx/Y1CPR+eYajRRdQoBwLQObEPexn+/Oxy00wvBUQVX6dew+PXb
bbYASJhm58DcPno/BnY9RbMgUi/4eI1YQdfXOpWAIe0p4NpmzcJpN8UlPquTdDRMaIH7vShbDUud
3NIvBlhedDyiAdKfVgCN8W/qmwuuIN6b5ty7xQSH2YCFpNGDheY5sAdgjn3gNiG/xwZ2V8myOXqi
3EjZgTYxozp4qtIuVP6vYe3i56WfXzU84yCG3Akm6aD6FvyU+Edt0pZ9/Eb9g1hBvy3BXyIO4UIP
JkhtjM4bw0eoTm3JZR0/IhNPDQHqU0z0WJkj8oqBnHAG7jP6csKGMgja327xiMP50LEpCFiZgI4m
Oba4knN8cf0WjwhvJNXZtXiRaEQGe9EsLKcm53OBcmZe9VO2EZ+LHbbvpZP7XN2ihGHgKbh//Ouk
Ll3lcWOpVDNJc9B18m6cMQ2OpgAif2VsEvzfsTjru0IVVgk/EX2qIEDBwzLOljqcadm04/Ng8Wuh
yVpWc7TBHKtOhxP2w8RoI4wBqjoq5lmtLZ3gb+dB1zQXNc/fHMdUUiKYEnmPghoScaReWM/EeutU
QNex1qN7SqpLcE0vc+10XqO8kYUaYMdIkBTNAHuHwPitAkrhpGhIcasUU/yMo7m/GnXAtNkplE16
B4KaTZhGeQAvcWWW08uMsNETU1TsMMvYn9Q48V+jgl8Y3omTiO+KSRno6lVZzgvCPTFGL4XaT4dh
GNwumDuzd42WSPk7pvE182nFKFvD7rmdLuWrloAp2TI0mWHryohPiZlpodPm8/sdYCDOVB6I1A1T
c7Igrh9aRjXeO6XYmYjTHuWOxGhDWjxVCKOFJzGwLZdmklloJ+MuhhHOKNPsj43HwWAwjmRedSuZ
f6NgrUmrlLAIPalzmGVo+GugUEhea+eZPV3xx2KwcmcBKoxybjDYygvtkV8vUvv/2oWmgJz9bses
s/IHBq/GL+yr31WRTKNy5kKqeMs99elBPZT72jfMIFoZNFxTmuKj8zdYildkFaQPDYe/Kin0wM/2
uNtCS+jcj+1esjwML3/1YokPNK9gr4p2q8uxG1rKknPu32M/kanzLQsY57o+Ds2UuDfIeERmoVmI
pw4jf/osLvWl4KIjLhZPc2Kx716tCKt7KWlX00XcOgrmRP5c5A+15Vp3lPuRYAFyCN3CH9MeFdfw
P+PKSQBAlUvl8+FJaKk1JeWTh+Zy3pT0cj82jhbAOfVQunlHJX6+u229TWZ4EJ1Id6h9Ov0r4p5j
xtTnMWefQpypFe/JTDHb9MinQsiK+M84M3XGaFkPbESQlTEylsWnccHdSKRKxHYLAbVppnq6FbAH
Nn5Nn8aKv6SO/jqGja3OAOXe6xMmt17oKKnTf/pHYKa/IyQHyq1wXQ80FQol1yRlqDko+GTz7fRf
Mji0SHxMhmPlEmIwj4oG3Aic2OMfnGuLgYfORZsREDTUdYkvzkFgV293qNpquz9f0Gn6KL6UV7BR
/GCRsNpT8oEg5lJW8XaS8FDkLIG0raIkjGOL/jlUdlrQHu4CrL442uvq8raSpKJjOF6geAfbIHPg
/aWeDLhzno++IMNFulc4qYKL1FuYc/SjD+O0xa6Q+8ILMXFjeq/LID+hsvLea9DrNWFBo3CcmQEe
GPA8uKQ1y0rF5quIzS6NBx6FGfkQUOy+f7dzbxN3nfhGCLIb+a1ihy8H+X9UinYWLW+eD/qR4fD1
HrBcPMgZIkWZ/00CVtTDFEV33u3c4EUJhQA3SInpBAf5ukNZTo70500nqqcZwA9195D3p+duErr5
TzBjh8aoYy56rj45kZeKCNYQ/UB0mMWsAp8iZnZy8S62nsdOt1LpFWOaFACWCnjEGRgz0/YcskJT
/+WKhDnrLucxIDb+P2/WWNnA/5fVrMnQQ6wW4BAcrmK92X4lP433X6r9rMgfxWuvZTGUarAYAvyb
kE40UoMRAHB40h6/lmmrF3+edpNxjCGc3bUgoVyTMxYfQPN/JLF/VftoJA1c6+DU9h13aYLjy+XP
7SEAVXoThZMWbMEs1UJostDFtMXFxJgpoiyoGTjLkvF3oCABsgNif2o6CPcSLyKPSlDOuO+vinbp
6RC/1KIguvYBhmq9H8oM3GJSomeUx1IhAQvChamzdc3uXSuuC4+LT/sQ+Pu/GmAff6LmqE+G1sf3
T27gj8jwTOi2Xt9KPN7C3V+StHZJMzW97IJxKJe+rDHe7lhNbi83K6404HVpkipSrz87dvQLEnHt
fMqZ2KUhP6/VNne6pyBO8DUIIShxgD/ESjQg2gTtoHa8YAsvpX2At0Ku/NqvqtYstYe1kgAfHTou
51VM2rQjQQ+ZofupWvmsETtEDgpp2BR0RJFBAmZ7AJSnIacVtqRgdWr3m8Rg5HVLqzHIWx9Ug5GJ
jerNcmXI7jLBS3WAOWARm7bkqpmVbWvOYmXJ5w0RPWNWOykMdKimk0EtvECHuY+8Tn0F4oC4vRS5
t58Hn0fsUJNgdLoUPKVKMenQKtXmn65XPQgMEgpaW4YHb8K+aSw/2uX6kTh9Bhd3vZZJs52YahvY
eN14p1y3+r2TJFQvfOldcmi0utK9tq59lo+pMb5K/Y8GAL/SgK/pZrdAV4u9VR9z9f5RbgDEZtsq
7NW3VsfDfzuO7AZph91tddRO/Dsgv7t06d7UbcEpId2FarUs9IERmIZAWA8PPPoDvI2m8TN/LRoH
U26aXAaR/ao8RakJCHpSr4s0cP8gnS8RfGFY8tuL42RQKM5rh1al03/JIMw0F/VG20uY5uYT70/K
Kn8hl8mTywlYzlUP94s1zieiI8eljIMPg9vevVZfdLmcEumfq9a4pk6dD1+Geicbaq5Pu9FnT3pk
2Taqb4l8f5SRI3AthLeXjKB0QNnCsjCm7uMveQPL0ZDCYLFOJv3Ux8Gf40GVZ4Pq8ietIV8tE7mN
VThQDOs2xrgEoUMom1XdQ7/hjULugHvnInxLs4aVgnoIoR3aMwjOmH32l/s11kky1VZZySdOuH32
zUFcjtg93+mCaXUccruM1+kxKKrSU6vGUKhhiA0o1lH33wRVX89lDe2UM4ohPqVmTRgq1kRzuhrx
J9xPf96hVU2H9QvNBto7JTwFl+ISlAm1LdCG+sB2TtXubnMxHQHl89zOt5H2aH/VEM0eUY0WjNDB
DfxPvIiYcI6ig9ibaewPsBr4zByfBQzIKxNHcTUQu2cm7FfK6dqE7G5ITsAwSzEh5QKg70r0KsJ0
1E3afjA77iYzQWLt8+BYLNt4YPmPKGkMRjf2RQLs2BkHMQa5+f14ZrDxFH5MZWaVbFdEy5GA4S+/
aFNEeciznXZtdwEvOy9PJI7g+lqMf5FvyaGYjIlUp61RSG83rw9G08esDGYpySc7reHCXcUtSWsX
OKqQBz4FY5aaypZelPjWm5jx3G1drgS9klFs9kKpQ4ZJMTQSQvrHbZ/GpsDHWKN0D7sCb3HT5DGt
93dqCU5YRxxLTt2kSXF+W6AM/S3PhXakMPY2lfggcUAQLnloXzdN5TEUhIiFu5tlpJoDDNVmhwmw
8qnPjL6F0iP5FVjeZb6Z+9mmp4jW3+gbdotNJfwMQ/Iv6ylz5++ZdLhxUUfSl+T3VDzjhtQysxFK
kKlgWwCp4GI6fz8bH82YBS9WzObBIfCvz5+SATfPalhrqbKKOQ2cdOeefgTzGZoQ3uPKFuZiZJBv
6pq1kbrkFHzQuS0qyyy3KXNG/+iHZGIXbj5bw1l/D8+5vq75qmeF7qqDAGdh8QIAdtq8gCwmn96M
71NFNc1hiHdhhXZgXHePnLrJKzSLaArk1ogUoy3o1ou8BGld8jZoFokY3y/lNwx8jExqeSYjUKAh
AgMXu6N0xn9CPAvv/91aUjHQK7g7sYZaAVDAFZBB680ZisFhxuLKKBsjj3PvVL41s7loRg1W5fv8
9fQ7YYofQik1htJy5HWZTB+YO9IhjzuQrWJDtkJs9fqzedUfPMVTkdnrHluDU8lmNpb5vjIfO8hL
kut8rDIHYGVhR+NXByriRo3AHkK2teaziFc/FAcOUJD4Yv/9DdXf7AS0FoaxJmneFNCBwWJuebxv
kqHdn1BDbH4aC218r7LVYo+KWqa90uZHPf+pvuSKB4aKZai5tI0TnPh5/pB6z/O5z559bopfOUG+
mX4XJJrNGq1vMPHASCoD+L597D3bMPwtwMbTBsAuSxUN8oRYbNBqvRZpwx6uIKvF0VCd9u8qP9zr
KZtQQpoPuMyd2nsFxiC/iJhACvYcpzJJHrQ+n9Vhk3sUTUbsJcMeEWt/5M1j9h5Z4Lni5bGMeXSF
qDfIReMmnYgUBdhN0fUjNohuUZHr5ffhNkRBehXkkWetVZgdv5V2JsU1Gt8bnxyJHiDeJ4S9A4oO
NPZkPQqWQiwKe+6aQlsWCbp/DIhpZJpVp1v4lrmlRKDlAYSmrHK4RvKCseb51h/iVHRW+hxeKMp+
zemwNvAm5r0dWwnbHpNPXcbHRESlnlfIdZWgt4Sn882U7JYnCb2gCQTAB99IHJ3s2Vabys8nNWdE
IOSxvjq2wnEyZI/BjqRr1P2Rd7/QvbqUHTReCXy8+gcxDCl6IoPbWqfROZgkvx3iwpwM4PnQfO6U
kHrWXLrlDKIIWR4BQTA99FKUr0kduS2yOoahmS5DO+HWX6xjfpwkffe+TEm3Q+4jWJZQOFSjitoC
bY5JsxZBNC2g7miXO8cXz1QZa2rqDW4zNfP80aKldaM3N4pOShU88HvzcfBJCgDiTuN6ZeKNFgyR
w6ebGBi7o5hZMm6VfbyZFdp16ozf0yG7ghgPTqSrCIgVQSok/IPVw/lr/EkYCkaS5hx86iL87jbn
okeXYPrGsoDUg7XW1GGHHM2IgD7/Gy2Aj9RECsAb3GZjDnU2TIXUBEExUIu8tYQTrc3O0ejJs+XW
brmUaxLVAv9lj/cqdsj1gHys2nQC+EFmCfSeE1CxWE9PKo30/o9CMI+v8MwV8nA2/8PWzJgWKntG
WvPENUMNVX3dq9hSNJW1wx3FyWUau6fZpdMu3cNYuqZMOGlLByeupq3VXl0XNBYN5JHPd/6Q7xUQ
EeyRGoZ7rA1QadbTEgHu9c1Faehc4OC6WbANGWSHXB/oKoOcpR1xfNn7JoveKC8d4Rj3pur2dKXF
b3dfyE/xkv5craNWvNKqxmcmwQjxloOWmT4zKznNfwIvgAPEsgyVoqpmsP0SDkAOVjEAoZdZ5JwR
3LIFHIv2xpbHu+41WsGeqBwpWAydFtneFw1VA9lBOem2ZP1dtFBkbcM2RnPSgyZSMa8sAt/ltCMC
KyEi1fmQrhz4iD/URCP/GKB6t1fluAdDCj8Zow9+tjdmv6ZqW4hrRyM87b3D5vQW7JItE2vuen/H
NClL5SIjQRA88Z5wElZQj+rRzrrbwiPecMV9Z0//JkhftD7UjyaHe1t1SK/hl1eAr9t+iFF8RZIy
mBy8gZS2GvP7PavM352KbviRCPsIdjGZ4koAXBujY7lInKLtBKXaP3kpfWOFr1ciSerOYYdOPUYO
CGA+QuiZAR8+9+Og82Ln3evttvDbpKWeuVzOgMhNbyfsP+T0KEUJVQG1Wsi+3jA8c6rPy+KQSIgM
KMqeyZ0rWB/PuJzlHuvNQiSYkPydaPCYa/BdMfHoKWyavjiQCX9haXI+vRkN93ObKfIZLrVaE3+T
IdXUsKPGv5LM/h3AiN5oVmUM6x+Yx+YclELvVo0wczsl80HunfXp1Pt3z4n8S0u+FGwiacYBYaPo
y5k/U23Nf5u9tiqcScaAZWuRBzqsbL7eEkmhX3qnKO5L3H9RntRfpAN7bK+P0OLILwKtHI/QX3iM
RorbeNd7C1YITETu8zli9cC/9180Q0nUgXNLxC89RNdrofMBxeE7uzolLMD2jCvLdjIFH/sfFLCr
hwiah87efEnv8jPqXyvst6652SwoqH8bxrQjKy4mhDbqJlxHcXuXKRE9Ebl8Cbt4uT0lA0fKAygj
XFauKoTumsgIdEO2fq6lwmDqJepVubZaAsqUwZE0AF+HAoosZ6B7JJxcefM8Bu6s+TMPAHWcipD8
HiSl1kjvq2RJ0eeMC4ChurLADwHYN409gw339QJclos0iwww2yHRuWeqQiBUePQMRoYl2C5StiLm
tLdGOgHvqD0YO5OT+kOqHbEXrM38QxFqHdH9KT447pwlHvnGCehnHL5ihaB0y+8W7Bfhz3K69wGp
KSyhzR9YvsZAKuf3J7Xl6dDi3IOFoGn4ZKKijxopY9J+MWsCBZz7K9DkMkJ799PCRIECbw2vHJdK
fnSwlwox/EJCxL8r0aPQXbnUAUgfXTodOhHT4mcjirjeyzwkbrUvD1RcOFUkupMo6tqsbN83FYiw
xwj24jJUCRg0PQlLQGbpYnZVQolTBz1GTC05p0sF2rpRmYjdQ8Z2pweO7ksz4xlifllXDYR+pZQ7
bHm345gvJIEQOkM67379CdZI3pjslu6nkRcQ5TBQwti0etNijpjUjLfWjoIeA2N9JbxzWPX4P2rs
izMCwxj8T7Y5GbH1tSJs0aX5nstZcyuWCLr6M7IM6LTg6/1b79a0F0+dKoW8GjxFODYXuGhDnNzL
G7iTkp6R01hunNc9CyW/19+dUMR165ulXcxK5b9xpvWeLWt9/LT7/1EPYxUy957UP2SnE7bLzyfp
GDpnLvHH2uvxt0anfiZ9n3QLnQz3JA4IcPc3w63Dz63WD6zbp+Uxff5UtoPgL8AcIGblHtoy0BNL
6XLKbyPiY50tqUQbKQB/t4BHrhaqLqwgtGyToof98A4ZMQ+ecNXJG58C0i8AVNTRsjzXyCRxhTdV
qxCPhiUteV9/fUPvViP66+dFkOp+PfrnBALQgb/wHYcB6/xk+9kGrq38X5aJcuD5gT/ptqOkGjtW
w6G3+PVWD+Hzay426LCD14i6vSykPWspoiN6IulBH18xxHMDDaWhHonaafKggwIZJjieBgRYbZsz
BIJa14Q2BUjSShgOGavoRtyhTKn08q29wbKwpAwda8xx+Zpt4yUzmVnY4xJAeTXpRHuZ9RCbnLVj
+3pB2KN43wImQ4YH6UIE+cRQzUoK65jP69Xo1Lot1mvfUqisX3ouYOQrXfadXtgsz7gUUyUuQQHw
9XIWp8Em0C1SNgRDvIA5LSIWzBr4OekPsCsR39LMMVAAxuQhWQYOzm5yurW/55eM6BKMGJvkGxCY
apv/HzqKMngI2zwS2lPQGdQtms1wtElypBrexnzpCoOLXq2t6as5wa3ukg8Lj8+rD2qErP8S5QV7
c0HUENF5enMt5xmGy0A354qLMAgH000tatyVtDyyb/mtjpzcZCE4cIbWHByM7RGd145AxFUaHiu0
+rUNvm/qhceVZhREjWtFPZbe8XeiL8OwfeeEWzdiw2SVmaVId96fxzOo1onLC9gstac5Ujrz/NYJ
xw/5fuobnFmF718pu47/EdLXT2KncWuyeFbq+qmWDYIDVDh8w7frVKMzQkekJ93J2auWf+FqXnFA
mZ7dEUfy/yCu+um4zSpkJr/ViPbQAsDrkmWlR6qHZwFcXLMs/w0UkouC09OuxnGrlCu7fYc15QXf
0COJRZc0bIX7CpGNaU14KeQp35QoLPcsJ86eOkM0qq+g63hPSERRlyoP5lk09YU/HGj49fZq+Q23
rwdqGPuxZXhw4vgssYRXsen8DfZos1ODbZdjNLhiyNn3Tl1GZO2MDAHnfxxMCXVVe22YBjVTHY36
bq+KAIYF3EX+tUinUShjxjCGTXNQgyP7N8oKpu2Nn8tijjWPaWbazHLK3Wo6AsCaPUvGuFKJgPOb
CWCuTjfh6Nic5SThqNA8X1L91CZ4xPKl55eRc5dC2GXrQN1Blr4i6m3r1YkGMaUQmCi36Cejizvl
H3pvCT+kc4s6yIAk87eob6jGLfUSuCM81FNOtRA1FEDD6R7w7qexNgRNG+UVxDf6W8lBcx13C1DO
LSV0EHYypG1WakuK/QKWPe4rkujFTI9qW8D6CJvDi7AFC0Lvv22rHylZzAg+sfBavfBPYSvgHAPG
Ofz+xDxBV54ZWWhzEKHseYzvbkf6p3bsrTeQ9uppgSEqMiLwJsRJLcNe1b73GUphu4GLD0jgsmQJ
Up3J9j54HxrWRewir4Z6f0GAsD7RDQ09fgYbaOFBEkHLlys4xpxF80JlY4hRRWDUzwGQEIH2n7PM
AankuOcxEuP3VwQZQVrPtzUltg7Eab6krbkij6/USsYY3DgiDo3gIISFTrVz2Nvrj0b7ugyfUCaf
XFjJ17DzxDjufGl8hQTWngDHRXmfAJnTHQW/oxyz/PK9T+dVH4WmnrDLJt77P2im1+3eTkDxIs9o
WcSDFy74C2wIEwiqLuJ+7UMZCyJtT1HccvOwkMkk5y+pf1yXOt7yJLt3j3sSgVXOId6LXewQD0sK
VN6nEXH6EGxs4eUuKZR6X5qPvJesjkGwXaZ5S7NCUHVbpIOvkG7FkkFoF3CsYhObqxunryeGVO7b
/GrcIQMQ84BFpg2/AxJPEcfRwJZRbIHBrNOHc2UcVA69jQtNpAgJjBUixLWsAg/JKgOW3GlkTfSu
NFTIbi8oPNQHsxW5xxFImF+zMY+Klpu/ODd0m4WPSU9yS/+S9Zoo49rHVbgQKBY3rV11FUmTLEaD
bmbSmD3ggDOA2xJH/bWeDaoi5RsV/l0Z5jozH14h1g1GS+mcxR6g71Zgiees0AFiKIqZ3W67ZAtZ
u/e0mVNhMI0+6QtCjcB/G37DM1GZE/0qcSZCk0sUYhoVYONMxFfTm8HAtZNCjzT89DwA+Y6R7Owd
r0pDgIJIHG+KR17o9UPPdEM7mTpK3DNAMisUJNZa6sAebmLR3rb/tIWVIuFVPk5vUh+C/nox1Hg6
oui4+mgDA87iDY5Gw8GRyf3iDGFjfBNZ1abcaAht/wlvVOTgf1QGLWU/kq7i5AJA4IivtfiLZ1ix
Ucc3/VbzZ0u8nGHd8lTR+F9+bjAFNLzSe50crUzOt47LV3Hkc6fmOSWeuNzXvz5lY6ckJuo0OmGJ
BcBVpe/McjIjTjJNN3VfQSxf3qe8f1bzVZ2kSR53oHRnW4ZjB2b+Cu3qmhN6LROFCd7S7aQmBceV
vz33RSjju3627kXSMfa1bEWiF7Ix4Dqf3cZcVQ4aHTFPnSTElmL8/OKU6dQWk73f2IP+1iAoxLGo
mOYRqOIG0WwORCxUeXlsky4vdMzQq+xc0tyoUGfNA+umB/KOWpKPCAcRStFfk0XWp3lVgo57g3hW
sdSrT470q54hjbBFsu1zvlz7cc1qtyhwB/0aLc9uM+2FGZxi8SF2UPYyCdoI+rV10ISF9UvD5jRw
+1LGtb05TVqPXJi1m8FwNsR9r+x3QgHuydE2dmpls5ZP2hPdd9Xa91Jo3jYraerxOSimpjF96krT
Y2jZs5DCI4ZG+QmeZm5ePdRXN9/IhADFefcWp5WLZli7VAoBwZ7KwN03BsebVVnjgLtRKjsKKi96
GLUDKUWCYPLbKyxpYAUUX0uXVE1he7AE3hzc6JKpG/Lf5q73fSyGphhYo9m6DdZFErsEx7knp9bb
G4eS0XyWwqfMYAj9XuEN52Hbm4PsMoR+r0V9ephTsKxT67yKAYJeDCUY9Wu5Y+O1zlRq3fSUNOvt
3cHMS/98mkzXiCRJAmlspmuaINRarfosrmFQ39OmZq389Gpb9rukGRYW10mG1ueVpSjl3pvckiPX
VkRWgmCH3wxyufHQZqIA56MbBlWTgIH1Ieort9+12vG8d3Q/DOkKy9X/89l6Y6kz6JSqqvPNZPN3
uH1ageI5VFpsVFWezh2ReGFSy0/G9dYY278k8lQEIdhQ1/1gfegx9qQIt9PN5K13XJgtnhcjOPFo
BHYJE9fuX7hW+K0s/5+0bU5hzRH5t3bZdWi7UEukrhGvBD8FKjbnhzSRrs5JRJ5c8kcNg1vHSfSv
pG8cuAEwQl1SfonvOfRfiSJyXyRBPGaFk+K/BKaY7Hg9marJlPq7x+TJovs5NivOCtd4x0J1rXE+
zZPzXAZDfNcmQ2GoYI34kXvRizsteUhqykMaWHO3p4tdCDXXju6CeDJNCoM8c60yPdx2OShe2ozU
2nUp+CoI26rrMBg7t8tVyOXejD/FO+znwaw9ryawkstqax4VjvzrNgh1Uxwxn3d90FrTVXoOsHkd
Ew6sbKwfrINAxD/X3CWVpj9NSRrzYSLQ8HaWLIGuKGgzJHhz2PoUp0MI/9rUEYq6zPRIwBTN11X5
a7qY5z5F7v89fOu8a3RUaFCthBob1p7rCWeFBNgN++EtUdVgIv48+ZL3wrInEc9m/LPAyc880cIf
ZQjE6EncaRHsXdsbuAcbpkOWI5J8D73umE9KhOsU6mvSFbdF79CTIgMJx4ceEzx5XVCkmPeOJAcQ
hULIrx3JL6k50qI5QiilVMvZMvM8RD33sqyRSBnn0bFuHmjYL6ai3+iq9lYpDzoDtOtysMTGk8UD
KVd5cpHiTgRLeM7w2Bs61e7ADQO6V62ioaSMtdw+yx6VLt5Q0pbB144bKmwgpkDcCBbrNO10qMTr
M1sSq32AsLGznE+U5enKEybUMpyF+m0O8oAW2Wjp+4kLsCRcGs+blV712RfaEqnSd+Yy871KgHph
SGCjMSlsbRrHQnSasLsLim306BxkjRxfobWcf/jGP5BUjfOFLj/1O4YLP2wXr9ctUPaa5JVpsZI5
fb90pFjfAevj/pIdUFx9kPtJhnw2SBFYT25y+DVFogX6T4SnqN+QzAL9IFYKt41Tv1xyYK12t2oP
TpvpmKxdWknErdvw7OV+Gcd0+uih64MbMObVyhMJVZZ7D7u8JrPik5c8U0VaHJN7iRrE9BRWnK64
F2GwvkY5aHU9oVBP1DEbQF7rqnE/XS2de+U5v+lcBnUfAdtFRb7Oh5elTY6b+0zgqVcbb6zFtRTW
ZADldtRKEsFxM8xxqemsN8ADhkHrWnRDfjmkbd+qU/wPu4kG0LrwzkbEex3zLIvYSdZGPba62CMT
qW5U1vZNQ3SWszQjDNO4+CLfd8kWvTjzY8xiSCiFq2m6IMAuvoCeOTutI5eZHLi3FPu0iFD802e6
od87kPjqq4LNWzrAytwiag58Xr0Ep6gXnS6RIaUuSmmSDgrtEkCH2KDr5l6CxPxqgkBCLzcmcmQ5
QVbFRcrnc7ghyYLcGfVfHcm75hqjHQRJe4irHMXRasA+YcfdDeGTIjiMGf58/0cyJdTao8dQ7KIi
tPsLCcDClvWlkBQrL7ntjLOcS6wBnVjwxhSomR8tAZbXdB8WlVGGcd7nfx7z8WkLvcQN5P/hzqFP
66AMWpas34yDrC1507rtjDevALg/LxhHhzWiipZ7OJOwZaSLbMhsSnkGDAhToAqz1zMFqfYu+KR6
uCpwhNhvaJm1V4pLMuIq5wkPvU9eYzuBamfxV7QRWmWOmc/j9vJUgpFwgxv8SBllRGxfvMbRPDUO
PRrRRR8uHKQgBq6Axe5gJivZtQOcPH9/+EucV6ECcwdzDHyNijRYEaG3uNWoZ91upgqB+T021mtj
hugSS96FfwNdetzSyr/tlxxQVh/ntzQHQW1cOUnlkFiBd9n6XoNLK9vxxXv+XfGi11qfIp0YhRZG
PPspaT2t1+0TWfxyG6bAtrXEOnPAzy87nyVt/IT7qyaBPvYPjaQE16doeCNeWXTmjbHOHjwfYuY7
2TFDdAOnJyfJ16//Nx+aQNAwwcRadXXKCN4KSThXZ78H0FKocBvaMr5v1O7H1PXKNxHFXc1Dtr7K
lL4IaBemTqMkbM86SC9pVRepEWHUanhflmaFQTovXRacC3jVX3CsXpxH0DiymskbVNrQ1AKAUxVv
e0iO8F/8cJEPtOMrg2lXDLEfSrb3iAtVViuyak3fk2w/awpwO/2tw7eWoG+sQRd3HGmx8n5FHJK4
0gu22RlvoVWybwA+IHcxWLK5naph0pZq0fnh1MBa1sqKKlaI8jSPaGMZ1DtiGlWt5i2cIlIN/knM
AiX+UmOiD7RDKv6a/8RCEKwKSkdOkT2xQ1u2L7Tf+7YaTAJlQVsF9rvoLyfcYP3a/FpVsL/xxBRB
UI9cH53qHPDtLhQWxlMl5/8Uk5HED33bn+qQZGEuDhO+LFZCc61QRmLu7YeoZa0awyy9WV7ICutF
EULZdZGVCt7TtWrcYl7EHtewVY4MyEYtXNzL7HKMpJ0EQ0EUhx05pdQuFo9SynsXPozB3ZeISD/0
nxj74rhXY53sD8xqk5tsMQQ1OOr47cf0enXsvC0q/8hZOs+zRMzyHAXkXr60HcpSEhvvkoJmHShs
33tfF1+QDSGZBBreB1l1Jh9lleVjhgw/InkuT/H3kWkIjnKl3nD/gGpbeXpN8ug40cp8UVa3F6ys
p2iu89M5qb1OXUZJskoK6zNcYP8k0EWw0aRJgkl2F9+l3/zGEP0T94/NyD3VB0/Rh6r4G9vlw7MF
kRFB7Huj5/2DjWcofLB120T/yu+1EndiZdp3OBP0/4mRAIWpj4qRbiAYbbpJH1LEhBga5gDj35uF
11qg4W7WkoCix8HSSc2EXNhvYIpXC+UOxWS0T9HsLtIDjguTc5zEdAJgD8kQvPsWvxcx36eD5Xcz
H2SyYsCbE+gkpVnMtStIJOgtq9fA77Vy7D9KT0mzDS5lPLQaayjuVckGNXXsvcn45X4q9spg1WoF
G6fhAiFR4ntIXoX/qqGijNa53E3vGyX/JNDJ2AivW2WBrFNXCO5azdKZFJB7W5CFVl0bWz1U5qIK
Zq4qL4fCM7I92mDycavn2Dgi2VeHPexFEEjVfS8+jgi86D2Spmx1IxcWr6mldD4lml8VlfTKjF0m
IzdEzM+OJC6RBUK0w7/tDfxRgXfiJ/nIDk9xjyyvt/oGjVqkRa2pGvy3AsxtQpIfOYW/pMnLuRKV
ymDoMD0sv8y4uodqCelZotQk1x1iDYa97bmGg5bDIvKjI3CNc+p1vxXVAHd5BHUpya1efoM1azeT
yUKhYO7qTqtloHKXuE01AfD8iYmsiNWCpzVOr9KDw+qvnD7kpg6zc7Hqbc23TuVj9XD8V/yyvyAR
z+QXAnENKSqJtpgqjc6qwsve53m8YYCLyKNBnR+agk3x4K6/1mFXnY089cVJHrQqyTcZL1wgYCi3
kNFUhzRTnXY2vRjP6SlkdMFPbG+mCUgK6rXqM4ybLWSUU6bNd/7zNVERXiaFU4o/OtW1+/0BfZ3O
adC0vr1NriZ0htvOrWcEzr1+zzB/hbHybIfAfOn+VFCt05gK4leBkunjp7TRF8gchFL/zfvHQX9i
O9iZo+cvHV6mO1BqIbhAbfsdF88S7MJfiB0dx4nTmzSPPGFlnMn1VEkJEZNHnOdAc1h3tdr3MMFQ
9QYD176c4R982Aw0rFeQOSID9e/wFvjZAnlGcMjaCdSfQdNwpMVPH/Tzvg9JEMOB7osRGOKmFMZi
CDVSZWdkLl7qLtEOkOPO7MsmmMcoq1eN0JB2vEifBSBJRp8VwZSocPiI5Y9gd282OblDUXwUiIxn
kbCgGlEF2znyHkjPipVPSkg526vhrojeWSHX57GQG0/Nquf9ZQICL1eVw18rN8UnxF/vNtwRfEFk
Cz0G+WWRt/b3pvoN5yWipi7Z6D03iFQURMXmHjZaguDwqA7Dml1Oxbs0Wz5E4s8M49WZANDrs+NU
KPqcLpJ9a3uXGcLcvnGZPP8h0hEyA1YZUjvB3seCVjeZkUPmPdwiWowpDjX3nCI4q3CAUOFFpel4
9N7h/jN/h2qbbRjZwJyW53RPqVo/Xt1kcU7LIKIATZIdw9EecFaNg5b/QDCnlWVrlFupBjmPBR/1
NfgYNxuf7e4KOdwGhOc2tl2BE4BckPRAzw4yJPsL9vYjJvavVnFCYxAA6bjXH5t3p4vn0GgscnZK
rq0L9fXDwgw6T6/43WwCq1nk721zQPxXKPJsNyw39CmMjQVcmkTkQxwIKU1yhp68GETr+bGG4vDC
5JhMip7LHmXCIAhjwY3krP/vfJ1M2WWUWFsLoVuFNBB/dg/wo5RsF5+NVRxJgLsso67y14tnEEFa
yCPPRQ5ecNt7djg0gtwaOxInpJHoYNuLiXWbRUXSVr52GpZp4ouoHgPUhh0pvtCYoVLSNg08cEYZ
jQR9RwJBCAig2dP16O86NQVP5MkYbVsFTX2bF5bfhmJ6ir0YgbVXHNDJHbiIgxCqnkp/1SREtD67
rdtaYxcm1yJMF4oyxErN+bhjy+eFzBvosYALatR+4XuQpN1bFIVNoZPT2pbexZ58wSZXOIpBfhRP
rx7+V8Eke5Bd+bccGemV9IgLC+YT0ZAjiSe8ng6DmVEP5/wQ/633T3guZiWmn5u5Rfz81OQvj5Hq
QUQxAO0D4hWQpwerePsKZdfM5U3MdhDnLSLT0oyJ3WavhXFIFkkx7vid12pFKw1vfGAC9z2SI5pl
0gZxVBAHB/xqaVOnKg2jZgVBS1rOCX2GcUFR/oncmCSoHd9fLWq05j1uGCDo1vQi0PMl3ZDIghyO
/pYO85TVurd9QKPQry+WPVg2K999DtZC3Ejxmi60tuu8auIIEryMrxyu5OqoeIDUFFGgYMsUO2Ax
AkEUDTql1DjObpTYN56jtk21w5b0HRH4lgF1O3fVZQO0PubV1pJv+xRX8BeK7XYZNCFo7833m5b9
MuZw/p49tAGDeWHarEFlvXYO/KuG8suTDyOxDKNki/9wXnQM4UncdBzPOBgeyMZ9zPfwLBOA1/ZX
cGFc3GeEyiv6hoYkiDOCR/CCDDU3ElkFKJe8rqWPwi+ueD0vLhYA0w3niAqbRT0ls45mtm/Fsv6m
JUMJF+R+7thDtHJWwOUJV8fZnUGK0BzZr+AP3Au1AjPVG1ntT0kKrwTqdSQpt59aSUmcMgIt/Z2P
ACnSORXUp3zQJlFzIKsDD4sBztIzAWykyD3Y6zMtkr4Ft6dUQzgB+GQQyvG83RWzniJb33GCPRhP
CrpTdAzBIADW8ZkCPrOF99Z1d79M7DXiDgzlHqnHS7FA8yoSvtJBt1XBfn0Y7owf/g6uFbD5whaG
0I/1eYi5MSG2tEI238E0OJEQR2XV/hq7zzNU+hw+4GtggIBG7JqKUIXm2NFPTSigjmg5GUrEAEId
fb/otamW8g6Ka1A1zaRVB0u92r0Hz5S+nPpcwcTrgXos15bWVUR/IGb31WU4L7zKZXpTPXQZe6SQ
t4TB+bQ6c9shLbWf/NzJOKNKrAmKWku1pGQWFhC56SKaxFmhTmOiSTF7dhnjUtJexsd7ka4Osgvg
nMPqt6uh1sRMQAF9lVtOiFqUbJk2mrCGQfNXyZu1xVgD9dUBojmYByds1BxfwnOPq8UXpVuve8sw
BL976aob/XSse57vQlDKqiXVSzYYuRq2cKg86XFAFwGkRH0lvQ00oN591N3Z5QHoRA2Jb6IihgK/
Oq/sXr9y9RntM1AXm4JAauW3xb1QHBLjT7UaOuustlKbs0t2q5VA9/IEfyuksjm89I6aB9iOGEBx
9uC61kFYguP9XGQwybU4vKLF1MWP9/A1YIc4yeDQeajk/YC4C1ml6TZvPl6H2hBGzvsg+8Wf+8sm
cSxKOrYcHorwjvFfIxjtRRWgqG2XpwRpmo3uX0bBqmj3jxVLeQtbU7Ff5M+hybZFA8GyRQBMP9iQ
Q1eu/0NPVcaxiWNvUOqz9b5T7Q3aGmMHIf41qU0fUT1HR664CdFxqyHj7hl2rgz4JdTozh/JJlgj
JB2UZAXf/ffFRaDRsvEl9mOH0PeN+jPW3vwSLPcMEzsAPH4An5OkQsmPAwC4/zH5qWNBQt4XdWSv
eLbwB/ryGREE8zCxUA69e/A3ImrdT+N+UNV4d1NvNS/mr8mkhTwJuW/9LuNHQ92zXTFGx2f0Ryks
c+XSMTTWZ5C8uqGCoQ9Z3s5XxfcFL3WemAIzlz6Gi3O4MZjhjgWy5qMPtiJy00+1HHAoKafECQs/
e+vK1XkCHms3L9sgHQ4cn8wUBBzQz9Vy6WVfC/h+OYjVPWq77trD9MemIJmYHMmHd4HzzFdpbErH
xDNWREENVJQ6wkFY5HRPQREHIJNZvwJBkI7IktpIb2UmiQdIKk0Qsk0/SU1Ooh0kHgo1QDYlZat/
KLL7+5IlXvosyH07trGA3SXb3jzyfZfEsxhaSfkogyEzr0VxDOM1ikUJ7epnJ0aAzCb6uoann+sH
q+H/xA05JJE+JSrX0bFnXIzUe0w3sfasLWTnPPh+08mVMXH+dwYhnZn7CX0pg4Eyi3+ivaOf2KBH
EOTshdxI4J/RQoOmIfHoYVdZZuxd1AB14QqoVSG0d4zYttHExkw0FD3Vz6mzhINga6jjaHW1s8y3
9AjK03ga6nIxvt/YbRW4XntvGIkzLy+NCCgi3izzJzKhJfg7JOh/14HVOt4QgEFWZ/e5P69wbdd/
IWkZBtN3s48HHqixeKaoJVcwz5b2oZ8BVexUKyit09ldIn+S9I358noK+cnBMH8KcOZ0OsoayTme
7tQN1rdFSDfkX+zzLxmtXcVegSby4BeVw6ogqmTPdLTXA4Z9aUtfz9qkx5dKN9imuKG97SDC1NUj
zB8VrD12iKe+bZe8mSKu22C91+YJSPWG+8ccIIDPBsS7gaj1YrqGsOd83FA0YujXOwhJjKJAtKP5
vLxjmAu5Jh2lTYBKbWGMEHgrKuDfZ1nh5zAYFkYcwsWoObpwabj8EDcrRuAgE/7Z3VB4MAOI9V1j
+EcqOrK5ZeMJl8W6ML4C0A17ll8qxENXepz+A3f2uSQVWh/HEBLllyo95a5GyIPP2g1JqSEv6WTA
76l+9fT4h7aLD/jZLRuMT6T7WbdIuHnUJcmxjX+n1XJMwYUYIbRCymAz2dyzEZmSy7pN45Btrqgn
PRPAoaXXphILUrXpEP1YUglpmAmYsdGYACg2fbCVglnz7Fwp7ofQq3PMz6b4nUk7my/MKzUp78hF
ntvE8RVB62YRqBfD6OQeEhbj7RIv0Jrhe87JKVnvUWKTqUZToCcX2XgVN5XCPIBa8pjhprnaOGL1
OcoYPrn4DQyRGCQXLu5x17SnatLhEQ2IFzRsNRIFbTQC9VRxnp+Ci/Ul8zDyka1NNhVahNJ0q+DU
7QpU+hiSKh7P8TasLKmp2zSRWd3gGoBuG/ZrjaaqXlok8nfe+7icTa0TS654O95sxabWIvh5zSzS
AbzbhDOD0ollM2yNzPAQwF+Q+iAbEaG1HWXd6CtkMdiyV7+PllrmDmhWjnzAwRbS82khbvNyJUZU
rQ+Xe+yaLv2m2mXS90fwb7KVIWJ9K1g5ldiMMs+3pnGdXNTS0qWNR9vXlYvEcUe4PGRJBU656f6P
9JgWSHPKAmd5EIBe7/mjHIiwbp5OrkVdUXM4FPgi+tjFLfsinMVBiNGuNfjnL3lSeQvqhl82GcIR
3MJRrcbxpH2Obqd7B6KKO6P2dgelr5fSOWCfapdTc6xx9dGlBlRj1B9HB985gXApzlkLcOrU4uwU
ntSkqdlPPWqYgcd3CucS19VMtXjPzrohQJfNOqrtO0eez2TehW8xQmFLjHxybqxvxiSrd89EPt3P
zeIjG6hcDZ+ttm4d9xF5iaF2sjTN0aDciiMaG9GudyQilBcU5poupPOLX253dbvyg+VCiSXspav1
0DBVE3Dhrdve3+DoZ72S/CwBE6J6N7qsCeJI2LyMTGgbGAwr2chvZmverURUej/VYS6NjjBJm3J8
Jg9djFrjlPLDcemu6CQOAiwlUPkTrP6skziS9E87hYbr7NjWV6ZiH3NH8ahdmZF2DKzLy2PO4PKE
O9tRHDNAACGEToFU5nWqRvEU9KL8+pxjuHv9G965BsZswNXzbP8eZQ0wgZmc6fOx83vTrmDNPwup
TOksk7k9K3Ff1rCFw3fTt6HaM7RegD+ObygoqOxATCiGZATnkmVsSD2b7OJjhBKRfixbfvtoyhgS
XieIWfu+MmXwrwWf4XH64Gq1GgQBtQs/JunO1pq5keOFDbtP/FxgWFyjHcMQ6oqFis8T99RzAszv
PQlqHtBF9hyF7nb0YUUUQ1JJcAIKrZjUNYNWntMSCWoGXLEpQgHOGTrRFLmZ/Vv5L+CeMOVzpNDH
DxUz5ESLtOi9SklpAfjaHSqqA8l7569xDzftALfJleDR5GbidS3EJb/8JrVEyimn5i6YkMAc4qtE
US/D7oHlgCRn5SBvWxHMvv0Cw39bMN1ECeJ8caZf9w4nGxi6w237aSQV4KazOkzkKLR5cYGp1Dm9
fiO1YA96rRqul4rh8m6g35p24soPcwCJhYw6KC8Ujd7dU2ZYm96RxS4s5G2RfhmVtm3WNgBrZwCn
FhrC50jCVjfkCyAzCI/SwyPDGar8YwwVK+V087dGWeMyuhwulViGvJNM4ZZ4BYvaYIbCR8CTq6T6
jDTBycHqDgou4Bv2aocwJmGnZFNvgz1SSvu5iWK1CBnHA8O4uRykqbmTplJX6jWGTUk0FDijN4Ag
d9Ak3tRLrxNX99x1KfKeV5yefxc5ICx0RUyiKgsYgdDXysM5mYI5+I9KDheVSgoJ6xyAKm9AHSXv
IsJblDK/0ws30c416ciqvZqF3iWvDt6uE/FmoSEvyfF0NB1YZiDngZuCkgyr6MjQMyu1sJJlEqrn
I8pEeILqnkIMh5O5LzyUopwa2t5bzHe2B7ZibngUS3v7NgY1EEBP6znW4hhxspYs0VCgWYlrcJf0
DkiIY6g9Orqw2FEgghYdaBOBznjx95W4Obx0i9bkHo6YqtzpRIpkiSZn52iklW4FQEE8qB5R44K/
s8D4VxvP1oWMPLeCGQPqIeStIQT3gU//Hrv00/jhA4L+oKQDDCnkJJme9/QcJQdFvoVdH5Rtagcq
KddXj+7PLVy4ZaBCappRrY20OpPpI0OyPVtxqp+5axNLSTKtArcZGRunN6GC/QSNQt0XRBFaVPGz
96fIcSVaCT6MqnDiasJwhnC61Ba5T3MRipAqv07DAjYeXCFosYb6utCDxq32UNMQJd8UeYHCk1Ci
q+SuI1YljJBQs3uMWZg8TdOVJXekJNc+S8h08U2LXoZG0ZQEJzPDTfhdKQfmp/OHwtpLilYHhE8W
b/i4dgfZoBIM9AKo5Fkz6okT/KaJB6N3Ir5w7yjGmU12I7o+qdrsOGnn8sBFwm5qwsUecfonGJ66
1IF42RZcdVsZb7d2EVUuTHmkf482PvOAxy3frQYf576ZHZgjrQC+oOsDO/998KhyARGmFFjlVhcr
rAokW9bbTB3rJWwpe+sMX7uFrvWr0b3h67g+DkJfn7o8Cb8TPa4TluzKkAkzgHxHp5ZsHiEJL0mm
SK0b/elfl9XzXikPU9P69C9lqvu+ZJX+NqbZ5lSbT7DUiHNUIsEYlErPso5SPCdIntKf6k9xl6Iz
8Jri7ctHE57Z6CR50zWjSUOa7Bah7ERzroURwAIdiDBFPpqhxWekkcukcOaEyIvjykiptgEf2sHU
LpnPY56XI3uQ3NfrtFgck+KPJ0ppC/ypE1jNFi4PyjCrj7sNYJiTVDPSn2famXcOLpyV/s5qfjLr
Jn6XC7UauIoSJ6Ak5TiJ7R7HExPYzxAjwPWbL+2FFYYmUMj2PKI2ETdNz4OZ283KvsOz1+cfgfy1
NOcsf/6zx2VoERcuxb/hCRqA66SSvWAG0aK4X6c0V4j2ZW67rLdyKCZ1Ep6baaEKxeFNOcY1jAGY
k2Tjm9uycbcvJnj7+RljI0QixgEAdQArrxYanu9ge0g8vvBC1DZhXWYW/l6Lf7miNJ1tyAxNqH8n
4a8VMlqFOpw5VqyytPV1D+gCuy8XKHcS/Q8KE4ciPiFcG6BodXdfViLIJpt1DUeqWlvP3PDOpqN2
fzNZrE4Hyb65N6qD0BVjae5Swgc6gVDW37YiD38iEjwZ32Bqj+k8SdpcWsmypRJH9WEWOsAfil8t
KP4EVijEHR5SJ/0r8iDlkE4MpMqeHWRapCd67fZbfF+KnwM/4HmkYsFsIzD7aVz9FyA44Q+ufDM7
P5Y1hJ7j+660HvFrsfWwCKAUqQNgeNaSJbbcJgI4EyW7XHrQXNpMStN1SpxU4pH4QPshY8NyRTIJ
3hajPnvSqf4TIemFWY1vewNnw8zPJjjh8sTZPuxfAjLu8ejQH0wthgQAH4e6AAnRJ5F8mTMyrr99
tECUVIPnoDFtk4+EoasR62LwpSDI7p9B8U14iZu5N28OGfgNwMeRu6HMQ/jX5+d3xywfgk5zJe9L
Sfvf9QGu/TRu19jUHIauP1qpYCaXxfzjQbGrTeh0uOh5vlVoQqX6mnx3s9DXS/YAegfQrX+Djao+
VD7IiMqWHOlxK/HSXroHMwmWcH2FeeGFb8NU9rFlgYYs7aN4HbF0r9vFTg3qgz0d+3uhiAU1M4Hh
5kS7hSXqMacyVsJzgi6V2laTUPIDFSWvROfyURUhxRm/bgvjvo8cvVmmH7ySasQ3pXao+eqjAmgU
fYT/eEaCscIs74ssZw8clMAQQx7JkgiE9H9LV2UObAszggHlXitTSYhY7ZDotsUxB+P7rBX5gc7q
2rodRZlspzgPIv3glHqg3hAKB2iAZCwQdONCBUIbRJf0s4NmtTW0ERyTueyV1iqEvhnEaV5r4Hj3
76K/aM1SEb3/BLTVVjDL5FNEj1BazTKJYBLy8hKq83Y4aRgO/B5b1EmYeqxwr7LUU2or61eNQdaj
+bi8c7s2/1aIu6qW5BmNol90nF+l76YEPAiUlL5O
`protect end_protected
