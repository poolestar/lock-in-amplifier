`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
jeN9kBVWeZmJ9XOrLt5doMZhfkNE0hibaag5IsZny7wcSCbHzHmCrccr3rYXU0YpvMF4Hh1BBxB4
qEjIsd8Qug==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
LwFgAK9zAx2XBnmXZBbJMir0Ce+0RlPtWeodO23ubQTVvXh9vIIkmwXz2vZHwYBR36ttM0GnDJNI
gNKH5GdFTduCq7Ij5O7pD/bf1JGozotHDQiXdBT8okYbBbUMfiOYTK7DBhY/9m4BJVzzleNak+v2
7KY0iTRNNbAJppipwY4=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
1A6R7yh4xVuKpZLi7FbnhpjcGtQzhrKHw5usVtsuh8w5wqraSqWIq4JdsNUwuJbdDVU9+iJ/XCxe
CmLvrILhqsFDMNzCMh/u0KSAuwHr5z2VlTLfiwobomEki5o1gpNcRSHiVdL8UAdLx8r+NFpZmTDW
oZUZVB2BTRZdAeK6ZaA=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FvgKmauwQ6gQmSHzCBPMYwkdBkEK9mNkHSLmBTD9+GioqizgHG8NC3d4JFMXKgujGOLfXViq7MTz
NtF1fxgnA7qnWbO+x3kiXjQoNTfv4Oj9v+6J5gws2FauLayTLBlxIthSpTRXE/uVhq/JHUBDD9tP
Y7i/+OO8PUzo8co4OpJhZ/GRtF/QyVO5kyKgyfwYBcWmefeS+u0amYvxbtMwazFbwIGYjuPiyYiy
9Ai8qPv3k5PQF+mLABkosQRseGZySnDYcP/BNMM5mS2+aLXHOc8q2V/tTEWCzchiyEUWoVhi5jKw
LwBg3j47HFzzaNQ4/4qrgU33vYFmgB4x35A4dw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MEh5lfgaayixZWnkLFgtpYfxyUgCkjB+PiTS+xnnvbarCN4QcJAU0RHvKrTHcpXBTFiYDiljwqL2
5SAlSCoH8rMhdDOnu0MaekySCSI03TlTapiHS2r6ERxbI9XHw/ttTWFfwmsYjIaSCfmd7ffLq4BC
1fsulyAzhY29sMXeVjR2A9x2/hwLHgzmDyULy43LV54MAk/SKeRoannrh0KU3pUw8A2lZYx8Z94o
c5B4//wV/TuJXubjEJeH0eSRhzSp7GqyjhARvpaSiejiz2HAjqdFo7TDBsIhgi/poN5PHVdyoSI6
zw5ouOkmYCThT7/ioybtgFYweTIsC0WWFtDdeQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rr6p8CbdDU+FXi5rG+oDWTUK8K6+hgThbFH8XWrq7DZIXLkN0H3iGOuutQ2/B8Dnnm/S/WvD90eX
hNZvjMvroenj9JfGyBVsjMUbQefjcGs61bkKiB5Hn09ua0krokb3UjfLBImpPSnARmaQScdOImvu
J3BRHM/8F9XTdHLsZ1hYZ8AI1tpBP/fPhmysNKN42ukKjxRqICWug/B1tF/sTzqFJQsCmoNu9I4P
g39F/06VR7uvliAc+0M9TGxi7fQSllRykt8/j4qHyWqaY8q3x59uC5M5aKmes5Gxexnqw9UG7JuK
+AkmfUUM5CaegDf7Jw5NgtOKXScxjVGKYbWXlQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 214080)
`protect data_block
ndKclwschcjg2Ybomj4OhNT3PyDo06Xw4QbbUHr60fgr3CI9IBfvF9gNVl7FM1o6jThY8Q4oeG9M
40RkzEZ/DIOjrN3caNoKTtBckM8E78GLJKE2cnCQn3wXD8dv8EzS5ZX85iMAEO5tnU1a5+fedRtw
A6WZlsZidGU+hG/iFlGFOXRpru+/C84+BYCSi4m24MJ7I5bSiXRavWBxKG6LsWk3zfyO5JPewEx0
/B/jG0hzBDMGbY/d+q4ujnSB2eyYbmGL4AF5SPk4eMTwL4nSENQHJcV62rhTunggsLKWnHz1f3z3
1vQa/bxW2ReMCZ77OCG9oc7nFafyCU0or/uC/9C0HjjCkoxZWNyI3g9SKuYnjZXsxkvojX+KekKj
2tCwMiROFMHolEcXy+PhQ3mnvo/5sWQtQ856d/o9l28fecqrKzWE0bLj076Jxwk+4Lb1ElcSfzw+
bR9OYlc5pxhxmVCgfgv3B0ZygKyoL1dQiBE58QVZ8Bo2En7YXWI9gIrq3P3WJcH0lRnwkjI9HL+W
qeGNkAWkeCavT7kdq/hERm69OafUdKZj5/VOVlaCh165Ym4KkugJNYE21f+3T4crmUoJduKPTjzT
dZ82nhue2gc15at1zT2JbReB7vYqY5SztAdenf938u85ODLw5kw3Bydpkm4Ui8plunkTYEDfc4Fn
TEVEcW+0VdMrHsmaVFJgKARFx/fYYmPLF7YMzLrNKypB1opSg10P950kM5z4karVLOOwAQZYNA43
FC4ttpYwC/LF0OJXjk5uGrlKEIjMlu4hH5P3jBxUqXiRKJqI0DOAU8lcvlpiB6boqqZrLHgTVbzX
2ik639A4aCFdncdDFm2iVt7z8VOD6O6HSbjI36bc0ub1Y7oanJKca0v9btOtNMjAh4fJ6jUg+w8I
zMDqc6twOQFWihzextuvv76naov53g7bi4sphp2TKI9fHgAICbT5LLu0tuMZxZexCpbPtSYdOjXL
Y9zGz54esvb9mahLfdaoFbymy2pRXOWojUfVmK0nO9ur/oID2A7C7OOg5z51TZkPDCmpPof6fh+I
zM5HAaNkTG6LbC75nlW7zM0GgPE7hFKpwQ4BMhUYqJZ5jDrtm2lQTn1Gvu0dRZguFSZAxKY6Ce6m
5cnVcruklQj8IHR6nCoFw/n0Qup5oi+XuyUTRjxafyEfDwRmIoQgTakB0p33/QAGAQkP1XGOMHJJ
6rGknccpg6ZyI7oenhGA29L8SW/YbkiFBwi4H/8Arc7jehrQHdTalH6kr0q3W4a38ZPDglBD7DYe
FsNLvgqJsLqDXhMmFvQQRvHPmUNdbkAdRiC5ABD8dwYEPC+jno9PEf6m/BzrvNdg6Yv9cpuGEEww
LVU8UGTzNbd+zLFtZAa4V3ntD7HHWaoXzFkNVaAJvAdLY2OAltNaK/FMwFBXRguR0wTxNr24cohc
HPOyiCbM+1FqOOL8QNrjrZDvYaNThTF7wxmYup8LC3UB8SQtcBk3PG1ldupsznjyy35OVUVvMm2a
ECADRBLB2tlPF4QwIEs0m1fbZm8f1K0BG0RBo4xK0AVLUGTyOroPV1wjV3FKBXM5/3k5xj18LCkS
8GxidPx1nPSHBIgHvwZ1SyKQPnH3NyPMdSFWD1VRjzojeb3rpWQSXz0It106ZTAQy0WsY8VzfUOS
i1ZGqpnW7a0qnOI+Dk1FRNtkghhRWMrfKvWSnTt/+n14KFfYioMizOpk7OKyIg/0MmbPXZprOvgw
Hwy7vqooYhyw7qoAOADGVKynOUsvZHOsa+Ct3CquptmUu4G2AxFygmJWbGa3xEnmLZL2enjoMZip
T0Xy7u8xc0RquClmci2/V3BPIE/f9tM5Vx1Yblbf0KwXoGlAUXx7paqelbUiqMAY9UtllRnTdc1H
krTIoew3m6OgRzED9hIlsAnGVPE76+YyJhNsaE7rdwAlNxnc7e9+o7elIQSw7Dl5AEdP4gXoTgmt
g8oe5np+Os02ZJE+JgTb6xOJGgCiz9CFpiOuHYVrYSdi4OFeHoDxhcbY9yKrt2Oj59wJpf6bAlsz
BenQbchghZwOzdP1UuGjCpdX5DB3bAj05XjaTxAtPLmIm47m4wZuSIbWwzqXHFjhY4zEmHQXZUCF
J9CTsEaYPjwVxD2B/RLhf3yuWXKpL1mWdy6u/1ejW9eoobgf54F5vKxqjEGDFi1g+kuZKBYU/Dud
CyymAm/HnY0wpJW4nvR4FQmJxMZ7HXbcNl9Xl9aQ1sBokbyQ9ovBfMa2c+FskMftQ2hQP/hKvUrD
t4aNS7I1TH6S7KJ+5LUjwUg/rVEdG11K7NDf6X7aApYZZ1PahFbJdiCoeIT9e6g2fuVTZ+yRqz4O
cmqtp5ZDJ56+GDDr3Bo6tlEFvaqHqJXD8TwfgxmyjdE+9gc61ciHZpdUBmi1xDVPvRFuo0TuIhbz
ykbbsb4NaF4ibzh4fMpZwpfYCtd/EGwqcwafMFOpWr2RVo+MKUsJl0Jrrv27bMHtP+Efkpwyj6sm
3Lc0I4e0XtuirOdxytOxlJKfzm+mK9Ft+78hslcgBFSdTopDJa16ZCCTl23AWt8UIg82FqDNEsDS
jvlHFp5iHXEHE3FH0P+HW9xmlfFbZyTMzB2LTDNyReOZN2XSetxdwkvG5eE2JNNs1O4I+TTujzZf
2W4aaLYZMEYiiKt5yF6BeYc+LHUbdNUoQMhNg5SiVEM0oFEqpENnWnvpiGVqVhkpQETqOeJWxbb4
J4e+iXZRSiuBD/2SWZfnBA+kzfyLhSZ8c8oNMae/pdJYT4Y0G9qTywWLykzjcQy12MyDujelSk15
hZ26HR/dAhuFgms3F9/J4R9JjTCNxOwae/BLK4uH44Uln35iep91QfFmBj5yRFvpHxaLibxmNkgU
baG/ehoG938OtjVf60Tzbuz8USXgt0JgiVFZ3X+QuKwwvomWTsFt3iQCKS8SJ4848PmCx5SSfSzd
w1q35i/8oaOr+70JuZxtgtQ37DcpMO+ZElWOuXcTs5Pzg/0OvB0RZ/l40EmMvpEEZvTVihz6c0ji
86hbswzA7bevyWg/Qqt5U+3lAmnUpGjOWZjPilYUYW+Vbewd4c5wOmC89CQqSot7SqBCFbtVKc+j
V5/E0WEFJF68Vi0C3FppxmxSboONqrkVEX9LWpFLMCvFl4YqUytuORxNjtUI8YzJnc4OrQdFpIIt
KsFWq4t+qB13ivlrxm8ms+iTB4DDx/e84Ixoqw+ae9DxKX+PAonRt8Em7G2PxFxnmFjUI5jmLYoz
brclNZB0/Us3MCaqNTh+SAZPwk4up8cKQIQL/AiwyzJfKIRxIX3a/O3lYzIOR8/zQ1gHeI9Fv1cG
9HgPJiuQaAtQKl4d7Y2ZI3PLgKhIFlVeNRtRDtf5FYI8aqkydWPSx+si/9meWVf9uTmU/jRg65zc
kwpvtsuM/9w7dwZLeFP6zxyrt4gN4MeFeCl5HrP2JP2T4SPWHbmt00monmwkTSuk1heVLB+JjW/4
2Zse+Xh1UEupRZp0fwi5wE1r8edC+w9t5vPjTEQpYa7aGgOHMLHL33XPaRoFebuksgnZB/vwzaJ3
07cHmfBwl7OvWOcKBNQO5Zj8SPGqitIId90DkZudMp/exrIBdUl00NuDK6yDuKC6xM4Cp822FaEt
jImUqUZ3yUscjUBUmeIxANkQB0t7nAdSIRS+clvcau1+Q/Zpy+mCN4DZ7cMjnZF/+f9d/1eid47x
mCN3+3QLCJ1KnP8/NRLmeWjioNOtLdbF3gvwfVmgvlx3bLyKUoxdBdD9rGiqI7Mk6pUhU+Y+V/GI
v4gmUWa1a8lqpkaN4mxuvrYt7HMQDUQxbb4qxADZKv4d7jOD9sAH9PBLyE9rhr9RcbIEIkxPpclm
iRieCDV6DNUuQiS+QWjV4lmiUmZiKPRPE+rsSMu//MkSMR6qJurFhMAk16srY+p9kuwLkFFvftZn
kq0SnI0b6hyOCHn8955ojeF+EZGi8K9Ci1BBIOySIeI9CephNipXIYh59wLSx3T0WCIn5ldIpUON
BD+p3YVfl4nf7X+xNnasWAUEtDyPAlOv4OP5QL8+8TGOTQzVcNpOxLKA6cS+kZdGRTldPuc3DDow
iVLS1svGc8wOMTnLFsDE8UIaVwlHhNJCI6V358qBHgpdPFItp6+MMez6xrR36BwVTyuY1ed9tsa4
P7h/HraRRjc/3LCjAlTt7IgYdqlLainBRQX0sVZqKfclYv7dbriPaWxHLJRAMVPffrqTUtymI6Jz
08jKQOgJO/zPPMgSYcd69ByNIqqe58L8c6fi7MNSR1kxlcq7gdKAKLvJsXKmFzxml75aSzgI+yDF
5jcRFDSkSqSbo7HgFuHf/OeLVudkrFfgzFnRuI/RK4gMUeMjHob061niFF6tH8vxJ1YLxGVSR81+
GHyKbQp/L4C7jbbg9EIol3isxNeZfmtLO70HvsPYpT1FP23ZrW7s//u5itR7bPSNGIRiuUmrmKcn
M8dI5WYPQ+ufhYag9DFqu1XqxdR9beKbN1K9bk/paYLZJsmZwpkp+1kUAjGlXP8yQyJHTV3STClR
+O9v8ptJLg/181rS2PPB8aLKTtl+dRlswIbb17V+HViVF8ZJIhNaANw2j3RAqToD6Rkw2m/bnE6y
UtwWxzBHcDa/PlIuIIMa3H0s5NmWK9Tr+idZ1A/FswQyfjejYugFAWgTjveiI81cDyR6tnhOMbCQ
69KVk6ygcSvUOgGvgBwIYvOXtANv4LxiGWNwTlVKEg9wsiP72IJbGnP74sxxFeGxCiL8OQ7TXQiV
dg50M84Y9OzZm4xC6NDPFZeytLAL6DhDv8vNquMb0KWB8fnTMwf/MnRIZRMmZKYgtlSBmQpU+9Ic
mmJrw2HdVBqHkjqXrv0onNbvuDe4GkoE315/hGjlYjJ4uqAZAAk5MxLT5U7xGTUKA23w7ir4u4H4
QY/tDDimnCIPLZOXTkw9qQO5sr+L+73M+1QlYSxEwKcixUgMCAcIIOubJZaMEa9cZHNCJdccuCuL
+OaLzCizmCRzp7CoAW2vi20b5NQsEO3Xrb7KMFuo59p4WFjMqb6s74l63I4KuyQFZjSfo73pDdUr
LtoMG/IyWYuoWqxgcBS0mOjrA/sOoSMTYaXhaS64rzfwMofY2SEninb2uYUbI8OMekEoSVc6Hwr9
pxla042MeMUHjbWsFNLURWvQUt/54UrBf+f9n5oeCxVpl1UqWeRcwVQDhPPzmm4PZXt1IMgfYjuy
FceFgaZ0El3ZsL6UXZJc4lSZYogALG9vJo9l1e6lokkSezCG7oB/MSOZED65fY77GJ6zlov0j8w3
7aPMSpyVbWeibq7L+DnDMZYlKOsWaUqUJlvUO0CfO5UdCl8KjS3rTzCw1e6u9eIgRN31JVWVO3yr
ykCJdiMWjeCk/hfjNbawdrkYZ5orAzrLyUtv0iv7CZiHub2ViEzGgq2dMDkCmtoTQLMVXheN/L3Z
F6wU+MFSeOdQMSsKZhFYIY+4DTFRewI0yhTTFQIND0XZtj1pbjgCKNTvolq+M5wMW6hljZRCbDuk
D7vobNxkCvdmsB2WwnglIRObPr7Vy33Ron2FIb2YhlWxblcuwfnSJGyC9A1WrWdWH8/EcoPrbsjc
/q/aYWOWpOM3ZmFfbF0KBfwkfrZp/dzFucLWM2DaFZ68HuNshjgDuAkcqb4+6SAY1z9btM34Bwsn
Y2++J0v1R9eIAmyIlwOXZwOt3ZMbbb73vW9jRjwuDAeqC8duxqbscfxUXigBqqPX/+T2pLYNm/R/
I0dPUQ63xhuBbTqzpPUl8LmrKFMYPPO+ejHaznRaBxt/H2gUXx3PtOqM7hBq19CY43MWwNc6qDI5
++RpSKuDsoBQ7enzFCtXvA3F6023DJIPu4Pfv1wr1FjNf/H6RwEScvsd6arAuPHn8h77Q+rZ8K4N
2MfR3d+YoNb5J6VpEBhHLe3sCnHP2CulroICUeia2cU3p3A5deF55gsK9ks3GAw9fO/31e2Srva1
89ZNd9lkQnlwCrm9goGKmkTSP+RP/SKBP67NbFushtztmQ+WRZgBkOLw/RJX1vSqVikd2CGIJKbH
jsYeoaVAvSft5AnV4HWClM2zl5reDpqA0HEzeYTnrbUe0EWkMz7yDheVmYlbttz7Qi/OGBVZ8NMy
mZvx6McbZv5coAsqEfCQC/mARTkcUs+LLtzdqiELYD8IgmsnDVb0V5kr5e/txAyPfKmOLClIUSo8
2sWayjPZ/cWzneXVc4FULd0UwHSjAtswnONGC075/9iD3O4nQL4tz2SQj5gP1nGTzghcl6oawL+v
Fgsar6oB7gkaSXcpUbyJ7812SsXtLhD73jjQOlifT4MdKXteByj2uQnkSiBS0RjoUMQ7IZtyDjgG
0oFknXJqSxbuIj4mJhDj95P5yvVG2of0ULj0d9CXBQrd7zRjAoVxjsp/8YkvIIKJQ1FcWvf/ph+0
2Us7VvuEPkNu89CLNTQCsMTR8zfsQ0f919Ozel88B4bA2nM4lD1VbkwumflHMi1b7Xe3AIvP3aXQ
e29FcfeSVk4J5EYjm6YiBUwITvaa0F2mr4Hl+M9wr4gWKvj1WYIILC6A+px7n1q9S4ihJPS0BbOY
0BJg4kvcKeRWUTw9Wm688vXYMWlxDmTGuCUQoPAISIgI8QBO3quLRLUhV9EIaXc80b+E1xJndOeJ
SCB4VrxVY2PZLn0L+3/400Z6cCsI6LAtHWByyqOSqEM1tweea4etUxz/ifGQiUfvb1iVbTcf2N8N
qMCsbf3289gkF78OnQx3j0DnzXkJYfBGlZrlddZbZWN4emHKrlmqNm7lqK9hzJsE4Bct9zRr+e5l
P4PGViB3vJYyhB5uhmPM29undqWy9k6V0gBOPnIk9IjPojFpZ0CDBv0Gfbf0bgHpbp9S8DCXR2kg
EwAvCHgiyN6SmZIOoVN5M5XR3z8nzgzpDsLFJR4lJsjLmgyecMKwja9VVgLcUAIhWuQGxVrMi/oY
Chcjn6AJgdTDidHOOF/rpfOoDfYFbFn9RdQ/8yUf7A7xaYSU0+hzDLBoCym9dK9R6vqQN7KMIYCo
q0tEKkdFv4NACGW6cp9EuM3J1frW7MNUMtp95jGKnZ0C4JGwiwdU1EdZSyVpNt1SxLbjgSlk04t6
k+3KwIN6i7qJGwUYmJa/4sb6mN9wyzq3ZQ9LDayg4hkEY4x+ljQp4FJ4UXgP97lbbJ5zFNvYjTD0
LLCwCmK0Ho/qJJ4HJ9GVAHwIdh9udpQjO0g6Y/USwLY/wGj8WS2/j3gB9PBcJPN9FH+23PkI9oJQ
g27OU/v7ojNc4LJtXb2s2HrD3NMmIkRYd0GLGkNsjyzcdkmjn3J5IIFFaL3phjvLPET5sKXWOjtW
7451c5LB2RCIb0I/a1AfG3Bs8Re/FMCS+e2sOpVwMFZJqwqSXESNADHlesStR/1wvLBoXlkZ+uzd
AWvJ0XIqmvno0GN/A60wtZfAwgx0CujpAsrEeDMPL4EhndgOVYLO3F1vrEdrdoLedLo64Gu92+xc
UPHEHrkJunZsT1h8CX1R3l7JLtva8KENKMVO70ch0Ztb628ygGfKhCRvAz49pJNqY+hPeWsoaWmM
4syTG9n23vl02HTFk10AXHWj4/zrFLVPm3rsXE843+fUzCEBCCFFZc1Mhp7s/bow9W3Saz56iQ2C
bmz1YRyBUYt7OXFmWyizxAfvK4KTTYDbqLnQ3OHvJV+kDhr9xl45vhYHRKofHbQk6q8PReR1pXoh
4E6mcAM2XsfhAJY+oBcx1aeFRasUlGBqooZ3jKbPCTIUvAs3NN67JieFCjQWfwl1+BALsbl0yWOW
ixK0ePPBtCIFtT18yEiobQWv9+Uu2WakgLQupZqNNffGRHR31sm8tr47SsLpSfYjFt/TNls5kYxk
JYG8xG8Z1iM/wZj5E0PmPo2iE0zE5nibHi2b7aXo4u8MQuDkoxWgSOXJ5/A2YKoeCHtN1quTCN4p
294m+XrDcw6ksiRHzqN0hYDGnD+75lUrFwxTAm2VXT/lQadI56SshUYS8ORof+zBsBmoT9+jx/st
wMOnxXR0A3m8Typ2SXXTiXnrIu+bNl+tKjx60VtXOTHrNsg8rxeJu5Nr+/+gLeS2I8j0TUrSzM3J
E/lOX8sSZ5AmcVcWlEWyFk8KQDeucSwijG9VzcuIh3dQHwYoQLKCGom2kKHb6YUWMcE/b3sI4oux
R48U81hpbPRIVEp8Qp/0MWkeVWzpXRhA5jehpHpgt7XhGozQGcaM3tNEyvsySUN1OvrELPaNO9kd
igLzyzMj9IHPtOxjHx618GmkL8mrDW4r5kpVZfvwYNfjGW3b7NODr1lribSWMtQRGyYwTizWoHHV
Mze7IfYBF6InKlOkbjjBGikPKBJzg0TYnAxX/QUZHfaBrRS4zlDG6u/TT7JB0Th8nkgdbAJh+oVS
sFgTpLkFt1FywlGvx5aWsCf5FfW0zztPEZ7pDzeHJFfYk65r9T4aXHMcurse274eUIMntkKgiJK1
9qf6SIUrrR46XcKOOOhS8FdTt6TaQ55HpouOWyRe6PMAP3akUvdRHW2ObWFr1moCD6CaOZ5B7f+0
+LuzAtn0HWJWyekRCHBx8DO4CRHlJlbvUNR69Wp/n67eHvog47Emmxq4M0vF9unRFTwQS+tdFLAM
r/VHTU9iMlL9EGhXr+vCdGYWzBlbdh7V464O39irG6QjxR2KoIHHYz6hBfbFe8F8EG9K9f6hICLn
OvqUwREx5bIcz+pT4k44HszyLb/29FiDtt/lrOSdH9/4XxFwNBp0l4eGZfsRcYUW8H+ZHjpxa+p2
hoJ60cSXNUBP9YYo38dUFi/tONLp+qun/dFgBcY9rMGVf8NL06UY+IbwCDDCttWIaKTblCHnqQ4Z
ZXn6Ia5qQCLqCp36C9Zaib5AT03BhRubH5iL3myjfGCCB8+hGutDpISjxSZv3Gh+0Aeva93CJ/Wv
T/hIhDQRR6ReFvcVC4IepcUh2znBVoljtDL1LIKpE20+Ftf9zrmWw1RJGPVOTNpzxTVfgfJUMLbP
fL39KQBQUKyjwFwjTfO37F4CWIiAPSrPT5EhuKP2DGTXiU5mZWrvUTxqM8r2v3GRmfxz0X3PX8oF
HCh2EyPmlD1F7SZNABwDEUFHC+WJQKXUJQ4FaJM4D7cX4eddVsrB9iZKmZMq53F8J+B30qNGmilT
91ypY9IeSL2O3VpDap1csjx7eFEw2jNG+bsXTycT10+XYK07mFD1j+/5SH26Jyb3CuHniu5r4qPo
kvVYQJ+d39ZPollclYZFZmTiJ7X5sV24HNscjUqm0K1JnG5pCwuzsvYRZQdZ380JB6MOxWp58jbj
u1/cTKLONHdhQ3/YJpbD9D2s4zOQ69EM3AsEUoggeXZQhpgSnPaimVvYZdWHx0+ldSLgG/Vyodyf
tKmw77jKFGt0K1WxtzYFkn2xXt6oXbDvflNW0Lm/S/edtG5zvuJkYiWHcQk1ld9Pc10C7yVDqdOi
jImU6M4IUWCLdcfoT63Obqnn9g+SMA8mH/rqfxHccsI3F4x9EN65kTc57lFNKveBIyWM94Zt9Z7b
LMjWF3p3i5qNL+ESGWgD/iP5Bk/c1pE4DNOI1PoOfGSH2jfiW6MBTD+ucxyz4x7lzuhg3Nl6GC3a
sUYv/ArGXhcCTOim5uOAenudRLMjhFa8lou5nQAjXfCivhs7C5UKbRD73mSHHE7He3IJP0dFyHIB
U2lCQSK3lCU+bUR6k2t1aWZ29iiijHs6O1TFaTq5sUhk4Fhrw3FAUSd71FVBuVYjtKTtL4/sPjC9
n+4sQC0N9CSfYXhOm8bmAN5Cf4OzKReWN+eW5H3VFK0CgePN3FsOMeKolWxOEORi2jFWgB3yv8+h
MswEMp0A9qM/rrhObwKdAM7Wc7l6cHeYRkHujYWMVTsEjmcnQbdkcQcW9zVXZE5s5vOgJBEY+dyi
3jCOgdvQ8kP2vqhtS8hIlRoE68onTewlWEBSLRTqEXQgTzVIjG3f0/B4gtBHuxdYoZ2JQgj8Sn2v
kA007slNZO2rfS6qIKXSyzml4Qazu92mE1FiPT7NxiT4lW4DNNqhYKVOO+JgPJ8z1Rx64uks3dtc
DhlFWmqcIyOodgSelisjM/v2QALvHQxgknVu3WQ312akr1PvlnVw6vdL2HPCFnA2B+pgx2OAwRWY
rFrLBcbdFesRBULLcT9VPYwj42ApOQuynYU5oaVXSXoY33HB7FkxQkpkOtKXqQD+pnZDXi24Ugtk
Cd4Bl5hWb9wlXmZ8VGVa2Mpe89GO9tIJCvqT+Q6bHhXvfTmd2gc112iBmdRceVS/GWLLyNlaO+fN
nsb2k37TMHQBkgrprU8gXqeorkxtKATa9HnZdYsdgno3VOsdwoTm0jYz6mJEjwRl6sTq3n4hMXD8
kpLBQdXPFbk9BA9iThUViNiE9NrQ+WJsGGwHp1y3lsKxAAESUE5JClWNZEjLi+utDWSfP0vaU/r/
FofKCgBzWHJ20Bo88A1IO5BNz+lNNQa35P/DaemGk1QUFFTkAMbc931JR3uetP4Ye19g+GY25VLq
JU21EfboG2L3mtqX17n5czCbV3n3+uXhQuvj4CpKj5GheUOaBM6XY5guw8745GK9Jzt/fJ+uOO8U
m3PIE/BYgI1jan6sfn1hN6DStKtT7VZNe2nAjbu16sDWQbumPu9XsPDXe1dLIbWDFjM6u0mJDLp0
JIFL4OoJe12hJCW1if5DjyBy5V2c+9Ii5rIHC5EsP0TFnbpXSGWtgJ8X9qFp2imqteRVttEW2T0c
04DJKOePwYGMnjsfH3zzMauX0gRHBo0z8bhP56BUeLqQX1jsaaGlni3a5Aw86RQe9XX7YAH0Y3TL
C4V2NxLy8iVwOI8iXb5zqH2JBf5VAeHTuZRkjOKABit0rphdPt0QpBViKs5RueSuvu6qCET0Bm9k
oI5/b9Y9XGBgZZ2VGWk8Q4pNbdlLy0dpXPnngg9cJDoa3CPV9oaztnqpxbBo5MWeWpPGI3KUv0BN
CJIwHz86G4NLKawlHgRcrEiHEkc/aKhqdktroP1qYi49xmJtUZrygy/x/T8+gH2CyGAVtpQVYEpc
Ma2+KJe0DokDWBDhCQntLWP69lcQ+lMXfc3Fa/lZ+UnWImWIHyicZ6pP6nJbeUMn6zVMhgNaJaS/
Ou0/YKMuVq9WjiyRFK2rTZicViYcID2bw50jgqFahjuCcLhBjtbUmj/CQ6hzeTV05BRnv7bilU3/
vcSw+RYvh5mYTdv82/k9OJUSo0IGqOovs0/xWIhFZgJKDfqsiwtw2yAF29R716STSFoO2zgTprIX
/eTZtUGyXeExhm8h0B76DFwTGw41bpTTsnrDOjRmD8lIvpF0iXqYwd8cMpasqcxl1n+rA+48Sdxm
BJOCvAhqzBN++WEdAomEB+8Ly6+H7J+CNhtqE3u/BOqmSKanvR0dcAXNKB4i5BJs1cO9TXPSr/qp
+F2jhn0uidW4BeILXsItQBfwtw4ijL/2w6t+b4pYzIZ/a3+pZ03rUGF6aJMMrmQyTC0qBmPuqiu2
7fZoyKmvEvnj0mLDOlSEdCR1KrNuAzc0n2H/73rmST/h9pLrUEUIBqYLEG3DMZoEQvWvKGhTiL8e
cZDEQMgHLIv5bMXq5BJqS4VcbqGVodAbnUWmp98I5xG3gZG9oRhBIgZo9G0DBlD545FaXl0asQuP
oyHZS94n2rJTlhX1NZvmWwWfqqn0wHQbtHzk5fVNEXTEq3mxQcYMSFiNZ8hnnSuG7xSoPEgz6uRO
WFcsyHmUwIXKDZYn8nav7x/6BC+x9zlcMgsx7cPbr1bzbTtjWr+fEWbx6xj1CluDlfj7j8YUrH9g
m3a7dxiIMWyBHwUbO/T00O0k4sQicf24+7KKB37AMRPAR+MM5p3ITLOHIIqYGi7dTVQfz3V5NYB+
bSBYMnrV1d2Q7ooIyAYgYo1rZhpZOLf3kPNyiO898wUGx+1H8l2qe3wAPunI1OKNomIDe+7h0Q52
a+CeRkYfRZwYvw//1fXytQwHv1n7hJP6Ose4hoHdKzyTIuxbDgJXF1TQcCg4cukRq228S+WAB4lz
YPFSi98bdW4Sectp6q1LOshufT37+JKb+fLYGrwklzLG4tWc7gNSD+Eul1wLBkXl/NclDNQ/xU7b
3MWZV87ags/TwL9T+VLy66O+jvquzRpyggQ9jXuffbksVLwB80PkP96gfdk4Jccb2a3gWsb0uED7
OG0pEVplFLygm99/8lo/nm3UH1QaYE22/7Mwcxmtyxe5uHmYx74MlNVGEHRd8Sxb9piVbT7xQfBt
O4sd4mLkrDjrmc0VJWO45cDHBu877Jm96r84fJzCEyIxzZmzyaxE8U1Nyiasl7RJtLKNk4zzgkhJ
DTT/Uhec6o3F0MZbPsD91JGnURbNRU0M6izg5BVD2MA5yLWm7MBUVgZN2swwcWMk6V3d/0Dm+5LZ
t+Pe5T7GGFaofeiQx3yrn2cJg5jWUpK75Ko/nm9+5B3AQ1np9kVGVg2LYJtLz5RL/37cCtd18CxC
8J9gk2inwUgReIcHllMNxSQKAqgFvO41JPKz4nYA5RkPwl0f04/WaZdUbGZjMm6lxWUcapyxcNT8
ha/3pl750XO7bvoF61x1NATGTXTwPsidAJi/PQ61HU2V11I1LSAkdSHE4nPEFY8jWJrCR2Pok/bo
icnAZ1iYfEfQPZfadt+s4ZUMQsk8tGfFSuc7oXJFgBTPVnV92CtC8z2C/FoAzK/F3YIF64v6svlc
IiHreOVQCk0MDktl3ubx3HqYj+24H9TLwC1q5ggljcOm5bF1rRcXkvra0XH29mavDZmbkZKSkV6a
0uTWPJiJoiHfbu+yR4xnOBMSAQu8Q2FWKJJRGQuZWqpPZC79idrO0W1wiE3Jbnfm9A5RQNdeIBwB
5JCZI/qsLvdg7ifWndZu1vZG4d+ifPDcNhLZW+DiSU1R0M72CQbQtjk+FrxWQ5NBvLNlc1CDwQcm
6HFE6hrx8xBVHK/fKIYKMszSrTo2DMMWiPSvzrwQ06gIwWRrZ80f7ZxNKGhGiRWjqqh7nGaCD4jB
6DEBKBZjySqiKoB7S/tg9YTAg6+qWseA6Io/0SIIkOTort+6S7JKuCrwiZXwNujpwyOC/RNAWh1M
ZNhEOKUN5EauKYAKrPH9hxHm16V4p4NVHx7lPJPsgvf/7YgzPxgoZXlKP+LT+4KyNaS1tfs5MjWo
YPexyHwYwWDF4mjycgTTDThvjBlPdgmILzM29BFDnB6fwHxLJqEHPcsll8eRL/mGY84TNGt5hyht
phVSgbAx4TrDuDQRZp/yEl4fsf3ra/X/VdLq4yFFgWPhM1LUQvuQIkppXEMQt8LzHvFFW3ryMJ3f
lez/ZzkIlQvSuurXWmKjqq7m81n4hVwUB+lz4I8Q7GN3rt899Xg4e4UiJruGTwBu4Z5ab0e/NDDG
IyKOLQJgBImOjFCL1+jx+JBWlPp1mxV3lpTyhE1CBLlV3VTmPjDnPVU39GhiZAKPQxZXHYPy7lln
AWx86DjD6CiMA1HASI67+QaGcPKie1TST6j1NWvon4nwA0SB9VoNvOx0aOjOPMonQQ6VNuUJjbhc
HpwrOPQL1gfeMw9dYBBGW+1OaPHoncYgxU9gl4dIhNOVvPEbmV5D7uZqAxqqMZcZN6Mt+2cyqqrH
RFoQzZEXnYu8IU02qq5WBj3iQHOUhG4iv5UXMIsj79UQnVMHJEEzIlG7nPeb6Vkxw39lWXaWZDyf
I49mpIvZbDeb6pFQTFQDhW2heQ8VKw15OfJDh6iwDGeYFz3sG9kRIrNYTCrFYShZNGjx6jgxtoBM
nj0855ZSuQ5iEDhZQNyd9CgeQ6gJQIqksKHwBSO4XkMDjtLEieI8+enatpUtxsOr2Q7AYUUn0ulR
JEqAGax3Ix1gCK910GgSTVcWD5v5xoQ/SwEbYLuXCLl6jkwemY8vDf0hm2l0k8sRGKj+hu6tlhnv
Xk7CRgQsEshVfFb6Ys1TKtKlekMyE7/1VMscc+wwmOyL5O6MHxsbmz0qvKOQPMxgyrDtJJM+ryDi
3ubcUSWcfAxuR//rZfkPDykaPDisW2uuhYY70sLZje9o/m0S4Z30n/qxJp9B3e80Or/vhIs1ZssZ
uTQHFoJDf1/JBN5xhPiyUklJC9CIc0dEsGTPj3XlnYEz4aex7kbhZa+evOUO/3iX+LfZvcDaogZ+
OvhPC64JhbXM8FrB133SRT+/gC26jCrlNzQsNirycbuZ5SJDOOB3xeWB195Fm+RzkdQV8YtuoGGO
Pyz19AOzs66q4gzn91A7JIGtnF+Gm9rV4yP7FrXcgVnN2f2loKQlctuz5x3yUXH8JqGD41Y+dIvp
LtpltVGvlLIToG8viSKzXtzHrp/JTS3AsiPXhaNwzgE3We3MT5Q/wqN1WQHl4EFsKBYljN7NnaZ1
mNsomn3wqfFn6Y5SAHISTF2JVO+usCsJETECaNVzjnKtyrT1PRbluIpqlDG41h62wCLDkaEjZpQQ
SkXnratBa15un996ux33OD5pSNNCtv/LYyl3sLxUe/FUYQhqI0xmbnHjRWedrxaaq3Gqq6qTzlaq
PqDWy3KK4kldr4QEsnGFTc6f5wEhdhdH3W18GWt0hTMQg6EuHt51/4Jiwbl5uU6zUQf2H3fyejpf
QmfKfBubvoKLxqWwjpmKkmzOGb+GDrzIM8keGdG5UqEmDmu5v85viGigk2oTRN1X3k/hnu1zHdbU
a9tXjiS8uAPsVZvC/z51FDowkJ64tKR235uStIrzqXBxT6Yi16fBCIMqqUIKDKKqIGn8if81omxj
mxP4LBbO1MUPnL/GQ9tfHpaYe5pNYEXhdW7Hx7gymrv1PfU0MXnFqZOpSDYMxUfn7Fte/IsYM80w
+4iiVWC9LHoBr2DknXG/+6SYDhJGsimp9EkaH0fHqAhCsftvUq1/y8E2hOy2a3JM/VdYiTwi8npY
yJ60mOuWcsd2IDtHmVyQ1fBYE56+0A4EMJdbt6W1f9fCTSl8sVopn5/pivkd41Ewq7H0+VyiibwN
DkD6e51938EO+Iz+RPATh2aWKH4TVkFuuWrgbJms7RIbQ+BOixUBcDkGXCrokIYlxFVjzlqGslCk
8llHi72bx61MYS8t1yaHhvl6NnL1pFFTAgc6+SHb/2zWWf+OdNwmvAWeTzw0gx3xCfEQQR5yoeWl
N+qDV+y9nwddGE5pi9ehckRRrqysY/58cKRNJCUDuhZInpneQySJB2Js8D9B/VUzvqyZPlg/FL7v
3oPXacdERotm0er4seNIE/DsA79xIgNpcrG5KixLHIObjto/u0vfJnz989W5UhqIY4F+QcikXT/1
SLmqH20Rh/kdwSnxeH6IFw0gP3UkXDnQODfrc1oSkcmrf35pbtghBUscu5DoCQH1HdVi3f7LKTo/
uZL3z6khRdpKNl6ZC9lDE7MQphbeBLcvNpv6+By+nKvCRfd/XKXMByG/Ro1DNfIg6H4BeZJK2orG
LpTG7baFT8XCz3n7TFeC7KBeJG9rz7tzZcR1ftvT75zmB8AxWm0ozKWF8MsAPjJZcPPM/5fsWWaZ
qrq8EwcXLxu+XBX1+ifpWzyScIxhfn3hg/QjT28S7rG69S+SDTQDl9gArbHl7XzGwluBFKnZyIbn
oZSVu3pKVhTNAw3py5UJSTAbh2IfEN4wDvS4iFX9F8zW3fx4+QrJNrQgTc15M121IuBgcAetGze1
XUFn1N4KMOvcVqNOVnU5if4zwhNmN1O12OXuvwzbXfi6WcYNhb6r6oooy6ANsS2uGI0VfCPbQWUF
3ppbf63eDGT4CAkxNWP0gDGxKjBtJ2bSl5KlOpAo9IomXyWy5jnXBehrVfCFvqMyaTiai2aByVTR
GuluiwXdd29rkrdDVvIVFdqolzV7W33+y+6gw5L9b/VrkGj6OJPbSuciRLOBQvUTNZveJ6R7NpTG
Lrm6Ptmrya8dorC6Tfqasi3YMoS/WWOGJpBxA/8dPowGI6/vU80vHzRp8CrN1+frZa1voAZ8E09s
iCjqJkVpCpAwJkImH56XNcEzl4cKLQVx5Rfg4oVkOQs4VlxpGlUUZ/Zsvjxty9buWZpgVjGn9I3z
Z5FFfy4uFQ/xAZUJjFrrjoL6SEngT1cClB2JKAiWwixepGRuZeol1tNTiBVe1ngdbw7gA+yLyxWI
NfE3gGdd2ARkmu5otRQ5D6Ctx1AX6xS1bc9ne3n64YnmLQVG0mwExRmlTmHQQNSzgiC3sLYTyi4U
65TJbwsZH16ZB1iEyrutf2Q1W2hXzYXgu8sZfmITrOwMXo6BQ+6we4lud6f4sBuaEarSHUlp3NRQ
e1+Jdbv5xYeGQ1kGpt2wgs6Pak40xUfLp8nsCmMBXUYnjP3zIhN02CooxxQQbIa9gCGeA1YP9vL2
O0GfJp6BW4dIL7Yg9NWBRSJKRJDMPXfcfZpPWxPHv5+oSuXuiMi7tTE+zXM1cjdUdFX4pMzLhC2b
nON9RBUT7F9VrhPbZ+//0xnGOqxTqvkmNcLdqGJi5QT9JssW6VRZXCDsj+LFShoFQtiSlWnTL9A+
MU18YivBOZERNYmgYl50RH8UMBZWnCGnNcG3/4Mu1rgC70816OLEaGUHtZBLPe2JTlsgvk0bZLio
J5+ImWvs2GABRtvv9qDXi4KgPj7kkfKOm6NwuQ4F9WA7aWJtQPOSnLiFkzbnKT7HJnJbrgmS+Dqa
qgLD5D9wsC2oof4iUndjcblnVEQ2L2QQegklo+E4BsRF/A6+QcdwzN8Gwzvco7xHFvzr/jYehuuj
hVWGO9jri67Qw8aZgbxkX026dkiDRt4Vzmr08joAk9v1kPwFMIP3hBLWf/MU4+Ca3qH8yaD520sE
PKPqgdOOlckOnpqdNllkbmRJE5P+ZN89knLtzclCr6X3QVbvzgErdzikY/JeqIRI+NCYlCJyMie7
6leUkjVNNzoOsOOjECpUqU0iXQ7ApzV7y0572AQXWXxfF8HgZWiOa3sd1h5YMs1n+7ytC9vrpsq4
58v0hAczQTejYIqbObrPwVx/1Sh7Iv5sneDWSsfAQUS4XxQ5CjVc4D4gT548buNoPa35EVCMhEJr
17Gac7qkDze9xJ7voMLGD4/yiyJsD75xjKxrBqQoa3vw+/wbeRQa7FGODKJWzqKDE/Ez5jfqj6eo
sh/WkyKjHRrKuqoqCkMHPTfwnTre81533vzX1hA43MFlW95keOHIRW6FVzifTA31bxvVOq5jixLp
SX9TvJvPdQ8orXry6BJh3u21gqYznnr2uvxU/Ykls3tLFBKY1nFtcQbFq4Rqa3kYJL4/5Xe1i2IS
kRTFaADahRok6i3O8cDbau5Q6iBztzHgNKVUuYel28Yhx2gWqBPa0bnKfrKO44tQWQ9//4Oh8/f4
SIkTT5bjRo+dTlIohv1AhmDKWXPIxtPTY3KUmG+VD7lhT8OcC8OrA+8/qPPiJ2Aw8l1cqNnA/Ash
/pfqpC0cmMNGzYK/Yf96B7kCWp8nt5lBPbGnJEkUsu+1BthP5GR4pfvnoDJ3PndUrZbTMxRGp7dR
ide6WAEXyaR2Guj8AXlF1bctg6FYaDOaA6ufEVu6muB9cICa0JfXb550CFdoUE9w0uxu8RA8ygJh
8QoT2L3ZVpuas5tVuHUmJiOqmCiM0o9MMKkieQg36MPAVcl6DPyf9a00yrtv6AGOVsMhKgb4QDpH
ylp5YToiFDX+k+mFoGXvvKDlVafaFQB68YhG+jiYHccLZ5S/jVz9d4jF6WpKBuaAl7WwOsnP3uU2
5Tggk2iwScy1UFaBuwn212mt4mxb8NEEdl/n7hlBpLAfV10Vt3/5iwC+lVnzeHghIXQgB33hFRRm
0c2WDThh90zLzFocaVv8MrM4a+KNT3mJL9LVVN0xgnYf0shtT+0dKhgaVcLbb/e0nGQOb7jErdlf
DqxVMZXI0yBjQXBYE1qZm4T7q4HCbDsQSyTz53XTiQZ0rtyWJ5y+LV4STziafFAgYNh8GrKgFmXg
PS1CkFQ/sHkq2hu94yeGDOqqGUgcE14/PTJa4xjtWYwKKYwUYC1JZgCrx9EMloOufh9OqnnOFaZ1
vhqHU4nh8QxZ14y/FZK3pBef4HlQuGXqQMe/4vze2T9z84JRL1mSspPCT+n5/jKTrIqv1lK7cF1l
2aHZ2f2XQrnnoWRxoPDbhfxyhj3g1pzoda3xlndSPZROMNfc0RW/HV6okr3zQo6o6CnE4/0FYrjJ
TAofHtuYFjzH3dP2kycleLIIU3PYiXdMgdxGYUpN1z+O762BzayjKu3/iCxSMr3VzP0xvuqiAm/P
i2+jFBqw++TsU88H/r0UU/UBQaYs/2QnpEEjb1Sne4vp05CTft9AkMsvK7CYfKwaBzTqpgwqN4wL
bvkT1D7x083oj1Ix1XtYztrPle+jBgOkgcOe4LnGQkar3lPEGZmvq3A4OSzU0RVYXsr39XR+sUnw
W87HoZuhZ7B/x7Fts+NhbCUFNmrlss7czEcpS5sTedFc4kis8PH4dJATLUlrzUgNziK927obWnSQ
KI/6nxPLm/JFRRsBQFNgxJMWAWkltc8kfoeAopiudZyoJwFONMsS1sQYJ6BHqlli759ZkWJk4bQE
qt4P4QkfW/7W2GNb+lBe1v9tDEQieo3u289pS+Jv1k6ZHDpK926I8/9Ms6D/404Ccoxw5itC4eyd
kyBNxIerwmiOQ8zH8yqu1S3MlUQpy9DrrsbyYSICg2mxoSuw3f6XlZcf5iT4LuP/jcApR10BFdE0
RVF5SVUXiz6YnNZZN9PZFJNsuwBnK/2L+V8nXmpXttv8HpvvqwQw8+8HyYNH1wXcTt/x8GoIk9CD
GnJKyNF4hkQoBQG6ctIRS272M/hW5PSHMcluuk51IdRRCnQphEINZRin5+r2+BiZKIaQ7C44nZjn
M+Lz943VwhU8xBV9H72wWvf9jNrzHKqdIHmQBXSD8Ugy8RP96l0EAbTlJCqdWY7oOB88lH0cVjmW
Of5LYkL/4VQCVUF4KGPPJVexSdku0tx+yuHPzAathpUsYKMKTAnsSTtTPhcTkRqOcBBdgze4ztRY
v4v1e+AKHi93zv87OLzWsbMLppHeABCTCG7yRwWXlC1DU/IcOv3EeZdFoW6E7CFGx5Eph2JBNCq9
ML4aA7f03ntmJmhynQzHO/0WN99KeklG2CdZImkg9qGXllPuEj8LK9IzCqLmxHADHiwKyNVatSVa
rBvfOPNscEebKU0RbJ5OUFtvE6FWBH1lt0cZ7F8o2McfPZSVGToq3pXk8ZS/kN0TxloihxFUsart
12gMSkFVC1AAPOg6am4GfJjX1DolupjgRc5Mpl0OEaKZlKEiRp37/BIkUL7g0I1GdRgrRPyxK0Kw
PSlJAJXRoV+0M5pQ04WB8FNTENt0fZYXz5Onoz2508X8RHEo7urImlULZXMeQxX0cE8+8DLntaAo
ODbuXUcZouXj0ibTupRFS/Kt9KQJPdVG2xPsCIdFhckPTQzOWuWlouF+uiMlJdYpxFRsNOPJLr4G
grskLs2F5X401HJyAknMkAhMymdOP+uIfWAv/Rs5QJC2iZs3C94DVfiCd32sTk+4L3LKQeoIzbL8
8XTqEJY05tvIMy0v44+0puxlrw7RZd4R7dG/hp7aw0usHzcU3Fv9bN4HgncWP0Rn7k7AFmd2IWV8
1IMIUDpAkYIpxvRBeBicaMhGGIS43WcTYjyEwo3aU9to7kYyucR2FZ0UsoofNEoo2JbSwcBEqxFe
w0i4Hve0jMH7SYTfwQb/pTWYVluRhaKN3jQ6Y2eEOWm+Hy/OLNuimVbOAvEM63PvIGu75A5AYW/I
kDP9GXr1Fx3DSsBIAw5UI1+37Pd7eKQzBBWN070iAzRJwrj6ONZ0e2llcUm1ShNVQx3oVmgdBhsU
nW80ugJFj6CnV9cL+5Xd1y/xLsUBCJX+nlDrz1KLmY85h6Bx7zAiZV0NNAeTBxbpifPGaTev6foi
z1MZ712OM2y6HaZjdPTwoCANWhAwYhIFYc5PxLe9cTXb5cCRq09hTsjFBTUYfh9at1DF0pZMgFGB
RfLzNPNxsAMdphI+fOqbjB2pmBfvmv41ztIJ45Tx9iloxyPQy81HHCtu7ZNNkWni5yfNJqnrFU0A
Z43Yqu3e1FKIRwfkh7COhsHORv/2zRRDpIzgc2v6if7MTeVJ6aTJYZFzn701doBZHH7JwubbdBIw
DhINKZSn6sIt5emDduCZsJzlJktp840uB3PBf0sMnkcqCOhqj5SBW8jWncLe+76mHpc5akfg2DSz
dsjh+v3plio7bR9PXbHIJsQ2hXcDpd4hQRGombU6IRJWHjsQX4ElA7DmbItd6BtpDzfFtZT+o3EP
ffEVH231V3XKyiYQ6/DGUCpLsYs7OXS3XJZG0L3RyL4A63JcPdxvrey4vCN66cCRVji9/K898vs5
BwIlzUBIG6kyvkVFt7npe0nRbLuXEK7NTLvw0HX9VtLz6pbFQP38n0FXP+quwKcoAaASVespgAxy
VKNpOZOUGpSuYEFZEQCIyHbVKx7QI5TagT3Z/SFUHXey4CurjZt7IMQGnbRu1zuRSHgC1cOcCkTM
+v8hzC4Q4pb2ZBJrxX2guuswr+VZS4pwSkBotnO5ICYg2oqxN3JCc9AVkiZ/z5qzOJMux3lD+2UJ
KHfVgxzYlDgdQDPKvUgcQS6wSomUiPb/C+5l4o8VHwNLu78ax29gzCOJfVgzFelCJ8wY0HeyKP3m
tL3Zp+Gtl4PUnAorZOZyprcCg+ABWfpcRy7O/+/Z56BXvYwclvlXH/Xb7rfJ3+qLBF45eBbC6Bi1
jvwLbKlDpcxkzW1Nv57vMW1kdsRzi4/0tO2YonF4G4zM6qRA2kJJhi3yRfZ78wR19xc6bVfxFvzk
BFYOEiNSvg4mFDn0isDCr5Q87RcZQewluwTaO6WLjrTlP3DpbXlgWrP9pNBW1MV9xbNKzA/T/68A
Wkh5BsD9/50J9eSStEGlMPhpYT8+UFzfNtM+vGn2U3BaEL63FTLTrx9ZsgX+wOBAD3brU8Ke2S6x
qbJE4PUvLU+SNCGY6GGJGtSF1xBCRs313/7jYsaW33ZIjwUc12GvqRTLw7aC37yrik5quQkGVNbD
uP0Er69EDnFNcOJ2/8/gaUJ1AMU9tkw/SrKznBE1KZvZfsV2nEZMDvTObe5j0Bu6VrdNtvY41txS
61warMVr++LpokIB95yJc4f6wmL6zZCYj8a5hhtzz0oPsEIrQgUGZ+wih1DrhFzHLTYX880+reFf
f2b41SlPOl2qB2mzDHHSSwWKF4fwPeU9MNc6l+nKOeHXANRO0yYoHAuvFXL0iHj2kqL2eEbDsteW
vTH35+g6HhVhahvGbL9ijEip1yCe8yWEHX2ZdmfvBS/EfIVMdBoyrMPERwBE83YX3id+w7C61YTj
w1zwML0S4/hB8QIpPoDUyKBTWcS1yqzAIuohdqAY7OJLwzjbFLvATzqWgI9hzY5TucGw8kpgvxFv
xP9isEfh6D13wUGM86W563QNAf/7z1T/Z2vyYExr1/i4+FiPdiZvjU2p671lzrFJdYA1a+jwN1Q6
Iz8S8yqiuTsaHBA70lP+VuMvAwuSe6djfxgTV8swDpL+hH+9BAaB5qwVzpjS49jWoa8yB64VVVr3
U++8MKEMhoOlqmK03ZLGpulfAxIxUnJRgjZB9Vw9Kn2MRXqCzbmV+ssFa/6p7Q+IOPQk6aN2tygZ
0ApMCu2hAVlclrxvmCgBqrrpQAA93kgI/yXvnT5aD7X/NDHShBAnCYgJ2RTPkV7zDnTzpuQ2+e93
FHlPZPGGxgUYt/IK+HhaXBPNxc3h8k8zzilyFCGVhNFeVbvVZrS77ylMXvTNpJRAegOtpREt2P5t
xVqZOiGGicYUFhtr9lnY1UlSVs8BYZv/RPeJf6RMxre6ZM7iR3VfnxbZgVw5nIT2e2xCxl592Ol5
rcJHcN9KrnRAP53Cl70h4AdinDezTX3jCufQ9USVxh2dVjgoWn+eRhSPyXNPYj32LDlxO6nU6RXH
gxjnNbfcrItBpvI93GRmZMHiYFu8TA2rDwTuVIHEIvTy64ojzZsYfyC0afeg/nAlMFWBYE2xrU/4
FHenCinUS6A+Xwzcf2r4HCbbcsEOa8KPJnMTgSMj/BrrMECePC5xe14M/LZ9Dfsc0uu4NlRRyrgq
/OhmuJynUgf5ZggMGaK5kvndphQGWvk01YESO6VdqEfWX/P2peqHUI+mmaAUOcLuRCwLLrtx/Ydm
84GElOnWRcTkTxRnnKmTzAyYtVwDxhBHBBzfymQkVKnmceqIFGsEV6ee/FMAeZR4zu4eMU/Iag0q
qW3Qaruaajx7ktsbkElDWmM4maus8lXFzwF56lzWzXXZmsPYjMWcDpAWqP/j+tWPqw3oPm/CMzSV
t9DoOxc+pnoP6HJeUspMKhSNzbkO70QHJ9UxemKNq+yPod0CcoeYj4GfEodCiQdSn3oX8rjWCQ+0
HrMt7xtIzBpQoEfAAAq9K+yDZhdsbsgE+EyeJYXTITX10CScgLfP0LGAJ6IKbaY4FWNP1cS3xBMv
LKEnoFaXbPUMJnvnOmDNG+1IkGMWHc4YHeKVYbWgGDPjeTljkV+hF5XOFFyO0SvHuDaQZW7AyjWp
KAqePBN9hthGvePMOLU99eFqeF/QloghkUKmaGcrk5lWSKAck27Tj0POfwDdmPCIKgcKv5xEUYgs
SFH1x7E/iHYOIXX372GwLsMiXxlTEEf9TFiEIMRrTUOLb2C3IUh00/7F246YBjV5Htuzt/ui6Zy2
EEYVjYVRbZXqzyCOheDxU+M93+SluHYI+vBb742PaFBb0aCCqoxJk1k0Q4fy0nb1YP4PBPcjMJ9K
kE/UxLQdjxWc11/l61e34gggneITRKuqNyj78CBJzr0wrnom01xWPXIDhpAobf4r8HaNHdcM+ThO
iV1GB+ZoA6V7JhkUp25qas6FTjbl7GRkHUN0meORhE/rA1cmccg6FTORBqHTnIixfw1+ZjXnL+XP
t8OVMnXMdRIOQgKZCFU08+SN85A9d6N6UI5/irQlpVOFSRASjeX1kLeGlLaFMWSKzW1Cox5B+QaX
4e3soo89VTw5jSeO2Xx9N5o5kcqrzso3egaIXlIlxgzyxnHtsFarANTPvlulfLoA+HcXrdrHah/Y
KON6Dn/YIgByeo+ZpauH6cFqj7IkNP5N8LLDz867Ootr1d57ZTC9FLYcGzRU1NO2M4XMVLVV5zLP
niOXdN/o1LdNegoBYWX6c6U0sfTu2h+ezpj9wsydZbl/lxSwVDd0UczZD3UOZ7qH7NTZpVR/4/hj
oAuaJSOCmEiA2SW/AzrRlusPmNb5I1vBJ5MAyH5UU+Dpk9n+eepRu2UhYlArzLjZFS5ZSzbuLvKt
8eSPIhC56P5+ZbOvxzFtcvI2WlsZZ3k3ZepsN3hgh4JKbu8O/LJvbnPWK8R7+EY4zjhRjrSpkPwr
EI5R57GCUEYqGW5gy6/WAcQXsN6kGpMg0Dl51YNJ0sWH5b0aWUsPP2OgUeCgs4acN2+oGZCUE6Cm
5y2pNuC70qbFUSb/nuvan/RQ5uf8/vZj4oL9uOG5t+sdhCpmXQCbSzDS1U0tBh8Tu6FQY/kqjMJC
F2+v0FpoF6NxnyMMReZ7GOtqIRgQ6T85mIDPQEX49y7FzZKc/D8u+gMBGD4HoZOeap1mLZ9m4LU3
4Zx31Gc6CzFtOS8uyU2w2iOIWZshGJKGUHCcVcWDlBvZG/J7KGlJrkRwYRMwU4n78J+6gLOwrxdD
hVRuqIGuEqvU9gZ0eCCKBDKJjrn3l6Id2CaZg++LZTAXEbIWm3RrhZvER1SFBOXeUI2W4CEXOiqt
++1UrXQszbUTD8bCN77LVkMJ0gtJilvq30R0b8o5CnlVw7UFE6lUVx7BPBt1BmWWsQmr98OBsGli
57+ZU8uUk1JSq26YdHro874hQIjCy5ZYQBmQE/+VluWGpHgW8XJgYqTNPXuPoi/8qUwLNZNin5Uz
x33IHbUA7eYIj/El4wCeWRDUbnJwekj8W1RYLJFVgekVkwbCIUn429Jv/b4ryrIARng8XLjV8U0A
vwqvD4xovAldSmuULZdU09Th7HuclWWrHxohYUuV4Ab6QpK7e8qlJGPFqVQ/OeAOjSb2AP9cMdl9
JkSxGx7Ua0PYCbPr/O1ZJZPRIaX0TjyP3nzmpcevMKUsVxir7zY/nIYu8sc0lfC4XpDygEUuQJwr
mMLIe1sZ5+2zMKmZo0f8HLYoClTm98ooafKjsLR+vf1P59qbSSpqNaOPPN/ey1IQKDdAI0r1nC08
NQMTQH2Si47CF3kVt5qCDQmL8EEytUmF2HTcdysqWGRudMvFng07fqRRsc2+Sv45hWqQkkoLyXKS
Sw1lwR++rBJ7nRN4ZEtIFatft7pTCP9/KK0kvykYLmJSdnV0beUcllaQdq4t4eQCnkvc4Rfva1sk
rBkBJEsQ2XHbHo2CKQQoZBK+Yuf4vy2KnK4u+Bpu/fapoJJf5cfKFAMpFKNbRGsEu/3/ddEbRDKH
FQmAPM4NWYusSYD/JkAxrfJc24iatcbMxzmxy3pAMJCrRrTlsP9hZRXOmx6Y6SCNEs65to/fMd2W
9B+EKgBO8vHnxgHNwQOPmtAgNpBtGWdKQLwZSsPhEIVDth7COYPi3i/zx5ECyQCXBG12ypveKL+G
NbP4yAqWpj3O3rCd5LugxKiYkghK7j+PAk+9lClDvBzcC+Ms8Xc6M/Ww05qq1K5L0xO4rQPBAPRa
FSHeomcoxXu2RWAVI0hqccq/Kv3CzAKrsIrPUT962MHIuuJuHzeP4VQM0KWpBjr7hP0f4yZd2Jo+
xBiOxDF/n+ilwJ+919OsgAhOjtjljswkFSH2DjEkYn3yk89J69NTUzbA7EYssib/C49RHqITUMsy
nQ2nF1UnMuk5GNKak1uOPAgHIsLzYtn0JMvGaI6hoERbOd7Wu5YowODak7cuqpwXkid2shRDuue8
p1qVUlmG6nkzoho4zYyBRbdtVoUpcV5FOVce/uTkw2DvoLpo/Z+7BxQns7917bgBXjq03x7nzQOX
eQZ3+Jri1XwRA4CLmY+2Rt/bzGxJnhgI18iRvaMlS+50+3A34WLu77eDU1kEEat6Lh4ZCWYnA5gI
7Xj4qM03aLTj40Xsbilns56jaHAZQxu9mJspjv2uOGe4Gc2dIrIVI0nAVguyt5zkd5okkvOIS/G8
jhsDN7Av7pPzfNkytdjnfvHwHSgdj2tzWVtJf03ZSFLKY3j2mbjphFx5Z6yHNQ4hMISLr1dFukOK
lKKucA2h+YKUNtDL9sVa7rVp56O1exdz+pmzWFiZJ48Eo8C9YjhvUz9XpJXaI3VCl2+VgRdBM7Ak
OduvMTbTrtdZgoY+zhOM7A68XDf5DZwRLnX0qpnvhS9ZUaeG+COUUV3FiqpqGsvwd8QvpXpMg6Ut
ztFRYoLeaOoNWw6Np08myok560DWchsT9dRu211Kh4S4GLC1R8Zo703NhzfbOdTiIkAcW3Y2nNIO
22/x0QKIDurhwIVfGpviHq4FFxStEWaJEwyaE8Cvx7Eg39UCbaExENmIBqNjCNkuJrWxTwxoe5HK
HYW5GTNK+dIy27C8sK2jl6AMurce5NqwXeqE0uvgDios6nBgh0EzoBBM5DNIMSY6JY5w3HOTgfiC
sKbpHMnq9aVwZIMR+s/MhF7ZCHTZdGN7jwlTgK992BvYsd7uVhiYbVcmbYO9V3zet+LOliApwiOS
DfCW2IFnoYGS9UEgp3mNHwyoK+dhQEW8pGVP5bLITbcP5ahO6u1FWQJtiD7tJq4Pcq45i0LrYEC5
Gip1mzN1EijOW3eAS2Za+dZ/klSDsvWJ0wPze2qYA7HHedrQGZD1nh/wcdwpCdxJTbB63I0Bv3H4
AvT4YKphaFIhwRChLK43fWHx3UV7b8AfQF4Bi/VRowdcuYUBneLzyBWflcrI/kPjK27XtXl2PxTs
ZuG671Z5dXMtvKNHtJ7NZnWNH56zl/QNnntdAPBoYvyuxTyswcM5KSL5iL+AFICiWIRzsrYKE3RZ
Wjw+OBZpu03AhHOWWJRB6LT8b75UOnczRWSPKbg0ZPtK/waUCl5vPjU6qjUs48EEMc6S+amWV/es
/YzPNEJUsAIV2c5uC5HtATTVpP72y7mw/F5M7YInXQjyND9t86ufgUQLRR1G9v/72bXlT8wu2zo1
Vll+RFQ2i4KQHENd7LIkDLgVa7GcvIxcnE+IFG7CjIefZdrRmT5Q+bFKZamdEPnYWprXM9MzRsrn
bvN++NiVrnD1BO/2oHEChYfFk7tckbUMlhkBZgu2kCuSsxbdx5LN7Bze90VA7qbXdAGrQRfnVNQw
PSeQ4JokCAU8SYHEzWLIbsTTzXntXDDJpjDPiAbtmn+e56dgwcPVlUXofhC4+0/WmXRuwzivYQfQ
ocAqDQYjJYMJAi2/U+ksnjfHevUdC71/x+X8+tInAWQI/5Nuu7GzP8/a3AEDeROTXZI/viVj6XMv
2CoMTVvyAAwX6t65ZSx3X//V2RyrHJvKfgVyOi2OD9AuoxYvIU8hC96feckhh0azUmkCgCukGtTF
3uSxkh/DrdlsNbRajVDcgwIwun62ygLAQs3qA7pEGIBKSkkUGd44kxocO4+itFC3AxWjTCEjHvZ9
8b3pgbZXii+G7IGI9kAYwhssi2/1ehY950F7SyZCntZIjLL0ynok8403rShKUtBUPGJvwTqfxk5P
0URWvTZHw3Gok7L5SN2wCjkaoqT2Bz3En0ZZ4H2Fbm9xI06798VAnppgcj474Z9ZKd7HkpNzNOcY
Vd7mRP6LE6N5AqZNs/p3sUlk3AbePWnCuSc9IRcILcYI2Luq3HwqfhTSEANLs7NooYynk2CniZvf
g4ZPGIqO+949Zd+m9DmD9vg5ngtexHkFMa3p6IEr4aKe18UVhy8t/9J1woAVtn+Q+xcx4WTsSs/S
O/VOL3evbGYAM94apzBNzXMuhTQYeQuiUXKOgrZ3ql5CvuuXALROdLcZSXal66iXWf4RrkbkxR+5
/h/MkvM2FWY8Zmor+KPXsdJBKyfTIpZYpaK/KEaajEOGnON139orSwrW0cAnOtfRyWE0yujROpqm
u+s3+7hqpxYD0N+3eUqyvYZL7FQy9nsybKMcKJeRQowifRZ2LkVZ0ggWgWh4bg/jYkOhwIOaIH2n
TqTEP1KbgjEfMxe04bg9m3r3lNn0zsquk8mvzFHrW4fd+2HRUZQQIGSyQUBEMM11BIvwbJWL2HHH
g8uew8mrtt1JFctIaysDhJcEyiGBJ8bs/ZW2BMMtI1ChpYbrIwud9lPO3DRkZm4UwfGdKv8ORkZ0
StgQT8jB0sBkry8qCLCUmm45FbFeGK9Dyh+VF6EqKw8WEcIbFSttO1btclHkaNNux4wtOyrN32Mq
Nk6yfRaIGldG0jMaMXaFc2p3Z5F5np+PUX8RYVyY9VL9rBFH6bAOqdwKCroa3gJMteaTIaIZfALB
BKgKG1KUeBNxHyHTgKHvrZPByuhEpX4rZVRibnc7izwRw1rZ7n+iB29a8zgmrNB6gZJ4mtUpbyrT
FkGK/J1+NKFVpgzeWAyIpBoSEoK39ic7wnVDhcuIEkB+jOqHlhNtP9s2p5d7oh+6CW9M2StExKjt
RUa1k7Xa71tqoPdEd5Rs/8xobkLo8yry8y6BuyeZVBMjnNMN/pVB2BVI5ooBgbpevE2ehUAZ4yO/
a0VrM/Zco0JgkWiAurosOYtWto9MRVPXZq/89KhxzuXTed1U+7yi4YCMJ9/jwusNoHWOms0cmJV/
Aoak2OOK958UJhz0RRt/YF9Mym7ibZ08/lVOVNF0LTd9xEj2ngpnz6+RrrZx6gnTpKdnnkIuyVts
sUXYdArDL0hWJPs/Ah2s6ewkNW0Nd2ze7sSE8RXO1ZtsyCvuwhkH//19awQkaWntrhUTUQcujlZj
P1IG96geAtdAaA7dTiYkIXDvIiksZsIa537txbFzXv0R+4VBmP/Zw4OpzfgEwUxkwMxBwYuaZoPR
OX9CYhjUPMiMn6/Uf9OV3WjAYnj4ldSG8D2SWEXSyP7n3r+NSVvDsQ/Xe1kj8Yx7rws8X3vJHdVe
0Ks03SvL4gVLJxBzSL4jtYNnULNOAKX5lVt7iAf9iIKP+DPqyQGEWZCflrHnNJY5vwQJpLxNeb9Z
/kTzKLzUXytDLsuIVQUimqM/7zD1qgrpQRJufFAGo9nGFjxFlXQzj1xodyJDlUubFS4gPdxN37Bo
I6DoymqcRs3uMmRSN6ySW/RTiPzje0jjNv642lCJGMSboliab6Z9Pxis3lwEXnVNJV0kPJpeXJvJ
TlwqSpkIBpyutJ+gFSQ5yjRZJ/5LBoSWRXqKjLaRgT7oJUWmtsrBMHwBXc/2HobqqhNZWEWiUCDr
Zao82RCx5DEU4KwDCfKVTOB6eCio6OarHsY72g4kdRVk701H5CtEybuA8sWabIroEbwc7eZ7qNlu
RlrknSPnUB0iGJtcY+63ARdRWgepk69X8wPDr9Y3vOdETpa4QPjLzTTtC4PU68iAWpjnBCZc/w7H
IOm0Daa/cf5utJM8KjN7LSqbxGYlguWiqyMsC1d9oD+5W4TxQ2OqKFrAmjdC0BPxm1FoGFlZgmJl
DbsV468kemDaY6k+ATfFBwljGhcd77UH1FFo6Jw4KTWJv4TTtHPH94vnO99DrF/EFqAMJ3sdDdB8
tAlgEnd6omk5Oj8MJ6VkdjcN5+lJz45dKDSU8pJnXkzrNTDiQ5cNVrGc5j4SIRRqQ9TvCkCTAtZJ
NxW9MJRKXdhxg5uu5LlO3e4b78XSyDdDrBwjKm1J/aG9J9CE3KoOmtA81BEbE3IiD+iVpIVrfn52
wpcJhNdz30ipyGwjBMrRCb7+JPHorNDz1BqCP6ClNNw1OpMioQEJyvI6nEc4ePcaWufgdoqEnZuo
XR83gp+xQRKsFh1XR0GwPj9aZbDp9zUcW8R82kqauTbGqTs613DJgNtFfL7skPKRfwEzy61B/k5R
KuGFuapBHWpKWP22I9UIx/URnhk2rbsuCbDpjoUuNmULVzkfotjlKHd0vUsOTaCMH2d+OQ7NuL+K
DTRPoZY3bupvQMDYlJ4eFjGkzOUt/9ZYMFNgGgIn3sAHKjPYHHL4i9xvOWYe4zhCPsoVw7BU5BpO
RMHaOD5WUfvpRLaAJrsP6eS7Kbq3QIRf1USSsUysGsi9tIGV9AgKnCHVZQE1T460CVwcJcJYUCfy
W8nghJcEAqcBkZ678cEj8ibnf4+ACHheVlTyQog5HZkDu8Qn/PN9czvDWt+qyQW3Eo4qZWwT5UZB
N/mzbPOZTqRbWc9lwOtcGcLUOqE5vJSf38aL3fMMCgkF1QcO3PusZMe27jKBjQCfrkL8ZhDwQV8S
BJIrMRhkmC8g55hF/i6x7kZpPGjA9G9ym6fUexY7ivskF+51qLW6pihJozUzobI3/JmKqQj0Ayis
rt6Aw9ftv7jse/Yz+B/IodL5k3gXA+iRAhdyRAmQTWuNHDmOOfrSA8a/33k2VJIkBoSGAXX+fcC8
M2q5v6SWjCJZXZWPeErvTybTsg5kXr8Wv2b9NpasX2edARDCt7+8tnlOMBgNBfBbRlE+HsRegIWM
3D0nq+JATf5d8aJxfbVHFdhLP8HdB/KTK8SSifLHfyBQpAfHaJMVs+neLT2QL3t+TwlZ4z4lFjLS
VX7yQOOagbzS+Qw0zs41XFaf10VIAtRu7W7zvdmdKMB2rMqx/yM78+3BilOVwm1tjwVo69SlXH3e
DXqrmGf7kXmXA40wCp33I/l125FF6fnsCArS+a6gpU3xQliHgOFeWRfY8AqqzrxpGptS7WCxVm4k
OV/nkpKZ/cp12Oje/P9aL6oD3H5Fe5EFrDOtUxgeNQoNdy1FDgZjOYxUisGNthn4DEDeQLPdC8FD
8qKjWps39pDKzSvGMF80LyTsffQC9/TLuS+TicQVz3MnNowN1FQxfnAco1ZZ0kShbrTak41TQz7t
A3jLLk4l1iwRvAa0Wi/NqNoo84+EZUIG7wW7DQ+bFFR7X/6vMK+0s3mVPb7A7B4i/i2L4f7i/ZlO
+ZszWpg68SK+cbJUxbf7Bd7wbXrHnPSLmx5Zm3GuPeD8pvyyFVtbSntOxLeRW7ha4Et9c0FulHYy
KEetVsWPlAKkmf1gQx9i6J7IoatwXEFBMHAWBsIjdNCKKr3fqEVTA0Yq3ChEoPspkK5p3/1CKmpL
EzGdj27K8XYwET+KA6a8kuyStDeW0/90kNvoAuMy/DKX3piNFJrGhWW0tpLAtnBuDT5SrbZTDAFY
dsBOVaxG2vNv7gn1jBTB5m1gLd7CbRfHF5f4jOvtCetH1Pj9wQ+nZ6jKcawzEhgdBPmvEEzVm5YR
YqJyzQXyB+VdEyJ4XLekoLo2OkLP0zN44rUfI+appjOKBSgOrEEOS8JhmBO84II/auYMMlM4g97X
EXWGak+BIAn/siga+suYizT3XZNCoBpk/I9I26NfxYvtB6Bu/5T/QZH4OEeF32W28SieEnZ+682P
bHDbLq2DHP4ZgsyHFOxmVL9+kIDOoBXP77ZH4946a4u0wgtbsyQsbRRbATzuGll+OcgaRChWkJpF
F8fmjDZbZZJ4ifkklNm6aV6RP4mJhIoSMU7na8lyyFnl8J5YS8QPmiFSKcH/jN9Dn2GCC7JqC9Lv
CWvPejv4TBa9pyI3hCfp+wuHGlhamHN9dxuNu70bcz2fAFimffqThWGCOrMP/B+E95VZZ0ojdwZH
zq97MiqIkDIAiQb0MOL+T8EGzUA5CRWVafcelQT9XoqAe/GQ61fVpKSCZoyi5+aykDkwyG8vF9Ke
ai51EO2ws/HjW8oAXut1ElPhqA3GhH/o/VAGlhZT+0lpXBuUWaxJt/jUbBNVIvaGm5ypTEUNGIqA
MKevpPTsgUVlk7IFWMqCBvZpl3RvMcq/n8bh7lullMQDVcReDjIgv3uytmvzDXNh4RnolBdB4taV
vP2ai0s4LQfcI5Ru35ozTrZdIftHO9npGIJaVOOJb9Fkp5fIKTY1IIpHJz9AepR6YX+Bw4QSwCsf
IhKumlY6md4USc8snI8BIiTazmIaf5Fl1AZ2nczd0B1Sh2cYxuQryXAK955pEvVmTerxAr6m1LBY
HVNnCjnzg3OOkhYLNTcBRxCiGeK7Cn48iIDOa6IFtzL9BjY84bW/uF9O1OuQcflCruMuo2D0vR9M
ZDy27eUTbsRBqUpD3xLFPhIiy1T2tI6WQUah+N2OG+Ktsl84xw2fm00KwyjJoFwjJxh5+3exs1fF
n+jgnXuP8HYNV6aINdLPj83VxlXEgKCLbek+Gjtbj1Zu3BkS2Arormm5EmsqLFA+JYXRk/Ix0UrW
YahnSfn2fjTf4G9urJBdTIHfRuzdLXpfxKo80HdfzwAF3WV6eSymMRBz6xTLmTE+s/IGhbb8ndyD
d0XQ3dbXsEXSfSe0Q+X84HUCh6Tb8irh8AkfVA9Za+RfNXSxjL/nSspvLe+5s0mompYfWvXVXeon
XRUXBqOHveP9+3OYifRkkyvEm6m8uRryvjPGLSg+oeTNGkqPkEmIlUnXevjfYC42puhTWrDX0CTD
Jn78Pvv+86AcUaINO3EwPETm/X2ftevYn2mR+ocxQjbkOFwgF+GRAVbITq/EpLM4dvibVwvXUYFd
hpsnENMtcnQzfvbmsHWafJcThxCz747XuwkqMFKPdEuQuZEljAo4erXN4yLmz5M6kAMcQ5/M1jb6
E/sAXlo7tgOrfyHAIdeM6PYLLZn/THurgQffhgwjh85iHrUBQNDarLjspCd42H2HiBqZtJZyTmnn
LD1KcICGc9xHrhWptgKrM4s0EkWyjIIeyEUEJlB6BeP+JrfJg1rOjRIQ6ndEUtJgZerNHFyewAwA
Q+nfWDdYWGPjShrrxd+hhGn8OPrZGPN7BqjIXVMVSNaRH3hI4x2PriTR9bNa+OfALjrZhOJsFRL4
Pi2Py4Q5k4yM0mC8QyEun2bondLWerc80amiOq2bC0PVMIBsF4YCaLJnQy4z0MifvLT+qgewZzJV
48rHry+D3rZ6GUkfGXi/wDIiqVYUykdDHKcbMtaQC0XD0rLGgpJVMd8TdJeOSWVTtJtVdxqPa0P6
0ejdbtyFUBL9GEzKIv6fP/kVaKhksb2ZLlOZuXL225RQPd83lGEXj7rOTS0ykJ7kCUzbjKZ8lLHf
pgAnT3i4MJMNBeN2HYeH2LSd5N3QnoupZxiGlBLVPu3A24GTWcAymysa3xuUZMHbYXNHjR/j/Q5V
m4J87nR20Yi4GeAnqNNw0rHr//E+cOD77hjXLlhXV6yjMKR0Kfh7hNEuTf/stTLFohFLboVkZ76h
lgG3NZnKlbsAM6u37u8lAr9R3C9Mch06rFikcgNo23KdtKcvRfyZSSMJmXXoAS2XAgX2OkgPwWlZ
bVjVOt5hPP3pNW/Gg/4WLF+II/D93E4Xvg7gLmvZhz1K/+18HGPTPxJV+laT5nHK9ymb4HuTBRaK
WOMsCpp6VwsuE595e6ny13iFRxItpGn05V0FmlSyAiXsqFTcNn7bUA7MtjaLLQf/crIBPOKZzHPd
blofraPSVxbVBVs4nhGdbF6t7XQAo29tuFCMX99/IuZz09rYK009LvBDeNiNa2GiJRrinmP6HHM0
72oJJ4QPZ3bsNZKbVD4Wkv6t87NWxH8WdAgb2jwEfhsmGIbw+dZMu7bEEU6fhfGG7+BhgP4BYPdv
BloniVjPu7ybpuaThI4XYpWZou9tZYnwuerBIvY8HEyT9Pb0pI1t9qctmgrvHsntEQBvtKBEbneG
whysoInI7cUbxPpk6vdKfowNpSTfrcKMWzIx1LJi/TdrqdyTBHUHY2BFSbpHimVpB93l1r9CgEJ/
HLtfDIMLupSSdALsW7Ej1utvCfPASigkmKjp1WQnNNi235WUzplUuWUuXVPXEx3kog0Mzotf5Nqs
O4hrELTs+RbLUKVn0Yodfc5+7w9L42hFVSimw31czjozH+DyUjdPfprAM/t7DnUN9WY5iIyxy6on
OkV8iO+l73IDUnsbJjT2AsTqN4/9GahaT6BLCxSPPQBc+3cRxD5uh/kGR/AMJTCJ1fj++6VBxQc1
1DaeU8YRm7PLp3qooJN/QcL75ABPXv87aN1GInhXjhtQLqXSNOnLCqzKgUM8fPDcaZRcnSaxG/FR
epl0uJCAyssi2ZAk1XBIRaTgRm2wFWyjBJFGSw2yEFMD1kXHb2ajSRIMxVkkmp/7NpJ12u/Ea44b
vCU+JqRRptw9m5pHlS8Vmj2E14lpzlB3PAnuWz7fOcLSxBT/33fL7x4bO+8Kj09Z5l50nE65EKok
rALQiEIv+nix4qNpaZ83qMDhXOz6f6GirS+m6+Cqxy1zegrAEnvOFz3W79LZTwamiX9ivtznhDEw
xmMLiRnabigO3eyObdMD9nvlwz/lFLSdA+E8MTUJa7BJ3b9hET97cjWhRkMjNEbEJBaTNCKXo0Lg
DeZ7GdbuRozJNYM495MyKVhPtK7Iew+2Sz53rFjkPJK9h2oFe7HJWnvbOHNwNiAbzCqhYkLDIeVZ
3FxG5vq8pG6hCHP0mnVIK/nnI5FdTjm6FUWBzyg3/p/mvDWk5lo0F+2QnCJkZuliIvtdur59Z1IT
3ReVEv9JXeevNWYLUctYeN1gRfEv484sA5bOxF00i+ONr06d2C2JtyCyt37QjdupsL66co3GAKWX
eCH92Q0JfhTW9s+adst473FXZuBZa6blYvjLmCYQZG6geJjxZ9VQU0tElc27W6oGeGu2iHmTog1B
wqp9WGDH4NRoDr3567TE/AEqavEzT9Nmm/Y19gSqWAdJkeKb1DJXbRgqpHu6cbzcxmUuaKZ2WFQs
Bb70ehC0NpB/aTa3irdsAaVF65yzpP32VC54J0PWu4KG7sMuHIik8n4BXzjv4e3IECcOkzQwz6hE
aNwaKqQKbHQiBJPK898vlryvW3aE9sMt7wCgCkkyNH0vK/ansbq8D174G259Mv8zaoGjgyXcOD8n
i5mD+6+3ayYUIGP6mF4MUMg8PFAWmW3D2brLRfYZQcS8ql/VnwKoJmhr6m2RYg3sAje6xiXWonXG
Vv27iy64z8Oett5ChRM1TLzjaKpCcwgzN1vborwo8+FMNzDbSghDQ2ZZWFxK/cTP1NOWLLMnvhIV
DLBQmgtm0oFdqLAkH5fZ9UugPSwa5M0R4iP66ytTuppxkeDCKNaXVXJaCZYMU3v+uR4/kLrhlWkK
7EjgFtzIXOUFnCypG5V2x8OzNYE8W4R2iQQdJErKAeikuYznDnQD9xra8trxO9rbzDIcf30aifXW
6PO58tpBiOfVUJxCRvDLrBOLaIR9mF7Qn0MVJ/gfKBfOy30xHnpZ8AjarFrmSyF5Sf65enR5XV9q
kqJLvDuM8m7DylG/UJVMUHAnKa9LtU0U+JLFvrrz9elXj+8R9r/bWFfLWRdkZPr8IR4jC5gigYOu
sYejGaVizqme8rkjVBx1zinS7o8Wa8Z78bNiXxTGy3wl/TgH+WGHjcDJSNEYjh/5U5No8GPLVX7c
8s7B45qi3B7+hUrIf34p3CGYKgKThRNv9GflHC6ohZYIo+GHIqkp+eGFLDTv2Z58c3agMst8knD5
3f0YTunuriE3hgW7k9ijUFAfcBnqExNlwH1yDgXsBseU3u1E0+Kywa4i3C+OufSxbEoNwMNgjvMD
R3yTMTlyrAVhMQhe29g7JYih6bZjOmPF8s+ouNmKo3pa5OqRArW6HXSMT7jXNpKkHpWg3UeEeXMh
SPu2+O3zaZfiVVXu3Qld9cFFACLLkDI3d58qcAdVpQZB4IL2Ovu0z/gidP9dboAOuxBccPBmjOW9
t2XfrrXKDXEQUQbBSs7CsAm6sijWHQZg+6iXID4VQqsMXQS9dAye6zP90eh8A2TSHw13QWQR97e0
OWGTGOepnbkVvvNwRhM6KvTT0mu5t0JBfA6AOpbQIob7FWCt25MtztfdxlEQGKkYrHJ+VCgRjTA+
xGTLDhKFBSstskcLnXtB2Kk9fqKx/97UjtI/Cx1nbQTOMFjJePChjQ4FeXdnqSwSvj7NIbspC3eK
/3xinLmd6AvrlCapKG8Ou6N6MY2CcKtllQJWrDgkfE6UpjxgmlsQxBVFbMzvBznAJSqZNQH46BLz
shxL7f+ZY+qDbWiNOk7/d6gULkSaCSlCo0a226bWR6PCCoGZlU4Vu7+R+MK1JIldXodlF3Y2OFKS
b97dvtX7ZD3whYophZaoKbLmZJ4hRYqG6DzlWA2ZxaX7hJICmPJesh3IIgII609W0zI1fgjs5gmD
ebo6ytbmzEtSzivbSmlZzZUF56octpfirvQCfvsSdBepYpEZdATTy6rPMynq9zvlqJd9npkbrZ3I
ZHcxYhuF+PvX88bWPRD72iZlSI1bm/y7P+C51PSgegHFxB20MCh3T6cBmMcg5iXeVs1//+zoqLSK
AkAQBEPBwDLAgsV2T8FxtbA90m1EOGeFs58OGZRkHt3Nx3A6N1umQI5qvuYansxOwTpf3sPZl4su
JmfR7W8Ke84s8gKLomlzwMV7O23hk2RzA70ZKG1kA3Q4NWvE25NgniVZANlXMQ2uUCsgHzjqIZRB
prk4in8CfpWnYakahKbGQvTpYXHJ0cpMRNUXiig1UM8BI3+8H26+g2l7gXbXLtssHDgzFKuJxz9p
IdU/hGSKkY/+MApA5nKc/NrrPdunREzdg7lk3Sq61cY2mVnc07+T5dA+Av3SjxfchfvzrfJ4wOzJ
SH1B5ppIyBc2vJkyZinTZhehPA/HfP+WXlfS1ox9gYlw9P4m0WF1mLY3g1O0roAj06W2B6TURIwF
qrdvsz42kPgGJoDL+EeeKpxeBoS+WsESmaDT+0G9+RxrZKULzeQHYn+lfBSebsxtpK3CWFFV0ILX
i6foz+6i7YPh1seNFb3GUdDMFQsIP1sfsROkCGrw2mMxOIedw7V5NrvBbhyyAU/dI7vDS7KAVXT9
e3Uc8zT4l/0FBcESXcBCI7PSSo+hQ5yJs6af0Oq0mno6eWxaHtOQ0SIv+L5Ua6bu7dreR04bepc2
7wN7FgLda+qOVxFs7q4EhyKOrLomcMo/UQUG8G4XCpbAKmx3m1rATet2dSGfv92oIdy8qDJHP69K
34iiL6RYMeIdQcKR/IXE77edJc0JB+17sEQKRuJmQjk0SFjZODDTay+tGNBEipOQ2T/zaOHCRCMJ
sMhOx+4ep7gZqbx1aqUkYhPTXxYEwsUr1xK4rIpSSRl+fUwvrKLQTcUuph04d67qCnbqP1tUryUI
hVzh8058TaA+rgGHa481kGW3CgdZspdIK7PFFcjTodOJ3jYK/mZ8TxueXC0jFKPpipM/H2CZrdRx
9C0H/30XkQa/MFoX6nQgfOrdFuAB6lE9EMdmuqF02nui+iDD9LoyMjH2tS3dM+B28B/0EXg7OEzD
WhighjGsaTUAlm5TNLY4qb23m7n13TO/SuVyzGC0lIpeqg8apNFsBYacPDCvLIbzba0tSuQCDZQQ
5XHdxAReJ46pf4vH3lPJBFkvTxWoYLHILqypig/bCoDZrV6g0Wxo7flxgtAiAzdv6/K2+/RPwTM4
wkLbKjegVGI/bV0g65PR4Z5OSECdJ9+e27enMmqfzdzANwub832eLV6vETELMn+39ej8sCN6lFWO
CYy2O147fMBpFRxkcGQeVUTdTkE9ArgaJxB67vg06nxmnfArvTawhv/ToMuH2qOqD/Sy109nowF9
WhWd4nfthpGPAQaMIQsGlu1BWdOHXkeeDpzFFueGVRqUdvY63I4zUsVKafoaGO7cFYu4ZkxKgabQ
wZ2F3sjXgK7drtrzPfDpnaw4C6zjEYeTtqv+qAx1TT2U7UCQBXBkwJk/c1xW6ByHK/xfENPYxPLv
dh8tLJ5lKIn+pHyQTE/PyDoprbNRX0rG+FBldEaP4rsjrXwlxdJ/DfNMlh/FgPUt1deJk9V5bE8y
3iHrnCeXh4HiUqtzckYgYH3SGCwKh4lt3pxqnWda6R6ls9iHPSx/YqBXv8636gsEHVkiaawBKWhK
Yh3FiF2mQGgE9JB7OhxXabcnRnW5zwVi5F1HEUBPbxqBC2O99iBx0UlJJEOsC2woin++QdSJlijV
/tfSu/g5Tt22c6Wdu6kKyJ0wI5WgK2r/LThrAjSvZhITWrvzGAvPV+9+kf1FmkUBXZ09bzY7FTC1
Si/1PTEe4Ha5zrhHHwiHua1i7CSa2+sqEO9hQDc/COf2FvQBhlEPiLRQxWRMvFrh13ftU50x4DRU
oheE8/ZNbqEP2RX2Sg4mEpRgIXRsMo6IsbAuQ11GT/WiIhvIeaeyp9D3vqw/X4sz+bF7oTAelQE6
hdVVpHeXmROw/X5tjvOEGwl2dmFojFnY/EbHz6X7ogoT7jWlaisvLuilzBc5xIqSk9kweITo4Djt
pdijUkB2ikoEbzhlYEKtXjTS4ucpIv3Kuyj4WNSlGFKKBE2lLV5+QkYPPRiswMmnwIB6DP8BV61z
caGpdE36tGKpO9TKZW0hPS7UQZwJLEunfSfgstmqFABUmkjTx9/43OPDmLKndSfiqLRC3coVxXHy
csn9VfHc/vEhuRwl7NhDPlHGylSUXrGAsltQL7OgpJJHD9zo11w0iA+4L2AzrkQYd5OJA+Gf8Dad
YMnT5PIAXQcgOJKyZTDTvIw23tYnybmtpiaL9njekq7wlCbip89wpdL8CyMgVfNfN+jWd6jI8Y3t
DhaW8/yIns0PE+kEZ+ej56MofwZF3jmyybJFV+YYTidDWtONayk6BBXCXjWAJjtBJyn2vTuMcgUq
qATXxQheeNcBOpvWMz6kvPHGI4tHmqDwvgsf/hIbaJW2MhOpyoY4ezwKndMCZ535uVw6o43GskN0
Col7vk2bERtvjWDSCepBskgZfBKZ07515NWZLlNZ0RwJdXH3aW4BQpRM3s7uc7TCe1c1FVcjmjVa
dpXP6RwNFpLpPRFXDELpocHosioJ3dwnuB0OaG9GGE5MlgfCQC22aAaRNmobUJ7EoyCoK+mhnqPW
xcH2HboLmbfdqsKrYKV1X6vvICiRHfF51aOZHof0FWfMSv9L1QM+AOUYRFkdxPtmzc9G3ddzke2Q
7v/ByBDWYqnpgWOoFLxTttiBJOLL22CPVN9KDc+jExjsy4EbQt23XGdjqQd0b+Un9fa41yxA9tP5
ZkG3ZaSmLZbQdN+x1Ye5wUK5383w2gmnz2Sq6iQxNdWhDvV00RC9i5ngfSEoK5pAc8zTCEweq2wV
cpWrr5/HcAWu3UpNrZi2UR+AcanpyRL5YmJKUF5Ep9faQILitkXwFRxT3kPfRWAnX4b4huCNii1B
ay5GZaptLZkNrnTSfGaZEAffWsQcIePU+MJ/ME0AJrZ7mSMVQ+0XJ+Tx8MeYMe6+N72X4HNZeQj9
A+vlpRtx7/si+MVqZcAtLspwXZdJrZQ3K5rvtqIyc5H5Rv0UkvMLOy1L/VIsH18bWK6N7dNy0Hlt
pHNYpApY2Zhh1GZ6z7sVgYAe1hIhrrQUIlhWlGu05CyqWSju7yOG3lGr2XwBqcjh94t5UQGuO1/U
4z6f0Lix043aBIzs6B66GPgIYtWsIEjyJjEtwDwWpRMWazYsiM+FVjIhvSUxug17tBXtYAUtwvN9
CZpaJvSp0LvDeW7o2WjCZmE3jexJj+9P4iuzjWoswQWSfxSjrbyTt4HC7XHReMvgzt4CfBxjHOY1
cXSpba3tHsqyjntvABMq6eOIu55v1qW5gEbqMgSsivAxO19vGf6V2hsl/SVYkCCGDf6XTwh9C+hb
NsWrNwro/aUbh5lHAWqVLzy2Zll/B+na7LXWN1gTYCTBSLTop5R61BsYnSIuG7GwTItSSM8kIMF5
+mQ7hD507HrJlp2CbhGF16gfYOIkxKdHCWAWpGzHJiljrYnY9qy/zIxGJT6XmvbONhXjMx57cQrS
xTtm8n/NkWYWlhHb3wnyd+Pe+VHJA+FqVIeT2vjJFMUo49m203/s6AwrLviFDK5l1ZFDrKz0wrio
2csFnDDHRA7NBB/L8SYtmmscCw8N23cy/J+QbJJ2niYp7oU4QbAXVHNxaOgr6e9Ex8i10XFvmM1X
PfPnblC6I4HamXP2f/NbsdRZUTl9J9uSyF9y5A0OaQsjfpANuGj8B1fwMfufV65V0hMnH6VpNUpi
dhnPXXbBK/8j0yKIEn2z2nrdbPPG2X4ukeku0hcyFzEyqFCXbaZhhrgOQwzDboDjRzu8NN1PJlAj
qb2B2w7edeBuIijnYA+WcdR2Q0KfYbXR3fltMLm9ywGqoy92LgDRIS+Vx1DuqOpLL6KpB5XyCKAS
gbU2tEtNMrADKAHdlGqxbajwG5rW6IcCksv9fVOiEpjCe6Dga1HFusbBaLQsqMLKMGeCwttPR59n
MuC29y5yZt2a9tWxSP3mGRsDREZbIo23XF//BIaAo0KW5nSi+Br6sU22++s1w7OaC+hoqHlFYhXN
rZihMT8FfzyLYKCoPp4M9FCVKHk0exkQ621oL/qoduGXG7el/F90rgsT+uKGvns8Yti4RpmHtUBj
gnvnVAIkTJi3rn9p7ZvWlJB35Z6MldU6+CLSqvP+e1lnyamF5RrJ7bw/2CXaoUsS28zHV7gcHpmz
FlRomXTrkuytfRB8sIeZwZFGgYn3mYOv3K4nTYJTVjwkZdBRXAIZbj0twLlrhWyI9FcaAq+hCPOw
NYqcsh+E1Dk3e8POx6l0lXPXDmHP0v34k1/P8RYnp9PtzZA6UF/rWqWhHUMrw1W6OCMa75AZ++1c
8UEQtqTIrJdEjhsi7bH45AXY3++I1r5SG+J3smqWZi77nYlqqK9ugzCZuRD3bOdf8uM2Rj6EjdC6
eTpYXq/sUeMkoEkNUZXEiVjwfneVb2HB4ZoOgvX9COddnnIfWllC0tnhERDIKzohU22aAIdpTRGi
HfZ0mb+GOHdCyjThUFOtvPIliAb7ep4wvARq/pluQQKTurF2ifLif0zHeK++aT9A7GXX34KJ4wdw
FYi1byIbXRsoAl5k8FSLS2PcaWbzDnK4CohvWWObhxUs11EYZCMLcuYSRyjYtt4Me4dJUNNLAtZK
3YvS3pDcY3YR+SibiuZYpCuvptg83iYbCFtku1P1OIuZEhJFOh5mro/syuPwbEPn0aDWgKH8h1UE
dDcp3nAYwdX5ke3FqWc2NyklSIPpglgKL9f/sx/1bv6pThmvDg+eaAlamQHqgUIIi4FyZHmSRrhW
jE11v3Uw873XU4NSh1XmTYyr5ibWsGRPKlapLv024JRXe8GK6znT8mxGKZJN9FAxsaLHI54vlFH1
aK2IiJCEPRobg9qWqcSTX6Gd+YI/4uSF2FlG0Yila4IXh3I1DdydFavIFYdfjvFEN2h9WBNMAwcS
1+rCGYU+Mm7Unx3y5kp9A1gi5IeT5yqmQfPrld5bUAWVagFYufL5694JYeC1AEuwTYvitA7CB4Xi
SemIgsQ/EPMvHu2SwI2rWjaEK3yK6eBnvo/vIpbIw6O3ugNvbLWWtuvytqHLSHx8Q22uY0lovHjM
LZcvs31ofcUJ7lZvLEGzQbKGDVsa3h5lN9eLGKyrdDJ4NW3uyktJywD370NeBsWKWqIv6FVh2rhd
B9UhHF6eaAeRBdc8ChLjHTTSJRaTbhmS5t8b8NGSfIZri/eK1+XrowsrUj+HOsseS3vh3Kk4gzyV
oqI5SKHwMh0fPguLxaDrELAHD2rDhaftupwWgrkLiZJZ1hhV9/DmRIXhTJkGDjglz3+/fZ3FEfPK
3wHfbPQ+X4zumzIvNSyn34Tqe7dtZ15gUE0gd+4o4D5ixYEY1+dsRReQuscP3vVnzVD/38rOS0/7
O4ZANSmiZHOZykP/Uu4QvOnr1dVtvMhy+2h0d6rMzh+MSwyE7hrJGeDNhl7PzJvVF5Ci9fE09aaC
t0Pr5IRm4FFgVNsXowhwa9359aA7G6NQcPTYhp+awlQXAX1BonpZlFd2MjOT1I8EI970EB/YL6UQ
xNuL5/sS8v2zE+L08olZLtokbirzvFX5cuYYGkpsuUynZb4TyTZO0ZkTYF4pcsRORnYTJW0PN3cg
JJ/3XEk5apaN7eNzoxPDMCBb5zNCi+L48E0LRE42bCCHyXi7l1+wsviyepGFY13m7fo8AetsrLQK
IGDxUxd1L6pewGQWMHR52/FF/aGf2uT5+TDAM7JleJkYv05tYInhUmeXybONNyT1H+IXUnYnVqCl
77iXvFiE51VhQCxKuI71kJWVhIlsWXUGQKGepLy5bSs0OJAHexSAFZvmY5oD+VN8qF+RcGuasluj
NcG8wt1FIH+MiWEYsGlaZqRbVbtONND6olF2yt/raWn5zMRsJ2dh7kQzLw2T+l9anzZ8I6DHlK/V
GQD5PVh49CYixyjR/hk6geGEgctq7AENWgzpzcV0ZkqliY7e3h1dS+YleZ6DsxkJ9yziYYSXlRRI
xHHxT5jEYqLqth7ibu2Ox0NZR6pst24QqlypM+ZwJrAsLEjFW+E878nJKH0+tnCMvXRT91qazcqL
kkC+lYzW5ZW5OHUbFSoFD7xftxNGRDWlfNsXZHuzMSS8TSHA5UEsMo+O6Nw2ZdkA8r8RnP3LcTxS
EtRD7Qxm12aBdCiU0wt9euhQ3pOq3zL6IVohSzJmRYp8iNm5Av9lX58DlcQHOvRKteo1214jco2F
YfQEvXnzbnPjjASNDj64RiIGg8SDhgFjZZBYdw8r/cUmgg5SIC55icomNr7ut/5kyP+DhzP+JBsZ
RtdnngG4yoCfw1ulMV/I8kEk3YRp/mryt9xqHJdcdmLMv9RuwibYrmly/Q4leh2IhxQGanDQEtzD
HkmWBNKInKYHxNK8VV8q7ObI+Q8Tbb+bVXt4VDub7+Iec4v32bvqoXlrETlCi9xGD1Pi0U9czP3g
rg0d1EQtJxbjlzQ22YByiicQvwqv097cQ63cTLBVQ2Qq4nneoQqIiio9z63dLlNT1K8gC16mQjYu
E26Jt3Yf44xqhl+SZIpiuVonMOQIrysvIO4aYVFp1oGEZNJrkX+jEuK9z4XEamGAORMEDhZ8TyT1
HN/nfRV8jwlAz8eODP1PRtXF7HlwaCKvcvRuDd9iHyaE/pUuxiFUhoOx50Slz3eUqGmieSnN/vxk
o4LNCx/EZjgubVoXn9UPZcH5Pl7aefQJd152cTAweiAwP9dsviELHMDpASmvn4nlsrw+2TUBQ9zA
GrBS7XZyv1x3OJZ9apxZf8tpfry+czJjovyurdIiCndA8kYum77GAKZUerhdBfwiMAuihmNOVtD/
crQT9Dwh5uuANd4AyY7bGS84CQK1oITHV4EkV7NosFsz9Ada5XXdjQLHBbzXjSUg/rQycKexWAEY
RrHICULXlk9JEWPZYomXR9MC60RuxsBdKd9YAhiVDiFoiYLayBwv4Vvff12x7260jr5fX7qzztMJ
kv+41rU9h6ViyyB49h65RFcKTICTRApgOH3OkLCUglRr8rCABe80RVEMAHHA96W2SYSVfi9/YzaI
um4yYOOlUTHnUHHSNI1JpugOTJPjYpSycezwCQqiCzP9MQiJ4taSKpyWqvCGHx4+34VPZ/dcoqHH
OIzH7FY6/9i+rrONRIMv0XknwPotPCZ3tOr295bfGb9Q7c/ZqV2ir1oYBWzCb1jifMOU61F49IcG
1MvHE/SPJ6/oo1SFGZDfYHzDqA5+Lj80+/NqIqE91Y/5hB9lhfHa5q4/yOBph1bIfbR4KDc2Oq+K
IHQc9j/Vi2AYGLMzhgxwWw4yuji0qECulXrXd+OPQpF4tsnGlG8DCVKwfHn02wABwTpvIE0U/1hd
bgi5+qieVcGRmWWp8HHOqFRGBM8hRkxFRyoicKaC3D29jyfEJ07JfiWkQy39bOt7yYpAtQubfowq
J40hntCY7q8888SlD18rTf6FUoinusWQvvwmK9LGPWt7FXGFz2IEV2kQKPTdSQdM44VdNXAwSv6z
DKBCnpDRuwKEpMc5qTFnqp55Iza6rLLLDRFr9lJuOenpg9H5qmVt4mzXHuv6FO+KhmoMWRGjz1ci
REfig9GYKJpxcjyuo3Mz+PMDU5oZPWa9SgKI31y6y+t0NA62yT9qEktc4zCHSgAznilK9MmXMYFF
VbsdWRahJ7nHQeyGP/lje1cN8qsfxR8HD/xWGWrOuwn4fbhZcKfU5vSrlLE218v4Fd49dXva/m89
1XWoy1FEkSAyed3ErConR8CHbcyNywGE5128+K8SVqzIUYwRR8aPwXH+MT0ecXhnlEyN4XV9Zyo4
kamGagDF8BAswLWi8CB+4K5IocLjFRBwUkZHEt7CQoLVBg9hV1kqvkcSVWHAXE8MM6MmXbrxVUiB
U/DGj/HF18SiRr784eKO88Gm/4o+XLJnrsrd81c91RNGIP1vJ2QY4i0mzivptBIoEhAX4hJEHc5L
kgdmduig38KiBS9GL36n0OGBEJHC1H+2gqqvgB2mC3YtQbRVDsPwKpCZX00ju67UjuzeIaV1HtBQ
kVw13XDBFrVFzDpbfaNHcRmANxiNNq39Em2mJ5Wmb4aBRKwRX9L+IXaRGqKXO6JDgxp+kRMbXvjW
b3i+8PXT2ySEZSWsqioI9xmPnIAG5LF4ka1MtZ4bqKlQ1ta7E/lhWjLX8h6ABAMSyXJghizW5K6v
E5iuFd/e+A2QqFzaGyUh+L02eKyv1AbdD5TEuFHA6dJ0y0VH73mmHkpquEVnmP/ejGvb54CXLIzF
OmMw1ILhFl7S6NDkYLX6l2ZcMS+/yAYOVrBkYfsAQJwmZCBD19szPOnBuDPpN/4eWrM3GpHXRJQf
Yn2SJctnIBQMejNnm6cwH8n6+GAyP6FfaH37usYjaHTFD3j4zAxx1NiuB0ckRQTzp1kdh3UVIWDF
HHCZb2pklxA9vvai4E0AmB0L4PuFRBzKgTh/+RMwaQq2ERZT0wccW6pJ+wNuckCd4ft5qG0NNu/d
1etxx7uza7QEPZEjmOLdg4iu3KTDifB2eDzJ0eWpXMdu/qH1b7GaD8X/asI5cHPoUdKSB0/w6Cee
UbTAkt2O2uUFXERNBZjZ6TjoLs0IszvbFponw2KO+KQK5MwBxytYo+ItCx3xR18yFn6JcSzbRkTz
tWzvNeR+R10Pf3cUOPGdL7lcxAJRGhZL16WH0kVGK1Tf1U8iajZeaj1qCqcKQLN5T2gGXZ5RYoek
rOA95VFllHUJFqsoXx0DsmeYmMfjJd12XI4v16Dk/qrvolQwODx2DKGZYyr/VaCrlB+kwXWZe83C
qYW2M4uKXvqBepi68L24mVbVmRwFun7lV1uih+NURpuyG7OTdFj5wL+URQOOT8Nruiv12tEaE4xV
Mc7Nel/dUlc3fZvHjKpwPptGX7h5+j5dC/dAc5SL7tPhcBX93xSuBVNV3L6Ko4xvxdACZuNjsZ8c
mhwY6YjliT8KmKiXPDdtUh6M629zXtjYSItmm5Dtje6T+vtVgHMgXPWmHWrVY1PDbEW9y1I0oOuH
b2csehhQefKgvd5MOxJIOjGLiKSiOAiE2TIIKGsqXdQ8ijTumiiKMwC2f0U2DIaIFbl2G4ZpFuFw
f4mIgHAnmUN+9e+qrSdN2qJA4FlPp8V+E7DsYm/evjouMQu3V1W0CINcVAWZ7oiZyk2xlFPgZQGt
txhoydZci7Gz6LKwKDfZHbV9PCpTfAqiw6m9mKitd35t1DsIQgWZ2tNTqsc6kSQrL9NAtztJ9koQ
ULcY82xDg6VTIvAkeLCtbwPOrAYryHy2IRYTvUoMWi6q0sSHkIQy+tJq9DoE90Pf8/Xv8m1lzVfK
u8uJQkoX/VmfO1TiWWg1BUTXE3znL6rfNQqLnNQEbmrr609khT655jPbd1gTR/ONZdswY8X8nhaw
9xjE3I8m59r248iJihtMn2rrt7u560k+p93fVaycA8vlG9r/rHhVSiXbJlZPsO6yDlYqVva5ehTY
gcETyeyH+aX2vvS1IctT6buZLJWVo/NwJhEs3WHfrT4ap02PfDcd28zbZR3eehn+ixcytTmje0qU
ZDRLSpSSyiyzmNMf860dL+maODJBYNn/vEZZOc+wkUFk8qK8pK41Fd1DtMpu4gQmhVg6M/wmiPiN
IQ9Xm8QghNQs7Jb1dWLOrXasqSN+BZfzxg2bN+0Ajbx2xCd6Leg0F3yINSJ5PClxHNzQROZJ0AYj
afAplnOJ+rrMfnRHt2fq04B3WcwgHnvYzupSyMBZsLI+1Q2NkDWMKe3SPS6Vw4hHGKy1Y/BLywSY
rLQgbXMxnairQPFoQgBmq+oaPeR1483dwDtXD627nljVIave5liUS9QPVIZLHo9Z6zPjtkciFOH8
PrS6ggRUyO2ej1roJeL62za7IfbuMCGVdVrYRkcxZVnBNLQDRc4yEb8LrYpWnv3cempYoB7XcM1G
g3CnHu6f/87V/nJgJKfJbapkLZmY9ss9hcRxK7plsp9QfJcvD/p1cVmsHgHHi7Ng0o/j1+lUY4ko
IL+rmEgzA0UUKj6ewBu5zu04B7f5eq0lXJL/dOQQDvPGK5kcBVQmR+ZzyWT+9rOLme0AmmC4OBaO
PKPM/6O/ApNzVHffyxJTOlinKPEbpqfBr8ZZdfhJ+k/WDaeo4qLg5GsRWOGjcbTSTJs6+zpGUMCq
w7QxarbsDs7NZrIHX9YYXpoZZ/aMKyDSFPt1tTrSMDOw0nMZpbsDFWKtRDwRHTEIK6MxGs1L2UKX
c1Oe1KKfon1OrwU6Cw8RcQK3ciTNdIz5Vvu0oCuarSvmButVutYWjBCP+pTV9jTc43dkDcDEE/GX
l2c9qmv9W59JC9IevHuQpkh7kYpPuBOaEstQOS83OXIux8UwomkTP+oMx1H3QQGNJ+GHGk8fF8BM
ueV3L6LSYzDTxbx+dHe50HkZuN0BLEW202Yamrb+jhQlEcCYbl0G1teAb05QU1cNYJvhwmWJ1gYO
0BtrNgPmHGW3twQc9JzwQ+9q2h1OVUtIC0TQqpksz6sgxuOOSFKVBbxytKWKwIEQUjzJOAOTYexK
rpL7PUgbRzqvGYeHg3XB2L2P6JSnllhsW4eqByJ0KPaAK5q0PXjW17HG25YLj/rJ8lrjdqFfwKie
EUIviqj0VdJs37Wh9K/pTzDzDjhYIiNM0uCCtNdULX6dqvDUWoHjsGgjL/QXImWSKxRyUwAA+jIZ
HCrCQikMdnC9wzEoEBce9Uf9jq9v318EtE5KKw9KUXzV9jn/cM3F+GS7uHEMaUO6BMKegah1CM4A
nEhjojNX2PTfaP+iIoatMBbr6lE60w7ImNq9+wK16lpU+N1w/+d3AYlstZiOrg+1LhKoaB80Y4qT
SyNIRGGWtgJot44+rU+B23poR6wJqg32jTJ7kqQwv5AJlRITuwP+KThQcFtBBI3TPM9TS1ktNhar
mYW73I9zl6ExOpLI0+ZSWJklOCD5+LSll22VzsObgLSlXvUzPhICf1YzG4qu0FOzbIIfxAFUXFUM
NRRjB3F8H9TQhtmNzAlhY2+9FNa7ol3gXTXOGpkCfbtJ6Cou91X2Z+vNlXwfXREU+eAeB8eExxKu
2PsF0Mq48Aw3GLFeUfeH2XKqR4OSrkVGn93h4jk386I9vjmIiBre4rhQurcvf+JD4hpak4hvS1gt
3aA8IbHdQe/rT/qhuvaqcbe5sS51u96ZXyvGgzZog598cYCu7xvwRVgf2dvUv0JnW3XHqvZblMHn
ILo7UnMxs/7Z1duywJJToyvhtYqZLUkImdAGD8VXgu6jpcsk7Uuv1Ey2CPdVvgMRWsM9j0NPjfHc
OqZgAO+dRLNfLYv0KbCPaT35stHkoFN7jZZgeoxwoKaWWhDDJc2TAwURHQFdPGEPOfZvyvDfPJ9S
9Cfuimzl8FhJiOBlk1RfyifEl+hsHwlheS1+aMvJTuH9LkOLMBSFbP+CyU84VLa0/QHM7LdU2egC
z8/pvPvmQ5ypPLBZiVn5wUr0m2VxHhf22kGn37Ke6jNgwnSzxM+RwG697qdJMu8JHW6QCgon6wrf
f0yCVP1y4kTbLj8qhv+cbw9XTIN49mP3+XYxu6eSsDEwGQCKbt1XyagKyzuG6/7GYnrgM86syOWi
TXeqYQb3ST9zZV4X+vNWIE+0Ot3yX34FzQ4jGmT9Lx5ijvTRcS2u7FwwnB3hNZWewcin288qJxIa
e4B4VsyVbAFTBpfriDKwI+wdlCj77UH4jnuiOUTbJFY1qM02OjfRKAAcRaWus00ENHShlTJRDmaL
08DIQzZ4IoUYRo7D3LA/dwfSWgrXdzn4ulcgXfKX/CVqn3Xkuy5eeDWf9tByKeGxoJd2wHCTN4ae
2eKh/e91o0dc8o4JLBs/W2f4qRFPeMIHTjtwvaF4pM3492bYqFhyf2FgkIwwYVRQTL8Im2k9qf51
CtxrjWccIRX9JwM4xd2KHNyJEKCoQIMWSZLfozFDXoU3dTQCPz6rEv9eU6Tjh33zJZzsYQKeDCDy
W9hRPBVbB5qIj5G/bbLPxgDZUwBwRTsk+Z8ISNaUSGYs6AATJ5CGnd+msWhO4csklD7XJtTBKDql
yZhvhpLL0CJUrzESnm/HnT0y8rtNP16jBX3HspxiugauXOfWDDDY9dEF+SVkV5Dcj+yEnWPNjiSn
EZIw8we11yAB/Uu4kJdIzIp6XkxLdJNB7oGFHDe3tbJJvViy0F0fAyjm2JBI2yGib1zSZ8LqElFO
FZ0TJezJ+N/o35SUG32Bvr3yW5FRLoPx+T33lWfG1FwjxYTo5rc7B+nc1IAzwU/RQeItbycQ2PvR
J+A21prYDnL/U5m/Gjdvpg5v1tESOmppPMcHnDv2a/HDD+ex3KuRm1Db8gRoEPPM1bvfX9UIH9tr
QYyn6gR3WK+2E9xwXAzQ8bF7ODqp6sNO9dmQiy3dbvOH2PV0oVhBzUgIsiQhEwXN7P5Bq5O9aScf
akle6qApH1cELWuQbhqVVGH+FxK4NLe4kk0EZRSBkGoKrrmF/mwRcT92uk4SrIQDxAadQw4SDgWK
H8MoZMOw0QnWRAWD+kH6xuBM1NLDbCgZhD79eLNHzUFU9+zNcH4LRsN+cimWex7Gy7sotpMyNTko
afYshLAOTaS6IunUbi14Z0Fc0Nao6a1uxn3A7NFSIKV/TimSLmTEWPg8KcYx3bGAKfaoKsAOkFUF
ozWDUG5Epg+MorxpdOuxeCiMFVJgKSdPNcx7sW91EwroI7XsNc44G1oHC9Uz4lDU1R1ZNs2bu5eh
iizrOxhZ9hvX4nEEE8ikVqGEy8I15JS7mEgQoCWJnt7N8cucaBLZH99NossrDijAhWSIpNiKGgLJ
mtkQaHrelaymYsh4ispA2uvmZu/OsSPtST/eYcil2J3qAHk5wKhVNMv0OOqKshByE/zyk10RRMJx
JbhJSe1/XADS0LHkj/wivTEBeE8ULBFvFph/c7cc4nH11Mg3POnmw/cv5PkG/vwkyXcxEy5pGHf8
M9q9g+9hl6AayhIkWpfHMBuOGVKzy4Dn1q7tGASHnYLppktQR3O7XOKjSvMQNF8TiHjOvHnbQ0JY
7zsY9PdpIblokYnv24immHtoz8U0fxH70z3Hqzw84FgLpHYqRYFQb3QMrMqFl3RKPsNOd9pLHG/d
3Zcf5ScJ3vMMxnDG+Y7weLaAi9ynRqt+98QWogfcG4eltiWBJ8hgcMWC1+xR+h81xQ6xHzB86xgC
hR2dQG+NNO0Nu1Kvp9RtHQAOncAh9h1f1gHNjOwJiNssd8jULu91ut511l4+zjMDE2p0FW1aSxEY
hcvInUC1wYQT7VfbAkiEsp2J+1ILyKYalDFgWlYivkw7iXxsJ9FtnT3Z/OjPcJQ8SHQ9d76yetJV
McejuqXFK34rU5FJhoBqsWIQZtuMVcwwRGU01jO2q7Di0MWMEWFPY15u1LMKZpVik8P4XJWca119
B0ut0XGuPtQib5q6vTTk9w2gbPQabgM+/Di0OMt+Wzu/NiSQZG4aEhCDCFYPcTjH+sdyky563ww+
dBYQobZ3wwxnbsDCo3K9YF1AicZNT1hKLck9s7EbVcSosdZnwaAgLWjylYYSXY6FU0m5k+GfGydc
tC9wY8CONBE9ffujdabTUlGiSvKpaFO1Q8+ggSRR4ygeW7OQMuO1Qkb0VCqNpYThFpRpHkB1nwrj
uHDli1QFtcAm4IL2FJd/jEiX3os5LwPWjqr+FMAKt9L+b9bIlgHU/JK58dFIk2XS5Yg5oTDsSl4s
IGxM1xT6h+ac/YRTHriuviZelNfQDj2xiV6JcRBtAlUdnYjtECMgQTCHZeLZ+/pVNJrlqrO5jKMx
oUCPblfPwM7518CbYyzc0qoNbfxYiSrexRfPQmISipBZ9ygWEBVBbODo15+sX+/bvyleOU9cXvJP
yK+9DUhtxkAdt+ikJuzxQJzS+beX5+fR71I4309FLGtqdFSYps8xtPehACYu8AxvzY2yNiaUKeGE
rkP5RIlvVgAdcHCWSlUnBIytJouagEDqtWRehW3TPvFSSdCH6r7TFBqbQwyT/InWjS+Nysvhy7xu
mecd5ywyviI/ymD5cDDxYYw8CRjFET8iNSXBEsBtpXq3PfnCW5esQ7XBNxyxSG4E4V54V7khdxrZ
YV3MVH7fpxSk4oDchn0WJCSf3dE232cwtl4GC7SBIdYBFchcN9JvXt0iNVKJB5vxx7+oyRHmLSPm
QHc0HblXb0Z+lJ4ZFxsqy6Zi+KgtPBxWx5TMUzi51MBjIQQMBGlPx/Z/UUckqfGM9rESwsOL2eN0
qHipoZ7jq5cBhTBBj/T9tts3Y5RO6eXBaxCrwVnwgVTwTJ+/1riK8jOB/XyzGgbsTcEE91AcZq78
uFWk5qhBk7EbcjNd5HOqXbPqZj6bJWWUjbHUqRmN9AGgOPdScjLw2CdM2xSoYMsnfUxpMFpknw1G
mHDIORzMJOn2o/1FOAUIThlbi2XPCBxMYm08jPGI7eVS/0MTzzOVQhCbr/c+g7PEMGzZRsPQhdic
1OishWFqxkvwefq3xSp5+B/8/2pX0Cy4MuXY5yM/q4wWobTcnted944TxV9OSuLtusIuRX0QAvY3
0YYrU0y5FxLySADOFLDfunbZ9U5yoqtUImR4kFnm2c/RDxm03Jod0WOGxnG1sTthUnZp9BTzBjCU
djczDpPlqPxVz5nENR6zNf7Ix6C4MJwxqPvyAaGDBSPgy/zvj4c3GnfmC5s/dkZpZL0EISpq5r7u
8GJgqmdPRO5w69TEw2XAnjlmdVAkaN09IeDX3l7FFaQf8Tonl/3dShZ/s4ALWFN5UK0npr1f/Cw4
1FaQUV4uIJ099BEwtKN0JS2fhwlt6SqNpa20wBAywfMYGGzuBa02MPRitSi6CmhJNet43HWfDdmy
ZXa3oJs1Bu9FxoE3pFdWPvot0/ayaGjU7JMrpF4o/RGsRXx5wZ7ykovHUGNtceJlYiHxzEYl1n+S
zccQDSxpPL+JHSR3i6kSKRDe88c6Oe3OZHjr7D/a8BRxwls+fg377t2xfWlGcVuKNIaxhobqo69r
AVImaAClRRhf3oplTwrgHWLXYlYRXiwP/+9oqgKIACKRBNAI/4q6Fo7Tq952ceZHa+9cauEziivC
WMZBZWwudCAuJXB9Q7oLiTQPYdWkDnrkfQDdbQbCioIMdw6uCxAnntplPaMtWRTXEb96PDKbQxC2
GXgO86UHQdUdv5gKLBf4IfoL7HfXZOhge0i9xDBQjR85HEv/+E9UhEhTEcn43QWfBehtnfoGVT89
hw6zTV59+a55jKsKEAT4r2nsn3+ZtDFmSRP5l/xEzao465vzYSsB541Cobz7e2FNP6l1Dwx1u7z/
u/LgFfHDnYPywwFd25Uj9BIcqzQP6UTOgpb8jE5lpyrI3BQi1ag6HQHnx+B2XY0b2QnqIQjah9qi
SkjeqcKUDWbhQCYnhzXNFTttqgUWMTDCH1hcfvWRdPmkpKmbyRq5pFfWtrOfEqDEf+WkmAN8ML9V
n0tFi+V4Huv+XeGn+ccSVLhI5qu3i5yFm5r1+IOrZTk8Mo7go3sS7cFSrjiKXsWhpFXdbXsz38I6
wPbeoTGmdDn19Mml6UhSOQzyM4GrrkV06cwJPyqJVmOSxGobRGMHw+XX/FOLTiG9hRJ97oO9l2tK
IZOWK7FFTP+LHMa775AalzqqbL6knmzK7R0YzSGY0W964V3PcPEl+LZWG0sqhxl6VHkCnahu1TsM
mfKD2YgmiPu801DDmBFiNd2yCbUfDFW9du/ucIvm9bIooHithk08zRpeTp2Ne9K1wQyME+s0nFDr
ZJu3XQQodv7CDr9PzBb1h9vywFtIINiFrPYWT/2MA+S9+Fg0maeHKQgadwkhPYL/Rrecl8C1eVHY
mqKZMzu+T/TrdeRFr0A2oVQklVYIBeRTm3kEBe/pX/Mj9fWaB1v2+NyV4Jn02VCCm98f7DZA1Eem
2n92rfJDEzt6xPXpYu8bIWzV6euNeNFc2moBdrQXJ6UfYXYpOp4JcfDU6VJEQQIkusKQ1FSjMcqg
S3PNTtJbB2swkxvmWUh9CKz7coS6ymAhkld20u0sghXaXioY8wfz6Lm1dRIP3YqFwMvPJnzqFhEO
dbSVFpNQxsISTZUkD/5lAwHHqoD+893Y3ZH9kKn0sjbkVwbEyX/pTVEqVhUBwdHyPDYLValIHn4J
z5r1gMNvFrgWMUbpt2wkqh0TjRaJCY87m/VDZ2KHcc52XmHpsioa75STwBxGq3gqa+myUwv/yX0p
YNis+4c+eN6mqrcNBfGb9MN/wIHvwaRcVf24IK8MTOPv9Vs3fKOm3/d98N2KXGK0wkyXlT7DGvgW
ufErpY8fpt77IRgbIjFr5RdQu7zmhJelPJQhR9ioCZUKbQDevN71U0B6P/4HPueFwxRG7WOZmODF
3YAY8wyxgNYm/abQcyBh/saf7W8pi4aV3djlIAuGlBgjaMIF1Heu1FJTKQxkrMPk0WvtzSZxSKd1
qiHOC7ekB86T5/mDH4Wk2xmMtAv00ons23KDTm27mRqunX7fvli1jLymrFgRI92ytRNkJZSBybtx
nREwo5JHnM8b3sQrDCVuqSsvqM7dAdhSKto5xt02zHNL5PXITycTFlz/yq31aBnXWRik24CXXJhU
Dsuh5+N7GZ+RhxPN5yl0w1+bxGBCFw4wbiEw4GMCDNLdn57hhBiThoapVifkp7tQOCVOaacccQQq
YUtRemO1ffluiJ3IBuVSHBjhTSULSaq22WXbkIdv2Rwd7XLLblPYAJjoJKlilyZE/N+5pPZPILkR
rpwNvaaXu3NHn1ThLOmufjGXc+538ZBGGJr25irGd6waTgc/Tqc6ZlzaaNBacE/kutuDlFYtNH1L
d2jMc+fMSB+4aMIVkuySwfpxksle17McC8BufkKLFCOUGrzTPqkwfYBUTBpVPlWzP7J4fWp3GAKv
dVMTivVRWEzuqPuHzf49Oq2ruZSY9nJ3gYVlrUmaUg7I3T5vyg8E5eiZCP5XaMnlDPNjye36CeHI
FQ4EK7rtdvFFLQWS+AoBgVEIRhPthUGNVgKeLaUNiaOBwTtSEeSiqsTtUracgLxW6enUuOxwsK5r
SBB6ivRWKUXSj62wFWdvJwmI2SGjMFPYqxz7br5gp7oI0WIUTuodpyvwtDEfeBOxXoj8sExrD8cA
5/XXXhka2d5XaR08NCU/U/2IYqhDrmAJgSgmHZRH1Bra0V7QxRK1Q0k8cASMZFoC59ti6JMY4Ybg
G/5mFnngJUZ6QuqnGdxRXJaI6jsJ2XA+zlp64uR+bvzgLafhPRCGFkxIoEBOgiGWTadLYhYunoYw
4uTXExrwpj2T/lFjBUEdymzK8H3jTiArN/P3/8XwkK/FL5ALrf0rqosxaaAWZcE0kwYzIGsac5Wa
mn9iDDjEBiRKDTWgxIiZFiX+0emN/83IxB9/rs58zu5dzu+hBaaQbvDO8emfy7HF+nSnQSsN3JS2
lm7RzlyYchz1fHwSydBEvly8Pi9EjAR0OA3djDWQfXsTxb+qQcTuQnoca/3dTjPRQrB+mxHzNXCq
mZRM92RmpKBgCrAHJUkFfTYQKvT4dhxsAJ1s6MmIVLgtLeOugElA/+RbOfZZ9WHw0S0TpS+en4d0
03urvG/gYH7UeitKtHTl9aejuW0ffbhlcvI1YwDuaNtzDZ835w+03kZSvJqrTBEQg7g/VCk9HGMq
XAFcI0392b8fvYe0O+yiaTyVRW9DWxWzigS4yi3/p2ZsuVts5I5YzZsmwSsSKJNPAYZywFMTsoir
binhHJ+OVNWCTi/qx72diSFG62IBj1DaIYzdngbCdV5TB/gZ3p8rdYa5+Dr6zmCbJk00c8W4KFC5
rFKrnqOH3fYXFVzNnwTA7Lisf3ObaWvnTpXBUpIGoiH+lCE1eBdnP/3abyIh104LWPed5gP75Von
9FA5fjHp37eBT2jQ2+SR95uwx3z/lj7BiGhVV0Fj8YTMkNgWEICzEDbI3bPEHdzhM6FQ0VOlRi5z
8PH6VeQdYgK9AZLWurnsu6j8qOlqVesuS+PjJwVb/cYNV4WHlnrkUir1xcVEtKsqKSaDjI6br8NJ
wZ1f1s2rJtGEb9GZ0+Qhes1+eMENIlXFLHuvJTC5yDdcPhB71JGYdSg9QLCjFZiMz/EiOjb4Wa/c
+5NoYfHRM7DZqsU9Iul3cs1o1o4Zt3LyiiLEqWoQK+xb9Pr/yjGv4H3gsX/o65z6pLxuoaLAEVyt
/nZUSD4PF9p6k2pv1mSPgwil0Ttrxy95RKjTl6TZuqkvmwGZFnk+B58WfMNRrm8IF80bbVPlnd3e
Ez/w6++MboY/AB8SPwLGqEbHMergVY2qeHMETtllWMTFtDjYrod3858cPNmjO6RlKmHSN1TTf7u1
RF1JTOhlxwaXgIoT24+uW/pvl2LICc/1uNS2jD2qqJnu6s1r3hAXb+K7Xd2vGidkxbL1nUWZ1g/k
4QX5JOmBzu8bj2TQxHqXXIUaIOlux01aHSvgvSt9B9SNso2IgSuZKT3843sy9VlM05r5Ba9E5nZk
qEUlFsImG3xjogijWrbpuj2j5GEVK4rmPNZsmtRe4y458O8YbfSAF1sTAkU2sMnQlgYTryBi0dSs
7L0SyaUhqL/iFPCKQd28E4iT4GsJX0wsYoHFMLUI/G3NQ8DG4nI6XxPxTl7C9+KFCz8Mhj+qCx1a
ZwordK2qiDRCwsNG55gBOaGuK4mLzUnec7x5rS4OT4hj85i9Btytbr3DhUcw3NloRZ1pu89+kQxv
CABBSulj5uYenywUChJFj6NWLl6ikFlx4yspK3Ve+cl7jfIfS4lIEuC7i5fnPBjh9JvB0GscminD
aj++8gCVs9FGM2HcW+U+3Bn29s+SWM+RS0pGQyMWXZn+QkmlnXc2vcwYQ/6xBy1HE98AKKv26SWH
uckvRnv0BzlcBDqtUIMpeC7jgeYCz+/k4fK73wdIpj5Jp94RNXwOehyr0b5nu4d2gEj3cbE0ifvg
T2vsW+EtcDPN7D/rGeTgPedVG9EK9eAF1nh+vcr5MqIFtu5muyD20ZTtNAeSMqbh+G/F/WNaFBgq
pBAWIXgvhVSJQyC7e2WGDpJd47RptH8T/Kd5tz4GNPDF5Q25/PW3wdXzeS+REUGh/OwvOeEVRZFA
8togzj1LXqXs3wwfOJGnMhcDJ+csb44GG7mNdZM2oIDtsbvxCH7M1iC6xEVq4aux75AJcM52u6OJ
37C002hbSZPVAqV1q6Yz/TCe7HKcemmNaTVOZNvfJySKmbcdjCyXSAPuTLjB2jIaIPOj8jqraLky
FGsY+ZltDr3cKcWoqEfsZvEuRGb58BPgN/fnsBySvSmk8r5MEKATsLyAO6A6soOoK6gSqBJmbaLk
7+7qMfp3fZ9SBGctrU7px833Us+7xp2yPzgwo4o5RYhUkfYx8Z4AUcM39wsE4N7JB2AMCNZ8lX+k
AswSTnVkWAttgvcqn6nEm/sb6/nfsFviSo8+WQMdOQFKlELTCyxzw3/AU7L0V7gRC6ghYHBMXX9J
vR6GJCdyjY6eew30DYUEEjrjr32mcCsZz00rD2AsoCcK6hIbMNe+BekolehLfeOdABwflCUK30E8
dyfde2fFfZ84i5kJ3zpH6AKlQSijLBDuDT5pt6u/J1zWkZ15nJl2t6rklLKmXcRAzpexS5No9bmL
wUf6QcPD4hoJ1TQZpPISRWI17QZge8b6fsCxoaGWRRu/aE/iwmbW+hDWuaxILWRCEI53Shh6aza0
fHu040ICeH1JkHLUoIrv/rvhhsdnlBVhSLiyCMR8l9RJRxDauqHhOR5yaKqXrzRi/V6HeaV9DB0c
dd1vQsX4EFHdr6qIUzGSDjE4pP5jHmpmQ/P8sEAy20lbJ/d3t03X6ryLFrBV4g9Ky1qbizQi4Nyw
VAkChV3MIBmXkDgsW8SSsqCA5pIGJKCTtvwe+Zl6dl5gmQOuu0y5u+SXRtfawzjde50RTNSa6vVV
FedYIN1rFfGHZoYyCHIb9rMPtmFzEunUrnTDx7bXKj1vBxCEiXf703GRbMXVwhjjLXSCWsM2l5vD
wZAkyCwidYo5VtD7eDsTOmn5M1E7gBqDr+aduktmLQL0tMRFU9LMjcWAVLe8F4TNfzZPnNjTt4Kz
2KAxEMhJTOuyYIAurobJeN2I/MjV1zGsx/eCvbCkSz40zNBOIzhHZG/ilYJwSjAfZCsgd4Sd+8xQ
hwGpYAjQVh4nJy9pCDWuvE0l/Z9jJW+b7d71i5x2Znkgg6DTuLfSw7S24rGxTYDaHSPAJFFtRnaN
x41YNHn67R34/xtDF1n9RqILinIq+VqhggNY58EWbKq3ZaVs+CRvVGZv1ZGhDBd+hRBTrg5kCM0R
vZWpM/wKyF30RLHIcsnYr4NxbAuXt5++V22TxKFQBcD9tDsS77jOvUK0de90phDs/55g8dJygFx3
07N9ZAEUnN2FOt3ApFLKnK+JMKx3mA4DHD8/2RNW5SAnc9PH+Qvz83jxbyC9QeYmlFJBdOva5ucx
pnpzFvKHtzBdFML2iC92sHh6fl8y3mvIaKsnQePubdAY++Sr2K2Fw6mTP/imzMj85jzdTek74TAC
kzDd4OWaSm5P/83dxK2YazAjPGuPVY2heMdvbhHI0IowskeohBcGMk2EgPZeNytabVr/rNYEzete
4+HzKM3a5ldkR0UKYXRgpmf5kCmltsOmrZ1PJevNFBDhpcjNGOeoN+Ya+kProjvPpO7wkVqUTksl
jKgpkECcndJLxak4CkpmDIfYiMzm+cmNaVcMIVs30in1Om/2jwbcOyv2+E+E/XP7T7eID9jFNiHx
XfSrjXf0FIgkaImk/1fulABTXrsSF9M+bgvq5nbWxqbRRlOD8wfO+AEdzGWXD5galWki8GeFkVPs
UGu0IJKBKqrXqmvScbU1dHXtVjxCsnyZ4NqhD7pKl1NeYZBBQvB/N+XyqyEgrptQgQDSvK6rkVLE
MtvKA589LffOe4xR+l9LuFx0Pg2cVRl/c8IOZoNlYGED5dKuU6kd+6bcpbn3xkToPqNPGfQSgNfa
COK257HJRwgHCtA2KuZyNI7t7FigDkx4E6eT25hcajgsXehuYwJcowOM1LcKan4Z5xjledqGc8fD
wq4W4hu/aArI+pau1ZRJ5XGC/dE0uVHxy6se6AiAo79BOuioHbuCk7Z0ser+Ld+CCYs7lWDHrrh1
vN2z8pj+0r0iFIkEQV6QJbHQOEXNcanqaHwiKMjaJQdIJ8iiQhYaibQtKa710N5QUoJmMwDMLsJU
0d8AGGQLfr8PPzAgdJXwQ1S65nh22MJt4YDwBRxbEuvVvMhb3A+IJBFWTTX3Om0OaU21Ikf3eXBD
OMpl4lzBZlHREc5hqYoBJ5EBgCnGJGWzsWk/r2ePKLTim0gHGwc4Pmc2Rc9nuaRVYsBBfqGnag9w
+VX6w3O/Vx/rc3seqYAb5lX6i/uRXlWezWfQDDOHpyaNtDgetEnKkdMQ88Eh9J0x/0YC4M1DFW67
j9e1ylvVgi7UMa4ISV0XxNwSvQBHAS0zdlerAtdx1SHYEgsxOFcbaTbWWQqT9C7P7gSiZjMYPd6M
gJOEJZzXBPLdXQ5Wwl+Q4Wk4P5j7FXHfWYBijBtE1Ut99xsDkwxUj2iulPtvExdNT377/wZ9S2xz
izO7BGn4aINjjD8ZMWnoW7ryDJPj3vNgJVNndjBoGUMEJs5JgvrdCFvvgxsSBqNyU2nFfP5cc3WV
3PWNpBGLqlKI6lhoAQlpueD3ZbaFSpY3cgUI56vlMBMz+8NKuStnLN+fC/TJtGCl3Cz0iVSMSw3j
4qgPizE5EEdoBHgI9uPqeYwepCPlKLN7Ha1fwY8NtDRGX6cK3la51x7lt+vfYMYw3H3Gn2rFbrTN
EHy495l/PdVL3cczI7YGoc14l9wE2yYdnMXg3uz3vM1OU2FTgAqqmTjhO5WRP+ckw7UzQuLHtaHd
7U/KKOJrWdajSVCT9jmJGQr2grcLbUQ852nte/XqK6hYOxv/laTP3kfNPztR62ebFfVWaNb2qkob
znqs7bFyax87l2kcHRFVrM+6lCL9P5PH0WnQUDJLr6corRwPVOuMobBrLMstyVhBhqsSJNBjsAad
WF2wWRFpZn3lKBPq6JmjO0kPrSFgjcCIhBOXHqzq198UqRWpXJt1tyJLrbZ40/WbiBGcQsNsZwJv
WzN4yA2FH99HOkb+DAN/FQkeK7LpI4sefH7WXnfcKHLo8fW/ct6ikkFje3Yf3QCG6kMSL2DhCtAE
667RPi4Aw2xTAPAwm6+RnI7Mku1AQCxCaLZfZu6lqQwP6zPvg2wqT89KKuQ+v7WTbmLeUmvKXMFg
yJiSlvOK90bePYxs8aZ0OVFrVYXy72/mWetPG3q34m3d2z2nfpJV4xcGnWtJ3+uGB4fL2U1apQDn
el9oNJyf4aqmHomghHkRf5NMLGsKcfJ33drLOVLez43FgLDVr/Rqcb5vKWS7CJM36jjOXQu6qMwD
8rczz8DcPunD8VT7g5bf5d12axrYtGoeAqWzMT/bsfx63DBEMpVxpBx0le21QkqRvyqNnpFug4Af
0tctDAQUNsu85qpNg/YLcUzD1WuQ8aGjSU5McxHfwaPxnNWo/Yt5lB+chgfXf91K04L/Ow6vblpK
yK3YGn4MPjKAWtq0/pxhF7VAPsGZoq1CMlvtmRuiJDk6OJWQSbMoSYrZ1vmTnZWrALObBLgHIu67
3w0ohwJ9LYfR3gT0KQUe2PYAkMwm54d/yP10GiajoRRB+0ApVnAmaEH9/CL0lXZDK8FQST/6D/O3
ltjjU4UN7rHz3REJ9aKbyNpW9TuDNo8Uy+vuNTSdVcr5+XDLyV4ur2wy1uBgdREmIncQiAz10XyR
m98A6Aq7IY0oaZbOBusB8hXzR7f+b3YM0JWxNv2WZtCDQQR21DI+xlZp6vanJT/QuPJcDZrhRznH
3cM9ueK1P9Iath+1x14X/KYztELoUjgOuBILabapXQamtouxJz5XH2DoSMxWz2pzNAqJ3jfTlYCq
RZMI5dyMLm4Zyc0DiQLnAXxIgG7ZHSCQlgzdEaYeUd/dMR4o67F+h5vYPFTIt8E5W0sPEB13KGVK
AyuaT8ejFQwy89qS1SP+5E2XZbtAabfgRCI2YvfV54BmnLKhEiG8P6eq3p1nh/eSXmkAgd/Z/aSU
JmDk7gfcyYmz5qFY9j8qTvBcnxfFDktvH9Ng5NGQRwgNkK/HwYHNAmWOOzpWxphfYY3vCyVJ3GoG
OXxG6OgPDSqFLSNO2v/PZx5HQ3qn07/12y/Af5UMOoD9SSfEogJl4Gdjj+w3QwCaLDCA1RLR2a1x
17uB+1yWKLqUWNGOPfzzrty9TBmg6v3ih1d1RdLq9mNF3JbNm94x9wousHbEcHj/iJsLNWp5bST1
4uoQ1EywrflO8SyacxUwPhU6Y4CZphgmaV5qIbo8OekYNMRW2ZeUkZJlcjA6rLab+qNRiUTlHqCJ
jv0k5X+l2ZE2USNU5KKUDgHQd7wYFzWSM+L4Td/6uXP/AxVEG6hK5kl6K4meADnESphi13f153f2
4NtK+Xq6FhWMPLwb2I4cO88T6cOBAZ26w2KvcyujXLQXIxzXkwM/uj3GlaNn0CkT03atxawNQaOx
PwSY5Slq2ikaRdhGj7JdqiOEywk0aXNPlLkxww4d0EbsV8BfUS4kzjAKjUM7+cS1+FWtV6ih7PXh
9nMtugXJQImrCjmfDAPNrVRT628Zo9FYBUfrIpFXI6+dV2RCUAN7rvLH2lhPxseaOd8k3fCMf5tz
0wZj3v2Q1UCsAp/gp8un/IIg3EtQ0oO2khepa6VfHkIxmw0n2lalhsz1Qj9c0BgE/Rk6+TnpJtmx
20F7VflvoWyqimG70LVId2zPdySIBOyRhUaTFrDIPkCULD3mh3EDXzDCM9RvLPT63OKmj3762Mrn
o8hCVgeDVvFlsnPYJPFLVgZ2ZSeqXn0Jk5vomOryKZToRuN9iD/cC9cQ00hksa9e4ua+T+BxpChR
ID7nIjRUK5hXNL5fQnac0Ott0a6zg3Da7w5Bjj2vGAqPFYGGxgJgTsGQt7yfU9InDFpfKhJ23zAe
rvJZn2Wbn1j2pjVVU0cA3A/iBGQf4qvpee3Eky+W9nhY9NLbzmOP9Xao0izurMGLbYq6xEx2w77I
3Aja9iBBO/ynuG6wIrjBOIaE1eZPaHE5kIE8vZ5qpsDuUgzXuOkHQQXn7rrCJF4ddPJhfpAn8cwr
OnLx264p+zzCXjBfPOGzMLd3hinBF3kYNmR0ZHqOO9sy+kFcPxzkywnAMmFtvKAQGKgYke1gq9o7
su8edHeUt8mpSxGpm/9JPkL4/c+m1rHBXaHVYmxi1O55cwSACEdZJ0D5oroh0/GLG9ijd5dhlb79
WTa0/jN91Pd+x2WhzzJcqvEgz/K9h4nwuZFISuCJbfiBbvAqrFuJt61wLQ9NSs2SDFc7TDY2Or3R
fQADZH9TzOD78tIjXwrzgQ56nw32+I8hVzYuqVuKug+AcQaufn2+fpNUEGmkA1tKaHXWjiKgptKY
klf+SftFZhGNcR5oCssDHxqN24lzgesUrbzX7+7Zk2aTtdSlouJIXCsXSnpUnt0qon6aokplZSM+
JNEF1jCVxElEwHTj4Rx2NZuYQQeq4Ar6qbnDi+BOvSe/CxFr7SbzlentKkkwFwf2x4yPSz84sfg7
hr4yP4VsPOcCgbbj/JaZ3PvM+y5g9/ePr4qCEIrunPVWf7YzTjG7L7FhT0RHUSfJO2MBvZe3iVGv
CDfo7RjbPLplaEv7Q1a7+PvlTKtNdZMSi+TFKHesk++6P7SIgXUq8VyGW1WHqzAWcQco9NCnIQ7l
2tCy9I5zQmg8hwrmD3+HmaF5N71GoMeoVxEJ17TIveKMQzNzp+zuBjoTYYM0V1QOnPGY7yu5e19A
GRsvSN6JtTwPtc3gOhA+S/IVoW/pbVWQ/p2WU1h2iFRVOR2B+nkvKYvZ27YNHWWAetUaR+O1tpBn
n1YTyZ8Wvb2qDj16pg2m6DaTc0j1yibZpRuQIeqj2v6ONMouMB4GuncSZe3WaxAFXkUW0jXBpik7
i+gxhA7cN7DFCvsUQLmomMgYZJG4yrMSygGdH9X2Mia/rkDH5ZSy2UzRXaKeoRwmqDS3WMbXgHUA
/NW/Dyonwu5WKwwEB97OkgBMfbCUI3K/mSM7tC2tSqfqhmxBQGrfdg1n4EdQM1ZAhW1zH7n9GImQ
wArbvfzmpeMVFhuREgiAiYxxxxsj+PVoCaNPQ+g60Zmo3RGDjst7bGw7xGGQLcLaEW1ajUXhffLY
TuNJqZFroB0qdZWR8ggd5KrS/SbPmGZZsq8WUf0RoK4AkY1Z7/a1E2Iby4MsySmBMVBx6TP1A9iJ
Kri1W9Im2b4yuKTeACEobtBJKjoRZVMNpaxEgvf/phR2hC5AXzDjKDQY5rnJgxiqD3/bhjdsijIq
+tJDe1VzClo5kjLAEfYhAMZz58gxteisUGZC4OL1Ce11hOh9aGlusOPVLdOCAdbxhg4EECHRbHDx
2ExvQc5djXYacf/R65+iV2RvYVpYTvKcs8ejBp7g1WGgfE7A8CVtIpfUgc68BMnZgvsdtYJHRlSN
avE19Rw/vjn0x8ix73VqU551+k7EBCxrmBFtqnMaffsMiXbdHqFoHSv9ZrMfx1OzPemiBiIG6ddA
N/V3p7yQirgw+JzKWVe2h5OXc2ghk6X4koTkgxoea7yBaEBOwceg7F93nyEPyAAqFDNV4/qZ7uUb
HtUmtgh4RZbu9fnRivm/7qhG2GpfU6gLSavSqF3sKaWPSh7SR9hY99rNwrhkZmlwXX5VwrbNtOo0
L0ue6ds6dBC3fNKBS4AGdWypx269K3u7R+rh4MggBhAxhAaK5B3o7tNvpppSEsJyt1zql8qH+PNB
wMnHBGAUatK4/1ee7dxEG/54pfwzFoXi5jp7K5xgwVxybCuBrAbXkxFJGbzONP+6LrR6v4AgluYo
TQsLuzNd0wIMKx2XcyNLaYMt+rdbqhmYbnRlhC8X9rSZXzsjUxduZ3gTLZUA9JOfYUZw1wRIP57P
GUKwqc7wDSD7Qp/KWti6N5WtBFn8OgDErt+Dj88RcTCVtbpwsWHMOTLa0YsuymAKgZWtEGUazC9a
+Ou/QrVTEbv8Akrcbdi741vhDw0dHtYY1Qp2O/Yf6mshWv8hv1rtUbMUsBtK7s0Jxsuk5jcOFKWx
v4pVbcKTJUuQZDFSXofuPQmC+yYppjkLmKBFJlUzWVOG658//8lzcj9ucvIkJAbMBcW0EgqxAKZY
BajBRPu+yKbh9D91a87QpMmFUaaO4Tfhn6H9fZdGhrHkc02BUPree2KsiA4JVPKXW3KOvH6GUPyK
blsDyoegdSQKnPwxQdaxOMyOUZwd/O1LnCyFhJKFCgQ+aoXDAlRdT5xCd1LM4c5bKJuCZ7cEwVT/
IZBk5Kijwt4cpDD5phvkt7TnBOSPy8BKxY3xmimPWfvbMDN9jimzACQaZ7rk8lrODcme49a1Op/c
pC5BtJ+WTPU4UTKceqK8gal7GCZCb4RVoqq5W4ABzugYpAExQ/LSegeU7svdc1iV6eZu8MLm4CU3
n5N04reajo61kYkng/ERfVAITP3O4W0GoE8FE8ocbQgMterDjI5pyl5iwZbH8hyH1Gy6cBd4EUC+
BdEv90kxF+4sgzFoE+JIQ1pHkXWWZIZwxyn2Ob79eDlfaJtAlhd991bIN8QJugHMKL8GhTRnoax3
WnnfG2QHaiC4Cl8QzCbxWQY713YMXURyz1G5VcsQnkrtUYjbMkZQesvdEIA6XxUIz+YMJ3z/X49T
MjxzzMFYF3aukBDm+stzODVFvSaGaK9RMS9VRep2w9zZFitWuC9FaryXNvgoGaJUzHNOOOga291F
gE7i4MnxLME2L+Yu7EJqNvEEqkKZZrqJmU0D+gxnwkFDCQw3ti1Emy6HDx030VXZttxM9h9ILMRj
NcA9hng4AIs+dG4qH2QLLcLAvRtBPu4C9ASj5QgiUXBQLAEPwba0oM5+kzMkeRBkYa7lrNQuZ0+0
askVfemk9uly80VB+LUbBSHJf77YMNqQ2hz22UcR3mHn9LvHmOomkhc58czaYP4/gNUgBvAnLiRt
EAoQE2Uj6YWb7y+mpbwCvUfzdWnWpBHCknJFDH0CInM0SJKpKSf1DUm+OliN99r/IL9aelaplaa6
YGaWDTMtOkhHrnFrvaATkdUM9JRzAgwv1KRHuoWIfiz6tNmhH0I1B3VXKqufBmK7fzZNkVTiGmOU
LxgcSbVX25Tr9cQwJtwHfif10q3647gqfYXzZCRkWaNbDuh6+B+rQU2s+3EdjLw4Jt4l2kO5gTLj
EQOZ4hFyDNag3wn+bwkTYihYWio3UgcX61zbfM3RPJbgWkuW9xksZF4X+wotReIzF1/L8KJy43OA
Uess3waFqf+pCLwWJWz6fC+9k/sIDyygjM+xsIeKddsUxbeMYLXKvt+qXp1ZajhWq/WElv3dBTAx
15LNqtqOkTXD+CfiYXYNfrtYzSJ2yR+VPbOWI7rGHNzD/3bHFuSPAITQGhVRhAMr8jr9BmR13eBr
+e6Xd36FTBYIUfHiS4PR15LInJMmmfXX8ugJOeFSz1AJfTgoH3ItMgVHsLkiTJcb5Zg0M+KAab04
4LZWlySydDNukRT9yLa806bxrJsjSSAVXcZR3pOVQGNvpc4/Atfh3xfC4QjRVB+hCr2Oybd/Oo6V
yiOMzDD77ZqdP0DFYR9fdzmizxVJrMfW4G/Z9RtT8d0DOyIlQhHmAUpfaRAGlePoXSPpZcjDSMFn
8V1ezmcjwudsHWEc0Q6Q2IfLk2saU7iDJh/SJU96w0IiLhE8+8G6JS+S6TObH1IZfpVOZ5xH1mxL
7mPgkSrzg2fnnolVbj2Se98UVxpRQwYNmTin9QsVlKjXf7V7hZMkd6kfc00X5yoVVtSq08eTw4hI
CbP1wW1HqIeSo+9OhiqB7rQepKrxu4cD4q7qQMt4gzbwK/Iyv3grcJfjzbF5dLclS9TCfpKG+KdD
7XFNOhGXZ4wOAOCRK2Gc6F+KRiIxP+bz8FBXbiu/x35IRfuhYYpoLPFBb3V9QOetsr8K1qpy8+Nn
EDvWGxTjLz4Hc7FcpdPpVhJOOHTqxf41bOFR9TlQqZaextykrVCT4aP/5/VwH9xdA82dxutRmxuO
kk+ffVb4QCba/XWZvRUV1jPQv3X7/Rv4BfsTa7/5fk/azsTNgKYv3kHR6IaIlcItB69axJ4Igsah
ZpnMtgljVtqZfWv4hHAPH7TYtEfIvJzkRgrmrBp1rxD8WHbFLEzNUjjwEEixaKZipYZOhNh9CuYR
24jU0s6z00O07SZGJWU8jveIv2e36jCEwwH4wgb0HxttNrtB8FCQ7dPHX9iFRonbQL69apgUWUFI
xv9u01x98rMPscj+6r5/RtLtpJm8ifBz/zj7iWvkI6U3xWsfBdvjbxmM5dSazGrk0TMWp7nqiCwX
u8qqZlWwcqvsCo6J8hCPOZ5NW3+bFpKwH3gXnwgNKDlQvwU6/heYyGECpB8jHHr5H9UoievzMbz9
5krvEvb8/gb4tGfs6wNE1Uc6jvcluKmu3YPyz3PMmPexTycqxhXCVK3pzLrQuSIDy8gr5d/276FI
2waj90hPScEcQIybDj9Yycd2ytbfkJAtf0fZ67Qts7bvVBMNYvnmS422OcYsUoIrRubAaugGzfbr
TRpSRwZ9rT1AxG3gEWAO9CImxgdV+/Ds6wxEfDPnlXLaqvubXkr6apviGUA/Fbw1k0I0p5dATMdu
/WEqZxU0Z9jM0uI0KJ6LB5gu+H0WqMLTAjNqB5mBEiOLslKKuETtdy294PD52SNtvJpTgtddYJ2r
QHl0EW+/YGVpy4mj2R4FJFopXZIzMBxEkK9SmN132KbwPIFwoZ3o+OilSZqr1zhHkNHtNs9SJS7o
JVPdnj1L3UevTUc+KhZuOgr9A5EXBZImhHOb3OErEmtkE5+AH9ebnbmzDqWfMjNRoLYwWfVW6TLS
0PGIaOMyLZ6v1x40Q/o29sh4ql1p/UZz7QnpT4OR8Zj/4gUKhJ95MxlnDzFvOgqkAEAnoCX49RDV
W0RdlnkG17u90TUclJ4eha+N424IErtBKvh0bjeE++w9RL0qBaFI0ogu86ko8PPz/0o3Ew9eUDQF
EHgrW8btFtEQhnZ7jJicORF2WgcW9MyryWJkRCZlpmf6ItcPiTDP51tNDz9JROBY3ZNzmWFds0Y6
b8I4cy62KJ5y9DHJarsh/cdHbR1/jnBvFF6gnQgvJkqkqGcKWB7pxkJr5+mpnkISUMvh5/72VsVU
GTCJC9mcqvjpTpVQy7te95DPXIdVJtMIjUuQiIJhbJYntxSZNxd/Acz5z9GamEDGcQNVb3I0jsmQ
mUGrT36xYCYcXM9RbwN97JSU5XPg0PV0tEMOQlnWvwnGvEoDjKLvDXS/cO2VJWSBj1wVK3pvUYCi
2sOAULefKSpJuq5S6kk478yZYGMghLk0il9OdFjlGv9xLlDYUWjpTm7yN4xGcIs1c1gVCfMx8dgZ
SGqAwDzRG7v7lBv3esxnZ6l4J4J3D5VCYJG9B1GF8GyFbf49r2Tu8KsRADdhUYI2AnxzRWDLyFRW
ppxyUVViBYuX1UGsINF0R40AQyV343B4rKYm+Kuevp2GlRUIKvOQnxhIZzndWTrMB9oRKr0K88hj
Z/K6T9EgbWepBxPzQZflKh0f0sB06wyA/LDuXlzMErGPuY6yRIc1Fb0ZR0HCjiBo5HegCj+t0+SP
Wy6vJK0mSTSvtLo5nSeSI6cMKscmriuggqX2Qado4w5otm4VJ0bCGe936/VzXQUttnF+CSzeKrPX
y8P5VKkiEryDXlkSwlMtkrnzDdYD3clQ9Dpig/NtQVZZkpkUT3cek2TJWf+HgpJg8vV1TSaa1YS8
co29Ifa/KYqjdev357GujydOThDbadfslFcWfOLq4ymlmZNr58Dcubim8tSJkFFirsGIVB7mtfS7
4Vq+zEauXU+ZbPfmQTxX3tzu8A2sr2eL5TI9pM0IAm1zisUrGN6ng1/kQqlt1E2bcJuOTiRr9DXN
8Q8CYX/0S1m3xTl6IF6l7xmQ8KqoMoBA9wtom7tvDUPnmPk7xgJskB/jE5FFVUrJd5MbR/4KEBk0
YSY67F67dOdxjRai5Sg0l42Hc4jhYp8425kFhCTj4vQHciXTfLDW2MoiVQFHwKNwMVuGPO6JSH/e
Ha77nnOAWCXvt7LMqVO9cQDFbIRUkRn2Z2w5EIEQVD8ZILfD33IlyquhPIrjoEvPHPI5SUpjP05y
KuhzlOM1F4XX/gTHkFwADSc2guNmF9J1pva/M4joDN0qjo8afKGtNF0s6Q237znzA2coVWRlM4MX
kj7mBc5nF1dl8oCDmMRy+GieaTtodWwanQKwszrxEpbTkyuBEa/WpKJSEohmysDmhBuSEA96D/zm
4EGUuUER/5fLzk14TvzpIVbR+5x6AeZ54ryYB7/L9ParRjz5v45o1pSwCa14A3JX8zaWhbIUmFYx
10VfU0otFccyHwxqkPjIr3RFOpZE01knKzMGOq7a9r6nlYqL7Z/dhhGDsycPpmCBtpK4v7D5/B4F
+Um2CIK2cBNxsxSLP7Xf6F2tRza8iY+ius0R8ykKobJXB+PzJl/kk9hM6JCXMX16o1s34zfM5hyb
Jv22PsG5EqOqNHAjuoPQ/TLnMGuLzhnhOpbz2hEh7iRPOLssSog+/7iK0B2jYKvCiCIRhZIlSm3d
WrR8D6HkSIgRJq1tDNefv8PM8YThJsZOMOv6QjGHiv5/+fYL5xcgiZgTJyUlV1niotwqvTQNj7tm
n9hSpNPspZM/BKXT6d4XIZWU9Y4XrPen/kv86MHJ8EwO38PTWcTd/06ID8D9Kg92dbS1ORHW7Wiv
deJeSAZR0ye//TF05KB/77COQPxmK9frj0W5O7uFUdbgvnlHjtT5D/hr5h/uyI4Eci4N/dR/9YYK
PNaKhbrQrv5H/xwOBMBhN7c59JiVoLZIf55cFIWCEckbRoh2cd8HBrkhJ8P5M3LShAUAdg1YehcB
TsPry6SU7ADm1o4VBqj4cnvIr4GtHOM2ZRHZFNNHkeDWo6+nUyQyqEJHex6sjZGtxWxwMptv/hnm
584rDgeRcmM5yn5yc8+H7RDDQ7clMLqCLQ1bgVNhSiueo/L8MUCOCisb+SdnYwdbUEoWA5vDdicv
SvP4ty03tMTFioW/iIyB+WMqL4oxH2s8vk9vt9DyH2Y68ld9VKoZFcl7SlR6ZAlXNkZZStytT4qY
wzxqZCHbmhre0vWCxPMTRkEZXHVSRzYIpgqkgQ/sYGWs0dFdz9n94zKYCn4J+TDDFpBj3QR8lq2T
0tOMXaTdgIgJQOgIR7TDsZM9J2Dh7kuC+wWvNsrw0Y49Sv37gXwXxR0LaAQfODOie29xiQina6RX
O49W5mxdQ1Zus+me6WXzpHnZ49/luGiH3cEC3a8gtxWZnWPD6nhE0fEWVsUonBZdj29laQvtzQmK
zK5Nf6F24sJ14rA4q6e5oFDRXlUELMCUbhqetaJ1QPS+DaDoPublITBt7m2gR38BnolZh1lvMfTe
jkDNO009t39FpF5O06CK84erHp6QqsXhMemmmzG5dS38lbR4H4AoDlPSvPpgj+U0HATSHtx3TezG
82GZbYcb1/iTZq7fcQg2V6Phs582lvuQaNLI8f9O/zIXA22f4YDens03v9plOcoBPU9PNlHeqmKq
iwRdj68QEmcxIV7cCru7qIktvqqxQ3fqtrAwXqm22hJmlYTA1vuo6sEW9/F0BjXDgZjsW42tfN5h
eDoIUbzgIHgJahyuuidzc2k6d8R4MwhL6hXeNCNnD/Ip2Z+Yq8ZZ2zA4uPvg08z0CDxLjvTsPLVP
wEHzTk9vqVXGiWUC7Eb+1eByMnrXsuxZsRtd1Lp0HIX0EzQmhTozSGvs1JXUnCeDMEfbkwnC9xVY
mrE5aZuhvzcIFrTfcmjcLMrb2MxY2Tea1JbTNedvAtoMZu6i+Up4ihCXCiLKwsMHHdQa9WdNBkaR
et1zW+miPfWUG+wFhn/EGh35mWOqyF7/xk/Hi65D70LMxQ0akNAo9vgxGyV+zYkRvTyWu+aWMSC8
98QwZvSm+Cr1WhDB8TCWlf3nEfJ1Ip5ihlR4ouH0ednWQVVw6bqPxZ2EO86/EPVUjYbUBYPC9b+X
jG8RO37nAyqtodLUWSfiFV+napm1h05x6/CwCEAUTHiNXp0QOswmK+G8Xa5xzAAhHUDwIF3ChCPd
Cw1byE7pWXrlYcBzvhu+krxSU+X/eG1k9okGuE+oBe3q48kbbtAjCUGyPEur3j89PgT1JZ2GBAnL
M0kg6kDcIMDlR4GyOiVIP4nhet1lElQzXSEy350zdIdd/dNuMPmCl6nUOaBGK4u51qhu8tMYS7qb
yfQhF3S3WoQ1e4JqAnLhn8YYDMnP8lxM2puRZMeRdjSXvVxo0o4bVAxpz8NGPVAaxfsj78DD7T1l
c4hfQkLitHKKeJWY71gpE7QAI5pVCiJeC3nPOmE7hw6cMb6mLMVYj2n1h88J0KkXjRTo1ROQYGw1
zwlfnVwystDBLvcFPJEaaVlj57PGdHzoCRvGX+VZw51Q3ei9OcyYSWisQA68ggtkdpCCzxUmIlm1
uPch4j7u2TxmCSuo5GkFMq7gvn7Xr6gGpI2qcYJjhfGJ06DyrFGcSSCFvAPewu0L4rePWkQdQvh/
dtdbwDYFM7ktmPC9TtsCraNAMnsF7uY7gbA9qs2unEU0Xloc0vb/ldc5G8Dd9FSpcBzWSxhuiNDD
UDDi7qQ3ZcLpzM//rad2794CrpqmCQAYp6zJWGdQFeOJh5P3QQRw5QSfvzhzfJw5On0Z2g0K2iON
zB2UWNzPAJpbigp0Am6X6E7kQEKL7H5Do5Xjfvh1rDUMoSUZaQkLXeYcZ/zVrI6ODLMIIH/QsBup
fz5xDM0DI4mZqtZOm1fN83MwaAuY7RxNm2Qc4wcucYRAT+eL0pJAltYgbqtgfNPicVvHNtiCUkID
9buUIdAOm6uKHQh1hwFEBcBchejUtJ0mbCVfd0OOfyi3EpAEcqctUMtj9qkC4NQT/PPQfir+KjaN
7hLPMpagcKkB70Y9FOcJW8jZ2WApX3CTS49BxHnjA3yc9XfS5+gDrslmih+Qy98QD6xMP3gWOsj9
ltAS1flR0bzPcVRgzWXILDHIneMRrz9mkdtKU5phwXkq/ZTYMLhez31RtMkagwDX6tiVHR52BAob
vKfsIJqi4+kv4ep9TUVGb6YeAVFhrKLQcHvTRFOtaMYgm3FiMPBDnBSGMk/ajKUC8jn5aFZGRagF
d+O/OoDdXnQhgzaxmKAasbAvINkeStQX+JjFg9Jlw9yhjnOXHFgFbQ28P5QvOucvEWQtNwk3ybBc
JIvohz8AqgOuKmHNajoWJGVzAr8FOGFlosIfT+m5wDFaZBvvAC0Qwzlmml8ydyQqgjoFARwkZWwV
8AkSiASh85ThlbL13wXmm800DMXP6hV+MUpc+02fT4one2mM2BaRLhV2rMj858HvSz1diA0YrOqy
4eZ2gouqvh2ogNqSFopNb3l2POxgEsuLJn3Kl//Fhcbu4gnAjkkD6kPn75I2Gp07WTUpljRkZMcO
uFJQqWQu0wBAz9BAbKwPCezSc416L1B4rgDOTZiA1uimKJsmikJ6uEa06Dem1aZTXqArLpmIO4HW
u7c2MRly3GMiRof016jajnSg4SYMk49KqXs4yUadsDb+tvsv3sVLhuHkcOzN6msIzOOH+H05QNvc
k09rVr8qy5kcKq47idnHFvLKZahtA8gBitsDvv1rSlAZqfrmHwNf/3PntwGw4sdivAZhf9sqjA3q
8XpXwxiMzNPeU4zXFxk6DtJk5JbKnYhCFFUlgP7pAFW99m6w6C5Ja0ukLYwkLJnRMPOw1Ne5aSDY
cBuf+jz/+xMhxIg8ljzS6RDRV33rToNAGDCjOGJURI0fRme7rGbSlvuxyfa1TJKmGSvonqNM7wrh
I8tz1vCCbRPaBTEx21PhD0AmsyRB8yZr9yqk5/uUWSJbsj2pRmIlCOLQtfw/ePF1V2qhhnf3gIia
eXhm9ysGSvHDtVePAW3NDlA8GNW2ofywt1HwnHp7d4yk93zEjj9dTglo7mrhgPVHgGaEu/wbINqI
ODmSB1zXvRHcrho9jSd+okgtQW34rndGjTy7GznRvp+qrTNGdPZ6JnG/RU9oZddI3FRvwWeFqXOu
OBy5Frog0zq1Drt1krAWSYSTfQMQluh7uwfEPSe4YQXZ0vJ1lzYRImrrkFxCxCYuiUxX/anyzHs9
wUhuLSosD0AjsbXQaoySJ8R1iZzyBs8KVozthNHXSxeUvlSs+7Xu3qSBurfdlwi2VD7jm4UE7QWG
RaO3DIe1+E6oyj+nhTs0wELJW+oBPid328cA8KiEiYqQC6z5YjdkZu7ssZI7yF8GpOTX3nyuZfnu
0nq7UeKwla7xpkZRk2/vBsYIZSNcQfdpH4rCK9JZEAN4NXJMziuWoUFR9X+tiC+QQrr+ic0NLFy8
4xuPOQ9iZRYE3dKhFwW2nzy7fD9hZpSnNPoAzBtLylcYoBW496VlvmX9DwMgpU7403UcKLGnDPSn
AJZJAdmFSxxQEQl7/umSu+qHNjG8/Ks47OC0TZSlZUMcS/+/Mlyf1aO1/pwDmy7A7gCxYdSNgmwx
garmgc2S33aNgDBeRHjQLCDEQSB8pfrcTQL2jP3x7h8x+lDdjwUqhPDxT2vskMC8NHIAuvmDC1RQ
2lDLqZQ+o+KfOciENSLvGrofWWFLvImKhD/xTNB+312e7C+Yt3nEFucEqEmgwMKstrQvBgmK27BT
cJQ+9itClYhbEXpCulEp0EYU1IXQV6+z5LK4bWwgl5sjNhEs2c9EWijLzc1kJONLOU9oYV1yroYa
5GBASn90sgZHwG8HFMMEtYCz+gcjr/o9vQziKw0iecrKJs+OuruwdgpMwbfN1YFYVo3MFcfcvlGb
shtrqtIwzagf2R05obGmvRQ0XriHCEwrQ45KRj1w/d42IZMuShuXV3NPJbTjqvB7cXkv4m2sXHp3
0MtfIo71DYn0UvUzrjFq9iFRrEWB+HNXPzaJkaUoKM64uUCZXnShRqAdpSgpy/T6/R2yxBcqARU6
atBSUzoRJJpxZDC1/7BebGaCTKx11hOH9vN4nYGLrU6wvcvVEh3yNa2A+zqVTtcLx4DDCBk4xnJT
WBUEMFAx8FIBHKQEaetpEe/s3OQZ6khxKF4kQ7SRClZfvwMYKxVsSoHSuXRYem7Y3LjT/ClJu6I6
TFSu6OUVWandt2PuvkZ5GmxZn+gTN0yLHGlb/SSHAes+rcC3hk+Gw0Vzb/9o3wb24AJ+ruemrRg2
AY5nDznE2TtedY3axDlIHCnOdlVVp6uWzpqiFTgypsPPcMbBC640wfdXqrh3v9An/A02qz0G8Zs+
Lq7IqesjlnyEquKb528w1iG7H226nBKDXQYj+pQddZEMsKrJA6857tdvd6GqMdqJX3Y3u/j7LZKG
I1r9I5hlIZTBDpmOyTJ6RtWcd6hyfpcm9Tc5Aff1E+rbCF5IDxQVp2zXtIBn24uQTYKpdi+CSJ1+
YsYurrr7JK7PgXIMHra50rAWI98vgCXXIIV4BvuYNGY97Q5CZF49vMlAYTTJRg6BrvvTVnMkOVk4
cfCYIOUJCXGpc9p7V3qsUPPdaWgaC8B4sAlJmCHeWxEOWYoEunHMqCXrQUDcXYK+t57aagDE8v5C
jOVG3A13mxtUkyHIic7vIM/8IAly2exVt+pJczAyNf4GFnkWL8LpV0XP5F7ik++Ix+PV0lShyuyQ
UaJ2PBQBpOoMAZrOvJQmAvGoooS4DWBh7iL4RtEMPrYgKLF6EWegsV40EwpNUECwfrIohYOYNMHg
1xOuQINEmeUqOWsXZIBTUCdH1l0Iok5cRycnbuTxSH8KpcagxxsbpZfVD4lgThS8MuShdK0Lshc7
VY9o8V5vbPtXm9kvN8eu1CFiUfLaf60blkdhkU5h/58RpBbkIyGz4ABtt3K+z0kqjafsn3dMvt33
6puuDzwJSAro6PAmSkIPYVPNUDqX4tUIwgptT6AQRiE5lpXftdqWgoGGdbhpxfwSHHKb/QPBu82m
raxN4EAqsk0VjzKaaJQSzYiL8rw6WW5txQUSKAmzLDldQP+STX0N5eaBIiZNOuAHxGwjijhOgwHR
6GbxCHCles2n7o9x1khSF3ezpS3NlDMQVu3f3ptHR1xG4O0yZ7c8pMquxKxoJCmbnUUPzoob+ukG
CJzOTCsyHWWL2DGd5wvSqZ7dwn/6xRLtB8wQVXUI6KN3ZDA8OI6UxagldC5mHKY0cRHM/HL3lxyE
yhEh/7YZUJe4AiTPkIw2JwjSDZ1IS+yzLI15gkV+seHOXKor0XDdTYJib2W3brfB8p16/A6SH5x3
2FQbsRfFKDKy57EOjGBkd5vi0QlDsLbJOkC9JFhZEXQn6Rtyg/lT/3JBR/jYhInUfzOpvSoTlGq9
7kHXIXwG09Gj2KzBbkTTxOYqGmy30+US0KFLL8Rg79Migudgj40AM7LZkvSAsncDKcDYTTXMpJWE
+MlVO9rv38Kkfdn8iBbou2So47Eqd17GekDHSIfJsHMWfd9dicmnAGaFfFviJDeVMzTjOx00wVgU
YJD+jhRyjKFU3bCk8csgAfgP7QrbkzB7fIpDg7inz3+Ivti0a+ApmeNTQ1AVpmCT6UvnMSgCeEAN
lN01qQqV8xbSsC0GjJ+9O24mglhLiRBs/a58awBUbQ86p8Nv5ojRTheA8FSJ7D0H364rw8RqmGt4
ouZoTA/koOVkDkTwIpa8/ruvOXaRA1E+nailsYZTZCujNnvFqjwHlj0qtRdtRVhnBoMvfatpivmj
AzYZ7tRunY10TzVxTN86TgnVMdWlHBXy7aPzyv8SS1t54t9naxe6ZAYIbmo55T/LtBnpz4Qc7Mxl
1wWlH9gJdlQq2qgoKuymaJIWT9LWxGvfYBuyxrnGa7525sxck0QTbkeDv5RTTcKMdUP86XlH9VgM
Yphts2D52RCqrT0q2uiTnBY3HS32/FMjKKkDw5kGsQjE1bMd2uHmQtd9hEF+NQdw1unb32tqOGXx
uOowy3nVFmdf9Xlx1XwGEZZuSQWRx2r0mt/CxOU3z14xjOXnUxxZI9J/sgMWWTZzrIsPJsnf/mKb
qHx5rhAl3BRO3KEOQ8hyLgFO8n7UB7KYHUYTId1ciq3ldoeF3vf0n/8ZvarVBcMgsX4NbcDyC/up
8OKgGS1p/vtMSeL/HpdhhHM/C5T8XQ3NQAGF+bTBAeeiEUKAo1d/eGH5NhMZ0mrK92nk+0Xp2hkg
S8uT1h3sEEX73MwBNET3kdzHkYWrAuDJEtLA7nVHj1760dxh0Tnkl34kuXysGAJf3G1Y0Y7Gegsh
tizW55HttvzCeTevkd/LB1tL7UAGmXpaX21/9bLO13ZT6XM2QXM++4XlR66VUD18FxApAEHH4Rhg
vhEHz1d5L31isgC66UXJBvpHVnriycYfHMYVN/eQHyXdIgqAgjimUAWV7raEa2FwRg7OSZebxIkv
yOv4Zc5n+PQ8PTltp+Rbp7FXmc0v4ZzDQ3PzYsMUXzQekMwrsZgDg9qViudv5Z0RFjbpjLIwJoGO
DqDmLYhQUfoBzxP9wmsJF4RiZ1irq2HtlFihAQQRwToEaSqKtxywYHjrYF670FCzdKJ9AJO8B40E
YLAvvHqfq+oXB9SPv7ueAJdsBsnoaneRpGk/OYXdhqBTcvb44uwFCsVNjxLRNqpMdd4eno0s4DW9
9zIJ84i+iQ3VBA6LsDOiQVZ0kRfSygC0XeFQ55eT4CVjpuiDgbM4jpKn6LswtPguQlsRk711Yagc
sdLp+8ShgtB5Gxa0m2iRsiwIbDj5+vIayaQumArP/arBrrTCy7zL+8whH2v4ofLp4x3RxPmC155p
+bwfA9O8QBYnodz51EMQln10wFAxW6mZY8ZYENLAW/x3pWm24ngSq6fTEHewxj2snxhsAAR3Eycf
cAQfDcZYyJW8CIU/Z2b7o0mWfjc2I/0CQeNFRKHvqCx5W6A5TidYDLfzOYFjOaGnFozmYbnSUZbz
ejBkPIBfT4q5TcRX8rQYWa7kfiCcYKRO1OAz0Gn8K7ZNhlIORzB02pjqbH+rEab19OaEEPEReCeu
wuwFuRNpn72QTHswItgjOhFgMBbGLt1YuMEcBGEgjNZjOEQcozsdSZR2nsElSOv5raN+x/DY6YZf
xs5DX3pfe7SnTAAC/MfH+OHF7sP1GfTglgDPltg8e04xR9CIOV9GBj9rWu2aQtwgx6N3NbJsgn9n
0eismRy12/buAD+Pv8J/nrDI822AatC9nPDtpjK2aZnuwb4W2ElM3CxcO9Gf13cKe8VjeAWxuiYv
ghUc+ZKLDDUPxtmHOYN7DIyhMK7hsVnqYOAIAjULxX8bidIcn42awAcGq8rc/b6V2LNwUCfU43Lk
Nz9GbnG9o4se1ABwJVGqMYkRkkmmkS/pO27qF2Y3viEZNPnvUli1mkucAkVgdzNeApff3eF8owsV
xKI+z3y2BU8u9AZXgsGSpUN2qGztcEOry+mkZEq+F8OPVjG0ENmzbsFm7VVLojGIT7LCp8MxV1qh
ro/lKDNeA4RB+mrBHeanhYmmCBcZ+pFso2iTEeFzPK12RkrLX1iCG3uA0jHAavl4NNqIkWRWF7yh
FkQvRzsfgsDA8PWDjV4YZPlXnT0fVfGPFY92XlaJwJSCoD8QhJHw+SojAIbksboNOwFPZ2+58qFI
3BrvsTADEvnhh7ZuKHFr/k8gL2asLb/XDtidgKViigcQE7+GddrJnsZSO+AEnJGEKcEdVY4OLBJ6
5PbuedVtEHbHV29AKxDb/5H/7g6m5n+H9R7+xAd+/JZqo8Dd8Muhbq+tIGboBQL1mnRH8fAko/IZ
7balwN84wlfuy0WN9unx+wk/ySI7ngdTiUFucy+4eTELiDcBkSM3r9o/OkE6+moNJB8X7w67xyZm
evsts4qPytVtXysg14VcqZTxXiq0qbbSEQtR3X7tSbVA3dbKHWrqqjTeODmlFk3WJxqAPDDHGNJP
HDa8Sn+AWL9VxyRDCQb21nTawz6Glkzhplt9yWot6Y1o71Jet5wF9friGbLlukK+qiJSwsUQaQWu
q+GKC2UKBbTq1aS4iTYbLWMXxOVqr+3V+6x+MeFKOjTc5swfeZ6xV4tjYggb2c/+dB9HYusBYpPX
sRbJSKSGTNUJiecTMx7lCEjqmO5NUIfMeLEQ6NjUJ/kKAsIk+yKG2YGt1CzC7zWriTOGp8C7LFP9
OZNYq6XV4Z81Zwhec3qcmmMEOBrRvc2wgQ4tXUrlRPzA/xUmDY6huxUE7mBWCj/rAWu60JIdIaKF
A9fWXDUWac1EeMiuVZQgrvlO4RSmC82kBPov04w7y6/YyHc1f+hDvEin9EJpgQExik+U/XyRVqjj
QA6VXc2BRMgKtIRhgxkBz1WMJhaWkSvpxPP78cqOJ7Cd6Qf6l/xmuPY+Yw0MGjw/F5E4TOqiU4BO
Ln0TT8CYZyupqR34VFxVwN/zz1zPye/VgbW++pyh1TRRTMn9UX4pSlQ1BGw2F+QIPsyzJCIsSHqJ
5vr9hJR5iAZjGm4WJ49/OGUqN6axrHQbPg2Cve/QsWKapChrdmxOh3aBiN4H55kqCoHxs/hN4xLa
DOFF/rhfaArFtmUg6klSVCdPlg/sqyiqAaNQ0A7xLp8PnuaNcoTndWNqYbv1+vGBjne1SWAU8nBm
EFk5OcUq9nMfQ+ifAPzMAcTwS4iF1dFJfnsOBJbYSdVxz0KA+E/EEEVxxAIg9YaNxcsoxyvyLN1i
7mN+8lFrBxRKDMFgW16Sa38YLWRVfNKMvOD78S5UFq54VejdJs1C/n1gkfqhyePFuN+iHdYsGYKW
qdxEpR8DJhBgLVY8kvUBUoZDTyhdQjJiPXxBuG5J8AvxhoWf9PDo/AMxGmx5LSibLfoTrKnqWL0l
0FSUBw0zbc+CN5Fi3BmnZZ6b1RQ9Y+vhPgZQoKi7JTIzG7+CAuDAGbEfAhAZzLJQydAsxybLTU78
OyfLOaD4NVAD+LfO9GG1YOCW/4+GzkUJ5Y5OrcTjwcu5l/WfNhw1z3e8BfTtiSqsB++oTgoWekyV
EhycQE3PSnv3BafhQTNHGBPp7MgLwyzcyqNdtUQL4vPSz4BIppZuFNof9x8jN1MRo3qoq/rEhXzL
5o57xwfNzrZdhp4uTdJQbg+cFYdW3k6o5o1/E0QNZCaMHq5TaUv9oivDXLMkiXscc9F32GhytuAO
KkqBgarE3nBT7G7FHM97BB5+tb/0J8H2Paye2ikZaWrNMJ2zMU9DY+qrFOZUZxROcnXkLFkhFCCb
FEAd9BzayqSVDFQihmU+2ENgwQYYM9pMKAdFL4RWG18XVICSkpNss8lvy0/M+ws4ZGvzHJLu/Ig7
OuJ5L1KRuIoNEK/GhnSNHS99H7+4V0Kf5acu8/RZBEK4Lni5Gp1Aj2xVyQ//m2BZh8AJ2mtcHphb
/hlvCrfyz7ID0Xt5Z9xVLN6/OJ8QBGANe5zyvw4StbyN9nMyT6awXS1UJK/3nFwUPPas2mYmDQIZ
5gvawP8bkOHP7YaymetpYzc/yJBEdZdHQMPWUDAX1zajGS/KEittd9Gv9sN5wpMfDpGd1KciADN8
7yU2rSOFukJwARq64xsNNp3LZaco6oHovFzrIHGcuY55U3V1iKJJnkJeZCewg4RwudoOVvrwPwK5
/A7h8bmGZQoJcxlLLAsZQL3K5ni+7ladNu2feKb+fhuiiZEwPhbXdaB7w3B47MUB9nM+K7qwkR1x
d2ZedWiZMjmFGRdPMagq5wp709J6NvslJACoaf0g28HJvBqnOFOdQma7eLcixgiPWzZjPWoYX7Ms
NlbRENA1CG96/++a7JLEjrM213IIJ5G0sDpUFvs9ebBhF5bc8LjPjKkGgBOJmqB7wVShexv3prJN
khKFbekf0L5EPcElcI838XrojDXik1GBOmfMaN0+GC5bKTbzkfGupXQjRAeSCVo+suJgUAkTuPBV
TpUDW54Ti0Jdjs7EpohoCn0+0S8aKLrA5n8bOYjKu3ZbhU+UsW7wEXMb7LqHyUie/ueE447D6TD1
wWdA//vbhDaux+PLjY5MYLal+pcpmZP8/KW37Y60wasPXJSDhaAx7UzD+P12Sj+aPOGhO4dKRGEU
/Uzpbk68Kxye0m3KfUR65Hdc9qopSOpoJJKR3wm6TPw3j11tXQtqlpYJkz7Ruz3JbiWt0/OGMKMl
FOCFoaBbbYLrkk7R0JVxYg8WFeJLRdurzRlC+htKtyNSb03WsscFQv7TlO13mfHnkqCHmG92etB1
LgGA+AlHeNDfgjF4GQ9W+X3Eq8zkt2hMfhNp/ZKJ/fyePvddEhOOTFyclxoko/6jJ80J+m7ws1Z+
9SaqkQLelDCCt1pbnkSe1jn2kgF3x0puQdANv19v57Z/cghaqcjrFtqSo1V7j6JjOsVQWIpvsXH5
woVbj5agig5WYnpYbq+WV76N7iKsS1P199Dt5N7/S2/gIlqV2w393j6Dr38d8kGD0bW4MOiF98Sd
dyYgvNHDjmPrZQADDVfIdQzHqrhQZGQzvqAzL4i2L5na+n2dF8oxw3o4C9StuxwR7Wg9DUsg8OiK
NiOBeN/+74YUh2ORlHvBwFe36LHIlGQbmyojR1v9RmgeUGkfpZip+NbEuAyR5vkKC2fU/7ykOcfq
vnxguvImdZqBb9yGE+ugnwNyR6phjq/C6WkyIR7e9QzznRKQC08WndHg3KIYhPJPt664Jyan3SDD
RHvcYoK5tr604LV1lz3WWn6m8ky3EXzqeDXasG8OpPe/6f8tLzKtySE3D6jvm7NzWGwCHMxbxyv4
BgsGPNAWnW5kJBptgJvM56P9FOHubB9s52uZHfbWPXWBXKm66ENRAIRZiPP6IoxJjx/B40I7zmmj
xDWUamRr0mPxpkvLON5+9AYQSs9bUef8GWdsBWlTb3kAayOz1WKEN4sp0szemwlapIczj4m6ztgu
so39IHynJFQUAFnu7z85TPju3NwJiaalt8LkTTvJJqjnBVxpL66RDbFU7U9/+bQEFq4VwvfrmZQa
xXMGBOJQSBkg3x5JkYGZa2v4THV9lcrXYZrLc09bQE8JkfIGPsyOMiBgpuveDyQzBNyjGM6hBH26
Zpqjph6D0h8gvU2/oIObTB4wbG/wWL6LqWPHI4QOsr38MSLt07YeZkbBt8W4os+mCVncANXIWofg
D+eqD4qqaj77qQ7pPmB7xOHiRS5NsrhW5Gu27KMW1WBMWoxURTjG3vf11RUTNOMJzkq8Vop8wVbp
8BqdMT7ZZ0rLQJDKqEJr0yaNAMFEwkr0SoxF3AFIxPCuOA711XLAZ96kkXzN1c2tkEzwnByinds+
OZ5FIpZ/Ne8RTtq252tXhtN+jtWxubSDyOK2n7uA2NgG9P9j7hrgxyJf2B0XkkfKKcKjBsK7+Wea
QE9aZEg39gdgSL6NCujleS7xiZa0GgaJy2RaTfrDLfnLJIRnkltAtRWhIaOfpGKEMdA6fSeMhd0B
hn0kmzLTLBPE+xc95l7yvnCcG2UtS8Cnoex43u5fdpxaOrN+jtk7BaflnJF9kAHxZgdxlo/Bv7JU
28BR0OpfWX+Ea6T3d8szYD+gQV2txkMNsyEHl1pxASk8q5/ll41A6zWU7+c5EfQFE9HN6y72+csx
slAR79nOfSsGrjU3v4l7AwNN/iLZzl7PEo7vgW4DtGfnY4QMLoJxIzZpCbuos76CQfzH8VXvkUd9
XlK2mOvfqZkIOLiLie3K3eIH7mWW6kT02pa5jgOPz6Z7H8TJFWtsOjlKtHpXjAE1Otdbe/e37vIL
dj1vb8fQOfEsFrn0vmFMWyGNN74jJ64vMhs7O157E/TT6gGod/WV710iAH6VEUlibrHT1nOCaCOz
1JAiJ0aAGJMfOX1OJjH7Bnz7GD9ZpItQETWZBdlbfrcgMbFIDKLUqxaIcHOEkboL5siYMPmg3Yj1
PRo1bVo7BPgo8Lq4n5ojeuMVquyY1ZlJUkE1YFsIksSTa1DIeIh6eaAfKGR9BkdIuoxj8GA8wCuY
fClPQQ5NBUaoFyWh/8oeORuTApmfy1FzXRW37BP9/RhwDE5vutyrFAY/YBrTkOTNOZdzXlicek+y
4ghnWEU/ZSfVLOqYbYvtHyvoAftyCRJl6wLAzyKTd95ITOzFgDyeS1sJ8LjVklCq8f5/7Mw6X6JZ
c6Hduv39O3SVepJ16trjsGUpMeqPXT1HigJQSakhapyy4FN2NxZ3Or63hbJETqtIwrd/GfO2zcjC
3ko+M97RBKR//1/atgGHRMPjPVgzmb3wJxhCGALY8t5zASgwKNJsctTa28xcr6weWEM/ud2CarMm
Yzcs3/lvCZq251SWTkum2IIW+p8am/6NO99kK6HGcwVbYn7SEzpXARWyglU8EuolUAawQFhsrS5n
hQP57hJ6tmzKzBO1UZwYHltGzMsxEVi6d5wENxGmjhHN2yYcsji5dWJOMQsIumkSUfYCA4t/BmZB
3iS1Y4c46BR6cf8ojwvGWl9AZ5p5cbPpTCUaa2FSgWfOtSKM4oZ9xp+vb4HxorRZioyHr5qYXrD9
g1YO8VODJrFIF2NeSD3oK/ERrcy7q0LC1oshCbtLtWXNTkgDf3SJyaTUA5gZRFBwtoRJDIqzFpjJ
OwEN8Cv+B0LpuqPbWJotkHyP5GWSYKmeXQwuwhkBYSVTog+UG/VTZ615SWstpOvmAIM9HVywaC1+
zmPwvfFQIpIbO2IqOGL3vJX/TOQP3ZVp81yaEQzC3d06+OcFMAVCHVUcDMUp+9yNbaNBQ7Lhda0y
Wgj1UvNhfAw8l6XSZgTtNpvV25lFAf0r9giozSn7fZiLwYAX90UmsLXbbQnYK7x4uAD+en4VW5aj
lYkHr7P1Fi4sHlaRvsmJe/9SvVngR5i4X6pM9yBX1OPuNwcuw8BE2ilnPNuis+So882N/jdTMAzy
fWXwlA8XzguuMJFkOGxWgOH6WGuav/SbZGbPkm0BBlPhslY+jPzfbt78OGkfSyxJyL8SnkoFEICa
IhVLnhd8uJiX4KAh4BPmZ5imOicEsGTFFTuiDgQygSctCNKqLEEbq58jVWlFC6KYmwBiqjdximGJ
7Q1TuHkeCAW9M45ANrrwo3rNJa37f0svvDPsuG7Lga/PTIxBNg3V5O50wZNznmsx6Y2aaF86bCcB
OA8VpEUqBX/mgK84z+1N/2HrtP9plNcrlrfS6aFZoP1TyuHfYUzUi5TBr6IoqoqR2+AJWB6hyon6
Xf467xUsnZ6k96uTOUxxSAlcBXSJI0CI27L6ru4yyDIkFv/aipMHqZYoWBCUBtgyfddXn3YZywu7
d0raR27TAfkJ+dNbUbgDbR7Tk7JvVPzqxT+QsNDg/4Su/XBWSuw6971dLVaYzKrTyULSRxG/qigJ
42BbUzP7012yra+tODDf72znwBBRYfAVOEsTGBJYML2mcpxRlKVQnE+bmtTcHYTSlBDnQznHpixb
jB3PfW9r9U4OP4PtdiAnba4zSIzHawOdIz+D9A4RG1aWrQirDCzDwuLUClt2CQzYpAunFlEWPOQH
ip2E6UdV18/CnRuvu7JJX7sv7yWtjJKicRF/rKWzJz9K+ou4wKI+wGL3XBt5MX4zJfvn/G/4w2JA
7xnMQtKucN9bDD6MNvZBUcO5Drzkq5DJ+bQJolklMgkleEM+7OXt00kiyE2LJmi1hh95cMGvwuwZ
fKNDwftNKbzhqTyrLcZFZpt7X07p2hmyRYqPyXmPkYaqAYt82UZXc+ZaG288fgwmJU/iKZafsNE+
QB83BeHbeSYc9maQS4rI5gJXQZ1eaLwjSmkFYcnjGgTRo2YUVUxwKYXn4mBLmUnjpvdXzUhVZ+nU
UMG3EM3bVt5+ygaBenlWI8FB/ExVltxrCYZY0+rhFZzBeSZJ7QmeQQFnyxpdfCRGfNtVjSswvRug
g+SGWbT3wmNzYTWoCRCgpj4LQzyl3WDqM5Yo3pWXYXNKwWbvEkqAjwlTdqdA7jnfn/0//9Ecvzbb
zgkcIhWAHjqp7UDQ/8/5lKz+9cHYYlfvQ+waV0O0AAURbRzMk86ajNcXopQcr0iPlDJ+9wLaOG2j
fN1VBejNiP6EUMaGKOM5Bxzshr7HVZkHiwJBRvcbHPyqSY300k36AiePxSjDbEnyjYosuX1UPE3N
sQgTN/lo1whtX+lhHm8NmPrN1E0ZLlk8uq0ef9MyLiXlB1vUnbwx/+ua3kDyk50XiiQ87hLQFXtS
+RjQf7EzxnPtee3EVKSx99OjwemiMbau4cjctVCLcDSUT3EcZJzkKOV2qB1UsJNm1wi/fM1WYhBj
ePVuYZQj9hks60ANKcGvU2sFgpWLyIDcyf7YcIyJnXiApqLI/USqqnqU7vYMnu4X1fXMqjeeBXfX
r9msN6iOUgVr1ahRnQpDk87tBLAHE+ztgy+IW4RkGnzZMIazTWtirmkRtdgNPEEpa+Wtnec+xDnW
Fs28WSo4IShTBAgf1Uh0d7Pt22UgiXFm7QJa5j2swhJupGibER+MSTcd2TZeNV/kmlQYr+0utJmI
l+zGQIE0ZTPeGAMHlAnD2r5tBWwMAEPFCVfJDdcilDsDffj01Sr1R1ep0Po3z48lFcpKTvP+u+il
0wQ5I2mdivRVAvmfh4N59DoNAYIxCupMLFMeuwo9Ev3uzSrabpXIuwuahGsuCYvzFKafcyhdBwlc
eYVwDzmAiHxrq6Om92Xmjxhn/VNZT/NoTVq5ZD4Y8a2NhUbapWnKcya9/3fosIHqua5xJ84AUPzv
BjxsGST0pDz27kxYnq8d3NZ6D4Bai5bYw3uikW4S/RiKI7faY8tEGsn0qQ7mffeLzzD4eVU8HTN4
h4K4v5xUxDevFStbcVJpXLAQbvC0TL0WqqTaSn2DMlWetaErgo7niLOzgWvChmuQmQ7gt5hsv/sJ
m1NWeCs33OOOzZI4oAtQ1eTLoXuURGFm0nf4lmGxq/G2gOINq3IJDJCIekCa60x97nDMxwSELMnd
lQTIolZUvKUUU0MAhBds+qEYKKI/9atfOm/CE8Iu3Kdu4/RQF8M+eb45rK6lVMl4WtmmposPYqh0
5tWwQJxrsuGnPBvFouPKJg1Z4v5VBd56xNxUPmXAXHLpyu6AjecWPoemJj5OIN5p8E9i4sh5IpbH
QMrnu028vvP0qBuCYeL1qJy1nOGYp1KV53f9tFoemvdniWG3eQh/y6JDFIK0O9EBA0Xuc8tMnR4v
DkkhDEbbu131LmKYhV6IR0uK7VPrUDrZe7vv7/s0JNH9jpLQnvPa79XwOpk0doGOJ/TzPQsCRl/S
t9H59NRba9ipeIvO61q2Rf1Ns4Cy3Wi4lN16Z/KhGv1TrfWuM2PDOQkhBbFiLI43lFfSQgOLempx
l80Pul+eZUwKzrfuvJOYj4UF4gqhp2eoUnrXL0nm8IL9DFRI7N8hq8aca7vUwj5PKIJ+ECUc49h5
Lk+zbcuHEn8n0CMAdVwJCh95TQC3Chtlw1N19Ih+uBaMVxr8CQ3jSMRFrKmWA+fHCrlo5O9TXWFI
B+0m3Deq2NTWIsJxtr86FagP5NW1LrUWA45d35LkAefLzfZawY+7hKxdjIbh+77GXPPKNK5/HnCJ
jWhJditdKrzFeXV1MW92i7tmxdui+IPEKWuKuR/CYVmxmwTaCgjRLhnd7Dz1XbjO+6eQuKVXY4hC
+UYl9TtRm1XeeuOwLvZjsnIRKuK6/RckBnTNbOZxjF8r82dg0bMqYIK42wQAhqT3uvCXP2fJ251W
zt6vfg4qA2FdE+Xm7z0vQ91XAgUZXz9eRrxGcCMijgHp3DEOtM55IaOEjUGL3X5rFklZtlRkGvE0
yU6ya1+vnfgBa8WkBDjEyaQZkhmx0mHB5D1WyXLun2BybBrpEQa9BQLu1ZyRwWUky1bU6ouILKLk
rHuLo5f1Tsl/6yv0IAfSbgJWeeHaWQd+Z6sbVd0qDQ97QwUA9Rt5aPhZuyEwHVLY8ANATJPLC/P2
nc+eEKUfxRM/14ErkPFgY1ui0PfV0H6Lvts81oiB08JPCrQX3GekeQ3TJzWynJ3E9ysyZLL2AWvf
saGKsjXmotwwGs5SLWhP2anu8SMINW+IQ1vR7exM64MY7onNrUhwUQIWP69Ubr18Fyt2qlJwfnOS
ggtZKgAO7C0L91VVJegZ88o7xjx1Za5NT1jPbOhBG8zjIBDvxq1WubNoKjSBt2cQnofIq/Az7SM6
VgUIZIJODHaQ/BJDktDhOCU3Ehmng/LqFC4XwdPShjiekJAR6NpPu7omKRA1hwgbKlXRVmH6+Nt7
pN/0UlosYAmNOv2GhUcgUTzxJAa5CUHWNgHz6Jqfa4U+Q/sVbo9NnhcPWxuBKiz7UCiJ2veTZQ7P
pUqHl0dsIG3qoPf27oaOz5W3pEnmQH6mcQVwBsXLv2eyK4TvleGwTBkbRNsCBrQP1cOriCcAveNU
Gf7JRE7HBdSPcAQ52fi+jGzbV3uCCktuxTqFeaTW5jL0q1Ow4p2luSmG5Csn7/dGFsi7m+2Rxi2X
MN7eYwZAZVgc2h7W1lPihrNRVqsE26RTvo280BnLk/z6Te8A4fd7ueCEA595vk/bhiIbjyX9bBRv
a17DRyFHX0MEPhLP9WtSH9Gqo1Js48WEkqELu2YKAe3tXVOC/3DL3CxjJmE8Lzw76wGlJl2jjI2W
O3pE7CnwZ8A6J1RsWVwEBRkC7whDeNPc/1pZ61QqK6GENzeB4sMAZqkGMmn++GoB9FL7VXa1fxlO
E9YUUXoVkIA0GKfa4Ta9XyQGeoUYC4lFf58Gi0Wm4/QH6BXIVRSRzaqm+ylvGVYKBcnT1YfzDb6V
XyFxb6oOD6a9a+D1LPF0lrRxXi6sUIde+ZMsyO6YtyfbhQA/zZhkqRxBjT9+E8tNuAAkASUW5FOv
+tsdvnxof05fP5fKZcWub+KfDUL0hs8xK8bU9d9BWp+4QnxgPxZJixz+JCPma6MMctZaj5D1w0ul
Hf7JsD7ZS0EFw3HznOCFEtXXnnF2i07IghD3RMD0NUghRCOVwgD7RoPM71B+AyeVyO5o32E03OHL
prwdt3kQCdIXQuoqrVHotFDz2ERc0s85qwdz71gYPZi1v5UHdj1O7jL/7ubqpijhAHJD1ELhn25I
4rEmAbFesFz9fFTpaDyHJE7TOBWrJUJI+/wci1xU26Kw2jHVJroK5o4CM1t9rOgCFcfIR/fTYbbo
SHpwOdDdqIGHDnY3npB0CoC1P6bUvlsbIIr9jxDZBZmaGFwr1A/XRH5r6o4PcfRKrLIA6/6IsXvk
4Oi4ZRbTgKxV8UmyMUBAII835DBXm3oIyWKpvFA4ekk4lmr8apVTq0oppU9MV1cxFY0AkZL+Iyuo
3zanhNgQEIxqEdS3MLpl1g3JnYKDXPx5Ss8hz44iYwpUn0d0JbsPG00KH4ROQSEtQxipJVQjztXu
T1wXbNnmS6Wjt3Ld84SD8dqqGIPf+IPpbalLcvNVNuFTj2buJ1cAY7K63HkmBAZs23an07Nvkwyj
JYkWkmzAtdaFL98SeA3LSH/4UScDg6sdmuul2n44AJ0EL6OSmZ4gEte1QjcFAU5romoSVWx3cCDX
tJWTbgd0B1Ib3RTyE+/Ov/nn7um1qt9QiGVwG+vDqgCU00fuRfKpHnkfY+vi7E3BdBqb5hBPeA0j
BGZO8vFUhV23VgGIrC10fOudMYnFyKytc85R3C1aev7/davaY0qHNwwet6knn78BJ76Yi8gc5F9G
f2Tq6cN607Nd8BRRZYMXunqhdNByQ7mp/F/1wDta8tGkMH3et8gMjr35SOkq7IV/neOKGDbC4Gn0
DuW9jkiovQiMm/N/z94jxRgysiyl5HyDeQqCIjaJ2YZtZiIZNxDgWx22GCUcGiLKSx3rd/Gnn6Kn
4NZc5KCOpYvIe9AAtNy/TW6bdjpXL3d5ZLiZjDyHmjni1KgVl6NrcJ7Bpeo3ZQzMl7k8fXZ4VBBb
wfhSgBiw04PeVvGgu9mCHIGNnjF4D5ZaIbaoXJoSQqpdM/Dnt1QRmXJLjisfF1got9hteGFogGev
RvY8AC/061yfpT0IVUAR8Wo0EXrufPO8dOx1sj28UX/5jg9E+MCHwneMLM/QVTRQqLQHPqcW5vup
Yr4/AnyOeIyEQyJL+hBs9IpdPX1LFbxXbG1YRC0e3Az2PQYHe/kAROST3sf2w98PFchUxd9QlXFZ
m+MLPVIRHMXQ7Puk13OM9dS0eQOMQatCuh7BzSaxXGJAxaIHaAE+vK+Ww49KZ5ayHYU8Ks6RTQIz
qNkSPyR6x3EDrt2n6tlwBXXXmyrefXyYHDcS3DT17YdSp57ji1Tpurr/P4soZc5blH4ka25Fw421
NOpnQ3FGJPVxQxoTIUlIZuE6DJ0VBmYj8n+6cimOTr7IhneW5nNh3wuSaUBp4TTek0/4a60zLBfY
rZJIRRIUptLCTfXPM72z/O74SIVWNMRN7wU+naQAm7UlCFhpB1whlQf8FTjk+X9qy2cRx60eL2CS
M7J4583lLh+YiVkOIwmYYzcPy4hv+Di4jpYB+V1smRF0KTfbndXpnim85Lc86l0IjrNBIZnHd+zc
lQeOnFMsFD2fU4+aQ2hM0PMOTMUYMQ/g9L2kcs3EGcbDEds+89n0SFmvMhrBNzZ8EQF0c4rOK6kU
v473xFVN7nCvRruUaEDFMQZPQpWdfoXf9gGcITBULA8EV4y7VWXZhTwE/V3BFs/lbqlgjNTcOD9i
q3nLYJbqIu4gq23/URqCUSEEvw0+XCDO6bnZXisrLvgyVAe0rsJ0OvP0QnKJAihsb+0E7H3YWBL4
DW5eK8Nl4dlOeNP6oTSeoxdJHLbOkRbutyRCdM0rF75II33lM9WpyfS556YwdmnomFoUrKA7y2hn
iitLGlK4q0DGTrodhv3SUJrsR0L+BYX5r8xOR6m7n2tTzGNkCjEH39yJT2pJme8VdnF3SNgjGGUH
ZYCqc1cC9hf/iplojBiJpaLefwSeU/tSHqWHbbPD8gWpy+zBm+Q2kvgmS53anS3WY7k4R0H1hHEw
I2lt0UOchJ6lLPiiQv/ndUalit333zPwDB6yQaIUZMhvX7+xQXbC2yrrxKQly0ozwwkzKlb0tycj
9rRZ4I6fByU2uQ8cZETdRRcIP1Xhp5o9kCikK9+3pcktcJCQng7S4wBJfpoOpwp00q1GcZlpPSki
8B/NtUzuD9oTKZnmid7cuwu4/vWN6BrTleQzhEX0fdAlKakSGaoVmPtW/eW2wiBRRfPHzZCfDdi8
uwRHhFdVWCWftFCSAwpaCGlMBuoXJxqpxbXkEonAA9aWXqw8UICrwQt3ekzGoo5KlobZ6+1cDNKx
L1shHBn2CcRgFZPEdwXnXoTPs6weZ8DY+ya2FSonE/poQf00FqaqMHi4eJjB4ti+J0/ljrxEdXKp
15lOs8Rz2AO0I1vcY08l6VcRmOfSa6073hxHy4VKciBUW8egMfE4wATqldlKOrDSw9S8Hrow4Nn9
sfw4+kq5PzbF0pa7/gtZbCN9Pd0T31trF/iRcZMPMigD3Z10JSgO7GZ6+lQy/FqdIm64n5Pt0qTK
KhjZuq6kRTMjWy/Hp5EhIAFr8T6oTKjS627sSLd4O7reIbFK/KxaC+sYBMqbRosResQ0B92X/A7/
kV0FQ/IBOs17EIAuhhtzt3IIyQjdUrQntYnY6isaYnsO3/BdxvwZmU5tMpdwJAtNXietAct1+YcS
Hw/Hw8KuOfjxV6WmnpV7c8MFFbqgniF5aaEh1NAHC5AcEJ3OuADE5DxUVIA8lrAWJR928F1irLcW
On1/L6GqHdnZNc/RS9Ro8ZX0M3yIVx4/rFOt3ArVkc9FNXV33QeEcFNM/JHSEoI7sdt/HidYr/Vy
rp/PNAJBK2MJIeIk5fXZ00L04Qbfn8uFd6kfnKB0gqXYC8ZO2vVDYb9Dr2iT+TPoer+1Ep0xtn2H
Vk6gEJ7kwGb1Aw0XnyenCldnm/091GpBVotce2JGftdLzFR62cA2Qf+nqXmNFcBC6eMe6VmuJEdx
pxrGT2DUHSWIJhpfPhLh7ClOiWrcVk2G5vJG3RabnEV29NnliPuQKxucl2L6d7zII6/i7KBg7XIE
8NV32r/FDRAVpcwztf843FtaOZtHr3M0xC/2s7GAuk0OD3VR+LUXr/frtCw2zuWg3C0cupHsZSMO
448uRVGdXPdvU7yNiIg5Kb+VivzTBfck7vhlLONgLwlxKhw0TFnoJTO/i4HR6BZ3lpTm5Cq5m5AH
fLyWJS8jHN18de3igcMce9gXFitsTdFx4aBOc92197o54J6IFdsZZLEXAD1Z+j0fTQGPKpLQU5BQ
/9clNURLwRkPFJ0vZr0Tja9jSy/E+sDrbEqjiszP+dEgPnMUr4btIm9p9rzC8n0YFfIpQPPdKF56
SWoGkD9Teqwp5OTbL4KBkFJQCZ3Y1U2kOaZsmarWQg6WxunDqx7Do7Tja1d5RLz+21F30vY3DRbJ
C4ESR9n6F3XIIQfc+Dq3VoC+Di5ZLhOQoNs4k/Z/LZYytWvn2/5GkGdfPC0uZ6hkDGdH/5/GH/xL
dJ9kfnaQ+BN068mbH7yAheQcMwWNApnCz1Xv9iYEqWHktCSV32os0D10RimcENX7dk5gApNyQO0H
dzoEFpuL+tBa/Z/Rri1jVpNtMcb99AvJZdPMU0/6S0oSlYT0cEyn6PeIbE0r6XXZMoXHIhkpEMmC
V7sn5WFEvodDfxYQoc24UAGhHl5SrdQxuoU5EYur9rq5dRteGKMkIX+7bXgMFtPEb2Pf7N7MiUV8
hD3HHfvZ0B5JVci3le2d4Vsa4+hnoXV4e2w+5GoNTL8b7cR3m0HWmdlGDG4V89Mm8PxP9ASByYhz
kcLkYWJKvkF6CK7XNDSol7l7+rmkZbTdyOI9JBX6WvYb5E7NgRhyK7vIOJp3OHxzrXR/cHZ6l48M
kgtOdr91EZjqTl+WB1OjezdCsCzPYhH3sjfSgHUzxWOWcGZA0HSrTduyck5pbQBZUHeqDGtRtz9V
dBM23HQml6qHUkonfStUuubJbcfV/IRGl5CchoKirLm+ueyHoZUO9acBFWTuB1yktrDmiVC7ixYK
5u2aPpb43Q2z6lOn3RMkjdodITd58fjMjsY8innzSdMAm0Aqi6qjakGKje5wQGyefjDek2NhxApv
Z0ofPvtiquNF35ICpmDgnOPtPcKYLKkiv77H9TeRxa6wxPi20UFDV0AEB+8pEVkgTG/TM5q6Q3hL
KNfjMoLHIZu6MlcyaQ1OefS0YoNFlKwL9vr3TltVR2FbijrZ4W4IGnYQW9ty1G8whusJqUCWdKLs
XxCmZjOReaqOUk06WlJz9cAIEczErTJVnsubjT5sSI7TyD2vihLGH7MSh2QTykILIV0qZEzv5hW6
l1eGd3dgR6WD80LyfXS0kCGYVdx/IUTo5/t72FwlmgLAwKQPdtaYhd7Dx+dbz6vpvNPWZgvk7rmi
+FwRn4MjksLl8zjRG0wiruw+JKcy/9nk06eAQ2ihpj6XjdRPz+fzsgb62/7YXSdF7xs8AoZ9zZTo
bZRrWuBNkO5FNnqIcOuU/6Q4U3XabfHklLJaZTARQBveQz6kNLlNW2pNWmSkawkIQ+OlSMg3CIGk
BzxTuAMpYzdQd3hxBbl0ACCopZHQZJZtSSC6VAkQAY87jlzwl8RzOYWu0QBP1IOoN6AFduvTPVNs
9tuiCAW88JLnGY1m4Nic/U8BmBV/A/zOpCLRisyI1dbwBaAzAEw2vSn3AUUPDntufBqQwW0Y6qZq
qI5l9DdSNRjKIQvJTURXACC74Sijf/A3q21Z6FGV9icAqaJVfOkHFjMAnyUupLSUdOjJlGXHj5v2
ZUaJDjD6LrWX6RhaoViSURDKqHEDnle+TWqKwsypoPbivuXkVJRDyCLfCkMblkKSlLkeaMysMnCv
rtXz+Sx9XBHikXfdeFyQwnj7Ni9ca7axCw1HOpQ2fudwA0RGiKRjbgYtF7AnNZxZRnHD+S/7BnHo
EmmyYkywsEVm57v2z175/o4h3s/2e7UECtN88ZTKq2P7adWsXnM4pdbr9SPpkxW82qsD+Jd47gif
Vz5BFU4k/efMXBXuVLrYneh9ZXW6PiuqgRxh0FmeNSKXuTJH+/Naw+tiFialkxqhdvODt3Pp5I2R
O+Vba8AoRGuTY2USlA5R0IXiKk1cHADj0h8p7tjaO7+KvfO9/9bgEroF1co7T9sN7dxyxjltAPvf
kyjzz1RsJJ7o+73Dhm22UtveKjHekE3Nj+kXlgIg2QbAJpiK4hxLwjqe52jq+3c3uCyXjG4KeTkv
Z6yO0p+krKAfhbu91qcuGxMWIs6rr4IVa8uQ1HEZjQP8wgUcFwbczlC+op5QD4H8uVHN15/LGZ+k
4LiMbqA28ZNzeiz0jB4sRl3VSAcgloVFihq9eAU2wQvnIZXhGmYl9wmJJnYXqXEcKmRgoQtMwTXZ
a+jCLazmhsk77JcPB2+009VHFqqHduLhuY2PfuY9avDQdIHl69TRKY5JoUMd8xAv1aDmBuBB65+8
pHQs+q34taNEgn2GBqKU/3L7E0GwiTdfGNDKF4TmaslqWiI+5Kcb6bXvnbJkTC/VH7WC01An3R/W
+8Uac8+kCg9FGUZ88qZ27g4zLW6+FYMdB1qwuUvlKdLzk+U98X1r5ihNZS+Mj0M96tGk4bvzJGHB
7/KjnSzA8d4i0tsQ78CXzWnCK8xCX4yDOMEXRgf6Ix36RNsShX8oe8EhD2eiArjcWK/KuVCZp4uK
KynqVAOsmcn4Hf3ESAnj6VBGDssYWJlh6prxzq0b6NWcpKrDe+0T9rE2i4TQiTWhbEV5Y/u+/1hm
YDtlrn5g7IXCAj+6dfXWTGGBX3mLyolrqTuRKHSh01WyUV3T7H32eH9WPPy1PMwwCIfZIpNBAsH2
vBBMZbzLcg8wFoTP+MQX5NKd/vcIvh8QymwWHf7sjcUTGdbGi8Zz8ECEeQD9mxOv8HrAhtpjEZdY
VdJ6oCosRcahBziGt6oeXUys9GImyZXViN5Pb5c6SjpFhBUcRVTFUIKeYegD93oCAiF5/GP1+nEu
bDVndbP+MhAO3aPN7sAEXqeCRNvgAN9HPxqm1IlqyUpUJRG91N8C79EjRdC/KwnmWXkYQcSRZlXK
z7GhhbK7P0NKTRrqgG7TE121KpI6Rd+DnrmOt7ugNFtPAr8ocx1eaLwLuOzhwky3rDixYhM6RP6L
uZXqA1IutSp6Bp4BacOpQkUpW98xUrVrY/HvfB1fqopz2FYVTU+xAf4+YUkHeEpNXP7lFzSgi3dY
1j4I9jafRfPfGrlFIKH7f6uTFeY5/9TNd14DEkBv/7XvdX6mwhKKBgdIZ//CYIiz4K849JPAbtpQ
BRpmiVX8QHmC8XqkXqDmTBds3+DT2su8AjjF9xjh5MrwCdRvj51VSw+Suj+njS6UcODn8bmiXTvC
7mrmvqSdifc75ZV+ixgViR0vQiRXPKV++k4nRvpFU4IptERTR3h9umitg13ICTXB53wkyyVx3PIS
5kgTx3aSeZq8IvhrDwewT8LpBmuQr3FA1B2KP9ku7CTsuKH5l8O6ZlStFBKQHyyCfPGP/n9H9GnL
A+3Cj2r2OTHCv8U+GJwKBMD5a+MJdbxBWUewQGrB925QvWYoQlzQwNoNMUQRoyKvaJqd6qZ6sm7m
wF/Fon1GQYQ5aMRnI6ItXLe+kbC5rWVjedYjzSvTcKat1Hvjefmtqt9OrK9f9N6Rx7lsCSerj3cS
z3x9zgS5lyJ3C76nhPvYEFK1f0W061jgFdOkydIiJQlldwiV+nhIwmYLfoOmk8VLODEcFHK7nY2w
F9IwYB/kP+IXUQfj+GiUkRX+NlPBjjGjEG+RhBrq6gj1uXDEj9LC4kuWrSWR4K633jUgsflwjUAj
Zn8yMnHSs4IGtJn+odgq0dJkR+jXxdIoNEJeZ0B14THVVra3L+72i79YZBmCqGeLZZgTtWDd/A0a
fUmb9RJIG8G3lWz/ewwCaWbmy7soeiWP3cRhtVCAulT9NU7/osbk6ckzhQmyGHPiB6b6unMnqfj5
i4ky9XEGn1SqZUCHybvqR0Ozmq3beybwxPlpadoVxe2cxTEG0t02SGTnDDzygr6TI+HO7/4CV1Q7
AnGkErUcDzuogyAKY0Z7zZKfe7XOwojuUrO+fQtpHx8EfNtRCvFyl28qTScno0LUOHYLGf1epsPz
ydIDzqnCRlGmXzi4g2zA4hAF7e5cnRm855dqnBySLG8mKmxBnerMn5R4Zyrl1TAeUSyBTVJKtKFw
KSxenRhnciQVHGwOTSVTQNWDhTrFDH2yNej9OxqTy1Q73TtR8IuX5u6SEuEO9hqZLacpvJBAUptu
CUmvW9ZVuXltiaxB28aG2FfB/UZz8VzpnZKX43ivSX7EX6d7zT/EXsKUvm4+UsHtD7EEZWY3rsZ4
uNmiqO/aOsoTHVtJrPXHWA64zhtHi/Chw9lcmr4bvNmTHmskV9a7XrkW4fv5cK8fTdsTw+g94ksb
4tSqL/41m+Z9dghygxgLUv6Eu7L/OLIJwxnuJYL+CKeYHp/pisITAOLG2B8SmXHNeYLn1L6GhcK5
FG1CDEKkPaJO176oI9/sqZf3nRDuzNmCc9e0PHVhJIb+BSKP8/+r5ivqLrLse3KMDb53l3MXjjHJ
4P4fGi7jx2ntVQSdtkJbinopfwWZGxd7PX436CV5Z9X0pr/91UO2BRn0qli/4AbhbOPwPyzO13v/
BgmiKr+r0DhvzZuw0YWrCgB2nwqkOdqO6rCksaKzC9J8VQeCGzY8jbhVsE2YFCQa4k1lw4rBNLDC
OO0vsbZgiP/JZS7r5BM7iYruMU5Q1mVypTs7QGjsGwH2DDrN7Hna+zJMtl7vphSrfr/B0OHwMmwB
+yycIYXnCa+0xrtL3ubKQQESHQfDbkmoHMuXk3HP0W3udYNOXij5h3jVwTtQU1NYENNo9AVIoQm0
y7O+cvnYXfEJ2EkI2Vh7icIgoAXWFp+7BYoR2mTYWG6KPz+qp/yyNQlNNE6ssJo/BB6nkhpIDK0I
lymeCH+mLHzMDxFfn7psL0gIVW7wrVxHe7nyQ/h5TGkCjiwE9CL3/qX5c5/MsYxZVOflvv8GJz6U
66poiXdDzozT7qbAGqCgyNPCL3tGiA0CICvy1MBDRoDBcErgzkv3HzSdeA+l591MTiYPbwH9Qlhv
emRDpUlBRJopARWUxiypSGsx2r7ueXuyTnML06MIc0rfE3YqY727mOJ4VRbcTTW0rZSmlLdI1LrE
V2p1hCLQVGpTBMwPOJhBgLIT52HU2Wljwz8wz/YyrkSijaKGRouZmSELv3m6pOwDQKecEoZNUGiX
aaUYUgVKUOGRpdTJIDg0N3n9oS5m0NX5kETkXn/es8AU9lFH58MtEhzjWKfqnkck4I/cV+EfJjm0
GjhLP3LE547I+KzL7ZbZBN9Rpu4pG1kOLkUtJn5qsTINgcxr8v8XIckHSEUMzbES/oPh2Pl9NLsX
/j51jF83UGip5w7+/DTDz8Y/+mv+DOhvvnsbkx0cZZsxgO9tQKRrhHRMbxciIJ4poL8Zwe1rkAKM
ukqh4Kx+a+/8YEh1RPYHSxreFx5tT7n7GcKuOK9WtxtbkOAoOHD6gnQXkBeh+nxezJqZLJVzROP4
U8CgM+cNHhuMGKCrcTgVXqwio1+x06rZ43hO42ErCt16gR8dO8yB2FFJxtLndi/6E/lbDN9diATg
EydUkVgCAti7EHb0VDPyNT3uj1wouhVpI1+qPVGqaut73ksrK7YAifoxq7Om8hP9ddMLGDA0jvwv
yN4EPEDy221UUEUM4ldOmxl/D47Lj2cLLmdkevoytb3lPK1GETt2Mrg2xSUF9rcrcyoT1jFDbR8e
u9CLsPySWcx/+dFrVE/hxW3HH3h8bFFFc7ITDepspWENs3X78c9oh0usN1UyAXyyHE0AkQmM8Wzk
XQ1WFDFc2y9tZvFvvL95ZwGCxu6z3RjrxzThrNbiIfTDMhhbKnW8g/DL706RDSkRXz+n4QBQmKnj
DRxELkOlV55QI+x9KjzjQ2hqIYbWtxFJ+bkIansUaODE1vyLlkw9nNe1+shX6LMKpzkXgrqnLUT3
aMXDhjpWVPia0xYsH9XHHtHk1Vr+ZWpYeM220ZilEStLzE3e8xkQ0gVRfpxjdbz45f8jR38kJdZ9
Y1QDWitp8lcYB/qTgg2R3TfCSZeXUlWylXeXKpTRZJ27st4UbuihlDsz42BOfrADiwiE1y0x5ci+
XNM3in9L6yAlyMx4eGLWDgTscb+07BuD7z/pyBr6/LY+GUdQp57Gwqhwaomcx1GFWQjlR/jmgIm/
nj//9dxqvEeTpH4vemfg2WXUNiOkCBH4ImqDcY2le25VyvruuEjA8oF+p6nPHn9KjQ3zB34+zjFO
XeDQJ2POhnGNLHa98F6ZZpL+ExQioAjv0dGzKRcqSMd6ODaL+bHY7R2QDgLvbn9Iu/cE3Jh9OXAw
R/Rt2daEknaAb+yO3e5ZvuiBvQxMIE5ckE3L8ptTyiWEm1LXUIZcWvYzVhxGTP03InJ2jLsxs5qE
pHd6/rIs4bUXr14cs47Jnid7PanfLemTmF7UXg62E6Na5f96acHvmbrW6vw1inbAwgphrWz+6KMP
7chZV1LqtEXAIvUG2U5ho74bevYmjivFZjkGg2AD3e2tpIwLgNEocskgA/fCJHt5D3Bvslq1sf9Q
YuB55ppGYclpeswR8Ul40jRJwsnjQs+m0z2KHwbAZe5rImBm+E5B2blaZzXkJXlSgdwT+WtHUcCy
jc53FfjqP+uqxMjE2Y1k41aDfvPvDOGsOlDhyEBRiIXWtLq7eJFvKQasWN23dfR/gZ9oSaibWb74
y5WP2mYtsiHyjnFgiahF/1BsK6K88lIKJDkTeUiBQZiosQ6ycZw1xVERB2aCqtv+4eSLOfBltO2F
mUPD+0pykjJXaUqFMYS6tmlhXIFa3K/xB2cmiRgAJq7tmUAfBFLD4n/TqiF/JkAPRNw32npmb3Ul
1vJACP8IBvjugoJSEPbdPwvm3Z6Kc0WrRYEHmPosYvwfofKQnfQvpwBtKpMI8C4bEbiLlOfryogZ
X3cJcutKpjDU4dmLc5hCx4paen7qVuv4RQhivTdWuERcmhv6iI01bORRwoPEQlwkx6xDnNoY55HD
Y2LxUqMEjxAWgfHc71kAmCXFcmSMdCN2o9MgdJ00IYM9Q+jrp9ULN8DgNZCH4kfidEgkOr2TL4z9
T43LI/iN/1iUZeYHzuRaWyfJMrCq/3kfM8O5ia3ODcbiQEXmIECwKHOTn+HTfP/ppFdLwYqepEnn
0RA5iNOI1zeSq5t/UZTVBMnvhqx8Hu6Vj+0BL8yyP9UhdKJMzqHg7VwWECIIT0Mq8vmKtPDEhHAh
U3Do1ZJHrcVsrMGKojRziNeBx7kAcMSgNcG8ORI+gJ16FoDoFc/Ec9OtsZ7ffR0fhGl6DpRjaV3V
6fFXjMHz1f9bP9d43Bu1Bx/1Osn1iNc5HrKZI//zDDDhzHJbN/RnE0hxwc9KyDN8vNUvNzlpJ9Cb
IuC+vl10rID8Umz+8Xdm7+Cy5ItDSRDAimp9+H4fcwbhMqDXutWK5BrUYKdY4OJCgO7drDDPhEnZ
zS7B0oLPCldio/dZEMbUhs11BsLqmleLwi3yO49Aro1I58txzps//JI326CICWlDv72zGVMq/qw3
iXUdR1WqKfx++kE1eaP9IX1NnPp9OZA38BgjmBtFIoOpof0y1ohdbAM3KYLySCrzZe/gythVQRWK
ikxOLTg5WyI2YDHX/JkkeD0DeGvgfh0KjIrU//Yt+3mL5GeImfPW85TKJ9wHAIikKcRr2q/fy5JM
bsGasP+a5q2yZ0JOHGyG1ZfK5OaxBiingE8wVfAP7MMCJzl4vR8zg0EznAt9y+sygEr2YXHaWdn9
BcCxeOiSRi5NXleAlvwLkzF8L8MzmrnAge6qKLkrgqT+qlfxdEb9YeeegMqlOMnL1Oe7denxWlUT
VTwrqLGagCPfmXZg0/v4iNbkSQIXos75Aqw8W9LHYGzZ5q5PZUge2+wV4hk9fCH4Kg4UNtaCwYy7
+UG+4xm2chJPnHf5ZvZCtOnTUX0OA09N/wWUmcINfRkPT2m6B7V3+I8WQD5QNxdqj8vcmHyGcSnT
fPvrh8V8UtuoIV+oirKJpX27gdE+p3tfJqA9nktIwjs7xRcLiEuThJt5kJwtWaCx/g5Gz4CxDCsY
ev14b5gmMdCSdQDHEAY9i218OyvJ8CMsa8ZJ3nBRIGkOvPzDxSX+Bdj6ctBrg5n32kF5Ondpkp/M
Jtn8iO92Qf98k3Ab2maFUz5s3dnKVYGMGM1SlCYuVCMwno2v31jSCWooDrVXX3snMrkhRsO/1rF7
jea+lzcEdOZQp6zLRGpRgM8JEYrITiKyu5H7cfer5J2saJHn7APNZykJ3Igdqx6leuc5JaX6zoSO
gmP5Gw8SB8bycCIh+yic9mVOT0zIj8TW/09LOMWCrvfgYj6NtgxCyd3DLuV49ly3ahjKMKdd1Fzd
SO5oqZmiLvlmWXlHAz6DCUBy/V6PILqkW0tkOZOCnHiSF1MwFCkTRBF2Zz/hM14hRvpqHIiVQNv8
pk404iZ6nrZztcGkuLke1quTIw/Eq6sU/5SzOdKjcnVnhdl+p+N3lbXh7oTlCcUJ6q9FcoKHLWwy
SiNJwFiLo+763tswwQZiQWN7OEWn/jiiTnNKRJpTFr5cqXXsF7NN1fS4pp5XssQFOEqGmVJEXymV
AV7Bq1drZLPs5DxrNWcz3FYIfOtrqUbYgvW1+TUgxkUTYYsMUnM+QV5vw4X9Ql6dKtShcqCNK62o
5G876RWFJM3mbQCGNQu6fxlpzn0iXcUyflf/x542C7YQsC7dLR4CeKnDFLyJmDZS1qME4JJcaqEj
ReGZcDAEEZpVBnJEKzfjggDPY48Mmx7+p3VnoHzez2G5zYTmnBfNStf893XBFOHr397v7Ke+basJ
VO7+puZFDy9kcYeubIiImE4CwoCOnmTUzO/uLKVPT5ZMck4gBI9iIoADowIjIcjI2+HXhWeDTkdR
CiaPqgNCVpGnO+aNkqPhH8Wn9msFVNlaP+Dl+Ljfel/iNevkuUGoQJ9ZvrvU9oqKX9lIHIb8iXsP
aunCvpd6up95pV7JKxo9ZxvqCERXzZ9aMOhPjWC2pev/Lonn7zhi+Pn5bhD0Ty1RDHkFhVKe2Yp6
kafRthS0OE8BCpZ/L3+9zOpQDHpmT9Ww5X099J9tmwEFBbb4n3i7CpdHQcO2LKvN/yT7oBcdaIEb
S08mQ12osKzK9OtG6Dpm8VEC2fetAk8EtB5fKuEWNUuGmY7bFyzzDq4QpuVlbmQLZOB/x/HVQZ6N
GZWMic14HmpNNNhoXCKY33eRTmK/YLqa0DVoKcMvwHNB75itE1Nc4SjAVYjqPrgaW9/CsyRou2Ri
VogcQTieoQSLEqiaceDqBCbJB2lvQPA5lkskw6H3iBilEot4u7aIFNAFqZaEY729FAqtE8ZhEKLL
mzHlx7IqOLbTGKKBgHcWz+Tlq3CXUCRAz7hjcZCFoKWPjK3YJ1y2VcMcsy1Rz7BA9dQ8UTaFYjoI
estx8wYvS/Y6t3sGlO5TeXwF6K52MCQWo2n4QRp2h4NNWCahmapOJmOr6Z1kh8Jg8vWAfqwf4Y3s
WX5DIAUNrSfMUVsBA5PO3O9mvxWfwf3wrR2RktqjGJakjzk9BGxREFF9JzRXAy4qA6dydgO4Dcfs
UNKcqjaSSZvQHjoJ0naR0QUuI88MJ8AuwUpW/ugGSwHVIylTqJU3FUsaLfqS4XlPttuP0LqsIguJ
7CUNjh2MCad0ne0PGGqaVKvm46Q99PPo8JLOZcCXtLvLRtSbjvp0a6M5IH6dF36f24/NHDEwHYCY
LpqqQ2biiU0OPLj+RROuB9xRh4Inp8KxHnVDQtNOF25DY9l9u0z8EL58Dj5qaJfOddUCfmvvoIg5
HmVK51ScnyqpExK7wogLH2qPD9ZBEJ1AkT/5WmE77EsR5aEHh6onZgrepMt2Jrx1lJ0BVdvzSixo
wiq+ulGWqJj/+Ufe3tcl/HUEElgIYJaxuusRywhAnSRwRVP6WgbtYtFIbS0p0LNB4k7anP8rDzSO
gJZyaHdsrDAQeZSoILVjZKXMFU1l2b8PVgtllh2sJSxHPeiNk8ptprIdznTijOUa4Heow3ePIPLw
5ihNnCigJTi1w1VYhRkJOZjUOMqRyXvZf3c9Fo24O/qRkQH5NfCF97ZCL/CDaNxH2s3GttJDXtX8
qa5xE0SRvQj4K00z79H6bmdPsOSrDBCJTEOAVRmVCsh5O6OWcqlNrpatzRM7ZqzhVt0uRshoaDde
gEKmFIr2UL89VEfj1igHLfM6S2Wr3Oi24SsvhwwytY7C4LHelLqG9abmYaxrjoe0a/GReFrglH0A
oOZLXUYnpIOAEIi9fRFrfz9rxm9aHRdb9PpE5RWXbh4WYLJC/Xljr/89CH/ROQnWXw0Zd0geW2+e
0arOAgujfkvAU8DfyBjPQN23+SCjW3RE+vYsebAMNWc16X45JuOUmrkqdQnBQogK8lnLqg1WXMEN
AamVbSzVxbrGvbAc7LeJCRZpyeD23N6qV8Nf3xK27dcXuFSVXmZI2VxMoFtRYNFSmPtqVCGvwjmy
WTqIdTFrAW9IVOivOjgBKcZyc+q/gjiMgyYyqINUGiHdX2xamBg63Eim/6tZUHx+C68R0F48YV47
jRFQKgeTYvSP+nI6dIOIk9yDyxHtg8FbugXOclOlG0bmEp9jCa/t0X03uDXnypVnF1fZgWXTSA1z
Xi0yLKyFORcgFJcKyF4dl/7DeIiyaMcQ1aMVgJf14psxL6bkGmlmjtPTaquFPIgY263GoXcYhuNB
hJ18k5/hkgcpT/BFEux41hWmC/YzSLvH9tW0IM4I9gS+a1v5L6wWEdJRN56gLT4V0YRQjM5c3911
bzGXXb8tewTJqsGZR5NkvfzMWsWKXlQssfI2/gJGW63yUipADEU3ohB2m1bjsFefL8ANmXcHxrXd
nt4cI8ofBaDXOfiETvfdl5x3NcOVVCcbsFKlQZ7UmGIuKQ/7jnG+gI7d5i3k7Ey40jDTNbQzv6Ok
9SX5taCq7qemRE5AlBlY9O7Wxr51XGieRHqfLYApOIERC9h9lg2y06fRU6AgDI4F8QdFaY0Jp8qg
jazYQtLXySEUJNjdGzuCb3p5fccI51zekY8AJhRfMFiZ3prUWXX71THfWILezy1cDXXQK1cdpBFJ
HKHYZUuz/LEIy+C305uDUMoEYt5jTgI65wrPfBgPfqWGb3dHjoWlgq2W2IvRaDZ+rMTlDhRdAHf3
ry9purv7s3MVN2IfhH7h2oP5PFA4ksSp/h6rKQeb61hxoyDuGddCKBePy5YeSWbYPfpp2N6cDOLG
g95MOCTe/zBQ033GmaMO8uyXu4986pROnGISLEcnIjOZ/UfIziCdhPbwQXqSWTQanqVM4Oh2s9Po
R9UYbdmWCp40T7J8Q7dNsEQHvEMDwqc21I+0s+xNRNL5MdwBt0iZb/PsYKBJCkmacdHkNAS+OdJL
wE4DPAmvORcbhIBfyrle2JylrMOZW4PG0sjA130FKxw4EktZxa8hPgNed+Vjqh+ExOCPyJgVA+mZ
SeizeU6e8iEFmSdJQ2c7TDXOJY/vU1G0YifZ2YUy1KNUbVHYs4S3lDXpoFFvOrHHbq9lmXzJjXB6
VOdyK2FLZapPWmLtKhebvzNgPo2Z+4wVjLQyf+NJBLfpkFfTIchMzOiJQzYc4vK0dKjj7eCeGF9G
3Qiaz2sBZCSbe8Co8jWS6/pDZjUfwj/fLjBHGyu+6eh6iZmhA4288XQ+FRhwCoHVtt0IaqVYXGky
4R8slko7f3tNTMKIJ1fmpYPPOw5Iu6FCehg1llt+a/gxnzTVgryHRG4XXH6/7/LWhf1PcOelXbEI
rw4vhHWuVo4kjXd2BRn9o/YxVDQsFU6q9o+8GLrECENLjlNkMBjsasjnfdE+6vR+hvlpuaBBM4Tn
t5VSXvV3t1H44WqULQB08zAmCqDJymFNe6at9opJLbQc3UPXNoQyQw35PctQg/PYf+s61RVDgf45
fVkyV3yNu+wdaBDpXEU/0D83gJiD3bBEID06Dc99K+rhh/boi8mmsoZvqsjfLPP1rfNmCqNj2T+C
pMg0xnct+QoELekgaeacxbreGIVac1o8m29VD3cbwJuEiZY45fYhzpwPdmL41VCJAGchf1cWl1Yk
02Qdg7xHvwu4wHkE/blG8cKHDlycTzxL55OW8+uFttG0ow15FgyRbVtH8FkyAQ5F4EFl/DpqTiuw
G7hhsAMo52aFPYapGI1Fxlk+Z2D8qo672xPf1OIS9Cbdys/3aH3o5EiqtFaGHZ3DE4X2ts2oG/lf
PKLxZpgB4qh+kcHx83ZkeRoN7/p+v8obBlna6eKIkJsoyL6fMyepsCMxFhIJICym87c+xLIkJK/a
wKWKdIkNGiibs4M9SOJ6eyIIjwTcRf8A1kXUCBTZGDY3dBdVDIZCvqJg8S34rt00vKsjDKNQ09o2
LriMGBAJkjFy4uvfJMA8XugPW3mjy4zq3e/jrOSVFHqvqw4o9DRBVIJlrpR6+b96wpHdiyHtJ1Z6
rcb0PRKEsbtk5yQqMFpbCei3sUxIDWN9KdjLEhlp+hbZ4Ltnyg9DiCc98UbcXmgW/kuuGfDYWIW0
IiRgh1PwxF3eF00WN/MIw3CZhqlCjuHJdGYXxcgyvDjjsMKspTXjb8PGGYM3SJ6CaVAZ9IvVhK2m
sTHDhtr2qZ1l5nP44Ze2G7xZFHcJbeFJ95CUZvedK8UeVRiBrtxDfAmTYK0OIAvrH8/I/++f7GzN
YhUFITWWVYqP+p8Cgh8k6thyTaWmIWnBp2GKBsBXl+Q0n2EVeeoXccek6jVKjUASsiKdmvuhjIKr
xXkQ3jxrQD7XWaybCHCM+XSBeDZpwxycx3xt8CVlXX2slPuoUg0ZONadtGdgFp4h5WGjln21Sb6D
KiQkC/lnoM07iDLWHB4bwK+TYJCoeDNMNiPBKpjbDnfKPptBUzITDeDm+kL9O6y+59cKE8Ydqt9+
dGDrmONvZlKznxhODJAJw0DFSOdpOc2e6+489jjjHMTpS2czOsIu8axm1kz5MDDVEJGJtoH1hIYu
3LeYbfxB/h+v8z+QI6MVNmL6rCHLUZsCQwo62ww8QaRNBNqpPvqt5A9+aMCx9NPmuwNi8T4lo5mZ
aq8F+f0fBe3hgIZ8CzcB0yElfBSJyI7GLsBlR2WG7YGAiffnHrswL3KYzmdxHFCgPtn1ly/RZNOT
yvctWNE5PuQy22lwa/L9eGPM+42p4zk/sAOk/NxYOYBa01sVpr+PZ6L4mOWJu08UgP3zYuDA/1sB
QSKh0CiiCDXdHGL6FhrTO51abDFg54bBG2yFfcIN3DUdrdOiNk2DTTUFAyv1sR/75mTgJrs+Fxou
aiBXVF2kePbInPpXzx0RvAQBXP+RGffbzltwZCKeFaO6JmLJUpLw+u0DLvniMoLqFirW9mT12OHz
7OFMwr9lKJe9w4AIOLjn3m0W30rn6sU8Us7905TEbv+P5w907dQjP81Z5oLwsxWcXHC99/6ilEt8
6LrP8vRpmTuYEAHhffGWkC671fBO9MzARnTJzkGVAnyMm9Dnh2NqOCO7ByFa4ZfFqEhVJgqgjj+7
xWfhjyPFkqsAtOs/dHoze/YpaOD5XMhbxZJYXITMLL6eSzNjvu4ynXxmAqx+UYtXhidg5Z5qO4Qa
vLAPKtxHMGJIg3ZRKqTZMEnj2D46kfpXa/OZHE+CNXZGeTOePvd7rjbfMTQNHkCfreY7T/P/qBus
sh3j/IfnGqyFJP83qUp8fqA1CStdvYk1Aft0w+XUpU4w4Bnz8N0bTH5UiivP70NQ+0Ln8UerFuV6
YnIfqI+V9lWiV/tagultX7b/5he1Txx70ktTENNHxzGu+ptcBO41khWZqdWB7ZKsvNWdfYqnF4sX
fM2fBLHF/QPdT9DDLB+nfZlp/Fj9VZq9GpT96xXCYY8/CmbbEUL6+PNevLMxuoMJYTl5RMP905uK
/JzxeTOE94Z2WtyAB3Bwf3bIjLlB/e+DwOy1UMvbiBNj+cj0r/mP4Kk802Rk4ev61bDCf7d3jEoh
DNeuvFNj7aFI7m8WobJbxB6st6/+bFVeKw3egLE5vIIi7IVk12SKOFAl/dRuPCmdzJmUIuWxWSY8
E+1JatDV7PeoHRx6UYAXQZ8SIC9aT608TXRONrbuuP6r0H9D5qoKx15xWvukzEKlBqXwWNWTiv9x
G1ILCJoRHl8A6HswMe1CfVsc3V2jMfMfjcCMOAvxvKRrbP2AOBJkpkX1y1Bv9rNWZfNRy+bVvN5h
W43g1LTpnqboUF5pad97eOviAtNdW7kxl/fI4jFkHhswjdH61L6dV0gqSJ1ANaiV9YkkHvVbTs23
aso8zIgLuM/vTvthGOU5hl+MkHsVyGdrbgUGO8FUx5OPB/hgM6UMZYHMc8gs7HKDlVFv+lLC8YrU
3KVDrcheI/uSF9bkrgMM4E/vL4LrCpnObiVvGBi/40PM+dUuMjv2YEO/3pwwpRJqZ9sgIGa0B0e0
Jf3/TtsV27LbPfzaubvme5Bq+Vg4cT+7xQrOVnhM4th6yqkk06iWM0ZsJ5FjiNTwLvVAfo0CMht5
+6kkGyjKGXZge1Wr9QBuN30ArGH4qvQ0Sg0ZvARrLpFMqTHLJxDTY/G1uccHJqBRxQk/usIdUHqr
TgK+vQusVTdn4+SBegiaWKnHnpZwQajCHSRKpJo67rW31xtMXNZjRKViLvJb0VoWGbzKBvELs8Tg
ViUCNtWFjaHSktuogEgD+Q1pZDb5ly1iKcNPVW2Nt90xY6uN46LqexchXSTtCgqMLnB4FST434ls
vhM9ps3tLxtt3JVDNGbRcDCkg9GSQK5axwKHv0JfafhS33ZFcm0ukV3QHipR53YpR5bcXhyvPgnu
tQ1QAEwN6TSMpaJJ7odcrt3WGcLU310zmi/z9ukKjPElSPuIH6CLuiaRmYuVSRp9HneO02uXcaXT
QVdWjfPO3m9CGdj037l6QrUEIadY+42pV9mQaNRURa8Hmcm4OfWaY5dCDqL1fyD6Iqr/QQqpvvM8
YGCmYrdpdTgiP2gCm3acdqEAMAvL6pM/LkFaEMV9Jqy5n0KXBtn9eE8vz8/XX1lfV6ZSyEHryqvs
itUIOYfNMYlLeutmiWosHH3M3ctB0kLzzpufFHNKAV0oxc+dtAAfqKX/R4Mjbjh+dbY8rvBDwNPQ
G+E9VI3PBQGxFEhx5ujq5jKjpX8BkIFrtmEU8HZGde7NdFbROdDfhAXZdmLL7+6neGJ/pTQliQ2y
yCQY/X9sLDB4zNHunhPFoZYgPdVeClm6iIYZ4mt9ncQzEpgEVMmaRgEfsI3dnD+12Za1Td0GRZYW
i2IKgNnPEugfCGkrK6i2mD+rDVeAI1CLqPXQVDh+ENu3nhulFD9kJYZ5BkxE06VjluGEUt7EqytG
NpRBOgdLwthDihJD+VMGSo79m3orS2drsOM2bpR1d6gaF7oS5WTAHk9x1SQElyS072sj5lHHSDqb
IhMYBxQdOQPjQKdgMmmCqSCKkXVxnCq1KRnB9heiU+2TFZZChFAXuj/7wypw+DnOKH0lXc3dErkv
zR/8vqcu41NK3RwLUzlMp82PTo0Mvt8vq7Y/34+w68uAFesoCsv95OpQC9JvrhHbMI3f1xbDgd4u
sgop/+K/fHqIs9HsW49sFWCIZ+P7n5ibmtTzDXEi66Rpuh1sPh38l76NEcyMiA0v8gtnW1Obkxy8
HTfWLffAs9th5zySF4nJoC9rMKn/OzMi2Gyz3rRM2Om6bXuiw097OHX55UUeCdt1KSOTf8viAQg3
vITzujKAEJdnVxN9ybqc9JhPXS4N9bpVSfQ2ou5rsxjuKC3303XTqGr0vA9JfokNNrSm+6dOVger
SOcPykjaaY4s6epXcqPgng0DUR2KBczSrDm6Wy5KXXiGyFzP3j2d68uAoqzufu5D/x4mSPEifRAi
nJH7jKhKeE3cyW4hNuElgqBWEbyWDd1rEjzagzptz1/ufjOQd/rx7BVmOsoyBgHgyr6Lo0hH656B
9/ZcUwLxhd+vUgSSccI4cJkZNqnhSfuDSH+PucfonUz68QTB/F7RRJQdWU4F4AB1j20JZcmK8ekk
ooxjbZ8LPddo33yjAsOognnjXOVjpSzYUIACcXuzhrozozr/SGBuOZLV5KawNP6NpKbhUwZZfny2
ucQ2hmjAXl+ZJOUD2+1Ko5irkN7TekAPPJRuyW2JKOasFyDQzsksZNuYWH5upEkOnvxAtdOm+paZ
LU/jzQACQASibwcLJOMde8zVZjBF0a5ABapitaE1ZRGysNdRsaXAfY83jWN/EUe5y/5AkT/gIoOw
Sjpyjvm0TVQZhX1LQtiDK6Cz3K527Z6obbXNvKDQ77Fg6BeihVpJ9qAFOllIJOb3LqFK6n7ZmheP
kmWUUx2MHongph/CNFLxBqhlumSJZ5lhPn2YneplJdYmAx+AhDn3wbiE5cnDuEKzK12aQXNmY+Pf
XlvLjYWk7kXzeBa0HGS+za3ycqdy4+vuf3lHeREopUpk/SbNt9AnVN/CJELLQH3+89v+uakOiqcO
5jlPQ14E+csE96zv6IdLHmMh4E6IuxGWE+9uRkYWJuwcCZrgYIydECYG20b7kMcBGdUX5h/7Tv0N
w5YFychbmXTEUuT073PEELfzQGlzxQ+o1Z/6m0GcS2EveSrlNVhzCXPj38AAakA4rgZhsrVKcjMN
fNGWKwWn4WhIsp59FlvQoMfM0uPhXAwMh8qHwI1ytxZnTGRXe7ji4ZU0qnCGtJKgkT/jTaGp+5+u
ktx+PLdDABUchH9Cz9vR3rZ3oJztLCJe4Goki7sUVDyNVioujgZbge4THdADHVAAL5KpqNeaZiku
OJOz5OLo6sqBr5Z8YFcKlrlgB2OVYIPUGwH8KxaZKHuN7t1LytOYruhh8EUXVEPEitZHO9WrrymW
W1o2VG0qamUxmUfRjRohEgQznADDNWttSWqVHdGyraHkUxrHVS46CX4XpNySzbRyxvhwcB+nWIHI
5ZPUKv8S0EZ6rJqjWhjGKpCcCkrWlQ2zL4v7XMrucND9eDiB1ofrOaXDvrx7+3uVWON3GYLUaBbs
xynFbMx1Pd98+3TsjhyvCIIbNb7GpEbKRTsnC/p8jAkxM01lJCpn4crOSCIarBX765m+UnOk0Ujx
ZPNK4JwDkT7VK0cD4efq9NJEzck/qgbw1L+zSG5tUYw8xYctidNVQn5LI4Yp3PxqEXKp8ZVedS9M
RJOpn2fcECKGKCCrZl5tzpfP+5iCNjiOQrLRVlmNGQdse01GrKX3+6zHhDaDVE68FWPlhtEd7cAd
f76/wpXHUejV1l38GUUtFlSaDrOIIUWpp8o3+6Qey+BW0Eq6YyOwQ39bCEKb7UMtoWfpNrWEIFeS
nPxX9zDEaVaMctStVktmSuvCgpl23cscm/m9kRrWJsNYISOMv10b9Kw4F1LYKIjJEEurbTakurb5
YmNDMbEx59oV16zwzVkR7GmR/dle31EV3mMbPax8ACdIy7yopaYmB06GCLZYymPdAMdvC55KE+9U
a0hYM6k/NBLSzdAldkB8OGHN0y3/Rf1A7CALKUmEkqhjTSK5LzWv7ivs+uGBKGiAeoWDfTT1Ecco
qR/DV6GuFM/nV5kRpXz63GWuGP5yQAmEbX9rRRKxILHf4rBRxnFeaBMaPnZkK/sdmOifTcOR7Pf1
wHTOKHCLga1TouH8tLXHerx8cQT5IwIEPnpuk+2PVJU90GyYhlhrJz1PgwotO9NTRAptoM+8u1kH
5Z0Wv4HAim2ttqLOVFOLCiXa8E1ULo6hwJVUzBgEDm+QTa8Lhqj4ZgUihtG+JA3va5fbUQr19OjW
ATO+xbwWI4AL5LnHLm1ZiMrS+TnJ0NXU5EeUBc5VzsOoKXl8WLnFY79o5QfSjZ+6Y8fEwinIzZ4T
6k1BQ0FdQpmvdUrZyFMJK0kxdpvD3chqONTgYLugQG+1UGkxyVw3JyAaS+7Q1P/uUePP3D7FKebb
GHzmZzlSJn1uGBIaDcXBmqoLaj6ZngvrXW4h/N+i9ZMwJF2dT9N8BtnLMXoHvxRBvwD52WYIEfyZ
5bDjEVn0IlMexAIiTzmJBv8AGZK6Wic00dHggws79Y+2tOhXScRr/LHUBsCxGnHkj/1dHTCTTWeR
GQ3kZJqDIfJs13/InlnRKpm4ZJxHAvheuny4eIXR0J3TGewy9Gr/6ZRGDgxma65PPX8gmMOfxdko
4fJr+m+e/Jj5RoKojR1V+qHPDo70ePRWh+sUd/ozhcF169w+B+dJXB/qtbBvl6fEOWzjBn4xkZLO
BkwgkMn8j5yYn2kB8att90lnyryWylc+Fy1BAgOZAC3WhtSigrjkYK5NLZOC1pUO2Be/cgMhb/np
QV5jc0H/rdmpLv9FTULBrbtg0Kzot1jnLTUdEjcBWJDuQRSJDVCFDsF7XzbkO4oi3zlE9ZnGetfR
70neVkvQO14tsOLbPjT95Kh65s/wuxmmH2ZU1OEFolmii1FpFUoWTGT8MLqt6kI1x+66boKi1aQf
y+M1EeJOTDLw1uQofbA4PHI2jdW6xiflK4b//xLHIGVYRHkzDijGFmjpTHD06qmrpQfcTQeI4R5x
PTtgaZiwM6Ay0cjhQGApM+UWYO3dRcZECJbKhqXKVQ2JprdSKPqOvFQ5gPHKB7WsyViatItUlhny
9kkfmMDvyS/OPUcQAhgMTv8VVAANJZJ7GHGI45UOeFYKrBWGYWakqKPdmx4oL5bo4v5zLN0WopQn
cFVssFlTVFMmLpO6PJp1a10HrOTcJCtFyCc29GmIVo9qIKY4oOysGktq3qsoFOAsL7yuEkAr0ing
VfjjBDJ06FkF8NPsbPsip6cWRurLL1/zRibS0QKfO8q1DQOhsM+RWVz0wqgSD+jaC6s33q7VT1Vx
HRBSEoGlW9Fy1C940OWCXkpSApnH6Ydp/8x6D4sgvW/Ye4ER8JSett1vmVviNSAVnBPdKQtqzosi
6h6k+NZ1QVy/AfqL5aA+qbxfZf2+wX9L0x5qDQ4DWQ9WDVO3okkB8liLy1Tz3Gr+5sAYFilFimCk
Uwz6COKa4o/FY1D4Mf2rU64+7IcMSRK+iCLc+P6doQB79/eivccoiQbL3HPLWw2zSiatsrkpdAtw
GXFWWBY12wvoETS5IDQjldZvHCX64gKiSzf95WVbJAraAotcHAvwh322oq2wDaHyPNZAkWYH8OrY
oDVEvdYpVc8V1sMu1kaBxGeKm0FfYztCjPD0Yfa2ZaopvqtlLzSVdXhb+I7t6eKUS4C2t2YJQqTn
1OEYf6vw3GcbC7Jt1Y1yeaHTHOP7cfF1B+gtBfomuXR4i4hN/01Oloq/DQM4FXoeR3z/SCcabLMr
MftsTkmcf+rajHN7LmTXnCSFZVVZOkF6TNW/fxNBtor11iCl206gxvz5Q2/HEs/bCRjMdrBeqh17
gNFLvuABiRXmxybMqOwcbAWdv9a+XCPb7wapbBEnvnxx0lqe84nJqAF8sqGObC7rGP/w94/zY+3B
CWSUk2WhE6lGY6i3bmdk30BsOm3sdklt6/q6SYN+BJvbI+b6L1PLE3d3A9L0NSbBM/yuhKGCq4EG
GO38amlB/NOlonJ6nUjjAee1uFIwl9ErezOBwxyOdQrbNGRjvI6IMVx3cN9hmHjk3YkHRLhKGkzZ
qyxa3fnrCBFirLtKTNJZr78l4gmjqOW71tcoxKgKmmMOwNXSYP0kNK4zdqwtXLogdy7xNxOdkXQU
mM/FxTxVSrW1B5ic08DLbmTFJmRp79C4Z4cC7KfuH1gEaku3igb+/LPgilNl95m3YcCtXLAoQACQ
Ka3L84a8LHNVJBPp0tTMnc7EeDrdgD+JKsJ29JZ6rRr4HSdBMyM9psfCKfI3DNwU62qrIVzrIvzy
zbWxcwDctCgeebdw/2Sy05/YZ11Z4oVfGQKKQe8PkF/LQD/K3pFnYImQDDB2/jZx5Cdc4Rj39+YB
XtElqTIrFUpNAQnD2jRkopgSvLbp6C1ozsg4DelI2LU9Sz5vfqgcvIETut73vs4WqNpv5fbtvbaN
lzBQYSvwXpr7PvcnIZMmuHo/DOAaCwahIlsdcZLcRRGIyWIThlvy2+2keB6toFgCjPyv8IYXwZm7
cQMo9todr9pNWORzk4j3O88Ta+f0bfYmsUJTuPAzk6ySwdB+LDLpHuson0hLoEmBrSfmQUaLG5K8
QKaQjN5NHnKBgYGZ51m3cdf9jmFxSGnzq2CPuKj/22QIuPNje6g7n7lj5nwy4S3ACEuVZe8i98OK
Fu1Cn+eOQM4LvnGt2TR/LzvtZgUVToUwOhUsj6LNAE/xxuZShpZ4L76mBOWmq9kodaCz2EEtzKkh
qmrP6nVieNKNHsU01LO+IUTHev2zfjsatNmXPGgxdG2Ice9hBGguebjXx4YU2f8HxE14YN5hXjqR
dV2+Fity6G/Doh3104XTgHgNYKVAW+wcHG7ppUT/P8SbynFD9VCnzvTIaDzYOkvWGOQl41JVTacC
1ldAslXuENNvQTz8xKjgNpMW1b6amXodxn1+Z+JGzA1PKGP8oq+QDrSY+lMG0htYwFoee2pTkPCV
MeCsT09OImL5KAuOmp8hfB8h2v4EGRbwztqqU9/NAx98dgIGWhAOhAgylCMKTOkpY+l+5kxc5Z6M
ALD3EQaFJAt2Rqjnka+jxzs0KtZreKrrTKWChmfiSgcrjIAP+MiHv7QedeiUY3ApY99fqyUB9Vii
Wx2kETDCTnsTmnSRQu91Y81DyQASKfzMeXsU61oCLakEJCGSHufgxQLiV7GzSoTWa2VuUBg0B+bP
w7sO//ZnkWXvLUDX5OZlvZGGYZumnmkp2EeWpudyeezB3HH+BfIzrlMyAn2P1A89zXI4rafeyzm4
APvl6ak+NRkjE8LOpnMuzeotTWs/7i9DrUIdIVgxv075MKAXX5jCx22msrIZmZen7BpyVmxN/k3F
1LSosSl/wuprgnBL7sqXer6DBcSQ2ARyWDWz3Nccvl8sdQXuIcq+hiXNodLyG2hJQNQl736ckLIM
gd/6mRg7JN6fFSLmsRI+vrmff3liDIEQzrHIUNpgJWbTV6ZXb2Tlhwtj04CsTkzO8UcYLCrYBcpy
em8t6qWt1eL7GoH2KlkyVVFUG3WY7Lc8g1+I3AB/lGZZFF4Md+rKZF719Ni45+RdDYXGfgO8TQs3
npYUR88pqqwPzXUK41bzWuHE4D+0yb7VsG+AKdbnp0ylMDK6rqUzZYxK4/s59k3lWEXESsiq7x6a
V6Uam/VbWuHOTUj8tQNLIj2zrHCvMXO5sz28t3ncwjj0Aer/cBjqHK75ztDX21fCFO6T8rIM3sWF
6MX2ovP/gHpZFfJOJ0fKCQOxbElTg48dceO8ldjhdUDJKtPOcjlxiMa7xPaHY0vrLpKSkr3NoSgU
AVKc7Uuop8CyAX0Z/bza9Bt5ecWiEdd+6R1djC85A1n8ajzrPH8e50wQ7lmj8u91OFuwgmdvY3xi
UcDZbYcBfv9waqqtGrfWnzRyDrlxMNFvkthMkA9ZebmD+63HnkzkFlWdSw08wHvtPWlj8CBKudPq
UN8mlbeptq6rHwlTOewismRP/dJWs00upeU1ebJpTuUt0uZYpyQn50KNEJuMucoIYa5OdOxVYr2X
fn5Wi1BaPg4cpPFPO8VrxHBWz7NgkPokHOGp0DUo+9xrjhE4GgMQS1n2A2P3bKo2I5YOqKrCKbxF
+YpktgZtVhNcyYrFoRkks7pEX/CN5CFA9RKKzKZmZF7WmvMZBEzdFEoQK6+wu/FGCD86pPt33pzF
x8lcfrFOQY9bgD4V0HSY/UokTr6yhUcIglhYPXWmyYvIZBK2gzG4Jk9st/4fus9wjqHwBFR8xhdc
aTRL4uxkZqEI0H/hi7MnJf+OdIOZ4Y/K6aZe2uCAPPVT/siEA4rZVKPZz7bMZiLW5TfLzirvwYc4
sCPGbycBYMQQni+ZDntGhhrP4ydsrx5wGZB5nsVCcfxnpal6GUYvAXK4GqMGjIiG0X5eIFG7NfDG
r8R2Gal9b/h8tyRFaYmZh7m57KISWrj/oMP3XQ4IYd79DRtoYJAWy6iyzlLS5NuXUCOc5lnit8mO
8UoP0eP7BHZh9LFUJVuWikSrsF313A9YJib3J/EkEakKdWZtENc5F5m/UXpRhbgADnBSLXgyd/pS
H2TDz3TV8oTOUFmPFKibYBwuAxxCJMriaP7cbJFx4JI826U2EySRwX+PukjU/BHAWHVBD1cXTlz3
YOuBO5zAK82rjppLAqWXtHtZF55DOspCQOSRKLhaCWAkP3Q84rrUL/xudBA+aPrTFr8vghubshy0
DDJgZvq6G40dfcbWj/8ECzOSJG3eu2NPpSqGdOS6Zg+VMTreEga51nUdZ/ME53wEIojOZ5i8soFM
BVwRBhkol85UigTm2ztXklgy/YW9K1aYmN4t1Z05HGpAvQOP96otXGSNhAkgGqSQkbLsBkcLX242
UacBQK3kB2R9n7WsCHxkoKK96VdMl1XRl+abUTeLPOOMp3q9TyUY3z1zdbHin9u5IhTMY8FnfwGE
EokJthbaQZfke2MXDqHiKjf3YFGNiLcTQ3n8rX+1Bb4l9ehnRKkF/svqqqDFZzx8QWqPgfH13BdF
N89wWHcNwQN7Uyb7H+c1pSDZbjzDW95a4r3ko+/BVqit5PvCiJEZUUIGBKKn+ndFajrgISftEgNN
RWVxnby5Cq48GSRtvUP1YPjPtMpGZSiAjI06bsWnF2u+zmFKC8GI88g/jADf/NRHZdDCTVUeqFIB
c3+yHmP6Bxd3F9q66M404p3/iIBhHtDbtQnyJSOKBkAMu8z5VFF2ezEH4GyqCVpYNnALI0hEWdlw
kbwaD0hVQ96HK3r/2/E5+DfushrFit/L0CtVmhGt3h8h1LX/DiAh5FZWX0rtcdxCnXGVHSr4Tglc
L5szY5cZvhSI/ZNkWNFdJztgkVDQD+3vI2HlAQp3ed4foWOJ7o+md8bzBC3caD2xCOel3pqMUNy2
Q2QDyGXxW7lrIUiTiJO1bw162pJfuGHWK59x993LNNwMYryaJtbsrkFqpLSEoRykD3GtqqD6C9c8
it2q05yVX4hNroZQ+qQjOmwwafNPLPNmNiVHeComU62Do703H0KAb3UI1QbEwktM/+iNv2qKCLmQ
bmVOzOVx8O5xs75ixwoEEagU74ihJnqyh5md5O1l3F6nULlQyNvMp0qMOskUXjxz78I3ysKWCICa
qRRfcNYM+Iq5Rn2ZK1fD4zxK4hWy9UPN4d2vEpg1ytIfVPKTOpWhx4+0B/5/AQLIiSlSD7R9N9sx
eWgLrSBsUmYZbivVDCje0YG8hlOa9+wexIrCqDBdAgllpBSf36EbMNXWwiD0gZPfEGKZZ4QkWFBY
07bh/DCZFBUJd8e/x7Ut4y60s2LutmPNiZzIoXWe7Sm78wPUsqB89fvD/l/bT088x0OBEDixtLF0
0kHNGs/58CuHotEUKpeYWTXX9ZOmawP6FPlqqC9AZluDTprB+ytGmQmtFJrlj2aeEn0HPC+AaIK6
avtj8P6T7pt42OCgpQdwSTkdxt32dB/GXuAv0RYco48uzEw3qARrIlSDyBzcNjGkQAsFbnhuNkqr
ICCM40I5a41yf0Ezt2wG+T6cCXOR9XnpF8yJsHqbTDnNXYIC1ZFIGp4bpyWP7fPByT7C/G5M3X8U
bjXxDfqWzDjq9FHaOGX3OvCnFJXOSOYDiGiQB7l4UCt/hNr7hxT42AzAjok3GbqnE5qJofM9WzWT
JXiDshsJZ+j/1V69vPC66oXP2JVcf++kyW90wOynsY3dwMSQ2z27Eqc5FohBNk5eVrh3CbgLRLJq
I788WelPdHtw3L5eMtZac74G+gpc+uzV2px1HYWH1Sr6BbTloR8L6UmTw1J5jL5RQWuHuGTPJMHN
J2q+dnY/XfIu5wXfyQU1uk/mAzbwThllCFg6o3UvjpdwTfwpO2bThZGfkozu+hkMc0qpyvdswhl/
wA+LGcZEmDCYnIg8xeSmWz+h/h3P5I09bbmf3ZKPogThXj/+ELV0EeTGApPiIzM/c2Vrn4PSfT3F
uf8iSMlBHz7kL71YhIDBHLcr2ZpnSa3KJEBQq9jG24ebt48qkSacdcjHF242hOKHE0npene4mRNv
Y7iKTjISzXfnS8nPyZ8uZEqwoXUdG5mV3MfK089BhkSI5/uaHL1wDOJ9F2NNuJseUH9tzLw6BJpb
Co9dT/argMQwDF3N3kFmupGVIfp9G9xdU/JBzRfvsr9LAxH36BinG8xEDYl6S5tN0/necGP0tmkt
rOAH7D50wA0fijpyCYgM+OHQoeDdu3xgPjubRnPlIXLb2SdNbkrr6qMbXZuPGj/9I8HsIBaD4ksI
hqwHQHTUQ3b5k5yFeZ/6GQ0IiDb6Q3Kzxp7rR2qFlgbyBCIsl/Px3NpSqXkmMGid9gFVA1yywQqU
Bq1cEgyq078pP6qz8uzozPfCAA80NztOOKvYq5nyj/LbWPXo/hh3on9yDHfK6C4xnIX8QS5qshbP
ff3VRkUHT9oV3Q/fCHUFLbmbIXZt8O4SjOqSu1WMHnV7szJkyUQa53AXJL3G5nX6VvpEPgDoZWIa
3DaNTTFjdwPAdBap5FnYkaGuwdjimB2McPktlxY8zCT0TGFIjcOgr/jksVHLpox+ZWPa6RFuuSpY
YA1wRkEaI05495H5DqGGbyR4YoGe57M8rBdyXik+TL6nKADSPMo+bhFVCOP4YdK6wJKaHdq1d4pq
WbLSSv5CQ6Vl8v+UU5wo/QD4uQ9ZDaZUrI4//hN2KnX8klstnqk3n4VQNSTq058LEndWN9FTJHtb
OBK+2B1Vim+G8Op5lMl0O+Y4QIcwoRp9NNSNdakSIGCCxCAPx2PvP4l0xOhorDCnP8/vInM0wLm0
KCOyM+P12e2vcSuKmNXKWv3+30ZT44ghw4AoWpd2PXwRt8Bacyc7UU6k+l+bmvFyeXAM9TN4X2W6
sFtt2ptbHMfplzgMzCON3zaKAI8fl8Hlx+HkeY8W1wbzQ3/uSN2nbCY8EKRbC+X3+KU1QzDOu+oG
CGCkCaE1mErJFXNPUwa6dZystr/HKuP/bUItzHJ5BHLOBq8VA0XamQAFEH26yMRJPHZ1jAXILIar
X9/R1XWnVaI5hXVuhzGiG3JsNonK2Mhp5ExgORUx/qLQ7LM3murF48d7Tx6j+1PnneHwvPWBpcIJ
qsoQtosQ5HIuSLxy6LDiw5h/xcs0TpO78vousMisfrUga/LAoqFTZ1DSZOHAyVTADJ0m2K7Eg5hg
oqKMFAfs41X3OSYlMf/asq2XM/7vfs2q7ey9+HsgOjkcX9axlIBsxnlF8TM8cF2GQZhJJAqN+aEK
Uzj7kP1X2ptkj9rWufO7NCBDWWd7qfg6oYCxMmykGOlmBXvDUeSLtuuz7ZZGyteNuI0O72uIQtPY
cTOXy4uCjmiwYCfBonSeIKMKZCSilQc/KfscjNxl2vy4MCpNkYXyiC/JMx5vHYzuTHF0GOlZaZGr
LrpSLS+oUwvhMmqCvRLoPQptFyrS9hixa1aPh8Xc5ss1e2D/iM5CZfkYALmXgvkQleHYvcg2uXha
fc2EGm8PtNyPaXoTLq39HFSwr4St0pn+xblKEyUQhEdaHQuneZLtv6hEyx2Yiv+fgacfZdJeqMg3
9spif4U07nhrkGCm/lxzcjvgsOjyC7hR9fcOWWXdPKoqQmMdQ0eNPra2JxhJgFOs70m1Hsgk6dO5
vlzTExREOrPuxuT823OIlXFAZcs8cHVtxFw3FR5yhxacgDtsI4HuwNLQGNiUaNlN7P1Y1DSIqyd0
6vUR44V2DvY7E04foVcYcI3WhGto0IuSZyyBy9ZQoes6xlHU+4VmCL/1LBSFwQoqAkpUa5o1JqcC
2bIDjZwJ/nMmJfw555u7uY/drjPeMMXRg7m2TW/B75MtRCJiqGZ4RsDs6pT5fqNM3qsKS+k5xAzf
LKPH/d1yvElz7bzXxgKRFGHttBPq/3gHUERR3GnEwZpd2Za3PDKULnRF1JQZ7io0PrRdhyHD8vq3
5K0ny9rzZ4RLC7EbWzF1X55pI4osS5BQUvNFS8GxB+1TCW8DsiBJQ6xev0r4rvhTxFuF+m5D+Xs9
w2/XoNT8Q/qmB/kH4/ULjMGskNPiGuRu1R5Z7ZR+RDk+tDOBBZkFMkDphHHGbMkGgm4QipA58ky8
j26vwiz2jrp5D26746DR1k6/Q3gEgyVOVRPlvggB9orbsTbgM9Z65QMU4eX56IDHScApksw0ez7q
p6zBeOeM5ZQVcMCtLtw838DzXHoAJdeP4qpKhnr9BplPfyNOJDmlhoUaNV82MsVwg1+78BNN0nWn
H5rU5XZcNJOfQcyUjQUePlGQnE46i9SgIWCIIOeeMSuJrY9WUvXjZJ64ocyI/8WSwEIodKInilwU
WJaqWZDmVXx0t/Y39/zPn97+pV8p/6faKKtZrjPqr3PdcB7dcGNz7cjpIyhH9QGnyaIL/fcB1cww
/mmK23I2wK3raEZmOleaNaQwOXKjrgNLsDShGQjt7+DSdRJC4ay5P0DAKnoirw86OKenAwQrbcgX
eLuHoG0KUlmE60cPtSkl9c0SEtmiSogml/um8C3PT/0kbR8mdWXNCg9Dkd8+nIyl4ld1yN/b7I6K
9lI/aOBtKy6T40DNoUnBIZhBlr3oBvNGTqWqxnLo0o46qnaNLf1bNPlpMxryNoOashokwz82N01R
lTucG7UTfZ/AhYMfmpouKUNvr/0uOA7YmTtIsHEsCYr9kLE6qjEZSPE/Qsp2UjvQShuSDLzVxVUt
DRCL641CAHhbqKfbwb7KelbDczUqgpS1aMHoj75CJ8IPy6vE7+c0Vw3oy5hopLzccOH/9PSNKdxB
sim7UB0/PxkBp+UWeYovzNPA1wDsgoUMiF9tnENWIkd1gRRwWCnFTnZ9w22P5S9AaK/6py/F4yk+
B8E/FMQHJqT4FHTJDDbAMBdlBpwJa3S3saljfZqfTZKWSYCbQilPwN089HjuSv6Hvajl5HmJfymm
oqOh9xgDVcy4MEUT1LmVDRP1b8EZYNwbTONvCbC2oDKV11GDr++9kdBsNNzzqFn3HbN5RuKP5Uyu
jHBzBxZ3NAIMoxNbP32nrxc3XB1XsfH1n/kVDK4fM/L4ThnJPrqfTWY1CowGhsLhib8zzE8qq547
HRp5qkQMhsoEooA1xjCdwKBiHBZlqihwCpDicEmLM4JZrPcJn7GjjGw0/mSDJdJ5NpNZOcyu0i3K
KCPdz+Q81NrrkuervBTOks60f25h/WImM9lc2Ek3RsiABdaBUVC+r8zvfjAV1eaDm30U92XVioAz
Dlr/NAylMNnBF33wrb+m+IztzJ/S40bXch6to937IHhDi/davOrO5jpfIArdbGrrgHSEVvB2i0wS
R5WTqvS0pks0SVbqkdKb0faUFTaA5k+VSSxGHYdCjMpokfPcsq8FLMd5R9wUT9DizZbAI8shT43q
pm3AUoFewvTzo1WsZyRaMESttgZR40lu0joBfzwtchIBsApscBKKl3eksFYUDTscld05mOrgRKVF
od+cryZvYnhXw4uaT43grqKdNlTR0tCfYQmOMzeGKNSkPH2X8O5hDS/TvNSAX3vFi6s21DG/kwMj
GexwESPqHJegPd2DQekjQdP4dJUmci+SWWt188kebNj10JZyhyXx043Rn0CfJk/aljoOWcNeOdHB
aIq4TBk767GldoJIz7Jq42Rq4T7CqpE+y44GKT7DKfl9qNrtd3qv2qikJzUWgFGc4H1J+ukbFbg4
KeMwKEBPhPwlU5B2OUgqmBVsvQ0p7ZEwiVmGxBaWy4W5sLRWsXqCoY+gw17JPDfrlk8l/bANv/lk
fMtUIZLWwo5+bYIKTYDWkwl5WC/JHvnhuJlOXbqwb5LmvTtVh6pYDaAn/HuBdnSC8ouUSJr3JfsT
KS/GOiAEWMZNHblFic1IR3fdGH2NmV7wAPfufZQRmAcW4ZuY6kE76MZYSPTRqSON8iNiJALbkv1t
kbPX+e26NiPv5qidjxjwRW4xrkFj1BIA/+/MBxXwioRmJ1baSsmI7wTM2J6BehCIH6mWPzuVgorE
XDDuiUiBvMYLXp88/by31rNph1CXmVZWb4/stJD9Ts9URs8Abz9m5e75vtQDwLaxNDUY66K9GTSr
WRzsR1Evwd1uMbQ5Q9jkUwoBR/APLoEh8Hm5Nvi0i6YLcRyjKaIdGNBu4S8VKalafeC5xZUKFH/2
R0n9NKiRI3DeCMn9uBUGfMnK26E5b/uIIevwU4BAVx0e9GT52d4+3oGDcGHd5dhIqDejD9wI8pmQ
VdGbqoDS71w0ZtHfFwHvwSURo5L0As3dH7o30ef2JHWykEUZaroj0HF3xRRVMYu7WyraxQpN7+ND
2h+FiiH+811uLlP96qpjkUdz/tR26e0KrDuXE3vScTX9ukoav/M8TSc2l84Eed1aRZMklwOlq2x4
q4arcjjAz1/nmJSEkxrQhLs98R3KNb/8NiSt3yHNBBEs8bCvXWDHFLlqYq9ChLCSfmdW3z4Lm+Qh
i10L/tuRdzBo/WRj5LqSkFMWd3kxim233NChkDCPMS+zbaoUKzXlB0JrtEggMUPO/1NrXX4yQCsk
0cBiebUnCxMwYh7008+ELRyEUt95SfLVfIyAcPVQUaK8zwEyBS/jbXgjCIE+oP2YsESBM2Q9fVZH
XQBQJo0WShS+FNKyvxkZeVdWUVDF3Qn2kaQMPJ8luMkPqjgxUfVA01uWNqaX16wTCedf/KU/veKw
9W4GA/zJ9NXzIETg4tigEUm5uZCrwdruCoSIh0Z8TGYht5s66Lt3RE9qTfLXEmPHjZv1Kp7eb3NX
fZj2s5JbGr6P00JNPPKHOShRpsZiujHNGqF+deP/J19bsa4YDhm8hr3TSbPoX+QI1U6tAE+eKImI
VAyZlBSlnSjdJmdiR5S8c4L+1HnQymYWs4Kmn40i3OEkc6h+Yph97c6AneE3T5ZIb/7oXICz8W9L
xdTZzMalRnej7j7AeuPIkozKL0JiDVuxtg/g0w623yHiOTvPo7A6WTy7R6RvUNlPa7EbbZzFhVDR
0g9p8PStm6Fp0/8ZJ6EbAyv32vulvY5VfNe1ApZAdXeChpbWYCwKheJhM5fg+wZMLVsfc/pQOiY+
Jp6hkQ1cUo2YBVFXmyAUmhcM/dQdt5OSKuurWDybZmvPafUnd78J4rCNRgwBxPnYneYFj8fHiIfw
en9/nAx/TZWrraG0GMEwNkCCNzptPW5h9neVQQYyQYntGQ9IvaFT+8fBDsF3dcsvLzWAMymETvN1
G/txczV0r/FjiVVWbAfcW7yOCz/TTd/vE/ilySuUL8xypqNuZ2qlmFcWYZzxb6x8pLZOCJWHLV1+
vSudF3IFljGKHuM7dxCvPCVI0vf01n2qTiynCWFBIbsjfb1CvhuJGoms/JthEwDxfxCV8b8Ap1ju
oNgLPC1F94u8OChUxAmoZo/7ezZLMn+aRExYJ7zhwnL9w2Z3TOw+wyJbBokhATbFZxXSF7TwBnAO
2xA5n1kcaLmziRg246mWY7ZkSL++J7UFYZM8yQi4EswiDeNfAy6dvVi8p4i1GZu4u9Yzxg39jIuI
fPz5M9wJqD6WkUlYWBe0Auq/uJ0/eWHHBLL/Lt5zupR4RY+GaaFFGKrlaSbhfPmyEppi6QJuOapV
4xNn1TYqdo5pL75MJ5JAeifBYYLlVeerKnKh6sWgyFvitm1QefmY/rdy3kXsPrs83XWX5TpfE6Nn
QABydA2QrwB4AfJEur2bq8pMRBlvo1i8ZQrw8ZK3sQiqwgmLRQCK3HlL97RK5h9OUbJi8Zss0H6b
eyN9OpEl4k8aHGmzkjoXbN0Bu63eoqxt5yKoNjXy/PbAdKveNGM9In6LdZC3qCl/g20+ezGd3nHn
Nl3UBeTfNbOf20gPFxy6qYnnqmAAYV6ZF0K76MJCmh6TTmxSwWtCewYqqGqaOyhAPGeTOaK984aM
ummNAT0mbJAKaQieHsdKK1mD669MYSaI4N9+GPC68bwOOm+Iw3dIKnW3SDaikufO7Lf6cdJK4/ua
1zbAGAUUzhv9qip2LAXHOMJzNgz+0ZJCAr2k7WINqSzA7/9p+hBdR2lUCma1RUaU+fMykHY/eNbj
f+ygUqR0YyaY7k8H57p6iOZ+Mxr4jxfN2CWQclKijU6SQHqHhNqx9aK0t6FZs4GnREROZpJzmiaj
JG7GGthqN7OxwqWkp8gGvdZpOrRl+S9XeyFtGuLN8d6d94V/kCjVCgZkP+Mv5h5VRkluxNFdczOO
Erz0ekqkzkfJTSnDsFSeXL4m+d0Anp1jqCFEisCtFGJsSkSfXOhl4mVYgFWAFIIeB1cjGbJ5gmtG
OzvTgOAoI8h04nxpeGMlcKy20bg/73LRrZRknkNpRZuTYSn5M6u0vfnG0GPFZiDiSw2wlk4H3xQD
sBPEGgO++Geh9ixiJMZGCKZ2bWpaaF9DZjO2cMuT0K2rRKHiJUx+JJ1tsuve6KIKnubk9vSStyoS
NRo0O7zrargK0RKJF4IodOLvwhsboAy0xk0KAGZXjmXgCz9j5UQoKWhBa772C13mbQjUB07ee/5C
4W/iMZYLvsy255D5xm2KzfSRYlGDZEwSEJLpT26PpzGLC9yryVlOwZYf2oYkSLEYu+gn0Ge9iaEE
TE94WxJI73yDGio99fO+Jh91JwZrZyQgM76CeNctYQj64P08I1XwXE9oLPRP10Ihv5ZIgIaWYU7o
gGL8RsBbDhJrmPgJK7JAiwObtzFnvBoFnm9mzLttPnaVEkZQDXhko+0tKZF0uTyq3KlhH5LveN0r
jLWX9tegVAmnh003sfXeKiR5qap9LRC8F1NlVTL467VI6+C0p4M1xtrVlKloqIfRFTYGNuq4a8NS
D5leywXQNYsW3ptpOSEcEO476YCsBAI6l9qa8M44jln+w9BInL0BewtjsNnH+Y2IPeRVNAqP5OYL
4h44XBB0CBWNOkL78knDHFdTB/pVgnPKxPYCCGMrWyDUYwZyzI7huc4PgHhOlIoKFlbhnH9eKqh6
x2Ap4je+4rk2/Wf794PAJAZCncaOR1IoRLZxnA3ed673g5W6D+Ey5fvonZD9ZbaIl/reCsSZPhX6
ZqZ1G9M8iH94IYNBZ2RZ/6fuzrkUhZ/PSG75VrAtnBTtcIvKkbb4yeyieJad768eU+FWjhcVl7z5
7zWZvWW9LH615zG+kHJkcFZ8/XmkUNAHHYnv/49+MgsfAZDR5ckKi8655GzDrrxOyNVwyUBkPhGm
1PMvbdr3N5yplKaxAFyt1thdkbReuA1c5EwJOOmiQFTs4qPI9lsysFbCazBMMhOCGYSyQ38XMX4E
EP9nDBsQGeUcGZtNVXOOA1pyXpWaWP8/ddpgUlpwb0ULl/FAINytI4LY/Hz32GNmcYPB2Aap+COq
jU6B3gt/7Sc1PaRdnHBSiinUlNkSlQWL9i6o+y8YGcloP8wLRsjPftoa6qCDnyUdnzJvhpcct18C
RmsMmtRMPImjvsqA9WaQmCxuzxm4JuJzSwiY/B3O4CzHs4OyM5obRKE2tvOvCaAEN2dvtqdAHI7d
sogDjPV4sRYkwa9r4pGyR3w0fuKql8rEEmo/qmI4NjmYxYQdezffk+2M6RIjAHG+4NVpuzyNopWM
k7j8V28sEOkMQFaMC6aL9jq3ygH730v9ZmxpvJ0kniMZ76Ec210vtSzZ3BuOImhn+Qmlyz3t60FQ
ei147Z1iGXSPVL2Ue+2HKE5cKOkqC1ifFI8VwYujSAk8Hod3V5Rwu2Ex0CYE6oaoiilvSqqdA29o
pWRYB46k54thVTioQpCQmzySwEigZoVk7VBgSYE9EOrSPRvaB5xL+mXv6uIzHZP1yUnK+qpzejyc
paMBcOumVHXEpRXitA8Gu52UnMeaK0qEtsOIvDzKBDzG5CXulqqXchSSlyBMMvOhtAB2ecTkLiEK
ux0AA47+8RRxOJ1+mpP+xR9RRPpdE/qVY4V1jXO3xpL0amXoSnctmxplQttD0Dpw7w+KM7jfCaMc
Z8qFQvuR9xEAwiFUADLC0fBGHUbcT1EOc1yft6fkemIh+ayCiYAgiGmxHsA0T9Q+YELXaU5fiGoC
8mFqr4ajtD5U6MSZMTuPkihKm6AnW/gSqivF5Wj4Nbz5FnoavqIklhMMHzP4DQQyddeAvUhnEHYs
aMyIR+pj6tXzWJQi4nWh6NGljDczyghDpM/Z/u7QmNWsFRnDYhbL2CSf2XkajYED32ETOVSIujvP
PzFPCYIaigrtnPv9lUJ1jYD16pD8JA5vV49+izcAbFLYJus2ZOPI8LsauwOUpgnJ3aYqqrXV4Xd9
lHQQe91oQigS6s4v6sc/ejLzPwJNGsmT35rxgwgIDufD5NrkK4k8P4L0ezvM1nG4U+i5gI3jnskm
DEXhSbvahDHlEqsVLODxqGbXRTk1dXD6FQj/iR46T1Y7Bu3SqsTIdOvP3WdBTYPxvYLXQ0jxJR7Y
PflLGmvWBLa7EOtZanZ2imv8PgeixfwHiS0AoYMWqWfFe57QFFafvmAlvu7SolxnEpvbr59pjA6b
7/Q2Ur00RoSrj5UPG5XoTjsikpXE8y31hORXOCRyPO0EhWm18TFEWwFpbKdWDRVamFCJVbEPM8Ao
3AGV29B5OriaNo75PxuqAL/mF5XMpWf+FO9UpHSeUQqDmsaSZkDBaAomIVNaOrqhgInWEfEy6kba
mqvFpbetSjRLaaGpQbI0QNaL6OphAWFcr8hoMG6P0+m/Gqh9CoF6kTTa9gJ34HV494g6H8PhrUOI
C7INYcHbqMoiFzt5krxb8Atx/9xLbP5eNeQz+h5YuSIdrsuoVNvthfrjlJRRKsmKGayuozeCmb7X
nvOVZ9xv/B8rnmEXpr+gazFCAqG2ZJR7xI0ce/C5bD+nUPjXdipVyB3BQlWsCS1Gbk11oLFEPpVg
nIF9bBM0HNsw62W0YVY5vMEam++6dwk8eGuhD1SEHhG/cl+s0eEzQivSaAAdvXvzHTFyXjUl/XR2
oZVvJLNpOgPBuuSDzvCQjmCRT5CUrYhv/u+krzd/OQAjT/eFE+9xUe2F3X12oXJD6Csd6rya7NTv
lz9PVa2vyCMF05uY/sB3ZM5XLwN9zb71w0XDyY75n6YYLalafE5MjSHUa8pOCkZPvqIhm0KnSVF3
bryOdDjNZpefy72MnYX+tVi3GCYyJhE4aROpCLIe7gsqisPypuenORmilIVhquemldNWDZDOph0o
DkS8SQlezjG3o7fkmC7okA3vWukDjIO0JIH06oe4U/A3ZKMmQcXWYgVJ9DeOeZHVnufoOsSvyNT/
wC3O8O0pCcbjsMDc53F1vAZ8rLsQkeWJWqaCl12vfAwhJXBhDGHA8V8r8vYHFhxhcJcLRIY8tGwO
EjjaKvGzvtWq0tIn0dBGhFP0rvafV5l7+tjuF9VE7XhmgyRWENAQAncNkyFYgDmLS5ilO2z58+NV
ajz4iQBEFHqbU/UJYNohi4iySRW9PVB+9xbkvDYXDMvViGkkkTOHRt/eZhceULpApCiQLAzeLR5b
qmcw4iMM93RNBnEnq7DVn7kdhvnSVuyD7Jyd9s7NCnM/79VqqKeL3GORKHzppkEUnLeq1b2gZKaH
GrfB4ezxLxUJpHM199VkOqjxq5sRB0Nlogcz92X1aioASs082DQmSXLiMoVQRDVLAxX9MTTK2GQJ
fk+XdgLxESfjVK9Zu4RfbBNcgsyxgIwrpdgj/Aifzemg2DDYVNTZ3B/k3uk8u1W4AILKxA9Nj+Yi
Can4McrBdbtJmEmD0y/UTh5bEfhwnvZl/T4Sk4liTqJEDVMbO+mCVx9YTwqEtYct/KI7Mtricu2K
xCfwuIhmW+zwuAhQRkfJZeXgKRBnDLtzm9VpdfKtXx8Fjta07jyc3ALxRSBoBUMrS+E7V0TYMhF/
+yPZOoeBsGPQCqL9zn886g95PzZPXCUj8uvf8ehxg0s4jp/W8utBwVyDHBWDRTn1EWbbk7vM9+Bo
FKvpRgvlDrsWNgrgY9maCHfJtKkPWcM1Ab96hiu3pA73ylj0P7otYkeU43J/aedKpDbu1IYJNxwR
QQsDJ9hsLgQB8r12NLAq6eu6q4oyryrLnwtiqdEOVFSJovwgfYfvdchxQXXkOs/n3vKI9IggwtmI
Da+HAF4hSKv7CCOl8/ilepB2IZGVXp7i12v3earmncXkmv0xvr+UyQ7QbJrZvkbWGnhGi/1gannh
AzxSJlWK6aWFCxVlBnBEBLzz51JUFt4MtBjdwGitCWz2MW6S/zeh//R8saEcAeXY8pG5eXWT7xTY
tiFT3xyJYUxfV4ADS+m3P6cARpSnJmPA6Rk65X/2qRGIl1/a66TjBNrC+Pfq7YC+tkPlHAFxBbV+
IE5RIo6//YCX+Aa0yQChfwbHG0VbaqvOyAaOdckUavWGmV2PHO3+ccwnO2i8sib8FEFwxdsj15cV
z8Gt5bYnKNlI+UoWtWRqVtC4Lf9Iz+5X+kGGDzOiFK1ko00bFNbDg31RfLbYS/SbWnKRXdV1Fkv7
95vAjzkZXAYZ/+E2/fyftjTYZtBARd9o50IIy4rk23JPgChCQnG1w4rVC0mqjLnCMXa2TL9YM8sR
rrgYYNH+9kJqjJcrAQeAd6NHp7LRhdaNskgqDdi/jbnpYS0rfQ466PMkBiG2N/wDeEfG2SMkiP1y
pcy2EWWjSiOpAJou8t9LFTjGXJFA3fM3KLduxVW1+o+eI0mcpImELMRoVJXkX6mU1DUNC09fAn4w
tIBNAQ8H3X9UufAyXzNCXbgo6e/SQfs7B0kPFy0vW9QXhvSIJkuOuXu3bj9aVSksvQ2BoDFOXhlY
pIHS8S54zHCY1q5hL3zaUoSW8UxWnLPszmn4vwrAX7xe62Bv/RJnpjs5YIx3YVdKaZlxWTLIMRlw
8h+7sK9US34ejxvqLtwpivl1N4grBMEz98BcxpJf89Nm0KvW3W6tzoqkDTbjfd8Zv9Z7zXyOAa+L
n75LnhCzDyXRvnmj4R9U/SkiseSpriMaABZIqMzbQ/xEC0j68pN1s37V1IZCqPoKe1WQ/hYBf+9/
/R60/WypPgXxaErce+NbRG/n86G4ZQKQYlRzDFBIELU9doznrXw3o7uscTXC/cz1bPJamNU7otO7
EFlFgY9jrkJRfPr/NEZCIWDRa77Ot4ZqRDCP4bEHU58CjPt8dzk4K3vJuUPiw7vEiowvjSKGudlq
9h3Q32V8T+T1W1ZaKhOeKGnx2YVUSCScoXQez2WFc/ov+Z7tp3JxWK+XJGWUxMBDlnQ3T9elQ36Z
jYt/gxo764Ong4YKGkF7PBxMbhrAG+cre3ee7+qw8XNYHpgyJz3oG+ZzhqUFg/k/uT4+eXUJUKHH
2cqVtf0oroT9mxe9n9jw1dpAeJGkwKhiFSwnRhRzPOeVx9LNQJVZrTBlImWCHGaoYVO6DHEyTUCs
GRrCv9KLpQ2kp0Nq379N3otyiYh6K/2h4i8ahgQUJ8yZ4TTgvwtFmVXqqNBXpyhxXhKr2NkuEpY3
s9AhrWshOHs7IOpoGExhOup9fL05tSB6LV1JLJ6UN718LFB8yVhufjHbH1OaALvFEcx1IbIawHen
a50m/ZyYwQXhBHB8pcsmYTvJlvGnGYIM6AywO+eJJDu5ze76gJ2EQAIiGrWteMZOgaAc1DR1OtUS
rQd2iB1KZ4qx2dSh2dq+7YREImkEKevVu+thiZsoxtBcDa0X5+9Oh6z9dsfP6rH7OGWNSZScsxIQ
qXOhV2RA29MJP9GJKmGaB6gZxcnVaJrv6MjOzB3/A+pMqYV0FkcLL6abriqnth0yTPru1jzRwvZv
9F6l7Mg5618B96+7EstCDh1v1C4sot2Uf39TVrnPDAPvwcQh5hIZJhDZvqiktVEhqc/IOI2vV8Zi
a1X3xEbtlTw0dUGOOezid9GhhLwjxqrMBA0gbaw3Z0kbZXHuRleLoxjpCCaADvvfia6FwseoUKMZ
rr9PPm5Y6QKnjLrYJCFP+syPOwWhCxDlDgo/VA4TMPvWkPH3/og05lkUxZVz48D59s3hn0TAlfCJ
c01j7sjWzbhM2FYejTfx6BvhGAH7PSP5q46NyDzbhldBPqRO129dvYZZdb+lVYaVwrj3TpFBF0XY
MNlqsZ8SPaW5vCDOxhwH/zl9+KmGhH2AGqCZlyykRYsrbL8lhL0cS0FZfjjeIf5WENikHk6e9ks+
NuU82vkJfKLyqaztYg6/fpCZ+SAPAYYC/W50JhY6g63Q8RqX6FaWB8COUxBFVpY6B9274D3IUB6h
p/i2GkAaUH6gt2R1SND5bvBMnrU5fzaMZwwqfGopRF+XKWd+wsgv7Dj6ufTXPqEm/LqmRovSLvA7
dPVMZI4hF6wW0zAISgMQM/RKW7iPqYV7EEZTfgw08j81r5ejWSdEMtwRawPkIlI3fvpC1P+Dx1Ya
XktdnnfnlwpXdFdlcYebdgsmczsspYJsoNSWTfo9b94vPIP383NGOiyEhCbEkD7JwegD6fM1ZHRt
iZPi5mUq6UYD0sL64m1655TbKW6A6iX4ws/DQ4TY0yZq9JpfdFCfqU43C6YC9JoJwshYP4Pzcfr8
sOKuuoqPKDnuG3e0N/c7w4bw1xajPULZ6/ZEf6xIHAD6aKVPBQUstyBiMnOpShw66ZBeRnj2TYhU
3R96cN3f239rI188oOmvKE+yE4SKTdCI6MPkwQRSOQRQ3M8GxnKMT4bmMso+LByHrOF5NxkWeeB/
2IMD2PwCCTgEqVDZDpDCUD9QBX+lCT9WBMF2DXOc/U2obrwhAfirofVuBWQNFTOc3iTnIbwVch0j
oGl9opkwDBcEG95tz0/qWT/Kv2B7vbES8DqSmPzSqABA2w7swLGB9cZu33TkZws3omhu1hiqB5m8
EY+SWpxh/7Tlw7RGcPX1kPgJeQ+EVgFHr56S0v1na8WXXGMAMXutHp3jDOxkOp0z0dkvWgBAx+kr
No9RxGA+JnUKH8760xC88Pf2aWq1C1BQqJlmx/JHQUWRinTJnm8n1SYptCN/0/D7c5svP47bY2tx
DQFTzLlJZ1TBLF2W2w6wv3OGsw6EFeiE+XObaPp1WuQblpyq/xWQjz90mUSop62r1UfXPXnYSkp9
CfN01syAp71tvdMKWcQNYUxE4dnpcmrSdnqVgqpAZnPmKQSj0lRrdQSeMlcW1mQVz2wrXGmfuWjN
Pvv4OuVJG+ztFP7EoNb5+byxV7hFFK3kAfEFHFrEkCAxJZPTyUUXfMrKyQXsrTSwbI32thPJ2rXc
HWQCeGoCJDB4904ol0txVJ5zYXC2ISFn7bf8aXeGHSD8mbc0/5GrSUqyg5Zo4/c6i9iu5o5mN8q5
dKVbv2J/L1HSgnUD6Tmz7vyby/+WL5AbhSvUMN2vUImHcYCkzlTCFOBprqiitt8+Ozr7eNdHc0g+
rdf2lPVDDnqgiFmgd71R4LUvhDOWHmsdtt3jkV2fJlbpvg3j/TxN7jmlVyNkwBY8OTF16/O9o3EJ
GCFVaRaq69B+QudqsZMx58fau5FoJBSDniNnS92Mch3tOuFY9cr3yJQxGxdsTvbp94q62MAd9yMz
qkCtHfpVwYw7oDvQrp+34aUq/1iEclJ2cY2YVx63eo7NMUPvnyZY28vBW8cNCYPoLAdNNReuwLJW
V0Ck2/CLvwEfBajdd+VQ+72JNDKJ+M7f2eac4cfuIX6Qfc9YDeofOxLCZMPjZh+2VSGZpSE/8OpG
luSU5CSMVR5e08FH8ypY1FY/MNvNwn/r4q6FrSjjWTx82IWvWtjpgy0XvsB+XbH/M951YAekM9Ud
/sN557o+3rB9/R26sZk81h+6JUGXvqnbjJBCpoIbiB30DykV+IjlJ+MJ2RfFDM9u/TR7PhPfpel1
tasnhuVit5VBO8HZImdQDgjytEGGd1Tjffu5WwS02Pv3BKuGtp/GCBY42gRN7Yz/YF5Oqt1wddrL
rR4z3kaeBR9Ke813Lh9hg7qQ5OdXdadERDs68E14eNB+cLwGD4P9QgVVtUHWxg4njKxqQ8KqVWtR
rSFc8s5R5shuQKWxt8jQPT0EMp1xrnbM0EPiaHvl8BHsalc1RwriWnKYRrlzbr7Q7CWsRZQ4kgdu
/cBMKvWiXYxXt/pFR3xBN+cGcXfdJUj/ThMx1FeII4aYzSdI+1TzIAfTRNYICjXcPDFRVwAp4YHD
QSm9HpHNthyMSneLJem+HymCh9K5yAwKfPS2S7XPAoDs698bn3EwcSSbpLryI1ZZnznvvH+zp1nN
oC1lC6jWK2dhFFXcol/jJ6dOj7fmL/iAYo++ywf0DNvpvU1DJTptXBHmqxuzAqt2zBQWQRcz86IZ
5xLXChf1JylgOEXY48DPTHyVkl8CfVJwYdN6Fob3TwyPsq1RZGCtEM2bK6oPPDbJMU8mIdZWp0UF
3tyw38NAcO7tJ1gpuCNz0PDWrlIP/Kql33ybxDMuOta5LE49QC7uTgsK8+WF4Uwr0SxN7tnZWRNF
s7MkQ6qmULzuWZlE+0D/gNbUdQIukpWxINbwKHX+V2Uw09w6tQJhu/lH/xy97mfB/eC0z+aV1Nwr
z3VLVxGRlz2/MJsIHXC9p7yxd/EPhk+hu8xltlaYVGcOAxdvbgR5PnB5ZnNKRiJrvo2UWen2sUwR
GgGh5j4OkXf03TWRI9WStzluRyKAswP17Ix/3YsL9wk3P8YdV6/Us+re4EQCYhPjfoEnRE93nljb
5eQDPhCVzgY8iOglkEPVuKYupcAbJ8kfnUpH6NgAqQrlJT72rQOO+0Lb5h02D/eIC/harEJebNkj
GYvkoDRPxDv/fon4GD2NZXUXC+drAGtURIzhhbn2MLKEfl3IF45hJ9i8nraZKBu4lW4gvdAL2VKq
SWiez4EANZtErUir+pQD7mRYxwZe9VkmSsi7LWQTW5q7chzXxN+QYk2mWH1XPyLoULihXMywm6Oz
o3VcB6h/7y7cRRqxXnliyHKtEYgNWyWpHoJ0EYVHIdKwp0r97VVclJ/Hk4AJCVkcA7o6hz2ZY047
k7BkDAjfPj5Xm6qbCHxD0yVj+JZR5MRm80/07GBJdIckJmYa1FSnGBxmmDeVlubljjbmkM1RWrf8
YU8X3GL+KpMqtvELYa5r1tz/GYHxoV38B9UDdH8Gs6cHWHvJePAzZFQsaRNq1DS4cBP7nehWQD6Y
/6hfB6Hj6AzK47/ry2s5x8xT4Iw+DIkAXwL1l8kyJ42XpTBFeVwUzLpqEPbCdCKPqOyTq6yTpSY+
EttITJZOnVLFQft1R4KOJ4aMWgg1MzL65kR2pigqzda+WpBXQC4MpDpTTtqUJeXeGH8v+5Sa72Yq
AFiWusORmXnfo81qzD/COJJWGdoEyy1FJNV5E2rrbj0RQVcvXUoB/Psyi3EXuW48Ayl6KTIufM6g
yFTjwvutuQcl5IKXvlQqkRLPR7RZKeeacv2NHgQSuJjqUV8rI7PRaSdJ4icSCOjCk52JoIDEpiDj
zqpKgQJ9kS5YrTRJE3v8GNhaZ7bVLMlef8xinRxCh6fHQ3du3e4lzP3KcaGn38lO7YOuxI2YWyUv
j+1i3MFKaeB6N9hr2AuqkICt+YEoCPbtLkcY9O6ZEdBOtk+9kXcYtDKf1o8NB4YSw4Pf/qQitCGE
PUl+5KBodXXn4ELY0/5DmSnJl8RzxoP8m8e4c92tM6fU/5rlwlcUZYEyCaQBgB62cvVbhuxBaq8N
2MfWnhz2S31zx7qk+COEnViqWCeN5UOCoFqR6l7f4VPP1Q9zy1sDz8aDBSztIRyP4eqmcH09bOHl
GU2a+FL05MXVWCCP6gDiUDAYzE7LsLzjeUMpS7KR6YRbKqAo2DaXhR4m85S5hKYp0fMhXMKL8tnF
IFJQB15U4zviA//LGu2w900GoS9+17bD6KyQO85yi9IaIpXQB0P4UpCSMCMPIxdC0JeaJZ/+8pYV
cR2shG87pmZ6t3YXWmgsnLLGxe7ucukv5+sSYCxaSnuBvNJqSUJ2KtVyRx9dBUe7vNjnHYT7nBly
zHUYdL5oQvg+5bY2z2krrenYpgaVK72vSlHnGlZ1fQWaxiY34cV3DJsyTdEBXB1nK4v7VfmCZcDH
gzs3ejJ7sz3jPwDfYrdIR/uc4HsZlo0DtZbvnvSLs67WZ1vuPwCCQnV6L6x50kSeiWlElRawd0Rn
J3mqpELAXWZdUOk3Uuaa064XUwVnW/CJN4IdEb3X+bco/2xuYZSphumvAwcOh9zM7OT66Y+xLoRK
S+OPteGRrRCPFOMtEX7qg1HdhiLRpkNTJyC8JGQ39DE1HjQwJ0GnRM2S1cR7upCew7ZjLV65rTdK
aSSf8AZkRM+aNU1bz6yk1qDyJTAIPEej/Wp8U55J+iD/ejUOuxQ5Kt6/OEn72Y/GztvffYdxk2z0
b24Ym1eLn6ZsxyCobfsU4J74Y/Nv9Kxe8SKp4AEcQVEXjj/w9ZFXVthhxUij+JZ3Azf4o4LmOgx0
nM4cT4ado94YdhHHIG8pF5WDqAr95NHnRqSH3kHbSem2W6GY41W/bh4ZEm9k3Y+jdrx/VG+zQl+g
oqTTwXPmlvYgyOHqAL71GUMm71NO4d1i8UVscnDgMdbLIpnLLFRS434T+4OGe7ippIPm8iXDPsx/
HHZaSBc8aEwIEi5Z/yXiJFxGLJMavFMfDfwF+xy2jJujLY2QnhjLIGMoVnvDvt2Nx14uCGs6IVpa
I7Q3AUQbI2NjB2wFlBy1EMrjQfXExw65ru41a/9l5bEWO5OK/WMEnSXtOq1CsBBks4zdcDBhoXff
TP3xp71i9j/2kuxMNi9RDAjoT5ZDOl4+qD6pKaO0qbSJxCn5DkojqDjT2r2zvo4FEp5BLWr0EMzz
nkVOTXNrE26ugNvgp1VHecqxy5wfYg0RHZJ0d+28ZHKp0K5SArkdrpc+SBh2+IUjm5EQGvkAfwPp
+C+bsFotGHYAPRQNpuAlpbFt6V41wziNfQXdztYGDLvHdTzK5uz8zFw/NrqfAIXV0BNoFLLC3lNi
YPBdwn/OUO1ZuBZn2RfIhuVHt9t9ib7s9dY1yrnstO1JnRB7aXetghg+PKEQ9Q922pQTDmoo4iP4
Daeeb2zn5X4uuA5q9B69p4THY8KovW5Z9p6R/eYhoclEPyQkCFxjQSn7kYMHtQ+EgOTKOccovx1O
2q+MnewzE6VhwBLzHigoTzQHpuZkmoPA9PJstm8oSf/HfKQIQEvpdITYGyj5Oph8zdcmX5AnbXM0
moBMu/uIgQgb8wPwnIpFzOPUEzNDf6EOc1/Ug0v2WQ0A2+CvvQ9lccuBLxw9q4LaOzRC6EpqltDl
8u4brDeFjxv49mPQD9TVyeNu2n+oK5c545CKyq5Rw8WgGhqw8uGL+jB1nYPkgEDPz43p9BM3im0u
a+mI7S8jDH5ED8FLQR7wsUr3/uGeQcKYA7MrIp2RRTkn/sn4CSkuQ/v5COiPIWniUmTVGptBh8GD
bXRPPEy/h43VxEmBhCuCunSkUWfgyOFOblc/aQh9X8o6MTZJpTs0xyyqVGGQsu9JVUlzWw/v+cZq
9sBByo5s7P1hJwd9uIqqp6H77VkEeVG4zSwtRdxP0Bv2PiFmoK0yocHgnXK03EO+KOd1qLOxY7f+
F4xBJtA0rxHjRXvR57qiekgXXlZdnaE+QaS+2dd+Dd1NmB7n0ruCwRYFwKsQ1wbjZQ7lALKprzuU
hBXC6r8Yk6iKG0CV3UyMpSO7Q4Wzu3aX0TlrbL00aQ8zWpOz6wEJKbyyU4owILR6YIv9OQgkcXbr
iVjkQv/RK0z/vriR7bKvFeKj+UBhld3wp1j2AF0dZaEO3eTTBs0H82bZCZTBikDfNFBse4KjtWvr
u4cV5dxIIkP1MQMpezV/6R4wp2ev24yFWoh0eS1t+1BCuPYXdEAlM+4L4AcRH0iNQb+wFlaBlkfE
WQ3dCBT9Yq5iHMtW96HixL2NaOVpCugA8tG1XJCKOWOWUGWQA3bmiwhjt7WCqHjzg8VvpAGbVs3b
BqgyEeEuMh7+re8iqRobKsQxoTz/CjeiGUCJVRdTUuLKO6ncKVlJ4Ran6VmS0QYAXOM4mjpQLP9/
VcvKWghofp5tOXz/5+vM2u8vdXuWMGwq+o3ORAl8HbX/RjV4ihRMmN6SPdYwUYU0c8ZqvmuIxfhW
Qas9nqDlQrW1bD758+yQihav/J3mp7TFSnMgC4W3M5NJk4aJU9I9qchb70p3Zl26aHlCZdpx8Ito
k/78imAx6Mjtkvz4/QkpQVHLyY4reqf9fIbmU4oAqnZyhaRjR0O5/CWQdUijn7sMy1RvQm6PNpEW
veKfrvv8X1kFYcBV/i5kb6LmbaTIi78apWuDfsgAUNBW1JSaAmaqi4GAPJWmQxLrRrQZaoci85eW
uwbHJQKui4qigrYe6bOxhPU1uYDKkxNOI6L5cb781mZjFwOYZufQB9r5rhj1gR8AxeDw7j3guS3y
ZYjMp+Bs4sGb0pE35hfmJnhYA3rHJIIfxwh6o2bqq7creJpAZKwpqp/qlrPRxoQWwt9w0SKDlYQS
TTq3HxEDZEYSs+aq38Kkr/d+Z13Vd3+d+3SK/PoUTxE3bmFsJ0P6vnryQs8FYhQ8vJ90JHVLEtEo
pc5WLxofhnqyQpKlN2J0Ag4OQwlnW30iGLvPzrAlAWpiAe9iKPwrtD757ONtOeV0oetqzv2It/Ad
z+IhuBNFSguizhbZrQq+FQYV0twmQn+zfzDRdDquOeTneNMJ9VYR8XgMWvX0Nh3/0QMa0K+HO8TU
ybTSoMNmiwiHHrbWgSh07icZ00cSNzpIMfPrmX9XgxmeovtxdbKuc/s4sSbFGCvm0NtWj8ZuGGes
7Td+pFVZTDImmFW2tOi4BNFvu49aNRdeC6sD/QvtP0hqI4S2HKdnFGbvAWpcYDh4wCdhrtoncNxp
ygbFUc/lqwvZ/yayKKO91YQHtlAk8zR3Rgdr9WO982rgO5H4V5JyqQWiRWQsFNT6PlTjFuy6uz8b
uW5NIEQyJDT01YurxB8Y6unfrLp3V2N9L2bf8DYmtmiDBycKlvca/cW+xE8NJuNq8YOhPR6dcWXY
RW3oI6Z1kYgxABhWLnyOT3lKpgJt2o7r3C4KFim2rAjjwCgZ+7R+C4AuHycjQKdBctqpIOLV5P2N
3PGWsRYTbCDwhraTpBKs1P4aG2J6qsA09mU7z5KiqfKNOTWxqMc/i1HRdcWe4IWotqmxrQ6X7MIQ
aiuaYutA9aHwLoUjfUmDMtpaggD0Af+D8eNvmP7OfbKtPzUakMZKPffR66l3u45+QQgMAWEb6BM2
45R2+UBx2MlKsa1lrHMRtmTTktOZ4o4mIknwwiy7RFdH0P6ZiFFuXcE1APoRPoV0ZLrI5oxAOxtl
u/pQxZwf5pgS2XJXJwy032GVaEXBzjETmyqE8Nl6uZkkhjSzqgPnq2JyHE9wE6OzYzB2mcuf2fRP
L8wetPJIt6B7fevw6Jq5rjsZXZRIj+ygRCO/Q8OaWXFZFLqWCbyxhgAio2JuNNvZmOS0Ws2EPopX
kIfK3wrtZXEtlztR56wU/EiSV7PyEptef0EOHW3EouuKejRTKN0qwvDle2iaNZic/Edeexs6p4uG
fAXJPL7zJrhhTiOr4NpEumwu5S0B3BPXGXBgSZEqyjI1wCOy+8/kAOphNQBt425I3gg0Mm3YD/Bw
1nvO8WohNQfV3FZnsRNBD87kj/RIt6SZTXHvHYcmeS6B1bkQTtixbLAKC4UplamxAL1RzrVagMeR
KpCsRRFgrv4aJS7wIJ8Q1HycTRSCMpO06Qr3TAhB7QtmQ2HL3H5m0pKek03EKFfeE4+16dJVP6dL
EAN04focSZMLORURwBGk/tCf8GYYcdwearAZ+Q4jMAUEsyoVWLHQdOmowPsIciX25B2K1CaU0G5q
x4HIQJeX3O91L7ThUEAAUOXESkYyFBzpGz7mHnDDQgzPeepz7O90NxQM4ubqthMx2EOnwt63kVxg
iLjaKWJPhhQx6jFeEMIPp/oQf9Su9Y38NrAr8iCNLGXTYywPNToK9uRs6roIjhzSCGISfLVr0d6f
OR6RwVQn80kw6kCJ2/Ciyg6ukrLekgo7rHujgPtYg5wxZ06OlkbVCiSyI+TLB/napML2b2xBTan9
Qp7j7pU942popYf2BLwpYPYe9Eydl8ec46a7DYfMheIp0oKYiG4iwxQ3vu6bBG74ZqXAaDkJBJOW
V3AoUewYCerHf8c4glLeqjhqaarBjgRzy9kfDnMmXzGfT2TG0PZ+YVlMrbRG1s3GXceMGJ6Y9zSL
LqzVFlT/ffIPPazyiQAAtMFR6qXNni1xzYJn8Xls7pJIfJYlQAZfIEmHiD5nyXCVKQkE2n644gj1
oXh9u2R73a5+teEZxfcDxdYgY0zbmqtDuR96tdKfctr007V/LLXDe1htk0RZ/3P0L37CC+iOQWN9
mb6EEc35BRW/1nefTf16RRsbBh0X111g60nMY2c0qhg8a/gTAbtwcBhcxTQFJePmBjE4fW03FE75
NzHQFum3bOW8ZMpItGc3iOf6LCDdAGZ92iLJoM15D03aUpg2Ffh3kQgjpky+fmdmEFxbFyskMATJ
+YBDffHnb7ewiQkuJeswPkqILpMHpWhgz3MyZyfeFWZ84KCm9VINjgquPKU7zm0XT59Q8/fXtCJV
LY8aHgEFwjeX8fn87TytVupe9CsPZ6mNLthtDBBJFpRh62AZof6OdvEo6oKVrmY1znRJrEr7JlCf
sQNp+YPlUqjI4A3+USdVnCUdr3Td9d88biOuWKGASdiXe2QJdtBmAL/ZoRNvcseZwl0EbZSmbS0t
t/3Htk+4wHfagxuOWdANsJ8RAFLY/q+LdxnnKG0koMOfcX9eab7avBYtOiolZW+Z1f3lfshN56tn
xSbOL4/yvfNxIpc/a7qfiErRh9M0YnLK8NmdZZ9ILJlJEm/FaZkn3ulDdvZ9/d8CMIK7OHCqcfTc
P5dCW3vqoZ3+dHfI39rH0RdBu9Ebyo85TsffQIoFNWGHSimB0OPDLtcEaYshHL8dsWAvAo05EZNS
h8UCc2nMsguOTQTb7xa/qzzKn0tphNR9N6sstFimumWUldqL4Md3S2eKK/b6iE/MnFh3GvWJR9Qo
lrY6NbXUxBcApqrmylf3ex80d1ZKNVbUozZ8JKDUBhgCsZAl1zPlCTz9doSROC1AS8OuBNZNpsWp
56xYfBdwiOH5RUB7lVqpVumk1b8WU+iAGgEVyK4y/f+d0QLgEtXMPVjcu/XZtvCfyxRv2mbybc29
CyDMx4M0CKsmz/FqbFvtDLfzrXZIY09tYQ8acB2X644V2GCh17nyusHlyMVvhfH7Df7ILsV2E3y5
Pm6/KWdQd55nXyUijQXAcxuKL7OJM10eUolKhzMyHT8bby0srYdU/icgvaEofD9DVKf8mKAsfn7n
tN3B2Dr76eMuVP46K27xjVzk53OT4+9tn0r+/zom2Oc47XFpsfjkSXdttdwMJOpSKnnvuWD5dj01
jsupmsFtv42kabIJmZOSpQumK6ZuNgIjRIA4CVOI0IIlrAVMdiVBBROvR0N0GO8QB+5ZQni8AzpZ
Ei8aZuzB+tRWmTI2OB4pKqA6k/DjuEYuzpn0Ra49N2e7B0LoAjtjoDCCWEm+3Vy/dGSwiWowYMs5
jEtFCn9PiJdy9ZvmqWu6Kmx1BFMTqtBHW0WW7PA6Oy/dwX3yeZYN4Et4Q5FHbIk/4uRa5XmumozE
x3qi6jwx4+WChoa3G364U1U2UVbcHoTvs72ImXvrnwzyOMN+USWs7uDjQ/EgVWKAsTCMYE2LrFr+
H2Ju4yB1g5c3v+Ix9mJRulWF0+mV8jS3p0Qh8uqWM9OSRhZthClu5klYQUAOAEZHm7J2MzH+ux7w
yCk4ThcuKrEpvkMG3nyLbjXiNXJR/eJSNr/aAB/iUq5h5bQILfQfTUBSCEqmVF2EaHCCDUQNM23G
vzSdQkManpzjmO0ZCh8G6Cssh93b6MX6KgyraYAPClEa/CCbKPcDGxN41UFjQV/ZUACEni5rCBHv
qN9kWOSxNBXvFz7NUDgIj7fkR/lrxXUPNCz+WRHfLOaDBa2jFkhSSCc5ZGUMSJ+xVWEqwd7CdIa/
56Yjo4VxLOTasO6oK/urgvV70JDrbMFzcUYgnYHtyggsn+D2ewMYJCAWVkW82ruVXj+gKy/eVxKW
l1lpcRTGjVq8MS2//Jgoka0MZQsPG8DQgth1SDWMPlDrq8umouOQIpWxv6rm1CRAk/TAppMoThtR
KIoDRakle2197wKA9wje8ij+A/IEQyAKc5R9+8LmFHcsLwYOaSDpmj1gLHdJim9YfZQyR4bSE0xn
3oWp8KoJMFtW9jYkH2v2mZCE0eGD77wiyBaHWVXqcvfzw/owxsw6ShuuncIutxxGsyCoKaoNylmu
VEoQNPRD1ZIMeD38bL8Q2PaJ8iF5t7Wd71wV5Js8Zwgz9RfqlyTU9x01WCC8mpk0Wlp6e5PToqVb
ZwqQkF+xVSEgAHn2u7IqzjdwTVa0YlY9dr3X3TLRV8H/NhREQXeuztRCCHl6kWwB7uny6Ze0ylv8
bq5sp+o8zNm3E+W61ncHSS5edCF9ax5MBoW1XzCpgWLy6eXXdLIaExji+s9nUvzRr9crGuxZCMw/
/beAfLQK4wQuBgjsv4IwUpZF5c2rZVvanhWwDVFfJJVL6ngJS3ULaJzZ5kgrTEUrtSdQHdKSvuA4
mK0a0X+jcodEZOgtTsj9TMO4YyKYlyCAFkcE3PU9grTENNqRjuZCq442R3ixLSvdGf4RfGNSNThL
tCm6zIF/j9G2q5fkZ7cRnrdK2hICq6F/qpogagkBlooZZBM8UDjBsJQQwygYXDH6kZb7lw2r4s1o
Npyh93GnvL9afl+msTNcq3m45xgd7Fc3ZEIbUoYa0MXcgDz9V3jJ9d8I7s29BxY9c1KZr74ouZQx
sXorrletn4HNb0Msh+P4zeibwe7F2+pfKbqROF6wbyKxLtV2BrByZ96/eKblI6xvoLafSLlp2deY
NUBPRuYjYYGKypoqzXQWRpGl1LfeHMgB7FbZdU/PpExde2g4wzI2u+7yh/SohqrCCMpNvdWo+KwH
nPXfepYQbeIzp6PU4siEeVxmdJYKNGzPZzEgt+fmG5ALtaxqF4Dhm3+BqK2ZaELXYWbrkgnOjNMg
fsGV6UNpS382fN2py9PERinR0ATxBE13nwqvOp/w7oNN5VdzZWDtA5GAxVb1831+b0o+Xmyy9p35
0OIxPXyQjgRpuhHSI98EGhoWNhEAjdV/cgZo6b5qGaLrwBu72ZrF9cx2cctjhX1//UgE/o8Gxwic
mXoJMAe1xsJCxDMB3ABdRU9xwajo/5yw2oi2ZAtdZUifZyLWGGC1QrvTwqUfr7ELN8+pcM78hRka
/CvlBJiWRcWHwyqZ5lS/8ZKorJiSEPV0zZa2L17N2P/3MsjiWoqWeZiXCDdyAo11x//ZkKfrx6Ck
vf/X3F1gvzF+NdaFsE/vuZg1sNN/+4OCDI8KC/NrUkX+irlqHZZ76QKrRmpsM6hSv8GU2HYfciEV
5ts4JeQY0rVUjWHto5mWBeLSzyQYyEc8X86TvLffDFhmwDi7BsVdzwEJqEp1tYq0fRVmgJiuPDyc
4m2KlYxy1HaEeQO0j9/0h7S9TGPXRAcLHp8oju0b7cihyc5A0Wh4jaTJPhXXerntr9hKJUQS8zUs
yjQF8mM2scP5mXfaTi57gCJoWkijGc/MBGxXn0rAuQrrmaORgt1sB+QJAun2cttVdRkfUE98bBEG
43RfMWw+ZbAURQe2+u8kg0Qs+xnBLwOXJcP3ojDLukcD1iRzu6Q9XyUHH1ybscI0IUzZxrxY/oX1
LaN8MytbrXbrJprCTrHj+0k9LwSlGfETQoHROHY3Xt/ZOx44uLUcjgd/ZQtThTN+F+By+SJdQY66
2+Wsyfb61tFAFar2RpUv6jjSu6VW0lXAzIiq6AAUMbFH8xKpR8DPelsarQXFN90Hd+N91rn9pW5M
FAzRk9xANTHLxxBK81TSxS8hBbhIYuovK+7yIorARTaAY7K7SmnEy6Iwr0JnWeL7SOEsR/iGOIlx
azB4zeq9PKkX1QkMJH0EycsQZWfRjujHSURpdE6Aua53ZV/S9DG4/6EnRe8F7LlvzILypNSCVtT4
irwf3NJ06qNjylIEEl2g70R2Kz6PtSKcOSEsABx/7etqzaSKKFIeXnWHSi5vhEQhmQpAfkS/DMBt
nU0l3QbzkWh9ORaTWjLS2VNsALWkCG7CL2V6B2ElZm0cTct6PtVAGtYFPEKVduSS2Uylc57vqXFO
JpxJsTxG1JAI1dm7qF1EgfHPoXoI4bs2StP+HfA46l4m5fxrUHlh5/OBR/mtj8cedB21vvT4Ij2m
JNGFF4Xnt9OyDeOuvpG88W+PT7V+Q5LQ2XB9Yugo0vA+JtY9bV1u3PicDKbPc5l8FT6qcW2o1Yog
mO/9+YH7WxBIAvSI0huzoEeQSliBOii79oHG7g2aA3C9RcuC0v/6ELNCxagnSsceUZYF5RuWCKiN
WWuGziFer0SmkFy3sebntE/zQ5ZWcJfutLYZHKneO6IYR2P0c0LpDhvbUar+/Yylp1DRydHM6nyG
hR1XDzs2mW+7XQL2ZtESGguc6DSdTPH2vuOrZ+q2d4ClfSw9BQH2iM9AUAI24ueAdVi2lm9/8dg8
XeB2ikrgK11hMF90Mocr+2VLEKJmUCKE80SLXHsneC8WMBWBCxgzhc9T5+sX0nS7Gs71QP2YPzgI
x/uqt+ulA8GzfcPkuwMt3jcWJ5PoTY+wChaFu6NEevXhuw4urnMmObe2c/hmcb7fTuEpKpAzAE6L
tTGEnjQiCPQPCD3OtrvLuwRd3Wl70BC4cKff20LbJBPtU5ya7ufdj/QqRFQVhPzVJswFt0LxY3N0
s9Fa1jV/LdBM2QI6YiAphXOmZ2Kn3g2M8ktw+Tc5dZ4epzaGA6W4ce6WDDrnmHXA1dbwLVYwfZAk
Cmpp7aF/P9F9UzCmaDptxLZFqMvSemHhUA9f2SDMkqEnBIVMhiMqp0e5MopBjUGTSjKwkS0nC1Jf
gDORzbuuKuFqsZCqeZKLhO+WNhneYLD/tYZax/okbRGIE+g5w29D8qPv2ZjSrf5ndQmZw8asm1ef
GeVl9OW8yDo4cf1cmgxieAkvicLH9tiC7597tIcTGvBGUdVjahi2xevRlP4+j2p0l5kVDSBToRtc
Bv8hkQWWEubCIrwUITRSVVs4ed4jymwx699OQmHwozcOn48lw2Ya/MI1DsJPhkH3ZsKjxHlORAP4
EI0lkPgumNpEuEH3Zr9TtXnbZs1lL0Tpc0z2SRfcqdpWGC/y+bT47VDZ5TY3sYLOmsJQM4eTMcHr
yAaRWnoGU0vtmGRAlCoHway+jdh1AyiKyLObwu05sQPebYB2GMn4AJmFTNeLEyU6H8PJeMYrO+aZ
LA2OhQEuzcJvaMjI1Yry2UjhM42kilWy0mj84wdOBuK4eo2P3GnFRXtvaKPxwzDpO5QTFC+B3cMQ
Y2camqZiG3SbXKJklxT/xT5BtzVrEE7A1z1Ab5jKCLJQGQwM8LZlvRyiibH5uTSiHlLobTzp1gws
rlE5lGmqtQBtmr2rFQijv2E778gy0eNuaUvJiI8gJXB1thkVzskHE6ck8iw4XUXGGAv+CDi9cXQj
29ToDva1zhoe24+tqClEtYDiraJB9zM9WfXONXK/Ssp3y7uK4vwXUBMNYsWGEQcIekvcWWYwvYsk
Jr9e1fgOmGLZXb1R2U8wAluB63vVXUFh9b5FtAENlOirVSZ9SIXQS8Ujk0eVovVi+vy1AsCFiM+6
JRDFJQDQhsum0Isyj31kYrqyaxZA1kCq368bKoUzRi5bsFVXxtdhPuRhwgVem9H52dT93wDcEHvd
Ht6wffFQvUgSy9h4fiASk9mdt2VW3b557fH3t8WeIrUGzOwhGFv7QVm4DUGcqyK2VzvkXdMLBWF4
mfqelXXiMF6iSIW/k7fYYVxVULBKUSCnTTv2+ZusKHrudACJVfDXO5O2ax1kbxVv7KqclQvb6cCd
h3g034U9fYNR5+jXIh/4OK5Aqb6qaskXab38MfELB/MOkqflwVL+V29azIK1qFKhCDOieGLwpQwa
vWnWKzDYlGaSTyhyQF0E145xVSQB54XDTcgXGOl81pdXjQkVZjWYjrtxhd+5J0p0xDTyHVcW+3MK
LcZ4MaGuRfhiQbYYo0PuiUHxIOb/W7jVjXHC2nlG3pTKnHwxppkiYra1q6mkcqZlUF0QmB+ZieiG
mAVn5I9fjRh+9ayQ977URVyEhL7GTBVmJVbTbzDHL8aG9QqR1+potEkRDXh3BwxYZOBe2bWaWBRE
VI0t+DRUfSCPRMckIj1TSdrzex0pZOO74gLVEpnarqzFUSLKqhRATspc2P2nAZrew+82sGHrdyUz
ZhlSUyFZBvNtwn2bUnMp/gkMY1+z/AONNmdogdOIUOSkEX4vxe+R9QC8X0OLhyp5YgLJaZALvO8u
XAuE8eblPvF/UsbVLJDIVL7uRMUByg043xvCkydAIinrvvfj3vx18NBCGmd+/3K2ICob3sE0Jr6H
OgqgZfw6Q50c3vpqdk645a1zDg93GWPHdN5BbO9KL8E63Pph6yKRwT4wWyN3ECs05YhICCMgq/CU
QrOkPfjZhgIILiM3wFHkTg3tKYkq1RRC3Hxp0AZz9twpNkdik17gCQPzUVrS9ORtveybn9giY9yk
rMAKHT/3650DczYB7HwHoDu6UQnMEjpiskYxfoP2n2aPOrCT8WLycAxcgWWmIUwHvhs8kBGpiyW8
lnVAdhDoIGrmq+zx6eB4E35HnDx4X3nIbgbHraq3MLGOe4NXy2HLKQL1vnmm4pdTmfPZNymmCl/b
AgAzW1SFXqnapvUDua7G7bt+yx2A7VlOyoOwuElsZhbsD1hf02N2YI4VZ3KQXLxdpyTnmJbhwA3J
sgFgr/8h8OtLu9qIPfsPjCHcYMELxDitLKh4J6f3XdQr1FM7jQgUFHwbE/KAXKVT4Aqw3Z7q/Ck3
FlJ3Eag0tyLfxojh7XQ1b6qUsf8+9tuM+QGOnWPTJYLLWfZyTOIBc1tQb4nntscVQBPbUbcWTo4x
9EjyqUVWRypgXngEKQvJfx4J2ehQ3CqOBMSSUlSuaELx2OAu9uim8VGJVPDrwsstoYdOYSVbxT4w
VbyDti9QrqL2ovZvyd6IXLWKsqVgGHHlYM5ladXTNRgo1WUXfNtxuW872w/OLvioC7lmm1l0s4Rk
izwodFE+AUdk07t7gZb0IWcx5fdHgBpnDY5sH5MqxpHebMMGmcrwVK+4fcOsePJeUpbb3bE8bE1T
MeyTvYOKvla91Fh9MWf+W/7bZ25ZkGHMfzIJrDdZ28EWvbJwe7CH3zn28fLJGBpzQ7F+0G9+DRan
UOy5hym9UOzQenuU+YwPpv1P2QMRyHXmN0o4pno82GfItw6ItJ2BEHL0HpcV7wL6pMFbN0/eZehe
70Os+v8n1rj4ABTZUp87/ZxKitHUbSKdHbWVapKAb413+K2OrqhRs4T80jEfqDpQEWvIHZ7b0WSb
MnpHsF9fsgjrN2ofe7SPoP9yZdXcTcwPLK8YghcrK77AIYoPlOBDTan5mqhOtb5HwExDsvH/n9KV
YelK9NiXofVLk0oRskZoOx6D81kasx3keFP5WIhl4pGfWo7S9NM/TLx7pEuoHENEbLjYEWSezcVT
dTni/nGSz3pLGJiWn4KI1UNfKnIks5rfrUtOAIq3q+M4qLjQkCZfMCbwZA2SFYM/Cm11e7n2xTjB
nmJ91luWeUBGRC4VqA13TYq22Mak1Cjy9zf2g2/fY6XoTpTizoumGvfBKTWjzwmHSoseQPnm8f6+
DcAZ3020vR3uJUOPlMrvYPzI5IHEyheLhkON+vVOy+pTZQqGDKmbnV9axsUPIpPcmzWQsJltg7M8
spwf4/B5X9mdgF4qkPKIAIEuhKwQF7VEOv3h3lhT38nrjZfgyg3vRR8jk3YLNqUWH5VLN5ex3cvr
LRoKMCIxrbUlGOSgKwv0YXzsB/e6P9kGkdFucL7bZ8vNAet8encOl69oPqXGGDvLiCP0PyP0IYsz
DPSD1wIDx5qD821NCaKHNR3QZnQsJi7flAkJ73cpilpEjh59axK1/gVQCglTJ/IFxgh6gEPHyX2g
/mWW2StLfUg0xQ3GWBDQUB2aNdpxYKK+tw2RjH8HjQpwZNzsBtDzfBLdGo3SmDluFdmMp3xH8Qbc
q3ucKxSfpm2+1V8NcNcaNxbmIfF5S3ed03FZtyqGF4yEv2LzWySlK6r4c5hmvfYtGzygYK6cyFXk
1Xx13k/8lK/3HGaH5zZ4ScAsgB7QqDYdn2QsXB5HCjgq5w6oBhJOouloZD1dgq+FYyA94TcMxtFz
d/WPUIzepjWETqGqV0FKcSoSYSANRQZ9YWelR06S0wrI7rxrYI0mu97YwYFOvO22Y1F+N88y48Ao
s6hI65KwL6xo35iAUMBNOUlAXdiBaEQ1JzL5gFJvjJxbCunSSWGirvYySyEeIBzmGDjZmeDDeSC7
nNaR64IbbAS+CXE89Uk/+Mtyw0EZz2iYUDlTYllyv4dydf+sM/D1273VcZoq0yARsX/y0kUWNDho
8DaoWfjyhPLpUDEo0tgTuI0igceqxPXtuBNxFShvghdQDr7vUqnRZmEC/Uy8bo5CuS5xE1MJ57j/
CTLSjuUj5ysG4qhq5RmX2VDznr9VMbxfRL/uC17318wsndYH3Iv451/+VZTmmsizGXf8ZkbJmaFe
N532yYnGRqpOW2sgyDbx/+U+UcXSApvVah98DmTg1CtxqmYwTmdUF4WPH2bM9yfohsdr9R0AJp8u
Vs7mX7UjzKRK5rRUu360WmjFyNicXQ+FRI5EVz7CFZqCahd1g0T/SaBPErrmz9Af5Seq/djKhxcK
koNCItXNkQVMdxYs3KoHQpQlJVsLOPZVgfU3GHi45Y4aw5ZVGlhHBeydx/qPwTcHRCwmSgfggNJp
BYL+oiKTx1UShf/7FQXMX4ThYRC6RxBxjPM4nsfEMFVUsHO2/u66owt23y6YTHf8F/1Nxdzb5Bx7
JLEp9vVRoKdbAP7fG0GPEYQ8lYGr+MjBqdYTtbB2fL/71X2MtSslqOkWRuNa2Rc6gKBu+2/ZnBEw
tX2VeLhIr1rOlwI6gaOmJ2Atb4aUV8ARBDk57ifnvZ22wzEdvHH9qWgLkXicX1Hatx8d7uXa4MGg
hEsQCPXG4sR+zY931ixvCrYiw0Hdf12vwuiPsi/CowrNdC+UXzvl3ClvgooJPV0VEd9G2y4LTxMy
hf67wrdNF/KvAev2kdIduzQ5JsT07nf7ljZ8EeFRyyyrbtjN0oYFptkCYP4ZJY6c4MmuUgvwDbg9
3kBqE5alNQWSZ8c6KHV1SsPvt/rK6EZo+ciaE/+u9WhtQysOC/iIwg4ANfGgwRRSIeUxiTadzB0J
HvAv5G+pMdcbm7qDLavvmIGR4xSo5+QzGyrZ0eNkZkWUNNPDakwEdHhPrLVlnsBsBxaeCCjUDrqM
dU6DzdjM2JtnKdrRQJoTNG8L1FZS9cDecHI2A7SufhbjzCVP4pjgVY5Y8bqE+I2SjP0C/WoAf8pI
zHKStiuRAbzAtgL+faFAAHzYsBPTnPz2kelb5kSlMoMki6H7UNVO+cMdTUbfi6VSd4FJTt+44dJb
nJiVzyA/nUOzteSkgMKqxs658vOc2AmjEIP7LqpDSgGK9uh8QzysWGynqeHwxfL7ASL4ixJBYARw
HDMJ4zTJfdvBkXiydCi+tgRaFjnsOUdiedcNJOzXD4blab29MiuXMKGiAd5+XEUd4aS7BRsTsYIO
N3Ur6XQ1HPnWH0BKDZ49nThkEjmuai76+b4iKuJaUq7pM8iADzsMWqmxon/zOUKOZQFzhhC4YXFK
zbWA6/+pe3Bfp/vdW5aYWH1ik6EK5/LzCHu/A8PBC/26qEUUwIRXqC5+RVpjVfLvVHOfwJJ+bwGa
LuF7KSbUwbsoMrUKdsVkdGHw8Hnh/oY74evtf7oOH6uJ6xgvkIRft83ITH51jFRhFXYOtUoG34co
lEDCF0qEKm5Q2k11++ZQm2+qB+VPjdxaybhsA89eZXXE3iXSmoDhQEwc43g+LznyA1uulyLAO7si
aOqKJrHkGRKaKn4xzYXPvCDfTT9Axxa5iQsy5P47zYlFhBSZYBwqwTcrdUSOMac+Hq3r/21eZWLC
E4CmQVwWXvDbZ3HQiVoFqG4n3kRCOmIkTShPVZp9h3JFRe390itkIx9R1RiGV8ZfkFPQ9hr1mXEW
pobI3FFkO+SejIYSzjj5tWLJy9ha3QmfRf5QvxoVFgjNOlv2qEYX50XepHNTwp6UvAPKaGVVVU7U
kjt3GvBicOwJ14l3IXwQZ7736bE7aKgTh131t5D+vuWwr8+aH1OiOmvBCv7ZXag/hECVxfd5eFtD
KGbsBRWgSsp1xtxanYfLz/KuqFzYYnwNLE+pkUmIJa/6XEQfj8FHCJe+2Lx06QH9Qlw6tS2MB1ST
xgnVplf7Ank+aSMj5Sddhl0ZeZo3Rsr3oFHAyXHkxaZ2K7ujx0LLvY+f8iy/UT6Goi+zTv9rNPk/
5bhE/FP+Tr/rAPBCrLtzWMBfJfy3zIywPk3qe2Yt7wBrV2O2vlSgG6H+RVycyQUjD+W5IG6EaAvf
sIkoP8wWjYaauJm3Hp6l4Ubk80Uv0LDPT2IUnyjRLxJqDco+/bighL0/1qtBT4qT6bTfIYZ0gPX7
UxLaC3ymBPWr4FhekGxrMzzxgOi/53hmgkQb4f/dOlO6qYXmb+2PEeiOMZLUL0ei0lmXME0f5eWU
MYk1RAWTc1IAlg0d5Nqgm/pcz+Pg1UuYmUyRVgMNFNBAVTBQLTN/7ZaPQbRSUk9G+Kn0WOuN9kyC
07ztqn0VLD5xubrRb9nO+ZxQ3QWZ1ppjOqZpiTh/S1vCtR2W9nA9Au1ojLmjqVv4SdMrG19MEE3s
FNC7Ynlue0YWtZLWbydTyczVcGXSG+EsK9t9Qvhu4EShZINbSHD1WGAkA/bXfR6CM2FHvesYuRfn
tbPHwu8WEaezwZp7ju00kN2bZHCpj7tmpdolKvMmpLew+VSB72rSS+yNkjbe4f+JFYp5WaFjNiS3
eKAfM5tXOt4FBtN7LAXljSssqW6ag5je+aiAruTmcpX9NgPMPOLqS2l+G0vKX9oDWSp7VfK3Vd2A
TgD7t4Qjel6c1e7/pd3+bFB1mLKU4e/DmN7VTxtmfX3p5ySu2kzWQRtSVnKE6eCbfLubYv2MOJ6I
f2JCyB16dcBFic9JBAqeIn4GT+gw/25/e3KmB+u95eqGJ/EWRiEK8kjpAuIsa+ul1uYNKBCcfYLi
Xx65bwJ8x5jfrpZjjR8VZBpkGuoGQ5g3ItXBsEtyfT2H/aEE/DDMGdGIHoq4XpUTDxgOQkJ5Mc3I
/Boi6DnhRta/XyVh7r23327KQhuO91u4vc2MJWEweNtdUrOYX90MLo2Ip4FYdkStoDd8L4L6RAdG
uvc8A/QTf9sMsMqY70VAJ3NFsnNdalcFs7GP/428eM/Bq2/aimudaIpcCICY9PymNPMo3Re5ITlJ
Kj5+cXv0fvj950KhSCZsCXrhb7NtnEexUAZfFnC1O5czaLPGkLJLhATn7nr9fcQMRgi2lep/mgXp
dzBvuWKlXzgxDYu4i5AkEtTTY8V54jw/Gc94/21X1A8+opg0fLOEDwApt1oQkGK74CQoXrNuULK3
Hy7ne0l0qdWeYzSxFkVRuceTnFPKwe4Bf6YfPZrXcs1Vg6olzLgwEVB+Xw9cM5/ujh49rfcFAZeL
4fWFYcO7un1DNHSbmBt7ErLhvi83YCFpxvdYzOR0qbVE6PpnUKJux/P0u0g7kp7SwYYlKQBTJiCf
IVu/OISHwD1Ndq2uHEXb5ZiStY5ySq6Fmd4ILreYniB+GSWEbmM+EKOUg4EBhmDsk00tT/aEXBCy
7WbCA9aKpA4+C9334TmsgcQuG144lGWauXCnlxTTk7dO7QZOvxcZyAPpSRQ4QOFPYiWw5qO3+K4m
fxpYjXnJiMR3Xfk5vfOKJyMkePSvfQ8/TwgJmjPJNMxk+/qKR/xHUFA2TVMEVPMHxkgbg6aa3u0a
tXoH4Mm33xUOlV8RGNupoVXkZ4vcr/XVJWhFK9ZVuKpEVvERyYIWqS2jL0h0tJeAK+CXApkPru7D
Jfn9QKlKCFyrdaJZVAyqRn2OBoUX48vk78guQHLJaXYC83qANsHM7xXl6yblOWWNtoZkWKMlG+CZ
B4g2CVtZn6ZRJtKCkNmcLRmmWFbPanMHJ4DFOxhVK46nUWB41ZUTtBPxhYhPyLXlNsV2kAbv0gXL
yD9ITSx9xkL2o5ZEwWh8ZUm7aWgvSwE2lFcPannNw65/sb0S83Bf6sFI7Zj+r12BIPfHdXlod2bV
k/XQxJs5Ug/JLniNHpN7iW77kQIPuFlSCWMuXtlynNU5d9ibiGMoEPC5YAR38zBFB+H8z5HNsixG
efO9BgF3Q2v3CVfpiHvm/UmoeUtKCV5kGBA8nF8VveO5jR9q/8kpN85J+iw3SqajUki2nHmcPyyM
6HQYU/166PKlI9a7gxrwW6cEWNiclDbqOovXuV0AbFXFqxg6urW/1n2m9cPfVHrhiqI07Ybhr9QJ
fFRn4PXy1nJxUY3B6CYEtaqk43Kokv+UKrvJxVs8uVIKr9MnUPASTmckjeADKcjieHEgF0qDwlP9
jB8We3AV7HEzLo0XAS8NkU9T6Ba6NJcEgXYEOiOdxXYgMbOJa7Id01sOJiZ/guOKPDb0JS6Cnh35
4WCoGH60ADZlQSV28tw3lFOT+/O8Y0SUT3bgpXC3Cnh152HrdURAqhQ4BNWbe7feQa9pRRtJaFIU
tL6KujKezF3fFynp8XO8HDcsdKnkxIRsmINOzsoxOsPGDYvswAAwkHiUwTGyvCHqkSXz9Y86U56u
JeZQ7c4R9zUja51LOQQIPlOnb/ypQ/XBvEYqc6CZGia2vehiHClW1CHv1vzsWHQswQFBTfMDBeK3
PjQi0JUIQxq7F45mvbfSF488KL3LrhtzEqtpbBRyL380DKc8AD5VzDbOmVl5kCj53GY7ieI+DkLA
HLJmmG2wJj462WSVJ45+FRXd+xLGekw/MPNEIT0CSpX5+pX9fKrh5DT0mN/ek6J/o9x77y/fKCf3
djozNG6s5aHSBfI31coKXABseb5y0LRf5qQS6E9+krPPDzKa9s01+Cvg2GO+H3sgwKc6b2pWAneb
ZaK24OZEwhwQCJihfr1rgzQuHSM7+NeBaymyp5E+nxKAvTIbl3WSxuieAQo7SS51tZ9r5QAK9SjJ
Cm3LjAR7GUAjaBVyCaYWzXBa6JmQkCfikqrROugNzDZRvj5BboCUWw8pZs6RyvlwkbloJlnJ9RzL
OrikSndbKJWqvPWnhoiobswb9eRjasJuMG/5y5Zr24innBjDoryvMiqwfMb9TbRHSSrwa6KMcWXo
XyHHtYfH2NKY3G30QloGklqshUsKkxBujlQCgMTqleg1M5XsRz85zQhs/dBS7OyYUeVtT9UTYVUo
XIFf8sZ6biTZHXI2JXTmqD8voF6AsGq05jlG3yWefyYBvfDGPvAtu4PLpwd6YD+LmETmIWPWg0So
bDI2iRuhqw46NTHYpBaw7pAs8jSZWGNce0OGEcu8EPr0aQdKA5YkWQuMI/IAZUvzrXmu9gEDLgD2
f/1LfHdiaGYhyU8QzeAAaMLQQE0+OkJ5ilCqf/yFuseqVdrpC5RfzSSJh+Ru5Gi7iIWXSoC5QvhL
dXoCPWN1G8+nT2c17zGwtBJ4nuA7DVN69g4sJhwRCuvGYnLhup1OixsQRiH51tGBT+UANO1yB6e7
jegRTH044IGrSHIEvY2ZguOyiiKMo9AXA26D1DvJtCupktR8tk90uZmaMGbJSnRJo+BJr1cFp/2E
zc3lMyQx2SDzxAhxc9u+GhGAoNLVQdsbL8mUIdWIgoxmVrYKo0PCVJ5GBTEIQpyPuHHM684VRrI1
rfnXmgQC8P48RTk1kT0XJQcc1S2hrRbrOTsaSPNS2co81UI7jx7UoW9qyLkleL9q6w0KYUrr2F2H
R8WjhSwBgykwilJeT485GYD8AjygJSiU3YvjmMTF9DYWKxFwluenKbZ6sU8x8oivaR06y5dmHEj1
X8sGZbEd08G9C50g3PswULNoft/XCSX6pfrmt/j2VF4NtzblCbaSvREL9mGsbOP1uMdGs/JZL3uK
mqGqzf+rxeer3UiSk1PLrKJ6SWm6JmCKiKPmJlritaLCo3y4Pct7On6JNWyWktXeppUQESRfh4+9
wPVuugBb5Pbh1L2wrncQPehTrirHzauwVXcxBXKxnoeQjpKUL7HZZKiYcect1tmHoIMqzK4oPmi4
tdyRhk6Bwav4ajoRea9h6dlqjFwS0h9XSTfAPQh60KQR/QnnEPhqowEjaQQsyUoLdIbJpgq2GIqm
dA8MMVAzBHIm+D7wgvbqxoDYt3Hz3Me6zVG5XW8vv4es1c3X0adHlFE8tCqKU26bIF+FH9bvAaHx
EUso32qAiDNASu8Qb5AjJ8I/Y9H3j8tLXzxgDIhYeawPVmN2VlrP0ILg+BTtmf5y8PM7tX/SwDIm
QLe0Po18Izs1iCCtlqD/2zXLE7aUcNZ29QRiJOdPYjtnt0Rd64ClPpTrrtIsOofLDD6LFu7NK3Nm
LjEbZVtzAflqI/9s9KQyKAlibO5ytOApmKt2WdupHCDBJscEqfhJZAh0YbKvOpxfDa2Ex/q0L8ho
CJ5/8D45H7R2rQy9mSMsqYrxxsoplT2HiPAL0iIxqICJLpFaUrLyjBnsoJVVdPipKgGYK3gg91VK
ZZ8zCtyqMUkMXqrCMtPnjn9N6Kv3nsCQQBu19d8Hccc3ZgCmLU6tOV+vtUSSfXDDUo/ZkACDWPSc
fCSbMvVKa4+a+LT+OqSIjk+SbldQ+5N/O78frcqCpmVDBdhnhi9r8irimhh9pVg3n1n+afdenQS4
UOZDbJiT1rQrsYNH3pAYp3TjYHXBrPk0DYd+JjCzBlcqEAla3EIdfunaAE5vmrIctQAB493cJUKk
SildSg8kWGIiDYN87MgfgfquRBndyjoMGP34kLNkokNjQuLUYmiv6WGG5dlsOAmYzQ36QUV8E5fT
O1SD3RDHN/pkpVx2QbqGl+N0TRR9bXdNrvQLFUN5yUwIuMSpNIIcSPCXj4MsRJekNazvf7cQR23o
7PkuKqV1RiNL0WeWHs9OCZJOqlwMn0UW9iRffJJ8YXCWxWlI3HjM01ZZGdvG4Dwd5pN+F4X2VkEb
3Ey1LgGGGWVVXRoAiEhNugTuUZumjMly6hlekRMp8p1aelmr1me8fcdB9TK5LbF61ovmfA2RJLOL
1wY8kcfhqzFhsTnlvjkKjZQyHZ3Yy0ahhgPjUbJNENcuqQzilYqIoyyXjg/anneLUFuILwjbPdpx
M/qMagZucjAnoybFaZjWL9P1kLSdSZm0xfNlwcQZtz1RI+qxFhCKKgQurX1slWkxAt4IZlbU6Jbw
N3mqYq1TtRT3XOEq7O6ilgIRI/CW79QBM6K0sF318qcgOwEkVGHn4xtV4IwAGU902jlIEfElJukF
aZIhd46j9lmlbrKtu4v3+jz4Kx8XkHfg6vPvx0ORz4/PpXEAOlIaB+j8++ZVOAj90iFOcQbA4uOO
Qr6teeZd1Hc16vWhNQG8kxkVdSyIM9BaHBU/YR4tWUz7iGSLFt6JV/XNG/bayuj6Q0z/LIGue9kC
uO8P/zW1V0b5GC1I7+KgfUjKUgM/ZyKsT2ThqyN5/tuzluYK7MPnoZ3W4F8kULrXa2mobGR5iJAb
eZZ3+UKswcI1IeF7Ksl43+ybsW4rI1AI/j52ZTecxn1liW1wpk6gUNahnqtIERO1xGyScYnu8FCz
NM6snngObBrS3VoKMZw1ulNpNjI+xytppWRAL833WiSie+XzU3iNmb5dfWYDBgEXnV6hGwkCRB05
PlkkJfSRZV/Q0ZhBPlIkgqIGlWAtAFbodPFtjkX4pTsDYFVnZDLXNrrgloRfDbyYZfJYBffDWcz5
0MCWtZh2fOERsQPYBgC6jcuX3IgeP9e2ZHel6V9ACNKIvper7fvnq6x0zJIdnAx8eKdxXMJyMEcY
nsBCU4pnpyJxZzXZ/Zm+3LUoqHAKm9UwLSiQFC62qKm5xXnUvT/fMdCZWAysaVr6hhTzVoaXHO/6
C4/PqO4Hp2B6QLXZ1iEgNYhynEkl4psRDl+bJ/nvyb2F2KQdE5gt7qJm8PBQcOaivWClCCZgt8Zr
LBwFjjznn3MTVeJl4HITCXvGeyl+pqyqdT4RYmEUF7eKJ3ipUIDpSVIvZECpIuX+zLQ8UOWa1EWO
7Kk5vQtFz+kco+WnIkq0SdT9mdlVcaf0CEeAmP3zoTBt6QWR3OevBBYf3PRWODs4JAl/cmr5RP5d
CMpe/CqB42YrPA2YDLFP3Uny4zzXpkVL7F452HNM6VYu8vUjty8CTgimBCntbpginXeH7xsDz6It
Ka5kS0sVsPAKpxEDs/2clxdqqDBRahHPTW/JUWiR/jU3tCSvi1g1IDGsOfFvK4bnJs9hg/u5Waop
2D4wb7vDFoEIrJmk/xfJ+QJiIgu045VtumNdIpvvd1s5kmYM/BxFgZHvdhzbkWJZC0dcB1qgdsj8
nCs8vBL1ZPnQGp0V3Y13SnIrU3kMR9MmC0UqZTFEAG8/MFL3AyKNmSXB9Wr8MrblouC+PjP86Pmv
ess9lDIiaum5M2o+M9k6PdYROaRBl8w/gxqQoaz/rOTusQqiCbp45tVX+5WRCkWlWTjsCp4H++nm
2mjbnES43I1TvQvmUcNRZh7hxlFEtLhIYsLx4rtQIp+qEDJpSj4Cr3vlXEv3rgImTWYULzw1yG21
vSzgkVdk2AAEtKgtd29CjvnfgCZ/od7phA2dHTFGxm2TIPnv4BJ6ppcHgmbVdr77hWt2XlJpIbQf
QPAT0iDcFu7mYnrliBxoP+dOQlAB/aSRDECQyHT1FOufJbkenamvcNzxurmMzLKhK9uPaCmWUWkm
3gXWF09uosvZhE4Cih8KnfXHrtm3ZH4v8iwVAXZGYJ+mKrRpdFA9SQMFPcXWJtQEospmeSoQh0R1
GQrGjq0yIgQVcTOiV53ReF5WvR3pBk17xsFRW3nESPFq70ASQzuuBGp3bs1kIrEbPLKK0m3+IY1e
OO3t08i5YDaWKCaS6saemc2+A82a3TXjvZjjGh016bwDskDjEgUCqM7VvyZ7TaM51m9TsKscBWzm
vNXcnOnBMgXxanVv51ujJMXP97FIvyB70wPsXoJQBrSo6BClUwmH1s7vLKZjaXMv6JC5JQ6aUNEO
kDjMobb000QaQ3kIuicEd5Du/t3bwk5G3UqpG+BRHlFNKfG0xPUzyL0NcQFJOH4bc/xbWAgpR2DB
FszBBnHFbIO0/AGu0DKgyisLSaz42Oa3VJ1kE0K5WzutKKBaZGpj222k1ku5vSG7LYN4AcOpWAKn
Ha7PH9Zev/ZyvfOWm/uAatYNCzdCERtw4vu5LPq7f2MNyex5CE0ZfCr+PM4ZC+1RcwmMYrtPs6+d
F3Sv5DPJ6hrjB7Kezen7lKsacOldtgztqY7GJc/hGoHslhyZmz5zyn2djW7TB3Jl0ZzibmcB5GLQ
PjY75WmUjp61nQTK8cdAftDd5JTrB2wMvCsaTlV6LBy4ZtkQ5DvIZrKZFeU81zWmXIlKuj1DDCAx
kpoIQ0N5Y2AmeGRBu68/umZJGmR70v/cAgNCs4POtjiHdD+Woff636rz2TVkZ5/svq3TQGKPq9v4
dbodB2Up60fhzYo4U5IViq/O/aOCf38WF/LhGKsEIxnTuJGgcNvV4ev39pqB5vo1TNcBRbhIIMaJ
ije/7E2g6/FhmCEEgjF26Tncb1yK3ahEY7fSvdhM4qiK6ytIotG9xvorR3frtZAPd5vzaRBEB2A7
QU+pMG1NJF7jbexY3b0R5nLEnto4il5OHLYNoXMEe/NjRcSav7PGnB66Cq4MjPLQT/Zn/WGg0Sax
RJAuxX3PBPKLLptCvSmi9I2Qq3qoJn5v4Sj4EyC8qiV8Te+fZ4xBc2VjfIlbva9/2sinq6ZN4AaW
Svg1Sc+F23Miws2x+KwLOUa7gepPFuw/509Y4AKIGJiOhdkizRUC48tBt4yHdyg0NIQwSsGEsPZu
84wbA95YgkpMfr8yi0y+aPSBeBtE/8JeUz+KufvUjmq3jQa2ZReZFTYx+WEQYdZEI1AQO4K0r5/M
htMw+pOgy7yrq4AC/EZQWyWAtUNqIun+4avadX7wWiN7MnNcZtux/lu+7hXp+kTYz3l0pSORDGCa
pTit4oyWXi/3s90ljoAlOL/53Zkvxp7La9AukJiAji5VgUIKrby71iPZRgpszpaYbAdzivCC0nRJ
4WVuTj1LKCtqXKXvC9AOTmPWIMtd1DgECwPei53Lo/afPL3LTUYNjf6Zq/GKzXvZ00HtpFu4lJ38
yMDFx83xvlFdcAZltJ9XvYZpMOHXOpqpZ1W7MOkjoAKk43YbX1ETp5DZ/sAiUR6Ivs7NL4FG9TY8
o8GvrU/36Mb0i9aBn7pYACr8BLFuNWAvP2514koWmTRn3t84cqVpToY43DDB3pKW4zT8kowTrn4c
d1fwGz0aFumsYgq/ZSIl63dqgReZ+b1I24IQeyMw1JWx+qzubT3QHIAynn7m/jjXcOyrDkX0c3/b
VigY5rTNUlQcWjXRSU9PJ3wBLtxc6v2qG2JrW5nmoydJ2iGfHyxbDZcY51kV6EYgdhpBw4yPvi/D
IBnXwv0/PNrhRYIJGAR4aCaxTqZwiVkMTKxQQMRkacP7nGvHJ15XDcBp3f0b5sy3Rmt8L+c7MlXu
iv8faKdQfx3NIHo7ZkWyS4Nvrkv260S1qEx3hvfMIcOtPC5RcqmS2ikHVYNe1Enw0XWB2Q0F5vBh
Wtw9p017OzXdaxHu+RT59Zi809WVvneqXerNbLdspJPPKdEYWQcy9zJT+AYM7QljWQSFxAkPHpeL
BNsHHE6QUaptL6hekmA48DDy6DiC4u0rhrr6s50FIaQ503wYSmMCjAmrrCvTDUGyBLZ9/Uult+In
muQ1PLKyKoIFDpSgcxef6DulmfDCZ71oxcJ4qFD3TzfPgXm1BLtz3/QvZ4L/hznyOBC0q6zZZ6x5
0wDltnprr5UNu0HqLD2/gj38NlrkEEAtqSE5M6zs6hmMjBHC1Z3b+J6mKLNSx9wVEYYe/BU26leE
Oz8LRyC+zs25cQBT4gnd9wkmaSq3B5WWplgHf7Hz3dfFpf+fxPJI27yUBztD+IT0q5aQrY9BiItO
v3ZyVgZDXoaCw8NmqimmE6q9WTXyDi+IZar3Y/BqBNWTnC/IyzEad+qRXFXT+BGG7VYpm+kv7T/W
zqYrpUxkz36EN9lOWqqAZHoFjutTYIm6+vTiDU8aW8NbajyWGP3LOqEfr494taJzmD5A3OINvBX+
VlNze6NwIkXvntDqz1zPOyKUF9xu7QEfPjd9XYe2Lwdx/8qoIIsQsLcbEERQBkKQxRUxfJbEUfEO
JK8zNZQXuQLsF8efDtd/m6lpM8Etrt4CUnQjLpekuVmJfKId9Y2NP5Qc1ZAE4shhq5QdeEheeQ5Q
HRA7NJKqB1I6gKBKjyRNVAqI3Ky6tRuHz/eQofUw3K9RITSg2rEXnHwfsMs6bkgxe5DySXlYChE0
1PVqplsHcjySeRz3zBeKoyxO/w4VpIIftUUsmsgUHwQbfV1fNK0oqxpelQhil4pUgm/ZzMrmCjSO
rQQQqFJUXrQ9z92MlcTh+nVv87+QoM/uIVvvBZDHPB19VRS/FDOXgGDzr1vR9NFmEOhTxiObA+EB
NXkR+ALy5CoJOkYvHIDquVPu9k1d3rv76awzPA9ajUjmoX5KekYYQKK9LWm3epzsEipYcqnkB3Fi
EFA5MlUn7zG1bsNsyyxXitwqqN9DTF7B3/IpQk00wcTrska/MrmMX3V27ge4Nztx4BNN5SCnjavz
QVjk7z+FeF2ROIEafngllGXFZvwBLFlURgIaifB/pQ29q1Pc0fRSfW8fPgEG094EWpZ0bMKWXI/u
7Mo3D1BZWnTMKTLoVCcLfWEreCAqIhBu/T9RnNBsgZvlMCE6QpaILMeHX6plsU0DllN/yeEQTkuA
IopvbW1EI2ol35LxOP8t1Hmz9vJGTQ4ORHddg7aEDYPwLk734j20scI6TS2RxkPBjwTzIkICom5Z
odCoVwrezYVwABKVnxM/78f+YOnDY7OfNt+J0VjbRueTQog0TDzqF6cKBUxwHTS+W+H9CCE5gb4q
XPjh3U72OrO6u7wesmEh4HvcrktGqDbuIy1Zo0Vvw90BI6VudexeFDikZmGmgHb2NHReCvNokYTc
pY77n/30DA8MVFB7sfBuY8bJqpRSmtneNEjci03T8Om5u3l2lYmC2m8z6UqiXOA5+1fmVcQTC3Ud
4+zk5RIEvpDwf5DB3oEAhUeSj9oIjrEEdq2/YEoUe/5VswQarfE6PpBrcdBTB+RXhWKVWQM0XUee
DQ560UB/aZy6JBz/PrBAWfdxzW39TiYDy8p9T6DfJJLy3X4eQbuLBhMC2nF4wRxFhF6GmtIPP20Z
7s9EUva0OTSyiEHLUvNs7RsakLwYzl/db6eaD+XaDza4JGlCVQ6SIvCtcaUc1Ar9tYHny0ULYnhj
Sh0FkntIh1iuqoyKUg/jaI1KMeqoMhxLCZonE7igyoY/iMXoE85o9iBEkPd0BkBVf8OxuGx2mK18
fuuumbAXND8xUoQ1ESphrIPaciZSWQq8uXSPGWT71QhB4NY0Z85VZ//mFRixOZiWRzX01WJ/JeMQ
O3UYd+AEYtq96R44wcn/Yb6ED1WfVP8oXY/tkvhgvFZIY+MY6EMs2BnosIUaYsX6fdToHFXz2+XJ
bZHByQWjhBOuq8tY88i2UjIDoZOU5zPKXwPDtGMcdJK6iabJP6X9RKL1iIxtCD9VnxHFRYqXNTbl
kXwKvSN+AfKO/Mf3uYVRrsnzUopK3K2Z7AvwtPk1fVfyQq/T3NQXXrZVtHSDOEonOii5Ge8ev+ui
49rSSc66Zb+SOWfkpYrXbP0z2Bmwt5l1m5hI3KqSSAc1eq3qA51rDnq68du7mB7se2tbPGARupKq
w0Uosc17l/4uxpiOOtoYwKFeAQ9qaO3VZkGPVktwlbTgEiP4I/ACYYMURs2xjbDUleLiFFjjJLSM
MIYyj5kGiyT+oBJ3JiTO0yIonSQQEIyAZr8aKNfgladdGujYI3DBmoXgiXKdxTiNvWmlmI+4972W
TNWAOn0q7qc1Treb5c2HMMXrLWRsxrXZ7Iy/V28A4XUDlS7lDKP4H0pRlw4LyNcezphLiA77VTzL
1cnVjUANH3Ryyth/GdjWNZgROtf9aXbHgOa5UIQKUvj5frWg2estfIsRvZt0VBImzfEG12GJkb5V
T34tYjNmdMuRJL0n3VL62TyZF1+W4Js1+zR0aYTDQmBMiEyiTEOiQ44K87COABZBYA654i724ozF
8VH3gvfhpRt8+LhRiEdEl1meq5CpJOrhORpjH1FAlWJpH6knDZiLwV91qMmYSBPh++UhvpnSv0bf
FEdaTHgxjWF7P0ehZdywCT/h3UqJs3sT/B3T9uoI+O4jS2PaNobXj4zeRbhzVjNdlWwkdPQ2A7e2
cRsoLXtRFrRds6qWRhhcHD/JZV0TLmP8HTovXL+zt8yuXcqnGKXNwBX4/5wCQFDeZdXnMtXoKVfH
1b/PeZ5zlUlWIZvZSwEEPGFIpPH8NfxkAo7LOhx3SeumSxg0HHANEwc/VcTvv60pgxz/BXxTuqLB
SEpOsH+XNKQXALXMLmfsJdOIMrIVIIrF8/t5qpVtWSEreMVva3fLUNj4W5SgKsFZkpTdVT9RIpg2
W2B2MzIoVNWuGXCmjcJkYEImZl0cXIyAtw8PspaiV6v5KwjszzAkwfhEPjMkySH3/dcUH89v4nRJ
/EBEY97+Ewu4pkUCxDunmNk2w8TZ+wkSQksAQouQ7Af9ERlRt6kx7wrGu3ZEH1egCWHLZ1IHnhHt
sFZgCQnl94mRbQwO6rmkxtSdPY6sjZXZr1mcepPYFWCqqUmVJ9JYmc/rtpzhi+aCIB+BDOmXQWM/
+ThOltnZNtUhh56QWKV4l44EEUbfbQu0NEmqzepWGElD1GpybbjhWAC7rHXmlSCglSRrwgQ1YzoF
86CbfKH6GJft+ujrjvSnOIx/6y78VvIwWgVNpHoeYKAKfxhj+mBQM6GuT3u56uk6hBOS4G2tAK7Z
WMc1gelc5ZaCoVaHAjL8nageSTSiSbukpYFkoDv2Fhev52QwKAQ4U0j+9ENb0fjlL9o4GsGoTnXy
0DzizKAb1A2BGQINDqGw3sjmFPqOZDGurqy2w+n/uHhL3rEHZoCCkX/bDstYZHgI+nmeYZTDdjPz
Dai3PkIbNfChYxxg+5Gun1y9PLR+JH3iCrFQJRAs4+ujohT10fHHWaWL0hcFc0Ab74rsK91D8VXv
X6O55V3VnRUTdmfvBNkCyW4quC7YvtFgBIuITnie40Ra+h3kFmR3hse3q+xdarPSI96gv3tjXtbS
dvr1zA6cKZ3YhRiJyJF7sIOe892xTWy0/6xxidOVgnGDjIN9/KGhjoj5H/3eWrnHtAs4WYVMKCh3
JGZL+kPmfEwA8eEfYgearZZ8/DT7pVEGZyE6KWe2ewilmS4FIMPJztoHN6Xvm/nsKZr3OgN37pku
z+uy56n/GrxbvuTCBOg/yx2PODOxpMXYdjmYEm61p2AUbCC52ooFTLKoIjXPKICA+F4V1Qkkd/pl
sxGD7Q0mMrHGU+q7T6PpIaQ+tZdn/ZunuHkABaG/vokF0poYH9KRwYhGj4ww8vGW8DKCbI0l3gep
s/xVgfkuDBYtFOclpJynNCcu+AdXLkjIfXuw/BbFwDSvjF494LbIZwa0x/wgIKSRxHPCEam7JEgB
ZR4BDlLjlnr7TARJl47JssPc4LBi773RlpRIK7QJELcf3RGgNvU1oCKoDmFpq0WumlbY/DLR5MP3
+RdHfe6u7epQHZ6LEAFylQ1VRupGHq1zhvX7W4Q4XRRuEKFMW6QfiDDTX3XCIQn4a5GsrDXSGT94
lhv5DJI1SW+lSUwr/d3Jux8wxlnEH5XrduC6XLQFgZZ4iHvEyULEWJPBOC9MIAF9Lk5x52qKG9T9
8OWy4Xawa41fbOLhyz3GiZfyFvEUkbjulB7/oxh5CVlGrgN00wTgwF9VAiu1HEUSHG4AesbMImmJ
nZSdN+ZFH8z6Ob6o193f4WawO/XG7w1oIBXi4qH4e8o8txCe7WCawSv1O4cQ7wvKaVnuMOrhb57a
DhMqrk1ezHFMXbd/WAkZ6xm3BAPYj90Pric/XrNw8FUC+EW46KoAWzfyuK3JhAngId+z47ii4HoZ
ZTcOBbpgps55jF3TNYTdSqIN0aG1UdmDfEW37dlqrQRSCuMifWgGmW8TPASchHl4pDfZE51SV9P1
QQAxH6h6TkdhN3seqiLT0RXglj1Vi3b6c2H/2+8I8xHQYP6aerzCHNWyzmKWZIEeGVW0Z3DoklKJ
7RjBkAOfZFcTs0ljPk5cxA51Lh8PsNobi5DbNa+wACayZ+lb/2o1CKRJnktoiq1uLGDffQ5ZbXvu
LeI2IE0FDN7So30pHJujuTL2XrSZynE8m8w51f3opJK4RG650Pq3jUSPcxhZrJjdoI7lOS7444K8
fcxi4J/NDK+U8gKd5g3XzICTLmWIKlh8KVqgoxf2ENO8AD3PaXWzj8uJxtg3riVeFircCtfQalRb
UJw9EFXKP9+RT2L0Q5sVZQnxeSLlwRjepHa05HCuJUY9mnTSTJYklhiGT5cs35w+M9Z2Qxaarf3M
BzR5mqWf+au9WDcu/+sFX8tBviEWHtsRjxisXPtiNTBLsuVp+nFBEjqyWV4Zlylmxp3tnFNg0MS0
yIzv07Nv1gaI+EnNfcHbzwjilxxTnTZPHiCTgMVweIb5hApqmyKveFy8hBRXBoH4rwedXmHhAeGP
YQIqTUNDSLE+btPHXdaYDBdCoQQUeRZpbvH7bnaaM6a/6ana7eSeB3v0JucauF47xKgpMmYKtV6O
/IklXgpddN9Opfm6ocNIekIdNf6IzuFMTrYykaC0f3K21oYBjdDOyoTCRkRPn3gim7JnM1XeBPVq
gN0s0DyQsOCIsksaKDK3/24FjhOPmBbqHFZQpy581kQRb/DQWqX6Ou/9kwUvk4CprM9OGd57bJRg
hfsaeve4CdN01paVYdJ/S4AWusIUW+Ga1Vvn0lZ7Pxq6pN+B8RaFWLSWAOzsynjYfFtbZNaBsXU9
C/yCLXLAi/i6ymfOIZQtyGsW46GeTGk9NLphg9bjTqrB8XxHSe/KetjFEm1XWqk0jhNXu17c9xop
RWEKZIRj7S0Ic/xqg/nqOBh/b3RGuYgyYtJ4WrLksxlg+3n567ZxXDqCBx/B/gFHFN18tcoC3wC3
Q7i2cODa1UZ0roMHCDXg/bdfycVRrXYrzyCBIOjRqgDbNQ6KQyfzhtwI80xlqM/0357UMUI6rSXT
pcJwWV/cIzLqybdxN1SoWixr2zBuHZZz8v0UqDYsnGOgMoYhAAa5Q7rhQPR1gaLCpznwYFHkOh+j
gDkNfqZBjR5FbPSacBvpo+QsvPQ6RHg1kXmiaoaaA3UjWPYwxZlKerH0ZW2JXO5BB1EIOAOOKzRE
LXBNh7sZBYLt15oiPnIIKpWuP96NCcs29zjRJ2Yj7VXmI9xdsFN3v71WpaQC3TSOCrHOBqSFqPmO
s8Rjrxt2oCijYKePH0eHARcj7UlsGnNLx3bE3r6rdNBgV6joiAZeSEsOpO59XeTw6eeWKhu0wtQk
h+mATvEfDBa/24pHuial30WCU4lr56czZzsMZAo2l0RsMP6hyrbNq8HpxcPuKnim1Dcl3+4mv02z
GtV2ag3j3PwAwNI/CCUEbH0i74zUh/1RpxtvaPF9g5vjFlh2E2cAqswVGSb/1EXclU3oY7v9CazB
9JbrYE9EY7MxKxg/2N5mIJi1ZUcmAFhmgjIr5qbdmqns8E84yifoQeL5rHE5iJz+nhDZk2VdsP51
p7feDN7rcpU+/wbUhccsgNyP3PX/A2ZW5Znll59AUGT7aQ3V2ieNg4xoRJW3+YZDUIG3kUltXbAo
jkyBOLlOFpJOD26YquBrIjyaGHcU8CUQdURMxPUdvOrUnz8F4COjUIQ3l8HUsxRJ9QfXh6EjO4eB
aZ+eFsdsbKZPQ1abA/yUYGJlL1mSX1x56yJGB/grM/CvqD3t1/C9Gplo0Ystro/Vu3hQKD90jPVr
fb6CO/mkGe5cbsGUCFVYajT5QSkG1eYFXBpc2ULPdrDCfrQuu2RnsAAgJncvIL8S1BIQ1xKfLF12
G1z6REYlOKldEQgimaPmXb3wGEcTCsXLX+D2RbxF/X7knWLHpTLrMgToGUYNhXw+yp8f7FlppxRt
vCx2upu5FPQ+rQYowXSURpaC9NsbjJcFgJHXVoVGpKKehwsncjWpV965ULo9PXUH7M8wS9V+x1tj
V3tB7tmvakT9Te9DhKNfm8uN99u0DDWVjELfW5BQAvF2we4jDI6v1mo1WvT06sjS5FoYEFX92gfI
grktHM0kMXA/yNNpPqQFADJQ7AurFCsmwuebrc/ujZsh5D+3mJMzPL50ylPcbA3bO86YlxRNlHgj
d5jZ5Ti6bYF13FjpgnBufKpXStBRACjA0keJCDuVYdlaFqrs/B3hIhW7jqA0Mw99b+iEJHVes5GO
bClsRJ7nK9Xh+7ZrVwtq559Nw815ii7LZDZXa8P/V36bc1i7K2F1Ip8Dt6Bpp7DSLruz2HyZONMn
69xN2TW/3rNtAsQMhgn/Vhx+fIBH1k27Xcbb0thiEINbxb+WncVV2p7mKqU417bHPBQf3aH9hpbY
hFw4jZcYstYBuGQVQPax7mBhJU8FGJicwvDAlHmMX8ukBEdHtSB4Y1aVpRb5ukn7XIQ4fBuyu5IJ
yaAS+vLFbOxMCYlRPr1tzx/WSPte5lHR3tFTOXnlRbJeKHpemo71Ji05vTL+S6zYn8I5X6fUA7ie
E76YVJXAAX7IWa7/RN9tPGv7zMRupu2jJq28WIOj1U6kx2O6+Z1ldgNT4snZxn0TyQ1MAC3IrPt4
34YayFjm9bDyODua6r5wCc5boDGUoam0rXIOy5304rXDhU3pYU+2BMxsH0kIDw8F/SfJXKwKid3U
fh2XKHZorynXSBK0m1xAAgFC7D+C9s9Vy9/5LOhKixnM7X4315enZQdMnRVuIkUFMmhjgpceVImO
n3xR1/VEbBRqsTOGT9ElbMwEQbDZjohZYMlRxB2DCLdd1e35cjQl+XJlqYByQRrR/a7EqqjCyKFX
4uEqSpOZRvX0zOndtCe4slOIze+Ii/IE1W8EWQ3MPt/uhdl3Ojqg0ikdHNdGuV1ItMnejUGpMXoL
O8a74vaPSk0A1SQZeQRhG4HozS0vY4Vicx6Kb3hxH5EdexZVgSS4QAFTMUIcKAWjgh3tcgZ4R9ix
K/piGOX/pkTpc1Tf/7qhsrXz7HCIpzN2TtodoNEogaJhBCd5QEl3pLqyjEGgNxANyBRwAyTnkAlE
FU9XRKMvQ4LSRwjQiEJSW23yEoY62YuFqHxWGfIaR6yi5TjvutaBWv4evLgbung9VmBqTm7LDK4d
AqZAzDR0T8Tvqjq207nGDCEkP3Eg9i3ZFMt/A3altOzRG+8eKQbkSBNPsk/fvxx1zu5gbhQaq0fD
wvzdLk7eVZJ67QXVIA+lx/SsnF1AWR+cL0DjeqKkrMcB0IvnumTbzZTlK6PBg5vmnj3JFoMnXl0k
3TLG87jmIspN9oqpRoNjqDVq7dmBJ9F0TydDXwdrs4983I+/k5xQzSM4CJ0942amXBGvVxWhCJLm
2zRHxAdkQLochgwfzIo/zXDvoJljLB0GbCDThoQAi9lpscL1u8qu2f43hu3POTZ6GKIPGuFZ7j0h
Z7uaDXha3ZVIaztYFrD2/OpE+ffmCcbyP+s+myWjvQyARDz+Edw8B2qq+ZltiD69+tgTk1KwVGeE
jYanxdnbBYwspw95pVya/2WsfxCcJsf+cz0kvM2CR5BS2mWT7zzfHnoIn9zo7mYke0OCddwNkWPR
/7lYQMSl/fUaynNrnvGGbXScIJWgOXEvZKoK5P3Nv3571dneX44XREp0blQRa0f2SdDerg63Gf8f
0u1udjUm/NUi2pKYjnMVi7gsOCwngVa+nVWOLfzA3A2RrhToy+xNLNBb9PCJADnVp3CPYqXJiwMZ
YTv+tZCwsLLR35EbV8PIQolGLQcKjTopFgGnzGlwuVJKglQfEtswfDZVk0PmNEjvSkkLn9mHdfjh
yxdVwygknsf4jYZPOlrbJwELCwXAECHYUmUzgHhS+S5K9JtEeog92eG2DgVxoklrWHn7ALj9jZPp
CGKHbJZomdoFskbMceUd9fELCas4gT67fk2igMQBSzZP/QkV05nuXul7ip//iRebPV0aXQ2RvJg6
fCjubJjozzK0Y3dQCWDmiUnNRe7XVzQm9zlvDH7cRtCYQk+Pa8Jyl2vflBd3ankM973Ba5C/lrbs
mHz2j/FwlbEvnPQoGB5jspTAAr4s1HspKt3OMpIatWNftGjk1JILkx8jDaT1RuuAq0CY1roFOaKT
q6dOAwjM/48GoHORYvsiFpAVzYTPVkfNFMQZQEFmnEAn9cACjQ6nyrNRimcVnkGt4ANoJ8AS8rtJ
BUOsGITNsP5WMzUnSYAlhdJoXGkBfUjPov8j198l47GsRBe6qEcvUoE0wZ3aD2sBT7vk4/iRMJbk
S+EFpzV+Y5UA4g3wvKBWXFZ7pvkKJfkwme+tlAR22dswUs2jEcgL8zuDugpDKaieP/X7z4LbLokr
LEQ8Z42q86CmeJxbnBwRg2kwPwOSHjb27JnD8KXEzt3571u2K49L2TLVA5n0dWpAHkMdLvhRtjkb
51k4aDqBmNhzef6TyM2iWVsCjVJqXzlt1jpF6gA7v1X1ySJ1gFXj7dGgUCmPpIuRvuZtHh5wn7qg
8CohdZJYfIeejxIJe/HmmnBaOuV40GaZwc1L8wyeMFCU8pGpSgV/xapXhZheZxr+Pvwq0lwtZfFJ
OyerSeZJ+wnSWk6uCA33WETPpGyUJhEmtV4rMcWMlc1XMiyALDkE0N+mcSeR8XBU4YvQv2ypSXPg
fC0iswikBYn9Gk33sok/exX01Q6JMc+dW5gN90bO29q44K0sOxNXz/kWIDE2rnz5eUar8qThe3ZX
D3LPPMIVobgc8liSp03/WsiIh6wX1d6idFhz9QclVxls/C1awAjdKo45lY94q9qZnoLmOdwB09t9
/PdsuWiIrXdtXRqGNQcCv1DQYGub7TykExthPx9lPjtHFB6G0pOuKfKhNZ5tNsuRCGVdnyM1B/qj
VXQD3xnKDAsGHu5wKVOsE898L2dBnwvIOogfRPpybKJMvZvyv36QlGivfTXHpxN7bEDL2YgSpcZ3
cm+f73234k24fOWvR96Hv2DMUX7rovP2nPUjnvYqxiI9dVjhBprQVeEaJ3OcsTt90Fxj7U5q/7d1
nnhGB0EdZfq50al1ERsIL4FjBoBthUK+IIeFxx0fXAy1Y1xpqQPBDUf9AEsYYIm6q8yFyPl/Vnze
mjyKUZsHYA4XQBdTd0ZMSFYtsED2hDUABrnOy0Y7WDpMRxfCo9d/b1u93XKJog+xkjfBYuNizZMz
m10yAd6a+qi3GP+AAzcJ7hmpr7+nlpbRQsTL6SIQRrUHYWKa7UchO4bj6+u0T+dN6v0WhFC2m0IB
XmWAtbUzjFrnIN5K22+IvSzJIn5Y1fVw30sfYGkFSjDG+ubUXoyVrQC6YekaWYqVAgXKkPuEbnPO
mTVVFGuHp8FA93Ph6lsbpNd/8n/PMVit5gJQ9py84AQlVI3URJRlR68RKrqRammwOd3pdNd8ebvD
PIS9h6mV8r/WNoQ+h3MSfM+IZWaHc/ONxffnUMdZOPBaLR358Q9DgV3XhTlgtEG/skQprDzkScK6
uB1rYHAQ4D1pH0yY367682Ug5X4F/Gquy4TaUjBY2zaLN1feznKnmAIbLzS9V5NBsLEfZ11IegLD
SATVRgtP0g7TsrIFAuAMcDSgC41vOgChBSqZWPs6vGPp7O2qVuk1BX34FI6jRhQxmkR4g6O9z9Sh
Gu9RrhECAj3Sj9mGrdSOhKI9T+IYnnFGHsa8t0K9LU5tSUHtI8f0KGFRvVeyxkQwfEW5xbQ/vPCe
kCcVAvYmQYr0xGYHNsv6CKCt+uG7XnuUjj9d+e0Ev9bx1gCQbZEX3y1dIBJg0RCLZt5QFJ1BSAEh
1UxGCK8OTu3bxobfQy1f/GwGhObZ8lRXl8Ul8xpfXrfxDpD5ffgx9SR9ZcL8KHeGE9jFpJo35iJM
rBZDeWwZMS8haiBgxeXQoNrVIXIe7k2i/JVO/83cD+C7qOzZW6x4E6Yj1BuVrG5b6U4og2WL2Rh5
k3bFZikeJCPiV/zt7AuN33TvJCSCoUlKVciAF9Ds5pv9B0xYm1kvDpHr72Or2YdcKMv/7yXV36HH
WsLd7F+bPWMcU2sgRGh0EsRc1MloEosmLDp7szRR58Q2bw6yTS98Bs0qhgL5QybNr7ODbRJJQNVI
kpaJgVNaOceAx6D/EkKTTcXeiy98Tt2e/aT2v6MNOYAtYOaIC/pQFW27TkoPgKKxhsA8v5kn9HbI
ntCSIhHS4gRa/SGcY0EAclh8C5JC5GojbDIR875ATb86iExcY50R717oG9l7QALJyR6yafz4tpBf
TWwHsBYZK+qOvajeeX1SSpfPFmo3bMQ0DSuKDAr2F/Q3JaxkWcoopvovctii8dRSPn+d8GH4a3EN
m/IvVecRjy2UHmdSdV/kXAaLLF/8rK3SSfs0eHSzlIG/N3qilnLB6S2Juj1HmzEGulXDERL1NPaa
k0GTJdIjsn2dVtLhikRORD6e0q7Pwz8cIqhI4ojVK8MBXpjMpdbcNIe8IfetOqO5ulRpBNtPkCOp
czbRxwKwfjaah1QmvFY79Rqzkr+Yw/dSCRln9NBw+reQW7q0ocCV4wxZrjrg4302B7PFSmxzaSkS
DJduyBJSRQxDrClpvdledBfpw1MljZcUjjgyvswqu4Sb4/QyMIHdwM2NzJA3l1VdlB3KxLhK6VhP
Q55DNBTGD6AK7mZ8pMKI1g+bvg4CljdsYHg3UCJ6YVXK560UsfzCRR2Lm9P1PzcLiI1KWDAEQa7C
8/fOQb78LaQMMlYsEn8DtCVcj69VSykD7zO3REI5tRIxNz8m4O4BNho9mk5X7CiU7vWhu2VFFFBC
cRsekwcAma8XbXsDx069hVbiMr/n059YeNdV3K6yMe8GOZTZL6WAXDSkh2BVeTtl2OTOpZg3s28d
nLZISqImHB+XRBv0taok7m26LSck4g4tjZzrXPtbFRC6Oj27G5d2B5Ksup/6bTUHuvs/MZsy0pWk
X8S1e2zISFr9XtYg2La4LFWOc2oYAVeWgPqnB6/KbuUkkB7M0tCnn4Ts21CbZqduTYWyigW0WAFV
mQNX7Fz4oTCcMS07KSz/pXDm85s6cEAagqzQXbJ5HxBdOMXOFjmOgSqKJBW/mhuNTbUe+r22Er8K
6N/MRDMkehnmNIpt7vAmaQ5fVaip39zFdmcui3Y2Qop6+oJ0CWhK1Wd6MI8UGWcxW+Wlu/6/IONR
D2eM+ZiQfTUqCOL47XfmSP8Gtb+aOHH7dV9Wazn00jmoWr37sJpTZoII5+ZfIdJh1wqV5f8vIneU
QnIYobfPb1X6Csfy8AnKAGd7xynsd/FXuaIMCuQGZZ8JB9lealUKqfbUl1ZbppwiOgRkjuleZXH7
2ymTWH2U3QRDEPUdWb9G8+34Bzs7UwEgO+hfXF0YsQMCyposwgPCxRzhoogF3sd0YP6OlNFGyVoh
dFR4h5e9Nxe6CIBpm1kGw+PeuFHfbxO888Gzc4v/xlVaPabHvxdl2sXUqa2VWJdc3hAUpnD1y+kS
TIUcju91lu3+wZS1uPRPBb42/CJv32MrfBThyO6A1S/s6ONM2egTzudsZkNEqdtignF9jzyWeld/
LGgcngiAwtynT+jeDFaB1IHWsP4LQDYhtvDuEqbsdHOtXgXaruYfZ6W6+rR4q0ZcoAYhMVj8iGQH
WAPlDQFY5KqwCCKRGuXrBKut99xPYOsN1GebuyqtPgeJlr/nu0492R80UP4Fi0OOhhQJt7it5qJK
J3Tn0J48zFpQE7Cj2x02PRPzvQu88mhMRVEv2tREULRPjJ7jdkegnNOW3z7dUvqLrjv3NM7AvY6x
K9gDD2BFP53vztpk7746u6NZ/6o2KseBF/d7fgdp3+719o4DeFRrhofv0zpLmNqPvuZxYrSgkum5
TbCME9SF7nL1LAuz0+pn0oMtfVVq2Kbw3b1NvnFGLkBjLGjnRTBNbpVJZoeCpv8tl0yDk3zHIpvA
+Z6TbgtEcsxCjAkbHd1YkwfYVHl+aTa0R9sKs70soEigRwsyy/gLwk/gAkvj58J1WaxYl4PiOzLR
x9Yx5EH3h4dP202YmH/uNwqyfNkAuoOV+iahRs5jGTtWyasY29trBZlt8H8LcBwndNYoDNeJW/xd
TE25N0Wuy1kUr93Q84WlCsNyyXClKueRdtpqqpninLOnxT50DtAq65Rs1FTGgQG6CtT7l7ipjbSD
Rzgoqo62z5B41m8vEioXqyj0sDTwjLaCdmGaAYB293RFn6Vnj3R1HBll6UI4srF9Qi0rm/5r2zpO
0H+DHovUVBTz6BXU/Xzw42wI5ZKd0arcfKivIm+T65UIu6UeVuCIu8FcaXNERtzs9zNvasOml/P4
y0NjBCf+6trnwUgVgURzom9taccqsodPLOP6Uxig4xGFBOMLkCGqwPoTVZ0bkkKcgR++VVILTUBQ
x9zZWp7WyvrJHz4ooNGKO8zR+bfVlXo53EPojRVO4Zan9qWAho2rLo+D/1458+FwxRSv8Hqnq3/E
dMI/g1zlrAHPkrcXfnmg8EiKgoZnQ0uL/zSrg1AcrIiPJz1QqJzOQBt+GmqWymPSJhzt5LVhHmIX
5Guuw0Bo1ID5fCD/UJUhDj+MGBA4GqVVg3gpeovWuy7d3u+fxNtew5BRZ7uR08cDhn4WtBSAxraw
5iSOAtXZZnl2UbKma4D0+67Qyw94nxST2vYt5oqFEfv/Qw0zYHRPM0SmG44KC9plwL2Su91uAaaG
I/GxK5Ad/OyehSd2O8aJ6YICaBFeBI6l2a7eMn9L/KLNDtXEpu8QNwKftrJ1o3ZJAzunKYfy1P54
EvslBLZQvKdd9VTzPXc6sAdQr45OiVspMmih6q/3KoFVIi4uqeBUPQczA4TQU0FytKS//LknMr1r
1F9nBl/cnpCb2mq3x1MkpgjcGpn+Hp3QEF1TGNQrhQucTdWSqPcTlMRaumFfEoFJUMQTwQi9/lpI
vWU9Z7OQ97omWOFPoD6kpeaXpYGFJPfd8bjR+VmM6C6r2b0NSO39bw74nI80Ca6MXE5NUJwLxzZm
REzVWa9h6JhZbqpCUeXKnMmsWO+jYVJQNSfEYa9yonR4ijNaUVRZj6otezEui77+yDA3+6zyn3hA
/CxtM9bu/30n+XLkSUwXVqA5ecAOGnRoGM2Kk8gEe+UY5cyp6NqCOyKy97XGSuJC7R4U4P1WfUTD
vXrMyW00RvcGGLihRQ5CrrLqiaPplqMvQcq21w6GuBWwiisJCk80yBCurxBr34fWmF3NtXZlkf4y
hBD7sMAQMfnVuHPMiJAFGvOuL6C6Qc964nGw5qSKiQ5ABCR+aK8Cgeht4dXZMJrkRoST++qpSIC5
gmLQDdS6nqWjG4NdprEM/IheIX80r2qB0sKu4xsuhnBKpJxPkIy79APQoEQOfZ/V7KSA9yuqlyok
tZtXbUbupNUPKpIclGpQ42Va4xaQdnhjrF730FeqUY97V4WztCk/A3AFgFkLNiz0yrTdJ+mEYSln
Jf5wi3hIVjGEvilaWFXXikGZGwM97vDRnvNW8IW0CjfwesKEfGKbEOcG9CuC1gmtNXQ25/1wF/9e
bOTt/maAxs/MFDAWRCqJ5jw7tS3A8cOjtJIF1VtgryTz6kJz/dhIQV896fq3Koh0Pzcv2teU3tTk
ZDX2DPVAFYW+U2AYkzYaMqqWivgmL1R85eOMXuBdGEwx9smNgNhpbet/AJ2pi7sDELRCKQDfsqRn
J4r0LrORC00NCpmLphS4Or1x3yGL7mZzPfJCFNsytO4bjQBN+nbIVOBXLJ8KCxtaL6O8hJvSqf1/
u+w/LWb0QQiuNFvh76qgS8cnhkRvRIYj4OgfYDxwtarA9LQQaWfO4Xgc4iftosrpGU04k6FIcp7O
41M4KQc8CUq6DD4iwM6hhDY2V+w+QJFcxITPiIF116QoOgmnOeefF5gWtmp/LM9FOTK4NEJQ9iEs
Ozesnkxe4WUsiyTM4/wBayR2gsjaYfIaeXjAIICw8PQVoOP2CR4uQIuDYaYRl7C29W91k3/sHDEU
w65b6meEXb9AGnPLnRLj+n3U/pamJTUZenEIbQnxraOMGimRACKLblJrWxOQIeNAL5YD9SV4ZVv4
L4Ct+J2Afbd4UJXzH/mkyqfDzFrujK5UwK6R1xRSx/wkKJdRABiP6OO4YCUFYjumJD6pMIPf3DjW
hoe+5XwZ1NPZPaYjVObSPfH4BZ1QopNb0+wW+sm46am2BSYlkIX2USNN3SbLju+XRDnQF4SgdGwC
+XtqooU+ff5oPn7iyruTsI71MaMlEQyGRrjsSSTnUIgzLgKyGlfVcncWeQUGFn2drEUx8UyafMTR
UTQZ8ZTr7K4KdpjjiWT1SoIxZYKzD6/affs8KUb13+SZuA7xiUwbjVOOPZOeND4K+vHe2ESsGwAl
/PAKFD4x5en0fFcatTDvPpa+Wapccbv0AR1iD2xxPHfgyu/fzg4z327ISTc98GSD+1zArCO75izw
Y8ZRSV4xusLvAaLCdmKBEKcjZ63WDvQ4wlCjguCJqCTsHsOpZG+qkJTNNVuWWiHeCpHDe+75ic6C
EcQ+GSZp+gYHkCE5CAfgTZQ4ay8NCBXjE3sM2PtyDuN9DqPcxXf7/xDbCvgfUFDJ9p9WZiwl9ack
1PGqi7Fnz9Y8eRFE59mS6khka2eq8uVGC9+PQaTlp6Ab3xgRaatF+cjGmH1HNV6SoKsLAvExZkYU
MFankWFFlPjf50asZSRGHX+2IXl3Dl155kt7dztmOlEKVjWuV2YSsEcb7t2jw8vu5gupJPrU73iu
LKt+vpvePOz3aq++B7/+4vitsSdCHjipyRGls1h/bcZF2D3WxVUnOzzODik2hQiyjjDQfOXvZSPm
6BFvjnZrMH8RscSbyB2zD36BXQlnmkLIt+hTUvwTP705Pj1Sdiq4PE+R/QRSDEe2Dp/OhRhaZx4c
5d7+XikssY5wqGaAL1VZJ70NdTjxdgtMl3KbwGm/pB7z6JpteNvFSh5tKL+KdI8N3vEfLKpW1ACn
BfHlrXc+xY0aThAnpRjAYzYesEucPChLglZeRHAcF1PreOk26MTDMUOWzv7CZSGQuBASoIrjOJ3R
O+vFK0mobOPNKLkkZh6C/EZocphHF5bDDUiJhOFpSnvXbi43QQoj6D9gibOG3HILayAACdOLUkcT
hbYMInlwlbwigDmEM2ZocsV0qc3+yfr/qCpkUUr5K9ihMjylXW/AZM/7Ytol4yvm3sTKuJT8yaPU
AUzhPgHoE6OkCLsmtYqAAvc71+V+gn419pnsWIW9zxaJYB+fDEo4cjhhC5+sGwgiHY5CGIAGiOkO
igOfEiP3vmEeUU1B3bRFQi2DCXvCKM4GAdMJJb6lOI0vkbkoIcOggf5XrpkX7qaLTFxZYfnlMfWS
+Ydc+I+V/3kII+MxqUTuCuwV7DkhnYc5X8lIxn27Qg+7tFV9Zc/N8h8TPiUfydMxWRJbEXAtnO1o
os3k7cco8VrCqcc5XY5TomiI9E4yxJG8HXKpoIgesQ7YTrlZ/dHQcJdafHXQNad6n3VJm4XHUzVC
hJQ1Ajw8n1QVij3GvoOCGbSsDOlylxb5ikU8r0wYK2k3v3pqQlvzcZiJhOGu6HjoI3afycRnqtrT
CsrLmF1gpQj0CQ7ZzEjH9XGZda69mYmpiGHsSkXS4lRn7iKdpwsey5Z0rE1xkyxtxfdfkF1kUsRz
doBhTfUPKywlxKQ06zZRQNidMIjq+IpZ6FX7OSeAASSGdbAT7K0sJoxh+W9XYTouDLhhBt3s/5tc
vjN/kxZL/M9X2Hd7lT346dRfE45smr6xUqSo11o/AhEuP/K67s6+xZQgeeGCSZKGtNkOqEl0Fywn
cA0NaBZZO67L+Q7vUuKZq7WxnwfSyeR3EmZQ5P92iT++rkFLskUL4aRZUdHbjXSwvO/TeHOzoRgS
USOtBxX3DTf/J+y9TgKmZZW+5soH66O3vJjyVaUVKwn0ABDpr3pw7LyUUTJJvW08UXCjgLvkxiM+
LZfFhQDcsN//RMiRozJ6CzSFlH/0kjwHmXhXts1jX7ULpEglS7x5epe8fmJqZVVDdilp+sMKTEU9
nWIPUXbHXQEOTf+5WFfhtoir11BUWj82EvKBSIRlgZNm7/tRD3W4l6MsFyxnAibHOKcFHcniDNr7
qexGVfJ1ToTlgrsrSk7SoAfkEyejR97ulHIEBQ8qb1NSzRtW6xuHw/6Vqnp+GWqh35xVV4NFSaPQ
0ta3l/CrXtTMZG1dIKkjFCOUI97QqX2YFz3dRXBiqOBW/lsDtl0bf+Ew8TtrRMOLt1xcAoIBEPak
79fMnPiHx8WwPdxLMio0Mz4nSPPVW6tcAyYY2ErEYEFa9hs6zVfrN3yJ7bV2btG4xOA7UnvCi7Pa
YJuPX2wVWTJWGbMLER4hnzBD5Aw6h9bZVKB40s6vjZgBOXA2kBsZLNi2oQnS5NVUpjz674zJDv8w
fyxqecjMxjYwidokc0/oWqaWKjVzDoEJGWK3O8HiOHY1PK4pqx/1ocVPwxy0L4OrUVEPnMsOpTwx
MrktUxKIOKOXycwVCKwsIuwvKcQ5G8bzMGES0tDTEw5GEFQiP9PxkWQV4L90naWLQRqH0TLVaf6F
6KKdY9lB1hai89kevANLn5EA5iWE9Fj1yJD0ih+dzebEfkobx8TMdDhQm+cNMPtCe5TTA3F5CBxY
WVZvusD9E/J0OROzbdFMquy+S8Jg+O0z4WdkeoQ8imvUGT1SUw5M44FyNsS9g00aZbcCSLZoXRoB
pSTGHCIqdjP2NGzyFhiWHoPWORwTUffh6eDKcl4jRXKHJ2Cb73HstshzYOvX4eISAucYTr8jEhQQ
1YQaKklqejW0Ae6wS8Brr0UFN33e1kGJbx3iyq5+TPLUVPakmwJu6w/v0MeMd4QQ+7VRfStBtW4p
5TlEZ1P61LKIFeKpm7RjuTQwUUBwlFoJmdE5doAEwqUbcJFK7C3AYVUQbQJZQDed08Qw4gTSObzG
qr8NiR4RZVCaNkdIowBb5oN4V05Vkzp4Fv4dNL+wJATWfhWeLC3pAC4787nHcIUynSW5E61OfsS0
orxfQ1AC0nCB58hYVqbGKCCVWgQjPnak2bnhqMblTBb5TijfrHx8qg+t8cMlbdLIjauUhsxEeR/A
qlrPXOLlMakCrvq2ik1KpJDJcJhywDhjzmaBQLhnEKJ26riBvbOf2y2GWbQRIEYy1Qmi1FCKbv/j
8a9/CBnVRW1v3UAYbIjckNmE+V1OaxBKlzwLFgWtsrC/OT6dp35pOS+Voe/EJns8m6lrm2MCzL+T
4tdAEK12Z0AoH9UFDnDr6UT1gm9rYvEOBII//u5aHF+XpQZZNYutKBEN7CD/t/+QLiKIIlMkD+lZ
BMXTCLgvJC/Z2PTXPVFTrVCOrnetMBU5NDJ0XpR5AF3XkdiqG2ydMH8i9KifC8da2kEqGnq7WlOq
/BC5D7aKnVKh74CmTQw3aZ1KsLmhk7QvyTl8hrlr/LocBSOV7E7HTsP/V3dy33kznkbfOZWgNH/6
bm1+vfdbK0i+xAyRvwMI7f9KqnPsiVX0be5hIp2k8qJQ0UM66Z1bjY7XEpqZmZSekDgxthuuD59Q
uRxHzuf5uNOc7BkdumC4pMZUS7h2skRuiRxG7QM3rW6yA6zTQNtOn4iU+qcD1WXGxTPHM02IKRlZ
NWM8pe0mNlbA8MESMuULP7ZCFRm0T8aDdTbRXqDAJX9IMlibm3wuTileElYf2BNyT96M5mpodF7u
n1qB+qLYA6jWldzOC1f9Kabbg7YfTitkj+EkeZdoB6gHZJTXrvu8alD0B3zK4dfVV1pqVbqhPNhK
/1TFzZ1j1IwAeQc3awDwJ9Xy37R0TfLiipE893jeLfN8CZhlanKuBMdIlXL3yB05UqT0WMYRUryp
wmPjZ/w3RAVHp4LaCudOjIa5KK9YFWYS/f5Z6OOVSzV03sfsVkkFaZnxDDdW3VVNoXTVdxb7CT+r
eGrrmUu3UP9SG9d4Qw1rmpGulrHfnRDKqG7/Qr3cGb/FL83KRSkVhAYKePlUnZ7GjHcl1NptgwCn
PcAGYwrvU+Wt+HGWnekHgrjcaC1Z/hVPiNCpog80wGuMFoa7qJilZD+v6zsJ6dfL2DnbEJQlH0ZL
JPtDiVkFXiESJ0QAlDn/zguWeOo7Wu5cekF4D3FmQg/DVPtRvA5Kh3ubJaN7rnEqm9qd3H53Yxjl
khSNTR26xptQL0YNiqe0NiZkL3+a6dl7HZqQWPAxVVZcJDZEYvjgb7d2ky4Vx3LH4760y+JlY/EV
inp0iTWM5h0u9d+7AlZUiZh8UziRlMhqD2LW419ofueQj3PuW1Tl5ZdCG/peOOz3DunhB5INSgGb
egbFmxBTEDWf8S9havRNatnV8EsNFxiH0rX5kqzJEaiJKKsNpd+zV/oKsSJllYXZKm4JAMC/5c5G
PdRC8V6Q7lG2ACVtXyjjlDl1Ikk8wb3T4YWpaYR8NcZt1EUeNxS0SlDxUO9HFcmFBSyCS6Jnfh3I
R0EyOPqoqma+ojJZSLzGbB2hzIo5JiS7aQFAdDsdlT1nQp8tvh5w1WCIoo0zeF2NhMB9pNiSQD0p
MiHZW1bnx78TTgXgzcNWDAdHvn4Bb7T7v88zRtWum2vAW8lpPuVWWW2dFfw/WH3kDj3Z7qOt0gZg
Lnl9uk352jFhSCE0GMY8hVAY1VTxswRTrlyGhzfMb1eQki82gJiUT2ri1+vdSRZsLSuhhZQ2kDBk
jJ3oGnEWZxZ1aERYaOvJhBJc1PYEbImYDrDLF5Lb+pQ9CFzjcde1bojPktxMcZ0rhwiao7ZLVJwA
+ec+DCkVeFl7H9r23BcHVMHmX0dqfZ4ZdQEJLTyC086LxGNEIuxs4FUKGh3EU744txvU+mrfHoP9
XdbiscwgY3TC30I7VIVOsR3IbqIlFPBKd6JFAehkAdNuP0npVnM7J4nRJShnwWl3dtjxpqAV7FtP
APMh4wZQrh48mrMdUhxPiZFym3iCm4UQ1NqVlVeoaftrsCJTkdV9dAMSzz20YiWGi5s1SpmdTi8D
eUk4sJuMOJ0MRG9mv+fHSbaiou6JNXwvfiBjDh6cLd1y7LnKte2mAlWmqV/ABsNlRD4F1VzLPyvf
myVgrLO3pLc9HeI+CnimjrIKsJFwXnz2vE/kFMWj8OFZ8E5a3qjswnXl+khk1CfwoDtocUO4blgB
VioqgVLD7aGOca6sEpw6bp9F/F3kBEvXIpo9iQAZlWYNccq7P3Ocyix/IQWb9Jf4vPJK9gtpAMkj
yej8oX2mgCuMPhY8kdh8zLPmn8C9N5cQe+NMPrcE9CHyYF+zIZGhKSyo5XPDCekTvsWLoOsjY2If
Rk8VwZ+YnWVmibIRSnYwOH43hRmpJ5+WP/hp8FLcvNIsm+jLDvjsCKhF2Iy5kcQZk9/hUnS4V4b1
US0Z8Ml0b+oqMet2Iqx5DEsVQK0ufRYnBnDEtwHAJaxCVOJYgpEgkYXSfAO00JvEHAlplBGop2F8
z+o7YXR6SjjekwOOy0x/j6P4rqt68FlTi76QeMYRSvFFgvxRHdRij1uDyICyD+doBCUXE9MFQzQL
lATIVURPR8YbYqQXweOwQ+21IjqbxXYBm5zZsd/gerOpHjCxsUDxzVX41WX3Nuo4sAEAzvbjDfGw
FoBDHS1TOQYrb6lg45msyqWN3lCLzIobipJ/0IMs2EknNW2TkQeZnMkCWUP46CHBsgvdSjex5kNF
l2XinvN9dugm+UWcwO+2hSJLjJzDnfXMAB//t5OHsVu5iSbyhqam2mz4HS1mx5CTvgvrCrB2SNDB
SmuRADuqMx8FOQdsZVTFGhzzwPp+UXpXhGj+ju2SJWY2cRNty71e2xqit5TcR3macOG8lZdtHOGC
LdJ0kSBfL518I4gfOtW6ju0YrWKV644W1g3MMvjSLwI5v+rhUge12hXRHuB4nZNosszxsODhulMX
0Lu/OuPbG/Qpt7OLrs9hjpEuIYBe9bTC9WSMcTms+3Ym6IiMsq8OA16AXUbMkp0amMMZTlsdciqe
t+MRTCd7RxRGVu9bJLHxbqInYGZ6+1HtC6Sz/xUi/wcLY/uV9DUw0KVYrKd5+DccXxrzmfE91L+v
DhG0H/bV55n1HSCuPM4R5daKel8Bx4pPdKIyWQH2Jf3HxVjsqCO+6yOCWvR2To4m3fQfJ2RCb9bz
lDCNplXAKklCfcFB8JnUN4aYs/0JSYSJyyg2fOG14SjH/u+OjLvkJYbJn+3Cxa0wir6luVkKRs6T
edEbXMIbTienvPKC9khaotdL/PU0hsFJ/apTkfyWV0HAtgp9Sjb6xbJlWzx23dzRxgwVp3HtJpZY
TZ298nUuKKWkTKBDfkiBNbFlU8sW7fubah+DwnAR3SjPTBzXjt6tPpRxYZZ0sB2c+FsIUhjUu1J0
hKvF+CvLo56jBeZqyjIAp1L+PXkxWy1QMd+KpO3G96TcRRpee4t+YEQz/Kqpv4HhX68YdZIUy9i8
9f37qcgtbAl0PdDxhiOHFyaXKIZGXtqAvfFN7KEf75vCOUa3JjBml2f7amUEu30BbAclfy3NXcfm
RgeM3h9KjyByJTtbNvtASn7N6BHxe0WObhHPbq7GzdRvDg5jYQj7ziLJCC8dwHxplAESb3+LAnvJ
8Xsdc9vJlDzP4EpcQsmExAnG5sCYrkyu0XjxOoQ6hx/SmAsAHFWoGuW+awX1j9jOD9hMBSDKrde5
aGee1k07O3LmZoAfvdrFdzgIPNFYvxVxjw6M1Uxikm+mEwZbjiEk0lsnK6X4bKgaqVvLUc+y6epW
25Prfs3d6TKjiKbH8VRxfJmk4uwfzmTfIhp6SZMYNfLFJlUzG6ksJ8nK8r/6qSjsTe/HFC1FW8Xd
VtvqEm5jnEnsVdlPCO3nRbAEItZEwJUbErih1vAd3xLSy67+h/wcPx4OblqXwBS87d5PKqA4hsYM
1vHenJ+WvdlNK7i9aL9Bpxb18UhF3WumJrns7OOjfWedERczxDhzqTPNnnatHNKjlyAsSpt6doEa
cewz7p0PtFvReJg4jCfFQHf9QnJSxXuHHIaVeYSkO00duzeDNTOrCBpXNFz6m/KkbCj+GzFgWhPG
etJSR8KSdW8oJCqPxgzrHgD1mapXv9/E2qfLT48KrOtKZM9AKmiuchXkoCxYaQk15KWgFBgD2MAh
JpjaMaNv6dBHnUeRd5fKumbzaOdHYP+ORCBOpgXIgKUMmoLi0nAcF/tVQoio55Lk2h3iuryrYprE
ryn+1BRbZ5i5qu4og1BOkDuCz9FSrrMqLc+LgyotHgo6bXKHyCqn+edlqAw1ptZS+7to6mV+KwIr
X7JpmEaN/hXK8fYmpl042kQ4ITfqb4k0AHCc29jqmwgwVcQErHiQhpYKgDgLiHaKBnXZpxqQbr05
hcO6IMeMwaQAwaSh2kt5z+zqGUL66f4HL+ZUGL+IJyLEf9uTRkRjR9GuLedy5ARRRRJqRTcBFC4Q
fH0SNF7DrHSGsEosLPTwbvlq0GTN5223pPybtpV1GHzoWHHVCNLA0h94dtV1VdjHPC1kkwECl+T4
63KZRb1AEnMz1LhMr2S3aQp2M6BtB+lyoJgEbuYuFnqfFBy0r4lrDT3SQ9PCfANohGG3eHc3LvMD
B48gfHzU2nl8Amkq+pkiZAIAY2307WaXCnN4SDK07LXX6iYKtAX9fB5nPuv+sjJnVN+2AQdI1NjP
gN2NDJhSeUHksVBuDi81B2aeytW6tktSZ4Jy+yqTWcWDlRH7L3Gq6ovNx5sDHpcGMlpZZB365KTt
VWgMD99AWHmybmP4If21rV45JL4NJWAIoI2q1XzxE5pDvcIbqM6XQJvbJNtfyogJGHh+mfbiJfoU
7Si2Wj+0fur1fe2yi1gwx48HvWmrixpIciD+gHa1PGIKhMUCz+I288aE9KpGUfwgMWWcWp/FCZpB
Ivo4MMUhT5XgCWRSAaAKM4BkdpJwMOqe+xH7yD/Ok7QXlea0Gfu2RBm9tYwmmSIR3pwNoZxDPYGY
e7MxdcoxySHrC0GRZRO3pX13RNaPRDqGa0u65GZrUnbR9qJEpupzJLpa6tpR7GNiEKPiGjOmBovy
r0n/AcIzwxL1sXN2lGbeSkCRMjXE4/ha7vruOwxHaOEWO+UE/sutUoDilU/jtBm2VQq3fY6lcIph
SJSyJy6IZhSNyWLaPNxMqZUeQL/YlPAtb1NbhulTKRsOQ2MRrTTAwWx/ZkdL+CmA/p/YY/FO4pM+
jnr2IsMLl4qbssEtbkB80uiXiiLpe4rvglqYfLX3B4W7RFBRhvpH/QqneWV+J7CL+ypAdL76XjyL
T9HOdi4SzDyzWBws/DRvSCVGvG9IPeSVwWXk97q4vh6r/HghJTKne31qi0gCTDIm/G6Gb80kd5h/
AmtUs1bnwr+fbbvlM0QrygOGY7RKAmF4rHJJMO53Q2VBzaCsjwLnPiRH/TPjbm4i1HyGRpe94JuY
FS5f9XY7lRSF66fcfl7nUGYaCAgnEhHFcwW0hVSs+vTgvpcXN4NexE/YpPF1GuTFQenttly/GGXp
Ol8nxzOy42m1YhvlIpF85+4peqGXiNBUgDMkM9w1pW7yhuDsJOECiUk9lnkzKGe5EMIFrwmympZK
rEJQFexZCTKj6yqTnVMEz8oNMMbmsipmVM1DBnam8JLsi0IR0uCOaMzIMeqWFzi9vYzEYcATqN6B
9+pCH+J32wtF+GkqQs43ee8wn2KOdK+vcbOwJ6q9LTpjGs/3auzoEjnNxOKfr5s53mpXwg3EecNG
HiynmlcsQ0cG13hq3l/dvsRddjHq0g/ZEGJ5hVcpyEiCU4rYcx28HKbSblYysMx4HAAwf4dQkgcW
CngBIGewVwGJDZKIkRWwXoYPEnzRbwurznfcXokPFxsxHnGzVA+pwWF+EqCBlRHGdaN7NsK5VQVE
I1CDbcdBQy+15CWYnxaXPvcLBAZhhNSmqSxko43gtOkHx7YloW+nc2nYQ/MtZ+BEVukU5LOMeKnz
Yw+GGU9b2xavvy5UvJKCmvFHyQpYDD2eb6uNXzTLpVAMHPpJ4F5SL2bltPAaq/GYSHLT/T3AiB8T
JLRrl1Nud0HchBoeOyQ1gtauqVrHVoYIPoxLyBP9YNqXG/mVrJTxNXaxIh/QKFBddL7/uyz28O/O
Q09XDwI2BcW/Ff07x9IITOD6Dyb4SKC2mu2fvJDZd0nD56IdqmT9XStGtYmZYwfp+BqJphivZYeN
jwPpKHsS17rPJm4v3zTeWb6CoZ3ABiP2GK702trndr+CvoQYQ3JtCTaTvbyUyJHjhzVAXgiHsLbE
q0fsXAemZpbY2rI8tlWhTFfsb+M7XLIfPljVMd9sJ4C7UPZBOAuM9ufwJeouDpz5TcnHdpHOZMJi
0Y5Wy/9di/EpRGGIpiVNqi1G97+6rkHP19RUQmVtAYzNvPISfOe6M4F1wbXC5ah2HkEPi1IXnpUU
NmhDhWDCyr8aaFdGfqMuSngGrayUIRp9xvMRHJibSD6ZacFmGb7P3hILrcCuJhblgfNXAnftoaLX
QZK3gcnVzMngcC7RG4iexpK61bzrvOWMPNc+Fdvy0hAmNz9ndCjmlPaVhB8IjzHFHy5MLarMQJBd
F4kpHeGudQOqiFBnylZ9vI0hTnts//YVBJps4hjHvgNb4gttC4yVVSm4OXK5Bjq1dxDb9Pok4/Qs
g6BodHYNkEOEh/MIX4z4q6O4eM3KBXtOKFsjibBFIQ20Asz2KmRCtQB6WpRb5KJC86c1LptO7UhW
Xr6vIrS698zG9zvAoN2xmxMeD7Z1l102UeMDcuFu9Q5+6jZTf7EU+VYLz/LtdQxgyV88KRIgo95z
z0mwmy48u2lIDXlwzpvuqh8v4sLZbclmOam6YVAH8ZP53k51CFGA2DwcLpgyMq89aVfqS/+Bi+hE
Q3Tv8/fXMS8akrQyi2nlEXkWIiUjXJEjv3RR3BzAzyTsuy7XSG5Gf53mDcZpXk9h8xxTHSUXbTR1
zfol1l38tiE+bRs5TU0CKgRS5LNmZqlLbjwuMXfFqYGqCrk0EktSucfaNC7SD7tFogDGE5GE7BRO
IU0gVzNCRjV11qadR9/DUkZ4PvZwVrcY8spfgE3ws4lwNFMvvKtgu3NfO5PaJ9I+e0GOF71cJupt
GgILRvUR3yv1ZLDXjMphEwz19Z4nEoLm9BHS3eEou43V/N1I9bifOfDO82+e2Wi1KugsCvcU86m8
rNpyhU203qv2AfSYaAhnk1q/6I7A7t1aldB9RtpCAeRuRCe0DHxJjq2hC/eMXk6nAJIr9a4XsE5J
+ccYtX+jn4xgZLAQ+N1/odZ22IvmRXfKVaNIu8fCups2VBzeognpNuDiHtrezBiLjXSgLrNbqA6A
ziVxZK7mwUqfyl0ANHKrGu2goaFdTYdpkp0JOr/+9bOI55H/413eDhsBfl50jqIk8yFUJrTh2hRr
LG37Rla1GPBnVrDruhxHuJrdLLmJNndBLFcfMXEt5I7NnFrh8djOnsI35qtZ477fYNULLT+7IzQr
YZzuC9Hj/uE8tOD0Fm9ICKHjPGqIGGZxG+X/NaysGKyr98TmKx+Gi9ZIFCZLQLADRpK01B0hJEYY
T6TSLasnXG86rUhvtxXEchi5CyQMN5WZBrbbRq2bnFCYLAlcQaFXXYjYfPUeTVuRL2lPFocFvRvq
1frP5vFoeMpeTg2LzoH2HOzGq6JFmsKFj1WwXVvLK2XRhnxr2Q6WVYyfnEio3QBu89Cz4Szimijd
CJe1Oe7skGCfJdyX4sv+ugGjv64u1RIdKZmUorS4i3JdDFRVJC141WNRtMbBwmJq5QBw8DpsbXYo
ftA/43Oa8vD79yNPwk9i7I0HlnqM5XJ0NjBhX1BHVqf86zu60y9xhXZoa4fTLp3U+z1S/uHC44c2
JSSlmKZck1JZSjoEUKhkeT9x+bswMkOTU2B2eIdbZBFi4yAz2vvpyir0DrobydjnMXndSFayDofs
YUzyoLh+4S9T5e5HMzG3sBFTImc4AMw4WJI0yp66FfTDn/K99KEaqMpFwC/q5xXlyPathXYouaFj
69BqKX0yYfftpBkcJkP9yZ+2C7ovRipObYBEDpqtDEqqZUiaVly+Tpf6VEWsIBNeVocfRdLtecvZ
Nq9+Iuvei81aruc1IOjP4DQC1vXso9bnCOF3cyID50V3abezEHYQuv0tYRwFd0583usm37OebAY+
FQgfw3BI5GiTbJ/xC6ARDxI5TDtO5UVywvSDw+evS3O4m/nwgQ4MRcfQJVSo5PF6hovItYXK5aGj
on/xlcPAjxwoLMp3mDldgSg1baAo2gwqR9bJFlILEdNfLf9TlYhizKVxzZGRLV+Ho+lOKhOHBJ/K
MHjhzwdgrpRecvvsJk30kY+Gtnv9XME0MUopw+OMzoQ4GBt4peKpciC7CQeuVbM/K1alVCUmkSFI
6ZYiCAc1zb0gcftS3R9dRYNmMBQtu3VZJh2VUGmfh8p0tnrH9HCYS14lyb3653CGuAfST++9umlM
0CQZsSe5KJCeIbUK1AIUBvL6Ac+R4aUnLMOUoNkArfmz3PaXsmcaEx8Jep/IcVvqbLcKWmOQOC4o
/+L8FBdBLOWwdcnQHLBtpeFrlzjVI1hjAOj4ZaKGNPgk8gyE2qLtbsM+u2GTuCcXxjbycfqHhQ9w
tr4aD0qzyqVa7SGpMEdUBGD//QfCTmD92XXuLMhsgFLkPIpuYS8Ki5/pbnBX5llHGkpaNqDYuFyP
fT3ZVrdqxlzam4HZdajo1SIvs2Su9TYsECsWkjOHkntZ3/d8jTX4aXHOsQXQdCax27DDU30u/s/a
qMIHoXEv6NnkDADu9kQXJs/gZzLjR/8zawhp068CGnWGGWJmBroM+EV/+I2NujouX59yVjPoYABv
6i9CXseNnHzJNm8wxGfFmsJsNqSeKfBtFJ4uVxTdoWVbibwV6pPCni2VgktRsaM8syjQV+wf3sqg
VXd/IvbAWozuMYWviPCHcXzSzKkHb808zsPRERwPGxFzwPI0rCQNCdZjxLWQXj+EWFv+axPCLMo1
es0lwj2B3/1JYPROnqn86pHJJ8caYePNNP3BEK3HOYMF/86DmVZsi0c9POiyn84KHNWHnikLOC4a
o0RwT0GXutCUFlXSZbB59QLYxxyhuLqmY4Mugj+rSubyOSZPCbZz2syeqw/XtAg0K8GAHht0evk9
9sE0TJvPyXLoOEylQMr0eWbAk3XnIXCtzw4yFOMkTZTN2sS+btPQDIjdihOji/FsnYHcLJ0uCZVu
xotYWWEi3srxWqGj7YlSYpLkKrVHI0PJyxooqw3DWKU4n9fD5WrUdtBhVcATyIaOVk3WtfyidLpA
DBU26zHbQ1xJa6kzl+o/kQfmpgAf2w3/V0zgtpEFRt0DJJATAwp1DjQKgNqsjkM0yDDDsOuMUPrT
ebDpOLXXNXAdK/jgZUWBuoYZoLga94mmhwfd8nK6c88cIa3D174jgxQmFzvoYwVJVVtcXOQH6Q9y
x9r7r9sJ3fPncg85mmG09MtGEofbOT0Dfqmjo0S4gHZz51Zk5XMbaGjW2zJdMBFSJJ8mrK4u72Pi
JCJsCEXaFqPMoC1i2zNVLkuhmhXfQs5Da+LUWlrWR1OHjfJjWxRUAmjdgujF3Rr2WZVIltbQwfAl
fV7/HEGKPGIoZjz2imFHo29ICN0Gn569UINBr6+fXsgA5o9uay13hcIGNhx9MU84HXLlIuhYZHO5
hqn6hQqwDf05hl8B4NzJZzUZeRTjbONJ6wZO9/IFNfeCuGUXwqY85pRdcYHB5YwTOpKrimP6naJn
UKwPGmQeZ6YJWzgyuVWyz79dZqtfAUkZP6uKbyqdPeHXAL2EIwdzcFbFAC1/GYrKk6XaIK4JnufY
jQ3eveN52AcXft0EKdmHlgX/kt/aY/98ku8eMwBEWBQYDUb0Ww3CnC26aHSYyfgxwQJJpRr66tdm
K3nLWAlZx7W+fs1Q7N2asnJM5efloPD4RrW2OEsWq92PAhbfoKTHNSvne1AJxrhKRbHHsPoLRWBU
nybbw7fE78WiTH0O8/sgXJbnO33YrNP81kBkdemS5bevzZhxAeNH+nUDQy8z9V9iv1U6Busq2WJw
7Sxv4e/kjEwyT8mys+kBTx44fIZEQRA6UxAHikMea7cXhDZH8OtFJdkgOG1cPiEZB05jLkBv3yUf
t8gxbEEQiuK6EDVEClyEBZf6VNRg/AlPW8gvV12dqRkHUscpnHOuc4fa27Oh5+jAad0nGvHjVt+S
ZChd+t5ofujuTG7nQEnjLgy3JYsRcWT3bTqF4dfB7h8zaJFqWztibFkeCA7rrKT5rYV6em/q2Nm+
h7AWQ9RTkwT1jSQklWTCtuQlzfbTbmLUl3Eryqi/y0cf7q04780GvsfHNqd9QFA3FHnQ45OwqqrS
ThinM2Ubsldf0uSTzkceEETszSSCjmExpOoybV/oR/WlZHpt96K5qxOgzsqYOgqFVGO51SkWS6MC
yTwdNDzktdOAObdUGXSiCWWuWN6+bJdleGXGEGuIdhde076f2IhPalOPfkS4uLIZxgPz4Q4tMiJZ
7QSRYMmUfaBHZIzFK1StEnX9nwp8JLRSF2eBX/l7rP0lNX3VnXsgAg1Rp5Y3Iv7wj3SPZaIBfz1R
TQbT8SNzc1hjJHZZGgfAglMPLwHaSYeQirZ7u23KdM3Lxmrgah9OGDCg8LumBi100zlVNKPTz4QH
BYNgV1JUMazM/jDKIROhayi7bI8zAfXLdiI0kYUoP+HSisjEf8978CT9VpONE+WpMdQYtW6buiM7
71vo3AedtOW/5dfcXF10YzZQl3s47Z7jxeTZmVQL/d8DyE6D/QUHl1s2j07uZWIFFUxg1KrvASdA
Kpr0uje5byaHKMzPPBNJeHso49xbKUVqyGCuVm05yDjflYvlkY+K3khTvlahVA17EisWG9ZoDaE6
aZKdkoWyDZUEzY/ayUcultNyPc/44yP6bes0Xw8Dzd8SeLs0lKHxmSDDCnComugJAwYzD91yo9kz
vXI2oaGqhNtYMGU9yt2yMzxMYB6Vm5ax1Efc+ocNa428GM+CrlvECK9FXI35UfArLZAbT0vXTqgo
apYxvwwTsiaydfFdDuUHZD4+RiUN+L8kN1fy2wRD6IrltZbUMY/VcGKgFBiZRMQ0sAoPXtWC0KW5
rs52uHI0BTjmc2DK4IWT2dSXuUHqiQ08R72QeVgA4JI8YauiPtcE2RpN2H3luMniiSOXmgumG4mv
z5eMrH7pD1JBRj6+aiThQBGEGmkw7DwYXULwxfhpdEURzf9z3+uCAiZFxM+XYkTL+LXL+A1xcbw7
+Ek8AFZCJkZfTbqDxeknCGkk2+rUb/t01bzZiHZVDCkcygKJLk2zyBndqZhMc0WWzUszMLOrpPIc
WI3zvj6S1vefgMUVLg/+gGcPZn9Fh1D34x93dGu+DoTm4m4wW1B1rJGeyyoXacJi253zE0RwdEdl
L/VSQagACcaW7P8PzsSog6T50KR+CG6vTDYlSkKKbsUmSvIJGkD+byng3jIoV4VUl4JiXawabOTn
/7eotOPcnd3kmEfA2403n41fPCR7/N1CHNDQ9TZ+UPAC2vanv6h74UkoZBV13Bie5OSZP8ZBywvZ
3HOP9pdhgnPODgfJorD0m2DIi0ylKt0aHtskJm32kWMmMPHXjZHa0ex3Y/KLqZLII62t7r+MhzrH
Tt5tB9hoDU6ri0bCvZPK1Fl5esVz/5zL8k2aRlLzS+dm6XWdIUme8M4iFrez0xrunf2uEXp2eYXJ
rSaBwAHDPJF77+vTBVYdJgGWjS+et1TOdRE0tf8hI17Y6rkLsnM5LrP0+G7TfKuHwPBjlbaT8TLJ
svmLT1nIuSMl9Ac3X9JUO2b4yVaM12Yogwyq2pwazFGhRvbG4cJMZcJOBQ60xULnOUOzNcMuRCB2
41iioeKRj15USIyiJtxo2fI/mHtIftNhBGzhASA1sxsxQSZrY68udQCauAA8/ekS+RZvO+3mMnyc
9S7eqou/Z82xsw7fqcHBwP0K/psd3zv9n6h6XcOja7gf41vcCoYdoDZcO7nPUV1MWy+QU/vEFwc5
fUVui/+jwMupUUNrO/kgLirFHFEFn5vj1t6+BCl7CM+c/kiIyUWlKr5BKxhwK20akj3aPGNWhdmQ
93VHmSDL/mMJsxz0aATBDN6yX6ZnkuO2yqul89SArv4l8WhywVSkegANXbDOMDfPwynI/WVk33qa
FSJB3vCmz9DSgDyUt4h9Ago4iDoVuGZX+RV3sMvkFEseHQZkD8X0knnFLroFV10PpO0k0cq6mj6Z
EJko3ocHs1K2hRsEd8cCmEz1DEiQVhUCWmOM0uyGV4R6ii8qVmkOBy8r9Yi2gtfBgNo225Rj6jcN
zJpYWjhM4NyM39cVQVgf5/zDgj0ifLoIY7RLl7XoUtIq407Kv/U+HQX4cZXPMP6qfQDA95hVmjEs
FKavtIP9e2/5Er8tCU+KTbUkVu3L6k0DDtFkiwVLRz79fv3LG4xxVpTPnmPXvYpZM400+JKDGUkf
XeC5LDQm2JvEgdPd4rdcMECqOXoyLgy2KK6SyK1NJxyzfoa+MQFFJsa895pMiQ3SjxzSweE+aSuc
kzyWKich7ZzUY/4V7K0j//Jdtihxd7Jb6xO1SB+4eaWU2T1AMlqst6oktcHKBaJKQbsTWDRYr7Eh
Z1BRRepnNmIBnm76LGxuiwlJ8M7WbEQHE5KoGdL/LM3YoXGIonHtLM86NThPo8i/TB2bXmFeJxpT
1qk0nV2b4suFGYGKYVzkY6xXrcrwx2OLB0NWnSWGvMqc2orRhYGSmvbJsK+NLZVaQtSRjXD7aCxj
OOt72OWnQOP5B8wqjiU3iZ3q88dm/oVdhWczYRkvxZ54yyjtkvAXsLdfRejgmVpV1RrJIaBjCrKc
99clhwPcwHfdXpIP8n+wUxmk0urP8qEiS/dI4CM/+ApEeV5u3tMzayebWIq7K4bs/jMpmeWCmtMT
95r1sRxeobX+TupoD6M+TWlhA2cuRD4bmv4eE3hDEVwV5huhsZocNxfVz01mfRemKhSD/YM2r41H
oNsvQOXW+uOI8Kgnr4TI1zxHMcwUabc2WrXo1sC80xo55choi+oCpoq96ydr9sHYk5sXw3/YTSto
2NM3LALXZ7sFTydBETXaGf+qIfZcxPoufAIlqQpkm5AMBhUtlzW/dBIeZphOsEaWs+EtKUk11hEk
0IxN2qstrEAeMG3HOV3h1ibgLvRRVduRyDOjrExJdEPQkSMcXXFW+BgtTkspBeYoTwxfOEhFVlsQ
890k6qSS88pGNfa06odEdZsg0+40JrI7CavG1WfCrAbz+GfKIks0HC/f+G7Jl5EaknycG0GtoP5j
lix8xR48q31dNC18bFaY8ZZGBYvlN+eJqlmQHnUOzNV+a7YJTqfj2U0ebPovC0YYzgYxh3NCgVWi
Nw4IZ1gUnZbmhemcsqTGkeP26ZztoVHMnzWow1D0PlHqL29E6Y/5Bnrf/cltOOFrxnQV3vyTCRFy
9vcwi0IztJOZ3h8i8CwC/FZ910hplHkljGcZpA/3GSb0jDKSnPYNe8CMK6wHzjlVBnhGobT33pgm
hiJmMaWohD0ESzAqIUrtCcP79/IbgQFE4yoCVQ8UyTIlgGlK7EZRKubcvYq16nuHHCjD480BYLCS
/BpF1Kh8/0h42Qt+9jPijBiCn2MfOYK4HefKNTqxK2TTSXZ+spB3XOodyFETnw2newDsAAIN6N5G
GhOeXephRom030R9Ptt5o7+egwCh1CGCGsDY+KL5Yx3jIFhEABAN/NfLLRa3hNiJbQ1DOuEnDUx6
vFZjrpnMCQ4xUr/dEATWT2Sw9ycHItfrzHC/FI5PLnfEfwgIvtguWH5gxMNXI2gthsYMt5UrEYdp
SbKG1Tue7HYq4S1VBz4chKuaAYlATISxA/y8OYFfDtGucY/iNAgGCDcP7eva0i7onYzYOnStSJdv
Y0ev8Tsf8z1NO4gF8f2pSdHFNQqkyRmn+TcZVhFzTLznK0FaLD29G/g/xyhpdIFSFI/R4YUgGK0X
NCN8wYlvMgLT4A7iSRFSSQFKz9IcGlxH/qtO7QIhuP0XPJIu38WoEfj9Zft+jRkr1jFzQ4KGRAcp
awNzYSMhRJ+UzRtLF/DjZMvf9P9qopsLMy2IwPXrFoUm5LqgOMT1+Y+WAhHxKfRffg54fQ7YpfPP
lMIqUWC66YaeRlPU2fctm2nfHIQr3VUjNov3A8RSqzyioraAlsM3cnUmgMWC1v1l4mKrKBL2yAtr
syDOaHxtgEx1NvIagqBlxWy/5MhpsCIPrhbxyP3fufkMXSnEuEx6eL4w0KQzBFfH2i40Yar4ryYV
PiZcR+tQXgzcGyUm6nnldwARnnUNEe0nJRt7lfYt7NAXTm6BGufsgMilXCiVGTkuNlN/OLfUU9tc
E3jEN5Xu/Ud+VHY0VG9QKW0JrizGWvLtpyEt0pk5QMvi74IJbnwOWXV57ze84bSp1/GhYj+5wVgv
VEqRhU0V16/ih/TW+G2a15M5UbuIqf+otZCF27Aulqs1c1WENIYSfzdFCBj9Hj+/Z9G42xFR2sMF
ObIHFOJ8/BHYyfQgrK0m5ypfszXCIGBgromXYw5J4/ERVSzCvF8I7T9AbZOsZwfY1REX1SoV7veo
p55Gbwu5TL51/ODJNHB9nYbh2DXoy85V8yO8hnPPZinvfX9OvQnTaAzPdxZ5/aMYMyUTZzekj/AX
qX50gxcJzcIa4zNgvHAx9h6OTMCOJ4r9WUJZSnL6l8I/KjVxV0dtWyrHVTNiLG9Rit03aGp4+h20
JWfEl7uWUxKi//Yu08SZVIa34JC7lbMpfowbGbQKNM5czS2ZvJLXK0A74deq3JoWM4ic9QUQl3Yn
QVKgVhPQB0WAqAHYtLfn6f6KbKU/XkPCPQ8np73z3HdNFGiQBrsO/Sr7/9bwfri3FXkC92AnIIix
PjEPERJ9WLJDPKgpSfrkucfJIVYq5WgXkpAtFqriHTfCZ4N1NyvmVEaIARu4n5F2N8Z6d+9N9lrf
xgs+uk2ttqGBYl79AvzPaECRCDhhPk8VsFKjt0doKLQFwV06EH9dW6b3vqlA0PFp0l0feIsaXLun
5S8mKNl0efAR/5/Ly60BXT8p8cCN4SJ5yRVXnG8iESSBJtx+NSdaOaJrTmhMYGy0yH6DZAtRLdJ5
muiE5//lb0pmqMnJc/Ofx99zrssGV5hZ54q/pb7Gtr/o75naZoeN3ijThkIuG8xQxraojCeHg/o2
aTR2exuAImy3Wutyd5JFAEWlPnZ8fQl9TZYlSQKdzwMvPBQDDN3Sxxm9sW0Ona6/9R7ZJp3XoXXu
3Eqfgd+fq+ehWUQU6D43KkngS+cGNfZt8JlwyWzHVY63SrZuBmDrDQ4tocCHuFXYXe+Og/Wu37Rr
Pwev90h20wp6Fkeqof9jzZ5C7ym9IyKjDtUtXJw2Yf1PC9v+lFFq15AiO4aiCB/sohCfSX6k/jQP
5vUoxarJE+CQBfD7zZeUqMKKf7MWxFbmh1CnOeX1Drtk4+me/ANDLB5ikQHaGmnJDR57K5EeJxyg
OTiFD6tmtk+8tiCDpeaX7Zg7rJX84bWnAjXUIDnd8gwVHRHKyPXQNvhnC52uPlQqPL1oPCyBLBw1
qVrgkTbEPgsKL8MFHSI44yF7ngCWEgSe7ciXszrXrRUSN8WLDfmNcHhGJWY/mbUV21/fIyp5OMS+
tVN6pjenko1Wo/eo8Ga7deoQnXmrOYYQfgsf0I1SLhikGVsvaSjtfBgd0X8xWrGctkvbP124MCXD
M65p7l2Gk8FwVYuWqLf/2V2rnVsopSiE2NhlSnMMWApVAvvoGl31xS2wrOcmCtO3v0MeJnmhZA3s
XfwLdIKqjZ1k6nGRQBqDABDdYupL57rk5H2TqlBWPWkv0I2BxpVYVV7jK+fmqZVgylq01qVNQ6OG
0Ty7LZBq3i/7hyZndlqbqzA8Zp3xcaIsDEsDavdUv0Rp7J5oveQ/5pMePzLxyK09eAoVAjPY3vhM
YbEg1lQhBeKAQiEYlZTU3heuAXpF7bvKHiZmAUgr1oFow/vdf0cNfJV72ARu2w57d8aAxYKT0O1j
M+SgA7MR94sVMtWNM71G/ughTuMzpq5ACuE5/I5i18DEABPFIJX3C9D7zj1zOlF4aweVoM6YFdX/
+r8FEIg2HFuHuAdTE1qEsPcXhnfVr7ZLZ5QUCUBxTFvq1JRBFZROUcswuE+lr0jfAdKSh+8pj4lQ
oYBM8DwXcH4pyluojlB6X/cGku6HtJSI8NHhDPmqFbxOvDDZdNYzm+/mOX2MMzMXNPTopXSX6hqe
fZd+ph9KmE6h+2oB6sx0iyVXshWeIKPViG6EQp2pjmcSEKjRX1BprizIZcRqowCcYlBYebhtkoVi
dbB4Xnyb7DwIe0D5nRCT4RmPIu01wiuTApX1FHL1nRyit7RS4KSYDn+3ApJMvrJsdJxvvZEqsXc9
GVlrtN/cdu1TEVzAEgDDDxzkX9D8/0YDv9KNs2GdtCkCp98x2+ewweeHbXJYtUYpaSxgscKcjaQo
m/UpBe7OFoqWXCw0Uo0eyG6uE/BHTp5lgrmxi+h0mlaR076sHt9p5bGpburzZZLzQldoSVri+UOe
YN4yuSgAJZPSqigffX91iroc8P7Hb+r4Rv06C/SyMiZGgvLQj5cBCee0h9t18wnGrzu7nydrj5uo
RO8hFBVAIPT7j9pEMwgyjuOUqvus3/eVBGorwRrj2gKAXQknz2fOssBHzEbquNw6a1XiUUyhzo+2
17aYJyQFeLVaSDcl3lTmZCyJEWbb4bdvsB5EGWH7sBNkgI26YuUwE6txrodOLEA1NTh79qRJJx9M
DAdyWdkM3lt9AF2sR5EvyIdNUYsnTMvAHvunF/F/1fsnPJCbTXBu60oDeA3f86hzkSaGTFC3ntbg
KHBZ1IJ/FwwduSCErRkfT+KGMltTZSKALpi/Xz3XKO/YWFFcicRjGh0joIPHznMtkS2Q57DXk4uo
xWCnBo4EGzxyc19piWJmVUB93qB83O1xkOpS+I3pYolb22KstUIsm4os7lkCb7KjMuUqh0sXSD06
GcnBRWIll7XFRz4YK8LoQBR7s/mpQ+LZIvD4CBRTcENjwndwwwMIlaH7TdiQzfdhvb4lDjbv5vm5
CGmNMHD2LnpDo8aCpvGM3T2ZTkRh30FTAw6wqjvQRYc7UIYC8SYRHIFcT8bv3xGA+G2XLawIfG/N
7RUhGsFTFUH/cjs3TOY3mr6sbQszw+rV2W05ZzK8j+Mv4XCvqZmJeimMMHiSEnUXHBP10RRG5Yuf
xpbAzh9Yj/O28tkkIXVSxpbede5lsEli7/4EKMDt/NBTcQBIbZqpCMXUJ7ovRaAtfR0Itou6DYOe
BIcBtAyvNWCZ55wfcJUQG6PlDmAVp1aMi+HDVAxxaWB1/dXypf3wBkv7ncvkRto+HUEVBKEID89m
t5SPUyQQLoLSyaITtgm9Oun3526p8j/yK/rSO437RT8Fo7FzUvlVQxU7WN2G5hneLMPTpvsk/+4i
amw2UCNJTS4Ga19xX+JH0/isYPvxWGWDmcGqSMC7rcy1oc9q5b/FsGkvHgVaDKXgWz8lGQRdmhw/
v7ptaho0M8ZaNd50L2cUVREPv+3iZqGVFrjyEzrbOUUZni78QxE8z4zG6ZnM+IXFpMRv67PKRM4E
gmALBO8WwPA3bTWdnZE5cPhPsuag+Dya5idji8hv6zhJrw/v67r+GJ3uJF3YpK9GEmGaixjOqwBN
BzL9H6OCopRI+JCWdEohUtstb7sMARg+KXbPAoTKMoZNZdpmkRTwxpYHed96gVwq6cCS3mcXUHVb
pWGJ/XTsgTCPCxAnZCL8Gb2TttFhpAIswGaT2d1CsGDOpMGvveORWqISfCL4KEvZehgZa7WZsASy
3FJwAmtV79tm0XITmHuJVKG8QYpVONyrcTr1L830ElGE6J8x7L5GD3a7PBcOvxhsVv4IVC/x1to/
wcgwIAA2wMuM3i9H0YftDcq4o3Pe5KEeU0JCER7LeTvcsAX7MjkUZPdWEFiti2fFi7IfXP1sIOOv
l1Yhn5dcJutI8z/B1iKGCY0Mi9Z/3xUo9qbCKek61xx0vMyJ6gVecq+k6iR9cQl7XUsc74rOtr7l
e8tG4y+Zh6MIr/Ip4Nm1aT5JWbgiWZoEUJnXebtiU0sdPYZQC6TXBYSEO6WrugvOJZ5keJlFnf8b
CFn4hEBEGM95Vr0kHwmNpa5uLkNYtsKhp27IMDVntTLRPOhwqmjxvdIpHZwUTlFTCdP7hZmUL3jt
ObB3MDf+ISR6LBMKhZnUxI6ufLhVN4KHNOxAs0QRBUPe9RXzhtzMGD12w405NHhjf6aguDxtbIZa
RqU9g6320Q0crps9wZUQv4RTVyeS6ntOE3EmgERiwklA+bLAusrly+5T2SIY0pmjCVWN7G8ngXpV
tZMledEUUQ5bfsZ0wuD/Hrt/Wi9oAyrd5BU/f9fuC5qVF+QOFbPJDo+9eWgsC8yUOYEgGzUbNmYj
1QvXoy2WwYNLY4lJi1r9sara0GPieAyCY1yxh+dr2JzcSBSuEOgb0X6mrneN7WGDUqDEk6w/jQjX
zVIgFqKEc0FBHjEmr+ii46Zq5BRHbqOb81AiH6OtUEV37Eg9eOjLVPLMxmEFcqBFwzBYXlAUKGL6
0+YfnLwMA8DeqCvnoILsO7do2IJgUzVJKEhgsNL3w7HrAXPjvWGNHqZtHaN0r0kkO5O26IciH8sf
lgPIJ2Uq6UpBQ0vHux41EIwTt4yKR2NfRoDV9eFFj/dt3YWJIqw2MFryKFqE3LvkzrSH/xCj7MAt
wXRysmfqvKIxGV+W9PZwxzwgoD88ve7ZFR+gJKEOuLJrEPRXiaVL0yma67lJhBbRUvEz27rayfpM
5LE25xGY5xAPz2oRSP1YnTUzvajFOi3P9CbCQdNxBaJLVwBLBG2yk2qbZdaSi62Bu1sRS2LUZuTS
Z5Mx/4A8vUx85FnbumYSP+bEWL5AmlcsJPnuTDgRvmzCXQOLjpcWnTbBbzXKyYfRKdFUqLpBDFTn
eVr0UGN7WhFmotAOKFycTSYo8mtwdUajqDXpGSvW8bFMR1DxfVnDvr0qdwEEDXBF8njuefX5KZmD
wbo7Dd6w4JtP6+7108tHBfOmU3Hfxysnpf2zW9eaqzGx5/uaawK6mkCanJTaQcdRxrbfqmD68Um9
NpRi+REMtjZks4u2bYkkgT4kKu4FySc5faVGUKXBjRA9JCGkOABqueVaNYURh+DsvNYczC/BxIfv
HB8Ifn0FJetDt2bi0SQTPe4YubVxEtn9ROA+A/LmtNhjKs3Mka+7TZbx6EcNSHDNnPdxuzf/MGY1
Q4y37GkJw/o8uqA6XZ92uPp3g7VDwA6J95cCS58jSQdeDntk7tYo09KAWk0bQFJLsoTmoopBxvkm
KJmukH9qRozsp2iPcqMvYCrEq7nuekR9Qmk9tn7DeJct8fMRXggdBmCSvYsYte8FTJAvIw5JqTYZ
7dzIg7mjAF1w1ryJIPnijy7UhIGfueyiAqNRqdEdJap7OhepjFto4/Qiefv9FtZpQOu0nncL6c3c
B1iDfqk2BFfwUsLpJ/E2R51DRi7c1RKvhVb+pQirUT9fz1P+8Alx9oQBAz01KjTRDEM4QkaVjBHV
uzHl6UkNNl7xDdk0gsPjituwRo8axADBk0BjzuAE+sBXV1mzwdxd7VZiZxRhT5e0HwR7egV77lub
TI3u/5t9rlAgzNWDhJQJydXJDSPW4YgMZxvoWmugiSK38NletnkQmFLLcUyQZBryF7ApWr95G+tt
nsMbnPFVkScJOa/w2Hljqf5QgxjOa1gNph6Rs3Co0k9QtAl8LQzsJjoX7rGMoeUoP1O7FgoRzFfI
B74fK+le4HODkO7iz99GK++EXE0+m81vlXFSvA8aleAbanMHHBqYOOdh0FYl7e3E+aZ71dyx2ObS
xlQ1NjRa/NBuN2NsxDhklMUf7AGJHKEOfHQ665ozYwPzeGo6wuLtnm6C4llNyaz6sKm/p2MV94WV
ylpr1ELFQzocMaCLQZisWbW02grx1BCAReVCpPrktldtceZ1C1NF4LqFI0J9L7+UUxbQbk1CuUFg
3UbzPdYDRJ9kJr4SBWkJc//gRRe0XCvLKBK9Pb5FLwQOxwky5c1Sg9HIdgccKflJaG5NubBbksnj
BTC5MDQl52vQfBMOFOpOfFJgnTg8zGJX7R2ygc7g+/HBbVOdD912hZQUcVpBt4BVFxbOwOAzJ9li
DG7E05zrS+pcbbu7DOEeWAGCYXr2ivesiVXGF4diIVMM9L/EqKkxbsmntAaN1iQP0i9p1H04SvCI
orCeNT7eMF3p5QJUFxAryAnCQpkOag2THMP4lJawtnumV8uC4SJcI6053gGs7s/dNQDZfoD2+i90
6djwUG7nWcRAcwMWW0USyGt0+VZn9BS8AitJlYMOc03QSq6gWh0AIk/jp0OgGhvw7qKjf2RJoHIT
HUJXDu4IFOGo67q85ZYfjGyEIi1RurHuBtrbz/N7ORVyEZaGepU/US1D3n6Ib0jDJZO6rDpCyhRq
Kvlsb7qKuamFKZRWcnzzaObbAzs+nJFxIMlkj5VD1Zjp1e+srE0rEXOAEa+efCMsoTLLY2rNfk4b
pGhttfsTO3w9mLmvtNZvxN2RxEZRjBW101H5QIuGfGziHyEHmbDW4O5ILW03MyiA5PPgYQE0zAug
CdrEmYTeF7cJD7n6wSeSBAkUnLuf9xhjSJwuS5gKSZvuJ37gs7Dic7g1YpXGZ0QnmZXALBCac5dz
7XBPMlt5Jj5PzhnrZlXJFE19rUPOjUR8i9V/ILZ6rZef6/1ancArZsrozPfOGHKS7rNMGho8tnnu
WXaD6XVdFzhamAsxR4pWEQOPJamY+aimEyzm0TgSfj2XkrZ2sf2aWVE++D5tDY4n6YtCmcVNXTuS
iNWi0aTOMoA0KhDGyg/GqIXxnfS1RVddPtdtZUe18ckJipiwZCFOA3v0EL4RWgcsKPs3v6j6F1gw
6oRmYYkByRN1A9Qp3IwpUXklCBoQCRndvIxMca7NQ2QyCSAV6hbu562uDirEGBBOACYYOLrHu+pQ
ZqJzzPUH9gQetfi8JCM+pVRUh85Y2LDKnWfNnAoZ3mCoKtNOM+BLNJ32MTHdoA6bsbAgHtyrC/su
HCq/dPhysY+r/4unGQqd8zR2nNeAEsVyVJ8aghUyLCjCKdMe5VaR53GPFtGrQWkFxL6trT5tQ/28
Fy+ipzem5Ex1qR7SOc/Tei24sAX8ToBHJKD8wDp76JntOtVbemYj99JmIx1fuK68kijxpVqv4WU2
xPclmxwzsP8KOsFmMobj3RROZTfUNU0jGqMEBGYDpwnORj/OFVZyBfOOQ2CkSQw+6fNsa6OmLHuH
o8wl3SCzdyNVJWl+gVYvJrBLEQ7ovKHWlJSc0DGjtjA0OGeb0riK4NoW5xOLoxRhmHN2Nhh1MVjm
eH/1o2WkyVqa8uD+4jxQ0okI5H9trP/r9DyK1SOOpyf6pVgws5OXGomxdfb20ltxvoiUBanX74LF
jkYqYR5kva1HH4ifiTTaYHwPM06h4pVojA/Z3xFnvndZc/2R8YSb8YbLP9ipmBSvPlM0a0NomCkB
nZXPOQQcU8cr4FuPIaEgy2GCRzMSnX30AuTOb+/+SoSoqbWJH8YlHMkUNSyUgUImJ/ZMqS6TNXbm
vZUjLxz69pVcDNQp7bKJSKDvLbgw10srJz5HnDYFwCsmxTghM0DmSnuJ7Omjls7NL2uqX88r4iry
ZgZLt6t4LZ5RXYF988cKnH59jLWcUusMKBeGclXY/UXDwlIhAthBz7Jbku6Nvhb7XlH3LaPh6omF
CGMFvBmh3qmpJTMeKxfOkADyLCoXqBHdrFypKn5odw03KW/eqc8Elboe7omJLQAKEMk/zWm792Qe
EO4t2CrwixouC828nTfKGXTmdwSLoSJ+ITM0UQdVaJ93mqyUS5uhW6Y/G/MbPvq4pC2Z0tK76VO6
QqaSyAyV3MRS6U5cJulYlmKXvGlB/2tIzF7yyHChuwI+4ga/8vWBqfn0v/gLL1zRiMJ4i0qJ1cme
YTPISmedg+7OHfE/6QgSIsRqXnIQ54T+XSwb+fZYkOfcWt5QeheSl8Rc9FBNQn+xsfP2FUUEMJYJ
DIX0ll8SxDjS4UNrHDdyHFICzKY0s5TBXUr+lrGBVFSG6/+fjk1X39I5u5So36PFaBSNhnrjSSH1
9h+ePQ5Z5u6CFbJ4IzQ9L0E1z3Mr05Og6qoHdbDB50RwBRmZ1wH2QMgoxxkVQ+AFleAaN4AOg7OO
FUEAYPivZFLbOq8OvNhwwB6j3c30f0W1DbRaH0Fpi5W5MasDlHVya/3w7/ivALVcHU6SWZsrXvTC
AXVruOrLs4WSnQ7/Sw8NA5/VjhZJw0hOMg0cTnDhBEb2Qm02mrfqPwD/QSRbSV9rfofavnX+N/pr
+nETUsv35C4z3jiEX1eDjIdMOCUvGAIHyojXo1YKyAKibI69Phq5bxDbwma+4zCQB8zTYvRgqzZ3
p+zzi3qbz3yT0e/RsXIJQbP91OV2mGpm0qU2KA/rtgmMf+lxyOeLaVFNvEi3UQAVDJ6iQ+bcd8Qk
yi/H6qemF/fZIFBxwyDzyECgv1puFVj+c4TenWEMiAbQcV2DGkhpbQTKtZxGhoV8LjxtOsiG+zWA
PqVpBrBkBggBaFI5znilBnWff0W6TNBWi9/M99nkaiu4AQF6klgNfc5a3T6qCbLZm5P4tfr/d2UM
BEYWh1IdK3gp4LssIlqNKVVwF+j2aQfXb7pr5Lg2PficXA1pd/M9VtxKW82F9JfPTpitjeNIuOUQ
5K0UJa9msx0h9jNn1Om5syY7RXghR8SWAg2vphQ6LVse95q6MFhB0adeJyNSaUULLl0pESWCO4ZO
UnNoUaxbft0L4oka+Fl0Gv8hOJggaeGfNh7xqKVZRnxcvNqMPdodwksrDURS1IeKe5Hn91iFroA8
l3j+epp0IHYGlsbsbcNkwKow87i23bFU7KW8WAYh/pIbgQBkRxBO7sZ/R9UyY/aMOOjTNtFruOnB
LcOPuEroxQWeIEZ8814i2i9L04Z3nZe4RkeChTCgQHB4uEzTHoT1FkViSVp/thro+FXyxA8OJ8Mk
2E7QrYIucH4qJgL2+iD8cu/yWm+nLxe3LWtANalawBGV3ZK0WAFEvM4nxNNHGrwZi2CB47TF8gAQ
8W28rULM656HY5fe1LvWfoFA6Vp29pt6eQ46TOr2xKwJ7oZGIaIww1q7+oO9aJDZoWuPolm4SLpL
bwRO7BrmNkNsEtq9tWqUI4aJRQ25SJGDA0ftajzFNEEyWIyjq2g69dmqE5gG6IqlYKkKSOVd2yan
wKEY/6KBDTMTpTiUy3alfplZ7e0L6DIf44D9UruhSfh5n0SlvFVxlfX7TmuFzz1zIoDhCVXKdAaZ
cMe5EzPQlNi3zNvuqQt9Trduos7ZnwDSLTQONFkb/Bs2/EpVtNZN3N7Hlk515YSV5ifgrfYRK7zl
54gpan1Pip93pMUO4jEf1ql0DS/4AZrJt6sxs8/fu9TLMy6wrSuyIQph3fMluEo1cjVznaGCqeQI
VHxAmT5C5niFSa2titR+HlgceCXL9zdtG0mptarp5hbHpSJZnux1BBcFk+4OBCjTPN3W8gYISois
Kli/8wh4Wqa3L3n+lu0x0DMsL61GUxBYdWLDmif+OX7tf/9SyJFMr8hWrUBW/fSrmvKFzPBzq44+
SF5VIeAm5YBl9nWnkq44KEiigRC6y6FBSAdwX2Z1isQwo+1zCZ/mg7kCFsEVF9b/bJsHMUjmGXeB
y8gARjgdxEMmaAiqgIMYZ097oIFsB6x5hOek7rqogmWOj3yyysYdbXLk/DcNMbylddd96AR0J1Df
KS8jFbZJnUUXG3PYXcPH4w/hJzEJowgmFuGAzZWwaYB/Zv/iXtg/HpZNFvlOfxgS7CjgaJWxC0/B
TBnu+4D+MMtwT0rExIhsazJPwfJme0SBNV0rhn2kSHQCjwH4NtDUGij32pSXxhTAm9lNXmKkOKto
zvgw/tNFxNb3mM9SkaUfxsVgxuoHm5R67EFV9dBee4mLBBRAU/5AbVxU7D0DcYTSs+CxKGPRcrVK
T5h+nE0r0bw2EuIoBDF+sLpqyA3kqV6oKqy0KRVSXYzRJ0M1uIYuuztV66N68yZGb9viFv6v9W16
31oj4P6J3cRih6bKZfP6RoRLDVn9WlKV8bRomzPkINSxKOXOd70Wrf+xwBrUHiZsFeeeEIFW1D0H
PRJuDXsonthKywkVrDzgxZWq6tcpjXTFilo/HBYJ0cYpzjyd2shwqO1IRzcQfHcV+7EtQQZlANgB
+qcYOykBHUUn+JMLsPB/cKjygguuXfZT/QcmQv9IVXgfJFgYIO9ge8ZuMD2H8RCUp1G2zxw5YjCb
NCdBlCpSM1hIp5vIDhKtnLYpVattZhRXld0Y9xTwXWanS42oOqxbo5vnxlruz9gtuCOKeYjxT/6a
0mWmeegHzqxMbnbHuti87v8mk2bjmDOpXY5K9ZBQwB36savhkUTFOnlIaMNM+3uy3U2JstAIvpXs
qeuUZUPCyautBVVB5F9F7dn0dKKjZCIpBLAoBfWHXt6Zhoz/vZWM6DlyWAPB4uXPhFN/lMw5R/Ax
jNfHzYtbD9yahXzEgy2v+qeZJay1BnpbINNh5wcDCOBJNev+e1zCNyscJ8B5gefw5JtIGnqprStU
ygu5Nupovas6WP2d88MT4gsZ6ogOHMR530hrLET/ZdIqGIm7VRu4z+zl+HEEROIaJQCPQh8MJ6LV
ZNE8biOegPKQ+NZPo27/qkJwrhuL8SnhDMoieBym25bnC0vOsW/CkCn0iusvnp5D1VkSuJOpnLiB
k5jXbYDFmQ7EyOrSovBLZOpxAv1cSrB4Y+RIOMpA36mf+DOsZrsUufyj6gUxAHkv9sd5xp7JuJk/
4fFdFbkXPrvQV+f8S2iIZQWLHB8jRGXS5bNS7qMVuemx8fW1lnCphCSFew3uvJQ9xGF5Qp5mPdMD
jXsU7XD0i7SHezwDYSEsfn4mP/lXmduZT1AEhLhu53X/C1a3cVtTPIK4AniCP071ODE7ezOfSoha
fbNJKBM89hCgOULShyMRSF5n8UP1bz1ArSgdEEFEx4W1PsUJXMwpF7dc1ljdVygnMM+10eG0BF2W
rrpJy6X3B3ZSsQ2CVWvSMdTh73VljkOFSr2CF182k++okV1kogg/dPF+vSFli1+ekoxhHIwlWI8U
iwy0tUi8G7IzGLIaBBy1tuJIY/8xmS/JpV0+RwhtLyowUR2G+K4nog9QtaN+9YZbdGosvd/wWdfz
azLzp0uBNGdllifmMXmjIC8TfdCc5yIriauv5p0vzV4lfcrQlsyuQOKtzJfRbpmtUaukfzurIh/2
WrXSGAdAYNwlpmUI7g2IHzaIwKsptKn7oPY9ytIZfZ7lflqdntWiGWsttwGmte+UE2msWazcYFOz
DNleBUCC1qZoZLurBxWxg6C4WQSzqcPnHG2S2v/tZlYHxn+VrYX5T13tg/tRlmeaAZ9T1rcm2I0u
Gb+ZoEL1/om8wrM7F3eu9TYXdlvcId4uH1pDqvXeEDH20wSCsVM9MGNRFmmCgA5QN1yQ+R06RuL5
QTcYIOSmnCEJqIuubzDtWDPt5q5mAdWWbEI2yToPE4+6oLMrkbOVyrpngoFYAHhzWObTo0lKXvKs
ncjzQQBrvHZ4X8h8eIaZhGpNqC7iO8LGuTq7w5FMV17TcJDgBWpzmsXW18EAINEXhruDIky91Gdi
xw6GeKcOKYWbCa0pyDje7ThUktRPe+tX9KLmDS9WsHT6RpffxKaN70RBxl2U8i/YfeTovA5+CyMT
grfekDFew9ykhkb5J3E4E+Q9nCstnnlDlhEBL4z9mdtl8sv63nmAIkmomkLvZUJg6TbH0LRPvJNW
aOhc3LMM0tsnbn5t/K69U2HSy+D3C68vGku5T9gIHA03Xcmr2U0wfsZHfaW+JSWCJvG44aC3p3rm
JO0Bu1eOeznsjC1gzBBO8Qx7jZB1UoU5EPzOc1pRA19A9aiaJ6/g+jxpjUIlefdADNhirrdVwpFv
xDWxwiEqNuy+Ws0HjD26zM2gcfPypaijk6XRpA0I4rn8qE8309/Sjck6VWS+ksmcj7kHTMJjVOfU
1vHSK/lVnMpdSr9huLWTz/1deYnz+LnWMv9MOQXdJb7kkZDBvrNJ1J+lIyl4f2+a3Y141HeYmfSe
CV/uyBz4lkbTfDUEVHRD6FfbItP39LCw4kYN1zKzISVK6KJgRDL3ynjYOxtevsoujGKQ4cjROQHJ
NkFV657z+LekyA54frrPnSUBwgCNgcSsOIDNXyAE+l5B75W1dSd6sFT91CnWRLd8ZqzCEZ/QdQxV
JJHpFdQcg1cttC8ACKHcJuCiEgCmcXpUwVdWRbPu40w/kMi3EhAL7xxgLbrs1gfynrvcUO1D5xIS
lIBuGpydworwCG0CecPxGPanIjFPJSP2Qi1LlFW+eUlxZRmZGj/Tg+nzRpD5Fu/TDqUEJdq9lDxf
0XyLjRo2232K09Y66Yxd/9E9Kz4bLYJ406PSqUAgbyQvmI+qSFZ9HYXqr+QICCkNeQU1w+wJT1zv
a27l8IZ6/36/FHuc5R21kRx+1qvT0Rv7CZiocCcSud5Gdi5pWoFRcoWbalGMb2IxiM66mUWCOnc0
dAnkCH2HUczt7wxv8s8V4IvnPDFys90eOTTaX20LspFPdsrxPz9YewpGtHjnLXK8/j89ip+fligv
TTbJrUUKnaDGrJ5M9+Yz232tWw2n1NJb5ZSu8bciz9mqbvOOJYB+qsBH6cq8HqeikPCbCvqnUNs6
lz5CJ2ZggEuRip4yi+bToLq0YtsJVv3hwZani2yNk69VbtL9PyelWJxCvR7iGkCas+l7W5lyBN7F
3SfeyPhFIVzEdpxhP+2U+Z4a9Jogjgp1YQgyzt5v6NJjiPa8ocsA5eiJvCFceyNQlD8TZ3ExPwKk
n8Dnt+pxX+jfjSJPPXXum6SFx+CDBuYRzuxECFk5ZzY1sWK0dKv2ckFKYWVa2lf0HqTieM0w3mSm
mDs76meuP7N/YyhUsNMN32YNp9uuVQsBGdS1MyycVwWGeGkeTKBNF+b+SkYdDS1Z5TI1sT3o8lmz
TqeHFLR/0ip+ZEr5jNB9DG2YrzZ2XImLilITkUt60ICzTToVdZj657fTXqSYIalAHGv4mdBKBuDe
E4qZjxF9lJyL/xhG8vcPjfYNv/SwaGEQFUzCPv1p6oH7HjvLbIxMcLHm8AJ1skAqk0uDiIuXQIgI
au3tnRF7PrMBOM8j1B2lEkBzJUJV+nRicuDarHYIntdXbppRYMZ60FZED6gv3ofJps0tGEN7AQcx
d866N6gvPiorCATTEYZx9lGz+Eu/grojPglQg6h9JF2Fx3QdasGSv3qaiDgcb0wEb5WWs/6ozmWG
sJOW3Q0IlyLhdNWx8KVLgmOwPIuBIQEjDVmTMV7qZujJAfs8zmgChsl9u3t6Ce/7kqagp1Pn6bEW
R3da8Shn5bhyt2J1YxDN2xMyspEbA3bnDuGDO/mcXXAfUf0VFTaaUvzdLbgn20WG3Qc7cuPmXAf3
VVmgdPIucNmrBm1yPLEFOACng2Ul0HYyGUlxk74kTBQISn2owdv+GZ5oEweew66eGxfMiy+4Tpjr
lusXMOPeTIhkhW2ucCX1+P/nSiU7IQzzGWflxTsc3z6oEnDLBZASExDPpKWyINMeB8Bb5gyjJIUP
y5B8eFTu2OpnNweQ1MsTXYPkN5lJWZ6EySrtb6ysR9fEamDqEjW/XAy5wmDK6rZFUlskm9nkCjr4
N7Dh7xXL1hukVna3o9ZD5Z/YlZO9wNzFCo9sMWUNoPj/BfFkGiJX0WS0CjO6cvi2VB/aX/9IYa+2
nMqsNBGAqlt7PakmO5ihOHrF1Tux0+zceX1eU2zggBOfGwPn1N9jcRGbQzVwW4Q4/lNKf7S/dJRW
xxdMS/VC1muVPf93HAoILg4hyVvWBmDRrf8TVXgGcKaQAlM1EEbtqtdkzcW5EkHmWwufEfQfvYS/
2OXH6f8ZK4AOumucoeGBHTB1uQ+GdFcM2xzbtG5Nicz0rAH1OX+9sOf8doecXtp92YX03LQepj/5
FyOTQxC4ycpthDcE8Nqm2GnbuQLTFasvNBteVGYrSqu7kZRIUXNZRwFrxjlhOr6w+9uobpuQD3kl
Xg+1r57iFg52CF80rc40Z/1fHFfsQur6ARLwSy1jZ4uTbbd95remhjTVPV4YJkkNV9WGUh7/Zrmo
WG0innY+D4EHN+AxOpj43H6AgrP6tOJW1UxU5by06Hgf6SzK5+5z9coUZxUaZ4qwhj+8bK4qnerC
SKDD1Bkp7tn1GCEpuv4ArLSVh22iS5qnLlXr753Y23hZ0Q9Tz4Lqo+bmkdHXrwHuQ1ydy0Tzd4Qs
DNtHYlZPKNC8ZEnL2PMC7UbzgKjzF2eZbr3x9MuSTFeA2+YFuaaMEY5z1yRI0XN5T54DzVNN9XxV
Zdrxtazhv2r7IIoG6yW+9kFaAtdgSDLnLIvhpUZWkxfDdG8VOvtaCevgtrd1+Xqpsi23z2KHdHDj
pv+9O5CNuWPQx6I0zs/X2h1qJi69hcwBHD/4/Yx1EqMfNysukViFMIFCzELHEBWRXvsaxnbhyS7R
T0x+FPP2ZHXW0oGsW2fAQoAqPpnVI0ToJ0tOGPsxInHBMLUaDW1HpxjaVA15xJ9JWLI0zVvjrsmj
wg8IUtjhZHllN5UqG+10l2JOxCacp+jsUZIKsCGTjGHXRcHd5/JZ3uJjSMktXW5AmB50XCBkdA3G
t2emzHjHR+Cx5oufNjHABTUO68H3tI1Gq5oN+2PPRi+kuQQnCc3GRNBBC5WW2wp2kYz4LEqyq/Re
30SV84gPN8yPaCkv8x8YOccinHpENTkhxEhPMWYmShkzcfCq0NzCEzJb2cL/DoQCy10Dbgbziisc
7q/6ft9dD7rm5+9xrciUSRNLuf1AlJn5AFVbYfSMfS7Zc8DokqzZ5V4GHa8kJMWxiX0MGs9LwsiS
OoM4SFjscY5MxQQwi8u0P+4R15b3pZoYG9U4g2iTMN1UglI14mMtOlmOxKSloLa4lFtNptb9x2K5
A3g7GWnCqvsl0SRfbUVBot9iD7kBEpJ+j8ABLYjHwXwnrQCeD3ipxKXzXO7851ynmw9J1lhskKMn
deFZzccGdKgnoLkpMsAymYmwi7YE+0EyFtV/3PypnEV8Irhg6p9dctNS5jyLpxiZH/iVwIFRChnf
cG9zPeT5O6M77/Myf/tyJ9WBOuAIpfSId95QcWOj9gBnYAlNLKEeBXsh7T+GmKtZ1TGkcqRQo9nx
hfDeGUDBfZPZDYwSdO1vDgWHXyS7wI6M+fz9ffFEU4rEzkz8v/Uj4hpQajhXT1aICvKbzASTLID8
i6L/jsZRfLSbebPMIuygZFmvU1mupfE32K5psBDBxs3OYlTo8nDe4x17YMCPW8YAgaasCrZysBMg
o6SQtCw3qE0SCou1i85ftUsbxTp/HG4LwNOr1hk/JeSj3t28bLmlt5Z5hU7XuNGQVrFKA6GwFLGR
eO1aG5p+qTNNceNlxsCr7qN6oyaCgql9n0lKSu4Kndv96dRa7X+7/UYhVhPcxOdyQC6RFCKN4n7W
OJb1l9n0bMyHqNaJ02oMh+ASbfzcfuHQiujcbcfQjntLDWgSHj9emydF+Blp0DcFXq29WqwDVwGr
GxEbPojTyQkHLu0/8m3KvpnANm4sKseF/o29CJdfE3aLu/5nx+ycx0Mi+FLcJlAwMPDvWd0oJFLn
icZBZKFowBGIj+75TjAP9FCRlgKQ/rgMj0XRYuO8QecGBS8nHNndV7MgCgdASpGP+ntGi6rbNpZc
ju+hb40+m9xyYWuaIu8S/TtKrJkFNlVUQYpHdJmhk411a1Vf8pE1OGhmnskoQEW+6BZ83PCbJG18
5QuXfUMyN5sopzdy36MqHYdyOyeti651zjnpDrLVKM7n4fDaT4gGIAnoGRArOrPUU0i9dXG/Ypw4
JGinJF4iiMp/A/TWeMilIr9UTWjpoKMI5KGQoo6H3+HVSQYv/6ZmMAbnZlVmaxaErfgnk8mhIvps
5POHiuhEyZbi+SX8rS3NSs9Rxrm/jmSpIQJ1pCs1vn9WXAJncPu4852b41GIIGz2h2TOioZZY2yc
AaK6qXoBUxVGePcUC3/gdsp2A0H/EAVBzlIrzr1DfFYxuO2NgIvi8O4WLoirl5xOSlek2p/I1ZeE
tLzowCTH08fb3L+2AdXNTy2Wzmo+eicGS69aPHqyX6NAZy2yr+4XvfD8JtN5sC79B3JXh32qT5e/
lLDhA4iFVDA10vDH8YGj/ppxNrrb2/vNzJ2j6GUwGzgC4XijwP/htX420VgTCDg6jt25dN3zIvbb
YtGDlBBR1VoDga5qwIm9V4hjX0D1hBJ2ELGXBrKA5SHxd+hdFINgHyGzurbUfjTRNtQcrjEwmeNk
BrDPG6SLH2D6YAtx8LvQG+L7BEy7UHWXKUm2sMMUiFiBGxAPFPm98zMoIjeOEI1/JP/BocclB3Ep
qaNB1j+rfD3e8jMFemXfAMHDjWU1csBAkaTzFhJHUotNOjyawFM1OYYD9Ud4Aym2aWimQLjp5zGO
Fs6MywV5Aj/fLKrqUJEDOX0PkA35GIHqBAv9nBQuVoa2wGBz0tXDiupLNAtyxp4MWt0LNS+ahtJp
zwDP4vfKgIk8xCcm5U8OGAybwww3kTooTi1XaFIewSvkCACgVUvChyMfrL0SPSOARvR6pUlFxomJ
Q1TnV39aq34QJ+yYfUSrI/ue1UdQSvFvs7F1RQIM0/etVLa5Xz8UAxJojbE+BLG5QmJCBeA9IlZX
gy6s1/jWrTSMHnIcam24Myp7JXVfWwMp7HVl6Lz2YXLAvVy86bbfUEketvpHa/kMcwFA1wLM0NfK
Xs+50bNY7PZdfsgt73HXJQW01wgGgXGQgQ4vWoC1AgRXko7GlSR7UIBxdORRjBuWx+DCKCFl/8Lx
ttB4s2BS5RDLEVu8AEnlY/Ob9kc/gmJ30TaWPMZX7QxElnQkxdU7RY8hmr9WOsIzMWY37EFiQGhE
wcv8yXm6H4FK8+TLrjO1lbrdCAXrx3lhzV9YA05BtzMklMpukiC7DkKEQuAtvpUdjHBbdaz2iCa3
99HEFrmqUzvyi31vN3+qsZKVBJVKdU+U3cO+5J7Tqccq2+yLOepRoLjwIYdbqgm6Sgk2qKCTIBn7
+5JTXC5uTXOpiO7NcOuqcU8z+BKZJc/1nS7i2vaklq6hY9k8ttp63RpFNlOzfS/n2vaj0lyX3wNg
oKYbPtXU3rlqSA+IVblYZaufEnvsTTkwptq6ElifdURR+3xEZ55qf/7EVshJ60HO355bm3Sq3awQ
JDxkJc8cIY3CSnYqK2fnP0tchRpYz5QQyfdVMC6+BTXeGmLpLciHqV6pnThhACGsly9QTKNhK+3O
sn0NH2EdBS+NGuFww1RFcDEgscUf5JHbV7w5bs5CNaR5tpe+/lNkpgvqMH53VbBOOD+iHSpNEyF1
1nb8DFDM9Byl3CVNqW2inMbGy8/8vDdIIZasa58V4szs7DAuqwHhX47TG3BqL8TVH1HXxiNYhTU/
vvcSgxowhVvyfUMzIN9pW7i69f3rTfRcto2znM4hDcwKeIOrANweBt0QF6Hexa+eMv89istufVVt
I16kpq4fCcNQ7aBJCmBQVf8slzHe1MeIGqLBEzSqx8gzSOLmZm9uylPzi3ipRFRguA5MaR6v+T53
AWruKm0PmykzBgPfd6Seu71GWdliZ4BGJZc8uxHg3w6hIZl0iY6MpT/uNAsWzqBmah2hix4rjGRG
OLc7b2ZVNMgBQFeK8THvlNLgkqa7iIxGD1mVG+yFUuk+ojOQerDYv/gMLIFeziy/U9gKgVGR1CEp
0zVbYXIk7icbD/v4nJLH2IdW1ad/7Kju6zQDTv9SRbRqZZNYGrSvC99twRMfULckeav3KfnU1SbA
2QMY3RSBhb0V3FXOPQkZRVq9VIv9Sav7Y8W72btjdFJ1kEdj+u4GfWo1rIxRYPB2wLiqyQbaEgOg
2n7xcQsnQphgliCL5Di7dJnkTbWbgqM3B2FOQ6Y7tHkxI2LJpoO6Vd8/am16re9C9HAF2XQ0W5nQ
fnaUJ28+Okyt+xEhCSNVEPzP7XiDsCRDuKAltLLmgmcNJD14Hdd27HzELs3E8rZrLQmM6ZBx9/kA
HSFbbeuLGcQJciP/PKNqn+4tuI73d3m2aO/wZT5sUJk9zO4lxFwbTCej44Rw72YkJ0okpZuX939s
KfIlNVAYB7aL2B9VMsl/sNjuKFqsDnUFyeMvO2KAY6yia8xWcawTDUySk8DzaE/f+bMI5G2hf1kw
eiE3MlWogrRdP7/G69uss7GUhuF19tcc2nmA2n9k5EsXnoBx1YSUR0QEYG95S+aD1bY/01Zyn1qi
YQPu5xYMHOdaufoRLey60OcwxZ46LXHUKZwYtEuXv/bAYBpDhhzqeNj+Vm+4Yv0nTc+78CBqbNCs
M+zihFfrOhijQZdvCPpnNAfAvwoH0hcnT3r6nFu/RJxW1EaMhydaKsg2DuR1RET0LGADAWF2zaJf
0WcQWVZJpHG8HJSyGFTM+uUzW1PgzlFZgwj5H/n/KYdXjuuuDUDIUiR2MuTyMrs41zqETyQSIYso
buFO4SoBeV7oHvvOXgfdlUixxFQhpFRFFs+RMRNUbvdlbDiH9CJzPcQ5/nVkIZ83kYGqfyyAp+gL
d0VYUfyTjzlBeGzLPYbMDWNwIHLQce0Plc2L0i4ErWR19k/PnAIIYRErtJH9o5i5187UP+pWBBLj
mrAW2TPp1R6oU7SdGcXg3TEFs0TC0cZhqTXCOzWhv3aoet4f8/W1ewKcWVZ7fNZgvIwZgklKpeko
W+ERTkFDQzN+MQhjTGy2R9MDglum6GiRqeC27pYgrVhFG1KxRRpB6hPw1CfW9qgAioIMCs6WeZVD
pJOsCyhM/Bmkmpj89wlmFgCa1v5yCCMiQY9bifAyuCRqDfyr3/E8DprbGrmzoOMoVJdIITciavEt
wHsmJ2PC0Kui0iNfKMfZy1gXWNsgDLCBmkWBz2+cdXLpvLKVfcMUATHYhtWcIpDiCz0tqt43TcfK
NZJbS9L6cmu8QxWXH1ZWcLssI2u7tjWTY3h0GaWay6Cs8kDfGotqROG8oc62+pBekkRNcZyLfyGn
aYGcSi4biazIXBLb7fHz+UBUEOmV7sMopPyin1r2CRFKz/4cBFm7ppSrymqq5dGjPNDZr6zMoDvp
QCh+dR9qZYguZwTZAh4XZMGcvhnP6cgWXHpoMqix/wtC1lp18/A74UQUCJq8Zl5YkuAKh4v6DrMy
EodXmVB8qqwVEAdT5pzL1RQy35Fw4DKNk5SQy4iPI287Y4wWgNlz3zk7lppNNpsohEwXoSRXx78r
aeGOZxo4zjht0V4UGQ+T8m4K4EQ7gHrnNbyIYa7Xu8dpByktaaJjiclBnhW97gGO3dRrVrHKZAu8
ad2RrfJqJB/3xi27zX35vtkAyPjtbxoG+Q1nBDSU3SQqkMEzBSVxioOBAqp6h1epyIuQXbPJEC5r
WqT6+e00r6vUBumS8LTU80LcwHREVEyU4X4vg81BEPnSxkFbNmR3itPdKEjm88Bfe8nuZCOiCHIY
LRSt5KSxj8vHgDuVD0mGFDWZexAjquze3SCP10vyTi9rDZblstkZl3JDnRCLCCfC0Tf5hdi4Eb8p
jE/B67JXV4AO8uHTr+EYlF2MyVmD2Q/z/XZRlssh5GWA6sYJfhXu8J1hUDHFkbSaywl8QCxFpf7K
XXjAmfDIVXkENkC1cu0PPzwJnJuzjsffxPLncLZIHgnCNd+1ZaWT/NkpX7ZP9+8LEqttSVHNh2ee
E69GynQKUkor9BhtX4zkLfvjKmBdf36buU1iaJBAFJr6dyiulzbYrS4j3N7E8qsVZc/0YSCob1pL
qRRdYA6DAjNKUjcWmt4/RLaKq4eZB9HyFQg2CbyHi+f+aFZFhq043TmVGFQvmbhQojuCodaLuh4O
yJba9gKs9K4Ja6uAh7cAwZ75k+o6BB0DQm0xjzBqg+A5lSQEZqN2fUdLYW11QvpID2AYqEhWB/pX
Tt+IOY0N+awymF/dVXe0bSVzzN/WR0rD0vscfoMJs4xmDFrSJdxhSvrn9yTgMA3R8wKYijz3SoYq
9tQ0fgouayH+csEtxoMchfbXbh+ZZvwkTLVXpZdj3SCWxTISxd53qEWPviuu1tXE2ptSoLssxY6y
shqkk8f9Uq9a2pQieQhn1ojZ09xWU1TUT24Xm1fTdgbTIb9xxaRB2a+CeArX/EeM2Ldd4TYgfZAX
ylvUbJaqd4DsdihcsOs1Kuivobmu4puDbt3FuDlF5yLWPVum73kmQ0k8jqvMEByH9ZAKn+Z7tPSV
w0zhxrHceOxlF2nazdfd2wWRNJ4VYpSlmUHVrt5XTQqFIAMLICgM/uPuGlC0SA45z1bOPd8tF1kn
OsYv6oZ+QaeZQ9gWQfIPKiK0WHuCKOFDgHg8KeFwNygkcoU7lq+oMJUoPh4PKxe8CkLfI+HXVJep
HwqYQufZ5ZBcUNEDBIdifXP5HIg44oB7zqcT7c9UFcb2MYKjsYU0P2EKpDRYxq+KkhwtXXvroh6u
BVdIN8+a46oPS0RRcr+YnxOoxXrnVttPu1Oaxn8SkgmyKfntfq4rC6os5N0LYHf734F9DVBPD/iG
YMn+Nz493dbUWwJjfhXDSgxaAiMu1Tn9LVuns3J4+ToXqnQ/FC6HoRKB7TMSjzUtyaTgDM87sjuC
Wp9Yys8gwTmMz5M9DOlopFMAigXEErKqfBAZ3CBP51L1CDs6+hkb+nuWv7t4IUUM048Bo/2YNuvR
Veb2V8UnaGj/Pw5H23MqI3P4CFWlGMqfvzHqGip79JyaBti/Oq+hA7XujCpn70e1lwBE7nC5yId3
K0tR0fYLoizUKRZcPJhxHva5VCN2/sLVk22tTR4P6MyMDYy6GukTwkVr0Drht/p7H8JQVZQCL2kr
c7He3ArkTq6rT6SduS1G3Kg27AK3wsFXC5xfz9v2r4mP/Z2WIsZsOuKDerGq4zFo1i2wx1G0LgTU
dCJjoVbJEGJzSQ6eoXUXyA+c2c5756Ch0z4UZVXgIVCcU9Kqs1eHA5nliVFaWYOH7zQCnZNRhyUG
njqQJ97h44FpnCitjsrfA0eHLnHMxHnzNtAB/qjpvB/mj7czaN+Cr2Ew0qFVlFXVQE5J4Bneqprn
iquyDe4xVhMQ/blYIwvWDC8+TQsxVmylFnwrfO5e8T0jkYCroin7AXZgls2h9L+iK0U31gY4yAUk
F+7M+DutpUa3K4T3ed0tkmNtEYqjp76pV+uQRRD7DZXCIVpB1E0z4hErfo2x5B12q8Tt0WG0zopr
zweisbvgebB9OVxP6RecEWsMvT6rgdx4wk4dAxR+5bGZ5ewN/6vKPeAorgIh8feywqwIE0EABSy6
bsvtewnd+QgYA9c7+YeS08CPNd5jH+v+q4TcbFdt1LWRpI4Dgyu6CiHGofcHrKszEFdrKY8SK8L0
rxZiLRkFJu30v4X+VIn7Qv6yFUmpeG0uICg/5C6uGRpX6z9rEY8JrBP0jl7JtiLlXc2An19iLYOw
XMmpHURNkrD/M0N5I4xZ2+8vzNE1eJ+bEMrGL2yok3/BRallt18/CfY6s3BkOevJAG+HMpk/P5cX
tdbG6AZL7IaCD6H/glMcGJmU6I6rS4q+dz43ND+wXcigUnR9dFD8UdHXocJV/mWl3nkKurG2FMN7
qHytwd/uusXRVpwmyq6LUdWJWR76YyHEtZfIC9EXCw/OvnadNqlwZp3+bnzrHDB/m+C6OZ2YeJaK
FNnjvSjbEXAVusWvS6+focK6Lb3ZhVacQ0aLrboIyxqKTRNsos/zrmX83+AooBO3el1jO4oGiH/R
kvGu10CsnLAObuE+ZCvDSy654i2vIdZ9jz4PygKbW+J4AFBnM3xEmGd06475qPeotyJg8TVB5vU+
59jzIfKXCtaFoza8F3NNQEC02hPAd1IWNMVx0XvDRoFPscAnn2DFtlybn2Q6I5RIRGTbtJE3Eaor
FG9JfFJGr77pdWAFXUrjiQYofnobZSWdrDEmtCsFilTNvX/bZXo0IQ2xe1V4UNH5eIcpdaGo0NqE
aNOgeQI3qr3tJ4EDOxuBLSbDEIEEGvcEmXHvV9jDXHTuZn3xEE2yVkNQeqqD4ACmifiFda4L8apu
Rgvum+fjdVFWKnu2HQjbfudK+GBlRvD02DjrrRGFe61MKEh2HW+pdKtEpDt7REgEFDxKJ0kE1aR5
OTUYdh7mWfUUCQ00kxf9+mXGq17MMNuv2vGnoAodV1OOQ444+fJish3b+GEuY6tXJ0l7DpCPSdqW
98YZJ08l0p2bDMsW6ovllUtiC85/hkZR3v4Cxqc0Db0KVrSNNitfRftw+lPypn5/EVELmICOVsk5
kQy+FQOICCQliLjRhVdUCg8gnWITdhg9QLEuxJcYg1gqiwCIfaJtKAMulKybaEeW/AtVvzMWNNBA
NUDezWBKSaes7hkKA/VwQj906wdrKY+euMCzOlIrcA9fnPYkAoWEpoGIVBrPgR5CoIJ0Dnj/WUDr
Z9Wi8z0TugqSgSevnXFe1b6W31CnCI9VaypTgT47FQhdB+0xSwfktZUP5hIXvYhm+/z1CyeZCtp0
1Qt5YHLEqSJPfYsSN6fih0CE/QqucboC6bgihcRY0rcPqfDVAhRl028Sx+qZ6OCQDX90vVkFLVAQ
UkEVE/5NQmF2/V684xA3HVNTkadhQu2svgLDve70cfIKW9tc4o05+UVVjRcazijhTIOmJsonCoFH
p8+eTH9Jt7zYHJ+oMd4OmpAhWMBMqvce8e7d7gL90tqw00WTMWQzv4bWKDrb8kP1XGxxZXBsMBDb
TECxnXpKzbviulT8//M+p/6mZf663a35WsVFkjEZzdT32ZwRQHwM+eneIaAOt+W/Kg3ILJacVba3
ifNVE7iFDDezOFGx+SJW2XQMHs6R6QTJfSEcNP1qDVTptaRbHLBmYohLWwZCQM0cpiTIJmYWe4jb
tK7o1ojnKkdb3BR3E0rk2kbknASMDkDvdqtMx+5v0/Zt7BEcXYeBR5GTjU9MFpx5k/kaHz3jQRhT
NaxS5+PRzjIqtzR1UTYSsr/o6z5SvCC1kd0wfs0KeZogrro4fQ/qmpzFl4587N9H4XvJVTM99iXA
dbLnRgbFetcMHArbZDRC4/uUhlZPISHHb4AVVGxSpkPbPOKvxla4fkwKgGisc0rROEABPTuzPSMY
HxMZe+jf6c4FjvOHATaGgcBRSKb1ShyflUOZ/A0fLwyXMTeibJro5ZD9agrHxUWD31zqueNlbQp+
8zXmjLX1/1ShZeAQ8ZMuCSRN8ikNCb7gxfTl3lBRVr+lwAuJMC5PfSQrFghLNoOexoP0eWI8ldnk
qfk6f9KB+2xEAn9dp2lSwvQjM4mpO1MWQ9t+MKnFHGE2dCd37I8GgBiMjmJw05FOZv/5O21KG5C1
QGY+cTcmvzW7sHm14Jla0C6d2dKJOdXSqz/2jMIJwPwIeIyvTOJVa7w2Mm6GYPIsb/B0zj5L1bRS
5K48+fzhVdPVmAzL08mLRFHsOZaH503AvfJN2u6R6WMsixsxRJ/eRc0SL/HN3h3H0JiGuaeV/Kkn
wYLZquSx6mTtH4HvEmsVX/eb4wcszy8AMzejDHWe77aBldWFo39qNUpxRExJ/XilS7J43EwSWjY3
/Vi0kPvYkm4n9cTESTkQLiNZ0Z/LFBytrofYWZPbfpBd35dxyRkYUm3ZMWpElVJB8+X00MmGLazf
mCMpkovdChLlrXma24JSVglJACiJkM3NN115ethR6kui48Cvg9QoqD6nQpiIZX/lgyQJf1QqSYeg
n2WqfQylQx8pfbwaHTUhWdTw4sYv5Ugwe+mmaIpW4pQHa9d5b5e+FZd6RL9kcPHgQKHko3NF0iz6
wEAReQbfI1z6KHqmagvdZJ09iv3Pcsx5hcKJIcDI+Ud5ofVfgMFXPeMlSDpj+/hTCjL8YzF/qBko
doLCq7WAjv97pVkYhBwVnjhmPkq8UBhWvmJJxzu25fFt+xNXyHHc4c7Jq0atfNyWRTl9yGIuWdJ/
TfS0FPMcLP1gNHGyYTaXPhEbQejHs8++0a7UCZcCPc1nJ28mUCyaYfyNurq0bPg3C6lTEDFwSZQf
7wy0gucKB8jM0f3jq2lgQ9x7l5kpMr4vF8RbZGESuZb4UbQJ4Ha62NijRh83B3HpoaWOgAhOD/3n
pxj2mi+nNgnlzTs9esl/GFMw4QsBYx1p1tVqQQYSRuW+BzdPDsaEbs8eDwDPr+D/Ho2y495fJCMI
5A2dCHo6FsUfRDRb4CEoyDFugjeix+/loq5igzy/2OD30RwkO0ZBTDTBC4PRhHPNkB+406waw2/S
JziU9mRzE+fN3kbFaJuNjbhN9mIKESyp/gs/tIw6Zg1NmPJ48pWJMLpESV+cTzTFG1cmleXzNgHb
M0Sz5QG5FIgnIxWAjot62f82leM6XSnZQ0+8g7J41G5mIqhyM0+qzeiiseIa/msJ+eg5u61c4I5V
RTtPuucPM0eQd7huByrRhwtOx30/OsRdutYGdzpywqpvtlMY6uQNeJWWLbWhe5E//ZjW7KHYKMu4
uCOJv/qERHla/U9rNCh+4iUStMFVF5VIp3xuhMeLN5p1s5C3NmvpPZYE7+VLElAe/1aBuUvVeY8s
8cbKQIRrmhbDHt0TxzKIvyFUbjgshu3ObtrQeiKhLlGhm6mNFsUaFQ2sGKwJZIOzb4cgTP46WEvQ
g8rOa7jRd9Nn5v4a7uFFfvAIyFx0J2BO+OPyfew2hGoUBOna4kMkEOmRQ8d+eO3ocnUqeAATPW/c
iQaGV6R3ABDhfbeOhg4/msHpEsvTh9WP74ckfi6fO41dKem3RsR7HDSVaLa5v3TdYCgVMkrKAxJ7
M5XaYf1GEi7pNVRBCmXJ/lbfDjHELl0tWzlixg1apqZuSj7wyUcI+5+wSFrfbDUyoLUFY3/VvVeY
3nUJb2pf1BKtrnz46XEqy3dt3aagW4gakH+CcrSDmqR3VKjOag1e/sKrQqsNGvcKfoWg8WYYKHIY
zShHNEwPK/roHeJGzUqZPBsnQGOGUVqfPv3hpc87digQzatPk5VKkklagASrBFIWrzKRLisW9Pgr
cifOWQ+Aof/yI4U7fDUqQVw6wIi+dZYWxD9rLYv4b6BmCGoXwUCXPBQuRk2mOpe3QXPLZexy0ZDj
1wZx1jPQq1u0z8VxgWIEjokU7M68LGwzUED9UcEBxcyS37p9u2qS8M0wu2VZAg43JvcjyzhzeT8b
ZR2r/09JKK3iItR0BPNrMV/f1sujmuHKXPYIeCESzvypCb5dX2iK5RiKTB9EcS5gMNZG5VhQYPJX
SNAh2RNde1x5sV0FeFusNhNCi+sDMlMkOjwW5psdr9jDzfEYnJF1pgNNGz/LtTqTJpbF8J1V4ObO
kUBjYHhxRa9BD9a3WK3fVuzBAA5ahSV/0fj69rTeUu1kol3sXSQp+/Hfim4krs2Jza3iyKbffGE0
D7MZ5xWYuOJJDivayx5qD37H65zcV1GrbyTFddZ9U8pDUdDZbcXXd5aeOsem6jGpJ4Hh1COh1idI
BijBAlkQ8Jsr0/rUYxdPubAaqtkJTp80hDbv2awvp0AVJHP31aMS8pRpwiwYzzyFz9ruWYH8yN96
luGQZGXMzMmkEN79/wSjpeHf7Pdfz8WnL0aBX46kHHreY434TpKOkjjcxgAX5+I2mo/l6m9yxbDM
SxTQgH+PAUQLKJ0sMVROMTVgEq94lV56U6orEGswIQ+pFQy+of4DmK+j8q53d/uT03koeTTvdtLJ
xDMMxbwhgNKsWPzyabNe9yIvfoFdqjhl4rzGqoy8xkVhyo9CmJ9pqAXYbSh0vG+VZBmBOB846OaE
gk44yoAzhMYCH94SdIh+hft2mK3jZiakrucb2m/jcXBBiOO4GFN7oZL3IBzQtC7tNQRM88I1Qyn1
4OU1GYuTiyvg3xDTj0wt4bbvPD39amCtyWHnUnwkpNqRg8+q63lqTPnkc8ZTJ/Vb9Th7vPl2NbXA
3f8V3pN76CFfLawecCUFhHD0mke7txndJouyVWYB51GEZvUf/8FKfl80b70VIsMykUSGQQJLS7EQ
cbBHOgLkV0LZKIx14I3BY/eLkMXXMYVVfpTiC5stgv46S9x1zN+rtcQtP7k6DlsGm6UPPfNWuaq/
Q7G01Tf2iBzSSawxnu3TKQV+ocEFYLbAoiYufi2Jt6080LOGc2T22Q5S1bfslbp/ln6GanqvFRLQ
JSgVGolAbXa5v2uI9GZDWdp/ukNWNJUFkqm/mG5xkYtJi1YCkC6ybdtAyViiaf6XdrdZcgrRUnwp
OG8y6/oUe8pnVhPgai7+DpNDlpBeNoUM0mGqME9iG4tMo7qfPPuLqKr2CocNBGHUmEn7bjNJ1St0
KGRYhOqCxghn+l/v2I4bEvpd0mXFCRAvk+kVbDOOYBbdWzHU6ciFt2TC6PqzPjNZQTiQj3+LLyVx
cLvlgO0LitSNOLdwySC/Y4Iz/vJB4v9TpOBD3ClSwlSjI+jeJZa86c9Uez9bsP/RTxM0ecP2vCSK
DvPuhm94kDLjK/JdLcuWIqpKNpzS2lwRXMO1Zz4Nwa9KrhkG046UhoFJcwX2FFLccNPAvHIQ351h
Ar9ZdTwhCEiL1QGnPKRox6p9URnWyFR+UEhRFTJEPRbT3GN2ah62aBiZuOiOHatPGQTQCFloDfGv
39gFsyJO71D4zP7LfXLSRlaJHT+i9q4SiNNDE0BJaGxwq4J0955dbJ+4z+/5NBL2Lpg4wCdVYIJh
KaV8nogAZo5meh44lDvX5e2Z/QnMXwDDYuyXUaRtdSLgSlIDL4QIz8dQPPpN1K0t573IiVhzZ+dF
ab7UUv6Y4ESwQ8UogWVpQblkxqKLLeVxlImWrG3VUEjA76ZySWV/LH3ypXbFxP5j7Ys45mvznFIf
5eAP+AKcp4a3WbeIVf1F6WehixI3dWqswjnUZ32T+9QRE64qK2d8h1HHdJLwTEt4yoSsMbQ1jpvO
9LSzN5wFxeizBJvyJli2v6Ceatp9XxzUemxiTP4yVn0VfygFazWiWCd9a9AvgpteoN14kF1FjKcf
LJv0KUpY2QFXKDYvAvNUlDybaPQeYdlQoF8giqYReeauTMxaiMPTVyfn9UhjUCtCfjjIXJl874ah
DHBdCaaeocp8Vh062mwyJo5CjluZRlJ88lV4SMvIzD1utfvPjWDyMvBeDtllyC4YhP9Wn8ojPDga
njsPrNwHB7vpDGeVE70ORBJm32Lr0t9s+OC+NbIREejEOUPwhXCDkbzdJ1Akv36zLZ9vxEGoLcHe
bunSmD4o3+q1TQRyDYjhjzEFND0MAnISnOQWBfuWjVWyZU1GP10Ai8Zk6snlM3d6tpHsc3YKYUvJ
zAFP/blUPt3PQrDDX8yWGA9b6SIekboGu+5NZk+lJv6Kng6AIu4AgtBZMHOxxFVoH9J1mL7ITScK
NuVQeflbIIAY1elPlKPmPi2/0mHg9TQVCXhJpBjBMjcmGmZA+YcgATebWoDVMj+CE1Bfxizyg8xq
eKByvWp5nm5cKwy8YMYp+UPEgA09j+5fqq1zeSQbgSBbaypJZCeqHef2xNX4Z3rPSeZMJ27/HLKs
lERYncOIuXSVlhXT2NXVO6+lm1GRkv4b37n7z0FJaU53btSrCh98abMuwqRd2MNBf1yqS08gqVns
GwHXPc8GYyVIHrYCFOxGIZI4SO4O3WvGuBckuziiL8ldxpC7d1qhBGtPrs5hUbcagCkzD4ek3gUD
iG1ENmBwn/Ydc3HVc5GVLhB5Seb8SLbk/rDncV3gCNzm8BlVRPCfneazpurCEEztS2rXe/JhYzRg
3C/lJzQmJsAs4aS6QNdCGitO9L+LA3plybjf6FFzJjHLiQmO/HEmsSz88SBsZRkRVmNQ5qboPPRB
wVjLfTao79HcbQKTgOhVVkQhlbNpKzRUcOKrniX4KF5gArq8OVR4zjvTiKwGhOB1jwxOIaScCt1T
GeFvOhME/Si4nJSlY59KJsySLoeuM+VZcoYnY/RcWXso44IjJ2Peijm3CkTLrZouawhBq2oky/fa
0sxkjfX0GapNk//+LYVpx8qwVvRJe69TpG0fOL/9mIdzdp33C5NVMjzMhgk8rKR9c4ou3ZNWW+F7
R79lBoEQpqkgShDfLbuTilfRp6Uz5OQ9AMjWymyUMjgPhRXOAM6deNSLQQ+deAUCYikvIXg6ptSy
pj3JSwEYCyDzsXcJ3WTMAh+nUB7VLP5no78AxoXZk0VcYuU4TBeDeyDSOT2SHxNenk2cK18VA6oQ
QPilDhOBYiZDKB/gcmhBGL2mWQ4mrx0uMIp3YtvhzEC5V/kI8LpJkYltlUvImhEOrUnsXpiFGWCY
6/i/+zyVwY0Mdu4LCQnoSo4ysIcdEqeIF70EjxPlOX5j0G6vKKqHMumkpjZfuBhEJsWduvNDMSV/
MfBDB/6NjjDGjjcBG6hgZmqo28rvd7QVGQJtyollfkwVtI+ShQbsgzOdtoCqAe06ZWw/Q97VjBRk
kMtKTb+Qt5Z6h2SjvgTII84vGI9Xch6FfaSABQQgtTMv3Sqns/vSEadCS4LZqY17c5aQ7Et5hoLd
cJUn/p5wlRd2pQsZgMxlAYDAHyX9x5U5WSKEvre92IcIxf/eJJOEDrg+HQLby6dvC5VyYpta9IF0
Ss8/l6zccXYwncYqWTfT+GenpFVw+un7ZY2xBlQSKvbCjKugACBVzeK9NRQMtFLoIjIHK9qnFTPf
NszBunW9y8KSz4dNJOCisQWgv3JQlmHirONDo63Ng63yoes1S8XGZYXm4n0InKa+6jl4xJRfXO7c
6Q/QYjQzGE6RBswgN85tMHOxDyJGUPIXwf7KZHjhI3CmbfDOHkiwlaEVsIKbD50b11/E4KxFX34F
tQG0Sli5Xh3NVzEcekjkfMi+/7fX5dJBVMMkzdnV2OYncHC2kFrvLhlHnq45DJ6eCHnuXMWNVArT
TBPTfI09z786khWgJt2827xMGt8j/Ey+paCICXPveRQUItO2IbPD1/k31s1LZprX/i43TTSIICj1
p2icqyv7o7/F1Vb61p1WaJVWo5tq8FtURI8KU7vN5jqhuW/72eJraLCvx/gOebxAPuZrUay2iF+5
HiOg4u5xmRsBZXIQiEnzz3CEb0xVVXFQ9pTJz/1kUR+V60YQMI1taHm8vtCxQKEOJZJlSskSrMQZ
nTmBtSBjmtqovXtUgzA4VtvxYk89GboudeGPePJKvjm0rJOdHKGWJZG5Ls/bi+hcZwq0Gn6SkSnU
btGYTN2+yolLvV9FTfhr+G73Wut7NsZTWcW9N9/RjKABadmUwAigakAmxWNwY1e3m5JZtuOGfKP8
5bcRbAEjPYXHxf21QWvaEsV9oVTruStS4h2Cxbxrty5YfF2qEC6md+xwbEUIXxRa2xxdnYk12osN
bBwzhqvrRybYu115e+A4KumpYpkYCetmGqg6PRblFTMVI+HyhDC8rhG22qqfFc6VJC5vy471sskI
orYxt1OCQwuMtwn3UJDPqPmKcsdaG3+HLF29Dh3Ga/YeT/pG96lbotqt9ixR1U9bozzjrGg5u+R8
iyM6gsv0CB579lZvKIugPqRGRvfilE0WDzH01rxcQvG0wde4YjAhbq8dXv6fjhN6r7h0F5iswikP
ODPm3/CTkgCflJRLM0oJa4FcwWZEjUtKyCM68QnVn6nPfO974dYIklErRGTEn6oBjJ+dE24l6LPt
EmTZ1eUTZJBFY/UlNUN5w24zxS6ylEf3M5rQ8sRtXzGn872sq8Sp2MpvNn1JxIesayiOo3h9g+lZ
c3gLwFi7wtaZYwjXEsG+FPeMSKff4rRHEEAd7r5PsDOZItY5NNDUpWSeXSXmqa6jklEyAVs6uGaq
Wl5k54ZP6wnxlsNBlsb+zG4kAsHqG2uxh2tVXwWgK3fCoU/dq3y9vM8nb9RGR67aP4gQPmnihthu
BqyPj4C7BCpjXrGbPcHpPF/3pf9a4SH0NJOZ26mthpJaVHcH5P84ckdSOPxJPrcZIbhc7rGW+dHu
s/76PHS/nKIQrM+VLNakhmRA7Z/MopIt6Z+648Ka1IAjbVQHQsC/y3uQUsFvtTD3OYGMRjGyD44u
MMeDSIpOni63FwwxhsKlzBf3N4dQ028vdLbctQdt86RfZ8H72VFiKeWyMijOKLdRjVsu4sKXZtJq
4iLdmuRcrPddDwswTY7WBS27/pQXItNEAnmaiWaaBS6JjrLtqzO91D5aQwNIRUdW6x7cEEJkqsb7
QMCVHqudw++WTgJ5ZqGsB21gQ9gpGwq3icCLyvwFgtgJrmiaMqofK0uxbb/D8yVhpL+c02W4q4VJ
/8Pnm11YARrEKDk7IY6JMbgc7Gt3pz/XVQFz07Vc4MlOWkFQN6nJllflJxTG3sVqWNsZc0pCIYLx
IwE7T9+xZVwbLYKgzYZzPszCIGhFosT1ysXbA4AJ1ryjLOb4nfIkRkbSMURIX0TuGmnZ6ouzlqk/
GRFUJRk2Ahf4vGA0CxcoPJlJbgoVYiTRh6ImfXcabtXPKhQPTk53rm1Imjao2BTYXOyur7Po2lfm
SIZ4hbw/NgR/sK59Z1vMsSWmllfoBBMqufix1kbLjw1ImCWnvcO6PXwUwC899Hr60CzNC9cQmxcM
+Hznolg8ikbp4AQKHlcD16EK8KJ7szccxo7bjTzcZmgfrDbN026LMmBsU2nDe6XiFHv5aMFR6zBv
ZasouXfbvBIADF/ZfOAJ57ga111rPDmiX85aI4RidDvsbP/DaRwx7BLLXzxcQKCX9+9DNdV6EndA
v+1PwCHBzuOdMm/Iki2GfOVoIgc/P4JCjZYbssMlQg4WHzf3M2//eFMh1cm4TTDSTocmvA1gDDHJ
Lk+MlUcxLyzUOlLPtDoDPgPRcS7/dHz1xaKCK+Ws/rgYCuYlyP1UXkxnOvsNd2QkbDy+r20ckrtL
dUTq3NwC8znwNHw9KG1Kir0SOOny82ZDYcHCsMoB1DlDdZk7jVIBYggvC6/kKll1Nd/JsFfckzw6
BODWmDoIvqpFVvCHtI5nzu4O0EEmVw2ymIQIBQvNMdp0FL1xCJFAS0Ds4SVEzLpgbpIdFrSX2f7I
CDkTyzcY9GhN/BpyEQSn25qyMhIHDMaMtEZ38dtIFWmjLhaMDEmWRb/ohtGn5kfJUve8A9nyM0h3
zRvDVIhkVosmaioilpWt27vlCPbcZB2c6k2i7klxtMbytjeM39lYLyJ0w1Fj87rMaLFNGMKioshI
3AI0+TtJNrbS4/TjQv4ig88LH9+t7C99nNcAR4+vli8zDu+cC4MGAyNmn96OaUKg/T/daPzfiskM
AtttrazPpBmzb7/u7J1gy+/NBeoGHOwh78zl4nJtB+6OWo1WAn5eVEsjwp2kkrZUQA2yCvFK5lwr
pAkwL4Ub3S/GUPdCjOe2/qXpKej7u8/4oQcDqTFOOiZU8BjnVvCBsgIvrWzyUwZjaQ9/3PwwZkgl
Z9XmE8C4ihs6YIL8tR1fWvoiFz5oBY9YQ0mq7a2mJ/WxzmYkPRq0mFWYFNTiDoG6d/czGuT+lqeP
nCKSyiluQ6KDj5C476aXLe5BcgdLcL/syge02Ozevgr4pJU3unUn1+kmR9uskYegvRY+etGYEAVy
eFcci2FlLeq85nSc2xCpY83P5od5gUaAnq47xx7FGogPaaVJEdgo5M3FtLDv3DWhzaw1Q0PsaSXv
kFi4bfROu7ihdNiTCDTsLpV37RhVBOCjLSSz4Lru2BU+vhJlWjHhsm3Vhv73S0eVOvJYLLizftc9
T1bXkIzK9wEhQcD685KBjGPPkT0m5ECOcbCuh1gfoylvreh85Fe2HE0P96iesnd/3tq19IJWQRu5
9rWc+o2ou6U+xY4iVq35fDqqlW/Wc3akj7J+6hPq+DOHscX3VQzRxQObgD2+AjDYmlHL3tr3H9g9
/FTNi/rNHEycie0e3hkQEffxQKwRVptqDpZd2N0I/mtlLkmNs6slWSDJ0xLXLaQQK4yWefJ+cBAe
EJ7KVhqa1BhI0/5BASVXXJiWILs5aTSq5nZsisxKDutPL2b2uG4W0UTjLFVEithhgDnnRS8aL4XT
A0DJbm4pMaCprPGalXA3CNP2DSVn8R5+Tt73NfKqndZJE2+gW1yh+NRg78Bc8b+NkxirMJrmQEQn
Oi4Zc5w//SVJE3TGWzc7dCo+XzWG0IlyRSwBcGRbTw7jXRqJbeJNd9LJ96flQ3uWo2gOwWUUy09q
WftPpEDLLl6zP0pv3PxUHcIJ6PvsVQbJLncFO1OSSf7svXZPPbwKZrjr3GdlJN9T6Lju+/wHZiWW
CHsdYvNYf5JhKakl6N3tUHRgf3rQXkwReNe2OyJuRAjq74Pqh6UgQ1cQp6Oml7kxJQ9dh4GlZIhW
QQrfh6xhIS4y7eHwD9wbH0f44D+OfDuAOuRME/75eWu8kVcXoESPrRWaykyS0gy3sHu5gqlYxOxP
EyOYrQw09F0dr+dz5SJAJZTnV0OqUd2j66nNC92YHWLzMZiyke/OYlymF6R92wrQjBh9gS1G5AuI
ejqDa5jcOeYNNrWzQqWlapmGoEZ+ezWRuBLdhgP1+92fJRm8wM8fNCd0sK+MvH5dwqHaCrGjK8uz
5jSAq/VcrNv6aulMt3vkQwUiLCZ7EImdvzYNvF0ioPhsm4ZSCRvuxiqVC+CdN7QBCxFFx4KtPDTw
zMf9BuVCLRDeGCBRn3/EI0hCtd1m1tEmj314XCioHobVffPEPPNoastya0CvSzmN1ZNCL9xp+OIb
fiTS70xclWFj6QXTJb1P5qDcxiA/vlWdvDrujncH8yass/RkYSLQWRb4zQVl4Q8/QvTga5i3LS8E
gRYXecrEKKAvwS0d1P16xj27s5TPk7vMIehIm+NN2lvVwyDBiYPsauqffInCwUxQ88obkZMyzjc+
q/Yllv/tL4QYKT027TvrSuXI7t/DjixzkbRrT8QSXeXnX0sDCLva1tAs3D0ad9f0oDXdUTSXhL+B
pp3OjMABysDoCfmXmR1pZui0YqJmMnFJcXpMn2PFcMGo/HCARxQp4yq0c246YR84I4thKJjGK2Xl
J3QE1ZL412ib78WIQfHqmDsOX4yOGBOgf+shWbGGzMfNaMLF3vVDFCkAG8HAwLGFGW1YoOhThe2L
SA9ypLBtj2cZnqWw840fp1qwALzfRO8pbx8vFbvBi+NNlE/jfMW2msBUnTWJmAUAgkVIMpSa2gDy
PXeZ8UMXYoHHIEjPb938Wtel3vmTJohAk9xljcpl8eOo4ctnkMXINUTX6eKkgOX+LqqR9ByQuI+H
w9M5HhQafN5mAjYsEP882W4r7h/hYaCMQgDWX9gSeIutmzeYGxQ7HY+xRZkOXNuAI1hsI0txLgk/
MUMeRMb6OzB+E121/t2WpUO9LijXo6z2Vs8xaeqjH1h+4bd8JDtEfiKqe5WPEWenK9wi1gh3frJA
5MGKbU5Xr61N9SXhqWzUHwlvkXPjUe40I+QGUcnwXNxYt0WHyv4z8RO075VeMhXhRlTR9CIdlDLA
cqV9cnIbnNT9fHQgEl4f5jBPQdrPC6iWadT4vyjZSBpfL1YVl/GYU2v86o90+PLIYONNkb/ZoBBK
Vsaz7z93op1WQ3S/ercT6XyZoK8KHSQKdMWJzaq8EtPzGZCEt9AzFwB2niueAoaVQnGzHw3Qk0ro
MPPRKFvzK4OYFBWgEpTiPyMf0IMrsHC471R26RYINg6rgSN0VI6aJlyw92Ykj3C5ApAa4nOlIB80
ItT6+5dcWmPiuFZJ6qgqjP6b5As+7wU/qnavaom0A8LqZot2pMMiulAOB/tF7lAogIXWbtStnb9d
ICV+Hce32LTWYE8rRi8Zz1bEEzoVe2MU1rEni2TNyOSK0185CKAO2I0+EusWP0/9yxOgvwi7tM0n
m9GoCXdYZ02z4l+pv8F5Et9yLCdYpg2fwDwqhu4bN+DCxAtSAeHmx9nsKAcOGm8HdUOA4Yz5LijI
yVmO2HOqDeSCJ+it/zm70TgloSmp0gAb076soVkaIrGHOYmICKLlZJkeVcrGvIQ6aCLhmRYKxJZf
Qoyu1jG4k5uFueVhWWxXD1Is3douRC/73/Y9oWDKVRoI2PW2fwBWIaU5w9TQ05HECWUTZ3CA/DpH
sbQtAgaGfwwHqXQAKpfmK/RpZEDusjLajuDIXNscFVk8IJrtbotLCLygq87F+H9DZOClBoK20roq
I5bj4m5N+prdxec6HnYi6ln7AyiDGRs/UdYKyDA47gX0q340on/x00MZ5exGjIx4Wm0epYpjB0u/
MOvToxbXxv16dbdwaLnWdihR7wAj+SfmsyKXck6IvJSYCyPcFPrsPuyt1h/J5qePLWEQkPJemYrk
S2a/7KRQ8MacUt4hUhD43v1pP2iHReVCHWCxajGoxsNpIJN7bIlJhGqfHDLlFjVqv/5aHIgXmNu4
bdaK2QmKojyjDVT0vqd+2jhS56i7xnRpH7BIiwwEbQqMHoyfO/hWDdw/ERABdA52tRGdrw5VqyJ9
smiT+srRF4+Su4ATnH7bVXYk7hns6///9hGkN0i3rpkFqTECbZpr1IBClDgFpYziuLqJwS36dRQ5
M3EJFPXbiOdjOgMJYgz+bMVoOeE7cq20OuMvsihEXqmerga85ypEO/n6ls8rkfq6OBeoemJzppYc
S7Lc1bpMBpwojPzGGhrjL5Qplkx/w2XqGnyInBWFbVStA02LbMYf8n7B9NDJC+150cakvkqvJqQz
bxqRCA4PyINL7vVShb5VSr/QJA9aD1O1IvWviPWDgksSo0WGqU9BOBJ7tN2mErPBIT2opsEDc2dF
Ng/N2H6hHUNM77OW6gPwqod5q9zK5ogVNLMG5oJriLoCn0MwclR9JNAcLJiDdV5pyo0hkWjCJlZs
uVz2jDQ6hfQEoJdowZN+v38kI6C9x7i2pWHjXyqhG+Ym7w7Iio8X7SQZLxd5jNmB4vMQJtrvVlna
lYs7wLdzDaRdyt1K+ygEkWg9Q/i6gc6fxRMEFJvqotyxpxOmHfMKoHOU9TxwueetD32hQ3X4DC0R
ptJsyLmRJkrHRK0xl7lxXNlaOcNDBQ7D41ZuJ4LmCqfgCPjXM8SzwHdDbfeSie3WHgv03yfa/dPT
mydmi7HJj/55C+NJgQy/coKjd+HM39U96C4gbee2ZaTTgKu7sQ6kLjZydu4oiqe8r+EQnPCI1/34
YraPJrfsHcuZHih5Zw0AR1r39hMdz+GY0qDLdKNXcpN0X2Oj1pRNK5z/ucd0KrdUlZMQkNKEU/U8
7gcG1kUfo/p8RLG6eDhtwcCFMIsoNW+MU+QMM3Z3DbsEIHVfR3HfERfj5Ag/yZqn0EpKb3UUjv0u
tu3jwdbDkxD113I0+7MFVOZreY8A7uJJ6IFebBngHObuw8NxUnYqfh4rMUgcv/m2XgKmwq34gjBb
1YC/nVkSvPK6ypzQlhN1uzoHebJUkxj9uk+5UvTZqqyuB07V8Lq9hIOZlo/91QWuvdS5ImWGJYJz
8vpooTvIEcRuVykTGTbHgUB69SHs2YgooTKO4Th3IEYdPKg+g63Gq5EWLiREyw5KWvenelxBKqip
3NWwit4IoENE7GOJrdvyalkoVWZFFZfBleeUG6pVCPxhb1rcpZgRqfkjlvYeH+fL+cUMLs61TUdk
sEYt+IGhXh9VMmszPlFVNwxGJyv2HSM6w3OQ5WDIBTHz1ThqK/A5Ogh9kWe5OrcauMfwxt0OrCZ0
AYLjxdFl76SgdICmS/vn26So0poqitc9OCGnZZaybW176gQhzoLFrNm3t0xv8pkroxGDg4QvrWlQ
I2uycKlsjlg5h54s5ULmvGe4x+UJ9l5Pfnz8iyyiWPFK4K3HrPwJ4IDUQ17v3MsPo9ducODaEG8j
kTWG6WR6pEyrMy8PncBI57DvjjTmnbeLnV9+htMKEaIDVQmIjrEYVFRLWv6yn006Z/5iCQiROlkz
SYiyLBa29tUEOZtI2Dya5bIfVBtE5lm1D3qOJLugixBH6bfpRUu42lCy0pe3f2Z3SfhrAiPAB5HK
806tzDakNz5fyriLENZtXwDCLXjbULgq5CV8kcEjo86tWAWaIANHK36gcO3p8b0wA9hVDTfp1Xjt
ZfyOINQFRw/Xf9uNgvMZRycUL+G6lnzUOTY0nStTEkgOaCt0KfwVXddMls7jLazZRZ1Qky49Cg9F
0apnrvJSgUsbh43bYhq0TnDcQhQBA3bdAchFYvqGiAkOKtVQt/kKJtDxpN5XXIq2pMbLL3AomsuV
tZ1Ag+4MGUkpbH/d6p+r6NgtSWWJ3zxg+k3iecPuflqrPVV2NTAhZjVPE5fmLF2qJ+86vm5Qdt4K
uwkPcvGPW2q6ElA+yRXzd+MJnmk0H13f+1dWgQCYaUrtIkndVgHQ0yp6dpCJmNOSryQdKsqczY/m
dzanN2MDfR5+kD9WkVYhhVRaQDLH4kFeRwNY6cZFNqgQcyU5/5LSc8wBX+sUmyPtJiTBozPhjXLr
DK4ADO4qSS9GUxPAccGXCOGdkLdwlbmZ3C7tVnb5URF7PRKBcRl9+x/br33ciKhlS+3+CuSn86Zy
CCPetQjj6D89QyH3XPtiLxX7accrfvkr7uuccpoCkqRmG4eRKiza8Qj9gktVbXV2M3e7jwWTFEqh
VcpOdDDI55ypaha/mGGz7t0yrAZxMfhohQVd2Coy1xFNd/TW5SKQDAk8khqzCResPu601+EYKfjC
8sJoY7/H2W+aESof6ETQZ1VgR5Tk7AQtNJsMu7WMf5AUCmy7ZMQKjVo5Y4iPS1lehV1pu7k24ZtH
hZ6HqRmFbixrMGOwrRNHMWnoZ72T5KfewFgCkU2t3CsCAC1Gz9+lDAvZB/yytpyZhESfuLOhi4in
+OmCeR98GysQS2/iUHCI96YPMiKrrWsgW/75ieRIEqFlt2AkaSwbrfvJsB+hyF2U0hp8RXzrYIKF
i4CXYUkbuabeDFEgj/3xYMxAfBHOvd3EVQovsAUsAqEICRXDU2w/WdqXzARFivkU+2Cff5zVBF8c
bVc6xmM098jyZYrqmr9FEm/4k+HB4ALqxNHZVM+UFMe6CG66mRUNdbMdSPonVp2y4pbVz0a6XRCb
04O8uVUJRiM7Z04g4nNfigfbzYLFPYyx3VrAyICqatgPNB4UfjSbSVOra0671MEnUPJ6pDxX6IvF
mNTB1oZ+fKBrIc9UeZluwXW2skB+SMKetNh0s6Z8hGmDrvNmU21xkOSbWZlTHQb5smewyPZJeFBH
fmo3MfesRZvCDBXzgerxnOwOzZBG1kS2heLB1w24LLaDFwSn38wOPwdwdiZYq9yudleVgM35XNT/
tXSH5kNmp4zek6AgsPQcH4TRkB6cdwc++ost+PRlXmrRJkSWmy5c1cz9T21feYaNf4ZDDmSgG8AZ
ul0NgH3t2ltp2GNADCdimeXYyT8uAa1tD3WrWrfDH3F4WE7p3dO+R1jYw45au9lf0d67m9jO88m2
YQQh4qp4q9s366a8nD50zOW9879/ka4h4EcH938tM1m3ykwpnOhCpeAr0wBPjxgV1kuMUYGVlrI7
Dt7wlxQYn8Cygxs9XlSYzxjCeO6bLMeGRLdaUf2xDh10kRB7VHieBPoL3AR6rT6e9YrhopoQ/UKq
ApeegXdDuLWaxzl2f2d/ujPd22VYba6syt1MLSRQeXKw/hYsLG41mI7aGRYIhNIDehRPuGbP3axC
TfNNSWjSD4X6kpJqoQ6LqryZB3ZWiZhQR1PeE941UcOol+DPxpQOErGTTo2sK03Zln2TXV19PhvL
9naUdGjLxPCgT0BqX7jQDlumgq3aL47uHwkUyFwJ8nWGC3aikTY0RqLDHyXHzkqy9u/EVSAY5rnM
Wd5Ao+gRVE6cY1fPf9ouWBf7e7WgTR5xgCIo9IzLFxST/Eg76mBcOo5t5D3KK1GS6Vb6GXCQITvx
6Fod0UY70a32CkptkEXu8WiwfLP2+61RAGYX3kwzs9iR/mR0z/8q1EJPfEyoKqQpXE2XiD8PMFRS
/1SWqq2C11xY1PbuciNrDuba4rKabzo8i7WLSnQpndFWx52/gcgOOlT0Y7bJPK8WjCIN5BI3apsW
++jgipLqrEkyhPwFAHMeC4OgSMJeSyJQW7deVjrfGHzLEmRcRDv8Y8auqSQYsRrKnZDnU8px4xZe
PaEm4cOLr6jX+F34kM5X5ii0A8wDBKyjgiz5clMms91NIGrNOT1UFy8cIx4yQQX+4sDYSC2UMZOH
65f1aLRSeBi3S9WEeu4nTHqS8YlaAwjcjbw+F/Xn6j+kA6/B6hDr9N/9fSrs8iEPYJh5kDMhNsk4
+Qa+Jl4ornov5oKU086a3PWZcDcEqGQ8/yDVaGxN8JBvWWr82p4cpMAm0O/DRVZZFuqPq6Accb/a
NfGLJm4R1oBo2IENZTROoINb5342/Fsms8/Vtcr+Uk3NF95UJ2pgdET9PU9lZwWUd6umsapZtQ5j
+RnWAiQtE9wkm0ClN6GAwkr+yO3ycPoXmTUPH74KTD7WaXh4Z/qimGbjZhhibP4ucuhopQKD0Suq
2JqphyGLY1qCwNoEd2AHVl7lAHLLouBDXlSvyb+mK9Jz8F+dUxL93Ibdw1RLlUARaLEwUH42kLn4
oHxbe/oDNtgeMzIJGWjQUl090sXjANt/d2synk7IB0xjX0/31rXa7cPEKfMfy/C4ZbQ4LDE1wRy0
93c6YTuMfSjqR93qYVORWHVyTJ6CF/Um9tfLUA73Vm1zeWMVtz+beAFkw+TW/vdgu6w6toFrWAA8
73jDJRs4GB7L+V/2P96vDY78sUV6DL8Q/amagJ7jMd4+swpDMlRp3sAYl2pkRjRyiVbKtuwQV+M+
tsgYvkT8IJWx+jjzLKfPyj5qRkmzb2tJrQnx2FYO40jAlx2VJoL4HhIJZY4qfT09JxkkoKHu0Jx2
tPnvY4ETgDRPO7mgzVjFApI0UTp22B1gKaMu9ig8C91eVHC+tO6g691dJ4Rb/FQTSrDcyvV7be0D
8f7McQXjnSS2mC9VHCcDQBXw0iYRToM+Dk6lyGcUN0m7gSZmeVoheq7nSnqoKAuvhAv8HGzEvR7C
/UzqHzR3axhC36iDdqo7BGrgOIIvnDx861DkP2e7ssqB3oX4kfNgvt0hTqUxlHtd6WNmWWy89XdK
tPkGoqF+GBN7VYHGrleglOsy2TwtuzX5K4q5M/kaZ9VXb1uoFP9Sm+haIMCWnzDfmejeNHwx3xW3
oVFQCtERdV3bSOrccVK6OckJ8H/vl2/JmV2DCvtD1o1CIFfKeCxWep6budFJGlKKipppQt9W7VBh
Bp6uSHLhuwlBj6xZJ1yPpwcp22E1SU2+o9swBXnIrIlDDVWd8E5IByrD+lcnYgG9jdm2W8CcBQoU
pWk05afUYHkzKlsYvrO/di+MQwftCC6CaTTSwq7mwZLOZdU9FjJDI5CbbOVXnvybGTNmhx8UX4Lm
T827WwXtZwVj6Vauiwa5vfuBAp/lSngyrpurqoXP3s2+hEHkmAjbhC3kryX3Tx8sfS/lRNN+x8sl
DKK99o1sed4d4dMQjXgQRFdh6sVqUIbtuKI2MWm5TJL8pNAhSFEvNUTfBLTF5Psj1mjjE5FzxfSv
ovKVTsqq27SuhIXBLuoYhfVg9ZfJUM2lny2gkf8XnGNqSy/SnryBUtzbAgSE5meil75Y1/lFq7Y6
+qthdffnSA+b6o33yNb5pLXU01EZe4l+x9gRSYLvivZRcgLH15MniGYKjND66wIlG3FDo61bxrA+
W4qUunnWkmmvDbmvbsmK8GLPGSsKzusf4B0E2cK7sAKjervq156/qAYLXi/U5fMYCQwMEwvXnSlu
YHPjC/37uJpa2A2hO5Htr4+C8li1LuzhsJIuPMN8RAhS8pap8nMx0MAkpyuEaTsVXd9LYCz4oHKI
+2p6Q7upEiiOQvo1Eg2PrBv8OoqPm/q+Y6CFAsFIKJJM5WheSeNctoRlQWvzj5S1MwPBa89byWYb
0YeMMt+yoyc1Wm/yadNRR8REbHqaVG7t//hKmEaXkS+2u7iURyNMJn6PpTqCV1Rh4Odv1nWulZWT
6DyQrm+XU2G/qZ3KH78xvKrGOjsKnWfjcRWIPDaBYfVeQcXFL/dgdYLCTtATGxJ5PYi6P9JK+PNB
4bGT7b1xuYtYZnzRAj0lXIvj6tVX49XXGW80AGr5eypgabZ+UXsr+TYVa+1iNgWjkbLyEwGSDHZB
mwmb1ZOkucjvju+iQVXReIQTUow5eCfJJieS5CRO/a8Q8qDpz3BwY33XJl9o0PFPooN8apUXFJHz
14Nr/M2uO31ZwP8KnZss9RIwOqi9QtILWqf7z2PsDq5/XgX51HOHdQvrQe11bcbyUG5KA+9c3HpS
B9O1QUYk8C9BXV+6uOS+sCqkeJPqr3NvKU02+/iCod2969JR1oyeHigk4j8rnOYuhlciAUJDHT65
iRRF6vPB6nUyo7ihFKw8wwmUeKaaP9BHPMytk+1CfFZib2i4Q+Y6a4MMBY/NGcY5+kcbqg3bVYWD
uQfuj7IOywv7wCGQ+AkfSGMkvzQ1luRgpnV+RY0AO8FTFCtzVpWTnmjWWgxtCzcPLkfm/71MvJfg
Bxk0zJQhP3KUQYi8dVtD+EmfnsFO0uFW9/GtEfcOtpV1nFptiRxQXy+AFJ+dk05Wu+Mv93w4NSCe
FUN/y9D6DNbwx5LKwayLincEe0HPk1DlOIUZI+xSfoKCczEGo0mhmyHEBkp1OVUVRmu945b9fRWt
mxKbIYI3EzK+elH2r+psYKRDY1gbL27FYoWDkuOm+DkKNTHPj2g0VP90DlnSVRiAhurbETIJfyHb
UhI/opf5SKZZt6q7mz6gbe2IR8wLX7sile0LcFlRCMdrBPwjKi5lEfITvUtyOXe1iL2sPM88Pnon
ch5dEveZhVodYy60hpzV7/jqISsLO6fvEV68HKwH+Eork5fwMuZPUFqcNormYbEr0IkvN5fAIsgX
zDGsASdXChJ5DCufrWH6fLR55oiRQvAALi+90Nk8KMxgQJt95K8bb47p6CPk8H7CVDlT42uKnn8F
wkhx/jGhBi9OAYvaps0tNa4qq9dJp8CREmsO7l/A6qeR+Nbyvxrsh1pPdEmNVifztIDzi6gnAVAe
u50BWAMyULVadwXZs0dWpl4DhE5PlNeCscAAYJBWrH1TC7Yw71ghBGyqOkOvoHP66Zgz5GLqhYNW
7TrLbnATbiUpBerkjadG592MNGZla+WNAe5ezk92/7Oyatnqdg5ZDNkSzN3NlTWeCdRVkSo53Qdz
9u6j3n/IrX7afsVJrsCXzVscIkxdOgGblr5u6HzyzymXwvepr2yLbmZvi/c80pnAiR0xIjuXYZKw
RqBIqaPlMhan8n8x1TqBMvA2jMdzH9mfn21eoSNF7MnPxS/scN9slGA7Kn9XjBu2ExxEOqDt1bsW
7o/tsWF5R5W7MluFsZ3u4F/Q/+tAaTIBEuku0X2wKuJbdp3DhUU8G0zd2IUICVBBefaxCUO8Ompc
cYYFcuFRHLPrrFsSPGJytBZnWcPJ0HkmXYkspBccXn5KHoUNlffNG4zEkP3LkBR9a3ktexUbZLZz
VzQROrxxRlQe36N5X1YEf2K2wPjHVPeZ3oADGzl2pQIqFm+nbd/cA91+ucMAy1yqDNG3nJ3vpcXD
cH14xMqndehIJcbI2ktbt+TNnfcYsndU97l5ZOcosu9HDL4tbsvlVSM8bPxeDr12+q4nxAoAg+5a
IMsqlihoL41iNqRE80fL4lUaerZ6g/b+Tu+lyQgA5Ioho+kkqEq5aHxJPhAB/Y+zA4u5RF2vcWk8
TNlv0eDiba4Hm+6HMF4qNj1rUgAHXMDXbw1PcM+2s65lu2540LT8DFgqSyQh9azOadjSoSC+mO1K
foHvHwzb9IcRPL1R0mHp1kHULlUlEFtTIAgKXO/lREgS9lr6kMClejwrVQUEHuRyIyouj6VSoj7n
yYVO5ljUb+g0CS+iO55MY/2rQT6h/rkcWdFZTg82gvM+naUYbPIG7S4S0mnMg3riHti1dDQCox2R
M4RUgFzD0bpi/JyfYCjVkZargW7xURZ9ZvxZt9hl224zeaT/a/+FK9H7dw2BHbxVZ/SHSFbKZZwq
H0kzzvhuzI3IuBkDJXM8tbiDoNLwhywVaDpehdYNkKuIsv8aBs2spS+VSCwpUJKT78rj9kzxRfQS
zomhGNvRfEi/IZSe1oBitYKK4jvKSXV05Jk9AWgNiwXuV3BPp0ECsC+pemFB/m8JRnS8LkCfSyou
7uKJh5LH0vrpiRjp0bFD7pUHUprQ2z34Fpf+tJ4mGBAK7DP0ME32/AefQIXNnaD6/jk89zKeiLXi
Se/IlF/djyRVXLuTB4KHbAVu4alYXSOeF6CfLS0hSsEJv5d9tYhtVZyS54cRocxeLVMSpArm3o9V
v1JXbr5mc8MxEcFXbm5oJqCsdM7hOcs+B/AEFv1dVfFZlAwprvtgdl6/S5KogQEPrj8YM3ItvdA4
hKlNpZ5skQUEGZ+cFBFmtLeIQUSL7WThOpXolXW+3pP1ngQkxW0/jI/V5rHTTBrh+6utIqXiwocG
waSrxxlhvCVM5MO7kCXIRgAnelcA7voh53inkRGpO6QMyHVLI3c+2IhPTI4wjVPHBhI5ih3QAibB
+IQu00qimFz3dAiyIo4ESjtX1CVT4gpVb0dEvA+f58Pkr/ZM5S2wd6FPybmDUZwpkL95pe9vkDJh
su6gCS/QLZETZ+i3kwZvotKBwCRr8lBOLbnZas3zQy/dz1SKjOUri4N2N6/5hp4QDgs14KmGjUE1
5YzshoL1KKbF81Ih38WNqbgL6FXEBNQ061iFg8FNsnC7cbLsslagmy9p6xa1p7j8Rx8ZdvBdjnS7
XJ9hRhVzthsCdljXqTE/DS0OZ+Zc07ALRrXmaWCVenQh5TIxFmz0JGbE7gZqjypWbH6gsT/LYOgb
BgYeiEAlgtSdi8Gds0TWIMJkgTqMTp6ciAw2b2ImJ+VtI2C+PVtkKIpiTBac5C02N1pUQGGO7isU
DmgFBNY8vQP+Xsjl9c9knfxik3mP/hG+tJtwkOmXmmXS4BXip6kQlWiMjYdY3MrLMQh2TZqKLt1c
bmaQVKQhAWDnzGUXuSihmXyye1bXO5zG8wdFOz/CimiZM9XJ6SL7EhfWHglOvMu3pNaZScVzy8Fk
VEXQhXEw7lj3mTPurOasCkmtq4RGAUcpPrwQeajTwjMZwZjpT9R2Y1+c/Lvwtnfmdaaq2gJeqk4V
MdYKWP3MODmrVVrSIDlDc93h72KiVSvQwuTjk/XWezzuvB7/nolxGshqYRRpgQcGCYgX85QkrGyQ
m16Qdgpmhuaow4/cXUkJy1PaMJoou1WVfHdBbWdsP0nVcrpFm1Et5xS/3Rk9vtQL8Jjqo9UwF69F
ar3TzKzEuLv5e0ZzhXN/9zrCr3cO7frdwxo4Kj3F4TzOkRd3GiZSK/9NVpQ37xWxCHMQ5ZCwRRbV
bRX7C66lqM8EkWm2IveotrvIMgJN3N6elkuAXTbGaPduUZeuMGwbYgyUzsJ0/dHv0kDzMERELnS6
95GCHm5lQ42rnYyu6ZgCMNxy0G7I8hvzlyPARsnYbtvUmfl+4AlqF4ZBmUY8bsbeGkW2O8/ufW6/
T0TQF3kh44orReUBBLvjTHaP4ztPDy4b0lk8CXfZsJNoVuqg08GQRYsKuHzTnHF6qXoBwOl9AfUT
fiBqctvgPGoLupuoxVG6o48T20NTDpYzyOfKorfiP9uGD+79175T3rehIxED7Fyxx/Pkka/EblDp
WMeNzv8fSv+z2WfNFtJ+5kPvjk6klt04TDTZLG4jZNjGjr3YYEKgOvGNr85pL3QgYXdiQAgQc2wh
iQxb/TClkO+YQvn8L6c60I27CR9FVMpxEGjyb4qdJkhIeEv9dVDbSVtYlYeHCDb5wwV0xLZKpkcm
hsJdUh+MjJ0n6lg46rjQHtSVK6d0XYwFkEDhWJ2voH5WD7BM96gEwT1u84kSSlHuc2D0OEBIY9pM
KYjy+IJrpIF+cXig1Dnqxkm0W/uKDi+o4zfkbAaZjUi37v5ZJPHUGx9hgbbFdIgtHrkP1yyGMuS6
v+3kyKt+4f156rSK5JdHQLP/PLJ3c0zexE5BWHm9u7bkbpWB3PxhJUH98f+ifhyBubpPu1Aodtc0
qfCrCN4QG96jtQre7nlgcFmHsW9eu5j51cl5soTY74OR5ubK+jadVETr9xeRyLoMFAzUWaeXgA0P
SUkc1d8EHya3IBMsvYhqwhUel26g5iQ6eBnW6fAz6DqM87iboK0cm0Kqf2wQi8SkbV4lkYfhKunx
GFda1AEhNoWNu1Wxk8/cqk9XVw2xqDBfoUYDznzkMgXNGGBnfjxWjr6r+rcG0Ds9J1wcnHWu8U7U
0MQGUTjySvNiT7JFO6112vd3fqDihHwAytndM6V4oN3L0J3U7txffxR6tNPwZSDbl8RjYZVSoMNb
2LOi2HRTpw7LtPgAlp1FFBvwOCg0/9a6P+eNbJuoSoxBVTXAXhxUd2OOzqYTitT/AU/4bttVqo6T
a17N8xijQL1SXGGgzqFBZ6zlBol7xT5P0R9nZb/fJKYM3uE0/fRYdZf2K76cj2+g8eI4VmmP3v8Y
1TZ8r2AlOQKVtwL/mAbKvkPIwYN5tR2NjAyTBVKUFg4TYWYW/RNZJqwhorv7xn75u8qs5eA7ztMq
15qfQ5mYclaTTaNBodQl7PQEAfDDP9d7lWKGJ9LIr+GbmBQfIQz4k3rYApolLBSfPa5c1d+bQ8PX
VDNdNQTILNdaflaqMfgn1xPr3prb3OEqrYpq9ABRL3rMzoalkbvA+097tfHdeLMZmNGB+TOX4Ghl
PjTFWTmTYNryQEpTv3h1nWp+aKkEPl0iwul5p1QEc/MbQgHmgn2Ths6IHyrtnbW8b6ozY0XETEIH
6Igtr5GsZLW7t1yIqAQmVisiz1VEcUt0Bn8mAMVWW0gf2cmNJZczsiHJ/9CsTOs5c+mMwZzjquS7
DjGTbIYt/1HCkKn7qa66VVQtxmkxECvfZN/SLeh7l1RaRYX5lUPqTuOI5Ya3YIDGC1dLcjtRkT+C
LjFgVOKntXafcj0fcsn4Y1yVmVZDtrO5CLqJambxaQZvABHZRKeCmOqOJDkA2GXVVAn8CUDgFMNO
eQPdr8F0bwyFAoqZtk9KIRlqS4t2cf0zCGahK/SVd+MsNyAf0lPhgIrOu7zH/vVub4xZ4X5WY2gP
YqIBnl7tUUXjECUu+JA2svTqJbeNyO3Q5u8bDpYbh0tNas8rX5uXglUB+7Zvf4HcYfQmBJtK43j1
RppSp+ICzZsAqNgP2H0buSSoGg0HpKBw2IFwPmaYFZTIgZVBcHPzx/8H88L+KFepVgJA5btbE02+
OiloI/+WFsUa1h3jBx4Man5R+eWJ9hZGUi4YNf0e4HKjXBJ4OM2+BnsbPp4ElrhrGBzsQ+Kw/er8
XvceKXrx9AUDmU59sRyIUThOG36LMXDlR63gKFxWwlmbU0szkuyCC7m66ltP53g5XRD5lv2FVlKN
YoSpAj92jXkcOwF05L9E/H2FfPaIF5qblgUGq5lyqUASYOO1eRdpQnwEUNkG++jQ8uMfIlOwPh5F
d84dXTGTi4QxAnrRo1jlXnPTaJVbAD93wM60P0C/9FDkCVPw7JS7IQEebMcGzZywLUlZFMQj5dd2
0+4dHkuK8AzajLrWNnEtnENtDlmPZUbhZitZIAPVlQypz9/LdulRcIrSLFD6+27KGnOFXFb+zndW
IBa9Xmc6804AwbFesRB6H8yAEeq1rxMCvPqkuRWySdbq3/ulWdj4zq78N3RfU36dmcJCu7QCCBZZ
KTkQQm/aH6G5Thub5BJaGhVvgLGUB9/Wsx8OcjPF7Gv1Uq/7ZHE+ZEoirjyjLOYWkhu6Nf6IuFE+
CmFzMkgEnoA4YibDrAwzXIN3nWTa6qUVfzifp3nrvmVNrr37ajKckxny0juBjaywUfYHAee9JAg9
d7daGPV+4MeQISYHho1fmqYPO+Bb3Ivxxnmh1vCtkaZDwFXIJ22wGjubeX+62QJiWGgsM3SSbuyH
6gZFF2JCdVPXg/2P0tJ7RWhRMAgAdp+UUmMiF7Kgn0flQ43ldONtZvIDQzGLVCU+F+2mfUR//uas
Pw0iuMxqxuYPLeiJAgQ6WKq3B8PVo+7eHlbY6kV/6Mvdo6g7Uth8SeKtjexsMgt6cWoxdmQpx05S
36yGqwYz0Dqlfz/j/zkp4QRqypXCjJuWhVFbuA9e49MSFdIdVVFxJ/pHrN3s+ZTtsYKjbB6fFWNp
hdV3enQPxrYzX0RNWkyqhh/jkYc7/QqmKmSaTTbn7M+ZWLcxVaD2ofGnSsmu7wB8AuuaEqLyiq31
cCy1keZM2Y61zbgBke0eIGfxqEl4ep68z22utPhT38MIeg+rT/ZtZbxf0y6xpycfJF0nN3h2zEbo
lEwiPizJjP0M/zSr5Dvkj52cSbPvocZxvwXzoTWU31pNLQap4FA6yQWLfWhJ7tdeE8fMy1EWpk0P
+CUYxWjFyhSXZu2t7aRvT+a2cuZQYb25DQ5Yp274mrSK5EyHBfIH2McwpyilnhobLgPr88uu2OWo
aoUrJ7e3FjTvM/wVjVnUaKscDeaWEiZC8OAhiWldVq91bjZ1CpsBL3YiBuIc0WgXxE3pEwJoqOV5
5eiB8QCMlC1xiKmtvsT1lLzlPnE6Qc1ZvFjI0yN+RAdx72g/hkYYTsTFhPaq9/BM4GhsUw6RBI+A
fKjt5iuOK11/jHnuWwJzbpUxQXJXA0sYh6XxupC6RkElMiEa9TF4HJ8zMxPBGduGcshi/4d4W+sV
+VLEHykjLjCv9vmqnU0na+XjSV5oKX7Vi7WNU0AkdIIdLgjhyrNdYC7x+Ui+17dCLtO6dvzuidCW
MEiVi8H2+aeHfcp6BZApNZj2QeTiywJy08pgI+kygXsHZj4S8Z/4iu5N+K+UzYbjswc+yRg16YZc
mWgtZHpCxrigmxdfkzywcEQ1yYrBbWcgSEJN27YwATz+98XX9sLTFLq08vtO6duHUa57j8Kg0JsS
+MU+QbwYCHWsVUOjKCwxmUnCBv62RIVurUa95O4knRI8+uJDOEpYf15M6FO8TVcZBhdZOkF66nFj
rwCYmcdvcI/rFIntARfEgutqXK9Pu0suQthEEBnsz32vmyN3cYxyFZGrC/i6JydzCE60zVieRuBd
HAaY3TmTaLzR22vXCUyEZgvvox1AK86JXSKMVx7pCs9GBoQnrJ/EOwZn3B4G16B4HasOKC/FQGRw
iwkL043fX1jBJ4SARz44YhMtBP0fXlTs5F+eLxgKN1JXf2yMcopOsv9hWV/aXVXfd7bKWPdeZoLy
z5m4Jxrj3IZL5xVw9mxCvgFL8ACEaUZ2VG0tFvO/ylUOgZZEgQDfJtqDCqSfSftu48kPJor4TA7U
ubPiiCW4b03ah10HpC+pVVLhvpQGbCfR5JEa5FCbdeUnJ6/Sf8Qnw2oyMUkpkE+PKrlTkx+VP/3W
u0pFetzBsL/Q6WtwhGhkLeChe1Tzk6XMgELHOuYOIrQwrrVRZHdKDzXfEk7pQb1QKS+DpiVCETqA
4mUZy1pMStoCzTQrf6RctLGW+s3GNc4Xp3NecZQ4S/1tDZYT4DBdsRe2m+Z6bHM0YJQStWif0M2d
JyiT4DOtwYtwsSYGdP8XwE9gSn1OiaIWfUCMDCAUh1fJ1frUGpDsqoSVnVrTGyTrSGmOQeSXTB2o
qeP4ad0+Euq5Xc2rCZ9Tie1wlkI23Z24D+RK5LBkVizO1OTvguYfnmfOZA00HE3FuxW3t/v3g1HD
sE+3QhIwhwGpI5gOqMeY8zX+N8bvIHFnKuhMCihicKvWj0BqDkFVEXpbHJTFbYemTbNr/L9Iy/we
CVmWYJFluwnjbdMtvyb7OU+TuC9eKd9SRMQDtv+6dgsQjCJ9iKR2eB43Y/tuQ3/iu1luF8CTDK2m
ayjmTHn9owM4ZySKOcMzXt5PE6sxPX0WyqCkfQjXfdUMtEMW1QbpaIGlpZEfI0DRBhMopeSK6DSg
xrRusqKpz3hrgLJ6opttHTkkDkCP+6gNJJBDH4tDZ1NO7CJUnG1p9ZuFD/VS8OfRXe74pR/5qcXR
hhsVBYQYDwZE+ArHX1usCBvOXmOuBM3oqdII76BtqL8R7G9ZrfoQj2Cw5adLpYvLBYn5PIPpen6c
8WRXG23NVUND3l9vHuS0inGTm2G6y2bqAOLDXTCk3Fq4WDeUtDBU93R7deDBPFQbE35rH5NxCDVk
oxDDJfYpDwXRNZt+rUKTc8CassUGtdelL7sqfx/isokkJyrvBJbasFsoJPMZn6yRJT6zpHnw+pwf
1EDtdmoq92uUZ1EherdtU0pFq7/5BDf1rEpvrXjqlWpeMkOpcNttZyd4OzipWQ3FZzqF0cUHB/2t
EiZ3MsWg+w2ab1eQZglBZA2CzYIS0PfYG0inNYC2FbnSABA/xHpYQhdlaOXQoOCDvkCI19CP3LdO
Ofit3v0v4PsbkagmdpVS5pfp1T+NAf5K03EW7SKCPhrnt/63LWsFvGCNwTn0FmTYn22LHxLIr25o
C2BRpbkGTZ2jBfBh9LpsifjtA4kbhs41FiYvr0dwA9mleS1OOQuppmgFZBrYeCSc1xsly809bVTU
ALCIvEuNYmHQPiN3UG0oUDLJHYPdw38d/Uu/Fao8nLKIPX7Fkuz9enj6WUbyzTeLUal6c55k3iBz
XeF6LUw8ZQLbQM9tTLGnUmpJkkd1t2REC+ZZ7YHRjPEsL0wadih5L3p4fRDkRlw7XWrTPnVe21At
q8Rmwk4VwFGD5BlJU5HpaN4UDr386SL0UL5GEl0GJe+7vVH6LWLhZGjGSVSfHWEj+u8pm/chOb6k
Pa4UpUJDzTSv30BFR39agbRx5dv8xBatIutje1nGV/aj/iwyDezexVf5TFLB/LQ/ZX8YK5krEsZY
q5Z2gywXQb12F7RYZ0OjxlSRMsdm5hv2smcTL6YPDohcPFpT3EdhG6Ms88U/VSUhmvPQ3Brnry1s
P23YGxN7eTvqcK9D7P/BJ2Pu+RH+XWdWrMUkIHYAdMwUKEcX4C9omRdOKyTBVEvRd/cq0SphUlh4
dBeOLu3BhYguohTyf4t5fqe5g78fg947sK5K5ovMtUEgqUzLHwc6M9aeV3HD3rAt59zUifHli5Ek
LZnf9xpU4W19p/gAA+zH7m7bWaViWgc79hF/K+PZgUSt2WsxOGwdQyRfasGaPdaUVZSoj+IdPICN
2lxf8JRT7fp6CrqxPF6UBCvfv3qV9nJMx1Msm528qzjOWmUzX5Y1VPNn+5XJKjK9YhVAgQ+Tgpnk
D3F9NrNkjMM03Z2sBCCLzhh5ey6fOdOyDFbIAIFk0/TP5ehl0TygAcxg96uRltIEW/T2zp4/06av
3ZiwO1Sistbuoh2TS83j+fo/d5XRIp9T0egOryEYE4jlLvKT/0FQ62VABhr4+i/W1de9tjHCKTWP
cV90WazmPv8JPndNb2WTXooDyzJPYOy/hE1Qv3X27Yfm2S/0vLz8hAeNmNAC3fKH5xOdJhApnmEy
c0CrbjLy2Do/M+SPeb4oUAcpFKoIJ8gABQvXfNobzpmf7QuoMzt4rrUNXHxpLSWESWQOpKkYu46F
1RXjPBT1sXnXpRq569NLaJPK+fQ6gwGZXqZ975shvXjUg/WnfICkqEtD+cVovVcxsUdBo5gtui/7
mtmLZhwWPNSk19H03+rz911PbiNZ9u2aHQsGxttsvqsG5DH7eNi8UvfAqEhAZEgDNL3hpciyWwpX
xtwnPOF35XuGFk4q6h4p6qQOYoY7zEJH1Qiqh4NbN1zWlXwbIaTNUi6OnY1SeWkzkSqmFPGmPgBT
alN9g82OrZTrUiayX2DvI2U7XCAYdX31MtBZjeTAT68WQh4wwldSRpCd4ZWCzbvlieu4qk54o65j
REQHzirOQ+Xb2RiQxGHpNxfx/FP3nnemjzDjmxOjX0VRMsRuRyzq6+/toKQ8UT9aIf8kfW7wPXI5
AunpO1DVjUpFFAjS3Azcio5U70+ODZg4QNHktOOgfwzU7MTW+msMOvMqr/tGOBgv+0MvZ0ISP92Q
FQRkTPxXVJQo9v6yA4S6HBeirIeW4zHbVY9R8zBc2M2q4YTVfJ0Y0hXlet0szN9Eo7qUwAFyCBJS
UMN2tNav38DZb2WpzfbbGH38pgdcMGUd2DY3tccKe7mTZFTkwi42MKYG0jMRXWq55aynC6nO7t9g
BvB8qbivnxA3r/yrbho3egn5WP32n3CwqtHNKf4L7DmzXdQ/98kiBy6XIvJUD1LmXsoXrm6EghVY
HZWaJ3dFy7QbAn4co2SfNbHBGoksZxVFeOefN6VgBzFJ7Rea4tWDQ9vZkie1vSwU2myZNLRzJLXs
7wiNDI+Vf+JcdvX5pJi3tk33beUs/b9UXK1EfTPjgFhOMXCeDqiyQ4hqmUHSYJseGXR6f5vvqYql
W07zA1Cu++75kfBcFwfQUcT0SbPmieF91pJA3g0EsXIZf1Y/eR7xzew9xkaoG+FSVLhEPAx9Ek7K
SZXKY9C6Lw15jt9Yl0Aid20F2aYwb2bup3e5m/PpOH5hGDayToa8lNJmV+dexXVCigY1LvBW3okA
Y2kQ67GjqMJWKQLga5DRJaPk82252aoxIcvkI9nOUJe+NJSxitXlXDa/t57w9PA2CfBsVX+wCL/4
85CIwqO89JkiTUQjUZKoKfI/InFYtMCJdlrFdSIwlqZJiwuQEHxucbnGSC2aJBz1LyVvr27U017q
1Dhape4GTiz9Q1cdQ3TXJUTVhRdwfDGxaufGDNs7cOZ/IwY8XIYH6uSG0urVAV0X1t7WHBoKnsZy
2ZMQ4U5lQVu/Wrfqx0HXjyArtZYYGvTEBbPrkbUpMldgkw6H3Cwd5qfLiqIetdGnqD5/6R1O1y+W
SwFf1WQkynkxfEjoO/1GdS1iDzQ7BwY43OI8rPcFYdqL0Uw5lsfb6/5x0SZdfwrw92kOcC56182p
WAbd9dcRVZ0cCoybGo0vwzsRUsT97I+HYIS8yjUkGt/4wcAX0ganoWJ8onyjTafYhyMQscMSaUTa
k38+EG8Raw0Ci8eRn+q0cOBdwZaNf4WyQsEzaNkOhIF0fOc6zHHNgWUyPtz65bUp8/HttM939cLm
m7w/AZmnyOQVKOSkTs0UuhHOXWHPSGlFcUEX7rhRFRAeSE3qukw4AIZhEd3ryEx2OS+bq6v1MVLR
uYEmFXTPhiNNxel5+pg06wpP9Sy+n75xvTl7/O4cPo1kmaxLIdCPYfXo4NsOVoHx/sgr9z1ohfVq
TlHUk1PFpgCqrDHrGantf47/yXrqBVw4Rh2ObVoFX0T/qwhm1Qz2V0myI6FoVqdM+D/bAy+x7U6W
EtMgzYgJrm1wuH9ZY3+tzvpN3s6shmEoCeus52Ivti88GKRUxDOrrmWQom9vEU9H4CN3qnIlyTsj
esAx36BuP8S5ll1Thn/Ykfw/E1PIJ3zeH2cZzzJXld1uNkm1/sH11ijzPBmSDurtVH+TJhpUdUm3
2eJMilBF5PipIxgzj7oe6m5+BcdB7+bI5ABk953X+tjpmhSA6jL4uf7hzGkHnuE2G7vkjSGTS02x
1T7L7mvnzN7l3DCV3t0khfTcMugSvHLngYHQGezKhsyZQskgBWxpA7MLB+mTfUo+VVzwo3D6hD6j
6nacO+r5XstX6Bbn4M1LOkTHAgYU24foOkI9EPjE7/7vSx80a4shG90ZeoyQq/nIzq18gTSB0bn2
noLRn5OlnwYVJGoTrC7ODMp6kMfeDsz3pp1dxD7logh4OgbsKuvuFdsf0zF72TaaGOqFjqhHExrP
lg2mLx6xdRFuYS/ZRTmrJ0RhLYalCDiEdmdO25uvAMbKVkeCu3OMX7F1/LLKO3xQmD5N0J6nKgFy
Z9MwoFk+GCGZaKxekqQPYGpVyURAFseO7xG+2qAXhomvkgGyjfC/keA8oK9/Fts8UWT6/gvWfWsz
4awRgkrKSqhf4FOtj7UUQQdCQ2OWvF/YV8FZwW7VnwE9vOnIE+62DBZqbncJiiRGv3QTI7AVE5m4
rkUwI2O8XmcQy7QId8sV8MPSmF8HOkgXStxDJf/kiPrtaNWp/U+wL0QDy/YrAlfHEEaAfkMRHXkg
AamW9eDPYI+gwHst0KQhEoyUXRxJk2T3h+TagcfkRSWZW6sM7S6v2S4OWf+pbJlEt+A62r4jWW1G
Tr6vdckV65kTU6PfjcusuF+jGksSy2WB39LGY3ej2pOklvU3ZdFxic0UOdanqraM7u5md8IU88yp
4Oi2TD+c4bf3fFBfSbFXtlSA4Ruy3kvUiXEUamjNiPx5maAezsL6AgWOitCyfjszs0wcu5UVJjr1
4D8FHZt/yCU5UTGtJYi+p83w6jp+rHihv3u+fh0eduI3A/1JBAJPyzsDcbWg0hcTJjSrlz6fl2V5
MNvFj4v3QlPi/FxbXDSrCgr8N5VsTkpbRr1t0guwzH66eA5qQnA3K8BvFPKOIhRqAH5Fyj4PgC5f
AFUzhzivTmTWmJRZtbPHqvhOGGXTOE+jxhCAz0m3Z0kHVJqDiEH/U8BL60Afe8SFAokWXujRlZAi
qKdRmlGT927XUSm4Qo+vY8ioIbkMDnfZFWKIH8VSI91rT01ojolfF+tRMAk5NeQmt0uRcijGnb+7
YpcUh7EzMnzwJ/bMKl/+khlz1MaS9ByzwthSkAV+gqTRZl4RVY14BlvUxyN+6Wb9HZm4j0HJ0Epk
hxDrO0qUv+R2rHoX7BHqZyCBedn6Gn8avMLSYAqSrLfwm1yoVDpFcng4dMrHPpxmScin8KtEkVz3
IaB0tjVdPPLbQSDKLxwCMiMTeydLwhqxqi0BbiS8MYWVEboAMrSVy9+RfrzMYBJLWK3vGJBUi17/
InXXQ9FMm0A2ijkHcm3//SyJWRJsPuUUa49yAPL/WoJkHsPhS0VKu8535IEsTO/wog3JNm85MNMp
dE2sOrCpGqlvzJcu7X63N455IT2eb8L0J0nnsuKUZpRzJuS9nYEAD/PdxDj29QpOnHVdq+KBqu0Y
V1Mqott7vj0I/3o979x24RHyaGQFTxRkEcXWQ1i1UlE3tOBz7LPCCvKgmqn3XPXEmsWuMLVoPtLs
mi3n/j57VIH2+DdaMIpJHEr4gOk7+ZnQ+wG2H6AGsuuilkn6NZZxybqQZxuBF5oaSIti3tvIHEnQ
t60MCy4moJecyYoZXOzRtUilCMNRrG2FjrbrGnesnlHjkTAYr72EkBvhnMZBvDJ8s2P+5/wRCgHf
mlgvTkjv/+5XtLsWV9UE7MUN08sPG5ePtXAut00X+HKyq3XpepjTGpoGQkTASG82+DB6TT6FXrgh
GWTkSRTOZ66v30S/AOdgOo/m/CRs5g6eUwMeaPRorZrL3MzGegJlm27ngoQcw8jZYLYjLqdmmF0e
RWDV2DriVjPVxI6qG4xisF6svz4mksOJhlU9ne3+in7OzlPtsqqqvszG/mIqcpJYUQNAa3yi+xK+
QK09yLnpg+r2wDmiP47il/0Nrx6zP01ROgZM+vkOlY+/DBtD3r+fvE3lwLBuA3F1w7PkAnWaf1L+
h1DVWpWPmhxKcs+i20sHzYc2IvgAAa4cpKvMlElYLr3+giGzxqPUcjzCB+94RYRHztBcDC5IuxPW
SK1rBz0siRr9XmrIgJPodm/zxfgnc+32dzd5byjV8HvWjxVMcs1xZlTrIn8QfImLOwIBGOquX5G/
sIKmnr28AdQUBWbdCYn9GH5aogZcrSygIszKusz9t0vTuLXq5V+onCBI7jrPz88FCS1lKUsSJ6M1
C/R014C0jPAQcrYqZbdm7nOMGL1svm1UUEpX0KNlOA1lNGHw4fYKc6GqE3xMbrXoDfq6NUBwqaWT
pLCqQYW8ObWegoypWymYXFx4iADes/9yjm6W1T6JdGjQWx5MPENamW6hteFk7SshZa/P570SU15X
OfLPXB2nZK3WPD05ngzhCVl2uUWcRXcTi1udTR+mldpiAjK9KSMjjVy+5LN0LiZkX1vUWIYgwOMT
7A8po3UPZN53+XXgHeGnBsOKyqu8o4Fczzla6CUYGdhAxuO3h0fvMXmsQIc2q6fo4lH9ldjegmQW
yaDAlsk+a0dw7csjZtoU6gIgq4/BSaxmoBqglM3sqX5GzsyCHVu6e/oVLJDE073yI6JRBjgjDRIo
3gr2kq5mVd2JSqEQlm1TVCGx+v0L8Aoykbc351+Sa9gpKmUWjWRWcUUww0zwLYqZImLGdcf/rv52
bW26RxX+t2tQmZEhjKLYt8/T45dPar+NiZQ7Xo3d6h/rMuDe+c8krOhpY4o3tFEgR1yFqDiurnN2
4m2lp4qyi+gncDTf54CAxkqVjNk92C4MU092Wng2A7y8M6Syy4RoEbdRMBAdMFVfelsUUHmh51JS
IdhrdaTl9FRgA5GEUcOvvWyt2HyvuDgNukhH2qXNLR7RyksHrVKvp+95OAcal7vxmcW2EsSAPrW+
VaeHsVMNRc5R72d1IpAJwnovdQEU4L3DQHNLtY/nMht7BfEBQXQLMbxZnxaeO/O9SKdP/hYwofqE
YeMpv84k53e+onh7RxwkhvGRmPXk4dP1MmlAO+wAV5PsiSAPY2L+qiQcS4LdcIk42YaHA/0554/H
D1ssUof3bo1/gfszbcCgeNFfBQt2yuJr14Om+OF7LAqRRPkEs/dw3M/SugWKD9sD3unB4Sc0mPhZ
TxOINKfyTVFIFidh97QKUdkQ1n5lITOeZInGXgh7dh5XkpkQAygvj+Djm7w5MP9g7JPQPP213wwS
Y7/CHjRomcyLixKQYvmRomE5hfAmQCdTJxc67Adek+GfRqRG2znOagfLHcWFKqH5bezavjnZQS6Z
yZXLbxLIqTheW+P4E1nejkJHc7spYA75LN+ouJcXNJz3UItojHvYazxKgzJvazjXV0XqsPfU/v/X
kjkKDU2dPX8xnmwtvKNREYlx5bmNHKMY9C1osdSUbvMvzXwyq8IVt4q3WXYkPbDLzpE6WM6NnMs3
tVgGOhacMJcnf66s21lK+Eph3sgVrBIlAzM+MQWq0USgRcSEVM3LgwrnyN5Jzsw+YBf7yltIOURn
b3IngBWeAZEEzqUD6vdsOts2Hn3b1zo/ppOH2WZnF6TFKBbKZcH7nqfOs6R9kUr0ox2VMu2aMmj+
H7ipdfAnVqUadSV/nZ61dvqvM3O1zbkm2isBtn/zG/W9ShzG32dJ7+i9yEFP/1sZ2ivHxfiGZzy1
fCjEg3VBXbWr2qKxux+AjAHd+rcup3Ff2CabXt6T1z5PMQwKW9ZCEqoTxoBlFiVJl63EWdhgqoR0
Dd3mR+Wa1SaEExslIc1rM4eTcF+GHopjZmN7G+5MEJVq8LWrlwoElgd5Uz+AtmZ8VyZqQPzqaOC1
qlBMJqR20BpSgvUtmfnkGfBMsyTHzmCXgL6KQOwizeMrMcs8dTfYsUZRT4EMjAHBiGnsKvPAtMOh
qwXncRnNZZ4b43xTQpxfWGbkw8EJxPq9ZuU2INJIEdjGznN16uEcQJcX0mDgo4HNcrqgiBqnW8NE
JgPeBi2B8Zn4/XA+Ojkhmb0yrGKek6Djbj7KrOacMNJbyqDqCWI/JiaH894ZfqyojYq+Utu9F/+Z
US6dzvTvc/9jrAJAFGj0OgYttry6pTx/4RnuDr1FLP3eYMzN+PoJzLeP8DgDTh9p+qowAy4q6GW2
C6EH4m1MyLLSbAUyReGrRM8uFl4KMD1bZNs3b4fokZRsAYFU7MH0L2L92C/ewHKGoSFF1pi35f7K
K4aNPZyvA8iLTqyw520RMwSecoMzixKnoV4xqs4LEhVeDt4D27Zd0fVBkBi2rKz/cUIlr7U2pDFX
7tiEujQVSTWDd2bcUKys7sVysqsbfnxUpAzUvjsfrV8c4YpQnvPioCIGROYvOw8aBGTWvLq09Zlz
ghItxib1FKboUBx+naVLgMppvhmVQjUGgR5V0m5o4J7H97F3LH01YqEd9XqoUTuVmhBJAYANEImU
Gni1wn+smLM3zMMPMuqaed9Fm6cSrYnVTFYj7mVJGokuhR0gTpac2vT0v0oNyD9uzKMCsWBm98SE
IVVDz9Nsjg41aAw+KSD/zqvaB3a8XU9r90M1xC+DpHEeE+oRC5TfvjEj0+oPC8aM3jkR3OIgr/+/
/BI47YErLRbS04pBfz682Goro98IF1og4ABd9pWJQEbGcdaiTJGx0kP3m1yVRL0lm2VDzCkLJQL4
HMII3/kua1k1BG6bsn0MN5EhpUKZFvM4J2Ty7YBTeGTRqWbpmBCQNLVJhzdzmJbS9CFSADBlzWH4
JU5j5VDffFN1f8/dIXPBbmnewpxWvl3A/qkxY2jxHJ9tvTMqtzEmy9LdAabX/3nsuWLT+WNBouxz
79oU8IKdAQ+nyUHILqCwNsEKSkMGmrtk1N4SyprXUGJUL/o+Gf4wHfypdsFfYdNYVtXSi6oOoz6z
jTnbQp9RkmAyaT3+5vFTm/zPM+F6SBpjx66F/72uTyEenWFeUZHXL6+hY5qbFhwslv/5zLyO0C4f
TwLOKCwaj4S4eCYMhz1x4bOMH2HjkcGbry5CF/QEFhT9tR8g634FGLsMwogY+xET35TDGI//6Q+5
VoqtIk/YlmvhhPFujsGFy8iWlt3iudw3aPGSkVOiiKhgBjhX/hWu+qJjRRgkGuoBKbllr/YdpFXC
59mdSTbsh1uNIIVvDxuwS5P6W/SMnwxKMb9/fCa2lUWHKCFnpsY3jSPu8QMhTNwde5ir+dkvaj7D
YXP8oNRMFdkVbv7S4+BGxp6uN+qmDmdXLpB9wk1g+6cpSsYVSxoBjcKXZ3lbIfZOR/a1q9zGu96Q
hE8t3jia7D5OhS0FBelw31w4+XBUV+rFJ0U7y0Cm70R3k6m4kllJ1mIHP2pAGJ9BJoCS2vvH0S0l
QPMbPjmhvkZT1L+POWhTU4GNWUj799k2w0umzL1eh+j35Uk28jY9cSQgoLCkZYxudiGpH27FrcMq
hT6EK/yGC7Oxev+Tt/Qboemeu8A2SLeyCQkalrgVbYVHYw1e3DIuLO4YykB8Yur3CQPWqm99l+Lo
B46IGOQxklcRfwBSpvohGJYRfKGU7qvl+Gvg2NWbH7ifEzVV5je6aK+IB/UtBYtZgdL04KAz/XBi
oEZ3iPkGXR2B4xTTWcG/C1ORDLpKiUEstS2v4igxj5G8Bl2oW1RG28hJJPiedvhGS9HB805Zus01
ahJCt67VbKF3f8WrszpsGkOwJpG0zloLybMzpzTzbe39D7cIx0KDUhTZ4S3Rp0GFJrUd8iJmUnpZ
fzGsgPIWwD+QQcfO4mDXwKn0eae/ej/L+0Zti+WJBFXnb4R/kaExTgQNz3bSBdeoxDmcS63J07Mh
xI0IIXYHbSeowGuCyGyH6WRPMo/QRHkKzN+m5amVd3Pybvir3Y0b1FTnpXtWTEdfLLmLztu0AIZ1
mJLQFXySeBRNJoexxR//JaZvpswrRXbmo9HxUBx5kiUZVjYFJdA4ZarMGiGcVXMUI9H7V5WVQt8N
FF5E4FtolhBde+WyN1YOkLIcvqSjx7ZkRmYqSdKZh405hmknpfEskLgdaeyh0W0VwJT4MQNwoNC1
RPRzHadSivDq6BIa/R8kkv83OzdiwryPVooDLOFnf/BFB5meaKy52XFhdUdmXezbPrHBcOuLWBUN
FpB60ekrwJZGMubbvECVM92KH2YYG/nNFCGZHYNkV0utD45qXa9FxtqK0a7liZQm5i9T6YCwiEKD
eX04xWL/mhR3u9PPObFeHfmzUixwWJoj2+h22DQlH9VNfr9CD4u5yqiyr2qQOIOjM5aHDCnKb6vL
NZ43aVbxj+ciFSaiYAgJW5JxVb9Yx4mtxb9ErNxDbVDKtd46vQaWwjSjECmvn2PZCBPKAG7oWi6r
qEJZXgLVSzoHrkLzrcF8HqmA/6wA6In/ZhOMQBeIYvy66oQMGySSn863eOj5WN7WE9vLHnKcNpGL
Hcbs5mTun/CFG0L0d5eBtFQtmHRvMayzbuWqg1MchTTB6Hljl/jtEt69tYVX+1gUoG3AWg7W+WiU
gX7+x6iB2wu+t9gG9c3+IilY2NkcoQQfSVlX8AdR30RELY+WV3X1RsZKjQbm4C9dvZFIg8vFg7KM
gpuAYds3j6ynaHDgAsg/WzXDa/WhydEvyakawrl34LD8j6GrAbkF0FOm832H8xcLeEsSmtyleMYy
UR4L6sDhtUTJBD6lv2C82PxOUVASykAL6y32QIq7kehHGaSoW9e8U3X5S1BoN+4zjIN2ozx9uVmX
94ObJpvPT7AsG5Jknb9S3csAnXNkGouvb55eNVVRI26ZfpDCLcFuXqCAQwHpmnFABJLeqbDvQ/LR
M0Q2hIJSNHrbHPRJy5je3izkI1ohqqNNej87SsSC1oDpzaRQOjSE+b4WuzhUSqK6HDuwe21XkjZe
hlZupYndNoOeexI9c+wxAvCuGc/hL8QHn8stbDoCoUwEu8VpuQyyzUPyOcK0vZyOQ4nR1z/6e+1w
qkq+GDwiBYvLl5LUSsHbhTm8hVnekzZbrndE0EUZE2oXqiJ1Ttj75MbLyE//1h/tbPfFj0nbm8wQ
Q5rmOaY8XCGSHSvcCZDuRSv4vBBb83GG16X2YuE7JmX47k1YrSQni6/4HvOy/72vPqfx+yt+K3TW
Tg/TiH1u6t2MbfFxy5uGcP+HkSo6dPNuZnAWFSa04yineCB8+Sa/3XP8hGa5uBIMmqdCZt3H3dPc
HhOF1RyhZglD4+MZx5rKRy2D61Sw5mz+/KvZq43ROodQ4IOo1/3CNgkyoeX9pue84v3QI5xPfnG4
aB2Orcw8Dv7GQxg0PB7FO4NF8t6zK5xCECdQyrMlKpes4/v+tn7D4qqU6LE+9yNdGSBXQd24r+f/
xIfzWuiwV0uDgi4FB6f9ydbQegKI0sgWWTeQlEC6ktuLBWAP+IjdpWFiTKC8nr36cgxSKwndEYtz
w600wODIKvip4ojOTCVLmqwT1G2tzbNmtZHhHnQzZhTKrIS+v3VwfgolKB2Nb/tfop26FY8JDlOi
Qvjl3dTwftZQdtYDZxXlfBwT6VMj+2thefSPI8HxCoX+KQFxZq4yJrnR/jWgEvsCJC2FTCBEVuGk
7Td5zwNHSOU2qDibDFdbE/DfeJjxqtG/44Zo1wGJk4uwAIfrGTN0UKv2lp7OQx1KG74gJWafB0a9
CukDt7lveS3Z5GXO5coh9UPGT/Lqqm2uW4DGfVMad1CXPrKYjPsRW3EWqbhI1wn8WXC3W7JLVZmS
N/NxPJXtrdnMl2RFAuqyYQkEkhun2jtWkPhWsT+KBPDtBYO054fXuI5Js31P8ZIAXCVHZP/n1yGx
mTI/dgOfyEgQ8awL0ljN0NLU9BeHCfysKOZKQE3Y3phCFR5WKZflpjTDcmrCUNGfh53gK+5skjio
5hhXVVBFlgqoB0dJtdSr34/OMq6Ue5bbAxZaKwHF9MHTO2wy5mefZSEzmtLprd2R2TpU8iyBOOdM
rN/7MhLwIJK8E8pDAU3a6YOo9kqhJI9J1s4C8dRHsQNDS98e9gVt8oC6BwABxVpQflCaDt54DSn8
NphWlBTICb4CpNgo4yYdVBrhz9MB2yO1BVgYU80DK5HID9/Bf1IJ1xPJXJH95Bosz7MWTWBLdlu4
EwqPLrUftF4woslmX/13eSvHOypGUBPgRhQu+oKqv3CEKcCSuxsfJpLfVosUoQdtC83BbrkDI2mg
lIyyxpyVibB434HclHYAIK39herFFo1KMHC5ytGKIYudUAQQRKY3fZoM3497l4AEp6SFxXvYnLMY
wr6jGwXfmDqyTI8pIw4m/75AZdCxC+MN4PnrprWh3T+XCmaiYqHfZ8MzZfJhMK2mewH6VJSUtpaG
tvWwH1QGuj5MVTdeXc+1bjGve49Obm9X07amHxhCkslxP+8wYZHnZYbJMscUVSXXJi4U9RPLV609
WMeFxlJKn43XLrg8+43/+D+80/pcNaVVq7p6JNuCKXACL8U4vOBXmXbhfIzy1edtijOXbDk6t4bX
FiDhPi/q0T0oApiFmA0eekeARhoGUF/Aw9PiHjYHAsuzrPVa+2h9c6Ms9PqQJGONaCH4sWkDrNbg
QfbMZMGAApHaEBGWku0EA3YULdrfccksrI3mqY97eqjQX+s0Juv3VQzWjuHlyrd23xtO/g2Tkdf2
CCcF0mqJY5VEdQZnArh2vfLtTMAMLOUx+JfKnz+6pOtqS8x1SMVSw2eH8ebWz6td1RDsuTQN1pLU
Cu8hYcc90Bm+du2J15y8v7nfTUsobSla0niDW1qJwAJoXnmaEHA4RighOisF1JzCnhnQcizWJtil
vVvlTVUXcHNo5vLNmH1a54abj3Y2t+CctFM2+q0Rd5hub0mi4luEyJ3ZjVV618ueJtgXWLP3fY7O
OPf08AL3vlmoF3JR+DiQCWEX3WgbSGLTKJna4wevT+IwfDHn9L1J7fLODhTzAyzYyTBJB4zHnNs1
gPQJiVOBaUSThERYBPhzCa94tfrJ0Uo2b9hWkFqeI2TqlhTi6HpxgbvthIV2Kndejwws8RIRMrkv
dNQReORwWziYI7kdB0MY8aG1uvyekM8q2otzQ27F32dYXKJacTasRFcWdAo+Kv5yQell3LWUgcBi
vqR6q1BZX/yLAaRjfU7Kd35vlAq+VlYMWl0ZGLd+LVl1O5FDZp6dsOXVmMgIbJXHlrmUaMZRB0ER
cp/I2iWE7oOOQDrfnQFYaCO9LJFdW2uChxD7HbJ2OI13IGuisvXe5kZmK+Ur2ut5zXRwHmLvuuP/
h4bHq1RgxhgAH5+bThnuXf9yBp5HD3ZcJslAAPn4v9KvO2sEGTwKsNtPNcT6VOuE1SC2j6xVqNlq
/aQGC09Z+AvJViM1C3w+6lXDUbYvO/QmGqNTG2HyH72KKzsuYT0eS396o+iOWiL9g2SM3aiFbknW
9hoTn7cuwBfg/tJO6+XLx8QYtnjE1WHRS+PSFanKMejO7lQxQdoOUT/PdD0z0TX6FgQWn1K/fuk+
6UzYRVIP4i5mEFpD5epbmfG422fJKd1QcpvJIy8m35IIXCc/OkITIVbN0RqVR//yVEqy9FEQ5F8q
1l1CzdIX53dgrhJWwXez3JqfdEtB5N44NO2UomuWyz54SJIRjbHsDSM9U+RtIl77GAWhrtiYA1q2
+qbhdGAzwRi6DHlIlWr3/yN4HxgKvCxfMuHW8tr4mViqq9OEELWX885FJxNRvi4dlamMUALtgHYJ
405SHDP8FsAanwuKu4bIeVhQwmW+s2EqXWhslYK3oH6ngCWh/2DO1+7DzdZ9m5+3cjFe2pFFGDRj
0T4LKxJZttvVC5+SCKeo71L3Xyfh6BONiM8px82FKh7x1MLapJnzvY5dB13v3Ia53tZ48KvHUB4w
iCj5IQQVAOZnePc35DNpxRBt2mdgrrSIbdiDMc1jvYu/j+oc16RConswrE7BeFbwP+WDv/L8kq7d
ZGk0MQ+ONpkaDGvm2/NSrlhcQtcTXbNfIPwEA8zHBcZDBSM6CS0hsHJ6lwuZuuckWwLT8k9d6oXX
gQO4fprKVpKTrTAE63Gj0CaopON7Yj5Kc3ij2HzDvbQWnPV4SHWRsoMABN0fge4xEjdcrutNRxgf
J0IMZpeilOtF+5HP3iaJfeOb00qh8p6wssX77gzX9Xz8gg+EYGNieh75VS4tynNbOxoa9mroZZOS
Sr7V1vPCE6kn3VHsIOBI1vLeFEsOfXfl6bbtaVzV+DpvgnLL3ZsUNwKGl41Gyux5aoGXphGr+NJ1
RS9bdMRGVjY6FHnXvdgkyUQt2WHffTqdOL6dceIktqS4IzZ5a/lIO5V1O5X+MciOKhBLUkRqlltW
Uv6GgKS8wV0n1D2vi3mvqEoLxmoJ6NqgVFYivnv+n6YWkan07nu0a8soVmrYJKzFLPRc+usatkmR
NxRsSvpUQrm5BaJc0Yiw/u6HVnSa3aOGQU91qgm/S90xb0IxdgQT157lUYpwU7QqCvdOWTnpfO2n
dh7nL3TMnK8rAa01Kkst08P0k+Izz510KOrxtiqWBIXiQjjWcWHZagfQx6t1QZIRy8BP65lH4geo
uvqOV6ov0EN4WLMAtNvdC+9tDKpycMa9VWQOaEHd0kJRQsWaSDNNp8NrayoZj/UE1XE6HKBXaJrG
9ky4Y2vS7YxIZZZjb31X3J3S56DH9EZPPi+iE9QIm4Zh1/5YEuIoo1afZVKVxzaJOGGPtI768uZx
QlB7EfFi5hlzsWeVu7ht06DVo2LVHZLNMR9cAEQgFxrwrcJI3SQWkAk0j317Z/D6VXILnuqzO+BU
hG5NiU1ogpON+Sy87w0RxNVp8gytTfD5/bwYjffsy9ZKiJoOy7P/qvdZJxVivYbyXJVU6vxQzHlO
9SnjIco+LZozDUsMCQZiS52aTNDJfMo4PGRzS0LWufXRXztgUpx9CX1AZ5IorBopY8voIahzylf4
xfxY7GCbGx+QKqYpu1AHc+8452kOezr0Egt6sXcZi71Tfak5oQu+6eQkfSXSTB5o7EKZiLsYtuR1
++2BnZYG005uCVQGXlTJznz+xcVABpc2EN+CfIETrz2b/9Q72YWSDdhx+2Y0cH5rFv7fOt0Qg7t/
WjWzdgDQ0ze50Ouf0zyBy+elT7oXq0ipBBdUgMiO9ZRbSq74fsxgNfThr7420qEEn5VD4Ej/KpJ+
6niC5HwfcxeGJp9EQx95V5FihL5uxRHg5KoykpaQurd5UOsyi0g/+SqzddFrj6JAN4egbM3UFlEH
NeqgcDHuV+ImEPi7I1JD5iOeRgehb3KPo250zyUFzqiw6Ctiyo607Fr15UlgWT6a5aXUhpOvmniL
nF9szeNoCfHyZOX3aDqCP8NN528wzvWdw+/3NpEZxb6SLZzmucgOyLRgDlKN27P9UC9jlI8cVoIX
6sd0jwLjOdbUQgwFE3WkwUVxgqsqVTGyaCmYHQ2Ytb/P2c4oWUKlQE/EyHab1WyXwMGVUaTrHd7r
VFsDjZHttsxvOOfEu29Xk6wROqh28pU9gInLh04K5mljoi5Xr+BeVSZTgVfgfTpAkMsvZqSHRHSa
ir1AW7cAQD0yVM2xmdpUtG8c1pbLUruxcDTydwDpsLycTIQzKAgfTDSCkGGCe4s1jjvZYmbmgkoH
rul7RCr5G/vLhADgBobMbwGnb+ux05CwZIQFEbxn7xt17wV+vDV5Mt+ihmT7rnKipvW2ZfiQthIb
OKBcGcsCtsBbHarjjszWEwBtDxACgybD0w0JgZT3rWG1qNUAXwSVANq+i6AebwgEW13B/T/e23F7
MR79m39rvhIMPIg9PYWvRKUzSRYxcsHVFxapl5JLxXPJnNZ+0/4y6EGtQ9Qi/0b2FRcOjDrObdlJ
5yBINjDh5ZUyKn9+MwhVPvQVw4XmTgPP/6yiq3D6jnQQD4vtYf+389cjRXc0LHcoKbhhFIdVQEbz
+aHW7R3+UFqcMyYL7LbJi/u/574zq6psMCOb063LaRNQkStjNRYkh3QValjKGf79dQQ53WalYN7R
HkSETyCImMH4W3EIFH7QKWpdSXBZ0byptpH106JvSADfHm8l87/NOajEa5Ib6V7vpmYxwwPZ0Bqa
FQV+Ik58/Dcpyhnr+3JYpmSPTfWrr9RkI19eTPp7eGPs/SFapng5AMeSF4wQzA62dTNZKXltCToP
oojLF+NaS6/It9rOcl8WWn/ddVqJEEpCIITXu0vk0dTTFnf0WXv7HQcBuKTKI+EG4DP8BWFx8kL5
o8WJZaFbj5i9PSaZinhircLwXzst3fFO/Bd5oqp3Wd4XH+tjw/7AIlzCcHL+Ab0oRtLAyNLCp2Qf
+Rle/AF+uieFeSSSoU1YwASW5oEespe+2dsjAOugmUHOWa57SoT499SSb5+zoGXebXfU+hkvYqJY
zrV5Gs0nSCaIICvn2d75xM/WT4Vpk9Lput5na2OHhsdd7yTqYgbl4tdsYasxFyvases7BkFZDel4
nFxR0xWtD6km19RObZ5PcZqmVA1HzqqPDId1pwgER6zJxVs1n5uvTUrGCxcf9gff0WHFo8L1aGyh
DDcoso3yg/2kbJ/iB13OzCSoK9OlLhs4DuDwpDHyRo3zg3+YxwoLGk8L+ob4Efq/TIJJXTZCOlz6
uDwti+98mNFqSG18fOjZVWVo/QpUGEFqlfo8t7sEZd2B7ACD2VU2WutONTWsf+bCvdITCbaoIe/4
cXbut2HFdH9InIVRD5ZNka44qRdgSpbLCnwLzUl/j1dHELDdXmNrFpNgupi64dCMKAcKo/vPpwUW
0Gx7Uuw2o2d6E3Gvv/5tCavvm6sraAocJ6vX8GwTC8xaIjrySVlASTs3VuCUWHqBxNjBk8fJ9q8j
ewMOfcehQpofz+4yDH5qyKgD6Xdr5WZ0FF3WoeAOH4cJUu/Mckvz9JgfTrmOMfpA3eNyv9D4pPHD
UCrUvvmQuwNL2ywOGFdsKtIDzkCQIXuMvneaYE4fIbm+m0KZxAL3pHZOLubrftaXkSLqGTTqjb9W
pNmL6gRWadiDafao+z8anlzl385FSRYivsF+s0LYfxGLcM8U0dSvdyYjzTk82iIGlH1vL0FPavVL
ykXGrUm7joGBl/WqD/3vod5RoKpHKpbCKgrFiwICQO/3SSouamXyqJqGqHQAw3ZMRbLfUDEimHbr
FoCvULyUpsa7ba9fuIVypSjJHH6qezm3gnVwjFp+biTBxK95EVxiY3dv0svPX3ji7EjG3pgzmAl6
Qh7ZnjP203/FoB7TceorZ7oQHj1x6FSaOwC9Dz5C7NZ1bSXP+GedkGcp6j/Xc3irXprRS+3Qcyv8
jN21JHXdA9zXnGalK+eycqY5sdsUZ/anttIbEb1MukuL9KaKg5nv1R4Mmj3HsV6qhmjLmDFEjM6E
SitQTkCubCIVHrzQYcMTv00XnbW+UWxIuHGposLhxny1DQ8rkJ25ty8CcI3XBgi840yB7AWSp17S
/3QpCr3r364xtT8m2izog/gkf7OVkwmgP7S59K67bZUDBNgoQXFYZqSY+MFQKSjClbobHHehgXx4
EehtUImFXuZIUA2U8mD7BBdim8BMaxPnXo2gPWr0qlv71rNz2/eg8SptLpWFUcuNE7mkmHOe0JxD
9k34HaCCNogFUrvs1A0x1NBICIoA+f0rvf/5fmo1UITauynR3g8YlkmUrzYlVbEwtnmF1A1A0q4+
jRquv+STPWD4df1JnG8JjRqmUzMAoKpfCIvaN+m/Ya9Hxo/wxJQ3EElopfqKN61MyueeTKUk79Fz
Aj508JSM69gGK7V4krWrLwmmg8wmT9z9UqO5UHau7GR+cXr0VXRqvi2kHTp+FYVhRdkNdRvxNj5E
Kgbsuo3f2BO/uxGTOuieFKurJ41kFSYtuD+9l5LFTHTQEF6NNEga778cm66IPADK4NO8IlX+NtPJ
JL/uNujSxaupmngD5/KC2KlLDmxs5OS0OIepFDI10cRfaBoie0l3mYXixTkPkVUCR4e/41HhCdDK
krte+jHb4xaAorJfXIz2dr08B/7ZC7vUVIswKKb/QIFBsdlaiOtq9scGgToBrble4xj4NiHhovoh
qYCjLbs0oWuYNEAbMHLCN9RbrNUnPVuJqQmn3+5LYdb+dFQcA4j4e0Ui/NcpXpwr0lf+6Fqo7BdZ
vOPA5yfEEwnp29D4FBmxWW8mDnY6FMeFM4X3PHD1AySgJuZCVwtO3VBVFN43++2mldTdAEajoRKx
NhYQSzgVal5QVxebRVOBQN3YR/XjquAVJfP6tNb+JJA4zUT5uM+jUML+1bPeg9usnz+3/iMrbAgT
XlZ/NdwLxvIRj7bqwDmBq1/YZujVWvfLvydqnghzxRq0gOcn63pEw8eVhB6lSwI28wBNR1xM2azp
mBT9xN74axJzJbuHLZENVFJGNJtWuzBYbo0foI3POpP2VZX78AlLT9V5mTuzigdv+MCtb7Rr6sdo
Tpbbdu/hwnhp5AANWn8meYRqiz/qKQutoT5FMDb9BdyCTQZhuYDIJdgaZSiiWTzZeWwD4kUJyv0z
HlnVNsSI5qVwZMZ5DQ5JAIBZtf0tpqtP7goNZ5vbgn3Xz6VwHSqUuJejA4kINoVn4sOZcBKB9nJl
cjr4ZodVMZQ0gj//4GJS2O19md7KEzyT39iaZ27/5DNnV4IqyWx6y+m0k+Cop8fBjsWst68rClOO
Kq7A+xQ53G+tCAup2fMEjwG1g2+EkjpKJ5kHdnJkT+KY/acBMNZ6yaPXzfFtwUG341n7a4ktVQVG
PXb83YN323IPOvgePnqczfREdFcKOenn5fMhRllbLVAzeio8D7XYafnXOgm0GsUseVrhXRDP73mS
QYZl7D/A1oTA4oKIdX3ysH9JTyrI4u+/73Qq1A4OxoLVgO+zXVZ4mGxLwyjUp1bVyufqUhlft0a6
0DmWu6FmoBRpy+NgVkM43chznJf7evMGbrl55Ox0mHdAcKxUOYLInlYbj/qm47rT4/pdqanVs4up
D1FI+++fcnhTy4Rce4w+NaaEWIHForWJ/l5IzIsWjmtQPXaEgzkVt1/0q2HLYneFOfDYyqeEzQYP
qwVr+RMPYbV6SF7a3LZYwQCPmuR3Wx/TE+IGEUefMRNZOvSXhQKuUVl79ZifZ4GrRVz8lty/ZI+S
FkH8G8lcXiTLe48CSAYOy7apNu5osKtN4R+MtfmNjHkUMpw80/veQifCBfzmzQAksoD34WCajOIV
8bDA6V7KMbOBai21nvv7cwBgRDBB0vW/gdf+ED5bWF3FaV8jTTRYTyZkEcy+2YBVwxS2gNBsvlx9
Cd9fijs9mD5bv0+HDiw0uCHw6GnAuLa+qsx+uffSQG/25/tfUk/LhSfL62Sk9xuVOqmuuKy6pgTg
4VQlGholRq4H/06QO4bM/ypHZMkC7xF5XjVKoUfj7EMKqmDBCMJA6RQHrHZSKfAejJjM2JMVRyVB
Wt7SpD5YTDCsKdCZNf0G8/0tCf+EYrOtcKrYoSl3KXItlT5P76a1srWE5nokDvFiICz339w/MBxI
63qMcXVhNC3R/sac7pl8VxHG0jzGVFpx4mY7dxb+3AR3kdqdp9/kv68jGXJOnEdcQ8g9+L0BtV5D
RXE8PSrThJkYpIMkBKw/wPRvE4qcfnht4vA5wA8+T16bxHXFQiDQGKRdFYPU4D01netmAx2SwkS7
QV9ao6+eyx5AmAObgdoN1nLGzvofkkCJObTYLvuGudjQ6Ehg/+91GRGm0JbrvOHVQmBUZo+DHXNJ
/3k7SwvEJZqPjSxAlPvREbtOnH4LduQZI3PenDsDTAJiyr1282j/47alleyRO12GcU1Y92U9KIHx
PLLjmtTmwXkoHDZreRCB/btj2YqRkP88X5nFGj+I62of+d8E5m4h/BHA+kDGks9dpZwRntNPfge8
ecgvdokExLyRzKwe6zf3rK9t+mSK7m9cBiNKRFefb7hTcmqSP1jfcrwIvTPSbKIj5jaA0lD6OuyB
FuisWDiZgRbyV41JvLPShtg0CzsjjFU4tlOwr2oodEKFsaJ3xyCkyqj8de6L3KLUxfRiN0v5yc7s
H7nJNF9QFxMO4eg3pmDxScHKR1Bku2EAA2szMon4gPhIsE5x23drqTao/C1KFlOF8RkxTlU8pjCe
Jsj+2XQx+1XtkbZjTttz9Ho/y9k8PwbAubSdFSDeYm8PSOWiJm4ijgrbz4eP+WcYZNKEPIyrg8yU
/U9nZnCNDiSwOFVtSZFAHJBbUQnEQl80ALZR8baH79/gi+ZufVtnaEdlu7QDAqFm0A5wke5wgM3R
CkOE6mVQetpkZQm6sdtHZoK7TF8TTCG3ZnNZYdbQ8DUyII0a5OqzxS6tkxL0BVZgHCz0rpxguJE5
EQriXBWGvXGCcbRPf8xNHvVwtZco6RMFajpCeUppeAlR9BW8C580wizJv9hbVkVTPOEW1eS9sTaf
Jh9wJNpt8zprMI78ZfvVw4s6+/ZOj/MGQv7v2CoUi6Yn/S/Fep9CJCjppKK2PpnNK9B9OcPkC8EP
78Q0WQViIhHq5g7U1/8EsjqcIFiTzmHQqhIhi/9wO6swEOowW64D6+4o3xjU+kmsfnCgHg+BaW9r
wjD4HZ/07A6D2OSDK4YcxBC8E8MUDyR50KvPDoQBrTbSzzMAXP8luY4z1KWAv9h/I9jgbkjFxyBZ
rHvTp0VT12lGUqZwfbzNeen36lfDa1F7XjtTmEwqbX8UhTXNrMF0fbuCDQCq26MZumCkayyGv5Sw
Bl8ktELKF7Z4sB35HiLVW8W6geu61ATPfRotXHrX+VqR8Ce3FZmO9RgGJHZAs8d+qQgRk0QWgTmR
QLrFDdwAS9ehS3XAcJIRlhnG2sHXFIVDu4i1/MrjXmFmor72Irqznj04DzZdMxbwqBckE3a2A17l
GIuc7m5F8QoRdCdBZRSplUS23d0juRwr9ncmAms/J2Obd7WoizMZ5/p7U61VQS+bsEpDOfCIKxr6
gUYHSDBl4XDI7idk8vzNHpexXkRIoaDcreu/UaWXSjhh7tf7rKfbS54OGQWi4yvInlhM/W3hRJAn
gBMPqeKZUxjC9l5KppPAZwERvgIV0whX+94XwL1x3tDtIhFV5tMR41+1pj4OeKOrCix62nqQ/15s
0Fk+lwRYfOfS2SIubC87Kzx/00VgroLtcOqksPQW93e7inznMjuLdMWnbXv8X/naOknmXQb9Rw6j
NkwYUL37MPkwbvQp0JhsvyqvQx8b6T6EjyomTDyTP9LwjZlWozNmnFHTk3qsy/yDWuASt/ABnRD0
1y7PM6ke89M1MlNbtMjdRjFkRW7aakqY3mRrPMMCJ9EsVD4c3Rz70tHtzhGnvu1FLo8zaiDDdV7A
vyIEb60hWYiNp19oYExEqIFd+pU7qMZ7o+d5PQme3yOeGu3cuo2xGf3dvLXQmzVz8Uq52MObYoCM
CNqvfXYF0ydEjNx8z1ZuMOB0iBLsIZ6dXXnnVIhbnmd1xTuTq5x73z03k3uRY7PI1o19kcZtv3eo
uquUkR7Wpjyp6U5Xzq6bteIRONsmhlySkDUCEKS5TD+bnQmwK9zu/5TdYUlTJuSr7B0CQz0KeNIT
uxLGd/A6mm4oXzA4gs7TUvzjU9RAWuaYZfWSiwU1/cHqRs+pY8gXO4sGCHavp7jUvZc4ZrbKhJgB
O26mbTMZ6OReyAcYpNLE+JAMDxrj2JWg/8j59Hv35dxJ0I1uIBeQH4+uD+u8TE0vjLmo2adlhHHa
YyfOKgRkt+UprgwOyFnRaCl4/CDp0HzEvrS/x3aWIGtCGlAEfGyFlG/ZutPAApPZ/ABFDbciiZ68
0Aq+7z0LKZER+siBzILry9MThwI53Y8QQ0xyI6tN3QuodjkguTqEHplMZ6JyF2ES5tkq898p3EPF
VwbCVI6WJqRRtxAvZVSZKxTvq0qvmR7JVHlVjsDK/OMmZEMW1d1ro78FICITQ7S6iN6fjr8YN4FZ
VPhHBnJJdS9cejcGhsfjKJmZ3vBdK2HHdzdp0Hs50xTGimzlCxwvyEcft38+9oCMdQct005t5nVJ
Ps90+QLKztttTVZkC1pH4e/LvQ1Y1KY+Vv7dCWIiKqx6Yavu2JnuqcPnDM+LClLWnlTBoObyeIrd
R9GUWL9bhQACSGyicP6HFPCdYuiUIdiqtNknMggmtq5AEGEhkbOkZrfHIy2E/ID2x4NwcTb5MMtw
VMlonHhSzkIxvLVjiatRI0Mu/yCefkla+I1J3Mi36X017XG9J+nivipFheYN7VrJJRsZIxrqSDKz
RUqbvCoFnH9znLa66xp3J6k+p3HQxQ4g0WrnrE2u85NoqSN103CubaChcphJ00z4V4i2uAi4X9gX
4bfR0wm8XSeSj+v85Ko2tqxxgNAnGywhtDAqIuhmN6s2aMtclUDVIVKh9L9p9Wt8S2SKawBKAVjt
L0WdIJh1x/1jq73hrbKjsYPh+RbCtGClNzR3OWfYunwv62xgs9R5j6j893yQ27NeJgDyGinZ6AqU
qAaxtejyV3Zpvwfuse2qPozUD2zeShzNtzby2/oCs7Jnz9dZJyrx64GnfrvDwOOiG7lp2DGzsrAp
t4tY3Nt6YzKD+S83+f1ueVxzjMOenXLMU2/2W7iEQioTKIU1AIn/qJOAbzX6rBXOBDzI//BGjtia
cPEWHZC2WZtnt0zLadxNiAoG+CKdNeymr9pzZpBG4Ij6aujCWBGzT0MIVyzKSZzKD+cL6XI+6e39
CO5S8XblDBndAzjYxlQkOteT3UABWIJfcwwH8xynde1SFp/PVnRLSEyg5RCp5dT09/57gxGapBgB
r44lYiA7TH0Ie+SnDNqvDlqQHSGe3EfuvOTJQit4Bib5Cag9rqzJERuHH0cgzx/LKqr0BTpW6SnV
Nfs22vIhDWpcVO0r1I7W6yJVQ/YzXwYOn8h/c4t49nTiEm8yF37R3Ky6x6I4RJg2rOhpkbYKXsCa
u8MstaLTjfBMj1ODALfclihJuHVrXknOFz8cwej51QifkUFgKUtO4IFLkVS9Cg1WiRKPbo28w9CA
fNIh+uWs16cGmDgbkAPGwmlEtxuBv0bdoWf5+h8ff3IwQ3coB8RBV1P8yZZwdoRzf/5qbn1aBpCd
d5/p9EImyHiJsldBZ4/qPep0hOlmq0qs8pim5VQ3esJwu6oDMJL/cbzjgzSibqc+81EMzoK4P2VI
nRoBG/bcWmP/7koRcBa1WzsjFT6v259XuO3RVUnOgvc8PS6O2Ux4JoIbN6gaus9RERAU4odZ3p+q
Lgln/G9Yy7RVkb29HG+XNOmD3/gJ9uGMzN39hmk3gVXPTpPofJU2PjQaztcrKQqflVir+aQQgRBG
gBDecgqcux0+UE1Tucoj8VBsbDI8RLmYBrq+L5AFzfnZLoF4wetDkbAmqf1/hsCEgHfxDHhQGn5u
/On/kHvhLotkwnsFGSD8TtFhAQnKcqBD/dvmPWK14AWe2IKvV9SdzTbDsuf78i7Glmt1oYL+j0A3
4Omq+LP8HCMH8q3f3xTmTvn6FD1e9WSmsKoS2+9pFjgWsftjG2yPURePSnEUDygetxHR1oiAw85j
gnVtuTWJDtrpmSflNAZi8h/ns7GbjXSeNvgakqjXJ7JGmhAa8EH0G/JjnlYDUomR5hBUERuI1Eov
4I8SFs/T1/lKqAU3oRDAU3P734f08mnyoNooCk1dDc29Y7Qncckog0DFqiU2nK3MBiv5D0wUqcel
+Gu6AznUv4Q2Ju8tvlyvfFOfAXmEyV5wvQjqeip6b1fi0ln7hs5UGN8nz8PNugViVO938PzeoNuq
QDVrMqRtLaeSe1rtuPZwaUlgm2UXvr1wU2DutspB+72fVtahYOT1RURtufSpao4HTy6jJS9STVrR
q2dNK2mRD1JZfFRv6aCGO8GeFxbF2Bb3OqvrtmYkPVF1cLK30BLx/9QbNvuR7xH8HuADlzqPU/vg
kDKfmfbM6bV4zjcgeSUjPLWeqUzeQWgeYHYeOwMqND8zuxE+9/hCilfErrH5PkvAx8plYGddVDWK
5v/zlVJFl/DbnEx1G7mYVjyTt+lBV9A1NmrqbFBdnjf5ZpzGuR3PTBhiQBK/OBc+6hppMTE2yQ49
c3G0hJLDjJ2mzuRfoidiOJ94rqEDQaRS+0H4e6oTdvUaPWCOb8uB8aBVYo6S6ZIp+6DsZ9F256EL
u0MNA1Va9yvM/WKiswQ7N0DN8WBkE9zTxgo4zy4ZFC9upzfAmf0P99D5Q6TdXepNEZf6GSspvhxY
FOWRy6djoZwXiQlFtHVlCSoRI6G+hJECGBRSneBXZuUgX9KKEOmxIilZSifU23trIpeFHyGg9WJs
gLfiT8LU8LgFwQnjGnOQRTmorjlo6J6I02qGI8I1xdSAfRPOfXWtK13gOKz3KvmcQtAptzFTVAC2
MxywSeyTIxxbrtYlKonP96dE9TxGBZv3a+orwX1C5M3jxyefFHykXXcuVgxcHbRs7zuJ9Z76xoMP
vzkhrzyp7nJ3/HwFgdoVH0u7e/LquWdTrZhY6zjsNFc6DVaALQ5QSQBLAKBUJe2Cx5wqxm8N7/y1
G8eouXRIWDYYGJUysJsUbridoAVtfO0Vqejrnrahjzk14JHXYgbZ+vmWtNw2BLe1PMBwZDzBS/Es
8jvM8j7I6fffrkqjsMq1Dsp6PRlPwc1+WsptyAn2pbD/22qPA6gT7B5R8pl5Isw6+7GoUe7SVUuK
9wMEYNki+8Rd1GPxk7YRXWNXRU04f86L18Ym6fL1K3M19wm8vCUmy+dY+55nom+SaP7iVrSQnfra
MA8mCJ4Kj2+tCCGKpgcV7qyc4RDh0HbpvBI2NofCjZogLL0ISuS1F+4MSBV69DvuTwaoXWJ/QVj+
BhBYQbmpqeQRknPJBPIGJS3KP/pF2TDKOgFaApkUwhWgD++quxJ0Kr2zuJu+u3yh99lZC9or7/eb
3mdKs/ELkMKchajXHGtw8tEdZG+Hy6mEqMU9la9OafNrjd9vI+EcDyL1BJzYV/kiBU7Vm5I2wZWT
YSEmJqOT3SounXbwZv+aq4IcDlP5EFafo1qRFjqpiA/pRiao4RCnzpBRRRguZJ89ZqnCo1J/MPHN
j4kbL/LlbwTCWKJkR9JgBnPnxMsrCv0JmQ0dCDfLuSO+NC+rj4ozHYMq5c9TbJbPE2bUj/KXiU/r
mP3XGz7kmuw/RJd6mLDDJO+Cwa95/Q5osLHUUsI3eAvnw1+YHNx+Xn70a9yxQyEPMlwm5rUA2sS8
gTwlkCQKi7xc4Vn68zyvgWM/M+Yud/3/NGSR5FP0JwEO0j4slfUyEOBt6Zw5PHIfh/n+146bQqFw
d67OXC6mLlTysbLFa1CU6PEEvSYVVsk0ztjFq5qAzwaMSLmqkmYc0bq+8WU3viWbbhhd0tBu6fpu
yYaMF6zwo3xsvEWTdv82IBd3DG6C7zaWh2iB2ZPlTE1sZxntSVngjZ6lpHyzw3KFt9beO3oR/ln1
J54hiQGwWj0ujNDWy4mc94zTc8eoaV0dNKs/WPPUB0eLXpeGH7qxmDOQ6ijFxSwEoD2KcBb8PMpB
G0UrMGWSg1Q5TdxeNhDPrvLgcNeXJxTwBSCTXb/4yDu521Ylls4ttlVWbUXB6V8cKy1+RZE+HL6w
1TDilXhups70xwLBPWCeRegj32OeSnHPDK95wLyCQkaCqHwSoIZ6RF72RO2ZGYoSn88Gd+/p6Gyo
cMI8Zay9xlhkJytYLYPPc/6LY1LLcCHdd5ZgSoESDhUaveLYJ4fbeSaj6oMZIZkKgP5ZQ9KVkoHS
7D3tXwrsBqH50jdg8sEWjq6zm2rPtn9WxRMznJP8ZD4av1DEArIvFdaioU80i1oWFfdT00PUxTci
svzUYKnqJompRAWDOZsUZKS1GvKKBjM+DTi10UzT7z2TMwbxrvGOpifCphwigIlGnfUWB1aDTCDt
ObN7iuMfRTfsn6lAMIFScboVxPqDe6I+Ht77BJ8G9DZcGYlinY0jVEQ6LV9IbuE4czyDGG3JcUJg
KVrTdVAO4fgYrVPYb6tqCCOc/nBFdeZBkhhjixlRnf5cW6q/nOz6TEXWu8dpnHinZRi69VjObk8M
b8zj6qL4/UKmBZ6OgPtQh6R55cr8kQq2cvj/CbCDQx+1Rj1R6x43i/FvjIHIYm7UxTgFZWneIv+l
1Ak/kRiRHuiF5HrY+GqMS+kwd2MXMYloCoClPsvQiYAqZNVV6bhTiEwdaQAJAfVJ4YSAtwko0aVY
e+b/+XH0PD1Ye/FpchDgonYwTEQ8RKEMNsba29Ll0yeitTLScdWFRMaVOekwITKJGyXbEobPF28O
BazLDjpDrvz6l6xQHjnfDTg8vhOOyC3+/QWgI/Cg63LJFyKISbO6BH0XMsJHC1+pBZ04l3Wr38y+
IvTAuFqTjeEh7fwpl6mFCCMF9q2IOYGjNGDmt9xiGAdp0o3My4vekhOp+7fTzfmR6NoAp1C3jJuH
GQFYL4nkTI6NkIoMEx9KkXKfzvTucMXT+P2w50WFsJyVM5D4grQu/wDU1PobpzgxNcjgEtPpXWdL
QW3xHkg84LsSTeOUEJh8/O1/WiO7y9A9Bkfw7ImKynFmnxlGorcllELmXiFvFxddwG7T7blKJ1An
QG3DFKKZCVZMLg8bQvgGkNG1NR8jL6nhRqlVsEQwunRsj8pkIOOmhnFcfpt+w7lIRbfcpnhDE2lF
CVB3GUAA2q2L9ObCz4TKdnPbCAaqHDZFZUWOK3mwOj7HqRky0q0LvhDFNEe409fe5OFUYussRcDg
uaB4pXv08xiTATLec5SasRiuzygsA9fF2k8Sru3FdCFrOaA4UYfYmSJH08K5NjjhonIi4dok4rG3
vNqSRfMBo0p/Fcx8gTJ4dPGF3faep42eToTw2yTibEn2y/I7x5X3H6o6Vmaxb4Z45L69HmI2Q0Ap
u3F676XdFtP4WhH3/WizWGy52tuVOhsM2nPIyXePDCUNpA2nBU8XpVDslVSew7xnmj4dg69l5ru0
v7k6knn4LkzIV2lr3dVlHxuQEc+tN42Dwaav2t/SwZjLUoI4YQhQ2+rWwKCC1BaHhfJ1tamNiX5J
zEXPZMExwn3XGhtFfYY6vhBWlgqzuXIPSALwWxzJZCKmEiVzXCaTVAYv1yI3wihO6tlWLDQxk3th
nVSD8ST1LimCFG/AVGNDb85YUdHnDI44KrTKVivpxfsiyVs6By3+kmEm7wOrT/oHCg6WjVFsCxb1
jc5BH3V1jfbUfOopqYG9L2G7mE7CdxwgNn0OdWE+9AuI4lQadR4jHb12j6FQu6clsXr1RwK20YQJ
U9H6zHbU3jTpr849g5Fo/aK2CYpaS/atRp8U0lrPcepnuEjhKefw4N2fPJGkEJij5FIEORJVYxJJ
Oabv73EIvsrcWnL8TlgXPWHQwJ7wYwRThaVUZvxkZjRLo5ANaY6iVrmrDCkp1Wy75ueHrK50RT1M
V6ciu22yPbnm9WmBKgu5MQsHW4ci2RF3JWye+J/AzmsbP3Qan0xJDhUZ/xp2Kf0wLOSIcaS+lRpm
J6bbLfPwtOEgdodlTiG7R9+SJhtuBM+dAMfRgkDZYbpHFrCJoea29nIBxhz+uUXn/XXDkVteSiB4
hsfhQpTVJG9dQ/GzevE0llLuD95Zy8SxdmYKy0Q2m/F+DgsROZELGG/zxzySuhvawcXgy6m32lqq
RTQPrAbPN+PfXAURNb+QF7Mai6BD+iDTaUzQ5dExRQcsQ5hw4w4C0B5wk7ipc40czyyClf0sPYrC
A57KBo/9qanoMbbV/P7ZJ72LpxqT0+iHBFqlviEG69AvGDaV5UsLIkSrWQ+CPRG8QTFiQNZAADsM
U5CrHpAQq/qDSOiMN4RmEpr+WURvHt3a/2bDcV8HbAMGDJvlyM6YymRF49lDh5Ev5hhlBYo19YRt
62duSNKyByExxrd8PjZk/U5rCjggMrq+VnBQxQ2umwcbbzVepjuB3gQtGtMI4iUTFzpgaW4X/PC9
deJX+Cx1ioRL6rjeGnqgBkbNywJRjbvUbn2pne+LMCFoiaoPStbN83eNrn+TjsKFfKObgjqy/KfW
ANMxQHe9ecjsCXDSU8jKUCbQP/MkG8hwN0j52ek+tfAM03h41IezDfqtxUPYIVEZAm1NuVYufrO3
0WLXr7IO5E69DP91ZXP5K2lHlXh4fq7ac64q5FgF3/RAhdUdaKXVJaYkWfXhrZQGvZAX2FAaQm69
kO1wZkdF5LlisL0jbN/SlJsiYEAHfqjIzLB35ECBJGecUSo+kdAo7nRd3/OGwalryptMc0nFGotH
ZJYzuZlTQ1szjdws8jYJhEeaVqUDPVCYPXRbZHsLJ6+fVy3xk4RgkI2GNfcWfQJInadt69OXCHJV
F0O51xhQjgWSuxyzCEVp5wQUUQ1dh3vVRJmPE43AMxPsXlsg5DNsjL6ptIZAlXaZuKD+D9hKICjA
xaVQfo35RpKWEyqDe1jqbB4L72Ajx1bH+OkJK/rVvQOlQenVjOyxIOxLXbVzHfBYm6KknfA6f8EN
LclWVlX9BSxRFq6QBuvW0/XOcBWols75F/J5DCwTczRF/z5yneWOEBnjGGRNwiP5cIFvAuYPNI8R
pGa5AUDLnoUWdy/Eoq7zuYbTy83qfqpsVkwoCpdIx3st8mjBkWrwpC1npFOs1n7rSVCaw7sifKeI
hmYXdntTErnDV6z1FtJYb6hf8zSft/0au0Df5x+Yqdi8q+r5Zl1hVT9iF2daWUT2mJwGD0KGGdmn
uMdl9G92XpCw0C8TGSLwrJ4psgTR/mG8VeLfrnkH8YdSpK1150DMes1sZb82A7LhSG3sORj4kZou
GWsIr9xqD70wVhTk0UHOui6QI1uHXpnGkGglxqf44kCU0HswpNpgAC0SO7tW8CWJ/rD4sBXuyzuv
2p2Q/4BYKqwPajR37cfpFFi7v8vfcHHoDFjub/WvFb8GuicgZ8qyV4EZ2vpL2ChpUGsWVcajMVq+
TwwnKNePTPVmLT5K2UEtMRH6VaBPDSTIko7fIp4K+XWLHMheRcOg/U/x+5KYDKiknAXBmJhWg7+q
S196qaAzT6c/RowTueQOISgNibPhaUO9BYrCNz1MG27Pe+Zj+Ms6nT74Ud6XNtle1pP9LgmQFEz7
vGqrZvaN5nZEyZczEkfu0G1+/SKwQW9u19q90730LaXkHBXZoyy6+A1FOTU7tZM1zwUoPyN2WREU
9y4cPbBHlOkTx3dTCtxFqI4aMnoXBpMPBIOW2kvyp7jEF7HtCysy4yeYtUDiy7z8vAFEXCOqIMnd
CSgxSCEd40OnTPMrAEgiJvvT/s3xrtAtMRTRcyHUS+NH0FkddKLyqRXZCr+liPj1rkUGTSgOg2yx
6lr7gwmBRAXzPhcbvR9M2OR3Y4amU9Cmlit/ov6b/X2HNnfL0/rFwbfO23K+GbGJ4GOJS0SYZoaQ
pH+oQb4SVaE2hnGJUS0f2fmRgZaAKMs8s+YbRTIti3cpzxUI/gxt3Jvs2AbZCS9fe0ZCopqnIMAR
jDAFOEV2aI+/bwdNqdltoy3foPa5HlylEI4I1yDirj72u/teqsaQ4fWldC8+9uroC2TG7oinG7xO
6bfs/g+PVhoUALxGP+GSdQwCpfczEfM9VISStVJX2SW92qXAZBwv+LYHbn1lAp51BLlOqv5jq4C9
O7Ihuh54fPSBwvVL0I+F8cMlcwIXvX6xIPu2q2WvaWIY3vOGcJ8+T1VlQolZrvEWfsw9kYTA9KKI
0gXZFtcBZiVEqQ+t0VINCtEXx/VADJnVaW3MJdbCcaEU86sxW71NhbS1+PUvQ9FgIECBdvkRUCmE
sun4eage72jQfU+y33EMGArLKVD8evZWLBZ2wJmNktNBxiT8VjdlJJs1vwpE0ccSGtDw2vPh5kSb
sqwoN3lmxKGpYkpfZW9RCAkLiXecGYmx8HIkjmZuBWjAVOirZTkvlYOe/N2ItG09E3+C81eo6KCY
NMs46FRv2Zaeivs3onzKj6ZfZJo4WgJ+rzj5V3ygwT1zbvp5qPo7ezfEuxMxfsSg8/UeiEb5YxzX
x2SScuKkk7GpzQ3WjvHgisXWFd8Fi1wkO3lwNl+wHsSS+UD1yFuwdLuX4EEid9YHQB8ZVwk84GRv
c+9S6sCQ6wHjHYci73aq+rFkXxLx2lFYw6lCyzPbAeaFaASoKMQtU7EvCsWP3PXm3xc619cOAzGA
qEq4rlJCEWlWgyay3BhK0te0F7o6ST9u80Y4MwyvWuRtlVCMbESuf5JxH8t8Cz+ZuDgXRQ6vV9T6
+NIMXcdfqT3tLnkfRjZsI3o/um+DtRW3jzmCrYajIf7a78ppMB6rFIvyq8pbiDGqB8GSDcuyUF82
6t0H4mZ27kNzbhOetZMzFPnhjOPFUvD8GeKw4R2H7tbnd1dZsEV5dlthUyhNQz7L5EL2YTaVdVac
sB3Lh1Bh78spIcUScN+2OdPEQnFxtjamegrTVANkF9gMS/2Lo9EIgeKHY2u9aNzdC0/O/QxBErY9
uubD2pCs1ZU0OsMj4WWllyPZXNp+zOvQc5jn7tHQQMc83Nm1PlRliorClYWamq2y65+70Mlp/LwV
0aWBHiplCF3jxZ9fO0Akpz5qCpjMrAf84fAlwPQS6+JnbeSqkMpuegxVzYJFCLB+WsRQXe4dV/9d
T/xfHA97OsrVnAr1ODzM9lOPr9a5mK/czsYk9uvgFOATuZBp9VY4wkbjUx99LKHhJmFlFOthmteK
SGFNhyOIc0HRNkwMRxivX3MoaXXyKvtGuDK+u13qp7Qjqnd3hAAunK91im7i6N4jSzVlmKJ42939
ZR2Yali6qdFOGTS8iVtL0AZCuM4qHNb3NQHNtF9IvlWpcjl90h66z7fATFnyHY/qsWagqjRyh3LT
ElC5Om+yiJK5QeQdyHNiTAUN/hMbUcjzZC8+n9882cgha9sGMnz93A+GkJXzV8eChr1vb3tbLEcK
0QJzHR3InfhM2bNpQl2SccqDLMv3TGH6+v9pN3AeY7pGzuqi2PaitBjECLSTQ7mTh/95yDvwXEgl
GWF6iPUaPXR4YIVQTvBpLdYoRhbGB1zEWEDhtKQfqGqxlGTVIH8RGFrgmjyD0lmTRu9qccLKidtq
a24UqsCfhl8JJSVJwDZ6kBHCOyMBgVH7OoOsAa4VN6uHuD0O0MvwV5TbWqBGFR1biNDHBxhPVMUH
G5wKv9ed1bHCWirEa9whZ/bJfaO7T+W0K+fpx9TdUsmU9K0oLJFiPI/UlGMRVkcmjB4rlo9iL56j
q1/T2elkINuujkQ8cwDsPOU/w2pUDsNLwGNb+K/U36eP2ZB1K/wBtLm1lU9jew9VnnhP/YXYvebA
kETDlByoeF09kMOLEsk09DHXxKHQ0Ne6TR8V62cXIWrl1UlVMOH9mJg8/XUqc/kcOmncfxs4Di4S
O8IFHlCMexFwXpxy/A+/N8HatYXygMMYgjYShJ+BziSruqxkJEuvkIlRLAcD4cdQvcwT79Vz9x4x
daCpPzRwcwK7mClpF7j33FzFTq9d8cfEsIO7VF/C3cUp33ja1xVhBb56hY+mQJZbr31DWoiLA29d
JUvPNPlDHENgmYE2P3cUKoFLS8mdnjQjDIQv9gwddBd6NY7jh7TBktmVmh8m7dFp8RniL9e+gIuG
QEY8dVXxZOrS+dzwUcyW3jQx/8ScnTTtOAt+tuKGRqhTfe4olxEGdpEn5v7aEwsXSl/zrJGpHBkN
I/aJwJ5d0WBsLm+8Rcnmpb+5UUorPtoAGLaCUH5MAdE6YBkFDaVVRa0a+BlyQCdl2AXKkjOcbDg4
jSimbRLX17/yHBvxyW3rl/VtnCGIPKmkXafbDfQq1riADxOnloVa4QvyCHPFHSsJ78Ta4/LUMOWC
u5L9k+n8sVEmaXdIpAUZ4tEFDx8mWE3OfQvWoOgSpQFcdCZ6RQuY1dJMkOExy78dbwJYEcWMrBzB
c1eTMJy0LfY68Qt9fiJIVk3xk5c+ZwKdDYKkfGEvAOyXztbwn+4BAN91zQFbAmZtl8Y7AURNchmX
odN5Bd3nxt/wCjie/CQAY9H6/8kIgBaGTAHrsY8HsqWOq87PH5CusjiZGTJz1aSizbigLDTR50N9
ZVi9uMBGmjxyNXIg5kB2ylCyBPEVFQ6s0Hg2FjtHU43BxbgOCUlNZ89lWOB44PPJome7eGTNWfY5
zjg/UOLRU7cI8cM0w1q5V5NgLwuTKzq5FqI0aJ4PQQknRGmEmA6hQUe+J4RK1sIDqgDnWW/HNuaK
xceIBjSlEuPuI7pDeJxopCFti8jFkIrXxKhld59x5+dJD5lj8jRyJZ3OjLVq/GF0tFWlfdui78lV
BgRFfzqUYVGnydjRSdbi3861SqD7ZmOyx3WHzCGPz9n0MOjhBzav/I5bBrmv/bdFLYEinqsUCSos
8chCEkTvj0YXCVM2fI6Q5GKPIHdUAiapNs6zo6sdna4OtkHOLFnlYOhjL2hMCSEi0i9a9zul7eO/
LrI9yOfEcey8MhMUBitrpm5pYP9X515iArpbtMhrc5s01DgCwu3ZMVoWoJC/xJSgLhwTSIiM6YAI
xTQDoVreZkK/xspOrtvF94Nm2/xWXaOqaSMVTGTTmZSknhbMvBv1O4l54KaIyg+3jXP0d9RhPilC
Og05UWWeRFGw8l6oUP6Y40SSiHReUsfMW+QCal7KF9yaEn3QYudOG8sDkw5VJfLWHs/cuvH1h2NR
1T/73yUS0kz/crFrKuN8ADXIwQiantIoEGSU94kgkCi+UG8cb0zzzW+ganstWbxuiEqt2utcYycf
4kqGRO0iWfrONBYOHYk/f1rzVYUQD5iRxdr2urnMb8niF8UtbaJMghtxn2WvSsvZdQ/4aafO+jED
QHXI8EkoneVMHYSWEU5g4iyDxo4Gma/DeQRNfamAn9EFz8JiV2RnR++kESa3ScC31Kh5q1laWfq2
p38OMU0w5DoO81CNADXrmLloWEpDkL1B0BGmttjY6MDEwZF+jHqi7LkPv3n1hKhDnQyU86/ULuwb
fgCu+Q7eRFACx01XJsQ4pEwpruHyZJwSmqYqs/gTlWp7BVYFyQqbKhij5SpmDfhxNIzOoLAVZXh3
5omqv1ChTo8eWvKo5+5WyxNCxrIAMBbzmNgeljKVbdMaQ8MDjmJw+AZfSj+mcG40ryknDQbjTh05
z9xK187zaq770fjmJTA+YwzE2Bw15hW7Jr/YlyEfKffKZSfOlRio3uqC/+Ps7O+6KCVSsY9HHJ2L
oH3vkDaNP0t+M9XgL99RLM+YtQ1ws5iB1C17OsTE5bnPrFf08DxTKyFxzrtK5FB76Cyws6XL2ClP
Jglray9HVnhPhuNY6iB9ik78zESKMD0o+uSfuR4jNEnuPKhXc+qg/NmxXZTA8uebt56XiIOv7mGS
/fPIn/RWeuka5TicxEej8m/MD1JRZdeuCPbJXl3jbGI/5BIG5itplmC1QFkzWdohBDsH3RMubRhe
VZ1rDBQrvNIJ/1PPt/sN914s5+m8/74Dh76wu6i0Ia4tUYhQbjuVEIrDBexPCPnkfl8CGpgBarGT
6sHJDmdzcIatEEZHYQvz+NPTlxTJptAid9srzytOR5Q2JD+GSuGN75Pa4ImWBrW7sgsYg75I2FjF
k7/iacuchkXzvTk8G/fZxSPWicldLSXBndMh2mxv6tBZ2N5TI5G5xxg3NYv4NsvrmiK8xYxafm9i
telv8J8yOhbqcQOSrEzc1Akoc53Eb9OpArV+rOTVHlTsX+CZErIw0qshYlLKNl+aafUVDuGuR+iX
hj1iBuPk4tyVMoXLDARoSd3UhaX40PaZSpOJrh7v2cqHg3BalAiXlQRwcBb1DDcBsP/ipZbef5jg
c2NhoIfkeOcgPj0fGve8pOs+e+O8JfVRvukHjALycOZLA/1M5MvSx7W32lag7rPukJcM0znzZN9Q
nA+1m1owsiSBLktWtretKNYt6iV+SakAr+5zcwHhhvyK7iXPwRlADuq6rgR0lyZ9sQjL1g4rhYWw
ptQr1F0GY/5l76p0UVgRC2rxQx+vxa/x+byvYBXQRX5Ty3VvkQR+xUjFHXZCNZHlJoSbbmJWr8PZ
VpUKtQToGgGJBQ1EiWUVUD0+3ko35PJm3IUC99sG/E8aZXWh64FEepGWy2h8aZLQEGLvrYcyUJUu
E4Sg9uzCCbm/P+uqU2x72wwK6LeMdvpp9zkPaIYQV3tO6z8cIdsFNZgLGzIOV+eIytAmXj+vDtHk
qTH+E1xFKzhf2YupdHyL1CC9plcAJnyaWkTLF5eMEt49lWJBT8mrF/F+ZvUSSou5I72NMoGCh8aE
jEKWGVERFne6ceWvQywPPsC7km0kwmWfvnPNF3qTXPwKIj19BTtDBvynm3OMddt1Wwf2VcM7EVWt
eXNxAmF+Sj47D1O6J7lYfK+sRawXh11WK36QWje5OM1XHZVbMIcTFSpdfFyzuo9bE1g7IvrYMyKI
LkW4fVeB9Uh8kGUTfdSRs29Gi7VFuCZ3n3yPSxqVvLeqKZHirG74c0/X9tc5ZOSHFM1fuqUvHNbP
uQtvd1vYMMUKr4R6HTA1pdv/0pbU0mtWhEyCDJxIQ7Zy44+FJ/6CjuppWul8Gq6rT6TX7lEkWDf/
XFx3U/F3ZsTWr+GXfB1Gg3votSovlENCWUKRlBdM7uWI7q37J2GmNWUGYVP+n/zy0/9zXvP8FGwM
lnRP3HFC9aUPHodaNK4pZlWIeKTNRwHtP27pcMy87lURQ+EvtiybDjEsvKJ8OmMHavs9rK56dy4v
ivBRR+F6EvPY6GDV9m5xfjglZRryS3GsclGrk/Zb1TtJptQs06uKeB0iGId5CzJTx5CNi1SFXWu9
BFTMlVdZPCM8tYreqEXvySwlwcxeM3RA9nalz9BJA7qAIjlZMHZIhlP+vQmm/fPaKPe9wX51dmQh
dOI4WURAr52HpezpvkNYy+c0+nJDpkaN5lF1M46NnLF5909ug9tGuJr0K7JjFVVuLNlb/JfPGkIn
ge4ZHAfRP0fq5/puDhbo0Y026O+RIQUpX5eOmbgZ680kA9s2Y1M+NWKjfYQhurzUInWrYqtKvOn0
JJtr4tiPal5220PEAFqH/9/0cGxrCTvxAr6ry38xeDfWZJdrrENju14WecT5JXJ3rbx1LEhBBaL2
k6rSlqsFzbuQy6br5a6ban47M5I8rOmNs47i2b/MXV/zOHpnrs6QimEhACqZZ9sQy8dVKxETn2Qj
y8//0Q07TbmQElmJknCO9qhpwdCW+iL3ACFqEyjzsR8W2RO0QjbhZHe4eo1DizLBAxVP6+qqb2TY
p9Fk/Ba++OIGo4AkyVFfKFInnFFq3MSgcKaGxLkyEgSKbXj8LmToLdTapQoxWhR+X/eWid38OS3o
jsVvLekKTvVKl5VDQrBhDrao6jL+dqm7iLoPE1/yOqDVX5QgMuskZZ+2YaE+/ItPXxzcdYygRRuA
cH7QPvAl9+XoR7jo9n1u4MwwqFwInHwVV65qKtP3+C5wzeZJIE1Km8E8MsMgj9PM3jd02mrFCLy3
gCtWB3YY5GHATTQGK3IqWaU4SIm8HKSlUveAMyMZ/fOZNZZPUNRyw8w/rZa263A/+Tb38KMYEIOf
IpyREp/i+85XxP6p8AQuTtZaPZJaU8v9KBLFZ/oOSdOdcqE0sYDYLVSDYv+hXOkMHFyAPvzNaruj
qlERcQeaew1iO2iwxM06dD+HRH5RkJfYH2JB0ldl67uLSwuVBZLLWGB44xHqcMzo26UgZfn6ee5k
V+gm5qIVHuqdfOwgzHv7d3C/OcoGi6U89h7YTb2YPYs2TgEniEpRTKmiOMYK+2s4nYiZNgbKhHbS
y0RFpJm3gDYMibFYz2LL9sqHJzdVrDrhDcmMlkBwXUnBjA6+wJRMX+k0FJ+HveLYCqwOXAxGwTzd
RHyjUzpQCRWa3MsSk9eNgIX/YZ8hrGWt//Jn5O6Csb0r6WwMPRllr0olnwTDOvYYDb0NsjGufYUj
U/XnTHyRssMY0MaaDE3bq/6MDyZZ4pBTtFuE6Yq5JODQqka4rAoZGswBberDGmgIrxxdbCEB9N+B
BLGWoAZg0ZlkCI0DOaaZnGa2laJ1jw8mYx+h2764dITQKuJ2dYi52Yh0PZ6qmVxxB0xVt5HBBLLL
AEa1wJs+vPFRIScjuzeBgAzlaYH4XejeA1Zl3NFMUUfwo8z0yyvHxqUCo8ilY+BRpGrJ8fPa7q8F
FYHwSAcDqkJ+kbBqh283aLQK2ii1hOMsS9ecWHtlyKhjMdWO9yWoQHtvPUfZPXwCo23yGHK8+UAX
f0WEnfAIGXSPfe19l1wbX6wxi24phdntAIz/8RVhpuTzbzHlOUcCD6+NGNvJ/EapiNY8npR77p/0
rq39jqNXUNe7mEND31XHtPi0vkUkXbIiMyClq5Krp5RY+wyfudTO9LOOT80e/Cr2GvUvjf7BiSjO
l26/qi/Ll8C9FzMANYnJ6dlrOP/TjhZuoeOHNRc9UGs9N09TN2plbvqGFOM8x44KYpwR61bTz0ni
g87bneMC3RhuFvwc80KPouQV8QYHUXbyA7cby8sFKsK6K/8CTpSfHu+SA9OT4cxfucbKcWzay3Mu
J4Ko9DrpOtQnKVsraWbMvGPF8y8zFEZP7aGV0c8354+CM/qpV90tgC/PfuYZvxt1S6eo+YNInWrA
Uv6+78u2PoLMDB6zKvVly9LaO2HVcMPdsKjxY03yy3/cUCpjBxl9e5lA1HMinQrocd3Uh4cxDlPA
iNiMzHG/E/4Jz3ZP5TkbRBnppdgeiRPB/bxEAyoCd7vuIlR9E7vBOvpXhnASisuyaahpvrdcf0qx
OKAZgUisD8YuzUK+f/XeWLaRhiHYcVmFGNlZv6wRAE7JvXKSbMAyk7I8mcn5zC5HfFfvNEzerZyI
i1azzL27D6spIGRkwfN/UpNyKtz0SYltdSIo63tGkmYEvN7YytEUqETEsmUruvAGj4ZcZ9xUy5Di
MbHd7NPYyZDkHIFzlD+0n2Js60K6xUIB/fXsxzoJnKsx5qfk4sBRetJz8NlO/mPLx6PBGiCb/2Ek
xZdHkqQb0ah7yvCpZ7sqBa5r6Hv2rbvnK3vwVpuGiPk0kzR7L/snjxsHtg8fP+AucNlGoWWmva/6
rM6JFd4BYiRmxTf1JwVRJJFPHqI2XBunvYGFf30vw+lgzENAEnLo4OcpQgjcsNBramhIaLacXnAj
lfx7VpCpxVEW04RgEBlloOFA8pROrJHcg9Tzv46EypjkIO0Rsm2OxCVOSFqaSoUP4WmMOKMN/Zx5
DM0yxQDwwPQjLzVpRocJqgwFL9u4cP7o1Ztw1M2pxzrvyV5egg4khrGTZRzhFiMIZMAqezxt3BAv
zopLVslSf2HlCiC6J4IEa8TEK8xYkKo57BJie21X+SKWKG600vFTmt6d2eNJruzLAezYvYbI7L30
/PfTca557XT/aEIUAVRVH/xjGQaR090Gi2Q36opmaG+UQX5dmCDxLquUOu1WexgVVqb4xTtLuO8k
dZ2cgrTkBSPg3pp8s/CJvJoIm3ZcLC2Y4bPvcl+WtdJc2eF27QAZPf5GvW6nreI+Yo9dYT8z2pYm
hvTmSe+4N8oT/lIeeEdK2nNyGAuN+r5J/AHeyQTZhcJTsOaymkIe0tvhdwBeMjEVkpF6UTaX4ovy
sWRJpGilNKwGvRdjULOb4XMGYyNAMKRLGYUhQr2a2wVPKv9T/6Y+JhNzrF20Q9GLNR3sy4g10Ptg
ydnb1T+RiQDgqStX32wCX02j9C+68qzvZLYze/jKMzrSf4mCYQtuAteePOdNVQubtYrP2VyezNX0
VioLL/aqRemdrwfTpOFEY81JXas7ZaRpaVzmzCjnf3ye0Tsonchnn9V9jKVUWS41lFgim8bbYfUH
pK9+kr0OLXb6Xg1xf0/TL02/ccO4MVyfTpzpPbmHyqUSjTkWg+P0IAX45W1kOIzrVW+No2KMj4Jj
FDu4wMsOoBqde4PWKHRBOqUFpniOiwolSUQDitFi1S2mkqGF5O1z42pzKLOX2S2jOt2lHOetIZji
o8wCHttGxaDe37llLCTQDT3iB5n0nQzUpuRf0kJQUBcMyOU/3igllU6D8rEuXDmXhaZgTg8YLUPD
KPM2zy60TjyRkrjpD2HNq/2SMcwO5LwI1tqNHZ2giti1mgRqA3WjtTsG5kl8I8fVP8gbFktu0QJO
dMxwLc31j30laQJ+vq3MUYGCb/zyr3U5sv9mFb61OJhobUdUNe2ASJJXfpVpwqMjY8oimj85+NWn
O5bPgK7OiO24jeN3CHcj9hnYCM4vidA59Sm3ElyKKXR+FHKZfRmKFirfM0+NAUy5lTHfIcht5GVL
eAEvHszklTCZqCB59iiOhRnTRVdvKK/iOnozcX9N8xnLeh2MD3PglEte0UTH86YkaSfNXeliBsuA
0CM4TsjymJRtNamS9KKtB394noC7I6lsCjEGQhnG2DUjkFhtJU53JFj+e8LgVE7mfhNjXayt/NCr
jBTu7GLepqHj+QxXBlrRaDQ6gfn+UfB2ujOYrR1IoNN7hniwWzjEX7DZEBswvrCKU9IqcIrmlvUo
YeZQd8XT3g3jaWNJhEVT5KJiRhPLSM9Orc3ZWJpA1iQnyJvUFQPR0XxqSZ0oTSPJNH1gxpK0DhB+
qDcnoGq/BGLN+awm61xdqqxIrYHg8iyJ/pL5TL0nRQkzrBhAyaDbXRwFZCZ6FRWsL5Tlr5iBeHnS
WsIL6X3j1LTdkpRjfl6t3UpKacA30oqkOs+9+2M/R8iCe6LDcAuz7Nks7UdIWeitfypTCRo25NTN
BdcjEgFuAoWozbRCfdVAOVPXMldK+DOMkpbPquU1LaUlU25VHMV4zh6KbCY0Wq2Qy/K45gvmXZeF
r2XUWyeWohxJrXogWMeBJCApbS8l7Xt4DmZj8WIybZDZRUXLaehcQjAySAIu5iGxCNlr2yjHwJiZ
eOyhhxmiK8n0w5X4iccpPOAnDfnWryIi1uubOZKUzllR/UtPykuHMVlq4YLu07tj7JQ3nEua4nry
IDdrHeWgYo790Q8sKQ7kXBamBrd4k5Dy4sYQgVlk725ufiYQMpmbOlDnH7souz4gUxmfA84TtG3f
1TiHalPrHBUUDTBNZBOF49WKBZpSZrscVrrROTqfZGcaICACI2mkEcV9R+RN8TRkbz/iW/0aVJwg
072FP+rxZ/GOhNSj5/4ZQO/klV0ug76FIaQdDm7a73u8zYP9TdThcyfGxq0Qz6ln448HTRW7Gmwf
pSzwvM7RbkrHjf8sEJf4NkPcTdUJyb5iM37FE9H+W5apLXgVPyE+F6MTyXVwwzIDOSL6/0RX3tCS
9e3oZEzWO0YDT+n0amHoUf/7aS1Uoyo8xIgxdOL+w2yRztCfyG1aDrC+0xP8ACGcPubpbUtdxg57
EFRYAxQXVzYTzc7Avx4UTsFpE408AqAaINl0yoOYyrbqaiGy0zDo9TaYpSTJUDfzcU667QWp3COF
ICH9oaeCqz5qIFJYLNHuYPIE2dtWGMjw+YF+J7MTfARufW2AOTQp8YyfyOQchNCxg7El+4zdpLOX
XUOQmNKQAQe6qYzS9uSuD2cdVOJtdB+Hr4Kn6OigXjPHU6JjQSjmB56ivZuqlyKtKKOJArd4p6IA
DTIUwoZCQ+y614saumR7MPlwHi16AJ//I6/GcrY9DfgpMg2bx4P4HKZUkzKXDSTe8zmsMDHEHTiG
iKsTDYe63E9/cUXfDuAiH7ahJ+aHE5xFZLEbTqyyPufHF4ZUa8eiAc+JRhMmXUAyxWa94hXIWJsj
NZ75EGMORAMAESK1bcAn4oIqdlWQ0hYeZ1g17dNhAKIAyFrY5CG446OAhaLLGlVFGZz26uNRaHA3
hBGe30kjIR63IZ7iwoT4baRM4aLYSsA9sbITllK/TxBPvIJooprWV22Y3v7sUTHbmi0C/0wXfcB1
B0FH//a7GJXGb9r/BqoSnJYR1Wm+KJSdoh9zDztmYlKGwTaYWiVUjxcW+zaY1C1UCKvQQfj6vyR9
h05SGBMrjdWAx0FJWyVGh4tOTtfdUNAw9JQgAkKrKiQYiT0pABAUdAJL7xbm66Q8MHgQdfJYVTjG
WR9JVSigR+ui2u5/HQOM9RKy2MAj9YpTyh2PHMy3kb/HkeE7LqtnR+LST15vpYSOKf3a6KfsFyqg
2tGo8nBzE9icURH7I0fI8hulLdH5YYx+KtTbVZ1SMk76tVyWLUe14M0EEQElqQRfHHIWwlEfGszn
WA8QtcUFAkL3U8E6vUT3EKJ6vZvIMk9cpSJqnxVaLJ/TCG05bPC7NyiCie4Kul5jbo7VKRLp6AKk
RL+UQoIKsbGT0UQZ9caTm+m8I9KOc+O78vSWvltk9aXF0OrEopH9CbXdAGgMVFzxu2MYLEv5q1HZ
uMIp+tu4QA/yTHGO80tLVoup/Z++JWw66MqIHF+e74W78IjQXUNQa1VrGcvMlhQCwUcyvSl+0eY0
N4fkVCibroM3CTjDPDnjIBfPQGL2HglddlsD9GRghxaha9r8CpOoxccJCn4aPuINHMqlc0tWTfsR
kE8AJrfgXdYy0TasTIYqWBLzEGQVgdLuH9e+xp1ucY0GB2I4vy2MUQCtVKVW8NjbE7ZUuteEWMLz
ROUWbUHbaD2Tr/UGy0quCY8RVJF66Y69d5CDFmHyK3CCN7MYrS3oU+Q8/8Jvp+BgMMm9md0vu0IL
bZyIcVMaYN1Ob1Gbsrn+hkHcLCJi3guksbU2XV5A4/qR/Mf4Veqi2QLjZ56MESsKK1pUK+liFOiZ
B+xCK+bFnre6OZg2dnOcJ+xU8ssmIDX68yTVkOC5JVz2oJx7qWnJ6spVvDj24Pj/t08oeyPi8/D+
QPAjMUk7lUvpt1udSl6wRi/1m1mCAI2tINH03tuNhsHGByZl0e19KN+NGg9cXu17SWhb7Ct5EWNS
v3QX5uX2yzO9er+SHNtCXpQKNm+pFSGXeqWHjuaEJWQhSyKq0IMfXw8YqEJVZRSjnRyXMqvOv4eg
/qobPMsXQkHF2VgAwE42hk/xDmEAR032zNOojwO1DEXl8r1vJ9qtn+vgNzLPNfXPyhHmDz9qmQ6Z
FfoVFdXhR1Smb+2bGNAafH0WpbihjwseC1CT0U6UOI1FWuCmWbuyWIon6GPDcTR88zFmY5WJFrgV
89jkXZRk6IKX4mvmtPwdBmQOUpMzSwm9WuhWh582s/mRWZ/Gi1pS88Vc7AskEvAHv8lXMi59dDRy
ai74ludZh2+1QbAQeDZ5U6E0ZSXOCS8FJ4vtRgs0/tlyV6BmmHNEBrsmatsMliuUj/FJkfOiiyvE
aJfLU36gKRCGuSbq1lysdCAO8bOWZqtsluNyK/eW15lE28RAaoCdAnlkydwPT7Syj2vOrb8c9R+w
o8aVlplvMin1fI2kO+5sPtOmlhd5MZIJTfsddHlB1TA4YznDe9rHxWpav7WI9bJ2n7AK/yYZdiKP
kZY3KvFG6R2FaN3iZm2QR7oCj/rP60xAFx//tKy5w6INwfdAFC6dx8OAyxw0qRE3z/2Shv2Dw/IF
IUgzG0qjMB0oDSQBL7Kv6mc0W/LXnkCbqCKtCUX7pX7HYZp1a7qlITDSmnq6bPzuB/QoFvWHPLTs
J8XiPBi6M49dcbWQ9+Dmi3QW3l0Smg5gc23L7tUv+1jULIZ0a6ht4vU+X6w9mZmgDAXrCRuF7t9w
2sia2N007uQKdY0MK9VzzPVJO/VCeWtsQkOaAFgMkfwgagOJ/10FFp30neq+NaZz3fHXk/JnVKcB
8tCLWieZ28VUVjWjZlSnMgu+gV/3wN9dYtfuZZ1/d1HAcMsLfPiQx1APBIP8ebxSG8j0s65uMRVH
TIN4HMJKBLkJq3NRmYFyjMd99883295nAdnc9EBigtJn0fdesygh0IHvTeRlulzgP+UUOoQbtNzJ
ulvGOCMDe3bZrrQ3aGEDQj2cZDGwh0pdPM1xVb2RwRVxoiaMj/kksau3z8Oa0HEQUAZtX+mkE2Ri
8IwtUUA0Cne9OHMrydK27xHRX8kDQJrUt28Q0Jm+3idJopoGbwiApm8ppdRvaMJKkq+AHLZydeH5
Wc1GOpeTh1YCMBLwVBWhzFzv5I2KhIX1CCatMjYpmm3UiA+kvX/7TdiwDqIdBYia3XaggTGgF04x
R1CthFViPGERxBhuoe2zv57VEQJAeh21gHn3AqUOQ/ylqOYRFhLLPgtKgPcPJhvGoMlUGVviKRfP
6FWAH2PwDEH02wak4eFJzknnxdePLzY/uh7JfHvyABIowpFoBTPVgm4uD96GufsDcKKgtGCtfhBT
Zh7XulxzyyZictKW86PTxmWgy4+ltQJ3nx3tjn7J5VqR3EXIOb1dFeAAm5VaJgQK3W12RQ9XLuch
kna4dW9yHEDD5T3B8HJ294Q0qVrRJYuv+W1TvTIYyPujYo62I/vW6Y/vi+ZWtSRYcUDjtNtvsw5T
QZbCLqbNP4/lWH4wnq31ApsjmnDZHuHVgapxSuzARDusLaPXEPTF3qrchoud68s47R0dvAyoZAwq
XqurVIvN/KAeNtaPZQLU2oa52HtVRL9/Ckw1oMS5E7Zz3QWy/z3ExrK+kwvi864wquNB7n3y4GA9
m8dbu1AkIrUcvOx3/p2bd3zubOq62D+XsZbX0I8KkN1xDAiAJmqRs2ICC5pieIgYZ2RIamcWxyRT
tqCQnDvqxYkPTBfZMzCDhigUbLGHF9xocLZdZ9jbkM6LZ2yUFjzVn4WoiGlL8DL8xqe1qtlj8bc6
WP1MYGx+qDvKukm0qx+amHKu1Xu9B33jtDqg4E7gMQPcQwd0YrsGecwANgAC4GJ9sghfMbUd1dxf
V2ZvDAm9FJM1HkhgvFuHToYEU92sPyPRtOrnSjidBPug8ZIB0v8R8LP6mJyszDkZgQRQquxLym4d
yimP2G2zvlfqVDPiCszeQ3jG9Xj7y7oDSfL6x5AWb3zcNIz+45smlvxxvXmW1ln1omx+N7/uv7sF
glwpqzkRKxgc17azB87x4ucI3qbXEVN1mxcJ2+jX2f88JeKLZ6bH7pK+Fk1FNT9Y2o+TfEPajmca
N3RJFVf/bI2OrXJrnEO6Zp2OkPLz2WYCufwOFEbiJ7SzUu3UiJ4cmvruP9OmHvuSTama0+McH01I
DXjENRFpTpduLd6eGqizqfoWIOmLP7oeLcg8VKyYDl7QF+ncHq25nGluNIui/jbbuBmidz/BTaxM
VDkzFMGWnn2ymBvVQRTi+92weJsjErQ6VMCR+/sN1pkcp4fhuFDFEHBzemjy/XdwZJ4QSEyOV+WE
7sdC7BRE4PBDM9Zu9VQrbZ1wHnTKlYdS+7I2RrB5CYXApKHsMhK9cNyNkb8UNhUGbo0oAexOt3xw
FnmF4KJzcS4vXbvY+X2iofDSc1CXtacm3pCk0ZryQ9FMlqeBG7SYctqcxWQCMJgElkCmvBt9Fd3V
Nrowhcq0a/GMDYhthBeqAt/pY24Qr8oBCMl1zBbSusOMhHig1uVK8z5wukyNFbnKz8uNv0ZnQf5X
8mxYQJDhYfpEaQoDac8r59L9ohNpI+IQXfTtuNdwAdv4jE4n34IgvebK7GaA2FLU+7hDv3Xd3ZWw
/CAxcQSQNnh20Wrob4tBJ+RxeUY9JEZdSP/jmSUH5VwBWFHwcy47rOQfLqZo7q+u2O1j2FgaXakM
YuZHKscPMTRUFEVzMAawES3asmLHLSSfptOz/mV/HQfv9yKECG+JEc2emacdkXKja5+tjUhmhAZl
pKUMIO/R7YOMzsQ6U9nTU7Sh/+USdWAgOm54yGT+mAbhPPUDB+JppH8UojSHtLNw9YKjY63ZM4wr
8ij1PiJCmAX5/fc2caJySKaozhEtU5TDuubRt/7yS5yBumSQGwNjLBuFPhuFZQTtROukGew1uzVE
bUAk8WPKOM0ydHlTJssebncxTw7LLyxb9COIeg9UnaYkvD5XyW2SBsiD2P2jblryuqL6VKaIRk+R
vvdM4xRLDOQLMmQ9arU2H2iKJa72vHdcMfTHfDXdlvPVyzWcBn1DbXvDmEbGtH3IeuGj8FMb7y4b
ThYA/WjDrGeT/l3AN0CKpFBJD5UPZf2K3DZj5lXBV90KXFbmr8YpjE+OGP1gvdluh6AtvQXBSfyr
p0/Fyb5+kd+sKh8lfkrqa0ICoJRaIJ2G+jR02ZfnfOWd7JTO0Csl82C98FgFQTOADTTcS9wSY+4V
TxCrVM9JX1ppknrSLP6+fOSk9jEANCKlEVm0Bs/7PCTDN7+RKMnW65ko7q1oMouMlhY10WC2lQYo
UdgXiuq5u5oRh3mTaqzBIx4syv21PAAKRju2IEJE4QZovUHSw/eNfvRE/dQAr8tOrsyql2d/R8mc
DIuGlj0FhE1Y+wuoz6M9FnjoKz4jXIQaLYDhxxKSkdzXQiin8hdwJadOCixkHioba8vx+rr2CzdT
oAD+1TZjHpfCjaXNB66nBz1sUiA6tiNfpYsPv/1THFHsq1FJ9DUX7nylTLaoqWKFVlzc7a305XZ2
05dJT2tPINRggnqKHmaBHiNnc/3RHtp1gjep8GK9S8u4CMOhqIOnYDYEe375qOOjVJ7RO7T5j1j+
PuDLpV29jcvNq1UclJf+pYe1dnxpC7amUAoZXyXPE1YjzCJ+wiMjZT0U7ZaOhGkyw6WVTPaHMLUZ
1FCKWnRbuHq0dKGwrOPEhB77WQbhpjWN/Tp+IuUgaJdNsOX+bD0DEi9SIsGMXg499xRU/LBCTj2F
oa2IISQwepIto7DGNvrzIj9rwfTugr67BlXNJ8LzOvbdicnr5/ndvbrJmBVxHFHohvQB23y1LySO
HiPpkOKWVGQ0ZH4rmO2iQ5OgDWhAnYupLu3zI7Fkk7vwVUkncPuD6HKOU2j8yoGAYio6zUfO1uVK
Tkcl2Dnofyl5QjIggALLdI6MmHEkr87D+E6QXnz8GzzPJP6kLryOukemif/t0ZkKcGYpbGuCNufb
b0rmer9g1u82zko9msGqvXTTTRxs5Bxe+HBM6pzW+8CQFrBumj9hFg+7BwE2v9ijuXYza3cauxEa
Qra9Cyp+sBU8oBbA86HC60twkU18tDKC1eRglZCb7M7dRsDMqC9p6kA1UEsZb6OeX1A/QpgnwFor
r38aXVGCLO2oWb2HO3ay5rG+Leg0cBrCErtQmlTST0VakpfvmKVCle1oyp3Cbfep7NzUB5+5McZc
eLDhynKFwDaat+H+shMaxu4ZIOtQpt6ZSFeY0lcVexx5esDrC40OKwl+prxncjlqg2M07Mk6uepi
SQd7cn4OF5aih+iG1sk8Fx5FD9l52z2uys/W1Cj0gsyfjiFxROAHpK5jqFZhUcWtjRArxp29A+yZ
ZMbSI/ZJhvCCleOhofp7Xr/HMx9XOgJSSTfrTFtR2eLWCFOVMgf2yoUdScUe7s2TdTu5GaALOCuj
x2P9iOs1rtrHv8U7w+Z/C5SjLoi756gduo1c/VaU9T1Hs1DrLGfgkoL+zkuGMrf7p5mNZkW3R67X
n9X7GavylJ/lP0TeSrzqkRGzeC8WzgCAbiAAfUkqhDjKHpkhjFU+T/xCJIFfuxFaBgnv0SiRkYPe
LnsRrBypyocVyoXMVwnK5yKQ/tu7dUKqpZdFVc82pkvYR40GzCUBJDldT6iWyEQohRtFJ7WMBOlJ
Y4LCGAhFMVm5vZ0oKcyjsM7ZCMF+atM49as3LN2Bgk6P6oUZv5F8/jKEa6JlEq2IixEFsh9IseOm
emCz+r4Z8Rdq6T0QaqgwSetoZ6p+o+09ktmFa6qnsPJFEDVED6l7iOfWDcoJCNnOruXM6anpIAVT
7uuGUABGBLie79FVlegGV1ILU4+TEwc0p/FuatlX7tRFmPFoBqi4qNZUgLibjqt0uT/oUUHvUK2D
+Qyiq2XvCzYKZeoTlHIDWd7+BCEmrHMd3pjjmqA7dOAwIdeY/uSU7saz9xxgCePX7VafRYhTIUlZ
AUbh+Ag3IHS4S7JLVDHXWCUV7lUphJTZqW7/QO667sSDTGnF7gKvc/y+ayAtUrAC2gPYAKPvTiav
KqFkSqJ1kCOAIVYGCGx/etHqaj4Tx6jiEiJjL5qv1TSOPcxuwYWGR2UZ+KB+0PsagSFdiqQ9PgGP
G++zbM14ZHbpTTBbPGhFU7IPw8z1XUEvY3A02wNQQ9Nag0pxAD3Up5DqY4pj/TVpbOxH2A/t/Cmf
Sp7+rigziy9ONQ4ZZc/ebzAMc5PdRTlubAoUe7fZpVOjRoi24CFtRyzxD+UoXVSoP3wX4ZzfKq4H
rTT7Tj+YWpsqokRSCPLQmUzG7Ez4LgYicAWxIjZ4oKYJUC4TAEdniHnk/nQRCnLXq8ja3ByVeVZz
jRS7+3mfOaRarw6lhIFYd7cMhOlqksk12dWqsMoHI2uQHshKbJ5M1cmycsXelxp1fii2YRX8tzJ9
eIblPPV+KKEhhfb+Fu9mudIP/D3/MK2Iu7nGIq44sfREteXlq9c9vP7AdnQcb955HnNmq4LhCCcN
cbzt6xAC0nekM7tvxKaycZ5yuqG3JRv4QXE/jL7GnGIDzYJzO7srnduCHJqg/uemejuUID2bgqwG
u3IMz85AqTIG8CLhRM+30E5uUL9UWhH5nIn5eiVamNb2GJ7/kzhAJeNQDcXNMV191LrUPUV1SuBO
VeMgPS3OCyFVocLkELDipvYyOrjWVSK2n3PrlyhWi3AXTknkWZunmnS9/YUhItOBhSt1u9+FgLu2
L5+nPCEPyAa8HV+RqKhbjDqGq3jIVXdS/nRfORYbsR/JyW6CEElv+7L2BmTnmZQgJZTPzK4lLHfu
tmwH9NSNtipjx2KGzJOup8INBzEOqthnjh4FZxi3KcgXTHquZ4AXOHJDUxalvKH1PhBZoHe1eHPl
XuYZPIrKpE28JRTJdFxyV5la7kyIF+MAqIOJ7u28G390VrXw5y0MgGujXNgEMwsHQMnSs41Rf4XU
xITS6pT6sxZ+4mEZ6VGgVJl6bDjJ9MFXD/7JzGNwLhws34vVnGs8sN9wU4gaPWjepvbWWbui57JL
nPyonYO37qtrsFMykeUkQ10wKdZPJAtPVQ9sxC8QOD41Do7bUJzO5dhDghP5hcVf270oPxqK8n8W
GXSLS8uV2XVc6Q6ncirdbxfqPMlRsnkvPQEuv5Jn2JrRkA+jweDTcb16uxDPY8Yibz5xz2rflBYG
I0XWIPrlDsgWW0XvT0RcIohOqbOd1B0Yw1ITXaLSigquHnCk2zqQAl9kONCocOgq6KCDUXowCpUU
VG4mpuophJ4+lrVIfsV19BQrukqBcrtebSYOS+00A0gsfuJYCHcxaNB3xE2o0EO/bidMoM9ghWRG
kxV2I7BXas2mltOSD0srusrtyBsqCJsXmfpf7lUIr+sCrdg9Og8meF8KD+sLrfbHtPSnqHL0vazy
oFzzOt8Mgm/EEkiWHnsj+oFsckHEXUrcJbf78fZWkWtZgL8Ttfn+p693yCqyYNXW/B+9DhXjvgSC
ZFnk+gsOpyp9qqQXUUtD8Hk4ipMaTuTPOxjVpRTTC7KfKS6gtL4fesV/klzcpZX7Sg0QWqAKNqFE
VY4w2FjN+xTQZGhveEiA76m01BtaqSc9QNn9g/zNMVXeuBIDAsLQBu2DW7N8t0BlWgQ2n3eG92YR
2OKgOxLomkqUT1YIXeTYckOA4JvmokMLzkFAg+R2S+emIddUCk+4wrGaBx7u3jZ49c/tWhYDjjDe
8yJlpLe79hEPpherJX6NJeIXnOcg6uQjHUqck7n68A7FdmNb/JCh98CUpb7WvnR/7cwV7OqRBIU4
58T9rtpYFNvzpRdj/mS6SwIF1nKiQxAmxuSmFKbOu7rkqEcpV7d+5P81OsHB+TIWsAS8COX/qX9Z
ctrS3U/Og4X7AsES5OgON53wy97N3OPN+uaMn30Up82PXMn/uLX7IlUznjnFEXK5Zi+KDFyFcG69
nwX0TPqOmzKMh3xd/0XhP0yAlYKx4HGqsUmerVKZx7+8lK6hmlojYlt+fk365CqP+uf352tbAmxh
KUttaxpXuak9A263O9ieHFE0xDZzASF1myZnBGuJOpYT6IMzLBlPUZeJfpWJBVswjB1DklyanXwU
vAF2RdQD0hvK2sShtUsE3BkOxg253Sf7ZiH2GshP8+3N8Wz8V0u8Yw5wxZsJG8TXwAjatRBi63hs
yyB+s6uboa04A5uy5jUVDReJXaRzIDNx6HBsWkxrl6L3Y8UzI71OXnjGUv/i/8qj3QQ2E8zkQw7d
8mof0gfeqk2D16Mc0ZcLKYPlPoQC9TgmSZvTsEq3Hp9Ot6leiZp6gd08BHFhRRB6n4FQBMoTVrO6
LRtQP5OLw0+hwSOh8OfBet+rDfUU+yIVsdSjjRChsnPgoSxHhTgnmvY4q6eVXE3O7RiM+CY5fyd6
MJDdQlufPu/VQ29qjJmytw1atpVDdA5yr2ShGSipPvbECWckZdGzjczkt605RkiX8CDSCJkVwyBe
HASQUmo+vZJs1zdUvaCLH22FqW/G0ap2rLvVVfxWqph/X3rZglfh8jYaJx1ePLEnbeMCb4vs1zx4
tSEQryatuRcjbQw50kcQaLH+Uxtw6uGAQH8Mh+rn9ieJIpVZ6ZNr4m85tClccaVvz/XyyNdSWcs0
lz0OFR1td02SMs/igyygRuWiPH3Dyz67Ww5LgNQotswlbaEgCESZA7n+ZQm52/Z+8iWuPappKm/p
GDLCriRBBXZCsssuBYeQhbnxHsolSP4TPUFYldV46PhjfY6na/xMIuN9DtBYzrSzrzt3wYbbnz5G
VKJBLkE/cuj3xS9C/YMcljeUTlEeR5rlyn6MKzJ+5iNcaX6bhJgZSWeGqzROkEkfsmAzsMIQIFa6
6tP+KnzgDeiFCA/gTFbPXX3x8u4jCn6xQYH1zhX0+qExjVtJWOp9rMEfz+jsvIk6+Yu5Ljrjwp5U
+Tc/QDqavYZmPRJ8zudHgXZA84TPQUeWivfjqD6qoi3p1R7ixmbUnlJh+4K6nmV1MeJSWOxlVDy1
mroSnGRIiSK/uNhUqaxpzac0bx4dF3aLqjRHRXt3MbIwrTaorIyCAJPbNC+9C3egqMnIPsSJGrEv
bTzUgMenhXSWsL+Md2ltFZMwtcqPMj+cGGzaoBt1WOW0fCwMq3eAEzbSqrdKWNRB4Ag4n1ZU3mNv
6ZzCRTL3Srvv99B8SWTaBeiGs7NAT7ND6mK1rJhNphEEyMvt5zRzcyQLuG1SVF4tY3pPHQ3CpJfq
pUfNAmrUvYzuT1gh+RuVoTF7sKTKb2kKMBJ66o6+ttXD9zL6k3YHSb0rtd+/2eX00tlHYI8GDEK1
1e8Qf5qvRP0/UmP6MymHVKXFE7zFBpUJW/rpShp7bfuLoTSdunNoDrt8fZTNKIqMVTBCipWtJH99
bt7bsSGCMgdEaIyGSKiuIaZtwinEeFI4szovGm/V1A0ikOOWQnwbpdp9LucnoC+ojO9SrVmm7Mzr
w4luFjNOxROuiSe6U13jxtiyPctjM7454CD2+Kpco+RXOGZNwHpwtPrEedHaCBG4TkJli7GGwD2i
2EIo5ReoegV/Ob70DvlILg1C1c8wUPGTijacM1G0ovtQJuXQYTHmRdpN/WEkmXgJKUdcgbR5P+H9
9Y/xXsok/4hnxpmR7Ym1AeAUCae2BBhbePLARGbgvG4XKtM+YfHQ3CEH+hwx907Bj+b5zqy2QJjS
NlbqEgpA12FeWEUMfoKexTSmGlfjrCiWs9Fq3qdWTlIKTZnx+ShcUJN8hPBbg2nqHb0/6VR4YeGl
TaEdq3InYijgYWleV7Gl7/04avD/BgEr17ofGlOQFEFkVhm1agcSRXIDNOQ4KYQPhA35xqbd93gs
2yHcj1HTnwgHda6sxsbzYeiO14fhGBz0Hh0KfyODlAPk0KeXiigHQKjiLAuXmpTzQeOTzr2kEH72
Xvg6DixyPa7cLVQLNNBdltzhoT+y1PnpzIknGH2u/GWUao9q74WCicLMYwlS6MCxRT1xHfQROX4O
NC/TXALiPHeY0uOQAmRCqUXNPPCjEaVlgYcr4aBt/0s30MTsgpt1hnoxvqtTdU/2Ie9KlGSVFT4U
i5ay/htfrF4uqB15v3wXaiBGe8iXMjD/wd9ZnFHc5Scv3u0zyVK/pu3DhC92Tff07qVMeZXNpKW9
4lGP8qet9nJ9ytzvzwA6o1hFNQGO0V/C8vKm504eDHJJ8hpJ7r7lCff/aqJsTvXdEeq4rIP4qpMN
W5jWAvj8JnHDDXwYW710uT+yS6YDK//UK50scYmuL/JQJ/ZmbvrjBD7UezA/QncIlkg3FpxDVa3V
M49Wj6B5SS1NxeRGTJSVr/oiJ778LFTNmsXm1xnqJ2dOKTEy1WRRR4/arUjsULXVCpPMkOSZiGiv
b9bsZ4QtvFbhran3j9y6lme1hdvGXbGdORFEBJzdv5wYhIRHpuiKG8KhQQ57exb6r2sit3y6xrfP
gFYf870tDD526xtHKbYPVdCmMPfT05Pvf3JplqQakutC00u+gbNNGrBX3L3gHwdmoHfPYqWkSQ9w
pEidbgucHznoksIzDrY8vlMKPYPPy/lcGTth98jyZBhwaDgv15cuqccUmtPBCxS7cxFkAtpe6XXO
K26/Edc40O94mqecw0QylKWo0pck6k8cAXMTyOBZkLvfVaislv+lF5z3ZdyvoczItWo26p71b/t1
yd9Oe9PRZ8Kv20YhkWkJ/4DLy0JFbfY/fbd+yISlAi8E7nvmvwu8x2lEWasfKmmmLfIu7x3/7kQx
eCVetuaheMsLGsuRhm4BUnfVtc9hKTtXn75jbfE25sNnJyIHoF71OUb5UkfwbjpvZ1/40mHDIroo
PokJ/VVpSCIaA6d6L2F4N/fILWKYhnQCg42mHUWbjjipIRDUS8wGkVuUr+FikeDJnWUrNbbFwEiz
OIlSKFUBQBwrhZ7ARw8oYikrbMrSiw02xus7/DsHKl3bX5u5LllWndm7XCiC6IW/+tPAvFRQlz3Z
5338RoXOXqfDsZQWGsxAYoJw1J1mtyKcdiOpttLbIHhasZz5MRhWUKZCe9UEBvv2Iyl/MOyxUB8O
fMlz5SOBT0OCUoJcrWr7kHTJmto39kKsc6RKP1BBlgYhiXjwH2etDc1kjJK2VS3N8O+FMmmCmTcp
h1zG0dRgD/dEY7WNtixpXKTod3DGI86YWlwImOLueQZqIsFPcuEgzDW7o+0uL3cPBgPrJw6xXNDG
8Mgc6a6FKeCHuMKkTAT6BWoZcB7pV64nf8WKk/GCY5U2y5d6v5TXHmq8cyo87QSzrh2Oc6PZK947
uzZvZtKrocA230j6pb4rgWN3mlRFn5kmRljnebXIjfqXFM+uadpSpGJ0ek/x0ddMmK9+/xBf9RLF
4J9SsIPzAGeoPrVyuJLSffPqEniC/MX7Rr9JGwO9WC402swTdH0G+Gc+akTlXsBQ7FK5F98bJ++t
AxDtC7y0WwLPnQEKX1rrA0Pu2k8k6iDp/eUY5eBDqSyHONDwPScu9HZwfGfNHYwDo/1IAS0npy25
6zvm8rjXlwTtiBzmZrHK7dsdU5SfoJDZRN981L8GKVJ06NJYUvc+8+h/GbZcqlNwPbcNTdOmFWxj
cZKx7eafBP0hKPAqq8VrRcRQs1kDRQhoykgJqgZkfKNF5Me+EWQwhvEpy9qwLTMxTMxQMrI8RggI
94zanAuAm1geuoO/Gl0CB+UwNs/knHb3HiyZsfBxnY+N7KuiyGPmRonf8bqXgq9MtdQracBDbN3X
214Ha/PLkKnIz4+olhz3L6NqMHJpFxwqNXA8mUvV1uKF1oKx3Y9CryRwzLonGk0mthj7WNpgqFof
VkmgiHSgFNF1tzYQJ2eEnJKony2AIemGVrlfBjQMT5F7ZzsRylaUo5Djp0837cMZgbpvrccT/8yy
LD06LM2QNnJW5zAABpL9ycmr3uvnkgiHPZhDFYtdakKVXaezyDoz++5iHllS51PkXqpNHk7bkvwc
itu4plSpZ1d+4qMxXVd1W9l8Z+HNT/ghXhwEZkk9Wv1mNb0Lnql1Sw+iCXtwzPJGjwgR363GS0KA
ALGc+biqMyU2LBGetfQ5rvDzdL7vEGwkr9umhcdvQKkXB+lxnS+wL2jpnaG4xUVwDVv4IJGbYPG4
UOE7/BmoYMD5ZipA7PwhZTfsXdW0lzr/maDov1MoxCmRQqoKM4SJn1Mw8210Ud4gkKcinFQGlfPS
UpCETxnlYedGSODDcFChCWAT1cElsDlwTYxCbMmhbPcjRsEB6hG5uUJO1vDZioKvfRpbHycoXvUA
ghs30DlXslzrdHHd48kMwOmuk+Hinf27O6qLXGt7Xj7qnnO6oSIIeZy95WAc8IVhqWhubVLen04x
pbhzPopo/0t1q4JKlJ5qoOxnooHyQIunSvEMpO/0+Qp5RXoLgRhMyaicOjvumavbSz1i3WJthAKW
bP0rlodBw0iKEHvsVlBGTaOB1wql8kEi9Z7uCIClDHSqEa0khjXtbLgeB++3e2BchHJ/RqyOAUtN
3bMr2qMQrV6lJBeUFlvf9tWJYh88sERCFRVsaMHKmhWsEhR24BbZkgk3GDrT/RFF2p0AaoZci7ED
58b18I/m+MbEIBCMFKyvOFR+XikECyGugiIYCFPIT+Nr99PG2LFJiQow/lWDj9bVSIZWhPkVtrqJ
0ywgNh1kK4V9S/VAp6t1XonrbRkuk4NWb01eHdRIrMdF+m91EdnKF1+9VJiZ/pa1HC4RLDfaP8V/
mvGG28IGU2UXAA4yI3l7oSi6eWHBZX0xchobYjpLg6Vgg6E+RP8U18svzzcw0AFxfSeurC1R38lM
EDoKsr71RrmyfYi6nju5LVIX/iGktwH6ObDWmqaG1eXV/ZsIIpTl773rwaSn4ddE9VYBd1YXsgLF
dWpxFO+BDLQvEYNZJVFhARZB+WKq0m4F9FACg+IQrsRyjbHZDB6CZE786wKeasF+Rhaalz4td44r
Il+Gv7Y1dQy3NIYb82KbLfJ0FqFmkOIHmYztSi6VoIbRao7YD90/ZRhdB6TO3MhFUFR+USrfSYzm
4lTy4G4L3cKycghyHAzEXrFbynt6lzRWXziDolC9OmQkBpJIzX3rz29TdoWCZJUd0eIEb2anqlXK
tNxlXSl/CdJTqw3+lpgD2WPmTycxBHfFuSMyy4DpmDvoSwVxNMj1+iUvxYtAl2R6JCTAQNA0z5CU
QPI8gIE3uGQoyn0Lc5jFH6TXZAluFg1IXdodqGEf5CnhN8DceS5v30HgaJ19GG6IY0MyWk1txNag
pprMWYMsG1tWtSzpDqXaNIEhrR3R56lBnPQzBCtIjiJ+IRK3aDayvhrPTCbZjO+/4kre5KBFjdET
Qqg1eVSnymIIuWngOWINZm0gKBPoYFnV+J+TomgkzXOrmsxWifVQKd2//Shno8c6n/FQ2zNnRwl+
ok5kfSD7hYLmKuXwPIuXdhuA5KCRi4BLA4LDbAT1xBEXYw5b4DBBsYz9A4gPOUF3X0lGHWlJvyL6
umA7AcBecfbZZTvGQ9+9J6VXA+buA2rChhYoi0vvrwmQmds4oElQaSffyddiFg3J2bltwpIiA23v
Ba71kuVIX/njkmzJITDZuNQVPJvx/lSAZmmB7diOdXXNaJyBv5/rQm8ByFd834zwwMZXhISH2NmH
OvkLU1C20QBodfaUI7c+JM2jNBItBAf8ygDcvzzex1Hz8ukYDeTE5v+E5/5YJD78MI48gNjb0Ymg
SaiNu0HW5BVwD/QiTuUawvN6AmcM9QT7lKz7cC7pw7ECn1Glb6CZTnmwRqtuT8guB7BW/rAi9F9I
a0G2cZQyHn0FY6zwe8iRutLCKaye/EdoCQ6T6AnhIgf5budyJlqDAGxEKONlmhmkX1eFukXRiKJc
DxbEg39dNS+zC9iTCj6XRhVO3CoKPPfjFAH6JDzVTjhYnTgMdiSoP6BYuGa2ymonXED5vw+aR/eo
KEb0+K6yfAJ6X1n1R7jTVRq30FWj3FKtovOuuzZjIat1Lz6XGGZIbmi0gyi/2ftz4YAoEHuXXD3l
yP1YuUhv/i49vu3L34zJRiD+x2S/EeHW1NyZ3c1qh5lRWUG0hdB26Mw6Ivmfdl1C67NXdVdj6Gne
N+8LJTLNq1678fZmxZb1mUEP790DymeWTIMRpK3BtJY25iUARD6hlOC97YUe8B1yQj8bXDc9jJ37
+kH42uewRZqIJsgMTi+wrQv3xJt2lJA7h9pQZEKkjnrBoqu4xJ4AIdqxGY8Lj7eJ+13omJLW+1Ha
N9rrTWLAKtTbE9wTbHVTRJc6iYgltWlSI3u4gMuZF6zx+gGmx5sw936D1GcPSwXZFbEygvjgDIfM
O1SXQaJ3TFw9xH4gtdh9vm1ldA6TObFDRzJkmlQS2razaqyAfkZoU1E6YDx0rDarzNBWzNkt1fcY
5K5zyq/p8U2/I8t07mvfPM9U5LlIEog/JLyvDvkZbIlTFDNc1f5B8MnvsLjvBljIp9Zhe2sGYd/1
N7ul0mR/xC059vdlWTHf4Xk+ze3Yp4JIn3lMzWrpaDBt88TVuHhxZwldO0zFuhERYC7MXt1OW9Y1
yke7dzD9W1UTberNX+M/YvGnlMAJ1nTN6ZGqz6mxCuHyIJuGRo7dByJ7dALCexOrL9zpIAiFc1HG
sXhTzkqwwsld7PwvjIlKGyvqhFv2lgr7AwTBBWw0keaUuzTqqSkHbMukuBcOz1kBdvRhjqlhvtw/
tcWIR1g6O6DRkeQmmC43Cy3qUgGCZu5Gzdee4ZokWFytvLqorKk1MVrrNiGfE3AtdNEqhc7siSY+
nhQ4oCHRwSSMaF5W/Nx69daMniQUeKVTcl4MAir483FkY4/FAU/o+QZDd/6Y6h/h/lQUTUwh/JIK
nDzbL1ARwSLe/A8dHeVNkiJmwvTKndASemy9cyjUCJ1gtyMvGHqtAoJp3UcdUajHL7r/m0NHLdsi
8TEtCpO3c7ZMP/IFG2oCD0D/W1vucyZTlEWWP532vqs2fV2c9y04r0bXtFGBV4sAHS+9OMYPhmS9
9scXBreK6XZLSqmi3TSvdK1UfFq9/urFzFOTcWtRlJhzmzuiNeYkrSTPi0msadCtarB33TBXhRMz
OqbGnvSyIqIsnKetImqiIzzSMLr8ESxtvi+hNiu78ZJ8lPU+u/OK4cby0NPd338Fqs6p0uYAgOoX
0slL/3/Xcb1kWU++cZVK2/o4ghlLeyxiEIe7S82ZVEOayEKLGPKp7Gt1DEDQBzyx4RyZNONRZeIG
oJ2A8YsK+Iz33df9sisdDEbgvsITKRSc2hPYiYypyb65Bas0ivpmzzsi7FOySB4j86aECRBAtOzY
jC6vP06hdVneUhKxDoOoy9eR6l483hc+8MJsLSxHh1gnhmBdMBPoxY5o2oMhrTwxXnMEiX/QegPK
DgBz68FfrvNmzeHrGDiZ7JhxadydVlw5YtEASmZSk6jA8LDbtl5/xK50p8VjqlqG7+T567ah6f4z
YbD+7n7xsWIF2oZGblVZ0dVrBBR1dioDpgmjP2WO406VncT+I5ggjtDrHYi/40OIvnh1aMUqOH3e
64ExOV6gR8jqO+5X0cIbPySmXzPh9tC7GwqfsNmmgx9/LoSWJ0iK5irtK3OdgEHP+hUEV0KThLyc
9Md45lvFlGsLVvlf8mlCdeybWU92MELpjyMfrk1ogj3GVEkHmHDRKr/csYeVhL0v6UUpkKPsiEIP
7HgVpCsz30WNXI7j0Db86ysUjXfT8sy30JzDaja2Fj/wC23ZAwtkKuJUMR7fiiy5lFnDXrIi7Duz
xptEibW5RZkHnsgSij8oAzCmSD/e0c5/vodyAgPydtZBr/3nFO42qjHoH2wFLs34gGg69o8jKV69
DpeDWJNJ7uxIag0TvThcNO/h9qvD0ijZANTiu7AqPFgdFO0ODzDyWSi7nJA6b0T2xwXOb3bcmF7I
4W7vUqi7Y4QPZCR05hyWeu3jfbRtLn5pjsxZv1oiOhnRUvNZi0rCa4AL1OytP8PkJdkGj7nln3XX
RTDmum0JF5aymexys0GsTSeB2vhnXWInr/hodXhRSMNTD0A2/Xn81gHq3TPXS4yZWjIbSsvZIT3a
O+BsebX6VwJg/xuHLBrQ9KSebmT+m39bEpQm1Yi+zEdgf4eNjxSgwyr3aqEtFjWf/ZphyeN7pkQy
/h5+KeJL2oqWfifE/wHMEQBpQroAk56x0XVL1ridkJK6613o3Xikwb1eawMrR2HXppHnDqbpj7GI
OUE1EM0nVVqGWonIzztGg/5sO26XUTfSVGRsBITnCCCGsdyPiaVxMSX1hK0jz0S+xyqlHn6GA7bE
+VGR21Tn10qcneFQU0mKtPn7IdBhJWj3OLJ43ZFQc96X97++zpXfS+GNNQYLorPjjSQSaU3sIm+J
lUxfHBU956MUPGyWWAExb4H0YFtKq6JQfncNXHC6LNNTDcibX7DI1oBUS2a8q05PsAeECYU9Nri5
0Wf0fgCBRGy/JDdLLSZvDbWZbjCK7zVReAgwRdczdp546DfJEgtgDQZoH/5Q
`protect end_protected
