`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
PeqAACiKacdbMOWs2XqEaCOpUVm6letI2uGLDiD9lX0yoyBIWN0n2TcEOh3r3UNckwNHImxwRo1k
8kO4TiYYhA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
auZzPkb3r2HppBydOd/o3UXtK6rJTIS7GYUl6UfoNc2fuxKNxuaX5fuwuO2C/xW9Dwhj6txvdXSl
6P18m7eILIWtScQY/zFG6rhvGQKvakLwLjdAKDz9A862+2PgGCnRM2oAlF5f2cOeaoejq4NzIssM
trMP8apt39JggmVZdB8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
e3IEv7/wkdd2X+qJoUq7FlGbH6ss4+2Kprvx1c80iL0+RtyfFn7gRQ7KRscg+b2pSX30CAA3rZvD
CipsqO/c9bZqj5VfXOrjBqJgQUrqinfK3Gj8SXPHczpmxpnKjMxM1XpBs1v+GuafN4/8KAQ6I/7A
Jq/CcecuA7nqnwT4KVIDPnkeewZOWMG0knXp28/+fOLVIYeEjEvtOerZiTizJTtPwmRPVBH+5Hql
/CtHgmxLmpitZvSNmWW9DqPhkuyODcInEJrl4b4SGqksRts8kQ0XcHH3B397/Q+FarsF7xsdta1b
9usdtMMhglSriQUPZrBPHJXV5L05ik/uuXMlTQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
LnIK6f68C0hy0aeBngl05Oyvlp8vnvOvN38tYskLxxJBl7ej0TpYYaSJOAL2lQ6FLR326CCaFbhs
xgb+zjGCGs+DNfMLn0hgRkl0RBaX89Xm/iK5zeBuUNRjw6QgyyQJYYPDbwCrfTi3xoJkSoIOaHFd
3wNNZCBA2WEnHKz6aJY=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CeNA35IAS+fDRdKelCkD/EK+Ucq+I3G7pjPDlBGYhFEdN5nbyHo1Tmux9xdwRIy9QvlICCoBH21L
SGTVHtQEB/e0aTmfNHUbwSEwnHaM661voBhLiRTU5qQpjAS9zNbKrA5T251UZIbuV7LOoXyp6Wn7
yLcqDCJ7nNnXP5/aFaTEPJV72kevkZNB26SVxFU+ysrxXeK21y6rHIU8tS9pfwjRqFWl32wBNBZy
c+7uxdI/r4KVmipuD4kHmdb7eWXM6MKrMSjlgWvKiolj6goWmzi7SRLQT+U66YMNp8BfQ4XlcT0c
X8Dx9zPFetvak2ROciLf902FNilYtf+vhnmdWw==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
c7btEZIH+CfFksJLkG9oOMqjkJg8WlX8pEmrfA41RU/4n9cvzFdASG+OulihbL7e8ZGDk9ye8tF6
4FRVQH4GOMia26DiobkTbtlNCIbQNYQQA0gZqATjTqU8oSo3ORD13OWR8ak0X8/ikYV2tHfqKP3v
AM5v8u0JTb92RJ73Tu8S4JX7VYwvRstor6o2UOK2t5I0EVDSm0q3pIekgq0RtSAfpZcEmIQbR+vD
Qi/qtGGFSRYICGWxK647oJL+o2/OS29tL4cj06NQV6MlPIUUyt0sgT2hr6dPjCig4QSycBLh5w9J
KvMskGHNUDvoszKAr2v49s694p/o0Vt/btsOkg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9264)
`protect data_block
EflAiSgk5UuDa3iO87+I4FtQ9n7oxGrEmJAz/UOBDusDF5JIspoP6YeQPzX6BeKLeaBB6wFHX66f
G59iwNITmHbcGn2pH3AzQIiI+19vr+fPsEriK0kiOocMKCX9QQuaehpXTghf1CCfCKhVAFU24v65
n+BjdU+LRTPK5VNkBSPJaUerstKXidFtDWzax7S4T2rFDX8FZ5aCVmTFrjAqGO5NLO2tg6ibXO7f
90BWXrdXapsimKxwcjHY9cCbA1c2Vt4OjLXG6thCTqgkZpwOqQCTkSrJ5nJ11h/C4FgFlJ1ZPV1O
ublNpxINTEP/Fm59U7MrFmr0jAS7oQhKlZUkcHdtY7I2dziXZFu54uPX379xA4AkPfQoErQdulF/
sWcJsXMIbQFMUTDU6XmmrKPXikGYVPOQtbQ6nE/4IO1FMERl+UdTDxjrxhWfmI7ORio5jbjZVYn1
50m532QYBbg846dclg+xu3qipKRoOxMgB4hiHrQ1OYWhgYvFDFVdjWqFZDoq1HmUOmt7JG5JSvT7
AYbWTFhaqtr1ANQ7J+ayuVHS1tl8s/XdNIieHThMi47lTTdYT9o6RALqKkIhvlP4mwmITpSz/GYz
sx96rtKdChFNs2P5Z3gsyzwibp6GN9oDrEKJw3XngKRandUVRiGKUMMW1VSqX3GMMseS4d/xVInA
Xyo0xbR8WXTY8irgAzjEm8JrUM0OMvA7ulN4H5YRF6/JfffOoFwBmM3faeX9AtCj/bDRuue8+aIt
JL++qHvCBwbS40ke0FyRNxGgKfnn4/FHbuYuHeI3kf5ksC/1fWCYcyKtn6OFNlEmeLCZ6j7KbeuN
Cj7Q+bzNhdl/Wvts0KEJdRSDqYQNmm90wTZqCmS4Ip1Sc4PIM9ObNQN9KhSi3iOrPuwK7yAdn2qI
DMzirsfELMX3Fx7DbptshVg7kLRQmL3PTiWYHWuKh2E/gNZ8Zzh9zkyBEeZRaWi9bCXE/+jG7sqY
Yjt7h5cSYlGdwlopQug0fQIlaGsE1SD3qdE8PFanXHyiOe7XiWV+2IkeUwtZNOucwfxDnIP925X2
AoWhHt/O+8+443QSoDWcra1mQ7EUdYi0ojDuQJ7I1GdMbL3BJEMAlYiFFWqKbA7o44zsgP0kl78l
IbVt4znlaTLxZvTvPDA+ereobGRiJxtZjoWcYdLcE92Ua7V8gbyeSivYU6erb3kpcgoZfUuSI7LJ
OYFa2mR57DHMPhRfrKPzCCdqf4y81qEWiHKUqS426YXBSKYQlyw/4U0w7oQzfbugzvl0ecPOpUIR
lcFwDo5WslEPb0s7i87lp1D9TZlfPM0luY54oB09Ynm69Hte9NyRKuRZRfDPTM3Tt0ACVETY6Xrx
0/mmwqeewZ4WtqZIB2pQWmIfpmt7xJgHK3MCq0B6U5V3tpIKM2ncE4p5km3lKEa5xMM+aXKB5tUE
b8hOOyFZBVID82EcXvXHoP7QYF0ClH7WHu6S/wQDOgUR69QM7cZPbPOgYAwIefSaprTtqG37Bhe6
qZqxHVzk0w28ghfF28Vscwd5R4xTeYNYPQSezGKejkJYpeoLXfDKXDbOkS5yRed1X4rJtv0p/AU7
DcUJqJkyxy3NA9VZX1OWPfj1TkXud9vkpl4h3syodD8Fnw921+YQl64PRMCz6cFY0AgPZTd2++2b
yaxAsiW4ldH1ftdXhJkGc+OVe1XUgiHNxdwg3QAY63W1B7NAf3VQ3jcfpji7IHrqVnQ9m/6TqNv6
uGa9uqubq9vZ8NN5OA0hyFkaYUuIKeJcofCpmFYzNF8YzDMumEr65zmkAzHv9Ubt109KODjqiJTO
XjGNltZ+uPbi9Rt0r+mtEriP6+Tout0pzqBI95Hj6v/RmuU6RtkQ3JycBAnXPZXS2+/ZEYE2gt38
OvMLrdtsoz7OVFcyJUNusajO3jFeb4ExB4KR7I2RQgFKCRmpN5c3aYs//Sl6oZkPGNRs8rLX7jgR
j9QBlWPlDmKluXr5xl1HoUfPWW1hRRbg9fWyADBMrIlDI9EmEWxO9ldD2UnR0cLmzEB5oXV/xo2S
h6qfJX0B9Uvu/KwTkrjcrNfQx32hoHGb94h22aqxy1RcAgVE/UpqDB71wSMzzFCadQCMUbIdB5yr
ztyvYHaa9Sm1XefvS/JUcvnPuhmjRXggjJURSksvfuD88cjRp39r63K6ckA1fwny8/PSuVvyooaa
uLQ5yP5cS0UPRekLXGu9Qs5xoPnxGZn0SD3gvr4wR2CJKOeryBbJBLbnia4te+nMSQaqhTUL1sBD
Gqjyw75iyO3HKIHM6CMcfhU+PfpsdyFCru6H5tXeAm2HgFjNkaBxtVJKWQdp1ASPwYFB245M1nXM
XqA9cACcqvRZqERHsx+TLZTSnZhnJKA8rqY9pN42YYlJRB2UchmAUAN+fP9cypCcMGC9g4tFCgmI
BaPS2B7QrWm0mg2ye8BN2uxtbsMZO0pL0DoLe0r6/HjwdS22VFCW2TkqsYI8gpzeptqOGDqDN2JA
Cn7jcAaJpuyFwFxSadG17zLLimAwfoPej3TZjIE0tYSOf7LbRBIF1yC518x232VbaM4ZRwDZUl/A
VzN4556tB/SwwYidFsEw0s+xZWBXtK5ZFOQNEQwROYtEvCR7b+Qc3ClDBI+qQGVgk3sXIpz6iayu
em5CDNwNc+lZ63T3JCJFN7vgR9dvxzIK+zJVJIvGcmjcN2lYEs0MjCf9OJuA5vB241rfz9uYXvxW
rX9g8AtTN+Sjc0rh2ppozIahlVHhQMkAR64Yymh+SBG3YYIsVx4oxL1wWkv4R4qrgb88z/AgcLxw
Yg6qlsMx1OXTu7N0lvS9B4zGy+V4SnBdlaT2CaRtvB+lagKkF8h3qUR43lwdcQdZYRs5ked72XEN
EQy2P63sF+pXHWEAaM0WUa9AmLp1HHK5VQVqhNtVDovPWn1Gh7zdSn0DN2Jm3urVvzFfInGojpFf
LNpxAGdz7UHGFyH0goI57rtiSA73UD2VnaG3pGhlioxvYnqbX4yLx1WZfqHPe3CT15jD6lfedYRN
oo0Kdcc5i4S2zMKaQp7gss1H9z2pLJ2sMIgygjUWApS5iIdWUJjiTM9sE16+Rn9USaAR/vSFQHoP
Lwu0lxc+Q4h+F3gHKiyeuqyANPdr25UNsA/fMoWqtxpoFpEoF4ItJChCglvQ5bhLYUBnHShPgW2z
QQqLYYt1gkxWeGvkFstTJVSqCY3QCfCnrqwe1kjgGgCTb5o/s0pCAyoaA3DGMYoP+1l+yaWddwh7
mi6aK9aKscCxO9WD3Nl9cwYAW+yAWflTxo0ByOuFS75F7U9ZVlCeELnTdFnGaO7y2vJdOOsj85Cy
qtEaU9+rQcgMYCarIFKDxUCjnSuZP+p/WX92y63zYnlXyJWDo+4bWzjGv7o5lhRWvgAGVWtnmkA+
FQUyGhPiP89Yrbiq9wtSbi51BhZTzd+4MVq4ur92K+eH/+ePZ9xp4KerUlinOSWMaaDwYdtf91t6
gTqJApf0Q7r7EX5lYbSJGZGoaDWUEXfGLLLeiF0EUw9I4/cqO9Yfb6YSG3N98A4wFfMRSYOB46vx
K04P36+cDMULJxPiaxQiQCGcXR3A1z126Ea/yqmHYRgDJIPflTNukzZYXB4t0de0a8efeaqsJGDE
xgAM0ugBDW47nMRnvKbxlhRC90kuOfawLFK4IG1MYSgQuRUPV39+swLNxfx0EI0mDmXDz/8YNv3U
oRMZDoic7NtGX1LNFux7K1UCarQOMDJABxtDC2OcN85H9HD0nlP4v2CwUVcMot0ZWvCNb5O0o4L+
D2mSsAaPzdTl/8HntRbvn4UGOHOaytA22FicOaAhkRbZVXzZ5ZJdxDTId4gAJxIrC8E9pMNW8tAD
Nzu4/iaVXtbB8DumYbYWkYNQCY9yh+wtHV8OQZwTR+PZqIATakJnYFMXFrKvQmzmID4sFuirp0P/
jRnnbFLCcFZwS6a1E0n8K/jhMNaJb1O6wQxYxw79phTKcgOufGIxj7sgOxRXK2vMZXs/At6eulo+
72cRz4Q/2+b06tYhIByBlzrkukduSCD6sFTF/QUJWkPMxanAxMQMBJ7di/sLU8Ho+gqE87HB8gO7
PrPllVskCj6r7t6T5dWwM5bRDs7g0NUsyc6P2JW3a5ITB/gophxkaU8/wAAEc0LvxBWo9TQf6adc
hjoGLoOQSGtf7h2jXqebtXg6Ei1IkQE6xOy69lZ5PqhTurfuzuRyFIAQVdfSxq8aH+W4MqWinOLk
9RDzfIhYts3/se1uM/HBaF1l9BzYOUM3ls3/KR6JxOkL+CfvTc36gbhuiwJmif/mmQBIFK+xRFqy
ve5+Np+SQkAC44b8bfV89oUkz5RzVtRCPKf4mu5VZo8lCsXol6c4PD7FUsw1eyKNniuD6hoD188B
j0MJh1lOVBLJim/2/+G1dYwG5QwC/kJHu8smXgeYii2PK5ivlTCtb3CMxQ7miboQyRWZaXffSFQD
hvu+QtpCMS4yqUnzA9ceHe79ZkXfFeCDhjELnvcW9NTMpmHGAj9OdObTkVs1SSzX8N/52MfAoWH4
e4a9aH0KwxoWmzGBXYSysYWWvpvSswErKOMEzP9cOGkdltHNZJCk2FZwdhu/0kznx+Y1zJl22tdH
pKSfUwoIfrqvKO97bImh5GeaoRDyDZ18evTAh9/ImN7GPsaxR1ibPSZ0C7inX7VOqkDb5YrhDCJh
bTLTsmoSo6Qdla1Cm9Zp0pfeDqykw6O7j/alwsspE39A+sHJwdzJjPqMYLl/Rjce0GPYz+caX4pO
MdknVDgsjCM9HscVubtNrMUiD1JBt/HrdTpXeD50QzOHQNXtgcNM0ABSKWw1gf5aX2smKkuFUayG
dwmyB2D6/Ec7BjMrVZv0OZuxBtzNuRDpghI+rMd8UrkYZG6PCT8vxd22jhoULrrrGsFJJHw2Hxyq
4SEivIJ8z2qKelVyyL1Z5E8jRH9FHeQJgA3xt81P09wKdKe8X+L2mjUv1PH97XqCjgVc4L1yInp1
O6i1HL2QVhW1LJckvdIGALDFgtXXGOLReX63CWtvDZsrgOB9W4K1cCfLKj/e3N9LzclxhNgx5uhI
F310gGuS+VWviDjAtW98/Cy1h0lFwSBDh+N2AOFSWFud2fkkH0nLG69jO1c7IqhGxTq902m5iVIX
oOPuTWn02JaiaSmyoWsKyj4DTcAX6glyZvA4Sg/v0fnOTb8DQpOuqqiJ9rxLiz7pu1i5wvDwyP5g
Li/7H+WuM4OX85H42IwgSPfTRABW0TMztwR5LlBZRiXazfW3+L7VzCpCEFJX+lzsO9fQixgv7dSv
biHyklpDP3UN15l39z8b24SdaQnSdtKdgBGdpJlHU7A1JASfqgrx4OleQm/KpWbkNKeaQFpdN6yn
441mEvUwRahQroOPXtkvE7lZay4LnhaBpDkcOQHnHwxdJV+S6KBeVc2snttNrq0bHavStMYnu704
YJQRtWLBNWKMMy6d5Dsp/ARORa2d5++wTvmSIg9IJFARXZ7Owami/qt98ZolZr50TH8BjkKEON2z
gkjlWVhdAsvH/+z8nu3r9htVNkZ4heuDSvuv84os7SjDlRBQrakEXmPaOfVzlNfM3f0T4Y+623hQ
rfAer/dLyQziMTzT8rE2pKezqpSuVGd1uHxDV4ZKTNJtxEAz7J5jPVAmTFaECj5wESx+JTbMi1eC
7AXB1f1iqeJz0RSTvR1srasPTxFk2idsXg+gDjoYCDgD6BtmrbQbHnMj0cHztq1+zrqTvP8UFROg
zPZAjdZb6vSFMj/feicI8VcFKb/jQ6CtAiG+lwpj9jOoUQwqUqMokLynPbYeKCQq5VpPopRBInfc
+esWbZ5uQpX9FLn/lgJYlyTyF0XCg7Lz/dFvRRHG53l6vVF5V+fUuNkn/wP10N5rMLiku5Izui53
44XjYIiY/x19O2zFLaA/cR/9TDeIuOnd5WA8tUgEX1FhPfNdlPsK7En4j2L3Qj4dXAYUj1QeazFf
aYpaHQravyKz/sNSC53juF47aNsAlQ8tB5cvLJROEWxbvKSwkfjC3OE3hvqOmEas4s+WDqQIlDMx
FeP5bLxjCFpwg2uttOcKR5+vcDpUj/YgF+EfxYp07QHGgRCTXbgETT+lLCORXJJXwg6/MpuWrwxk
G0OAIHZwnAgr7Uh9jfG7TN7+XE7RgBXVsi9D+U7orGbmArz3eFnY2SW2D95uyaYxgCwqYfBb6AJb
LmhtXcbM66GA/VvqULRwSlV7fi3JyWkRBWd+RIGUL5t6FyedLFNqKVrtayf7RIY32ipvkd5/JtiD
EN42IF8IGcFolbkxwzyvmoGBAgKSI7plWkrbkfZiSHsdlPkGBnwESdd4W/26wM3VZbZ+oBtR9rnF
jUvxBWf/r4aOamGbSpOkgzlyXPDrL08iMPoJuG6le4aZhjGugjls5mYjx/t7DVSL2J4EH1izZQLK
54TzLbLhHPQoG1svh7mc4/9INLkfszBSf/HylBPAmE52NTQbE7gfIikF69ETjosHBfQoOxUsGMy2
Gg58pwzIe1Ser+v1++wn7Bn0MeMZ77eHgFh5UVTtuC0YOsdUrcTy0QKR+EZvY+FIqUTxJruIFtoO
gRxhwl57RzzzJP7Aqs9mMNa1n4uwpbk+9ehZQUf3SVX9zP4/vszcqyN9VSg0nIC5N6qu262zKcoM
dm/yh9TipLXw4nr7P/aO9RXjHMjqA7tn4VSaVpged+49H6YbZkpTeqcacEGEg241gGGir3P1e+39
n11+wkUNhi4E9eku3RyId4lxTHOawAAgYhTKN54p3VvO7K0ITP82zuAqEOOO3NJ8cB4C6q2iPJFX
jyF4vTlRbE8JFBY+dj2lnlR8PVTUtFIVBFzfJkjHIiBXZrwW8T79Xx8CO3iO1TsQHY8ypCz+Jyq0
jUpMF/hEYXBRYg+S7GUXXfw0Gm/RIz08hXT4ZWyiL6wNDq6HiSb0Jpl4Jy5Rw8fUc+43MjGlSnae
SZEzsQr4VkE8ygrpGie2x08l4+91zoZE1TBitCiiDXjvKhb6c6TjPXG90bERkAOd6WhlXjen8d8V
/aKFkaoD77PYKdeeU/3nac4hndvdTGm6xa1IbkCWBU/kFHQiJsPTt2d19ol9+iXrHXUNvA8KtHyi
hMe+1G5JDQbTGxn91Nkf4DVqHAkrhkiSByN/mv4PJcUwWg9MrWSflPKYHUJjGJ49poV0jNvbf0EL
VPY5jxuNQt60tbqnWLQwJbGBns6p5s6I5xaZ2fPjnFEGplBcJF1dDEVnSDM6g2YyhsRn4JZDsCz9
5TBWnFEFB8VheKTSOpu0uIbyOL5eZ+0gptMoUASXaFymutJX680mnhPQNbL2kvcxyOFlSn/1Ooxx
Jxqu0OIUkgHOH6bIZzOMdlvcaiz360mW+Gk6qdBbsMVkBUGDEsTDrxvNmjqUs5uXn2pwohXmAggX
Cw/DCyzIH41QCJrOiUUtoNzYumAP11BwYfQEjFaj0Izp0Euj5xw+UnK1gFbTm7AHqdkQmqtAh7Uv
h5RGa7Z8Avo3vccnYrTt/PCMBq8BKeNMQv771/mabh42D73dUCMrJugfhGHAqI0JMY9jZTmzhraS
uMz2GEZXTLrYf4ZL1P4SNW4O4m5+xtW/vHj5u7WVHyIwNCj2ver1P5fs/1uWRA1EM55nKpQIbwp2
qTiu6oVeoBW5uUma6W8ZoGM8hzg6TQRL3E8Z91ZkF5sRYVP7mWwCuOj1VdzZcOdiR2VCEr7uDD33
IEHz8/Q7M527qP0xs48gDuOEpb29Cmi1Y07k6gi+24a5eUc6nGWcqn9PCWSEr0mWNn0vG6etYcXs
sZfzyfZTb8nkz4rGabkwEaIlO2xLZMQJIC4tuks6jOlc7nE+W/liOUesSQoOyMi+JntEIyP2fXSd
cJW/l8bs2AfgDRiUJo598X8HmetJo2Jq9HxcZv7SA9zdHeJlN3PPa70T9D2GkhuF2mW7HESMxoxK
2SDxAuhikEyj0g4cLK0MDWmpwAHKWSbOX1o40bYoUdAR4jq9tXrMKRAaX+war1QNSiyJoTG7ZVDG
B4AGreIAZhK5M1mOMcDG1pK64h74CWb+4EJjhHsx0VcycqmHduhM4df7j3G3KIa0NPRWevuh89S4
yxUNJyGuEkTpDj6ETYecUXZy1OhtdnTwg78bkiZPXx4p4xUrwTaO4WIP6PUwq0XGyBuNwvOGjdC1
yTfhP1miDrgZsyeqEFSw0Oy69ftITgyXuqBMqrjtJt71l8+W0Ua2MF4PJwSEvykZ74+rNZMO1DhP
IwJy91e42Lse8MoI2pNg1Wi58nHep4qYwMzsyiGc9WXuwdcli6uxfj49UeBIiV3wpqnjJR3A5xy3
/iu2/U+bx5P+Xjz1NEn16kBOufrDqLpQuol/ED1909kdRXXBKE1FTwMm4sNev2J9jgdKpbnOUNmi
uWzjRjgwoFRdog6Mq8KNIEYdS1CeWjvIFWVCLbghFFsHBbJaSua5gYQ7sszdyVuRX9El84RYDhaF
k/tX8AyqlFs1sWhQmsb+i1j0dsmpTku5twy9h7B0ETcwxv6J3zJxAPF77NYn4JvVAS3nISqu5duA
MmDaTIL2Su22w1GdUMGfs5JB4H8qJjFKKHRclHMIWUtdErMj6IFCcPlG1Bzi5DqWgYm/GlL6eHve
ZbjBFvdmiA5sb80nwx3Tou5eD3UHJaKfukMApYN8h52MkUKZp8lH1Nntv+jEVjbr3xbrEDd4ZiBN
BVg+UcnP/keUyGQcRzt6mkyXcu5YQstAHTytwZO4gtNcyumU68b8KTIsoIJBPd+0eWq7POzZzyCN
HE6Qrm3Uvz+LYwsKQ6ItXiD9IPxBJMZnOOneLgJepa/brXKtWuAZsnmAGOH4U6Gg1H/uHb1GZ5lH
jZiSpCLScBUmNieZ4rQBsBF8411HkvZSdmtbR+4HqEe60HvWWp0GsrNpF7xwES6PvlMBHH6Cy1OU
nbb1pGh3yJF0bDaI/qLbb/XLFvI0uaomUcBrw9rjZK+hZw9/I84zrGoSJ+TXGi+oFvCfLxn0xrbS
OTOyFGIDRzq5Ul0shrcoDd/YHPBSJXwTKAfxlT0FlHmbI4QNnDDuGcs9WfmCf5CGkPvPl9Sbb95/
TR+0fq1gv5gyU56JwsmSQwAbJbKHl8cths1r8Sp7zhs4pi8wpEtEhpr8/G+5uxU7GK1w/wEuIunm
40bCiQX5ujSykaxsz8jEGRcF/46LprZCmMKge2P2kvOrtjO93Ul+XyjtHTnYO7O4M7tg/grrZ0+B
h8szVFMBN4WiWSjFVOTD+2D4LBnrLGh8/O+5AFZnOzdhWlMb4kzn2XjIWoMJ5UWUe82A4NAKnjD0
vlQdXE6kGnOu6L5cwl9O8IkHrA3LlIb4/yRmDT61LRwafmxqldlSCFpPlx0seIbkplxPRRk4BnP/
DjoMwALEgGBQ22Ppg1qPaJofkhiozhJjtbsECWK6rJX+xjtygTqwYe8fWsEImf3sdP2f2a0LYRe1
d3PBKxtcvgFP1zmcxV9mcthm+IRFoNeK2YGf7+iBcgkDsRu0+g4SVlHo/+X/VroZVfND8GLOhTJi
NYyNRE/tJIIhpNwGyl+aneUDb3HOJJp0Evfbm1U+iDgvyJMRxSM/XCFD3QnmmXtxYdFhVdktQWRx
9usWNHrbhmYqWo042crhR8q5MVyJU005ilk6arWaQuYQnzJR3xD7pBJzrk2v7friiB1iA7xLHiYj
WTbPp3NJ+ww2yp0ixVy2LLxv14LMLpRNE187Bie5yQ48iT7kaMfkHcj/dKtUwCoYW4MXMOn7bt6n
EStikAxDWUonIy6ZXiLogwOs9u8iuhk6TcpDkbFE+tftXnNjhdU16XfcDbCOEADu8DHR4zBLUmct
vDIBgVx7440CYpk0YYO33UKMkaKPv6hVNU3fsTL1LrQqu13TFdVtxeCkjcNcTWDEvnQfmZaHKWKz
dOajFebvXV7G69leAL+BuIskMRIsgVyPMOL6cceCJGownUiBOF/K6AP8JPIv9bVXasDFH2/W9Gv/
8o3D2NbVdX5fupXnAL5GB29wS4uFnL1WhhCSU4ppv0EyBlPUI6+TwxYBFHs1p9JTRJPhbxi4ayHe
Qcc0aapmQvFmycMLWBQMISTb+/LCc5+roCOI6IT2OAPCTXprbkcbbFFV8gKj4EKV9Vx5hDe0phhy
YgldHpAtYMyIoY8LxR1CzuzDT4uv6ySe3poLr+81jSEkbuf7DVCmw4ePPfN8+b3nqisSANF2uPAx
nrRNy4paEuNw3C6plHYtXQ12Yv0+ELYBgttiC9EEgbzRfZxyXIY81MXy2l5OIPe6a4Gh2XTn8wl5
diXxi68V88ueuspC/pRJO3ivpRiW4Bm2a2V01qA3rpCQ6hTmRa7zfud45poP3sqxGLDo2VfN/VWO
3+PqDoa7t9qdUAe1DBFO9nuaYVSpIl6qy3d2BOeS/PE+RadrZ5COT7p5J93vRW7Aij7yDmrIC2Co
U5sGlRvtycyCZKBj+Jec8gpFlwhqzEyNtOk1EWrMopp6JyIP6wSAI5uaG3ZIDytTRa5xLXWOD+bO
dG9Fopw6+qA3zINDPkU6vZwIyipYX/CitM5menUtFkwCj9XXrDqo9bTynbH08lyVW2g+KZA6upkr
GNiqSvBSXvFWJgj1g049NEUsVnicNYTZUIWS8X1r1CbwxT1CussyQgcqIQ1E9niu+JmphVMkE7Ss
x626SnL7RhSIZWvXvNcwEEHphUauHZUorMs0OJ5mod/sDT0knMk5vm+cJEqWyuOUNRUolLu7V2aw
HOUVt/k2DZhuZWvqAXlUtAjEwzJm77i2LXPcP4qvJjHw6o4AcQCPOnpVfz1CSFDcT6f2lu1UYEoS
ONReEB2li5+WS1X3+LH+4RGB+D/eI6RY57ADFtpwLvoHfQSQYYn2CryYEj4vy20OqnviM4ibJIGF
OtlWgBOlKU6fWiSJD9XIh9buCtUun1B/pDU1kJbrwaTQBidQQoWq9JcJMSp5jpIjr/2jp4k/Qb53
waXgPGpI/B36XI+jdK9k+/QGTPhzAoZhKdvg8mMntYJzuIM48IOvVBGbffhZxVwXsh2PXeKtZQXo
ukMMf2DGsZQ1dvFfNSKfccdmbSUBtgZtW2h7LQJmQKHES7z3/vCikAenRcpbdrG+3EoZvJtHygcc
ILdAvICKLbi/N4u2BxTVld4XVpN+hmlTsHr8eAY4aqAYgLe6/hyNiUAXdLw9SjRWSBVXmbwidzwG
993mCKYsHlR3makFAdSsLf/SQhHw5a+B29tpkyxtffPcgzT+QBhrCpefIK06sgsIApecNgn69oW5
b9uR4ipt4GUFPy9j6a+9qm4U7wf9t2EPPkP4plW9sOJmKBzUBQUgRQN3yksHs70bBYMz8hKpyZQ6
iw+nwfo8iVQQks807rjkpb1OtP1i6je70YFavqWEV0yhL9aPbZnh7JaZc9sciKYDwT1pW98UNbRF
I0bm5/qyB7TyvJqSTJTw0cRj0S07QME1zGK4bG8rDFYf0JAY9LQFx/OBR5za92PEZpLGjS7XAdVC
EcF3OrsPT1nJCdz+MZ+mZ0awHmlZzvIqy3H1uP9ahlT+0WoyjLI7gpCz5ZEOSlFDDPlPkRCXBMyz
RXlHDeELEjn8nXnWrqlFRgwX7GTHy+YpgOatxK17cFcBwPwiAEE5dZUP4vKMdLUNg10oH0rnb9eC
/f5NjsMTsnULlYwcxO9zRuHmEIncJ/QbIudXBJbuE3MGMgFrKwLEpZhdb5/85uTlaLZbKkF5np8y
+ZEJGf29h+5769LqKaqjyfJs7Ubhi02ejfkX0X637x7wnNXvZqHS69g/G7Hn5zJGWOIirTEWtthU
e5YvwDL1koYDccKQGUJAIcEZdj9F7O2T6zlc6cWM36pwottDzVTVnxd46pJUhqgJazJDdb6feILS
YWQfEpyUKNmr4DZONgVbLzK2ai4FZewFpzaCsIuZ7hQKL28GpI0e9jti6kELNUkym6mIwwjhfw2u
AYWk0Gb/Fiikxr0lRecVUOxJy2xDKKDvxeF6Usqen2PR1UhvqTkJ9xrg98gvmHodMPelRlNKpfrE
wkliR/pnEWSZIv3SWHQHUrWdYwF7se+d7ZchgAGLbpWtGYSYIjGFqU1lq3UfibgZHYQPa0q6g9KQ
4S7NTqOdV3cHX2beoZ9zzTDo8S08pFNthREWxEyQ8/aVprp52uIG4IKjFywOc4RggSNV4Tz7n013
/g/rQQPX/hP1P4ZKTDBWS3eaYYMVF7YYmehkiscNuZLz/2Ul1RwmGrSSDxarM0znYVuMG4DrW266
TwQSauF8OO9tbGgHwG8ApUqe7EdzKQVh6gEsQV9g
`protect end_protected
