`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
NBEaMs3qf2vRCt9CFTGP57HVPZ3VcVCIDCMjXDvQFwX/EmPbB88zO7+RCFEibKSnL6iB1S9uRUV8
6fkjPweJ8A==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
kTW8HzSs+TK59Udtx2nT0jkDmTeoDqv9kR7OeIAboT8M9FgxuRhFueLgbroU3svS1TD46xwgjO67
gjud5nWulR/xxnqkG5XjPbXC9RS0FxG90EL87XW+/vq+VOMmh5Qm7Th6oA6IfcClHONPSSuNz5ez
EjyfMffr2SJtq38ZakE=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
uQ9YYSMvQJDTKZv52gFvzo+bXLpj8FsCE7/Zl15EjVcMpzrwh1dR+fDhWdLXHoFmtEPYtHUdVU2T
7cG9Jz0GHq3MfhRFJ93/MRu06Y/L76cEgKJ+Ojvibjq8RbviK3gxA6ijnZ7LW1voPiUFPWK/QERz
U+lI9GDjYIRepWe4IkU=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JfyN7w4w1mYxh/nQyD+Jk1BAD1YQkJDkWsj37Gnhut+k++yBH/pu3yzGsEfzw627nLpYj44BqrBl
AXv3ce5dfl/J/yqcmKdItSJAPip11eXnFDR0vPHZ6z2Vd8rPI5l39rENGQLuU+QWlNoSMPH1f92X
wYGKLJ8gPjFgwPmosASaiG5JMxsqwQuXH6ONZRK8zp1tQEFGv9ZfVyVMfekvuQJ8+z7Sra6BQjOr
i5MJ+cwyqOwv+rkZl2msvfENIl54Xxowc0q+cAKlVH/SyPntvhalXdVNHvBEu9dRAk4dPnqjlrTe
B5Aq5+m96pfONqv8kPqwgyfUNG6EkktCVigYUg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iQHmyIgxxlgJ32N2NAuClrJcxSP/FFuyNYxcCJHEZrwYdlX6KwZ8sUoJ/UxAPPzxyyiUvuVsE+Gp
a042I5zfBo1vSmsLsShW7r49tWICzld4PXwCm3rW7hkPwcGa9dId7xg1yl3ub0srhvb8pcBhli/a
1bxfVh5blwx3Vx32jWOm6fMWKpKBQawvb+RsmX+hMCsw4IE2lRuSwS00FsoMxkR95wvcviObCgQa
KrN3ili2Xr8IpDiZW5yiP6R8npYI8La2+z2kQh0jFrAT0W0SawlE3rB/GCkxZ8KLST3/CNLW5p3T
6VSbCP/kVOJ3Lqc6V3f5OJBrZ2qJAosHKzjUdg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QZOleoOE/U3kW4+Rb9J1mBPE3ap7T5ZkRXRYHDEf14UtoZXkuILnTdXG2hYCNYR0tM7b6Scfnyvm
MG/YovfRxOqawHhIk+BJ6+QyIsS9lgOdsOzSAweY9l81dyrkTgZ4UG+xzydnWVLvZKrH+Vr7jln9
VWgNHmtYuaDMCgXx2CaYRfdyX4g0isygcG2ujr1iyneSg0TREZSvjMUpzK3Od6BONp9hBynnLakX
Kc/AtT8V986EKKGglNTGNS77Xp2/p6u0MPUpWnPJnPYBAbn4TzFgl8puOZyHgHXMivYWvHJJ1uY8
cME7QLv+iwnVVV9BLtmO/rSOhsc6uN/Mkc5RvA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20128)
`protect data_block
Ov8OnsmDbSus8ONAYOdLtSgKn93idMS/ZJWCRSoQWLOKU1ZVZnEI9Z/s/hPXZ5XaWXEFwy6PNXV+
eLz5dTViDkPSG2WktvvBOiHpB/lThc+3Aly57HySsZx/TBzdwihcLogRYZCjCLTNLn6M0V/dQKzn
BCqKycQH1CjFnaetT2xXHpMz7Iejny2bwPbgmVh2omJCExIgj7C5VP38FhhiZAYvK23jioczO0/t
hTrVPx1dXEzIFXSzPxoOtwQQtmQctobUHPciBWUF4IDJKsIHTy9XPPawEIfw4l9Wb2npW8Qz0fA1
QrmuWXwUj2HJ9f5nueOd6KqOzWaGz4zUUDyLMn1TovHXcOfB/W5gmkx5UFq6soydh9ERM59ACxHD
/64jm7fOkNUXOI2IKbbBX1IjrNeOIpqOJNqIkkEB7LgnFXlV/kv8hO67MxlDnov1UukCGNog9pD+
vwBAZILj6w//43N2/wZ0YsNzV5vwtVxsgWC1ruk2r3hVHARyQzch/YqgeiIRyZmk2xrtGkd7LcWb
0lQAf3VLpnze+qLx3Fyq97MfLIqK4q6gQlnjyuEkIUp/lg459e25c3pFfrJ5SCcIQbPeEDWzr07P
utK3EJ7Ee95E2A42OGsyQvgNBSBPi3KpCFCl98baDTbzUjfPGHuVnZUmg9zRvZyWzXdvhwVvSYMQ
+kwJugWKANUpCKvLezu1CJDnj155zwYqSEx7s9zMv6Pt4DCwJvlneOfwzCw+P1VVA181ZaRNl8Sm
kjoDb27ln899wvBi9YGqliVCyiMJgIEzDJ2x+//qSgzY8orHMLzTeC3+RwqtlsEVRQyJ25Hbt2On
oMsMQ7I82OyhmauD+pLy62MlaeBiDYIlXtF53HzpRBy3R51UBrCALPTnxB0+Xee74zlyttSEeHTp
AJ+pWDVeIcfmux9t9Iupm3rE3AzyHBkKr81LccslzHL69s7RBstgjTRzqoLkHMVR01YPbJ7FwjOM
g/bpZVdF4WWy39Y/jBXTANFyQWDoZJd6tVRjNITzWJaGmhOx177pnk39i8g4n6bUp9zYXG+nISvi
75N0qdmqr4kAnHAgCN6p8bstBKt0iA83XAP8Yp5z9WgqTBR/je4dLMRdYooXR9bS42iBdWLFHtMS
xppDpNyaq01v9m9px3iYOGlXoDkc03CqJ21fPIkQDrN1yMK55sgWZEvpsLNyS0p2nvcNq7ojepNW
dyBDpyRGnrPitKEybKUzr4krbyS5+8TfMygRNlv0auR3pkkx6OAYcvCwuiTw1mXoseaLLxjbWwuz
GUu8PL9IRqKCrL8si5Wp7Z0X4OvTD6VsmRaFu066AG8Wx88N4jK/od2+mL5do8S7rxCK52kvlwUl
dxZSGvqayfjq/Eafsl7t6rRKzmbf4VrI+pUOEvguVwoRaNHBUM6l+ssvdvSLAf7RE4DJ4Pj5BvJv
osbb62jgsg0bJIvfe/AgfJSO1tpBDCPiLSbIRc6LJ+IDWqaKQOc5rZfGWYdRndDHAlV/WLE5vlfh
8yzGZzZy3S/RyjKmbsvyk0FSB1kAdfU6RhPKlR3e+TCsUZG2ndzjiB5jP12KpPCzagxRYLbxkPJv
+ZDetFHecd17OcvYjHw8rlFMJ2bBi307BNnFcNL5IPyf+nFw4U4oKuUpMF956T0M7u6P+oj+nJYF
djFjfPAjybBLE0Xse4OBtNybLFRvKcBdpGpF4+3AE0+OEei6/NldVZuYuXdHw6eSCafRdEskb/yg
f93s/XD7NxGhyENEGzxWFnnTBZNuhOvB5vOhIvEOF4C2abD+FPzATDSzoSVpZ+k9lM+OJL5dXV1I
BNIPcf0Dilws0NzTgoWHUnDCLpcSVJKiMn30qVfwxArv2W0XvNmT6HQIENePhhWAXpDK46I2/3y5
juLqEEYE0YHFXxqH9dKEWC6UAJGe1Z22vLkJy7u0VrM7yYZmv23PlBMxLEgVp0Kd96rtx5IpI5My
Vg7wcwiWmVwRtTCIcxNdovKd+vwUwzYBxm4Z7nRiK0naHOebIJnWMsq68wRKjIvlYTiZ973JCQZz
xjzE+eT+o9nAgHvZolW7lFUB8mYAGG0jkbmNMvQnLA6IOcbcUQTJ6rsMUab8iTF6eCBg+g6ygKqD
w/uspVYACLWoDvrsS2wCNd3/GMnL0wIIb2zS2V9OyhxkWqc2BepKzrVwRBcUr7zrSJN2j7Cht/6m
QehV9cRhmUIaPJUjpP7fj+uIVIbv4ckX4Y7bfPniX7GiZMk7F5l10wyxY4bNMt2GyG2T/FO8FDrV
mqw+sfn5PkLeEgL72tzVifRYeo305He8Skdp0sWW46s1ZaInjQciOfIstjgaTWT76RZp2FTgMzm0
vHtTJBXIuEb3qc4SlQkIMrrL246IAZnj991Y/IS6KUUtltzI2WdQlgaVgFE9Kg2QE7RAGYmT4VjX
mE+meKQAaIqPo63aN9JXKZF7M/dhimAnHN5RDYkJfHR8qCoUFapVniAXrh77RNRfZbWQ7nTzuqxW
9tmICCRyhMoU1Ydzx5rh+hT5simyUTsJ0Rs7dHGZ93fvuafSkE25wch1Xn8G5MAOI/X6LxKV8ByH
503YCEULlr8xTT17opGVgpEXYWb3tcvW7I/frv4/rfT8BhhpvFPdoQGduslPLGkM4/Gcl6Ft4ldk
34v42qXOgcIKh+sW0WYTk8MYHfQ0eXS3L16RvRir7s3a7UBl1v6Tahwu/+qYvDJ/terGnRfn4iNl
ASvfbRWytyGfPUwxeC/vT4j+16uPsCWk7OWNwHfDdQJWRqQvOHNEMqmX0j8NWABKSP+/r5a7kZeM
nhKwlbBt2t0MB837YhRBpTTHgBN0/ovQ35hXAn/SfJ7OP/tLc2FUioiBFVOQYPNWFExlYzPKLUgV
DmOWjSL8bqUW502a+N0sJegJHzULoAoQmlRtxZal0uLiUyOd7ePPR8LVNZcUg50QHGLFkeymlkTG
jiB2qZC9P/W9/s/PgN1rhEzlwX9pYE+kZ3xUXZtmGLGhhbsGzXWmy2OjPA2xC96bt7Xg96A3VU2u
H6pv/plxf4PwoemTneEcRO3sTh7O+w5v0t7kquEZHs9SRsxPU7YQit6BfKt9WXfG6JVmUvk6oKiy
G+RnOlMf6dUV/VyMvuW+6gjHl0dt05w4hQhSaqVafvuryg9EkxWbIYLP7QciF2akx1sdJlNM0rUj
gQTHzC+1Y7Yt8gnFVzvHEAlnLWKIie5YC06aH1gVerYEQMd9n9uTTL4xpluzgSA+hKHBWAjhJLuF
lPE6I/UULchiznwmYanWqyL3qkhyv+8+q9o67RyMWDFI6yG99FkLLQogqplllbZveH812TB27bh6
Je0A4au1eyDfLfx5JxWpDVFraJcuAv9bX7A+coekEvGrXXDL3HMnrqedV+FBoK5yZIOh2YRxWyPQ
VmzH+C+QHcmxUsafu27uN5rRO475Uph036Gq6nUCx8DThJQqG/zhajH29pOyN+XxKBb7DLVNXabU
uIL7eKD8pOgM9uPtu4sE8SrMDHLUEl1rUKBlTY5SxmcMdMFkqxsxzWXKN7toTAcPBjkcMpEDBG2b
Cg1li4rtx+/3nVpcaS1wbMa766RD/O6W9LtYTPFu81eLFGLkOwQ2WTCdi3DrwlRx/I5gQbbVkcWO
ktDvdn8bnUOW3+BUkCEdVkxYOts3LYOJDFX5c3vL9uL8UbuYL+dy/g5aLnrKxei7ryll3NxmVz4F
yAwlbdSCmdxMZhl6AcjmzBZ6r4PeqgMwaqyK0O//qCp/JpOBq/5ssGpQzlEBxHUVBVljrBGEUcku
B/HpCWlF327p14FgRL7azWRx4ka879733OMdT1Zf7uVEtfg1uE90eJ/TH6HzM0Gqgr1PH8QuEQlx
5cdCKWl7Ih23r15raHXF6fi8alux3lPzml9Uc2HVWYJvgzSlR9rzeFNjpo32zPXvN4cRHF5S5qoy
z98CpbKL9oiMqPxJyuKb25Ywb9pfoTbqMyfhlORfLrdaGZdQd/8uL7UGmKbegqZyDpUtY5e3TNiI
Y1BTySB9hWaWEaiDDun5AVJQ2aQnER9rh/+DA4N34xbybBfZiDkiGiit4FATYl7+SxvJWTdJ+URS
/zam8QyHFjJ6JL9UvMnpfE7N5J1l8li51TDok9Z3bEOXfZF94ZaA7bvhFlvUIANLKw30WF2Rauna
ztCi4QJdPaw84PtJx4RY8rWJILv5D+e0ExGuwB81fIR5A4nnQooXuA/s/6MxfNhY9j6vWuczuWhC
chhlbGRsTleFbP4e6TkSbZ4uUk2S2J1NaaibkKLMpkwLF7swyzEqzk7RDDZJuAkYQaGeTb2ooF1s
+junIUrXZjFHpQ3olWqZXosX9ctBjtt1oQoWkrHvHwjuf73Z1c3e6Liv3BrY3jcpUCKsRMrTilAx
uh1+LDiWfNHaSlc7RJFGLBtHnSV8OQJ2CxQ1Fd6aqrw035ntOdP8CpxwNLTKzE3S0zfAgEex/w88
eKPSotOH2nTiS4B3BeT4hsg5oRWvMeY595dFuVVYNX+lMHPjDXcF8wZmi+p87XzsnkeG136V1ojy
cFgBVmBIkBvzhdHxvYJcvLD7ZyJhJu9D/qXDnSdfXIT+nHeA43H9ve+bY1GGOQCRDJKHXf0cKgHx
E+vZ6ECETiw42JOF0LWeWens1XaSsDSZWAGSiSvCRSbFjIBWr5vTZHekfBed/vKBD6h5F03BwOER
f1ynvKOmxoESrya/qHQSV1nFow5hxur3ThpvfcHJTBKtbyr83EcTl7WNBjTfKGt7zDNyZcBBHuUt
1uRteZPh2kZQ2WVre6J7a3bRtIMJmGNYrMqYwwO2N7BPO2iwlw5CWO5QV2ZN6CqDAyaQ1tbq2lZc
MZVf7LzBU6RJwGZfLuhdnBpY2mbJKPP8mYoooAG12ctrg+NaGfHzO09YhNVHU5djFfJhd/jjzG5h
QR4gzeZA4vLmZYSsBKmL195cRwYvJq0Wkg9ZqGwjOX2jdkVCyqv4vV6wyoPRO1qATmvwuNITfK6W
6aGIXGgdCgAsdhDsf6xKOnDxTYPJO8CJBxf8XbE7w4qN/+ks404Ui5ikTqlN5Qo+bSrm8aWCpEVz
CqrOoRJI/CowEeamxlVhg7UIKKCEYJU01Z7gU5DwiZzt8WhdQ7dK2pEkO0BgrmRSzTyGDtnjRDCp
nVghid6X1azCnNwr1oCwLkZCIKrG50U9XARScd1CvdyQ278edYWJ/lZKhVTRC3sckewvpER1gcvR
3F5ULf64FqcktMwx7jbw0IZvX0FserAyvVSyLjQkiOFoUOaeEmhcNdP6VGpWg4Pmx+hc2Zg8j1Lt
jupsJvOPxi5kfM2molNq3UKm5t10Fp2SND1yybX7vnhjdaE+95aePSMHCOtCx0Ooos5nRYn3dcc1
kji/WB0SqK14zkzgODOAVJzDVp9l1UaG9yQhREzYt9SlEBN5En4wxUX/Ik6KFC0WosnZw9lf1J1T
8JNgpXk2wX05Q5twTnHJfnNAvkh0L5wEpWEvGd/3x7CY3oKxxgSSteeiWnP/U+6U3anRuOyvqx4A
MW83OMEmGyC0KQxe6MYxOv20N4KGLdhvAdXPzrZAJtP7PKuP80jSOg0Xy81Z4VGfXH9idUr+HBZl
mfXjfoObFWB3Sr67IC5X1ScMNUSshcbdyzt1Miglu5IUxrrWG6xg78NpMB4QL6fs44xTnCh3jSX1
AO1EufuGeXpOxy3T2bbHVbDOY74YRYW7tagpmhbKYZgBq5+FAhY22rXZ2kwax3c+mxSN+rlUHumI
hJT7LmNdcQE9AJBHrU8f6r7nBY5PWQx1tD5eJ7reEh0YyExPPlI5MzTmhbh9t36eeMhnHsclzpba
8JGam/wdaQ1yPBmR0Tz1FkhO6R9k0Gh5X3L9oSrZjJtuWV7+5j3Dx6+p9FZECVxFT9hJyEmVqgGk
H5JojpR5fqbd1hEFG7dnMbLrv45la1f0LDP5cmE4fHmfTaLcosmyMgrlPg3EzAuymJtxsz45uGOs
k1hC0PKXFFbKhaXes7ERlW2qRcWs7X/BiNIPcZqiA7E7ejms6rIAsZP057GaBme6goaH13HupEZu
lkjpckqMVJGvhoNLYxJ3iYxeTOtxtDkoI3IJeQ56sP+6gMxUkhJKt0GkjNAsbTE++VbZgiQy1y0S
1qknh1xgqqT99727skbcIH//MxnNTniQC6BJ7AaU+7SkYW49JE5VSzpyHMDfZZfPFlY1JNUyKOFV
xLnX7/e4NS0Kw2kzgd9+ZWsF0qXT1guuG7nci6srTwuGuCBaJR1ReOFkIftupXx4SIQXcY1vkgud
g2oieGHLOVkqc41LhuUQXNvA7cpax7/VtQKswevPtnMzqFXB1ve3ltZGrBe7kAHhrGvJU3kWu2YD
S8jE8UnbYYn4ZuH5Bpg7nFBZg6+hv1XJQ46rfX36KNPy5iBElF1oTXokK095X1gfJXrm5uXfPch/
I2yDN6OllQI6KfW+LA1eLJN1kQ1ZkfhkXC18XNkpQbiZoYOgNFP+eLFhGvblJOoF7RRvWAimt+xg
6XWIWeCfSunx0OegZBuHGh5wn4FWXSg4k7rpj3NwXbzWUQf6UjPDapLCmbB0NsoZhML2Dgd5xwuW
DnQuqWOXeVNB/WxbFtKoBbaDsuOxqi+dQAKQDc7IaH+1hshlGSmBUFyCdl6HGjpwp+r0k5XM9hoS
icqsMNsv0TLz92fPrdc7Y0YFJL71IYUta6eR2GUzc8bFmStFt7dWuhp4m5PX3i6e7ZRkGgjNCuV9
7QJlxGH5E8S7Yh7XvXtJjX9tHBQFM9C1T25wli0reKYA4hCYHI7JncpqzZcv4HO/ktRmm3ixE9/j
k95KcNWyQvxAv12OsOHkpkW/UoLeXBi7KlvQpnFmpguWzklO/6C6oCePE2/mlhxaM5grI6ZWOKyN
o9GSgQdB29hYf83gKzewhCTxBwMzKYE5urKH6XUsu0Snkh6MVkAb44hCxUXDREnDjgwqB9TBDBaf
ehYzXcFGBZ7fnoFNrli2viDdz3NgehZC6k6yXLyTBdJldhNjD9yarSnXvs4yDeFo5OzSCW9CKOyx
4hKZ6sXsSrdf1UQ1LbxcktVoEKP0OQHn3Pb0dvGuEE7dsKT/c2PqgiF+LPT5ZpUx8Cwf+ws1cX7c
TXPeNj4Rt7HqP7oC8MYIh2eL5MPZQVuas0YK3twpNGdYbixFeT/x7NuW4xW/L3O/o8IuppLSWY3B
F/85mrcti7NHOt2Lg1KZyy/P4Ex8hrCdlQkgcY2t8soh8YX7nblxwmf2zh6b5oJoJ+WPrEbcEkdQ
UpPtF3OyIscG33dwMXIV5HBhHb3YKDE29B12EjDCa/4wdkB6dY6BHYVsY5fOukrY24dZK5yyIvwV
OWoe51OAH2N4svX2OOWq+kHmAGpufAu3ugJtFwOMRjdApRAoFBAxVah4rcsGN2TsuMr899/hrqnp
P2qHRRYtMMLxYNO+LRTp+EqZA3r5C5dUuFkOePHCdcINQb7UHk3hzhE6qjKcqGusSsh8XMAWuPyA
WvJzJzCZaDBhUYmrGZZLLrJNeXoMO/CfRzbMsPQ46q1USn1fnxYeIiT1JcIYKw94JZZMvZn0rb2E
zTyHQ+/MBKflxDuyd3eqRK/u/rtg9O+9e6EhsfQp+8HVYvglW8pfsStFWnpNNULLp6L0iOZzKrsX
AculXI0WiU6/yxVK39cwMjMNbdfgZoM77F4pznASrkHNcCkkQ2r9/ilCQtGFFB9uNRhqxU9ZeFQC
/RmTC7Ddh1pzlemUBftcEGF3W+YwVeYZ1c4/qwjTH6ejwCF/SuqXZ5HxNsAKaiIfkU5soJ/0a150
+vc/SnXSa6UPZ+9PPh8w1XUHcrwayEyFQrxNWVR13zdiXq5bxSdGvGW7NZZnyt28iQzk6P4HfqLp
BxNmpYtCx6M+psZThekDvNvk5JIex82TXhNePYFzKcpL1cJd32CR+0dWQrji4fqLvFOxLxUZ6PMV
gNpdPgaprWw4x+7hUhixoj+qjucsABZ2I1lzoPvBOa/Omb20Xr4NpXCgc7/pUXDGfBBJE0fcLer6
BFsGFxrQuSiNdkPM//vuAHM7tFvSrEjpc2UsyL5tHWrau3A8eCLH5lEEB9psJ2x9Psx3PXgZt3c7
GOBDI5Bfrh32UXwTqov7EfkcdSFOWkcOyScQS7LQMNAvw40faWxlu4u1B6ORanVtXscSH+4RgLal
A3cVaVUTyfk3JMtsAtQGJb09BaZHxIohvrowV3TyzwjKYheV+wDugPZH5zmAC4Ss3c4Shp/zHtlk
63fnd2VdJVmfoSaY+SFBBapb5uMdJX+GJ0QHahGKncipCM2kg58vkMJyTPoQgB3UFmxRCos1/0tR
FRwPqMyf5YOBUQ7YyIBfP/hatwpP9r2YPw43ZN4OJu6JAQEiolZBa0NwTjtsWvRkAyxduyfhviPT
lpsRofXFQc2bmwKG7bryxvFPXd4jiOKkiFe0ZntPMucOKR2tWFmJfX8gOPDzxvLJQhWgzCDXOXrm
sd6lR26Gzqhrj7ucEdrzMpsnh27jmwQYXKNpVDMjoDIyFQeyJPpPZB7dXkf2SnAyH5rP0F3vfhBC
IOA76baKODaHd5J8oeira6SCVTvQbNZK/TKZshAlWl1yACr712G6hkv6K+Xc/U/YT8OhL8WXW0vA
sikLBLccpwz67bYURI6BN8d3M8C/Vlrxt+Gm5OeQKMG8phiqDdeXUZVyB89aKM5jusTvxUMkLa+W
sqJs9C+GdORvUKea8WUMgpGExYFjlVyI9/hLe0egbo1fbbsehOAx+TPWODxUKEbOpvDOGfFBv24D
+PzAGvYKLgo33xnMMLHqe62tkhIQmL9dYoZGaT6z1zeWXLIScMyvsXmVcVd/YU/egSbjnWMttLoC
JW3gKANCkLAAALUiERvahwkqHD5ttg2rPd+pKsZe9AWHE4wu9crkdF7jEfGt3wmCjwQH5wziau5L
XnDMA4B5N0q9WyIRuyOz8qw/gB4iK6flY7Hnsuc+CYhkuzroDm6cSo4Zfju3K0ql8P0kWVfhb40m
VIWAlYI553+hxIqYY8PI7Cf6ofNVPUZAI6jfLM/XHbzHdnCFozK8WErEKJ6soXA55mNHWMcicrEO
DLGd2n/N/STDQocSiuoim/unctqDpoFnvpGkodN8OPxsiRIFaROkz26WKo96748LXfX3TsYu5H2J
STTqLwj8pJwMIJxMEnSSqa3AmGw9iTv4oIec+dAa2lhtPSsTKNIct+vU/xEWRRFR40604Vk4ngUD
lSNJeEsjuCak1yo/oJDZ2KtgQ6RgYsQR6OVXfxbxk7YCq728AQTKSLdQcr3rzZS+6Z+jP04Yofh1
JwGqYlOUv7DPNR6O/G8gCcqTotrQUfGEMrJKkumZCMGIGCD056ZA9aCRL6hT8y4wEEj8bDwrfV53
neJ5CzjRPg+LFEbmvAvSh397noDjeQsWyl9seAj1E58PfZ8CsLbVGEdAJEXq3TQx339RvYesKZLB
i1BCScxmvkttWWacbkZyVr3GM/XVG5/YNZ9aXZDwKpQLaD5e1UTfEVpV+lxQ+oBrc9n7L4f3sB4R
i4dDwoQEVwbex1/krx1lBl4eWFpSXLfQfscLZJhmNj+L5HJEKMv38r0H8HC0KMdiCVIU+Va1fa1a
WSPrWcnWiXE0aEg5qhJkHUqh3YMm0AlgzhdFNfiMGqUKKxYlb7NeeW5R850CTKccminjklEP9OBb
DWEO6y1br4qMS2lQMzv+kvnBC1Rvlk6spdkG/rKBuXUi1zHw4bihbSj4BIMstI1Lqc3jpPPMsLH1
/gOLvHeSQS0lZKop93hVFm4fJPCOAUcujWrAe5ZnW+bbY8AQPyeRTGHqKo5oNBhliWwruJBlx8CH
r+EGPvsdYb9ITkc+k/UAYXAJjLZSDX8csLHRKdTKRdswAyJkwVI6mv8SaXAH543A20wEo71WbMsY
2tjWGfX+Hhdt2Fn5dUkd7s7zaBg/yDLikDmTdTDNMtuvRuKy+LwHqLD9K21pQ1KhiNVO4s/B7FjN
DDDu6mKJ+H3X5tKO8p7Dj5O6fydWK2bWbmuuvb4QDG16YtKSnFlGzmpIRGcYe8upbZjslqlld8Z4
MWsGbwBkGscLwfBd9eBp1S9OBigjZxmPRlITJe4xTQdyEg2aX7gxofA/Ovu4HkfKUpPdVvsEYDd1
XwugovJKEBWh75GNY1AJkHaztz/q4mkY49h9UpGnPsDD4v+rF+ASLwe9W/L/lifz9UsD+M6bM9SQ
y0x5tGSnpgfYTGjgVYnl57LDGOAvkI5eiGnKwbmXWNGXH/EsnrRtZee3p3hae+OA4pUmEWV4qfTF
ziWjqjGVXBinYmo4s+NTpRvucna46OeqMQpWCkUl7nXG+YFELa50c53eb8vk9dYJPcO3ca5UDINY
3hYWlQNbWgfHKpRrH7+P0imGdzGku4xdmVoQjRKhd6P7RjxKTr+rxDZIYbBJ9VY6yy3l0WBcsvOa
u0YUTdZmPk7JoFQ8OOh9yNf76EJ2GgTUlwE/fqxRAzK2eCwWmj07ii6ENk3+3tLOZTqZJbK2Q9Ti
u4mOCavltuwAmCAbqDOJEoLOssiGiiNwIVNMM/BWChEoafn4GXR4JenHkcGsulBa2hC4U6NUs5ao
DBp6q9RmE4bqwnTsjCnXw1Vqs0vX+KTiWbm5Kt1sXP36SwAsRWNGzPSwoySqlbsWgfo0/L5N7oGn
HVAdrOySxREiC5idaH1mgafXBhLbaR+9KITGrhDRiec1N62ETKO39kYrlvfrit84qNCP1Xdlnq7A
FnLila2TbYX8GcjUSApG/eQiBhHdQzNFdlPAOlkuX5T299Dw9gD+ored59qybGx1QGH2ONSazn8+
bOpPfghzMiJzB14AwwP7+ttK++OTeoUkNRHqbu1ZG8Q0rdLl1acnTyJtEFzpOeT1mPSqjoRMiYsP
+GO6KHlsvZFdUc1okMXEptfVy5/VbPSOimF6hxJXkXzPjTfpGkAs6Ul41keddNF7HbSLqkJzRTEg
TwNoAJFN+wjVpjJQaZcm/uBYtWmABlMaW4oewEOLPpLYu8qaq6pDXG6OOVCo/f4otUpRnjriyrii
6VAKzf+0NobF5x45ST72eatAIfsHLg/xZJlMaqmJU/Ub88OZJlhUfblNw9zTW7dD4WSClLZRjxRA
3IvpzE+pfa/sPcMa4dmc/GSYlIbhxI2UGiA8k9mppfSlk6dn5Cnyk8QIU4l9PSJJTMdWctqPABrP
luAxEAltRxIKOMV1n461RMHn+CIVUPy2hpRItfG74X4ue98d4mqEgTMvGvZylmbZkQnV+jSelhz8
C/xYSu8CbogjROwe5fF5T+SOJMy42sJeWPvLKvAxcd3w4LabA5AHAPR2Xs/sLDVux4vLfq2jY8fO
EvPThuPs0oQypphlRuNZsNEo/9xvZ0u+4a47OgGPBnJ/PycCu8KlgjT5IVu5Qz7l9I46JcXsmTcN
DRkDG7aKWBQa+mcyIYAQFPqqkkqrNEFRi31hLzmRfc6+KH9PXvBXkQZHj95+r2jy1oAhAh1pQInI
tCOkYOol6jpEdGCtTKbCrugqUntUeE7wOMvXFmEG6QajfJ0/lYRONiK+kFhWY2axKN4lSgwrWEI7
zai16gbLRTd71ECvvCa3vDm3brWIeZr4MMf7RzuLWy2FxiLBxPPjmVAtT0u+sfxuTcvMD+6hIE+H
L7R+e8M+312N4v6REWD+ZbNd2ech9DNhfuefa2GQEGE/CkyrGv84aYEvLD3neoYADHDf3tbXJLys
qcCFZmf03vHmGFySQEPQnNzej7VxLB9fU1SF5u5Oana3MD7VfWwneWO8BxgdTwrBeuHcVQLADi7I
XfArB4/I1coTnWT51EOu1Y1uERp2YmUGq3Zn/TUB06Xhl6DMhMOJd/011SZu+40+cd+equ6ERROx
b8gDXFhKRgR6vn3Xi7roWwIAVcfoJ0pjpk1Feel1fxBnoLSTD/BlcpYUv3vt9+rzrxjje9UR9XCt
6nijT5sfVUYLnTzDXp67mAUeazY03OsO0/xmBaE9AgXy2wC0aGf55mGmFIAvW8m9i2KETla8gFHJ
+Ei4q1aQunLwrCNT3FCSvZsJImpCgIcNrBoe57TGwKhVidP2VWLIXatrq9DEoUNkj0RChXDMvVwC
FTvJKufgnY3Ye3pkhMgHrXuT0u5xWcXuABbdjscM71s2iSRCiOeY89kN3XPgAfcbEF5xTjMiuqHe
s1cL/Cdz1yfS8GUY+WLjMZmSt0KxX6AYjAQ49AdIa88OA5Edzyuup2zNthwec+J0R2QwD9yCXRd+
tMyrcy0SJijv/HZFl1qqKjx0eheKtF11kcSYgDq7Nvlj6tFCStjZ6gjH0isqPXRpp3z+N3hhoOMA
yMV/bXE8Fsi6oDU/Wr5v7dUU/Ji8mHKap+OZmWwaT+2ZBCfV1ip0PJ3g0dRLAvZBKhqfw1+V7exd
Up1E0hppuaKyxwxexxr+bE5WVx08avNsz4rUA440uDziRw3Sf68P5WoZDz5nMpo/aTrt6pets2ZL
RGhAOtcHxRVibPb98A8IzLiV/b9HfntygySyNbjdxW5KtAp8EFNiCcTaJmzpoYJpoNFqKBaG01EI
XwKbry87bKJ2oykwHc1lZJjUQQ+Na9GDkoBa+ECH0e8xnDYpl/MTmQu47+bUtfDO8vSQCaY6o3Mg
yOS6RWdtcKhe+bLMLQOvxR9Sg/7xXEZ56xrVUyFvx/zMYv5NkW3XbskuNbi/nBNQ6Jnft3utkt1k
nMhL25sVMzlqwLVHj/Wtd0omLKQNdEfUhBC2z41tsYowc0FVKC1YBZsj/ScBGuyPdimoQy5y+k3h
Wn/AIJXJ6nU4siz8mvNA1ZOlZa9PzxyAEh36tqW6giDTFLSRJWYbVpkwfGf/yS4gxafmU7mRqV+R
qxCtSqbEw628jIVxQW/IJuzoMWDr9W4HiqqAWVNIiVTnyumoJukX1SUFFhYMcljY1Kw7JlsRERez
8CI6SAbzZT7lMhR7t2ahC2J6877GP6f73EAK4FKhPw2LcfstKWUEHY1iC4IJNnwSvEQ7fOj9Quif
FpYGYXEQHDkQO+SjGXjJlFSJ02dvMj4Qn72i4tUdW/F5sGFpSIHjJm+ewsR6EdFTlCH4jKwPYvij
u7/uelVwcYnrwb2OPueMlADixre0gsUWxs12r0As5Un9Y92HWmFKMxqj9TOimR31BS4P/EQVqmBP
oVNzkcikFHLuDsgZQ0OSvEo2wJobsypydAjH0T+X52FRZiFfkSG8g1AjwqnOeuAZIGMG1aewy/BB
T1x6XLBpstYNOrXdzFVw0vEX0G9Kbdo1ytiHEnWEZiwpNAVZMgYcg7MFixR/d+FMBuz+fIYSZ+XH
TaKNbSWO2rPWoGtfpcxEoxms7aEeYnAtfuE8fB7UFugiTClMHHwBuzRHXJ/HSYt1b8axMfSNWusU
jlbUDrDmiyZbxl2+40LSN15X77IJyLewQiIjhmo42EF2rbt4UrKKkDB9WLP/nb9r/P2AdO31fkX+
ngHOhnrFTNvBTgKLGnfS4XrPpiVZ8VV67df//Zxx3JfVYT28Zsv1uGOIFl8Zyx+H5RQ8YTYzUp+i
oTsFTzHnHOVb2wZ2rAuRZS0ZT0CctSQG4aH8mHxmGQBwTSAGQJ1zhiDZ6APOVeQeUR+0A6FrUOlZ
OGdat2in0Iqez5e85SCFLcuAJEeZWyfo3s6ityfuufPS+/q6nxEIn+iJv1BHmYmRt+ETKZ/2oYw6
0z5mJbvG6+OllvOKhndK9hxRkdk6w4eMpFln4umED1W91BrVyxJuSu8PDTuJd+QlIZDVMrSu7Yao
jldmBSIJNDpTiHBGQQoN0QBlURhORDZQFQJEgU/vBjIn3DHanJ4xjmQJ/IBGkPbW/n86Yz9mfz1s
SYpiDbEGch+9zw7d0rnSbqxs4eX2Mq4YhMTaji4o0fk8P6X3xDZwJ+RDuG9Wo+Y1/3qTjlxp3OSe
1Dt6+oeTvWd/7KCidX8N3+Oi71dWICRL5iPTrq+R0skr05/2IJxVW/wxzQB4WQRWIgX9mK/FJ7+v
zlRFC/AHV61qUGMOF52Yi5HypNAehpeT3Kdj/uCr3cpbcO9e27bXA4GtZ6j6G8U8YCszkLAl6ho0
qZD523LO6YUUc3yVpZcAKj7LYcpEQav7Q5Z5Tj6l9+HQ1jFg7Z59RZUgUBbWoIiJHWvX2+xNHssR
IIzJPK4bMpIERDVRHarw+6IFkCm6+HFWc3YDWypInoDx8zjdJp6QJTip7cHNOZTmnkJZtdRb7e4g
Zbc3YxdfBIkEHINaRmGAIoKt+PRMhBfGQRpi4sfd1f80KC4BquBLMsk5VPnbn8/5EbPq29R43S0C
MUr5mGLOMHTa+pmPCq8aIcgfqV+bUgOTO27uT7QPcMtfeqYbInkS+1ZslQ3B/fi5oXCgTBQqMHMM
kfPamTM4mNgsdyX7h3JKz632f4x9zj3W5ulyb87BYUFi2QDJcgI55lSjhwjJMqubd3aqGGlSV8L/
NSW3N5OIWzlswLB3eT3RueEdnSke11oud93v5eJY908hnszqlQYrnWKVmVSc5E2ET6VjECNr386V
nYipJo929kLhM+m2AMOE7NFAg4qMl4Gl0qY3GoNN3aZyNqQ+nnQOe9M6QbZnuQH9TvqjmZ1MQbEr
dUlsQrbGlT6DXAi06ism2GL6zF1Ca1Mm2iezgP5AWaKcTg2bxPucSV1Vo3q/W+UilSYGIAjIvWES
ub9uyQYOzpiqWVpziHWRtXpRgepzL1lR8mCX5nApgCjioka54CedgIY1C67ai0B1yziTNJa0ab0w
Xd6aVVrLMlQOviiVvdkP/48W3g23fCCG2TRLpZw03C0wYgfENbR86aeEAYjVtHkCzQF7+Pf81m6K
4XKVNKmNhaLXfZCO5EvMB7NYrC/ltZkTqmO/9ef8eD+1lwRkj618rNuB384ANKwZjuhDnhi+UDI3
7AoZacyCoHK0R4ieMp/3kNSyiEzwg2g/GEMTSEstHfWmqVQtsvafjPWhiybSqLrZ+5vYkWFBcbI6
AbHY1Xyw5zeB3UzjckE3XOmPptDXE+qjvFIaMUMoWa170ykhxX9mBAd2YQsRf2pjfWsBikZcijJT
91WkTyISsc79MwsjOlUTkOt5C6treK+Pmu/3xlalDCODGRPghVONtR4F1uDw0QMEiO7Vi/t8vPOd
yk+k+N+dDyuMazCCzixxJAFWcia9NASH/hjWwCM4f0DMXuUgn7INilJhkBNkq/cI3DPwYWmeXUVY
y06Hrtn6N01boltVihhULTv2ZHosliE2UKDFIkevWmQEDdD9UFTDBs51Gt2rPt0rZI3fatUop0SW
uREcASDguCN8PhbeWcGwFPtqZplFnesYR5Wz/X8tVEyytoyGpPQxkHPWjDy+tdlyYwK1UwL+Xnhg
doxskHCpCEf9iWomvvwEIXk2F30MkoQmmudBCDNr7YcM2LoUnO8kFDR5t9PoTOJo1XZwNH9EdDyN
1+M6Iy7TCfm8nQOaUwXVQN6lIf8zk846MDlC8mvTdpRUETd2vloUqoO3aLdWZnwvPOZKnZBzuzNj
4X1lEN5r8O3hSfWzKOZwRnFk7Ddd4ONqQZOPPBwZ1t506tHnd583qSmZ/fh0Gw9s/hyKNUQdmFp0
gSsa1LmxT/oUCuT5F6kRJGgA8DQCpX695aLdYdLBorfM7GIG2U5CAdxpihtBSYkOjqJCS58V1Wrm
qdNr0ABUNOFZQQW0oSGzppC2pcI2lO9ZkbDSKDp7eJcimPyMf3e92pjGq4pvWljKVThPD7FbUpXt
JHvw3RBaUDEQfFu42jGtWLIu3OP7Na0iuE5XcI4bloydFAPFgH9OpK4utMMAjYvkLVimL83Wyt2Y
gAZpcpZZJIa9FoB5P65mY9rlTkOfr5hbjZXBTTL1Z3NYNel4Ht0EUhPQEHO0jB8uknhvZcwoS8Ac
jbRyoLFNNXYT+3mzDC5BIe3P6o1OCR7h4pVUdz/AxIcAgXV4amb9PU3sk9VD+gnJ0AUN8sVurtgo
aLz2t/LCHuH4LwfIuV8Gym3LuBtO5gnx6g0OG3WCcU2uMDMrx3iIPyaIG+3BxGeDcT2v8I9eXzQ/
w5M8goCOPx/FyzIrlKl1Oi3TSbu1W715zMyxNtiqi/WPWLksT3HE/9ZzgZCHsItUMZi0ncHqQMwX
w96DiOcncqj8uPSPh3HLlEQIyKxI8TsecUA1veKsjHfe8s+Zq0ZuoY3eBE3Jc24oFDrt1bCCyUX9
U+D1r/t5cNkAbEab6WQi/KSJlJI6TcM7+//p9Hm83riMJmnqndcJNY1lffzYx5QZVbQvYgM6OaNa
+iQAPb23yeCFNfbd3KpPUTdVfXSFiaoZLd34NiJw3y5fIn3UytmgDoEod0Ks+qeGZ6MMh5weLjUx
zAAbh5pfj+7TgcS2z/YcwN63es8HVqE2kdQaMoIxo0RhAvw9IU77EX9dyAFB+3EXXN00QUPpY6B9
akgQGN4z81AB6r+Kw6K+ZjzVEyMWZ639QG2ljs+yKne7uk1TdPXnys9ABNa0yXN9S2vAv1qkDKzs
9gpPV5F0whW7GUCPvDmaYhgJYhx+YMGyJQuu+48ZPp3axQzqi/535SAnYE2Q9BLCS6CNvtTooxg+
JwJNzOl+6IgSFkxaGe849csuErY5SsTdiplVzyFGPeNoyPmFQYPxSqBf0clOoamLHEi/Y1kKBFGD
O7fNTxIvLAsXZdqJbIl5taVGd2T0sSWqRmzavZXB5loL5Usp7ShQVGJsn4uQsaQAd3jroVmooXA3
5CeheVBJYLBE0E8+y+Y0N4ePok8dAP073rDPmhjf9naILH+FtvOLrytlFMjr3YSp4lCbez/DWQH3
eOvd7apKjvca5y4pSL2DnqhCkvz3UJTCdRluUgSmDejNbP1KQy4wtSggBGBQf/ht27KrfsfriGK+
M5gudscnVbo3WZRsq6aqUjExY/WmL+1zCK/R74VH8vdsUyeIuxZbMIU6bynnqQjWGlGAsFyWqHTZ
nGoIBTSRDZ3tjTcTX9VnRqqMbEyUU25wf6B7jOfmb6A5pie58CPRTXpxprO+bnHZj1lENNazfqH7
FzwTlV1N6Dxz9QTxb7KKkgizhlC5L5AgyNgTQLIv0RNTAHqn27WSJMVKmnLYw2fWMoHRLX9IKEnl
M4RoMdBI0ipE4r0h1KhRIyLt9FeZyzoq4Egg6XEV2t+uAZ150arkrde6HGx63RGnJiM3hwbnDTb2
MOjQHcWyUU1zkYtgfHvjKcVa+eYLL/LhQKDh4/XbDlBcq5o7ZoRuryokvqHF5s+Ao0sUMon3Gau5
we8rWQJ1OqRNjtcJx99N99Xr35PiG01554rMeZd5rpHVkFygWHVcMQGAcwnVpnjgW1w54okFSFfh
BgX9HQTG1v8802uCwarKrLGCdT/8tMRczN8na5Xc5KiH21FiEGVHVxbMFMhJKavIywLEbFziZDuK
UOwB1KQkySvRPdZ813Ul9gGB/bYK8xV8WEw0zY7ZCtR9u9llERudLo7ONxNj04lQLmwnHLCifszN
lh44pJghEEYNf9mJauTuQy1HRxGbfDE0Vi4aCGexRRhwagFFxZ8J9DPyIXpZMH3GFDy8lFuPrW+Y
EiWSadgwqqhsjD81WUZygsA4XuyRMogoSEhP4mwb+k+yGovAQtoo30vPzvGD1CHjiHdnE34JkxM3
5cvH8/sXerkL4wiCUtQZ+oyhsc4o0Vu9KVaIDYKek30UglYzOQSeSKqhxGLDQoihFln9mrMEf6RY
OrLeK0RbUpJ13jtP4q1X0qts2GCBWwWbnOvLzHVKoaDBQ5LrHwy/IeaEPqT68AhenlVGOX3785w9
3lz8D+40u0CrUzhnJB05ccR9/R810Vml7dBUp2zwTNQTQuKYsvzvgCGChsq8WOJld7D+ZkjRrF+D
bhEsxT9DrIj6yMc9Zqhsjd9AK3v+KW5kikOfA4mYaGSgAh7uCuQn5xGkESBiB8SwFuPp/qoMTwRS
+VWzr2Pc+WdlebOvOxtxxKrgAgXm6aQwUmzNQa0Ywsi/yMGvr6lTQ63mIGhP+7kZJPOyQuyB/Lk9
ljoRtr59rRUWLX2kA8mXwmXuVsGTFQi31XcHwOHMcLgGr4ItpPd9TCmeFdKF30wiF2k4L7u/a/Iu
A0mFFo79EWogygyw1jVxjkjTbihefaKPzoWXjf36sMgm1lW2pqPCPNDoB5rHYYjugDPZ1eZpV8G+
vN/qCuOqSCbPryZ+6g5MyMQrIk5qv7AFESW3k9pm/02lMaknvYhEpwQXudiS4ZzxW5GN3ehKdisw
6yWqiz4NRFnNmb2p0z8su1ln1feYMO/DTxbbDDzPlzl8gJZGknPzvsSviHJr3A+uTeeBDlewnq2k
lVFnY/Z50NRWSavOa+nidp3IqkeaTqbS9GU+0+QZVpGX+vjN9oyfkTCZTTl9iUeI4v6WPo+ptfx1
DgBv34s/Lt4ARz+zPIG4TuNOujBtzl4Kq7jJGyLdgatBSTzvdZfBXgrErTPpehOrOAzZSyGhMr9l
V97aBYNUV3f8Xawu82H5wTUwdA6xpiceOXbhV2z9x/tktfSZUOBq6PzhUQy9l2bHPjMOVwjQvZMc
xWplmDQQF1H+jyEGR/qqv+yDOd1e378U3nhSyurldCcxKeZSIOpAw3RutVbOmjLAwp1+UTTuvagX
XCH9E2NPq5HAQ/sj6Do4TILJG5sYqDntA/7YnWvepE5/4KcLtWpoBBU04vqKAyHHF3hJ+OBZyvsA
ZR114lQu0wKsgkdvUCWeikWGwXxpfF4GSszT/Y1yD+58A6DPrnH5k6839nhORWi+Z/BotRZyhzMt
wPsfJMoLHBdVafnS9XMeesl94IxVOR6DtbtG7MUqD5aXf5WoML9qPyraTVAQ2yR7DzYPCq4jO5hz
5ZRP1C+1rvEh2DWcc6uCH5epYgjZrRx3xlWW1XkVZgMx57JQvCFosAFXx7DEKgZfNHd8LKVukgBb
EXoE2CjOnfpsFuI2lhHIe3c35Fj+KnOH6Z0jmgD8h3pw6pEFn38SjTCtYtyvDexdKSgQ37Fns67f
s68sUwiYP8DkgkQbkYpWLaK0Nx37lUvttPUk+E9PbtSZiWL2JEJ23a9ewMGGfXT7vIh4P1iUho/r
bBDcFCxMznXYS+sybO6uG9Uycc+JAZnyFW3XXxBR0zIgKc30MhtwIU0hXAz6woM5YC8LzjUAfQ1i
9tHWqJT5aoH89sBW3zSzYe0jyiYYV1xfghJWsqzG1fdFGgdwseMQgNPeDd0agz4vnO1vlaOthkUJ
C2TbBt2BrhFgwhFI/uzwcB8dxAe+FdV3irUQU3dg/Strz5DekYWPnPF4wxKJ3FK8jOMvdq8vDbbH
laGtvW52ijI1UzT42RYTDG2HmQahkbctYwPvL7HEaLEu7HGfTSWqG1zIPCff4YGqOkXn8YMNMBuY
X2YgFhH6Boxdd2bX/R8QktaFj65tv9lh7s/OAKhEbNlkComnC1hl1GqeEtLIsaP/DjfUlFwqd/Kv
2BF+qByjidj5SXc52+ubyLzugRenCX22o8Kv3OxNJhD1N+fG5Q0Ada/CAvjW49gZkasjJ9pk5aue
NZbkDqDo8VjI/yf4XCZCl2AJu1ud9bOVp/o2fKdWMLlOSDu1U0C0StnmaPDeHkM6jZA1e/yS8I5f
PHiatEM+nGTnVOKkNJQARJZQxqB4EvAydMAlm6RmZwQF8dGzJxiOFlzczuy9V4T9g8VNrBVPwKd5
TovJBZe3lROA+37GdLhevq69UgaiF8LuVaWIhrnwwM769X4+HR9bs0430xlDxT7AmGYwNzfS8/mM
Su3T1Z74VTQVYtUuOpFuEMmn89TSXwkX+HgBfuV+L9cJmi3hzMtd75HCu8Coy2MqJD88ECbOn651
6H26O4uZ6qap6c5KI11ClcZI9e1UUt3svFYsC42PCEyuxvo/sD4PH1b77nPLq6mO38WTq6iz64lr
D21mc/YmDzO8mjti713ueRn5CaomgHbB4d5iAYWrQ9nfX+dfxriICzwK704XWCDfrenh9sggTOVY
o3LPFM6CPY1VwvBxINbW0ak7sKRT6eLYi4aO/gyDObf8foDa6h9jWs+EHiSML7KKFN8kevQe5MtD
2wYoFhB6FZWnB4yH9JeA+aIw1Aa/9R2yqF00Xxxq3AnnqWnFb4501if/CABeCWvcZkfWIQbfnZUU
makIJWz2LEvh9teyUEhWF0rThHYA0DeedOAgm7JU74RZVdDw9gmJrNH7q6mRSsVg0nu2joFNnlRC
agv2Amm/ckGVdJLnGKXYV2dUqNT2G5q34WGsjJd8kvqlUHLASJgxziVApS4v6a1eQJjHqjKwvLoP
1cyeMH1kTYOIy5DbZHU4X54GNRTNdIpJA/IxMpV3qHwWtINKCYb7rzdlhohOIQZV20eS6KtdRTlc
giLDq/4VSL2Bv0KlDWsqEJ2bhyjQDJ04nii0HurfrYFGBTC+xdwsYZz7+wMC6X6jsZupgsvurZ9F
QErZzpP4oRnvGZiDl0EicEnLFeUsjzmUyzQGsivJgSf4ATwXGJGN/Rh0CcL7amQmeXN+ZcBPZlfB
qL4Z0kctdwazaHloKA5BK6qt4ffH+sRSxN8lrclo2ij1J/zB68hUCWQbjssS1qtZhFvGKtZNtcJj
VpZq5tUeZ3e3A605QHTgNIeWjK2hum+DK1PIwpDI8wdeOBulcbxK1G/hClAhdAJy2zZD+0H+D0AS
fLRHkvOs+UPAp1PzyR/FZHUtmlrZzDn1qtgQsodDQYUtjwxaSnClD7/F8kcEAE5zx1c70lWl4P28
/EZ8hWS+Rjl4376uL9aDwuAZmwgK3Avbk8GHZMG66pauaEqYEXG1HUfdVTGZQx3cpDFfRaeojeKz
6fplkRJvx4cIT1+TPpFJL3FRotOXe3j3jXEeIWWI5dZaJbi0/TEtMmzZU7NRfCdIPx7+s0JGZpsJ
55Rb0ZMjHa+dh4yW+cxcnG6SYEzaowyxq9515oDAIhCQmsZhtldnenY7qsJUkFe/iSnIuOr6P0cK
woX2KejVoeSIePinLpYH6ZT/Jv+ENOh8oNN3n5SgT1S8OdbZHYx7aKHdeEOdBXT+puv10TALrP56
QSqYaXC8j7/9PWsgHinrUtIt5qAstbi6kn/G/dSxVT8Ux+LTKvxTT9cZyjYjcoTnvBMLwCP5tIH4
a+sG3cPPa6/6jrHnhiBAEurpV7bC7qaf1Ast3gXfRFPnMwEEl4q/8gk7vzCDI+JYsGwRnKGoDOjO
CQFespzjXfwf1Hv/jBkxpItXV2Atx4uBNIfPARe++3ddbIc8gQfVwMn3ZtgXypB0oNfSWwoAKW+6
h9KznOF/GqfIh099LWrRwIPbPgQ6XkwkJl1BtTpxKH1ucf9sj7MyQ2xVKwpPGR4I+oYQ1089UW3N
HsioTQGlgPJEfrDxomAPYhgqoX/Uhj38x747IQBVzGPGTAJUcGNJ9bxT1alntFz/7z3eIBI7Xpbl
+5VnGp0p/Hn60D87ChxRFw9sch2lpkl5JxacocNxlYdg6A7TY9mSAsMY0iUdTCsi+cPFellmVKle
ud40QcBaoqrLuAB4g7zOS8cFOnYW3FlgucvUhpcRpfvOxrTWOzvwvYLQtGuEGEv5R4ZAe8ui2bxP
qga4O2B4wW1B/zsGA2geCbjNyWyVx+lnwSrxHeCrf0XmIFmwAqOMTMpH8aUsBKi9zfQ9zwftnX/B
4oupRUTw8lex1Sxurirp+jOyLY5p0BY5Mw22SJD0eu/5CVd6+7UMQibyD+r9FtI8JXrJipq99krl
aLZTo6FPmlM8BzPPMZSuDgrc4lSWB8gMD+Ai1mdmikYyE31lGfdN1wDHOIjCekhtsLJiKCIush4s
nV7OjE87L1ZwKyMy6tOAYOetozSFKJGxSfz+Pja17w4zspa5f11al2w4vuUjtBBj+Xugymwa+0sL
YYlOtDr+1k5TbQB24qHnFldxkhth1lDAS5T0G0FiiHQqEMBh9MS6ZsKr3nEtkqwWJk6wzf62HMSg
lqRgGkQVx56DlrweuvBHm8K8nm5T6eEbfEqgfEDzqBJzeJh2glL6Uom2w3XJjPt8USR7c2g1udiF
9TlxydY7RWX+YoHR5HHGmHWdzfBsACts84nfLG4SozySsnZ/K1yVtZXMiQBaMWklg0yNmF3dx7/V
iDu7yHJZEjgLXLQnAlzCOhoANGeg9jUuZbug44FO+j6NqDL5JFzzvMNTzrhn3xHH3J4junTMugJZ
j/RSF7m12ICTlP5cbUCOCm02KO4Kiyrh36Q93Kt5LQZitYCrKjFJ7Pkq3weZCzz2fD82SmH5JgaM
s3mBzl4gVlwBHS2KsJP/YnX6YOHL51pT1QI5GDJBoDIRKhKot/hMNZzYKx4o8Lpt7pYK1JSUsy+O
c+yUOur3xkSpzKuDs2R4IZR4Wd8+noLR+xNxbVDf4VYvESJ0jwn5pQEBE6c5zhfptlaFaKkoDJ7s
+v62aEnuqlaRonXQ2pqqB3o/q+1OM5eUIqG+yLnB+eQFlvuwdQQ+DQEO350Q7dCQYIBl7mxBxPHQ
BgeCNYTf+s4cejLd6krmUNgoYU0VcddScf4IpnlpNUW/RvFobIIecJ/HSyrK4yPe1liyrDFGyF3g
U99p2PuOC/2qJN/Bi/yhCMW1ogWU7w7ROUmlJJHDv289k94AgTT9RllExQNxt0m1lglE40OO82uM
NsLOL7Xor30N4QJ4xsNqKO/Azimtrll8Lsvg3Y/OD4broOA2TYS7iI6Q6fxg2HP81g0gVQ25uzNy
m3D2DP5iFkn74uD2Uu16L6PTXyFrelTGdrddpzljcKY8CgnLNJnvsXS7kLi0R0DSvhTKsfOVg5pn
q9nV3i5NDzCDfwIrqYu9ifdxWhoxzjnALX99yAhOj8+1LEeaM+IiSPp/uGUAZkIhGgEEaaOgus7T
8YVHtU7YVRLQVwgkl8NE134wn++95N1U8XWXf1+I5yzKQh6aNYIJ8kG+x5a3elh3pf00k7PP0OiI
qZ5H9Q6r7UuBllz1GReVCU+YLBeB2KNq/8yHIdzPKpCglkaVHG4DY7squsiFFhXqgEgLcTJk4K8q
qSjQ+fyeoDKG27KNGqfbXsvjGxx/ND/u6ynQsKUDkOgmqVckdvjxv+A0+QbFbdG9SdD5JU3ogdE0
iVQqLwp6vor9rr8kKTkE5SiCzaaXtAd5wGLf/mxezIm1nyi7yNDkzhjRUelvp8cNPONtFk4TB61A
drfsy7TtQ+31OE/dewouX88XdjYDbv8Pp508i+4iZh98dctyijL+QzrADHBj14Mo+zDBZ3a5k/6n
jlh1leiwfeYKrUPoZyPMVRu/SlJbgX2A5NCOwsXJARoeQGQ3L3fQ5RobQYnmpTZokSFy7Vxx+mMd
twRm+4cKGbtAk/d+JhIFaipfxUXL8w3kdRn5yJlecw1/GCA+RHjlrH2nlaeGyYNeyf4eigend6cc
W4WZQX2whavK3tnoy3Jj9RFKfe9OVQY+4WjWAh1CN1+5Jjm9e5BM+KeY2JfvN03MyjAGIo04vUrJ
HAzRSzxnN359+WkCNj1A66ILYA11ygFTqJkjAJFinI9nIy8ctVU+1G+wlgzz9bqXG2TDRi9FUmRS
YugYicWSQ3hpBJ/TnQmvTxH+L+9IGsErWM2OVW99PYr8XIunTAxt1dcwvCET1ykZ4I+s6760Cotx
URUbjTTfZv/dOq0z74Z5vHwa34d35QU5ZtptihZ2Aje57ufYNDhwQa5o+1FFCjhY2MvYUpIaknN0
PajjefEH7JRWv37pVLgCAskuYCOm0e/OfjM9KPZZxE+RE1Gdm3AbQGGBXcbiWuWhWG6sdjw8Tjx8
O/I0G0HTdgZjqlbF77+FqBdpRiVsSzyPEXeZ3Gv8JGKm2PQmhWJg9Cvb+KmkuI1kRRb/IMj/diRR
9tDVaocOagM2SkzIGONywFi3R6oPfi9jjYCeyarmi0CBZ3i1JDlDGSdWAu8cdxq8S4Ck6KLY2/z3
0fPFYWH7NaJm4zVoKN22Fxc4T/lNeUiwFm0w0myPSghPlIR08ddnNNoQpZ21MBl2cM/53so1PsVZ
igt5rqEZRPePzvvjepyUb294oDGWMz+NOM4DpzfPIEOwRe0iyJAFsCd308cOSxofw2yZ5mhK6Tr6
GX/t4Y8W3HI3Ve6ATzwYKXj2GeDHhrAnV2/eLuDI6CUkaMsLUMtGd0/i70xdvZe4ZIplMZsSAW5S
uRgpLlfNfioFAdkNZLGp28KxqWYOfAHGOUmBUDpMUsB5Af3FF2KjMq1mOU7bCYRC1oLOOLLdz4mY
O5d1O0pnIPTgJjIOf35NslIqVUY6KSD0pankUJDiApgAdvMK6kOEJ1noXsa8L97bNcAUmZg+Ol1C
tts9b89BcydQbGZZKgd0kG/mB08YxU36mjmpYlRL8sOUa/MEaKqg0Zno15OSRY4qbNZ4ggOQ+QBp
hToYo2jcaPEYVWiGZv0yIXHiNh8v1uy0+UfcRqY7MT/Ma3ArWZxYYh1ifTk9sFI2zS/OPSdpglb4
/PY6NuaqV2MdSxS0WBZCbNOPM7JsAK5cLYs5MrtDbrMYGcZTI1DFYgf6Htkmm+Zj6b4iEBS+rjRe
Wp2RDAoLOvzdXmw3cGSrHbQmxzDqzME0c6Yd3Nne+f/9XGHb1totNLQSHrru7GyLytfPTD1WVPxz
55FtRIioJHXmT+bj0UgDu4CzuqqtXI/TjsGUERSpz64g9f0BFQZ8MxW3+xp911YpWbbMzuqhi1GO
DY6t+xZG/oj+sHmpC+F2aesEmIrunlJ21Ty1QN5vU7UheaF6mAD5KPScvuJlBheLoBKl3kvNy6r4
eJ/o89QXfh9hSkTI7ZLtXIYtJ+QeCxVrS0ozrP6FxXdf1Pxh/+Dc7/xbQQu4/XgyeXR63fBVVkXz
WUdVkMYq2/yj14uegiqq7jEPzweht7l4ZujAuDa6kgcET7wWEl2tFK+WiSGGJ7oZDRFDipuXvpDP
mP8lcfxjfsFFOsMILJhAa7DxuE8mcRoJTPQoMC23y6v5t/7l2U+fOJsum1ZToCwwTNbDq3I+sM/h
3ZRyUYAAkwivVhIuuWlopWiThLz0F/MQbaB05IsW/yFKBU4CTPMQn/Ta+CBJ8O2iAwv5eekQW7le
URdiEiyhOWi5XWDkygJDORR17bmIHB2c7RXhYRxS1N+dRRShaWslQIxXeOf7vp8vQWAXO2UAItA0
SABIgiVdSnwZodg+5KY6iVAxfpcHD0s73LVFVxBC+uoWkiWmffuHajA87/vYsGfDNad5RE7nDVjL
4Ck9bpeV03MHd1nSYXuyYqq1DImC2E5a42qMBvoVBXse0kUzjaEQv4sX/WinfEJRzCmbe0tbn6Jq
FNP6RYBcau8nmBUMcLYmI95RwHfUqL+zJGP6we61vB4JzIRaa7T0mPrSYqrVn7/DI2061SD4GJGI
RBzLlqh9aHYYH66xb7OdNVpn+DVLhrlWg3phhy3RwE6arg6HwTCt8ID30xIZlth9qoAGeQXfAIE7
+i++qeXcMO8nJzKM4BwZFF5csxbtmPxgEFkDiONS1c03cdxFNZp7zFItP/WzjsxrKjlrevMi5uSB
nnPqFErzhBlcXOdFoB8kBXQH1loug9tUs6uKsWXpSSGoB4agA6amNmImueQWTT+4D2oLvW5TS7i+
Q1qcamTTUE47z2TUFqOzn4UBVygAvS0WjG3ZG+NXi4u5FgbIRio/w5zDHHMnKPUQ/h9bL4mjXD/E
bo0CwtuzuAdH/W1P1WlD4C0gpTBZumgFKWhpFPTBHBy6lxrjSwljeC8qzBktQUclUC8t7K8EkVBr
uwLasO5hVnaLtAzFgyZLeodBTWPKBbOvEHN0mVNUZ8LOlxNXTEOn+pBGaUbMPEawjdQRdlfc2kxm
M1TsQw2U4qI9PP2BCRmHfMoVLYO+bWhvWYK/knZym5SLBn9G9zEaBmkV3TwIM+IO9kyi3IE8KRoV
IcDOQf+iUKxLlWNItypjHQXr9AKkX72tD037Ofv8hzMNM034jaFGIeaJZ8cnKvl4v/uNihyQah1Y
GkoBK2BDe1FWpyyS1PCCjreGc4QkHyAqLVx+pS5E1d58BigvxnwXi1HRmPLrnnbzGK/paiOkPW75
bE56FrdiVnD+Z3xNPwrNOux3OAmdnAvKqA2B1WqRyYzXp22liqJ9/CrbDlVQtf9vQENeGPx9RdtO
kmRGv+a0IUbxfjGv/SLUPqPmpHwgCEwqlxvbxn/0zU3SuBK3lDdPkbLnQegG9JiTqgjWaScA80zM
+U6MXrIzQTk0YVa0wJO1Oli8oshppp/DpKVRdBqLedlojo7EyCLSZgxTebO81OmaPl/O7UZzTySD
C10apGV9RVkjcC1PgxZwvS1WCMhLoFRmDk/a1UM6iV+P0kI1rjwv+jQzzlhYA7UJxSqCX4WwN7Tx
S+Eqj/EaIv4Ypwv0ZGjgzZiac2VpCqtAHJ5TkIdz/iQhz+Pdv3oZlDLvEN0ZLvuu3I9uVDLFSPyw
DQs6Noy2PU7WzLVNrhaAjCVTDjn5Swz+Z6ts/nSsHVnBxSVx+RxPxj4+2wB2BGArT5smAtFJaQPT
mgYagqbXNxeb9+8JogBLX4HeHaSivbstTfdqVJkwLAZG6bWRm3pdSS0GaRnAMJaBJ5NF0MmkJdCz
g2eWyHiOZ50FoVurHCGXErZm/zNqyFJX+EmkXXxY32pTrEugpCpeFUhdzsORW6IFEkmqMI1tWBHT
dVH0dsC3vECICOBwk4kE/cknCbrNV8eNsteOXlqNiYBNYGo4QsyzM+PIDtv924iDYVM0MUr4+TGs
xzLIHihmIg==
`protect end_protected
