`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
qQPuRISTa6yTV8jVnjDSkAIpWnmjwx3kjaC0UCjHjlxURWKOpytjCpREdB1AZ3k2rOuDKh1tFF8z
nITOmdZ+PA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FhyfW0Ufa/XiVrqmx03BtroBYCuU/mp6sR3FpSaGqyKkZFDoDRM/ihUn1g7Mo5KFKFOSABJonGsN
ySOdGYVbpdRsg+OrUW3RdLHpdOFpZU8uDR68eu8kg0+zwNjbrsx0HbvIeLBtwr0KoQQhu2pBS4o7
mud2ji8nl0taVyBozi0=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BE2ncq3uF8tnDn8h9h5fHM742dMiNCfhsDawJ683Nw0yNiSjTQ+1d/6HbLM/tVbYYXmmcE4vOkkH
Q674koQDlJ8wgf5EsB3kCidNIx+3gkuVo5nM1zxATzpwZECCJXm83EQnDH0Lv6xY/E9Yu3j3QKGe
+7xamN1cUjgh1fWgZsM=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ud4BXsJG+kTHw65pOwWDRCb6uxLWdd9nVaHEr4rkDstKTWriaxV54Z5dRu1HvPL5yid3csZl5XFu
Dqt6IrmXo5DGMSE/fbJ3/tIWfsmL7VpEq18NRtSZf+NsiLguHJ1xMfSMr93PXkqN3FYvQTV2lx5R
Rh16G0TpvTTy17sU1sJYtmrI1AwLDEOv+ZF7K9m3CUqcSylWDzQSikoB0RarzW289igUg8+5Z31D
oqM3r0L7QkcYsnW57Aid2cLxQYI5RWvSsUrIJI1mGRNl6n0jKx921ScNSQMdLfe2+GECAtQDrVVM
gFAPQsUaNLZFH42qTJKd5YumFlRihpR2lJRYkg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
u57iRnJNC65201+394O6893mBhn/gX1DDYraiwctabLy3auAGT0lhkyBcSKHCVSBcnA97F7TrPv6
Vrw5DVlmCk0ORpBhXNgMCbU38+FMxsPE9rR0yV2mdTHXx8VB9E20hL599rFWWdRK/Hpy5y+/jNSk
FHs3zI9MPUzpQTUWQot8qn9ytAI/F34u54jpTCmeTrde726xdwGDLqSwa34CS4gq5jC2MvL4XbWn
5lrObExedvHU0nQuz55iOFW3deuwcJUptOVLu7xtao1T2SzCY+gEsIZD8cVv/IL3i4xjdgZAQmMT
k4olqiQEN+P/sz+tMSCknLWhaI5cPk8fxGQx9A==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
N4ZPkdFwfTQ1lL432dKkSr0WfcgT2w+0TqO/8gZgriW7zwcrd/NY+iISaE1i9Fs7OFpmQrowLGQu
uH50L8dpIcahExL8zepWhTPy55u1DDTRe98Nx+AV/o6cN/RKUJ4o4sSAyVeu6SJaqLbMk3ZJKH0h
POekpClZIjwMygSY51H/hIoszQ1CirRsBoYpS2LnEpIBfX5zusKBh69V9rwpWTTku+HkO+vyeWaJ
Hifp22CiFzTBTyGscknns2X2jgjH+lpcgN4rGz9skAFqaRqb65f2HM80biITmgE3dh2UbVBu9Fck
wbHuIImn+BU8qZkUUBcLw1JPYKhdfQR6mfTk2A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 296032)
`protect data_block
PK9g+yub0axHWqdSITxQ36eEOc0XHuaQcwDfgPQppCb2wrgYVIRzmb7uMyTMFEPVJB1ZcdW/SWou
zwj7n/fB7NseANKOWCZ/w3Q/aOVXp4hH28hfuWZxsUschg3pTTHhz0STRTjuCHYyXqPlF1jsnlnU
HuSXeVyskycrFY1y91Dgh/GDogzaTxM2st6sMpIjMf4u3sGMGC+WjySsA72FUPQ2PumTKZxnF9vl
49AiRHYmtX4MwW2dXEzYLUvgtdcIVP2km+EjO8o308Tkup8X7YHMJJt16pVUydzJRpDkyAPMuYMp
ysRWgMNUHC9AwBUyGYOoiGOukO2/cGEL/m+jE6wLyQbsqRJMQAGVS4fQLCLRm4usThgkch4P7oTk
YW2sFjfEsUZTK8pYP+cwCm4brageGV0/FAZF+6wp6Yh6svJ/wuzqPakyzqIVDwRHwhZ4ClBGwaFv
HVNO9s+uplSAdu//LLJrl/jxhvFUpxt6wWVdu1aGE0TRIxhXRwwjDr4hWkPA6UhTyARQqU5QsFnR
swJFssSOWeNdLnZWYmCwArlfPRot02s9oD6jZeZbWJLLDvP2QIDPOMnjBENU6jgv7DSPKnnEsoe0
eys+6meEYQ5XUHy4wwNWe4KCQULfbyJU9ffMsszKu0+aFpI2Ux8/LYmB88OvFwFq53ampmjTqTKv
uoizOBakt5jat2LqeDTxMfPo67Tc+NicgZ9ej2C3d8lsG4PPE76PSE9XKKJn7C79ef9pWXTlFhdI
ketDrPwKjzMeDqtD6PcNlGQEBKBafT1R3JS+wlUNco95fTavY3RdwKnhhOT10ZZKGEWC/xZ4U2Im
0r65NKsbZz5/PF6yVBSy3HXI3/HaYpmYL5w7xFUoVFqc2Yk7FWz1rPkcgQolZfclniBJP+LIm96M
NtejN2SFSQ+qWXyPIv5mfK/THq0hTIMc2ivBbG5zhVYCvr4p+Ei8sO5vqEj//ePMDpMDPnSQcNFF
2TQ7URsE5BWYk3VTI+eZRwD0JSakhIgkyf3g/KpZ3LCUwaYSiyWaYeGfMVtgC7OtEgTxL/eoTdGq
gE/rzy/1yXkY4yshcCoU7eYMiEhdQfSv3Cu1SQAsMYybsnhYTONfTaCZPh+kAwMTfQsuV9FOhQR2
tm66lNjNjHjyTaw00lVTGOoxKVoI+X9BtM//btlpoxjb2LyJgcQkawSysyH+Kqt1AiVOzdzUeNS7
ftz56JmkWVSh3KWpcFeKIBzl8WeE+4YsbPmjnzXcQ7hfRxgWFnAx27Um75yOLrt45gNy0I6LZVwK
AQwoIUe1ICluKfsPZKe6XDUjF2hfwttUbK06VW92TUQdYAyqrj2HD7SRI6cefQz284q4bpo69Qw8
Ff+encXMZGe7mHYAr5Fs9GwsAPB1ADr6umByQtJEQvage0wNIc3gS6feUPdvwnDnC3NeRl3h3U+B
6F/VEExNmT6CKowguWu6SZgxS3dTvL7vuOtRiOzFbAsGs95fGpoocy+RMBPOnE1zfrNo58vzKDTr
B8Pv3ikEnOqxIATnGy7T1SEUrd95MNHxeFELrlsogAdT1PrSwtRWYK7EgA6fshxJssmfDQFiLmkJ
Nm+kRX5KafRTrrxcDOgsjtPhlTY51XB1tjMbYuGNLu/KBrg9ssoXdmLpPgq5xzar/cx6ltkBql5Z
U2FcHbDhJKpGvlJdv+7wVcrvB7Jx/zPVcFQZT2z3s8UxzgW3Khff40LlIbBgjaqau4GshUKulAKz
KNUMiic56dGdHsj2RPvGr2i2KriOmjqhlck7iLsLEAOaZ1BLTOuf174xKdvqOQ3ckbyGf92Bfz9n
Za/rNvqQ4Dr/9DjlEdgBB1IIz4GejKEWeo1ndpACfACszC+cHPtfnWdfSQrjN9+0KE0Pem8xSbgv
b3s82tyKNkHJGCJNhGSX5T9/xZt2dZ1smsEnqo0/bonYBQAEyD55/FAEC17KALZ9kCdKNeSfvANi
dNkwPcQduSqzXOIkAr39sRttfmOjbLhF+Lz3ohFiRbiamsjCpCsmcoUSH3rUHapcXbBMfcDP3O7Z
YTu0Mwk5MUYc5F3WwLN9oX90jIPVarrf3IqK6l19yGrUEkEwJGeF7Njf/bcHCKCLrJARNvZ5NS/Q
bpVN9mmk8gUsYjKBg/FAjQrXmmJv8ueCN6bOfig/Mv1ot8ztA/KHyrcP+oNf4Otkg9fYPavA3i8c
dUQOZRJTRRKE7SzG/NE+ThwvPt8ZAPR4sZjhj+zA35FUGhLO7ekFXnM2c2M32ZEt7lqupywYVehO
LVnxHZld2aQRmeWBLHv0q2mkMggifVCrlg/Ix7Eig1TByv1f/F+hhmn+TCKN3KUql7lOdg8OrVbw
S9F5HK8XlP5Qhfz9TVdALNxf5HOxaaQJUOVU36hw9/ZHev2g3sfVwNOm4REizX5Eguq0xSY7FN5O
Z9pbNmMQguxbWDiywtxTxKJZ7FobsycJREo1wNk47KWkaqTG+w5KjKL1dqQyMRcd7vMjugH7AlBg
AEYG1Nf2b/BMK03eGt23HAqK3o7+2ctqBSNB6Egz9pOamn5sjOqbHBKykOf+QgYuG/QqQ0sjZJtH
yFjpvtXrhSz3uYqy4cylxou0lMAK2htFWpIT8ofz+JxYwLvqXjPThb5xCZjU/2GoQiqHGUlTe5Cz
AX8oSEkr6LGjJfAmXvrEzO+AHN4mOsW9NAg1k1nblw5wjwhNyXsuRWkI368CMFsspVNyRy0ho/dt
ZJdmMbz9cDx+96pbTYHfA+vC36xjsw4CFUTriPcsEp6FbTo2Lo67OeSw/yF4EKME0mqyDf2hemP9
bBrt+KZHvsl89FnPU60EOXh08flToEpnh4CEN24dXUH+wDr0NF076bH0qpIC0YVlAHiWRaTbzM2b
TYmgu2R3tD0phlfCsdZIViAgnft14R0eNu8XV22d7jJbqOofItyJpp+hIMsOzSWdv/dlA3yOhizH
hjQkJCeNOEt/TX/gVTuV4z9Gx5Em4cxtZrljEFQGNIEIUYuQ2Z8h4P+feQsXH/xpN1SBZSHaGta7
YUMznt7Hvv2wLiefmcl8uMxzoh5nozBavqn01w4q9U7PsdqFKM6F7ltJuP0kQziawmmNg+Qn3+0U
Hpw4DmjpvMW/azzPGG0Pjb6NG/SDEoACJbrMa6jhPUZ3ERrEzaLjfe3OLAcYZf1xHKjKhy1FVePQ
Ucn6j6NjNC7pLcqvg8E6KhWEi6GGm/r/h5LamcOMjs1lKFb2jQecOHh7UIjQKcwEhAgL+BOiZ46V
s1NI1QAyzl5D3etoY0yNXKqVeZa7dt5/0Xi0yCRxJYaGUfp3kl32q/c2shC0NHU4OELyVg++LdNn
kP+cbD9z8BZSSmJlje8DzvuWtxR+UD+dn2mcQg3RQWajK/PxGjdhYSrVIce4RCSz8grdoCzwClPV
JU33qtI/s9m/txcfbBd7TKOchqxIQdiyuBFlLgqY5MSc10sWqhQs+6LLCOH23EjMBTS0Lfl100Vu
tZTkoYoZATy2yJOwTybdWfdmBmnN4VaFU/vrdpgHlIPjThwaCO36tcqpO4ESXNbi/ZEqMWc6EC41
chnIBkv5NvN9ElQnTMSsVlu2M0DIQAngtBK70RGl9yLLH0/LuXK6Ay6aaVSRJy7UgrDkbdMuoia7
syXN2xy8fW4hj6MI9eP4J13Ll6ePlNwwwv0Pe33XS5duqzChZhTTlV/gMGAItcWSe4LmQUGw0JFA
9SMScSs9pnQ3RRWOkc9axGLO7ogDdlY2SEijnESzFSZHTksR1quiNxIOyo5rn6F5ABQek+2vFH9t
7mZY46Org1B0dMawjSjxeWhf43YqgoQlDCt+G31lXZcJGiGQC1+qe17WmK0XNJ/g65AjCKaJ7Xra
WnGDs88U06kVIsmm969/3yPMbRAataY5fdTsWrErDf3H+QgFiHWWUrPmegWjj1aByvagp/0PQIHU
D2H6gp08kdEXVbpwEBVe4tEfJnFdXmmr1O36qp8u4Pza/ELW4azlTszkgrLqATAlEq1kqo32i9aK
CVlQrUSEo/xuJvXcZxvaklUfBwcrcrty790FUE9MzaPaEjomdyvlnioAyrBpcX01LOX8Z5AVwOz1
BOsMddlx0f3c1zr+08Qopi3EUUEP3NSCOao0j9ZGzgiRWlh+1Sd8GdLXiiEUmYM6k+2d8LhVGQPq
wtM2mlHoE+PSw0InYQA3nlvZJoPR7ClHiLv20xhhWFeOtunZKGIU/zMozoCTLQVXjdajNB2X+G2z
tImToh80KrwDJXxMvIG4nnWjhtXY6KKBOXWGaAgdO+pfyzrW7rdH0tSBmM/CroSRswZwkgItK6tJ
tHOwkwc0ljXAzoRpullVI4fzcFWLq9+1Ejrgdod/5VRYh2WZzTjxFvOAERw7raIyYgd54NJuj2E1
+bi/Btf0BH/xQoud5XVAVEhBT5uHyt6vWV9YoQTt0tWeFa8rjyZnSaSqCH4z94Lc4iDJtAi+xX2K
p4Tu3tysxtsCZigCDpUbkfdZ+SoHFJcxMdmYVdCVBYDajNFH0LrLoPpVuFsjYBti7wE8Lods4suI
uxPkiQgQCGg5NB4T88TJ3xl22ENA3i/AZoXaVEyJVbk9T7orqwAf7fYknIEy5DF4Abs5FtdKwHJ9
BXW3xjRNcGUQu5W0FkzBtHxqEOR/UOThhWuTkBhMFNEw6IBgfm9rBcvwEUF2Wv0jZOfnuIh26kWi
i8Ccn4ZpySbhPreFyYYRj49G+xDJpUrj+tYwpBGJyATD2x8ro0zMw5QDmFjxloSu0+Ymvxv7F04o
ln6/pwmrGaZ2rh7NB+a0Az+SJx4iu38P1mJokiBT8Lz3n0hRbbM8Xg5UoRE1mtUpW+ByDAV1Dzrj
eM+SsygaR3Dny6585OI/HRqkvoKslsdtBcZjb6mMo6mhAhxOQ4MXuoBsUwWZpcKuzYWghR0hLFrK
QMErvHH8zxemArlN/tRzEfJ3+AiedTUKxpCDxXpgOYvhUePhaXV0iOvKrcC0DfGyMTiw+QuO5w+3
LU03LiOHc+dxouQ5hyTrw4rwVheppIB9g7KqJBQ+fxR+W6DLZe+Za70Zc8SOd8KTkjMZN7/COy/A
GoZkmONfJlIE4gNy8/XbtCtR7Sofgq7ylhCesO8st9+R1fgfjdToILWhrp6i3EJ4yyIL5kdj3JIn
Q5pSNzUuKkpAj3W0HDw0KZkp/5JLNcaukSG1BmZUrReyS6S6lNyjJvw53c1wdT9+Qf/j86ayhmAY
6XQooIsBFS8kjst1Y/uHVDd5/2yc4PNNTKlt99eli8eRTo66HgjfbLrf9dTmy3ZEIcetzUQuZAp1
5Qxt8xsieNGDLVOyGKExTUPqfWYVJBV8VZOzHOPDLjCDnzZFP70U48KjWfwX42hGEzVsMMD5bNEK
V9vw0ldVgCzX7AbbaS1tfcY216JUuLCaiRRiarxQ8qNVy7otRge75Jx9NjJAbFIR6JoWg960QApX
Wz9Q/lFsGzb8aGgYfmZo10tGFGbemnG9WmUI0FiIPJ1g8EbyJ1YNr1udrW8HyNwO+TffVxTu4xpe
p85VA+34HNjIj4+mIz9wq+KdC2VnJp6G6MWDiKqWA6ddf4mYnfvpGDXIxUY5Cyvj8/Ou8474Vj9Q
qfWlmtmyhpgThGzUlwF1FqNj8yRL1BKS0SJ4HBLzSSc7Kw0SVCfXIdI1aEE/8cC7Ei3kl3YUSBwx
agnuYndE7b+KaQBH0ZxS/mXXFLhXFvcZ9mEJ9W4JH7cNloPRE51Ky+++rvuhLIxLzNk2i5OlNixO
4ow7rP6cp7RWVMvcf0yracpFzz3b0oFwRyEa4rMwE+4zQiF32oFbgp0mXPLNhLe1sPgB0rWaUlpR
x8/zEf1J7ez/GIjB7VRNkJY73IkaxS1FSyX89qADlBlIbK99hgusBCkzFueBcM09tHz1f0KhRAHY
0VGtczZMv5nqPQU70cX8TLDZYU9qgVjTH+y7qROraYvjecUH+FMQBaovy3eOZR4UcTLFZvxvucIj
U+u7TJLAiXafNc/BUzVY9RHmXvjoas4Tmmsttvx7EQlDTeAhQWHK74G9273avCTFVY5+hQO6GT8G
KmZNiV8aY7xCm6+Si36deG56AMw2WPsSEMzH6pTxBh+xlr22/9In0j0hhgEEzoQ3/n2c6sy0ZgjL
JkGgm49eMVmA2H6Yil+YRivZTaHRQVIGsFRCo8P1BKzcD+tAUMQ+ONaMSJKC7LpPYbudwpUsVduD
6j10kCsh67Bf6OPyws5drE4AJ/WyeJpd58zM2Kbx696cfu/5oQEIvYli4TGZbNoXaV/b9e8GtbUH
D4dgO+X3t6pdVMTzO/xU85qz95edk5QgrMkESl3tIkTWxJojUYmMXDqx71KsRv/cZ0o9hRB0CRtg
uYxyB9zN6+7A8Rw9FLcIl7pRCkdl+lRPnOjUOVXg3GOMIzym9lbaW3CaVV0GJS6f3eguTAiQLog2
JZh4IxvinxQW8H+LiF1foWXGk9hVp1QNSz+wgAkaWjPVD7D7fJhF2x2bYTacMib4hHj3c3mcV7E6
pBB0zh9Vh/HWmROuMa8FbLGdUCWF5YSoDK55HQNJ0kZnADsBEQM7FwCzZgFFJ874AlMZrDJ53pEw
xdDGNtyDX8MXcmNwDzhzMp6EtWUp0VTp9G1Mi6py/0WuvwU+1MpYymnalveJxOBcDhMsX4fYy/vy
8i0b+tlCS+vTBWzXID0Q955z2DPCvFuQThvQW0hyGvNtbCQzZtfw7g2mmFWcI+KhyvKmWyuo6FpU
gJStfr0izf4ZzUgpZMJdyQbbGhwaKpinHgS9B/E6iCW98iwv7fgyWzBsTaWDxQlTu385YyXuyN8r
bHvjIfIj7DADDRnTVARRLNoFqo4Ri3vo+o4RjOgePT78zJKlFLQwBjY7VT/L4R1nZXbKG9dq+T1z
haljwHFOAK0eCMDrzijJYrP66y/yIYHYyAYoHiNf8Chpf60Lmrmr/ujaiwuSk2WoHJVBBW5D8Ele
OK+JxUD2ad6r8IZvdc4uWMc5JAmvQD77mr4BSiiZlFNBj0G4DRiixAvvkNbRuJ9/iz6xtI7GVe+o
Tk4KVjAnpuySQgUd5Ia/fDKjCl2a1WGBXHUatzk7QWBuNXnpHjyA4F18yqSgaOmh39Qz07pobvRH
uf2IWthP2ecJfmFYss3Ye+yVDBj8I5myR6zzUHJizuzyAsTcFq/j8mZKZfJ/56hdRRHGxtTj/4Ig
gs6B3rbByKGD6l6JIY/tx+iENrPpI0aIH6y15uRnLt9PoAq0IHRb/menydnIJPHBb4Z+wK05Q6pi
PI5/KYWX+hFhm9ioa8bDRuyXSJFPAoKelzESEXKsyaZmhrUAKyXR2QcNjw2iHQ9ssriNLLRYlm0+
I7VWbn1gNzjXTyeUDjsXOyNE/96hWjbzVF8DZIH/Hl7+mReVjvRQ+CZIuOnDhCuJDU73uom3a1sa
717ObVB3Ko1jFlCQ4ChEdcmYmXrDpCel8ppqhPQ9naCS6ut5cOoibLKq4f91meyjE3vf51suMVRd
A2wNR6Ikqr7ayJ5C5jv/AUH+IuJzg7lYaVg1VHkDeV0a+ERjdm+3smiCwsakfWTgut96gqLTm4A5
Sx8k0HuMu5CPh/+1vo+zqMfJ7pensYkz87hCY26Y8Jww9eCUo5FsS2FmtXRPeeL/bpOZsLF70IOb
0L2UfhM8a+Do/Mx9EvvB+qdd4rgRvXgrfd/ASP8NTPAdTctmkzzzTT7TR9PIX2YbT5jW0uAuc1fq
7Kv4TsGzh0M8mXr5HZUtH2c+IX3qAirLjdfgzd/32cs2FTt5tenC7IKBpKuCpwRMIFxPjyt+vKsM
6vEtRUaCJM7xtqm/HG7XT9tHrFNDW6S9DLc/DXjahRuo4Oyn7s/VtR4aoC+69wPd+0B4+Ty4qsRI
8VTYTLGmOYPYDjhLgAeVCZDJtPHzQeuZsYRFVgN+Wx7EoUxkGLAxorfzG9vDDV0AADFob2DtnLJh
pToTVX9mfl78lDvf7Lw721Yrzt9AXbQ/S3b2AR4/sWDN7/mpDkpKhBwjHQrWaVoQ/dZ12SA1Nn03
yuxktaNckDFPoJkyZWb/Wf47EJsiyznAQDD2VRQ/GFiHlcA3A03gQiXc9XlWKLd0HoIFKO3h8Uiq
ZEVgZZOPfp0autYwNm9ynmbQ5Az31gYiiIPE6IN3vsZf/qm7rbP44OklOl9lwXpTxbXrqlA/lh9O
MgnnuDgL7/gBUvhXe6c62aWHpTY9r3K2teH+LF1giptQJA0jfrzUzcev3LgW7VlRmNoa523gaIwW
LJTIib39SGk/QUTwKG3PQewMh6pGI721Eu7eGDi9NhtyJGfK1rn3Iy1uvXQh3O6qsjahSFemly2z
h/E7SKJ7M1OaGEX78zNFQkxU1+80SY5O5RJ8e50iJJ0Vkq8A3mMTZLMkrA8vq3Z0JyCTnlMjqS2R
bHp7yRMj2oorkdRpAfT9ZaKl4E4CpqkxOTGrPu+YkOyMFdbOVgQZIuuR7Q+QXTV9jdLsTDrY8DIn
M/XETFctDRkhCy5llGnlo77JgFyviaUXy+uc34HiQFG1rX1r4Cw+NJvGXV25zQVehsAKYCop9xj0
x3s7rVvBgC08jIj6sg6gfWwmxJm5m2FGtuHqXp8+sq14EAWliaQPTBY5MPxnrxOWY2qVfy1BmEBr
GiLGP/vPra5iJT7f9s1GYXIF/H4ruq2F2aikYA3Vvot3agyA1W5c1oeB/cHGQoCLSa5zbB5r9rXV
ZDOza+XNe4XVUnoZD40uzWRgXXXCJl+E2G3QgA5QKKIhW1yfe54vdZknXpwPdm5aY0ydJIHxT7wI
teDSy7CcunD7zBQ1lCVQMKqhIHjA5nQO28MsWzWRCcL5ilVjiDdda+XPZaKynEM4QlXneR+W+nYs
WvEuXKs7Gq72kzkymOEwDMwm4H7XAnJr1EpJgnfDd5Fj6qwNpUtF7FplMvdPoFPsR5n/xH4XIAzK
9ZpTW1I/Y1PUDyG1XjJdFVaurU8xBFn/KSDl/eDsiMZvgkbtyTVrS/ylNF6hVgBnXyt3piiG+SKW
BxTiYwMAOKYNeCPCgS8/CY/Kl9nYgsMDk45ibIyYrqtNHMSCtHxzBkdu3APPrYAWnGwqe54kekYb
4ZGG+z+UuKUUBl0Hmzias/xcbthMJkIXxwq5jev2rFuQsSk5kztx8VBdjmk6q2eP3qpmUjl1fJj6
h3WOigMfevNMVEYlm/eZF/Gl0+FERKbwgJCgnnP3k+nSfKrO3yJ7J0o7/J2jVLuGcRYvJz1QMNFU
fQRg7oRHAxfZSpPyQ3AI7Hjg/k88427JwVGLKKqi7/T+U1QnVFjFg1WVdm5KurPRcu+4hCm8rSah
62jxTF6P0uYRqsE3mKlFnzFHp+z70CYWpGWJ4ZZMMxC+hlb9ZGMETnMJ79OPx62HyL0kTEKSbprW
9xsBn0t+t9K6FjlSSb8aoH6gK3xVT2levCrA9zHlnmjrV01Sfi0dtBq41hqiOgvfsMVkE+zY58OW
FIq9ZZN62mFsVPuZusJ7edGKWDuVqTckbtPKPypuzXQGaZbh/m8e5LWIKizZJXF1mqdvayo/Vqel
uLInOxqpEbSqTh8Oz+dQu497BzerdVQdG9hbBhGF+S2wZtKgPvli816OZfSUiHSx+EdBRLqIryBo
Bq+pcxUOs0T6FhgSc2xiJoh6xWQxXyaM5XePmUuWxRoaJQKU5WAUYHAr5+3QbWkGyI5E2/5Ta4B9
QPqW0B6kocjV1rVXn/KTijbMmrC7JgcP876aeCNTBGOIzdJzb55Cl40o6nwKqlAGvSnpAHvPxMiN
6nPhYuQcSlh6F6G2cdsgLbwG5LPEdk997YIgimbOLyg3cJJvx0Z+pMOU436rqF3/8S6COB9aQ4Oe
Wot8JheRila7VTsH/GnuE1zccdXGDu9uTz6H5Eo+ocHu5ltgh+axc5lSUL28d5fYFtDCS7aPrDuU
7W2drdp/+z9JTx876+67tmT5DEDitkaTTtZsxf6ezphvADxzgJ28jW3NeiN5CVPvK1CEK5jzyaSd
3TAANrJM5fBTxqzKLmVUx7yry4pBphplHyQO3l5tSzMN7TRP3Ib0Irp0moqdkGbBspeiIlpeXRli
3uC5Qq3GARuN8cAMkrmZQzGBYM/VnHV9ns9XQ83uRX7KKf1lBqr0j8hVSl+wD6xWsGCkMwKqxLBR
Z/C0RxXLLLteczAlsZQzwJ7juweLY+TEH1EOba3Rbemnz9JGKVp1wN1k70bpD+BVW2UYLYQLuK0c
u8HKHc23BeeJi9z04aPvfPrSCF9yAjRRCRplDIqx2YFITKAYqOXmvYj8FFF/P2KN5KZkfGlj/lyl
+t3+AzwVCOHAehqqfsuNs4EO2CiZl/rvpdSiOdv1tuAirz02QVyXF9cui45QqhTc5KAE9524rQX/
115MhFrodrPLew44n+y6+RyvXI8xzesM66xPLuJU41tAIOmGC/HQp9Jq3hBHskXWwz4glR3T8VRi
zUxVysSTPH+5OIBGG6vwjY1NXKMgUVyTmmUHYDVwv9oaL0o++azYQMJsUiWT3XwimtKkuagrrZXW
gH2BF7GWmu4Zpa5r1b2hmgObmaokMs/LQQ1kRrDUlmZi+a1aHZIQUxZlKdt7cqB/omR7q18U3CNS
tq6vv54g15LoIA2CmD5It1X0llonLE1u4yTgUANXFciCUV/K6Jso48xRRt7Sk7nNyGckkXPFa98Y
GKmLUGW6SBP6a6mJJVWa1oEOMImjCVcLjnZ5LOMKcBmj3u2h4eKzMY9KhBsHIbquPJ1TY1CgKJcy
YFgjJFWLm4AFBpFacHNG2jNR9dU3OWF4BknlfdrGP59/rf52Mja+jeseRcE/zsdfTzK2uhStaUUR
q79fhqMEB6QXMPtGQwx3u8D1CnW1qfUshUXVOtWXWFECxLNx5pLi5Ef22P+6hUyw268XWAKBUuBz
8I1tC2UqC2eX55MJzMZFFwWoxA/Qh1+ewWQUs+3Ky4+WvF8kMisEftQZyZ8AUJPH4BsJCctD096i
3Mf/MT+81FJOGl68qwRs87x8cYqTy0Pz7F7k1ITuF071mDi1SmcqC7xuJwOmskRXjABxBWl7QFK7
JuPvPokmURrvV0rSNnfBSzrZ8O8mfUxFkO0JfXVW0f/R2sa6dKVjbBrcxjFzV/xcPsIh06rXRpiC
g8aGsMB8R+KkvNV3b1vjarjPQ3ayPPZPgWawf+tyvOZmdLXGLdvXPcG+RVlNzhhe8yjzj2f1rNnK
cLGzpze8CXKV6le5asCNa0LrdlYrYqPaXcj/oDOzRyh/Cwmja1Sn/+Isyy+xovHvvYSANKp10zv7
ywz4o6JUi/ni8Dmikq62/hWobCYmhQ4TlmQz8plYsngzRw0I46GEP6mTJwMRKmCgmqPHf80J0XWf
fZHlvRWrSSaK4ko99iDQcojR//xYjan0xGIukqRNWAfHELOKM6rvEurKLJUL3ldkX4V7djV7P6qF
pnVe53ZHPJeIIVM2s25Lynd4g16EWuoUa02lKtgvk/ImGt4Am6oNS2IG7IHStZKUjm+ONc+u9G/1
4mH+ZMA4Qnqtq4hDujyJZfhi6SVSLoQEUL9zIDEIWdO7rzPKGSkJWNxHlYqOAHRs8tAUz0j3Ytah
Aw3iFlls9ExEi82h3DJ1RjAKKgIjoGK+7dWwcm16hNpgwONq9MtzHXHGHdpX/N9tDUEZPQtC76hp
lbLqhdaTkXZIUA3W9tVUJKm2hQ4ZWY2zSdPSOJfD1Y+1UX3NpJBOiH5d+IP/7H2ailihly6dXKf9
R6KOytEtpRyIhQAUcJEIzqgDIo1XtHuvVbF5YHYA/jfHws15sKxtgbcfOGBwZ+3VAPeYQo2HB0iS
rqMssm2lNzcJiw3+BejDre8WIwzESSvGJX9gCW9BPXWQl3wDTQ+4j9W0c/JnR7eJOAtkKG+nIpqh
14m36xuRn5I3xtG/86DqrlW422OR54dujFfRLRZLfcOLPqsfgsV6W8GIjNp56yo98Q1xdJPrxA3s
r8zapRa7/xrvF+AoNb7AinxXC+hFWFdFn/j2eDodI1i2bsvspi9gW9ieqkWdOXopEf0mnSUO/pYP
kWbyxFUk0MC/K6kss04tn/sL57uDOPtWZ6VNGrOu0L2nNFRfRoqY7GiQWDJYReXK7zOaRmMLxZTe
eAUIU3ZS3xKQnmrGbOkaGokqoMEAE8D9WsOInVgafUYqITdPGhnHbDwaMGJuWuLvW9UkPdNki3lC
AWsxtKJiSLuRt0O29SVjr+wtCtmwFMSDUaYMyUO+fZzYW2cDmz3s0jgosqvgmKX0OO30FR3mF77P
3vREKdD1vj+VpF3jwj2JYuqbQrAqvxACHsQgcIptnQDMw6yvXyMDAh/CCP0pRBKNpwq/KY2yez4a
ifjgiNkm2jYUBd9Euz5HtSjS73cFkJSsYF9vGChp99Zq2hnFLPm42C2tuLFdqnArg+zWb4ooilGJ
FArIgKQe8AZowTvSQb/I5LT0YRaNMQRz0IWiv1gKhLNPJ4gIVPzXiKkdWd8EhIRLbNW+FPL+BWsF
kpkTr5x0haRYcyHvsmm/O/xSavXAlWW5yKLsYUkPPAZ1op6YxotKpVWzexRjMjZNxDkOepDQYNml
L/iMI69qt+548QTqPL5xaRqNBSRQzjzvZyY66ZAt+kh9cR12UC/ngRy1ijwdvaEEvcOq/LJ+EKIi
E+aYYNNhoG/qFYGEcB1SGXuxhAsb3lp0YsgYz+qs3uBKChvpfrDuoa/mbpbvhR3QZjPl2bg1LLil
2uRcA8MBtzrKn8OpLOii+o51zZdcQt4HQngkCgMZUDRJL/2p4ltzngjNvqgskyDvmx1NoLam/mCU
FJcsgTeiDQSldCeYY+lxQMgxsEnu1aKRiLrspS2sjVF4udxgE6YOx2xKBfONbgXxYgfXllNPB83Q
nHybt6lIufBgpeGfux4+PWoFjiqnRwPv4clVThQo9SfpI8U3fBPdYnYUnpD2yVEmbAb+wS68bs/+
XesAE4MFm/Dsrxx10L8y0kCLGnrGgQyrzUyZGOhIbr4CZNsFvHApjDJVF1KIeGmAYOT6GjTb4Ptn
2qpRK6vcT32nFrheZ96YrBGYLX+6heCmUggNnGf0LlqG3sqQAFDyFVg0GIkyqRADjxxzfF8VKWgU
tjh080xmy5ju1oJrRCKmwz4DaxGgoVYUDqGrm2enAC8t3oMKMSU0YPNSAdSGLmVA2PBkYewn6xWL
NLT9g/LOP6ZRoA6dEvH1hlkR8lvz36NUK7/VkLR0WJyRlNcUS3Fh1v/JSPhPoaRt/DLGHBQw0N/W
pnSHf3ClvrSmgz5nT1SVT5RGCPZphZPqTLIiQ62n7QWcfYbSjVa3Giuymcc2dM0wN5Zfi6H9jUfs
aMgJSaH3fZEuU16xLkNVn68oEvLCz4MCUX8lnbOwnjlQlf9S8NLNtfKVXs2pXA3yStudxonFo5xc
SVRBpw7IK/o7Ky75OdXEjeh6DYUjW4+zDchRSvPMZYhhUdj2HVDeTHkxpGJBQ6MLuRwLEu1lg8dD
VGkM3UPznmyPEVHnGSodTTrGvOnD+eXS7W/OHHhXjAjf6V9Ia6i0tIEMMBT5rseZznh7IzIAanUy
j8u2/oCIhhSxI0JyNqE/h0eEFp2PPL61SaIq/LIDSB26lzBIyGVUgaeCPRuj5MAcIBo0ZqdDGmbX
FzWV/1M2NZLjOJEAgwjoeCIZqu/mb0OKQJ3x3Ywn+4PPLEnapBcBcSbPSmpsmjViyhYedGmi2+mZ
c3QMEyo7Xh9X4o0RXbCVC0ZvDpfx005pTWhdJaqP6cuN780eBYUN2Rbb3/PscMVgAPiQTUsOD7gY
U87EzDQfd1LNUaqs+YvBih1U9n3lcaMH6+D/dZTRZIWxB6Lyw46LYN8xhbswC8u1+ua5H8S9LlVL
rLHEGB4bBKa05Y7RnWTc5jqwC35+q4TwHJsbkyn2eQrH5MGC757fr9n5UCm+OB6MFbu1aRfE2LnN
ddRkcNKNOdQ++Mso33+n/Ne2Bd/9Rj0RWSyYfsbb93sE6/r8sBnfck2zlR2AytModYjrwhZsUBnP
hvan1GYzQGJmsRaCxpGRi6g3XAGPyhJ+7fmwHW7eTUjYii37vElb0AmOHLIi9L5fTDcNz44n3ZQ2
UKeRKlEDg5IiL4AWzOmtsIg7YahyDWkJwGOd/T0uEAgK5i4LtN6ENgLwBoVRUiYYQAV/YJqsj9+2
yGXnk/15P2X8NoGH6+H1DEQq8UrHKeGzDg+xC93Z9celEsplWUHllImjfil7RuAHiDtQ9p/kebh8
CBlPPkdnHvdfcmHFt/3XtzfDC/zPJhldIhJK3ZG2EqZGdkuVZ6EkjwoTxkBeJoFd6etPgMPJjfVJ
pBfbRDnXF/4QUKJY6a3sLMiW87wTQY6x+aifq5UIZJ9gQH595Lfl9i6VuCwzLufF69Ns5wzjwjhH
51jTMkz/wUmyTkuy0vjZYzfhjuua3T7B+DrsFsn4JDV6w4dVF21uh6VgLAowdXtB8jZmAQ4kFy57
nnXcf43KF3iRRNR6emWo+al4anX7RuzkJoew29vb6CxGmiekyvYUJ9D9rRPU/UIwcSp2MgUrLyY2
GlhGvUT/wtAA8H7XYncvSyBcnbzAymtLitTg/KPJc/2/a5NRhxfbJizEBl6CD7tofPGkck3f3i0q
AOaQdNpfX9iUQV56BqJmMEmoMpTNG8442NS27oHT/3QdNKoSVq4p/c0TXO6AZpTSxkrm2/4AFT9L
DisFDijwEt9cwuqUb4k3EyNg3h9YU8hqour42t5xCy10opd7TYEDwq6fp4z1grbRq97G0c5lZFH2
gZMzoiFl1dILqDWxpiib1bl9UV1GqV/jU/w0NJuDHuQZNUDFp07g9GL8HtuIehkTdPdiSiKlXPFX
Tvdh96sH6dOw1E6aOL3PlEZWCpgmBAKG51ZrNi58qzrDxfYrOQZuBgFWhXxHfqhSlCGscnX57IfZ
teBEg9ZG77qCcLTXeZ20aNDjxb6/8DYtLDrYM+ZT+vV2IP0yny19wnqvkxHOMV5UHTKWBhnb6ZTX
r1VxXXTeW40rtUEAP8zPxYn213gOt++PhqH1noy/3WUeuqgBiw3RvO+iyoGd6g+km/Wdy8snLwak
T0HQv8MtKJlQtr/9ro0vb6lzEd7pnrREdoagpI8zA4YhJz07YG7ALsM55B1qF+rSzx5Y7F/zbfi4
6k3QIe801qxY5SIhKE2DasGZIoTxDN417FHovJprbZQFO1t0dwW5sp0/J2P0wKOzgiO/JB36kDC/
vBAg+EfJlp7ivX/S9gNh4b0jqWeQ8MGZXds5KKGOzqUxCmIT08sMXRhGUOeTQv7B+2N//H63XZUW
x9P1NoBJNXb81pjt5qDXWoxI3nyxoMVTqS+pcRQsF47yTdK3z5QhkqRWKnB0jW9L3twgbccF1Dzs
0XsH2zozyOhvvr06cLHXo27+dAnlDkAiwYiJqSkU9GUJFwfuIMjU0UKik4AyFweNhUAHqD6No8Sx
6JrhiCJACUiRvEHmKKIX37V0sPaHQwUexQcxY2zNjFe0Y60rJRsuP1pWfxC+jqCrVESzlvNwNE4b
HXdMg39PJxNQqkeGrxyI+HxG0/Jlz60VxduZlWnZ/j8yPqNePAzSPHoaqN4zBnTBPTixHETdBhNZ
gZ734omRMOy2bmif6RO5zYnKYIO/mMUMkGP+5+CW5zxmBnYwxdC89G6NJfkzJia9fKV3Tmyq/bFG
gurV/a2IoD8oxQ+Yt0gdcG/tyLYVqgA4SrwkODhb3geThsT+7bb6yz6afv2seCQKDzifXMSupgRY
X6tWNB9XbpQRBCN9Qb6LwcAUGK7F7BoXxxzYnZRKBRd3lBpHIltcIqMfL0X22ISTEmOX3AHbjAAh
jFgMDkMdtUueL8ViWvwziR2nQO8kqY7N/pG1ceT40JsiSlHgG6Q+9toWmb54yBai7LB9ENiFcEGQ
UKAAkuamMcmUyRO1abWJvZumE6OA7Oio2HczNcIIsPYCiPKGLJDIeAr4r2Dh9Mbsz/KJ/3EjYE9s
dGlYQOClY2DtwZDacvYM1di/9KzBUnpPjoSsfAXUNIhrB61VUrDRU8zK1UOrf98zFNYJaDnsEcf0
rTcAy/zWxw4+7lg8iLFHxo+qAcdcydIqFFgwTOgg9Fv2BRSLFo/mlBPndPz9novuXRCcBjBU+jTO
al9WplBC5xk5oTxL3R/EBeui5uXSrkaP9WAn2c9XmJUIpZc5/5MSfPj7KairU9UdSK2QupH8KJD6
7InAxlnfYPcUbftH0egE/u+EmKxfWwNQHVbiRyWpG9RbNfisiqDVRu8j4oxcqaQqxMLDic7HPHFY
dxFUCm/SkLVKcPkbTL27Mt+c+N+TTdWvrQzbuvZ+2ZIM379zMl+Wzm2opmaBAiMdNV3vNAQGsM4i
jr0cexqrjzNpJTnZ/BnAgnsn9yMTP5FHiB/yxqIEOsqLTJ47zW4ZrmqSyU7FpxwO3J93FZ/At3rt
Q6DZJWu2ELWPFBip87FEPzgETKAoimuVx+y7/QuJ8EDmRxD6Jmbz5QltkT/4igH41WzKIX0TrZ4h
QjQOfsN/x6yXDud56wBfu5w3ItGg33mPt2dKJWaAqR8dkx42lj3GD/jiTlg6Nqlk11k15l6OoMme
KzdXZiicq59D0UGSI/ZrC+pv/kM17/svicxK5b1/rq88QTMSyAA40Mc+pUMZ5cmy7MqfE8S9bZZx
maRTue8lToG50C1n5gD69Cc13j2gjols1ZyASbKtA8VmVJ5kveV8v/AsOFyKizsFESms0VK9dYVy
TylE0iqsjwyBAfRAvNNOnuzhA3qBPyrVFwwrKFPpt9LYC2/yeepFfYIGgLI/IpzMut16qgl1Idj7
duB5LtUvz+hD7VSogccrtvM8pLVQ7cv59lY3TUIjcFM/NP3lm9OhiFpYFM20LjgdIuYubwRffjOM
9Ws0XO6cg51N0RIEm3t8tcNICDOQCWfwBysvbNvOazUJUgHR1Qftnsdl4LJpyuuWNvmw5T08hSfc
rEYPLjoZ2FaG1NNe1xta0CgcF7AovH31Mpyv3rJnWrL7OOP+q/0U/qG3L+pstMqSFsx6kRY3d9kc
7OrKxcqQLwYm6dlKOJkwUYoJ6NSHW9a+GINVe136+V0+TAnYqLqAhZPfvI2+9uCcYWibBdC7ITpD
KelRs952lI5Z8KdmvKBo4Cl0VcIhvYJhA8yl3mq8hwtsbaVD4MjQ1dmL1GO/4dNQf88EZnqfl7XA
sihMioehb41TlfWioXg0paJ8fFAqJfZrhWrCGzUAJpjnlxtH0GCzTaxE9yD0GwqmcHVzy4hBajbH
4LwLxDK6rN1qV5MhkjDi3Lii8oHPn/yiTSVL3j7ZExWklLeDcPl/+t5zQ44NXnAygPUjA93s5QcR
KSC4v1QSdoWX7ktYWi6yKETKuaCaCBLFZ9NXvKB3Vtd7xyW9JKOdwHaDm05GABvBMXpdTHu32jjQ
VWBorf/xgSv4Cut7bFfmm9xHh4ZpihcKvqgUhOBedhDNMKTHWKhIjuQ9HRmrCrzOYJ00JLZigt3R
3XgHqEnMv6Wgc98n+Gpy5XMsIDt3foHCBFIrQVRWao0sikSwk7GmOREhUkOUQv+CBiIWi4hQXAbM
ZJmezjzPfkbfNyI94CcvpqbWias2dI3a89BEZzbDix7RZ73Vowk76Om7EoepWXbldeDAtqMMIDwB
LQ1Sjd/yNeTjZim5+NoeguBj6yBrGIqZkdGEZ8qiR+2JYZ9UnrCVXt9+dAymFWZDmOA0+92Do4R7
ivULVfOPGxtxbNox2k0KE9CKv/FjsZwuVbr1xLKDLs5mMIYra/vA/CVgTYccqhiWbAcf7GdkXGAu
fWDWmcAPIfO470LWgQ1DxQJlZK9P4f2yk6mXsXv4x8AYDAhePVzyPlD+6oPi/Kk5822eW40FJjP5
kvN0Ghrp2nmOdrK8A4QwQQxZK0AlH6wAZNQbuNJJlNxapBIcwpAAhpIKulPpuqwuOxgLvLG8aWTh
Fh6yhIjbq0AKcNpfsvTfO7gdvI+uGgBbt6UWiIAH2CX5j7aoBSbd+aWqNMQ7ancBUMIkMU9DtDVv
Jl7r47NfwHcUb8qO+hkgBduM9p1wM1C6KQ/Xr7OZJBgI3NEWXcVP2V9C845v93GFxqkgET56TBP8
CYUCUdaGloa9h4yQyWh9BnBGkqmhZ0OGDw9EPUTsvJ00Y/mcrZ69A4EtaBSS6wOX+D8UiCQexIPI
IZXJ/QhPQ64g+Ekdwb8kcNQiY42nKS3phGccLdG3zQ7ETaeJkxTzfC4QoaOZRbpMA5RDpNxCXW5s
azGCPnsp19ZP0wcM2D7LquI2dEZlhbDUDtYMIIXHHyjVAi5kUXb/JkOjgiEin6OGaJYkxoKI9d2J
EDHCi+QFR6/p3IP/wfRaha3zJWILbJHlT6G/kVEqeZ5HLrPiH6Lgm4d9u7q2rHzng7/IKuFqywAL
hijL93ZY84sH9JAIrW00DGzSNNxnoaE8eSbVCNtAjCiPuGKeppzEYp2P3VO58HxDmwvBGr7Dpt7y
/kQc7YCDMXEsiFZZIPqVSf1lgCDaJnKq3SmUlvQyktMHznKN7GdhuFdTG3awSPbJe401JgN4ZD92
1ZxOuhZpvBxxEMANP/9qduWldHn4B6p6TD3SyUXG94w1hTK7a2hQS9Kzhh5mdaUUdkvRYv0W1PH3
BZDl7zmpPvbfSr9GC0k39iv5lXYgWCFvR/KrPZqg+ZyeDE/s8Zj26BXf7f+qanR7R5WXf70Zirys
ljRVOEBdRXc6bCyEcXpPCbCgqN9donKs7HQAVWJMKr7TXr01zDLRCOYGjJMqisfHrxgEbvaNipE0
vmuwX+58jcDb55vF9GuwFvDMU7175/ldypdCN6ZskdNSW/wmeRgWpR2c1AKAKVu7lg2S2E5LefNX
YtzbrIWeVm0telN+SLvUotOyxB02dlRhgT21ubjwZ0fYA2IL30fO414dggaqSzjEqNylP3+f9FL9
nchTy5TlzJuX115aPz2x8vLmWrFMbIQioSyJrQ6CmnC33KOmkdjNJXrAfH8zWmKRGDEThDd4M1tM
wSpPDfAG8LXkMyKsUZwG9jk+SnRWawcnvYJ6rOLEiz2zVz8VR4SbgyZ0kMR9ZtY5Y41M8RIWbQ8W
nIoFI+afP7OqJYr3ISYERAk17CeZp8br5VB2Y/My+ljQNqANfjtrY36ZK0PZ8x/A3O0rFpLET9fV
Bkcgc5yINYsgc6O9LfJe/BVBloxVAo2NweEv1AGXX4SrVQzr+wO2bm/XsBvP2q8txE52/zYqZwte
zROgpNaVrQ4Y3ED+37H3EdORbJaNh4CaSgp1Uecec7YIWinMQ4fW8C+M/Tju1WTn698VjJp/XUXH
cP05AlMuPL+n1dEbinj2NCRAGb72Khtp22qMWMNC9M20n7w0ECHUoeLbGfGpoqBDn7cUIaHXFClC
y+3KR9rpIqwIakfD3p+M1ecBsyL1LUFQOzLvQvJhUt93yWVqcot1oP19AWgg0mCc+vP63inEIy0F
OcD4BNFhYHHYU2nV4s/0cJPJdPFkx+eHUj4XKO19fdnfdMj37f5IQGkoMIfe4aHQzmw/IjgA87ck
9I3m854FyYorJFt+5vEoGg2Y25X9R2IN3kl562A/KmEinFZZndV6NlIQTOW484erQIrEllQOVb41
JSNfpkA/y0vSGsfwdFHALYz6oKiR4LVhlDNeOl2eZETmqph6F7uw54x60Q9R9Sb5Pe6s9tsMLolq
nv2tLk3nWYdHCNNvdxioElRNtebdIba2pQmNclcIM+pnVw9dZvVCAZZBwLQAvmNzfbjLS+S7pyZ3
vXBhOHE/umjUvjXDnNFXOSCLdjPqU0rCfvSxPCVSJHNmqdoDIPT4c3YbYX4K1A2uqhr7I16UdeEY
yv9hDkI40SKbEe8+463MqsXMfZu1wIGzHW2LGhTES+Gcpo47jI1yI598MBKNcr69bpVt3JIgb1SD
m+GU/OZj8+K5UoH52azgC8MqdFmqr0CKbVvgOhWzCFiIpKOtFfTxa5SHOS5mNmTl5wElSCD6z2HN
ndU1QesBclfuKZ5alO5ePdH2GauF6zjPtEXzAbwWPeESq2TTANzLD0JSFf/BIxPSBsOISNwoo2Eo
P8tX50bqKS5LNvwK6jJ8PC+oHfUyoc5TkGQoLT/4KX6HB7VQTTuNnLIzpcEg6coU7+E5bsrtmG2p
KJXQ/VEH5Hg0zvubo5sl4qwmadsZcZWIGFtO3u7yBFxJ+nLv6GcQ10tWTAQLKsLlbHy7peSoQRD/
jSwtFYYDBSYNrKz36bUkqB4hgsVrRSm4DEy1iXlDmsTGgyTpJNvvvHyjOQumxuLz8RtRxe8t/+JH
na/+5n1/nPMhUv8qMXfjblZcr7RahwBZBifGerRsDwhY3+WKSBzNCbCgP3NAK0gkSXrsi3ZMaLtz
wx6OhaFYbRf6cpAGHiby59VW9KbNl7T/blWEr9GZIUGTcVBF93DvdzQU0vjkJneft/W6NWjpsM4R
QrMOXAdfSr4HN2K64Oaz8WwiPotB1/uDvmMk1ECummBiqBcEO4RB71uY8Dui4Dv/ZnCb0t9uAL/i
Y3zSXEDk5tWlaDR7GRuA2AcPzWCj0jZEMRmtj+O+wXk+f9ARExKbapdk2jdA/e+W6DDhBS5skTne
juH6bUL38u3orKj5WvbWbFkP4UkTKD73Jd7uc6wMSSeEP79aqg2xFTbycQAVSL150/9G8al9CZBm
F7oHzCPvSRl96n2N+jz2yGduZQ4HTzM/VKxtifAV7x2RuXYY52L0YVgnN0I2+a9mSoHUGvl/jFMv
h6IsCeD3vUcjHSpr/5sWnZEEx0yba3cITzAQ132ckyYLEt2nKZV3CR9yr7HUYQYSMoJUQJLVjm07
k/57BT5sEudNI/28JfYsl1PQEFUngTw9hWanBWOAOp1qxvnFaWV1ha57OWHph7cOg79peBVrH+V1
LfIN2x8b07DV66cKzcEM0FJLokEI7JGyLJSdBUFIoTuGCz0ITal8/GnZXj6gS0A/liHwhQUfzHm/
uKLXodznxpIJMDu4XCvpKj5sy5khrJgVhFBfBkU6rMpjyn1l9UTZRuBfm2qJGUX3/UhgIDerdWo7
vNiaUwfHGnc1OkmMM67PDGvp8VcN4O9+dwYMpYHep4HlsLgk1ZJOHkVUQ3blwI/4vNfoi6MbksH0
yOOQRhuDBbhOfmisf+mKgzH5cClrHDLILo490l+HAEBwQJMv0Mopk0RQAxC9JKUMlu0PHOn5hyVO
lXsZTe2V5lj1dwndru4G5PsstfoNQ+UjdSY8P80aCxYbiGtF/Y6lfJhr1YmBq+FEl/st13U7ijg3
JRLSs4QMTbC5y3rsAdqZC6h6FEBocCEH6vJhjkrSNaTcP7mIM9hUBAqEdXbsqVHyo34a3E5atRcg
ezNFVW5Nr8M/VsWV2azqtp5q9cIYuXrJ10mGBMlURqbZf4PQKhWQ9G0B3830//KkyYz8Ca3kaSuf
Bh8FmIoLgc5y14xeADqrB8YICuwHvvOQJqvA1lyx1hLu00doxFvQEUGBI/GtwoDpbmb1R+Z1nR7o
3d7QM/AFxwHDCFwJiPVMm04v00WBYjbXUqulkmzazjNGXDnOfOBelZB/6Z31lisqSalLImQ4FVmL
RooOKTPstMxOwvk+rZcSrt3Da2TPPFAitAUELA8BGHFluu0629CMS4yAiL+Bi8GVRid/Fo+VjBrv
nz84NTC7fpT9CC9urvuJbfPfq6Dhu8BIkKbxUSSIHQTFowULcBE0+e16OXeK6l31a7VNeYmPZuWB
ijNOr1deJDfVKlsMSL0nLTi62mPDmdhepz/GCsxeq/QXl8o3Lq6WJSJH5AwUz+DsiW33Rg1E0xUC
q3AfsqncvolO7EepFMxJkenTXht20YA3wVkUTrrVab4fV3jm/MaMUcd+gm6NxOGDkXyPuMPwVGfn
gwsI3y1ipkYCjF4ck5jpeWz+HtsYfMsIM6cBLKGIx5a3eRFdsUzgJpbOdSM2MPaWpwSLVrQREX8i
Upkof6f8jRXXWlHDpeHu0DObJ6S7yrYElAH0/4wfgZSuidn7prCeZw2b6Pp3XFF85mDHKRijLSA+
Ij0PJKrHl5xT/ERnTjOkkfI3xa4qlwYlnazcl3q9YXy5csg4tFzu0GGi7nK49J/jiCiApGKmQUKW
x5LB35wajGcVYTChqOlH7mmcnlHJ61lf3LXJ2/LRuj9gljbUGSw38SX1E8BhuHLFkD/1FDfCCqeJ
X4V/elkhChLUspLr4B2l1MRnEBVgWonQONAh5MJ0+ixuyTEtc/YDTCtun1JpmkTIzj+kZGu0K+MT
S4oKY6rQ0aQvXPCEm/CPuO65sxWueibS67WrvJOS6AhsL1husOFTJ5LB+72ao0LaKTjjY4MGfzO4
P6ajVqOkh/QWg0U2tSNGj93CGofJt6vnRIkhmqItviZbFHi5nT0/GIKk3uxnnXkVVB4doHGFmgNs
Yvv3IFUbY7EEnBgfmWj018lkBzQs2hRxHKpvKtpTFf9v+wq6ktZQ8qBcB8hBeIww/Eze48fH2fMu
TLe3ZEpksuP0R8ptMchNBRDzqQV7udzzjbGStsFGH0BoxyjVShqqrk1Dek5YL+qkaMrTJSHJgwp/
v5HyOwhjJd6quMnIsTOdlNHrzoQ+6u9YFTLxzlVLSKvT798jFBUFaI7IZbTUCdeCQx4wUfjn4Mbx
E5GmW0L+/LEtRDYlkwBW0lAjdrlUYtDtuFOjhspBizfTSfGpw9kKDdsGMXvDsM22bGgGScO9j2R8
jLtr4oXZ9P0qbY3yRjP4+DREWbfvNUnPUbGyPilXJaj2l+bdbdvF/m4zmG1I64HlURomYyQ7kWhs
cC3C7pPsj0EFxne6eE4T8t/i4gvcThAfKKa/XVk8f2HPXw17kbpXYPArFaxOVLFvw9tpPxYMeoF3
regDs7h2cs5mur6joJzis/k55gxMUkH4fSLeAE1BHkh01E3QxGAoooLmSUXg55OOGrVg9iRJcqTY
EpR6hCS5qQcMSeh/bmtcB32bbafMm9dFhcjK61aW7BgJ+DCkXTVscVeAGNqtoVRbh6Wa14ffG2+O
W1ML7yaZwUx8kIjxDULyRaIlP1BYL03Wb6sK8u0XcNYJMkgJuZPgLG8Kmo4anpu2c37G51J2RGDp
nYi7XULaedj58/hAS/v5KnTYtDasrfy0E/wVBSZQH4BWkg3oXnn7CFWZ0Ju6OloXwRKv5cyaqNbJ
JXAdAZnrLyYE5GhHA+bX18W9PW+1qajfX6GE8er6IgM4bYTc7oAzEITC545xDNtlMGGx4K4d+VOS
p8whHCcQt3loB0EjaqztoWaVAzQWtjDXyeQlZ9XqxYJqGF9rBKwQKHzH/JudMCOfIBYrtx6xq/ui
6WBLN5FDFw6O2ZeAgQQ7u2zwjYyLvZ4cyl0U3Yb8wBMD6xhYR7HB0W2H+17mcDKlnDKODQnZj4fn
C6ikNHgsqWmxRdk95GEkjhJSo06aGAbddv9/PGAV3E4ww52Do2k7aLpS2w0s44FWH0nIVvB1U5iv
29tohgMlJCcF17hOB68+f6tRGXePVqVe1+X8uRQrNP14DOIk13fjiMf31GNgPmxX9MScFKY/Qoin
Pif0M4wlq0wwfgiCcTUJlTzUex7wjpyQiuaCJc5h9BdIIFhoxjDcvZHhDRidKA417TMWQ8Ye8nws
qF9KomKB09n3OVk/ydnr5QCWvh8e1P63eJEZC+PZgzbPvgCjDLVAmUbqNnUCcVY+wH0n/BnRIgxq
/N0z/IXa0sX1twdJSr8dafJ8Pu9v5U2uqtQwJCtU8JOUQSrfE/mQ2xVW6cDavITiJLnuG788kVAw
izuKxL6Gh5RRYE9KhxG57UPeS0LaXS7aG5B8hzIrHyxK37pb2Kq0xzB1/Z+os2bqmq3KoNiDw8is
0ekhBw+8hf5XuTDQOgdx8xdHv8dfN+6du6RFmByXyz6RZX3wPrEAnTFF7HtpVfXBfhAOfWq9z5iQ
Zbc60CJ4yfZ9Xtxvj18L0tHrGNMY6lEtHT24u0D0wNF0WqqNyohgUVqx6u4srP6HBa096bxEXDCQ
cEbOH1oB2W9iNZPLOiwzKE1Ut5QgIXbdarPuiUH3/aTPcPRbZrHHVBg1qQbanykcYCoovWrLV0ma
iMfyIIkfSdTZA/Rplia/klJonN9/p5yfcEsTNYcDMZAUoEGJ+yX9UHJZceSbklvYCP2Qju9LPMCC
p/QdgZSPxXJGpYSZqCrdXGoNzbynC+GKPoHttjM7Gf1BhIZi4og51G7w0ZtI8kaJtShxnFP4iHTp
nwFeY8PGJ0ZwmBzokU8hY37/2uPYv3yqBARoIeFT+EvKTGVe1pCzIWoxb80vnLB/Mdjz6VWo7iQx
rIC4ryX37UFgWmXIp5bP6bl0woHmml1D+TyvNKBZsm9lVZPgFMyTV+ZEakqrHWoOPLrrODqMj3Sx
DRiVmwC6au7l50hDeDuHTSrvrDcTvC5b4jdlCES7ZXI8Pqc16b+ogx7PulGUs8rMMiPlB+9jtdYl
lxloFlLP6n0GTun4mW+eWYn7PqcpJt3eAbTjZ6J19o8PRL5O1abZIwJO3Fl2gWGvXT0EVOXiK2WW
/gxXtDb2RSnbDmDEhXn4/+ftc+pymBsdC0T+fPFysTIAP3isJh93WCkWoeia3Lc/YGEnwDNI804v
orXjW2xGEGtLKkxKAt3rk4kHD/DmxM5knPj28Rms6RbXGLwKVLGIBIfxBNnpFLhBJg01IYTQknqb
sLPk4+b8QiygTRyNQwBN1qnbYbmflhNrKdpgO3W32/FDiIjwHnUTP8HWRV+Q6Jsljirv0MGfS1k9
YqAE0D0Z8sjLI1TxkXMYrroDSE8rW12QircfDl7uRMXMOn0VxQ/fTxjSQQ1K+eXZRp9BwkEsoR5X
Dkskkh0Rr0q/4C2IzZpsY6HAvn2Qoz6n8TXt4h6PYZsH5W572en1bt/PZYwb9LgKRrntb9WcvglX
RqLLKzGu8HScc6wv1IlZH1Nk4CVkO7R37+5Ua9DM8bsJ0RLstg1ATF3vvZT1HTKdJHP0J6Rrow4m
u0kzilsqQXaSfYJpzWnTCvLeqsuhCK5CH52YkKtU1fhdB+ZMTwlM+Q6sUiacBom0Mt/W72MZMYcC
oTCFTilHU9dOlQSIKnGyXWB1zlUQNUgAUkCeAVGRoGO2pdmuuAGfP4uFypiLU2xhz4fOze59fGlu
6WLvI1MSkH5y76uhIGPdwOBoG/YKYuojn7VClfzSIiFDfesHjq44edyDVhABurDFrEEL38FjNvb4
n79PJijl20Wnrd+ylUBhOf6FZ+gnsjvcjELkBUAXPZzBwnvjzRpBkw42UWGr+LUkTWdIjq8Zsgba
YfShGco6pHWgC7v9sdeaIXseYoIcdPTc4Ct6GB5YnKTQA1OdWDKLIbxktS7Smr6x5FUEoZqA4rTj
yZbz+UgX26c0jOuqDwZsGVbkdAJjkbbekB9UirkdRKmTMlqOYQj26IF8ORt8k78ZB+DoICXQ7K75
buUpcF4dJYmT7dOQPNfMEnn13fRgz1yJOcWYMpzhmIhou3KVEBzhJt/2x4TlSdYqPhUKYsMJNgUp
4Z/RY/VihNCn6SzCWIibZGGsgtTWgA4ufpXf1f0TqSRWu84U91SVjMZrS6xVU4RAvXg4jruMMAY9
VAkDxror9ScLdmYS8bwXJSSn9xQajmffvRmo8ocNq56TNf6YLw+cOA33dY3NBdfTK6Xwh/92TMP/
kIcU4HewNo92TylaRV59/kSY5sVT5AwFkNV0aHiP/o7dXTVWlisFQ3fJr3cnJFt/EkNgiBeUBhSO
j2S1S3z7Gl499BV+X7voF1faPRQCJG/J3XIeYOnTDV2dODvzn3seP8IwMWV8TZ+chU7nWfNgihom
zcqsfvmQH+c4DJsKolP/v0x8sdcvsVgLzK5P1w3X+2PhUC1WeXcz+NiDIzz6jC8yKruBBx1PLNAn
DEW4B2G8yHUw7/sGWXF3lkDsFH1HXUTeQeap/PELc4necWTMMpbxdm9BOYjeze4dwSVSnpElXFqV
OYc5ZtZq6HxZaOzSIXY3iXMiVCmOKJW9B1YxuZOTpGi6bc3/FRnuW4v0LLoajBJ3rXGY0sJz6KJP
7PZ4sQ+Eczr8WUTPxnlcuarPyXe4RXcjYhTBV/ghuEN/bjPxRQ6mqiBzH0WvUYpEFvmvJGG8U3RR
ZDfYniWYUQZWEC8PvPpPBBDEZ7TWZzmZ+zaU4Diu/wapn3p+HiQqVB2z7kbVmBZm5L3Ug5fcTI+R
DkFExM28FanX/L76n8WitBdDybZIaJcxYWNqfxfng2V+svj9uGgbE51Uh0l+zZJZUJYK/I5LYVYF
JyNj/ogN0tT5CXGQHLmR22KiZfIDshJQkJga6zYeM7SqeMQaIZjzZRWdHlNvXchYu50fHbDWa66R
GcmWbZUSX/7TTpseSeF2lJUqRiw3mtd03kY7laqfoQfIeeuMc42MlwD1L7UVHTgSmK6PCi7IPJI5
SGpQEe/Tmf/tzmD05nA4y9kCA41RzVmwWrvgGR3f/8pIee9OFRVNsIsqrTHqfZ1+nj/uGq8bTYv0
N9sE2HDfBFlE1msX5SL0CnF2KNiOtTf6MV7uYt7fi1Ay/VjRSpx7qDZt+f+5rgqrhIGZP/s+qvxO
v0d5uTqDJXpKeX9idflOAYd/8KJ9o6cW35NYo3DtrUK2vfuetjcMyLMJ/Mtna8V5hnk4ruiATh/5
obiai61OXtbCbxX1WhAsld5MtRD5HLPXruOuPZQfl2pFKMwck85txNxNBLlAJwS+73btamx/BqHp
O3cIB5wrLc62K9MCtOkthzDMU1REATZKQCRS4OTMdeZMpa61gru0qEuBLyf+o9V2FZ2BID7mjig1
PUfUZUeC/iJ2N4G54JMIBCdLBVS1yvH6sK89I6MbooSBYkSQVNbl91ymylqJlGUU1+w44xQK5eDU
N07hxTQE1ho3GPo26GetNCUgVJp1ljqWT7wPnV/Tx0d76REFkn1nbzFYGj0mVDBgPLOCYFXJQtQJ
zu+SFVK8ovmr2Suj+LCPsZr29YHunKAl8InlZuvS/AJzpMVK15xjCWrA4zPm5jGGwd2cPXZXa3ei
/wfalNSnqRxcAaJ+N2fjbnKjp8gdtfUqjBNzQqkEI0fQnFzvGlVCDO2y0C0d2pgq46sUCCwzrmOb
HysP22gkiXINDp6jUowGu+FSmxcMM69PqPNO++DbPWNBjoYfVnHn/F5GnAJ5hH7cgbATo3/cX0Zq
y4hkgulxxXbz/tmH351n749TBV3d7Vq7/j+5kAlnCLr6wgERY5qbo4I3FEuiJ4jO8MKTJRJsaapu
n9p7lnmUpTWW8C63uMmL9IZ2kKwfT3kUirg8T4R8LGCQdPs4RxohkNKMJDd3fYMWtAUU+/PALI7x
eNoofaNNCSJ6d64EDX6BSs24NSZkNAOAMHaf20NMQvfV8zsrRlHsi4LEpbnTrmBh4pkFQ//foiiZ
vvDbIFgjS+mj6sAPi0WRQHHBZjlPWhlHeYcM5GlsuUCMFLDroFBQzL7whn49cTkOUU35wR9zrh75
B2biezdAuQ/NUXEeORxebdO9rqCYQg9quNR4qG9Sw0GPCY7ZCyTh+G6dTYvQ/HghZyBiOef8JgQD
NnJPETW71w2nNhg7YlqrCggDryYVdagdDRiBmM9++XrZiOHU3q+EMKWSBQpVAQjUizOToGCKJ2z1
Cv2DC1rbvV0KcAvglE+j6WAgucvOlZKWILQMo21XX1uLuOumBJsi0mhdCBv8zOidnPGRiNyxocna
mSW4UBK+0Rn+k2nrKF+GQeAX81SmLdyzCRgv4S+EG4ixtQmeNEyFfpOjRW9cAmfCfXUeIp060/B6
A1LS6xQX0xCAauyTc/48hwxWegxOyiWrrZhRjbmbqbODx6hag8nz/SjF8j/8Q8x3EyjTihVBNLRU
6F04DgPDi0mIrHexvAnIxEo7xumZ8F6heF5eTeNjK0urquosFj8osIBsiyC435BV7/duLx3DueQ2
DzzyV04oZxODRse6YTYqceTeCbFntpNQPPxxinKisNYTH0FFkrlf/7rmvnShWyx8ZSTClvjfZOpz
14oKv5TyLhWSufb16qlp5a/YDXKkYp/aI+OzXQAnFH5hMX3/dV0NAwo1L+hnUjH+sTzFTz/Mb5QD
3EPYSOkfBDlvikIolRtfbm3h+LFhb28/KXFONCjp1fSX+c3IrRa4w/Fvc1nmWKJrvCtkoBUHAiur
QAdo7WBxojZjMi3fsGLOsfARJZXfC3i1lDcqUXmNv4NNpkEoTM1o/cTjv/VCjGKrE+1S7pPO3QLG
b/IBjKl6IqwdK0x728z8HWujav24EXpNGxU3kKOIeFLnw6ubqu987yZAG4aGA37iox2sc9/toh3X
3QAxwoU9C8pTX7T8q0nchRw1ihHj4/kdj0ypz+4EHdXybx+0jm8llKE0xh9TOzMygcP6SsCK6l2i
3snAjjbFugBEyuAxw4qw9XxqTsfY2MLYODTM5tpjvJqeOwtz1rYnKuZPY4x889obOMbMBep6P3Zm
t6BgAMPAg1givZ/FxrgNY9zio6jkT1qCRMdfdRZBA/qE6UStQeYAxNSH7/iwjX2H+or//5AbWsd7
V/KwWEb7iq/x0s7CTt1iBwnJa7xjzg8SZxjKRzqUY5AT/WKffakJCIUOUKKwQP47QWl6Pmo7Nkh4
3Bmk14FIcDqrWvTVTdSNpIKwVjqgub+KN3WArqoDKXO+cBVv4AeUjTgX97O9scIxCanYggd+xsHH
k9gSlHh/Kyww3iUcIajRsHKYZGWDqT6mAL8fNErGVOZPy2gs3AwljaLQKLCh53TPGyMnpomXvv1S
VKCT4yWb0mSQdXhRwVIsLjRtYf20h/GVYe9iV1L4nq7kutXgtgc2dLWZmVeSdzLwqHbPQYjzB4Cu
f173OA6hwlGIxJh4a5i2jbrPFDNomWI+YYPp0r+rTB/+pTaAcH0XOpdXN3282sLcaIQaGNf4EnZB
e0tyl0Fb9EO12Uj698JJOuL+3yKt+rVv5SraPjlt43HM2dMwy/KCUMbvjcyxA15fuRg8Cc0n1MFE
mGq0fUsfMmGL2GCp5IB0sCSMPqq7UlXxgwcf9uXBXIp+OjX3lhAYR9eOwcgI/6L9PsSGqaPf8c3C
0xGABaz+LYBbGG2xO9jsXg7DTZXc1JjAt+sYJyYBwJhuytYeOw1mgXcx9gD4HEt6Zz+mkYawKMsa
J1PXZLv4VJOdqBtHVuTJxOK9VaJfk70/xn8SO1NRL8C4u98q/d7HzvpeUSfd8XdT6uA8HZ/p1qL/
mCKVcxdn0smzWMkY6Lrg/yO/4XOUlAxo0XusFnR8fQNC8Q6tgsrjc7Yh28dKNuc1F9c5peM47d7k
JZ+puRNrbhoTtgixU+JGCRO1QKzOmMp79x8YyQZYEJIhD1GfqC6JSxunYZLKVU54lSi8ebcfBHBv
leCXjMAeGiMHVMwalLiiy+grtN9fCOOki2pQNbkyBzEv6CL7pY9/Egh0PI4dAD1zL0mZhfvvv+0a
Qc+ryDLMCs5OeGD0Y8EgnYNR0SHg4TCeRaYMIh7oLQ9PgGOjNMItL1EsulDhbFOdFckxYzKqvgGJ
RIPK8Y5C5NEMKtQvN1OL9uNO82LRxYxfC8FNHd1SOIk5l06W6xquYFFmzKrI4w6av3NDE+v0TjwY
0hwQnjMtlOp7eNhiGOhmSrDsGsytKYp8++Ihnq4uyOmmji3uiBichCyNsT/QyXvl//cVgBGLQ/h/
i87Y2fGI1+DqsFoszc7ddfdATiwlFJC76Bacogw7IKCPgJ3tttGZinM8rIbhjw44MHdf2Qp5ZGNN
Oi7fgrQe9L2TtVREqf5ERpm+Gm+G3gW+cY8k/WXIC9EeSUGJwf5Sv4Dvxu9dPi3YzMX/G5MB4KMY
kVyOmon3YzbKoU4poSmW6jarPN86Clv3ZphAjA1Q8i1A9xe4qaJvqH7QL3jO+4xP+edq6911HFtJ
0sw9LgU3XVWsW1e4g4fWZhzqp+dk03zw6z20ykCVhIRJaOYU/qYphwgPkxXXFhI3d1dTZ0QcHP+W
FQ/QtT/IrErm8jmMmRXMNHM8m4F74yWnuCNFfuFayWqaSTsclj3mXniNPag+eUFAPDVIHKTAexxM
Sl6NmxrZuo23UmvJIBFuS+loPK6m2deFhtJ25P99q7a1/0K2I/fggfLAkf7+EBUQD2A0w0HHiq8J
WM8x7fVbYlVCb8MRL+L5nF0Je5LXc5o+SBqCmfyoHtSt8tbiobQsmesA+LkomtIXjRhZoduBlpCl
KK00fSEOlxGa/eL/JGeajV8rzzfjc0RsOhNurnHzIgtRREpvxyDADsyQTS8itiueJZz0UmdEroFf
TutJNEkFBLKk4a4okbPSITea1thdUiPPOvD6T07DxRo7HlhzBOzj3tjUeku1t62IMITW8ghkPkcz
cSnKTc4sR/8VXcUwJDr5SkXUqCAAc7vw42DvA7u3GhlL44uNVE0KaKOSOtsRSKEfF254e7jsHNPu
xwxw4o7/VGf/PlCXFddynYuLE+5H++mAvbPOu354jDOBboHpS9W8PGFNHz0/QBfMw3EWQhU8QOol
ShOjkQxzWhZ14LuoWMZPkVHbxfF6hkDUxWuuSWkRV4vbjvOZseIEAWbCtIhX9oVKcLodScj7joE/
7Xaroqh5J2x9Vk9r13AfgYmZ0wUFH4xc2G26YPz9ewbD1iJuIl4tmbDCK9iT8f2tVPGBjievd8/9
Acfnm6LnKmI65vq1IdqctQMCszYQ2/tb433HJaKsM/GeZNEjSls5lcr9nshmrZFDLwheCW2gUhkx
bcBEsakTud+n+CgsAv7XXbWsqtd4b2EX/1i0rJZqZbR83gXJS5Mukr8mE3sQEMmzCuIEVvzsKnc7
up6e59iW1X1cr3b7z7f0fr79ku01vxyvkWJAUvmFdWShc8GvLbW17+bWVUZIUw3cUDZhvVHOxUFY
JdxIMzPvLDhV+7y0DskdylXXsvAVwFy3+zTgLcPK/YzSYudslJ78SczbD8spsMYZFwq/YfrspJpg
8u8ezJFYTjmjQElus/hhY0uXzDyjB5jUgXnrxYj4Fb+mt1p5IEYzsh+GEF+YPJ8CxzXm2OJFqKpE
GSCQt/ewNUBVCq2ZBv79Zhf5NWbfQQqlDh8sc2+oUl4UzggFf/zgb9p5bvia+oqO5DVN5D2UPhjE
iwNtTtv19bQy8zlJjGKMakSNpobOm3C8pM+n9aAo7S4KX+hP3yYkMDBocI3JRmOGv6bHmWrYTAS6
Wvkx+ui12zPx4gJP8DG4Ied2pUEB0HRzIxEkKF4V3IwDWWa/DVk1en+l2TtfFqDj5SbhKMV7b/Ku
iAtsCI7Z3HoaX5SmLQ7jnfpQ6cbHOSzvKMK3eC+VIEbMxz5UWV17tQ01nxRI1+pkMLirbzLrP7S+
klgXIpEspvmzKpuwCPSRvR2q7+ejCo9qd2eQNnR/+wiMAt0xBsKq9ccX3aIvwuBfgLHmxcEbLKN2
fC1ha8DPKBRejGd2rHW9RYaWyG8NbNlujlNvd4X0ijqEpUl3brwQc/wdN479JLcgO/o1n9qxdoTu
rFGkRSSmIQ9ZfoTJT0cBHuep9/stfcU72HaUCfy5/Syok3EBSha08p7aEKuDSVhjuPXuPvNmMlLE
BWvhwmdquX8SBbs2mUVQANEVCaAnwdkNLjOCzn5SD/d0Kjmasaz8AkU+g1IA0aWg52DzsttNeSBW
0YZnmaNr/twk6yw8pg5gBBrxRPruceCOU9Vw8tgionEeNIsIz7G91d4CER2XX8xpNFpXXYguDw2h
AGdRz5kpYezLBiX1QHB2G6MwwEIUVRH5DM18ZVRa7GTNud+/7A3tDMIgYEtlvNMjxHvDQO28VTYn
sTwX3ot4xzdRxb+il5/OLyU4bkj3PiIDCOnCmH9X7mtlimhQsXOJas/lSqVT13GtKUATwemUtTuQ
z4sOCg7k6Y1ragEdiC/JMY465QBI5TSvfchQO2wuYkl7GpDqjT74tEJ+GY5cgWXnVAYpIIlxEAGq
AKPtK4SNcCp2xMizOD1Cqre0oaJIWDo9lxqhTpMBtZHaAPfSWd8hfmJYHnqMyZFKByR6YiQNVd1/
hAyjiZ9hxsFVtLvKp8tiYZmHnD+GEiZ1HK2zMf8nKu+h9OcO2dPE6AUCClvh7Jw8vKaXeEhalK9e
sNaUeWdyN4HKemWV7/Ulzo+XyChxk8fubGXenI9Q6lRpfjA/UELsPjM52W8B/6bxZ7Bm5iwFtYW3
JUdGKGQJ3paDoEVGJqSkQ1q+7/xpnCfvKM5W9uQVSCjtIuIuhifIKMCyD4LHqcAab1SrpoZjocEv
ZodaONRhUmSH83kjyBGh4RaxbDU0TKPHn+vFEyygA54bXWnKn8s9ALZffBYVgYaxMu3I5A/kKidv
mA4wdbajZsU34wV4J0O7oNx/RxYo9wT6yH88oKY4T2nUBZ+5Bn1vb/43X6FYhLAzj29dk0fN+lMO
20vdnUMtEtkB20ANw5g0BnoFk4vi7wG/wSecarKLKCBONvphcoTphTjV+zvO205LCFwzfdIFHmpm
bmEVypoARHalNIUYH2hY+o4D1Fm1VpE7tS+0VExNUsHxtZ1YZXM8QduwqLf/ne3bPm0Uz6MSXu2U
iKCDz2a0nUJdBJ2ZgotEbwHYBo188UgmBLdL5OnncH/GqWIMlH9eqtFDVAR/C1Fb5nM7xvbwQJ1P
vlUx4dCqPJWcjX7xI73fEPndwvQL12j9+8ZBWs/xsK236pnDeew+lpjMlQ4pxvtOI0dz+zkw0P5F
/Rz19HZtygynEl/EkkEkNMsGNN9trsyslHkCpCLFw7+6JzBZlJZeF0pq9fw6NZm+FH6UwrsVS2eP
0tgDP1JUYRU498jheVAUA718S+ut+iHTiFClKdxZ2O3yWnYggUnp7g+QxBPg6723W/PV95i8tkm+
fZw1Ax0KlJ4qafjMvIC3wiePlU8uJykv8hUHdZZYgj8hQ/CoG9TzC1MlYYaEuWoYAb+4LrUTJfK8
1gkf3OgBt4M9Cc/k0Pikqci6QttzsQPwUDtNaDjE0B6YsBpKkEfvdwnKmMoNHqB60FZPLmQR/Vzu
ViOsBvDLaO1cSgRuJidhhaVhhF1sVYiMC9ncRhVRoIuaINLlc9SMeE42eV7U/YIRW+mOVL/bzf6i
2EMD6EIqPYbZuBlf86QwJkCQBD4f8O1CQgUFaw9k7uqrnPf4OITaCZoxC3AC8mHYHmn3iMpGpNd2
X3YIx5IVLdqO0GNIIPotW4a/+WcXQohixYFiw2Q0r0K0wNojAVFojNr82qJ3lTtacw0nAnIadHRZ
u8+1ePSLML4mei7udPoP1meMSZPXEjxCiyTIJYp9p07VgKJKI3RVLA8zs2rn1hYsnErroCVPvRn5
RbZxUSI24icizPGAatSjTEILegJuD7EHBjfpB/4Q2Nxr+YHzqrQLVfNl9poEPYI84ILkJs83VyJ8
XPkpZaUqA00BRlmgzLPiZ2Z3AdAuvTuZzU3rs2pWRguqc2i1SHKXrKgUR4ZRy6x2Uh6sIARsQf1z
z4Bb5CFbe7IjdAOGYZYi4Ault471vr61NwU1RSEKSrXTAS21za8qgNBsd4afw0ya/U7np9nKNnFA
4tsZfaAAp1ku8uz04W8UJs1Rb4oPgWrg/B5qRnYz4CV1Plh9vSgvWeBcRJhMSlqr6sA2JeiOcGgo
62MOfwI/HnymrF+sdSiKpdJHxev6R9emuexaf5FktMhkyJlEyLiZHaTfSCE7QxwI7JzRsiswCMAe
KIVHyvNtUrSNk/2wQF+M7hITbO3b2RPHKi5YoZFDHcNrxXRWus/y51i1aAA0uyreqWaRWoBae7nB
eo0czuPGYj4BMizT5n6d4bump6bQptSB73tIi+zh/RSdZOHSkQCtvDo9xoxAKTPqiTSRO45p2ex+
aBqo5wn8ksBvXmLKeOm8xL+3xweKfKYdgbKJ3EDolXvFD7WrgTMIYwZIZTGW61DYpKS3Xu56FER3
6ih3YQ/LzTajXv2ezaNk7dFN2I8FUK0SoJ0lyy2F2gTn9SzN6/KZt0iNpHhRrCXLeUaxsUs1d28A
OdlJachtSVrgad4cBgFpJbbyhKJJKBsw+PY6VgEOZUigJCpwbDF8pZO1hoTVVPNh8aWqleTm1WWB
FJUm9Edt8yC0zj7TlHzHYwdHRuVjqfSZ400L77sV/wd+1Kpk6a0hP54aKpR0nOx+OmJc/tYlA5op
XADuzn52FoFWS4bqcnb5/oLv6Ojre6yRVRRXjzrlQIcCxQSYgPIWTqjt4vj4p3aYDNBKSHiqjIEl
QjqiIjJe7QYLOF0Cw2i4K0/+l40hDayELuMcsA3NuJgqe/PVUk/rp8xVBoBW0iCm8tmriphOY84n
H6kBn4pq91oE/fz2jB67OhhJYnqnq+TojNx6R/+Xzoa/wFJ3RqL5+4b2AQ7irgzehyY6/3Sw+/kD
mWgVFL/C1lvPNPm0XYDgxKRFgYC5pp5HxUJ1hdsPwQqtTOxynL1itV/4dQaplZ0L7f7E5xSUgcOK
eU9Pw27whUHaKLtTcMTWhRf8KPBZqt6mSY/jV4blwAaGPsN4wDNgdEAGK9WSKKzjryWSi6KNya+e
G/gnqSSH6N4+W8riQ5IbVYMH8U4J/CI+dheXSUfty6VnEOS5pyF7yMwOS0ul9veihlYJl9Y1LCNU
/0/hSzgvA4Q93FJsIPjm0GNXzrdV/OxhyLqMl2thSJpCiZLV/hlhw9nTVt0rs/dsF9mAb/YpmFrh
bfCeza1mG6X354sQIGcKxiIFJWiblX4lSnhnmSrG9GeE9PCQyLhVtMMXGe6nBqIKfSuz3sacuYA2
tIJ4Y61bJBM4iCMu6wfLKxIb6KDxnJtC5Gze0mVqL+ul9fHBdOwd3cOPokGt2HeqZAc00F/Nd0xe
C29Ccd1xKp0AN+DKisap8NZohDbFTR4Lyj5bEz34Zm6UK1qJ/d+cvUstdDkqcbPrNdVSzF2OxNYp
t7JULhNlW47k6/myXGNWuS2XRUtDySh5wskS2KzRH6J3CNnTovkhdcUQbcPpW05BK806hy0/r8rU
fs1Oz64kD0pJt19MVVEtW5Qrcz2/cKr10jdnALLwpFubHN9UMm2l29TQhbICMAbPGiZ1ltd7UpEf
ZdBtr8ZmjKb4gtvMb4Frq/1UqqTkE0Q2jxcswUI6jbj3eOT1UyZZnbar4NXuh82NUaKjac9CYwJf
WsFaHu4eXzEZL+6DqIR6/MOJzUM9G3EV0sOBQztyHXB8/FxNe2DcJuezyN2FNaVWiGv8vYCo8SdP
k/Yc3d+TmSYVbnhhbOVGqzO/jo839jEji36p4VdiSNrDYoeQHjTpdQtAPWNIk/wtV64uI9easSWI
5L2yrsZWJcA2DomwCbFYFt2lxWsSb74noIrrnE5y0bwF9iPUaP3thi0d6TZADynVTjuJBlsgNtia
62AgzYzJ+8utcLfiO4yzz8a3DBARXszL6F1ngOsaxFZOGVoa22P5HDqVstoCG4kxmAQIiHI6Jt9L
uoy//d8Cj8hDa1a1UuMWXXNiauR3oVtNTFl+OEFAwlvZt87zKHX7v4Zatt2RZHOj0BwXmqr5CHHX
cfeHUaTPqmrJWLRQAs/Wx34rwxUvuwPJ1Ah3zfXxgJUChDryJAn6FWm0+1qg8TE18apSJvq9EE8P
uj8WeLX10frpYZIAKFOcJSwETjKDG80J9GkT8wn1uczudT9IsBmvQfQYAelLJzcr9WEPCshRpoDG
taU8ux7v3lqGYLvsXaJghVOlIfMfGXY3XThwc8Ol4Cy5tSlvswCUMUp04FLeVjaPGlj8YNwATPpa
uDJoIU/vff1NoFmLQBYtm9vK+5ZMdBvnzV1+BGfblSj87VvrBd9Hatq9ioMYnj1Axprh72v++3VA
k8qmvPR72Hp/sz8fkPQj6zs3SStVjdgi0XofSSBnQCPPNp+ngk8wmEIzEXD9wWTL1567SW2AkDSl
HPiwbMPk42dXYRsUuwd0Q2om8/KN9WJTqhS5q5yXcA4RynNTM0Ug8UxJTF6sdlbjqKDx5X05xLpi
wfj8UlKdfjhLZ3FvxLfJiIfwi0YqPMREEA1C3jEe3NJUYNxqcZduiiMiCQuh+fjnJZFX+zLRxV44
HBjDy2BEDgQGC/cyoiuTjbQdU9Z2iZVF8gwHs3rFssGjXhhHLw/d6Q1C1Ch2rUy5FAuxrrueFak9
fP/e+4TZUFVydC5lU28HjArnTms4ts0G/5vbp5D6tC3V0A2oqiQgiBFW3a7+WA8GSqDdiAl3RpwE
NChhFCyPUKdvoTOauo8/Dr/glWdmyu4yzM4K/ZO90C9qjtc1lYCnfkiDEoyLmUvHtMNX0x75LF51
yBl7XzlBbNQuS82GHKhNQFWS8VEHuPZI3lxOeqpNYN3kbzA+ACilQ6Q3NZ1Q6XWwjO43Td+pvpVf
Eg+L7xmY02LBYN5yjCll0kX3ouu+/QpCmLo4h014gWEOsLk+GjhZDt8SdTAz+wQuqLiJeSQ+3EdN
S6Uj3RjUiuU37U8yzkUez8gY7oEioiAYoNnFq4m9XckDj3cvtUYjacflDXG0bbvhuhPmN7uxP4GO
ii7wdbp6bccxWfq689HUbWKyIM5FySifAllNtrGjVvYI7/j0O6ZgDv+B2HFh0E/D44mh6+22Z00N
FyqF5PIyRKuntp9xiDgoTgzlyDmempPlXNc1gkrDRI6G/e8aGYPrWYeFqYRHTcp0lEIEO4Vm5JkI
hIKoYqb3ft/6vEPxoPJhl4PvYs8HN/RoRmYlMYly6knL0I6Bv2iLZZU5i1z1ophxJ1vv/midYzLt
cLWjIAcI/wrrVBlC6YlTGo80avZv6b5pObyGIZ8P4ol0TbgDmn5+1oHP4HXzlirynFZzVX/ckZn4
7v+Sear7rW4qnapq4UXxVPWRdv9C+Z7c1YNrFJOPhd2B1NZkn6pDmr58on7/2CHGGLH1psqmzSM6
ZGKZzid3QktTxsGlAE7RLcwuqjbWBCOhwS7vOsRSI75/4ThxWWrUxr7t815S0ymwn4dO01vTWHsp
tXYJk5184xZo7trG05ZRmkSmV5+ygJUDLlBQgWo2na2zF/jm/ug7ktt3tgc4v0TYQRdDe2g35alD
z0TL+Fgz35hFnHbKL1x2cA3mtDt/4h1B9/X7a1nJKmP8u0GhcYp/R1etwNAyFzS+0ZoJ0GvpzxXj
j8s0qyOyR13v7isCaPcbkFtKwIjxLazFqGHtvUMPSq1q8OtO1kUFZgcFgXfLUdZjIBep7ohlBTMN
gxgm1aiyighLQmUhVDyYwtzrlHa9kqk1NYRV9LsU/ce+2AKkpSG575MC8bEP/YDPP8fft0nimQaG
+X5+yr9truFbEfOpffnjxXhi2C0QlbAocLS4luK3vvxBPUenM7hdSOS9minIGZrF/faIsV7ba1Lu
RIfPEOFrMDcgx6+JS1pQleAEwOQJqn6aVtAUhMt5tTRhWEWxMimKBeeS2WsKknEKt29NvLkC0lLt
frYX9iTusZzt7FSdw4/Db9c9O2xKGSk69ZESA+u8XGg5mIwK0gQisE3+HGOXGa+2CEhmoTGAGcIG
kw7Iq+PTA1WGXEyB0o6/5m6mlYpQelrsdrkbJgVWdnLg/gniPocbfadTBKqSSmVIuoK6VmfC5u5O
06pemGbU5kFZHYWWyrEoWzaAvGPvmiDcYvhn4UsRemvjePmzf+lYBtFPMQqZCsb/H12AQRLSEbCt
lSkIs0hh42RzPBLn4wyxHnmu4X5xq2T0v2gdYakTQivAfNOlkRHypXcuJxPpWEAu6Nf5VIvY6nHT
KZFOxVH6gAtVcudzBK1/Uin9cIKUkdGARn8VvANF0ZDWeN9zRaTw6Wa6KTlkGhjMjAoUYedDPrRt
+FPx47dL6eAtaGt6xKu2kB3+/tqCl3CSFmclEvhp4LXD0Q/gRiriHWicL7X/ZRp7jpUMB9zUHVSn
UtLJVBChfSxTk0A+3VxbxpGEbKoDDeIRIhljaOFZOaJ/15NMNyon3UQVSLD+RzYGrtuoY6LHnfFo
gEC7Ku5cpB2Up/BACIdKg7DZK+D3BXMHPywOY4cioaUlO4FMnKMuC2ovg0zsaq/ZFKfq/mL8E2Um
ivBmiyfJSDK6XVjFa/2A5nsKmBsj2psM9coEMN3co0T2zRfqXO1dFpq2jXpucG60LNDfBwZ87AqA
eGhvjwuSVSE4Z9b2pK1LsaQt88MrC3Jps+eMz1jg5Wv4RV2IhBnqF5gQtUORC1PrAgQA6R7c5ps/
UunPC0et89NSiWStl/WB4SGiYxL5RfABmonf4m9gopnu9QR6im/NepyFBZybOanEogBWJrHS4eho
7NqRphAKgrf/LBTV7vG0sWea7iuoGKBFLjnNRmaR4a0VgfjPKX4iL7G4gtVY23wo152YTnwckJJc
KAUmY9Q7z1cbctcvXHQO1fxlhccfEcuv8zqNJwQDBGR7YlHR2Mq1LfypCkvEv0ZehTMqiIKTDu7Z
3eeGy8mJZVNq3wgxhwZq1cxnWf+7vQXu0TA4a21TWfCgmbhTkOlweEckJBsLTr1YwGKjrn4am7qz
sm9k7VZeW2MLsodtFK9GWRICLAhdZf4f5znshXb8CsB0NzrQNH6IVdL7KCxCJuZnNjSVo35JK7Sv
Htdo8bASKEEMw5OKoT2lnQ7lANjwwFSBsRKP2zWWiLqCmF5BxwJFkM0OVvd3coPkoxo14xF5ETLH
3hq7AqRjia9eTGaGnFicjq1enOUWkMvkE+P15fLqEubnm/LYM52FpPLbvDRglMrnnsxX3d8erI1j
23z3qQUfMBbqmFvLsDVQfIVyoHsfFamchQaRUqH3EpWcj3msRUsDNfFgpasZMhr+1GJevP1AO9U0
ETQI/+v8DvvOV31ZkWna0tsf1O6li2l6U0hMK9+EVpvDetGxQfZVx0Qs3eJVMXZych6YWX8AA8v1
whRfgM//767uUMHb4ldj5//Wsa3GYYdRaF4c9RxMOyzmJw2OHviZ6HW4/Rn0jbYljwq1s9iDuxwj
XdZBmJfYWvnY4csuQfAV2ID35ODD98yA5SRJe7t8SyVZavP+3ZV5vS2mpl8yzIHEMTrz44tOLzrw
aHBTI+ussolqsfxlLGiKaPc8B1Brtl3He+fWwaUmCUFECPS3tAh2fEGfG8bdU0yOYwONatPCYaNY
IkcbabXttXd3jhh2NwHWG66B5RFjNdJ8VySx5DI7l3OHCkm71e70pdwO9vHS6k+9qngbEDkjIlLB
hPIFE1vrpT2vlAFvE09EAydgZJprK5F5HQVAK3cu7L0jnrxZ8oiKSrkQMfxOpEXgra4MbSAJoIMi
VpjDC8JUNuA4ZDxnl+kfpY9IARExhEbKjyirhLcDppgRZsIY9lMcibXolSH0oODDrEUElr7dxlMB
HeE3n8YO3/7C6gJWPZeYEJ7znimLjvLzRotmAsEsoynnBxnT39lFRNleKcetGQ9b+sGcWUrsd+V4
YSNYwUkV9eVFYwYPQNi5HGjp6gR7ZmWiQdpaKrjBffoShYwlSbP9ir5W4sZqueUtEWOkqn5eiseW
IBqY1n0Lqv/B3nq0UsecRNg7eY7T0LpSm9DGwcbDiJk0PLFaWUzn7Cds3USXnWhyA6v/CfF90Ck+
JRHV2hES1I2eMvOdsstpUV+GdWBgOgCZ/Huu7nwx4UVhn8MbkUeQGCg29aLGG5zknA5HwmfxlaoO
J5shmzfPNP/biXFQ/Ri+Z2l0ymcD87289qL5Nto0jZXu5eNIBtJQSq4olZ5bUHWOWi5BZn/yF4WQ
zFLZmNiOMHmhLqhx+5FcwbjK37gJ1hisR4bA4ZrhP7t93dy7QMBymM7pub7vtldGch5+jRyqTJnt
/wAAzjcNBr9ODLxKEA5IEEKKu2V62r/zGi8LOAXUBi8T5lfo8QPDx/EaVyKpEU0KPvGk9uKr8jer
xRUYf+1rsquorXThQ+7z3kBYSZzaa8kj1gq9iOqmBZG9nfDegF1U+RmRKI8rK6UJXQ+qFyDnjPjq
4aoxr2kHE5ML7TmLmGoMzOyNXKYUDqJSwhFm34mj1wu3ItGZu6jrPostgPpag63kNH2pt67e9opZ
GT3CNDbAyrOabx68N3NutGyTocE7DfTo0+1sdsS3cpefCLJj/w9nooaekAnWwt9G1FFgI0WW+wvw
3uQSctObFc+sgciUxgmPhLX6eqSnOPyputV0MJ50zzHYc/Tz1J1ERYZd9FIkc27TH5RXqEqh1WW2
xbJ/z+oqDyazOImXK9MI2IEqlHWzfm6v4PNZYLy7qfjOw/4pG3LHRq+p/npMGHXHnP8B8zENY4bc
PfY3RzuJOgB6NxbPV6fdWhmrRFf1PI0WluQtqUXG2eNMarwlBiwHiYYKUg2Cd1iR+2MOsYW5y0KL
RNeXu0EMNvpPL5CxXX5Hg2n7kkn8USVjbE6gtR6HQUY/Dd+Q26PNf4h0Xczc7Ecn7noDw00DFuZk
xI+la66n10Q6fRyl/3+tJpkvwWeCDE9MI2MHpeGCPZWmqzJxwLX09k1ohls0pYQuj7oJQXsp1swa
wyeVarSAtXzvMvTMzN4DL53kJOwTMLXerpeazA7kW/t9WyPAT7N/7db4bxrahG9ToSxnoU5nL7eb
nhJ0EPX5YnwDqJE1pRgSxz7j3MIoX5eNEeJKrKcUzhKdVKDH24tEq3Fu56zngh4/Su2ZC5ucSYV2
cuak1fk+qrFFf48uT3h4DRbC1H3tB+pB8z6Bfg1BNSaGZpxcSl3HgHVkidFWrU8rPyE0ye1Bp67M
gF4TNA+cqI6E10ix2Ot0WX54B/d4K4xLx5/D8G2tes6wVxXJhMovTMp1BD+tjXjAH3s2khJYUCog
LiZj2oHnKMvnqm+VOAcOH3t6lI+fcVaIL9bAaYu+cR3PJYo3k65IDNNe7IWhUllUGi2/MFmKRN/V
ljMgRsr28Esovy0f5GV7cB+omjrtHg2S+1/6r2ovJGqHHtjI/FRwRviCBHcYijMvAIkJLQzrfaB9
X5+yUY9k61ViRE0DRNFktA2DgX6xaXlXXHbNAKH/zfkxHg4yHVSj2t8zNXwvViI7sL6Hz7G1KprO
zYckrhoRn7yNJbkbuzahorIHDPejQstO1zxWFOHhTqBa9JsRjVnY7yfuhJx5l5EEr6ZsfCxo02qI
XK/sTnxvKIEOaPJGltxwoO/mOq16G+DYxp8npbLxHbgVsJxiUNFP9FMH21rYNd95vJ7oVpNuw6rb
JQg21FtdXrtcE+F3iBaZjfVwi2OpuOmcnczwtaEN3tLn6isdIEMePOb0x4bS77rGBYDgVEj/irsf
7BXHo9FCXJxiK5whPyJJxuxMLSJ7tt5SdCAEZw52gmYMg+QWe6o8zih5EQqZ/8YjUGGZjKnAOvV5
u2Fpn2JOvXG/eWR/Pd4rmOXwqT0IZbJIKBPBZ61Oqo62AcHI5Bpp22EgpLCF7HCO+uCl3GtouW75
05ezNWZ+lK/IjaJIV3EHtfFgXAj4mN5f0lPkwub4BsCz3UWfyAXCgZJZtrGocrMwwk2JU1J80S52
7gQjJMn81n+dphDFcpaLXpiiQYmZ7psJfLTukHx5j1Fg0Paf9iyyl87i9+ul4ddL8GMpdpWtUnM1
ZehnDtNypHyqBtcO4YyHuOS2o7Xbzb30aQD0gATovO0xXjm43gO/qBSZshJJ47w9IT39sbFNUVpo
6x2ofqGdVMUttk/5M9q/J/+cfOKr538yayphH6D8w4/jl6I8q788sCj17x7BAPAWeFoKr4TOvO7o
mbx3xAl00FMwkZCofeBdloFw1GpD2ikYrsDtXJpbIw/ef/KtCIzfBebMcPoOOlc54jqFxnT8J5hy
sVmNliYoRQ2pUM3Jej/UOdvm5vO3x3V/bCyqrvWase7BjgCBB0YqB1SZEovKUONYdfTrsyv321wW
h6iNNR7hqOTCDTxnX9lQRuCjlLhx5tEdm/KIwMUfkiauW18yWF5UPacJ6Ei2kGNvjwXeksq/cUIX
YjBAWn5pEkbzp4DsfHlHGKSTFI5HwJxRlCm6/8F4H8AzQDowik7uKZItOEUaa2KcUQT2AVJWrPi8
rWw1TzDEhRi5hqqHvgp9uO5ktaIUO3pwMRpUUWfrMCW8dohwjET1DM5uXCT951HvoiTwL5U6YLEi
FVAXakSeaNZGNnw552UERpTIFspBz0pgDgb9Bj4U4JDqFfS3UGQsdGgcYA3tyLfYmMrFZR8I6z/H
uCrBNJbQgHdPvuAxvNsaSldk18cgSdl1fodYpfmZFpsCyl8OL0s520sp7H9KJ+f3Km6s+I+UUB4Y
ZPnrHsWTJZ96j7XtO+iPaZX+XJMmOUFEXAJPdK2xCcvv7AMP2ejS5spOcrF2QXZVyGQn6RuMTurS
Pk08BwiO2d3c6HBgaHw6WWiyGdMoqViFDpP7NJJ3PP3i8HnWp34g/dGB863cpEIJr2+rk3n2+SO7
uwwam0YJ6J3HZ2kuPWBDB6ek46NP92UVe9FsfgFXYbMloV+2rDJLS20bKQ4XxVBnF/VWghbVIPBn
Y8icbIAjFxrKlYQdIoYkNeI8adwTebmE3UKUyoZAaAKSDy4exZXzOQMkD1rcJZp5EP62QmJCWGrz
8NBa21ZVjConb4xqVgdj3uYie2Zb+Cos6T3CfDtKn2LgV40vdrZhdRD6hqnpTHOLG5JGzdFAmBJm
KuTurU4yUkAge6j2YpQ/++jP20AWe4FQFG6fUteBuXA4x3wp2/3q0dUoeOvj1DtRlMyZyuRp1j/l
Dk+ujpeexNF2tgxkyxWBKCICdIq/u0xCSn2s4EaMNeYKyFbxzchhiDbGkV00S//Cpd+2+YtNEIB2
qjgKAwURL+9hOeremT8tCgQAonX7Ih8KAzZrRORctO/h3igCXW1hv+4S6zJBEB20IFECVsPaGhln
RCQYFA7OV4sn8jq3oF6CZjnO5BTG+sy1ftg6LdWFHlDCt4KZCVcIOkThc5PQAB32XVEqvVcx6ZsE
MrFnnnw7h/MKObsql7QJGiitP5Q/D8AAPvvyF9fInQ7k/VhoE5JcowaoYGUb7yQsvpILSibmtYuP
vkOb1YDlX0HKQD3enQ++IMQruRq+hgO5P8CjXKCM97S7T6IZ+6IPRtew4apeqNzaBwiYSE3u8jqa
q2ByAGGJHqBaXe+h61Q9++giVdvRi2Gw8zBHM1R9n0s4KD6ftRvXD/KRJ5Sh7oWNxqC8ulnIMhoZ
/jmxFHX79DE4X/AT70RGRTyaQtl1W4BISFY7VekgJkN1Mc2Hy2nQVBPdJL0IoYbPX2C8P7L0ppzx
aKJfPqhB3yUe6wp1EPbL+jJMOoFteplM0/5QW24Xq19GD1eKIvgyatg5Fp5GiCx0TkOzgsUg9e5m
RUa0TZuPyD/W7xKc2nIEpXmY/TU6tjAHB/vIJz841uwqk3a4s0L6NVHVKcxe9iTRkA5uLP3dgAVo
Ln1C65e8HOOP76E0YIXL5GGLXHeujYXVS4qF50wb6rPt8sKSu7DbboaLv7Xh+/yPqKYy4LcW9egj
9/MKRTdYj9t8pJ45QM8L6JVVnKE8eMoiddH8aQ183C5WGk5EhCJH3CAycCQhfHxEmN0LVNog9/GD
A0+3ftnBHmdceVycps5l5WuJae1R4CdL3KXMChBgifpIHwiAjD41sxJXzLSQhwzbZ2v+ljFjX4+X
LME48CpIkmmKIvo2MULsgXRq+Jot2ke0YcJ5MvekMCP6AzLXD4o5bx7KvMLsrf4CvTBH5NI+HG4r
zK2Ymaewt5jJA8rCN7Vdds0yPAOzGRxa2LGQl1fKorpxHD+SJMpRS5G3r1xoHw73fSSwuNiesIHy
RsndwyRG+EyRRD45ANp+bFOvHwxGMABWW7xOJN8dRTPtCOf0VrWpRLj9VgyGc6g+6lniNHymdVod
yoPN4lLwEJlOnEWYpjc0zmEIUfzDSS+8WFnVBynYAg4gu/ZwHUmhsgYJlHp0Z6fGxY+Ks9PjVMEO
R4y0lQSEvqi52KItRSgnk+faJHcjNj6gxS2puoImvUWgPoruZ+8/QuwqkAgVMaXYzLpAH3qGkaPQ
KIyWHVT75EfnvxP7WNCLpkTSHiT62LwGqSFKgyduv1WZphyeExCR7s2HpKxBuYowFaC4EeJUYDD8
pCLj7C3oLRhU59ix6ueyFpwBZAx19nF/jO8YyoQnu3hLXGbmoqo6M+JRFrA1wqSf/JytgfkR2BNs
UKe25AJ+rlru2eCcazchZapYP/2UOibmdChFGl5buN6gc2IDtbegD2fE/cenPNNfkI8UzEIhqrnB
sMZOW/UH0enreRL6JnfB9s+iZTSLqsBHEu4EA+gJgaYhdel98KEEsEJ2dPkOz51Zc44FvHH9LZfA
mcYfPepB93P0i9uEGOJpGcHvggrtT0TYMFZD2Jgwx4Za0AZ5slPSHXvIeBtiOtxgeV3sA2jZ3HzF
Y/g6TtucPViG0qbzTOVjz0YFqDJMqkApZFfLiOfYm1xiKLhMusWl3rGm6A+wpFdxkjTMjI1XllYR
1yH2niVh8Rzp//MDB8UV2TtcYVmbZTVL8WISeqA6FTRtBeiKIMpC5Ex5dZLX6Ccljf4FwKIKDTIx
h85K9Bz1NvnrhFecDLe4UW7nuv0PORw/eYsE0wyIkLSJvKuCa0/HJtgDA3bn9JN3+6Hp9kulizU2
dhj1GSir2lxREqIRcVQh89fCRYiWuKj5JYDRtB8CDwivu9bXoOa0Ua3BE/dg5F/dgOtPYCjpL+Gg
qdzCIrAZNHj31kRMew8eg0MoSt5UlQCsX1CCyIMpWOtkYyf+eER2FQ3PrlBSj7jQVFdURrPKOi8n
yXG/Lvy90jgXqPORkB7nMKIcb0bJhuzasxosVxx3SC+8UR7sdXRrtXIWOIRBUbNHt4eL8NLu2mGh
bpiqAUseMJJFgOPoysEXuxDONxT1p4MnR4C+myXki82LeKmU8bjyCkm2t1pUiA4t5dGogEKqPYi+
RA7r/idG8ce9CKjCxhPR2HmXqropCUwS7QZtM1Y4+Nn9E6FXT4UZBhMg2iSgPNTNde3dyElPsW5b
xqs1Kt6+7Y3AYGt2C6Nz4wbmH5exyyGZz/Tt6fpsvZChP0EpxhJPLxTQq+qJgLhgueKOWdJRCHr8
w3dBMUBJutwqINrk3SbqCA/ga6dFdDDbMom3QZHDOWSXEjD1wwxGPwofgbbN5i/nXMkTNIkXzVTJ
uBGx6DlO2oCygW5vnQfUEaCTRYNqeEhcmgL6+dbrV8sdDqhFAKjS+wY9kzQ+STAhVeXS7Ydp9pZq
ClUgjtHbLvnFV6I+xSPhmyh4J106MNkDlBo0M3+kPa61PARDlG93Dk5CkK8jWhMg5MHt8XLfsQqW
yx3FNjN9AQr4rqMwKMmtofG+0rSMwM/WFcqkQWSylBCE5Kxbk19FWiFP/cjP5l7Eo1fc4w5iQeDH
JhaP1yxDkqEntaqM7OR+PxvgR8svJQ4VL1Zrof6hwtdCbxwg0Qj6XUD5S4S0wTkD8oXIEGXaNqwK
6yVXz6xYW4PMsdVTLsTQzxME+GOEeWsX2WfGAu2XhdeZXLdTliU3IYKOPuNWF0cC5uHtzHvgiN1D
xA0fhxoTbMoctIVGqOfPALf3LjfeXZ2Q52hAWhhW2/BY+rBit3O7aZJTdATi8v24fOi+ZrI3W9yg
cu9M15A6qDK3NKF4A6C9O+JuySVRetrE6vR8KLIbEepywoU+Nr1XPjQw8N3BVL5rQqapwZ5WGdGi
vgGvE320XhJJeDoxz29NKNxE4FNxXqtrsYedOOiAu/dBNRs+T3lfqqsl7E2i+oF3N9TsPfStTkOC
7IToigMZzx0Gvz/vbcOVtqFXSLCTIibbxe0xTYki2kZRKp1sTCV+TSfrR9CxZ9CzQDGzS0BIy/9K
NK2zeADnGQG/CzqC4LBTm/DHydEcC7rWCI29rNbMZgz7P7SYKRsTVR3XGkYdkAgjkTRoi/4tgsYR
xKN0tdqCVPIxCHlf29symvBZJdQz5PQ9BuAwYpz90mMGAbBtD1mimM91cFPjuupcOQ7nOT3hIC+z
v17fnyJbed3XsYL8G8TmxAhAcs9vH2NJEfzzvsZfqQ03eVJ6Urv5fijnWZ2YBcZ3qpurh0DC/Wb9
GUiMCD7LM8nQApgJq392LJ1ecEmDyCpL1aS54jFjLXSdo3vA/wxRqPitUg0W5pTfH15QQVCDeXQX
DyO6N80pDTPgBRoJonMhZmHnMrfAeSMLC7UAPOyPoIuWdVligstLkDtwvEKuLoWapK3mXJo5Blxx
GuQTyP4nrWZc4HF7NJ7QogGfa1aCDgfyk0N+mTWIfg9CxESAP/eSn+cgY1ZZ/TNbQysykRM9vwx8
lp1DN4rocxtnfa12cHfRXPY/1sFYtK6lQ2kOYKTiHr2U12i/DvQC+K0kNdAkZXs0xrEqvyXezPwj
g5pw3H2p4CZ7niFUl84gpunqVn3Y/WCb5aEYMeubbO8vw5NFthEP9DIyljX+ZX51aBG+966v81yD
FniJ/ZnQCq+3BZWDRbNt2mouE2p7reIS/KIAVX31sKkOgyec/7Wht1hKfsrwlhfsBR+XZKsff/rH
WxUr90t0MYDfsyPeeTeo90+MDbmslZW51wymriEf3QaG1y5FM4d6y8L1PzS31Vt8xeCJGwrzuSMy
SCsJcO7KsLE8PtrH1NdUBSZAmHdIQ2YnTVdPmbmN0/N6L9gzipxhVjhgteZ2Rvl9P7A88krUa73N
OfXpoZOAaZ1o1za2bBpLBC+6epacui0NNmlR4Z1iR0HPFfFmA2lsZB4VrMYjMS1ZUM6JWmL0HqS3
02m+rn/tv9nQX2EyMztEXRQ5mu/jsez8tnBmUDDuIFYRiUH/ekdo24GX53lrGFkbp1chXV+lX6v+
v2OkLgavO/2vzmW2yQ0ar8Jxvh3WtpRvZCOZfQJQeGKj3fwJKRWRKdNo9XVMgi4yqQddZ87638ks
RQ0mKpxXXMH5IW/R0jNykoV87QEPsNiwf/3Ar7zUKQXG2raJdIk8daiNaqfMdRivkL69qVWG4N7o
2yRYfcOvd6Ymmq2o6lT35mIP4HItG3MA9L1Dad1DZypMxQYc2PQRA3nqmlhjP7CRkxUFcbCrC8Nr
mreZ6mrxux4gvQqM5f/5SZkl5cv4zTQYJA8LJc9764vqAbXG2I1KvawH6FvobALX2+ScTU4BS4NG
XcMrKAXakYX5MnLI1Xv+EXZG/fcWsBg0goC2yvIZCzFmNdz4rlw3Ig3HhSh/4mKzpDL5YUoVDp3e
//AWMk4hRrZ/EWgDgXLEnkG8nSvuR65TNf5U2I3HArR9R4cxd+qGAHafsu6wgXlkyghnTNrkwbDQ
5rM8UiX7jO3xBWjafHLf3JfUwxtquukzI9y0ckgeOGyRM0L4GB7s64zRGlu7lzkgy6drzcLHPsr+
ZkHr+pJX/9NOmBX/AQIJP0CzSGLjQVVkmpSHwU7xiXIqAHWqk2bA8v2tqzufgC3HW2nWvLbxU6aa
oQURngBErKPXDpRDrJsphdK3Nr1QrDp/dfJ68962v3TZvOfa1x6JspwqhPC2eVh95CECRV7vbZtA
bG8+oH6HHIp10nRYNnUkg2j/yzWYChq0T7o5YanM6I+QtxRL0opnT9f+A1Pnt639eE/sxiU9+M+W
Ozxikz1OcEqxNX6z9mCyVVDHflAX43DxZ/Cb/ogrmH5ohfkbMai1DAB8pAGo5EXsZmMxHxVDzrFH
onm6YeAw7q6vsxQki+Pj60gK6vnsEu6DM5O9H7/kB36NKL4ql5Krv/elgcqZSGTRpUn+zmMVLxPE
X+UvuwWikk8MQfSiihmO6tktUIj9XS/3DcHzRyBWzkbKJrGqxFNRlviUyQ10OVuUJojk6HAtvGco
iQ4fUz28Jhphjf7atln3eJjht23s92tRv0ydK5I24Dwo4ShsLxmNpOBOuj0Y4r9JHYo1rGehIIMK
i1M4Vu1o8euF9zI09oWPWOr4OUCReGlE2DSNWrxSxhSTM1jr/G6YIAMZWYd7kTyA/4EwYFeltWdE
7mU2X1ksofCPSU/jmmch4XuTuRH8FsYeLXQ4nWAr7Fzg9PHcQHyax4gZ/Qc2qYTpL0rLoyvzDqoY
VKi2EoBfBNEGQElT7jEsGaPU0Vu3MAk/ujf7ZRfoz6wJthQfhJ8XXuEY0OsbUiWYfO8CG/JQEZFV
6cD964vXcO5k5kQ8kvA+ou5ab8FMR0w2rsE5LviubNBBucmy+3IJDGwcGGBOX8SB30JDPpECG0i2
8n/gPw4tt75xvQp/yzMXxFWAwNobmxz1fUlV/sZoWIufhZ/IKbO5QQkrCN0kXZg85HF8ERJ0zAQE
osiFWj/ICTPoj7go7hLStpyI8/irVclFZfkNk3UR4pXMJCAzR4/PrkR4R13Zlin2tx/eMMm2faEG
Z6pTdFBoncQr7e1nxduSWb48k/LUTB1yDa4tl3X4rUke/NKrB5yhKAGyb/iLxeNDJs0tA99bX5Bu
3fuJ9df4q3kcFL7kuFlmKRjyRzeW4FjA5zI66zfkpe00AfZ1uMDEU0olXAk3rq23qfpqrULF5ITa
ZcSjMzyGzky7gpaV3UwYnu0G3pZt0xhnXRn+n1iBxPPKK7ZNvqBwOsyKP4KsiqynX3rLA9oNls8S
7Nin9b5h9NvvTqBaR1HiSE2H5GZ1A8HuSWVtkanlEJPcAc9xBoCde+sqABjOc2FGAyhLTWrjhmOq
5eROekS+/V6APoc73Ml9D+CBcI4cPpbCaREdwpYs3WQcmgahGmXy4NbIErug8T4cCCbrffhia267
MND1BMJ8mOMzYejzq+NjilrMutqj79MAT5XQcFRzltsSJK411cBMc0m2guCRbXncC5YbFTz6kKq0
2okrvfBT+jyuhlgPc33tJYF5qyLHHfSypKgbn0lSnNrKCmGOAprjBgE/6kU6JPKxxYr5lf+6xgUT
2Sq6BNDuUVUqRYgN4aWJ3YEVBeNwvqxsEay/wCU6GqmG6LfTPeQaDnCf1iwnhzdt3zNWKOxJhnoc
um8nhfDlYWBXJh4XU8oAmzJgd616JufJn3nsiod6sQjUwKkwubwXWfQgMBSq1NkWAQ82kUIsmu0+
if/xQEtZPRHsOVOf27rk7yOGQYcJn9uU116LAK3PBn7rpEGAABRO0lTPYS0A9tEinSYR3bsKf1Vj
OqdZTvNpxb+08p7lYI4hauBV/0Au5lpFffmBL/AVZx2v6vTqINaCLwf7K5m0um3KJED2c63bXc9F
0I4C4hBqp/4eBTppFmlFjQCJyrVtLtlVp7eLgKHNaNKCXBZh/oLWW9t37Rk8I450vyyvoLrCfvT0
iExltLFprDwFUFT7gf8P6Px7UCU39odZPrGtq+vmr4sPmn/OkXOKWH/q9XvI85gN+FG7ySY1Rwwg
ct/oKTKC2weebtOfBazxGWeH+wbWqY0PeVC2br9aIe0kPHIrLATE8QdTMkG+B/UAWzwQBtsE3CNj
0MGt/yMiL7CsbbHJ27uh1++Q8A3fga9gmwpUsg9HPpVlmB9cOA3I5owLwKvydhGogy6Oq1EI7FsN
jIPhIjRGtqlQ2QmOhWSuqFF/QaD36gS6l+7vhNKw6OyazKIfqEal/CENEru2v2sRJwkiG8JR08hd
nb+Z7QlqNv+GCKBvDFLBYknQbwQJF2wocJbOoqEdHK0IYZ2wGGABIyaQubGZ97cTeW6GB5eT/kcv
A0LWfInQtTxMhP69tZtveq7AVmM0MsJCBSEKUjQHiBurspvt0d1fzNSHRik0j5wRReSdaVjwtVMm
8bAWhcVvN2BjdZZwxOS9IgGVSUHwztXCONit0q8HOc18++5mESDoYIvEpQjPI4SZHN5WcAODLUEw
D5inY+q8y0rvdF6+c2ReTu+foVYzb5N4UbDxcbSj8LHt/c5sTEKOLAbZgzUDYhlK8MMe0mUrBNl3
4yYkLycMTR86jrAS7XLnUWjhFiLWvgm0zJzwbIXrehay8gtrYJMuiaLe78b7lwBLd+B37Ja955hV
Zk1feaVrc4vIS0dKO70DsDuOEeMfSpRxpqZ7ZidQ0rFH+dZIaUC1EMNsC/2XI1+mM7NLLFh/K+wK
F8bke6cNBW3yiEveuo4rvQVdgo72NgdQCLLcbfVYb0n3x96vidCdFazLejL/nUKiIRmKyUeSB6cZ
a5707xv497Nlz49DaU0bQVeQMynCpLikQzulabu55Gl5CDsD7xPA0qOv4mkILKJ4KxCfbKZ9Ggvt
Cp7g27ZeUCvtQAhqJs+V6HptE6+v/UOXUnJBTSP/3sRsc2xDKvoK1RSdhSSVXbHKmtayvIXr/qZf
AQweVqXSioPmxN04Dr7BW6MqHDP5c+eshOlOuS0HQjcxcsvlKLjT+qmXDd2UyISiBZm/JhG3vGxn
c0o9zFk/ctqsKdVdWpn7qQztFh8asnrtEMlUI9j25dWm1Y2RLbbL5lMD3j+H07fojuBaxN2tlU/4
PltFPGhK7bFuShifZaqyWa8eNVt7NOJ80AQOwsw6RHPa0ifPMCKLItCT7CS+jj7gbNK/nDISjqna
llwEbxZ2YxG5MdtrU50No6JpcD78C7oVVUcLnj0vPTs1xkOqAlh/N4+k/+CmoBd26S0mYvgnY7Eo
rAUYsEDv8akwnpXE4/u6uU19ZVfhHsls0G7yJIp2e+TdVMcuKL4X791yeIE9JJjLthBFrwxJNTMh
oN7xwgzHCHjbI8wVu5ZSnycbaCkyNk8qpX1aJipKfYigS7Cn85dc5AGw4GlMftFtBca1DoYtQPSl
1h/Kn4XliBZz6XSF87pMkaPTYAt1yNLZX9JLCMy1AvB0R1GqRbJwvSYV/3AB2KTcSqKluT7ziFsi
GBi7zi0l5lQKPQxPVlx2qANhUIQUV6Cwxp5bYEc0q6ngbu5Lc54mxahsyMQn9ULyFwk8dMf1m0Jg
dUSLikT8HS6bfMdzJMiqe9yCVFi2e4LTCPzMOpz//xEXGoFFTBiUWA2+IQunCgu+fqy9dU105Ww2
ZtDbQvWPsG1Hnp5AUppWNmbmWtgHspMHriyIqgOEiKeV+wgfs6/BwZK5tf2VwxrXmEmlHTz+Se6W
BFHYzoKgTOQD9dVkS9HcLpKUzDuqHmDFfiLcLwLEozyZ5Li5DXOMHruuQ3YWgAULO3RWVA7VDGT3
hN9XeBNDG/bpu/k/WBdCHOvrGPoKirl2Ju/2o+Ck72MiTq8zYcvUQXn2xOA+QIWisi/+aKTBoFyv
BWwO8ZE9RzkI/ufCPVdN3+DKPELDQKmWGYCUmxM24ShwvYfLaenknZghiBa4HnOIYscGptMxpFKV
LcEekyOs03/Fpfbyp03O9BaTjCUY3t9HViciCAI2lc+8P+nd43ApNtyeqwKGtY6icoyfLNR+nCdG
776InpfNobJvPQVstsLoNDAdAS9KuqQROf22LkcN9csDGy48P4IHzbi4Q2ns1qfN2Oev+Qy4T27G
FaV59n0O5W6zuDav30IYEMnj2zAA5RCGKF7jwMYCNL8XwHT4PdDFs2BzFiLeFwPe2APHKEbX0h5s
bEefqacB8XhgnKjYDdnV7KxEXWhWi/eaLxBUXNyKXVPZ4GYWuptm8dXmyTM90lrcysNGl6wNbNPx
Op5hZJd7H11AqAZmpLgForH7JyJnpx+lNyvfbrjGepwWW64TY0pzGGi5ffQmT80o9PSRy6v4POzr
edvCCrtUdt+9WJPtUfcgn/oqtkIkFeVcca1NLsZTbS0ANrql45lSlljiBeyB8VdbXkJwvjN0TH7p
OD8it0OuPNcZvtoL8hixHeQEQHOi25meVhMOYgchH6fPNJAGKnqbDeubnsjrspS8sTbz04aRHWjs
jxdgnJb7lF4Y0Gd9PguDIPzNEI+gwYlpsybnhnZfN+1N1nm/HFto1A62OafcNUCApRZ1bsmSe3zA
NhhOSlhkzx9gDsKyd3++09Cwovy7a+l+q3/WNWNPiZYWylXKzp3iCZJjKFE1pp49FLOC+Qf9NF+I
ENjaRquKDZV/NjSXzTL4kQxVt3fkNchpPp24wolyxkQinBBhsCzL27wNYt5vt2nxcUMSwpz+2nMQ
jOJzLRC0kSQDfhYYe13NLWn9SPW0ibTOjYt28QblZyxabKo1oo4WOe6WgwT2BRxTZ121vKo/T+oM
Pv0MFeKZImg5E0RdUr88b/hOIbok0/LjOZv7d6nqfsLTBFQBY0ZT7cvSIb3Gf3aOIDmpqqFgq4jG
zFCphpK2P9OmQUmWfPyyFL8bwOWArJDN5H+5cY9pxLODMhjRpX3rZ3wpDaoTKV+sAU2KQAHHtx2q
qftPHJIH9kh8/JX8EwGszKvA+Og2KmLGQtbEJQlwq1LAO7IrrHCOOcZ0V5HTJ47KVo6CNtwKaBJF
r4u9zp5v3gzLMWHngXj0sxN4JkP9jycjbQ5o6xUtLptLsU+NEbJascUkz7mLtq3FGRIkWkWr05JM
lhCntveK/MgYNchPUw+T8+NOob28s4+47m5kauFguWIyTXpEFTYlOHce+ERwG+muR6ufsS8qKKFr
nSZxmJxwsgxYDuLCNmCS0Xd/5TBLzDtiIJITKlBhynOAbZTd0ZZsuHZ8x87LNM///HRFk0hsLrpS
VVkkj8SPKyKQmPc9Q6ZUEOIycKVERmfDUJgKKrznjELlNLLqjfygqY9+Ubkl+/XsAurd9H+ONedh
V6Ap+CkG2vVH7qlYCZB/kWtePz3DwEFNyUuC3voEQc3CZ2K5sfwSSKzME4vejPGXiis5L0MUIm0k
r0pWpVpIngc8MgqR0IL4V0IRny4DvB5MZqyEQ4YhVlHgsIDpBVRksBSUdBNXOeeHSf3QjcvgB/RA
SFsATOei/aR0QbVMiADdmQCiVQnA5hSDnWB8B2KNcO281bPwdscQ7UXZBrR74pO1++/PYZX5uAnQ
FdyzbFEPrfL6elo0o678v6ez8jj+VO7hEV4ImZk+/Tzw9sWzZAzzVon2+3a7ZxUkpR9QwORqguuT
QR/NDWFAmC5TulqKW8yqf8k/5wgsRMUMMK9md6VphBVcdqbikB1k0j3d3QIsIxh33irMEDfavsfm
wunRowLMEnxtLq76igUI5DN824GUcqeqjl1ugTCmrvFnmA1pXbnvYfirE4uH+J+YxdQb6V/gnp9K
YgsCqV8m4SzpN+s2Nq8mgbSspL+0KTtusgYVNSXyrXenZSc8zKyp7bYc+yKvgaIYyT82Djy8njwK
7AmyY1Bm0xJkx2MsUExcZse44LCmZlvcdsA/rTYom/dU6B3Ubpw8y/xE1pr0LjH/JUXDG+Ndqxll
MloS3ikp00HOCKzHYICCv9YiAHs0N7s8J2T9RL4iQszRTd1B3PgnjeyzMZP/jC+FCoIxkpUjRbob
jrDB7rE3oLp+qnHqHmTc9aq/PnfOkvDy5imAA19WQCmFRHzSJDWXEQ95IFK8nbKK9KCuFNj5cVc6
xp6hTpkPN81dEHaIJelsYz8j/MSkXNWO7WVJCHOfG6JzmpZ8inztHldy1ymakk/7tNbYO6fFN/Ev
6hdev2Afb/tGYVRNjxSTs0gITp2k3TZ6mE/Phlb0/r6bRMAHrvQiW4ChwdGOvCanWShrJqLuqJbt
T1Dhz/FoXRvdv0CBB25/CcPOrKCkgGgls2lN0fdDW8IjEZzeb/2YacUkhl5pZpz5DQRjkC4FwvQP
uLgxJHZa+M+XzVy42Bf/aD1eq3QwgNReMXCSTDnqsV+dU7Sgy4IpbkD0Z/Chu4AADp1Zy4zQP8SJ
ZebfPE2EeiJtWdvdkBOL3tkWPS8GnnXEf0UuKhbFGBuUHrmFyG0DtcnncS/GOPNzybO3IaVJ8bm7
4ue2YWv0a5yF1Jrcv08UlQMxOpD0dY7B+YKJSuV8evzWin377xggTC34ICR66nCOjhAGzOognxgJ
spFhqgLaxwRY714L/mpLpxZaewh9R2S3LVAKbPd4/uQfgx/eNYJjv8DMrkgCLe/8MSVjirSDuqhM
A+d3tte+CyebEvzEIGg8+nvIC0D9Jr+xSrNhdJMk+omhaopHgqdMK7US7lwRyJHNH7m7mT7pTfsJ
FyjHHnE1Mg1lgNdM95dJOLZsKztSr15b2YnShBVXFTG3WxiXMEMVW9iZQNoXUGPrzBEgiCdLn+Vw
3/ofd4S44uG4GdXOKGjD1YrQEtPh958haZJXv1rhpSJUFSfCRewd3DPLY8mxPdgTxidb2ckAApFU
kwM0i/cZaGK6XsBdxGKdStPkF06R+EQMYcq5321d0443l7hK+Rw9yGYm872gI+r1m9D0bIGtoGNi
5UTHMGcx+N6L71Ov21+VmDHPkO5hpn5ghQae9gV8gg35XWT1DBWk9PeP4eejN5h1A5oXGXg2J4IX
vKpx9A7rKqvbKu0r/QsqmSE1AG4BBoMuozRukBumIQa72RkMo8Bwgr0GV+iqaok6GC7ids62LHzN
RAnRG0nUir/oNM/A+8Ist7MjzLiEW0aP2PXKnLBMD/07Zs5/WDu4AbaDCkLug/vl928ChF9OxS1x
A5Yo8IruP4ZUOaei7c2+fGoqisP0c5sYIPf4E57f4Wai0p9cLSjF4ZjaOjpg3TYwObkEzo/AViK1
1/sPKVZCCoFTZtp6Ag6kJ/bohx2JzcRwYQ+j/arL6UdcSDwzKcI3lax3zL0I2aEIWZhmvL6pk/Ek
5pF1ypIIzgkVr0WT+18mazNBnJ8q+LuoRMXDdHGQ4DaeZ2P7khF5KlvYhQgb0LSS1qV5ruEtS//f
5wEXOtG2eAYRBpcQGWwxGkRgWwNwwVyI6Bf+7lmr0ZCZ+FJZA/8XJGZ6jJH6mh7xTQQcNTn9BEsc
Oay9dWAdIbK70uIraKjLj84Pn7ZjhbKGvzCPY4zhuh7MSU4zYT7y/q4b2eSX75tI2esJ3u0bBlXE
dzD3UuVJSRGcV2DEUaHLXsyBov3Ab3UsLz0b2HNvQLWw9rRo2xJjlUKcB9HCT51zbUXjZFGfV4Un
amvMFoDadC3mxQ3mkY2pIBq6U0nBwz9PYBCg+rg9QT7aRevFAKw2tJ9gtPzBQJg3zOo48H8/71xU
UZwvddqX8m3dX8t0sBWHxcZSenlQOmwR479MAAjJa3sOcjoo4F8jHiat54nUHokbtuMW4iv9LYtI
YiFVFiqaQN6/EPvXcJ6VBcy3gnxF97cx/hdBc3FMtLj9wKPrp72S0/LZDjN1ypsCrSnTfj1T6H4h
ymufsNifWBy4txiiM/INrxLMxi4rXNtanlp1KAWKqNxlZt3b6PDBSTPgjQIc2Q3Jd/ky3Mt6xKJJ
X7ryCAXvvKzQAuoI0i7hBfqTVBhHZ1FY8Z1BoBUv1rZ6ZLTxuXqTx/5cpB0qKMAVRZkCcuGx878j
J7duhqsQvMWnIOQFWVanmLCe+4D0yYXjAsTEztipBlsF97Cpe9p6Q57avpaFFI7Z+w4aVoztssvg
bNtbe0A9OzIx1aJBI9KcxHKAiGXsJRn2U8C+f4Z/KsYyXnyqmtxCr/sYkO57VMvvtq8wJ/5LZIt8
5ZXqmvQWWWnRrPZIJEmftiCa0tV1oe/4gINoehws7KVwGfhNdDegr14rsqhAHYms6+c8tHj4KFr+
itbYxi6x91gVOT0OKv5ytTqX47OQnslpZR8eWc6YZEHVBEYFN7iUpTKyWMtScQMMHmldgsOkCC5q
uoUOZLU0qzkCvGhiqc+N77xvSgWXLUAtC6ZB0IAI/X7+AbHxcRTKcQtNM/3TRiDYJN4DduEwi278
FrS/d1KiZSuc2HA6b9/NTYyu/4KV+0Z6PvBvpdY86/VtBoxl5OyM+ZK47uoj7xuMPP+VU6yhWnzz
oKdzKzx2MloKj1q176izioPENiUVABFWXVHzU+1+H8MLztZvk5IS0lbB2Pfg0uQmuqWw64rc8I0Y
eGxsVfVAZQQVmxNEumanOXCIXvj4bCO4+wH91y1h1I94NgW4hqBWrfMXGM1ouj6alWlTbccgqRhm
veYUq62LSxy9/ywfjfvYMQZqtH1GnkAluh+glZAPo5zhJGnEDiNFt3ZHgq74TRYSheT0HyK05Ra1
Ou5kJ4ua3zWvnQUEjyas33uZ7GxDJgDUwDMMCka9WP9golOeh2hj/DI2T++yC0V+KXLylFGdZLX0
h/sQ4ybF8e35q6Z3nfN9ECkAqRB0YCXZBiW2/v5eXKj8lY5LZqmaPAkVq6vhV5Z3rjCPWOsawVLy
TXrzPQdivQ2PAtFgqRdfXwVMNs3uXmxeBAgCJyyuWJCfdigQDTq4xWIWRgyQuB5XMkGTHjKTT3p8
9nEz+YoTgt0LhQfew3Iot0QybmyRUpiLoGrWOYZ41d/fv52x/KORWZMyiRQbpi3ojPmdbmS5MINs
EvvcdKPzNpxIhnXSye50tboDdJd63nbsQR2wjeJwN3RdrznbcnLKcJ0LHbj7iYc+i7YtHXTimolw
o9IrsftnHxR4Y+SsAec47BRBvsQDtb9ihpoTRpaqpmNwoVijS3bvkD5UKnjg2Wkq9f/sRIODtCdh
VBJEJZg8Q/TZm8ebNtaejONVO9V/AJpvLOsfxF59HzewX3acAUSDXK1Cfn53Mrz5Tjd6Ra8b814f
QSVswf6nSu92yt6YUnrmRvfdFTYdEfyBaioPH5VFpxkeCA+M6Ie7I0NEhtzgz8Xy/x30DDTz35Ei
GeEFQlBACjbEE5HZkzB9savAEUrHj5CDxx9+YbexvzeL12uDN4NvkO6WtiTK5crPoxR8r95KobB9
I8VrfOdW+9Oe9LWaP3Xbf6RAtvxj9wEQh2qHI1k6obvU2c3jAPCH4QIZRr7zrCh5aWIIyEXmFlM9
0AQffOaIhTvVwCIkkXZRqYXwy5zJ5MXcuXrvwgfEdQQZ8mOBGMfdyg5g/XZfB43pVMthKaNV7DzE
Z2vwVmC3pm4yYMkqn+RXgtAL9+2WqqeDL7xMRXkChvbBsjOUog//MpCMRw3g1xOMZMaIry8zTaBQ
Jt6J43Gew5V3SNmFjIfLjXsHXsihBqK44Rk81jVjf7sftT5Hls1aTxzVl4+w+OxfCLaNgnz2/wxx
2LfLla9GlG7Bg64CAExTOuffUswkdRH1t1mCouqBKL7VgqRr6CcnM4CqDiVNQDr7RBvv4zZFpLlo
mAQMO66hof9cmwK/w3AyzaDCpSjlB836hXFGO2oW503NVxCJEe+b8wu7C39cEN5z+J4YpvP7t3F/
Ikj+xHESN5KVFRslaoMYJZjlNmm65L7gZJBc+Rlvgdh47i4o1ADlCONO+dH4aPW/KvW2fuYKGqMn
xu31pYFhntm0lA0Wp8sAb/tcn1aXYIOUAxsTSEQkxzg36hQGkbTibQvMEAo/e40TWFT97zfAhK/U
i4WqyxBW7Ox2jY1OAAFzZ3h4Yg5vIbqAsfv1MFRLQYAe4tRr09FtTR0pfsWojjM7DX+iAVITG3Xj
hJYyFRKr5FGOmefhD6UVmVqtfgZ7B5/4IpOXqMR568LzLimnmzc9h8s6YFmuY3aA1AvYJBcPovgO
PmvfuD+7jUr02kEnVdW4jhU2+z8HT2G27jX2lQENrugkeisXy1f9ReZgr9HjYv+kmWzlSK99VupD
wr6ODq4tYwnrCZp70fosM9uuYa0P6gebmz0b4csLVKCb9A5elqzXXfjBUSxvrIS39w4N5148O+dm
5iFHLLAu/M9FllTE4mNcrXMMJnTGKb0YHeFcoX1p3KmKKmVGG9xcwt8NRERq5947ghDPCk3g1hhc
P0HqutXtO9ovx5vbsroQ0ra+ftOjwbN1utTYNZ0IyLGwp4zkcXI2bdNdS2aXDVk8cEODTaXB8D0w
TsBBqbZY642+4vAp3ypzbduBbHNCBg/kqd43PveiYllWWQqyoVa2Ngsu7H64VnWRoObgEFgQNINY
AJbb0Rood9G8u3hbdYjyuDyD15gma8d6fdc8o8ftlipQ6hbPj9CESeYzH342KMTZ1kBNf1YxJkmR
LDKtB2Bf59A/xCrciGYdkA5xcoxDanqKCg2al3b7XPHXmEaO/hoc4MaQ9HQD7ct5mFRvEHQZ4Y8/
y38d8Jzq8bEzhFs9NMpfZnZ0S1uomvB4aJekLPSwuUdD/BWFo119Kx31OVaMwzhfx1qyyIZFLu3P
ABEJR3roqPbWf7yxuAo8psAYz+arCQxb7ocmaYd4gs8rmPa9oh/Lk6KPjcJdxTph+Bj+1XHqRHpA
EwWK+kPdrRIvf7R7PyhVHVFzWM9ZsL9eqbp35fqbMEqH0zGpoEXGAdN6Fvq9Ej+orUApfjWDwKF2
NDBDQiaP67r1oLDdSAQms1zbBzbc9LtsJ2mOCm+46VROJibXKRxJG0hmGkFNv0h+w/Pz7kpDx9YN
bXRIElQWcJ/AJiJTP4T6C/FmBRc7YShsxaHN+8VIU7LuXZ88ATjGWTSME5+b+DDIIvkvsR6DC579
JEVJPxm2ZSqHCLSu3vbHGFFF3OulP27kHeY4+msbUqx7kK3ZHeUNifSP41tasdZcEJ1r+b6vV0nb
mxrjEyRl+21q1Agcgl8F9dp/OdyR9i1zE9w0SQhaCqLFwE1oCQ1taGMq8+DKi9EdzU6X33/Ga8Ig
TzFHXOjmqiy7q8i0x9RRouLx0bIO0TzO8PWUgZ027NVoMclMDGEBIQZEl0KlFYQ4UJlAjTYLAAEu
cc5KCnpFQtkyxgclz6DQVstwVhNo+pbjPJj+5arntepitSU765V9jeJZmsh37pHplL1cWH0N2kMG
kvGc0V2fUHKYkDpXRbIWX+JGR+EXdMzCPjjApwuaqIs94/tvpY8oL2PCh1x5+fMf/8AG6qD6rMsl
KmFog0Wl96nTyTAab3GVjiL4+Rml4ETqdUKTh87fDMkZPqOaf7ZvKI4N9ilbt8uubKgDSZc0eQiF
sP4shu7mwqCU0Jb+UXOKmsZIOk3qiTZbQBRd3PDQSAcpa92re3PbpasBIsL75MOrSnbNNBHesE7Y
sAEmUvDOiqVeExvueZ0WXdufeyzEkOnxNGwLDo21wm8ez0mILHGolcdnSRbDwtlzvaJSvLliykky
kY2wh0t2Tnucj8ZVdaD1EJa2GElso9N9wdfZaHpHkO3r99imH4tWxEGdn943z7/kgCL6tkXqmnbg
46iqv1Em5WjIIbQQH1EphWpy1DUjZd5i7jrXOsY1fpm156C7TPNlHwiNyX863wRbZbIzdUpfv2pa
+wowx2GBTcntAIfuCLhkYWuv4TLuljx7dxwoF/RyOKKlckHuRWnoC1C/h7UCXmgUqMYgRGPnZKFC
/HgUNler+O+CL+ojMq68xpB4I5Qv7m2rxOhFKn+ejCkRuZVCgBlKl9ZBm9alwPqkPMSswjIwSTc6
F6wHoUTlBzoebNgnROUZIccwnahss8Pdn+o8xZMFgz4a1f+QUgh9ZhvA/TYNvwyZbgTV62dLnOc/
IzpJlIK9ftRid9+fk3gQgU/z4PXl6zaBQLrGjVl2yjyee0qny9gr8jTDuSRkfUNa7TYL0o/XxwEq
ijS0pCcb27D41UCLF9TcPExymgsKyDIMxxHMhmqA/r/LCBNd3nkVa+Yt6qRVUqJqvwOt/1IOksfW
Kfw1ACmUjiZYYlihn3OqMsunFxUQllHUcwLP9wSdoGlyW6REFTxUZ9Z2p9JdGtRrYskZGP0HlZsP
zx42CNle/Uh7pf+Uw6WvNfLQracXw/WxutV/3i+kKJLF7GcLYV2zwfa19GB4KDipl1h6pHjGxUz2
46VTL7VNq9fcpa3RD3t7nYVIYm6uWMTkRl0q6tE+yo0h3xjKMXh0t7MLLbAn5gVDRs5inQrFCgEh
We7zETHR5vwNsuuQ1wYM0Z3HKlI42/4V2aUmax9VeY7kJ98TFt9Cjh+huZ2m1VzmdiE6yQs5YmMJ
UVC/VqyDzBivZKSXjhl5JTVvcjQitvFHw657gcTP6dksxzCf53tLlbK9KvzRbUKFn0X8+0+MyliS
R3rjd7dBk/x2nmfjKvPgHaZFEHhXxdbRaYqcFZneM6WflC19b99NNnfU6RQksTHN3hom9pzqo2do
Dp6CWdSUktnetrXkxcnhwozxVFIOMQdTOMDKO/Lp78a6BOjmVP5ILN3kx1AkStXUfPtcasUvCcc5
n5XJrwhG/+vOwwXwlZV5Vy92zYZo5r7OQEBfgoUGBwP9dIFxSj5FsqrLtKETWJaOQTNbFOXW7jHV
D8If/KG/i4bp+6U7s5TjL5U5yLnNOR0Vioa48xplUqjuhFCjAN8dmyEfq9nX1SMs7alpD7gfuQ4R
UUIq+V1NwUOjwAxUvone3s0b4Z/Nz93066FJOC3vCbrt/LQQ2/Gi8hd3XVtzzDxetxDT3fW3C4cO
OlQLrmhvKeiH69ukScl9U6xRKsXUNn9TIYwqIXltk6wCx1EFFu389scA/TyE6uD/K3WFFQbzMPZc
Lx6oEUk+3uFlymiScEipwQ8AVqNl0d4hZveUP/TzHjZfBv1XKo3BBRoy8R9yjGLKd7QPMBBrVonU
+cUp39EDkDlbeMsbqzPE7nDc11Qx8u23GjWDbBP2lSc32MBa/5q1DNM83oyocd/cQCv3gIZpokIL
Dyla+2nI2tp5j00GVmBrSRF9M1wTF9uXIeDKf71JQqeupo3XVJoju8GWgfX9cTCKPhR8gLCJo8VZ
V2pyNzg+v7pCttJ2X6aNgNuo+xUnJSCOnGI2+p4LlrqZgw+6Qv50s+mJoiBL0z43WFZhDzaX4LP8
F3zWzbvFRw6l0RXBmptJ5qnuAjxaYywTVvjb62/kDyqnAzOJUvCl+VaJ04uo9yFWzdZf9gxV96cQ
w9PTVpk9ss3PRQrUN+zK+FB8JbpWpqu66eeWESPhlxchgb2O4ysLwc6yNXIqdVaGFC60lWCpmBkq
DtThkXIZD4pnk2WPxXfeaKdkEA3rOEsOslt0ygXaIfm3ay6uygZ5uRQMloNwVb8lqQTT+MQOdVBy
OUKsEJw3SMPR2Qvctm+Niij5Q2yBmLEKB6CJJ1XLiw45HvyYHjBE5FDAwVKgA2QqXxAPY4ovW/Pu
cXtklh2F0H4jLydTScxh6zIVqpEUpicFrdaBAzl/ZzKi+yz+q7CQ8//nxa/gAl9PubhXX7aS77ZL
A0dOstVVYaLFWZcWSWhlaPBwp8MR7UUq31q9xhqJgRHyE5PogFpElqpduR1AKdayZ3S0z8a26Wik
POGgfrKZo9jQm9puAAmDjIQ9Z6Qpic7/T6M+/h0rvYU2+OItNSRJFxdodKOCH/6a6WZWzfdUSrCy
vDqec8qmVzd684e+GlHU1qu89dZTqhk1te41Bqh2aWxDh2PyUBzbfe+ZZWX2GNI9Ftj1zLpBpZVt
CUKEFFItnYLtKvGGPYEUbAbrGd1U5MoTbkC0C5gWDIYf+2V7qWPVV565ZBPjbhUB6ndjByt6JQiS
rpWXBJrdlgVI7XXipPejA0T+k45lcLnTycry84KZtDgmKmozyDVC4X5hjdnJV9QLEybVSmkfOHGt
Y6IUkMiuLcoaxFWiwHYPH4RJB48ejickPbpnvyQECVGZ/jaAhMCX/nLyRCrtiF3kMfVP95YAEGoE
FivV4r99KWSNJdovVxYFhaxl/e/G/MHo2mMhL8CA/roFiY3GxUcL+xqeEvae54ZuOpj3B7FHJx8Q
6rHaCKkdoS9iKQQoBkSt07Oe0PnxpMaM/sP4ihuQUtmeuDKzRUb/Mid6C2MTxGnF9f00QoYFzcDF
CuoDJVyO1hfF8AWGj6PJugN+hsTJmmtgekDPhwSlVOH1MAs1Kqxm0CEsh9Xmpny7TWFLDX34TeK9
Z+13cG10Pg1R4wGpzdS14v1LKVmus/JBha0A3mQTGoZ/mzBv7AItHw8cl3TxRSeLB5ArDXmyZQvt
1Eo1/4PLOhucst0ydXBWv814HTE8sumCTfQKdozhkiw72tZj+Wm+mDUFZIkY//1uOxU00MSJk7v4
+kSpdffRV47oZlOU4//XrKolRgQkvUhxzy4QiUPJrDaQD9GLB+IsZqqyLLN1DAoCdLah/tVT4vlx
6UL/zgKnyNbUcGOb/CoicEOh6UechO+SODeVmRDz2htlgCPYUSthVGTlCBxP4AcRXShLRNlhA2fx
QjmSOaP8mI0HFFiWZbifevSEmVMZ5wowWKxUYqd+9L1jzOS8zkSVD9ueGdWe9r3IZ0tB/KAq00aM
+8k3hZFALn/1sQdVtbC1UuwpoM0i8Wf8I8IjdXoUy7j2LXrn1ABs5ZTvlp/HLDVluPaHXNhufBGH
hqfk7tZSvJJvH9NqjLHUX1RI6utu5dKpeiQziia2fsp6hTTEZDDr2goSD2LqjqUbiuoJqjgPTWg9
RGoBgH+ZhvZNYOf2W/+wUXzEe3tFdA9g+Mca9EzFnsPAaO+1Z6avdosGkNqFLN8tN044baZoc3GF
zseht5PbeqBlkr8jFrnZlngzjN5+dMf2/d8eBhdNYVhZ1sdKSQeeBAnR6HBkhAtwjCqMr889SDYg
ZBzB9yQ6iZr0XTgBV+mQtfWNRiLewK+L49K5JwQmK2wjV0wrOb3b2LTJeNUjianN2yIFgIV/YH7Q
A8Tn5SJDcjp4BbLBkUKhXUd6tYradYsm7jSg/z8YmiJnBVclef+zvSLSCQjACp+h6NK0X5+bydqK
sQfrz+jrlv5YZdcJsZi+LWntKJKTZyjvZ9k7nPqCWZAQ+yZwuiJxZ3eVkSee2wY3z9GdoGTs4srs
haxKoaxdXEURsCodhhtzJgxVxM7w5bzGK+NLEGHTn4xMLT7TWKpQiips4Y6ryy1h5T9ZKRhDqHyB
XcS6lvKZLqUCU1Sl6I4SDpzrcg6h20yl15xToly4WISzB1jdo1KrFWKKwxOkoTZ1RuQNPMiLRqk2
L96CN2VHjpSgCbTNBq7A6n7Zq3qxw5+08/epyRItERy6SEhKRDWYJpVgRVPCS9BDE9xbp2oNVrVy
8U9EbqkDhFhTimfvM04mlIHHQ3S1cLLeVA52Pa3dm29msc57lp6gA99Ff9hfMgamVc4zZCgn9G3G
vdeOUmVDa4zdHRhRGJ71nvo6BfRSYe+bZJNlIq8POOLUbTKLmAbOLD99m5ueBsGFFm6Fn4v4VsNL
v+iAJQZ4IFpz9nNNtByov8F/dL1WYt3YFg56GbUjj6nWDkLoEEbvg3ErM6iMQkuQKavvqBnrxgtw
7wySbJ5LXMn5A2s5OZJn06L4BDYcOfXc2dx+kBWx8ndeU+ZySzVbH9t/2JRjISkMESCjMphydw4w
K931+JFD7bjJXxm/HNEi9lg2C7RQgmsUBDxfKdab6dEAE/PtmNwHLhzuDSADvW902zJpp9dFC9aS
fa2Li34U7hgBpMsCU2SyL5pN7x3OXktO89m3YvV6y9VXCutNZ9fM5TmvwKVTKbTMvIvu52xeKZ0W
+wlDL1YlsqGW9NPw6WPls7eu+W+w/V2YQNqmBYgoLjmjN2shQ/0fqUBA7mcjbWGFxaTcNFAhhBFF
s1a4UYYeZq5uYB4vwgwo3/IOpLX6adazW2Ru1DBSk7W63ouJSLgzZ9H7BWKHdhOleA9qBZuOQaob
IDXcOxnNn5/l5fh2ysNWa1+ei0iM1tIJIWjfIEVjgARBVhRmxvCL686my5oxdc75hxA05tqvP/lR
CNtsmGVcbsEWkNtLmOFNzcDzosc1zWZIZCwuY/TGG3rOveIOWGhXn2rmBo6wQj0OVyGTFeD8fh8Y
NVlIoZxX7ngOHTsnXPZJBRaSVDLdobMcXjb9r0AxzJJEswQP5YVdWmRzYtlljxhloE/3RlFEWcx7
8H1o0NHVekXNKsO64SUN/RjnlCyLfkTJj+LaGB4yGSW94TXrb0Hl8GZ7iYEtbxyRCH3Rzd3/kHRE
//bEwk8jDLhWHHWgDgyXT0YAtoqkUv4LdvPh7Ea1IL87tXRN6YDdkcCk/UWcYGQjsqB91Xy+4180
DxEH2ZtM6g2+5GK+ItGfi0engZ9RJ5v7H3PZKVMALkCZ5a/16ie1UzrDkrE1P07TSJMhQ7QK7bY3
QbTZ8BLo++f+Bm839ryNULk0RhTNXIklmSX3ePgywDUpSuSEJvPXPx1/ePCwhma5f+6P5Oa3IXUI
D15tpez9vf7sO0nPHkYkw+U4TpogX87YBN5S+q2VLEm+HlsnXk0vsZa5dLzpRazMevGu2+WN8DWZ
chgb4sYqsPOJzgN1geuPnyRakDJ1uzcRRrA9ocE2IpCQ3Zjde9FOo1IuDvC8eoLvf3Vm6r0eB1l6
gRr3cbtR3zxFENo3M2YgXaD0nXVIKridATYT0haoAOcaREUMTx3FRplffXFbXdxIPlA4z9GsNABd
MnfRlB+882C3WxpGcK+xly+ljJ9vrApgVLRnTwBPZxctVP2RCHCQRGZIl0DZCvNUDtUoCmU26Gr3
wpQNcoIG4LoDDezsWkJXUgo1aCdlGqYFPRG6TLmvB5/by/Lnq+84jf722EWQdbuvl8LlJnJYmi34
47NXd70j2zXWOb7l1O0BVLF4B47NoSJS0grLqArdAEa3YUJXh9u3L1dSh5ms7ECN7vbzOgGEfh8f
zoLf3L95XwVa4EklzvfwJvxtPHY8ij2ftAoVuzi3UdfQKyGF326QuefoEaNNV0rKdnav2hdWoVS4
ADq34RU+gu8gi5yngso4P3Nlb7kKWOytbcFYk94TNx0wzr7GR0gWHUxYmjVeYaYhx+YnrL0N6eVf
zpYBZ/S8NDoMprtX0/UMVglA+RqgtK3KO98rHviGVVSpQFY4bgAGouC8hQgZiV6dXUGQj2cXQfu3
FVtuxuA4LY5UelmfIl/YfGz1e/5CuSoo2Pv25KU3n6roqdPzEqKDo1HfLYlB+/kUYudDo9P5Ske8
fhqD0QgKcdDqy3TxQg2nLXOBUZJnd+YegFXrQKjR34lzrZk50QI+MGPa1J8SLM9FTh2N6EmY1ODY
+z8b1OEKkCeJfwq4ZJLhSxpV+I3ydvC2IIiUJZ0LYIKRa3zgUjzhp/G8BhjX/xyhzQo2LRC8LLr1
+H4rDyhkurj3T+IrjWpIzEp1AZPDiSehDD9lBdv3Vrxjf63fBsPOAxm7P7el67JALK+3AElY/VRf
CHQu45gCZEsH7C0qQZadDR/ImF+Mc409kd22u5cxbr+D6AirekL7lnxqjsSPK0AaPHjkbjyZdNos
hzQqLwbyU2CVUgdSsVHOmGLKRej817STSSf80TWGNQyttMft1MNmHMYf64KSzkGlYqKd8DdwPoIg
UIHCS2YW6LwHV9akxb87g1dnakN0wby+vQPSOJwndEnFyXtkvvsXux8bC3dZNDQ/HPe/ROJe/RGy
4z80/FRdKXeNpLd03wjPcfRJkt6pO0ugKieGN7A2htIcDTHzyRpnUY74zhHxdaDWtB073mIwwyxK
AGY9iQYrsx/yM65iJ8hJL/ohljl3soeI7oCKl2dMZLBuQ7ydk2nFNr2yHRIBzNijUzemHtksTaFU
PhsPtc9ZsvVH5o3Q1TiWTJQWR25cIEZMQBhn32AnPdkZyOerAGlEHnKx2D6/2yBRTRwluNtIMx20
a99RTqyJ8f5HaxUk7AokU3zpgJMUY9wG/e+i62CWaJHFURbb2Yg3bknBb5Iy0N0GncX+sduQHSWm
HCQRn+FLuW2VguN6BljYgc1nAzZzEIL6DKlR4HCb+0Vk/a5ik+htlrjjC4zgNdVnc88ZFmIq9lFA
e1nzgkwQAvrrYBEHD8sv41dQVxbjqZvFSeAcp4CnnbaDB4T1CzVLqr/nGswbI32iO/eV7niABCYR
WTXQ4JSP0ZmF3jOZkc7EUnvdA5zagoi0aluAO9V+jydepyJnSpdnrARhW6CRutGA8wJZjr8PJ7HJ
acDdTDAwqP85CQtybyDY/pbTJ8te60ryaNdaEH/ya3uJ+4yiCrBETbmk0qNHkOxbCpf62chULm9E
iIkJUzMznNNMOowKVsf/QX3Ind2e6LLx32Ip3lLUy3pTdtPdD+BLH6IpRdR0FOxsniARmIipVhNJ
zk2BT6XJ4GQgvuZQJZLKdD4ptg1eMH7vQYkfuMRVlQmLlg4kjXi2oFQ40lpPhrzijpiIViUvsaTD
agT09rK4SJrh9hh8RUORLKG+wtrLzuBCfnGuEypRa1j9bkeOuNWV+4Yo4EBeRxtgZjgvSO5MnkK7
YoC+uC8zhrZvbF1qiIOIgxIYB+JMJHbCIDzUxCgRbByGNjQwSv0TiuwROshhJBxk6JvPO+inVGkB
4/5s2xJthKN9Zy6WxhBhrtFbGO5YMMvoIjU5Ep8DVyY933bASfznWRmLrX14fR8xAWsJ4p+AESaG
7Woq7Qmmt9XnFq7j1BiggwjER8f7Iek2ZP3x9idB+U8AxBoguVfv8Ynqv91RTjJUJ9rr6YGxvj3R
GhMvtIOFKkGl2NPHM7et+LUPWfuyR7y5iSdR+mExnillA21YKikn505Gm2g5Iir9piTK0ZBrGZjn
g/O0KghC6kboAInEFjxU1Js6Ntwkrt1+OYpAkCjMsj6q4bYAoY5GdlOIHOohiTE89f2xIgJauQSP
dV+hmwC9WkBMcIKg6IEjETx9c8VjiZagO561IzZ+RRGBwa0avNTiYlAoIUILHdU/oWEU1cCeaR72
nAO1E8jliYy9JAoFKbzEnrXdPpUWJNGUUK3E1HYE9UCCw2kdov1cLhEBOizJmYFFixL4YlIV3Hog
KOryFPG1sj/aenKHsLT6dGIBSyNZfPB6epbNkTAlEU2PpiGi4iHFdGJw4Pya5mMn5FhIbrZ0g9wz
zPV9G/PsvWp1Cw9uzVd750E6FupegFZdPLgrIO8Rz44p/n/JXLI/EZdvue4I1aN9NKn9r4z9Irpq
FudRt8wmdCj97DyJtJQ5cGgwhOGFnvxfEARfiAyoU5VNK+zWh0Aaxco08wh5CZS1xOGekOVXgSXy
Neb1OKAp+nJC0QIM5oxvASEod/iGzU2I0phIgkEqlzbgYhcvSyzsAbcsbYlFfMhz0VYp2E8jAW4J
iwONrvlCrFr/tvZDlbvkNICSUhvrupG8Sc9eaFvpYt57ES7xw7BrWYLruhAMa7op7LJX5xT41wnQ
DgfZ8Meb8SeNv7dSSg3Us1HgURLYsoWPdeI+lszUHphULpGPQzY1RTm1wBKaj41DQrdNxsujSO4f
IBW1hU7m+V9Iq6lD2Nwi5cynyCdCDh9V+1PZfApRaaGjrzbTpbf9NzWwuTfq/M4BZxMhVB7/WduI
1/OWoeFJ+5abNBhcLLgyVLcPTuGVzX4SN/ojwPa7BfC21WdBFjbNmb1MqxYItF9LvhtGlejnvWm3
mJymNUzRKWWEmnrW/pFvAo7tmCZ2zO05rtSNU5jRYDREw1wPmzLyLfhxEoJMeLzVLdWFEvHGd6hc
tFc5xlgCnydvzUfHMd1vGECc+vJhaWVolFjOSo/6Eo+vn/NW1m/qyE155jzwPEQ2Ab3ILX0dagbr
sZuQgcvLqMhXZ/ALRQt+dhLzOs3OEJ112ssFXQc2sbCJyUhNx72xeF2d09CY2No3obvHH4whSfsC
Ki3wfIt28wIasTuQ1Ns7LVDJmuS91/LEAey6R1haspIYP31qfgZsPe6A4EgNxrVwubFYKOW+lyFU
OqpAIVITahPyVoonM6MrYMk5pjnTYL+S6l37FwJbYcnhibro6jURbSCAitBirOQMPpWtxZ2CyKsh
fmwsNB6p3NAH1GGtKAZPMnPb8p1d0ZYikd0bANMHW/grSGVeDSVgYwEKQ9s0P6Tl6Pi5NnBgvD7M
EkKIQqmx8lhKGaRhVzqUy73ewaVJKYngxt49+NcmYATWxMe6s5++OPJwTHS4hfvXLinsnyEQrtTA
83k+q7dbQl1AAG2RcTcIyKCbwEZ9aSujdXCl9vQyRskUxIRGxlikZLa+jK3D3GL2nzZMxgGVX5YB
rj4nAK3w0f4UrEdNA+upILIj3A2ow/NgmqX8F/KYkr+eQlmwU8nqBbGMuTf523zx6gKAYq7GPgTZ
+KDS19mAfEojgYjllfb6DSRGR/9Y1XRnQ6Sb7FAGt3q8hzZFGt6y9W9SfdVrGyyJyX55uIeN/urV
/8ZyBftZvUzY7lDbPSbZdgHHFeL90RBVrBhC120C/JMODqMoZ4muXhnVvN0ptIfklH+rtXk2mjzR
C9ig+NXvGIOQ94JlPBUp14BxwsO2pYvON3wgyRwmWr3T4AjW2YJWgINfie0cj9LvKOgdxheRnh/X
91SMIQZvXQkOFGvuO1x0+AZCaKp7V/ZFR0lKdtWno62BG1MGWteh4nbR8rL36V7XcJfhdnRBF3D6
sjDFvUa32HZ/8gEnQEeWvQRBlMJDJuDKwmhAd073aHHCYfQhT36xNXgxcF+nZwiHMEwjFSPij79M
VW6eQGpQVBg7PAVpf6pbxPJbfkPvPtUHX4pphOKReao/nthqip970/aFeHtryZ57N83dgF3Icmvm
nbzaR4kwnJvXQiKggrZvDLw0PQ86JcjSsqH/WjXsojATDfn2ImDt997E4tHiCLi7uOlJUcZFWagJ
V1mwDthtbGtHBxKH7NTUSqpFBULD4cAAsyW1m27cTVF+Mc5kOe2K7v2+LBso98YBJDIqlLjle2Dy
Pu1FS+3elkJ/N1gajheFAl2wGtOkg+EuOvmxI5dezh0fqvr6wG7DV1HsD5KQ9QSGVM+Q1WlpKiec
maUQKJMS/UzKFnLNStibI52vkyrHFH04f30YHxnpxJIfk+xs3iTHraw2G1p/FSA+RP5LW3q450WO
OCWYq+tmItkCtrNlYsjQRX+wWKv/zTmtj6t4PlcPYl7eekwu3ChlUgfeFrCEA7hqx5Ju+YOGaatB
48eOLG1TqxtSTx23olJ2sa+RUuz68Y4bm+NB4DgWHZIdwYwhxZWc562UeF2dRUy/X4Rtv4A5H9Zl
KuwaMvmMk+cJ7ccEItKkOUaTUdceuTzJUbGreRYJ2+1dsHX3Inn8oK7ibASK68HDs1sIQu0Itbc/
883naVyBCfU7Rdrs6I+AnS6eX7PrtAE/SIP91W/8chLKmeKuORpVzteRN+zSqzOcB799iE7LVmQa
y+H94nvygTZ0Cj49TGnSd+gYhgceFkH7cQ3fRpgeU7/5bzETdc+12SHjKTh6oXMRuWxCUA6AuNU2
h6MsK7gEZjVyNbfLzJiVyfOYPQ+9iaH+Oa1wIuZw/AZsBy0cSrvxM517Ng3T9s22VuwAx9QInf7E
Njsp5jGmaQjOvCQtFLnT7DLTCSN2kpLve997CElL6dSQz8Xue8fnjthd8oZfdye1SZ2uE0R1coGZ
n8W0/hlOmbwvIDy2nZYCtXrwhysh5IrdjJrN9mrZiDV3UE+Wyj4kavh0gVVr+8zH+rF4H+NajEUM
1GIF0+pKjUserFrNH6HTDXcVXvyiNQo2tz2NIYDhLdKZ7P+ZGqadjd7ncU+DWmZYMDJK/g+U00C4
pHw33v/Eb7I8VMOjVLqgEdBZIP0/Em2q0mgQmyrKOMPC55N32GkW7wki5xl5PmivDyzCz1yaSV89
hi2pdvgR2fL9I84gFfUmYwNtMOFoFAr1KughRDDg7pQWFOcHSOD7E47OzLS1143MUBKvKtpic7bH
G2MgW1FVVIVDBYL0P9lXZ7/uNFpkjv9XySicXL3J38iegfb7TCNgJUthVh+0s9QY+Xp0J/mv5ykp
8cXJ/8UnVhNBc71ATEyGfYrAGZ1iUsQNcM7uMmaCyyRD/jQikZkk15TCopLq/0TBHVLtLR+Ph7yM
T6jnoetdQBQNuIMuVWu+Fu8fclULnJLuCPPPNLjnNivA3ju/aenhtvWbRVlNoWzyHt/rf4CIyedN
wEfNzbVTr+ZuTv+gJhPzB5g6UjN7laSb588qJFHYToe/i/cMTeEmciSZEz+REUYWWoyv9zIp1OFk
6Dr82St3fwyozzLKPqn9GuA1xr3+Z1Dhy1nTiuM6F6jfOZhFgu2dTursgFzOEeyRZc3toIxjz0Ky
LEYl/RKKZaFqSRUFMyYwJOzkXJ6jflrF8ix892UBtL9QWK3tcDBhSE76h04V5o6J1WtdQvjYQplZ
lGviuvsX8jfuEyAOkLq33TLq+7E35n/9V9HlrP9QeHOJi8QD2V8CL/IJiIlPXsMerKmziIjjerqO
dfRITXEpzGUbVZ88nMg7cXb2tgyNhlxXPCUr7cdN1nNRavfatYsLbmCOhA4otvL0J7agV0K5G0qq
sOOB8A0dZnDxiUJ/sBM9AdIzb1ZnLULpfICVHvnZAxj4sD3XikkRJLdWV42M3FYxuRG+KhJm1LwJ
vRLd6ES62gCIgHTS0ZCKPyJN2FhJWLG0YBYIldOHCnpM7GmKScR6PYxDEDv/Vmr1l6SFLcaG/fxT
3cAetSUbPnoSIDG2EQ7M/yoZ0iUEDa5DbhMN14+uV73bUvYqpgrA4GUILDtaapDsmEQJwrqy+P8K
7EZq81riUdYSM/wo7iwJKkL6rNtoM/yKrfS3I9KQsefv2pkRDjWpuQIU+OE6OFsW/uQ+X4qUrAlu
XGIr0PHWZcTwmjhkK28KLVewlJH2UfUfTP5b6vPJKnTeX3lhmIn8SNjPe2hRWPuF43XlGHevpSr4
0goO6qRdB8yvNPoV4B002/kEwo89LsBltKn4wJ5Ur/N0Goig/WCpjRHasBN4HjiScizh4ja9ZfTu
q6P+OvLO6R5tHJIYFWtGYmSjKjFDvmWh88R2XORww6osyh342qEGA9SYreSxS6Ga7ZlAjJVEo++W
8k/0hR9WyPJKrjd4gNJ1d11HtsYlxYp2QbacJeXRP5n7NckxS0d/G2uLKC2mIMy/1lZRRX/ZL3cZ
FHsZj80oYk4R3XRYbBi1Q44FWKmHTlr/n65gMbRckv+it3Cn9v8+tZZ9EbmKsqt2UTYqJ4Uoql89
zqb1pG/BXqD4WdZ33/h6NUMWWD5KU5PADLwxtCEJHN3m7tJoD30eHCtkIbKHaHQcvizZN06lXm88
yC0TPJ8EYPwWFbx0doQEzarCnNeknfskiK+964ft1+iLePgWcKkSKKv5ZUGUpHUmjzHF4SutWxBR
tsbbvsorrxaF9b2Eo7Na2F/HtnQF83NB4M8AG8BkfJVmfsIIWAKAxgUEIExGq5/iaW5eU9Fiml8I
EAPEX9X5quLwVvcIUlPFsGGOyTvwGM+BKtFyUbYeHbQZ3BE9bH4BJwimai8TrXNxs8573fuFXc+d
BaZ+L2AKFvL/1YTuFRAP+hGWAHujZXG/1q84oEGH2QzN4CnIz0Ddt4AYw9ltVK0McPLaBL5RXmWk
hYkhmYb36/izI183INBRtMPiJyZXiRqIW4AobHjaTmZdxn0CCr6BozV1VoriwqNgv23tuUKNrL7j
qL8d/x6WEYcwFk5uch+6D8ve2l9v0P0bTMBNQq2HgAF15WPcyNi8e3LFRBwqOBE00/8FYrUSin6n
GGCSP2bI4jQoFA2qLZRkc0m7ab7wxN5q4YxnKAn2AkF/Q0bmCZsAvO0kjaYuiJiWKLLuOpHZJdNm
8fyE1s9R62Ga9QNSDjlznd0PQ3nNjgNB+cJE1t2Kl+fJzLqyfprOc3vp9cQzGLofIj8KFQbEC7v3
4/CnsA0phBiV5VcvGnAlmHOOmSx3JRmR6v/ntJRKNewI76Lm4HvXB77tVvX4zN4t71ameOKUlH+T
YX5VfkRQmHgnHvo/Ug+5GxzmFjb5yvJyrp1ZNK4y1I+oVHmwSpHZ5JPh12yCGhc+Uf924mjCvhGC
RtWJKvY+SqvOPqnPMIcxhBnPJioKoqXqWVj96TslbOg2nGDgz9U1FDJ0rVcmQpXcUp5I2mynpdhL
4Ihd0FHa0XFDQZML0WEW9crzhQcFhT28xMlAOvLrRO+W37X70RWGQRBFcGGw+v6RXiK/4orD9tFm
5/EcOCa7YpEZ6edrqS3eUqJJBtrcWZHvU3q+OMeEjdEtPENFdwTUYQ5IaI5RrKyZuDeTgASKag1J
xc3UqPv82gxFiV+YJuoLMO0YIieMhp/85Tz2MzjOIYjW6YX6qc3x8quWxQwkqs/qOON1NvWLXC6U
G3lBEvc5D6qz65mppwtbc50EtafYDUsyreI9jBpNcpxIpaJnXuV/2zNaamCaMmyUquHg412F61d0
iQWi8Ewa9F0ymiRdiM40Yd5d53vTCfZMBhN5k0XFBhUCCVE07XVtbGmFRL3jJ8PtHT4Qxh/YujGC
a8As1QnU5oxnETxa9FCIWnFExThKrPcQ+TBAoka6WNDb0XXbfjD5KCGKtZx9AmZBhKcvvWh54LrE
wv67X8ieTy5cMW3OzP3ywjQIiNz41yaj7nJUU2VY/koEcgBGdRPLvJZGr4tZ3hmaVbqsStvvjlUA
curPViHLPALpxUoER1q/lgfMPzYMuDSWa8QoCwfid1/KKsSmU//9zUSdotM6lUEd7o9gTWvITcWj
VkRiqE8DW0KQc2Tpj5TF+7qMx5H1NGyomZE56UgjYpoAj3dZhBhD4FZV2yUChueLbLly/anSskm9
ioMXMPyKDSgI5N7bvBR64gnnortuj0U8vZgaMqqaraBoLLSvPsdI6hTP6v6eT5uUK6GG5Vt9HV7s
WvU6cGJpGsbeNADixBBAb0NdT4TBCeCGO0lBJGTrI/Mn47PZyd03zwmWVxtUGcGxwOdQ8Ki8ctRH
tZrLs9E61GiBaF0irkMPS7iY79KQxrzhXmeTS127MNfhtP3s5yz8PnUI0WJeYAijG4or7UOlepgw
9d3v1JOnqxZEu1Asy7xQOeE3jbWtTMecW6qzotGhjbyAIWHAmlZi+mnBz4cbZHQpdy7ad4GLAnPe
lwo6YqkK0dbF/b+2EgOT1wCPWUW4XFOx8XE29rphwWdBJyApskOCCJWGIWKjGZMS7oJvmIm9Cgl2
Z5FrVe489qHUnNWmg3qBbKttN+XtafwxlEAVSq9m+jLvO+PJQHwgILSgitkz6QIZC4RZH86c6IGv
r7njQiTC39fx20+GRohTwWk/GnCUTj3ExGCLgGEAJjZHIZTE4Pi2BP1BdqbVDCHU4zDmFxqKUJ4k
DEeK2rjkfg6+erIinHQh+Re8Hd83HzmeptJ2xBq1ilAHEQBqONnoyqKv7nzxof9Ms9xIILh9wqq7
gBwWB5egFkwd8iU5au+JqO3imwTikMt4iWcR7mYMVOjeFlcccR0CcfDixjW90Jndcr7Cbgll/m/p
dT1PyDOvwINKpG5MJ+c5RdCJXm9uc52EfWe0zks/hg9Mty/d5FtI+jY5ZEuJx1Ahf4yltlL4xC3l
0VQQLlmMiVBKnzdgmGk29z265015vTih/Z/PM27amxwgemtODJjSOKreRHbOoNlLJGAQHUhfC1k6
rQmCL0xK0JUj8kNw8LFxNtdFmHcznGBQkj4NOPwqnaDf5J0Dvmz/kiLq5biUxGTDyfE+huPP2vc7
CHABOqp2QjdesC77fU9SUUi6XZN5HdzNBQV8z9rW3cRqR+Ox8XS6iURctsJOuDGEiuWJb9ovloQG
N13Haat5XAF4FfsrfRLwPPYGZD19ShzjxUwln+Wm/70MJaWfplGIRwuSYVmEbrCQBYkhPElvQIgE
QYhl2+pYyNXdn8BqEudaEwAaTvq8iOz/8tnEYVMNjFLU0YzX0CM3mSTGVWs3H3NeZtt9yfLIeOKv
hDNpDVJ4j+vm2aFeYyDz0T//qwSgxyP/dD6V8H3NEsnhMHGd6s78hvro7Cjjj4pips91x/CFyxkS
ooO+9YlRBm9TkMpKclBm4ihGewGpKZMAkVAT9aDRr+minkmxUe45/kpS1X6E5hp2ORXuCK3SQIB2
1t1z+fF3FGp3iP1J0DpYiZi5QjfqDMsS+p1bClBl4yrIvD0dNbJ106K/ShD3lYNXUb8ZONgHqJzg
typoh3X1Mq2nl2Ga5VjRLpXf7l9QcvFXtFSY61HrrtiFQAzTyWVEjrT4xHTYbjqK7Ml2El6pko2/
uZT7AKc78S2lSsI/xRVmcI4fFHdl02Z2MWN/unMJt3WLsF53B9eChvtFtR9vOGs3QZsYOp/0vXNh
q1aX4IyPOsBwlPhAfiIneDQ/n/pUVKnSInjcWWYRs06aWFdiGnBhsNyqOp6lQmA6RN3q+NcPtr31
8nwvozBQ29t6WhB9t0a5XCdTGQSCK9ZfErDJO1FCO3KcDgYJv19tLYBpBdukXls/MiQS4H0gUfcs
7sHZ/L0/D4NNGWlaMmGAtRkPe0puZtCSue6HpvGj9Trz+O0wIv53Jmcm8dr/ZpSxY78tddZ4PkMY
CF0YDQucSgtBpYSltonHuHSwepfy1ejmmGL743XR5JtHNR3cEthGYFpRnrBdnrlGE7oa2G40SdNG
2zNkOqLB0Y9DS4Bm6b3aMil6JOrpZ9U72SmcJBYgy1AQD6qAEYwL2lmN5spRbPJxLmTSouqDoLY4
3GXyyoa8nN7gBTKLBU8nSeZZCt8VCBBOQEOpBf/bB5PauaFthfxC4ddQadYajd6ACweaE6fjgF8Z
GeIZ08VOUA3+cNOVxCaZw9Ab92A1T/NIzrFlTr5ODLmT4WKaEmvxKJxNDRlzoceQLk7yljjR3/7N
IoksDoYsG9pcWpsr0L4v+cmqC6HcV8h8mvczl6gzvWCF/zmIzXhjqQrmHcBp8/Zrt8tmqqEgyad7
DoyyFMNpb4BUZyahlAkspxCX9DcZz/p/nN7HOeMo8MT3QnGnF8Za8eqT9piETYVVVLWFO6YwEzs7
aL7brv0eG8SqNHjNhw5ZG/uoWLypuonWl+Q3Bl4Say66e8UcfL9hrLAXurWM2YJZX0iMnr406pt2
DSJARxtodME5gkpkwoDg3ecIp/1XtvwfwZSSvXBHnNOqbNwm7ylbqrdHWr3fNMZpgrSSW9O4tZAJ
AHkXsvkgT6SYjZ98G1feVZa9VXUz/CGp97AqJg8vALCSlhf1wEiq46xTpfZB+vNjVmCsqqk6Wy22
7wZYw5S3sbi0hL4ZJ/9EVcq2oIvULDOOiNU8WPqRiTiRVheFxh8V4pef25JXohju1XOlgUxNVWN5
v4urFIuCmxKtwnASZnE0BYcIQRmwOSiBV99nO7lIN74h9gZ9+29QaSvz3r0/t1vqa3MJt3mJXrMI
sWPeg9rKffiVrTmeKpiApZOcFMYUn1MVi/lBj2eqVNMRnY+eGQ/0y6l9mcEbZKVJJyd5Jfh8EaSH
NYEaYNZgNZ4SWbOb5QUqP1Tkv1qiSY920b2UQe8vTeSF9KJZaqQ9NwIMcF6YJ8aDgYzm4a86ThlB
Y3dr26AIjtjU17OvFqc7NgIObFc4MqLaICD6tbS0IqwpWFhKbPwmPxXwSs3fdzDOr6nq+jcYgudw
9iYnY3ar/7bHGkyVid5bGUjZTV6On69ZHxuK9Fqu9C8eZ5H8FdFp4FO9+2OHmOBgV8yV1Hq/wyTb
FGlky/M7vz8f+rbgPhYkS7rzGKYGK0KDYlqEkKk2Dgg3YlaNUESgZnF4GBOOuHzJRYf3ADmQnq3U
KS/SNTTxLEMTsjoQvaFc8tdU/eiJuhfGvClUKILbndpIOoxAAiauJdPtqUJIuUARXgzWc5zU/4jU
UIEJ7KC6soEP9d8uIutStSVzqb4ofL0TM9LnzKJ5WQtVtILgueIOssaEnFwNCYSjY+uh8hxsp092
o8bUPWpaLNQw8GDyPAAfsVl3W/EoS6ZLObak/sA0Erw4e1JhakZdQm5jrHXb2jEGGt1avW53EEXy
LMfMY3OrFTVAAGthOp7VWdIv4UqCTE+s8aI33wU0a8ak9uFBNR7bTS7AOBoprf960iCnBxR1zAyG
cMMjk5ZE7dptrN+UIieFqotS10RReZK8hCfl/rxbPM9HGZ5Yvd5p0DNcAw7/95LtQ1iD54BVUMNc
Q4AmshWcYrOnXi/ASiygpVMPezVzOtR6Jh4bTARlVm5+isHKbVHyK1UJ23DMb2w3XDshYFWy6FdE
DsVaUq/kmycG6gRuniwTwp3/OsFCwLzXvVdvP6VtGjlTZW9+0J9+BzZtpO8ki9pVLHZLBlelyemM
/0zW7JvsSi49vz7j0fILGLctvSdOUJ89jiEHHO5QB+9Su1EXy5hN0L/b8TneOV6o5EDGBAJzh7uA
aAuU/I3i4naA8Wdz35JPWcYGltZZkX+G2keWS794IutrK/vyfzplSgeBCCUuOVKQ1BxVjWlsPqIw
FASQ1DSJIo6jydUzm3jd9+fjF7qGBtC1b0wj4BxQPFX4ZA4SR5+EpNyGLbeINjbJeBt7MjTSjucN
61aNK84VWbwxlSQeN290uJ42hx0dV8DhlDaHBysWFhXOauCXRoZ5A4phgWGAkr0iIVp1TvGkEIj1
ExnZq63GpPfNoFHS75S/J2adwAXBfbXFK8VqwfIDM8jtnJsvEItoI1tJ1mcofGCbSkIcVVKu75ry
ax1IIpd9ey4/E9FHJL877oVxYYxvtA1Waa5YO7pDocvV3GmzX7tILVrj+STtQOZ9EZkWyIpGTRwp
Aa+p2OKOxWEvgMV3FmWeYVPIab4BZBy2H3nry6eTU0ouIypdhFGFpqjssuU3wx5mNz35eLbqKHMM
CUIGT4oZ9J9QLbhnBaX7zymypYqF/qSVqr0pYcuKwql504estHGyakWex/o4bhBpBzS7ATMMIQxr
36Y7hyR22diTMD+Jx6T8ZtMzIgDZ5pUVl6FR+DYT12wvbniRo9bR65/+6dQj8kigBBbsyvYkv3WE
efhjKIPtdYgdGzGc7MXgH1/0QvFhkPC/zn4oWE4zz3/W9NojlnjbjiE/acgPpxBjQeyaEN8mgLmz
X9FMsbtKx13nuR4DQfVlITICUmyDhWyiSQZ4yEy/ueCJkC3SKzdIahLDc4HTbgfj9fJglx0JFYmp
arNVxQaKTYM/xf5by2HAP4lZnwTGr6w22wc1smMNKwPTzJ4i1g4FT1/lz/EFt0NHla6N9sJox0K3
r5fYzt4EFHhatWd85E7PeXRS6Y33fNM9woCUZnEuTauyx0EtNb8ziOEKutvlvb0fyVv1VqDuMW2Y
QrQs61emBR7akMOXQXwrsUwy5MUpSQqdQQoqD1mGRHsEj1bLe0BhgxPl85JtdDQT9t5z2+1A8J8R
VULcdj5y+DAI+0KaWkytT1HWk57WytE7NFQwmXahBNu86/JLcwfRlnHTJH7kNVTjvFNHGg/w4xLp
LdZWH4nnG6SDqA9VS9sABAmqj+97U7UjcNcgNZnKAuJ1gOJSInfcAEnzz2Qxmv+EoE1lLtW9tbXm
Y97kDYGsGvBum0pyDidnejwlnMLiR6OXJcWRgqA6Y0TdLcaesR5mBH4QxTC+uWow9sKY1PY63be+
zIfgNG+qGgANV9m+Isc1uK4niZnzNcav6uNfcPGsjczC0dyW4iOPNCJjniDQznunZxsYflYDQ1nK
VCiaDKnc0VKLPtGqxnH8t8Mp6tp3nBfGm110jjseOTCyRtVLKsfYGPk/AksG+GA2wdRjj7bH+EqI
4vued2U4wf1ofyzkA0T3RNPkYcRomC9A4wcSmaWxICW/iLin2qgvadrr4AxcL4uVbHkws1eS9zgu
Ke1rtJh6hKpD2hSrWaJVLtVsMFJYe/4wHWm1EBHWxn9o5wsWXY6aPJsHta6iVxoBClRws0z3dqRw
zajR3ar9uE6Y0KjZB46k2FjCXR2N/pQyizr1iCVbywdEIQkTtcThTsUmCVNW/7zMA/BCAyOXqd0N
2yBAZk2lhlMwIs7BZ+WTI4X64Zfg2t/Kx+PDzrqfrEk+j/8n+APDzi8lCREvV0z/58V1DtlRFkxx
gnlmcU/vu0asORD9+xlMCR/tJKFwuVdR0ZO4D+mPEfK+YMgjUij5VHCmxvwMVkPATvcOkDE7EAH0
rJa1f2Cbn/Y5K1O6NCBhCS+FgOsMcj9E+QdJxIex4PLHIR1gKDfEMEjQMUz2qZM3INzN9ywj5MhX
KCkvP7xpY2f3FAFzW8Qa3iYx6TttPuHfyKEp4Rh0OuGXe01rQ/K8ie3aF5D78+v46UJUMcXCIyTu
4O8pwYtH70g74hBDYp0EdyNjXbu6d/XgbBT8IOjI/M6S4cL4HkHdPye7nd65UwFonjiYYUP8wCte
sdl+Taso64zrKXSy8ovqixBnlIPh8P3hZMfOzY5Za9PK9OuTQsjoW2ACBluacHT6kmGdMT5tt2gK
X83zStK4u+bB3DQyo4ihYNQEVMkRWKp9fy4pZ+k/jTPsQKiHKpbCuq9epc+izwSJkaAhblO4kL+K
ARvH5tCbGh3DTNJePRUmJz2CpwxtNznBUS/3mlNZOETkZMdBY8cdwpGobTbGwRvNkRBNQgLBouU5
hS5J+H/PBwyCDUhR0/7y6pMh33aPZQg3P/1TwlTpboBbQUUiEiKJbG2NpPfs9LuykKSiDl+zYN7c
bpQDVJKQdKTh7iYlM4DHOeTHHIqZhIWlkjpsD1TSM3NYMWsqsm/P7TrwHUC4g+vyFH/dQnSfoQZG
OpjY1PSDHs5c5hCmazXSXcrGpVmTiu1F9zktvGXu3EPeArUTEV2w0IzkztzNP1BaQlMGP3RM1xq3
5kpnmP1imeBvm6XECbX+e7G+oOwumdzolRNyS17OP0guo/Iqf6XchSjOgNj7az0tTrp5TKpBZrZJ
Gl2nI9dBt9cy0Xw76AY1pXj5vjcEfDWx3oBQqxGLckNuY7Qz9bt55ZPKr/Jb6AyBwjcjiorQ5dbL
PIiVO7IPSI0cHtE8Fh8h4ri4YDU08i3ev8IclOYJlEvEDH4cb8Ba/NXXTJYtezOhMJcyKBoC+cmz
icS9r2gvvljKXKvClGFlz2SdoP6z4cNbeXssnVNGR5e9pvP7+VhdnDKteXUHrwYCJ8I/Y3CKp0ZS
FSyal1mcjX7PdDZdLCWkoXxGqh68krTiFu5JKdYhdIQVDPlu9hH2QdKTkOMZ3f9jO+JSM3pdkfQt
Ip4Ty/xuzO/kEIf1XFhG4K7uRzRYpWM8eb0htxjKdVA5S+jPOMe+GyAqzE/my6j/4lhlEFc3bjjS
mKhMmv5NuwUJrLpWq8ZOj/AripDVHutZ+a3/FjtbLBrSOjdjYBHAivxTFzRx7kKsSoIFy1+BggYX
vXyf8+aR5L+WFHvH3ClzzyIZ2qKiQ/jcxUICnSc3MYsDNYBdFEBz2MCeCDTiXkE9ghzdw415/M/n
hU5/NDCqIS3CkYLr4vJWVL69F+cf7nttsY/4ETZZ14Vv4iCPfRDtuU4FJAfY64ah2YugaqoC07oX
dF3IEzKrLRhPHGGVEG9KhzQd65ehv9mV8i+fjoiewe6cabNWkGaBBeec6fwKZ+RuALZmmHaw8u66
yWo6IFuWpfJfMkURy+X8PfF7N3J7onXaVwQUYWatgKDTAwoh9BjGRKbKkDGEhzOjXPkULRIhbi8h
9+uJVbyRlyJh9ojWGLssP7A2CXA+/w2MbkxsgmLYLkhubxHPpXIW7b44pFXxcMsWfEoRZdboiA+3
z4hQqqLhzhvrYTGIqUtIBYbpa1lQT7hrzSheZUMjPbem/oUXZ+rWZisBTdKC31FCiXLZRCZQec0T
p/aVRSe8+wkVeEGRfgiLvc3Kb9kgKSvTczno97kQzJM2HN2kQJB0uYJYC0ZFYF1zPlvIL9cZ4WoH
fTuDO5uL/6mjcH78t821P4Eb3KsmdKmOm8xekE8tTM0qxAHw4XP6sz6zGnSCe/QzuteMlrJ3h7bQ
VuOD7kylEA2zFw6r3sAGJaBGyhrwhTknCyHeeF8plD6jKcwO7XlLJsFX0tBzvpjVrWuqHLd1FRp2
retOBukJst9CHFb6rJ8F/F46+sHBy0q5laOZ0uAQ/Lk/7JbkgUM6L5eCD1do2URDBXNZjZ4QIOE0
RoBrbcvEbTGS4Tsm6RGvnETf+N2nTAbMOhCpNqq/p3HAmVLI7KyOVBMcGdf86Ktvo6jflttYDDaM
PGhBrEgW3ARrRNaCGAPGWe87K/8O4+dpgsNrnTDrkvgqsM90kkPHgFX5fVYolCtsv70iDPZ7WBHC
eO5Y6isJeDZp5ykyDkvgWNbz4sphVfOXI5ETqhU+mSJe+HKK126d0wIw7d3a3gxWHc62cYXWYBcS
t1p6vdkbZq35V5G4YimdGdJ3I88TbstLwyaSFJOtqrHzJE8tk23rK1MBmwoaV9U+RyNn1HL75qVZ
sDCGcib/FEVf2NMiFjFyanAT23UIM4/+baOgda0FY8ip1n7kXW1O4l3BAlV0HZjLq5yLon5+dxws
FqNrYH7fzndiTctR9MSM2CTxcgkuy+6Q/yoX5XJuaT7MphVH0UwOF6n45NloGd6R/VnHVacTw7gW
Yp+PF1HHr/zQK8b1gfKwfmfQgHOfXYxWQIOl7KXmMg0Jygo1OzD/1CIoq0XwDLyAQou02lWP12CA
uWa+lIDWuLnA18xzqq5QTHUty+5zspBvoI4rrRag/ruQjiI8Ka5Frd50SR6RmZdGmA5HMlfaEepQ
4+cyInlpFFvtLJoqG+cqqSkWFqr626u0A36HpLj9lbrLlASqzGnR6s90Z13SKZgFfTQND0h0eJFp
4I+LHvENMHz5rMiAn7jbOR1BCZoW4wS4FtIQfoHbgEabkr0J7aBYZacVODwXWMj8nx24lj7ZeW0Z
u7qAXSTyqK/KnSoUbOlAemuHYSGJQRlTV/IT20SztOdStSbkyW4MKDMQ3wT7k61ApPrrRThOpsZC
g54OHCP8uLkX8E3qz6j7j7m/GiLdkRFWSUfyJSrIsl0m8aSU6ypmhfhHocdCEcQ37Oh2dzAqBuhk
2sUNMdgm1gALIOFnSvOE/EKJ4rHkSZoY6Ys2vD776pi2cMrrLVI2Mx4oDdXV/pNHBfASYlEgMB5M
YSWZ2PGe1lm18bkQeZW8cZUZ4/6QNopnK+AmciexW9IQVjYOhy97Y3mOHkjsqInteuBx+bq26z/W
Z9zweHeUcE9sKyNVZ8VynUGaXotoJMFp91lXL9l2I2k7vTdFh2fOeMufCcmBDolNLA/SzMiMYoL1
JawIwSDlt2OTLBKx30V6Gkj6CJuLDYpVXr46WwQJXGh5J4LA3kA6WYbzq/+4yIHJzobYDCCiZ/Q5
g7Q45jMkaPB+flMHAffpSesxKvdJvIJO1AyZwxJIUXJaNcIBawtQWyeXEV9cP4PcG57UIwUOlNLf
y1DR2Q65j4g1j0mF+eajv9y4y3cKxYpuQ8ALdb2nGR62dNG7aVMuMFtwYNk+MQBsWagNryYPuP9N
/zd6xQqb/AXw/tQ/CRSK7XLntbqs9ayA+CTfIlxc+3Hbll+nvlSmNCr10BlA+Oeb1vre8DJs/36e
ykhxz1vifDQriGHOu/AqRhMCe9/YRGIgcsLtwY3/fKNJf++fkKDtfftKvUdLUvi899WzSTVnBsa7
Q+7A4J8gFmH6nW5ZyIhIfpYMmxao/mCk9dGUgZ814Zqg/SJaR5gcnXUtMZBV85qa4EGv/poGGX+3
kqXOykKuJiefoftQ3AoTx2kWhnE+qhuby+El0AKTRxvx5S0IC7IC6/NENDFGQavVNd9W1ZuDlY/z
1a5Yn8/MSOe+Jq62S4fADu1qcWfST5UAylHimkr8rxyLn3edUYpUDdKzrTYlGqxcYGOYE8QPMhaJ
Ied34BsYjVOWg0deBwvagD2OGg7beyYsQFxpeIFz/ZPvAjpM0tuz4OCjadfOYsyjmb0ynlt87VJf
NPYaOmUDKRF8rtd4JCLzpagWQOfXmiZrdZKrj0VsS+ohW3C6YLWDTEtUTvQ6OD/l9GI0TKbWp+9O
g/sS1GBsal7xsndLx/2zD/mxXnEazv1EmcJ/v5zQWecFUu0A44oPhtGj8RUioUdUSaOdCVaRPi0+
mhmvhHaplXfiPPhjJLledGkdlAPj5lfpbkBtfuQKJm7i9js+eGmmNb3Uh/Ty2EBgwNAP+hBNT+mh
Ya2/20h2DsfAxhhhO4DNLErweRV4aqfv6/p12lGH6MVvzIB7NeGz278I6Sm68Ie3utTCbQdg4tiE
QOGpGyKyG/WYJHi/dTWP8WBb/xpUaVBbaRkc90SFNtiwcA3JSzI/iCUOyUzgJCEdb2klYFXHui2Z
GzDFKIjnChoM5YQMdLQmC+tl7LvRQXeWpW8DPGHcVcy6LcCnq2BArg02MPy4C7UOM2IBnWx/lt7j
DkhQ7lhhmTI1XwF8vsh6UkP/ftP35slKq3DyqDflwIChh79E1y8ldD6BBDd5/gAeHxqNYvIP0On6
L2Nu65w3BkCJCT8uzA89K1duyZ6HnyKhOIqvevdRHg8+RdmINKlM5i3ztjHFoEKfK81YnmSpL62R
jjmcLFTQz/aSplwdrHuhRleNwKvOQvOnSphmenhEG/KeFyhI5puVbvR9SRxScBpzPLPT4wAh5cE7
IyHsTkct3sCgcexAGr4forzObO+8ZaN8PacWQ39vhwE9lZkqNc0pYEaOvudV7r0B2q+jQV3a8vwr
sOrZ+0+fOVtvJiQHKpCzsu6qTWVOE/Pk1tnINa/MnJPFfGdOG6JCfuPy+yr6YunQWZ2wZ27ImzWM
6JM3tD3/DGLN+gz32Yv1x9mKNutI010BPpfI+sz4zMQQdc4VLbqBiVj7Y1nf7AUwa2nUskMgaYhH
9nRPFs5NzKncW+yc0y0sSnh21yMD27Q+Y8cJA6TLM0igcKCRJd3jXalqDmwVT7ADBOPBUcRyNljv
gnDa9eqRt677i73mMUfdWG3sN2ORZvzw6v4+VM4EhVI1GA4n1PxDOxuZJ93MHKpxcFwsjr2T/Sun
MFOmZ75U+NNkJF5ANHOiTTTDd+1xze3swRdDOLGcsqYhHx1UMhItysTZxrWL54MscJpYYgBLcUeL
kCghVwcB3ISJ+4Efv5XnlJVyeualI/UoJFHhnfFTfX1pYgGMYW1MA6KU0JdfPhKUW0ukKUDz/RE7
iQySC+osfzF2g0+rlwCF2drSDjjCTCK9/+R4VkOdLHswtHpT3rYuuqI56M891A+G8h8syuT7IPTx
Xw7nSuNhM8QYSBN1YlDDzjnfg1BFxdvHeWt+lB7dgqSmwwFd7WS3iwJcRtdkn/V2hOJP98mCwWZ9
67t8DgSHMabNEK1m9KxhUZCQwn27k1I8TLQElXNOS5olHZqkl7Pe0KJnXt1rQGX39QhkB/GbpCUu
Ke5aam4fnDLfiTOXFaMnk+Bm2kBMKSPQO2JJHU35m3SRxD0O3hpHiS2lG0kmvngqj5tlntVvWMdR
m2KLCZQbK6cIfSzfp3Z+xt63PGEr6cVYrIhtstOk+2e1/Lte7rkzGaIeEZvFGwypZkmYGIPixB/T
fD+3s4Ar/rq0oMlrpNiSlu5FgIlfc00LQcalamX5ldxPpp0y+rJvf4V4CvGKjokchkOBxqLQGzen
UxABg3V+xgLdMhbMNC/NEF7f8IpqlwRtIQ0CemdXMB4tIYh5aNMSQYkeVn5+hBD5j93C8cz8Vla3
2pAyS77cCRbOklA525Yu5YlXFwWeY19+PNxpaBiKJvXHovab0lhqqSevJqw48gJSTVqZ1KfoIlRH
64N6zv3z+qqa+Qqcbrvfv9J1Pst5+5PSrfqQ4852qlTD25YQsn2gnmL+tZEYLD46MZ4AjNnpzV85
iuWn9Dwzrc8k7PBo2lyHoX/K58yO4kd2mp3a5cU1xfg2Ezh8HpvPKXVAdllcYBzt2ZWBk26JnoUm
SJ1zYyuXUPEVQrg8fhstjACmL9/MwAalIPul+Tm6IrdwMD7011AoHIpq9OfJb7NvFRRWUcFGE9BE
FkuQHUxihOib5h8J51c59jMxFlk15MU9maKnxEK0/TW0mL/oC5D9XObAJt5QOwjxETrBifrtCFhD
57sVzG85vczKPJFyN8FbcwrpfIzzwm+889LdKXXKAdjtv7Nrrw6WQMIzIOdVl2eWTmSzgisWKhAD
1GVCU+Dc3CRTZyeNtS2J4FDh3f981WnZSbGIOGyYA7VSMPKxTzcaNiKfqYiHt64Li8uQluvZoqL4
CNNdltZd3Tml9XxcoCvaxBTiF87DQJl9OOAjTkD0Y7VIRiohJ2BuDbym7rSxion/3YIcyYOBLhlv
NBE02/mDIdxLD2frVB4tA325Uw2StjKicvp76OdWatRCarPiYaYnTmF7hQqcnrA636iptReby9pM
y594bN2/jKIIsDvqp3hD0Rmlui8KoPIk1XAvgoTo2YdssjgZr306ki0vx48xXs/qCuy6bB9h1qQ6
is+K+CuaZl7KSIk6z8N31zEMYCK+bc22OJ6k2SHrP14+LtDiaxhpBVJ+rx+UdZzI/OSwh8E2yfwh
vMiZHwp2j4E/o6zM+HrBvwwlf3nTnNjEDE0WESeo70UufkKB7EpAA4mI+RumwYySwI3l/Gn2zZ2B
YOZzxE8QgN4TKVcokjELyJakjMUx5xXeVHZHZxKZCA9K7De+ojTJ9y+uctwlB40EMsiAuAdyD8og
WcmFfSuq02L8e56/X6dg+jfdyAptaEEr/pIZYh6iRKEEj7NyqH5sZgxSVF53TVFtyhgBLQC/4VNE
LRuWFlCbjoYjGpb3l3XupRJHN9jWclov2fq7G0SrC8nyMC2rbSscChgfrHJGI5KHO11uDfNP+t/L
ugXjFvNnOKEvqb5IBPEJH5mB4b8biXOtXp2cgPP+YJz+u5Annsx/OuaKDmxm+C+9vPJVbySvP9gc
O9kUGfYDCXfeRqjTKICT2brZjQgz2G4+CZ+GanjkluY/AlZoHTNSyhfLCYqSwAsHH6a+Dmmf8VrQ
951+I/3zAh1Twhhpa1GFt8JVQnK4ToPnv2s4gDlIH51hUw1erZ8v2uQ+oQWnFpkMKq+RowYfC39H
H0cWjCtxsujBL4LFy100cAjmT/g4GENOrZGTiP3qFLrt3B7KmoirwSi069pNbZprNdeQfUcSpwWp
juxyMPsVUNglMlP7CzV7hctXuLsIyIGmvU5JnnRlHpiTsPA+gGtf5C95HD8J38av526l2XltIX1T
w8TOOSeRmaJm/gMii+G2t/SOfWdgT9igfWzce1wfGX7clQWthfdRuYLEC/Lo4zmiMglw9e4Vx+QY
eo1BsBvxnMd+qSnggLzg3U6+WGgtP0eQ6hq7vpP5zddr/DXXzLWFXIjABAJo3OysxCwS/MPEgA2m
UBDdF6KAbgb3W80/yZFxyxlpsHn1onG0QWprbwC3S7kGQm+GYoDlNA03CRMGtvQ/wV7Rgwl/I4hk
w/gOJbHtt6fMZa8yj5sDAwh7el2s1E/kmM3CfpmzDD5zzp6CaWR0lDlyY/kBj1C5h7Iix79sbJBb
H/2MvXV0OEj9316JkwC0G3169kkBRrXmX4ZtxUeC2v7Oy+DuAZPsj2hWfKQENkkpnCIPtnWiyRES
jlyN71miiH9K2r71OoCMkyOESpqVV0aTagFHdAGOPf/Y6tQsyu5vb5WWTDHwg9NS6+dicWO2GbkO
G9bjnZ+Y3spd9w/9a9oEpaWhtj1hMSkl/PL0ea3Be+uHEtaeRYbrM+YD0hZUaWK/ScoskD4ELE1Z
TbIIWt1tN3Xl8lWabUq4fCOcHSbZC4NgQT+xXQyTWyy2bik+bvU1vg0c/L3/yvJwI176YLVFeFIn
Ds2D/OJeF3fYWlEzMeB2T97Pqv6+FepPIaMbCoumLAmf4iAUmhmtaU9f1w0hW4COpFM2L7oOd+1m
WcOa/5R8L05T4jiQROvHYLEET4zQVbFQo4WrUVYfSQmLE+7lW9r1m7W5qvofPwdph+6X+grXN0gc
boYF3i5f4ExknFznfb0cGLG/B73YBEZ8iqA/gQvb+RVuQwWUtfpUK7Junm+I2CWpKSv8umatKfkf
mw+zTylVXHfIhva7pIDaTDbzQqj4/acvhIi71kg9O56VW3gGrsUZEwwm0jhA61oRc3VV2ItvxUNh
V7f5mA/5jOc3aDsp3WlgdWJJ+PQSsJEARAMQMBZAP7fgcBoVB5J1PvrDw6pVqv1t7kiiGaNZ1hwd
7m/pZ2ewKDIwYVZdyfKyYxFydYgXwwWvY9fHEHpuqfUUy+tEpifXJqLchogRiIFiiMnN9PgjXdU9
O58nhIcaRqXhnwZt6Wigi5mACeyF1HVGTKLv6Z94gsmsibWayX3nCw6QSYHdCiGFky02YA/DlovC
ua7E00i5Yxo1uejHukTEM/y523Iw2dhCHXfwLO9u4jpsEPSqHg6fCiLBZ6YCAsIvfVitkVAu8yZV
71ilPZzrhbXBTDVNFvcLuiUf4LHo7Hgg+b8rrswGrhd9X1HCBKVl4Vw5nuPpmPvLcZdnsJYspW/6
PZUvtm99Y57OYpL6IjUSUTf/W4XK0MGGdw4hdfbIjWr/ct6WDjl5F+LAOn0qUE2Vd6psopK6Tm0o
a1GlIXNPftZHtmhc69ixSpGRyTe8/D+Pi+83/5G9waofkvRsxCrU4Mwp4eopC2gdbnGeyF7o1VB5
lGUoHht9XiS9cIYRXABiW2hTVj6qi7oh95E3z7Me7FXaSvo0ifQV1CpyBVwkRAyEB0VwDBCVkoIZ
GFbbY/6qD5P7EjPGcZKpb+VktCOexwos2lxD6rPRaK5pmVle4ArE+9tIMJqOaCf2lnzx4o+LTiXj
3iUGXkOpYdcwRkEl6AXeOuv3AAByH/H2NnlneFd/9B8ccme0AEVHrH7rMtRzutDhLd2gE6SCrRMO
7Tj4kGw3QRCUQO9HqVXJPq9AuEmS2Spifny5jiMaBPEOnXDFbR6e6QVwRRI4f0q3KQrLhwzE49FR
bqsA+vzo7biRt6PHHc7wapLR9mAGyGfbtWc28/i+uqHsR9vAjLVGVGODzzemf2c0Wnh10+c0JxSE
WNZ8xphKBZ85dmUbt+uR3Iu9GvUZJY4Nd5HtNfESvpvrkgPnGkFHxeKUW88ApcmUvWNHe60rLHs3
hJGtuthIKy5LEHzLBllVBzqj/Rl6fFFlW66/7uJ3XFpIl4hTyoaOJaCDD0DmJLsiU3KayrkOqclH
vGPK1wsARBIbWDapMqNfhFONCZiVvxzaLt+AAU7ioaO5kXVVZ6Tv16zQoSZDDFMZMv1b46tlZE6/
m7KgbAXSdmqYa3shWkYyDH3CVnWnQdIZRaskOtYNBX5A04cmkVz1/xkhRelexRh1flmYyJjuv9y1
YwAiWoP4kXyxVx51CUv8yAKhBfxsT8xuuszV4ewRsodMraQdqwFH7s+hj6GO5wkfQysHx72QkeAp
NY4pXxTLfA8Z4v4Ei9mguIV+t0i6xJYW9Kv7b4dIoZGxZ0jUuYyHgjYi86QjdpydYd98q0+Fy9GS
C6oeihsVcLpvxMWN4c29k0zJNRbex7/b6RVPI9XWxgnZb12TU6EXE9yllm04X6PNZGkZOqRybJNH
9ez+mvwyFm89n6N8nKYfSXFft0blYiKK7SDRJasqtw0lPioT0BG/fLDrtKYR135mHNBTIcXS10EJ
wXsPKhucEl1Ed0iWhjCTtGr/aXd4BFwqseo2+uRO1ueCWd4HK5eUnoDdX/BDAAiKxsWmWCZuKD7u
7r/Qay53L4FiXPyEd0aTu5Ndf0YKbvLPo36kqgpU9r+8AJQFL8e4IA9uRSXl6Uoyn6Kx4AYy9KQl
Thba2M3bA5BF5kWWKkbbooi7C+DQQR/ymRTbg3lmnD21IDIFb6J/B2pYBQf2UKhpWPjDCMJUZmkW
D2pSWGlZPJLXCBMZoF50owA3NfATZasz6a2cGPF35k8Yh6QanxtlMRT5sg/0SIOURsbhEAQoIJpS
TI2BX3PvwvYV7nYzWr96TDwYVyZbhOoT+RpMyPvxZt6xj5uSryuqu5NN3wxiUI9ZbwTBS23A6oj9
LNnZCpAThJv09Dcqpa+Ff/e1Pm1CE9P6bU+00JdAaubBL5JSfC00Pu9R8Vy4M4DawdCGS47+j3iJ
f8YZwr8VZoNmYOB2bjlMgeWpVHQUuzo9sIM2YpWmH4lumru78MjwUI0CV+Na6p+n8+GeB/as9tcU
QwXH6EAU+lG3UCgSn3eDpC6rEJOs4GmKi6Y5MHoZtAU+Bp0xmwfhIXItBcLiSYSbWpsNOZLQXyF4
cepWibj18VhzTyaCGIVHJJWv2SCwkPU8ydnglzNheGVHX8utBytTVYE1LJCK9WMWYzFvRv972NBF
BpGx31hIl8cAf9RPyBac8/7jZGNRdrM0zqMONN8Auyh16EbepSFsNTHiOFZLDAtYsfBQi1QaJsdQ
uSJ/XUrZcDM0zInlQqvhJg3RLLJ9qdEVGu0YcsyjUB3Ubyr+Q0ML8B/sLfLqhjeodjGVCYcqzPuz
sB4GCAlIP84A2+yL/uqiP4On8ozX55vXfaZXaL3Y6EzdhHfnDcAwcvkgJdxwnsIoMM2ByCS0ApIm
j3GdPXCsTmmAXJuOr3/1tLx9uhCn+0CoKBrj6i1lSR/0JEAtF+flcMMlnLcPwsNKaEwtHd1t9ZIK
bvmpRZtMSZlDBYYPpy8SQezFGpGG2ubHuB+XN6E7YgcZRQc66DRs96XxJrdZigHj4qcT7mCFbYsp
DCeamNj91qZ6YCtQ91ohz0iM9lsLJMelTLefvXcyumZmXJphf0jWatxkx57mkHzT/+hLdKt5EXER
VyDOhD9QLWCEI32YCUUxdu+SKqfa4Wd+iGr9UBxHyk8modkjqoYfZANs7ED7fnFTTVasC7+2ZUk4
JKcT1B2JF6xCc4100wliLSChMv9weC2vyCrP5oPkUaAfbPjkSz72MYMfyPkPIhH2m8jWbgQJ8xzj
871QO1v/1TRNQBjCgM0JM7LhdVoBx59RJSZAFny/xuL8Ms/ED9u/t9GFCfw5KXCwKtkM3Fqw2o2g
5ZozDpdg1+0/frOMfIoVFp+unrVHdsr+uI5IE9panrzVDIrt7nnhKRT0PDEFqCzUtZXK9ded1r16
LFZQe+Y5YuEz9LovLthZMItN6CX9mMNyQZbKRKYyNTaaCJrU3E0lKOhW9F1BKrt3ws9RJDIUPEvD
q2Eqny18C+YxGSjbr7R3sXybvOc+7QwBItMSqyeH2z4MbhWNFRNbwTVskQ6+NxfT2cVSwQdHwwtJ
obKIBwiB8hCC93GkOzl1tn13oYoO75ieXhkEI4QAnqlQ5xafNNG7kEb8ZeqavDvooUsTbxw3Aa6Y
eOsYTWBBg5WtouQQ46/CHNgS9DXc4gbn8VVt/i2UadPr9oILnqL0JnUdg2Heby+iltiyXf/DaHI4
1S6bYf6tS76GxPU0CZcjAy+kyz8xgv1hJB+xdz22d7E4zOYZJEaaGqTHeEg8uaC7RR49fFsopM6Q
02E1us0gnjR/s5Zxvb3fWtU8WmCd4WSlj8FnwMT+pu8hsMS9eO242wfo+Xkam6MWH73Ag9YSiBNA
VnNLiTh6Q/AHgJ5KLbAh0j2dfbsIcIv9VukxjgRuexeiIunKciVRiQHl4FVqk71J6zraO2VrYUo+
dnNcQO9iWWoVbIMIVLhSkvfICw8cdzLuKwpobfa7UmUi/ovFP3mLMAe7+iWbty/Js1lfsE6ylxol
qrGh3XyUDO0hYaYWxiDQ9S7CCbtHkFyq/CW2lZG2/x/bizD51m5HQL/KmqkJRZOLp6JcV673m3h4
5PfAw0Znrbr6AD+upwohoedoiVn3pUYITrcn5TbrRv+NZ2VyVYgEgJeLlPBvK+ptQSlFDlyuIdzf
Rg3ZgJBh84A1MXejgEfUrRKHZdnX5/4ft0p2lL8fJar5cxyfdKTp/5UMEnXZAVIX9kSzqjFyLfHb
mpHXWLSWCvVsM5Q2iWmut8ztHuQkyRe1i9Pivf4jyY4nvzdSh0SS0mywUA2/RUbR6jzbcCWfZ/og
HUNhi6zxVhce/xlQQisFBDqp574nuFFjEo9KZjTfDNov8VQpKgo5Kjz0jGiy+bGRAq3qxHNLNQqT
TQCX0pQ7JJmI8agx/OKkAISUGzvoFp/9y1lrkPMe6lpbaaSj54BSkvVD7JKb6ep0dVrtpYr2CqXd
dREQLDvqPy07Z/bULm7Hxe2eO99vs+U6c+E6H/uk/tgpt1cRgGMRA9Zp7u0Qal/U/pZpdLiOas/x
sMrT2EjfvbDiuIOepl9ZSMf/VkgU0tZ6GUcdVzF4pf5NUYm7ZLv65QauFMWxEJ32QoRvHcqzh42W
APQ43hqkDoyYgPXYUeScgtwPawewY0eOEDZnPBYT1YaCtnD5HlrmcAsS0mWAiaPaQrazq9Jm2L1+
CVUDg4zcAArg1aDWLzM0EPztArkYFdhYwR+QgFlQ1heDhHsB62a4xhhd2VuaL1ru7iLys7aWOJgS
qepJHAIS49gzSZIzsSZknasx8Th7OxfF+cISMawWgz8GtWw1A/3Jvhquq3dwSmkgv+kl3mKhQrct
8/vsYFi8do6/ssJ3FvP0sX9GRLmfxl0Gjkvw1T6ssoiSdqdms2DW+aLCl5uprHOFTwD/8EnTwAgV
Wsa/uDWLwpf8BCE7LAQaa3AkF/LinR6wEvoUYkj+uIjtNdKoGc23vCsLTI6t1wl5WaR18TA97ABf
Fnb1GtQQwqz0dfTQLDWkMNeObJyvfP/rWcfYEsB2Ss4P0csWxDvlM2aVgha394bIm4fso+ssGzWc
s2KGUnhM1/LPVR0LURuvmH1AhamKc28FBqR/xV++3y/xj0l7A+ibfpleftYXVhJtna8kUQwbeslh
y2QOyWYoa+LTie8s3qzp6NDiYISSD76VfxcPn5E1mtiy5U9jgd/2Hz5EFy++F86WPWMmBM+PFVfM
FInJBvFhDIOdvH1QeUYUXaG1zyFXK1zaf58rR8zFlGffDsP5caZ22Lpv2jCnLIPu/P5EVai5Edra
VlSFVfF37Y4Sm5OGzM6wgYtmFAZHjkjBHyOUjipsmN1CjtiFB7WUAWOa99NU0pobo1CuKsGy6N9j
JH6M9TxSy3KdqUaDJa1Ztj67HOEYJQ7Xjgw3yl/wmuzfdC9C1ST1G9//ofSJEbhBb2z5pSYYoxqK
aozE2iHThFWizyZk59nl27wMDLtOGVxk9fBllM30GqbNvUE9n05Af6FISg+oTqt22hj501DsrnJk
vfTWEzH24RdZYhwbOnzhqa0dRII1Dp8348xiHR8l7/w3ZKwaIGYv6pWHfPru/BTrLO25eLECyE+4
nSeWA9oE5VfnrS1gVaubeBZ2UraDj+9khkDTvCKezv4DiPqhQIB3cksOfLSBR7PpJgf1hQazpCxV
0iC017IoBZP7n9TD/HvUkJrfexnN+Y67ndsryqRGc8qO2G9WltonTeFG19YxxuYuqWlwSIDj3Uvj
craLzQFR/8tWei6huzcRhFPixOjn59FtXPMioaK4DEJQtd3htFBUOKGb00PiM1nVueN821YjZoS3
IO8s/ZPexKHqam4WSB6X70lLhWFPb/l/EZoKt+LOLNvtmDZL3DbZ0bwQ6dCaICv0sLgdsChoOOsT
1oQuOfwTtFtS6KD1Zdri4y04dP+7nKNvoSas+7E5i+3prMss/hsHldjaw9GT8gXcAo8N2CyfGtvq
IqticRwa0JvdUvonkls1uyBWYER2NXSzrfYGxcXtBVsZP3G/G1aZ6gl6yeUZSrVllF7jIGBpEDP1
8mAWxlhYZvK0XV5rcPc8UIju50rLaZRbGM6eFMt1ZUtXjcmPNMWLRg8VZz7rEaNiP6Oeg/q4UmJo
k3UBqYD6otJ4mZdVAqGqB1pK5M5ZgBmY4n+biyj1++g4QauRt4FlREqa7+nc1pQIaXBMTwo1W0hK
cEsKF4fI/p/F6NKpbFmbTXAPsQ/LwfTyHStLfwQk6UaL/xNGeO3QHBa/zblA3PNhzb8xY+uj09lH
vo1PGiCyr9sdF0iX4dovagasWCnNadfIVtqk0hgYknkz5Az6zEPK/YqJVyljtm8dhF1DRjXNd2ty
HdSNpzJR70eHAQVlII4Dd58+bFDKNLUmKaAgdL5XAikUJZr5u0WnfvQ9fqenoiL2lVwT0N1tHVOX
M9jMfD7l/MIYaO0qVZw4aKRiQu1MXQwVY//Er6sMSq96wPWvwViFZrkTl/7RASJUgi26vt85L5dA
wlaFqrE/LdHxffRcRQEtsO9sN9h4XqAn7vZl7nvK+3F7fcHj2hRv1jShjk968r5ZgOenT6Eceexs
tnFHczWTuMooUwlRCWCH1HVzZIg67JoWzTPO+9J9Ujq7/4pgMINyIzQVEtNTCq3isFq4n5h5bgy/
lFhxt/bewDgTyhZmtB+SNeYgd2l7l8yuDdcIb86ocnH6Ah8cMMrjI+Z5VQdEz5cjV1Xjy2x9ayHO
tkNhpxPhTfrMrGYXd9lrDtZhnjjOfBMRIoA3N9TICVGfIAjsxZrlZQ8cmCNA1mLOC1UFZPDeX8O0
1OmusIbspZnZZoPvndZpeIVxCaBNHC70uVdK8uIYXTgf9jDoDfk0t27jsDcFaKLY44wRy/9z8Fwi
VFyl6yh5WTK2yEYrzSfblqJ4UGHc2xHy4QSkIbu5MJzBUvjF8BIiEv6e1objt43Iet4xOY5g8mim
vJLQR8e3pHe7mvKg0vgVljPfHNhMU89TY2+8R0xlZVbI6DM/T0MmbNoEsWnHsa1qJc+Y2sUc0uFQ
0xIJ6pJBPLADZc1XE+/x66fFhpQAmf3Uc27dB1OxoBXiZXMcPVQ5HgsSYaiXiJk8vMG0mmXcuTpJ
Uy7/0libE6IPoGgpHUprwhb6mNb1DwN0KYpEMj+aEcFYLrkB8+CctLuPUw9oeQJfGsUOw+Z4tPkS
9O2TkTgQeIFSO/FFecNhLMW+TM8S5fAEIHevUo26veKR4yyU6aLKPc9x92rg6RuAjgHcLnNJApTo
SGk38dQCI1uDjshqwiaGfWYeZZtArGo+j8iqOsk2tjIDwHGkzUOFYK1TjKJ/S5+76PKLEPm4DlcZ
blWgxcCT66MbB1a1aZbaCTAPzjuGThQBXeQ+b5sLQ9Wnv8GMbrKqvTwQ3GXu6By9PmFPRcAu3+c1
gpBqwWBN8fBvab+70DruyUi7kjUUG5d4KW3f8ZAp3ERNeVkUu20YA8KaNMIufT9mVaKt9W6NS+Cd
9LyU19m3qCxfvqhB09WdT5rj7wlNb8vEnyHdhk7OIrwt/kOINoqUMdcFa5xJXed7cgduDH2QudLQ
QQX0k0rlKjfZBQloBGYiVYpOu2DMm1a952bVFg7I21RyCMlCCR42PQsqlsQgt9nEEkY1aw147i2V
fv4KOmXqiN9BmZ3BR+Yvg+6SC4lz/2Jw9ZaK/qvJUgxKnezXINo0l/ckqi2D5V9Y4Hhh0F3K2oGz
ZO+GbMqV2MzCfAEd/PFH87PN7JII9KJSX5turY8116vYPFIwUhAHSOik+kh06mUJGBWEqoB+TEWM
k2wB5pwk8JlFiMTlyYxXkjlJ67MfWX5tbGhN29jJoOMZg9eLJlb9zr9isiIDRzGWUAYopZTm5N47
tzfmiACxFZ9njGkIPimby7DIZ5KCdkScvUbN48YwPRgHRN2+JBDF1LGiNY/8t00tjG3UZSwhPEJT
5xvQYq0mhzZCi2Cs1wQI9Ng5gmyI5gApXl/0r+OEooMTFlBlU/Y04iI04UgvNTVDtmasL5xNg12R
9h2BZ6Vssd7XP3cEXPgsKnsXcvqXVMXAAbemGla4vP4SZP0qaS53jV1AzgwBSgj+t/P41jMmpAwn
Eivw3IhGCPUSPgnj8xyLsHOiZD6e+GCSOKv6bXaaAbvErmCdSXqpolFaRkWd6zMU8ihyWwCXnF8t
Wmcpdlzo6fE9PFFAbgBjYsmKd4lW6kPrxFmvwcX0f088Apq0ErBsdRXUcp3bPereboIURCfB3Yo7
+7ht7wzT1FFeLORtujuf0kQsW6PTQez/MjTNfzll/LaA1Zwd4X86NBX08kg2pwl0l69SAqwbqkfS
gSx827GovafBjPdZHTZY0SD7l533Dk+nENxKfrRPTJkYFAUKuRhEv6dUQiWYW0aSkaOdZ7hiZNNr
67cOvqn0wt9lFLzofmrIxSt709FAXNbdtLGjx5nH1HSl8vKA+XZMgsK5Vv43XdY35E3Mnb+dB31K
7eGBCoqCm0O5xTYLzh92QAPk3Jpz+jmQQ9gfI6lmWAuGkroV+aPTVhxVn9tmebzeTBR3BRUpcIOu
3MNsL8MV0vdrf71zXih99iX2tHhvejcBPuF3WYpZQj7RL/X9ei8AX+k4Jgj0dFPHpdsL59BQL/M2
e3Nf/saU3cJ3k8VYVzfSpJep2C5rWpissodWMOGN9GivqCWKJ/U2WgisuAM/0i460CoC+UbH0UYs
DgbTeTop27mvKws454LJYKO1bAcKyVYNpPQAtKmmz0Q0qFfGJW5BWRoMqWz+s+RmzwJLhIAvw9FA
zifIw3LlbDIpdvqbcGwWtr3EPZD90qTldFZxxT7Qszi5IY3ANyXUp4jiInCOWsqlLg+UaNI++Zei
eevm2u3ywpyJcyWTlgEIh/ne3DrbuS/NGpUXjLI/8FxGdZrU7s4KopBGhwh26l1ZzLsWUG0sCeeq
MlOeaPKhy6LOEQLmvBrv7qqxKYPAYOxYMqjzJ70cmQqv0DZfQj4GoBtRvtMWm2lt8iM57rHei9j5
0D4rbmUYr1CO5LfZx4z3Fawli3BjlLxULJZUBLOm7eITSW7NfZbOWNRCFPbE3sK1MeSUqyHsgdjb
fRCCSFjjNT367OOTWIVC81/oj1+rSJpCxNpXukfrxBWxGQuev+AFFtXkMiAj+IM+VfesAsh50Dlb
bxNYPh6c1Um1taDgRlnWIlUn2di75K+nkWz1BElhiXnXcXWqZRkW6NsICohd8BkavWmSj45BX4mg
T60/XphvI6RXOjVUEgGdq2gWRElYY3uFCw/cNu+YmizgzmeyeEMPf8n/46Vr7TFyh30XAp3Ry52p
49DfVw6PPfpMuQ9R1/9a9jonKSXvqIKe83JfUbrbPbbHC8nHQ38rrhc2j+w+I8vn/5Hoa8Os+fSf
L2vbzvO7vEoWnTZXhkbpsTOPYJqOPbEq3Ucyig2C9Gn907J0VaNzUY4DnMNRw5sDMRRWTlklQc+C
M4agPFcioFmE3K+H22O2khJPAxqj7hfG7deAj1ZUJadkism5lRvdjYsK+l4slw6ULGdqGk5+jON2
mY+lXULlMgE0ELiz1SJMvh4Rvxhm1Xcty0/oTavV8qYSBbf37q4rLCuSs1EQYWu4OFWk60m/Qm+k
zWLiRt4Wa0fLPmixV5XymcOz18u4Sq4ITAfHOUGeYDJ5YNqgvedWVZGLflO9/auZcJpNtWr1O0oC
muNGMytrg+wkv57VK8Kahgg4BKNzoL051uI9A0lzBmqzqStsb3PnYZOu5+bE3NVmm3+mrFjZYTVu
0JKydiVZNVtTE9lx3hzXJwubR4+lQUeeq4vUVV8a537pA5v0LcMj3gehkM+kgr1nDZtNhZjt7Q4u
vG3r4CewCinHUY9rGvXQKSuBb+KqI+4Zm05H1yjkINVovTjkxeAfB90A8vTksPM7fvUCsloJa4Vb
r9Jp7rvjpVj4p0KZcqhZbgpgahkql3eQ3YkpuEhipCQftY3GvOGfKtbK0Q3wQT+xMXetDLLWlXWX
ic9v/C9EYlWfpugZejQDJZ4/oJBs9pnPZpfglLBVG4yCbUvW5/z/tWyvDrECOFhcoyYaP1HwhBXN
OpNeRayYPYAPlmZskBzDDbj0RE5SLj67aMeBjO7Rl6KJYzFJx7FIjCN7AjrOZ1etkm8oMT3uioCd
pfl9Tq72bRkYaaBQI67lUGJ1BncvBGUJLvvbgde+HWXI7XqMwWAJSISXVdN7oPLwrvqL6tRfGyqj
+dwhhIG94mNytkI2WREPaCJhpA1bGUHNpGk9H6bxAVoXGAo7JL5xsT3v/0k1QlUvnp2p0L2u5PoY
CaBHHZwWaJb9q+y+v8upXXXt49SnCUtBSttdy0RYnOXK+Zxg4vMhN7q+PNNZ2S3/9B9ZgaYHPJmj
aONpSkLXXEUx/tN6ZvJfycx52Sc8/ftrpnKffdXpb/od2FLbKh88eqdoOauL2cEQWcWaddEQr8xQ
S0Dfm054llmd3aCeWFkBwuO3H+bAD5h2GSSPAV5v5rB578PUM7TE557pD4M0x5Dp/OGwncnKBWu1
rQwp+b3Y/2wAFWWfR2CPhgohEFU7iRCUknch56Is08YfR1PtauAqQQqxj4TG9Byu2If9w2Uf547p
cLXpsxSaJdvwAiYydQ9T6xYzHGQYnynm8Dg1QIJAvBIAx3mO/bbc94BX4lxb9ZoEBx5QUrndf/0i
pgdGp9mwdlZdlzB5EVQJqSCuYjxIP07MfU12VjzSBXx4Nr3qkLEYqv3Ndbs/ENLDw8rQNNjD6Uwk
+/8RJDiWZ3OvQSBcjuKS20il0vDw/smtKXDli0RL2KPDhHAM/DXmQwlYFbIpZjucINQZ17Yhe0EF
bu5Vs8jMzVbt/c7vUFX+w4fql7gD6plKkTLCzn1yccy9zleRhrsuRnrHDs1gmbiLXm5PEZh72wKO
uzssfFQKMP7+qt2SMhumKwvZTnnbd+sIgVR70SGMQkZ8/X2zoIdZTKF47Rj3+AQjJBrFZINIl+ca
judcCK04/hQ/Od35nC5yDWynFsgZUL1pIC+gs8zqGkpUQg3EePugSS+FxGgzh2rZlRHLD5Ynf2y5
x9MtwK2z9T0Gu7M/tIfcnyL5HCJ3EtNW6ikppPPrq6OzHFypooPKCW5McIownqm6kEIyaMW/tTjt
rkAa73lsfZTu+7EFJ599ojti3ljFg580BbKgoKItnauFrT/qx7YYHsORWJXFMz7uUTqTQc0umC6F
UYtqseenX9iEIPETuhx7MElrMrScu9fXkAWZx6aC+tngRayr1Vq4yDF/RaX7NXPBsyjf7RfPJ9X3
mTt9U77mYu1h4bZIUGV78Jp5x/Sklgmh/RPeY+Plht0X6MDOCNtEaGNx7lVw2Evxd849nbsNMr0Z
lyD+S7vA975CfTJ/gqcmHaLHPAkmiZB+WMY2m0F123md6cvJm+9xkVH/8rXztLLBifd0CvbKVYdP
GQEuJu5YhelWzjNVcYCYgZHG0IHv1Csjk1hv3QwH+wN/PY+VmY+TEFLFStBVE0q4FibHKC8SUk6s
ubwSDTFXlkM8reo/h3BvQep6qenhPBQajh6DhDemqTa7JT2742R2c37ijQ6pjFf0qz1npkCNaOZH
u0Khylg/eYXEvkbRj+0Htt83joWtLXcb0Fe2oA3H5RU0f+Xk0gLFIDBxFb1KxWWfhtpETAt10cd6
pGBQa4q27VGp0DzE4t64pMO8GdYxhLqhX6lWa0afeBGwWS5weTUhTWS8fg2M6pvk3kLPRiDtyzRh
qrKemcAj180LOF0qZQnzqzGPmUxlwL1RTco4cleOBGD62sqGcGkLYge2qs1KUAfm0HwyLUBmlHty
M02crDkRa8EU1+9YZUZ2KGIVwpuW/iLmWUil9yPM41mDOSQLKOhnRUdskkWdwjQEEd3PiCL3wZM3
q3t/F+8LHd4DhL6rg+XkXePx33YFrAohI+Tbcwdmh89yJa+h9ND3oIlWkt7vt4Z6yDnlvDdi6ZEA
Jcvr9SZHKzJNQgs4NeGRLlEt/KYV27L4yAVz3RqgmEhSICWmrqKwSQOqL2F1QuS+jg5uMaK9p9A+
5w8mHrvT6em2LxRPSD2nyzjfZ0FWt+HyuBXNOQeXibwaBVc2V64xjR6rknvhSzFJ56jO3ZtdnKYA
it1tEWmyEsfFUlTjYWcxxOg+/9Y9LxI7H9Kdk5iBLJvRWBN4TmcSx0t7B2KkCEcqc3BBSDi+tCUT
bPc/R03FFvO5iRkUXkjYtgat7IkvlBaAxT63xNGskzQfMARDM5EFWJdYOfZQUFWnIqAnJzdCW94I
MbqvL8VEYXys5csxv41mwWHzKGRxRkx3yacxMxR/aD40ES5sIQXVK5zdysiCDlVUqJuY9me/2CAy
610Dz4l13Ziz95Bht04xrm8qvW892none+it3o6r3HB4CvR6mfKo+QPLxUeHJ+y70q2jOSld+hjy
hIJtumFqnOMTDtWBxPdMHi28sb9nwkYpQN6n5ap8/fL+Hm7YpuZyT/eHQTPLqJvn8NNb8WZ7a8eP
0BqVIU71Zx6KKGryLYHLNK6qmPq3r76iI4EpdIFO8zAF01saQpGIxJpfxhnLOr7I7t8JWFTzIigE
MmApzEmrqRjKcYXYfp0MC+O3PvMIWSjL7lACwf8+siQBAKBB95YUzfMlSQmbHpGeQlbMmfEiUSvd
PPeZPFFFcEHJqppfdiLEQCusOEU/Y3frTSBeENcV02m0oFnqjRMlVn02uwwVAdHWw3DaoxQHbJK5
Kl1cj50JcMIKl1clIqiuXROGpx0PJZJVI6EcoqqC4WlbokMCUkOq1bZyjFfb3MqWzOwTmjGv/Twc
z75UNzD+0xXV0swqgZBhd+f5LdGS4caP9gC7UAzMmAw9rPOT3GNN1PpEtVLZDY2SHv/Jsoqn2XZe
A8kPMS/czF5GgW05dRryJIe7ugp69MfkiREVS3wE5+Y+gbm/0cWTcBTLGV7N8Ix1s9zdkX1i6McF
EDmm1pYrZvsy5PPaO6Gr0Oloydt6H0dBO/mvkZnj5W3aVg4+zi4kb8Kk/xzKfEVbzfxlPsHBajQ3
OhPJJRrbjG+yK9Qsky9ch4SNOCjaIWXbjoKGc+5Uq4FfKI5x8v2B+klHiYcdZS8F41bMTxttMoYt
IwfVt/Hqc374VtMSZ3rmNO7YX+qJp3JSvN8KKaUUFhKtZnGBQiEpe7UrSrtgp3FZIF+zGWFuZN6c
X3nZxXOLlPoRqGsF0PXld7u4eIhnGafgYFTG+Z6IHoYxEMv5DTrMdsKjFhTPBbcod6wVXOFDuikK
bIxzbJ+w3sJFGA5WRRweFL8H4H+66Al7ksrifxSQXrakspUucCb9a+TmB1SVFC1ozy+LlCThbQ88
FpHlVxG2Fd53d6c7g4pN2QEcwc7Dag6zFfViWO+u+dZ1+vn88Vg8y8a3347lJNlCeGwQNQsAhDoQ
8ejYDCbgkdhiw73LRS+qdDAq29MlGytuTrHGnERmnclP8KIsIoLp/e8oMuY2fJ5yP6IHBajJ2TGL
lu+DVSJqgNt2bnX00N4zhYjPTOqqFfU52PQj4qAx5KSTS0Fi0LTxKMgOztJ8hOVzzESGt+lU8ApP
r1L/1Xj0qAFUZdZXdXgYxAnAhgxMOGwnXb40g5cKlY38n447FUOu1wXhAVECzPhb7aB9O+oi+7I+
EQYIzMJxfHg4Hq3/1hs7kR+OEutttQldLC8McJnYKrI4nVm+fQ9TCcqXFnvejceLr2CLYWqrG/mJ
fTGUxKdimaebMObIL2rQbPyx1ccQ2y+oGEdZvlLTz7MolG8bayY4t/3Q8JdzRWZlGxO1/AOx21U3
cQXI0+GMwXJXDq5RuTB+zyKj9bzIYgJIQ1s6cutZes73rVEvevauHPn712PpVYCInmTf8QSI/81/
NDOsxu9omCVS3GYFbnUWD1C265EqYd1vggQl90EDkx3b4LRTGo7G3IWhWXzRh+sC2ZiTWngsebMn
K02oiC2ubJxacdknbI6HSCdwo1tTTxuFZpztZCgzlmUJWYfaEUOMHul20y4jb9TnQX7TQGJxYeF7
seaNfhUUeTgsGnAo0CnUh4dvcom6LZQPoGJW5241Ehwepe686PnNpWaCVZ6DPurH0mwZcQZZBOuv
nKHwSx9j5Td9zTni8UNLcf+MdN21N7LbYf0YA7qXq4COTZC0BVaN0imlv4L98uw3JGmOB0ux2NOd
NYtX4AfEtv2ktuJznR8PM0RoUEp3jQA8Rk0dI0ycC7s/KONpxkj8vJEaUbFVOh9tWtdonFS8BvjR
DWA1oU7VsILFCRQyq/gCM7+iuN7JqxJWP/mcn3Y99XUGSVZldHFztFvIF1FfEErWFrMzKS/YNDt4
/TR8WfHR+AcOvFKTZ6csr/gRDShtOG58YZoumL+mDsp2RdbRyn6ptJPQOC88bBTqFugNJ5TjT0So
DjBw5x0pol9oLdLzf0nMKXKFAhxrhRGvA1gHVqa4L1rlAyNYi2+JboNhfBeY7UheKHKGUf9w+4lb
/f0vWZJQnrUVW8t70leLsIBlVendTXfcKK3W9yVZB4WsrQeKZRL96MCDN7GgK+MrZSHIDHUvCl2+
Rr/LuD3b5Z/4GX/eBCudCfBkfX9BxeSNdeQJkhZW+0xbo4X9PbIoqmVM5lKU9IYjMtrMvaQtmOQ5
tW67vxzGb6lGbxnhNt099kJVHU6oIKnGtORfefHF14IVYEekn4dQ9WyVhx/GIlKczSnrKeA4ToSF
7Ty9pbCE3aDGDVCltMAfZS4OWzWL6BthEB1kVLUGcE8q9cA1JkejGiIbAFnF9QVb/kN0sWzybE+V
IWT55Ciy0AylF8CwQMn4s9m3nTTHzvPde/KqfP82FhkcvJAAAHCswnYjeh/MvoJHtB76ipAtysAB
rXHDXX/MVlFmIX/meqYPmePn9QKlwd12mln9hK941+QWwZfMp0UGBxFY1xyM7rnipV7h+wiTq7WN
0VNyqOhaSQr1+IaoAmfurmmqOalWgkCwG61zQLGYWoI9NoiKpdH9h6OLHN2HWOklkyf9HKzN4s7e
5jR79exJJaVTERbLHeIjqLUY/Ni6JwfalfKTY955IyJ1Vv2V+3yhUbdoKINHuHgxpW+sROx7Rmc9
KQD4ePuuXyqYAdmSOIhB5duarNEzq1f/TENTZ4yEQeiide1ommySUdgu7SV167CmFatjfoh0eudu
1BEv+8gWcla8YnuLvY0iOUo9ZCtmyqeQB5/8cbiZLAUOmwxfnNUFJyUH7dv2AkUnvBdO4HxsIK61
QzZfeOwfwBkMSAaBywG3x6oyv++rzrXAS2lICoSRK2sX1VRtuLLPOc1j9QAppomwFKdXTG0ymZna
yGirro0Il4MqkcDZ0coeegMMyGjCIhZBV7wb9YVx/B36TfYVaJPxYSHFiE8k5L2qr66B0EUpZOph
U5r68nUlhNMHBdNHlcH1Za8TSBOwTp6nQ6btjwSDejx4DSFcpPGBZnNUyc4q4jTwlB1iZp9DZIcU
hSOMc5s5MDvtbQR/Do1zfmTuP+1OsBwyxg/ko8jysOJFhLDFwaxZr8YCQLFntXwvNTPzpwMoNCL6
T9BMUxz6id1bD/+WKGfpRDZDox4FlLk2+7WEjieMJK6p3v7lF/OA4+O2Ski5KQMnkKi0ORk9g4jG
xAiJTYdIk0bz5jDZN4Fns21akAjDijFUqp8Dh6pA1vF+CHJZ4q+KbQQ6AVYJQ+cAcovooy7VXIXw
wD7hL6i11yIJ7FsgGWIc5luJPiXh09PmJ/9w/IjN6GCqV3h503RTqjawtpp6fmeOkIqjSO0Crhrj
TTw8ZEN40T3HZpKwCBGpEEVm9+cLBfa+kGlhgUx2mCZjN9uVqfwJffho5ib4gcn0nPWG5vYJRv5i
1dm7gQDloOJ4JuLv6hONX5tdQWT1ld4XZdVEiNtPoD5iqOkPYNnvOqFg2idFycKS6AFC21RJVIAD
MI6cly3PB7vz5B1kfmL+l1bfUWBkKt6zfR/zzHKmvPnBFYWtjrAPkuE+2CTpd3x7XTzEPaMYt/Ox
WHRYdGNd6qsg/piYcNVaNIuBZ0D+B/f7Fh/BUrv95Pe85o+t64J6VqnSEScxNkzbrehIAnYjG3Sd
yJTzWPUWxM06jXtOG2f7bITTY5vRThddFl0y6JXl9Gk1cvDmq5ySszv1r/nydGuG364Xsi2vv4Ml
oha1E4mCWPI/Y/h8tKb6I73xdbJ33ajEeyxKZwATrxyKJxT2qdSmQtKEHwUnj/MM369Tp7da+eQH
0hx2UKVDaiOF8gPBzsBFwZvj48MnTtPARQo/LVbFWG+xK/Pk7dqlM7TjCmD2hkT4BnKHSrgH4iNt
KAkK8NCpHy66njZtch/AhOWCe+xIfC0/TS+XHvjhPPQ8LzlKx8tsnmvh4W1df2csA7ySM8uV0mjq
xj++drzcQ6DlpY5s+/0l42XDbUB4yZnfqRvtaXQKz01am3HPQfh044TQ+VN4QByYFfSStdvsEwh4
BkLYl3xkIsgjGZztcVWMcaAnRw7N6zblPHK5fElDNrrfnQg+YP8Irn6npNVnQuNX2/WIU9KgB1XY
SHfpy2KzAlHR1+nqRZ340BhFoluNWDItx+0405JtnotbdLnUyk69ke2ums2qDhjnO+ocXOvVOx1f
liR/Bi7+OeD+eNeivNjMG0JgjD7VI7wYKA9SUi52Y/io+UYFLsshVGY9xgET4W4VS3RxKir947MK
ZlXtvgEiy0ZDIu1QGSYrgKhEjZiQX7fctc7Kev5q1NIUKaNxYFJfqYuYZkkOc5GwSDRxa9JKmWxM
jyOyEK1+lK+FAdc8gX5r41V8orLWYsEmvS0NeV4JWIajou03FKB+mAuv5d7zTJwIt15NHHHtiwW+
zLYj0XBnDBFOa5i9z5WUdOUV0HQghj9pod9B+B61k03H2kAOzwTikS1OoKyfte4wi6E3rEjrCv3T
R4gz8Lwiz1v5I3UoeW0t0n6b9Vm2uaqA0RyGNMDQrBguugilPfDkLMaS8Ii7Xq0h10YxfBpkoB/j
WIFY1YHFc5kPPzIq+hek9APeXKwz0oYS49Bbg5uwrBiXZAD25y2sOhdnaIwtPgeXSgMLJ90RctJY
5E3k96pGLf1xBH1Y0dBfVwqTUpGru1UeXW9TVhNRD55/hoIx56nLmWM5mWsMSAldfhbA8aWFwgdS
hvTLUT751s7JeMjOgcuPsJJgid2fLalKPdVm/FYpzPAWPaRyQgxpI3UiY02CZdbb/IecFd5p2mbR
PdqTYzRca/hpHYEzs52ZDb9aajgZdIfDWUsBzE42pKWm8ZPdEXVIFRmCb+wIninbiHl1naQHstiv
Y3x2qIoiir1y6H+x8bNuk9SfZ8YC39PfAND7PUCkVpsAA+IP9d8ZMuJBMxwzzo67E0wvVIg2cqUE
2HNQE7OUGcLIPgPsYYAU5pvwz+80+w12J8s8r89onNa2o04ymt4ypGXlN9DWsz4Zez/S5FXx1gyZ
SgSX29SFU45JRub8CeBABqixMu1Na59F2iFA1ebd+9Qpkw6Kv1Eo9n0qvU1EuzqvdHLIf0UPIy54
hI3ud3UEACOi2FE4dLrF8CW1AFmbswsYN4z3XfYzEGsVLvv7Iedv4dcQvRBazdIGJYfwMujMN6X8
Zq+NaZ5qohqMBzjOSq0YJEB9aX1qo2wkAIuvi64SjfAll16VPQofGCwZAX6jucozu1Dy2t6Lvw/E
u9E19Hj5toWcFcKtyeFT7chmlNb90HAonY1jrfOk9EpH+Z6KxTdpnbBUhiYFVl0kPKG1jdNNbu7L
8NmjX4WH29rXwH48vkUJyAco5ZVkPMEAirYzzJJfHATv0/lMD2tYQiTYJpWTYPpL8PAuymGYwNJ1
iIqcbk5XMwtiD8oVlTXYU9RsIhUlEWTcfk14bKASE1MHfuQiBb1LgDitnLSVfYJLn9GNj/vUO8Fz
JpPcT5U7MTB5rjS5/7rxsATmMF5roxD2OzH0tKpOFa2cpLv5au2EC0o3LPp36P+FFKFVl/WUezpc
NrqZ297t41HPs1HyRXXxwIwxCnoG2TfWQbKLUxEDIj7o4CUb3TADeHnBXF4eb+kXMdOgn4NVDI4H
ya6snd2tgxl2D5jIyVCEGoKmPqGmItWE5bbCIT1+U+PR7KUnPsBxJ5/LyVq1mf/vSzy5hvovEG6a
jOUQe/AhyxlcQ6rJ9S6r7UNaZHeZmwg1lG0sBaYP9vF6E1o3sg5Ms5oZqQFsNjTeHb7cMGZCK6Rt
dxMSVcF39KpFEJgVmP4dnZ8Q4YCTQ/Paqo5MrsxDYa6N6KzHpNZ33HYyL2YY6osgmnrrxSWYhh+T
GLJv7jiRy49jNyJHcrRre2u9jfANEDUfaeh5mcojBBol/nzlsvTUL8XvILYLCCB/BE3l+fchU25j
zdv+EbOXj4xSzz4g4r78HD2wtoO8zXW8rJARZebRuYCH1+ZjBqGT29GezGF/gAlEqyTcgQTNWRJX
RttL/oV1XPJF6IlVm09cXKAvztNoZmxaMMLG9bP2+moRqB3US2Y3Zm8tPadtz8sbaVqKKRN6FU65
Ny9vIYZEYzD6/6oovS/+cCMI4JIH7bjaxgxg1Utq8X/iy05IVUaD2GfsZsRyg1af9IfJICRzi891
tIteXWYMsAwsoquJVpzfzDTcDR4oXRsH+3JZHanVu/9RlvtBvtMBgrwpLmCiXnL3K/5s5Yny7id2
v7wsYOgG4rgIeaVIzWVekBb/E61gwUL0nU8v4oWIOtOeAohDnMRf4ximP3kmwkjVCwe7AP61zmsJ
ums/hkUzZMTmVghhCRiv9tT4oo6b9oRKSR0H3zZFzRGWOdIqvOhxtxnTpzSNWuGrHUBoASL74fWM
c6UkSDfijCLEgiZEAo+KIPHLg/Y9U117l7mNOvK3z4VmS6s7iRZyojx6JJDOgNhV40dqcjxFr/QZ
QnoKE9mwrGEmCl6u6fpyEpWxl3nYBXl2tXWX3Oil74ID/BgwSlOTQzaM6a/KjmD4Flt2wq52cXX7
iwwThViQ7Lj5z2xtDqATX+HXsSzgvDZLCunoKlHS/enrO2ayxhnp/K1gvw8Ln+0n+exi5FokoQ8V
jz99xNdv0V5/xmTTRsa2fEU8pEABneMIyEMYesl9UPYd7bwOwZU0UMvzFQvXc6htPbPy6B0weJvh
ABycY9Krh9HsS8jnOVCxwKixhCnnTC75ERXnQ5pPwB4mG7sFwdB1KSWCpIAAHmc2E+J5ElAJud4K
037hvWUbVM9pq9S1DNszjdc2rOFEVqsNDy+PB+RNkzb06Z2e8dD5KlNIDRv7UIB/0Omie6t2dvLv
xz5puKnFsnhyI3jQwMiz9o9sbnWCcQxVLs5CDx0S3oabxGJ9Z5pgLzPc3EM2Zb4lbir25XIiyqGG
KYREl9enKRHXWv/uDewfs2K5cIFbbfdvsVSwvn7OxdivnjiZeXp2XiRzIxVagLcSSXpQdDmPlzgA
xB72mp+gBaI98djcuc1kG2AZ2e7cRHOfiiu2owebc6pc3/NUjva6yDjhDCAVeMMkoH+Ptyrgf3CE
Ir4esBo/A+NIta5lYfOCjq+0KCekf8Tg04CqB55k8sqLwCMx2sEVtPVCMkx8sOnw6S2WrcjxLxZ2
QWB0t8ozUWJRdSrnSsp8inq7iLK2Kucf6zUWA1Ul0D1+c5clbsY1IPlHv0PgVlW9LZkysbGPAo9P
sR24dp3iT4JCWdJpTVrVTEjI1VuS4FRBApWRmgiJqCsiGlo6G7fmDkkDImAhaawc9zqVKGKlnIkd
7GWnfA13yxUhuUk0mFxvNb88aDX1s5881fq9F7duY3x292zc0ByGFqAv7Mkx7zxwP3fw/5HE/UQC
kuqd4MDfeYi/gX2uWYlXRSjIOXCYQfjWCB2yBCTN20r6MOtDqUjsPhe73ekJLHKLY55i/0qDvors
RVid45wOwiNzmA7OGnSFsLNA/iu3dl4Hr/7njoHfdl3zcvW3VG8XNJPkVZrVZ0XV4HlGTEutXmcW
avuwHoP42iund1H0ynPwkg4w9Uxm4VYGxUqHPXKq/vXTKnSgcMtM5Jg8QNAu3wvYcNol/rsksYcB
kWs/7NQ7EfNYSl1jOgWIh1ambfHzkXo3yxaAgBZ2jsuSOHbIZp1QgWLSBQB2mfc0qjEahoF27HD4
FGCQH0xH2FIaFv00C/JKx3Fgob7GovRrNb6J8ejDH1L/1wxMUlyMLa2/c+dmm9+59+f9icdPzHrO
fhm7Mseqcn7G1kQ9fMB23PVNehrdmLwOq2JROPSW2IIHQ4X/tgP7PQ+QiOrkhgmjrzSLhHyIoBCN
Gkvt0H96/1XEm1dIu3dfNyfuwVRRkhNZjR3hpn6SzDiTB1dYwNKUve1Sm3KtEphJW/Tjb5jNJJwT
CSABMM2aX+sg/8nlEN9RcqXFoeft3hW2cM6RES4cUYirUKuOZNgCh1T7ZiiUHk041DPQ48ihWPh0
+ckUAHFIKoSqHySl2mpWP5ZKVIPlFIj+m59FeUh9Kwqw3nelNs0o4oS0hTXaXMf1xnqXVoDJT03R
PNmmbkq8pR8IhMySa7attec+efW8P6G/Iy0PJKhY/w8X61W2eKiXkdtq+BynDfqGELtawmQntdye
Wj8k6bJBWq/XVdiXIpP9JY65b5HIYCGQ0FJG1mC87KanTUlTKyf8c5m9c1GqvcPRMwam4iX41L6t
VoNXYGGLPi4SxCPb2iibFt7DW84Pwsc4gf/v4K9jl36mjTHUEUZPfZ2duVij2xQZF54LR44hYvUK
ZOBxq1sutQ/Gql2pjSRHKacoDSzcvEeVBx3T+JaQIFKdsw/ksxCVJUMZPOEJriGO8qxG9OzuesVF
lKwlwD6A+NKAohK6PdeaXmlxEnhJroECZjEiM6hCNJjLNdykrcBHlipEShAKKZkihlx9GBXSgZYc
TBLj6FWj1DXyPnvJuhpDTMUPmmoPX7CTuq65D3U9q5nO6gKf/m+Z+CfsC4EXN8zvxNLwP7MwGB9H
rXcrOboQKwDXarEdCxIklzzquPBwegedrfpX1MqK3W+jgtkVeYh7Ue2vVhwHwEuS8m1W8vEob4mN
N8auLT1wR1yMHoNOhdXZou/eYsFJqzN02RYSVht3r/Gp1yjLUi0+fAwMGXcGDhpKnWdqbbGK/w4K
sq6GX2hpQWI9u+DnI+ieUPpeDdAnAMRWFZMHBpWZxHmegknrK0FwgeKyh7SPdIBxDvTiny8SHJlq
KDZ9Ycetna93N9cIPqLcm4xG+drm/cQJl8oAuquzYuNiq0rg8TTJsPs95LUX+diGDWLYk6zI30U6
TlfYMXIEdxZ/nd0mZomlgrIOOTtnP8m5KuLCAwPDWlFMWI82b4os5xpaerlDCULVN1iGK+YhQoe6
zerwK17Ot9RaA/fDUwAVUp099ZDEvc2JJt2T3c0k0zNnMwWDF886RhAeZmjZ0btJGHpk8m3+5QmZ
cFF298x1yEm5BizWnOLv0cEtkAbfcc9rCt2iF9B/wt3+oEtCM+dy3GFAFlgu8aynikVkc+CNjAzM
O9e7/xvnB11GFtPppVhGoSJ9vEW70Z5gPCFi3M9gLF/TQaojszkj76lX3/u5x8ez75yJUWae4wSZ
I5EG+V17mLMjWXv6HAQs170zQzIgONCmR3K7pusiWhFguwecNKsq4xgrdUBXg3OtSsRDz7BbqLkn
4CzLGAqKvcICgMQQ9TJe5O4+EozsH16hisTStGzryfxFjes+0s9FmGgnjDEAW+8iJR4OfaGqwIIv
WExNxcFtCr2cUSFMeGqCPi9y3i80/Ny6XYPoZ0qDebHXor0V/T34Y07N9rgiqn4uDWAaUYQWrEpV
JjSkBGrxCgxYxPlWwQyEqNsO7tqpzQhstk1+EOVNETbV4YIuF8A4E738VmC926dAx+rpuV3/AtbQ
lrXUDXQpy2RAWY9XIywrwzFynD7GsjseT5y5jXCt2uIgWKTVADDNtD8MNY0xpVB+3V63/+GS7wH9
lIVnz3dc5R8vJpcH8PiPxnfDKD03flnkXIlSWZzoPiO1Ny228S9+78B5yCxoVJsUmw7WG4e99mjr
SRIRwTeX0S4JumkK02fZsZXXD0isjPis9lJtTZRYEpjYLuYG8pr7om7pYsFD7nPPlM00Wb/RySkT
ZFpQUjGqkUFxTAZq20dtqK4kM0bl7BAZVt/NG0h+IqiXqszkyQ10jD4xLYuR2gba41gzRu/jtFn5
7vqc6GnCiRcVpJUq5AFd+G4KkRe2n1xTHcBatOuRq6smPyYds2++VglleHuW5RyV1Gih/3OFhg+9
1MTRl1SNHRi9rq+dVuQU0c1PEEJS4rXwEUYpdo61WRCnLGY8cWRzFj4a2piEJWzWa+aZSkMyBj/s
IVct0phbSpaa6hUGBS3+N3gaGHoIrhS4WW0EfQk2NfibO5g+QIXeZq6Fc5FiYUO5mlM1MRcezWY3
PgnYN87SWhJKL8Eop4ArAw9afi/SmUnuPNDmdPJligV6pWsD/AOrMxGKvL2jWF0i8KAaSofwAYO0
JO2ugHtI2rNy6EmEvbdGKIwPf6sNaMOOnBZVatbkj3JsYnysHFhRisE26SI3RuEAah0CEocq23OQ
qogANcYOzht/KUCVVViZqSjb3q4/ZdsTEt7hf5u2V9jSCJhy2wYIFd8xjso55U+e0TzXNRQYadvA
TO/IclgSsaTJS6pQTT6IHdD9nWA0XjfNvkRVteDYCo2zv5CIcCcsqxReKaRh2x8LZcV3UGzn04sx
pc147F2R5lyddc1fVxM2D70MwSRtWzb+f5HsV/pemiMQs0TXpbs6lZedwyI9544LJ1+RjckIrBMz
DHnmKqRccaMyHKL6yRlmmwnQtrxAqja2cWweZtRfXqRo2lWdnjTl9lmi6mL8FRjZb3+boJY70Ib+
Fu0Y66w7LVFiLIpZenu1pFKGA/chDwYeeZRSL3aBJIqtG25TTaScr2VhjD84f+BXDPRlejGtc+sq
XlHicDZqG1Q/2/+y0JiC8U98hQYUMQxEFWml5MPExacJUdEQqOEqEKDE/LQsj1+SuxZgwTshr+X3
u4xXEabBIpQnHwajKKQCbTa/2r0SwL0n4YLFjKmxz8ikkYjHiZfCfjyCEeFfOvHme3FYOpP3yTlj
c9aO2R3LoFAhQo6t0XbTcTfVfjFoWxq78gagefeEl4C0GrORIWKxtOkCwDGQJuJnqjqCbDZfa6hO
rLERA5m9BM7gUb0yc56wRkYqdn9ctwvD9f0oh9GzPKJE217vsiUtkhnSOXP37t3dw1Hu2w4feogv
eoK5fLTk/tOo2sb2AiDRiEgI2VU0lqyRisAAUcYYUPWfX8RPhbDwxZGnrIRsSgSabTiJq9zKizlC
5P5inwKru2QCp9rBvUH5e1on10C5PU09kWX6e+xSMe47N2JdhRSXK+blxuCiUh3mc5Y1mUyAN1Wp
d1KwLRsPG86rjewp94vMqEWGlq1BRCVwrsY3h/fCyM5KTuOQ8QHvTBu9hXJchwSaS+PGi/fQvXtS
bMctCxarIaP999MCiDqB3HRHtod4S2dmxsG66ClWG9AtihfRFERtnwCoeWojf7PGyCAtUFqDtJDn
0iN1ZLm5t3LcDR+6XmMMMbDEKsoViyYtMtHc0yBOuRJ1ryttIgcWpf340VpSvmPM7C4jz2hfnrSg
gpeqB0zhGUtpQM9zM5B1cuUvScoOFO6EKqc5wXk+AIOrPpwOk0nVY2Ay6OBIQqLjSJEgevqQILtj
Cvl3MPYXZ88lvrRWwWuzfCFT16fNzr8tzFeWyOqyBsISoJmfBt9jkCr2iY1o7Gx3+Kzrp/ulVDsU
t5g//59kts48CVmISUaZDWbk0NzdGcChMMm8DJSWceqzZYeYMguPf8S/bl03AvwqcmjZTymDC5gL
zIyW5umFUHpiClVhbz67Si2JslKNlcfWfvNT47BXAnb1YydwCYcaQg3oJ7daBNPfonogC9rdtDX5
BIJC0b2Vb5IzDeEX/b5gMvIlRRZ/M36S4vBVxApI+Cz+hq7LhDasBOi5+V6mPvS3d27x4CYQwU0m
4mDzKn0vBFFKJdw8OJu2iWyhZFvWLnnM3BQlOLCzn0U5aZQKnWlnmfo5vd8DWwI8J9kFLqYsCC0A
nED6GqZkz/8mp29qCPUO4OJ1k/vrZe2HdXk2S6tNiKICnsD+tGmXlN/MEFaDmcA0VzHYBkiPAdHu
tUNWEU84WIIxZ2bBXjlS1/OnPspHyk741fWjNa23k9pRt5Btqa5segVJVqGn8w76s9Mk7u+CUNOW
ThL8AffNyYpCj5tyUtE6zjdsQYlgMk7AwRk6FJbrdlCx1FV2n9AL0/XfnZmKujhTNa15m2sqgbIj
zjJ/Lqo394i9G2nWFqYWhIHsHm9aEvIZ60PpQMm1Odb54VGbneyOCzeshjWCjPHbHSuJsdV2/pTY
QgUHaipnFypgj0+mPC6vaPzjO5lI0DUisYYvlb6HE3M6q3RkEO1Jw8Gpk/z2PD/bhIrK1Qllo+sk
YmVOBm/VHHYzdZEBS8zEHyAJGO77d+uG2f8/3cOEagq4vaxbundpnTr643Ug90elzz2KivkkYaR0
lilPPhcES85x+74VD9M/ncjzOroEqWiB3Vpwa0Z6ybTTzZLXRkLKtxWDFp+mRurzTvqHrB4U/dAu
17fsxSx6BQ7q/Ql8+oKngyhXOfd7AWt3Y+aLL+yUkRo7G/FlB3ERmgHVa70YS7or5dhvXNK4viTT
f9qyo+tGYTn3D/uScP32PfTlO9U27i1vVoUCiiE/hegsZ8Wjjqk8FLPpEeVR7CcLPFpXXMkBGdAv
aCZTJ+dyB1gWTTAQ4t5ZIJUuwkyRmIfgQKYP0ehbZe4RGAXhnTmBuTayEwqGPBG9GtU7+3Lsd4E0
9upcdvykTTthmreMVGPYGPouCJ3airKA2ZlK1DzDSMaeuDQ3Z8jY8g1knq1Si3p0/FIopOrDNE8x
93aYxaOYPRZDowE7cm2x6/m4g6y/hcqy0+pqh3rQ33nOYUBSIWN/MKtTC2Ets1ssrNE3eYd9+YwT
OboXtRgXD+WdnTgkWxrMQFn/pTpF6sHVYSwn1QMqHJhSxaQnHMOy6rcCsByAibF3/uWUoH41wrZ+
/qoow99wF0RrKZI9e8T6y3swQCEIL+DxrYMsOBpGuFsL6XFUfHoq6rOMEECmn/Bhuvs5KYT3WuMR
h+NlO5i2pkr4BF7UTHUFcO20oscZ2x4reFoIojIuH6pkJgu/fzCJXRixUKAODZV6vz6FGR8KGgqK
ePD1LSH7RVOwGDqe78lwqLAwScG8XbPXoDe/ZC9cf/Cr0kELKWpoC7XXUUk6YQUF2Cy+V1y21zlD
2o4arZu9OHuNs4RwrNm5I+P+BHAtnt7lRIMj0jDTv6LIgRW+Je2XTubCznb1aJl2dOO96hNZIQjL
quYjgMCJIOLNyysKUQHDM0hKkLDxGpO8wz2ygS53PwIWXk6eF/WvUUmadBTF0t8h2bHOoTO0EMeU
SzaTUIAxGgiaBUJQaoCS7n6P+O5OevBJaAAFYQu9xfMhM+lpiSLDyZAeELXFA9NOlaQch3nea/+N
1IHToZrzpWGk/OyRW+cTVd0ZhFcZvt7KRA46NPzulBTSCzbtExmt0QDcRj9vSO9qZymharqCkcsV
kL5g8DboXxrVuGjJEPjO9HeDCb0J+MJzNKvIsESi5FQzUipH4o0+OpbVI1LdTItgYsSAy2A8yrxp
R/w4MtCrpki9y0tiwy+9bcK7Fr5qb2/6amaPbe5cqB6MNgzhf6M8KLU/HYc7uZfDXv2hADRzlOUn
bIYtSUGVZwLLQpBpoDqhcJcgUWfGSjJfFcT6Rvl7hzwaTKhLWTVUA/oZMw6m0Kv2UEJMZzzYw/HT
hpoK2rZwT9gBNzBvHM3i6ZSn63/5gpvkFEZ5cyFRKC8k/ez82zNknuA1tP35eWmE8YGt5MU3WgTm
E5jnuQcAioVy+bAoFLXn4ZRc3rmmfuzdGnK0bY3LPvU36PfKxSmdb8nqoGd/f6ZDIv3mkoZ9quMd
fDnsucNb5ymq9/jiwtqPO+/wrjp1sy1+adq+HmzESYnNyBw4drNv+t0CnJISYw6eeOxMimYeYuAq
u62JvhaLYk83yvhVMVGwMmAedzn/GuxKqSqoxLiGNKCwloBWqrh6PSV3HpQyop9tqOoNuNuZ92Dh
wfN4mMJKuDw2op460FHl4ODaaXFVqep5GKB84k4fe2EZan/BQ+G9NMSi2ZBQDnfK0GuQJgP5xF5e
Qa0kwpV+o/f+Kdsqq8477bkPHhBtAcPVaxo2nNaI2G9oxvW+UIAKN0uzCnc0c35FiF5OFC6ivFz5
2EGeEMZ4hagvdmp7hQulVPHakR8Mna5EaKRMk+ax6B54Dq2dvDfPYpJvIJaPGRZotYGBrxd/baeb
3YMw3Gf1hNYFSLQidq+8H1qGXIXxiIdhx+v97SEy4PVYV/AQOYk/6Y1niEKlPs+6SNon4warLhSE
Zbdq/3NkLnEi12sd/LCGJAD1sXLW6YZCgB7w4v9vD4KyzEaSn2w8KTcF8Li2JgMvYTbByWvEGueD
6nWXlVcRG37Z/Z+npbV4NRRgSXqvURwQkeuNz68hrags1MaRFmSLVqitqzze268hjfsrh1rsS0LG
DQFghCYtGLVqEQheQiarAH/AWuOOaVdauHdWbivb+2FE5eYqaJoqoVeRub8bPy4rK7iiZYhWfu0Z
G1Kr9x4NO1UpyzQuBASBl2VOfK+yZsfMUp1XuFnNxcNFAK81i9W0hbSLIpU59cHHMDDV9FUsjnaw
a4VzOFeXKFNrZCs/TkBgZCYGOmt51ZbrgO6sAw7SgV+KjaBCsURffMizM8Vf90gEP9J225wThS+B
W/c3Af5kGGBOkHQGXPp6p/lloAvsVNg3nf7ay+oBxdc9L6fwJpQzE/igjkwv4qic90TtvSsrJjRk
XqrnuECOgZTya/JSJuqvJmQmT6tmyHQsIrKDHyc5Zvi8zAEuLbLRLPpMhddkHdfyCy30kF0SJJBN
lYEOFTybHVcVRt8b6Sxs93WulLLXTqH9LHockvmUNEexX6HpNReodXTO3gE02YorxteLZ7sapfW2
btZDu9+06vQpPKYltY6OnCVdPIYiE47wDb/YebeCcWdg6oT2mt7Lsei5iObxqQNgKxpBDS6Q4H0h
WKhNa/qbuFYZQiiXvqh/RnnzHDV7o1k0SEM1aNVoqBpvnD7x17wvn8UkrQte8yfr+zeCi87FYHcK
hvee0l6fB6gVqre3QuUQYUxrWog4M2jsoRaEKHxonQqVbdjFeLhFfiaiBzjhd0EafTlcIR/qXK6u
O3UEFsWMKgX0JnjHjO5ExXBga2PWtaptnq5dnoBUPNYZd5T/9WaH4r5NpTZMXPL7pnqeeq+FALa0
GfpltsfVHTVc/hfrp+eSOj1wlNeCEc/cqIkxDLRgLzBEtJK+Feu481WQVpFPuo1z+WoAt8/lvW7O
3kxlDtUbbSrWBmc27rOAI/y+6H0+lC76XQKK1hO6c2J70PjeC+xJsKkY4Km+ye8Dn0mgbbCHLcfO
29xQL23XEtqanG9Keo6Gb2vAXua+kCBce2gWBbyx6QcFP+3zl/BQY+WjDQPHXBnekbwICzDSdLFD
B9bZ6NHiw/Efe5Nb9DjqY8DZ7jrAuOci+067Ej4U+EhStfNmY5sZPkUMY/Z/ZIPLc6UNftwpLdYM
v/IDdBLtQ0V9W1PhRQBXIEOusV8c/k7MhH3awgtX6+9/8J2GQ2VSGomx2H0RF2fNHRK2XoDOaWm+
hDzn1sov1oHOzEKIgzh13DNDkSk6fSdNnjMZk4OhwpJgsgtycJbrAzPRcxoRG+rs+o65oJK40VKv
um5sQNego/43RnHsjhMu8d8RY0wk0zRlPTAWzsnVElLKTJAt60A2HvTu6QTE8LxYc6CdK4Vjeeya
B3XGlAzzQjdm9W3cmyh/nVsLdUToya3DEYrNyzVKuCeLcBjT2fHyJ49Nh0QXHV/LSF/sWu7t4WW0
NQ2LLw5nfNkU2f5o7L14/P8zmYsOrCCY/w66OS85qWaT9KpsHrlJET4D0G8KT+oA62DF/C+55lZV
plO9597CVU8CsFOntI3iUUEZOCSFmeabFOBYwtb+fOjhjrfQjZxruYm7hCya+FE8kj4YR4vc0f6O
doFqo7Hk5GZBqFJ6XHo4zgRIFgfyux2+kLCmw2N6Swq0MlyXZDP2zZbJpP1AJCk1mLaT72NfwXPy
+4FsWS8v7SKtEbFxO1xs8A41SJAUvV142dk0iu8alMQu6Yfj1VMtDQffnJsvsPp5GuTB7g/oQAof
tV01QvxLuyw+1uxVnjkLqFMlZ3y/t//i18sl0Hc1H/4Ccm5DY1LgyRok/sxzZ4gJkOLMIqnkyjou
Gahnffg5XHBt36/oRA6KHbqIt/xOiIh6dE+19ja+maNYLEE9Cqjo1wI1yDcBpZejMWeKwtd4bW5s
v4AS3JpxO7KGcR//sJ+UYYfxn1FvFzuQP/wwEajBZfv/9bWs7mTzhS0flLBIm2hEoEhzdn/Z1DlF
vtWAe8bCKsQcfIn5QrAh5nqeZHApi3Ozs5G4ssF+f+fBhVirrcHlRED+AcnNjDTQ9nYh/TacsCHc
urM2B9+ONRcYqkp6x4EVVdmkBTibWOKweYbwe/6r2/DuEcWn1GMN2iHU8s052NyBBVR/5HH+x8K9
PJSAJBHc5r6qlnu01tpEZ/Hg26SY3Hni5sIvP8joR973rXD6d+XAYgeGRLnplXs2iZNjZiATPLCR
I3FRSRHA0PyyNh5SNnPu7+VnqS8oXY1oB2q2D7ftnvxRla1NNqSiIbmQy4TNZy44BFs8oIYMBa0Y
a6NBrCNjbXNYsQalVpj2pm4Z7uVMsOGnYSqjdvd0llVSQ/IxOxCMji/T/fbwYndM2K+OTMKAyb5M
5hGZ5GRSVuK77twBpVxX5plHjSPp8nKRrHj9FLKNj3zbuVJ+9l1VwAvRyXceLNA9+1xSeYzaLMfe
PzWRAOIOdyXXLahnyx7eXhaJooI3nbpafpWkh0lo7teZAaRRynlbqGJA0ec4LErJkNQdXiVoMPzD
oDY4l2OO8hr/5iIVRXCT1O9y13wCpz1eJ2OL4Hll6CHxddQje5ycXUpPUE9xgSlcWBA65ZlC5k8T
x4GQFt6jLYCzmgmTUyq8jA0iEiqiBsckftuNNkCY5ExBeeL6NaYojb5YgQVxo2S+DGVWZbf3aG5o
KM8OGLUxmgfMpm4XRuk/clmhu5FDKGjMdRqHwlRJh26BfQlJgZ9Yhx4QeWmAdLid91+PYtVE3qxU
uUWQnYEc4gimS/qm3puJT97vDmi5GDMguGeEPhSCOvoxX/jZay/ooRhf/ElT1Q+DOmWUEvJTOI3O
vntW6Fdc0HY998g2HSQnqqREzNILLrexta9wBASdy7qNv9s2e2TWA5SaxywatXdJQzLNs28olnPS
r4rARTkuQ4RZfluA29Z+XJUEumcXTLYY8a0dCGu9mcIlnkOLm4b/Hoe8isKyXz3xDCbuD7o5wvt3
1Wj30Qs4Cn6umqATe8+s7ps/nE1L0XtN5B2ROuC0ugJv8f6Tb/B1GGK1NhWvdduwQbuX/W5fRQLY
Qiw9qvk9BgOhLQCAx5gqRELHlrDLkqn2zf5uLoJDCrsDAZcftcSM/VlzhZIfKPJufjkrWMF5CGoE
h4A+iPluQwdsW4c1xSALP+5bjGvCQDJ8yldDSFzHvZuiRxNWU2tK+v1Y8ZkQofAyPcmQrO+/di/i
xe9nHOQaHRx2B2XbtL/MPOeiHqtYXmCQTsT/hvbJdnP8YRSRQFrA+SW8UAuz10l9xYf1x9sRtSyy
eimOUIIFzmNO4ODLI4wD5fJzLOVWGZIgunzGjS1jGIC08Yi6vbdA/2Aqymr5bGbrQz6/uAHwK6lw
3MLZ+gH1t9kecmEKRHd2UsOPvTgKp0TlGdfBPP+DG1BgWpp9//H4aZArnv0b08lc1rsgiMkeTaQ6
WRRdD1gJ9mrPXRo1e/g9MlUq42RnUtvdnLreM/ILHPBEnvyIHR/CyDu/FldtUc1vgTQyGNwvmJs+
AiUkyuck84aBVRUufkl9gMFtjCvNMIlpZhNLoAZzf63NASbyady++VC7QgAZlKZt+0f4flba8umk
Gq8MReoiH4g60P64YNmA1qbOd8JD8GBA6W5bKbGikLyUCUJ7rvV/kIpkKdT+sCxs4ZOsrSKNtd8R
2TN/vMhMUvWap0Fja1b2sOf/tYXw7QA+GzT9WE2ONEzVQ4yLVA0hX1pmYqxtJ7bGYpKxcdrW5Woh
oreR5AB9n5RVhQZjxWR1DHkCqea2ALAVUBqsCgLaKgDviOK99LswdeNH6ZEc3mLmqEwCE9i5j60J
L7FZW1C2ZrakGgWVyw+fKVP7hfJH7jdUKVKQBIPoTsN1zJwRySFE7sQvj2TEEOfbbkJyXATs0n6p
T5iDlHlfNqLr/1eHYqtYK7OqCu8C2OarER9+WwIKZ5cKFDktobgvxPoBM+JwIgqmESzE0LI/cOJX
NfwRl6+kOlnQVxCCrGHkBnvRrRJyyZMtvJFtO7+U1RNgtaANI5fQPnt0knqV6hj9wm9jujxFuKw7
FX8IH6kQYnWLjZ0v+pg9fvxo11kRmNgQHfggxjg2ChvDSIOHV9E/WcOCTA8r/G2KKQ4+Q+nNi9xk
VwmIFFQs8+I70CF0moUFhnzYGLnpUL8j1kpO7SIx60bVXRPu2o7IGvsUb5S5m/S9aTVybSQT6YUx
RQiV055hsGkhEOSDK8klSdqk1Rn4egSCxeNYr9OYQrZ1mvqZfHL/nlWxcahoVa2M28Ckdp4bWfFi
7sUYdTq8Vbz+NharVP0CZhPfXPeWC3RjXzEU3kLVOWYlT/B5pfOIBCkhcLHLQ9Q0/47P29CdXNRv
ytekwZzEYqcsSnjifugC66iBEhZM1K+NigTL85GSR73XgQkmjwp6t6JkwdUvFdDTCYAX6LoVZFaT
ma2irHwvxE0Q/Zr0SbYFUqtuGJoyyrinZE5j11bY7qzccpZF3MsrGUgV+a6RggxFE/+y2xS4rjDd
6Tovf+DY8M/JNqRUGibQoe6um+KQbsnHcpTCI/u4X8ywOaEe+1zn46xx6WehxqjiJ05m1gw1FCZj
ewlgSxrd6et3jL1VRSTdnUEU2B1C9xmMKidYjPw6AtOPDn0WZ46LkBpZfxvo9AiF8c9cPZDhhj8b
iXTo3usVMsb4dP+5j/0OrsKYddfLFdC7NgQIgqrmulfe64p47Bo3/4vz3P1Qf0bp4ZMiHT5r6gJ3
BG1L4q6HRt1KU3sFnyom7to3wQEC6NskgyHJtQoUXFL4XB/Tdgo9dxzIuAmf6iUbLJy0pFmQSlt/
bTtTZeD3w4Pg+KxF0Gv7HzuZbCjFU1lYV/agfa4iKGxITKbwVPNvfcP+FtMLHWyjcOgPhEA1PGhq
XvcZo4UZqIovFSya5DjhD+4ZHII0rOSXFFCDC4Om4FcRp/u/XywhDsS0moFbOzuCxz7faX8zzhs3
0DLgygmpAohdsXcn3EZXpvseXOdpMJnRS6fstNqM4IV4LEMG7U/J5pZgQ0biI29/y+BzGTcUq3Up
7ztbUcBkSqxNJvRlRDqkU0jolNYpBigDLoLrHZdOBLizipGnhG+e6t8/iNmu307GiCKqmYd+tSPb
IHMU0kxRb9cIwECPAA37uRXPRm+nrj06kKeY+r5/i97+YHQgdGoHxTdW9pXvy+24n6UxcBxBb411
SeaP/h/rtJCAhjq89EutoN3lOVW1WEzBqiSYUaQe0JlclvlApaNyv7czUhDKcGqDk/CXzoEGPdG8
2Vexn5CQIEh7z0BoLtD2QHpKlVgAkETv8SDprQzVuXfpRC+4goDLR0AA3o708jQSOrO4i4JMhnz9
kpMkOLsSOe7rweHKJnGpTB9d6kgm31ckgyswbDRtCjOO2ZZjLADgpg5cpO7IKG56p7oi6psXPMgc
5Kx6FSi6KfP1x03bXDQNXYQlPGcaiEWskUyU62TNeGY2O78asbSckruDS5SOQb7YaMB/X2Tbly0Z
/abPj+z10BHGP4vrNqTFtuobntVA7amBFXF6bfn9kw5Dl53TF73qlSavgOrLawlBDgtKPuTW2umw
4TWttemqm7E17kcsn18o07rjybfn/EnZoKSD9p6pL57iFhWEjAUYuuZkQix4KAtgYvX0HHXMNCII
mE0e4ALD7a2JC8cvjWFfxO/T7UmmWVW8Uc8EAhqA3wYVYuXvf01FCrli5sWA7cxt29fS9z7R1j4b
fks8s1HvSmI2u0jxn2C1GeY/1sTYVhDbkcoWQAeAMMgsDrVAGzyDYWdrsYpuKlgkFqKmnRW7w0lI
D4SjrZntzIqz77KYV/grju2ISDcjG3WAJvJ+707moHgHDFCQOMrxpfvdDZFOeJD6sdNDQziY1E8j
MyBRI9McwhanpXPHiT81gWqPAxkBWxmZC4xpUsC+jMALB5Oct1e52isZLATuJ08ewRJLak1CrnZM
ttZc/sdKLDFxBa/KLnnAWsQHK2CwBCzuCsq1cZHI3mNKVFmlwdfUzapco8Euevn9Pd9T306YY0DC
+XtKk2dYED+eRFnWMtU5NaKWPDf/Vz2NVlmlAR+3nz70ngxONdwABcGMZIaHKK3HbyFrr5i1iLJK
vGZsFou1C3uGZC95s1Ty/pPgAAVnS5D0wNGL9p5Igp2UOzB3aOBENqqsrcLn9/L2BMRqu/OxBeIn
4AT7hl0Fa6aNS+rxndmUYdmqwNmdG03axfmKVO6S/ZLE3tcrquU9FqoYDkmJic6VJuk3en830T57
c44M0ZlMfaFjx577bpcDaKlYWp+g6gMZHHQEvwtFqP2bvpAxaHl7kZ2a54TOa3qKlzNQQktlhRB/
+/57UUsjMiAXOO6SFF1w5kfTCVur9NFPs6SazlVrEZeCq1I9xlVjQApazn2l4Qf7NCFFal9jx+GQ
HS5rVK+dk1dKSvGhOkhIul98kKUeB5H6Ej5BFZHuMOxr6BgmK0yTdQN1ljL8OiHY8ZHdpzUBls4H
ielCQnzHRXXtBb7bp2WncqzpwHl5JXXhp99UqiwEPTm2yLNNrOnCpnJU4PfgcB1xoVPqfMntd8RQ
eryBnZKDZm4RiJT8OIYLrPIng54XTSY0K48b0FK2fv4VYkEm5QrLuHeIhkXPp+8ZSnvd7ECHGZqc
HadXhUyMa4jTMCcNOqaI39rdOqotIWXOpq5CmKVaDoFsPgzv4i2l1i6w7DyxRAjYi+jrZkCSqRkm
UrmRKJohpN9GeaZ5SNGoU7A5/n4PtsEsnRsqpPr1KtxcRlk8qY5J/vtxQPoNzM4CnybPiB9LMiIw
U2edtbR7/5Y+B2Bsby57EcLsBaZZWSkG7VrUpWc+LKqxt9/M9EnqmlcDWpnR8smRGYyl2IJONYnD
TPXyRZufQB4rilx55KiKqbWM3S1Umz1PMvRgacXvZIdQZo3owfc0FOWtJjkKe6etfwyYWUKlas9V
RcmLoCr2snODLCLhdJxNH1SFKKVhT0dumxQxYxWeDSvpZGohSOXu3XNjJS17EMs6rZCZLnp+xu2T
8YMqVLuxlPMCcGq/4bj4TrT2A4+EIncZw8GthjCPozSXKvbdDDTmG/x+kPaJmPozTNJVOzDIxnmd
ohp1nkvLYKPQGMrI+mqdaiMUBcuQg0SbymtvWLZOAa2pu7zl6gMF/dGX8mNlJPxFFLjxg/Sphpop
0qcfoROkPFVciz3QUQ5Hs4wQZbIaJtBGcIadm8l+e9kEe+v+0aKlT6LumbtRFiNv0qkgpDtIfVzd
Ewna1SnWEfFVnjpWu9ob6Ux2kk+zVAXAAn08j2NRFzrGCHx5pVhTHI28emUOOTjToFAcQH8feFxW
F/9Nl8UumsdgmiRtBg+JP5m2NUYrY+JpltTod8jYk56SfZWVxndpthzODExXxoxLGhOxNBHAeD6g
VsQIdf8kgGP4587UEoz9CB4Cr7nLTprxvPKtxijnL/120ixd/fIoai8bGsp8IjepQI9xYTtgWEaW
rT3uPq4bURIQvO+nP2OTWNbX5GfPcfZr+eqlorh+IfTATiTRYEsb6PP80OTR5SPJD2F/RA103m3C
j4aBciyUebU52FU7KtREmEJ8UZRi+luQTlSlwn+F8OgPNfjDM4aOlzlXVkqhlTJLe07m5uaHMZtD
kcBT41lloiopmddQuMVfiKihmC9U4gJX/jmDVutsChrbbS+lkPD07D01a9lQ9bnwguTxFchcKQuP
/HHRl38VaFawqwVVmcYMhMFwltsT/bybBiOMsO4kOXf7B5zFAtDujJM1dAkJFGzfmB44snpn/tyE
vWgQ7StB7a85fQDBAO29N6egCtP4bdhlKFzCeK/OxyitCECjrjPf5hrkY12wqSOtAOM9Ygd0x7uZ
eMkREABOzSAb+x9PymCoxSOs7zQ5trASSG4uQFFFbFeXh2IEgL3zk90IkodrrNYzIriH53dnrbY1
a7F90U4A0UPEjjmNXtulEsTrcqLmhdFXxUHEOxB0bmn9TrCaOSRE2C6feiiedYbfJe4Jwx3jrz0E
XFiyUYz2ezXjW2VEjpAw/wcuVVlCLchfYGNm3WW6b7JxkIogW6p0kH0ZPOJ570Z5ud3ErH4xDOrk
xQsXN/E6S/X3545p+UOf4oXQoV72DdO7FWP/knpAIJSCYpfZn6Jp8FSvfVOXkREvIrSAKlCfhdiN
gmBH/UX+iHa02oZZ3VwL7hAXb70NxwTnf1Rlk06RmlTOF0m9+H2752wqCORba/yG0tUl/TUGAaeg
pRGF3TlwylFtCjzTnFaGUqKgs2dHRu5TY5gTO5809srmGFkbe9W63j3fZrP3ulNuF/FCUizxXtSY
M+UJdM4+EeGlBl1kHwgQozstUyfsU6pX+ok+gf6WnNX4WFGta9+TnYbUWQt7n2KofD2Ip48llqqo
ft3J3Z+GSaxe7PIUZmx1RhRLuKUJnLwy47bpPVZk16ajGAZvPmynhokgM9o4MGYw1cDt/tu0lFF3
E60xvbCxf5iKoTMOzFPJpaZTPj465HrbYXBSKY8k9dD/Oo0DSaMmPftAdlsFG9olpv8SKSgXibvk
lQlo6WidAZYlGoxbwfMa2YYsnp7rVAMyq1Xlmh44r04xASY7zCwEphDgclNqrg8rnsDHsKzZ7JbL
kRQePO2Z+v8vMyrT/7YnW1CvQkmvcdYoIxCjk/+/2uQnTPFg0OE0IznsEhoohl+ab1Pp4V7n2+Eo
fkObvMhAunv950pJK+LwGaBCIDDbNIErrktve/XXLHxL1EtZ41QG3nb5NIQY6DLygG0WDewfAsva
2J2DDq/u95eKIyK/MyL4qAush3eUrD/KuKEPdjz2noyb9kdqm7oKo/WlD2VCdzG2hNlQ9xfEq06V
u/PFbUg2ivj78m4REsfxMD4dVi8cYPPn9TyehD4uoWGS7tIVC5VDKeBWVXWKg7opiDcdegz0CGe4
sQFxTL4fPZkNAt2Z5Qrmctbyi2jHwTX0Y/4zfK+yq0L159YZQ79HeUmhaPwLYde4waqVxNeUIOD+
oqzD/50B1YRD+KwBp0jc/orryEvC6RNnASxS228q0bmUXcJuJ88j77G/jmR9qq8fzIQb84qfb41P
vx+Gh3Sc67mlIykT3ciYoiEnK4OCos8KxYL8vH9vWoVgcIqRGINwV9w8Jywl9nvZq/66iQosCuML
RkZxucGgc14aRqmpGfEeQsSM/TQNnYDrq1Sr5YlXla59UPPLIsV2C0M6zFnxvKv/3Un95WcNtZ1u
t0a8jYE2qppK3HuJBeuxy7OT0G4gWh08QU+kQBvWCjsGThvb5QVDhgcCDwoLKkPIBwEYcY/MdUi+
0QGJvuj8GEpDYRlZAKdsrYdVi8fBpV7A/UEOaeZ8RpgRrz3LoOm+0d51iunqxVTtYbTyNVngRHY8
DbR3CXKxMLAk+Hxf9GLoVe4M3p3990zVarvBJre+QQ8zKOQ5xaIyWk2YbjbGpjpnZ74KZYea8RzE
fHdCsTbSYTpKsQuMcgnIWVpTZxEG12c/w72+sxzZaJ7cK9aTNAr4woiUUDHVTX8cBDGWmYcmm5dC
y8AlZ9/kZvJsk4XdKVfaGGp95GXN3s383TAHG/TrJQ/D0ZmWi+Ta5KUk9CgOYk8smSDKGGipLgns
1sm8UInxYTBLy+747dNJnNf7hrU26+tVulVsc/H4rNCsolTVgitLSe+vwy75IIg5nQB8U4Hh2fzJ
MuFDnjeFhI6EF+/7meOpNHaH5ZKLkzdJ4vb9CmXB9R0Pj1HtimaAjUYwDPsuAz6/S0hOZm4etGCq
aTOVBC5hkL0HM1dM4nbxCqeHDqTPE80tjwqNA2b/7BdmA+TiAFMC7O2PaxaLQM4tiagYH/9ntJ54
iEQKl+lNt8Kb4cAJ+Uw2dlmwNfF5iXk0VKuhnsxJL3UBCzI5mVbUJCLD60Jtu5aiWOJz4WO4sL8o
eaeLGxJ2jZlOjnOsjiKJksAV89/iTnBZXaQveZPMxThruC597vRzahSn5omAjqjkfeyjQV8Q9Oa6
zvpV96Mn/MNI1wSn1W8ZR8fbgyfBejjoeXj64E0Zv5gmRtJo9N/UzZzAyjCpOz63/MlRQVkF20OR
ZuhZN/KptFhKMLiQRNMutT6edAcNsViekuyKVPgDQ5EnQ0Zh0nQRWHBnya8Wac8bGEpEgG8yjcXW
e3f87QlHAk5w9wIHmRu1TPOm9AKwcnb07hN9M/uRPBtxogQRpthZXh7Xh4i0rX6oQrDf4issk0i1
7HeGTqADHaBqiefrta7C6V5KpvBaGxDqm9fmfxZyh+1+tvQgNr7vbS8uN8JPHH33IcmLm1BcEE11
PuzDm3GTExbxYR8YY0xLmzJhRe4ww4OFBZ8YSFH83Wv4DsnDIURXaBDMVbIg8Ji4reFoLcq4Rzdu
M8mcmz8Gk85ESjwjrBM3s6zf0SVXztUi10kbqdCuq37ldl+az85+ev8LMiTL/zk5AAZZqg7t4QaB
7QBHIWdp+OaSGFfOQKLZ06LZH8TkT3xjf4OU5PAe+H5aFLLzB3YfsSYhnkbehfLH10M1NsCLeqWo
3hVq5oe6y3O4Kwk1r8eN5nSdNRicnWgVGe4vp43Goq0JD37+7MpnaLaVz0PWMGO1bUGe4C0oNSVy
tRywj+d4ZtjUg/BuQX+O4872elm9UkhjuCommhTrU46RCi5hcaMBgdG20TKiQngR9PFJEywtgqhD
rCTBQsR6q5E40JUfPxupQTQJ4jyU808nepV0ThY4QbCNdhO05w9rBNZ8XGR7Thfa1IPOat+yy/tK
gl5XcvTPFZM9i5jILf3shg4FDc+brGQCUN+jQ9EHIlRLQM8z0AnPJgg0lAjXMbhu0lnEXWthlSYt
qg3f9hpesat9ARf9Ax6Yv2d/KTR3g7w0tThtq+IRTU6SXVxYSqTneoa5Wp/PyTWgy6ZpnqfqejHd
h9+4LDIcPtb1fuz1CUAgQf7+QxPcrSXK8VED7tzuNQAm+MYBvwEHFJkXafzpE58HCX+tO1ouH6N0
8raNHcrT50mIWnecXfurg26MeRm3f2IGidkDi2zFuleYv9RIXF5Tn+Qv0heB1rC/eUMJAGMS9Cjm
EX0EfXJj80kYvl+Az8K243FUVHlZYc7gAgR+ZXTblyiXEx+Bn956D/jHay1bfPxw4GcgP9n+kWu0
NWhuFfMpwIhU1rUV2cKOLDMQJ+5kbUc8ln/37M5kixOT2hkxmMgpiMwoka2e1Y+zlWnv+YpfJp9S
Ps4JjoFyZp2Hn7geZ3zdSVBIBu1QNf7+Nwg1d7EVu73clKlmDTH9Uz6CDhSeYh/G4x59aM9Rf86P
3j0CtQNmdhLMXgjFHn+Jr57KU2fh3pqJOKbvRd07OtKCVt85hP/3EVPkTBjFCYKg4MvvELJrxQBm
IZ0GTmUSB6qZWRs6X/3ztxVArglRMekvbEwYEzjxeIc6e6zFHPgvE+RNko8mx5Jt7Rv6jYO1K/DB
x8GsyUHvRe/WZpvEnm8zr2SwYPCUK8+2rNgkLCXhfmOjoRJQ1Oe0V/p1TxvsHIx4yd/OBwQxEw0g
f43ZXrM4BCl4APftDw8DeXkXguROL9CQhgi1x/qse5wUlQOw77cMK2VRPUBKuKRWy/jyDCBI3rRy
ViedMPsS8ZwjVNJXuiLpkcj7I/HihrDcWqo0EU5UJDIsfRjCg53SkcXldEwZ+5UjFj4RH7FZJ9xz
bBdjVadQs+YMV6Q7Trs6hBvlYfTIX/O3rFknzM8hQy7OetEfGirzk+IHR7m10LMfmuQRa7nFI8U4
OgMrB+FmZn/D5NiG2qXq9zf28e2s0bDnMagu+hg74nxveD3EPIdcBtEPChrL+/gMeR1vlVMvXm7z
8rrFulGTPkRDoH4OZJOmLx47JiVHwn3GsmdiMmoDa2ghjtC/QKaz9XE3av7OeC9jNxzqeDvOZmrp
6tWspOGu/fTuqZYgVGgCy7J5yc3kCByFvxr3E0EkNBKcjpk1u08HN7GywK9XDDeKV4X+DRg25t3i
bfUD0LNJxTULP0/8DvzFW6DOFJRHcuGtY2EQkJWY5JYwaYmWRyWjY9M/oWB8ryM8XuVAEF0tmdtV
n0SP29JCApKY+Zbe09XLA3oHUjLY5uS2di7OpAPWU2sQxjjO8aQ1KqAmFjsE3INDeVU9srNGkvT3
xippD5kpNRJH59026qFd/JDaMwuWsITX8q4pYOj8j+49FMw4fFpMBH3pVJvOQuyJ5sOv83c6d2UG
ngojaHAfI7KrnfD221J1njxMJhWuskMD9R0C+gCMs7qmzbLICcxolwZie/hDcihMj1GB6OihaxSQ
C7YiGW6f71tsd/27H7tX/lNV0ykD4OXAuKISFA7o2mnReyo1eVJuBzoMVOFQlCjH4yk0vjedrzkm
LgZRY2Hytbq7HGeJT2C3Q0SYpN/CP9zI0H38B/Cce28WoMkthv1kTHtOOZBTASB5FJkr5HCpfkjV
YdFwgE8GjR5VXyNjVmic+lJs9g679FtXh37RpiDEurhFLlyfDm5/RDHvHgLT78Xp2EkeH0Hno8zv
Hb3Ooayi6NvxmpaDA144TuDc8E5elL/QdjDpdjkhIfeN8yDeFnWvDeUpOWD6or682jbCryxOxmdx
5Y9hpQBAiN+/PvKypKi5atdkTK/JzJL5Y+IsSLxUq29rWhsYIXMbxjpRXQKah1MFUn0/EmgsYt7p
WCXFCfUkzpCjpWg4gWq/mqi2mdl/qvicnQXHQ6Ijn0yXBXwDpf9DfzSDefeYp8pH/9fOkiyaHVli
aWiIKiji+QRzQi47NDPsCYYZZnHNXLO58b89ilr5onglBBUaZYojoRwz8Gx/iq1b91unLaAdUIgb
uc7GGKwjQIn7a1pujaY65DMIzslE9MgGGie9V98XZoj2PU8gT1LU1Jcx87FUYNN0j5DjbnjcErLY
txBqRA/PTThJodxYqJDtBQ+prr9eyVDxi1mehefR7p0VzLt9xwX1QMQZV5rh+SxSuME0EkoF79Eq
fIZA3tNREsP+pdxYeuczqi9KaqC+0bUyqiHqk2rTQpZXK5/K4nKLOX+3bupeZt1k3W6OBF0mbP95
850lxu36je/itH032C2BN1nkwZ/6X7gWnwoOvKZPLr4Y9dJ0ZerdBJ2jltno/h2bHTJ+yIedXJ66
tusKsYeap9o5v26fl8W1Ym1DVFh4l0MBnMO2c36Fri1eLBTsTgihTUgvGv5/Q144kgCg2jjsmigu
WmLXClth8brj11TV4YivPOyhrrqQACD9a1RI+iYDxNYP5Y3XbLgdxz2X9rNb+nhP0KUZXTnrs0kK
xEahSXqNWE0Rh7GBcYgumKGsh2/SF8asdYJ0Tb/FVhc4l2dJfNqy+BXtNFcDjM/0t8TcKB1O8fYM
JHpyIMydo8FIlkscU0m0qcXpqabQOUXrgyeiFvx3U2gjeZndgHD3QukZ87ovneP8w+Zx8c4yQEOV
jh2CIQYlCxNEqb7hdbwrwTBEhBpy9IutSKP1ZZH2Fxn86Su0umk/fvHs/Ec/TEsnKHqjZFxvtbmg
pOHXBd53S7+OgN3L8PQUHblxPEGWzoOCaaLX3IyGUWqKgwzLFM+2r3d2Wiv7KqLxdwnX3A6L3FEA
qRsWT0y33X9fSIqxl9HD69jMJ6kSg7RNJdxi/meFeMKn67gTv9JJ6Pf2sTAQsuAxuFGk60xw+nVd
xTViBn5Sr20yDziYkr4iQkNZEjD8bsrU3Bkk+N5DFKyRQINk9QLNIvgOHu4EKopnonalLz8K8sTG
97rZgR/8s7jo9edVE//y6bM18CdITFw0D5/evlbBmeQ/jFYOJz7QCka56eQS0I+4rPvWdCGHSTXP
OV/pXjGPE4G/sXE5Eb+B2HAfs+EQiQT7K2CFBUw+daf1qA68JV1lIO3EjqUERSmMRwNBlhsmFYqu
9dRrJkLsusEhXNcpbiLLjOpJZY+m4/qtgKoyh7FmBysJ99JGlItqMdsmvNCKbldSf4W52FI0dug9
rvFLJcTHnXdrJzU207VPDqDsoLGZvXwH5HfZnh8YxG5kHYooJBV67CI8zLbvonDUf3qJSPx/PHtl
1VUJnlRCnL5/Dq6xLBo9icjcI7dMEEj42/dqiQvZMRbX+3tgDWObBWQ6r2TyyIkRBB9Pe8IeGkxR
JRGGC2OU0DpY8QKF+K/JfvwelGBAm0VYJtt5aMdgJsZGHu6IzBorOEEGXVmi48VaEI8in/6svW8R
N91zd8LhcdEk1mF2/93HLapsCCxXv0fdkJ9iEACQ6bFjDWbGnlPEx0AaNJJ+QRqK3sTqHcY40k10
ttR1heD1wr7FJPri8AX2+boL4PilmP1a6/ta4wcxd3I3ded/OZHG2NGddBe5b4RiDDq3F+Ow51ro
LLOUWufz8KXqLv2z40TRI1E1gEnOZ0DRmFQRhuZ6BFpjAZRFZp5SEwAqluoZpFhZNDTW6eOBGFLY
0w0PMDQT/X6PoY8g3RKTCdWGUGrjTnMfvq66KXurzP4mRuglqKaW9bqSz2o0QinVnD9vmi2Y9hjx
4DF4GcWvVCNwWfOXLhtI1zq2uvGhSoOx/ZC3LqkE1jQWgnA5y+4JcDpni4VMy0NJasIKtDBKxxUf
qg3JhZDjhKLPTlsx439TryJPuVklqE1feKF2mBtPIyuhIVCjczeYoH/wwcChgBEa+fsjOobEwAaQ
I+HaPATKOKFH7l5Mfhh3rZ6G3Vk/SjuZWks72QpHqK3xQBemQ66gs7Fp/wnQhpFV5/MgVAMgHOJ3
VHY8FyL4qXT8cOFqRKv3CCCdQrlsZJayivH+Kp8a4y99RjqX48jcspZEaU2ElsPcWJFWoZzEwRzA
3ZaPlMtlqFiBknWmz0T0SruzSpbtXZIGG8fVbTrVkzmTGsfPFSa4wHeXf9XqbmAJMCXgt1+erHsT
0cw46WeHMN0JZlX3wJZ4VHONvUaHO9RKwowwBvx1nEgeWwSPKkoVltLLjvRVbz5Xc+A2HKqubyqS
b8hIpYCDQVWdgb6gmu3UO8WWHeXCbll56LFt98cBKrD9nDE8WNvOJ3qghyPOTzHOrve/s6UZ7Wow
XHjIlBH3oCv7MjwTiWu5CvHLzHMwnABBSUgi8F8CqWuSYk7YrJ+TxeikDZMjitfqmWCizFlfoaIZ
QNQPNDeGgR31QUqIfZE7TJnzSjlEjvuFoZJG2LapbWxSGZxCo/1Ceuwme6iro36UGJrljJilOcS9
zZYyoWqLif/XjQaufCHOKnUNGi2YZAzsQ+aY51n/HR/xamaLj3O7nIqMleFzjIO//tDNaZzTOafd
EWJoj4u6OMC3OQpk/pZYeoqoGsDB/pgtO7GMyNzydlqqje69hv1clXsLK6z4l/aDHPYpkkF55IAd
gNbdSf3olOvkPBwuzW5JzEUsSAd3k2Hi67+tTfBQh7hGs7OOXnwtUy/LvCdACGLMskGXlgm8B78f
wDatHrEw+4EHeptIeey2bATbPbabNWZ7mDoQf4zzWDbvgIVGB64VwLTzJOIHTc277p6iZhf7iDUM
CzJ221hu5heCoZFxPQYidB6EOBAgMc7UVezHyilc7g0l8dDVKX5Y40DWnGDIHmPLqtZ5gpzxWXJW
RZEMYEWOj0ZSglswevAvWyA/k45D9tDOiXwGGiNxw2cizChMRHMUtgK0aRTc3pFErnlWe0x7L7fA
YLm6zcejmcDqbiEvEvo4vqnbXewAfDwFMjqNWSFOyQ3P/lGCB9QmbTcl2S/cwS33xWFjqsLsnhMq
Q+UbZzy848QStIwamxHIjyP3Pqisdjk4i4H7I/jDe4fmDA+xN5o0QqnmvrxgfSCcPUeUFL7AHbCL
N1IPvtr8yrXtxclKUanDMccPiPpGbpZV6WdfbYfoTcZ6/YbtfX+cTV72f4dWk7dO4dWO6GLRLg73
ppVMclUQXLCXbLeiiJuYJjBSSxS/O5qrkY/6NKD3YacSSbgrv+etDgxIdZ8wgHu7Gm8FiAyimr0i
suhCCzPitrupQEmZ0cj4UZuBaoEUT4QDlb/IlPG/Dz2imxkxRRcLxh8oGcT2PhA/1YTthQ7TwsLK
yvWi2/Qq+d30OOSyULT5FpHAk1r27fvyvt1debiomUGZfbXXRWuSPEKFsU82hUtxsjKYeag5kYHT
qbs0KzEWpfBphFltYS2Ao1nleWQ7ygBLMwh3o/0oaG7yA4SreCeKZozYiaYqk+7/Qpz5YsTK/8am
EaripzKy4jh12BxqrbFRsiMKjQnfhCNxKtnSTtPWtypQkgjjCAYzJatR+MREKDVS7m3r59Q1sO5+
Y17tUWschswBn0xbA8HD5a2YTVjQACKqkVj1/TugMBCEPyLhvzk4mll/MRdGgEpGywowvn1gJVeh
agasvkvFf0rpE5DR8cm/oW2529T4kTrhK7qrJ9TeLNny3dPbie+d6wa058HWUPfLRChu8OyvGWgW
TcKGW2AC4i0aiR5cjX0I+PXcku3kjinWysA1iGdeJ0ZhuMqaEEgPMoRzjHAluu0X2uC7mT17LrQF
yHR29vr3ecuaJDZr/YTycz6ijBfroSBGwlH/V7GgUoQYXhDv/AVj7DCFc4YROIgER+9srBZVUzJk
xGsG+q3sgpFwLUCa5TbRdkYof9TYBXDdHGf//fwc9qKwNQYzgsuxoCRByvHAJ72YeIC5NXHeQWBw
niMLR09YwJR5yOx3w0whLoxmliYV7ypiTUoq8faxf0TuSDdytURLGOdU0O/8weSljhksB9/8iJsr
kRQgqe3RgWvyK5EWFz04BFfdmVKT9jiPCtBKjdqqylJApz47XA3wFNDEZBZg/DKqIUSouy51L1Nf
n2nZwiauMrkB1hX940CFzgJFyFIhNxC50hC0Z5uYT+7B0ArvTICg8xnCdxq7yb8QtXwJ585YEtIV
wAo9aQPVa3Z5hK21ufzqwIj4tsbT3k89rOd6VpdRtt1Y0OCK13wfUVVNXUgoZSUOBogibbp6SyeO
hfgTg5ih8H00e0lpTRifUnxGU04Vq4sb8LcNvRJtzVKEiJq4oqU0zssKVaGthajv1ktly7bq0lMS
natTQ70IWDo3EveJ8Odiip1VjDXW32ymSzlKskePgyREIevbM2Pd2zab+dKYgU0oMB9HTurXGWfW
ZuQniraybcm6D1C2hPqCvD3NpKzR4uFoEw9bOhBQbL7dRn6y0ImOJuzjVhX2LbFQ6LAbwp/g/fr7
JMNNprP5CWLwn9dU/nfkRjaRUImmesWRxkcXV2+rhkRbteXnFPCa5seE2PoEogcxI0t0A/voTvBm
1LUCmtxnnGH49djXl8PrTIGtSdJlEfZG/LrVmstlMKhfUKcpniLIb1rbzZTq5geAHms+nLjpy9fu
ZWWy3cLOWirhzkEq5hoQHKO/rEyfGs3H2kuClIdhdf7uaLowm16ETtW2TCoSJDyY8EU5nr472/iK
5/YdGvCBzc6KpToXUvdm6FCFLIKoo8QzSiW/jM3a9o8p5/22nJv03CnkthwSkDXHR9y0J7T2ackj
tcSt+vQGzqIfIJ888haVetZpdgyOf2FAdg6GmkETtk6zx8LXTsEx68Ro8+V1Ca019fnggtenPYZF
CU/bVqKzJqFIpzim1kEjc+A2lW7nIYjXTSGNZ5qhE+LHtQbdXquKvlmKB/JxDRrAHbedtXg5osoo
MgOOv7U0Q+xAJ0s/KSmi7JAVrq7MTyJtiHTDmV7YM4sVAX2DQxBaj0DSd8U8ReImwkCLYX+r7TMq
q1W5KtCus0uzZUeOh5eeucDRBsr86X5zyC+xDVY9RJ212t0Za/te5rOjg0PkDoiAv9HWUv1TsSSx
9iuf/oF2XCZ51QUzIOIpWk9uJfxCiaUbo4sgQkALy5Ft0qq7gwiAVsFw3rw3id7krtaQyhaoMFPf
htp3PmrUYoV9+OIu5oOOMW5ExspEQe4vwKtUcrMCyjm4fZAmJ3vnewn8xPJ70Tiy/qQYB63JHYhC
+1kjPRBQrZIYF6T/G/qkGbgBK67EEyVgWgcNnsz6qr7PsPRYDXvox1a3aqWs+z9pz4molzc9Jdse
mbjx8K6QCkJsM5aXYsQ9kkBHtfZ+aW9RddKgZ4IOlK+u5NFSTcqRDGTd+PLzmYhKAxL1xwxq/Xc8
v9mJDL7MLtSw+CQF4NKvtLWZx2Hy8BxqvLPP/CVp4pZqTKFkOrgkUJOAT75bmJj5+69BZx1OWgc3
7KMZeM1mecbeW/6quHOALlukVSD02YJkn8pSGEf2K7MQYQFWlPA0ThMum7raSSCsKG29lexVVR55
q+AoAHu2H1/bnHuh252CLuhsZLhahkA87zVSay+VvMfsVmfYzJUw0I1pntgSUxUx/MHyIsfia/G7
ZQtVYGlfwwy05KaG14bf0Neo+eAA0Gse2O23bTEohrIQbUqb/JsuoCpmZfPDkxhbEZ8J3j5UYbYF
H3a2/hXLETk+n1XFuS9qxLCaT7b/D+TrTuk+YW2Jc0k50WDNkDr2qRE9bd0dQrlRongAL8ozeGhZ
JqO/b0fpAOM+EmM/6PjZ/pQPqwSmEPWfLWNAaqxS0un9JynOQbR/ZEQtbwBOWulEkVYYU0jd1h1l
mxjHxpfMewPjFl4PAO1X+RC+NpHaUgJ3DnpPewnxEJrzFmRbqq8b5ZCjh7ybgBFJC8V3FVSMZMqW
ZIkqBEtiuCA0xHmas3+Ygp2G7Oh09KiwcKfEZwBpSFb7xR7xHhuDoonoNF/nbXvzCAnhzmky2v8r
Uy7kphFSKlsBP22oTyZyaeSPDV3WldZU6m4QvG2NQoytWyVyEc+VljulUEB2abS/TuptzcKNlYf/
zUyoMRPHjqxp1n/jGYG0Xgb1JA+pZzbkkho5jjkZWupm0OEupCovQcbHmra7nBv2Z2a+3Cfb8oUZ
snr5BYBhNxtorSeax94Wa4Ep946v/IiHAKrWf+cDvXtBKiimoG38o8gg6QgAAD8gZu85GsVq5L/p
eWVUxPH7C/NQXYzUEkIoA5uPlJ65iIx0x5XsubBSa6c7PhlxgQ4faxDhOD/4mxdT8V29emvQtW45
KREOJ955m+HREpch4ff4jucoN/zijmKisdtAcPFDxJTri3y/UFGbbAyFwAyN2nSBif0swFCO0gW1
Yr45cD9aoQ0iufi+i325IYCZ87OZ4iSVc7nAiHINe0yoDvp/UOv+ot+gZwol+da0fUEWeLy5hr3C
eTA1eBfOjPmqshxZxMpXC/U3tNEKJC9lBI0A8blsTpyEAXtPyrBgpqaaAalKOtMU5qIpGGJ6Hhhw
QQ2N3XGBanjCTA3Aw8Q7BnPECaaBipQsbPyL/UKu5xuD/97pGKSopIi9p5REq2YjOt0GahN61NEb
bgmLyI7vg6ZKZiCv+bSyAINmaWw7nlKqj2U5q2qBbFY0MS2KhnowbXRY8dWyUZA1f9pkGu0kPdr4
pUQzo2Ikt9eoJYx4SByBxLRjt1eTjS3z7ogN4NzE+BCfzL80LAq2EodaIf6HBAsFC3UhMvugwkD/
7qNuxQq8Y51i27GYy/ZG7gtbkByuWn8TzYb2J/W9T3WnvMg+QvGQ60tt2xl8uOQXZuN7GxuogNja
aOAIBylwk9p/GMobkGxBvTqzzkM6rrdQ2ePDj0UQiYMrQ0rnI5bEqZ+ry/NsCW975klP/+edT8rl
gBpqFyw7+V1NGpOnHB0Dlzr4ANtcDyeVgAefCO9+eOX9vuBsi53YgWWnank9UfFL9sr1cVmASO6n
aBWgRKMugMyDTvXHjDT7AYFGp2OjzWoThBQAIxzN+BHKqrv31SeDigoTBf9vT95adKE8sm098ML+
N9ds6lvZU3Y/gOqhAmXHVuhQvnfboowpZmJ5fLYx6N08sCgpY1oR3LE7G+980x9PRnKZKlRZzZK8
vJQPuqWk5N4JRk3zBWN1xTHHT9nwlUxRAlM3WiBBHae6wEeRW0c9ABh+tE/7ljZaAllPROIb2pbN
6iy1QHwXu5bbqiI7Lt383C9NKuSHycoQ+S79AV+jXRWHaqW9rCF2kWAN5jiReq7prXse/6pl5iVj
nm8anJVPsWhxIcGTvGyqtPh72xs/t5H/LDq7VPbyGpRnlC9TmIgT6oZhrdviR+X3Zd4cALGNO2MZ
DzRSv7SUkkDTlxy9Vs9nxDOQRGYcgZWRVOop2dLeMSW2Uy9YxUn6BhIRpFHsFiNRKLiAKckN0N1m
7X8TuN6uChVTZO/4fbxz785TwIxlyZXvwTXODurwt9iItV9CstK/bzycUM2ET+/wd9BwY7qg236Y
IODV8y2Ucx0lgX4TBElOSxGdHrWI9EamNNhj/iJZnSYPF1d7e46NBwPifwSyzloW8ckHNpgLv9lL
RYkCchPttrQ6GzqToz62b7q3Np5MhGZt2kO8L3+rcttE8/4niBVYakGAZTIQuOtf+axdZbpBtHPX
EZOWFROpdyluzKx4GgbrKXWLyM0ZUKZ0mckV7o+oOHE3RkUMv/koyTf4Mz0QhPvqtqV3HHbmdRRn
1w9A6Rqpz/Jo9azltTrOdOAn0ZDI1m6olzFDp4E6qKLYP5VBuOawSNA5mPHoARmAo2djccDhDcsR
wfDFEEXRfYqG/T4a/JSltNqW0yAL9/If+oqBYd89a/muJ8rP5qdYpby5rF3x91QvKTUzji7WQD+R
HAfwN8WohWqBANpvdy1jEFm2uZXadm/l7RN+x4H/H6ZvKpUFLtkMgD1yFVrgW0e0uyvYOTzZY3XZ
XzUc+TfB1CNGkhdnRz0S97g2LyrGIwrhGFAImW3gHzry5qZtC9hEVVp200Y3GumaxClv/w88MGss
dVOxKJ7YJfZFwp9xVThLv6hUHOy8ldC38Fi9hAiWbgt2ZRue2BCZRw/i3CyuSu4N0OhIR1I7LXZx
L5IcwwcJBk+EpIWVhDEo6fl3hrALxxe+SDTdUSfqPrwlftYkCWHaYdzV4O1LZtnkxze4GAuiSjnd
QUzUhQxNQ2tg/fX6U+wRLYUejJVf0cDaaj9PDUcQTGjXsgc8te4ekHTNfkL+HaBL/Hu2Gh4ZlDux
Fd7F2dtrFQE14c+20De06sBmPQHQpm1ztD8rY6NqQpxGWN43iygo/YmYXYyYTnhQOgDVCqme3CIJ
LRX1hgo6yr+ws4zo7FKIVK5TmLcjuLnTNVNBHFZ7mEmPaUzG+ufV7tvt/eyp1QmIoFx9IjlE4Z2M
jXVhbmjTwrF+mvfQikV9C16JkIMYQjhI826hT4Qd3YQqkJSK+w/Du6B7S+lUvBLSA5cMx8e6oARt
leYrx87y4ds5tR63By0xiHtWXija9v3yx2IM9P3sZjiXk5rKHEYnolVP8ws4ej94boQhznOjLdUr
3gV95VbFQlYfIiwUiVrq92IV5ZRf0ufBS1iWQzOA1EKytyXI9pw+a3jozVoGJ4YcilXjGAhFuzbR
2DA5RZRpQFA4FPR3ORJ0KY+BFVpe2NnBOLE9/DAFt9ptvzHgXask5D6l/ZsF6EE4z8lI0S+U2raP
RVTGuJ23eEC0oPunYRwqc6qLjY2jF1kYAZfckpLHT+EGXZr7yiN3ge8L02f9MJc5UxOrjeIqMJio
gWTFjC7zJJ+4lATHZr0vw+b3mlKuGIhdascsF0TKzDw8z+taXgD6M0auoKMbZUpKwq3Ry66ciGMv
0NfzQ8xmOMs4WGAheX1qnpQCcrs6oXHIY4tctTMBJLXlV1LnbobpPovHIuxgGG05Er92u7bFpC3v
yrB43+jqdGkUKXGaWQGFaPtLuMdAE2VmiIkxYqTLHFYTXbbIMsFiFdHixhaaqFE+2mk9I+riW4m8
1ZGlVppeMDzVCmIKWYbWIPjOu4iXAAXh4PN7PPrX1jeA+1eixsUND7m7jIEwl2yK76ja6vFgBm6I
rgbv9BW8Uo0R3hCZV4JTEqQSMvL/JTADO8l9Wo1lOLIv9f4bPta0W2lvj7pPDLfQErW1oT8KOzsI
9MKLMfCN47FmXOixxgXIdYNYXKBCKIB+2RNZaZbNZKMI9n0ZKng3JqFOILD2OH0IWnfFnKtL+Dtl
AwgIzhEo/qX1H9EwdXSAbQRnndWmJ/77OIZgG0Luobz62uf+3dLswEMlqVlUepXWm140WscfDsop
dD9VCF0QNI3iQtr7jIOemNFJBb5/tQKnEyOuLZ0yoOIudCUL9GhMvMqyKYZOvcWID7vlLuGAh8cl
tXWO5flRAaDpe+tAf3guznUuFd6wZPRSGPMg7RsrnyeQsa37jBGlBHNn249dbtChLHx1vFAR4VEo
YhTuMuNbkrBFWllXz5Rk7ku6UH2EOYmhT7oynLQjjbo5m9/YSkszLXA31drWTcbPigp3xGySHIQI
AtSaiqG0FZ5KXWENut6h3zU7uBjAQ2C1nn6kvu3qprYs0muQnTeepVQuQ165NIU9JPDyJNu9R06H
CsUO63bXI5OdgVMTo3RYv3VGn0RmlNOwI5oLUcGl0H5xd/Syr+SNxgcZqUR0A9uECZJhI0MkfbdF
Z9asmLk2Wc5A3w2LdjN8yOPkUa75rXkUzBmLQLOqOYnSvIuMSMJ+oHuD6QdwPfisZzl7hNcGo/Z6
z1pfxB2FIX5jNXXSheiw0zcq8V9dqgSRJetLnUsvWV6eZcoIIHGL3rkyo0oP/UmdQIHUbTm2xbxR
FNE/i31i3Og8BZlm9Z+Cz6HAUUXU3K09AtMoKDoSPjqO8VcGMVITstwiz2p798UJdZ9Gp7ZhueVc
VmG6SMudugu1W3kCi4mW3kXKDOEQDGdd53rPQmhXs8XwDmw6Cub8NaVtWdkyFJOE7c+mgQFTbTXf
IJb+o2qUurwqLmghM+DvVsfr7XpEADatdooMmuCqD1wwIs+6W9AmUwTJpMpIP6uIJNs7tE5LFKOU
LrUenvprE3DZhbygQ4ouQKkmMNz1rqpsPC0GAsE8Jk3MGwYrnasMjsAxumCdPMoo5Be9WRQ8sJhZ
kjIKLNpC1G3EKHyJSenrIHkEfR17AFeddntzkymVFIBo/7AzKk7G3j97Hc6QG/OLZ9Di++ocHJBG
/x8vFrbHzpkeepvv4/S4sosZj8bznT4QE0XH/FzcHnTxbi0x5eZ7RPzPf2VEgQJI/X+uwnvdAokO
S68PCsnEbJpZ1M14XqJ6own6gei+zOhIjO1ZyQ3/hZJX/M0aSrb/8YmQ1TysJ2zNZTxwp2KKAOA1
RXFVtwOqoLUmfc/bkdEfLewfnPU7gFjv/okUHQcna3O61H23ypCW9dCRCABggIca1HTrnX1P8Ikp
RIxPNulN7QgbBeEKRSLmGAv94z6eV6CVO9ylIJiMS1WATlOfLy1hdydIknvH7JL3K3PTmlTMQK1w
aI31oh7sagVitzyhmUsPDDX6QJ2fP1WdjtWwQoOHfM8qv703/iRNCTpuptPkj0DRUnZMXVG7BA58
yZdhylK2NELJOR7JQYmgyF+35KDHewtXBq59CUAVpjVCKwMWoMZyipFJU1vZSuqBgM5Gn1uFD6qH
dgdXc103AUztFr0+nE3xDnCIV9QYAEOYzqX6/NLa4qu0FRtwM8R0VsWylD7e9/vWZA+xI8gy/PBV
0A1PxQ90Lpfv4eDH+ASi4vVhVucCvqNvGV/Tp077EFVcZUAbUtFuCRnAWOuHDDya6z3hz0olXfaD
amnlAdBSnY9Ehxo+vD+bfuFZJJyxpUxKh7UbBJIP94S1iCYoIe/CO1aaEr1RKziE5rM6XazI5Nc0
ImeMih+tWpLcW0YWcNHNTjjX5Sh9o5GQbLObOCxMQA/F6f4qfyUIjI9sVTdaauzEZ1eYwqjOB1kz
bAzCKVyKiOIXeBU3DrIyuhckF2CsTuaWQA5M9yN1FKRVacLOkcqk6dtfknFDRqyYgTWNFNecPDlH
PHHsxjw2SvNH02sU2em4VXoACdwoLZZg5FiRJNJLIGfCI+9oes5hULm7eDgKBq+0HZ8NCu2G6BZJ
wvvzAMzAZedjv0olE5JI27fkzOjvSG+SI59EcPQ3cGtoCJ5Ct8MbtC+MgK4/FzuM449oAg1HLrai
x/b+HuIoarpEEGavPrr3tWVg/AMBRcBMYPDdMpceKA9OZ89XUWtL9a15f6XU9coukvmgeB93oa2Y
JazhGZoO5NaszxbbmmAin8da02t0Af61kfQj1nhDCU4q9Si+TAXpfjqXpfpscv6VVYyVdKdY6ZJh
nQIlAunT2N3f8r2d5/kBlWsHICdTK2fPWUDcO6bC9pTAyQMPbKZYuIVR3ULvx7jmFE8exdRyK0RW
/7TWEal3ptFD2QF+3vzr8h7UG0Rkdptj8MWEWdLqYkSr7YhNoUmXvn7TW2nX0hyaf5tHt5ReJGxP
ytPc8Cz499F6mxa46JZh8ppOxo0Qcci6NS4EKrEZiAPEuA0Y61Y0Trt1lM7E0fueC29apaEYG+W/
DQ3CXp+ew9I2hsz0lUmW59DujS4KoHWQik7z9ogZ27CcH23HLv8vxh9kLDKKBhHe2rv1vTamA/Nl
OMculJrCIddWRgtFoMCZfLqVGFXp8gwdC1ets4b3XZpAkAjLJZqMOUxQobA1RXF2AvyeYV/YbzuI
8e6EZP7C08zHJh2LeeMwvFT6jMEUtUZ0omNW4zsJArw92azQnW+vLKcLFGVKeY6wf+RDaVuY+xn6
ywoOsXTzq1tus5P9XUOZxKGIKcoGfvhLQHWlQcFL2N6xq+V+WtIyJZiH075nnmnccKyl0A0Ls1jr
j+am00G7std8KFWEZtcLosU9dEtkk+kqn2M5bmRuw4bQJdVEaldSA8aua36INwLE3Yuv9bSqlcyA
8r1WC4CV3yLVblvABc4LC1cLd0JxbMwDID7RVvG47l2Eji1BQWu06nADMAPIUMZ5vw6KhIG1YmEn
Kix4NWnxDbOIZyfIAqT0YV+C6BfttdT3SUgFfFqzhbkdAokvsZezGVywUpT86ifwk43Gbn0KYYq9
tu754J+XwLjEWl8k5PyJAWzBQ4ijisNkd01zqyKRRx713duBIHIg0uOoGbCFfm/uh4HkIR677d3W
DLmSTWcy1apHbQSsFZd06mXdELMfFyjzMdTlT293RplQoNIuGg/5qGeT4WKfRh/5r8DCwnRvEBX8
8zlyhEnelk9Mw9rtkuxP2GMwcLWiv0jnm9nKVcg7mHlvRqJ0mA95FznCYJwCFeVHfsdh4WYrqSL+
L9l3LsdS9P3YUZIQXo3gkZESR+Bl4zj3wYGiMx1qcQRORlsAP5NPDuL4MjpjNEUq20Pj5YgrWQ3C
07GRFRXfp/sMlBbBkwNrwvAItR7vZid4Jk+gY5rBKyUnTU1IVpSAT6pWNChZwdC++JRlfrRw/qoA
hr1P2qzTYIEsRQlt0u3yVhrVdjbkVIyh6+yip+HTw11xtN5N6XOuHNJrk9ZLU/zGztqzxH8IMSAw
UVGygjiBH1gi+BPHJF5j7dUyYH4yRh38UO8iupH5ILKJIIPG8cQVFCt8r7pBP3YKGJ+OfO2RqNN6
4axRnW9vOog07Ptqp75BbHyJcU5NEtVMg1zEN2OFx4+9LFoyMhWs/4B1csMFQfU2LUOQKsau8CiU
gGU5jtEDY8w57UYb9itAaJLjBhbXm8nPuV92/x6e/r5nHxW6qojz6u5Yl+ni0KUz5306GnQ25CVW
MX0988ynvDKKAHwItABJ/LOMo4UudjQkGMaUpndne/Z2ruCfTaUVv1iU538Zzr10rfWQxqGW56jS
o51e+k6Pk+bin+LiHXfq6YFclChsq1wJAatFgQz4SCz6HyjrZFkwORuGxmylfxuanMc71S/hzzId
cbQgQO0Br6rED/jY0nwt1Psfy8MNCFVgutRrUYqBQoiK6NfWHu6SYJGAS7jYC6V7KyX+lwJF7E7+
O8G1FOzWTgX25OIdhS4ffEOcXsJk+xy1VLZl+h2qXByLAdFhm50nDKV7dg5Rbjaphh9U/u03cuQ0
x3kybeuK2vjlobjsQfxMmc4tEPlnpq2m0AdvaFXMxpcPD3zpTIR0YGF/kQgWxvPNrOWUPNJNvcbS
hl4yQSmvlQerrfhMJGiPuVf6f3aAuqWYhFIeedNc6Nv6IMkqZHS3Lqz3xOmmVwUG4q2NfIl5qBV8
xwfLsjamrihQmHQGksIbFps0VEb7pvrNYJt0ayPO7reSzqiGJDAA3saP4cPKq3C4mo96XRBcswIk
jXILSPu7zIo5/wT88iK5HLp5gCY7edw6nuqtwWmjNYIsIVxyJqRTPwqysYc2pwd9ljsPPdUDKn+w
IYqE4Q80y7kWa4gbReJk8Ci6ogDc7szmkOZrN3YNhrbNd9Umi51EcNJCHGu0RUWDBtpv+cRQU8Yw
p4fkIyDsvOOsTVIxc8dTJa4E+/AYpIQLFIJYjKWLmffI1ev7IJytsM27TFZI2hOdaEsSv8j9uKs2
DS3vdo0oRUBehqgKFUNHTzyQCUN6jZHvKZdctFi25s5DaooAF0blZCOnSn7r3R4ox98TnUAG1Xat
RPoQXshHv00s1nTIOn4Oq6rTeWiYgsPbB+yL20VDlxK6l3uNc1Rsn0HAl+CDlEGGxY0UmGv//zLY
9DqxMskMW6mD459Gvl0CCyK9W7UbnYZ/VdmZWmKhYQuvctGOReZnTDneIYBRiE/Kjv5BwdP2woNR
wGOWrfPRjCqdW/OqbWvrqeU3650jx+0ycyhYQXipkV/BxQ+k4cQCgAro4vvkEzevsHiqLm8v42EB
QZP3/eC0+vkvhpqBwZWfH11MP71jNpj96moWELMWCMo9cExEjvTTjKxqs5eU82wFq6OpQZMoVrCO
CUqhX3bjUFV3wKXphWlcFk+Fo2CVN2+4SMcAYwLTS21A4S/nISAv671kLzTGAAlUjnJq8tCiUWs0
w7ApL7DdP25T8EoS782Q937rPK280YiAAHvmsG2OOFGoMEeNxnOshpllStqOgE4eDfe+OdJf0wOP
Q9axV++sYNYdfya08Z5oVduKQvDI6XWZ6Df9MWo3ofR+cyLFY5ifYgG+lfQ2Fu5U4+FS030zAME2
S82Gn+nURV9k0Em9ZERvuduGkAF/kNNSoLMtVl7feTA+XlZc4shMFtGz1IfzsQEkxi4TY1oThCGd
dh4Ie1i2gQYSoxINpInNiBofsrdLo21qLsdZT1aPJHcCUpDjSZz2EtQ5bHoq+D4GZ7NuPSnioTUW
mOtXaOG0gZTtLIODGRpUEHIjAPwlSY+/LH6FiK7/1XcvHvi+3APOAyLSR2Wl7AcqVNdXGbfHfn23
gc3pyms6dEa2y6AvwN4XLSKycHsLNW4RPmzqElQGs7djnu0tnrcGsg+ID7SmL3+3/0lO59ytYVD/
pB+z8iY4h5E8vDZvYjHZeiindnZ+rcen1NglEb4tijvKy6jqpQDVptJGWgjLA3B7F3X5Ib3faOuo
dp0b+mh7kT+w+0LF4MMHwLoaZybfg6TtNcBCId5k0cGmcBYep522YyzMfnYcbjx2AhSYfkh0Ixrn
4/Uf1++6H125zK3EbkWGbsNb0ThGJFChMd9W23cZOGU9pN5tWxu+SX2GgyO9F46R4oGemOWlcsNh
tzCZzHS3TcSG1w43bL6Y7YlLGbrQhDpcMwVnMfQJR84x97jWx9jic4knJMHTe/rkukm7EQqf0pM9
P41nwc9fyRPRwJzNls1o8R70XP40XG3Hb9DNrScZrHQkAYLHPgJa/JxYOkklwgZ/4ws0Cke7yGvV
GdwhiXqaHV6I+Xe9RWYLvajoGsbI5lEin4fWNCl4xr/BbB9e2TQUkvDQj10WZ91UAzxfKd6wzMLv
70Ri8glGXnb1NqZChfuAHNM+l3hXgDUTCyL+eMHBFXFHaSdQSDTu9GcgQw9+OIa9WPbnBKNVfbc9
laoctj5IOQscdljd/vdytsmDaSVjjlqBqmpp7fgKpa61F0CK8Su5Vl5FU3Ik+TIHhDbtFHAnqI73
Yax1gr5XpVcj3T95Tl93PSBBD1+tOpZsyjA/Nmyi8F8as67JlZwvCsuf7CmgPdXUq7X9zuymB126
oAW3Mrga7K+MzkVedPI46lOXc+9UOWoxCrvDeSER88oUAyuyM7B6y9pchNlzcC0XR0Rm2FAZ3JOg
/CL8SKuUjbJ+rQvQNqjU9hMOsuHs4jfnCDMJm0XzxMv986LZLFqKKpXR4EntxlC6fs7NeYpzwU6/
Ziu1Q7punV0nxgBaGxC2XwfsinFE5UhcvtUxn5dtk/L7SLIqdPbuY+zjaYzIaS0mbFXOdZzoDL7U
UEkxXofqzi8uL5yPYcUeMeot7c4K3YWKAJqsgCAcc1AxrZYcgoNQbR0VB92xBPpFYQFAbrisryya
Sd+ZhiClEI8ecquhT/zc+fIrWeSZvJEQetGLDureh+zLwLYfKPFN5oe+SNgVDSDqbuByie7hHMls
paNSlMGFigCeOuleR+g2EAfCtyAM81XBOHQysmFLfu/Lgp0vOGOF33aqI3Fny2cRD70cCfTFGBYY
7sILsSkGzz+RRTizOdeEanknFH6q4wl/Sdb1grdbgvc2zHKnQFcEBMqxIYpWS8YJf9vgxF14Bvkh
L/WBbS8jUb9pcFKJ7FroVZjWoETiRLThDR442kiKMq90VJOi/yZfZzXGIT5cUiiAYPi8aY7zSL8+
L8iomGp867t+RnB6X/q+M+pbooDnPgpZ3MgMme34mJMIxlTQZUAKRG1/ZrpQLYsPAznDoLLnXVwN
xKqPuUtQRFAQyOLKW1TkkHzXfe+GQynOk87gu86e3/ZRSGTDs5K9ua7AW6OA/70Kyy0Al1kZbpik
UvQHFd18l3jgo2ZNESECO9mS65P39hiEbBxQy1FETbf4DLM/yTK4SGQajEKLM4iOB/FQJZm/hrX3
5cT+P3eMjNOnrGLg6FOCh2ffucNrHwNFs7LNE6rIyznjPK6qQdl21mN05E1qo3nwkjGEjbqQW8tw
rxkatuAMuRUi4V+0d9e0ZrnLcEltDc+kiU8RTbQ/C8GvIZdTbf+Ht2iAdZeHa6k0vx8SpresKFdf
0fh1AqlDkvJYlpHB/gM3IszOboU2Zq1dLgDarLVdDLiwciKSPV3ISllZPD3tmExbZVWUuu/dzxY8
HxA65a3uvfpMwo7S1O03xRwrBVNgHGmA7ZS09Rw3Dgz9vIFL+9CLCaTd+/1RONb21AlP30osWcik
VROBIdnrU2YgGnUbc6Hv0ahGefWOBi99FOqqj3uVzoxBirTYbbqe2uSlC/mF5wwAKto/6ILr6AzK
s0qypLtH/Hq6P7NIjsH31gxahWVkfCpkxSRRvm0WkMhmbh4XC6sK661Sadrd0lbzV2HBs92Pw6Wj
d6N+U4+FXZQx4TDwq9rGluZH/hKMmkXt5HXTabNeC1PRhpEI6/Vl4bMFAyX0YxC8OJY62ycTecCG
Em0bXZK5pqsjNwuTd44Ut6imBGQoKCjDaxeeWq5C67rSob6XiFI2fOJ8dCcRf/ppbZlP37tM9XNG
0/teTozY66VAWYNFAqTQqReglpsw8vfh6TF+ep18syQp1TVXTUCiWfxsQp/dTQ6FNW01fMTcQzqW
TJNPUNfNoYkJB5wmkleBhkz+jytyXFMrQ4vGZ8PZRnzqmKU3cX87OvlTuVCOKPGou3910tydI0li
ZlJazUIOuK4XxCq6DtUkFOqEfmekllx3HBXnzmaeHW1uKdmOCYyb/P0pYSdWw/OV6+dYHQ62ANmc
/F2/Tu2k/zQWt5tKam9QqZaIf+CvFIJf+FsM9rC3zUncbgsOf9F5MCgG2Oup5zxSwvaxzZqcD9FE
ox0Po9Fd+hngHILEjyYAsyHZGMffU4KC+zfBlNUBEcSGCY/U32G9B2kqciEzk61d0copF4b9Gp5Z
poOstXUINj7F/dm2ayJAVue9qQ92g9ghvZWxYIwxCbQB/Uc9PQS0qWoWNcnwkhZ9Idv1w07LMx3e
uh6JRcoCzcVcFHQDLKL1IKTKFuDSYevIZ5J1RjkGr52TmQS+X2SgMaZ2FhA0ZT25rqe5mmMJzByw
rOI/nyWg0XUj2816vlplJrvm+kib8tZiiaC83uCaVMfW+Ca6o/zsufXSYPrGRwwgiFq58tZXfzyq
lAK1aQ5Ejagwlhzj2XKt2VToCBlNTYeQc2dvYY6/xQIAC5CYPX7Pefpl3aQ/z0vBmmkAuN3qaQpe
as/qx+Q4IqyCQC4wSR5v4D5k/MsoXnfc5NNFnWa24pMX4JJHOfPUdI3fFk8suX3ecgX/52Q0bLaW
LYpjgqeueac5qqT7hVFGA9vlm7FazLVgN+ZYUSFjCnO/vVJC3VzyNvexp7jfzCHbWu/nDy4sikYS
dp2yWOh3WCLROSv7GrHTB6TcnTMWJs9AbVlv9aeQMz75d9r5YAojNdn3zAw9NagKE5hpRx1ekbrq
qS93WRa2K03rMFR16UWFksvBoGOS27BIowr8UebyHgt53jFFXmqEdfsQKo+x3jlBHqAPte1HzUYx
0/jEq0KGOyAaNy6pgq4x+0GCSTalTlYaMmVGiD1SjnFVUSGcem/F5ADSEFLKxqFVkx+K/codTz+w
mpQcMBlfTMSwGBKI00GWVH4ehj+8g1F5tRnBeqxOgQNWgbATVD+NMEaEle2mkph6mSP7n9hfokUw
fN6MEde/A/gJJtX+0rogcQfnmmNqbUBpxfjjKb5o7cNS6Vg3hGSNQJdvizvgG9i/zEXwdpI/soP6
5tcgkSni28bUKpdYeaUa0SkAxlwAA5oRTVz048B9fZPMUEjlyCzm9aNFrKY5/f598YXUjkcHBrew
Nua/v8jNZlAr+unaAcoxXAcC5q0DWYJIzfPfsv9Us9b/MRte4HNuKEIJ10kRk3QzdWKZPxfMuUpa
hP/a8IW0+hgsJolhDQGA5xksxRBfegS9n3MJde2k6WcRdtKY+cZREIeY6KcP+Hs5mfOACsaW1YGE
I18sqM9ZyMOSN4XKGUBCSDD7c31YEIeQy4qA/kuhD/bNOuniNfuN18KWGFoOhGLprmPxwWjLRBIS
8kThSGFQcVxBN8OQGj8OcU3n0XJQfsokb9ObNjNHskdEzY46P7RrvriwUsAh91OHZqE37dkKRVaa
rOXGEFrgWc58OZEt2ZixdlGt59gNuJTuPXX7JGoy/G3clAjAHwdvJocpyLTSAkbz07pfnez4cDVa
SJElvej8lboc//oT6mbn11YKmVH7ziexxYemlCV3hWCTisw8VVBD2Tu7j2/tUNrZ9eDTAs3LWJVg
xsHknwgr8kMgsD1qfZxUVKdVUgkUr2DyITGWKT0NZyRU0ie50XYD+M5vSW617ZnaU2bYTJmz+r1z
5HSOn/6+ZI74RctexOYp/BFaHZju99HzRwbFrXRLiS6kPfQzR1vjcbROFenbq8hCo2h9385sQCjK
GVnGObjvf/qDg7EbbSD6mjjle8sLZNdSzth7HmmNtKA4hEC75iQw5ynYs/9C0dXLWUymdWcVQiQd
NrnjMbFtLJdMLQjmWDoYOca3wAzkmSXr1moOqCq/+WcudGhOeJt1Nht6JDdedf66iM/nLCvQysPb
VUXqnnZWJf96LkFtWUY7SD25tYSaD8mZL2RnI5wKC01f/KIm3MzBd6pTHDqKaygitVHQBR6d8sRV
qZWqRsGtJbgcIEauqmG2DGrlhDzOqAxk5+cx9Fll+lB2yfG7jRTSsqRoW3H1sqGexb6EpJXN44xa
W8VpScZPySjp7v44r/FKA0ONdhfT8XAnh+Nzz/F0lfklIhSuXV+wBEV6pl2bnHXQFWL9V0yQN2AB
SPuKX0P9skdyLElGPvK17NPpC1WP1gCkNVrP5dRkWPpgYe1lEF1t5no4ALBC8kXkU2rlwmn63AOl
+daAShoS90yaQyFyMPd13v38Gbdck6dR12ZlxWyokBS8b5EO+D6TalpLKoKTDLR2o9gcy0fHQE+j
JSwJ9EWg73ScTNfxkFL4/63C34DhhU0ojEHOUPwPBcQh1J3oNTrUnTmfI7Ur1DlYVSkr/WA9dP+c
2SzZIyex2wF+A0508lw+K/SdPvCOukzpEV3DNg4HRb6lLVSdsiFG9jXEpgkUdJlGoiVjxBB8VQ1A
o/un0/1wdvGvq2bQ+pyO505tL3KOTrfFWzqVUfuLzngIhcx65z/NT2wcx3nxpyrIKcpT+Tmpn5BG
LQbiSlhptucaqDP7rda8Hl06sdC0ctiuHUH/q8bZAhVeDRLEpqP1UzSD07IobXGsPy9dWjxbrulT
7JVWsE/KkEIRPFg3HzX/RVHw1Kbcb9z/y6RZ87McyoJBX72Lqmu2WQVCF/ToWtBzkEEGUKSXWoMm
ofENjNEiLTZNzXaW6+Jsk4eL+i14Wx7Wg0MuNLSa6JQrCWzzHu6MmSGZesYzcJauRVFyLtr7+j0S
iPGPkRauYmoxvofXG3DDyrVt8FQtvPiPSF+ajOl844nkd6DWEtyVLeUHzdyf9uFUDsbM94fqVXG0
dwqs7nT9867hLnir4F03KpaLI3cVSpZYJ2wWJSB7aFzBGmjynV6gEGSGLzYCMqlPgd2luNh3k367
yLp9QIQETXkvr0HAjSATk0TF0SqfMuK55rDIiBahiI9rqj6LMVvDQfcY2fzONkthaXb/ow+O2eFB
QiPokXGwsBYV3kHGbjTZA5yL2gNFsFVyJUNxKCln4qBPtszBqjxuJDWHtGRbyFSZ8dooaV70Xcm4
xTYtf/yEw4MdEE/0rQNuJERcWLd/3qHoMP9FmywPF1CKPsk483x/nGiCHbPnTiNiNFLI9OWwYXqx
z7VyUqicFt6aNxglofV/5JaoxLRZnGQISQ23Txdcf045omCKFvbGG2Ljzf6YBhYfYPBpSkn3QyI4
dl4RHcB2GSgIJsoY0naw3Ahf228Ehkk5um6qi8gBnptCxTOPdibz8vA6wrzwomu1hLW1vJ85xcZ6
mW/01C97Z/EtQ9i4v+h0PnstbYAkOICD7bfuH1sd1XqETYj+SQk/28nTZMUUw5WwhYdxEUoxxqdZ
/qHp2kuWyUDziBS7udw/9pI3fnIOLynnWJMMtMJESLOeCkhXhTFPUDQWHueM8/Sai2rGeu4RrvKR
uDpbQxt7Y4sizZizLAigtbOXHqVlNbEtC9jY9i0F6tBLZ74Ha3x1RUgV4luJ8s+MS4cqOCA5DWDM
y7mz5cFZ7aytnNcoo9BMyVGVAK3PrmjZCF2szq24s22kiPir9GHvEC4AQ4trGDwobaJtxSbTgWB7
W9umFglwSW+oua3ekFpESP92KFWDZo4XvNVisikO5BBj1di1rbn3ukiKWfmFUxCKFBSbkkVIEJG7
Oj9yrSFMiawsDDFc+e7Q1U1cGt4s7TX0+DDaGZbZm/rqPEc9TAroZUtxUycDcQpx68i9UbHoaN8m
pynveamApdnY2DoSUC7lIrCjvAcwDQ0qu0q/Q3EC84aKW0uX1iSZvW2J9yc21IJvEm7d/rd6AY3g
hFUxR0+WhJxb47NZxgp9csLYl+kP0TnUJWZ9seuMcYd5fBqec21UywoK0q197poPbQGfBOoAONYf
p5KJNNn8IBTcjMijroiL05dx1P6h5A1BeuXPyDodeNLDmv4fTZai+TJVRJLzgbsn7BJujvyw57lV
DxKiW75ibj7E0X4Z1r6OHQtsm7mogF4W2d5+RhTodvCvSL3fFSxRgbbS3DpK0ruXLNXAyrAVQBEe
BFOxMzFuxjWoNZHYRNji+fpsmI0XLgXB2gyVzijPLDDyF3FBinSqV1wKbpksvdjAE1U56L7lVlYL
nVLdxqmvyP5o5DV83maUZ6Z4nRepiPqKH5QKvGM8br+wCxn5ByT5WXnE+RYIeyoCdUYs9u6elf1G
ao1Um57Ts567PbDUzJVW3CH9mwlqmLZETRsESxz/jrjhAP2sGSraNkj3oGxznt8mi9N43IblUCk2
9m8cnxt9JOV3EOKHD+XZsF2C0XSP+WgyZRF8+XWBjgdnxGPDSqlO3xlfRls2NPHjwGDw3LKKsQHz
X90yXKCGUZzsyZbiP57oLFfmxO2bRUhHhwI0b6M7gMgkWcUBng0bQTmo2+auK3t24RKMtUeKboa3
zNc5Eer/BO1F6RVwOMy8gr8g/CPJ/Xv3vmGdLkIeqFEmEbzbnTmQ+3vrZ6x2osWzi0a2I5aXiMAR
g1O+j130Hy+w7SL7cXYyihK9rgjy28eVynnL30fd4SJ6qQdClr/+zM1scN+jy9CqET+/xXwf2EuR
66qeKYnsWr38ZF7FJfJIb3t1aj7iwSXon87BZQSEsHjdamAnPHxXPH7dXkNzhSXKIcdWyJ6QWRek
P4ZqVtezPjTsAyLFAdXOaLNPuJl+5F5Lcu5JaTsem8n0tp4z+rkVKxHbWh0U9foPMa+IEesHdQUV
9YrTYu/UBlPi7JktoIOSvQhafxUH+5Geq2qXXp68L2QdNZU55wKFrRGx5F2o7teVuHiRFjJQ3VUf
lxUQ//ujj4GNw2qZtolPmJLvN9R4qs0hmhAIj7/igl0WBNL1F/4If8Qcy+pvvF2SgfnH1zRa0u0S
IwnX89iljtltVXw4yujrTGjRgKpnqCyCLL4wjd8N/RhGowOxVTrCZxBhhMzEywi4wrIQaL2J3SYe
+AX2r7ZP1766M4VQiSLax7GRlMkI573r4CVrfRolf3oPXyiXecjlT9m1+fHN/YM8YxOH+qu5OoVv
dD9nRSvnvHFNe0B76FzNtnv9AcpSMcAGw7OQqqlBCEju2O4Yekr+XFVX/GeAjn4Qroyr2Ip9o28O
0jHw3ZmDXSKSZ8Ec+MchaVleQfNEqYIvmnJtQhcCb/AAxQjON4tyfvRnKES1rbxQ8zPffL/pnrCC
X49xf/qp3qevpeydsRtBET4ZpPCLf9o2IjFCf3XPizCyGxbCe5CuASodxk6j9rsIoPVY0GI5gLBJ
s2AAtrl4MkyDB239FLOzw9sGpcY/FLf3mtrF40H+fqT4YXk5loBO7P1DbIkCsT62+QFjpb8Y8ijn
SwhfceuiffFa6D5sYGA760KjaW7QLieNH5ihvP8w+zt8Y9DPdQ+wR5AgWHU0NRgx7bNjSbUyYPIq
ribj6ex+DqmTmLVIlyfiLnQolcOPMC/nEZ9qnLGLO1/7k8oaJRPNKg5XTlQwrG9ihEEL8GbmhQyF
9mRsWFXFVuolrxr4Z3/3cHa9JhGkwRN/Y4724I+9gs8lcWLWXbwn8yhyuLl0YRHABxhol0IsYMei
KODvv1XS9jmhV6/ILP+Pkb5y9BqpZ4Y0NHamHUN8nvuhEz3tN5Tk5hk1DhzqCPVh4y46nB61pz09
s02JSeUaFYEGfIjL9EfllzSVrbmgOnzWzWZSewU4K4L2Snq9eGDfkGp5Eg74psGuDe0W5jgVkiy0
/DMyLKep1iytEKokcLEhfNidmMVZXwEbAisLQ0hkDRH2Pu5Tksmqsx67+fIP/a44nismXQgG8SBw
jsA2QzmG+4APJ6K46cZc1lO8hHT7muWzBq2dS8TsDuWy8jXUNNvXwG6pV5N383knMSgI9c/wM6Mf
UqBNuDIo+5UjdLutdLR+EKmH4JzEiGCOjLJsTo64gjbR2OMQ5tZaIF+BhXn5mBNzywJC13QtTHsv
jhcaFtW0CkKW+tYkfCOKPVJfL5ukbA/aSTeHZmzIk+i5AHNRyRRrm53O4PIHWzUJQ3Urqi4q2+II
UdYVHB7DYHsgi7KZvn5+s61YpTM/OD9kVwOgIZ9Obw4yck3dxHAosPClz1bRxLUCvucjfxJmA4ax
bc6Q5ulFuQHQkrjmunq/Dq18bZKB98oz5GrR2sMJtdFGlsySKO8ecF4qlzkSRt7IrRY+anBbCuVQ
CpEbdg6v2sU96ANf9MwflSwiUwbvXWbx1rCbIY9Q+0ncIdo4juSi8VRfpMWKwgY/htF0Sws+6ydh
qCdlt8EiObMMWj9PRgP2gbrP8GKz9p/QfNfV/5JnZ3jRju1QmXbLCEMIjFVl1GlAhDjlHUPF4FBF
1JhFglBz8AxBTdfDUMBYny9j+p4HhVYYHk1TMcZWiufPKLqb1ChYnMYfpY9bdx6Wdv6gt0OWDffj
Iel+8d7UxbQtmVyckJSgAiyWk7IMWOcU9PiCtMYTrWIFCWtNlJE3RHDPT8pmuLNfL562mvftQrRq
+x9ppl8zkK/aUANUs7ev00SqHCi6R8Fn8YKnyQtHT8M8ECYMXYnPI+84W47PwWGQD6bq3ZYjSAXs
EKOMkSVdGaTt4Z2maSwdA6ZMr6Pof0txGtIoJt1Aqxih/8zUfYKMwD16G2ExKREH/as4FQSwrKaH
F/nKqJrTiKUc9GRAk28bbV2RM0vlkBhY9e5cIlew9kaVz/kVzOtKPZY/7yrc3QRv3biRFPkS+/da
jqGSc1VVhzmlnqEIeq1LuYSLJIl86lkrm2uSRQJFxLCFYNVIx99IzsSnehvXNrVnCmhQPgLKCJJg
/vJ5zjRvC0pmgz5bfBTSnaF/7Gq4sqG8dfHC0bZE24j/zr0LEs5koLW7OGVfR/9Sm795fbr1vt+W
Lj4e/sMxGzes6mbsKXvqtZtnrb+Lvc5FfmZOw+kbsDVykMPuYURXmY98t36anjMnqDhvSL5Ym46X
GAB7hiompQXjBTfbUbYHGnGF//j0jGaf1zQsuPPtK52K/eVbS+xaa/weq4S20+XaMWzoqqNG4inV
dpfhslUCwY9BR9GhiLlYYry+G3zDUriUJCHaTOtvkt3BByn/CTd+h5ksVzRP6ZSjO/N29n9cyRNU
ftJJnWg7ccomqNl/yWx3twC1UHmHgq5KjSnzp0a9bGhgOFs2BKCf9cr5VDus0g54jQfS643skjPu
O+kK83KJsY6HQ8ORaIwjlO3Bmtp0G8KR/h4OwNFcaBAJ0Nf6k8Pc1qL7seMm5vjROmVmVETqtddK
cIZTA/I84XQblpZetTU6yfutajiNeluT26EsXS6u6EoGuDZqW6L/3USOPbwnmMMfgIi35JT35OwW
2gVAF0IE60X6orqiyIEJ3BxvcMsTihNh7JS04t4MJagXTqByvYr25KcoDSAsDSI7XnrFDNEQFvSg
1jg6/0N1x76QvELF6bj110+QKmlvbhXWsHVkmnW20SuSzky0K70jQdBCEtFFvN4XPSnWmxoVwG3o
Vt6g4LwBq9KpkyZIFB9AjxxNvXiqRt5QJFecn42N19pnJK1gRSDhrziXm7TdeMiz6iSRlu++8uIM
EshzMrQYkP8rnHe5gmRsQvQ5h1edPO/y9rEj+bbgK5chtjrEG4EVkv1xa1DcFCbsGnvfwAc30U3q
DdCT51nWQCTxZRVlhotc+xIT/uAtI51zqDXrV9xznULm2xZUsBG5VUXhb4GS3A7RCTUz1PV7G8vg
7ftptt8xEbr/bc7VkO3X963gmciJ/xR9eyaG6nA1o9UYyKxGMvPJuHxpb6wpOhd7dd1f4WedwEuF
zBCUeyPVKRecouhS9EWOtGhtmpFXXE0bd+DLAxhk3xyAPfKu6g+ooqnR/L1rfTQrRQFrLdzKOBKt
2MJZ8D2J7eXsHYjjymGXvaV1F5gOW5yni7QAOITD6tRtcclhc/ijS4+IQuTn20zqiQ2YDLeSfkZA
ADjQpl3k+zdXO1WYRQhRJtNCBS+TSZHO+SB1609bz/mlM+kxx4+5ssLvopNY7WLRWqEsWVmC+62r
coxOFzlw2p1U9tuk6fC4XrBraM8sledX2AEv8TjNUTNOa8zJ8zvmdbBiJ6ZthiUbXpzXA7EDVD1O
3mErvOf44aZWB05j5BwMu3ortNHbdle9e70z1trwV1jJlJ2tLxa2Dt2uUxYO3ph7BcsyOH/HOQVP
g9XJbbTZSxXJl9hCWDeV/mvbqVakxufwF4KrlDQC2nBFf04PRoPgvo0EqQn26fpR9IgqgxNCswji
rDReGVp43CjOz1tLSE9pSRZyKrI0qVUz/ePFJjcyv3pqn+3URT2orCI+IvI6IvdUGP8R22h6w5u8
3MYc2eie8UgAz8iH78f6NSEgKPnNEkpnvk5UK8KWJUhCVrHctrvoKzTGt50iD6VsVgveuZf/zTEv
KxPPeEBoMI//zP5GZMoXnVBguyNs5CNIKkC13WIJ7DVuNGWvyXkEeNtGo15S15syGR7yLdEWFN9C
Tc19cN+L7SuheRKx4nZnZUrEXuyOYsV+iwT9Y6FUq7fY21rLD7+Jvyvqa/uiBk5mybPco5rgwA2C
7KNpoWVItRSj3uNpzKjmjRfPtuqz8Ddfd6ssMvxzfATUNLcmEur0v3dqW1G6td+LpuWUb9Z36QZ/
5Lt7VRu75yU/4nPld9ITtlZ1h3HN1cWTTuI8Dd8M/MM4DUMcDcSyKkupGn/aQHbjp52ExJ2o7Mpi
CxFe1XivXQlkdbu4zrFu5HI+YHxdgG1dXNQhb1X4hRZAY5p2IMZYr0oproX7hXPCMBkRgFVOBLQY
CKDMZAP/qY6bYtZR9FVfCWIiJ2lzGYoJRJJeih3qk4Q2qsmIoVNsNyNJN/obEHaRzf0bRk6MP8e0
7PrJe2U3IoO+zb6EewnunyxMbUBdvUD01ljjA33gFHDJh1AX1DmFdWNzPG7IfboxGdgkuBnHjjDZ
hGROJysrLE6kqrf6WqamsnCNukS2B98qA/wZ0gXzxvrXlBmtpg7vC0G/lHvN9s3T6b3Gwmwspi+7
MXtlE0K+FsyOAJANKcA2+JyvU3wE1fYgShkQ5mn3xhtPskkP7MeioWicDcRlgYhE+0tLEAZJ53xc
KOiYFMCPp53Zy9czr3DJHtTng7VcoovA7YPdmUfdc7+PTchmTPBeZEYcwTU1rr2KbVBEgbogBQSv
9h6RNB3j5EXWJbdKxDz15VjWY+x3g2MYrH628/TMi3zlXfa/ZOUlEKRRsvRmFYT0muwQG8hrJqrV
SaDXwfRnBLTCzwIyxkFHIYGPe3C/w5GL63HFrzUkJe7sTQzlPpuco2WIDRi8mpqj25Oor+33msAm
Sgn7WdFKAmJjf+1mPPAFQQdgqijI9M9ksY9IsTfXoteYTbIlPtkFL5bG4OWXNVG3+uzQLvkG+1d9
qzNp/G/Urd+WNoFEO8smJJ0OtscJTezPvKthk06CsxLUALFXJqLZdLnFPJ1ODYi8afui30cBRl0x
/DeQdoWVmfgx45bXO3tY2ibSsXCI7qaiIJQ4H+bplEMNoeMM8/Oq7rJf//LsDCQYP49VDDFEwx6u
tu8XapXmWyCf+4LMAAqRtKGgNuAaq8SaP0cG23SSRFIKLPpQ+jWFX/r8qi1g2Nlax35dZ5ZlYUiy
R+3bA3ABUo142Odikexa+dzc+H/xucV76lcd0D4qQAeVCEFhfC0NDgrbsW6EbRDrG0zxjGetPwzz
UdoPI7sRazlWVpFwuAOqA15hJLaNYnTNRiKHp63LIP/cUH9jBCURdsxgPbTat0sD+rwL3lDvhIDm
OgjPAV1+D930MdphIeo+VFdqlrWqJRLX1Ej6CbMxy7ElXrHfMHBy7/X5IP0bZxnE2D7ALBmqyous
wEYInulr0b1y6RCqki8e8eV446D2l9HexsejbpMUCyhwVuEMYur/DT5562th3vcuZq0Ds7gQS0k7
al/5FSkiw8qdM0NzyZdrCj8QkeNudQTwxZsfz8ai5+EvarW4FwejtLi6q4GsXTfhWZnQh9OAXUvC
+vCOX9TgEE9kuuxBBe4FE74N4WgyY59eknaomrieY3a25QpYaK082mbxcuSVpRkS4HPbVlTgRFue
Ael3UP9Xt/98hvqL7REKTT60CJPhFdxMNv1XtrBr/JqJXuAwiF9NFmi3/Hsv7FwdPGsmem5/0na+
mFarSI4qM2g9Syp8Hq556eKQNuJ5v2UDq6OnrG55GedP3IW92WkctVVdzHca1X7ZLqwDzjeUHovh
EwHj5afHUawsutibJS3pQ8BYIZSPwlONrDnZC49bJCVLX83rW/ArCI9FrwBzCp9blDzBYqp5wW0x
wQPuiWrRVlKgs/CG81WxNIYTUINTcB53y9z7O40128fEDVaRZYFyuKcbkIFgZLR956Ihq9IsCgM+
NvSNtw0Ju3h6TCm8SYvj66QfDprXi+mk7dcc68SSMPy1LRGWx/e+JgJDXDqLBu9b/V+Mjb68YxF6
mCLIwjiasBwrJfR6XMOeVrfBE/dyR3zDumHpHsV7xXZWQUUVL+VzZffeKCqUgco5kS2Uxkbh/Dzm
OMPZjxWhkQSjhGalCMCMre2RyJTkbwSxPXI9SAz0V/ANU9Z6iF5R2FkjQe3fyedaOSqLSME5TocR
BgqqfTRZ82ZKzmMqzzCbrWIgfcnhAK1FMB17gVWFwq6uGEurVZthtkz5kid7NHbsUEmhbP5JqAyD
bt6nzqSLG1O7VULRwkc+DKH1GADroMKyFIc96z/fK3gAzVik0PyS6a8WuMLjytxTz355Jp/M0Jul
WiF1xDqBh3wNDrIuU6m4IkAWnduSKUXz9g5XkXBrKdFQRQ1fCc1MWYeCbtFUxTPgR/uS0n+HiKaw
qvR2X1KOGPmWf+klzOTtUvRJKkFDpLCk8HhinxlGNN1aaGiBDF+anCV3TCUw6oDzEjetdUq/JiFa
+Epca6eWfySrx41VDxa9FnF3gzSLquiUE5V/v53qbGvhIFJiVxJFmawwC3fMaEyC05/IhmWrP/o7
Nu9x2gUyM9ipuTttCUETb0x3o8xZHhNWTi7frUX8FVHq2O0UT8hWqVF02DKUTSyZYciZm6vXDs3G
ByEmBaT/o+enz5hhNAsM6bkz2WSI8b8jMe/rpWlbwvCgKYzw8dTLdn73VSS8RNrwJAGrBUQjmeHi
iLwYVI7wvsRDezV8/XVIe4gSggPeqhMNunOwrIMuzF5B3cQNoUeonnKSPefTI34Bx1acL7/92aFJ
8aYQewOFDL6UBvp3GcmDZ/xN5o1hsiQbjDWNHO0PEp1tW7hmFe/2j9GLgjGhd4+1OW9daTbreMx/
Tkf7MC8rwm0fT9DnHuCTHmorSq5vwVVxRao2QCFUFlSbqkHOcSeHPyZVk8FhFxAo9J9KmbheRexC
1aWyjrAjh8GaKNRXIxbF7dxJ5FA1OEhXBYeI3xTPMYH9UpQVDKMmoeJ4yIqbqyMCOflPeXgoYobx
Y7F6A/zXRCHR+7Xa4WIa/SBUD4hooQiIEln4QOxbA0mkRw8L43LRXhcuKGqru15Zy4ObP+q0jZ8P
xcL/tFeMeq8CqrBo3L0GsK4wGagI32TAiEGCNoh+hJKtiIRXEQEp2/QaIwYSFjhm1uLFvhMMZvvN
p5U6dhP3Yl0rZsgdqH2qjkN9Q3Qa5io6Zri2S8+hSm5AUuCl9mhNGOxVVQZEmOfBRZByLQ/Cj5VB
BYa9mlQWbnMPwfIgR+FS5syJ1YumjsT6t7sf41eZ+enM1iJzVJW9w+zg5c4Qy8HzFo35bg5t+iE0
ZUpfEKZb94qbjyE/GuaZoW+QZdlopWoltdIXggNxEyUyNM8lhNf+1RH3uJ4+0XuslyCCjetaGSRq
1oaarlCouxuDaEEuVeg8Jr7lplzAMuLhelO1ssXma0NjcXzqPFrMInFMUPyjBraw91VRH2LYQ5eC
Qlg1hWYVkkHxfu7ZXl0K2/X+ZfyqtO+Sx7HN7t7dRvk7VVpW40zRDvVzROUNteVmts92/OFeqtkn
AnXfnv0Emfdn5b98jWysPqLuavcKS3R/RfXU9ssTwXi5E5cJCFOzvJxmOceFMauJOEMWIClIrPrL
moQRp3Qp9jxZPNW1xIRo5it7fdVp7hyBzyT5aO5MCz6sls7NqIEy75MoemoqfoqRjuTMe44wHRuY
8HcnbbqKdR5XgSCIvjpWtD8HY2XV4CNVpc/YYrY72kfhOP0yPRURLAVk25olURjgHWMLXgxLGDow
Ui4sU+KWVxAaxjHFiPMlm33+8PMrpRVmWfJFPyMj20spq+t4p24CaZkJ3BjvufyqhhZ5WJcKFBX3
wlprAwULW+OB+u7DB3QHqSbpuQRMzES72FoitEvjPwK16T64GsgOmZrPnR0CDvqhL8MF/TxYN80O
a7CHnx4zsVlDBVlsGslK4VPgdD0+7bs1KHerJ+ZoaA3NIaHJ3KE4tJIMBRr0BJ/IMgf8g05wfYSA
Ue6O0Xsw/Rixi4JlYkEVcCEntvUT9l+pCf0aN/njQVaVem+fK8SqEM49xpL+jQXjjCt3a5FLykWr
Qs0pszeguqiouPlGbV8kip8YcCKUSPZNOGpEZNnLgLhzybmnywKcCYKyohEVnmh73T8FfArsL596
DSGDokAz4bIN2vpbS0lPCxvpnW7PBYj0x2ZvIqM5oq8uGZW8Zue72/Ys41UXOKNXbE9+eRh2TJRs
OJn/VrxOFOH2jqoeXpnyOAl6sNmrX7nKiRcz0vHIU7ANzuzyhZ6Nwj+Vj4nLOtqliPMEeGe58foo
myoplKKhYvPE3hUZcMd/8ZJQxUgc31zJx9jDs+F6l2HJju87ZJbwtQi6PefzWEKjoM2bvDVU6ff2
56RVDPAyu+BHutlmsx1rg3XJ+sIEMAFnyPXFKKI4VqkA/pHcm8sdRXz/ifLYRjM8YjqoQSqWp2eL
y3xVK69ggIdenZX1pQumN0NxTzNJPul+kvnF0assWZO/SN6a2/GYL+6QaWZqMI3Z9mJx/A0Rmszp
E5+dLdoUVY0hwtIzBwp7xC7EaqyiFgEXZuCEn+zXU4nBkcKDORob5G7/JlqSTvnEFHyUeOCRH4wb
Mkz/mlIcuctYHUPsz3Ixcn53Z1cDCHf2ZBCvzeQjUFlw7pTSh+P5Tklden2jJhaNceRliB9GldjH
GhaR9L8OmNe6gEioER2Pil0PxCyclcRuQqvixsGrKUJmoCWQRKdenfxWrG4B97tLbY86yfLZ4c96
Klc/8H18YdgoiiXAhlqvE6Rd5hZF+IMe+Jjgd41cUeb6FToXqI6gAjCzaQlHYiRXbe22mwcKaWnw
ZWRP0RGqk0L35X5WFouvc5NYkG+kfC/lNAoev0X07hCZpxVnNZhzeOTPAOucpe22l86Ccn1tLRpE
txShVdVVTMLYdzqUMyHRmA5N4YySFG8IO5Nea+PoyCKhrAgwsPzHlmxVocs4TB8huPLecf1UMeXV
Mfwrd8cy9099C7SOlFI6iIe09YpXrwT78HrtXN7UHFtd9xjICusMqIzGpUp7133/FBfC4lZkyt+O
3HnmMyvK6sOM17xom9cXl/BgT2KpzHyop7w1kRjMf8uUtTZaLBy+kvI9rmtpYjJRHSsw42SHsUBq
BtrK52f1XVEvN6OP8UAoEi2EP50Fo87GbM9w5pxNByOPf/Uh5JBsv2icuQluqqvzCW1zkHHN6E6G
wJo98PqLfWWEFt3K2lx9CEmzBdsRw3Sfq0nae8HiuXA01oi8C23r+x+e0nmHHfxHV/bqaWEs50hH
cQLJzvvhM1cItvablFjYWrejF6toNV+j88IAXOcx8jk22dzpsMtah4Is2mhCEa11S7maIorXIife
5dfFiqV1ibSZIBRbwSdAmMIMJJVHjfzKdZJrlHY5+T3jDRrsG7yxDk9arUaiMz99DyiLr8M5Kw04
tZeIuLApCJdw4djFLGCBOdMEn9SvhyWbspjDOKO9JdSusGSMsl+NS9qwp1Vgo46fMyKGdtSlQBHe
DTENMdBxqppB8bF5TctANEBshl2WSWqreHYIAhGwjHKEsHil0/whSS/ybOoLe2gaWNz+wUbLdCRH
X0mo4QsmaDymNJo1Pe5NSp47HC2ikOkVjkMDyE3gQikA9Iaqv3CR5nkooNHkLU13kPp0vFCqO9MP
zaYNzfmjdVOvK64K7f2+ZfqTsbHq3VapK2WPmQnWav/MVU97Z7XtB6XjnvQu5VUm99rbCRxMf0Iv
Y114QDbDmZLfW5Z7b5mkjAogH2lIevmTVClpObHwNPbC0LtN3mmBrfGqyNysKtKC6flU/MMRjGyz
DxZGS1/Nj221oPFOUuNSBdR3Z4nkvlYUdLEQ4nVQkUoUae3/UnIHxi9HsCSkbm/QWoc86A6YCYon
hTe3SkuTiovqKfJ5Vx//ShYnLd1pV9ELp3Ay75GeLTCKWzSS7TVn6Lg5zDX/xDi8XMTCmyd0mLrY
XJrrus0O6m16bdzG8V8z/oi4DazGde077Zc17+Xlrq+UnvZJTK7d/zQP7GZ2iZBkQVdzCcVKkyvz
oKeugcy88LoERT2Q21QHkbL7ukuWjQegIHR6QA1LeU/CNmPfgZho7Wt3y2GTvvu/s4oSTjHjoXJU
EquhMuU8E2ahEa489uveHJAIlKrV8ftJwvP4KAKyzbG85oafLQRe7go4MgLUd4xSQJtKdkhm/9Gr
Cn1Idi8iYf0foEzAvo8LU1jH/MtYh7dbFcBcbru35jZ2J14UHUdvHp8AYF5NkxHWGeFMCKhVOSHk
IEmLpVkqQ0kjLKJAv7o04HvblMCRtXVdcNbxKZALWgeMuMoLsyMqgRRHhPlRifHVI/bgxb8yOUnJ
sX1rsHgJlT0FQgfWEZfOeI+y8UOfibYNSbSi4rmg1KLJHvZ+X5sHiacxTGMdPCUBogxBguk/CsbM
e7k7ZmUNdaWKJl63XuIVgIkFGshmWxHw3WFzA7Ff1jHtdOJ9QL7FWUu+f41PjobO3M/WeCE6zNlX
+DEo6GFj2zovm3EtMoMIYl/IEdRXo+DWYI92JlQuaIerxksho1qtXTQ54MRx9cti1TN9Ro6Efh8N
Ckow8oYZmkHrRVaOszub1FmnPjNTPY5Rcz5T75zyAPGJBiu38YnEZEXbjaqb/lE7BZKJIuzAmtc9
xjX9l/dH6TYsVOD92mk5i4F7ocZvWcncvQZsaAPgjvDOuEAVcm3NkbXWlX/7hKpJJVzihXMxU4XT
nsZ9i7GcErUPGWv6lfjIf9y/9sfybov362q0WX6T1xA/4paH5RI8FfVxDaW+PGoivwL0Hg5RR1fl
3cKYZUMtRT7Meqi5TepXFFLdKqrvHszyZJVtqWGur7aYeqBU2r+G0QCPbxHlmPK97DKlrWXmH1XM
DjsiFuPaQM5oIwfU5N9q9vTjIjs7EKPbI+R3WM9JkE8WGZB7qKnNyOnqKdItqG3VGmIfZK6unadZ
d+7aS+xv4ZV6BvP5A8xInBq5eJ+ZELmY5wg4U66j9J7WUvyjx1i8zyAtmo30rNaUS6rcKmjluGdd
5/V2Gef7181LLGGUd7crNuZxfjlS31a+O2vnq+g4RK5ud34vS+xKWycXczBlpGb+PjN8pCC2gAU3
aiSjGpespiLKJ+Waeur3LyEgAccahtoRlkt/SPNRgDsNwcV39W8oQDGGfy79jYIS7SlUstIJRacq
VawR/Xt1ascYiPWUhewuI4hfym2l1pDCWVLq/Q1AhMVJ6OFuzJXFGyM+rtqFaDcqnMNsj0zdM9aK
cUKXdAplkW2eNdY/V5uRJYy1iQrC+OOQoNRVgJcnFro6Hb1k4cg6GU11guwdoXRadGWL+5+v/QG/
AiI1n9pfXX1MnBSgD0ZPwhhBgTXXzBMhbn3pxMIrSZ1VQObRbMeuEuDaMxNMB+4Nt7X5cX6x+1FK
HS0VJeOtHFOxMoXCXJImQlOj8R+tdoIeiu/4lnNmaVN5naq6Fm1bTm7qBnC3k+qtzpQ+EcdCdWvW
Khj1EKjy3FXF8tPWQSLUMcNa/Bs0kC7wNlNOZAH2WbAMWCmicMJhEmjSAyY7nW0jm5BA/0rv5ll9
kNGA4e8ymps71guPwtcu+LyJRmDC8oXju0TreaR8MZxb6RXBApmkfIrQ6Dcg1vKMbunOnTpbAvvK
aeYVilxMW44oFFzba0296iRAhxCfWfAXxjhhgis62XZIykPdrY05/yns/+YYHOma3VgpcDFlCLxA
htrVcNA3liXaV4OrG8m8iwRX6jpWUKNADP6bs9BQUERCRR7FTd1rjeTDRGqsBvvEffyX044JQASf
K70J9z4pX1eGjKGh5ygEVR7kr8RiFEn8PqfZVxDFryp1MYN4a9Q0x6Y8RBiIjnRDFt6e6W7aCy+s
JFffCvZinPdUFhpGOyRZcSF5UQi4gxKZB++7WLEQboK1v7v/JCGmcbN3yD6N+QeZhq5sSU+TlCxu
tBx2kOZwGmneUQ4JERNUdHs8l6aARQbpfKxjh35mYvbENB9sk6z+kbAeeMbARWaCpxdirPZ2GyY0
4DEspeX1Gc9+xrVJrH5L8uZXapLN4MwEkrSoiLm+DeVGZZImoGkXBXEDsA/5oz3FaijusC4EhcpO
7bykk5J2hcp1lKLxht7Q7iLe9i2nwDrS860t/JzigqhXuQ/hI5IAdnVEElBeVKYg37vYJgBxip05
gtiFuMvs2nKYJH42vu4s4FE8sbgWNPwRrq1cZnWc3jStvftdTHIp8bfVE6Ld/dSQdLf0AA5z0CcT
agsXsYuu0dfVMbLcBEp2DKj4ZOCa3Y4e4ST7R9Z2/gOM7nUjjYFrtok1kSA7aaccDLi/ph4LG3rH
igwkL3FQNkuTImFsdlolrZwzq/8k8+W5jgU9vYTFR6WT3MeG7yNyLXKToRWqIn51e7vsAlG2uqla
sNKBl4p3OREV3r/tCaPWVKo8/XqwTQKtJHUJN9jvHqOHN7WFbMkwF1J3oC6F4gDIPd558AvoX1sd
SO+JgISYb22gRw3nhHmC4+TiHB2RK9vfoKYzk9EAFbYPY4Kz8daVxsRGSzdMsCAe6rJ3O1GL5n6J
WRi3MA3DyF6W4GLlFJ5xGjv1emlxaWvutYFsY7xQgln5fzjtTLcbn/f5EIgceRbnCwj4T1wMsZ/q
ceXuVPvJ8F50iRt1884YJG1pGmdJEpDF6TkXXlgsx9refQBHbG/zZ7cA+pld2Ye+tNGFz804JyHy
2qzqee4xgWiGJUhoSWhxVf9Sfg72FLMT8seBrU6Gu2Be8Bl4/Jwu+3nSQqRQFjcc4P2a1tr1CULJ
rKQz9GhCjiO0SwUXMd+m2ESd+TKLEGjU0yTqEkVfKEOgHV72qcJNvznge+dQxQbtPyxjzwdPX4np
qBKWQzxJP121HK/JmZuY86njWQ3wuvwQ983Vg0foOktQQkhS3X0k95pzIeTlheDJKBWAQZJPgMN2
YlzqLsKAhAwPa705ZYy6ME8T0fR9xKsUVr/RxLrpAICZf7Judo4EO+BsbZFSx3TLfPo88T4WC6CE
lD9RP7EzaNijWIRFx923UUZQAKfpxm/baRCMRc4cHdEboz3t1dBhfvPCCXeE77P7xnQuH6N1ry3N
YbC03GUHqnEgfwzTaDYRBkgzLdhHXRVf0txBOBZ4Pp65PpBSmefS08lMMtKUc909OyZIj1Qdk14Z
GVSWBUgQa9YyBYmNQHmUwlpNI0uVLXk2y0+t7uo9J6XhlnOro0x+DeOYu4KH33zF+NLms0JM9Ob+
zSqOLwf+89MJ7y8/uQgED52m2R0Yz7SZs+DVpHDFmQtFKFS+3y5sGces0LonYtYEX2y1EoyLX/cG
p9v/JnISbcRbMEsbK8uX/agaXpRCMkMZRxE+dsRWDq/1eOTAEYg850pLmt8LaDhfYwfQz1j4QHKl
1S+XF8eigz2JuI3gwKhs4RoQqrjN7SDXOtJh/iJdyB4WkxWs5Delys3NUnJbIT9gOqnGFpjlCytR
YSJ+7bzbJB+6WiXi9gwq0//bOjLTAXcii/8I5oWtY/9BYnVBef/qhGEus0IITSW1NUBcGJIR16YB
aB2j2gxLTW9YqYHqDz+BR3dupHxawOpaIZhKEIq9rHhLueKo/HNIvVjE5hQvWJKX6lzfZyoHMrib
Fi3qUOshAOvBz10oF8Gf9fcYxL4b5yODgicKYOiELFZRlzrSSjk6G/gTHWaNqFCf2WikE946ORE4
KhxRh1eWF09pEx6h2AME44e1Rn5eJAjrnT5OkHuaychbUqbBb7dUMERoh+5stzmU+2OzMXcDHQQn
qJi89crzuStkgbOM9wFVYzTuN5tiOASmsAnkHdNMdQZlItUnFwcL/8ZVj+qYzrczgVYoKWlfI0Hq
rXj89uVTudd5ydkpSU7jo8SsF55OEYTBTRW+eEbmshi3fJSjFot2yNsEMbK3ZcY6eyOnijDQizzG
jX/qZUqucryVmSuEkWyoFaC1dnFlbRls+UQg2ZGjQBNwnfUWw2Y2g8Gnqcuy+MszW1PacRmZRUBB
j9yDIalSMM0o/SNY9g1RIozJwgxhFEsSR1mPBpU0qhzymux/KlM/RwwC1/o5bZ7uR4NGiAsSSkSZ
QVCJs3QaoN936lYsKtIRGAXF4WGahX53kuw5KJGJ6w4/ORKVlubjxWkEf9TECSWU5xeIWeyvkQ11
OAU7VVvqa86Bewv9DOjAma1LzljfGWyuyr+0OHAScFc1+MawMEcUvWDUudU1bPNHm3O8UWudrKQd
C5PFV2KnL1Exg5VxsIwuLjcgSs+OW6wQxKAf4xWpjLFq9/rYRT2XrWRuAGMvt4aQbpsErI9+FEMT
KKrA2ifBsw7ihjw17Av33hmq8aCd47RjTkoYCRJtr1LShE/2vFRFEeTct65x7XgTE2AwEG4bJfpp
rueA6AAA9gz7A3oZ4PX9FkCAzT6M1Zz3G4GIKMs6VmaGKhxGthyAyLTNm57pYt/+MYcf85HB4Qi2
s1xhhW/v1xF6k+2Hy3HAWfyX2KAUbfPT+CNbeZujU9Sl1SFlw/DStVgNlRIblU7ib3FAb+9wnG+j
UzKd/JH+DPFNdlbbximYJNqDyZ5eJcu/X0ErWm42Su74+6OTCRNapdp7+8imXCIC/RQHUurRa2w1
1eAHOfdejctpkfTdfbGT5WDKqJvmWiIa8/BndiloDdTreQJvVg2s9CUyFXQPRrdfZccsfpdJsgzr
wbrEsBV7RDzrdZQbYqgpsK/3snqRGkg5iTq+GZhb9ethE56ytjAupg/ykDElxDhSGBvP13Zyglaz
hudSwQvB2I8phItS2xuA7uPVKqSV02L1bh0+XCmOnFtjLIyq1p/RyQHGPe2LREZTeIkPFQeVGBYX
gW4nUAl3hoITprMLzadoAuMQUEEl9x14GRrGowoTep7e8RdHDUu6aDyePrftFN6UZdtBNyVuOeGx
SuzIi7yBKcpGe1GysWdd/d190F9h91zzLSr4tgVkpPuyvbJ3V/vqTCy1O9XULSjzDaWcnCijdHu8
It3HSVmZxea4XxYW2asSTZNClPAE7tAw2GAu2sNNOTS7IA+Gx4h4INTRHmGCRAqCm7CRtTBW/TjX
u6ZYC4pLQyAzmHB5XM4AxvmcM2920aw4dGX/O6f21L0Ny8ywakixi+HwmGbxnutOA7NgSaQ//T3q
gSbPtIriC7koiOLj2r1v6MjjzwwL6VWceZTzDqd0pJ2nrSOaUZGCrykJro69DZ/4rMzbYM3wa5BY
MDpJd8I+7k8pA6zbe6xjc6ezLfS7mk27Jo2L9VnMtybpukp8x79f8Q/+Rwo1h5Ob7ERu85pVt+RL
ietjf4SDvS6KECF92np8BVnjhtc9IrTh72VQgADQzfBm9uCpbrkQOXF6J75Ld0K5bGpvdoi/fLBp
zlxdKqx8sSlyDKG/P9DzgKS4jcVCMlDS2kFCDPrsbkCl7Tt8oN3gWYo62Zt3sc7auSX3Mu4ySJ7F
d4Tj/0lOdFSBqiCCAadEWSOluOGEC13R+RWPCTDEiCy2lDw7H29Wnb2ywcMa4jYjU6SGSkkAHbWq
DQCIxGrdFK3kP2nbpuZliHjXXsY8Wx0PJDiP1UzTDvYTDKGPrHtYKEFK6FowuKER/SKqtpIw1sJ9
S2c4QzBf3wLz5Ub2DWE0li5es4Cnblot19SU0sCgKK9P4Kf32ZKqCReFQDqAhuiVWQ14RKGb9fYO
/QHIPlFdABs1BFHI4c4C/grU+q4UZJ3ZtY6CG9PfRgSauA+o4PAs+ouAGg/EwvP1rQMMWq0RfDuU
Tpo1O9tYwcNyB3cHHxDrAyNpxbHza84dB3C5j5eVuS2FMOkxGYVLOCTsIY033QHsX9774iJrwfAt
oOaooVmBy/zPvmPxU8OPz3ZxIcsPlBUhZ8TvJ3mb4bUhRcADspUE53trOTvC0gjTQdyZwihmxmZx
nshFlr6vNxp5kMVRdhpPMDJU1Ac4rDaAFydV9/oEblfRAAa4iBaEGcSnmBoxw/ijYX3R9C0WFx+b
RiurpZZel2XOLdiCtvnGFMfZSE9Zommdbfl0J2PfEL93KkxlHVbsIQ+rS6vl4SJDxF4os6PAheE3
AwILYDfbrOAWbbvvqf1VZROyue5FFKRiJE6p/7VITSwpio7viNdDkpdy8QJt1DlL5irO/p/0wGP9
VH2mYZwRtY9ASMgF4n1wKmYfcx1qrpLEeHIety2J/KjrmsDa3IqcXeV1dn1USY9opKzU+LaSD2bJ
oE2bJmCXaYa0rXLBqv+4z/vPpjG70u3fm9bHzW/+jQcl4U5V75j7ut/tw+m4vzNuvdCctLH77Dlc
cDTGyrdYYtCryRo5aj35jWs/g2QyD+3P36F4Q9T83K6B863sgTPBEc0SSpTw4cZmMDaoWf5fGfab
BycqGmM+wwK7BN31vSX5kKYhib8PPVy/oa5SVufAzJanTKpAmr7W3fFFbGNGgxFOSEg9jGOV9v1U
KinqsrOlJ9epSjZqc4mW1hscl9qVk2a8HjPfE/YGaZpwSqZEuYY9Qi/V+wDsZfOuPwViDqVhi9Hs
GtSsaCzdjDevN1Nzw5MGeRZccx5TR4dSOtVDUkJ3aLxyqX4LtlbK327RXlfYSt1lRsD4uZU+kelP
OvO4Tfw0bWs/rM0XNhu+tXdm0/L362osC+Hf+ypwMkU7KObCBSkK3BRQ7XWKosNvQZ9bZLsoD/lt
PHbhmjIIr8wnf/kO2WQrV/90+amMS1y70Tl2ZphENtjTqT/TdBUDIPydxVGDBfKggbw26aRLYzM3
RjpGisQgmnv3cRrM/WG3djPd5h86b/7Km2AhwllDxuT1b7UnM8Sbsd24RvO4li2wgS5cPQi7l6AU
fc7jrKlyz0xD8dTwYnHHZbjjWtk4+9+IeVggHNoVL2twAFlL/MoY9flYQnj5VXVxyMxy5QUoKsw0
tTvrcpXLs0/pTAdPxkWBeP9g6SkrrYG5jbO/7TeghIjHmZnMR5yogs+8FbdbWrstJAAs8DDxnYqm
anlnJfBj4PfXtxBRcLq7PU6ZGtBmVZIz70FH8RBl9G2KW7pRrWIaLiIuk3/rtGLKXgE5aPtxGu/R
DJk4JnqIx3pXh7e2oC69eCrRYD3MWlqqI3ubqo9PuF+bSFy4tVAnD/8r4XwApq06jImyLi3BPuou
TJQONROrbPxW5FhxUOJBE+Cdw9u72P/E4HYxhZPG7M0vSg2yF1u7vlQjLLVC9tlGo+NzvJYJINLE
bc3xzj8oPUMmDxubQXvEXZbNdUueb1vK5VAc9H59ACypTjwpfWI+PMJ8Iiux3UhpI7BNuFcoyKiU
sIVd+7Wj/pT6e7+aE20CKxl924vfJrpxdxm6cPnJ0M0GCtitllIGlH9snD0PzuTvbzuNBGujiUfA
EDgS05nf3X8Hrd9XH+YS+Pfnw2O0lIXQxeQ471xp1EO70MxcA8rEbAKjB4M7C90a21iedYHJX+av
xGTg0qBlerakkUnLNfowzNv1dno9MJK2K4rUnrdXZ2EvEuSWLmL3QnsbsfKAy6gEQlbX0oxual4v
izlKIzkRL7hzPrvQ2u+sVpZJuaKLK7vo5751vypFuQc2GjVPXDWsjJf6ti7FzGZzkW6cpEbAXpRz
eRu09e7QqFzozD3PwL+SXURdmeT3JYF/gMWYwPg/MXtVtHrjWM53zAIR6+9uPq9pbHWIe3QfKu5i
G1UhKACO9SWwfQnLpaYGiE0WKutwyFyO3TkeGf93t8E7/r1cTc8bIUNpXEZ9i2aDk83Zs+bCtG75
rwIfB4g9BaRFuomKPhPKTTRu3hneBTuFA+R+8NMs9Wle71r0XZHfyT1Pc7HqSSm1jpxX9uOY3+79
WM44Mfe5fodU7tOZBZBGXa9bbNCG3q7gP5+GJiHPj6VGR70fEO75R89rUFqovGAEJIMyNFgssyJx
8aorcYyFCBRvoiVUU2+xpaIjQZVgklw6ApigHPxY635GGKKfzCFxopWAlOZOlAm5lQOvHjLDUkLB
2N/FP6VLGSt+U+JZ0DjxunE5uDkxtTO1z+JLK/dJwBUMN37gtowfdg1rG0XFFKBlSklsj//JcntI
zcQ5SNlgjVkCHNuqaaz+HUH/66XR9BtAiW4yJGWAFFs/N3GMH8AOK3IzdQuTONlkh8jO4mwHJTk1
pcQkoyQgLGyeQzTrBD8eilexIKSrO5unKc/rJWIeju4Qn+WOKYu3UUz8kDtVpDPlZZs77MuQvv7q
ytKdk1X+iJd1CH2id8FkO1JlHjoo8KxlU2W8VbhB8CFUp0O4+kCNAdpf7Cy0OWuDo6gg2Trx3nzK
C2X7vnJ3zqruXXbnwo6VrT9ju1MYzff5yMHuY5qHzV9LzNxQFN4nPklly3d9B8MXsLC9ztKTCfXl
E3WOfQdnoG1WGe2iumIieA2Kt4wQvPIuXzAJhVX0rNObyWfKguki/kYZR/AsbJOiRMeaCTDx3CaR
6aG3wiDnl9VyHC+tipEzcQTlydclZiCFUAt9Pi7lgtWKnHy3ykgs7iJRzFTDA579fW5PjssNS6N7
d3lbajBzsoAbof4s6qnN/J5FycNya/sjdvlXlz64fV4vTc7e4SatE+2/xYLwpSbcq/3eFt/R+uGg
6pwnp8kRWhUxIFnGtBt6dv6qKbZ/pdV4SJ704QVDrcRYHeUXRk6IZvl4/KapV3oVOKiol1HIYXET
JkvHBlA84JFtm4AY22+jR3ZPlKqnFXthriwOqPnKvBWtwQdT4SNaZrLR5ZBXaNnw/7uTkMZskTQg
nPM5vQ1g/tfJpCzevHnyeB/kZZfsys3NpEGopKy062QAOQDyyihxp5KR/O8pv64BSLkoFgajTvv+
8w9XryPVLV/FJe1e08XX7rtz+nMjXVcTCLd9u1JLc0k/LCsSWgbICMGcjdLQffKVmm8Y7tbFAEiq
MTDigUDJ39wVfvxiO+MwB1zGRQ96JW9aIn09VYZVXR5bgf4URerVhpXLv9x4nZsDcSF5M6f/EFEu
SkaXmnSnWeFeJkSCJ3E3whGy8b6LrG00zpu7pv+abjcdRWgpGuKXWb82mr1ZkwtoxT9JKlyZ3Ffm
cRFAMafbcQlA11NvWIjqAolSsnMCfLTLjo3oSTM1ekKvRr8aWZyUsJByN6QFrz0zOIwUxkviO7EZ
l8wlxxfbCIqqQ3o+Wqm9ctcH/XQTUSNqTRG1k5u1R1fivKablepNVN8I9Af2r8PNx+OUmxQ8muS/
2CLMM8GMjntIXsQBkJoeRcFjJJxJ46orMGQ0BuawXJ1lSKD1gMDs/AIBGsoQ+j0CaF+pj0f2LU/Q
1Yf1vh8Xv+shR45RqdI1gu6WKbVz5eEZkf2bBgv4+5RTxXiW2sTz+0CB5V5u8+59cO1RgTjJMG/A
DLszT/e+7DdYd/7y3txvAQuGRG10MBCbvRqN0+G5A9RD0T9raBcPYMhscpxRDM0dbOTnPOA2LbUH
UPI3CoKGvfUvrlxkkmtUCxN4wYxxIMhquPVH7prFXt8sMeKXK0hkufjpZqIJgfWdkyCjF1Ju6hlj
MGaEv4cNg7VATB3NmkT51DbbbhUMvZAivB4+mwGpgYcdG+c5sH+lB8B7KjHphuP+mL/lNnUptpH1
IAENhegrjXAy/J/NDqtF7IlzNkCwE9OW47PIbzvBvHkC3qNWVx79j99QYAi8kL78iyFFYoBrFzMo
b6PGOBEZwyZW/iDyD1XkDLa6sErDnZE0zY11C4B1vOXxp40MAAqoKANtxs0dPwjWh54sfckQE4FD
axew0sgNrSCkiiaESdFQ1WFo6IEWl3HtjuS4oBdXGExYuwEWO8vyo1jwsMmuxqaaQ0xAUFK+2Bf7
Gw4rwaFT/z+sx7qAHqs4lVS1ed/BDwYVmj7ySXtEkgMPU4RhrZWoTqaR6NklzfDqWxTfhJ+qMpLv
goAw1sxH5UQm5tQof3cxJ16sgbpIBZl82SueZbj5mxPXSZNXGhe6BYeSgzKev0mI+FlTK5mg/PFn
S/RkI7Um6G1zCIaTbwW9N9L5+dFU0h0VlwXTHAUBSoISr8ATFY1JTnIn5U6ymQdy9/fkWN5e+CMz
87Unqd4wfFtV4Dqi2EQ0LvzhBJF1fEWoH/mQuoys00iN0aW/D1j1tJLz3R2uolZDqspdFbNHbW6y
huX4DQ8VW0Ak6r9jrTIcWKRzzYyln/xoadSZcXVmUhL/K3gOWZHHrI+DPJjBDL6ZzY3aETNdTspi
TkK3lqwB7Ew9tQalNJKHB1MXGP4mZoKIRzDeGOVJypWEwMBSquOXENFh5XBbqGVeU1UTMKFfg6c9
l0D1CZOCJu2OR37ruIshoiAfuYYQpEvLLKnsQuXfEany+Qe90tJBzXdxzmIPvW8p86yT1yrnWlto
o9TuA3qIo4WBQzHcuXUTLS++Qtq/t/ZY3wAnODTG9ZcG2UcOyiEaUBjxWfAEwFALRCX9xmmp3QwV
rS4Y9kXnmSbKFvDy/8Q3Tr6NPNEn30X3GEeizIAzMicDnm50SngurLdC9Tb8LggIv7SILvANTCXK
dNyDt1dTLp247VnJyoFzZv1KbXJU+yPScK5JXD+7CPWoSa6oeEjHAR0/XxdxUXKnTIDDIV1vq0vy
s1daIojPEGphF8+29KUM+AxWqBRFhSrcwnX5kqye+SVIVNRVRxOQ5n5kKN6L9cZ0YKNZbBFtEUBq
rLAFz32El5FDJE31zbKSnqw+Cax0YLBgFSybzXc8HkunOmKjPMzKurCaWerA+e8uTKANmzxZRCrP
33rMTss99R+LBxgkYyKCfSxg63D5BAT/UVZl4KIvpcRzoUtArx04sm4Tk8m8zlJSl5Y5QniUPbDS
Jd7sgwCGhAkU0duKsYwzI4asCEtb7+cdWPdT/akeKlPrCBv5L+FPThsCM+mHQw9BziTXclnwgp+1
H/MNWE9Na/FNVG4tkUucOrtsPb71fV4a+TiAVFGxCLR4S+jaGhFeNaUzfBBuL3a1Zq6znhz4fExG
XFbkFUR2LzQqG8VC1mF+fASjODiXPaMs3bWQ08Qzj3yj+QgcJRUa59UKgFdsgdQrVaxqCjFxeJiO
top9+jcj9/gLeGn9dGORJsJoWOYx+AdX7wumbKyRzhnT+5f9C/FyW80w7KjRNfo4jTuSG3xsSsoe
Eplz+yFkQH18wFIucA0G1+vlxW/VWabJfgEfow19UxCur+9cXcplAHla7mkopnr02UJGBfSUyMXu
zpBz850WQ4Bxos4QwpuFMKoX8T9JZp0uz4oGruFsLMjzTOA/mYDAo/b+FnWUeJBF8Skvc+OYVWSN
ieCESXqrO4lmWm0tqJR7H2E6oAiygtGQBI/H62diMsIEpykFKrS9bBxYDAkH0s6YbMm2IIH4OtqK
blILgCVwv95ZjSRp1bTaIiAt3knnk229szqYhH/xUsTJd1G2nKrQllM6DcBUEXEfgNyhtgUOVxqW
JOVEXtDIBL9jVC2y/Mvw3a9qyMwrzp0pRqHLVZWwPBRH+k8X38TkZ2WXDTltofsThRPAhmfR6S5h
ZfCBxrnyYvBpShpoNRWKmOm6wlff8w9jjqNWay+t7Dg2CWIvsOenECRJiO4zJZFDZqFmc8JOjsau
dH5VmfJ9fZ7Qcy8Fn1Yct56PBe3MP2WpbjX3j/eGsYjflRlI0M5gFlD5Raha1vcO1B26FgZpotEg
3x9S0qbcpo0REU79G0Txg/0uk0r+vH51O/YeZPUusM5xPb3vMZjmlDTTiBmIR4zrhFOOPveT40li
hzzvTx2aXqxb6iwQK+cApQQ/N30I7wKTAq/o/JizRxfF7+p9EoYOQCoobNax11ZUc2dDNmqJDvBS
oftCpZ8GF0bHywzmgYEQHIotDzBcd/Y7WfZy0RD8594E/STLWgmK1ex3WWWJSvBQkP/ye+70iXXz
lgUHD/MJUiV//FucZo5aXmGEzGV/jqSH7pHASXdQ89Ryzk3t1yz/NjYQi9QAKMini04pvwDqskSz
2neB0gVpxzqToNot6oeVKkWjrUJvSS+EayoFSKCaROO8MHLXRmQ99eyw/q1S/TQFrZX3SoWZM6g9
9kIJjl/lNWlJq8JruSsf4aF2OIPVKBNshulI2szkBy/I2W7OGHzn/X7TL7f6oAJZ7DAtTPaxQJ2O
hbNBJHGxMzqSj37f/vN+0qgvpUGC0Th4g3wuQ19N/8GNbXHmEHLl5vzL7SmWHwrLaaONoIcxYcqT
iwzBW3cQiq4ox/vH6DSR/A625wBW/PXM0OxkShXKJJbLpE73QbmhFFGDDHlc43NBr3UWTObXiLZO
vOeSD0M6ioc7pOeqAF25Ki1BO5NYSiQrBWlrUfGmCSYjic9pHPt7+Ykyq1YOKCGOpeeQOSTA69wk
r95bxll9oqLsYpPKt2jq2NMl6YbBfZ1JnJdFQPF5i8EIjzPYM1xvKa4rIq6AGeuCcoyBFzuuptYG
FVAOwL3iHAipAyK1OzEOoPD7A4dXqcIEf5ijjPKGO8TF+v3xF2+ues4w40tJa9Uuo+IPhgqCNJjR
sgi/wdSsc+47J2JolAhsI7PvKiweX26t1jc6DQpy5aQIDVSbmam9UUV55lmKr/QNtIx53bEVZv3/
qpF2noe1ZBMREeShKnuTFtXrnwBLLH9bhwvSZJ6iCq1ddi2u7b6cgJY2AcrfaIBLY/Fawy7TRx+x
gNUTNbnQ+VrCFuUr++u8bwTD9ug6g3KsJkRO2lt2UgqJPWtVpqZkC0epGjaqL0FU21YmwlMebACd
wZPan4D+wTvVdjZxOcsKgkCgT/s07vzvwhzSQumAlK5ZAmP/YIGcshzBzyr6IHPYwp3VI7/HtID0
A5yFTqepxNXEvXEn9++5r2Gq//mhFE1+zi6x76vGH1qv0OlUOXjXD4YDvm7mh4vl5MSNAhWWwP/w
1XtUK4MH19Q1F4LLrzhj8HLjpqdzGt5xc966apaIvyCJT5TyR7P0A/F16CYizi2cQmp81Zw0whpU
t4lMta8b7F94NVArPw6Dr8YZEfNg8yhVlaZwMfMMNP0Iw05ejdjUcbH9n2DTycHPtkGxQ6NqqB4L
3G3avIvcNKGJq/B7+0DG4Yi0sZMB8EP/2Dll9MSLyiDnRU0iH4QTDirdAAbwcHTFzeDNuGwbgSob
FkmqNeauOMEqJ8SteX0cvCyN7hGRB524CopGH9YMGbCDneqa1OS3Z40/HMgQLKsGc0JfsGn8BEsC
3b8qEQBSp1qSXPLa860z+7Oj8cX4Sd4oLXZlrrm2XUkkFwHtNYTVuMX/D70FoVEZ14u6SPIH0G9K
hAeMSILXeqeuxrGzBT3uDVnvWunBuDc7T3vaOSoMjD4dHn/JFSLSIXM0TBL8oCZV+ILSraIfv0aw
byjOFMyUhPzXmQC94MqgH3PDLbTTY4/yOPSmaXoPfkI6lGHPSrcmBGHQUv5vHSTGf/xm3aYaVzkP
448pOklwVGfZWDGQgIOI7PlZ5plUb6yyg82cWsn+J8yCRCclyCZJ9hgs0X2MxlTPG51BxfxjP0gN
tU3xWDUqZZnf5uEZ1nyI3YZlOV2mvhUN7OG/cQqOeEomvMVIqqf8Gbv9F9ENKgXpTxdGskC/kLch
HXttvp693+WOjcprxBKaWd7SYCqXbbPMllVaiD1meBPu4P8FB9IQdN3O9fa6er9610Iu1khOvHOO
lNFfwolyysnYwLLTkXFiNA7PD/kzh7+/D057yI+Wqba0Se9MVOdaLX43v2XZpmjcQO+4eytIBRKc
7/lg/aMaQgNQ1gEtgBUHI8QU9DXbCKjdb69dviGx27ajRC0GuhG1FBQCNtVbAgy4ACQStLKYYrbK
QSSell3F8de0Ck5iPe2qYuH3gMOfARoViXUtBAro+k21tcVtXuFe9rBdrVhWeOm7gZg2Y8nilcWO
tIPFlhMtYdz0UkAFN7Hbd9JAYvS0oN6Jv7pq4q3VRBFPBfTmVGCtHLbVg6eZR6o+at302b68cMoA
oRvGQJsMV53pz0h4Ct4daxs56LjUlCJLVeQT9+bwxZF0VuJr9cwYRvYiJWIc+ZuoAxBxOU5j2bFb
rbGJO/H4rnEwpmU6RL2L37SiCGzYlnmMY0HNBLLMfq80eODAl5W+n0fDYfa0MLneoNAvT+G8Qa4r
+0WeFiqPJd7KXxFsc/T8RNIYxYgxuHP8+rEG3RUp9GZdwUZu8WqNn5Pf8Po6ZTYfplUBPGMPZ5G6
akRhBcyJzgk3PMNXms7IHa4hEvw1bDT9Dfh3XUVGbeJM7OnJCjyIrsI7Ey5tsiGFvRt85hWrNPAp
ZDAPoVcQB3TDGF30SGPtOZ4Xwe9UDFom6Zmm9r3v5d3w/tVopw+ifXXa3ygcDel+bNunBYx/aHW5
YuHsY1D/cWBEtTB0YFGUsOGvhOXWkaBCOktmlYT6qUrNl4GZeksRpTk5LyhAmL8O6xY38Ow8yidV
K5Qg5Npd6mZgfQonXzb5DS8LzjrLsw7CJeNdn4ZgkeEOaqZ+4fPHyM9qOeU4vYxRYwxKJm2xANz7
xis7Ipc39iUfjKcT3Qihhrcz7Xy/lb/re3RLiqUu0+hCVcRqy/DrMMWikdz4IulpF+9Eo0htzO+v
d9ds50VZ7WlxgsDfzWYdqI1ImEPTjyZK3Pm9ZsMO9YH7AkzsJP0ZKdExl2ZwboM3ciKt1+ZDbpfp
B8jVkYvTCF5Yl6orCVCrhWvA21zjWbcK4J/Mryfyv30DxAlbmMGbyhtQ2ha1Hdlgb+64BGvg2Rnc
fUFROfadSrjYnPmwZE60kVbuX8ix7JVnq+vCq2XS6s/ufBBp/gLxfHwe8G8lRuORw+is63BXvcxe
u+3IEvZhmxQ83v8cJBvlTnvwM2dE4Ovz7uxMJBne8WFPDlFtqBPuX7mkJWXZePsGZFR44Y02Qt9p
YmgIifuMzYquMw+HA9o/nRRrp9wJnHQcdRSMUXnUVBwwu3lXj+9pooLrV69yVWkf5b03U/slbEgx
mjpGTugbqX5lndAbNGD5h5BwufsNredpIvVkKJBt8O+dxK9KphzwmziLhxDjSeyi1GwzPJSWvh9M
I8ES+Xs4VmHH8/oLDEQ484xtVbVp6AF9h9E8LkQqa9xHOKFeMJT6tvY0u1o0uiEDuyH8+3oix8uU
xjHQBxvm8XPhLfkmpXwzhhjZQWJ8azJF4YLBCbYEGNcg4XSxA3lvp1Vv2zHbdtulw2P87wYWPrWo
nH6RFrh52Ym6tIrAUsEYixNhLqj+7195VVX2jRb1rV5181oe3ApR7CvVk8XbtpwlApqg3Vq2ZLc+
7UkOU9XPtDlB5YNNC0B2/F8G/aHU4+F01j/wVfNGrXwUR7CcBL8pt4+sksSrX+6hWmYOu3iVimF4
HFtY83vQV8GPSHG0wVM900lePq+4qGaQzmFMyw+oZy0Nz4UTGY0lRRLxie+MSh9ltw2fKKLBmLnU
jXIfS/vvJ05yZJkEGfvrPzBf2Pkizl3h53VOcuZJjvdfaiYdXewXc9y+EYyOtXysGUBrbaZmH7V9
pltLIHNpFpRyPpcE8YkFl0nAGmr4gCRqL9evGoY/rnPYdoAcRaVCyI31NgsegRfQhPYeKimsC7FR
O7qH0f0+KPlxgSe8xzFkRD8Z/ENGL3omHiSoWbK0j1UbWS5WOxNjI+muADMMwcQh9nYBvymIbQHL
VQ6X0150/h6cyYRbyDC1yHJ8ult0u+kct6wpEloCVMG8wuD6+JJyS32mweUMaNaVDMhp+4gGd2aw
etPjrknR+XCqMz97sDPHDIXlRvHYKMKm7rGrXzWYU9ZPyENdxDbMjRklS8932UIkCgxMISQdIICT
KG5C1mSW7BVBdV/vfTjzeASsSTjWLSWxUObW4K15jbNWDzDysJRaMMgxjlYVWDwFkQKwZVW5dbKR
pK73c7y1qDRsuu7BidD/1xHjcKwPWh1JepiGw8FDEbqwbcQdWGRMDSqz5DF8gTQnEAgZOhQY+TFD
Bc1twSIMx48iFBJgFoRpff9jgHTs2HJdraMY/KDwYbvGkvmIx/A85XA/vXNaQvT+dLIOW6koFxB5
v/iaSG7QFLZt6H389HEokj+Xxm3CEOGCPTC9j2Ms6q26PH8bJC+OiyeWIbBYS4AAIxKM9xFan0S8
wa3xVueTSyWE37GgNxBePr9bjZkHOA5IkBkcL2k0+1njDnrby5Vv0Hs7W1/TdiyyOp4oT/18GIgX
KSgv62ZJJqaza1JI2ay5oT1aFbXLL/aQ8yxrzv6Uk9cVK2+UUAjPMP2Sy4FS/2wdyAd7poTdSVlh
OASH8At0M2lZToekmJLcBMZeZb1etYq6SSOp6V4d4SfuzMqOtkFDOsSrgHv3Ao5C+McVNO5Tf3Tn
KpnnA+CYhe+PKaWF1szi8uIq95luZnUu+ph8XQFSre/jhRR4lc3W2zBGQ0pKfCWHaJ1KUdx/nTpM
Pu46WDatiRwV0ZVrxsFCnKJED28P3+XXWqJjuwH1kklAbHjrMt8LnqXboJOuaGq90CO0WtS3EFEM
zCLjOObfC7R/s5oHEy+3+A0PRFPec/NgTFUmFFd2BC24kwUuVFRerNs0BCJGIbhe69bYhkbrGtdD
1HiLYT+yFryEhFkCuFVnxfjhxSVNf+GH3BjZnynoiILkaKyPwCNG2NJ5B9mW5lSRwMgwqQMtQAHV
hx9hEvmEqkmSDNy0UJ9AjfgP5ppew0zaMeArrntLWi7gfgT9mK3kJFWiVNNwBWDtMsc83lTBPZQs
LsCoiRvcvYx/0XLuskSFdzjBxkTvCN7/1XCTZnneLqjymrWbaEw4USZoX6VaGJfdqobQbfHdIpnw
tcNmqsflb/Gggv3wjun+CWQBwiyA4BtH9LR8xeeqvr40mj13mBd06D6S/fcS2NSTd1Ni3bLnYXYJ
pzRuT9TC9YEbEwVqYnw/07uAHpMN0mXCzpLd5OKdUpnwFo81TdLtcg1r6oTWnUdqzeawO6FisF0H
I6sFCaMDn3q8V6EZfK6+ck9XqUizEB1y4DtsDNr3vXczbHq8mSFJ8/9XrCuaH2LfiCyG6kC/QhRU
DOIry/Xq3X8ieF/aa+95sInNuRtVySrm6ggNNrRSrMStwc4R1WE0HV1PmmNFrkxw+JiHHq0/k34W
aeo8PDMM9C4CyO/AAoH0aNOLwFIfSVRWmg3QtRZJ80wdlLOd2jMpnQi0TiYhpFUa0EXL0puNEezu
dCXj7K3wyDlTFbKlq1TbBFPF75qcQ07eisi6YFR/8htaHSWHYwhC1Jbypsl/9Sara/j4LbYxknxY
wHTym5xFpscO73BLOUX43RjRnPBHBDLwAEFUkAGiSKg58izH1kVYo0aKhFXVg6Do+bzk2bgFhjih
wvtyfKqEk6ffUo4wqjJQ74k1DmjpAkcDTviiQ6fIMdtXlJJQHAI5rwJHVi8zIYNFoszgHqrQDjJB
jtI01ZUhHA6DxxFvgp3DqFx+4TfbayHgYZIVZw39E6C+yaHHmv5JXhXjLM1bc4GuzCoJJ5o3Zhp6
G5OfqaL8I3Bw93LX9JBnRb/47T4FiMvZGgy8PTd5c1EkaVBxRyNsw68Bm9BfiyZIehvO3Ec90coZ
GUlFc1/owDlgBLhdgIn6WAC+vjnI1Oa9AioG+ZX5Mpu81wjWg7GtxZR+VvJ1Ki0QWXA7pgyyuKsV
HjhjJgHoeJL0iUKDvIq2AnE80rqqL1tw/Zuv5flhLY2oLRX0v2CqSNB4QSnX9usfZDcFv9GG7e2q
d5xexzTDfTeSoAf5r8nD8IJMIX0pk7nqo1i/NSv8K5qVgkU4AO5Bi3PhSDUvLpQPzLkZYz+hymjJ
T5LpZWSTzOdO7+XC9hLQe44oBKGYD8DyihXPu69UmhTx8tRCDg9/rTM/9BDXN2oVmGpA9+e+S0r2
dn3Yoc5J/iX8nhkeZwdjmlv6RuNSwXvkRyIs4I0S1zDo3jh6l4RHtmuqh9r6h/ipv3FXjmy+dRDD
s24sCwie1n5zXFKqP7FZBXqHgS6Ncz4AXoeZjO8k0bMBtL59hNIgSW6GoDojqRB+D9iR0dRRHTRS
qOlePlaHnz0gQd7f6b2ESO3aWFAAKMfgyvlf7j8EG+MKSpxnriRA4X8Z7jkbhmAep8W5z1D9HRsz
0c1JTXRz/thQAUWrti9adx1gaM4UNjceB1EuIc8yXQaPcAyK4kazLMx4gEk6vqudM8+jVmDWEA4E
KAc9bNnf/HyDTp/n2DnlHbzCRzoH1AQfHixTw3nXfFTa6B7o3gXScnXfZyxFBiEYjJTOsAHgPMnz
mvC2JbBQ2z5fuU8fxTSe1+bERElpHxg+tDIWkVJPL3uLVqg+36Wycz2DXef+fDk/1fX81mymNntX
5OgvikIe+6TQ+NfGWFAN/gFgddk39yxX0+1tQYRXo26hqMwqhvAverBgoL0Fp5GatgaH25GPPAeS
vxGMVJY1vQUXvSGzCFGdKaUjtwEwIk1gilXLfVAv6wO1FCy3D2+L8P3ZInZRy7jtJ3wtOvTnLjRw
S7uTzZ5leIaSgcSSvpHOMzQwh0N9XxKzEtFZqwat1fmlL8NZTrsRHnuKk6hVVLR4qvHdjAPmXXfD
psBD12FKVTgNYTuOlOHyOrT9ziObdjJjNDkcYhiIglOv+kSARJLu4mBMhs4b0oUgzUvvocCRhtLR
mVOpT9GHeuxwVB3tPbEjZLukbRCCggzE0JtLclEwSrWqnPaoNdFw8XxGdGLweEZSpNGFVw1KpidM
SZFGarmIU52Bg6jPtN4Qa3D8dzupQI3pHiTtOozRUR7C4bM3oxFjk8z3ks6tV8UFDvPr4qOSRDYq
Zw85brs9DdUILvIfZ96HxqoySTvKjlUR09FrXs97gc02pXdQuQFpi6zKZ2QKJXswoHEW39AAzSib
mx9M55j3FpS2watb2rpVA1BdtKZEjEu1w3uWdzUlga9AZO9fs5h3HDmI9xSyMdm4Vxfd1I/o1L+K
OIDrVS00lYe6Fa4+AmSjkO9XUE/v8ujkFPCwf/1w6MvYJrt1AhoQAE75jEXyyKm4TwCRLc00F70+
9wOrBPkLTNuTMwn+lZHzz6wsgDs493Lc3GldQveFwh7b60BA8mIOh1HXWgC0pZGxH3XfoQt33jEH
Ni9TBJ+cN9I5E4azF2vfeYLIhY41NT+VIo/n4OPNTdDJryxjyveQhYDg6ZsOkDyIXbvAmmWXE/Fo
kyvOHOC9HJXuNRij7isF8b1C+a08OvC3EPSSczJuvlI9t6XPNSF/Mt2l0rw/HGQagavO51+xagvr
NVhEfHx7eB1rIJTEL6FKZ1y9x/brQhf+QPhu6beP25FLoLDGSOUGc4Oq/BW8C8K599QxvyN49NvW
SFBfw5k3XERvmuO3P+5IY0l+Rcg4QBULL5mQym8e0rkAGi4PdGO5GbGeYLIGvNui1yTqrG49s4mQ
GSj7aS4lqx7xUl1MPIEVUlEyp8i/CIfNUaztmMl1TUCMjKplfQrmqV+4rlNp6u7ebIwDk6JyUu1f
3Dk8Su/vmqkep5AZVKzyUuZXCc1zTgAEejHDC8/4DqFPkf1YA+uhem4MCx7BMODxjCBhugBBnNEr
6G9fb5vjbJrO8tJ7YO6g4DZzKCZRXG6Vayd8P7nFZdbofsCkauhhnlJyyZFKKwCgi57692ycqif5
5aqTLfhgtG8d9eCsvu91U4xb9yA8jJJq/MFZhZz2Yhev9U828zisFHq0ZNeIf+sd1iIo6fF2m3/o
Ut0DP7LGkxyJvvkIJucPVWzJqJp+grAUtlokh3ahBWjZ+IkwLZtzjNHEAAjnV/HaMImpPIZI0Qfg
4nWMgFJYIUbgipuzRvW5VDG0Sne9SV19YKecaoMK+sOQTf5Lqq/Unm++74fadW4Zk8Fbnj2o5L9b
0NHP4LlJSxDt8Y52K01JMIWikj2Ztg6wYawhtpdwnR4gmfTerMjRRJKR4CJsSClQWDdgRPcgvWsC
GPPKO/GUoIfEBFuPbW9uUgSnZtOx1lmAoMkFHK5EVwbe41rysKGxOmqMcEks8B2Acim7QvcTWeVr
Tnl7EI/CSYpvnUSHuaPGBmGXR75rOiVZ+3Fcq2MzNaybs2r6KwlY7IEAQdjV7ARFRA//Pg+Q8TAV
UMnFALXB1ft4J90QFLEE8mmOlSXQ4TccneJy4LSsJ0CNa4mdh8fkd5a2rFbBFFyMpfLU6Qxqf6o4
7LVc/a2HS21WINmbYq3ElBOnKb4ZcWqf5lVzpIcXKFBrayMS2FEk9irWqPa5gsIvDSRojaaRHGRn
czVZw1I4IE42/+ChYWGG4OltcREz60Y4xdo1CptkDawiTIhsssgqqpPqZS/kfz6KNr96yAWiLjEX
d/41DbduRxs93vb1fc5jOEyjgFTk5E2W1F0h1uzwkZnlzeknhBgJaSJGdVu6AyvQNIca0OFK8gDZ
HndfgYiyEgH4nxE0rZwrOzd8B5YvlT7eq5jCfXEb0C5KhXqjTjqb2eGrV/EVHHkfIPO/r+Pt8U8N
dk8WA3Qsd6+l98hTkoQ2rbXnEowuxraVW6sBZ7hBWjSHjrYBs5AzXQXG11O3tos03P56TH0gIRs7
c5cFOGUmu59gDrqItoKKFjdWD/EBlFH9bEHdRy0rWQpLNoP+l2m5WijnBLI/lOADG+EUnj3BlN/T
wlifxa5W0pHN7kn7f95IOBukAYMNoas2GchWkQ2NgHTa+GAdhEb7Y6gB06w7WCmuLj1cCrkYoFMp
7w+Bt8yJg9yOmeAG7U831ODebHGd/Chqcl4XMnFpxMWod1PxJ6ZUFoH/DNFsy4Icky+/6UKc6/l1
knQ32xMIyJowKmA0OEu3gHd4ZI1C4v/QcqZbTV+3euR2FZoriGEEpuUfR7FKbJP4FzcCccjeIHn/
hajB2QhWZqJeS01u+kcOu642w0MLHToX1alJ32hZ8SrC6ph9Fw9rz/cXjwsqS5g0FikvhaWDr/u4
PRa3fB0vsRvfmwP/ZlwkFWZv9eXWR3rltJvlrqr2sYSQXgvZ86U8ZVC8jpnGfiCxhajAPnNKv40Z
Y+RfztskQZlxAFj6FSWIv5wWbVJMqy52ArUhBxBT7vL1c6PgDCLYs2dxNRvivRz7NATMgnj0xyPy
jJoHcdPWarPqDxyYj2NYsxd9edGC+zDc0v5sMN7+0pqlCYqru7MW5qNk4a9cFlErxHBGni073dNO
nmdXzXpn9M5cslp75XP5xlApGqVPpuF+fpTip28OqEXkf3wUhw1Q5KCzgzNe0ASesjDuTY7wPVKQ
LLp4YRtyWTQ8NVRf8ZLz10TJ0r6RF7BoHoqxMhjBYCm+E1Z+U9aHgJqxIZILb5n20N9VlFjAzMS1
eIZnxT+DF4uR6Ye0ykZybtnqRbu/Kmp7haAEz9lJ7+wV25NpBTbYQbUTdLlmb3qwc9SpazWqg2No
b9PNS9gvdKNWZw21lt+GyAenw4DnVyrbALRDp/PqKa+ZcFyHVJ+Cqqzak6DQpgqeGjP+ZiMSgjED
60byDtJjG66psJuQf9evfSSygVJRfccy7BkT+WYd+EGpqFpIItXdeRW2DbxkiRUS9jWPaAjtWBIj
D4bExs6axiTbtO+avq2w3l7/AYk6Fb7oVu+58fUt3B+hy4RGXTtnWfVlZ5ZAQG/EQ1dtQ6d+jjCh
l9lUs0prBPplh/8OHhTc82MUfLjJ1qwf99ozzOLBjj4essJKgK7dZ/puoaT7414Xr8ZmM+Pep5I6
m2Q+U1sb+jgVQuSqnPs6t4S+2idagfbniyiTnbfkhhkglq7FcIniZ6TM+WO1paaVa9yHQ8RdZa+v
OQpHjBey3pvAGV4aXDXYLUmxuKCy4lPorE7Ash7cLVXZl9ARE99jHyIevzUy2D6nDTIfZ9Y8oQqP
4504SfM1fY2yy38ouYqpBR589B86GTxQ/RiP9K5s7kkdFXFTtCPhPwOooaObY88247mLxAPnXWsU
R/VH6oUWpixlr+xgFuak+bJlGjlka5Nua8LHx08C7z4pC7wQjgtuwGxB3KbKOwbw4R36xQDoxndG
PGvpN3VUfmQw623+EI+93eNlABEKcQCQ4qxygxBrQhC0e9MwhBxXSj/S0Xh3r6lhqPN8TMXbpNfW
wXM28gMtWh55cuz/MYdddQ/mC9kw6rKkz7Tajj8FwhRCccW366Mh6msWL5SxlTXzwUqlfPYNsRzZ
C/AjP0hjHxL2rIElnSR+Scn6osLk8Tc82U/EPbFbCYiQ2DHry7CZYtcNWw/PaB0y2OvsK/pM9Zg6
ufgR4OIraqYkI41Zj5U2CD+//5S/hIrOolIKiDfO1W95CXHUH7V5LBAGrbhkKEsAUkSvvkGXu9kl
uFXY4nC/gRDIYVrFkR1iHfY3ddV8jPMT9grJ56BxTzxitp7ucxTMsaMbhNjqGuAJSCjjJOJhmpXK
LdwblGI0QTOy5ZlHhI/LnBN2GrZ1bdPMiTL7anKCnKHlNE6cg7tCh1rg+XAaLqc6WoIBr8viaUo+
Z2QvHX/q6pCaF0dbIwFwalur68wKTzmswCBlU4SjxveFMP1+XLx9tenk5hXY7DL4DO7shOlxU8oc
QyiG7Rdht2FXrAYbEah4gBN3J4MLXSxFL/FM7JU3zHEC5WtEvBr5dqEQ7FminnjgQQRP3+tulNi8
yVhMjpXn8nny8Tf9Epzdqlal4cy3N1clrgBexzmO4oq95q0HwLFhhR+Cc1O54N6y5lGuAx9kfTUC
4g9oi0M/wK6odTz5IahPlrlFEDzp1TdBGRZA6Za3PUaLEqzd04XmJ88hUEpTBgEwKkqNWQa2ueEZ
B7PyFFAewJ/+09nDU0iDZ1jAgABg5t2r5lI97xmHATTkipgP7JC5sf7NwFBBvfVo8rpTaLZ0Eyqh
qU1xmc1zFQcsLd0jZboKA7gAory+3rG9L9DJOBVdeRDkesXGXvUE67iCNs4EmesOKAC0LWU6mJU/
5gRzGm7hlm/zvXjYG3bivI8DPmkzPgAKMjeAMHgZhqVGkFMAHNzpDS7GKDqvSibOVFbzkTXzyqUh
kG3Jrpk7LL3kJMZdU6QrbtmR56M1ApafbGZ+8YCogOxW9J67m7LANQrjt28pgrdABZNFAq8cuy5e
HPDN4TuwDXbw+HZfNHmCSUkowKo4/ljKhJd4S1Q6Fo8RIWXJpKR++nh9UutvgZ4mG9UDgWZ7Dlif
mC5nemgd0AUAAK8L5hsyF6S6Zg8bNm96zIEMmsgJKk3EtVCJwW8NbN6HXe7L7l1XvOjASk1oVoIM
xxllIZW+PsswnI2gNMZeRT6cZkyJPnZwWWGYJPsEXXhuVaDewWYyalFhfgAe9J12eLQTMwm/At8O
aJhL9fNufKA7HXuMGJ/K83US2L79hfOnlDCx7Sw5UyrL6z+56MCuQZFysQ0m+qDdRiRxo19vIWB8
t1ZI/iBArEKxa2clsDfPWoxyvO+A/LNVWIuiUcnoULxuTlm0RpxkcMHit58lPMo8npvSg5TR9T6/
aspTxiXPQAasfe2UtKLmNIUJA7nYCWaPdb9kH5UMA/UZLV4hzOjrXGWedEFQMJBDFrTILndC7KXk
HMvFmBTtRCpT7ftpoHML5U1+GsoKNKIZ8Ce4A3cDBiaDkqPFXUtDe0BXgGVXHKuy7ugLe560e6fA
Ggf1l69B4Zwjyx7FFvbv8tPw+7hrJEx4OSBeo7l/pgii8mD9/RVUxMqodMxnlItxiDGf8Fq/7Vb2
whGwoUWTNV3+gBOvjazeMHJGubDB0fS5TIguQpHRUt00PT9Cp6/4Ec9w4OK8yQQPGz5/A9Qc13dJ
Egbxynkse02j2F6h5L5SPozGARmuGFpwno0nfBKrJwLyHRv5KTIjBECJusdAubb6odRLBwViBaZh
e4KkpBONm09SaOuuZoeqJ2kI8ZU2UL6AcJ1zLxyxipiPX/i1cfEkccFWOYhwmcM9gqnKvWXZidxg
tKspGcJIg9khG8238tp/GI9dkUROjjYRYlXcCYRGRmN5vjeuahl/RtTvA79BCWiBNLhAMmch10mF
nL+mietODI2rOUDABXv7D4NPTsbzrd0MtXCaWHODdJxTKJpqJZ8jPloxmgXTkfq04WQuDdtyjWRQ
SqRXN606+fJ0E3tpDIqAtVo4JSnFj7Vfcy7WIJXPDK+F406Mm9POdpJhyFKgDdjGGAqlVCLCq3CF
d3begVqn8KznyR62eK8IcwKOmh29Yz16PeVS7VYh1qalexEIxppZFsjHmXv7g48czDdrjACPUyMz
mzxzOVhgO2i267MEWOo7z4x3UwZ+1we4hFToRdiNREXzWM5v4QVVggmWamn9doCNhE/txIZ7TZ6W
Xo7i+tBIszqeTPC1VYZRvB1S+ubaBQ8l45zSOtefyaXAZbZkEf0b/vrRh1IrN9FgR1ipBiFZYUJI
ME0B43TxVcUWKOjS+878hq1oVSvQSW3rjPCoZxH7ASJcBaShRpYLbjQeLrmxspqHsw3BYIEvavWZ
UJlIBUJ9wvROqQUpQzVXyPYq8fdFlQiszqCW2+8Whp9wJEeaS8XLzyV2qPeQ60vSFppNh1Zekn2F
HfvQqfSKR24LkoxySSzrKnyZHb5On0XHTo/ZylDtxgmk/vYYdosFXAEi0g71nlf7lJeOJjmOMiP/
/YXjNv4Ig4O4D+81vGiprQPgO/t6ZoqUQVlr47F7kYAHWl1e/jfVjj4fxSEopWu1xc08K3XU2jZo
Y+se1BAxF4kcsgrfI0mQYxypUu6y+dNoBcFLpDfjTUaNfbIgUl4d9nm0yZ6fct54fxOW52/8pLjX
e5354nT+vslgyyPSC2nLLMy1QuiSHv3+J2lKyqGuG6zNjFVIv3EqbzXl1mXNmyojiO1Gp0pAq76Y
klkbg44yMwhNxfH1Rwj+FUrKrbxrD7eI8YApN534tkbB5Ln3jnN/zC1/ktMQOAPLVxM1BR4+feb4
0XZOE/X3s4YdoOelo5HDItWDcwU8g9upzET6aErUveKBZ46J+pAQo0J9UcgmpFJMI6BibZvb+PtE
Czr+5/pylhkXkkE9L9YtwAzGKcAw4TBEtVvzpRPXnnwSF9hCRSMVKvEyewWZSPsX0roK+Qe8bWSB
2WnkzWLrTtqvXU3DFX2hjfdwgnILH2/z3gVejT11E7yK5nKo+Lf22UxYPINn089Du3xkQNrSkcNH
8zfcm11D+b+NksSCh5FG+xEMQjlUIeA2a/wSu5Gfe0Y/rIT72w2qtp9JqyLdUOTK1iCh6LrO5Hc4
wlJxxZ7fqRPBfpCTKGjLcKcfd2qZ185IpHzLPGT/FFPZTdg03Z2DZ5Vv4ynwWum/EIXawI3o94as
4F5y/jvt92szMu5zQV//ffkGelu4GLtiG+CNOf3j0yvjn2xPkR9lpOFK0KahPMi7mMiGCc0woLWe
DyWvoVpr5bFlgVErckt4DS7R4VSXPdeCHOYYPtqVmZM4Dsda80uDfwpONCXJpSB4BJUcWDTXg5NH
uUojmPEu+Zrc7Jt173/Ys4kpXQOs7dvMAgOge5pw+7CaKnuwYXijhtBNoipVieAR8lOiQ73y8H5M
wD0PfzIEc4ecX0NKCUNH1K+l5Je/EiPYfsJvPQkwsOv6DokNS2s6ZFc4A5qg6e6TOkQeNsvDPeQK
fvetbyYukKNGDZs43e1GN01VKA2l8ixJVGviB5mue8hfr4hEzbSZ/tj1BG4/H/Z2i9p3MrJKRFjE
cTRpap9BI1Ab7xz3jxMJ4WHZZ53g0kTZfcLAmGlx8tt0KtsjlHBQU8BktrF/LlWPHmhViYTjIBkr
4meZkaHfT1462z/inDHY5hK3s8Jq11Nq+yvfa8Oc+ASYA1YcfCUfugL3VD4VF2kfiNbd60IOBhPG
ysSteNIPTWdhsaHZw42p9Oprf9Ex09b3XPQdvCCNsXMbksVBDbWnSdXJbWLLBhIkkoEIXdCkRYsT
6VXwmhiycXQzT0+PWADi8H07r7ErDYGEzTFI/wpq8WE46C00kJBOPCIUxn5nYIOTKMmXo6qkOYvh
fHRJN798MmWhQxk7GOWbXHFA2jVi3ggbO2IGWZ976MLnsJbvzB/BL7AEC77utxK2hd7XqdPXizJp
9EMnT+LH2CrXPSYDrpqDnW7DH3lteP8OG1Oy5uNUAXxJtIW+5V/KLQzUhVQFg+CzVqkWT6n8iJB/
hCxpY/MVm8x6S0rQ+TudBKKxcQv0cDMROeocwNhM1FAEZm1XHWi9Vneq8XEOvDuQ6h2VXid38+jl
ZUIqXMaigSlbjSflOURhN3B++h4wkJZJxKo7I3PCcTlfoJEPF9hIivtoDI/XvaXMXZ6DSqsPQZ1i
Tafkl93JVKmPxAxKFOKXwKKCeKZF/YEbRf7HuUNxv4up5FdvLBC9dJsWoo6EY+xf010h1B19ZFf1
J9bYvAdxLZiPO6Q8Ev9xjZGlrCYzWpXikT64ZsooeG1Ar2mepB/SMu6UsnXaPBnJC4/u9BlR9a29
/oV1SOtpLCIkP8B8a2H0FJuhhyXFXcU46vlg+3BZN0R4/qaiS9+aJx3y1MRUzd6Ai+w1oooC5G1s
pvL6m/6uZrfshAJieVB5sRWPEZOJti+yYsky2zjkofwgdsWUQ1lH/xT1flxZhRgX9DNTmgVtsVIw
Q/nKe/Dm7Vdyvkv5q/f2Y+GJ1Iruu6WlNra30vmgrrGs+DproC3Ebxga0XhsjqRwxOwAnB6x8LAX
Vv8kyEc41uAXQdGBR+9EjpN7VTppgIhKg3Ge+HOOYWyLf0cvDAJm31WK/2pUEPzznddI+FwUkiqd
Lfe9bTOATNz2Ip4/IeuJo5q1zsiB9iapVLEPz7Eh5rl3Hja1M6SUQdiUQ6x7OG2h047sZAnGfVK2
e3HkNBHfKfNn+OJhwZJJJZmvWISnC+vam3l+l03HBtdeeNJBzYc/ULI6xGvNxWmXlqVFxhmQBDJv
9D2WSNP9eXJUzaOaCK3zszZz+hjPJ1gDq8lJI+7/KJcmPIBgDwCD34LydqsCnPguvBYd71O57hJT
UH8aTFvrPWFAflZ/zI4M1MfdMaSLAi16EVtjQowGHW7LgZp/twampOrFD8IYUMN7bLoVx7+q9gbA
ILDjALTB8NlFjN0E09sZSvZm1tlC5Yvg2SU7RRO0WqKx0w1SFA6R0MXemwHl22C1+eqEuy+6l7Ut
KVxIWl+oQY86yZ8l3J+PnyPykQeixWCpSGRQgReunKEl9ov+NMGouSJyER5mM9uNhSdzuO3cLYZ8
2i5CqOb6EPCxGOe+woG77UmTvv/EV09uWnpfKLKiLH/gFi2iNl3mvnbTCuSXZ0ShfPtUzNL7rgd6
T52NMm5l3ngpW/aWUybG8MhIDoJyGVYlyQdWcARPVRRUvByQqj5RtgoD6QJdL093oy6XKMo8hyQZ
ou/8WazYRDnheXilkc2LXlRrNAS58O3JCzOoKAkRu7IPPbLtAhXlZsDffgB4NwKEgKG5KTedQKUl
N1iO/m8o5+ans4lmjN5fXjmLyG9Pynqw9ramFxVlN6NR29pGXBmGZYUlIMDABv94tUyBUcDRBUoa
wH/4dIglZRifz8DN2EbfP6Gk3ynIMGcdtMjiDBOVQBRKALghKdAlqqi5hbvcfg+nEf1LPkpYd6BF
Vim3EVaR4H6NjWpqA70Ue0n1AVt+STMBrpWbwOjJrGOFnb7rXg3mb9WzUumg543f7n1d6cwBEr4P
kYPH04gAz5++/fCgAJyoyXyNwhnBCsLKWEelsmggLU7BJwXTghwCc7xEvbhNqPRxp3Xa3+h437z8
bRMRyp9BCEIdcrmds+kZ7A9046egnmjFZM50LNLXwxHgWo9uaI5ssWFqJ1O0KwP6GRhxJpLs27Cj
LF7HsYEypqtIbH7a4lHdIl+Cts8BBXs85+L9981NwCIQNetikjya4t0abhDhBYn+hlDNn1wD47Je
Vd9+tiLf4bZRtR6Nq2nyMtvIWpQMVo6HnPVHViJHT3nq+/YAMSmUDADV/fEYg4BDDD2ybdubhWtZ
F1h+OoNJ4q3fONJI8I/lLqMUnz7fo0KaZGB3FaS5u90IA8kaOQ6fw/cZRXWKvCKd/l9CBvrEBZ/V
XOVShrLDwM9e28HcKr0nc7Cw5E51XPxrsX3s658kiwBBMVzk4zdopd1Xkz36fxlSqlbr7ROjGG5d
cIDf7xPMkIlBYLPnsYt9L66c5+k+Zg+TnpTUtaTVgsjxbvoHYGTeJF9Jk9l0N9nIs0+44Cq/GJtL
VU+c0qu8gm3BBmTLhfvALb/1FOPLGGt/JpokH+2wZmnWXyJEpysO9oJhfWof7qWhp+/oMspcP/iU
Qd287bb8hLj4e8grzIWZcQKQV1cS12OqUVri0rlX+ff7uqBHJxhw6KsM0ai8yOhs2PvvY8Jsb/A/
kF8OtYt48WxH/L5J3tT9uuG3jIsg+lAJK+XH+poap9ARLaKRr7KqFaJUH17it0uT29gUXmJHW2EB
2c11XxCjVkC8cEda7QxTiCQwnKubH/397v6CwDGop7YP6vhxN440b5QfeOQsxUnKR0UnlYAjPozc
+Bj/YPdsGAiGJgbCzccfEq2MY1nnAO/OTPcnjR72PgmVXIY6EU35QSX09eXNbPuv77gyrfxvhtyZ
UwaGNg5mLUadmbYCwmWWLwu1x+zFofmYMNRqXKSOkv6OIS7ZBFeZL8S2yme0Vy4t20zA8+3QYsYR
JZ6f8y8aq91mDzU7pmjde/s3wCzaglTYUNJN96w0N11BoUpjg+XHE1OLiBb7lmJtdmcZvR+fsczq
zSRi3iz31dvLlPXlaSQbyVCSRHQl7oUfOm9DrDkn57Fz6kxBFm706m/mV1azyoSHEFSysYQzZi0R
EXo0Q5tC5y2QDeltfP96pvVqikj1tMnb8/VcsBbNZDkwZB2H9LFyml3FFuULy+xay+wKsvgpXAjg
UYt7CHagS10+EFy9RsVz27NjZ4WjeT+njcSZfdchfzlIakA8szKYndYYFokTfziZNiZoiZNWDbbo
hMfOyffT4jk4gzcxhwgLR5Ui57GPoTtdttMCLdS7u8UOgSdfsexypItwZMglDh0+FHkQCjA+PFqQ
Sz+E7SgxNgG7U0dyW+oVQ5oubNvIxaO7VXg8YyySreIiA0DxAltMKAimaFmCzE7NV3tuXiJOcN+0
Hh72ZfEYDtaKte839o/pKHU7fjGO20xSYEViDEKtcQYQzuveM9CUJXli4aYj9oNZAL9gqKJL1p63
9niFkqEAwYhOYbwWo4xeKU6hY1EDErO2nfE+KUk90xl3aFYQUAKcEZxZ6LS1p8kBv7ddxrTkxFZK
U8tTr2r1yxh8Qzi2bAX4kvKe360S2EMY56eJmRbsGwwGahI2nPSAGgVTHDByiMDxLelDTLvQBrty
wPRDf70Acu0SeLp+zGzWURoMVt6OtgCApxi9updyFqMY5c1ZfzM0JDtXJN+FmfKr7d7tkDfos6eZ
p/oyZCjDi6YkA/4aN6o54nymotgWiQjOQMO7Ke+Bz97sFTlpgCQMabvpkJDjWOBVdhEzy40iZ4i6
Ko3Lc0wBQSVDij/wfKiatF2WPcSUv1vi0Ry79cyi1S+2ejk2ODJ4lciWI+bsQ/IssUcSHNMOW/9T
RNhulxLNlLF4/8azGtvp2/brVq04k9TCFQslry04b9YfrFIlhlg7KFOhCRy56tF7Svbo2Qkz8xCC
GlPc1AsQtp2sDlMBjRLsUORBPrjE6Hnq5EFcVRNnbQB/Qkn2yjA2PYkqzOoWrD8RBtphhd2O2/Nn
yVif6c4lz2XtaRVj1RNLDAj5wxG7frLhRe1wUqLKtPAbh7mROP8U+KkXmGf+ieqO/Svoi/qdUYXp
KA7b+zdgY4NdU7Ax0ZyF/v1Fxy3wB3w0TaEbK3SkL2bUcjOt9VM/bOqhE6RDKVH7jtPsxWR9mioU
YQT0bDvHrF2cvTwxqF40t/UY1jlxnaGM2/Ny7nmGSIuMNqsixkwwJl/Zr2toFtRBfSLdtiXYM949
puhDNANz/ldyD8oIUz0EUGWgQ8W1s0noy6b+Bc5Cd3Gd8Ihf5k+obEoyU8VBa0aQaefh0DOucXFJ
GmZNmgqNDzkUNrB7zaSL+NgLCTjreGQe52lusN/XkB8E+o8B+qUZKGxd+AOBLC0MQ5rwrTd/ma0s
WA/aty79o1W3M6tvDU22s6Hao5i9feFp2kII0FBnngr+WcuC2NdTncwNM1asURFW+/bwmhjWZF/5
EqlQCDfftXeR3iWTA1wjvNy2ImTIvBEN26z2qUca2ny27MI4Jj6R7NKEhgBm92MCsTQiwVvgpISs
jAovMyFDgrSKktVE54Zj/XNPIIzhm8dPTD69wfyGm3MmTwYFsYHFj87A+76QTRck6tdF3t5dDYMm
SOchC+7VBhnY5n8JB8ZGgdGXJBD8j2+kMPcuU7OqmWolIFBu5AaMOIysIlftZqef4jGCwgLBdTAP
YAuQGQ+o9kCvlfixHufrQI1BaeKhFqokNscPqP0l+dSqBMWrNnrK+jym7LtlYOEvZcQ6JE9vAvGZ
ZP9N2/NX9QmU855CAwEhZx2fZpggt/bErQXBVJhlzL5wCa8GLA1soAMI93A+MpOjAqgwnkUh5+qC
eVCEhxxvOXuYb/7yvzWkVhQjh8REBpcuyDaiS1drMyrdkwMAi19N2BTstsXExLI+SQhZPzbqmlG1
5t/qrUwvOSSR8+wRVoyi2XV+Rl7hQmy7e47p3qLR6UOWhHf9Dyycxch0if/9hR42ktHtrg8FMH+R
e9HkoxfLecAfMjBcBzaG+p7naIfyL4KaVsFEao9SJiD77oCVpfyS6l7Z4M4x65q0envq1UauF3QF
6A1M0Wofy2qeGDe6NOdFbczkI6SKIXn1Z/aKrdwMHx4E0iiZNQxzdqt08mYNGFg/3wjT8sV/JCV0
weqm5ba1TLsNbRS9OCkhiNgubrxQ77gJqT10T6P5p6pqfLAcNbFny2/G2yPl6AX1N9RkMU1lJgnU
rU7ECaquQQkXke8cnv5YKkVDTxMyPi4Qgc84a19ggdU2Ybj+ELYkJS1MIOlwmD/pbUPOmSU4/uHu
gnsVyJVglNYwZluZzgAlO5k28zLQvynqM+BhpxKPDfdlCcxnztW21BoyggL+VqtjIvcc0wNwB/h9
HPzuMxZIJE/QIojTx4uVyEn3wZDm0IZuVz51Kh+I8TlZdtBQfGsYzKZAxtLK0wLfsVbyF/ddJHNn
5/lB9ArjYjlq1WaCBiIjM7QM71NariVi3wr+hR/laLvPat04+Gn5aRqRXXuir6oM3UMmBLSano4B
PhieKBjgsArDFJkRbn9AtLQNM/WUzqQqJ4sUwooqT4w0rw+e/bstyk49L5/mN2gOK/5SN4iIVB6q
6SZLXgBrHA5g7702FiaxeMSo8X0l4LOqBKkhibnBHU4mBi1WmQd6w8VGzplSRPFrJeGKyiWdeKci
4HjP2PEPITNHyZQrNSFBeFQ8VY/0Ka9fIdWjVNsZHo/0ZlpHycN7H0Hx4hecYyzqpRdfMvwwqPsH
Gz5LyTULsSk7wwqT2Og8vkMOZQs69dxIbnH/gOqLPVbyvMWIx2Km5me0sfATQJT0t0Uh42ivE65L
UoZtgYaBhyrteftgqdcy22CJIjiYyscF7TUCstFEnwPaJET2uiEtF55giDA8AJaH0O8Aq3igA/DA
LpGfnXlUwx8imGM0X1Wsj2Lt1kma43RkOQlj4IYFRcKL7oP2XmxmSOb0z5MNBlzO+A8M8k4X/j/4
qY8ncLi39c3qUoNZucFXnb5qkleM4wv4tISJSMjgqrLTlWgBpcEtJCJItU18LMMabiXgqfupeEvg
qDJ/LEymHnhUqmf2eZQYmlsHeDc0LJCwEzcHQW8B4xnJcC1z2fsfq113CyyZljd22HwNO6rRyD/Q
KMRU7UsZ7LGUOSarEn6qK3VJBn3WNaQntUvQTjCtk5Ag1qAXvGvsb7zGYs3I1ETTefLqU514vY91
O650NkUgSxjA3SSryxuuYVNEzOSu4oglpZ705qs2GbFbip+r2Os4DI/OJp960B1N18yPIR5AMrNZ
fCqjQ8EV30idKSgcPrd1e0smkqWe+nYrOJylgjjeDq9e/VunXze2ESn9JBvR1mtloP142UTcykAJ
A1GLKlr8pt/wQWut/2lQWRZIulFV2wsP3SdvWrfzpA1pEqgZlcYORtXYebBXHmAueH5fODNP8ZOn
CG+0YGp56WDAoBn0ZumDb+CmvRU6FwZJiXxajA7tBsLh7tDGNtmMV1RbMya10/KE21Giwie+43D/
VUyHGFtFQApL/1SQCMJIWkVbTc/9xcj8IxixG3RzkcNu3vqjCrlSaT4SLJj63fdJBZMofNHUva4s
2a50jcPK9Ld0CwDh1qZMQgKGPVhd6uAOGp9r7LAihiZCf8V89GqadIBYwaGUyV7QIpGT4Tolh2Sh
uNfJzZiCe2MlOJbiBEjqmixfBVNqGJ5TeaQbcXGAPCY+tri4ZT8/F+uPzNNS88wqOsUPEVh8D780
i/FigwhCuIIkzMl7FCbs782m4U67fBgzCJw2MPYN2yD4xZrls9gtUv6BMb6lgaZM/13ay8slCn8l
bdznxGFZenYqCYMY5xP5f/0BcAb3gf7rezRmjX4PJj9OBKDgh+hojKe+7roP+bOkwYyDsKiOr3Zc
m8jR9nVjyFhNW5UAI7DMO/quucno2yLeUuJ0reFfMQ2TxSnesMbFPYXV6tkskVzVQzGk5aovhcRG
NDmk3VgtHeAS/G3iZeh1OWNAuzJGl0tMm+VvWmSVlAPs5S1qni1sET4unadOBJTAz8GmpL2Yt4Y1
3bqKtcm+nb8dForwX5FYxEmd4AnLOZq8RRS/wYfDE2pFizSdNjer5g5wwd9sq6lugvm+6txsvTXP
PCK/7VUfBQF+WVkyfbYBdwty/Ya0PEr0ESXxqXRKszAy0Cfx2lKMOS3Tx/lW11NCoRJkpRzL5XlW
Oe33pEDrdFzl54ZN9kNuc2PErPoQ3ps6pCHYdbZjSJ2qliM51I2tEYyVyWUJn9IiQg17fLDHNvi9
UYApVoZRO5lvWgmUyjHZmzc7ODjbfdTFKMnijZb9+CeP0Zw2U/refsvHlYfOprj5cK0+hBqmgUcM
/i2xnPQr91lGEjp6uleEwdp1/2QObTJvF2hkE/yhZ3eh5lPodtfdVs0UyUjAU60TtBxpjnKFOTG2
NRq1+oXCdZycGEf+PM1WKE/gqgpvUIPATvX3YWDsKzVREKbJjZulB1oruMIoMzT1oEhbtgZ2woPs
5p8ePkUADnClCSaP6v03bRS9j4PtMKkOLvRtMf3Ptb8wlVWMubZXReyOr2HXWGflImHP5uPcsYVs
ess+XyjVCiwPHGo7/3zag3Abr02kX7wV1+TG+a1hxgaYTmaAp0kb7wgHz2tTr1Vg4T0md+ut9PqX
OLkgF4b78CE50HMEB87XmslYLd2mMgSPyLkpsKesrYAJUHJqoaD7yahjNCKPE1/PSN1rQ/TA/FIP
RGipOPUgQ8NePxSoERXVZA9MvHsdoG3YHFKV4VDDbXzhsFzxifsc3oQk7gUTBiDVv4y39LoVmEWN
uHB1MM4IQrSKxtWkQ2c7zMd9BrlStXCSsdIbujt3CBvjA8ltEk9dVdCDjkO3RkkkLaxX1xwtIvy4
0otiYu/EQC75uPW6s4hczFTBWI14sUjYVlcPocRT6vk+POX6EMIrrWbTSJjnRQ4Q76C0QKyscqSW
VYcCwFh0YtNE9EPpfjZNpxLASDw7wfeodB9DQwiLoQ+WwqyqWlUgj+Crq0e0o4IQH6BNddl/yCtd
MgAncjlirxA3F+0jY+hkud1La6RUzj2FYOepaXAFGUEfRcb3dcoyFcLdEmt1hObKvP1u8y9bacIm
Nw0DbAZBqiku1xVS/+YTXIVQUO1TRY+zqTfs/UiptCJ5yn+dPWgR+aePYi162iom2CbJjYL5fQL6
Zm7/aLvcTHmBpdfO3astjKaPgexkqCsmDoWgnQv7Pg+sJBR4ZaIqjDdDEnDrR9548I7V8P30F5xR
/hRcGe3rJ/la0hlFPHPiTHqMMelvuaGg2OFFX6X/pEmwOx+/QeGM8doAqM3K3ANaZRRzJIOdMkAq
CiYuRE6103IXDg2qP5WbvhfwxiT3pdpz/OA0jkfbCs4L8a40k0MzK/TIZtMKQ6M04j9s+e9RMUCf
vCtcjAFJ1Vtc6wUIMuxlHRS9y3W04qZPfkupr8aVlWwK8qpAUyzDy5UeDiMMa2ehQeQTVuwB4V52
6yQPuYcQM9CYIDxfxi+Ba3Yia2peylQkT7pDNPOXzD7PIrQLLx3Q080OWWQ3kZDFWsX8hTu4R12N
G5lCy7Np1/6w26Kjny5Xd4GpZ3n6NmgnWudByNv2Z5vrsFsiXeHpSYQl7Lbs/GtQo9Mkp6lxhH+0
Ejx/hgN17Yv94D0cyrk3wSk07ZinT43h1Mz1UFGdErIyV2KKsSvVYLQxXJSlct2GPYH/CVnrdM/n
iEp80iXTZr7YaaOdm5ii3HYwSag4hlUkr6IPZ4CrT0QP2Rr06KsjYE4yCKqh5W7WIii+dYxllHVN
z6OBEkk8/kfnlm8SxPWncUD1ShdnWF+g0r282RC8BR/mfuItnU0i5T5+sj2tDykDSQ009ffxmR65
CYkpbLk0Z7qkedVb0kblEMJtJKb0oSlUuvFa/z7m8836glIMqYarviTL3xZGyo7n+mcVEqp8gUhF
OjDrSVa7oHQ3ZnP+E8WU3G5NZIccpvJEsDCHockKIB5ENwatl02Z8hcUtQwyaW/vs8c9/GJAujUq
v0cH6bHmMtLIPxKpILNpvldRVZo3bW959/Dn5gXx+jplpJR3d3QJRmExwHJcRoddy11NEFYK9MMF
hFi3eEGjl7g5Q7w7QshcTxpjgu2KQoqiheC1hrHy3QfkWtqTNgOGb7RHKjx8Dv51hvtjjZ44ChB1
lvQHsyPZEnPT1iE1UB+TfNJdt59nAdIAXO3ClHKI8xk4DdWiFjMku3h6MmESAl9l/W1ygnnnI4N9
Mb+8BoKf7+JNlnbjLg/P+GRmO+9l1Q7nzUQYNf4YRnCUVGOyuRMI4USBEQzY+r/5TTxndXoKgpsh
o87u0fkqoY7FW5mU/FAT01NE6deudz5Ow7tG/vnKhuaNg0nRVAtHpt0dq3vvTeOe/7T2BpckXaGz
gqiLlJU6hcS+lK1lp8Sq4JqC+LuAsIt204Y3W1Rpajw8CvxGxW7bFhNwEkrlGjSw5vkV8dH2wLkG
503N1HM4XSKzzPETPE91ztvD+NSt99q0ZdIk4lIcMJgm9skcMZ4hB30LT0J/KKh+N6zHyFvK7xlH
aIpsoqgLDlSAg59ucVz3n4Aku7+j0N0Z4rSNFzEK8pQJ3rFALthk71+VEF4UA8CwtWLLQCa80cSv
K8mYQ7rywwlfiKIhdpDNYhrpfpqwBMwUsIBy80LcvvX06anF+wtfUMgdq5pRZpHJrm4sW6/VU9/e
JrEoG/XZY9KA6HlCbGn+7+0zxz2ZdPu93fqthyNrhwvwZanMtrbg4hUN5S98E7QVylpfyeUBss9L
ahF9g1WQNYTElisiaZPklyXxOQJRPhOfVXv6zM1MAzUOQCWNu3qAf+b6wjW+lQXOVme4PvfvqY6m
2TeYsZRZSf6gso7lKijwKInDaR0k+mRVD6u727mlsK64hzxFbJnclR+EqIA9qAgoUO17GdXO/iUK
Xbd0pyObvAVVFqWMjRJD4t+GgM0JV4Ra6xfahHTg2b405BbUqYPsAN90a7q9/W+rFPNCWdXqnghw
z2JZnRdZEMglCZt17M4wv8luaGDbmEYW8sUs/skLi/vunW60I84nh9xgRxlponVyRbWsm4eE5cns
lGU7X3A8eufvmscRAx1zV9vEb+CHk1hdGFcEbPHhMJa56Lw4CNCIFFWfNv5udSWEGCekEv/6fof9
mkI93IsOJx4V5zLiK02XkmyPwHG5vWCa70W6SeHJvmuYy9TJq7fkUCdGnBYKRIalCy/Nji4xBivH
sJmQpmoBKFmra62lziGNvs5ChKGbksbtbD3WUOYvtheGREiWOp1dnzt1XeepDb+e1KOUOTz647re
L7IFinAPOlQo1s/DFxPY/c5fuzjHuMW5+gEzdABruRMHz3zqhxFwzzyCmKdH0LTzJiOJMVNnAB8I
6Q20aXyhtrehXgdrgU6jQ7nCpTJ/pMReM+j8eR0PySnH/gIdckAKarzsAhTTWftqrPGOrBpSPDU5
QGksCbJ5iUaqCTU3/fgvUfhdPeAaW6vqihERKd4t3AO7VgXlp3zosu23abZsDPcTICTmGXiGYi4T
UstbQvgqmK9AIyPgMuz3YMmTRt52PgQDqj/HVaLirGPlIcBlmirCjY7/TCIfZgzeJWPqaWVhqHc0
8GJqVk9gj/A3J/k3i3MOIPajf6c+AjcY/8XOCHjJuS9AOcpuU5iYJ5qO1plPlxJTZsLBf4Os9GlM
5I3DySIp+/M6SyXr1AdAhWWMT6Yfa/VbQEnovIfVxzveGmBeo5qCxoZsoU159uBlLvmUyG83y56E
EvGz2+fEg9yr1lfOaGvLZMKkuoEOWIgJz2yldsGk3SFgTyHNZxhSgEA+f6HaLpuS1soyW60H7JIj
boHJpzv58gJ52ljj1DOIVp0xD8bvwpruDFyA6b1smxphmvu2ik2riSAP4SewEDVSX4sVi2uc4HuX
MFPvKcV6+61v9iU1W32AWTRmoCi+Jyzt99TQPxPm/j1v9m8c/7A4A9BzRc+e+XQ/bieD9/FJxoxf
dyuWkCYD5AeN43wF+IQNiHldsGnw1axTV2K9x4TX0hE9QEOdHCZBA+TKI5v1hlCFHZ47+5tulBz5
6PX7vEKBkojMT2ClNmNRjOfglusSg7Cjs54N/zPIm94slw6fS/2r1bUYLkqsShJRgJDpJFFvA/R6
Z01Z9ag/6inPtrcL/Fh/dpUCFS3DsguySc3DXLb3g7UhHypnszVEOZ4JVKu63MyDljtjARZdeuNx
6mcGKrVT69Qj8CGNMzgJnX+Pq9XA3mcYs8x1vjzRYI6i3XcGUyxlHi50zg6A4xYOE77qtB23GQiu
OI71NfAbOCs8oNEndCIfi1VtkKhmZn6YaV+7Brfnfni8LDaAqfAQdyy6d2i+GgYukd7ZEvlCy5eP
G5EVVFOIKc/PoD+vdiNpv7bc3ptImRxS6ZGrXEuQBXHgRTtuqn3ObL1P0BV3d4mvDDCoUrngkBEu
2Fz4JTAx5Nx+g4t/REKaKjZ3jubQ/tPQvCtEfLyQw9EaXHYcRrJKxaEn6eubEJ66UWUtCn6QD25J
0Hd7Jn5dSQeMhsk2EeQjpGaC6kMhQEOoFE135tp5ikRJLwknvxI45n9YrsjmsymbJ09ekOpU1hrH
oXnHQzm6FhviMkwataxQOeeI6IFEJ2xklRmcD9wu0LpfSOaS1YDubRIzAuHbncDAmiDWWgABATef
7AU4Be7USSxXcLCL6jdnWKnm9+JXBL8D2sO6174cvxtuRbPpLCBNju1MQA5HcFpNChGl4/rFd3HK
luoPzci0zSX5BpNYuTEX+B3ZgCZOAfI7BcrMx9ua6BxE47H0DiUPEzp7wJV8Ggf6aYbQhfW9feJ7
zZQnr3tBU0kfj9ho1kzn1gfzrm8+fEzAvUfVjsAshM9Uu649EMjcGd5Z5lQJMonit/y3+gk5j2m6
utRuzd/uVANxcRkAoTfOL3T2Zz0Pqp+vMljhxZp17Hx0xDqHzV5cf1vPTjB69F1ZnaBiCtwLakkn
wXnEA2oIWpaW7F21Gg81udzjXZsVgz6D0jb+SC9a11s0PUPaHOozRoORd0VmWDWwh7hS8GCqFRoD
u03NvQFOVI0McBiUqqMPsz9Y0SI4YW//7iqzFPQSEBzTr0xgKskqYLM0Gy33jgzKH+APkC6hDBj8
Iy61xE5oLRhkgQ4IzJTvj3a6nPy7SapqwApI1MRMKfv/OoF1BP0CKayvhonLFCP+ucji3uYBMIR3
qJducUC9ZdyyBRGSvMUQwh6tNQCqAGVu4REtuSHHb91CuMY2Nx/6s2wtD7sc3Em4NBT8DjrARS8b
haUeFIo2KDTz7c4fkB8f2SCBRSNKTc5ntCC4XsYcncHbOAa+jHRf2h9BVtKfKH3pWosqnwpvIF6e
qvVx1qkwUsaeJq6++6a2wcsZkf3FVZRDmPzn4ud4WcK0DXxG7ynxLmRASm4X4+mBdhE/57SZFcxp
aWzcSObAxeOaxZdItgwh/RQ2K7XXtEg4XWhwQnbqGINWk8hOsZh9455RiRSA4+YwpiRNQsVTyyQ6
bdNhIrF8SWNyPKZNtL8jtzos8dmwiizQ5503Ht0FQzGzn44zEM8rmpIlnAPftiMVxzaH7Anfk9Xg
LJlpgVsm2Od1+IJHCcSbgeiM2qqvEtOV+/m1bP8kvUiI2x0cc9y32SxmIi5GrbGRe9S7h4V1AY9S
eH7Oz/KavxATlF5VNC47Ni7dAQQ0TJ9G689ReCcTSBR3LDhxclTUFjlL0hSoULz1MABPRfG6DewY
QDLHXbAX0OeqZN7aRTR3fUOF0fkZbZmHIQ1q+e2M6xSTqbx8EtcbQ2/wa3JrFaVKTPMEcoKq3zRj
nnEhtlqerA/mrZ0CHomyuXMnIOdCdZgDJkzCIcuMbelfw40YagH4e3v0ka8CXe8f9rycQvEL98l6
wC+NORu+Hwvwg1B/+vT+IZEKMZWN8AcgZZgLsNmuKaz2fM6PzNLufXAtK2Hqj8hELMxbJSC1Ek6U
bGg/hwDVcb50JZHrCYESqviu1//Qu/gsJ293GA1a2d/Y7R1k5dNJU0J26EGZK9t1fDm5VOEnvYdc
s+xYPwlw4KOtkcewpWQ8cS3HUEM+uTBuFytTf2yPOJRvtk86xvH4G4IA9+3zacAfod3uTP5bGI31
g2Z/oVbMivzp7PN7tImXR4m6iWBojHIcSfToVjT5s5Zquc67EzcVqJ3gZJFw7LHBzYPXZiXU5xMB
P9yO/L68KsGpoJPlOupb1RNInEZcbxulqzERPGdXLFGM/KqHRZQ2Aciq3hbsuHjVW1TC/hzVUgvw
gWAV8Rckg7luFRkO8grODGGmHxSmlKu0xImRRb+KEyi31uXovGAHAmAQKnVVdba0zFh3IsK+x7Sr
AqJ7XB6eWLPqtjuu7r4SRk/8CoQL6o6vNgd/06GTHoXH2jbtJI8yUQh3xDtj/WH/p4w6eSP0DaNw
yDJmd9c60AejOYmo+VAuw/JSFKPBAPcNHkCfRZ/33Pd8iZ7fAhiUu3EsdzGSpdRKOMyrtaXmKG1e
5AUlWPl1GHZAQPWDmGovb08ttGUVpDm/jE0I5C4C5tPpGvzk0cA2OgMmq02eyS04BZTL2bbPNCUy
bd5Kk8GpZKg4tVmXuUDToNXopH9RNjlbAb/cB68HFNiMGksCy3sevd07aXuQTms6B+fkFXkJ1qCz
XhnR3PIoN+vEBYJA51A9Y/A3jr39RKKTbs9ktiBlbBz0MC+PbSCk4tTit/XhHV8/OVTYzjwfXpXE
AFk99kPHd+M7ebCbZViWGWmE0i72oZjwVEm7ZEN/CpUJgpaeg9k7vak9bZZQ8T6kO26erDhY1hzs
VB81BY3uAps2p07I+vnZa4vw5865+e1ZVjoTahxke7eveMiaff5VjecP+36ldgCqvVG8N2Gm8Bcr
Lp8xnE1InlSH1CLMxRx0zMaH7crP0TLxo7FMCsSZ8wuefeaRFQJ2WPPQpVpOBHOdVzVb3Io13bdd
jFZBNDHYYR3fIKPmpOVCzuMk2H0tQc0AnezjlRtulYT8eR5GWvgi2+buZFEwYZaMInUvvWvEaBZs
nC5tH1tESVDUzHbnNzUsFLUW2cr77uzCz67hxIcZuDP/EAFMiR8sTcB3uPAnmV2qTcP4SJcF6kqN
2LCG8Mb6kJqaJGv5VbqaOX2pbQuHOFL+jFgYmdRLkJ+FtORzJNseVCSuUdrP7kz9JOUYd9pp9orL
oOrxSRZ4Vllef65MGg4xGJglW4rucLMbgi0q52eFD2Khg4v0GmWc8hhYK2FkicuzRb/9nET+yjWH
LpNwk+ptZ8EVrEfOo+wBnBFfkHSNOddQ3VbP+hYrVJS2MXLrOtAvhNHEue3yww+yorxDZCb/cO9o
uC3pzgrCZ8kR+PQ7ggvCLsmdIvEWWwGeN+rTYRJatlx9lIQCiLi5vLItTj3TBo68JEG90fm3uev+
DxY8enD11QtjqsdwdNgjgkbdVG2O2np7pITDjuV1VPCM7BlPAPnZbpSYGAt1bZPXaI2+bY+DgegS
cTuGGgr5OzaNl3IeHlEPFDCWtwonRjEcPoB30Z/CoBmsw9hgqMeSVmXSXQFbD7uZusmHrpAlYlPL
8NYB2OgTE+Y+DjckooFwNHXH8SFSXwkwQacIUEdIqLplr7842764L8eEjc0ozqU9kNG0BcwmkR0L
smiWnelDGRjkYjNxcZGX7HxlymB6dBAmS9yaVwbK1Xxv7UnvNWhUxriO2aX3o+Knpt1AoGttmnuV
Ln+SSj6BhAKDgWB+5r1xAXipF/GFlaBLSEVNLnbruATJ7p5rydm5iY84k1GEKTm94RHX6uS/LKeZ
qgaR+/Krp1/+fH2gxyvOXJo6tKvJJXo1LNMs9h29dWQ/nEdTaLMNlhadCw1ustlw3SIGVBknBZF/
uOsjO65r8R58128bTQmMK25Y85fhRWfk5gyfaIoy47aRc+wi5mZD6Aafd7FxbBpwqiQFQrEJAbeU
rWFNFJJlbKzsycn4AOPmkyW4JBsaIc9la1hT5CZXH8NMmTf45mMeEi9M5w/SI/i6g/PUeZrau+1d
ai/yaX5BPU6uUHY+uXzxI0s07tVzEYkSm4TgDNCMuwEz0ZJjioq/3M/yXig0cOoo0Fs6GbyWcLaZ
AYMs7xv1GQETT954bG+gridIewsHx2VMlz3l71kk9XvgtUZBuZ+kXXHwzNl09acQ6rqtbLoBkJnY
Fy7VS/AUvQG+NjNxbAhdWsn3UXoiYRgFqeM6w8ADllAQpIwe7iu5iyKGoeNWKkBHDS0bGQI3/Gj8
2kvxsO2cnJSHt6FwXRXWvGdibHL5OxmNAvqB3YoQo0oTs7+9hVOuXNkif9oCukYXZKZTicrCCvPV
HiRq/4tax2CeKwU3G9ulNKPSAcLiEZkxNXytHMlcxfIrcBbRcYueut0phKR+urAo6bdamwpx7Fwj
rEzlPxuigVBDseakZlAkkBVwEghoXhF1hMZY3+igUCFgcY1C5vwYUZAfUWs+E5/fk1swgRsCjZYr
UxxZnkNR2t6SVeSsXull2jmPUcuI/alWKhgoHf4meGYPUBsWuvYYH61nKth66wxAXAImzwiUvkin
oBO3togwGk4Oe0KoN5eE7YFbJDb5bRH6aQbpOHru9TVwE8gL3rhAFdeN1MRDJkYYsL8cfUPrxbZH
M2Nxk4wMuva83jfelxzVLuV79cSvu08SXoRDl4vUMauIxmfZmTeBM5AhU9G16YE6sLdR89xYC1rm
pUxmvkmoH5QFiY6txWpY95jJFXKuJ8VMevF3pKKDHOBHpAL1pTnE7WXNNT5vLdHkb7R/5ILMzi2F
+BTSkDTLZIjqw7Ij+JYjZkQ1+HM8ODBokabVMOHndNJjncUJpeMWBA7uIVUTBnzneFuuND/yCRRu
8VL23OnKJlRjceJJntsaKX8e4KljvuudJtCPizNZi9gEcjaIhjR/wqVBNH9Hi88EPwZOoXDNseio
vVa0jbxYhDPM/zQpbBGWvVOdp7FHauOLvZdboiShkFPCLraWf9EeaWvyU/NDv5wP6YN7HLFeu0Fw
QsT9HCp3x7qR11Z3Je4YNgXIB5A63TkHJ6b/uAeAWOKdV2CHZ4DKcfsQExMS1bc59t2zZ/6VV8QI
W/Y0GoDSnqO+wnpoSqGiCaDhRwf+MOT6JZXOfvSZuX/r3faf3WLtxU/i5LA8toaIvKXH7i2qi9ch
QqekRYLoxbD/PBSb0ARdA5xJUvqhwemai7scZtdGnaDkKzEtGx5deS85Ajyl6YBJ0Lj+8QtOxVnQ
r3rS6tr2UdsPy/ZMyfBLLQRD590TnnDZHQye5ZmqzP4jgHGoKtVSOaOx3fQ5kI6t3h3EmhVGcbm7
KrrDDPPl0hhp0KKQONTU6rZngYja7113c8FfZD9/8vRR0n3Jxy3Lm3QHohtXKcvIhghuxz4jwPKk
cjbN2YDK8VhSiUNX0Y77fQp+/LwzYDcSwqdAnU5o1YdwZlVky1IuLar4Zvy0FoYjj2TyrSSaUzfJ
7ihDMiaicoE3CD03la21sKp2BNyEecUiwTcwF7FuMKqOSkxIt3hbO+kksec3W1hBGM6yEpXPdYzl
dfFros3v3/Q53yA1guTZKJsMjzvi0EyFgixvPyjwd/nLoZVXzWJyhNQMYGMuYttqeJldD88db2cR
jqqgs9qq8mwO8Xv/SrJp4URFkpOm45jcirOnW/Mnk4qQvqikwMSgDSVrKH2mnVtik0xp0sNQ9Qsr
txF/MBvZTcRR0OPEnN1XqpIbzHuPER79ZiJbt8qwGnaWZGAdpZjbfmOyfo7vcuxUBs3RNA3Ymdum
x/D9TAcRk6z73ulqXjqH2M7xQcVSMQ7sAsqszXk99KUUVBvywzLkJlPjgiiu6W9TRTqIVBlFuybG
KQRkQ+u5uFxcMOidcYQgraPmOw/O8b5VyOpaj9JVg7VCG2mPz68txcXqlwQmwEGMPWIKJJmDAm/z
zvbhObo2TCbeiUoMJBBR30E7nLPflEekpgqi/5pB/GXKqKnojqjJi8HznfgboqOYcsnAgdJqLa8N
gFm4GTz+y/BcgUnIMtDe2iw9Cy9hjukNk75zkTvpxt1/mGJftMtoaSAXlhWpy8hUH8g9oHri8mL/
/b7hk0UjEWuEi2Kff4CPzuV3u3US0Q8fNhwlAwatAJEoAMMeen7Mcit4n/3IumudsfJIGQX4L5e5
nekvqaA0waHEWP10/fvMjJRI9ioq9leDjxj80KYgdGM21pfFeZlJdeaGvcuVZzE9pNtBWvsV0gSM
4VFU74wx2AXe4GokXVCiDfrZ8oSC3BJjqqroe9UPoVgXsbABCI0Spe1URASczc63jRExFf/kVAI0
x7eFVoThVaLBqacB3Ha7Np0tW6YpgZ2TVd9+ubbemgSP6ciie2s46ahl2R6xGSlWSwc6lLocXaDB
FVYJ1f8Ca0QnoWaSz311IFH9PWvRQWuBjzx2xHtZCSUiMA02zpURh/y3q+kJZGBTs1rTKk83FVNM
4YVYXV+6KRv+c0+3jpPt+V9gbJYHZ3o328xNJSk3SgHsYnD61ZEwmI7LlOReghOj+fsodUWQXBHU
jsZR9zIYoEMksPBIOQ4NwABfiUGPLr3Iaem09P08idhS/MftzvxYO0FhcyEqzikfILD+wzARitz2
8y0BgYf8yBzvx1U1AN+b/Wo4Zhdo4BGpgyOGuTIzXimS80tH6wu6elMcv9YqM4wJliBGUmbN3xfE
8p3MYM5mIO0CXpcEnCKX7/P60ZhatJokIdHMEC8HL0mNl456c/G/eRM6rcMNou242f/UEbBlnFdB
1SopbfV+zC/EmFc4EEu6zhMWbENl7yXZdCNyQJTWwLCqe3Q2pHEcWNwqBA04OQkDcCl1qFxfpZuJ
VLD91XCEkNxbCRALF5quKvA/XNLHAc0Corxe2thgUyltjHma3GFBteb54Sdq9FW8MtI6Hsv/OjO2
eZ/zRYYt2L9i51iuq5Bx2HbGTLN4NVie6XFURQsVhCd0qGuc4KIX3pzfYhho5Bj7JZYeNSnQ9vYt
r91WzD55z1vQv/DS4zch0D1TJ1ARFp1VH/L38Cg1cQXX7dDrC6tmMcEAhnFkqeBCGZuiE/t1K7OK
7n2WsmbhaR+MGNOnNRxhdXY1kxsDM9WLkwo/8rQMVt0V4pF2De/hssCe/VnFKSgDzM0PbINSo9gs
B8bLs5DD4diTr4HHe69t6pK/fN/CUQZhyD+vlf+dwkPY4sltutNhKLKKAF8gL79h5A/CndlGZxxw
jOaUxbcYgvEfAaJ+GcFagArfkqvu4qjBTQlXyWIM1HGP7n1+njWippBDE+UjUM1SY1cmKginrtX4
Ic1QnXuw1XiFUyTKetp4e7nTbPyjPQOzNSVhqDLzinPq8Q2AvxT7XbsosLcqzjH2mBgngjsak1pe
1+pLKzxrmKbmXrW7J9+Z6tBpkYk7FpoEEoMInbSqrduW++a8uhfSdkZgYdDcU9mIZDydxW80E8GK
L+zNUMulLbLMQIydpXMpRKCzdwXP2qoFP/sUkP6UWJ0OsU58Y1zCxXMtuHoXKJmKlS3k2hY+Ya4Z
S19xv1L4ayqHtBDJcIuR3ugdqq83YbGlUp9o0WBFCfaScUuG5veI5yhMWlxQ5+SGa0Zt/K7YrTa3
T4pobPAvVO2YT6NWkS8mvwOkBgtLTlYeT0ZXGC8fCTfsido+GfNcdQ3Vv2voJ0NZUKbzA7jA4GAK
0jA9Lq1fjuVW7H9xant3zIapUX6WyYKWgSEZq74XCeVyyvS1XbiTmgHQ46wS72RIWLHgp9SYloqp
8IlUbzND8s+HNkbzToJ64R4PRzxR1ArODay9IF8CcdcX/cCOqWxeexDE5HMxmW08x+rBTuL3PWE2
cwPRRARpZnLmEkqPYXoT0GF4SwK5onIXngW0TDQ/vX/cv0VS6+awyZ1q0uepponD3P/RU6WOO/cF
7ZF+vdTcJiD8jagqwevj92g1gSM/D/QrOisDjAd4sFdA0CHgv/B6i1iyzahgdYDx7JFSU1YBA7yw
a10DLMByVH2XtI9pyiPhNrJMw7RvH7oOZ+CM138DF3WXZMBzRAd4ChKXt5g7j96jFxgHlbza7CE6
iLRtfh4G+ogk3tZHZ3ZbdpJgrRPhY9dUG/i/+BsFsOr3zS2E7V3Nc2ih8qnzeQuFpPcSwStH3xh0
RQ/vECqqo8TNc4lgzXoGYb0SoukGw+LoBzXDQQmHh3QqjnKdKz1q5LqBq/iYsKFP9E5atHvmD2Z+
bZ1iDHpoqN5+OrrFTGUXxbRwOdl3Io6eiRUM63VajC2Jd9ZAjfKBw0CxRUuT2uGYQv0RK6kiEsfI
wrTdiY4lzDS3ZegDYN3aRdzkl9oLcznNwqZzDMiTUHfUdC0TsV930FE8oXLIs8af8UdeJDtAn8u/
L4z6nXJMrUD8vu/B1dvZGynEV5vHWxOPfWqDYgSPfI4dE1R1xqpEz1tpd8saxtSNqMSKKb9CrICU
bYKB99CgWDsQBcJvj6vTDhhJrJcvM+ymrQiHCGFRS1iyuCcnzIYVFBwi7A/irhCVjPH2sF8guHzY
VCRsnT5/LWTxy2DUpbC0VLwxqeghGiY4FZ0eP9N6TJ6gwD3Ya+lUPt9618E21vFPZGG4RXc3JRRs
jVPZ/yX1baLY8DLzCB57qNk8KG6MedSg0TKV1z6Yw291clOLMbvavCR1M6bTy0SQE8xXUIAec++F
5iJUyAeMZYLetXevSuF2L6KcbAUvxHmxCCSeseHAvdc2j+lUSiwSekfdAXaKaiYTZhhKacaiM+yu
xb+46aHNV47UsjEZfLKdLH+pgETMcaDOs3UdmdO0NcEpzes84hosEM6E3mVbsIgt//UQaE0w6ULH
/FcE5O88WoCKqNMLnEJqMu/ZijTBtYqYMmDlGdEmepNuQhcVxlfG6fCXQW+Kgpt48xOJVu8ilhR3
w14DkhL9OS1jsFTz8uqHkwWOT6v560tDcPl4S1NCooFUwp9LE5/Mxn9usFH3fP8oy8j2BbiS2xrN
EJmsD2Y5FunaG+EmeZpUCRfX8x4sZ5Oc+5NRKGLcSfUfHJ9lc1b20790RCjzMka2CKrlyTf1AG7U
z32Dr2RwE4SZStj5xHdMpd7sOexgqYchdEx2S7Wo7a4iuY1Q+T6WPDLumyO991VIHgSzVdR9QRoy
r0p0R13teaPjKiI7VHf0cuFmBgLC0uu0fM+6Q/ejht9KHM58xN9mVxfc5sJiLNviTofrJdMCmD+X
6LPVorFnXONFgrVOI0WGShu9BUjZgMK/hLJsMkLSLqtAYO2QdhRBGyu1y2oun+RjGn/YRYe1oS9f
Ib9gmTg1tFxQ4GYB7NIYrl7aGHB+xh6G8emlOqO1CGZkNqblDNygWBhznbN5K2WlbIJPkVkoyJoc
nakzUH2KYuVzbgVzmgkXcL7hUI6przdg0UF0e033XOQA/BnmbVNaSZ9LZAyEPbNnrp0OrwVo8+W0
1Xi+7NlW+DTxQCSOhAVAuS3BU2XjjrYWgSKgoClFxC0kRvz1xh6/fQqLaqTavCjs/XomPJYpuCSd
p3RUekEMMkkpXr24a5kRwpkq1dMusZcB0cWBH3d61YTs5I41Qn3IgGsL35HteTkygpGupprTe7+W
55aV+nf7f5y7hw3AnNvdZDAvkKoRNtVkwDUG/Ufop08Yk5vmmSMcp0YhNjCmXQYswgIPza2cgoDN
tEXytBMRhTIy1kjQClG/FovVVkUNOCYGhQI1Y1STcCyCvwg76dYI2BHADlDb5aAstDFLE1RpuGU7
0mNd9abbywWi/rm97LZe9rX43LC8AEJ2CO4Wl6ORi81d6FtVhDyVpVoco+4mcOyPrnC6iXDybmXk
AugwrLpD0UDPHpmytn2N5C/u1IzwoD3hJtTn0rL70G6Ggb8AbrGQLcVFnaq/QAxq6ekxXt7Rjrt9
lDqfEeg670xx5yCyrY553jpKO4Qh3uqgm5lKrEW71aiERTNUQn66CW8gNXjgnJywz1CTtlN6ED9r
E8J3CqmclR+wTKH+/vd8Wy3YTqa4yEISRciRxso1l1pu+OWdeXJ+GZyKyAXEV/5aG4kThAq8HkjN
VR4m/IGzJc37TDDlMuRJrJyG5S9r3A4bTha1Og+G5xtPEV+f+cGehYV3IcdcftPHWTPnkhN6Z1fS
jgoamFduL65r/SzwZxI0tzIWfmrZ1ClV7A7+ejYoVtneivEOoydJI/VIlax1ElCAK9pJR0GaX3J9
TNSn9Xgm1Ogapx8wHee1ERxXLk2eVV7DAbbZdADvZGRZhpfM/8mnK2Ge3SiSoHMYNwn64bmAdMLd
nAS2knmk5VsQNG7YOao2llxw2KEAxacmmBV03tYqPiTJ9fVLgeecdNdLGqzDtUpCC4VQXiGVp8Nl
VY3Ykhyk+58SH1v83Q6jEIYOdV5S3sZLCNoT5BewAt3xalcH9VVntal8ML1r6JfF+mfYA4Dr0uUd
OrqoB7FN/DMwtoeqcwVT6yaLr4Awx/HzoaVAhsJrqJ+2g6asgbMas2Eq1KxaV7GbK7Bs4ccaoh0J
VLOJDmzaeBHxKQlckittFDVl/jfrtg5Sgt3F1DCkV1fUT4H2ElMvwvJnplREBxIJFfjfDLS2Vcwp
3UDs3ueF7jwoQa1b20f7g9nXWCvhhEVA0xH0JZO6nOO88CSqDi7r8e2eWDTJ+Cq7ns96cE22/CU1
q7eNyXhTfaI/pul69mxORcBf+m5MQhZKSdI2rxY1ybkTE7KM9cCKZ2x1azFOfHj0zKyC3ZU7+ShZ
5fHvFQTx39jrsy21sugcFGGm9AtyCsG6/e6ziwhfLbczYPGKmjEsySQVGEYuY1LSYjWpCI8gJ28a
lfzTf7aQKkOrw/igpqkcBBD4Nnu9NW6TrteQmwWsxTbyoLIMxTA3/k7kGbED9vw6za/jaMlYsS11
rMlp5IsSs4BzEEv5ay495BiWQy1gzpj0mCF9InxIP5exVSghZ42m5HjwNAcAJuiZfdJJhc1s8Y4p
KQ1R3JFrBz2N2Hr6PhbJfuTuGlqXwYkNkgCgc0RJ/anesY9LhZ9y6X+mnXidY0TdPB4XoeHLYLsP
TZ4K1gPN0cpEmNv3ZQ9NuHAPss297P61QPZZ7M+WasAL49K8/Hj2MoZNYQQ+WU5KDcQJDVDu6SsT
BJwG9JHCoFBRdUS4y+m10SwI0VhihZTXv2eALz2kYktyb8r/yg+6pOmRJf8HJUn02IByjDiZYTIq
lmHo6K0JmIBjxi8e/JVhURnd7H+0DQcpcY6u5srXXLSwf7vYgxtH/+eMtQveo9Vq26FwvzopNw9w
GRjRYlqOuqZHumQA+nKQa50XmdQMXySaXG802L/d6RH0U5IoM2Yd8CWirXd8fPbjJPDDVfv9yIbq
x/A7eVABm412O8AQ6K0yOklHWjDL8zztMJTwG7tUxrJIx/XLP5pnEj+XY4oUv43bOIPXT6aq1Rrs
chFmL2cndt0lmByfPpQQZOMWzMM5FKqQCktsBFTWuwXE4EEveA6DV8SnhPX1vst/3TGlLM/0v10M
TAjuOnGe8xiP/g4N5OpkAj+LHYApvQ49N73NXjJZZ5Fh+HzaqtVscKUFmx7hVpv49mGwGKt0CvA0
e6hn4bUQYwAmSzT4ogVCXAazGX8kGpii7pRsUrIP50kpQkRqgVm66oFKLXwDvDNHUHzGg3aTPeF3
5eJ9upqozn0ebU9NvgbnMdvIQg6YCiFjTSEKp4845iqitcTR6huB5kiSBjVEh0YyT5lpTsI0E8UX
qL49AcE7ByAuH728JOOhWhHhEAdpkplossARbvIy6wdrShB+2qMPLGLIk/0LgMNQqnug7+JzHoxj
hv9bj6VFj21ow18mWtJ8C0eBALxIqW3goDr/XS+GSkI8dgatGI6W03KKVOhj6aclu0bRizMO09AZ
unKD3f2IOzEzp3F04AN5NljgAtBj9+BDdehojDfqxXLMohiGwE96bzioZTYWaM7ZwrlpnqVVUuTj
C96sOgSSz+G8r5uIJXx4sKuYK3+hLeiU2xr4np2pW+ujWpit8nW7WCY4peuRUE2Yjn1NyK/81lvM
u1xUc39ULZ9HeuUcmNP+uSwmzH4SZFokBxZqxq+t9dxXTTNMQkJ+hlBaHBzJ7QBJxB9T5acLJlO7
SHyO4BpSzRKp2ziNEBicXd7jMo23AZ2aW4CAz3aXMfIoXJS6n66SlUacn2605vixUKrAxpm3bdE6
nxoQ8KTawNr6KivrftPWafGC9vP1YzAuO+G+w3SWegHIX5aWFvwtUlKxY9gA3xAsrf0pqWUnDTO7
MHZTUCz6mNH+8yVRM50ZIHpi8yFSf+D+PbMf5rUNPL5sLCYdGVdyko1zsIteoTgULDGKB9HchS4u
LwctoYfxVe7cyHcOajcw6GYLEpnCaH8xbm+byiwOfb6wY3YMafVAyneiID0KW25yRQkMIaCPP/IG
GHm2UHC2lZzQzroztkWKRXMZsEdRc0nMQpNTYmMVWtvoWiF9eMSHCoDMEFCyYuZDGfPufASG6dpb
YFGkEtZeZhpFCbt/XfdRRz+NsYSk924IFfSNHafral5JGbCEfKem5Xhac/BQo5D/iztqrD6qlxzD
QMTsm9/weAJoRtEhno5Q2jGdURTnTFLlMjU4X9yOyFf4LqOIHZ8WghPfLee1Ou3VNs3g3n6NeMjt
pncAl+RNH6ud4+iz8hL2VXly+FWg1dyIr+iITTWtm0M4W5IWkRHhxs6h0euaGPfk/JAezqu6e+Oh
KpblbWxenqeWC7i811JG8pY6YIlXevi72U3nVlDHrqwWWbXyWpZwW5ruJ3GiyJS9kqS7rWxLcX4j
MqLaigovE0i9qatTBUJDDrSekD2x7kF+rP2jgsoG1Aa10t/oTmgBgrtWDsY+qfAnaLrIazFwBJi0
nkHbSsrNmAy/v8FWsY+zdKj5juFlW3Q5dLf3LAsYdZhaw0TMyFygwp2qescqXBwShON4aMw/G0vb
3mw+algo80PkuLbcpmgJ5TofWQLE9rr3K9U+r/VPrtmGWbgupEND3lsyHirnz+IAOvpu5LX2ovHP
obK9auvnSQdYLBwHWpr4MuykSOyrJj3IJIRq9GoHdoSP8OWG4fcYZLhUUg+AaXo2fYkTCO/q30fY
SI34HamvZsoeBn+oWPhOzlvEL+7b2es8UpJYt3FaRTEeo/Dm25fD3ufcyMoLt0SEKwlLHf3ZxUzJ
2SR+HhcUkaX5uAMye3u4r7qIlMGCUxhcV+oWjnIObLUS1wEoa4zim1WFVuQ+OVSDIJbjt/DQSYz1
m1vkSmsTxRRGz3S7ehFkfrJGsNiijHm4Om6koY+QKlTOAgMCERb9FlITkIuQqL2gd62JsvCbsWMv
yjZNsPA6jJdYVmugdeNcQJbXjg5914Atqj8ffvD0JSV0gcBOFqn5JpYjjcqsYwQFHOSKY1m0Pi/0
9424+gYtw3pU4UnWnj6FPvLhLNZauD0KgpHxwHxtC2VQOslf3I96bR6TwR7OjE4/oaPlN7E41651
/AtvoqJJeFIsJ5iB5nsW/ubWjil749WXaRtqE5YUVak+jgORV7F/C9RPNcLTatPzGL4IoRNxZ5k/
I0OlgdKnNzo/7LRJbyyljA65/S+kLJZ0rAMuwvtJ2PeQQcyPxD0dglUf/SSY4R37lomfyv2OfqDz
s5K4QRuxTbNUcUWK0Olz+Cv8xlL4r2aOmonJ3vXcE3bqMw6KoMh0SoGECrTD4iN5efxmFPYfQJpy
9QcJu50kPV85+eN2qX+oLn1/IJe8Zp+2wpCI7xw5Y3iwRxSo4URdd5TCVmE8PsBxP0egzKB5EATp
UlOElL4IgzPFtX68a4Ce46+Eho7DccS7S4omlFP0Cj++bh2GprlFdJl42lhX76y3OaSNxiRJ7fHI
AVQFX2fY8MyUoWCB3S1Irl7118wIoqkyafwXk7ZA79RpWsPcRygChTDWNCc51+dbwA4YWiIJpPIS
SgcsohIRPh2O8hgDt52omKtDD04BqsjqC7/88PJHRjfzyF8gT2VROkB/Z4g57VHs/AZ9P/r3zFSx
3mB5IZZj9wUJ7k3ovU45focjP/NUMXFy9v8qkqkiL82zNGJWRdGTy2MZSmfhyxaR+pZYr1dn8rdn
5xuugI1X92wY1pDN+Q8F5QLnYO6StlVcBbmxUIXTng1tFu0m0NivEptiq9Uc7ashqwpnrOWVvpLa
PjlwRXi1R00q+wc/NAkFqsKogFH6KgPoheMeuzQyK0fI2SWFAbC8nly9f+ot6kkyuda+noJIt6Nn
nkM12b+nGLM8AN8bpNzvM5apko+canlNt2nHqVeC7u5vbinmuzayUQ5GiL9A3b8KgLuoopyktFil
qlc2THZ9MMHF0m/IqU+RuAKNgNzqPfAmjDS2rcW9VklGA5HUmAc7SXxSC7EvgTIXA0vdAU9NxB15
aE2enYaJlNODFD+IrDA/YFQq77KaZcQCcNnPVzBMtMANaJGgwWmv97pIl+zL3twr62YY3eQCzhkv
/1kIH9VKJ9NmuacGTtds0fDXHymc4I5JXZi0pzsNAg1GcNrQ2PBTfLwo0F3oA7jXDbNLshy/wjb3
WsME9Xue3sTJiQZiD26mXVNc33RSn3EU1lph6EtSAbVv2oIijRhEbcuNYpY84purnxfTU26//Ajt
Cujkc0OJhtL4JJBL1ny+16/nztr5TFZJ3txQRdRmXhdgWfPvX1VGmq417SF9w8WHq5/rtCCBf7zZ
X2xjXrO3nEdgoFjukjDEfTj6fi6qWTt8ShShHTsh0aqAeDek8livzt2ANaWGgDzFNjOKIHf/8q9k
9fxaAPr6ck4KMh3/8/7+qpU2d92G8tSgwBH3WGQLAnVo6wS1s8V3pV+WuXr0KHbl0jEuQjiZW2lV
aADn2qSVaP22Elw2RI+FCp7BP3hnMsc2BakTn7aSPWhf23gcOFiNWOaIhAfurCT7xz/0fj9mLneq
+a+yPcwJRP8T6uZQxXITl7OAwhxIVd3qiM1Aplhgmm0I+4LL8wocNPH+EImk9DozUY331IfxNZ9/
/sHRT3RXzVmv57IlWXAGf1MlrjOSw47skrveBcpMuasCCZypEiUwG7LFOk5J71UMj7ngyLyqLS/F
XtNbkoDaUt6Day0K8fqpGinElLWOTZBtKmUrreLP+1AJpOl8gD/yf5qSXZ3PYseYBbYaiqtCZuTq
uUFMwwHIg6sjVxu++h3vHXai8ThkD611d46CydC46yPyMtO7GTv21Q1CCwSuU9x0RFxf/u68rqWI
Y+afQKjIlrJITSvdRh2sqr9f3MofQXBpoPx7goRD6q43yDCFOtGarvmuH91ouf7z2ki1/4H+JX4s
4MRu4JG0k2oiMJ/a7D/N6d+OkedloTmIyZPrV7e3Cx+WbIx/HIqAF/D/A2PX6C7nl3FDIeBcZXBB
qyfeAFXZaaW+uR3LzVlBMWjn3u1AIUaEOX2LK1h58z1yYHUrPH0D2KZ8hdnIb1dDHljypal42uxM
QxtH2e8HZdaUAdc6v/GWcJt6WIX4BQ2F/6PX1rc/nyHpTX0Clfb1MHsVETe8SoeOn5alf7+Zt8K7
txlBok2VMvRIeIaMldZwzypPVRmQ65PsfSGUucmwzC1cv/zB8gA6xdo2TQiko0pcxgiGbXl0+Dmu
k+QVhfNWl97kN4R/2/TBQF4SV353aftnDQ+JQ9l3zTr1pqWIbyb0Du5cXoTPj5hTgBpRPfVxN9op
9S0q/tQ6Wrbs2C8WovDSrbjstvr+EU4dNE/Fcygh9Nzv6tF4sFk2Cb5/uHn4dMrxNsDXAqcyeIes
42wCzBSYQedvBLqI6d75eolpR70a1shYrgO347y3UynLqKdgDCUuLgq3r18SFp/kj+E+hk7koEhV
MJ02I0Hfq24gZl3xxZ4D3qtL/C0dw8g3wj3MYAEexwnsiw4G0yVjJsgBP/i0wZKQ6zmklkgJ07RS
O+cA/9Xzm1bCUDqN0wdzY37AKwWda9VGfPOUF+1lH2GmBs4jhL8cxn3E+kluhIZjbEngP7QK6uhX
nx1JcsMoy7ygXA7smEEqabuign8VZTRcwPu/fb/wT4Q6PmMBsBSGJ50pVaGJTTL/DOa2HFk3nhc3
EmAO5GOo8RNjgROm3jBtI8LE38OWT0oTRNyVCM/w45Rw0pj3n9hBstXTai1RG+cytnEYE6x6o1x5
3W9fE7emNvTqdgM5PDqVixQWqrKF3E+E0dZ8ErFiLfS7zbIpvuvSvLbMpogIoxDK/B/ab8FLoG83
hXz+B4a9cZNg4bpXYLR0QnR1do+/vbP6Bnz+TAqLk6oG6VDXO/4lNLegdvA1ryIOr41UsABJLA6J
o8wjcJkJtHJ16PxKO/mr63nGM3DCjYjI7Bqtmx+rUgQM8dfQdWSF4i5z8yBbBk/Na8XFRXSfEbIi
25prtotiRZBebyLuOm7SrEqkseuUurYLCUKWi/MIE151ves76T4Sy8QQHqO2lhr+2TzyFgjItuwL
jHCHEc33euqe5OxCrksM+gJfQZYmPUcMx3ylrO3IXIz21M7Df2qOt+8iJ2A+tVcayvL5Dz/ErAmK
uUGTZ4otBoDzC5GFaGHJiEgiDrNH3HrVE6AYVoNE+u8i8iOAbMXXnbtmfanXvYZFujLl/vXCElWI
lbTAAnzM4xViky4doTyDGOjXv0HexHxsn1SsNDx+45DYmsdEjwstyn7SOiEQKoeaCZAM5yp7HvZ+
0y9mF/8nq/wSIyh5OZoVu1SPPBU8GxI48ZTVO9bFXMY7xDYtl4dJxvrORy7nd+nAVEVVNNPac4Ea
OWgK4PRy7bbKueJ0LyEIrjvGmqwGqU4hgTTewZ6rCQBk+JU+u330kb2HCs66/d26bbTwQquVgPTr
N/RDK0MdQQM1zjg0ccsgHsDybMBXZvbxFCLPorPhAyALYpMTbg69V+NM5SNYzqU5bn9AjMzaS8lN
IjDi+UE6NiFAzh61t9vr/AZqwz78PF40PEyqDD5CSj7kDQNbBbuEmmFYzmC0QudubSNOft66bFW3
1GA90bAtoGliZ12Jg9zxDhUr6b9cbqlihDteVmVUAcQ39z3+WFhCuAHUmDngJ+mCcI5DgE7+MISm
y0tqid41YNbDl5YXhvjWCj31uZ04bWsRCERPOJEsZ/8auWNX1RWL3uMwpc6uUhCWxT54l7CAorLK
XuOcQfGpGLuifU0JpYVyC9KOmUZfN1NGH4iW6ELuVFW+HaAixKUCIfFXx1Ksy5yfQhB9Cpz1ej04
EbPFgzZqdYPT6+f9x/JKXxvC3z55tMXh7TdWWkwRhvwwajtFzvlOrlAN6dKlg9MeCxSLaxWEhF2E
L1LkoeQZ+ZTQtYgp4pS4iSCGpyS2n8ScKcQyTXLq5mWKemRHPWszZ7UpOMmj3SCbBe/oVhPuer+E
fu5k5+lkjfpNFiK53hBBR7/EVRCDkfFJY1uCjDwn9UKK1NYoITEZjHMRdwrIs/feZ5IdFLeuh/s1
NpgtKrZqHpxmDvz21+hdI1hrldaoDpunh+nMjyaFnsz3aCfh+FZHRRJry67XhALo50INDZSUA3kf
uEVVRCZcAYQfmofsQUcprgzQvFEs/uLrCueZTNT4lf/DdBRW/5LnjxvIukyoEu4ErqHn5MF3cQGI
/vZOdEK55BoGYfQ4RblIEKRLnNF5iLADOUf24XMUp48G4KktNKl11iA0q0eaxnZNr7407NuhHdcw
eNKpm/H3CxR094aHW3UxVolHeLExFtldkJD2yhvDkxCUOfW+weHmyjX5izJLnqQAg1nGW0VApOHM
iv0z8nBH5Dfe8xHdw18Euj7D+Y6tdW3HzDGjkd5ylE/OlGQblWOKoQfi4uer2S/Fa8jOH1toAe1X
korAQG7v4Y5Nn8om1I0v7t34Lnk8WWdvShPFGaifQqeOuxjDDmGiO2gPWf5rQvB9XNhpTgOLO63H
uypocHAx2u/ECbFC3gDTq7RZ3k95ZU42gsXOi+/9agMuVcx8NTiZC5Na7kFlXerI8cNfTAHz5fge
fzhNUidjTcGG860ta+nT3iZmfv65MF8S9Fn3H2qncGNRiDnzA36MuEJZf2FHA14+hO3boKCMYF3l
UMKCxvdB8Bu7FJSlTCfCdlSAgzT/y8Uv0IJOBXwOXd8L+nvj6Scf6+P/bd2pPLyibK9TvhFFmWwQ
qFI6RwHnoRCbKFYvX+TSmrIT2aZkDrrAhGi2rtVl9MHLC6nQgC3zjnZ2wwnp9Gog8+qp5eFtN2A7
kcHu6oLj372Gnax4meEh/v17TMmlTOYfPER56rXPNcskh7SdtTTFft7w2sOAsr0Caj166S+1wbVg
i0YWlu5ah2wLBmxhkBeEPbP8R3MCdKIKVanXTkXZmYNn0ZIAOpZE9YyOFNINllBMae1uHqwucSDf
d0g1z7CJswfGKR5/f95FkAuxUNZy3w55hgd2vihO6EEUVwCS2migY2UQB82l5x1eSW5dhagaXdrb
DxhZoqxcE4Z7z/HPCHgJbsXwdngJKfyxOV7SDXcTyQmZCneMwsO3+d+XDBPO3NdabH+SW7wUdkQW
yjMTECM0W6dek5Dz5LF9FMyhdr/8xzGFf04DXrp1HvG1joAyJhFpsscyzrUGFhrdYPbPxrB1PS4c
gljdGTfk04W2t4tUoFuhdYRGXkoeHEPnzFzs75FU+ap3Dy3iLqWzS+xWONy6BdzbrEvL/nyy7x+s
MaHsYKaJamHDyl9YuKD1DKtbFp++nzCpUm8Pa79zgeO2wLymjF4/gR5SeDltaflpcInSGHCux2bJ
QJrjkpOIsVUIR7jwx6wKKkgbqdqE8hdTnm8mHedr21jt+ijlsZXG7KScRfQe/+XZN3uyVW6I0+rQ
OcGdnRdK0H6Hwvgs4E81fnjLjAB3lU4+oK5RkYu3esHOtLDKAWtjYWz5Rbz7+9rqjyDeztg9gFBC
g1x7YmQ+ne5ISR5EHHzFm8QVu3CYuFZaYlx5HExwX769Qe0kncuytpEMuOMo11Q1MaTdHjBO6axd
assEP8HYB9LWu8EO8WQfkawRE8e7KgilHfXKADvLXRTXRUb49REKCLqvtyrhMjrQvvDiIC1keeTS
XjuA+e/S+Ax4zWMibHMaIkK2/qSqvlO91iVDEocQoX+ULxINrigK5mLUfNaJBwgxBL+PR4P6N78B
KVBKr6MTWRzvTUgFaW2EdwwnXK7sS/IdMOh3WonUWrfLcy93WAaDXLJXb7vhTgReYvVh9LR/v2Qv
HMvSlRJcdIkPuPsljRf1oopGMmr7C0LZnI4fmHWS1WsItpq6vwWcMDwMD8vi8nAQosTQsJL0ZLCB
gDJuXtBKKxTj9ivPCrsc6aifNOcoweKMAHkUn3w15VpwUo3LQ1MWkzYpP0rHGqmxHCE72Qsa4Otp
aQJXpqVL/RRaPYXTQunf3rADPrMvaa01uX8qvvJuLlAMBZQi5I/dR/u7tvpfWGTLzp9EQ20PEo+d
vR42m1tVMz7GpgXVewU8drLqeVUyRSQrCt8Ap6YhigHTvafGmU+3M+x9RyAFJNUFNPsRA4jQLrVm
uHNF5AgexbjBjhYFwuPbbWL6Cy6drk33v47cdmTFlqur6cCqFcuzlj0BVQQOOIutkaFcqLZSEvG/
xAknEO2dRIQUbHeSbm9f6e2VvV+FQKSuXPaUlclrTGiTi5+x27SEDuyWV72d3XCQFzgg6e1tHGOP
uQpObtLAUlKtcGBnKyxXawPFpaP66+fBY/7+BzcCtmWzpvbKrr3nk6N8cm4ylU/AfvuxhAe6zg5b
8urCX6oFpRy2W6HEbJFKKcegPOIcOgovinKsljc8goedgqnuBrG7DL/18OA28hvgJ29xCkiugMta
EhO5xChHSH972+/GlK1TMdK4XfGtBlmW8k0ghzPqX7tuvLtUUoaRuNPDR558+/CFyFsn3diCWiwy
9c/CzuZucQSUVrxlRbY/U6Ai/tvtFg1q7i5LJEsGUlnGyiPnXEoul7jrg3LY5I1tU9oMoP/pgJsp
eEJwfeZF7TITXFhQYzZqwnxH9zCR6G/I9mTcvouDa1w3ikCJzq61GzoqBCGgdChY2h7hG7qJJIHD
KlTb8Q6X9KSIFvhwFv6Iq8ePjJ4Relyp3ehX+yxHlibmj4Tw6xsKmOCuiai9u7ufe7HKWdQ5jOfK
xn/+eycSvnrOMi3sSNNrRI6deN4ErQR1HD5KYzB8HK0oAc/litBjz6O92lX00294WNAbxuaU7Z92
o3+1pUFbC0x+eLJl4seXKGTkKaaCB23ykiph6rSA0y7xeSk4AlzqRfWFZ+UtAsu0iFe6nv6Yjs0R
OfkeQ8DQt/Eev82V28OdngxqNrbReBiguVcRciYzTc6yBjyV1OZCSWnnPskCP5UlXMXkdVOuWgN+
EPqOUQDHXEpA3NHuusNMOcDVqScDzDjVDOQlRn92j8WFlAgiXOC3/zSShfJ/81jZM88yFOBGMwP/
pKtfFy3nSanj9uG7RU1Flw427BAn9RikiTS+4G8XZzE0Q7RYwVZTWxyZy0f/qjPRPMDijWmzh0On
HU6R+x2AwPvVwDw125jYWZOKUrvPrx7i9vVCm9atA+AdUjo0kl+3QolD/CY3CwcexswIaMrurXGb
/pOtGIcWQHlRf0xFtjwSiMXhoAGqEUvfe11hX97EkltQx7SsOXAZzPemNpvpVQujOrYP8hO8aJqK
+5xI09a8ATY7vEuf7VXjZEbSv4yuJUcsWlrfKh2Bh9mw8uZDULxOpywATi/X+8PMeNP1wxNuLNmS
YPXHpkHOzNRhpy0Av9Xpg86qRrZkdYB8t62k5OaGzxIuBwCRzRzGmHN2XtY3pXQiOmDj+ujYUmCT
05AYtHnOydOtZJ/MKHDRd3UFFDK5IHIMZcIc+W7ek/cDWw+OSh2XJIuj3OjZqT8DYPbi8fIGVEDS
U+tcCdi1JqtYeNv6pE3zLLWG9EUGicDrgdAcnqb5heeAnuxJDmITg0xQWIe6XxPzg3e4rRJ4c6vx
541/5VG1g6RhWGxbVQs4blPdA5keCmd/pZWyVTRTiolJrWjNZI+5q52RDgHWyliQv8aqNhShh0MT
M6i2hwBXTDnItSvqGD6tBZhCTquuNM3GLgNgy7RMpji4ctuvy77mfcEvfaecZ45ZUD8y/W7H8eBW
JzNzxvp0znoLp60RWiiYMkwqMet2BrPp5nKb94Nsgd+XVpFwyLr9S9arbpBnhoTUlyQ4hfdbYNLV
jvwfQ6otaoq/Gv0I+VbCWiGKwxMS8571W2ycfkPDeFrL84H/p25AAoy6WG/Zo2/JqfDy7lgsLWwh
B26MomHyHvBQOpczlTuinG/ajVeaOz8zMvpUnyw4xmsSl+90b7s/ZtGQt4n2Sqi8uzINOTKbTpBG
fq5+e7x/nf4xAwXxGWz0ks50hsQNt1cBWJkLuJJQJ/eCWZw7t9vMuA6lXC9Ymz+W0ISSIlte6I0h
eIdbjlxsNqN1C/QnKOysavcrmhB7j0gedTx4mm68XZkx9DKFDSZpxJmaxT2bx84HPYEZ7oW0e+yK
Q1FYvCZBoxPA3kvcuZ2vlqeneOCBNw1t/lIJoSXYQLUaGf+bgFgRrjoK0B2hZ2vNfLJFVfJWzR8m
bGGyceDDxZQ3ksjdFWhHwacoch2MTt0XRUJyHamRsdanAjd/RW9VqfGQNiREQiETIDXz+ISurPV8
86rRoHRwecpnzRpJnsjiUhDyp5Nz2QzZeEYHv2mT7tvPZPcTju648zgI2flCB62Yh55NKVQ03Gjz
thzvWx7a1v3qYepVTKuEOF3Wi8rGFSSFhmfNiZ4qqvb//UtcZCuSSX0IG2bBbhffcTf1NELw+EOd
yjMAj1M8aKITR3UoEZJlZ32M0ZTwGl+7BvrbOvLH7l0l9IWJ/v3DujcD5g0oT/tsGeQmEcXqUm2G
Gv7aStlw3yJwQbCxFwThIDvJMRZj2+iiQjw3ICCwdQ9820+oA5Lil7vI27mPOpj7s2eq2r9OfTO5
PP1NwRQAGdKiCWti61jF5vctIcnwnxN+Pd2McPFZRubQ0QPOOWarA+HZzzbrHuZ1ysh+54KF7cib
9dTiqKkH0LZrT3ZhUl+/nZiUxK4sKy4gtu1cyUJw2khZkSXRnPv5e63S85bu1fB4q7bYcsqyqwLe
tcLc9NY/UUA6BTOy2m+T9izDXYnBb4HKa22KUQWR7kdABDERg2PFGVZVTyvSYDC3pfbJMJDwXbKg
yyKRzJH9Jpx/T9f/TQWUoC8G1upfJZdSbxwNUTCzKE8Qnf1LuICghNg/5MPkjgLAkWm4MOC1KaBB
DYKfVWZID3EOSQdxsUq1xvXoYvaZQXKrKKdGqyPMjEwuF9t329DpDEjYMYChbFfz/nQT7Eyu/kyJ
q6FBwB3v9X2GoHv1jMgieGzyyjTUdy1zdu57u0t1oNr3gkhcNPytL1iLuirR/80+F3aYWHFWbSaK
FMR2fet71H6yYRdxYHmf0NF3OdLr97hQoIG6MGruD4stqFTFmJKcEHy0A7/6PABdVsOnJfsON354
KofRxi2vxt46AtCjir6ZFQdPZHLVN+Q+pKT9xua1plN7cTpjg36n7zUqCotygbpcCygz8YEcFhfh
09lsM09ZczfWjuFzKDwlSQCO8Gt0h1Ce/toJXkydfj8SbKn7wvgxONqKJdKHH+lEtB/pl190yEGX
wu9GJSGOYZWqRNdfAs8j+hwoV3WV4nZpBlhos+l5/mLUSUXjOkKftNE76bZ2FrTBcKu48HurTX4J
v28tn5tIgSnZMUmPPEmjNmffjM9kGZKiqCdFYuRwCC4RCNSDl/TWZ+rw+egIkPUrnN6ZNrzP8cw0
xOKG5oURQ0EZF+eMOrxKnk/XeBcLPytkcw7/HFtmB6urtgX8HCTvhhy1irBehd3Fpyy4oZ1nkdQM
6qWaa5TKdg2VzJtG6cURUVHOJexlK3h1PPINJh6an03Q1veUoMqFVYuseDOealZyhLbHYvQx0dIq
gdE5bynoVCuggkU5fU5WrB7Rq1206GMEn5uQFfgu9GfU1XSZJ3W00MEfCJ2oE6jsbbTnA5F/7DQC
MAOb+MAx1L9/2oTHm+DZi7vy4tS7/8eusly3LCQtXs55KfPJ6OLUIx4k+y/ovubXV59ZmQn6m/Uv
D1ATpz2r2iwsz6yemVCLLM1w2v4xZdwtAgXRRiAeQe7MjHwzUOEl5GpGdnnUH+QqwCozjJ6EAu/E
ICGj1Ish1GMu1owz9ktyEsYQBaRw7tLt7nOTW4BXHqsy7TsOiRD1Ap5C4cpfl4oq1gFoEjZcokyG
z+FBgozoS/pdJQu+jgTVBvg3ZJQQY4N3yC/5t8aC3AA68k4yJCD8TeKZG1PcFyZcG1egeq/DjNV6
8GO8qg1Ekk8ORXCJiVWw2IYjT2lwv9obfuFw+qccOKUhRdIwN7DvSbmInK4Vn6ieUfBYwbyEImMF
EdReklyViwyfeDSNvay73jHs5W9Z8Daync2DRcxDpBH309Xl7lbZyeaT15sOK4byRSwBtS2+IChu
qC/U0AAcHmgVr6Bu2YQ7ugDk1+Zhye2ZEdMpCwn/9nbnkyBLTC7IOpL8Fygh7enwJQyG+hpQCKBQ
eV5d/yLaKcwws6eZyqMkB/0mQb4kmE8olSapUwpeHuM42faejmbL8Y1T41MS0/YU5t42+7DVz/w0
TQP4TS0v940/ljPYnV7cA5aVEZkFGlyIbHxbrx/Xe/oxfTXWtIqZ2pp7sWEr23dyVoVHGya30ZNo
SxZlo/0vJUPulKPpvbVr5znbQuZc8KC47c8dHefkWzJN51QdGD9DcslGv+Pr59Rh59psqHXBOrHa
N13im+DBl0valnFaMbDyDndwz9Jo/BilwKZICcUHrvkdtMncq+ajFYbBzrjKrqA7xuj8yMhndspu
ksX11vNyzWe/gorjahNmDRd/gb3w8Nag2KTuhgKZb3qZX1QeQy+lXJln0DglVUfuvKEC+NDiXAjT
m53vaekTsVRPC5p4XXMTTAuRDqK2rh6+rMuGxVNH7aJG54dxPMy+y8C4sn07carMYL0T7Zna1dMt
7ALI1YeuW0pw4yTyD6YPHNydeXmC2+XUvbPixrl79SmRMXjqkPrq+7yKy3kiPumhWcxm4et/D1UW
w7udXkisJDo4vraiwQuooijUsSlqSMqPanz2upiTSGmBlbvsFj5KhpmdFvLif+uTt45Q0HimCBE9
dhtdPCgHzeNULb8e/MlKZMD+G6QD0lH5BZY5cEYJcJyoY3Zz624RCj9GVpUub9mTGF5CLP6iuPwJ
Pu6uVue33roMvhJYT0yLtiQHQdnr8oJOM5np0uBuBRACfrX2RfYRiL5Nr5+sb2zDHNQVKaNYpvO/
0HggxYTa5ncKFlDqZzzmQu29fr/LGyshbZVsAlIUJx+hGmGDv9+Wb0pPIPH9cEtld7ZtUw1aS7v4
AmgsXR2z5oe+PLR1h4elHHww3yIh1YHb7NtMc9V4Djma2kGW+8SzmSTiFNBwng0WmSRmJNaruv3q
QU6E3vObpY1DgWgBg4p7n+Fh1Ma9xu1sNBZhfNN+0BAbt7ywafI9x5CgPukBPUoHmMtn7hQfjqhg
5HuFsBmzdVyQVvTKvgGsHVE3dLaJfjOWSgP+zCDfNJhzjmvx2Ei/djtLAT88YsRK2BfRME7Idt2J
Ay7J5MxVgR4m2gYN1fsUU1f7O+EnRTFKCL7toQp1282AZJA5bMz1n27SHFm5J8ksljNPGgZPd1nG
h2sTgZeIuZft3JFYM0MLtDSb97canPXTIFYPHoUiiZ3WIFDaoP9ZDxPSlgrUgtpaa8RTzAF4eq6v
WxtzNydTM5W+M49DeytyGaqaq7IA73+aEde1FVQPyGVcLCTZU1wlWJqrz/6TfjuexI6w5e7k0J0Z
Y8F8g2i4qGVqLO0n0haRuZV1ivooYxvzzcUM2eth8cbNhQ0TO+gv+nqY0CN6eQ/nstONxPg/+WP7
boPw757KAUGCofkb6iSU0cuw2uBbp1OCu/Jj6KUOdGhTBv1uw8XK3Of2qfKNokJNxXEtmG60A9Sq
q61hzbG7++7mifgQgSuMdScQ+7VGH0wdM44tG4R1TXDvSULBSAXn+znFxLgZ/FFZyazV4hFUqHnn
0mX/RN1lBOStumW36DXMX9F+ucmL039rBjhky1F9yy/LOlaAmtWY/pV2bVP58KFO+q2rWoT9IEGG
WSij1aMHpZzqRhp3J4+pFPd7/wtwzyilq+Qwp3raWNem+Fycesw9KzFqohS1H3/FATIKIiOrZn/3
BbgC0dy+1gpkybZxGlP1lmXD5y5OcJm7tiGhCUW96kNy9Usdba6o+6waTTg5e/SFUxwKFUk0LKUW
urp4OcVRLZqfipDjaDBMgL0coowaWX48TM/nzHjDqNiUeCLnaqG69L7J+1JNSshLTvnfmgrguXD4
VxzqCs1f7ghcoM220g/8GhBA1dI9CTGDb6/7oTkvueknC3sOF9JVmbRt5VYIcnwUXLUKaPFonM5d
dpAStGqmh1GCR4qjupTnwBYld4aL8ItTV0buyuk2m244GYHqX5dkLmGXMWlr1J8zW8HnDFMFKuLx
yFX5pm9TcvGsNpBuH3RuYLoooXa+IxoWV0qfPchevuw/CIvvlHGNFttmYd9TheQRQP6n3+iH+qAJ
bpPBV9M/oZ0LoX91Kid9/J+2GeCaY0fnOxBJ86IeA31NZ6XKo0XePsi79wKx4Iw35FOefRrwzvvT
jcz2Q6b4BHMz5PYcPcnD+/X8Pb7a5ezgEMp7APUFNGE65Zbtyl80HpipkjJp9r+xRdTmI9/Yf+FT
ZH5ymKH/07Wk2mG3ojEuxRLDMz3knqFNFp8/ul2wlUDiCInk8KxvD71q7r1EakhYhuBGTgKNbYZH
dXnelfD1YmZo/ldmV3N7vRO1bDIZHcFpgIq1zz2WWByXijIagyK+GtW8AtS/UHnsmcgkHqsf1i/7
rclL1D0Psh7IEpYyxXENHp12zCuke6nVBIVwtaYfXy8lZTCJKx/UO8wJVpXOGEgw5TwKrjq26xL4
Pzyk6FKmUQyKwZxvq6oTlCXwrGsGP4CGMGpGuIg8i4x4cZq3UeaaxOpWN6XoRk4hcUUZLNvgTzf1
yteKfTn4dJc7STff75b49xm2bWalw72mJUn8wxOt9weM5HiiHf4pPBVimllkBaaLU5fH/apejKrA
Mgj7WfpSnU6lJyTxpiVnlu4M1GWwCGEZIwSAWHwRzyuwI8+PrBS6+eR82e3EfGB8f7MAdpFXm6xd
0RqN7uxIJ8uXt5AvaWMH6riOw9l6U99Opn9lLiPHL/hk/JyBgX9WR1hgeo+P13PVUvk5Fqz23zJG
QjJH315Ks912zulYASDIVMFKVVyXa2Dd1WG1rZ7/CTXeShkW5wA0wNxQEXRpB8t7iRnEcSOuKIRU
Ge68XfkQ7ydbmNfMzpRd9KpKyqPMu2fworNL1zYVgCSg7hXgUJsB65fjuFgCHF21F1WPWdmLK5wI
24esYHobxTfsVUySv8Ho6iOIQspLBz2ujhvwNizM7Kp5DQuDEp48pb7vX45Av1bPxzmrvCAunBdV
o/Xov9eniZ7N+pdZfySAY/it4POw0dgdLOqk19f41UFezGDlv2BtW4jZAfg71cLOA88xAN2V+uPa
xIcEkK3ztVofoOMan51s9GXHO8M0ah0hRVQrOke2LbcQ/6r736qpWfzhxF873YVaZF3BnThiy8+W
ZxiFbzyO82/cRgfgkXTF12qLJLjrGc+ZNmp5iVuB/2qzfghmSxKlj0U58bU7922ip2pG1SCEw8bd
zlE9VsDYUHQhFLZbBVdbogQ7DK6GcyD0uiG4OgH0wdEIFf6UrwGZ5RNOa2uanapDWB+Vt2uZnHcz
HOtqxDv8lfDdPTpYbovNbzMkwo90uzpGJSDImzEnkvDHOJwZzSFRHtqmO6jF+srRrzeaSV7ZGL5W
pFpENzMyPZW7ioDO088s8ThUPvxCndhKOW3sF3hV+gErAyMXiLaDOyHIogPq109a1aD+brQemtE0
Ln5ucGPQgi9l3FRflmZh4JMuiV93Bn8jJJFyXwixvnwXRciVYCRCtC4I9QFCRKfw275Mes+PW9UP
tRrapjbgS84d7+HS3alFSYpKEBsKCnB4X0hfqenLbe6LqiV4oKTqIP8HUyxGodRm7Doqp62ywHmz
o6aWLkTV+jhFxg0vvzRIRrTuXdTCe5O+JocqIuAAtbhRKKAcyJrjNAYBn5LspzNrwTBDNqfQt7Ev
NTcZGwr9Sj4wmNbp9SWBVDK/B6OoZX0OCS0Z4mKADXtYNtBtm3JGASvmYbGdxsD1UE4yHfj1eA91
S7fiZu8hDi+bB+Q4su3x/6ew5q3HQ+4Q5L9JyJqPJMNULOZFGWv1RY6tFl+B2KVpiISGxWGyHjx4
ZabL/5z0irzEknRLpI4ifv7Rwj9Y/7h03U3c0n77oFM9wAtNKKGKOy9kasENIMAe0Ta1lijgwxF7
ylyBqpn20wrUPbIHst2DjamTq6hgwwq6CNgiPzk4V5SJMBkCca7xe7pC1ww7VqXRLg7Aly8x2SQx
N+e2HVZHAGqpQROE7JLMEQItzrZ4HHq8dS6kZFSTmdp4YPPErIqo5Hs+16PnoHY3DJwcNHev56RJ
oEuKsga/mJIDWCNHPiwwAETPKSLBqsSXhePHGRzCOnwG3xW4BCwtSxQPvudnjxPTc49WBjJmtcpy
1+aIs93i2Zf6PWRiH7bp9dahc4wFtUHOc1QZBjKDCNt6RF8n7ODjx36e6XwDURhrIKnuGkQJNelL
Xv0SCeAjwfJCSFqXWXu3jIi+bcSLlNXIC38mMUfaoprR2EzJM1DqAeovvYPO4hwKkPbE3zjGczST
kQmcFXCW55IhMv3g/Bn4TKSB/uz24tnVU7Sw4md9G5Cs4BJwfgl5FFR8ecz6yrgOwtafDclGZL2O
oDMiH1fQo2pGRRX47IwI5JgQ/JiGyfuaKSTdoTuPVSF2uldtNrik6JjCbbsI0NPT7kMPe/34cMTW
bD52/kbsT/nFq5sAwsuDwPVwq2h8R18LMHli1OU2Z65j+RJzvKy3817uTius4PobkIc2/KllZrKQ
AYOhyHqtnVPcKXxk4eEb9kBSm0cln0JYutJ78Z6oVvbDEGnDDzparIC9Ti69OZpthHOMP/lSRNW+
kguROM9ZIPAJ9gImyApzJS1IGNQt1oCo1QRL5j15wuyzL6X8gCutJC4noxLqr6kaJG5fx5xYJ54X
UPDmJB7qZDzcyaI5fDG9WLPTm8xwt65xeD4fqvNXSyfs8DHGt0gBDIux3Olm5lk7HVpX/Me1pwYY
cFIPWcJI9qpHKJTSOXztlJOfpTcjUtz8GolmwJC/yn8TKJ0VGSTXe3MGdPnig0u+YwvDzS9Bd5Xz
yOOGfCteRNxf8+81fFt0hkNsxiCn/aEpGl3sTdcJRsVzvsJrG1sceLdTjH6OJ4ZIeYqcVsi4jOTV
OLd10kyjVLvCyDyysWZ9cpuMu8/4bikXcGaH7xEpmmHFwW0FES8chL/xOeBpayL2CTpFcEGmLnP7
jYcl86bjvn1nVcVANqpkEe9Jyo43QKKVj9L+pqKDBGACbJyuia87mwJ3R31hWvAie7A2PCqd/wBn
/yJnHKykYpg2vKptCst1rhzxmOQBrS6MzRYbW+7yaKEUhEN+jQ4kSOEetxmyO7NfakTc3nsEl+g0
BvlVYZTwMpYlcdRhW9jusb2yEHnXNhuRs4aS4ZY02tW4g7zEzPYzcjl8hkRbxHDgO18F3+KULRvB
S8n1aTVtDsGHga1c8hu8iWbpKtpS01cwX2ky98+WEvo4uRyLUcsmrIKQA8WmvXU/19qtbYnNikZB
UkuSYJs1kqTbtct5J3cYhiYenuIrsDVabQouyTq4KP2w8ZJcB00ff9B8B/f1pV/VjTXVI3wGJVnP
/VCLqj0CESMEqwvD56FCQnsZSzWMPklsXC1Xrxnu5ph+mweTWkhQjm3GvSN2T+ul2o1iYcHtE8L7
NQIa67Ei7FRJ0nT9/lVdr9MHCzmNDzQX043xxjuN7uXePF+Ejbtz1As4ErOR3mUW14ZOmdzUfUhd
hU+DqLlROOg3NUBNHRZ+woSiGNrgO4RYwWSL21SerFTmGLiMYTMm9urj0HO6BMZErfKU4VZ/kodb
pkeMFPunjEhnv2VgdLkQnMtgKWI0MtqTN9CdwwXmzb7dc36WHmy/dMJtwTe+iyl5HyuoIrSFBf5u
EHZonrhPw30DCM0HbZzwg2kFqX+05wBgoeBaW1AWTgbgacPv8c/rf7rvL4TDf+VmfD8Yw3p8bTBz
TA+XYfPcZ0QvgZTg2wYmgxlGWJJZOPZf0fw6NPIZJD2T7DyWvNFUnb0pXZNQ+AGc7WeegGPO0RNh
sXMRP76lNsZdlv9CjA92q0FOnvFYbFr+TGaDl/5CoTTfmc8JKvMhBlTi5sI27hj3hkP36m5n0r3k
ioLCU9AfF/V9UtfXVeJ5OnfQQ+k3LO+uheKVzj4Ens0C8Ezlo0/1lPpcGAgTzgPwUZCESwEptacd
/MH9AaUpy4OI+11GgTlBXPFkePoz9l1tk8HNRC1WJnfJ9i37X81djcf+noxsJ16yui3btHQQYHx+
CLiSOIrGouFNVyMRGpWg+KDgkd1fL3y/8ttuv6c2Lj7Iu9wWZrjj04QcgL3XYz3b/j0y/NNhHYMJ
+WniHNOFUizyoYXqO/tN1q5cLKYN/FORTinOV8BWBZxokKjEwrfBpjGckYD9V2ofjapHPXkTyhiL
dFigMGtHkYVUj4TRqtlhEg1TnkD/PcoSDFwNyAfUQL6Dw5ShG0nEkt/nYqgcTneW8CxVMLaBXVPH
gUjJ9Ntg8aqlaxWhP6yj79N84xJuWIw/uIOPCRDYv3v4hTqHZ/Wg8/dCteTbNXJ3F1Ogv9cxH5OK
mlS/Rg+Ov20dGyBXKEjuBrbt5Wwp2gsxMQ6zEKnU6e0vyObif7BxnJ/Xzkl8yNfcZMGcX0sAPJE2
S1D8GQ3fNfje6BtceyslZXwd2iDZny9LHYV8nLQ5p2VV4/coie8o48+TGBtbCX1/NxJqZmP41elg
aQ962Y9DbB+M8x3AdnGwBl/Y4ZVYyUQD6j5pKoeCAnuTKcVB0ypV3FZiY3sXUqg8CzHWaNe0WF2B
nN/+e0R7PvEAXn1GtukEgaQXwMj4UJwT0hoSMqZTzP3c4vx96WZCOigXDwclrfG7udKor8ojv46D
Eh1g4u7509Fmu2upSgqVYZug4g08g08T6O2k46HIyK3w62/uRdLEZ7bYDjjknVdpUvR0igYlriOI
5NE9s8XXscxCGNSboYoXq1qwL3ZqzFFk5tYi3rfI2xoWfC24O1EWCA/jYMlGQFd7iKemQmAzkatP
aPymSVUPLGUyCfNI9qfTrr6xesVW/qb/cLGdwhDJB5uD26wvc+8a6H/iv3lIfU7u9T6iqQ+UL/8I
CvSN3gpFdgNrO7zIlb7UokZCXeq7Ft0f7TGkbwTkvzKgZZ1f+vpx6hvx6XxLZnTKAyDgR64K5Zx+
8sWpVWNmFaf48taPXflf30BCw6ygDE4d5NyOZz1eCeSZTMen80pILkfP634eBNWFhlwODwQz3mU4
kiMn6pxwlP4OOoySdHbttU7UmghzAVsi5jV195PXbZTQMjuxBmCgL3srNgaknxkIp+gSsjyRIibk
D89ORL0RI0pw6ibcDWebrQE/H1wHQehKLck3eLLR6t0fGRCfk1DIr6TA97HfW+NlZ2nfI9h/JkLA
lkl3ljU+wSL52dedoUkB7DFW+RLcIydkc9dKrna5XrUu/Z/849vOUQzS1NxveVZHrpNf90ZCiCXp
qyRUMEJV6jrxbHiFromIwgPltfUP2EqZaYkKhy0UdswTq1+vSAYNGTucql8gvMZXKIMacZkoDXsk
geE8eGDbRWL/yC4qYITbDMWvOL9gvxXtcfBYHIpUmUOz1VuXM8Fc1X8Mqpql1Np3MceyRYINwKKQ
wfHFrN7XfQPiM/G5wiLA2KZaOcbHGjhaV2OvWeidkHfJZEq9SmctWweS8jOVMk3OijIsSpNzFkWa
NQcAiQLlnqUSYehxBz+VPlqVz3nCb5jHjrW7brtLbH9kaq/CPsNH5tIGDUqVKq/ScPUbO/EJ+qwO
U5RNsJzTNbVOVS9Zbs0uw9Run3/p6uQr4t2G0UJ+Y57KrBwGooRdshyYbCZymnb40KkgdVTy+/SH
cPzxUD5afotZJbzhjvMtiZxs9lt0xMlnjzPbknMY9aLED6f8xSlUMAV08Sl2HMQAj86hBNPMcPpA
8c4lhCgcsp/huBCv6F/iBQrsh/OD6UP5NEXPb5ji527RHSsADWjF9+smGIL5YbA+cz1l1G8hwTVN
O5g44Q0hpiSZa0wVhH4CpK3hC24Uc/XwBljRkaj5YlxNSvNcz48ru1q+RWs36cKfMPZ0zeepTd6v
M5kY2p5D8uVUpSVRMuKfXo70e6+ML/Cyo+Oj95v9RMBkIFq54aPvlnC5NmxRBzFw36GoaCJOMSJ4
umd+2l1z9Vz9Gbe6K7WCwKV/MDMyhsy4tYugV4McrIqesehqRDuIem/HP5FwaDUSm3hacNhEKcNw
wC6d0NOBfaKvdnHIOWLHNLsfira3/sipJP3QnnWk2Om1j+AlKpklX4OGc80+AfdN/AP8WiMljm2A
e7E4zKzHZP2RrJjliK87/dzKPeWThMDCvxAxZ6vO+uwahGopsp3pnxMkKaBvxJBMMgCs99+I9p+0
4o5IejBWm7GZg5pa4BoVPD24Lwl1NVdAB44saQx7t8t+KYyaI6gsdAFD7YeLSUrdrIalcT7FT0eW
d707Px5gpZ0zF+gfaKui36CBBK4BrluJ4JJPR5LFh/wAl8bR6EOfUUTq61TnWJGKhrIWTfrPjsqA
ggSXGym+wo0XRbPI4EkE32vmTJgyo9nrfbz/r3z5gasOmiISnAhHTZMx9d2YL1dq+orsZ6o2Xext
jo5aAc3ZGwmSbDbwIbB5dPZIJPAL82fYs+PaaASVL71s3jsj6FWLaHR42Hw+gYlDYcG0PLjbHkbQ
qqBQ3AhLMq4fVx6LCljbxGMQxQk8yopP7vaS6DX/OlJvJ0xlIWY2G2YhrXNaMyH9FHuuOIrMjfcF
piS+0yO39y+6hDFG2oYpJeNNRMTLeAX9uEYXPZ3pyIemFZpINE+hj2wdeyqhn88ZfLwtx3niYUZq
NiePK1RhYWQxdzgOWuZ70D9cNYBkoRI4w6i+buZtvi0AK6r/C+YvcgkPWaKS/SzYPjCM39tKAdL+
V70Txri3Tl6CkeoJwfQqmshX6RAkGxoLE3NaOA0MfLCq+/HXApf7WpNyoTWJIAMOWxA8GOujy4fZ
sAC2CcIPdVd6exts+b+pUcVe9ZyLcnoVGBx/MbSD9Rr55x4MGECwJ+J2B64+H/Vs4XypWNOZSJOL
jok32Y2mlXIhhEJXjuY8AzVMr6O3/o0wrw5Ya75srMAoOmrvixV6BeahNBlUM/DyCVfX3NtceXUm
LheOrF0cagPAhfaXIRcX5qMCfkzVpHtbZ5tsF9AfDdgOP2LwPr+PGIZUtJnQbt0UKnlRSw2V05JA
JT2NpcF2oIx5HhkzpAlsCW870HlUzTsnyrkmOjl3QwmhXtYicd16mm78v2fwkXrW5wQJRHLOohmh
uktW/Sv5Um+Mp+no4t9IZtpztx405+GT5sHWZanAwtCCI6t1OWsxLIOVXJHhAT2xjyXRhoWSuMAp
HbSJBiLdKGMpqrdSfOBhiJSJm+5zh24+6nMvL+pyYZL0lHZlh/lG+7YF+EvC0Ily9yVdx4lO27pu
wt+1lCrojaQaG/sXEZpJxL5x8EGxPA+FrcsoycMpI6bqMhmFpoo1O6ipEZhzT2Z709KVeUEN2KsY
VusKbaFk3KtCKweF4AwweHhPLhCbLmC37JG3RCrOmqeQL6X3F/p/SSlI03kQcWMoEnJJdhoCqoc5
YR3A4A5nNPAKk0wto1QVX4EFDitjM/Pog2K6cCwyMG8OyNx2Uk5ArAtMce2hRT0+GXxsD9jsqjwN
X2oyDPuZk6lmmsWieaKyoQYg3olfbDddPd7La+ECO/uan0m9x8x32pb1c7mEUBU8vNmRsO0WeFDC
0jJ15cENHRaGx1mnBBLObjnArFECe1cCUD7L4Py+TRNEQavamNd3A7CTfibPOnrgZjFL92E5fFHW
A7PPT8VxB5XLz1/xlmUC79yv6j1yvoEqkW5li3VSUqkCYrje6PDMX6dGDZn7Xvp+HHMsFMxz+DZ6
prqhD4FLPrTVkj9988rea6g9FTtgD6fiZTbHYp331kwcqphLzVUG10D10xQHWDOYGBDV2dkjixI8
QHkZv3g1WnfDZ+DvGM35GAEtazF1fNboP/ZWbK5a0UaSObOUItNh3F8aRIJbTXR9rVyXCEiFqieN
LAtkINGyho7xVpQJbFL5o5t8u4hjWM2VGmynDy+3EMjwCwACoK5STsUuZLwU+3SJbjBxAVYIuYkC
z6HMio6fWPSZ2DybjE990zwgh6fZ7xeF2FIsc6EJ45gDg96kLXkwdgKJe2gwuUE/rMRAxf3++xmH
T0Bgqztl50c76JPTgVJCCkcOMDfOQO2uogRk4aWX30YqGYxwFE7S2utht2Pq1chi4PeFErT7rusS
UsuEhjck1AQHgIpYlKpjUYWAwAHNTG61J1Tv5TWGgvDPL09NMvnX7lZ4GAW5P4XQyDP1hBd+xASY
lfXNeemhBTF0itb6Xu+ODkDSrGcvX1tsPQKVMIqfN+oZ1/2unfCNIA5envaJCVgpNK+KC7bZRdeS
YnX/cgPSbI7MKvolaLHsbVomonM5H2iLTy6zVhx/QaBrtaZBL4IH1HR38wT7/v67n/mImaQm8JeJ
zin2e6HlY+wiDMWwAlH6pHjcpPD7zoRBOqhIkGWI9eHWbeN3LTXzln37zIPzJyuDj1ugP8Zsc3Wu
IxcINWotqeKJ/eMlzul3wPW4UW9guYZZGd+Y0DcQrMP5wBO/CGuF2Y6snBKRoLAuJkR7o58Ec5k+
cbvwlMaxRV5ii4K0M7EpSCt+hwcpmtuqYcgegXzCMAFbUgQ9QhONuXRgTZOa0cCySR7ZmgsHfngz
v+N2Vw8ZDMo0Q/2umuQr78bGKbnL11lun1kLN4PNUDcDhg2hNZGO02CExMMgBpKyZ/+QO5Htcm3Q
0c2zT7cmkU9BupOC3shu8xiVYW0iY8eWCYsyBDy+sbz7HdU53A/5raXMrDWwvGb7m4czGmsMxtYP
gG148sfcstmTweSqSFj99AIAQWoo6/V/h0RNgiYS+4qcg6Uwg7Dm3ZPEs8M8IdrWcMZ3Lvo5Cemt
1wkRO4NrkdLDMxImdvFOua7ScGRDy4U5a87WBcL0sKGlUz4Ki2LuxblYbojgOqAC6GDxuUg38/KA
u+BXvRlK8PYxAdK6mW9UhmB9VMZhRqEEpRmZXef7s/htgUPvUkOGqxphACfNRHekZMoeklHAf2u6
5WZsfpHQNQh5gRUUqveFJjPgYnvHs7wn81Xpw9L1GXbZ6b9bp/FjRco5wP1yoj5eXgzFgicp0ED0
HiuN6CYK98guP814SG3aqFIj+/6ovCx/8lXlKcjSslsx0S0DH0qXb8Znl/ubXGq8INeZ1mpBtquz
7MWTO4PVk4eGfOrTVpaWncmS1ucPe972SDaL7hVEqiAW5W2aSfiJZUflxK3/UGEYXp9onY5zXpUo
m4X2Y+CYhjGXVbFt7Qk89LOjigacZhXMFpMwk7vMp2s2nKrz0eolRj0V0w4qyXe+tkfrrcuaThcd
KRh+IHxPSgw7cuiEwunF7uGNlFpLCToZw5o8p0mgx1H40uhAgdVFasgh/WuVOT6SjoEjd0REAC5e
AQ/NLl+maSuo8SwPRrxKCFe8VqUfTE7dEAFQVakDr5N5LHmaK/NPTqZ6HR//d8VnDmPolwUiW4uW
I7xtvQa7ELICsDvK4ctWHYRvDy0CqpkXPUhRropc59WFtpuKlMUZaAp/KGCj14z7lYdg6sJgcd6e
j8EMRdXv8mnzj+dD2JFEguXMZlImXsv4bIfOkZuOXBwMuF10cq6uH1JA9k0tKiNV8l3uIjFb9Bd2
kw5n1ZemR2L17VNtF85EY3qbitSHOTu9mDlBFYgX/HOsH8/7JTQTkFK0c/aBEWEqdWtJrcCs6a/9
sHkNRmuDF9AbkmFifCUb4dkJPkDYIba3NqpoADkINXH5iLdy6pDRoGfGla6IItG1kZjMfKvwossX
kFVfX6riyEHwslinMZ8brJSg5QZ272Oo7IarbOV8wYoBgbFfZdTQbujWTgACWExzsxIU0NoKHUWf
031Rh1kgKII9tyi2ZG/Dwgg7q5zTqy8Exv9qTvdQTaw0z6jdGfBxMkRSG/LGg4MUeCgXnn8Hu08N
M4bB/nrCJqtA8K+ownrwroaGok/IMPgVVQEaoa3eb0uFtu9P4GKLCMHK/nAh1DqpSREPUBnVaV7s
9az6sWEmwd1OkS6HKEdEbP5phGxMhcRJ1oDvAQOr0ToSyqA/aYDLg1YALEQaVhWhYUXw3+87Xr7w
RmFHLsYIr0XltNiackFlTAm+9U0gW4IbjZJOpeyEwpE/KCr4AoKKq5z5IzM9eD9SQ/5o2RgyxzC/
phiftpyTzLc9Mp5HyM72HrMT/01mCDND9HlFmOMnvf5LPjcFNkCw6C97JdyYbEaBe07IJR2lhMpw
WvbcHX2rhMJZj92K3kNqizbbzeJgb5KTQ1gfnWo/rQ+1iAvNKmjnOkLUe2WrMUsmra0ewA6EVU+z
kpjpdzGKjCyO9HlkgMMFkfNMRZBrQKR1W9PQqIUoe6Z/dJM/W9otiEM1ppgA0F7L+AKPvYA0rQ0u
kFyRUIHjF+sSuUF/m3q9H9zGEZ4RM0nBwlflWn5UTyNK0kjBLkXpZoEJXRjhbyxle7lLpW2KTxJm
nCyP+Xx14yb+NFgIW9MfpYdKvKXGCw30Ll0p+xppsmkiaNFMvmvEJORD8t8LDj02b39J4VmjvYQZ
OO11LtY9j942ju7jMv7zx35ZFfq3DXzGVQFn3zBRQ46Gdbhu9z4sAJzYTBo8llzjx9CTW2wRHYCx
Y25Xhge+7lG/VsKVWVtp50smRD5hQspnzRAU11CRoPHvnOvAu3dF7lMlCqxI91HXFGAxymNC6pS+
BCcVZaXn5COijfl5Lqit3+hNhlxlZzAYzgmsBaifnH/pVlwuyvfdWvLh8GnUW+tDNj3bnWvcsPJW
zvWETE8JqBOpBW+rUJKlyiDBfVGcQMVooL7alIBChQk/R+drU7XYDnMrpIie8WD3vCwPd5nt/x3q
XUWNTnMzwJv3Xb2T8OeGut4V5q1lz82YX3Xr2MnOPh3Z63BOi45Kw/vpw2P6vU+kKttWvJxFyS/m
ICPyuMu39SK6nDd2cVNEpeB0TLyAe0TNIUqI3LZHRGD2lxAEt29H4nWTCDlb6bgOmpoa9aJec9u4
Mldj/GIZKBVZQA2wg8j8f9BN+N/MI+PBNKhwy2i4eQBLTNdTDfTi2NUKzsSCPcLrAOQi9PENJ0Uw
4pI2hxTNby6ghmsqGaGz8YaKk6312IJOmbeg3tI6OR0oQJoWCptvENPmsT6WW6UD/wGMWazr+wOF
YGe+QQRSl1FvT5W+3HpnT2OWLawKqegiWOHrvA39LC0tdqdxr1i/+oirL0Qg4Ep64n66GR+ZHVsU
LrMgnYG/PtJI7Ig8yHUT5RfXd1bw6RPm9JRU+LD/JacCNqD6B9lwb9JMg5SR9B5Y8KuFxRw5NDPj
h1Bp8xQkF5CykgUIOBLBht9iKzX0ofxURxJedje1TAGR8CGAAE6cXpNvWxnK9GtTG+qFERxTLz8z
KGqmafyw78By4KusAYRVMrv39B14EnAJaUTweRFkGtPG30ldwB94TpqzLKCpX7GX6Pr/eoG58e79
I6+uFW/klwMk63PCIeg5sIG45ETq0TvPdfCB2Hr4LY8Ih5ZjBllT0/zKqKK52wPBfMbHhgWJPp5u
qBluknCS0RLE/eqd7XAYK8IOViHA5FiLwNF9RyabvNLVcQZtcJVbieR2MMEZ7hiOCWpuv4UHqmHl
zSkOfOIEd2+VwztEDKnrDK7LlpYTe2qNDNRaZUqb6yW51oTxSm+WWxTOkVVd4KRZxxZ/VMyIfIZp
lz2z3lypB7KpUcj6PDsRLfcPup6Y1S/4AHgSpURBW+hW1lipPW7CD8a8BgNawO8Bal+FoyNkBgks
1ttoXJ6WgCDvjfw4DuR0e83W/sHMc6bSLgg9b7gGIOcRM1sM2/gIetnCOKAcTxyjKJtJ5uTtTwnf
Oevpu6THpkH8vh0DbGjLbZNRHNWypQ0us46KOnEK2Ow/zOrKkVT5xTlZXcqGzpH5Ta6yKTizfA57
YfiTVWAz5Q6g+4T1gbtOFBcCt2TzLrc2Q9gCg1neCdonREpZGOyhIeZof4jMctGeOSa5d9xqPkdO
vO+n+cgWxai/8DhltQt0h30sQbicarfSjeSoaiWvYyk+SdfBrW4R3RSJbpg1S+sfQlwYro030WHR
ePwE/ehV8KKmmJCTmBKjjLA4MT1NdILMAF9LXO5Gkjd9NVh2STRFGik+lfSvCceAhiboF/iH6i7z
cpVAxyw+QgVxVuBiP+K23XM1N/+fGrDcJ//HjxTBCwGt71px0ewmBJPrn4w9LxGKi2MsCFK0uHF3
9eWA2W6CLAe58rWv/DLkwlg0BLoO+CuXZLcd+G5mw19US6xLKO9FocrvQM2RfSmi1z+85MaNiWgP
q6xbHBoDAHGZ5YxKO2qTaGnS5X/yYjVQw60m60uRhv+lfw1ugRHR9zmCqwbta3waYKGfChBSJi+t
bCr8PRTNfjyHVOjEZ+DLPNOSejzms7AY19Bz3z9DQEgpAtwNANFkKzwP15U0B8+J/Aep/m9nMSSQ
c4JZBPN0knC2h7Ug2IdduOjzfHVsBos/TsmG8Wd2KkeoHhb9SN9jtWaplWeDNFLoRnU1r3oEHWo9
phHl6U0QB/KdlFpky7W0R+nIPFzALw5dx25n2Gbnbbu5BdiXPVxcLQsy+ZZlRT+33qslfDfL/M+E
QIWLPF6XglJ/zm/tlz4PywMhbv8z+d1B581uzd/Q3a8duRFrfBb5BpEZ7ps4xQFIZg09Rrv92SHT
Mimt0MHr4NT6855g+uz1lNhBkInGkde/gHqMVO1pJOB6FpORJj6mBRqqOjk8PdcNR3P8ljxSZrpB
G0Xqx8zr/ofX/nT/2zjvzcLu/Vcs3WsJKz3b1njINaalvL5/vpFeOPVLEGzT7g5ZCseYRzQfqZL+
E+6JNn4aqRbR9MCAFyBupEzsIL+5Yzno4NucKIqH0AHO8eNpjMDbUipxrFpNq7sNN3wFFXf9kxQg
896ML+E7pktM0wQ3Q8nQ73rJ3ATKjyo4JhP3SR+WgzmPehj20mCGhrwdeGg3FnzZd1dhC5pUK/mg
Lf93D2DZ6O4rrX3HQCpgNKLgsBus8gl8IEXEIOb1txG53eMGx9PjiaaPeXXoufnOJJdoOpbtZdGY
ZbxAvUDYlTDtfMqYXOBD1SSzkHz+eNkQsVZu4e2TxtqCI80fjhlQbPN0EYy+CVJtfug/Rp5ROud+
A+tcDP1kb4fZwbT9wBvpjGlmJeqTgUo1Euue4Js2NIxtcqrIUxrGjKo2bJffO3swct+WMaVAPwG0
EojdMH/6nrmqE/VcYzTAEDOjnGVRVNzeBfBM/2kM8oIo4rIeJC16Dtj3RrZ3uKzCgxJlpq89Aqtf
1mojj52ZtdTkMwDJF8H3AZ2G1Wk4nQWv3kkAP89pN0uAFHTajoH/Sggjst0+FN03q7ClYQyyk+nF
kd7K4SVZLhsIolqDlfYH7dh51c7aCUgAJxRfrh0ayhq9QPi9AhxndkrhPf8boZQ+wqidAtZfBnmG
6XPDYg1VCnmhNJqLbxqlMFCELGX2KhYj2Fa3JSnZHTqzepkuDeUUwDeziG6n+7nFkbD0THtl4kmh
EbFk6UaAlo0LgY1C94jxZLxSJJEM/w4lD55Tsf5FXcQje5FCmOeBwpnpEyexOwTafA2xoY9K0I16
bb99Zegk06VbhI9y/ZBryQv4K4lBTy2LTicZDMZeQB3QmDqxlRJpssVyk+A2srQ3/MLgJqMhN3fu
BttzxKP1GgE6VKhLGB/5hvFijq/VbutL9tbc5neE7VdY4th95ky81gSISZ2tSkCuZK7npFJgxX/P
YZ9ydubYRnlDg9YGKpQ3DzcPF8djebvmZD/Dc2cromgE6o2hIY8HA49/1D+Pd5fR0q5J0NAhHtRX
u9ODQ2Vjf25L5kr0RO6o8UnGV7hkjDzunEpUhnufDu3l5nwT/XbxtPqkpNgUAd4+Lgn4VqBwXcBM
dmJHqhtuSU3v9B9qeJJ8zHrX84AgJ8iNTHdLbPn3I7aFah4MFn9sGw4cBOYGkFVHLnxmpcjHp9UH
PkloN5FWKqvLo0qyJevoDsf38691GZ/Vs7vvKLTryj9Ndra2SuH3LPxrT3Oc4O2+H6j6eIoUhkJ7
hgHbPUzZP/9kThbuTvq8MIMv2JYN+xj0mV+HtJgNsGkS3EoSX6XJwjeU1pWFW0XgcGlFqca4hVfT
lGzQ8ksAg65qNwvEAK2zKkrMvIdHTO/z7svRVqCWxgBD19yjjPOEEBwrD0vBHNpAcNlnP/XyKXgp
HYWTZUPIO7yi/+SWS8MLvuLeIpu+6ki7bZSS+cRdjEqRez8SR04IkpzJbgLvw107Mx+LA7q5w79o
WPiVnD1eJgly3i9Lb56yVg8xYxJP72YVPwsgNbz57DTSvn1nfX0GgdJ3yoSeXyi8HjnRZ2QFJM3c
i+lSQzsfujto8tJvHKBIDsSjJzXADGpBE6MoppwaVjJdorEjyqkPKwrPaBZlgEE7ll7Fw4DB42Wp
aLazy9y4gkIR0wJG1VSdrN6cBtluuttnRkA9upZAbXzHo+86Ej+cO5+iGCDJ17HX7zhVn17SghkB
M+I6e2qN6DowTk7MLpmAqNikBQJeFkXdB7VjRGHZ7cr3f595hpxGhu4wpWDP1QYg/MeR7X2B/qOC
dGchkM19q6Sg0o2+SrkvWxEkrbGYkeGgOvzdrRvQyrmV/91hqlKTHlA6uvWXN+5SJnmQ5u+BEt7A
+B8TxYddKxq7ufk5u2yXh+QO1CmUVDORqF/uN8rDIwz0DK6bDqn0wNnfhGmUWwI1sOb9ADG9Urxv
E3cAQ8Ux+x6dUSrnMcezf/R78GwubBLKZNaphHZEBIdL6I6+VKneprfvZLagsFFLhoJOxZlqiB4z
qr31DaZpVS3pv/og5mWSEFed0p7zeiaOOE8ayVUaUx2UM/hgEc36JuOwTS2f8/jjxt+TE4WDj1bv
ciyWvAGBV8C5bpqW/BVtr70GD3XGFwcYPLQtncqxEIjF9HahTkdLtmT94Vjl9LCJ3Gf7bH1GLQiX
92v9KXLLC5HixQHBdR998IQbtgopDa16Pr/U+vFWxMsS8dfVZsGo1NSmpfaNs94YBRNbbMOKXn42
c/ac5EGfCReXlEUmtpQwila92odQZFLQfW8Xwd6uSpLInve8TxAoiAZcC48BItdum1Ghnii7Rb7Q
o4JcmtSlb4YrVXHSlUlNAlPujApulLOipED0dc/Rp6Dz8jy3CRsvVjsWSwoyBkvkU53m/ScO2Lmx
KXP2WRViB3k7wU48TSVFPtH/b1ng0Vxx2Y5JSTVYxG5auDKkvxsopkrIJLeVtakxH1Oi/eFVy5B7
XX4hAuwbWjn8r/Plj/01n0fF7oCtFmmgUDkMocJQq9VMsfp3sQB7cALWQbIQX/0JQf37xRoSjtwr
hEK7fUc7U8fz3K0AsUNsvvnBZ524ecK40vN+WhA1U9gpFjRBPF1sFQ3JeVDHIAl2oCpgziqBgB+v
7s6KVaDqm51yYtqxoUb2XsIp5MRsw8cceti24kiyO7KZWnRWM96wHOhXjUuITr2Tqg9Cg5YgMs6q
+hs5iAMM3okjUj3Lmfd4gIbpnQUFGTU9YAkQb86RLuM4fIsN+AFXveWiAMtu3xN01xbnrOZTIbbI
SA1Hh5JAeOeBa0yvpgACdAOhgecy7PWj+qo8H+FxCzmmWDzo9IKXrKD2G9ugbxaEYf3CzgYnCUkX
jNvL4qaK4ZHc3Cj65PssS1kiOZwbDTkMvQY3tsDUr2ycm8ZrZL04NVvTW3JoXNTX7IdhbW+HOYJf
y3leVEuEwJ26upImgd0oEmPX8VR3yv385koCuQddCpacuOv6Kr/xTVvuQ6m4kWviobeOaqtPfrGi
XGy3vIx46Z4Zk1mIpNPXcMr+6eAXDpCxcToI1xYqM6ZyHwBdpHXOPCnP+fhKCXcGfPkfBkvVY9i4
0LMt4rryQdL0m0QfO0G3DGmxLUJ7IQqI6BBzQHXR88KSJ92S1pPBL3cyOuI1hTh/THFSwBXXNzJR
LIQ4YI3yxXmR2Gs/8XQHAB0W/qct1NRci29O7J7fkjcpa72t6sZKjeIn3layOqdjZUrvausW2UCc
zx0UtzmC9UQQSYrCOu38FdLQQPhggso6drV+lcfiwHPdlQcDQ3reStXbFdVNdc9EMUWtyEIpdglF
eF6t7WvgB6Wi564G/5w1kGyUbZo9iYrp9M5MKGlWZ1xOSXk0lt8x/R7dI3rDwVuCOB1Kj37ZElRy
4jY7X4M39xLSqkM8lftM5fIQdW1RLwy7u3yJfNmM3TKKWaCj63bfR55z9z5U0bh4GqV+HNWQIjHd
xA4daQHimLf5QWGovPe2TkCMx7mviDS3oYc1zYg5PgUgcsfyp9aV0PqxQLET95ga4RHeX3Pq1QMl
aazPqn+3cM69ud9MrZbEdAqkE1OyOpH5td1+fRYfx0J6QWwqW8ihHoLnhpNlv2r54AqGGLyZ1grq
ml4bcE9mGMTWQFsaFOoDcUzbei3zbHBnVpcbrCroHHOJuCgehk9T9+GAMz2K+LPwoVsH+nxb+8nN
TyadmAq7F1Hgj3tfA9qetRKEvPodto8H7bSRz2fIScEsRAAaOhIw74txJjs3Djrrvv1Eyfx6CxLB
Zzkb43Jo7qW4WM5+GbbvSje2zOQNQTP0noThEjEeN3KAhRlG3GNTodMp57CAX/lpmk0+UwFF/OOe
UOdKHfJ4FKeJO8qyAeejWpKPy5l7mtyThWXiPiRuyDIvNbg4iqzY6XaI2kcFytp+WcbRXKkC3yu0
hS6EjqEM7p68ufCwr2hXaYovz3735g0MQye3CudfTjBkLIPjfNIa2Q53/KV405vbOFkrQpyGphpg
EoG4bY/Srb1nWLCd/WQHMb13epT+qNCI4lYbkN+9sMxngaG34Q1ZDMMCval9We/lT2A9HTixkgzJ
EdzKpySNvxPc3cnWdTF7BCug7xX7ptJb9BTCFl+sD55aqAk2X9pmHxSSWDL0j/naKtMngqmr8Ddw
bQMjoWp7dfNEyJTurL8AmHW+pParDOds5rYsz0oJd8V4c7lWHJRz+BI2LArEyz69+pPB4Q77zJJ7
ziXkE1NQAh9UgwWeItjkfYW1iwlTgXJcOfaeklN1YKNBY6y21jqbQKaz98PlYoSgb/yDnAEuueBt
lY/Lx0QRQaIvfRozX0TS/a/yJdcH6Bd2zjh3DWOH3VatbHwDzGAThHiK+XdBTM9OdvVGx16aeWew
J2e2WzqVg02KTTPDt1i6SNwQn/89b9g4EY2h/SFcHC2B7PeCZsmKefXvxW0e2kZPuhPJUh76LucV
eZw1E+U0KKWL4oNk41IZR27ewBV0lxW0jRozBm/XIZbBGr/BXP7mmGjhljqj1bG1wqq39jH4dWK5
5+qkmOPc9e6o0Cnx2ElUm+nfZ8KKGhaeizYVRqF9bqntbUp2n87/kb+IVdGKvu8f/50LsKZpbKpJ
Y+eDVv3OH/anpe0EfEQ/8PmNIvcUJYVL0X5INxQG3Q+/ozjCdRdRdPVp5k82fQwkm8+3fJRfONxw
J8GANndD9S5BuYzafgySsIP+ToXgjDBA8lhKponHOT/7rv1JjzAt3Qmbjn0S3Wytz6XVY+l0tKKf
eWpdp2LUI/DFwUyj8/QOKMLxlHmZVFFCSWIXpwLXX3g6IjGjO//NOrca2dKVjhUOOWqYhQqKAZJ4
Noil9EhKycpTXX5ckZp0uyzcbQu1KvYVRx4DH0EFMIhdtEJxJWfR/q1HP0OtZ1jVru8ETYIZjVNZ
Cps2KF7oOa4sQw+y0Ul8ZQomaHLvWhks0Pd3f/m/vPJMP2TzfAM5HeLsyFfV8qvTX9EtBRiyWJZl
V31SgTgS9TmY+V8iJztbIt8gVOQbV8ZAUBSVoBCCQrijyCgyafH53y7qJvKEyWmYgthYK74h311e
PUt+3UXbJ1KY3DWDuch7JikxlYqFw0SsDZZwAq27cocQIRS1paWsW3FEHLTdsGjyvy5+OqlqkDcT
8rkIo0J8SWYpzDAIL8hWGFbQumsZPB68jsUQmjTTVnvTUeJi5m6jrOf3dS09nfSXAmiXvmkf1oRc
XJWoxvB5u+wrq5U7a8bMAFFrKdJ5VeXb8i0kS5aHbSMZ2NvPPWFdrH2fVd5XKQqE0nXoGGs17fVD
VHCVyRX1FSwy4HDEnSbes0bI/me9PyZ8vB1QcwWwfP6BUUqzPMXC6GOH7S2U9Ruo/HWRvbqKAAek
hvHronfRxDGhvXkY3xlGDbT0FlHEORtRBrCbhFNZGR5yxEg+X+7I+P5dy73mGSX0Nd/DF85R2uNA
GU3NSI5WLEUg62VwMSJMSVGKA2usLTzUDxhc0d7sUFxcu7LJuakEvDL+IRro3fb0UU4OfI5scnqc
fip0aO5wOSgelio9wHzYUzBtl7oaNYAiVct1x0Mz/qTLEk1Gyi+oUIuQE9kYsNvII5znX0HVN/CU
mgOBdaNXocJMmTaAJsvnuCOVYOXexBFMf+m5TCVPh8/WgpQNPH0kl5IH1seXKrOW5hDxSE/VHSSJ
9N/CHNCCdpKrkgEysL7WwMb2/TKBX7J5Wd2+Pul1/JxfQLa1xT3bNnf66YF4BsZrPBQAAwWNsCT3
+bIN6fnEKdI+A2DudgbfSN/yBE3gr5+8EkvZUwp0zPYXVf7w3oQLCREjznFFMsfHWY0Uo0joyMCb
3udrzjS4ywm/LYIfgrtJw0GsG6d74lJrdxdzrvG61EA0xg9udbMwgaYXrou1px0hHnCKsTHsz7dL
qh6otJHtmui2D6hDg0Zw1z4fXjFzjdn2O2PotnaTYOX3gs1QFGeO06QMig+0rJahFAWAU5fw2X/S
nP5kZIZAG4NMkhx3HZys40Rj/RCOMd4QRBCrG3lw7DX24bjdwGgXItgPJQ9va1M8uuXBV9IgjJYJ
/M7fkX7DdkSKNwiGZSAY/sWcwgFB94opGbe5WdXEO73vQ9nHm6i2QoMGnxq5bFFspRjjM/6UUy6a
ggn2McKstVsMIMb7WxQ7KpPzjxHsx4cHlq8nSEDEvROMIkRQJyaxFM7tdMi6FSadtGvcYFJmHzXE
JoICM+npdSZsoyIKRzOKFccLxHdRb0yZgtCM0JEf2V2MlcNlRHQgAgdMLKihoRVViL3MZYSAjmm6
bheKC0PjX0E8VDr7+hS/5g6edGe/AHkifz1iM/SQXDr5CAQfjME3pcTwEsPcEM7ck4qrqSfwc2Tt
Yk6nlosziRTex6vXGNyKJcKaalBhkB5DsNv9Y/Z0W1ziErc4w9Rp7QeIbPaiOmYOuBqR3k7RIC9c
6L36EBVLQw4OhyOUFEjDht/0kt+oMv/Lv8Fp9ggH24fckmMNA1MlP/UHcyJxUCMbtZp8Ieb+hutH
79DCu28G8sArLP7kElJQmdO6yusgkWhkCeqT7EqI5TOBhKakNMNzNdPDixmGObGKjjX7csmBBFVI
GNqXguRni/3lJeXFZVJNGxD+G3ieEJ60leUGcl3RJjbhcPfjnvnyLwhsBzd6J4sVNfvgmsiln5Y+
htcUC1yyzzGfN1v8vK2z8+M/Mbzddei4yWXQ023HtdV913njitPTaviP23WSMbzd3CU1OpYWxMkr
1ye6nRfLaH0lmGGHhW9lSwz05frIqPg2SGKaWN/cKCInyIaPO/LaMK/n8VQheGvyVgzPTOraE5Sj
NlmUJ1ekdg+DrrqNYm9GliXv+D3tXpg21xy1EJquMLWYj4xg3th7xuQ7Zfze49aHbC/dIRalLCsk
zGXz/icL6RBvkQecXGAVQ/Tqqb0rjfoGqjhD8bu3B0BT9IMLHBTUtDYJVZ7Ek5Y1jHcUX2NVrxxf
K2z6HIyOanO/nq/hO/v8MiETEJ3x28iTkIYVrYgCgiUGPaShvbDKSdpPJEOuNbMmlZ0OaT7vfmUc
dDbA8O3oOOId1uQxY4+VxhWtJp19TYPwW46ofPBFB5xaXKhTI3DgPzo2FcsUu4FaZOOKDk879rjz
4CubMI0Fr82BKIOcv2x1uksCllMDVjN+BdExtKJVFpDkRy2TA/JkjQ4rQiMDPoitdCQD67EsXoD6
3qRqeOMvbqxEOLI+fKIVW0xkaV1o3EV0eSPCqPfqfC0FHxAWPjrt3w12evUc3FOpiHhFaEonIzwC
uk+Dwwa79UBTuHRUJ4yKz3G3MtUuRog10Jj9uxip+IQjAN5ymCJx9dIcTuLdlBlUjUKxO4r2v7+W
cAQXcloDkVRCva4ZzaLgjOGeNusnUt0vtAJCntjUwMEXkEIm+Pp/jXP91iTApeHkqJPpEsrvTPXm
uNspS5v0gZw7K9P3XY3Soff44T910NNqjBDNRKi7rJVhJS8+sgBqqzXaZKrFYELP4HnSNDSpXQPj
vSF0Co2yE6W+DvqNqUUuQJVr9UQ0gFsl9RcxlKqBWHz3LG5bMYWKscgTGuPyYXu8oZVSIEXoH6YP
p6kb0veA2twzmer/EwfwFtVYmfrFutLQD0GMe0hCR736IiUFYF2j7DMO3KX0SqyO5HxiW0WAiKY8
iXjsMBb3GesiVTM/2lBnyKvbGuIvLljtFdyB8Lhj0WDxmprF7DRCHH0czImalC7wNR+7OGwkYY0R
p4Q4AWxKABu+j1+cVXnv9fhxGHa/wQxp8FbHGOi6S2hN+OSnOaRCMvDCJs+WQgFxfVH9grNSBYzV
jWBi0z2VlRytQ7olssjBv6xo3B20tOboP+PqyNhAngdfx9AOZP7MBZPc5VkwjQg0A/MV2lO+ZOBl
e3NeqbQ/Sg+3mEm9IecDkp2OlYRTzHORcV/lE0WjWcuzlwRYvyFe5Hv33at2zctYqzt6MdoL7zJ4
i6+VypQlzdEPeC3ihC2m87rjJ94kkbidXeTirF/g1Auj5yIyCAepQg6FyBPqiqV/ZRIPQ1lbNap+
69yGKr9Hal51OQTz2Witm5UpHUNawT+8KB1f8hwev5bTVYO2kcTDoNkIe5d2ejOreeJnkH3ECyYH
YCTezwWh8YwLTmJb73F+zHCYtt8AQX6WIr6gg1ecBOWYcdx+TebV8tVKLJbUysGTGwf4E19/WbrI
SIJzWv7UKbO7/WOyzK3tcTePVWReY6+jD7VpBPJtSrSEJGteOoUiR9BZmGqXjliItUjIRMVo4ZtX
wKnFshsY6OG4iwKrBMTCST1T3zR2xuguO5m7iIZ8XkrmzWBuwl1D7Hxt1/efYIxC5Mk2x1YPIaQm
MIMSqJEGrHobyu/RwGuwKPoqxLNm9nY4FmpABMg+y4P1EIvO8WFsiF+idvFT2RYISLTBqRuspOzY
vSg7qqI43CtximQ8FW8DmTNksEWotDHjdH0SA+VsiIeJT2B+PxeAUlnUJAybjGip27mqrZT+qUS7
VjkKreSNEqHpp/AZGXf0d1RjibBd31KeKZNglr4Xk3HQNFim8IauhvNm3gYDooqRBUFN5MZI5p18
T1sid8AEhg2bFuabOwbOhBMXDLybqJNODNj3wgJUhsIWiSuH0eocuIg1PbMJLl6kVdY8WeaBJGlI
i6pLkOh2Gyj8JHk2BEgrf8vCR7LlhJVd5KBxeQq5je23b7scQLwW5iA1jeAIuABOkrkYdMvBpbeF
kFMu45mGPdFsDEl6pQGXyXJcDeGDiptv35hv1Jq4gw7S+/1niQhsEMoLvQwZ/CqGtXCsfQDZSuq4
6y2k0elWYfTtR3M9gNJz8obx+xvDgv7yujTJ44HU5EnsQPoo/7mQJGTABr6LPbthnleiTCozDRGK
aw1Bw4tSAfSvzxeaonsHKPeCnyy7gV1uzEI0Km9vJ54bY6ysbNjw+aNA6DECS+tzmhJcwXMTjzHl
Je882aPWx6R+TLucg/tmpIMGNsED4kVdb3XHEm4MJGqKPONKKryumnCS8h8bjHHFQ35s2FqZ1BP6
goAj9FRW966YCVjlbiu6QleXBI34rC0D6eILFQ6ITxoWX8sPnOqnDTHLaFFbyfeiCYQp6d/lRVtr
HnW9u+mWXegBPoRaGoldNeBjiscnpTGrjrVZ7ZZQZXqsQb9KdWXHGRV+Jr6LQXMPKEmlTnizBr25
WbN2WEVxVC/V/CdtrO3uW9FHm4BlqRHMuAwRhkJHNOb4opr8gY94JQyG02zG86frnQdfNWVfvnYt
0IEhP8pefk41s53qgRg2P2kLLs0MkMojNXfHPat0EzDKV+kI0nQprWt0Db7Uo9AJPbJgsIAzewpQ
aTLG9mtqoUJFteQrhYHzgoM+s/CtyfKiNftWb1zrYjy9oBJHO8866aTdGysr5O5gHxwnShQw9Q9x
MwlupRMAFL/knbhGXUxopeOdpJ9aIBTDLXyCqq//R+m+mpBBII7/YRqmYOA1grWlU7tRha9OD86u
lzUTzYspU4RoLGazVhl6PwaSiN6eE30gsQ0+JOH1TJgw1fMWBSKNg5By82RPJwE8XDtRNmrTkhvm
bMOwI7mc1PVhGrPzTAwnHTnDvhdzV/RmHsZZ9m7aSuMEBeRBW/EH4Wh1xifcBDZ8Xel2xwAw6hJ9
9CDFBkFkLYSzHGz/80e3lTaJDK+cuBlRxIUw8pqK9hRymTHovmyhqtq7ZpI9AHOoKdZbYvc1hI7A
CNqgZ7WBQfriOYKbsevr1qnlpu2bi1WEm3k/Ut0IaMD4f0BY0CDfmdbnWNkDzY6L/edUcmMdc3Ar
4mqdfqMOxUi+FleyZfZBFI2KPlDSspO6nWsYaRWmp7uWsXUAHDVWdD/UxXqKdUFbBUuR54FPxJTB
5iVOgX+TUHZvomopp4DR5svzoYn/dnyru7ESQY3lN6hKiwraiUVHWo3Ll4ig9N5maLMslAmKZEvc
/PRzNAhCoUdJqC7oER8yfZ8wMy1gPm9IwoKlJ9Em6ia+f22vHFJsZllK1ivIl6kLEq4yv3SFYv6j
XAlnaV9laS2BRM62ch7WL1AO4HPi8DURzRC6kmGZzLwj2Bdnufwnx95IW8pdTzZdMzh3rsj7g655
BKBemRXXwLy1p1go7Bt1iknPGSyVB4H3rr8jAhtlCM95WN7P5wMrNYG21g5hKFc3YPlVij/skZ2x
YjSwFZjBiIy5KZgDtCBiVflJiB6Jd0qsntRAWAfP4STCkOPO2Qk9Vnf9MJPcP6lB9UaugFJvjmJR
EI27AfT8Gp5vVPENME28Cg7GAP3FSnEMblIAQtEXFP6tLM/QxmlsVtVpR5xPkDfNb8fZ5t3z5u4D
mamkhhLg7ZhPU5yrLD4in7ePjc6936ussRLc9OhUEHZO7txWJDR9lm0rEwm/nf8KFger8pvKk3lj
ZkC1yO/8I2GoHONiSVmw5hB8UaCSUX17Gsu9AQVi+t6zwo1Dur60ciEHgeaZyXEiy6M4Z/kuQlEX
WIifHJRFhquik/WK8W6qv4uLYZlaXm6zfbarG4XSPkIJPsL5ERBFdx3bYN7Iuu2kiauOU1hba3T1
VlpsCtnNB6IH3PU3sgmZfJgnSUZEjbg2csLO7S8AUAhQ+DH0hhVj+3DMyqV7Klucfs/jAkDuFoED
CQOrZYs959pbcVgj1bGo3eRzQyrZNINAW2Tk+cWQEHPQW2PFj71csWDuOgOz8j7BnqhgxsxZT2dC
dck9NxNxBlI09JdH2K1PS/2zfTU/oTeL2oUPjAERijF1oB5Lb5OiCCc/UNgsfxvyfkn/Jzm7NrS4
KeLzanv7aE2FQHcC5t6pUNxurTEPvQA1L1ULzb4kQTtHairMgn1npCZNgY0A0TkvQj8qaKdCQyWO
1jywGWBPVR19RXwwkZhsRL6Vr20SdZeRyxRje5GDhxfgVymlLSLy9pyMARWbJZuyX605jcoqPmiJ
g7yEf+gaup9WDHRK7jl8hnOyPgOQcY2sA4Eyq1wjeGtRqavNEeMlYjsJC1xMWgrbJ2PWtEdRJ8dg
fwWFIOsIimr8Y4XahoVSG2ykoaIxr2LwtJhHIMO5cUh94PPkrPmXezGmFAzbzNGTVkuZB0OAJBDx
krKu9wE8/OJnGw5GLuznoUnSpXUl7L09Jk2sOspWeyy57O1+XAwZ5cWW4jzJy/+7h7AJoFVcUxRZ
cO3dKgTtpfS8e91P2sw+8dgek9NDr2tdFlYPSB5FUs7v7FzWXGu8l4sMlNE2fM7X2b1gpRU0zXYq
BD0mkmc7vZFJBxk2m4b9saPJLP7tubSravYQseN5xSFxL9vWQRjhkDWeFqNJr7vySTFt4KECiSYW
ws7NqXVnjJKIjjkQ9J7z4/+kuoYEDlNIkwT9AL5S7Da9TBK6j6tLbGXiWFNZKCPPFQfG0/Z6qP1p
zrDN5bW4EvLmpIAA2T5my3nQz8vHZmqrtqVzeySUlxLMZfiKgC7wXRol9HvkXJUK15qB5SKRK1jq
b3B3nGwseg+RXpDQuqbjv4fZPQ1SMkH2ZAOwV9qBbp1LiT+0SSsJMrXkKYBVFNE+kmI7UiAbliG7
pxyLa+PQ2R2xFVt0QfWBeI7roJ1tqiT5d+7lST8xdB7etb3nXmi0Q43ksXHh5qrGPdk9rgYvltJJ
MqDMB45tDdQwUBf4pNCJZAz0Ch/l1lo9HQ08qZHn7kz1EvJiUHhds9uT1PYMFYJY0WlvJ/yhe1Vt
xn4ckjOJlKzRTTpFkUTYoYcTCHda4HAZcqnTujmTkepL+P9PGlL93Y5AEtCLc85tIvpHIgObC2SM
Ub/NdCEiPDvvuIGWxx9fPJm4dCvRhH58+P6c7kBgOJylMzg7uJT/AUnA9xU/3KVQdfEhrj8DheVE
E1cSpnQuTEhEbbIqesDMsEwE0CrSA6qimuWWgbguV9ncWKkxuP7utrMv/3Os76U5CrxQs703GdxL
XKNkxslCpYk8+YdJCP5rKHWdZygBuORLHe0sCuhkKDDu1MIHbt4npjFt4B9Zl375gE1V6iQvZJSO
XghoKbqumJHK6SGYfIJ2olW+Uu8ix8bOzK3cpPsaCnIusMjRXdJRcBwEbeRQOZlkJ6O82SueMnml
MTElxzAEJTkqmP62JtJEM8FMDsd6joT1IKowjJbLijPXnK6GUtZb/OAjR5k3rsk3AzWHDpbaaHjm
qHruUSY/yTJH/dLywe2gEuBxorq1f0BgQvMZjpXsxC0nZj8Sqvh5Z5XgfSzm2aGMGi7QwKmLlKts
hr0w/zhM5D0PIIPzMjAqw2HvWFcl7c+jWRcBRB5cWVyJPgi5ylG5x6liMiIGkhDQreE8pTQUDllW
26uHxHDsOaC9Q7HKcOjWyV/FO6dToeFfik0mJQH9+DMQPpjOWbQdGxFxIo6Ui/Dw2Z2HVaTGGEUx
IiXYbDx21KhFPniITw7jFew0M7kEl8EcSuBqZQY7/6ZaSOpmZiln3PP04stN16zIuuY6b5c87BPX
rXziGSx/cxPcLee2xZS0T64d7CVzvXwcf1TgIK7OQfW9o+BwEsCjvrq05Ax8sdyQ7qeXjskS2Z+O
EWmB6t7jKqHB2SA8aW3jp0WYoJEQnOJc5GHa1uBBiKKXipCVwoVTCvHyHqg1c3CooqCNSo1VKRMb
5QnHNNc0oauaLtdUEyH+/BtNAia8PadaRZYrsp7bGqCi3kba33m51hsmeNOlmgL5edOH36Ig0Afn
EJWMfWhAvXUEGdQ1Ol74u0lBxCOHfg3W1jqBXPKLScqClz3T8gvUhXhKQhgNBhdUKLIMrZ9Ig7LQ
toxkIb0iizixB6osQtgxp8p0w9fG1dPZex7PU3ck40U2ZxKhnyaCMPn69sNKLKkMG1Hp01VX8xtC
m3hppiTO1T8NJCrWD0Oe/fvTC2aoVOYNLNllx7TvncG3emtEGTCiJli3sB3Jztwt4plC3rnRH68t
djLewFU//WlR6nc+ejJwdzEgfx3LuPJjteOVzeD9Jy8wl9tg2DIwU8HE0wEDiAsWtzmG9Pgw+vhi
gcEYYBwWueUIGArDvxEmru/I503Wf3jC0lnTSlsMUhuXvtDshJqYE0Nupa6LXQsg5nZvRK2F+5TH
pKVr9SMGV6L63xR26Rtp3u5B/qEWyAO7glDksVF2O2HS1IU0vixxZ0u/Ch5PVO6kNfL9pgoS8frP
wa3UmfT91OBaQXh02odovMaLqZqk0xyTp69QhOvLpqXvcXDouYV31O0Nl5GKVFRsJ4qyzpWwTIr+
mWZEusiM33pv7qooFrAA7w2Ye6lonmHs2dIP9cgo0Acf/pliYALQVM4Y2sFS96teBLBFr5mFwiCO
eP2n6yKI8PhUx5vJXVKNMKBfbkKrsACwMpXIj/FTnay5pzNMvZNlHlHVpNCpSnVXZP3qn+DqSAUT
tYioK15tyttTERZLkLDdclJk2NircSz9JhNahKDYjwErDLr3P7/3iyHvOyJa/hfAx+eMCWMtlCaR
20pnkPsPGlLE6y5zvlh3r9fVn5x2yh2MvfszLxEbUURleWW+7VM5pLm63ax5AnMHVF7bzDKDESPz
9AvMeha3jLxW1/jpHSfh9uEIWZrzQd42G0TR36rSll0++7CcKIfmngXR40/yboEgKfo3DTMoY/yC
aQbZ41zIQORB2sTz6+GOFhm0UsLxwfySZfrDheSdUSNb5H3aMmkxZ0diylKUs6MBEBVn4gqGBAgy
cQ76/jAVsxNX0TTyRGsevIDwjRXRJAQX3+TPt+NLVet4IwKWj35C5XW/iGRIL11JEi4gvt98Cruz
qY7WGOj+kgRQa/ECrw+ycxkrVhfENIqB79KL2qAAytpDlID0sZZKFO5YqYrUgZ//fVfmgViK1kFN
MpkJMPw6abBRXG5JvQy4701dnCv2DjxTIsKkHSBvKolrQr5rAwHVt552xvl9cCIliD88rufR0zy7
hGFjcqfykxxa0MaA9L7cbER02r0auZUPmJE1y2nejLIpcOhadinhI7gp0OPJt3HERlmMf41LyrAF
BA26TyiEiQHQATaj2btHwJrMD8DCbCPQh6zjBx2FRHG62WqrVx+icx2d3voMV+RgMownZXBfmU51
mqyLW8JZGItW0al443Zy6FmuSaL5A4v5+NDR91zTLlTR6b3B7h2tf7ra0/cl9GLQKzvNdKyuRWMV
aLVfk1/05g1kItBK0EMl0bWfaTkL/l/YQsx+NAL2u3Z1Q2hs7WmanaB1KQRsTwDLI4pVhUVvowGc
OllRLLpgZyqbrPmLC4exlFePmJz4HUzpwANp8ENLc1iHYpnEY3BlmD6lHnrjmYi+NbBSzl+pavs4
M7z/RQM0xt/4NGdKKVLiuuVA4NpX16iWUaODc8X/t5pXAOlkJx6eVr4M5UtPHGtvZ2mJ9bWd0pWZ
rcOVP034HGIDBs+5JKX/VGw+iwvdn3wu1ZW4bi33DOGuerQqUoZu/L7uA2dCqXQt3Y5gBvc/uAT5
Bv9txOz4eMJ5vxg4zyau5dlLiLGPCHI/11AoMDoHSAGr836xyPOGWWzbI3m3OaCgYx2rXlxoInDt
QtQwY3g0QgYrE6Ebq3ZyAnpY5OfSL4yPQMevYModmA4563zrVF18FhVOOtQ3UOx6RdtrJiPSRons
bETYW1ozwAUXCz4imG4fCnBclb5kc70hdeV7KNUN13AHMddhR4YEN12mVJi7SxvHZ6r0PNdXOrd+
Ko3KhOEbZXMwfJHxhyo/DDSyuYoNHBxA39NSNdbsUef6WF3J08WKqzfG4EGsWJ/kj15ACw1tGZbf
Fae/s8sMH6gCoPzYkbmPcfE0BDu32Pp08OszeElFz/kCC+Xc9n/m3Pj4u6ND1jPsSLhj4rSFavLH
mYyVYp+K/aeIfVbPQZsXaF/pE6p+ufeEY187LKWAy2a2haSz5ekFvyapgKF/ts66rp63Zv7/TPHh
fLpEC+qoBk3az4e20eQfk6KI2FvyYy4Cdki4s/MpMTpwnZPB02KFd5NvOnBOIWvX8qO5Ba7d6xwy
Bq53wsgE4EUl+MLkad4Aib2JHJjfSt0dziUkypaABfJCUMj3WRbLa8KFnzm+RSKfFBqOpFGPjWkI
ivV6ycBmsmHrVX1MZ9utHpMj6gMTjIwfm3deRdg5WMb6Ba4ebiBurMvk4FR5+UbQOgOMQUc1f0gN
/eJdme6uB0Qhrc/zWvLxNELTTgmFzlZkeOC96Oem88y4rvtPWalbBbp0HcGPdPshh68SUS9mMy2u
ihxbsAl2R1X/Ytj8YnqmKjPymZszBls2Ax7iqIBbrJ3/UznHzIQBe2Pt58jI3CwEPLVD387Ugxo9
zt2DSblHWuqZIlLLgFf702X6SKgH9rhBUx75k9IibKrp6SKtweB3c9REdJBVmKkEoT/b2llyM7n9
H+9YSRp7O86GOOn2OYqszPRSG9xik3ySR5jTrsiRtmQskVGPDcODvzKmEH2gdwzAieVJ6a4PZrCt
o87URioJxzV4ZlGjdQap2ak4Cy2CjrVvZBjHZJ/8fiEXLV5emx4npwgTxFADeqESAetnuhslQ8Gf
Csrs/b1+Vj/eSmXNi4sJmAnHrn5XN7tKerZ5/pVkWMgGgC5Ew6GRf3sqaZRiiC/7R2xKXU89r5CE
96jMMaYuOmRLdchOk2nxCY107dqPSUrSiuuCoX8SMLodZdRkLY/JmY5Rl7ODEdXHd6zo+OwEXm9y
NCRJeVyFLe+dnlRZSFriBNtT6oO//G83N1mf/CB6C2wXz4fECVwuwsZRbBHiwlAydd/vmEZXy3YL
tqzB8cC7/4S4EFc2PI9MvV2nvB84GLoBTRwmVssJkyMelxO0YyWtG4nunIppFq63pF76eUZK/M5C
3Pd7TGl7uj8kZUQhElvZDN4Oz1pMU2XPHTwBV7iKwVb12Q73vYRDa1+iqtkNxQJkmnFIKCmyJS53
XMjCm+Nbl+OXOD+iIou3q968e8lyFETEO46cdT600w9o/emT7J2uwoobQP47wdSiNXBk+CLM/jMr
kY5YYumAXS3sRvA8JDCNPSUrQkWtLQIHspkaWMsNlFcblsi+TVHpambEQOhr9loXTvLbeZIEE+TL
hkuewF/8oGMk8zBOV5sMFREaXLmg99OB/nUmkNt4o3ZvkC3H3afv7idQz5/iEDLDrvXmS9fzedDl
dI21lIkl6COlz6xLqdYeEeINll2Fz4NZWiacAqHvpY8ZOWM6WJ5uS/eHBe9OW12LxP/EN1u8Sf/9
AMfCe5rUhJXsJjr3ZeHPND5fqigEzJLG57iSTrMnTb2P59iPNlTltk0oxBECJbVm0+WC3KeVm3qz
hf+odj2S/CHLbbU/zEQcGDA96DQ2Aspy3kpNx8Uf7fnjC+ITW7iC6P4kNdEpgRRuWzUi/vVOM9iQ
k8jdnvCQ4o+o4rtLl8fISf5vo+e6CmGPFoTbv9OuI/DNkafqpAq5hELsjwJ1gr7w62E2JB2Wp27p
skgMshOgJYQ3LeeCnUuZ9bu8qJG/HbDKAWdk88UzDrscxGBlFiYajV0He0hE6Sr8SXY90leQVkVj
jzQQarCsbBG1hG6XqjCf80uZLcs6Pju7OY/6iOz5R68VijVnvGe1ku5dPqg/8i1+90SXiqaG0+Ir
98hRtQ9HtzF7jVaLbal5XacTTEqwEybxrL20Vh603pKeR1AGGdwZlzLKnIROTCn4mcI4Qw7WA18b
fDRPA5LLEKcezwmu8Ff1/s7Q+BzBLxyw2XvikntvVxJb8F/lg+C2cMTcqQn9dvfVVm49bdCGpK9x
iwmQwH5WTrQNtI82L0DYxHZu1RoxEGqUXeFlabTkDpu81S2xqJlIUewV6fNPnrtVHU3YGgs8U6xt
dt6Ea24eBbV5xYe8/EXw90uy/kJedS3ZkzfVLaNhUhhVSm197PYbSqtjz/HNwFa7quIjkUaL06mk
Y0LEGoEgXlGUCD41M8rWk/8n+4SP64e9hff95A/CjqZtppnPirdbhEaKRJ+KBjeQ/L09CHFyf33x
zuC+q9VDWf5WZ4hNT1n6NolDGf8f76vgfp6toyYaj7K75pGoSYl7f2zi4j0jd4zLSsfkSJk5FIRq
hDijANtoMRHQ7Bu3ohGle0sJT95ZTvmhcMSVniUpDEVsqdOfbAU2HZIASJiL1rRbcy/V2J0N7Ovm
MaFcmxo25E1i0cxLSONW5367sLVCiFCgEMmL1aI/sBxQoFpMA5iQh3L4JZBjDmzyoKzw65B8Vw/8
uqjTeklIIwyYqh4ToFMFQSKLYnuVVgMsZptka3rfiCCg29lKog6Uh62wdSAu/OuTRNRa8y+ZD/Af
Vx1YWJ+3q1Y+m5kUSefdunZuOPEAbmaVhvzduSRbtpMhlfkqmB1W2xQUOMu47BUhuSHRihiqEIga
B44b2FWRX6w0PcndW5VW3//7yFtSHkNSK7oS9jlg3s6IdBoaVTgGau/A3oZnqHA+w4maEluTSO56
KA61dnKQO/LVd3CL/YU7Lbl51T6Rl63yuq84g+Dk4RlEmweJZQVY+pE276eEZao3ZCXz2n8JXN/v
LctISVguvn+p7LmUb5tswQcMXVCbVT2wvTUsyKvgfQw1IDvju8ZsQCJjtlUHtq6lcYXUlfsN9FrO
NN6ldc6Iz79KvJpq71HuA/LN3KrUrb6rJcYWJwhz/m9lwTNIOUDcOScQZPy0EHGJ4r47Rr5qkP4l
EppN+55O5p9txTLkGgs7adOQ7n0l2AJG1KOkpWZPceixlDvu1UuskFKOBbkPRwXZUIKMbIcntaAM
8JKohbJsiQy1k37NeIqaHyqGbj8KulLt9hzn/AXrN4s2NovAYHr78U4HHyd+05fPD9pMQRMabqWq
KVRaCzjbVE6ad0okggt8wBuxxITPqc+kvKts/wD8SUGenVtrUtwgp0Ec16Kf69uw5iNTJUcV8atV
41eGNZKEnZUKZtY99OvJ3HCUJ7nSP/3HL5FtnbskXdCl6C76ny1jHb27O27omfXkH7pH7as7bmBv
bZCk8Dzca7RBqZ4UK7xF5WsVvBwD1LXZXAFgn91vbMW+duAqhOpvfDY+c0ybuTiPp+dgWykqF7J7
7KreM4gC3zTnQf88E0RW/6mt2pn4VrOL3Bvl2x6Ekawh4gtX1e4IgCVrbEUu9vm7QZ9eToqzDh+A
GXR5vzTrtTUQVjzQNGr1ckuaRQ/Xq/9JJZmEfdBcOuhl1qoc7vHLCP9kc5khDdsUaKAxDiNJx5Hp
xpPWv6F0toZn7s/tT9Q809PhVbjofo4KGphR11YFmbLaZAfZmXhLZJQgSzywBcR8yt1LoOYa0zxl
fTbZWodZBR4NyW0/qMWT2rR1ctgogzES4PDvDY62X8TY9BpNvQQ1RGQT9a+jDKAw+iICrLlx5gnj
8VYw8XMbdFIShhvTqlc5kRkBf6rfowLScjq0zdqsELifACy5Z15hR/su1mM3LaYTTL2GLbmm2km4
+JvdBsAkkyFMyvULb5wIxoIGDybjUGNBiaMSFwpF4J/UnvD2cVu21vlfd3gTtNU52FdzAZI+O5Q6
4NZkQzv4mT1WYYhYyEEHSAt72NcywiuG6vlxX3CkQBCLfdwe5qs7Cz9GSyicMuPEao0F/PQGbJGS
Qa9EJ8SzvhtkY2YDbiibWj75Yarum4YIkqEtZdRi1WR3ZiICgS9FjDyDJMgZyIL1a6jqMtE2bE4f
UtJ8ETVvSkGjTAoocy5TYVotAT0/3FzlFGzUhMiKO0KPXsErb5JpWJ3RLzxQgykS6kkKoLa02bd1
eIve3e75ZEFoKF2KNzvppg3qBjrOl5yN4LNiA26Q7ZUcZSjG1n4GVP2c4Ru5H/gAyiHSns16FodW
timvpVxZp/2nrLWN3LRxINNyK/SbFw9ZIA19F+rxQyLwOVRWSpUyG3RSQwCXhieEm7e/iNboqXCV
DpU2A9K9hKlgfRhbFcL4VwIBqp9pvmz2q4Nh+et7p3Cpbk5gENsJLsdELQhzSQpfNRL55lg3fVtE
JHS/zwUqMPx/kuPd6ag/R98loRln/7wOsO1NmI62fxk4CRyz70jaiyXfIXdwunxBnpA6DL+HKCvR
Ch4o9dCuOG8rQv+2t46RvIJAPcWAUvhzWI2wLKgJD6J0yPoBPYxn7Wiru9mSU8qz56fuVBXB6Kji
7myOaP0dVMn4n/sLELUXcHyOym6ksL6ISMGVd7f0TLvtcZqs1DqbCGMhwO59O4q7AY/Yjm0arnl+
YwWVQjPL2N6XT1DfB8KAzyCcFUFnmRSj0GC2CKjeR+7IqOLxPJYm++Lb4NCev2GHXx1kf4YHaLB9
lNdRupXxmepfDw0+uFP+lAICQskQ2CAqQzbyn4454w2I3PelbsSDkMs8lqQi6CCY7IhR4Z58fMuK
V9IYuDAB9OhYsIIu3Cppg7E9CBjQ9Rm3BnsAM41uOJwJJbynmZoL93Ed8lsBMginckeABxVaI0AF
QFFa94gCM9W4Drjcgh9L3n5wUiDct0IC/9wchHisRJJvrPJWxpwZ/RNqDhtH4XOYuIh285CIx7jk
2JqXe3xFsy4GLTIYhJ3bH/Vlo/WiMEJQtuWZ3OiFA1Jw6WK+u4mHsUSSBW0qnbmNGYaKCirvEatH
RwJaWqUeg5kws3HBOVx2YKsjRpO6rTe5c9Thkp6bf5BAAoHgA58CBcztV1Hd3Ebpr3BGkzR/7ek7
Ji9idHAdyYUtcfqHds5Eu/eRrZGv9F7TuDRStO/64VIyYpU5P1YWK6YNGJ7XmFYdfF/ubE5yDJIr
Tu3bWt7/LX51Htr/RaruSmIi+hXLOZbrhas3U8KjrNg5LW5Rrqw37wG2cjm8ce4FZtZkg+4Gb2a/
cF+iFrNSDSL+Zuv5RgHTs4I1WM6ZF3dfNf4aUA6jOhdMTGybT0r9jP7jvHo2WR8K9QxpoKn5eRWi
+NJUb2lTudo95nuqPyGsmcRvO4BtHMgD4jbT0HPH9Tj8QYl/eDqvYxk57xq2dYi+zFY/5Dv9dwEa
HkgZ9oJbJmtV+Fdgz2HuE6nhlk6Nm3gBhaLqUpr6KxSVpXyPlBBrKbO1x3gAbcOG4YqnJ7vmIBsM
e4rTL915pJpK9Qols4KEW/clv/efP8xtbTMaBkHSwdItG6vy7oJylW/l4HfnyblgfG74gYzxrKr8
ShK1Fl+efT9J3XzwxRXwkmYVIR+7jsK1qFJhNYUU8y0Wl6uBREKlNR+ZuSlpEsLarrs+YYm2dR3V
yZv5kmOXAPWCOpY+c0tk3pssnPVJG22+Ra6PtAniO8Fvjsqu05/S8pAiCSyKQGRG7C11PqGduuQ6
zd2y2Zxe93Urq562ZMa2yuq+reWg8HDRxWmaATS7k993boqBKzsHyMOdOzIev0OqL0s/0WD3VAx3
NQZBtzflIBFnuCVnPFGLMSzxcxcS29HVKW2no+Jb+UVrDDkmWHwQLFRQamHDJibyfqlTkzqjW+zZ
iHMQzvWU2+1jMJad/iBQ+i2r2QzKIhZlVlcnzIjzxL7JqGxh3ymicspmuOHgYtImuW7pAaUcqYCg
mYziBtIOEMIWjpiDQShCWupH/hc0VSVmqR/1TzR9ykW/gkgk9ysrn6rv8UCRvkmgVe/I35asu5cc
OzQVGRdp0YC/Ovd77pcUm1M06cxhAa4Pb0hVXTe4Qfdyn+z8VvROucytlu2BjUtt27qPBNucoah0
HRfC+z/DQQGhYuKle6PF/9vw9kI7RGUbp6hgzjXToc9G9pmqWiq8Gk0g2fcgs7QVbT9VZT9TMQeZ
5W+PIE07nEwDd9ebE7LvH1IhDeO+qI872342QMvr3fceT/2TSDimUWXzWaLGw+ExTmGReRf+30Cp
01ansSii4fVR5jvC2oiH4tfBmo9joSeX//p5ToHeATEGk8/fGE8hl5D9xgmBfuOMZd/dWH1YOr8h
NL+zYsitmV5iVnCv+venYeNOF5/wuDOwgOoWlT9SB2PxcyJhPtjmuEpadtSXVF+IP1ySYuLjIggi
PbMwW/O9FimKsSPx01Ol21CxuCAoAxbj1jlkdY6xJ7Q+Fsg9DGYUzo++OyT3SKTZ7KFSKENMXdoE
jrut1lZ/CRd5zpHOiSXIGJ/F8JNE6z0pQTNDCMnSCYbN+Br3yvguCF6WDL9SVJYs9C22SWC/2gGe
yNFxIpREKAq/7LVgZTaQKt3So+a/bjPFvkt6sVFcRctUH183Z8ohX4fHe/WGP72nzjc92rv37W2c
EWqNH24bnhsqWNxHeGSn5qt0jMjsufZAiC7luUdhs2gLaCLnAo5A45LuVzj3weSSksJ6SXuhFvhq
/tldeXpVCbO2+8TsLjDcRVJdvkkbdmHFqK1xdnFcczyVe40AtqP/78rweIuxzfc/s6r8gIo5wgzF
VL0Tk4rSLOFt+hmkmiiO3v2cbUp8KHiGP9hrODV7mSpsHLBbSDnCeCiDRuc9/QKQHsshZ4krf3dV
9raMoQ87pySdaRXA2MkU7y8B/ld4w/6XJFeKuNVouLIzdVifJ9HUmGsbopR/wbpNpADPDLfWU+Gk
j8LLdVN802nbRHupA58RYu90qpMG6p07wvRtSxVhXJmUGdDM6jRjBI02c28rhu8kXXWohvKIQhR3
B30IKaLQhBOyYTb2YuNh0zUOvD81TSODq8lkclKNSoy7iymgcmNKJdsKQ4y0S5qSiS4TCUcOtoco
EU6rRcPFkNxS8aQM9yK0fiMrNPbJ4aJK/UKEZ6MZaaxWYirG/nEZuI172WEvK/LU6SWWKqqjcduK
oOQXCZbagT2RdNA7QEs2TQtaVePHF5hTtRFiUXzFM+uTGzF/ACXQNw16KHuRjozrQw6gage/AZFX
wrvbtrQnabCqs/R69c8PmNW7ojJW09n61ymOyaNboFrO8Q1V2U0NbUY06UiJPBWb+FtiWX6OPTWg
EY9TTjKr9Pc+3axmZbpMQBN6w6y1AoGg9S5vtzsYirpfLpZZjXhZrTuzv2zfwi7hAe3GKfk6DxeB
OXuP62vljjbzoePa00BRKBulLrAkpaZY/Qm/B7LNZOWhP82nPCDWkAro0yzcjeCLtqldTuSbXO1z
+P6EeZ3NAkpmoLYGAR6j89ewtpKk4gtK/WQJs8UsuUEJQyqIChea35HShBrWaW6VmyDrNXti1Pg1
/bHVAjcweHnajiJDf6G3s40tb59bC3NAICZtmjTGOjzAn8F2fQz2te4mFwQmBo7SUQU+GUQbGNXa
MfuMnC/a9UElM4lb4Nct8BFHrDXefSCgAA4WLCsemu6ShePdenYZzdRIXpmsXp3xEryfSjd8IwFL
EDv57R4pd2ppXNWQbN96ypXCXRBMg2b3X3T2kg8V0gbWmAZFGhn3ZDOX3f7PpKbnt0t6tf1Yjc+s
FsyGJvcTRN3dxHG2KayOm5XqCmHorzn+DepZusIguSexMs+DCITR9mgQilotjQFPsDntMGuv+5AR
v3WDn2V1wdZ3QhU5fIDgzTuiDF68juT0PWdNYEr6taVlRbH56kGOP1T/Sf8wIiESh7ImCUN184J/
efYv1pwVAEip7VcCGH01hKW3X6znZwsStzwueQ9W7vLNSN+5rZBZSHJkuRt2K1LwDDpkBh/tDK7F
FbJn5n12iWRoZIqRRej+d0ogjqUFEIYZwv2P8Zq/P0Uhg4d6VLDPQ8BXG+R+QPsZSPfJQf446d0T
myYjhMLJhIx1WZBqWyWpE8U3EF9PmFfjJrmupoIcFcDFcHtyZb7wuSoIJ8QxfREHdaHPgmn4hM7+
6iI+WQkypDSUgDsQKeubsT3DNCKU+2qxgQx4PmQuVt4j1Bb+2RIAsg6Vf38VRJxH3O9JXiPa+AtH
biAzN/2wFLaimI3O+sfecGlLJB4LoXCW+GNtxXn+KR1CePqW+75tAXNyCKXwz0zQ8VrCxvk2/1S+
mfxVTsQWG20e5xlUYRlkaXbBYFUKPszyujs4a3kDus8jawKcgZhon8TD3HNg/Du5ZQH88kIy1638
vP45oGcZlzCdDUWDtZ7eCTrLaFI6O9+Z1mFzoiSlKbmbuBqf8MWfYTM3IRmYMVJ533qBPiTF8GAy
X8KOUrCP1yuOQUkcHXdF5TcX6cZAaqT9+YLiDJjjIftZ0KFCui1O85qRIUk4bUeKSzxYPOeYNjGH
Yqb3L4WmVGwAqaRQ2LMtNMTe7L80WXoHORZHmZ2od/4M7i9JmuIgibqBxiHDtGfDmRKQcXKsEEDo
wnhYcOFc3RHtnrhHL3KfgkWP/l1jbMclavaHPFvl6zvegISC/XR4LK0mbKYNzvSOL/Jv1XUN0L5z
m6QE/xZ7dWy2iY268dZe8paXT3lM1SRAGJX0N4hSJtNbYlT8LmT+9fbchefubKhqaUtZ1Hu2ZIU9
qQEBkybdrke2bXAty4lhmrlpt7ClrS/hBeJmLViJqEJJ/VxnPQhDj5HyvkPMTTGO9aVKetr5lx3V
exjUkSG58b0sqGX2r3NuUa1TUxYheKGTrM2bWGxTorN+Cx2adSIrZXAL2z0K7jQm8gNOA/lF7fyv
7l5Zwwj1v9NbhyuOBbP8dQX8S/rYC2YuF28+lgRsfFxpdlN5GgT36hWnrYB0u/czzE4ES5DeiZP9
x1raDsxlExQNrwrs5VaiyMDglcsFZsnjKJfdjHQ150f0YypShPXVbFAQX4LKiYaVRukIXYScC/IE
DDBXqjZ/S4wUOIi3LEsmI6hudJAF1GtlR7dZE++kfBBVmmsSwKe8SpUZy/JW/33+d06en+6+dtLO
vFwLhPneLBw31xPeXZWmnVD5pBOnobBW1Z2iecDGKRj/gQkSjwTtk15ZNaCmM/stbo84cYdWIBoD
+XPQOQIkRw64kdyB6iCV21weMA+jsiiPd6lNL5B8py5oJU8Q0sTvNH3oYqqrRsmn6x3D5mx88JXB
oD9RDU/XM7f48hJ6FfEUKQVmCqBr2m74TXeHgdRMVo0cO6CV9ATz3yZu60fu7+CO/nHaYcKoMtjU
3h9BSdZRTz4b3Y8G3JIKPlQS+oEoTr94jYMUJq8UZHtH0WvIvA2vSef0VYyLKKO92bTI3+dZAmCb
gKEuQ8Jw5MN4sSJCxdgEmgYtY4X61SsLYMKCMpL5c3/Cb4DL5vUO26cqQq7q7g2dQ3AQjSkHqxOj
qnEVV3bthVCaqtMF41VSqFPeLWMzzLYb85pq7e8cqZvGWI029/4SET1B7upKbVZnDpwQAg7Vw8Wi
mNUSeOsiAz5DAOCpgqRRKxffh7nu3p/Tl+qx0TNF26tMuFgWZf1gtwc4CTnaOTSOFXQv53OXMuXn
uM8Q1olL87NPvjVIbbheU6/vVBgAroQXJn54nuLuzKN5ijd8TlUIegzIlNN0Mo0kH8AvVnaZ43zT
P62H88OVjTeZCXCdcJWfphEKniA7p0nmgG6ecGFV4zhu5dxta7ltgyFBQJnfzerk5/NBdju+bTOI
jcdRvNYZfZ5XOc0MN/wMcsFDE7IRwFZqo8xcXZHukwbBExjEJ+DNQ+tgHx9D+dSY2RGjeDSQiTB8
hdRMP/urWPjrquk6xhgh5bv+McX64Afv89W+D/Ti3eXY1X5L6HvydP87KKMxZ/TX1/MxycNjkY7r
joXw+K7olG1ngoOxVWQ57hNg9YcRCmU4XALsVwPVCtvC2yauEtThZUupJZ8sfXVSg4/ro5UebksU
dKM0numqNE+11eCBvP18mwzM6TOqI44XUxIp2W1VODfyTlRzWm0ExQ5yyX4hF2Ge3DoKUiEbokwd
H9Q8xxtlUR7MweKm0tnzDz6HwOqOsdCLR1VBCBbaL+OoGKtVZhalspQpxRFGR72ytED7I3LtSmlk
2RkQ13UtBLkQ57HZ73c/FbJ1AAyyx4bolvAb70vnONzUFLeC+SHSr7k1IpO5rZYra+Jiw4NdGvHX
rSe2OcELVtCzJp8J+5tSo+U/r3nLEtOyzvtudz6mErczuPvh4tbui3rQei8M96sqeYmRpUMGyACe
CKcEwzkNN6qmYv0700+d4rxxCWVLugMaJ39dLEnJFk5CTCXEsY8rYjYeyqUtGUXtjgvbJvXdbouH
sxabx++IeEX8OZezAwB1zIKBcjK1WwIHt0CoxxlO+Lg0+0RXyElthw4qV7/ymQtYGfLFMjZt79kZ
5ZCQEQ8FiBwtOtLzSoK8O7nP4YoHyYOOQ8gwpzjC87+vmBz8P+nY24BrvI8q7OYJVI31Cl2Sjle1
EYnnnZ1kVaDLVMCxPRC++OCY1IzOFWVLbnRb26bXkw7QlW9V3YSapiOg7NF3BXbzzxJ2sM4T9TTX
/LhiliFcbJ10eQiY7aAHgPAJdbAAJv9ZsWONqos4jiIebfGAJ98svjRxyKHrgzELHKci/Wig/nTy
Oc+HaI/lq9Mb6TFzkMFZTrwqSXj4V7psmg8rXYsVjLnvx3e5rRSFhNxOnRj1HUv55xLubmOgmjcd
WTGiGqd+k6lkDtEOeFOpM38y77oevq0AB5cmSIFIYeKZEqIE3siU2M2bWVjBFuTpjS+sszb4t1Pi
yq/80P3mIBnpV1emHKSXxViqyY8n8SMhRSKSovIAUcl8G12mIsvXCU7+sFi+rXaDDl8VRWc59DFL
icqj7E10OhlL4mx7RvRxLifAfXnw+0QW69GO+SvwDx+UA/Fl8eUXAIHzHe/iRVjV3eIyk+iPVLUE
nplDHk5kf00z0ArgdJyU0ExahjL/7N8rk54J06sy3EwUQBvssgpXv5CKhrfivelWBpGdOSHDxqsM
PX634lXobAh+IEkp2E84HHG2MzSoy1xXy7G/EAzPzln8GRXtjhanZ/VYpJ8dc3qBH8fHOXaIpw4z
mhIexo0OJZh0YwIzyjkD0KZwQH/0JL1HkBPKEOxhScufloVuU1Ml2EyK4/CXrcLS5hLAyxCgFvAm
cibUFtheQaNNsCRqLfs1SeA06CfMz/jWKKgSmWgmbYi7xGao9hNLiWGYxOCPMCqUqR8rvLIv4EZl
IDn/8oDAsmDavA7J9t/pMNMoEuB1N0PmNUulA30QXG0RLPpV21opVAhmt+g1gB/dz+wisDM/ZoEH
WlklsljZ3II4g+P81VAMYlF+gkXGMv5HsTG+mbHT1lhd2wU64AL+NGBmSrVj+K31lTaIWxCoFuvj
147XDXx9AaxgzYIc0F7KymjmM3jT4iIVt2vU8oPF9ocf0XNLycYUlO8dUqZ7mZ/C5nsuzxZIGXke
0N/HoXFas4fQrsc9ff8F0tU/eODmY8ZqIk/a/+a74Ee1Ffli7lmMybPbBXghdE2oOeuqwLr7fxuE
Nkemf1cvmSYHQKIuD05Bxmwtxy3Wo5jSuZyCOlHqgfzDJU70ffCVpmsfo3RxaHLvff7dN/846Hry
9p7Za55d0JOaQSMxouBvsRfTqUfLO0u3j3oBor1QT92tVNZiew0xu4Tv11f6qJL45f7cp0atbgas
qLnvW1bVHOvrLjbixH6nuNepohHhYofzmb5TRCbK3CVUh/2/uNmEqvQd1VJDs9ylcCr+wvUYXyYB
ryolDkCwCbTqedwFjgFTzAkM689U+QR1JAO7x3ylBW3hZL9J+NIUWo0PpxrCqLE7Onhdms0KYRt6
p7ET4fJHjZY0ae3XvRs/ChQ+dtXuCjQFABkLp01dTBIBDEH2JLmAr/P0m/1Q6kfsiJWJGWuxxwST
WABWRDuviD/9KCYOgTudv0M/DP2UwNzTX7hu9Ex9LriScmYPssSE7Sje9xtHXZHYIKTABXUH+Ngx
nKJLrH5StNcVgA5ZcvXDL4YUgXzeswbOACE4LhCodYvBkmlf268OsjnpecI00zk2JZc0QmNvL/5b
qHvR/t4FjkmyefCEL1qH57GTtG2baXiBo247fBRE68+jAKxYylL9r0x/nKWOjcRMBDNQSQDFPOJN
qRXlmIPaY1k7L4V77gZ3yWBCC8sAbKBuHii6TEfKfPzNE1neKZVzLMHOoJJnvXREaWEhLnSEDFTN
6uEz+l8yoUqnXfxNartKke+qHwRmq0j/TkOeOuKP1RK1YXEUH+9N4BhExY8UW2BdM8XTlG0rV3zk
UIEx92ltyKweTGemHnbIiCumtbFHaLLoGLrpyBZo4VvWJo+N0vDxfwBAA47k4evBORR0DgbF/BY/
xS/4om3JvITZmsJQrayVzUZIz0n6j1IkYRNrjZUTdJJnLALaxtcuI9pljaKeKX7QZ3UpfBlv1ySH
lBA3d7EqbvUhqrk3uNA1+1SYLkrvjUt+4JlIWi4bnpRFbXYHJaPU/e4NsLU96xMSGK4kwMswnjjn
7UawT6OSpLwPUkh3drIzS+6o3KZ9TuWX01P6AUxoH784OP+dH53dVaU2kIBNcl2kQPf0dLg5JWcd
SfMGOHzI7u8b1JU2749WlRd9fkyKrQKsJWtWiVEPCYD7ybBPIpeawiLn0Grln8RKoCAhta43ybnU
i0bbePKjMypTU7sZQdhZrSR0cFNJbuF+h3dSt/XrFR3skYR8XiliNVo8G8sM6oAXjuZLmcc/I7Fo
nN5wk0QUoLOsxfEcyW1zkNiP0d9sPVj1ILc/WFj8lpg16gOXnfE3vMDWVNnZA6G8KSXKUuSFdxAQ
inBwmwN/n86icgfZN08WshmUrZRs72YK+ZpBxIq01BKDEqyZf60eWcetXNFMCnU1BZX8EKfr9hQx
5FOZ/Zv+J+z0VnySqWE8CdW5IQ9Vx32zWGZgRLpgvNUkf5A/fGPvmTtFYCxJEa0Gp6DJlCUSxSoD
5xCJy1Y5Ulz2V0Tl50dHr5KEgffyjmNhmmFl1VEleBJygF5rEYTAEyC6ryrBYqS9pAH0iETrcooF
VkqfYg2eDPIVl6o41vK8fBCO2PkmlnSjbo8gUURmZkJGxQgM+wMJdRB3DA6eInFuxxhhgJRsFMFg
vp86SCD5Yt1iiOPBAwadQEvPq3B1/xEN73YkAoIXA8b6OW4jvK3RKRyrTDilrl65jwvwOYFpv3IU
vbMgodDvDMd4sYzp193Ox5qhP9oblRHlD3zjb0pGFsLipPq7UnEpNGcZzVdH2jkviHEklFSjxnGx
a7PNihCynhNq/fsPsY2FR6h4I7NyM3T52d/SaN7GT7wmLBRtWU3ctdFZOVbA5r3VUCH5K6qmS6SF
aqqjHveRG6atXNkFPrsa45EQ0KUhYS1cJ3H/lnfdnjDL2Jxjh3vA1Jw6o16KM9G8B0ljb5w1o7ci
vuqiaQoE+qtYjDK5JLRRVZ/4OwsLM28LaYB/B54s3nDDg1Hahn0qBMJQSi7G2oYlro2etEXLgnEi
23BciLN2VOwyrgts1BLomfki4D0u4Y8RefA48s+feWflVkcrxMOE9sfACkTkTIPYNJLVPUpjpDVu
ZxK9jQgBYh5CDqKGWqms0a5wAEg5b2nKCtwd0G0Mzo+mxO6cNA4+PFUOliNDLCt+779auPS7TYUp
VwrDrRxAZQCcXxZYzC6SqzmqbjDZ1o7vQdoRJqspYT0ns6stV4C+ENJ3hx2ThSIH+pR5XKt3kXlv
akTnkQAx1erAoPn+XS6dKI3Tl3871ohQlWznhi9+ZxyLeCf01G1gPEqBsEYya2IWrqyu93YSmg2Y
1ZWM/haQUqaV8ZHozXEw9k+6fBP0aXkb76uD2KAgYRi6sEsDsk8Qf5cbHH+0TK2owbnsASVeCmeA
E5JODU1fnhJPvGfZcQ2J496UYxc/QZLzQ4uUHhnU7AAKNOcnXC4eBuLSCHsPRl4wRlXqG9tQj7aV
7smHuOS9xeOPIHvESvXcSoVZ4vjq3v4ZwZNLqD1At+BSfCCUyI5VoYuYXHura9Nl0GHixhrGRwH1
2z5LdxPcFDu1HtLeFVf5psr0Fv6o7DdN4va2XWhVH+OxP9FGjmhDGCq45Zs41e0UBxSui4lWpPtE
02YWz0XSqaua7ZwLZXsYOlS+hENHY6kcalSPaWq7WjdrNLrlqgxJSotb0X+f78XPqnO4CgLelTAJ
8rvG1x+KJzwmFFfML7eqrBfdJzRzJ4vupHHVZY0lND+BsuzddgfDCJLojwhuOqeW2ODzr09IYGUq
Ml6q1IEz3L/1K0S79Jlg04diW6SrAKhe43Y4shs8DknGCKOwqtUFmXDuMWiCkjHMrqQDRw3BTnmo
36ejOhHoRtq9Si+mnr955PwyNtXd2zLBSvZscDKUQmDWExCcrAVjsKlyzN168SU3EmPEkOs3aUoh
kNsGqIxmoOX669+xFpa/xwMgwqX/tDjVI5X7OUlOuWHBVJvY+7ZR+ufZaN6IedRWuxbr3sl39sWI
hmp0e8zUQliurxL3EG2Dd7ToeEldO35YKkugtj70EJZpw6Iq4Bqt/B2s90QL/LTyjMuO4Ok7zcn/
LOhNHE0txoPA/7g/UKlICptleWpkpCJ9Flx6QsYSlfQPcGMb66URYHzXNkCJ7cxC/BMkGPgyog9I
MX5PDiHdGA+5QJmW58epxsl669B9gXgGMIm7Z7GFRvnHz+4AgeluyNi/c+e1g0kKeqR8pJordaL7
UsaHZP5LWbybXJ6NMCiDhZyw6zDRJSCk8OeTovzEcLTqeaOUqaPARtoQjfO/NkNAaPl9b8vNCmsk
FH7erkoKD/yPJSeZvwjwTi1WYsKK8OXrHRNUzlwELWn+veg3Q4VImWKcDJqHLK673WwddOGpVaLc
gA3FlV6Hyji35UiA2yPbI04QI//4cD6S3uGQ6BngaoM8SdJraR01MqH06dFdjOr/7L27a+p+Tpzi
z2vxhdX3peHT7I/H1ILvJiIiPMlJ0tIt1mEm1IOV70jfBr1yjQD8QcLlrHXCrwJPeYrnbjLkydu9
RRHkwzHvlQBBU/pEOa9hP1Ww4fS6YJ8kscp1tfMUG3lPtq6eD14wF1GpikXUMwAeQu+ULsv5T5OQ
uidzDlDHeOtt6wATcsCULqJd6mCjW0Z0ZfUqjOlovzOvg/pBj79j7cv5uvAU9XilfYMBsSuRCw7w
R9SbFwhrqpy/aPjMeaJC5lSmWRqB6IrgbeXcgsCuSosjPeqgH3kvgg0f6L9QuEMgiwTNuzGBRc9/
+XMOwfxDXSPM5IRPzJKSs+7RII1sdJJxg9CQVtnXVmP9yKYm3NzEiZ+kxRiMaJrSGzskK0zSGTSR
JNMHW9IFqi2+TTm11ObiFt3IWgQt4kZgOneaPCekOCrGQhLD1tPKYW1aLaGvSgJJzq78MAhIE5Vx
6OTk9bGFf3wrSprZHEZ6vFyOmw/vCbLHuWKd+QyTB/Q64CaIevCo9EM0c/rnNMiVRPcuFoTCLksO
VeOMHLAl3JDJmweGF8YHGhScUXYX+fp/ungxU8lv9t2Yje5067Ova6eOY6FgaUdvPUEKVD2Fp8H9
B31REAESmWfzg7GnSVUPaVjTy6IlxIjmb5LTgg4rv336eQKf7yN1QtWAArj7Uy2irg0yWaBV1G5P
QmwcRosUJmczPQrEUwt5pshmC2LF8dk148fSrsiSxUdgakGsg/I3GIy0PME7cFHrtgtODKf0JhBt
kqON04EYLG/KKi8Qqb5jNUuGfAf7jAcPh+JheFl9aeiYfGCMZE+jb/NrmusPLHkd+9RqdAIOTLkN
IL2UVXWh0yksDIo3ZbeCIQkHIvXrpGay4zWPDPy+9L0EkKCpvMPSv3YqXFrt1CcWDc6Go0rzY7n1
PiFVsAfIazyzaDh/v/2VDwpOKWCvY4mIxMfXwmn9J/0298+6tk00KbANHHfoSai9YDqCvZdikg4X
JNSvmWZd3GnPNWfSyn44NJ6Wok2TrRmR/E1CNObRXDdPJqLyl0hLrF3WufoZAnCLqRNc+nTtjhRX
ShhrMfmCraQnQzzMVrBo02+qzjjVv32fD7P/LfiFlRG7QmMXa6+4LT7GeWK5h7nlbEg4lk7bAAyQ
93VVEhNKd3JW0UOAg4IsDc7Pjum2nTgJxV3GnPC7a0o71KPhTI/rX+5Zr+VJHMXNHnaHTnKFJhFV
MKQbuShIMXlVIfLqGrjQT3siNj/J6LWbOxulGyDsfpVt/ljHoDjDdR+qEsm8mLlgLAppq6F+KgPw
8f8J5r0ZEBIs46vCi5RZyRaO1bAKJfdT9lsttKGeWAErFGmpzEpzovB/HoimhTUtj0ddoGDVObQE
qOEoqLSdDf/4nIPJKSf2n6XtSArO65NHxagZm1AUp++0LmlSYEtgGu9iEYy/ULPX7Zbh/M+p19TP
UF9tIqD3UA+BaNpVMLLhpe0LP6Xg7eGuyXj+YN1DTPcjaC1lr8jXIE0mzPNuMD4TtTnztGe2tfwX
Bqq6UXg5TAshkEdK+zvLiQTYxCAcOkTfZpXfqpNFZz65vZAuQ/fb+oo3kuZj3ngoBljbtH0NJ1K+
jQ0VMf8le1s1Gj0/UzDPULjvFnAyQnh7XZEYVHZ0+ruBWXWO2kY0PmvmjC6Yg31UJLX7KU6KsL1/
w5SlwXFPL42XIJOeslx8lTZXfkf9NARSPS0GlCgfdyTULgeGvx8i2TKrlq7TsRWHUT/RWDmzjUJl
rwG/iAAHZMUwL4+0jZPeGmASmNjy2XVwfSAP7WeBT3F1ACA1gZ75Xg4SZGKSPYNpSE9/Jp6VrCnU
y8w/y5xXaExjAbhB4kqwXe8JnIk736VLeixL86GR0adMNl6aSKO7u7aVzluLQiUJ0xGZZDM+Ka/V
j+TMiI02JKxiS7078zmJ8B/P0YQGU4KcIK+OdUvPALx+4PbD2Quq1Jh9ULNld47u9HogCbEOgLIK
TBFLQIVTll/AN0Xbym8U/Hzxpx++5pK9NwNDHZa3Jq66j+DDETZBpjg6+EuJ0a3cn5BPJm2EK/Ze
s0Pl+VdrWRWlrlkweoBSq9HfuTrB2U5gkmLnZu1+xbdpWS1IWovdahF8hIJ36vA1f02mF0atuU3f
vXlbZecj7BJGqNLkLN4N8a8tPRpJdscI2Vw4Jwya4M6VE5XwDuACEJlpbfQr1w2BC1XDVMUCeszz
DUm3651f8kCvtjZjpUkvQC+4ubTc6OxLGFS37AAIUoqE4hTL5hL6yz2Yhg6IPpqQ0wKOT8pYAG76
rI4Kc27LDnUa3cZdB4p9zh5qQY5Ij8HmA7FXVdk+UnzEV72h+roC2TqD/tETu2zTPADmsS3qpniz
92WNcbke98vD3FP9BqaH9vQmDdpx5oYNr36f1xCN7nn9d1V3XhzPIV67SSN0SJ4DpYxUvNtMcUZi
m3KxfZtrgFI5kV9wXwxHo4v6tUwxEsd89SKvwlMg7eGUS2jyUd+9fDeX/AwEktjPk9w1MGkKpenF
FA4LZJUjH06fyOahlL6G+8OFNmFRhOs3lkcDiQL01By+DrliTO0BY6z0q1AB8+bU0R9D+cwsVXwp
CVxvbnhRBpTq9h6gXRlu52zZKDnGoONmQRexgryh82/TOOyCHr1GmZBdSg7OFDpfr43tSwq429dB
ODlktLpVC1KXqYlBbAYgiunUO0UGjdCJazFaixiFOawEMKlhVCj6RK1CjxYUJ3bQT799m2xD/ZL7
8pzIHVC3JeWeFoqAnZ5Mpw38Hl8baW4we6mIthGupDuoRVzln6S/98QKZlQVdZ/0uA2QWK44ZGbh
DnL/DTBew5yh45lO1kQSscUheKn8dxhfcP7iT6s4zixbJugRTYvRSco3c5rJfDfSGSmaxZkYnP9m
Loshp+/opDVGKN7CyPpoSgMMvVNCjAOiv/FwvudKNdqj0h8ekrl2Nrswzqoizvy5dpgqoOYH7wRK
olHHWl3yLiBOdoJV5k7C50fFa6NjwUEB5uABTEdiVhH/I4Dcu43nu6Rr//hrWWlPw0SIjE0N2sBQ
e6JRXPDqUdwvbm3zTrSsG2LNOvYugs1PEK7W3I/XH4SXTicL/lp4MANZS4mXML+9hzgq71PLmke+
uPaoD5LitJ/Cz29WPqS5Ry1iIVJxlg4JuSIhVF8CdYHgho6ox5RKR9VXXsFYtBogixZwyerekk5R
/iyMzDJ/D5RXEyJgYg6X2dt2oqq7yp7emGjM8laA98/qIp12P6pWGeG9ybI4oh7Eov8S6YEcMaij
GiGOyAdJwJYQzLczbwWaCMkMn+YW2m9IIFl9mXbLhTeruid3LAd8/7cM8qFfvzPz387Tgvpy/I3Q
boHdYbZLCOYt/C3/ujRlo8V6Yu+rUktsblYB52Q28QLDjXqt9/ZzUrGl2TXRb31opPrhfhMbxJbV
c9jA/z0q8JgRy2M5DKESDxA52DpvKbW7t8AEwVrSfvTxrjKjoe+loFbi64rjlh+2DzTTO5zJKVQ1
AJhZbEo3JXaeIIXfS4EHjX99daK/HNN6rzaW0gB6byRNPLIUlGWrm90Iw8XkxdLYuuSt4cmYdJ4p
Mpek99FNgPqDCh79VCjY1v3QAMvRuyHQIlkueosjwUacAJQiol7x9Wu37LHSL+yecWevupx4+IkW
IHLJVCKhpsueFF/OGSnQTAVw66toapZmpcbmzQiEdZhQG6KLC9wPXd3INslUC9eUgSSQhpw3MUXJ
AHx+MQ75RovyU3RAB6sFp6mEHUB56q5QOqvBX/H6TagfSz9cmnnQX7BFBGzgcsbc5GGH9puNSRe6
1MW9ULgnJ1dCdjhyu8DwC3phtQw1DwoZJWYyLON8BE2nEnWQmDn/owHodjeZgch9pZ5tVHdwU2D4
32HxSTOsidAHrjzWo1Buzst8ygCOOVf3UC2/6DFrPda+Tny4BNg6wQThN4Tl+cQnEvyjHZBhZfF5
v3amhX1nDJ6wICS6IstZ8HglAh2h/Imdfln+LDoiM0lFD/C24amDL0d3kdlMNP63QJtBWdrSkB/D
YkZZvYEDQXrTmrxYicedE0Mw3/4T/xEMjDphpaQoPRVWiX6Orr9fNIPSyu0YWi5XN4y2RKr7peI0
MWUTqNhoivtYDZlGT+k5veluujDKIEf/sqzqpjDAJGUgmZZCimyO7mNcn3tqyFps0iRQyzALIhu0
GYNb20RKShNMsCNNJovjhiXS0U7wIzvCJMDcSs/T9x7517ObH5FyuZyW+84z7EbdYbOE5TFw/WIu
kdBtQOoRiaw0qKgsFiVKrhijIyQ37Q/uotZWIU+Uh5O0KdhsQRbmFIFZNLoQpveRtQpdFDTC0uWu
8GTuixHmKiYGuIZaxwXUxYkcwsQUzibMIeiIX/NPQpR/f0Z2ki75ZLCHcutxD17mAzd0y5BCfcy6
xAlOmHR8Qb3pu4kHrYKj9lZgq6oV5LMaqr0iTTBHNoSRMmBkxhP3XfkFq+nMliDTwLFcO+o+HXuF
mO5tQvWIWel3XXPrXiXZoKTPyBaTuwqCyWXwGdPgdw9o3w7S9IxcXXvm7Ud6zN8eELJoFTjTYDs/
Vb656M7bIvGTyHNCx7xtSQCuAAFXwdpDDgl4z5prXBx+yGzt3/irTyf/uj/6l1aJoozJqdcCmQvn
e63qbrjeAKVapS3841WYnYJFacnGzH4M3asJcSjZMwP/3cKVNv6y5TYKREefjOQ5JKQL2CDr5Alv
yh1wuUoIip+Y7tte/cCGQwDs9Pctprr9fv3jhCX2j+1iHCFwxfPpfLNuZiJupv8PvynCvn7W2iZk
hgOTucymPVHHqoMYekIENC6HAUPl6r+6gCOjBUdoGNQMoSCJk+5I3ytfHliLVxfBO3t+PCgFtPAR
j0eVHHquHTYdf0YuuUgQzUXpHPbKpgGxR5yzeI+o5vqUTpuyzF2Wtb6MoSOmdGuNKyGotWbMHpqm
QArlov172bjKU/p+BhYJtTpOqE/5MS5bmlMNXN4gk8W5wNr5mmKhmUFoW2LnPChEEaMSq7IzjOwS
7VNRr63j1KcTlP77PC1RBBSwI4391E0/kqc4XK5MxHEw5ZDdbjLCZv6uLca+Hg2m6Xoj0MyIZIic
ov1/7qoTmpWYJ4a65VIHfqt4YPWIVwtw1mgQ7fbPwtExUalR3jifKY+6UB+lZQnzaxF86Rc7oNk+
y54kTo+WduaZBu+wVxquf8ehT2l3GoPZNfc/Fxq+O/WMixlPIwKWGslQvUMVM5QwREbPbInjNx6d
7nNpwBkXFsCFYigRoVQvHBGxYVza4RhEW46H7qr6+HY+lIk/eVM8M9dCcsh5ZuxxqIqIg/nhkCaQ
KhYBvO4qVGzSwP+CNLflIaMmqDKgJXE8sYEOBzHHnd4+HBim54XZ/4qo/c5lcEa5J9DrhRnyE2TX
i4hpWwi99oO6VuWmAL+VbhWqmCKoetxtPRPQCe4CF4fHl8bNeyuz5ar3q6PMySxGTpL9EwIwdO+m
d+OzLIbP4XoPgTsYNRrygLDxUsSpddoXSSJP3sq4sXWs9hHJN+Le2Etqz2QtarlUeYupdWN34RV2
bYxH1CuvikanLnvhVhIESockZu6MfVjQqjeNIhZ+Grq8eXfoWRAY+P+LhXRIA+wN/j1KaC4u1G4M
JNNt7e7G9GNcwAOt6kW/64U0E6NYHKKnOzb35VVFf2pMXRCqm1wsrjDuK6WEPiifPHR37JGg/ARj
nKX9xrnLYi99hWpLGleWuh8tVcptgrg+jic8B5KdrTfrq6oT1f0XXb3K1PlWn5f6cDqq+EEas4Dl
j1JWOGgy5v93nwXU1I+BmEdNeRkqQgustvNiyjwP7MK4RqY0kK2RooOWpRtYrR9XZHBteMOPdoEG
cz6z2IOEKg78XE6upJHCfSy5mo/elrKy+bH8Cr4LUBemIulkyABXqwxkJFbMP8+TC73OXADoJpxb
M5fIxQEOub9x0UuyDl55rTFGKp+q3okBHtEFlPH0fqEBzmzeS8Gl1/trnpfQIqD1mhwzIpL3ulPj
AvGOBUQqX4jURO6i8XHkbPj/w3UHdsGY+LSaSJNAyZNT6OveijIgO6iTn2sMTvucoIVlc0vNVWBF
IpUMgQA9WEaheWZxilBj8hDs8Af5He2sgwcIHT8OEAc3X++yAejb31OCLN+7tGPQ9xsOBr2BEucU
yoJdk8qAA0rhSzcToTRzgixnTLYxepcNgj2eiGFKVUXzv2fatqnjPJn0/WpR1tVOqA/96QlnI/Gz
gg6PpkY7enFVcB0qvcNKSzY0kJEakxYibyetayc6gUoyUtfHhcAjvFYIMdzLtP4Rcx226YrdmJCv
3l+iNc0/0rf66VNrumy5FG6RorEsy6c1xK2M7NivJP6maRNxjwB6Rniuz5AAMD0sqg+6WfEC6z3p
i2V3bcCYldzFiIuf2H+lONCGtzT6IIjhK18cr7GSQsUXczhyC2m7hPq2276fYHbKiFBb5BWvJkpH
N3ZcFPKAE6dZg0sdM3axH6irf5iRdAk5WARP5TvvRd4LdNsLdGyoSVbyIDUn7DSMZirwmy88o7Tn
AhYedbdtNjaAPqAK18UG2llJtjjJJHYdz567XZCn7TZ/jP13p6QLZGE/8o9nV7VXSOhgHjt+exyE
2OMdI8FW1I4oyrYpYzWwWAXt5w9W2y0p83iMpIbde8aqalACY7wwitIuRGgX/mxekiPagfQP9Rp9
OTajcImZ5HcS5WS4Oy2I5o3EsJLFEW6nq9rtS46vZQM/9+1v2S7O9AB4EWu61gUCW4xbP0+SQas2
UD5QVp+H6uBJKenMM0bAhZ3skHr2nRwbY1Fq92UsxGL1RkRMGSBBaONTsUgDKfDM4VVmbwwky6qN
wug6iUBOt4Rd6RN63DmKRe8t3nIUO7x++vbWSHDtgLdFzqUJsnKKS/uzvWNQJv+jkz0Gb4EoKRXJ
h6anAYcrT0guMdvXxXmmU+ybN1AmVvnmqQHVr1vlAueXcJqXdYTWySmSKEj1sC9HTgy0HPUiaFnb
hsG1wSAU/pIKJi4GaGosLvUbu2NdGtRxSpWijLdCC7dtyI9tbALQVyXBqEgco4riSeHVHA7e4Xxz
sABGRatt/4DGJ3U7M4gxu3YOTdwGYfDGQnbm3BvvvdAtrMHSW8Y5ReQBSin4X9OM7P6N64pZP30I
xUk19N04LyGpc5fCO7m6R0weulV2DzKPr8dE7nl0By+lsJ1G5Yhx83GrCWJ+8RBIA9HFJMczD/4N
1VlpTeE6MPLKRgP43q54h62jdbXDpWf+BsBMoEOs3yykfjRqlarCA96hReyKRW82g8fyFYLxYtoF
Ar5xqIHrR7zVHlU0WrsH89dZhKHGRc1MQObq5Wa8CDyO3plV/Kf2TZoiUFAuM7AJREecgG518N1B
l00BHBEFGeRtFivTeZbFX8IrtRVPN0mx9EwlJCXUj1B5+3Xed0Zq6RoHUvR46UpldShrgIsV+ga+
evOYGqGf5YBwKkngw4AqBjhoqHvQZz0r4dOnINWDQdKjWpFzNzD6IDtd5fDKo7nUgUOqvQwyKCJj
5uL0aJ4x265GTI1qMc1AmE08yetmW0INkegQXR/4btjmAZHtgm3a1WYKu2pjTmertxFrR01NjI9Q
TwNAsgJEvSdtMP9BHNf4hsReBLjbNGQd+HKqRQB+DsPnOAhTi6VDkuZhks1umDutmlHmshEV6/Hb
CyMKIiSt2cjv2yRVl8pUdneuoXyS+46UCRI0rxJMKx7vE0I9cLAu4xJMqlULUQNVewXyVJxoby+y
f0GqYE1qduX474/7wxMvT4/dSs+Qd2CTB1GG2wLsLzkLRMN0aYv/3HX2op+PmDVegzyNDaFl/fGF
rRLeIQlrwsryX5Wbcc4K7gU5rd7i2VWxuWfQf2DNaOlxQn53tY73MECpsk7lzVldedw4C5EeW0rw
ayEKU9NNBjpXEYJwNRJpOPhv78NkI/3GhOzKBYIv3HeHWFGCZ02kjW/EIBJ5ameqxPkl+cnBlInd
7Jf9mD+DgOtDSphQM2VoM0RTssMrZ036PJloqPYdlmWFVWoRlR6p8+lV/WfukbbUN17AFcxjM8hz
SdMlttdUA6Hz00tKQf7q/VNqCn1JKuQcbIMzLdikcNrAbrpz5CujQDv6aqHW97l7TDF8oM37HJel
ZUXwWEqD7Z7SRQyeAjEix6Plny2a93ZizSIXaJ4RdjwqnYQHoi238Utx/0hOftrRql6zhw4Y4GrL
3+giU8PLnmGXunbEVQs0TIPrweqQ1XFHy9kKNYik4GYVHWhhydQ+uaHPuVAIaTexXlmlHAXasVeQ
QXDv/Di5Ki9MBUFNR9f97SZXY+RPEwMc+4wUUGpuPOTpy2jdq5iiNP3px64k7Mdu0xS5txrejkAK
sHXDUywJhyPIrEeylz9pFJLxsFeo4IoKv5+b1VRyrc+3rYBWFqF4XP5ColkpGWt80L0LmQvFzP16
BFzKMJmctJKjj374Gu9Mrfa/ePcdSWujuIcE0KkNWPYNE03T3zw2y8hdLnx9JR2Fj9ouDJuY0Re9
WOB2RaSTgGvJzo4R25/jFXf0YAjK57wyeyDKax0HNDkHiSdYC7iys1AhM367pzd6lNJ0/wWwyi2z
FVsgwsCdlrIPfeTzEZMhEZiqsFwmaxmFjKwLW7T6EpKu6J2JwmjgSlaQe+NYg6ifyR88YS5rKgz0
qAqv5m+nGy+qH+T4lzY3WReE87E5do1l4jSMKz+uh4U6lw+P0ZFPiDBZW5KYZ8J9AmUFgz1qI2QP
DswMbC6/o8gWTJOb3+BFXbavIG8XRFxMkk37Udo4DFfZOOpogEKcznwKXNzDQFHCfGl5yNlh2If4
+4WDCEN4qkm2EEoBdttjfzCuFTHgsyqe0/DhMaPxihdLfySZUSqs+G4gQnlSgd9UVfvNCRMW5FH3
CnzDs3eHQ2+ZtKnbPPKmTa3wuws17earvEy0ExJIeRAI3wgk7UvpXwGk42tQh7x2J427bGue3iUI
18NsbESBTGCyM22GXhHE2aF+A9usyU4XgKLBGHNUKo6DlVjlsSbemhUFSb4Iqjlt3SUn/dOK1DER
TYCUZ5AOCuIzaOms4uN3CHETzGqf96g2Z+iNYrEid2k8pNhxtz6A0vgUdZAiRc2Ug0e4f0EGBVNE
NxIeWBuXhN7HUFqH8ute0T+Evr9JtkWmwIFEbtpyKDn4e7q10IqDF1xmTV0qVNY/bAtPYf2ymSfW
Zk+jACWdcJ9VN8Fh+XOjRvAVGWMOenReObqroqiXrwfGpJ1lrVlTqJHlFXQMVI5KwBGoE3/zPKgM
z1XaLNClcvmlMyyJtcIMMTbQADNVni3Khn8FE69Klh1NszhQmNKUSZ6Wge1O726xDzpP/2jLklZW
Eo2x6hRhK4oXQ6z8OMtWCTNEHElLLYu1JY8CzBff4i/Vl4GO4etyxpcNNvSPwXyWEAnGnfjVhm/2
/O+yyfPrEXShM3UfJh8NetHlxjx3hJNTUjQsha/5OaIT2zPsED1JDGNJSsRaXHnHk9OPUd9kio1I
rTo4tA3OLDB96W+YRoijz9AFoab21ffvmQyXx6fTxsTyiKDW8PkGOj9Ig80uvioUTXqCchH1Kw4E
eCDVai/G+fkNa6sKSxplEVLXGMf0+npK+kxMM2p4ganxpvIJi9jpdfgFjCUlHhH6KJlhgLJ+CGcq
y3prpb1h8BKa1qrHKd4BjnNRgnt0nmBR77TavMZlo7A2eAHF1eGAlcsPFqoKwdkGPwK2bsICVm06
rTZtLEysNFLqgrYvKDpvRvzES1ANiUaf9SmT6Mx8lmlQHWc7qkMmhz7VX9FjD//I8Z1MPrLkrKUl
BHTTbPc1+s7ZQPBuhVfmZ0EKMTqjczF2RC2w3sADVASUxyytuSX1aocpGzgxYYQOd7wfA5o40qMn
Y8PQPzvB2w75y6ahAnwWRzte7ZmHFSsNCiiVMYjL+2vqoQK9+yyLtPIBzHgd76VUHrt2+wUdqGBy
WG+luNvCTvJUAExGqdn78VdjOJRp0B8aV7cLtFqTjVN6KqZ+1KwH7xvNms4NHxCJbpMKkFM4ZMf6
p/Y3aSgCHhsFmhRGRxztycNU+a286OyznS1hvOBjVURTHY/xGRaTrDAWf7aRa+xy7sa25xUXbW10
rjfudHERegY4+31oUwfgx/UCY8otwOo204MsOUul5rl15KnuFcf/sFmZ5n5PeUxWZ3xLMAlbx7Mw
OGJkYUAEimiXSTWYyD7pN9G9dqNSk7MW6k6MkTYFFqFig+aQh6FEakgNZIf194RH9wIB31UXYnFU
23B7g7j25BCzvowSEcsNb0F3SmNQpEszEh6e5St0N+nG+/iHaN/1/bRSadQDgc/xgrHeO5qf0clX
ch1zznmz0i1fTAq2OGdf0bOHhv9oQ22/6iZYRJFL6rkkRJV0XSZ7hUBZCUweJ9L8Kw49VnLR5alg
EGFQNXkv8WpObDNYEWK6uW+R0yUkFfj2QbpVjxIEkdxs03eoB67U4aY907qhtrpBntQS1omiPd59
V5PwMOsNwCas/F+jyAB5iWH47bMtp2mgt8Wp1YIz+4ksrgrctnh/AuQmO/npBPTprgM5wDD3glZF
PVKZzyONyF63xjJjQW3oncBBr/buUr1caOqlIYsCQ9/pVoK7Wi49uT9Gox9J2ukSGkvZB2s1dmCn
IfUwIECn4/ullDdLZFSd57MuQvGRSu/1Dxew0hS3Xuto6c7YwJptst/aQqCng/22IwAjcWdaT6LM
sIPSpU7KZ0icM29HpOSjKIKTr5EPrIeJqZxXa3eAOvxIebAhKmnGR1NTJ7fQclGCTIH64pNU2kTz
JtBqRfuCdW5pfY88mwqrhAzCOpKPVYfH9mn+xPyYBaStMgChk/s4ODz09JosXoda29q40j6p/Ak8
VV6Zx+U+BEcAnMjRMQdYq6WHar8ctfG651TL3kCYJqdIKlny9VEMUpnzWTQgP4fZvSDiL7eg8Kq4
glKVXnxsT5RihFgICdZNORe/y3fd+TcHd+snSD/Yf4dg4OmuEbodj4L+s1TBYuS89fjccFkGGtqs
7Z+umjpfeAGrCt9W8cQBqNffK1u9Qwf4N/2rkYZRslz3MrOfgBMxdwWfZHXFGjesbpURcvuNJkUL
OzwEsh3+ccwrblnbyl3FeDrF40TeUFDXRpjvI+G3ZqT/T9gbv9dEhifOO81xoCTpaduJBBxWrAKL
zq6Uqs+4s1zsgp0hm/wqQPni02AFXwBkw7jnm/B1F06u2lZphZcofTpmEQpKYG3a8QqONrOq/Ku2
0z5qFdzsjtFz7vd4UYtQzYbLrY/2rBOacPEdSyRM2Mgxu39AldCTpAaKCbkz6CVA4Bqp1ku+b9dP
ZOUOIqncmG1dzQC/UALw0hvnRASS66FSLbiByJrxKU3eW0mB8aVkCD6hQz0Qms/UTqEBRH+tBhXD
dKS0n7lJ2Opft/HU1ubieLOf151zzFT5WQmw1Dc7ZcEdt69EOk8ZsXLNBrXQOjV3fLlVonLUKnW6
YF1xV2WciAhVdWObDxo1QG/8ZtOfpj7xAf2OA695pnxK9BlwB6B2hn6VB4b23wBfQ+8nePzJ2Gia
oYSnMafBOMru72yQq5AOg2OLnlkaMgdPZDxGJfdr9SEWXRa3iebvpSTu8Jhgfh98XI6MJk7PCg0b
6uS7d8tMwhGBVNai1Sqhbh21gg4O5FWMCnDhPbk8029pBIaNhqu1onStlTvxydaDOLa0VrjaKfzJ
h9CIBnE7M6RYa6z16T28tz2AXLumZE7sMs/i/DMQ6QMMNMYc+YLElFuYnwns4EpObYf/ZaUuzEYV
yVZ7W9OYCJ4zFkcKeBktkU0oags8oOOfXN2g0gcs0DqvqlotaKLc+Wqr3dGzrUVn5kETNm6Fz2Gm
Dw38Cyw/qTVF4r5Dk3edy6ZC+UisTGR1ISuY2WAHFAkPz520MGBaxD0Wo+uuBfgF0EM1Ct++qOkw
OgeiduOljC51z0IHPGp/60FW6QOuUrPpvMMyCjhV35P+Z4kDZXDv5TUjHaJl2k8ywAP7RfStMvf4
q6eRdP4UJfrbP1gqCdsjSo3wLCQMFxSsOhn+74dAa0vXGit/rS7Z00gMnRA2a6LfGjrRR+WPTIE5
njvsmK6f7fzJlrr3wQwjbYrTY2OfRKKORLYOInXBElUW6mAja5taS+yBx2lLF2cs0SEjNcAcXWhe
1TB6+i2KZb7sJsouRNLhVEOEc9k0xxcl7R7mU6CZH5NGeEqzMR10GambxZ4mAxjwLUoEw0HDxr6H
nLS94vIeU5SEAO1zZwkiwC1u6oZ4jhGnZLbawhGvPt8//bvY40rn2r69usuLHPQaHecQXooDjax5
ymLEW91ntuPOZwe6T7SsioKQw7mCQI7SwSjWLwBC99WggSGrRA16RQXRQG8tgwg7A6VoC/Fi1rfH
gv2SZhN2jiU5+rc17Q4O7ChCzt5cXuztgzGKzgZ6C/fmvFhP/02vJ3GINR0W6iXkSGBFQuhwvoTt
O8Ycf7RuIaYb+d8EeYnJJWFNOIpZurEQMOU9DmfMAt2v6wnODPF15MHoDX/qNdd2EZ270i0XrWaW
KAJgqwWEKdWStBDEVZEyA4ve8JFdCCnmzZyy796Q3OgiZ7tOlTnldRtflQoqff8sjaQgfDjbI1ZD
QWEEkucxyBxpd/QsS7Pro2Q86WoyrsyV/2mQR6jlpSJgoAWe00Y8t7ukSeIHpstUqZTK5k3TXzxk
KG78QliKJOL/bLRq8qcfbt7eO+pvx7BNn4VY3+K9fY/1rrOiGtpraXcF/MkdQ1+zL5/s4eO7FJDW
ryplV0Kc3N38iOPS1Qhafc5ZyJ5TtHggSbwMEdn+mVqOnRcLAt2IU/zApSixNFBwj3TdecJQUw3L
fFIf78aKYkJ9LCTSUeJwZqATa9bLhjd+nK7JRhL1fbbwV4Mg3/R33rWnZYCAIlaDOqLGtoPVdiBg
mGXIcYGX/b9mFoDOIl4nf/UJlpacbQ/ePDL7SZWoIqNcWGHCHBj3hg3zQNAHKAG7TuLwGhxHY49I
qI30yFgtN8Ba9tALXBYvp4fWTQJAzOb9v954VUxPxjk4Kl3k0bYR3m4QfIvVRPGw/hz2rwIVrLzt
wB0wcUg38Jb8wzfpOdAt/vj06agDRNuAkoY9oQelj0xNEVwWRH6m0EMdnzrMVixqGa7i4AnusT04
rJlISrkmrD1V/J53YrmdTvHlGxx5XdXodbsILY/HE8ojF+zssO5+4rxnuhczkzydBW/SzlQFXEWk
OuSCFcl42hDT/2fOUy7f7gcavE1zkJIK+/0HwkfbES8xrGUkkafwuVrr2HW1NVbmV4/S/cL60jQ2
pJoCIwaY/pBopNwQhe6niKZaM7r6TSDC0pMna3fCQ9sXeDlB3zWJ+hsDaKxhRVd8SUQrRW7n7b5v
i79ER40JC4uq6/fC7eNw8hrZiCjAuVbZtnhlrJw91AIR5qMh5vA44CWP6jydlgeSPqRvo7afE5dU
08vPDJQUp7Mx0JkBDcbMPx+GJAmlw1i7rfTY1DU/Mbeqtr38ctV6FP2DS4DwGcDTcqI9w0FQuda7
BV5ZsDkmXfkE141Ngy+9cCefC2Pya2pDYeHiJd06RnUvc4ODX1pPcnHx2DnDr+AzQvkt1R+XwclL
k7/XeNTrrmgQ0/Y3MLIn6YNLCGee0Zb2urv1GSc7xyiFBPySJnGqTYhwkbHizF2lOuTHxNTxD0Vy
uVyyzoaf7vBi3JLbKc2s5dQBOwLXW9qM0tT/MeayBoXh8SttlD1OfK2AJ13EyNAs3VJESb702FeE
2J3vspx9RqJjh4Ghdznz9pw5AGcbNY/+oaS77VGlEdJm2xWQzchCPNXDNqwrqQlPaN0/QmplVF8f
FgXp8Jt6OZRhGSoh8PrklMZXlYjqM3XevfbO2WGgqGLyhzuZ4Cml9ESlY4LhSBqc2anePSMDXcMr
MtIEl8Gae+TNR60NchPjIgjfqmZqQyIeU01lCq8JIRkv8w57HcBoihm/+2gyr7ix52ck2WGbffID
WzeQCmFDCz4HlEhhimUPh+dvCSZBY/CiZC/a0RhkPRoqC9tMCTgaHDLg7g4FEPdUMAuqHZKJL/6P
chqEgddGqxlO3fL0uBTs2No+3bAu+TinBTU7dMk3bz1tSzKDEZDFMvtlnnxAOiq6g0sy1QzK40xi
r5DtDJdFkbHYyopWVGkNca1/2r6yeb9FQSI/2dPfeexLXJfdOagaBAWRXOYbjRm0L4KN+J3BgnAk
7EpF08H+4MAkvQRl4tRVd7fs/WThS3QLeJYURyRhb49Nmi0F87fD3l6WnZ4uxbVZJaoBUNim64nC
v+gUCUNmwW7cDcKTuubc/LV6ixnXV4t2Qdmv+ZkrxJqz5TOSvGxUV+UKGvyhj8zXbrtDgUIUn93K
/f8z2tNCYpTofYYej7QtX1y/IvTDB5T/ZmL7Y1534mfkRoMJd4V6tNMsp+E/AUlC2kdu6oOQ2uvk
7pbqN2DhDTb3KKgf7mGoTsveVGVf2FuOe9BNY9FYvr9HZO5SqmmbvpoActrkdBdB71R7p2AoLdnP
sZVQene3SI02nAV9snqSnBjwlw0apY51UW/y7tRPXLPsHcUPzibolKX2pltcLZ9ck3medPosRzm0
MnTRrqUzL1YfDOvuSxwtbhPWYnPk8pl3jmqMzpDGfEaQTBYfOnrgweHFnlKqB+IivOSifDiXsKF7
ZgnE81kEy+oZdZnjUMnxEwlYjkeApW9OFdaJA3mjddPefnHl1xlImcfM5by/0lqlh6KhpH1psxcm
hbVEUA+sDiBR1mzam7MJb0HWY9o6lQsvZTI+jPCcAo1kqrQhsUPHA++aEPTzMK71vZUbdqYr7lnS
S98A6K3nK5dJLH8GnzmYx6eqGD4GpjGh20WGu4aOHWFqvXWxkuMBnIry7qBB16L7CteaVFvP6s5J
RO+EfPsQ6G+2BMIdfRXFGlfvTBbnso2pI13hKTv1FkRA2AAdhcX1Cy7D2MIS8mtEhuFSwh1GQuVx
5zf+M4pAe6yX93qjQMoI1/NLLVF6NnMm/kkRHnHW+JDCREa/ctd0blfPpA20Gk87clH20vgt9Fiy
/q6MhNE7SI7/33Y3UgjwQQzgI2h7LGzcoQ3eQM1zLNNfPHOWjHEY9HhR1n5guugidoXNxLlfipkq
Ldj/IuOHokM12ApiOKgvcdeckmfD4M2CM4e4vmAcgxHyViDVE5MI6fKl4YqwFlIVhDaBeEUgtjhH
f8M2bJerNeIP7Bbs6QrmQGdKNTQ26+XqimLFpC622+CElK811hYxEwZcI6Ty3H9ksKiqPed6NG6p
GbM/3Hcux3694Cc0aMVRwtWhfOBX1WoDxSq1feZz0RC5/cvY0aqELfq/c98p4DJqv5WMFkcJbhJE
1pIsA5tXWLPXRayB9ihPrPICBwAzIvKLdT21wnv8m5pRrs1APgS1hIZm4SgFMAqXlITxBrNjpQbe
WPw2KjrrYP/xqpmUOizz7DEfZEj4hM+kSQjZ83zSAiCCFvzKuIWyYagm5JoDcqyf+/q6xQaxVDMj
ZbFL6/YR9lXEThG43U5UOXmIaOiSYLnAKFnznAlCSrvdyJ0haHcOBQS1LK9B0zNe26CbilbPR1q/
9fS2wI1LwJj7dSNeek4rBhNYSeRJWiyF6VoDd/AcT4RKLONdV+QdINGmmgucbB1UUBxPvD4gdLtR
So354HMs41fDatMwPqbQ4uxgq5nhWCn+4HBUa/KOHIGIKBQNI4drTpPFkbM6J9At38/3SCT86kKd
+PI/pc5pBM4tm9bb0dC65x/xba2yPABDHOq5ckRWxiL7VsynA1iNbGUsIvkNf2KUDqcPnM2l4lbG
pUK2EX3tQbE8V5BmRw58ebds6A2F7/q7iDtisghOGZYq1Gz20fnqfiahfNMTw01ZrWC8RrDp2o9c
C4uzMipj2MqCJ6eQi4rKXb+ZbLrJnlliHnwXPvGdn9V4+WZ9HZU+YWGkvFP0COtquKsyb/ztpHHJ
Bmnhrfle/g8AIxfp0nH3JyOaH/3Mb2mRVU0OwZNoiTBk/j0zJy/63+0JQnGU/IDKxqAlpYeOYZO1
1HIe+gors5D7vHhoELzrl3kpss+OtZrqqICAC2bz9ClA/y+RdlHmNDJOz0pWf8fJetO5ttpyOTdl
qvkrt99V6v/pRobvs7RIVOFFyAclBsPuvsmhG5rylVz/oErhvURGDzcLN8yYEtGhiH/3+Q4GvglX
2qGWeDrEPUpEB3dr6xRiC+H5f1rg310nVGtg+Z1YnLZ3e/qjoyQpdRVn8JsMleWREXkgMKIUjWNk
llLlWnqPUztlapAB+O+qyOO4jw8FhgUDRxsf2Gl97Fg0VQv8nWbSVYng9PQetlINyBYa1NUZ+fz5
i0ONhUw8iqCgOTzeNhWd8JehUfrDoZaDVOysHhuUEfuNgmFRWxVqSlCKqPii7DdLi2kk2ieM/utk
fXWJebGyZhwBTu9lw3Y3zUl/tfLGIl45gDJ2pIuKjHQ+HUpXQEWkUxPFTOCqlH1IAGn73o8I+Wbn
PVEz11KoSsoTwrGUUrOMkBwJ9Z2KtjGVNROSvwil4djtN/7o7VGLwuvMApSDRVTXh40as2+Elful
DdxxUukaGFpkfJ6ZZFT75KIzScFTH/5uryQTXEQTOu+yD+SchFpLwOT88KC0AJLyYHIqFzlPWDne
K/xs1p8RuzdYPUnnCJDSferDnMkMrP5fx5nKztJCDulBdDFd99+5X3O5pI2OrZ8TFYFVJKcR+h02
yHFm/vn6a9Wd2DB4CPHxqckmt45dYXO2qBRFQ0fiOtZPjwFBtg5fzzCedm08g5Pet+kNK3uKuEtA
z88y83PrRrqo6V6XV3Ubsbanxh2fdiT2lcMr9Ds0kO0VY7L0NmR7thF/vgUxgE0nHS04+zdI5VIL
olABmloRLTqZUjcKf4qLt8RJSnyQG+vHqxo1dHaV/cqvIdr9Iasmt7E+BJVIBPgzXaDwOBzsUH74
9Z37gOGbdvpI6QgRVndeiIR0ua82zFVC503/WyWDwSc3S3MfutRweMxh//2ob48Rg/2eWqFPl2Ai
DpesSVXduy2G2VjtymUempHPs6PZ3UC+5TU4yIShTVn7KOld0l08LgOt9T3E+rZKJYajQe3XOayC
jXHTMdDeh1sv/5DNQDqee1EWZECcM0xO8lPoC5Pgk3l1njhcM93GGzq1MLbefF3VTSI7jQbBPeCS
BGqkiITcxfOHE6/AoiVG1sRFJnRZSSngZVElsfJn/+ji62xF/OE16LeUwEvMO6VqFfyDe4d8ygHa
y2C8x3+aTEYq6elRrdumFZKLXtlpmVueSFVIjdqthj4Cg7DA6YIQ9NM+gExVSEJNvFAZ4RHIq3Od
k4JfTcimEowcrCyCOPFj41DY7BnoLilH8Qv6vkg8fP0daRgBZx1tY7ZMwegzj8WE+2BGmGJm0g5Z
0PkcXb2Znq+klLH4Ubwmeo2ZVsuSicnBbIShAEGnqeELIng+IgQa2NNWbS5J9Xs32B612ot6GJaE
r1vVjaL5t/+sAa3wAiFFKK37ZdCahbDchsftOTaEUYePsSNgNEnNRjHXr6VwJwMC1EX+0nwd79i6
cMmQjU1IxEiu/baI/RPEydFmyHU4sKEIPU19r9tEJ29uLXfg4gJb6RfBqPmFMuY303v3UAgJoqR3
8U3hmHQIADVnRhDwY7DU8aeipZYqyaQtbDUq/Wat06jyG7Ofi/ZDJNRHyOUb4eWj+R3x5vXphbTS
Q7c1+C0X3TkkuBQnlW/qD1q0EGVoM9o5Rv94CycP1AqqETw7DkhkLPKuqZw/9QovNwwYx0dO0Ok4
wz9o5ajIB8VmH7hFA6ki/VPdWNCFCy5sfO6GmaTm1Uj7i6QiZfYImTAnHJ6po28HqgPg4JSWM7zp
q+oA3MWQSdSIyHtVFtPW6aYV9ImtE/ANHxHEm1u7NqxZj377IMB4zL1/mKpRDcLzpcNgePz5YawW
Z4nHb+5KDkxJ7hhcCXKptkZ6HiBOdG57snPWPZHNP3NEsFY0JEXQ0bgHmfS+6ALN94zqrLBthryT
pILK3QjyOdUT6Q2C1LLTwB4jVLu/2fSGka5984b+UOWd2uhBVw6Q2YDkBh9FHRTjtR/NY9S7ZR5R
fgaZof1Kqqyye5nty/01IDXeEr5S+m7R7DyeJ3blj31jxmnS+qrpqCemKnOUYc8K8b1X6cZVkgb0
QrjRF/3sZ5/alFiKSl9zfkLvnwPVtB+QPG9ArXVhurSoFfcqsuBZviMTgF7JCyDJH2tapFzPijKO
rmnPlo+ZvzMUtk3yIE9CndWtjP0kFQ0+Ia1HFX2Gagv2WPlEtBP+YXoAa5WfoHSGKZDS1RQ7SgKx
aqiUL3V7t5L4tuxcwncijJVljXqoovmjAse9qRvFf6bxVJ82pJWS0UYNBcMO4b8jDLGy9FdODtiZ
+hLhrwxzWpUD3edjjjf1+TOGcEIugwglvEI2PROxudz0sKP21TOYwDeQ+RRhNVGhzKRyO3XKufa3
Ev5lqjzHj3VH9cyiRrgWT4PEclRq59aKFl8q7jOoRV+7og11/1UkxETa7JfQi92G+3ggjweLGh6K
vYZssFaGJ5cltLILTihSMMnNG1T+Y7LoVWh/B5IBTs/MstwxmJ5ihr01tHEY54c8hx62JcukRNRr
flkIEEmjq73K0OyPjLANK4FomlMhKHr9rKd3SCTfu1OAqT/MTbHZRkQ5+KW+z1IN68sck2huSLvm
EUiBg22/4PkvELWtgdYWCOwna5uUtmxR69X9CLJzp6jFR82TWYx9ZtBK9kR6k+ALacK7uthqBtqB
ScaFooH9pdGu2r8U9klS2EINLhYJnya+GgFek3rDmfE3Xn5nfRtRqvRWH92kMIBBIMgHr6HQe7hV
xi63m+VX6rkBmibuzlXnkmAvtGjYUD3uP41ywabng1qCbzAnWFQJHpsxf7RSsT486DUaE1Acwe4G
aew8w1sD7RdU574noZYK6xXUPenA32YJK93fOgBq3AtRRPOSik3ukmGt6+qL5ofEl8alozS2yS2z
/duCri2509h+U4JKuBbFT4BQE8qSMWLxLJQsOUrTSa/DYcP9p0axrDJdBOGWlx7Lsfo7H2509FYh
vMjISYkswaagUq5OCPTXE74jGhwC49V9NriOVDUK4yzKxV4q19GjSNk0YxR16vdJlaBH2TMqc6L0
v3rJDiqd+SkLhkeuh78KkpTIkhmO8IdLmafh110uLnmu1DCNOjrxSgqsacvSzcWZAyUSmA/7ZUA8
wBdwy0kgAMpUhBDJ/DTJB60ii2eiCifGIdXUBoRRrjhUNlTyFkNZnPu5fnguwOx6lXpNpDlD3YTf
wSfcKUXwFntcK6/m5OhHeG1csxnLyeAiTPKPfzmC2PLCjjnEL2JDPFYx3gAYAy9NUZrAqJ7ETeeK
Bz8j+NT03zvEcMsR2PUvqaLluih5nSDWTum7GsjT7k3Fi8EUTdZwWRam/dZ7v9+X3qfI+cZMQ2eg
rpU+HKmkVpBdIJORB5lyrGPMC5bNIZbnfKI8183IOuAws+nOnvU94ucEf3WdhVFLpaD18ZPGkoSx
+5g4+uchpvT/Sn4v46jrAomM+T68+qY6YkKz5Gamf8VK975a/1MsNa95FTbSSHncbCBkWXlMdBy/
O8RY3hoh9GISwEycrISjyX/KIEW6aRl+R3doi5UnkWwWAn4BF+QsB0FcXfQcq1nLF8wMTbqfnUOc
PuAC/phm4osCEjIGKXzWnQEpID5NGPdlSY5HOzkVWF5bp/rPlqFYtCibiPyZPJ4+sbIzOcCveLf6
mxQMH8LxqhlC0Ju1izFzhw1Kl4/xwk6Lm/l9uF2YHisey6eDbSUMA/vW2wMMPFkmMGH99dGNwegQ
34IZZnuOAjG9ylkYsZ7kh2WeOJe5+8FpXvMTxi2cVyaCdm6J4EnyC+xxUVvy+DEsjBRhaDFNDzUL
ZMQ7vbnHhXxTbG7Dr2XjO9IqEh6LCqv9HuH91jW6eKUhr2/tAUFz/J9HsI+pxDmeZleR1uikeBuF
jO+cr7IpubkhRuZY4cZ6r+C8oqycqBHCp1Le4Lp5tSl5FhNzTtOycjXnu1zZK9CzdLKG7sZI2wvj
OH5vco+Rux8pelJfVXC80+lm+0goJtw6aDeIGeGtcUED2XR+70kfJO3Pm+eroINbnBLwIZPJEXoO
Lyfr0/SA9tajw9SnV6F1bEiT4Wzd1riQjv3FhNeTYUATpnqQDJEQGZ7DrKFB1/TijUoxWNZWQSzn
3le+ZXhVjcblv+mV/+O4UObi2Q9MeM+5pUyrji3fQwwLWehXyu1mNs2JUZ3FweVg9Y9kxy+hZIIU
nzeOPVVpe0+sXQr+tuidXNn0zQFad6s1Wjhyn+xcViBCFwUJCTMYsX3eyPdToCb95ALZ3vhQKE4F
7POLSo+hTcs2rPGg9A59G6scTyyD0Iomrg8W84pvD/388Hm5Js4ltitTduclhY2EBCnRcZX7A8qJ
A9GeS+Seosqvy5lQeIb7R14WkP222XFGqF/iEfa06qLu1teOvAIuJGGcCl7UXusgEY3qBYGdfXnE
UhRgIHcFVrfvDBWMrmnJWr5bLqmpqrdOkeKqnnm1AI6WmBhtrSZK377KY8Ukm68GJmbCWnTz7lDq
wqM32xUDJjGC+e6neYZRdxAW9evs54nfF5YInJddYcJzL/FIj02qeEoxK5RP0h8ug70SM5jaIalv
LgqL7NJJDTrnV1m42guVY3u9JXMSAhUyUD78R9CXXJ4Ywyrqdme7hppG9GfYJDqD2FUaIgOQW1Kt
wW8gWSWweALPkc+5SJHL+v8+XA/91eppvNVOwbin9xSLJW65Ll0IceGAGubsF4vEvPX8rNBJxg+K
Svhh6nJacM9lpCPp/eji2O9zcLdweWv5gLpiIph2sdUHY0Z1L88dLgZP5hU9SXauXdiAhrzVVUXC
8pAznZ1KO1JCuzf8YuVmbdE+tNR0/NX+rZ28D3/OAO68tLQblrPTOeGBN7yQvqb8iBCNuTjoFbo2
NC7h7AvmNclVoivbMGkaAUy/ev8lPHmW9FXcrGl9K+CBc/xrwrcfnYcw3RIRzZnJPEvMl+jgRmfv
cuBwIVVvzndhbNJR3LYyh6ti9aINrbtbUr/w0L+KDbw7Yqm4duuzqtNHH0UxHO6oH4o4LybAnxvT
lgO+XFJ+Vt6osl5unjOo32BNMlnxP0kSZazcL0h0rGFngBv4cAoqJpCQZlfI/ohNcdDsQMrC+6Qm
vBfIhtueqZTh+JoPr7+AUNCPBWo5IDafu/N8Xjr2jrJzCjjl5yRoZMggNLzuYi2ch4q63rPT1i6i
JIUHLEjISvLZwwW1POZhhpiQltCWQH+ZUeoFz8LNomtyaBYBr8dk2RgMw8/eO200g1LnFrI3Ynuo
ZkGiBDoJBvCwluluu09udj15okra48EE84YecR7hx2GnfDWDwkGQPkbFDoaIV0MxPcrau3FAVxso
zenP4BNWl5TdRd2bYK/YikuEBn7UygXBfvbU4cHgkUtyf7OrFDISvoaILgUJHFlx+fMN383iZu4i
MI8RgnabwN88uisMi8nbOpiUs0HCSDK9AkWn5xFl7AZhtrcZXqUh7nOzyueVfp3iiPqA5Ik+lTCi
hiNLVv7ChbxxomRx6tlMO3ztKHVfldl0bByHConmDFlgm8H7N6OjtLZoSJRVW9+MwGJEIOYNJmlE
VV3w3LJJ56/b+1YK0XicysKp888sAFPTDuLYM6JJCNEnCnb6ngbG6lX5LgbO/LTC5Iyz6NphbabH
Ebv9WE/JNDbiCwTTP+IDWJorbjNy9j61uUc4bt/MlRvXaWudnZlVAR8XV5S0iwl9AKrQAQIqHWUD
iNihYYb1/rSL8jmDc/eV03FHJoazMdfolril4wnG+UTLNion9naZsD9KNt31inr4Bdv6WOhPoyno
sw+tsRNFUfTfoipvPeDgOEVGIIk5j86lE+UrCrVyuI5LGaa5UIG85MFIypyvkfVPFHlSIz9T4u1c
1XxNm39B12KzW3BieDT0Z3xTukWlSM4EaXSau5aBSo2bwnhUXRBCwApssB/UuOyTe/9R0KAebw5X
+WDAkR/Ak6m44j4PADER00LFFhs9UpI7nKeLxjH60ggqquw1J8loc62vlqFO7dKyTsYyBR0aVeIi
i7QoF9jHI+H8wNgzom4MmznM7VaTPRvcQdgC49RcEKz1psbupj7cuS15T6q/Vr3qEu/Q6uZ/PStf
A94QUDoWwOMvdO1CAc4EPc/sjp3z+RVH57pPZEfVC0vg/PneazcNoAlWS5UXxtutDx0PbgliTNX2
zUMEmrGsqFKe9Zilys+mc1rLg69kywcxIrppMNi50cLQ/uxtIsEihT3AlkooX+pEi1D88Fy+q9Va
vKQUHZzeyZitJEezZDFTuKHmmZ0+N779CZi38YbRQIU5v3pV+jNqxrpsjv8AH9r9Y1cC+lKrzPNH
+VM7JE76JXGPc+FI54n2Ykkaxv729zR0JFTl+DJJ4VGdncIDd9YkW6b0UIIeHDd8jVDH2fbSEPz7
KFOhXNDdGRCAMwgPzbp6O9TsAttbd/HAy8SOlBKlVT0uDXGpiImH+mdJuOs7aA/T3T5Crl0I7d2M
AsPxa39ck/lYvMfJ31M649CWs6TdvFhH9Ar2P821DYiJqnj17RtZGF2jhYpOQw8AOhZqy56CEUX7
ecUn8qOhOY479YtQlQTonnYJ99wDc7KJBT8ihu3UcixbGpHR54FFIxKAY4GK9+paPvewp11TwZjQ
czOEFytYBx1OslSFb6cgyhH5FITI2BZeycf2eI3URPVLI9pvc1Q7CNeGkyTEAMPh8TxcPdMZmUQf
LH1RGh6yaEe+IsJwzuZ3eUDm7LJ7V9SrzRWkqxrZfj3R8rxXxPJzsX2U21JD/CVFLVhDgehdqUAF
zJnRt04NfgHMlliF9aE6MoVaYhWi7Rb/JmTEaTdH1vOIhXaXjK6skt2PGRYUUtfsBblHh6M/hbKw
tmsBd7wnhyKSwWzbgKNu8ecS7pCZTy6adS1fX/NgBQVvR0fWa6K1ibh3y80uBUsywKNW2dGEbV7c
w2q0osVzjzv11JxoKXPvRLpCJzhiErh8cp4U/z0GIS0jnSWF5wPOEu3ptgvzJBN/0/qZVIo6i71v
WVnEgx2d/0h1k5qq0dx/gXH9kSf/S/Mu/5ZE+dkKojdDmNruKwE58t6+dR4znhlFYJUWfcv+V+y6
PV631YaWu+M2PCzS9GM5rkEb4RKixyKih1fVbNjKHizYyCo5g+8e3otmzf9MYfh24kVTzajWZdSq
qQhEjtcqKMxD4oqtQ+GqRIwTn7GdC1gQiwVzpWi4tmMC2ZUqqOlGyhIpYH2z+0jXAmYPj0sXZxrM
aYx6mfSsSmA939PqRUkQRSq0INZfXDXNprPDEOU0TYMRqwAUIUu7Fthb9v5UA23PXW2AfQDhb/NK
zwNmaJQkvysP0bZRNqtHf8Uarp9klYtiWFfJ3f9zv0ZVu+eQPUWX5vpcH2yi3/BPoi3Cg6v+IteF
bh7SJLS6yE9idheJONv3WsHIH97IlQcFbM9++i2hSRGixnUVCKvpOVMO2t+7q4nNoTQOLExN5OeR
/mqtFHvIWfBzBDWeBxILZU2NXlUB3iTiSRrcPvWqmQ/Ov56KkADnWS2sWG5zMIuYEE5uZx4Ndvy/
FPAl+IdmCFNqR14yqFGeFHT9sizKlsKyznmI4RHeM1cMqtC4G1ttgPUQ4WblJ/rAUUG5NUs81DFy
nS8lVzyT8f4vQxWkcGf/3t69C1ZmZB3/BviW9cEbAFv65itcj8EMCrfmpyRfNFpmWKX4TbqylDJj
IcbzGvSJvkVr3eH2uoE9zoEABy7NV3Cr9hoiQu+brNmCb4kGpsZ3F5ZNU4NOOwcfKhzGYFuVKiZ5
AsNIGChjWr2hj8vh3N0cIsx/S9CMyy+k8nidlmKOVQdnwUVoKrwGnIZBzk13t/0I6sA5Xx/fR0lz
AuoLxb0n+gUcvvg+WnHBX9YTNTYlN0TGM3N+KhVzIo0rUFpJ58WUxIDOgynfsS8F7k+1ieRRcb5h
Rg5UNmD9VJvD0tKZwFRIq+1SCvdbIQnfF1vfIDP+tATwXhMboEZxnJDyw0tNUJ+dR33rMjbehPym
X6pZlNdgWyS+23knmvCTiJWOwKjtsSQrtDl1YxKT2MsiiSHdCR02TO19GyYkWydjHPJxDn09cDww
o/EoHCDKlpxjtVjPEE63NyjzBKuv/8BXTProfaUxNahvRmgWScmBYVweU65Aw8TfAA8yTDJq96o7
XNHGMGn8inI7OkReP+rIu7/wlSt3x02ItDDoiuO5Hw5SXChf77lCmuQKlVMYt0v5wN4VRjh6Pz0Q
T5wkFniDpjtYXE7h6c8BFzKXHx6oxVtF+siFmtLboTd6fRx02lxgFHJbdhed3QCTIzYydh8CIt31
0xRhqPLnRiYnzDOh3ZJEPvXiW3ykBa/s/k/8hYHvz0SUpR1XCLAz+VO+U/2Ejh4Nnt/LuPEObnu9
KFmPvrrd61UOutchVvQ3gxLOCd6+LwsBQLPClaDJW2XjeFQPJtJ+zyVl4J3bD8WCG8dBE3LF0a1H
6nDAyPsSKmK+0BiKpy0pWsaDTISfxftN0UHN1M2FJHnjj44PY+oNn8rgd+rX80nKq+rQ/QRw7Pc+
tZlYYFRBk5Erp74v7fE0Egsr1G64vFwWLa4j81CcDXVueZg/CYmsUjZ6om8MMRSPJRSVm6FiwPbm
oqyu8YYA1sWcgjWyM1jC61Z9l0zSNOtzdTCuxowvhupIRDIJdMNjcFD49jY0ykeKcxLy5YhN0Rt2
Y/KLz2SAxboAgA9ILxtVn5Eyi8LBRhvnUuV8hs5Qvz3wxXuM1dwPJOl3qs9guyq+Oa0KrwYRYcaO
3eWmV56EjUO+C8MERTABBz4y6rrvDoMWKQ6QDFNP1SUqbAHdqA76wFN9QV9fyrs6p7K2EXs5mzAa
D0J2TAyCKjb/uSTGEb7vxm90ibIiANmXfmUZDXvC6v12nVK+rmoTRNwvIl9eXc1FnBS2wj7hHTBT
TJ8/6Q/soWAJ6DOX1yGF9aNChl6vwYp61ufzVMDzZufP10HKosJ2oktO07m7jMPOF+W4qWyUVKzS
ihdeLeY1NcRuV3SWEp4sEi2CGD5KsYf3cxQwqeIx4RyHTMlNDjJ/XQA+D/JCef7Uhv0Gn+h7D32p
SjhQ6MCMQenFADhgqvtB+zkpR0+hmcizq8fX8gYkOu+imQe/q6FU9mbi/Xf0d86M8PLZkbdApxJK
awdvpqWzskUL6i/+wnHdeVvrSbHjfyITUF3XIJVBgYFW8lFFecPNP2EtbhU1qkbVe/A9YMpA0P1N
q0+YUAgalgdfeUZvLa8dXs0xUjwSLp2xsaI39L96jXsc+tUZrLa5+2ryhVMDHfPgrTlcqXkvqZm+
CZMfg55DMMVKIIW3FEQcoOIxLS5AkRaB0lHt1p59lL3GLIKMKsgKKoyWsWS2dX0IGTeqfhOg6Ato
z6iAtdXqpnYSdjtDpQ8JZmhRVBw3cfDRpPwbX/NpT+a3XMk7YLMJBVUfChWmX5lIKwIxCyfaANKA
EKSA7LUFf9SsEaaDZYHXByonoHQQDZq/wjNv6Cl/MPEnlGvqLbNyvgKLTCkEX8dfkUZjgXSpH15q
c+4gttYUI4gMeR9UqTQLr+gnltq1JrS+9SeX6CFt/596dK5J1F/ROZ6sqkYeEH4ngVL/14amAIND
TqlyYg1V3hYL2Jr4WaqS0DADbU2kbhryJBbkQS+OxQFWKSsS9s6vs/tNZDnO1dRoH2XWCI3zdRUW
0Ng08y+8jAricZAPuY0rszAGFN8mSFDSMuzjtFtGxKAl6V4UIt5qH0VzLrmOj+L1RplsUQNThFgv
1KMyR5I5ZnoJesW7RNqZEfkSTZYylYDwuoZLsiJ9ah092n09KOjnUVdDuvM0FtyelLxX6jpLisme
/zvxsbFu7UmUp4YVKVgokG7QTXnUZlRYfx1g0FzJjZMiNeCB7tDeefLJP4sE0m40rPr76MqORGBt
RLtkmXqsqXAnDmtS1Xs/tePydC6ft52sI1TumYkoJ/s48nIwAscCuPkn3A3UBpmAFsPYoozYom1x
Uis7DIla9P/zJS5Jkg4/03EFdIvhtkuh7qR7fI2P8v2/b0uh9ukV3JHk/ZO36RkRRIVKemCx+o88
ZYmnOWURU7Muiy7B54FkF9lR9ftjAiQjewu576mYx8aYW030WtNsVEswUEW/6GLs2uZK1A9jfhXz
ek49GSsv+UCVEg+KFlbeP053pjPFLuK2sDdOC20rbnXwLA0zbzrzHvwmzSTkyh1kym+zKdSm26ku
dY1Sy0T4e65siBst/9F1pGZaB13DAT8bNL5/y9r0DH16AP03UeCsImOIeMG9JfW3YOJgrBbiXvAK
8CKclfpirF9As4/DOiml4gXp+MUKkOi22pfeYnB5N+avLgq+8+/EQv7DhJJgf+OkjcYCFSNkgNgO
1Xso1QM+rZGvBFcY3eCbSpI8WbvzDLTji2Ko0MMsX7aZckqPvEGlF5WE6oUzeFxy/aqTLfFjBjhE
zHkV8Z7Oq2VpODDHVYDt7WnbCnnhGF0AvnCxkDWJOpOkAzvYHW9UcO43fFMh0AGJ9/l63BYzNCLB
JBCk4Ii7EBWYMUbjKnB3Bo6OpeYX7AtyUaEAIpWaOtS+iiATsZ+6Q31uv94DMym2hgrDFBE47T8Q
4azIK2VheADWXtmCTIz8PDXkNiiMunvcv6P9nKjXIiuy7wRJvSEiFHBgPfGZwvZ0ScGjI3uOemyE
SMQuq4XIVttF08qgy1U7Tj1PzuiCXLIGTO/OrxBGvkEQ1v6SGMwZvWIAADwnajmELt0xNjoqFST7
ge5LmzDmcVBKlE/DmhRhSkcEopHJritbGi1h1AIYoHCfUZcZvP9mA7U1GptLlU968NtYYcVgW0SO
upOX4gAXi+79D6lmBge5sNslRe/lfCERSbVQeOpo9s+BnrawTQ6XaPdK6dhME5slgSeTchhRFbNU
/BzcZk4u7+ndGreyah6Ac6kYgSQdMNYB0RSux1sUDf4h+Nkdvn3IDS1JTx/Yg61+dkZxXo2O+Gq6
iKrYJUDYr9bYxofLfQLdgwpftyx3QrdM+YzOsEPNroepQnh/VlLLlL3FH1TNEBW8ZFDuWG3PycQP
DQ2lFMdZ/rUdwJJGjksCBwi90WQRd8vXjXW+MShdYHD4DX4OR4uVoU0U2kDM52p/OVMHLIA3WCTQ
JW/A4qHF2P+DbOI7bzP2qQKDFreTHa5MQX6msJCte6jwE1etUPb1FUH/+2F92iRI/wTubJ0Sn9/F
W7qSpYXQ1RaRxd9653I1EdEtStrBiiKE63TSUe4Al3EyQ+azF03d9lia7vNVrLSNq8aK0ztXLtQQ
oO1tBtm19cT+1oHB1JJvWyv6YUu6L0WjpEuLXZJB7T85VfSCA39+MDqhyQmVFcU4EwmLNT4VcnVx
F6iVg1JAnNsUE3r1SAkVXGrZZEh/0PbJNeBX8yKbnuV38ATLSTFCG6eAKEdW9poMi92ZIcjW3VK1
ZSQgkHDoWSj7tgxV9XYrOOSy3QpnEjWgEls6R+bn9jEufbYrFvCzwb+qlnrSIRJHgxvaSAdaBmzT
57XmJKO57cqgqDTLEKeySgaB0Unspeh39QnWJNxSIegxTJ4YhoIRkMfDG9rP18A+FP7iniokvz6u
M2j+hYX2ZVOBAr82kVmWajvQi7y9TQbolGmqXgmuKVfFXLTHeGzbxmJz+gcral1/NIRYctIZn+6G
L63xxs8uP6Zjlxn3g/etOfcUIc3z3Ed17fPCYzr47Xq0wQpBWbMhWFTAivzwRMLhJZ8/1iH0T5++
XLG7Ng1kuoY2fkmFaas9CiG5cYbk0zu2en69hV9fxCd/M7SCIiwwBkM9fJn7+2SOQLntdQpF78Hi
vEKucc3V/lqZs9Gzkng7FqGUcKzlHycefRz3QFmfnGKymAf05qLIyeMh9AzLI6O3NsN8B9U1orPB
WWO3tWE6ivvkWJoL5HGQ1t35MadoQSW+EWDIGLmx0IV0GmkEeB5y3k2x54FFTsRqZWTu2sGGVOc2
ms9H1rgQBxVfjxhEkefKzE2r99iAb92KxtMAp1kB58QFDnTwlNCd6XqgkMYl8L9hw4QGVqjkdU7Z
tUhpS68OAkvEFhIsGFdWktA4qXDat5V80QaQuVRMFRdMbNVnqmPMf9ME8nSFRYf1RH1Wjco5nqhw
XRXqtEZKEHq4k0EI3rZKA/90Zp8AYUmH87u8ZQCYYnQjVFmPmNEKW206qxgN3vwDubxhgS296nxU
zXKJoUoRfLx9EiiPHTg75Nf1drjHU92sRCG3Fn/bXw5gGOPDJD39RH5qG2YeRS0oSeyJnhbw1oXh
TtHcAdkcn7exhRlqqp59bzQR1EuaN9TDE9vwjN64sIXkQKhgMW54FTXhICEiCo0MTNWRkskoCqM8
1+wzCJ7Ey2FRquaEWreNJSrPmVf8LezdK1eJULjxGQZ5DBokKljpyTMOYhX4iN37bQ2M+/6yTLRE
O8lgIDE1qtnXUSs68g9YhftGrlZ738M8L1nDJsiKlkTIwfqJ7UK1ab8CUZXwv/qAlueuFRjQ1KqB
KeGchX6F3vegX3eny4E3dn70BND/qNMkG0+wplodBOnWE6CG1Qxn8zY1JyqO6+XXiJCDByUZxI3m
9CKe0hqRL3WzNqUttNSBt8hzF6308pjjLPtvrJMUKpaztFVLsvFBUEQwuDNdMOWW0xNwsYKaCzPI
sUa0BQ3Lyp7swOBuMxcPgph0YygwmYXkwEQQpdx0VkXoFSjDna7l6cIRS5KMjZXUlK0Pcnyk5ejD
pzQErimItJFClGNRyd3hQrkc9WUh9KjRh6DpFsVc19Kn7c1hPUmIeJw1ufp/p247vSQfUgTDFjrp
5VFHBZtA4ohfX+v/rmdDmcayz3Zh3CMneziwYfyzNx8gTLHKMt051WzLxKgH7LK8NOLocuLfUwfS
Zhbwogc5aA3s0P30NUspb+DAybXEfG7XN0DPVxtuFg1FjzhN2oAum1Jnt2bbSqbSXChXDtBmR7kF
buJzE5SsY2xrmKpmKstG7CHvaLUQBEFzWX6QEahKXxWYZ/KNizy11on8FrzlPJKA/+7q3kzWnq/w
bsgYNBLg2/656wf007vvWKYrMDVB8kJObxtbPi28Gk9KY0EBzVDNF4gL3IVNRIAtdiHzTMInzzD0
t2ps3rmalQE4EOzO9Wh7x+TAARMOEans3h2KmS88let3SojOtoYCT+7/zO32bB2RHuMChh94iVDz
YckMPL6F8UZ+X2kSyPcvPzLxPl0tLIoK60woilleOLU3lcxsFhL1h+QfjqzXcFEidaA2ygY/1kve
g6xZMHZdpYNd7w/vZ94pQCDDRCeHFZdJV49fg3XMulGvMavj6TKgOw3Z3AuMGnIt1uqHYEfo240g
WH/xXX4VHuTLIeOcFfzugh+q6NT0sB2VErouqYhlC0Gm1hDYRpNAN7mWS1I34I5tDN9KNbX6ShZ7
CVISQe+EhwXnXgW6KjbdhpiTx8XAcznQ3eASoiAqZLvJR9S9nVAUacwuP3KJWaOu1KfzkLncGboN
C7w52g7nsYZiu3tBLPUYHuxz6VnMTNsFvHwoZkMPBwLobeX5/3oqcviojX/kFKSLfxpiJ1bUc9iS
SFG1sMEYYfeopwfQdwr9c26R9Ze7pLxeT4qNJBNXskPDd3ojADlh/P+0kQOc0Y5hbZPVR/8ZuAmy
IX4QtHYdvBiTnOlCwd3xwU/dT9Ql+0YnjbcZFNalOsmfU8s+j7KdOeUWsd503VR7z5GJLX5vwM7I
ikwCn7xTfBfC+cbDUdDFuKuxbKHpCMMYpH1SJcmgs3KPCmjw39/XJrq3IA06aAPuLhJgh2fTMRY5
mWCaNRRWDBp+Y6zw/wo3BAeHnNuNHloUI0SqaTw3yg2JmaN64jKlW/bSmyOboGrDKqrU3JqkPlao
sDWn+/Yv25pY/iyhsoNv8rCNH2KI1COwJMahDYJtqSaUKQfFirE5TJSQD6O3G0zva7Ox6RZ7kxDr
xU2Ws7JabhvTV1EeuaCYoqBQ7HzYokJ1vXDMdeqLjCLXYRk5M2K7jYSMITz8aOuy4cGLWlcM8ST4
wttfMMrMJXxM2Wzj4M+hIop3OwXaKnUwu5raY70EhRBTWGKKrsr0XfZrPhDvQ5mlTTfESjXaS1wN
+osjwkVvm0noDncPZ4N4XLHvYaa8M9/I2+GkrSN2jRQqQ+uAhwfMc5oDaV9a8elYivf9J7BntpR4
13vnWPW2Dy9yt++VzAt8emGLC+n0yOoW5ZimumT0sVHuEDx0vAlYNujfNuLyxJZlK2DUn+/4lVFK
y1t5gW/rvrga4SXTQqe7PZuQqOGYUJNasNYXHnxTke1RopWBp3Df5+WnGx9gZ9RIWUH3JRAKMBXm
vZaR692f8SsaqhaOnT+IlS8mrWBGrbHeI46Pr12GpaYPq+u3Cw/1WTgZ5Msxc7xYPSVVQ3KSd3jv
V/iY9b7QlwWjwaFGRXJNEDolz3gc2TekiijPudw6OpjTWNmwx+D4oEAUDYwjixChOYpPdfjILrZ5
fnZ3kSE//6qfHe8Tu+u6SgNAwYCVywgNJwbGH6ywnItSm1cFwzAcHVsHDO9EmuW3AXCq7ZSRXZ1B
YKbtMuua9j/hWsNQUb4aG+bOkD9NjlCtubwvtg7g7dmVUZXfG0ANxPsvODNKe04xjJts6ukzrPCb
c7eVkMYpVPTYY4dnrepGnLUWmVWJG8U/N2EMZIkw76VlsFSjC2n0TaUri0IrnYip46tBc0NcWNm0
yG4ZuE9qaoxHyOp8zz4a/Uo1U95zd8ON1KdWDPlFGmZKHiZDrsgXMTcg1aoViTCp5dNXqHB2SE3o
UOsaNPcr12qTsCzM3AnLFYbvcj3eBIVdlQknxqVdbS5kClRmdZp/zEMloQRtW3Bo7iYBKpX/Puoo
XLFRLQqle0TgIt9UZ7Z/o/s7MeFw00doDqkZgIsGRo95ScB3HhpXhoENmHtsEsMtDzEbj25UDApm
wlr+Up/UOPbv+XjRMTNBy4mPxIr4/DkEN4ZEQByA+1wS8O/ne2ltbtUaHBgItn4JY8DQkjAHxcBR
fsh2V7wR+nurMwCjwLYeGq6uscxJZo9eF7fRCjAe9MKg25w77xEbL9NnMZQXxVgremnk8tgy0lSY
AFaWYmHFIt/hwNyUeYJkZlpuZ4AjH1uyTUbGBj3GyqwcpE32OajKon0KpFDJDu8Z3nc3Mn0CyGWw
ZkDSq4hE8/BGDTWruTqqnL6IH+1mvYcU1I0DGQ+MnGWIA/y20ITUgVG/vuhiK8/bxlyugQL3X/iL
uDga5AomqCEE4RqxuC2uGN8osxCZ9QWvEKkYyV9jCf/jHKbyaFJVAq+LKg9Jv3eOh7xz8rgPLQ/8
RAWtuy+aIoAaSwqodP8EmwtPE/AcYcW4Panqdv+0b76w8RgTUJDAZOlgUHN9innTTxuo5+NpbMJQ
+I7q6VQRvW3pnErrAOCpa+8UB+KhHhpspgga7LrR8WNVtVz7dq2GVBjis8yRmr1vNkR7Ehz9BpY/
fJfV+1DR6G1hvZnewkrRZlcf/12jYPsD0xtgyC2ohZWmfnfcW6X8F0P1zFuP55t9hUUvZfwIs3JC
ZNn3cne+MYzgXvcTtjVuXGZvWF1XUqpO5praKWPyXcEVAI9jI3LRB6iRgGLJC6/Wqxc2nEQmn43M
iruqR9nbzJStncMTO/N5mniBK3huRjPqKeztuqEGA/v8MWLpLV22oGJ5NirZj4g2wMXBJTbd7+4e
GlAMWf/O0eiBCKjWTR9fIXA8z4vpKag2H7ydlemrfW986Sw80rraRdQFZcRG3IPwtoiWXCvYCwNM
zF/SmoZtfjcqgqiWQ4pBOyp0tEasL3vVthk2YOzDfzwqi6JSCkdFpz9SldIBhQT9ebuAakMA7GCR
v4wiIRXnV88JLkKRipGf6kjyOcpp2FwMnGbCCcaQzto9jwLNFyixiGuiIwkoVThJQANoIZ3bO2KF
riT6W4q7J/xQNMQfOzlhozifW8EBcXsK00Pwkb+p61HwKMIE/ezuaXWid7iRPDhQdfTJAcbmykfv
KzCrD2p6Y/2YQA/a0Yt8D5wJfOnLYRVjoA09CrFa+gHkn425h83XlvFD9/NbMEk1YBi6llYCvXYA
gw8gs9AXuRQVs5S3Omki3/Jzke2BKh+8iGEHvqHclyoUXsn7RvmOfeYKXKDFu3730R1qnd/w3jl/
j5i4JJcd95jEd/dZL4U2kzc/9Y2/ninrgz4pH09N0YqbtGHxe0opZdqUvOvWh2ASNXA8L60UGvwK
wU9f2V5u+yOgBrO5yXDO/FHDNNs1+3oVt2/kXw97QK0JRVE5anjYHYUE0DhP5YJd0Qe9XfzQnsBB
tnSAY/DNEK5+mW7h1e+ywnW8Ui3zIR7JtsxYnlo1i8wh9Xt70sszNQdW/Pr5jAsVsYp8LukManKR
Q17sQ1Pin1kQp1SCLBMz5b/z35Lxh/KswDSmIDvKJeZq4bhKE19IkrMFzMvGmxGygAyjwpbTwOlA
7J3nEASpuikPKZaFWB/cei3gPlMURSqsJkjmyD2q90ohGHYHSYvuJ9KVZNtiXL20E3UmrKgVxESb
wYETfj7ut2nl6nDrz8hmuI2UvxLsHhQiXXBiP+xDXYebXwW6zAhfdpiQMBQg9cM6SPajCa33UGXl
3b4P4n4mDY3QOBRc73qw4qP3BLW741rJ5wMVsM4mXd7r2poP1XAafVb564GicbsaPb19SNi1xaqD
71cgdMq6P6dcTMNohgwLujjE6QjqEwkJ0gEfmSk5NQ3GtGoDpwlMh1rzCp1nmgUizMPcJEzZTMzG
DYCMA/fwyOCxDWKG6Rgh0Gv4J0TFcLLKWQs7xdie93B448W5OKYLttTufqfX0CafxkcIazpzI6Hn
XqxXb0iWTExDmDL9Gmz2XzVof9AAJio/unBCVIIc1QTdRBeAVIDts5uycPIcsvV7Xg+J8Jb9rNA0
PgZl8CPs/qKGxuU/onuMyhZEZQybYsHwj26aKTImC67B1gfvlBBoYVUkP3t1ZJxKc5syFoIhVbxZ
r02XHJovXIWvxYcSIyJAIeLuNI6cPDNT8usb6rKPZ+llUF8HjPqtBLZpPxihOsgZAJEBIpRkVyVZ
Qtmfr2tn98PymhRPeB31+GVka51+jrtOANZ26+Fsem+jSPsQjPsldRcxEPAywVKGE0efVQR02PNF
yVi9rKfrq+wSuI3T0FJxioBcklcPK848+Puq5Jng2TbMLG4nFjSbVV66OYAIoOMUX4iK5HBkKXwu
CGPrNnALdwob82vuTDp2GI+fpeGNspqNsh+YlKw7I6FFDACs3ZVVdEWpJN5gn19EExJ464Hyjy1/
plLOT/S4So+eAuURUxKYaYam1EfGaq77Tpkjcjrd4pcg4F3uid8Lb22ULQZ1LOQ3Pecpax7s8xkv
rMmQLSUwo+7neg9g+Qv1Wo/MJx7WKPjb8OZunG3/yD9dHDeTbIOCa3vFo/gHdhRTZrpOd8MLZtrn
bqMccfftBWNCQ/lbfEwBx1R3fvXniTBZP+89Yf4VXqOFXUfZ6uk8PZEmBYnG6q7IMXpEmE8h9czB
Q/zfcihbEr+sDN6x/RsgcbJ5TvikAguUrOgp0xyGSO966YQZZB0gB89A8mr0Lju31E5tL40Vi/LG
Co2+t22IvOOiDIC/3fguLh39ESAS+7ETWAt9h4I2I+eeEFMCbH62sqk/t/gUOw9ZjYNT09v3pP2c
4BXZGFvOlVrphsH7dWsRsOTlfmwQ7tnKdzapBYXJG16hP74XwSGjo+TkaDqI+EGiZOJmu1T3siVE
eXSTUdVbYc2NS8zobZGRgmeOR5J3Maa9FlRFq2mZQTpYVsj33yy9s0L3sHGoGPSwm5/8nz155D7R
AZhoDXT7lYk5TpM5Wrnn7r8dJLX3ojnfcYQkWPF6fU/3zNEihRIbhEeGNFLET2cQh6STLmlLmCnX
0K00l9uFqilYEQarFZclE1IJlkv95jIvXOwm2t0oFREUE/aPMfnZrEO/RyZahpIcYDl6TQAwlOKV
t/XQN7T5gcPajbBzpLnov8ItTupNvmPxpVuCkt0qzyyPhSX49mNGV9KIQGqjPkSkhWuy8uG8vr5d
+DO9sozII03ks9zqIA85SXy3r4sqkLhOsEB96XvPn1pM+xd+6KXWM+aOc0bYFTvoAedSj6yVu969
bLcOmVSxpDTX2LkQdIqkKCwzZhHFCRn5HPmmnHbRptZfpQtDcI4am8tW347kYnOgoy9SCWn22iFU
wWahN7+oSlvTDEd8rhFe84Xnd4VvvdaQISgGJxByri4I+xnp0/7Ta/gVf+V1wX75yqdTlrcA40Kx
hgbF+x11QMFoGshl7KHTgpgIg7oTUi9UcHF+aiCTuLROuOVMCvUXTkCw7vXXzCQd3J0G4NsySUdj
0+p7sy/27AvXX7tgGCp6GhUq4BpvvXujwJIVmA6FARMO76eIEi2MhranfIslyVLufU67NQhY66a/
zwVGovW8ydd2Jq9gz/LFaUVCjvGv8idCn/9NCU/WreOMBNjLXHYWgQtvBKsoFk3P5Xh8E+4aAGEN
uLvIdXmO8AnGNtDgGsEVPUhqFTrEaR2vhlzrhAlp/4JST7BimMh5qurdi8SYbAynh3F626BF+9R5
mBLt7MErqDUIFr0w5LTFmTNZh5c4YFH3T5M25q44oYo84XeQN3/qDSSjF1DDtYkBMuggFKb16jE1
FVrE/Ju6g/lw9J1466LTHYBatG4uSd4tg1QfXqNpT3DKw8qWZ3NxnNIu75busNp4lazM7mfZ1O5R
8JuIhkaObncNJ5q/VFpqdz1jHsH4/2R10cjQ/dJlW78Wvs6UgKh0xSc2ISiL4tkNk27beoL1gnxZ
fH9viICLf/md3PoRE8YBngZz1qWm1jgk/xrja4SDZLle/klUushbarCnuzS9njOvq9vgAN4TnIEs
aK89sHtgZ8A2Lyef7ZnUU73JikYsm/iA3SqCsnHqrfku5Tl4XnyLRp85JPbqK9K7l428bhGfEv6s
6oUGv55XXy0jbWkFDl/Zxtt6TLnyUrToIMyik1Lldqov7k+OLd1bzu3cqoaMNPofNu59uY4ibeI4
LuvUuYmuPypY/hQJCIlGdzSf4zV+WMZYVdQDr9ox7q3IkNsMVkOLIhffNhN4PfuraYGN0ZuGO0R2
WNlEVMU9iub78Z4Z5XvlPQ/ELpcP5fv1lKQ+zrehuRDo0+QDbI2ANTnkm87zfv1jHSvYem1FSc3C
sUKoJ592pRwM6t8OsPaBNr8iVsaj4ZTIqYs0K8PhiVcQvP+rXW2ebbT2Md7ezcHdjmTxFihLogTB
y8uxqZIYjhdSTTD7HjwGJzbiL0DybcrDI9w+mrCyRtJirkwDA3cymfvnFSYTHDYayyRzbdZ0GUCE
FQHNinbc0crV2BdgZgONbf4CsPDH3+tqlT5+Yjq0g20ltEQ3xnUtm+WzovRDLNpH13Y7WlyD/ZVs
CwaIGyv6JPPaB79+pfFd69VkSnQqJxfXUsu6WB/+D7RFKodh+X5sxyRyJtvCU0js8RddeWXozPH3
5wje8PcM9Aesr28S+x1CNOBOrDaxD6QEsrVFTlJD2iCOix4sh5vMZGZhTZ+ZR2nAwqYkUXZ5Nshv
SwTi3qvCgOFyYiekkTEa0imeR0/XKaUQq2NrrOnaJ0ORZfGgF+mfdAV7BpJstVT28VWr4kkqNgY3
vn4TFUYAPSGnYwMCRD/s6BPGZPb0qNY+BJ2c/8RMuhKyrl008JCLefIdjY8X+2lPWPR1Qn3qQXSl
x2f7jV100b7dHgaDI2RJUVBPAg8ZxoPPsTSairzDfL3O1AF2ec38Gye814i2RpqxUseJsYGK7GVM
8TBuBUrf9an/JaHTtpvmVm+vIThItWT/jvBLmPZsm5cTyTgVpfhZb7gs7Dej8uGUC3uhrvxDuBhj
W2t0tI0YcejXqK/3XOWrSA3HQ3ZEsPAakXfp4ki3asDtePhcoNi/lYqZHe1iPnHCH4n6G3R0syBy
ekaFrwmOo3OeP0EOE63UCo6+ZNPhT3oYg5bSezl+KH6LW/mP/JuD570PMTsxzElc2ceHlqYncDzD
GvX6DN1d2eGCalqIPs/oIwgYUtP3DLTecCsyLqlIu0AAmkQX34hsI2x4g29C5PjgUBpDUiv351S3
gDoJlYrU9bdCj4r06PpRZNTgl3DnU2oJkDi5eWfVWY81LcnK9aAkYilJYTjF7Y8CVPYLUF+hSjPN
lrLhBSenKx7j8RiziAq2jUof60rmTFaIDL/+5ckRQW0Gv5MuwS91O+qBPQl10/dX/fqgX6u68Xld
4gotlpiag4qb1BI4IrwSge6uBmXMMNCOvU1U5APxf77AZS7DoH3A/Ig0FrnPPMl4jaz/t8Fo1UX7
f77mgrmxXroh1b1w6ELKMFUpXglI4C4r3mz6j9t33ngdLgWifvCX6vCCQB8pus4TgXQjBPm2OIYL
qjsQEgCeI3l513Z3ncJlBxt9edSVjcEmBWRUFNKahfQDrtal2UNHV3YvCPThei20cd9RcYSBVMMt
qWIXWjmu56pVY+a/cqAXqQrodTSaAFBo21kiDkSHgfumkH+Gg16e/vNgejOh0EHe8RZZT4S+S7D4
e1A2IS87B2duHxVAFIGkgM+fXR1jiKDypqL8qwsO3BUA+UK70I9HGQ1spwNVs+O8jIJ6O0zh9vCn
4Yzj8nJG5mHfZo16GIAWyGiQZ8pe19DTZ+LdmzBg1V3gvoTnUZi/A9n8FKZoGGZCZ3eK3ZZceAqz
hnkWd3emaB2zkJlZjLdjkc/xDkoXrD8RZ4z91MsVQD/DolwwEpDRGABT+/U5bz+yvFxFZHAkSu2t
8dkyWSGvN8OBIWa/8P4WsbSUeU0mx/lp2cv98HDlfdKcYL9ihET8ykHulzT0xII40rEg8qohlOKa
WupkjJ1JLTpimMyhv0N0rGycg9ywmqC5WLk62zT6NsHU9WWpx+t6h7zfkBxVaL82KmYWoDtC7+hT
QVcfL42j0Tpr7gyJKLsQHOXDTVe7HeWlh32t6kTnqDX7UKEbd1Sy/yxTuT6pI06xJtfexF44cJhN
1KbFHbEMqW3uNmu1bpH9dba7LA5VGLxLMbj43mGY4PASTgjiAwuplHSvpCvhYCjR9mQ7qBe89N7n
zeaK5dIUv9878/tAmUGvT4qc337ntb9QCR6WjbucVeQPDeDzADx3vb/3UR7d7cdxNLOOwNnNeDzy
HRm0cNVeE471X3s2rtCIo5gG4dKYHZYUOd5aV4AvQfW0G0Rna0IZYr/erOrtJeYiu+UjCQIKXeUJ
JNdVuSYB89QNofAMLEzQpdwaucZq5qK3Og6W0JFJRqf/8N5pW9hmyOmEyu3OIT8DkZhNNkETm9PV
zzS8RpDm148uBH4N69kHgeMSEUJBo2Wwa1m/VLdN/aTXVi24zjzH6okj7GrkxE6xTg/eaFaydbYT
LHhiWpMd9aZhyrPKUS1on8mwQJtzFSy4Rd1IZERamg+LUEzNXVKeH7Sxutmi459q3XBB4Rb/vYWf
gNEcwlWqQD9VdaGyDHxEL/cz2X2meMisOmMlOxvUKAxeirAXUoMiZ+KlBMpJy8T8+HRv3d5O6bEr
E1kxDHfRDPmnJCdRHLoQ3MHASwfFEM6zsEo8s5bWu4K6sxm5Fm0iOsEUmycNOYWo3oS4BHIO8VRK
u0OGMpXKdq7CTevH3pmdE9e3m3fwr5zCkB9FWZ3b+sk+R56bW7zeo4LPJXG3t6dsgKmavX1+ivFp
QcjKn20k70SkiyiKil8a3AWh3BWJ3WR6cqSogNKdO3vB0P4RyuMmbpyp/QzitcS3SiTQb59oydGK
yeJ0qGernst0IADE/9g07op4hAOllhKgZbG0Lx3dxjlbQ888e7IS9a0inQCyboD6EQ5wMLaw06Sv
n+FAkwq878Tb4FgjjYI7th+wLTfUngFj4bVzTLueYwz8+U+rWy+k1gA+/wz0ppPv14Aey56Ue0Ar
BI6x7I7cWmv6ECAXJU148ERdyB+9hfSWXHhq1EpDj7Oh2ajepBjw1lIokSPiU/LaR+RtEzhTfU9e
Gpq0lD7SPH3Lu/MD1BSJWHplxlDeSlMjpg3HtBIjjudI1gxUE19mcK5VoJAfnNJ7bM6q2InYx1RM
vnvzfBnfCgrYapt/+7y+4TIgesE7xhGdGhm7OLaiKE/Oy4JGGGc1mGK99/lDcLnz2zTfXLEYi+fU
FH4nAkEfe7rAkItpXlHz4CWQDn+RvptC0Vari5HwxrYVKLZUbzlaP6ZZjBg0GcbovPWxoRzNTikI
LASGr/mm/z0SecZaI0t7bCkPks0qvyUdDVEQW66YDzG3Wr6n+AxjAE+lcWO3r+EiowTwKl4qXUbg
LfXRNNKOcY2rnZS7mPx8cT45c4U41/7UcOscusbEmvgQxitkliyP88w7LnqGZQow49+xKlm/lX8p
jlcaqve3TGS4cJC4DPfB0HMqtNHWTKvJ8Gf2gRanVLj+DX0wEMkHs2sclNFLY1r66qNRe3ghIM51
1kgpw+MOZT6og1wPfS8uLCHS8hufI8fpmRar6FUwWoO+gsWr6eXeevO7ZH6V1hRFn5WHGy0kwQzg
hW+fCpCttFsfPbTtWU5uZ0NEGML49ozbNH+yARlOYlXG3jWwvDSztFdtXyE+cDDmO+rT32LoQRs+
9Kt3pDYYKPr7CvaBoRgOTNaxuQhIAtKdlu8r9ECGy3m8mnx2ETLFqI+iDfzhrgnX9H5kJ8p8XvHC
zXEwnDPScs9YfiUBM6Aur0sB6veORsuI3FVyKVH1c57TcqjT16ZTl6Xw4JKvCf7ywniALor/Fw7V
s2zWNzRWqzY0mBup0mu4E/jn80uykc2mAPR7vLRaZOIpQBVM1NrB4UxvYslcz7Ucg9+LLJabw/Ya
nV3lfKPh1qTw3afAL5h5+Q5ZB3J4AG6A5wp6qU+j9/bvA6VSTrcS22rYsaWjqX/9XhnZHc4wBDw2
B71+pIVFu9Hct/7kI56/7uKVGE1lG9fcI3uX0CTSESOUSxLnX5h6bngXjNoiYNTQU6JUUc/FsANx
nekRwMa4kQOc7XtAAcxAXr6jtUV2F5O+5ViXBXMYEUwY09xPlG0ixs62m70ygPxdDdlDbWpiE1Ey
7AgQWFPR5L0mIakVi7KGQ9VbSTkPu9Q9nzGvbxlJeF4jjhpcemJr2tTKWEd6KQTXsx5LhOSnZcK7
nt9p4Yzfe5WwOjqoOnCCpk5hHO4s2B6SRDxR8e+S8IBOaTHXRiiG1wto9k2IUiv/AQRk7TEfyeCn
fg4A+0DyvQj8aR6tDcWEjcteq1U4ETtOSMo6JQ6RC/XAPUQh+oINJxha942Jlpuur+4mdYuBg2C9
lbjJyVhivVpT+o2ufNy5xHi5ev9advr2cLA70gI9/SiTJdVc9gxO/JxWkl3FiEqEnshW1Eu5xr2a
m9i2LH8kpdzarfxSpPaI1Eo2UImbzP9oJyQae5j3ofJUOH/8ay4Qd0G6YP0ebwIBG7oWu0I0nOTD
aEdIYmjWGoeIm4WFSufakteEU045b06xNiaBa0Hj78tgf02lcPhiRJ1JImDuBYQo8rnDJNWoH1Ch
sdWl4jJrx2tsCKIOx6PqlY4FrVYi70dDUTWK80vGi5HhRtZolqvQcQ3cPaGt5wQ4NZod9oWRSK8r
DwxJnOBRK5Vp6XKJqkg5AOXuUD0uInHXRApD/cQTXxr62aDeyS4OWKb7TpAjYjlR0zMTJcxGr7He
bxwIiMxvwk0S/fcSIewMroSg3ZmVyN0vfKRmtQJ16t2SyOZLFwAZvRXlRi9GW6kCGB2s1kScPVgX
Sh3WXSsxy2pnZZE+8kqcWFDy9OEJv60Pe8m6BtFhhp3XzKvC+3tNZRcdmVQTrTl7H1+tTXwUeLZQ
HEtILGyRRpPKHks0xXbdb5fQ2g42hem8nrKkL+i6iEbHFvKVbC7aKXH7dk1xvH+RP4cD7YyHjyrT
RxlqEd5hAS3SJctxDa8z4Q7Vt+PxVnDwBSEpwVZ6aGnql451mG/ji9meET/uqnbLQH9LgWRIQsoR
WVSH2YtNy6Qh85v33UcTapkzz7Jb1mMveuE9V3b9LbhJPwdOh+LGKPzH6MWjbOt6r2fzExEnaGsB
/lbn5RM7tPCrrsty7aUGTD8fWy+0E4sLLGVKwlpCoUP232Rm8uR2t+4A3AaMOfxeRyyE8IFEBzPL
cy5sNId3cTmai2/e9igBXUJZmTlc9N/5AHeJQfBWCajRnCvi8HRm0bRq7eBUYAuaLc9jFi3Q+Sas
2W5D3bKs+59y//oeXROGfy63ZE/lpUxc4lI4tgUG4tLULBfAzcnpNynU6GTb5T6R+P0gL3PPKkvt
9WJ3y1PicWx2IqtrSHr8i9elewt3cm9ekyECrDxXGTkVz8bTbtfYRSZu1w9DR6UUQyFQuT05rVC1
6Y7K2QChKZab0ftJZabwUO8pv+ANx/pOk326QKBu5K2ryz8oNb7mL6fHzK9TBngjJEbEfUYcGTJX
vjcPtpfpAnf1/TmeVYt24XvBkHdx9qINNMKLd/blNy2q1G/xUXKQYnkRX69dIoLqNlGHRts8iDZG
DhpFI49G7967HXXzyIk2uaCipK8Y3RMZL2FtP7YQCnysSuplxxFWSUqfTc4XFc9i6YV9fKVa6VFx
uW38EGKC2wnmCSLeypCgZsuHrJlTHgLLgRYekr6hiVHxNzWiSDR/z4FfrsmW2IfW9mF2x2zVXEZ8
lNqugvWks5kh7HoMv38iV+Y2u/TO8q1OyOqjDva0r6l6mrnls2DbRlr1r2h8kKJJU2vqeSUNfrzO
zEMzM5kH84FeCA6uE9njB3WeX4lpyXKRdetQyeRY8ktWxaW3m4ns09IirObGG5OA+qqjYXo3tXsA
zlo1vU1CUOgSL8LnSZb2qo19JqkfVaSkceAh6iTZPw/Crr4saiDeIVvetsl0LyQFOR2xTj3GFRYF
/hWCrco3S9aeON2wmSOXwXwslSEHYdjOPs4KoL1O5k07h4/9AM9BZyYNBIF4drk8hDNEXgFviEUN
hLrmhmTY/dtqVn3SJ6frvyGezHGn7MKjBtMC0b0TKiDC5RuaZABdesZs2UVKmf6sO36yUaxk79Zn
Q2Mqs42GNaqsdmZZtjFyy11zWWKhedWUetrS8ACKbDFGhccptiPVtgC24K1bqRW5xeYDCJapl3L+
KA41qZGuazVibKZHWrUeblnlLvDHOLyq4UwPgtIkyJIk3lJcO5MkaqP5gWiOPgFJ8DGxcQbCwmsd
z8vuXEn+7xkasttbbIB2+8/wsAadZOC232DgxiEx83p7EuehgxnjR8AuiFTkGey84shAmoGf9dCP
PL2OHXwmeFHmuD+VCi/gkmRK8h+Xw+TnAqRvdzxkVRLJAa75iKss3EKfKp0rKoC13x63bEdNZKdE
aPMU5IUrRRpSlyWck3Zshx7gK0naL6TFgC4XrUiy3a49FZ+H9zjeH8Y/XZAs2KhvZtII6JQD0x5d
3nLMaGYiRv5fmsii0DLGsAnYj+sRrFcPrgd0OkXamwgxVdgnLRy0hHr0QLemTj5FXGBnbWIs9ief
isP75ruhQErqQKzRY1BZTeYY0CAwTt6VAk+rxbv0crrRmG0VyPnUWzitkUsPMpsBNplE9yy0MgRc
i15a31rxPvziYvLBYC9w4fQaX6fC04WHTfYrLOfAzyIb4uuOhKIZF9HoMfwxyzfVezNHTNPO7N6Z
sGaZd9n0QHsvYMEVQDsE6xLSnMEVP/t2Xrt+KLadv9TqFMJsQqfLlrzXWSja3AJy6bc/tDLSFdUO
RtYwg6rXaaz6yOHvtyQmgSiQK+PmuQm7l8UNPf4rXEa+eSg03jigjx+sxqBUr5wq2NY3//8xwGKL
Hen3Nq8HmnfGFHMJy+ObbMjSLWNyqwFSyuDwPYsaz1ojuSKHqpInYAByMosvc08M3kZXEb1PMrPY
dBfjd9wrJ2/pSr6WMU3gPiDUppzYpfc/bEuyvsQJVuV6dUSauPOpka4f0D4pTPb9YZfWpXVoGwc1
PiJDoT/ffAy6LeqeNRiaY1mJPC7IhGEKy1Vxxyba5C5j//aeWi8NzvYl6enplkscm/J1B0JJHc+L
DdkqrxBC2yf98f3Xf7CrblZtv3syUFQ0lwEwwS6PyfYOhXUgTfiGL3ZQ+3fnJLPyHCvNhwF8SPfG
r3x8CQa7vWU0v5+LobRFUSVuRBCX+lmE14TKTD3flMc0YUdDEc487cVUj9FDkUeddvfN0LLyGdqT
uu5nGy7hdrufO75fEoeI0vma8VNhgfGGQ1FUe8SOyXOlO8Zz8bI4H7OB18FpODQsR+8vaUfZRrCI
9INg/hJ+LmtxZbVfDyakNRt5beE7lhEs3xx62tHtTGd8OgYJWO9PhKCeGLA8It6vVCzS2T1f+9a2
D+loAp6XyghGrg1dKjpvE+8/TYnZDGirmE7prJtbz8kf0AYNtAQuk1lk2OdqybpxLRpvsDGnrZyw
vWXZxDO848z3W/jpLNTsseq4DviEgYX3D43zUhvMYqW8NjzodKGzAgFtLVFLFgpjN0ENed6jf9dp
8naAtzVIQpjvrvfvQG4VqoYapZwCSfu+lP8hwyUBuPj8wEZ+ghtP+PbmmNuawym8dQIVHqaBUINT
wTVGEe9vYzJEOSp20Q2bSKBTlWdWTsw2NB6191iQvSP2kTVj2r6ZNJ3+2hls/a/80shdHaOjjX8f
Lhs4oj1hK2h+IIwG8EnJS8u7cdnxtmEOoSYQGLtbbEDJUCAOPn4HoUoC9tt9fs/S8Bk5U0+gLirW
dJdJGJYHrmLtqum5+DGL3Sw9lGF9XFbyMgO6FIXOl8AdL5zNInOiFBExVD884IppMbds6p140tJO
21gInefKcd+9cDk4qv8laYehdG9FyeUn8OFg0/byXToYShKU/qx32Wd4tIGn1Shlczjzyw94KbYo
rb3GT8frHQYXv5GBB8w+qmdc7FnlszUlUQ6u+ONu/2gPJg7tP2ntaH30wadGPLlC+n8JXUNNstNn
Fw/519NtDnIPW862aNVZCmGnPp2Rnvtx29BYb7bDtTy0ta9CvNWdSyjEep1CT1ixHYZR011ncnZh
DmOuqyzZcmzIW+RuWJE934OpIsOk2Y2w2hxmbRdkxORIFoQbLtJyjq+0OtWVs02azQYJcjErw5pf
L4eApFRE8OTHJQkUNUc1CltTdoVdTYLD+7xdOLsO/Khs0OnSAnpMxATmDFm2IjhDZR78RevZzto1
CmAlwPNIJy6ejfIwbN1aiuuS+hN9qYSXBer7YrAtijz0uoHpCMf2XmlCseGvzn8PpCPyq1ko9MIA
wCpvmE05tlBXpN61Vx/8mnT1vGrDlUQ8bTZP3DclJk2ddyLh1/1xSa/U5gAq/lb9ND+lquqTNg0E
8kg4K34pRGgGodQs/lj6l3DtnhUEOgC7XtdC2xxkUW4/22a3EHeacmnK2hOkBNJBrOWZ6Bg/X/O7
8jxEzfWOQd/zsTBBP7G2nKQ91Vv6nTlMm1NGqdPkiBiHoWcvYO0rJCKytLRF+5B4rmbmtIoh2Z6j
y2xs2issa85xqQGLfHYWNMqAOrz1ZFscDKs4YzDg5fI/UB9S24Vo6A5dRd3OZ/Wd6xzyOEiaM03L
lXmxnYd/RVHJ4sHuENUutj3v41Nm/0uRZzZCO1VcpJ4kUzT71p8JekR3inZoKEmoljOE1Y5MRp31
nwdOXVtGaBMYj/4kAWTlnvQxshogcW3FIaC4L+eTmZT7wrSvTVu0j2dfLd45TRB2Y/ThMiS9v1Fq
+22miPAAvpvBeIoOBwBxusDAFa5kbDlRmtFev8eAVFLppq7qUPyWrmSQIlfjOMsYcJDnG+8C5YJf
6JteOwcU9FTd8RIKyHWuJBVT+UFDfpDOix/tbIrmXL8vobF7VJctweiOn363enmfOUB70R7ThtZq
rMrBwgHHq1jKnCwdTNEpXXSa/PFN8uoAa7Zpne0OMqoukRCP0cr+KFMXxJk5L7h2Iz3ChbW0UHIJ
wtSsh7Mt/Sp0o/8JZzR5MBXHFpvuVNgEDsYdtT1Xo/bzl1De6k2gx43pV+U5PVy0WAOuOa9kG/qN
3OUlQkt4ubEEUTlTYqZklQlEcXxpDXg+ocIKc7ghST4hVzDbsUxy+4Cr6bQ+UsDRuTXf4GNQcvcy
5C0ANB5horDBHPfoD5b0OTL+Aq0qNzkGsw3kMOEB6lOuvV7LlZjbNl8Knuk7DVPX88jrReOyFMMV
xRjNROjDAQjttAJ9zzu+YkwqetF7EgdulTTypxNVF5MnRrT4ZlIHBtCCPcwTZtzKcHrpjqS6jE9w
Tk/FtGbvcK1vo+If3Xb0qZEIPGSrn5X01jHsg9+aSU5er+q1iep6EMDeEbnlpMqs3mkYhsyQzKQA
K0t07IbP1aFbYz5ILZisP5eK3VdF5mSMCRP2C9z5GVpafWx/7PQeLXKChLu1HMuCjiNv6EqiEnCS
rB91xKnp+S4qN2il1E9TEDOc5ma/k/ciS05FQ7uEggyK+rUKq185mLaQ1xjNJnpddAbCTEnaMbMQ
5WCPRQ4H6qB/KkKUb9w3T4ksEwUbpyziiYHdkfJ46/BWrIEZx4BT1C8l6hFmah0BvZBptwh9Qchw
yBQau5HYupCs+tPs3HBpqeHGLhAo52b9+zMcjNLkJMpM2Mt2162himlaIbx4YN+uf6yF3zajvi5T
oGqya9LEMd76wbZ3v3NeRskiF2+9Ho8coq0x0wWktUROKXvZtkpD4Zr8/R9TahzS6JBq+TR633II
vWvPk417nySOA7f1dft1LLvhvzchoxzRmDiXVAYPj13jCgAQDsbRBz/QlnQrW4V7LCA83XULSI4C
9Wl3LsvOYrKja/PXjNZbpxysiJzYaUqSbxOz+1X8SXFvOnrNWgzxNHsUSQoGuJxIZK0Uljjyb5LK
sez+dvTtTvAYgtGA2PY0/g9v8iZEeJ/whAl1dhqhkt8+ddl1CpFks5vINYmNspKL/tQiqpXgObdA
WNOGzgqzzjLS/3vnT3dDPrRxHP9T9nQTRXV46Oe0/5u6k97b85hZcpcyfMcp0Cw0LPq++U3+CtDr
8lTPhifNK5NcDA4PEWuYTQUosTXFIHnEa9OzcFGV/r9y9hz6Sr824+PwZr/eJgNkYqBXfYhggb0E
n/9Rl1aVZZjiPaEnleZykcHLlGi+cxmAnKbX8K0qFFVFbjnXfQ27lhcTqfklcf9H52A4gssHW9hp
iTrP5X7ZtKkY/GiFRxcfUkfxWQPChy5RlwVguHNFy+8att5udG95hOfQcriPEIpPgzopurTj3Acj
rh3exYCeVe+8AzPVYxmC3cQ6BZMw0cAF1Npcs90gyiTljzzWGmo/ZJHbxETJoBovDKenbiFahzGw
5pS6gorGn6TSN1TA7FAPcJxKd15PBHQSKLYQqK1XWX6kgprercxiG8pgm90MwEEdn/ZF6MtmKKil
RPwMYfGbrTYGBkhd7rP08j4sZQemG6B9TQojZN8ad1FnhaB0dSYe63Zojo2a/t8jiC0/TuvbKv4G
5VcZIAjuvRdwqd9eIHQVvx172zvcOdOpwS0/7CZmPQg18Ce2RsKiUjT3Oe3CqdQJNwlTKj3EMNFo
iN+Y8/sCQVgjTjBTUSRsiVSgIGpCyk0eScKuOpTtBOWfD92v/OY7lsdbU4zhcUNWYY+4tg90K3LL
xD3n8kuS3ZBARaoY1PyfFVtaS7UrapzKslJcClclxfQzmLXFQ2KmO+qowsZs8OmaY7U55B9juzgM
m+PUNUfeMyb5IJxL5FK8Je4/74A+m3ks3a12lZ8nhCvD2Orr1Z+czL/K6URYnm6Cz0wzsb73MOhE
QEZK+N95bHKK04/oSDh3CYvCyjjf7IEikGobVbGXOvxw8fmz+jwNpt0AUGm2fZLlIsoh4OSQrupG
63rs7OhfQY35yBPQEJQEN5Tf/2XNBRPtYtiQeO2wHJa82hd19tZYogBOuPWijAlwhXTHx1gDyBnu
9wRZ9PwHASS5so5O5er6ZZ3L6SJ1myaXPQb5tc5SKRYPg0GUbwXsGARkdPoAcmkSHNeaBr2Zp/hv
B4XpeQo1psJ1d3tk0KfkZQv4rr7lByTy73OtGp5WNmuCSMOzmFBE8X1QI6DfNHfWmJvT0zfbeIkR
00OniWugn3l9qygojZ6N74dxbnQ5hgozXWdY22fBLyz+Eo9wq+GBh4ZoW4VDOjfUdhqAdkgCprpU
l8PVuVF62GCh85QyfWEoaf/10tx1pqYrPyLkOvP80CaxQFA/cWfgjaI5N2hphfux8ldruJvnzhV7
VzoYx83QOPSON2avoA1Rcr0B82uNSs2FJiqot0NnwLhKttzXCcDenhZlegwXFKhDSbjVHIeW6YTS
57Cfjar1Wgv13bBWFSruZmqgmh5qqI++iu+o0ur6JYxyk3BcgJz03AHFuLD5Jgw4YqI58otaGuPk
VieasesUvYckDWGEgh2M+ZBHZRUgnX/yns80gc60/rNB5igF7WO4tGXKsDqevA23/Z0EOoljDtGB
nO1Vo5trv9t2O9jMB2D2aAmhdbRraaCPQB+dUCUnvV9yIuWCpOw1lD0ZO/8PulhlqnqLpHNhcqwz
3xzrcwAbI11UiDBMAMEDbe7Idhj9bpmWSif4lGsa+S0B7JtAwFy3Bp/VQ/0356qMibM78lGgOoAI
tr9ZS4B4DNPzIMrlh+3AiIU/wW+1SOiW7X7t3KrHqKy2BuZI7zZwHQedq4Tv8ScAeYFmBKkTABNz
QeOI8uJWD3PMyVuXDP/XxvtP8w5URNgaGJh7w352FBZxQUiEQkGpa7VqvBqkd8uz8jJSKV6Oih2+
+hmfUh/9HVP37kI+9V8qzYK+E+sVNHILOE3m9f9Vq8xIeRijAMlFjTa24Jc5fuM90dDWIytUpP50
MCJQu+ZAk9RUoow45BRUC4WU8nu7KJ2o2rOOY7p3UVfCcuvsd2InuT8Lfo8AkH9pYl6fO7B8yh/q
U4NBk1BUVLRjNd06KTiJe9+AQ9i68y0EfIYkPRdo5eSjcwRLtRrKtbK1MtlNCzK8m3NeP1YvQlQw
eFhkbHvJXk3uzSzTcgkDbqzzSaQl9yFel6VAleyWaJolVt7gIzOHhsKr+Z5XACM4V9nxYDBZvN+0
bQTsCYD9SRpeItei3ORnhEFgpZFjVgUt5xaDYIHJfEJr+e7GVojSeKu6y6SaQS9Al1jZfie+OJHV
NgMOb34s+lj7o5pPeWk/vF80Fn24kOJBJ4xeGWklgSRRrZhq5trOeGp/gaaezjzz/mp4AOv9egdC
fBu/uywMQpgeCr/MJ1GNfjotXRmf1iBaCKWAF20s8KsM/3+uIIRGbWqzj58Oa4M71NPchdhMkJDu
Mn6jUGa4l/a+tjkMg+Rl1/BCWE5Nl1C1WGic8wXHLwl/RhxkHYlEDAFwu/okoSWT9470nN+mrNG6
fgT6QmGiI3tdO2Ed+GUR39HxFJQ4V0huAvDc/sq1pOTEhdR9o/jYBN96z1rlHOcFoC00Mc/rNK1Q
nuOND48UOkWff99VtIWDN1UdTjjlmuTHR3NCJ6711lJzkPLP4QsPkBzKm00T8UD7rqo0lhx8Y2H2
3yYEC3BoyPsyTTW1bCVY3gmZ5oABOz4L+Ab85UF+GBbYZJGwP7iulwPPAgEglN+U3AKNCF7DJzDS
N6nq2dkb6Uw77TIq/NxnUc5Nmq5y1x21QQ7AcYiNk3cLHNijaHYiYPL2pqI+glfTtrsMoxOGPVaw
lwoY0+oIr9xBUavcBvkLaDX5iHhUHtayimQV/fO3NYISSggSq7+0y0gfx1X3Wg305ImmsC9s9lCd
rZ6tX6MLRbblvaswNjFA354Yoj2f01Gicxr86F/fqJB4f1kXwaSRD2/VTJJGyWCeLf2rdO0eojOK
UoWJTw9M8oq9bdcpWPPzqpUCAC6jxYmIpA6dokYpr8m3CmZ6mvNdnAKiJRR2qfQIkERoobDenEYg
Ersr7k1jap41WWvxwCgKCPd0SP4zZgYNo8V4rPOgtZsKxbN+puXgKBtkeloq854DHHYOBwDdFicD
TAhNaQC16FK/xYlbHM3Puh/9hqVBy8ArKt6FCoqElwpBV/QqKq2Xp7ZeGfTOkk85f0M621OkErNy
hhh4mVY1629RK/I54JAYRwOjdW9mF8dI4XzcYFP4RMQJHtD5YKJdYfd+TkNz/sEAVN2y88C8Ut3I
3hW7JNV+g8ymna39dpWHLi/xTdgbvucdlWXWkCdO1+KabWaCQHgsyIO7sJld7bnfuOztPghiS8gd
4pcuznJbWqkV1jBDr6RqAx0f1FEdOWb60BqAPqUt/0+GC6wMsXY3Dyxv2ge8pHxpFZhrXNGL6lIo
M+9WZpeUnHaMSjXs9yBAQi966sOSf9kma3ge/98rlON46Pvo3Vz0oNHgrdUMWUriXo4s5ipUBpV9
P+NoRfapqXGx+OM8DSuGtiOzoWgQuMUw+IZDA7v8KFtuWbfhKbPfLMZjlyhbYwcAdY2h/rf31euy
SgEmhMEiuk49vfivihNiKPlrG44+cLgWYvvu5dQDTLuGRujXs4Bnt1E96i48wVa7+jMXIe9siNIK
NFW36+sPM7R+VQgnRWaAKlqBJj8k607/6Aza/rpCo4GmKtePxkbIz4fR0xUq41Y9Ya1GvrPqCM3c
Ey1aXNJeVgmlrDWt5XqWmn4LqTLr2oJVQCv8MkrshDtIaIyi5crUyUHkBpVMpEZD0xKY4PAsFu1v
RLYGccsOGdnlTnZHS7UX9/fA3TENfdGMldBe46ky79ohXM70jlARADpb7eAAZBchUtwLVHqaOdeB
VGZ3fAkdDwC2/xb32TjjP6LogL5VxXgnyP8hHm5stBO6SIo1d9sumwypph1fPAj3q5g8zc2OBRbI
E/OY2iVqfD5r8JFVWoFT7CIuQkC6VJv1icepFBU3+5usRaWG6HfmkpEGrAkEnz35iakS+u+yW7TC
V4sLkU3jC8V0EhybSKPiEMpGQBAhYv44uCh9nNEI7GEzNvM5wKPMBoYG2leXrm501X1ArgVjqRxd
8FsnkU0yfGcX1IkSWkprs1mhHhp2zHodNwOB9x9keQ6KdSHMCFlvsCu/OP8q7lUzp2U2BgX4U6Xf
mCGgsv/KsQQwcIpU1qUEctQRss9sG1/S8UAt+nqA8ODk6fHNXyKYDH9k5r9uPAdGcjR3U8dX0E4i
KCOBf6wScYGA/VPlOS2c3H4BYL4yXP6a/jSKW9xHW4RBzMpvZKFCJA1C+SZecoCMh9MjILdGPtgb
/NMuOdGzLE/dX7EbeXyk3Tiw8YzJJNKqHzLXv/fmvwDkjbWqZBR+DKrLpT680gtjsTmbYMcIZ7jp
vsFx1CKcJdWmALUL5rzrU1B8h+oe8Ahj/sJrCYsHnhWBaoGLgIvfCT2M46aoWPA59bA6BncmAhru
vpaJLDwAVgcuq59iZs3NyALMVJgpkZ1QCn+7NaIx4wifX5Q16cI8pB8FvTNqJnQ/aG2vjdq3azUQ
dIpm60v1gsAIumT6k0B8/6d8FYxbXMb8oM1c6H0l6wj2BauAplP93nWJFnAG9lMXDjGSmAlD+zXk
FRsSqdgo7sOlIW/SpUsogUbMM+fKxOM+QdCCSwektT//764DzFrexPLSaZFGQfQXWh+oVc2U7hJq
1JAw9yGTBGjZWTMTy3B4NU4G07cSlVxeoP0otAXznE2acYUsLDmYLnPOqaZDPSTKSwXb7dDSRZfH
2TUHW//4GW4706szul5D8ZHU71M8YIY/mnOd292MCgIfswtDtPyH1otjuF/ag58byJJuzvQ3hdFj
e/w6b2SZm1ERnSabIaWp81NsARowIA6vIJsFGfjtgBZm2KxtqEhaRulmvEu1cd5LrYg5PImcZrUi
aS553IBoPP3zDV51ghNnO713Ft/1fm7V1NSAtnTSBBLb+qR1k8j1XuNnHz6g/Ke0QjkLNPvZ6YpC
1eVPF2UlYg1nt23/7IVETwsGwd8hYOr7AKPuCcjOBTYB6Sr2ZewBxDqYeP+mtMTRXHNKX70ssk/c
v6Rsp1E+jPcYi0UVJOiyBvbeQXHfHUr4fYnNdG8sPSV6MwDle0YMDZYWZz+BfeozVbSmCT3v6kOc
bZ9DxH4jGgnE5Fs7SnoCZI5XLptlXUHRnVTNJb0/KgeT3um82cat1U9tm0qy4D1L1XKbi9PxrBqT
Zj4IBpyAgsG88rXRbREQb5JRG2xjPUitE3WeQGkMX1hdtEeQPDxrX/t/7UoUzEiSAXEyH7NTQlTe
dRLKscm+4pAlzaQZmn7+R7PRwNT6Zbv1y8KMtnd+clo5+7WfWjL+YlSLNghL8U/FwDAUvIWu3W8Q
gNYFMZMMYwZwgJJLWtKYTqIFAYCJGBSkvDxh5hZHOp1zbXBVv7S25q0tY8WlU7oS8UgMCGgHA0dm
4Tub1M6B1uzZKQicwIvUms2NbdATgQccdPEo4o2dQLfTgv6z6grOIH9jpiaUCLWbnj3w3MIgF6ml
ldXmNspFMDbItvxS22uRKJgAmGYx5TK9xEwR4w7luwLkz5sTvd7k+4E8yj8qx8yfo/p+S+tKrB8w
OUajnFBh65Ex/tNDz8Nb8zfn3eAdAyW9CN0J1lbkkWxknTqQOmCDXMhZQOvDJqnXVLlb6yyQ4V6I
hFAkpG/JtUsklTDF+f0Dc/wpF/a/x4s8eBuXU4HeUg08VGUEsf1dCdmTvBFdNMM7onaUS8GpgGJa
K9JLCbaSjsEgptClB96BdLiyaY1hR3WjqQ77vEeYCZVpiqU+ZHTeHkES/YD8pTUDzbv/YR6bTf+L
lkAFYHxLIUCEBDsM27kr+dqoCdg2cgpSuFcFggQlU4em0FOHjT03w2glLmfLMSmwM5CD7War9Dx8
CyLtlQFORsvvrQyk4pAOKN/F2RF1+zEQcCRY8XMetaIqNXKP0xFVUjaUZijhO0EFGVcAYb594Y3m
ItKVZkSBYgg9Ve3JWXoR258ttu8It3w/ubgjyOJdlKELBGjO4/8HZxpSWN6wQar2VLNsK7qEQF5V
iMHLY6V33tNPAxUAXsMl62avD5XXnaFQoBFyzxW0Lc/3Pu0j82kCsOr2cd7w3R/J5Q3easoclbtu
KKc5IJzDwUKfEmqxWqCWS1j0YysA61VNO8okAHYpe9H+NWe8iSuxsrUesw8gvuDTxSFAMosrWUTT
KZ+bQOUU+yzR7tSt8fw2caARKNm95W32GVNxs5XkCNU5tmlo7jlZ0aPLleLp74QlGU6sLxZ+II2s
YI38kDHMv0Qa7r5BcNHts5J9x7kyBZIg0kuBGPYVdQXZT0xOczoIdnKshWkx7NjTAAHfhYtXWTC2
L9lI/MfavA9ASlkiHAuHqVARxKo51fSQevE203//vvUVd9Ff3JPFKmcHusCuAc7pCbvisB1BTYeI
+zhAy7d9dmbsTxPCBhCRcewAjnzRC4aFjOU9bAJGOKHDAgq4nkbQKJe8fz7MRZulIRMOCg/Kz170
LlDr/UzgwFKecMcoc3T5w2PRvV4YB+Tu0iKNEJx6f9Mr1BL7bktSoJUK+62vIzEc5y23N+ItrkbU
7v+PzSy3aCOf0LipgZWx4eGWpDbUKcpDk0Gml4oFHICXSXMqLhwSPnlTkIbvbgXmdGQy7/2KyJqC
BDKGL+FhmXRN0/LB83BN6Hxne7RxwtkDxD807SsRFcYwx6G31eTyB1jkFA3YX3ps7ZEv5OVDUBCQ
lOjQ2kI39cYaAgHf8cjcGxnsrvhMll0hSIF37uty68TepulV4OxHn1G0+T88OqZPTFeCphswzB2F
UxD4oV+vixYCMUjLpst6DhsJsmsUCz8Dp065Wive3yXLlWiQzbpZ2XHA20WD0adnOK40W+MDxBay
j2LZjMjaDjKqNNzQwILHIbB0IMPONWxOD6HH3jvgVuNhrUzOibTT+AeFe4pVCLSt3DokXZMLTT2Q
p9ElNFjfuYT7O6lsaR2i0jBxgmrLEbP+6x5xKwNBOSMbAa5yvOKojPoaC3ES8h+qtbEdcjRsujkv
ctYkHMi8yzowZAnYC8znmMatNS2Fp44Pz0s2+BYN3+i4VvD9460L2vyOegLzJ05JnJFEYd3KvSBa
OWw7VVtboC5Phkp73HJ0ndtdrQ1XOVn8pbkOSoVKxV8TBFOLxMIgqSHGXAjV0qkdpKTkSaFPP+8m
BP2raL1vGnibjfQQruZ15WkURxZN7K/OnXxgCaLwpkfu3iuhRGmBSJmZVvCXjL/6WSGpdxL/beHN
p5ff2EZP88MCFTO9VsAeBEVUr1LWIOk+XtnVLyWM8jHB1ZId5WaRTusPSYv+Af7HJb5MqOkFbPaH
leXnVihCcQJb5a8CXVZSPD86n/pZ835+7B4WqXR2aIR71yeLvpH/Mq+Ix8AAK6xFi4+ISbNM1QoM
DaAiVTLSr8GgxYq/SvilHpCEsLrYlNYjBtbJZ6WFk9fOai8cv5AGWrefDc7QWauqDZtZZtH/5NDY
TlqFdKk/NFLGSdYIr07j0a/o4AXKYDH/gK3ZZxYVYtWrkyttfSKxEGnR2syLefd0MSB+nOe/IPEC
ScmFBaPpDilRDVxtbkV2zr8VBaCkB4NKysxc5uDWYnZnaIBj8SLZYiJ+P2gXAkwvQsSjmA+4/+sE
aP0a1OlxTc8O+ufcmgFkd+nUKyN6x5SWHFyAbWp6Z6ZwgLoQoQD8SfTfHSfmzOn23RJB7st5F+YQ
J9tSQ4z5YuU0P8hb11W/5tUxQTeqp1vwkrcCELZ9pzNDgLpapB5eA9/+WfEgqGlAFPM05OJOElb5
yd0Ims60bm7lpFaquP3H8uQIaybumuDik4eX4CFC0j8rDzp9WrhIt2btw+Qy8ran0iP5dGAWqA04
crZLLDLZBpaSDGStdMNMiyni5NxDpMH/54RgYXhgKnB0Wh33xwPjTnhsaRjerg8PgZNhV5Jg0ieY
bduOlfjoi5gcVK3H6B4Q1FSPnGGzZQf5cIWXHhj/tUPe70k2Q+yUJEalxqin2coKS2/OyEq0jNst
RHTd5DDb3KFe3oOttte0KvoK4r2Cnhb+8l5ES0XcfBEv/tuSBp61nxwCsx8vwhZn8q9EkrOKvONZ
a6m1PbftOh9Wx28h3NLuGKxuaKWvZTdEafm2D9XwPt7J5TGTyFjOE/B1Qwhwsd2nkF7wMfCpz6ix
dGnd9ftXC39SJbYHYXj25gwwYosg1GJ/1av9RialHSnDiiIXVLXTWYut7o3pbhw+mdIlQUMR8U2m
Mh8vBd4QtLdWhWe9PPrV5U2zZh3Y0nDvDOAfKe5YdI+0yNWYRA4Om070Hr8tTjBrJ1rgyzBf22P1
ET85OnVcoPHNJSYkA3AHVeCd/d9ruuXsafAfMYRhCWGZXHOJnZdpkPmjniny0NJV8QRklCURhbzb
av5yQI7aWz3QQnHrruKL/AA4OxTNruyRz215iLXjDMmJteyHb3mvndVOCVThI4Y+PojpaFxMVzyK
Fndnh8PxUh/ViTarqIwjmtoORW1P7wHKg7UqZ80EHmbfXvZnExcTD+INlv5Hr4CRjHHDmBaAIBO1
qmHHasRog3sRowsbmHoY+T2telQkW94xv1dcbbw/YPpF18uQLZot8pkeM1ayrGLF73BeqYrHt1ty
pl1UguvdT+efx1Ik9QxbkB73/ftXGqq8iDuLS0KhSL4NJ1lfLfc40kFezPGZmnaezyhn/9FURUu/
Djub3hx7gZxgZc/jeGxsBiUQEfsu1iphj/ZrVFFmgA4LNwatl5PlFCpDtjRO8QSBtks2Zw9YENGO
/6kdtCmHuupGiRlVkTgLaa1OlFz0Py0VWCksPIufkjmNCbZrcw+f2a5bVzrormdhSf/Iv9D2jxHH
9oYTyJBc+RHw7MfWgO64txy08n7RAS8hKN2rX+9h+1tfMvD3ZbcQUbpAe5kQbsucKSTFL1gXDPQS
LHiQznZEcqVkEUU0QWYfENN8CtNvhMg0OrnO2F+yyVBzl9hFVzmbqjwAmAoyM+r+h7IGBnDTNN2F
OY7SCG50KPEo9RfPE785T8FQE0hXoSrKjeKITzqyWGrNAMfSsH1YOLE2sacDwNlbBWphyU4pR1FN
aRbA965mblqzbk7cr8WsVLYxVfIs39qoxFexrP8XJSNAkR9f7eVxag/8YMgu0TeR0CDyJK1ohzJw
WTg+RgaVhNgc9BnZCQyvwTJ1M8QfZ5mxgUKw3tGrh9/R68qHE0bB1X2GZHJ++YrSqiismeR6k0/p
slFfzAv7DeRiFJDYYmxBDHesjx4i5j3cNcbuJSsu2LMs2ouX2dnzVfPvCMh5hBRXH9VRXCU/uLSc
dU3xvpk51NA/fUqGDN1QOpOts1LujY3qNVeJ9pcL1RJFPFb/qqmaLkwxkw4muKkxWYa301mmxlTR
lQlB06bWM6esa986S8IIsOeRceHcuYiua+jrzPn1naWQgmZQZTK30+dcNcgJLSOj7q3yQeCENSly
URF3uwqaIuUEpl30AycaFMoaf7d6xsPzmfFAONL56wULO9nwydD8fVWfx4hY4bz8SeZCtDCqnIUC
AxTGfZ5TUAWf4UAFUZj6MCi+EPZ7NKQuN4oKM1dN/yjWtqu4FN7Lk7E8qBz8+eVuPn+cF5cbdY9q
btXjSweVOezcEjgJg/OBwg9+Ma5BE9aDCIBXJ04ZvmijVtSh5xBhz3LvsZIgsF+8+nNl5dvycxhx
KKsy22yAhogfkfM90g5CahpBS0Fwgdn0I2q5z9HuyyyFyMXiP5OC6Gy1cvsMIhg95PqTzPq/8b3p
HKI8Jl5R76/VmIUdKk2UTXgtMoiEdX41PmadUiHaPqYyGlYe0x5k9+jBCFzV8I5byIi3YXIrZ8+5
WTOI/c2sYTA2vEbtrEyKgDJjOL1fXv4aXXyviAMImvOnL/H1WS1e+9sJ95xhE+YYl1W6krtBI/Ce
4lZacZJHgRCLEqLpTQKRWm37GjNG7I4ZUTjwYDQPGMzHnwXhHYqKjdSRb0TmmkfUAafLmpANbXqo
pkWS0BQQAPxiivq7llPPz45Iz6JudB0vVtWY27GvaVyLTyoil9H0KY85QrCX5wL9P55heu/bbiBp
J19UVJpzUHE2BdYjUWLhOhJRoIFcJzlhHe8eG+3MzTCJAdwzHvpwpBHQHhS67mtlS+ci6Yt2J6x7
bhx5DrsQjsv0z9i+w47Ow/jPeT96oAK/OeeKqkOSXPyOQwxGGG40yr70x0kcR86M4DuQxbNLa+Ix
gmQLGc2XC6rNDO5Wv3pEVyjVUvhnTnkOHuHZ+3cNWn3Dtw78Q0HyeyWbcoAJA5EAWcIvroEr0Aih
KnH1KAXwPL8D4ASWenzkf6uCFI4x2TK07VILMq0cp0CjsWmQwwM0dZtFOCVFGbq/EwOL/A6Myhsv
jzCzBzDVJ3mMetLY2EzjmUfSrOGhDOTJnzry/y5vYRPAiFUKkgfAggqlSiyKz6VugkNoXBa6XCn+
+vlTA8kYt78wYwOw3gIKQ2guUDHW+Tl6p5FsSqIxI0oedWDgrySW3Z+M3BEz6oANOd9GL4ZYdpbY
i3lep1sGAP0w0D5oA4YY7RP7bz8VSoajblopxxPKfVStglMzfEA17jVZvUF96vTL+2pCGo+Aaa6/
UbafZc3uX00qNm0mEcduZhcP+DNnFP2QsMt0pIU26PFWmUX3uEF2l4PpPJ/4xQwZ8IuXjuP/3ruH
tXl2gNfL4VUUngHpOsaNPYQxbH+6QOHAxjDUvODVIdkxBdb17MP3hHmSctLc1+wC7BDrTBfGqmQI
BOu7lHZgRUW3axO9tYns8uBSywEO1KsCS7nMGxPqqe/qN2xMgMqNd7EDH6tAaGmjUTQSdVd0ntd2
Qu+gIcg4sFicA37HA6fJOhH8P3s+RPBS9qPJN6ZL1DGELW8NPYakH8ja+xVp7rzIGS/lMd1EJ+LZ
M7PZ5jLjQ0Hutqa1OTnDM0kooG0VO/lJ9ZXRpqNDR0bdly94gTfGSeK+OVJ2+eHPaPvuDtflxQT6
CaK6/3zzl0FTwkEUtlVsi21JDknZdxyhltqOPU4NNQcMbl1UdwPMb6acYuoW+lQxGbUnB1pvUZWr
evZGed6yKEhMj/OAySJl/x/wUQFjr7g6SKwW90G1v5SiP0qUBHVZDCAW2ZFz/R/yAvCpb/d4Q+lY
FAIzoRLb8dafcA1aHobO5tu9tbb1hmboUojSjDzpYlUuEKKna1KvUzoxWH3k2kEE8idEHljssE0h
4PluT4Tax1GWbS7My82aSprKQoi0l7b0vdUX8viXrOZYK4BhyNOHRaW1HlwR1QxKBJXVLJT0T0Oj
7bGCyXsuTncEmHTd9dNoPLGoLAxKWk7hDF2kBCB7clmAwCZvfmiws9znZtHOdZ3nkCGMp7pbbkua
YhTSUOJW83iQKJ17eI8YURYMLAnJC60zt48+QYt+/lpAKEFW2Jm7m4r9OTSHNFjEv2rleZ8NVQbL
4QiQDYYATpj9KXnpk4LhKPw2skzQjWxRJq9B2lhlkOjSKXo0PwOtuI1jZ3dtkb7PBZhAaEt45s/F
n1ksBKituF7XiBfv0E5ixgIdSGweFCi8z6SsF3lDy4gsWdgx5m9JT5+zAzrF/riFLf/4w3wYV8KO
EYtk96MhrhVhpG4b0on+Fngn8i+nbzBIqIEIZ5a8kfRHuLnOXQZ5hu0ecsPFtpbAZgIeJXlIVbSS
HrHyq0ztYiXbbozb750qI2ZSQmpjRNLp18bo9Fmb6zLZBMD+Hic3co0iOvsymm9MIN70SoK41063
3TLu0ztFnqKQAh+SLWcZNojlkF8mjTB4uK1kAWervFSkRTOri0r1cqPHPWKfDSSDRMuxrGIGgnRZ
alOkhWMNGvRsNDqZ8S6bvLofdGPhrNwe/QhQzX5QKxG+XTq/wSkIQTI+OUeGTNARSDkSfQDOBGie
kOaHvw2lIfHuF+rzKO6ki1+YFzAEe4GUU70p7ZkMGY9p7e8vQ7HHkJt/hnrQ4tZJDdP6PkTRSxR5
rKil4jp0lyO00OIEvY1GXaB1MbgUTZncV231CXiV3RsOXdNgchIGbPP4g0tlW+TKHIov5dbWR/Dp
XhSqJtlsFWuaNnhzBAqH3AGvLq2/bp4MbbUwjNfFRQleb1Rj5h4f/4UtlPuDshXiKbzIcZpP87j8
LZYhEjzR2TjpPtIOI/lsEp0Bo5N+pj88x4Z9TWUASQxZ4BoO7WyC8jo+H/XEB6FdWh2aWaxOaEhJ
qITwfsbdWefKlSWfnzQUpnkybzCwOM1ldeQHESC+zo/7FCx3aF4Tj22E7j3AmoreNdwDkTf8jZjt
pmKOm1yzbn88QJK5Hj/N5b0pEMOjnm/R+nPZVmuVt9URP0pzxdicwxcaRb3izeupiqRPNmMi06NQ
yr1AxuOABVnhBDCYKd0ruMVd5YPLBqCOElDCo2V2d0yyx81Gwc7YdrRh34YIews9jIet3tvcTkcA
Dg4tPWaph5q6rnvzApdwhPvxXTCEivFwpoIMnN9zxMrq4ZIOCjOAdd6RDc5nsFpKWAx240/I0uaP
7D8qVOeJ30S5tv3N4joeUUK7giDH/3XGjX1E2TL2WIcfwspBFflcuU5FyG3PpdriiuxqJ3s1wBcp
j1BXWQDBGIvEUYGYR/AtN1n3WlWjS/X/BYcPWhmsHd1/1ZZ4Tn6qCAFhibUQ9NhwqnTUhyHi0HTM
Wy8QCY6FJPPwrF6iaSM81YhhgbSn/m/FThfJ9RIV9T2toO5WaenQne8qUxm9dYQZ7bYqIqL+CByR
cNgiSlgntJQ2LSAJkWxaWZqMUOILqtqNyn3Wl+6ldVd5cghKuwNtH/gU3GVt987aXqmPCETKp9et
1MJy01k4cBJ1ICpPhX3PPqbOFS+Q9f0Ts2tqyB30Jn5X7j7/efO7zxuk8gGIwe0DvpHlal5vFR8a
IRnNR3BTLL7Sq/uYioxb/PdpjhwQt2LyjIuo+t/fkpk+AidDT/uNI0V8p7cgWMhtBSzLY26R1OTc
UE2UcZq8K/Bp3mDoT8T569r8f3TUm81P6UIZeiRdf1wvJdGp3b6c/hn4woMcu0WOeB6rcFwVZJr8
D23wEom35IGUNJjxfAndHS9pboVt/3XEz/sUzWbtvAfLE6uzrH7qtPTvEP8fVeYARpwsgy/aMys0
JroeL5wZZseO3UCa6XG46nA39TqSTnlXD7NNCevBk6IJN9yc/R74D4WHGXa5L6hJQf3LSF3TvCE6
Kqh7r17TSD6i9urZewtq779mZK6F4Dmb/ZlFbF3Wu+O4anR9H5fXF0DGsp5/BuoID3hrD0q2l6ZC
ig8l/VbaNZkO6mRiMg2Hk1CAzPF/IjlsgqCHrG2eo2KbA+X1v2UDW4e4iQmDeXKsuFFiUyDaYYOG
hJOAYcY23M/4bdySskbOkf6J6OUYemXK0CRDJMKnAaeB2Ziw21IHAaqXE9KA0HLdlObMA/sdkw6i
uPYevkdaW7/Kpsbv5keNcPskMS57wWfRhwVeVoyEFFm7KMizXU4Xih5zTlY2Wsj7oujPPWdThC97
oHoqAA7yiD6rDGg4VI4StGAdz9xh8fYG2bcCt2SGb0CG/QzcBhSjf6IRt436yatDUmRDdzvJyRpb
Rzz1x6/e1fBfwNSi9GgPgo4ZP+z++yBFxOmHDOrRKWZk71RNQoGPtd8i5M8QW0m8A7JbJ09/GhpJ
njaLwtlXashNqwJX58ueT6uXFNxQZ06wbpsuoBFckXMJkP+wg3Oggi31OuXWRkajlxkTpAjMOZkC
46RUN+kfhzDOTlU1nrZD/RTwAFISsY20hKZoNbQagRFw/o/lpjpw+/lrcW4QJALyXnqfBBDlumGF
IjD93sgJluNLCdybtaQQHJ1fl9N7qNPJJBrMIFWKXW8/xP0bF/BXMP7Rc/Iv6VfXunKm+K7jwOHv
ksVINuAJGFRUxUMGnccdKVGoZUNIGSxFiadOCZYQRnhJqa/I5QlaDwRNjZt0mupFkDFpS/mSPibR
XphxcGPmzNaMeN7X3u7edPDPUN9neo9lGPisHzoEkkmTnfA6ZUNtmD9wRpmLQSOXyRAlaNyuNpOq
0VWTZKWuFyabuaLG30O6RdvyHnUvgA/NDaMSVfk1jsUTGrCEFxhFt2AuWv7HE7sg5PFJoKg3rJm+
NkLGYZc4cl0Pi/J1hrCOTzVWY2JvF5K1jIRrudMmAUO/4KVOiLYb5RR3z+Y2ggHVCq8w536R5UD8
8uxRikls72Qhcry5aKeUcKFCfGQTFhPAiM5iGirY9kPR4Yg5sj4q5wlmU7EzhJBsvTFLmc47+jTc
7aRtYK9FxvqxzAbRwoBSjqfGmNAQH/86SWmi3XsT3X1+XJRIGqgIjgibKShTDUQNldYCqfnyqtsw
GIotBTBhF6IdTN6L362XKWdIsRS9eTRS0fAsQ2PBIqkRV26dTJEHq6qeV9AWQq7h4hh+h/JjB2Jw
If5IGYe0x4q+hqFuAMtK1cOA0zMnImkR4RrvVHkAKi+2N28Nx8uKJbxZ/L4Vvbw6SgRMALEZ5C+n
vHYri/G8RioP2l1BPxVc9BX0UAPrYW7v0sSLqZDIbekSZsPSeWGBjYLaoj29o0et+cI+lviSPjWn
JsCHmOg9uwLZcHsqjhn3mfMpjd4tt6qRmTuH3h6tb0QjLnIJTHX3HPLwuJckAr7W9SuqkwQToQZj
QZ+u1QRwkQH6ob5nIU/xxmH0v0cJ4vQqB5FIq2WeTzyGKl5kd4LP4Yy3lLM54umuGgVpqNXk3P94
GpCM4tx42TfMjDkX22IA+HkKj6DmizIpALJ9eHPyPOQ8aNlWYhDZDr/y4nNVaJ74Uib9gMwHbEGE
ciGJtHEPGF2uNQ3oam4mIdbcZotjS/Rg71Ird2XNshsskf6VHlzHn5Tu6JCNx1tUVWHIf1Nmqx8/
gg6N125kU2GlCXSrDx/KFZT6KwVyS88woffgp4A6j09ZqdDeqCPjVSQH72Hxwgq2wpmubse2S16F
HbZzRGsGbCbp6nN0quPuQrfWqAsveG1NZUFst1AJeQRDzt+jqiw5juahZlQNdLc3WCF2D4M97IzK
t2fpCn76pqNdkH+WQ97uIxzB8ZTcMuMPbuBbk/EcXVsuENCRT7ByQYN3yMVt5gbqzsvq+G3gpggZ
r6y+DGHmDe9kJWS0XvnDqt0w8ZmR96OLe395Lz8+N3Gb9bHj4g8aq3ojt9lJcjLeIJYkNUMdOG3t
VuZh/VvIRnMj0zjz2iaYgkDk4aqtjWWINT4fjGJeMucwuUcwinW1YksRLs9+ksPxcdNbU+hTSHEv
N29MbvFbWkILpvWHEJiOHVUUl2YjtbF1g1ubfP1ZlI2E+kW2oOLo94loeL8IeLIaHXzmL962hlri
w5ygu7UXBp+den+Exb8Q3yOcxwNikGbeGJ/f3Jvk2XkKlDaHW9Jye/YVHf1jNco3j0ISl1jNSRtj
5f0q1V/mfvRJ3F/tfgxuywq+d/IS36xcWBpYENtuTnM3KBYmFF0rl402ubppKX51wXgYhOyky81t
QK5TLrWz5ZWxm7/VJNVMyqZYggtCIzWAXTpjUOOgHyQHdrB32BxmY7a3IIoC4aoeDguT+W2PI0vJ
/QJ9FP5ugFOMRe9wYBbGQj+3GYR3iSrN7fsXkAnM6Sqf8Q9HNqIY1UNrJ3yIqXHMCcmKnAo1LPT4
FrGoe6QSbsc4Te4q1KiOdyoHyqCrujI/cr5T5ebgAuXF/zW3icWPlRwaOXrDj+jaL8M2pur46pII
m9c7FLbXlu/hBud9TuC1FrtJJXC0xeF/Jxbe3cEZRMgPgTuy9vsZmPgV1ZSAwOn/L1PqiuU9UL3X
4bRPjlKy3ToFhJgyoHZ1x6L0btG9WDbM1wLnlPmw44qPxZh7+zl2q4Sa7dOPQkLWW4/zaBgUHYUS
VtRdb5Ia3UNVzbR9n4eIt2GDbJ1jqwQ0TfZgvIQWhENOpwzR2XPrcboWTjQBwK+UNhsNUpbAt4Av
EQX+JylNr6KX/oirn1yAakekT1KcMYgX7lo+4H1LeDeZ01jGOY47kfVm1ewVN+hbwR1v9OIHRrJb
AXsZyTWOiEk2+luLy8RvtNIko/zh5QZRgAF7GezZ4JA6081rcc1BsLWOPYRtQcpX9FxUqJ3dTa/v
2OcyF5/5J4Mi/wfhnTzmux+gBr+LvYL5exfQyhF7P0D8KxzZmb69PeF3hhSVk31u+NURBYYeO/0e
ciNkcn5hid/n5Xb92C316BVmD8CKwRAI8N1TMSr/fduXRpM6SaA1/yVHdr0HsKotWb/Q7M04f1l8
w33ME6Hj3W0H8htSXSiGhn1QonnZibgUggKP/EWJvNlpQ5N5FBdw28wXePNA57catdjsX3RQ43Uy
j7/wrj+dg6Va+hwGgcjwvF6dfLvq4r+Uo+7UBwF5jW2AR1hhIq4sFNoPmQogx0VYp4V1kQngN2hl
PZiwALmtEb5r1lfw4Bw2ND/fkTb+h+8r/mswpYPhJUE1L7SuqnP7M5K7p/hCvIwMLwJP2pNucadb
otOMsGZ+vebIo2/Dchlm/3A85OZTiA3QBi0cf8q9VG8aIdvU8C846x2fjyn04TKrkdFkYwp8X3qJ
fNZGOOC8N/dAB7iFKHRns4n/ZelR5InZrdAlG2ps9O9owlpWPUZzNKZAAsrcruepMagmpQgD3tEp
U9z2yNyQSipmftgo21RFW9KzkQoTG5wmL8F5lVqLtrxdZZyOWVLNamX56dU2e2fNpoFlFRd3QgSg
6JSCFBpuq3aF3TG754snyqgQfQk68rmTCw7u4AFYIDr+qHBIVjSE1n/78WMg+JYgiwVmAbh6n+gr
dQ2hMl9nc21PslrLcx/0KrRtc8TxG7oMcialwvifqYvkiLG4v4iKSY1CLD7Q3bRtR4LWavb52LZu
srDDPVxeDlfLsilu2spcFaHwp2uvrV/8Xo+ceNf2gPxGvuJ8OStb8dY+ubw8ejlNzpNlRFjc89W0
y+K9OAu9C/4WdiDu7bQlwEA0v0FCt3P40W8/NBU3pkGfTQ3wfjU1e0Psun3q/5rSPeZiPVVGHGVx
pO+CBLlEuM0jNfIfIu9FCA6Szzrrp85rovjirlatsMQW8bpv6oCKxqCBvGACc0mEAlQOVV/JvsxQ
Us2r+P6eRLPAd4M4aq88c8/mWIt+ZJNLIP70/g3Gptw3TrPIWbuT0VBEdbgZswp8HKEmHnUMXv7s
QFxbsPBLAf/F+qR17Jw4ipbx5ipgaq/y1gf4zNTDOqx5nLn8ShTrUxpMpf5pMKS502o4vpNNEkGG
JOTfynvsu+C2BJF+01xnCHkau2tMmq27qPS9zejTtF8XqIchOHCNWLjygUO6Z7LNyLaNsb999UmT
gvDolCeofoOjct1ZT67+2kotD2PisvwNh2XUmFftKbozZEV6+eXsGgmarHF3c/QAk7ygq3p/Yzpz
VfV6a87DGh28/oayjAgCI+xYaObE/7ImnFmAfguFjqwD/a6gEd5qTXHzegusPJrHSRKMvJK4y2jt
NtdZzXAjSnmt3Wvk03e3kM7EpFTO6b402RcQ5NnHvz9uGzDj/0+Nld+7N/j0IQ+sAoGCUdM0cnTv
p6dKBv/TlJ4U9Tp9iZ3n5otYpOb1wf4kKJkkqak0XPqB39h2L5ojzehUHK1hrAoNbHM+OrYRX+rM
4p2OK9hpwha7p/of8jFBef8RpgOWiQoAJstG5EgT5QEASYwK3Yf56jYCVHqbQS0i71iAJwp+ot4V
NawI5SggPhDzP107DxdQmRyJHnTCfVJqAcCZ8gYbmH37YYWawJ+N1WbnZtT2yFdZfiFllEj1qMYH
LUIU9fuZFRti5EiNODSVEr1rU7zS3/Q+HBdYKb3ZTJQbqKGWEr3xdOKPxLD+UfxVac1Vq4qxx0Ho
gJUTFN6xJrjwPT4XbVNh43sfRZOnHLYAEuXQXcYgxmRJhZNNuk9lqLLcqqVqWWTVTre46+dNNf5U
5w/O5sH9810DOcOk7zxwolnSBMjNI3asRgs7b+H/aSZDgWbpcqyA+imcdXO7zTNEZ3TEXUczTv1/
gTIL/bYE7ZaC71XvjtdmwKtBaXGvGrQnEtzyp+B6LUyKBmLhiZxYLqZ3rlMvnRWXdwP8t9QtxGou
WHHGng8br6LW6ZSwMJsUByObrKk8YLLSZx6iPoyt5t16W6urT5wsTf+8Ao8OAtEbtgixnALqCpWQ
m3YOOPPdfzEf/Jszz1qz4d36evFiqvcZomcZtzGgmpT/9inb4TEkHgNxwqrPm65TzTeY+Y7i+PFK
wlJgnJHc1DRgvrHKkGyoQ/tuJfjQAew2cnnSPUlNUqtVgO70rPQM2/1xwgWp/1H6mr0ouzTUBYBl
zOw0EUnUyb2qdByvr4tS81BCmT0jj27pnxagFrb7fgNDLZi/HImkjasmq2WS8o4DJ0NmeI537/x/
TH/RiZSnJinr13GDFKpi+PKEv+TlLj3LxsEztM8i/Bnf4zcRCmTYNly7Zd5Ho4g4qBrG3gNZw5ll
a920yoh5gFgypw3kZDw2p651qyDFFJ2lUksasZZhRhN+fC2D1wY61ykgiHgx0R4kYsR4a03IAbv5
0gxr8WD25QS9yy0PxsEqbRCBJI/AM1aNKa2A49pZCjyR/SsNPBs4YrxpdBChh/iHr7i3Iubltx3S
0vl1sTsPO9RFBGmyz+IJG9S1BQZWi9bJcE15ZSGHMPHravaGJ8EJo+KE590qIfIODgT4r566hs4N
hVkZHR+ZgWSq/6FnDjQQ8G8S27r323TdSNOdqCYiLMg7IjVDiudpWNdVONU1/OeUFKqLp8fcxHIt
G1M3ZGKRj05IK1PmLgX4bYXjrqjfBX1GBq6vEDvnasP9Qg6B3gpy1WmCVE7F35mJMGHFqOSKiea6
xqeA++BCm5xvVWPnMuTeuidH9I8QBgJHAXC8NkVYBwlXvLx5NSqSGKqv9cVmyLV2gR21Wo58giDo
lE2bVj+9/NfV9i/iGIkuLABs4iJtUSI1pFXUM0eDK+xml4/KyPBqWRkLad1Sfeoc16swzA/V8sMo
KNdIHlLP9/KRSOZzdeoRiwSTxGIdNNJS9MYOidHxkJfL8J/VKavhVx/rywE7ZnunRXjgziKKm7Fo
TFyr6WrjUAbEXFgtdscMnWapb3hPFGT8eJVPce1BY+PD9k9KwZ+JzT7rTur7LTGYtsuZbXc4WCkO
0YpD5UphRytWKrIbaL3bk6dhw1TIjFelp9SrEFaqsTcGnsX20Xyw/inKuF7/OXZpmaxmMSDXtZE+
zTScHVeQ0Zua0o5dKyo4fak2XyX6gtqPpowV9/68weXCxmmIoqYAk4PUELw+fRajkqleoNLNK0Cb
dl3HN7WhtTd/FKXPxPJh7S30kqQishl77/LIHKKvwVnr2q5KY0jm7GnNaiyYO1RBl15jM+jhSDnr
tXYg9FT/OYrPn3SyGJBUkvLRpvgkE3GIzwP1agXpgk6Vhu8wbdWPPp1vjuxH/gaLWWOsYAXjJJEW
SHmpPnDqjuaWZ0zi0AK+Bbe87ktjA6z4rsD+AnZIJ45saCtM7k2iafwKas/i75S2pCBCGK0SnyTX
FmpOKTul++2cO57blowYpxBMmS/40tLXbKIrVbJ3p1n7a462R5RxkNUk2LaKb3uqERNerjaQeLlT
fN+4To2HdCm4YMGaYauJJRwEFOwnPtKINORgqdt/Ua/DIooQIJSjAI5Rh/yL0zoLe1FvlZ1w/grg
W6zu9LbPJPdHY3q+dYVS9e0IdgMATpUxlBNS+5EXz0meOLv+VUiffjNECoOk5B6VQPrb+pxcpxE2
AQ4dHstNNsmBVbMgxyse7mLw6G6EvXw/99CxXkWQEQXugU3weRNC+mNsG3cxP4r8lJdRlQrE9ALh
1kPm7HbYItRu0YfJpwCqNuZGXv2ouh/NrBGPyQ53aSTB8Q966D5srQFMThVqKuuOOhQR17lFPbSV
5Yh0BjNceixghBJAPU0gBLJNKE/sFYgJyW/bf1k3hs8Pmbv1Hqhi9+9HbQV5UOVecqAkHbAuNoMj
AmbtJOZn44s6iID8R6ZMDI85dwO0D3icOfuyr1/Was15/XWmgIM3gzD1rEdIdKeC6DhAuXlNa8Kd
bkIucjAzVSlcAcgp9C1FtxBPFs3xCBUxy7OnayIafEg9lqOFqexiAfAN6F2Aay1mT7ZbMVmeI5Ra
yhhx3Racgcy9JJz5wuqKW7PnE6nKh88ldKdW76ihQZSkCJfSBU5w1bMT3XiVhYtIgnwz7eNQmhn9
5UpG4u1rSk/DR5AuFIOianEafe66TdSVR9rkHnxEPxw7AXSmiykubd01/oE3HTu2vdlhr88GCQAe
EEt4mGq0Ak1FLF/5vpdQsmcwctN89KWbABlg9NMM6MJUki2++0jHKpjlQNmspJRfxdtrwdFAhq8J
3BTSYmgAKnyEypQizro7aiXXOLxOejSWU+5z8G9GAI2A831f6dP3yO717rabzqm8xp6Ye07p+Qgx
UJSfICmPvtY3kT5yFLI+u7eo8Qlvg1c4I2vBBqSYgBg5b4j9LOVBmEz173+KsaiT3Pq+lp6Zrn68
DyPavVY4dEyOw8mmGMSC6DXnIG6oYAHIEUIgPsLGPV9yhKSS2qc4GVlOoR18/u+zUUJD4eDk52Ms
qrzfrquufA75sb7U/V1qA/Jquck5r0jtGQ4MyD9/EGXODi+TcoW3EnGfEAfiQF7hsFD5LAZUD/+o
3rEk6kaxJOUefeY6U5KOGn8jJWevpCEgMosDLPhxpffxcmowHQ8AtTfJqRTjvB4vdtADPjHlSzSa
+Gxo+EwAhH6xf345kHqfGa2O79Hbf1Rek9gXiYc18AyCKLg3A4s+N/YgTOrFtKHxm+bvTQr6qhsE
wUKDAUr8czVbTWLXSa/aADdeL8WlZNzbmTrDv9FxmEe8RwRIxmYvMqmN9IPAN4b1r+mEwcpmrtCM
dOBeJ0P/gj4T8yBU4ju2irARpcnze4hmsCP4etPQ0ZSBmjNJoDD9l3XH2ZIyA0UHO5PtV5yNJg/9
KAl2tv4mfptif2Vbk4GCDRXA3dcpIgK2cuJGZ0Ubl/aR/sgE8l6hpth8IRMVuLMztFfguv6K3wUS
OKhauUF+gdM6VFJoNpUzvkD5vYGExZWBzC+iDbP+mw7LqGqjDkOJ/drRDXD88p9alWc8c/Qtr8Vu
HF6SuvTcHW8AVA0H2LBw1fKyAZF/xuY1Sgf/dLMTiWYrmg/qTcV6xeCaFhK3SgQg3xH4kO82MSJz
gJ6o0j6DO9qtXzn6QBkHzzWBZkhvQV1bj3bYHoBT9YoJM/OPmygtKU4LzDhJSnnWa3xPYHLQfmMp
OqO7ISVDa+UGrJkgEJ/rjFTnqRAtHNhueC+mboWUeBgwNLmZ5ncb5D1uOnVrZeuSoByHRSMZQxJy
3r4XsufXupS1Bu7t2cPyDLb/jcp7S3T8TvV5LK/higrbwc0g6d5bxCX/0WojdFay8LAilhT1gUEn
JdtK8EcETi6I5pzo1cG1G5CsQ3uD7iZGWKbSE+iPsLr0L0PQGDnaKpYD6HmSsJ56Wq9RV/eek3Mv
8JJRC3maLQFzfeZkzBWdEOEQwh2vNDqu70wNTagvMS3nbgvGhqD3GaDG18aqIdzPKzR3bKwfeQMO
WHctevs3QjUJkMeYitMJFDNkyaG36TE8meZ7p3lP/Ny+Qaw763HmQpwyWflx+mKUqm8ZhJ9JWaSe
BU+0Jkln7XpSQO5gPJXHvhLJ6RbzMHK+4XvWgtENosaWCjBBHDXezJITzQ+bKjUQASnA+kLyoiqY
agB+W8ZXv03VYlbUSjDrBzLDC7jOkV3Z/Y03OrqX6NYPfs2GQ8umpJ4cfqUPkrIbNP3L+ftY7Qj6
DR2Ao6aja6zYqmyB0rbEycKigDwgoBpRhuGwBcLaZMbY8a4GdKf5JVYCLV1y+MKcf3cnXvYkxdhf
UNBjpR4sh9PNXp+XUTtRXZZwx3BAOxiFnWsCxm4Sj7/k0NKhDoAsyzuQYS01QrMudPSz4uPpn+uq
6doVM0GwI4y5RpWX3Er4VrW0KQI3bVkgXTQiEgnv5SzNVve7OQ4GvzIOy78lbGsrcbrJKOZiqaK1
BVTgGSLpmEoT6XMUZH+r1+ZKpesLPC5ObLy2p7G1R/DIGl4PepCl/iwiwEVH+7NM24zoqP0UseuQ
cOKBJjgkF6zeuZXUMFSBLxwEfTPpgvKR0zZhdu1g8wIHi6Q5t0y/ol96BzNdobfNRqWNfEHCqPns
JEbHHWtZXiPOH5+1udNevncLRwGBonZpBf4THJUtmm+SSfNH5XgecACuevokiFyP28Sh6r6vcMXU
X69zuUv7BxzGyC1DY/elXq9oF4dss6306DoAn/3+153mi+3ihueoQf6B+GTDP407LbOGHIgr66ks
GLzzvHwkL92PFiDGpHl8KjIpuwu76jVSIkE/7nZzFy/SOx7uQBNsks4ZQkmWRGkeO+9r+mxw4Ap+
B2R2S+smdv1qp63MnxszonhBOiY7xoT4jL7eOgBc7mP0C+Pc2P50XumflaL8e/qh0rU+GsQF2dYu
Zx1nX7Q1Pdi9NWFT+h6jrzZHuc9CCbrFPiEYNVsA5xhrLJPLlD9B+LAT8sHSkOdo+/nFwb2ShV/7
fHeh3YKk/d0f4GgLJLBnPzwXqqat3UwuITgYt3TdOuIXqwT6AlKeE17RvLlOlrFW6SuATW3DCQPf
+5IpArlp+ZlPP/LaGZIuN+y7kKsj04WJX2wqdUYNtsNEHXmz0VJloQuAojG8qB4yORdGXsOwmiwI
Ez/FWEu+V02JvmGrpm2j0SqXux3tB0lpKE8Kg39yGQkT0ePFLMLBn3jLDTclYIL405lrh5pjvwVB
ZKU9Jk8LLrSEk5sBgKwZcOocp7zPaUyPXZWfBjQAQwWZFZl2hLKObZQOW3otrGcclo4t0UUNo7Ss
wzMv0G+1K1RNcaGbNH0Zujg/QNkzgoYji5Wawwpnz7liv/0ZxIE9b5Tvey1qyZwmbJYtBkVOlr2o
jDXC9WwnXy0KtOtIpYSbbAAwuKAYZ+7tg0HT1cvvE6JB7dJfK0Aj07wskQbChTNveQU4B+PIXYLI
nY+D3nFO41rCV6/0tLiVelrpGLbMTm/owO0Dnj1h1vwd+yOncVmMzwTE9643nlPIUu+56vw9dqIx
ALd8lOytFenMtG1m/f5qpfuEHp8i4HQqFyrI+/hao6li2AP+9kD69/GfLUT4EgOiOxdM1r52tPbZ
R41iHGNVyOFLiJQyOirYue2P5wX6fJQ6rws2T3FKWipHIUV5bGdIdTV5ioEUHdDcYP7JRsr9yux2
yqauImgL9XWoOfis5smLJhTVQkqlrzVxEjHmhzj/40YYnUGLL5Yl98QT49l454s1i5yosLoPwwh8
1qYspy/2UigOEusSKIB5O2/RyhSx7tiiTwHiKi0+tHIjnQiAhHzVnpZbRoTGHeSdEzofwhAF0lZc
aUA921+/yRj2PmiyK6UGvtecxhaAQgxzFFlAtzll+4/M7MI+dsc+q2xRu4hs+TIjqzMyCKPY5YHL
BMMQrMRwILSOqVUndOJBOmdDgdnwdi8o3VQ+MwNSxPPeYsMW9RyfnYOAT45LdsqFboBxlnZDIDbU
8pk9eo3iLuXy++u0/XZwuNRvExSWiA7B1vNYmlk57maRHJY8zNMqzH8RmLAUCVgUHXf5yEvl9FBZ
w0zQWWVNCaXY34U+lwjoBcdEz3ID+A7UltNmae7Ukq5qbOL/5tfMRzDog1Ii17vUYFu/LfJ81XRu
3n/dLvLys0uxIToXQVIaAcxhEWzqGfyGml8PZZ6V87bXl3qmvEcCqUaP+ZhXknLzJMteqNBbfOls
eodF5Evo6gg6/nNoIuO4XxE6VqJTsdHfcIJEvlSOoJQ045HSvZLYWH06FGEGVUq/BZprTP18IbEN
CWfgBil/h3hgCg2BQzkDzpDBe/qvqDhSfMHRDemata8RH7lSpYm2uXmVEBZ+eMVQ1ZkeMF7ZiIIm
aczzB8cbSlXgFhm3G340ufah02oA45WPZFzPOw6no5USDyvGlDgdpyzgQpuYKYntt8YEL0pleXP8
ZLc53uk4WKMtoxzfnE4fks0Jwb0IVXkBrBPQkI68o3cBWuBp8y6ix0KRi+FGBVCnG+RwBkbQb7Sa
pI1VYZmYuwDTBfLHXe4lgrIMbb0MxfODJgiYeehObqTCRBgDNaRs8kxoU/s9qqedO8L7g9ws4S62
CMilKT5jkVYz991NhE/fglN3EdLsdAO/HSoqq1sQ+a+fIH4iePIF90GSQ0RuI7d4toh5hzLsUci2
9rDRNJJsn9XQ1IZ2EQHP3a4gPoJ6OrVVpqNQyY164uIc1LO4phyyuK2PxU/6+epsksGewM0TBsXi
t7pvnMCzHwiwN+m8HLVReiUswJkYcoWswXsyikTRKcAfwJRJpuOMiePDOG2tNeN4vMPPD0UG/weR
aW/sixle9IqogQ191BE9sogBezjIUgRoU1WHHg5Gru8CQueYxYowos2Cc8Yb7hKI/0943ilNRVFz
cH977wUZC56VtBRr43cYQI4TQdHePXLiOY2+hvHczTCCiFB6cH0BxehPCVVM7BSedXhPXgKuYIRZ
q1SmbBFQ4ZvDKH4ezCKwK5urOJK9Lanl3Na4trqvmcJ1Y/Duv7il0eBXpJAO8z+ligUk3W0fPnge
iJSCry0gOuid4bo0max7Zd5rW/tZH1yziMwp3pY1sLLvKRo8SGG/8dlIZFmnXhf4dBVOavqjyzXb
bSyKc7tnw+s78Z8Fr1Clpv+f+48IGvgYNroWC/AWJrT/EFPB2XcRGk0YGZwMKwgHoICTUT41Q/A6
oVrYXFk8ZSvKbDxsJ+R5fthEw6kOKCNU26OMnCRlmNxjjnIH7rNmGnQD2/XbQx3wca5b4PiwunpS
SNJ2ZQx3L4TI+SnCo1TEEiPixf4dhH5Ura7UZ9IVpM7maaUyHI2DHCH3JUiumJ4XUMw+8HKRUotF
c0oZsdripg2+hTIhSKGPUxQzTFYew2QDtxeVlQ2fjQeczAXAD1t4+P7RMyc6lteBobN5FhdrC5sG
KXUKyRH6PfR/P5YryCrHQMyzLDZryPRaW1kWHO3ysyYAYIWk9GCHV2icapoPxTM8GQGi3Y422CWQ
Is8joW24GNAiK01W2tRE/yY8P6SdmaHh7krleXgaoRnWa+TfwMpGhDcEKAB5Gdtwu/CZiUsAn7HQ
SteJyY/VDbgLCLaLd84lriBCCxPkz4dlSnsp1Pjk1OVA891CPTlRoPm1EKzVJqDjiCyEC6oag/SX
edb4YmRI7+0sgLZI1NDumR8zNOdo/fnklQX1BaNR9d9W1azhe8BIlWG0BPqVUG8FN0vWuKAoJhQ/
zYIqShjWsXIU5q0XB5Jc+MH3m6ULW3jZeXsDDpD18soJkdSJkD2D1Ja0G2wnnOFGV2sk/AZqYfeM
xq2oqBW/OafIv7xKbABpuy+JiJuf8W13+VsRyaL3ovMd2HKuGTPIwPtF9JuZR8k6bghf+HentRqh
lSKm3f+hHBsciVBjxba+sH+u37eN5/977o+I84GJm0WDTeSlmxSyv0oiJQYt5UXYyNgOmWAM6jCf
2uFc/3Lr+5bPAPHbOfraYKkSumg8MGplj23pysNxeby5MVMJxR3UGLZP9rY93AQBbIB+kcgVhDpn
OBfH924X7PrmestIxr88PYx7vvRb/Vuip8BLHIIN8L5zNSJj9IAWg6hopytWtnwQMiODvdMGD3Pl
LdnSAZXduG1YaXCkl538lyEovxmI2d/V3/kOu6pgrgM+HqpSBPBG38bkflPb2/PSJPIHOVx3GWkw
U6CJU0wi/l5o1C6+T4JjL+8wWQj41V8OIwQy4KnEmg0LWhm345bpFLemq8IG3GPV7PbbTwd74DYe
wRoBhK4DZJWskQr3sRndMnPQXDRPoZdv8vtjk1qhoORn3Ca9CE6qRAS98QJUDKgVLpI+w8QVfT0S
R2U1kCsZm2oZ2VpCZaF+ciQr0H4lEurgqFJBG344XREnzdNWQJXeuerBN4iZYqflMjLAoWDNmN6P
Z0zyNdvezHTM1tM3GbArWqyFnyVBK43zm34LYoi0yyp9WJimSYqfVmm/GgwP7g5YV5U8MUwUevET
T960LkTdS56d2IdCAO637cMNrAgCB/c1bxmtVENQZmE+KMkiWo9YK97lkOZOmFkLNUCRzEJs8qi4
3DtV6h6/PN6I9v0Wob5dT9RRpfpfOR3LrobF6iS2oWVdbyUZT9nAo38oy+dFAILq+auL8hu0LWNo
BURGBtzN/4PefOaWBWI6S+7oF4twLcdFGjTJhl0fpRbHeJCCP8WRqLXf9TsRwt1SZHVskL+0Cy+q
K161qyOvPEFDmXY8Xkly/rj602rsbWf7wMcyxgyGlocZXRu69zQK2285qgUR5IMFN0W+3o4XH2d0
uBfPmaUYkmi9B3B8MiPidruvtoqne1tevl5viRBuiZyIft+2q/aMppwmvPEzWZ0ioZt4uMcCOewj
ibA+RPztkkBYmhRuHtN5l7//puxVqiqOAENcLK3G9ARfWWzlipNtKNcdg9IiNcQ5YuebRy9gS2gy
x5VetT2hbbOA0q2nI19Gxk7S5JCfArksAKoCGyxTrIVz6ru3Ueb1OYu4+es91PW68KoqyY1b50YN
A8k1KzGqor5DIEJeHpFK29P9NP2pyvPh4QtICSxKG2e23U9JLJ6PCtyFr8m3Jn6pSGSbfbA8zBdi
Z3Q+XuKwePJ4vhYWbPEeRj5jNFJZ61rxR1ZSqe3x+HUuueL9RlGnEOwS7rDjiHSp8Gn9RTFqS02/
muB9t1UHVfUC0YnBXrpX1JG3xTDLs0Bj8afIOkWJOEAfu4RI/OgtIX4JA8ABJCAkI1OpQ0Ezagdi
hwAgBWylBWnZ+25KwVzOQjGoDtonnwR7yZkXhw9idjItuzJsad45g8CreWE+jHZFeMyG9EP6cRJX
yeQYuOmt5NvXwFk/XXCu1XmT5gAGyBzD5ycc2nlEvb47jbQYJiVVfasB9bzEPr3MaDuM9XOXblWh
6DtqqompXfMxFPT8NTvCBIbq45xphcp+bmD+UUS0tHMMGtDxVVuO/uNSbgxjGCtuGLrLoYswduGI
99eCD92vwLH0DOFixsvKB8eGPtvRune4wUpKWwP9Kt2JFjXhISRgklFBT6h4z2WfiLiGa/cHLkhF
YJItfOaWzvbLQDzwNqAKyGWsgq/TDFs1tKiPltkIDVdVLaCW+Hno2H1Asiq/rYKkGamGe1w2/IF9
fvwBc9QZGouQt664FBUNiya51byRR+0pGBaslGywvhfqtOz2rg6EyJaBGu6w2JzbKCS8JVGnelOz
BDF6FSZ3wwBLFw2xB5wkZv52mAhrYgWvB4VQJOlKAG4iZg6snOSh6eKPU9WXd/JltdlvJnFvSsur
rx1AVaq5xjTe92vd2lq/nhBYLkoleN/VcI9o5XV7USYahvXtEFmMVFzuuUsNlLgzVnZ2TNV27zxG
HafXjZM3dH4FqNg6YWattqvQ4E5aVZR9mFV50BlI4Au+bTC7FMe7IU/srt+8InCuqHUae055xkjy
OvvfhSQSPiiKmJhr3J8IfPEj/ER17rl8Fb8i6ZUD70ao98pL9IOlx5v0/2DU/2ivnM+rhhgJ3bm3
+Td9v5N8pVMK/cNHmzHg277sTJZX7i7iL04rU5ITSuopaSWhKqZM1f747v6IB4t0kq3Q6QrlYtCQ
S4jlhvZA+mAS+Ldar0+pXrnYBVniFLLp4tR5KDHZ0qrSX/j0or62vpgK2Enl+zolDx3rGlTaP1kE
g2GcQEBwH0wEzTH49b3PuzQ3UUB42Hlq/hoU5aHVh3b7Fjds/ZsoCBsvLgdPgr2c/A1zQvmoP7vC
jfFUKtSkabA6WYJnZ10qPXKwuhTNh62ZdZXsRakcfaaDbl8t5BOVOJDI70SEnBNJoD/muJTYXOGK
UiAH5kb12nfkFFvZPlfRmvSmJToePcHxOM1830iGV53agQVOOCCXefDAOapM/YprxAcEeyp3zot9
vS0JraJ3AH8WC5cbMWW4UqfqRGMD3uLUDki0A3mW0GzD7RotBFJ7TFcOaPPOYwnLRpMGzaLFyAG9
ZKQJ7b2L06sPtx7MdYD6Cp5GKZ7TKz56rDBtYYOmYHd0n2YlTpI66d9DUSCFNybTJ68YL0aCF/br
suygwX7KfWXPW3ETHScHEkaKDplBad7mQDWWpOvPx3DcFim2iGisN75uVC3QBvkJVAWsOeEr97m1
ekKEl+nRvjuv6jwJnVkPOOqPCBPX5d7bEsQtpbHF6azC4LsjQk0ANXWofaedvbtEIRUjFTlhfkKV
z2ai9osmjmNYWbCQGXZE3peBFDhZn/tbHhZR0D2VlyomjW4GpaCmQdmxQnUfSoKOFlSDSE3Sxor0
jjVC5qlwCBrQW2mTWjVYjYnCxN2GqRyKMZ/ANsxPqqZL/Mte0W/u5mj0dW3eNcAe1n8rc6F8dd2E
9cTMxEkee7nb+iIRVmu1hNjP03sAPN2Ep4UZ9m574GNlJUO039Wn186yQftrl1+/YRZy/P24mcLd
AnVkUlnHQ9Zf7LgQNiBhorDhAAF3M3xSvkUJV+Faw3tT2i7VYBQzt1qW/aCRRlJiBIM6wI4XWcVK
4quXuuzJQKxvxZX3qvEURiOQuZ8YfljOATINj8PZNdD10eSJqjOPQUgu/Tfvq/QskE8/w6vbWpS2
0TjunLfhzG1ZZKUMhIgKUaFOQ4C94QLoa1MNw1nNEO9S6PdIV8KCWSxa5VGSuYpiP+4joINbuFx7
dCX3v0v9090JmCQAk+dw9jSZYNNgRtEFhZ2ij1GsH8z0yU8JWWZ2tDeY/Yc80IjApO2IjsY6rVhJ
SeWWlAJCOouRP8Uezoc6bv/IIxF3uEgIyW7UTUeufjMHwo0BRyFnfk98qsk7iSRYcf8iFEMicD1W
S+GBiiI21V3IcYRbf0N+zhjQKLecLHRaLvH596Ax7d6qmlN+S5lwSiEMqP7oyzmCxVK+zZiuDCh/
vjzRxtC+a2KULCVF7r7xpSxbTBXpBwV7soG8QXlDVsemyoa28K+1LgAua6CvRMVEkiySuA93VUaX
Y7RhplMDz3JPMLMqkVlHoZvqdC+UKlraIrAsWqeZzwQ/d9hSn4FqrT2RFRJuoGwc2U56LOTJR7ih
WTa4hhWymjYurD9ZwXstAu7Qi8+cTyIaYV2RkzbikHY0lfnQpR1/1+OuhDraYVjKW9yEvlXTURYq
QVxBEm+/6TYrUh6xp+FGtIvzlGeXcuPZOHUfAOgj7PqcrW9AJsoxFHemHNpiHjMGDg6C9xD/7TYe
P9eHGbL8AgeW+WFPuTrQ4z97fjA0pK4mJ8OSxgRhdTpkhsCxbwikHReBWTPadWzNcp9zYIK7yS/B
YsIIkFW0eA8HaXKWdRo7dB49TCPubjx4w7nbcF7xgLiU2MmkcpsLjMcsBUxpQ2FjtzZHvoZ4sIE2
wFJM0gNhipGL8pH152Fi3TlQ+5P3Q3rVLwBkm53p/qGxeKI70UHueh5EZTBGbQ2u1zKBY1RZy8oj
eLveMLr0dHhSDNxZ5QSU6PuJ1t0q49s3J+y8u6FFOuHPWG6xesADVDd0b2QueNZMNZ/TPv8/VjuH
q44v7hEPXbtR3ONoJImdaFXn8HV9WZS71+m9U60xRgPzEn2gUYlm/qh8nhsdVW4TOFeBduK6ip1O
jdWggsZBV3u8TdMD1bYIVmGyLxonANJ0sYOobFQ9cDMBQ9DBaNTmzkV2+9BAWJBVqXS3ro56Gwuj
7T9jdn6XC2/slXNXTP0/v0iPiRkqnNah4iFCzfoWc6A1crhjG+zc9YlJKUy5g9iL0ZwtJWrUZvFU
mq8P6d1X2P6Xe5IbEu4k1eO4r34zBcjzxMFdzIBziPJ2qFPu7CjPmWuIg+Rk6rzBI9UW1IdIuwG+
re7eVG84hJmRYIpyys4y3I74NQhhEvZ25TLRR3ZJCMYUAq1ylL3wD1uPiR3VEgn1SK3l6zz8cg82
IuFDPbSArM5XqPVh02bS/MLJBnAB26TApn/FCHxtKj+mmO/6WivIeyB8Cx1CkSbxbWV+MzT2ZHGe
0UzUJfhxX8OED3aSoCL9ZteR0WOahwcxTlbES22XmEKgPfi3VHZ2NNZdMtdHUeeC48uFXavQSolD
mvnzN3kSgxZLEk7h/Zohh8GIjrpefccxY6EuDADJ0YNlhht4yqJBe0tsnmdYvTFaW/ZNlMWiSVso
Z7xq5iyIn23vPdEcklvqxKxQc6D0O8G7eXbTdIcx5SuRrIiesoiH1z4eAoUC8nUEpkAGBwtRdFXs
wSInI9vQb6+1yBVtnGYf6tUhHD/8uONaVIcrGuaGIZXKquoQ5E6iNe1/Q1gupEbtF/oFVRA0j/T1
Rekn+lxk3KNhYjjbJ+P0NN02ZZqToe0Y6/r1Zp4QTJCYpXh4JhRb1tLyOGpFKzVKW8kpOzPvUBrx
GFWsDNiY6d2fwP5BoALIUZccWNaBt0p4zMKaZhDjYm1GIsEmuiPUeDqsBGB+0DPDN3stHGGVL1RD
i6O+zlR5QliYV3jRbUa+0ZtzGfOZtxe6BL6S+ku/VNOyWkNJbx2UJr+ZWNfJxZ4MuNFLudCVYMsl
BrzeQ2Nuoi/+lywqDRdD/4UqPrCtWOBm4B5C6M/wK8EZ9dwW2oNFp8encSIV+Nk0eVQFe0lAtjMt
4aHC3INdvF313DkPRVvhr+nXWO61AEzIdef9nngpgnevhQVyi/1j5b+GgaTit9Ioz91DhvL2thtQ
fAzY6k9sCj2KBdZVEdAJcbmMfX5dlHE+m380sSizbniYuWH6aOZ93nJmp7YYx95vumsN5E5YA/jl
qrMX5rlUTWW0JedYrMUP4WXjoNMRaE6PLnT9w2n/+X4h8vfhlDkrClpRjPFx7Sp2t0m38PFjXl2z
uOb4jR2NfSV6HI0uIBofZ+mxv7l4L8bd1VSa6FoiMDLFBcKXkt7k97od0LE++du/sgrBidxqjk6R
q0663W/Dn5+qapEk/XDQjbNR8gwNBZAU5WnHutFqhMjCSxyiWYLWRB/l65G+LF49wpMrdZ6YouSP
9nJ1bfMcPr4S4NA/5xhkCVYV7Un+16pvhYno1WpnkHVCI2wD+Ac8exy+WV1DNFkd73dafPEoCMhm
I3uI0vlHEzrCWOFFVcmAeNEET4HDHmW5fZBjPu6GBZnT5mvgZJ3exOs9YTVmtunkrVhbM3dpLytF
E5F4BnnNWg+5pISvN2WP2b8JbucytHSvQSxC/z1Q6L0TlfnFMojwZj2nLEjPKsDVFpxmggydEOE8
b/3301hXr4RUtmqLzwVjia8FmTQ7XIXAQrPGvxK8RHi5MiKEtjabraGb6gylEhrvDDZ3nqmB0yH/
R6yXNjQtSy5xvfMxMWby0u2bns5RuzY07nt8qom43eY6pi7xCww4R2mf/11KSt0oQ2saKjQpDLkM
BcuS7IVSrKDbfoxMG6X9t6JDQzef4mF8VPkCKZljdo7k/4EHZPJ/bt3CogiiL4eOHB2nSaIjGMj5
6jUdvEjKlnsbs2j3xSdwHiTiWr5OlPTAjzEi79ylmG4nWpRRrZOhkziuW1yONOuBHAARAVwWmM0H
SE5l8DfrXBpJr3vysBceSSepPtTMsv9Yk0n+Zv0cYhmSvH++ciZ4lT+z1CNWaKs4XhlKwW8TUmMP
N3bwNifCgPqk0ab8poeDYmFOXxH4DqCOtSu1KUv2m7i3FNPnIE507outCOmq//IBX5aIjz3ihDsS
lYEsDhm5gHrZ7mWpU/tjj3TfmKBDuNlONT4Qi9jg4vwZ+6MW0uldF/IxNAEGZS+yMFR+xTtr64MW
dSC945t2y0tl8RY95ZD+u+jX58RgnjRiZcpwotdvaqnLDlmg38N/8MUZEKnwAFMgCuCPDVnIJIH6
H2z0bak9TJIUlIcuIkLUBqkmJVZvoRf6AXRoIjlUHFv77EnNdtQIBXGjZHZKj2Ij/qS1yAccoXw3
4PLt0Ilqmuj0QNvlCt5k9Zh7qJl9CzvvEkdVhr52V66A++mH9RMO0fYAVVhNjq7JTatow1M0TMlk
B1hMJC9jgr06MI0w/lmePMyeQYlu0w5+ouEfUjgucNQRi9jNtGCSHEKtFYZ9eMsjkiGiKfjvSEzj
4ftoRr7FRQpKRsCTf6ddCCrx+1zfUbw8pbUrViIc35DUU8Bsnlkb/vogG4hQI9Wd/v0UGCNNPzNI
BIz3Kd7h5AXRr57ZAKMxrN4gJ4dcUGMDEmafuhk47Huoxj2EqI9IbgV2lYWfZzcshj43GAVklX4V
Hxy9RLCkT1fo6MkH3kEHWvVCrzz8qxdH6vNlLu/rHdjO4RHA2K8d3Dywb3Tp1eimaLpEGGbkfOUq
J10o48gK1Q1pvPu1w0BNC3Sxrnd2BRMScvkSz38nU68lsM3LIzhg6F6aayLfvsF/7ziIUTUpUKpM
hsRU8s9BX2RWRwhGnkxBxp3n4UyW46vNJH67YWtyjkfl23EfoLIhVKh8sR5cNKQXbwdyp4RcaKwI
2iZA58lTDMOJAX0Uu8Nh61GSDCS1LYkpSzlSKPnx/DmgEwbyz9sFPmCplxSV/f0rlfWoMTTEnDGb
jOSFhG08z9NKuaE68FLw2j7eB3vd0OQJh706spL9VgB5sV2/BX8alWugoCpw9vFMuwPq9MyQkc1p
w/n0kVtYwhXC7B+QtK+n2VsHuTPDD7HktDyqsK0jSXKpbC7SYj4hae2QuljTUHtxkVSCQm6fPmpo
AE61Zovv5Kz+S+1VZ/ViQMTG+FCLhnGbOTnjsUfeiHe1/uF+i6KEjoZ/Yik4pFVvXEh6tQnsQ0Eo
PuKytCRzPT6TB/ZRkgvPV6mBcqiv9XSrt7g72n/8jWbwTXHmeb2CiOpPZaL5mKBjzsJ4ffvEWDvy
TdlGnvBZM9/o4HLGrb7qHDvVWUFmUmw3N0chkru2DJ60KRsSOFa86wBeZ3y4jZa2oLkW3vnPoEY+
WSWuge2taZYYzswM5P0Uxbn9UyQlT5hMfjPlE5V7tX+ntJVQDbHgn3PUk8fQFrCfMjERkr+Ms1jm
CfVEzeqQdRHKaYcgmXQ1qeZ1TiY0wm+KMSsTR3cVqt2RDExETWMHZqqxI6QcHsGbyjO780YAqlrd
gzcV2JVx8ZCJ3R1nnJYXx0mW9lTZr/Uk9v+KJcv+JA1YPZV+w+IiDdhqgXyu4xMv3+QxrYCeQ+1G
juYBuTh1FdIDwZd2EiigfEx0n5+2wVc6uMsj8MGc0BAIay2bqFbUDh+gjPortOC413/leEipvlFX
QgRrHx8dEisSqrR+ZVIgpPOd06lhGEOaewNfDa+tVoDh9eK7s2NkVMEysQyYFc9YAXaTnxTDnQvE
hdQG66xUKP9pAA6ZdnaOwPKYG0Y/HDFvJoVpGZYVDmntBQNFszQEp3Tp9WVHpS/gl8wxM4aRC5LU
SxRaHPJwa/Vss/sV4n/pVdPDL1p11qr9IYEdZUHi+NiyZlUrzOSjzqhKvNB+wnnejlbFgB8XdtrK
BJmGb1hbx0EKXPJCAOi2jj1kDkfttrxHrOLAqwGewnkBEWlHLmtD3ijx0K/8s5bk9Bo+dXu6ysLj
roZIsfIlxzbaKsBVv4+J+1c93dE14u2sTAs3eVZ+ot8f4FfPPOeU2rTY8lvulc+qgSeQ87e2yVtr
nPJfpUHsgWYcF7WWGBYyYj6TyTjk7tPMsWpJipjinoK0JsdiyySEqFF3w2HYhXsxiIV/xqN3FNmK
NdSB3YV5jZcrvqAmbJAFX4nBQMtiE5GYhJdy44NaBbLZ4sAdu3rNJHreojZuSnxbDPf21+pOcyyI
m7+J08dXBFz0g0YZagwAOIpgciLmN3QUv1z01xDs8pV6WpUfW7iJ34inZ8fK3EBxWSI3NnVhQlLM
qxVvDPArSRhYfsb5HGJZXYcTBoyDnWCAJD9KuVbGnr/tyAuRNRCZBy/m1OtxHGJfipRHFNOE4LKJ
MtGswUxYYmF6uu9b88Op1Q0mZ5YILS7qCcukw6+9PxI5EQ0ReXnDvyrN0l0zfmRK9dvZnx8mk3Ri
TcIKvbKkBUulWiZQvfl661cPyHB6CJkjLEwP4ltAngc0saeVSEHz0e2eZlFKL3WeBAehH0naZpVS
K7jTiCfce7dNfo1ApJWySJZyMsuBf0+abOF05qIzp+MO1XcJzbwbbrfa8/BKvVrbr795x1/p1ZLB
EqdcAl943OxFRCWi++JiPlK/iJ3kMjUoh2Y3247PwrP0/Z+OmQ2PkwzsD86C66gOl4PQWqjVt7wr
1NhDbhB+x2T3o3/9JsISs/a35qojCxvLEimeGdFIMjFRQcaXyWh21ETpmxlCTPlCbj5jTrr8P4rQ
zIDt9csvgPsL3EnScAJLbgflw30Yfcl2K0Q/KWl5XOVgJ0Mt8Ndi7itF0brCkIm5DNGqI7BT8OM1
0+jbhJSIwKn2bP90E6Wyc9UqdGx6azxckilw1WITL/wiBPnFyQ9NI/qyqf/RDLmxU0BOs76NMou0
MBcf/S6o9nClhCS2hbF2qANmW2XVl7d1IRASe0ohtfkXb9KBSTLHdLf2H3HraI+/nMIvf7q0acIs
OittUDemNcTU/FxMiPw64nKhJX0FwxZCHlDF+4TBmwP7ZI95rqXOERdmcThwbBnYSu08fE1gEEwE
dDMmNf7lg5qcL7ieq+TeriQzdcaW8dNvBGeUqv5CrUZ2+AOIOVyZR/iY60YTdY4Cwx+H+sa9lwBx
/VlG3b7xdD1BJn0/0F+KgX3v0TEcpRAQuOEQwSkMKF99vAIX2SSqPYM/S4HMrCwElTbdpzMsBtAb
MdI0MYNK7RjhPKUXkB/h0EwMgAY1fGU0ytcKVIe0UbaRi5pkN2oNHC0Oh7mL+LilJFX9pGpzwRk4
l7F8alYkXcQImjuCWqKAfIuC7IKflh8d+tGg4P9TpSMyu6IB9iVbx+VUBnl3O8Sn7RUNUD7+SSqX
2IYT97QjqRmjvIF06lVoWCuqG9iUnFrICHUektWU6xe427RmqdfVccMiwkw0wAg1KjSWRNQsMVkH
tGQGs+GvEOFlysy2mNvt1zOjwYSeS5Q+cCzaQDtvZdvvgheQkfBUEmQvyzDagnLS/71hZo0vjM6F
b9Lgr7gBoI7bBqCS65o1ad2rE9LHqPHS4N3+AlDGPUX0YsfhtZy/pa+dUTnES/2PR1S1unzIN2zI
thqbWdQxuaBZFDYf8MfOWqJbPJT0G72tZ+v8walD17QF7pDX5iUvpdPdDo+tXnK5Fwbvh+eq+eFn
zWcj0O5K5DjEQE+z7TKwUjaeYgr4EvVmQJmRZ3aL45wrx3b/6G1VbeHyw6tN8hpuZTo84hSXk0RD
YR59F5/3impOKQT077W+BUrC1HpqoyOaW7lNTjeBpDT9oVeSG+J52828vpQpi4ICuFzR4RQV6iGZ
hV9p7JFSJju5ajfTm/EdScnG2/ulqJHQbwEEjgS4+OaXJ0OMLiaKafUrelZjwnicYp/uLuLLC2gf
iK0GSWh4INk0tz7Q8JQVOR9QFl6iH0FrRD+5o2WCI5aCa6rcyNlAdoHghnalQ8ghLDg2lp59tpak
3f2NEUF4VpHPrj4AnY6IexWhIbOCPbO9znUIMF9IkY2RhdD9dKlzoM8mZCjxZnlC1JtekmFrLZ7t
XXXlTIy0dQyP5rLTkF4WL2I5Vj2mJWZWVHUWuLbNVGoUdKcE8lynx6prEpjvAam9+STtTV7gMx/H
/KBRctf7vx0WInT8PdhPq55XqFgeo3Ewy+c3dEyd46af2DHcmRchkNqxTDtzK+2j71E3nJ7Oy198
tNInCiWJuDzwZo/MKdpghaFK2wnocxw3v6NcfO4MfnK39eVwgzFNtqXA5XMkmoq4buW80DbdpdNH
kK75uCG4UTB4nMnp7omaTDK5fxVU4Qv01QwdNrDL+Q5gFQARhutSDVD1rHEZzdfeakcrlQTY5R2l
NC8x83x+JpxED+4OQrriQRO/VHLiXvBS3vmnB1bbXvgIAaNZN9Ty9W7NaUJsFewNO7/iI7jAKeI3
cY1vPuLAZiqvzckdJgDxiYkk89Q5L3yMlZPoZr82RGDnGC8dhwaSdNqrn7yONkL9HxWiFffYXLl/
8eYvIQakiGmeJUD/5OV3UTuLHtYoM777glqPUztpK15L/7FGExx+cw9d6nN3K0RwI1QHzPB9VnVm
HI98K5f6Kw5UvmibolqxHTVgM0kA89JgLeoKU8sIVEKX6YLFUu9zuU1L8tyOzkeIkbatdE2uIlNn
O1EI16uBOmDejC4Wmmf5DixeImWh+rVzqArS/XoPFHa4HuuWBlckBQbvqNYLDCFmvcg8fDKJGePL
+jVenk4zntaPmotXT29WZBTxW2PF7r+eotfcGxj36tVUIwTxIygT744HSUlbRw161t/uP94TV45e
bFCrFzwKpg7QQI1UxATaivE6QKPC3f5HUq+p0/ZN95aPttIwSUnuTXn8mip0PUgfGkK8afG7hO+x
eRGSlYGyJXEvJJLtu8gwo9WqaQkjR6som2Ndgj7CXFhHJuJB9892LjqrvW99+8TI9oFKxbJD7kND
DmzPLPJCYfhYWpEkpjD3e2do13pgGaivWQv8qV7+Cd91be6G33B/xBDm8y1TyHQW5Wi1wU21EwbO
Xmha0lqhQX1LhDXF5FKf929iWQ+wIJgIygbaQ0b3j0/XCihoAIbYAXfwOvaEfPhsg4h6BUFptm8e
N8EqrMrH/NiuA3FxEM4lzPAa0+ptsLdp+ELTXRwmh8tvabxPa3BJEvkKnqYXKrBQHh4zkQrnmwVn
5QSEat92it9CaTPNozrz5qgJ+tCnac+iMMjlXF+8pZe5DOJL21FzHU7tpoNzWp0gZ4yq00v3rVEu
quL+Q1juGGaAqTdk9XsUe+ZW5po+Ef9wh3YpWk07cycstYJBvv3yZeQQkKB7T9WnqCFpE9kYw4uJ
IHgLbDC0HMklGdPylEPLc9997Om1iV1dgdPoRwQQg8zAw3IPR+ZqsOnsa56kes8b4WzRA1WXkzFr
VFf6JdyR5O5EF0S9UNhsOL6PqCe2f3FNXpSSDGsLJO/qbBPGxJor6+vCP0N5Q6izeUrUerpwGfUm
xQleHrLHmJMpzFRBb3pk+MNsOF+NTw47b76uZDIkxWbD75+E0MNeahpDbUdYqz48zyOsAbu7bXqJ
BIyP+T/rI9za/l2AEB4SoIW1VNAG0QeY/TfQLM/GJtGSESLTEg5ygUMTJjWwjEsg87Iasn/Z0JRk
OOxWbTkOoaHn7CulL+P3ln0j28MYUQ6fh45IgJ+Tj082ANsygVHN7cjBCmhWawMzKv+9w+XDg4rd
PaV14GTkO6g4uj4lHpsYxq0NudZJzvTEobF+P3iKuOA+nxNeGWk8b2gXlJ0VqspI21/GVKN0g/tt
Grj5Ub4D3sSnWiibyLA9jgUl4DPkQQjs4Xho+Ka8Og7oti7g5WxcJJXzIILU0UbY3ZcOaCEXZqaJ
7LuEcMMYyNI9t3dSs8lpV2T57STwH7d5xZG6A/JuO5FcpqMiTHMswtgQOcapR6y1M9tDi3abppyJ
fZlb9Gskao2DjI616iN7bX+pqtOvaPtxgU+XnFFmX7PBTsUOKbn+nCgTQXQtkKRlxya9La+G3JbB
8GIpllfnuWrWKD1QGqC/6gfMmdmsJeOLIti9HSP5HVlr76tftc2tnvQtsh2gEu1PJeU79joaYq5A
jstr68P1Ob6DmouCcPCkbOqxvF6W73kNWu7dmWLNGF2v0smJxvzX83HL1o+7CxVsktvdcCdfScqw
7tPrWJoj1gImClL6SOLb/zERYUNAVKiabQufhQHsYcRGNbpvaT/nDSmSkfXVtntxgBioIaCCVsiO
ofKuYuOIVV4fVa2vKgOzWPH2kz0+FRuxUeDVc1xqGQGRgFfPcltgMiIWWsZvwp/DFOXjbw4oOalF
lWT6GsJr4fdQ/KNFkYYH1N9dIjzW0oCU0e/VMo8M0sIJ/kD0NiZxnZxF0tIIAy6cYs4jk0ccaO2V
Th5ladUgkR3Dbb011xdycf9Ru8lRVtkMUn32Sr8Ldpp0nlBXAmM1uQLAGmnu31YQBD1oZ+Vzkj3K
PKN9irXVP2pUatbVQD/sOZQho1KCjA22VLYYF2zBGEep7zqznQyv9qMxISkHVEEFOyxmN+zAVWdw
gy8qDBQSRQKCfDQQduyaTDgdvZY2vXxKt+vgXrWIKUpNufMh6Kti/OWwhQbQdbDfXNTIet3/7uSR
2Vp7diHrr9/q/4U9NRs8szl8MrQky54llmnWsGPXLoZQ6TbYuRO3GYbj5Mc/0AGKeq2dVQZLP76m
zqJ1NyzafrVbTw6bJdyplewb6UnXsvCzYCKvO85iizwbkThNibhLM687aMgpGgLtTDo4YyPDVg8W
OfqPdejoOg0QwkWRzRQVYOUIchs7Z0ivR24ugGjSqxHH4B0akEv6RxWXgwA8dch+3tTxlG5c0Ur6
u+6Ubd2djcGV1CWLBTYKscVEhV/mVnHD8GWGBNVvTGI/mJuPBjUdxPIl23FH+ypv4OgCj6u+RTIt
HqbF8Ed6GEQcJHLNqaTJ0uKpzVmLSz1oRmmA6aCuf+OuaZWKpXouu2ANQc7adGfKr0qdas/h+Bum
4jcofb6zr60Z17I+rmWYYjoLffSx9NDF7u94rW7PiqQyvWEeNaCv+Fai1Z3HfNZoU81ls5MD/88P
CgGu34oY722OHz+/jeOr9Xu8AxCR4jY95BKkOBGL0zITa7pEgEJleVC8oVg8IlA04L/Pvs86FlQW
M0rABgzL7Lmb7hhesrV3CU2pOzvbPJ/WqKeWOUGmLZhpKN3BW0MeKoh/HM/8P2oL4WlHtpCq9EP5
AWvbgk3NhOVgOdu702VkcSgmGw90XfG4blvALvYFPvfvPohWhmqjPW7kUeFUv0t79UlbQO9KWQsM
k2MXPZItj59ftV2235UGXkaTMhfCjHIB+5EIGj29B5s7hY40CJsN2zHqsFJGpgscQK4SCpKTGfIu
HO+jLvjjuUw0jDRtH84JgSZK3VTgwFAkK9SUC3s6YEXTwFIKHeTifeHCCPfcBNl641qWquXzfYLc
C/1a0QEbsTjz9+QfoS7I0tH31XEvSi7gm3qH+xzVQFFWuMl//rj4mS+ksNzjMX7jGJKUm9OfB3R+
/hncCawWCqywJpUw0KsocwKgpxezVzC397V5w+pDQ0Sct1zeBknuvPCC88tFYoCZwxSIiMWR2W5q
yl1603aznDDnlcVFx42P/S/CoMuZ8AKq9Q2jYFM07AA7WKvCEp4imHxRKK8hxg7G/qci7YYOpVh/
OoVSc6ldStzC5RlsWqNtI4xHxHEUSrTifMLHoLhixxVeHuzIlvUs1qZ0r1tgggeDZnd57mty4HZ6
0vawU+hbxPWglqmbbKcQpatbawKOR6xTP8ibGk5jSjzoDEhEGl6AEnekwcV5M1CB42G5M6PPUnq7
mBjuwju2aba5Ve+jMsSbSfMr3xlsmg2SUtTCXKjl/QPl+05zvHWul44SX88YmaZF6n+l3QjVa6tn
LVCGiLT/GEfQFCce/n6bwyHJwOhXTZIqWPVWSDGal9BZHmCoQKkC0ivP38jbRoEEVto8Km3vArL7
0kppW+5C/sBmaZ4OPfK6Npo6bPBEbKgmYr/atnZVnVtSzMUPIToQH+PHQ6vTRZFkGzxA2tAJA/t9
jGuQrP8//edNbHPjD2bPXoYluEi/lWHdwC4rKUkQITXguXSD7vwDwcbrdjYf7TRzlU8Ir34VY9Dd
YJYWfiTvXBX0QU0reo/AIgBPZ9CiK8SiiMVlw/NzQUCKA6uTr3EqWKrys4+MKGGB8TvKaC5sQsRW
fJMjk+JJzlkmTAVS9Tlx80vYZzq0FrQRLBRVe3MxBFvdUDlDxfU/kRjL3XppnV4vO7DmTSN4Nf3m
USEqPkSezruGtrE833T3fzO0i4x/cZC2sa3MBqFvDZcfUHHlvR0J8cZirzwP81sdKGexhd7koHcB
v/OrPCUgi0eynSCJj6XnkULmUxNE4bPAW5N2YjH9qt/oXe51BN4Ik1PqunDXUhStzVZZ3sl8Lhk5
Ng3Cd+eVmZa+7L+hIuFP+ot5ijCUjn9r4QDbwg92q3Ok1Jv1jTW3nqdACiP4CpnBBQh3TX6s1+7Z
p3kMWoaEVULR5ekJ82Qmf2lVq/V2SsHSpUUVfr7wdMMxo5V+3ad0Cha/kt1CEuG/1+fWGQ5cSX8K
KEkADmGApxtxiAIud1hncdXHKbC2kAnAjlBqL6h44A/hA1II2Sh0wi1zapnMX4MaYxnbRx3vmyHv
6VgLLOhcLRapPQ6NfSh/kI24esrJGklnbpBhKau+woHG0x5lT1jezeE81GUC401ttnzGrd+/j+/v
7lzaLMWHLNyQRRJf4CVdCY9McMVX4vn2k3/EfhjPrJ50nUn9kA8Rf+MvBDFe7jiPnH3BuxGvdlyz
1OYNPu/CSEqz8Sj041KfoZzVO3/7F3Ij/eal9W2M5kJHmqhdDRgmpqv11DlHCPiTpdFTK+CWSNr1
S1CEtiz3sJdKdUojSghiKn6Njj0xTqV1g5fZJpUCPu9En6z3cqMGmVA1/maOnTHnzfoFJ84OOAyg
SSrKndFvrSFvsHohSqUh4GiyPUnHkxkncxfxPTkjSKB3e4UGnC4rq9FPYLmGeWUFh7Ucq+hafdpS
+DcfnA0xbMpTdG33BIsYg7GWGlGYWq+BZWasj4sE9HlDgUmG6X8Lk+CqKlaAbsrO2WBbQszvSfhD
dPPq7QsMDpoQ7rQpp+/rzLZDmNb/Avvnmos4ulU/4nPcOjaaCYQNUsaTJ4P1D+nHZ/sysuyDG+sF
DUF07zYMNP6P6srALsrZ4VJRkSWPHldjuF0eM7NVtSmAiNmeyY6JrG9oIFWPp8yYvaYvsaZUXDT6
s+8XYBzs1HcGUio+tkUpWdMbEVWBqx6/okOnmMh0ErpjTK38hol1kPnQyWV4hytPEkTCLACM8hOg
AiQaBfyzOQxzNxBwF5L0ZP3UvouJJRT9KHn5qdwD2yKi9QMlaIo/C+a8VDgiZSkujEOWJNWHC+89
gt0/EvQ1IPvYzWBGrk5uueQygWvVxA1Dsxggyh4IjnRLNLCJgCdcw0lPdH9pfqXc1x+7Ia2Uez9P
1MZJ2cFdS9+l2ZeN0uuoJCEUYM1nD1+NxvjzelO21bIxlZ9NpzHFfQx7fvnu5KO+JaMK7APfztyY
wUhHUCURQUpWr+tJVqEjiwKC2BWuxb+8iDjcQgc+oJFuguB5xtJBp+ULBB5c75wfrIEYiTY2AruH
/EPTWyTZeklKo1t3c8MvB8LO3lDQoDVbUwC9V8+890r4ZNUKzMiv0TfoR9OtSeocqwvTPpToTmIV
YDrQ0CuRht8bdYFRFo+c+7l1nRyLHEwHxvRSc5ZGInnyCOlAqL3U9zUJWFaE2N4CNiiW0oL85n1k
2WtdfP5VultNcio2DKtjdsYRChc6XE0PcDN3p2MKMCKolTe50fPrnFDZibvic3T0l7p5xRFsA8b/
Rtd5rbkewlMoLb7X1kwbeoYMldlb3/9fAkIrFpQezEmjwvLaOu/utuJeJJtthVjWhn294+OkIqJq
LZ2oOqIDHtrogHJoDXaGNQrUKjUufHUpTMBUulEk89VIKgdNk0Emp+DtoktoB2MTzvoV8KPQtk+F
Jb3dwthmI6i4bFqVUYssq4DuCni79Ibn8datIcbmPctT/c3CuIambqfAJSFt1ZWfPYkZdMr/rYEy
17c1qzCP18a4Qnsv0+UJwFpBcIQUxqHLFWg5tx3cSv3l6GBoa+suLa7xeoabrWVNSLBpnseB8xjl
Ys4UZW+BPBWH5w7nUe/1XTyhQ2YWvrrlGuFokU9UYhNUZ5zIEMbqFOdDnp9iGuQO9onWDzuji3Yb
kFY6Sn4EZBYliVXRfwsVPBUX/EG5Vrx3HtW+H0rT+RXCFmZpaAit8GrmDBfaocWkkgeOtowNVLm/
JPrhAr1n84KIx6p/Clu3zUx11LvUCVnE+XiTez69JZ4jdhqTMZNSUlgnEQll0Sj2IWhOdmi2g1na
AQ2XF+n6jxR+xpqwM7mRyXwV2v7AzMW6vNAcj8HZeCReTnS3MjM1EubwgZfVkpsHn/S7kRTd2Yo/
E04QcMNMNMg6KTCQhFgQTbPehQfLhCt9U4qRfa9A4viON5XTZg/vzaXHQtYK0+tbBGVFgNeK5UNP
lusrQmN5DNIbxfSFbpufCt62sVPNBq7CBJEPleF32ZgH3AN2YHrBooaxslc5Raoo7i8F0XHWZlPC
FikZ25mVa+j7gQh0Rb+8ZlJWpHrHJj/BOJRuyU0kA3sXHEnF5wurfBHnyG2BzvhuQr9PiSkBEi3P
yFE49gnM2ev8YxO9RfCeD4FBXluztK0O9WnXZp4WlTskuBG7PG/5Dye4oDRK3E5zHR5r741XN41t
h6dQTDDpg+75kMdl1Z7pYIqc6aq8H16/BIpdT8JvKByva+RWxTKAtPxOpZ8d0fGWNOM/WsvfahxI
asQ3v621Yhm0bNt9a4cj0jAAdthVW/IqhyitnAb8mrxTvFMsFlPW7B7YqSUtnOXQpW7P+jQsRPs5
PXO6mTYuflep3R/jr3kxp8/yWMXFWDtHFTvD/+IK6YWW/RKp34MMkQYOMXPcLg4ouDA8ALS/yom4
8nkL3mTq5Tfobb0JO+zY0NQdmygtbe/rouDu6JT5GhqnZU/Hl8z8sQbR9liRlI6bzFs4H9pdMmFF
mztZUnYZbXBAr/Yf6PfbHwMFFG6P2C3LWlnx42AxAGx4z7HGivE1TxRbPMkyPDkjoEUCzyS9BJS+
pMzm9TzoWSAnINlPjwusMsMG1Ar4UkHW2wOd8sz8dTnVhzI1w4ZiZM3UCiQGVnr1TTBYe/838bq7
kDA4W4YfC0pOQKt7ef2Mj1FQxpoQ2qMORwqRM/sZO2LBnHdlX7zG0aRMgFFCzgLwzUKfA/s+c9Om
2YSWMDxc/SdSxNs+K3cPwedsjRXG4gMkSD1Ekr9lrqedscopX0QcOrpe/OUCy4DP+KcvxEv8wnv8
OLmkCA27vAZ865vSTa7WkG4BUk4tkmSmvkBKk+A4pCZGT5uV+r0GNa1RiKqEcW6rCBTdreEYs4nC
OmU3/safLcLSZuieHBsqvywikfgij7D54C6qhYMulr8LEvGTQ54YTpW7okOm4XKa5t7qJdN0myYE
Svl7DC3T4kAEqHOThrcJEi0/AW4YDeg5Y70IUubGZG90jmu9fOZhDpnZWdQX3fR0h78oq8uI3lPx
qRtjKcdfIJ+3UOJacSMFtz88o10iasFVG5xA3KHFvrsl8a/+ikRHlL7gkKtCPrUxzv0LYHexdlok
nKOaWjM+NBVA2IZ58EJiZrhtJ5lXc5RRWN9BIozpe+5GYQBQD3GcSvHnjO427NDh9jC9UX54xnUJ
9D4cEDzMP/uDwF9RB1huFgq9QRDEYU+D9vaaD3BB4jDIjy7vY0ucetMudBkpdmHpseWxnJCYr1eG
pZve/FR2pfOfWvbpmPYGoaJKxWSBQTPfQVcZaPHFyTh/LHufpPI1uVE2rbra/sHv04/5QVu3GG2d
lSUykxr9ZPNrbvhqFndQ6cA5XmS2eqI/M0bB6l6ojpqoE+uPsUpstAAweSxdZNGtQMZARgBrwf5L
7QqHpJE3IH036x5OdMKbshHI7Ha47jZI0dEONa0aXbC7fxmLtETAc3d9IT0MfzUj61lbEGSyZTi0
9/N6FbYdo+XYdh8bBalzmXoPgg4T62X05R29Bu+B7tWxie+w/WTJybhLTqFs++2Xl6SOA+S4+XGw
Oh/41XkC6CgSAh774cP6QoTByWZ1kcR99rGJiG8RVt5caMX8ilNW0LIMH5WecpBrIuOMtONoYwBe
pUZv4IOvhdsgKwFrK4R4OZ8QgtHs/CTkns1cW633/7jtwhHeZTZQjzvYrVjntNg2cQHEMTk3ZgqN
k6M/bQdYivCLMsRkoDjsS284FoFs6yuZE8IyK2iap9BQAnb1ZPkk9kVVZHrvobnQUhzq0PgD4cPa
0eS4q25BCj8JpWFvcSEesGN4fnDtXE5JGQBfD/hEvh7Faj/yxSMfgJm0CaNB1U0TVtz6MOVKjH83
J9XYDtb+TILn4lcGro4IHJ46kTpgeGv86SMTRGXAspzD8/ls5lbuXVbL83Ezg0cDLt6wKxjcyILq
oSGhSx4DEf7k5/22KOTlp7x6+3KHiVpVIuU+QW2BZbxqZ/xK2H7Vx93kBLBJKkbXj3SysKqN3HQT
nuIcCyFevteg7GRyB+SWNtvZzVj95G9YjQkSdIZyRlQ9yubaxuvzZKUfFW8EAuNolLVIZ/0OJnUn
UWqvkmsS7ctc+lxNmEOMUROOmzvnB4YxNJX1gHeBXafy6QBjCXlc/w0n8XMnRnoqyC+mR6oUVv5x
YwmsuSYwbljcRRk8C4UAncGxElCgmwuLr78q8nCeF09ZsEyiBmEmBy/HB3HleyYrxc3yyP576yB9
elk4P1+5xKoeXcGh5FCyAaGx+km110LmYxN3kVcn3oQpYFGBYtumf6XsUK47JT9ieheQc1Y7s2vk
cvHrz7wDZTUzNSB8LLbpLsCP3Vo4ZD2bOUJb5+RxxLK1VgFnO0cUCHu8Ml6ydK0D8DUec/pFCHAS
9uEUdIRXwA8JyCBmQToy5O8h0btIgl3b1UgnukeUe4LS+roaI4PlFYZJuJGlyG39bDwv99y7psHe
6GmCX9sS3Rp6C1DGXdWdul3WKM+dlras/5gv0z9iF7UGmDKUkz8voIKHlHIQGJeCiIzwEkf0Tbvm
ApVY6klgWDHBSInFi4Voaw66gU6FCzkq5ay1+jHPOHgV08ND8fCJ9tPihvLpmtsDSE4tmqrZDz5d
dFjOI34lZSlyo1m+oDSyCpcNRnNro6H54J6p7opq/FXzu+uoVNK8aw6eFbHFNjEHdKhIiORaCg5F
Q0FdgJ2f1/nRydowouQz0yAn/iswkUfvVFDuzZkwsDTFZ/mWBTAKmThqQ3y6vlmo0DI9PYlGtbQO
ULsbbeJvrfseugEBDwgB1rXl1m7u3ErYASICCazLORKWO1NfVt8fZJPXZ5t5h4fnDYruwwQhOG+Y
oqvwP+Fq4ylUAGZ1XkScs7zWlU+AF6LvgDxGc1HGkag+MyNGfTNqc9Hpt96p1Jo+ATccOuUIqj+s
PyG6JS0ZMJq8B3HMGyGmYqeZBgcphX+Vk3XI0wWywqQtBFtnoGiyze72ovn7pPFPErc9ned5iVTM
zx1SKsnvMrY+P9FLf2ZIpmwDPiQovln5adzmNUdaSdm/RiTyUeZx47RnLqSxiyLLkV2pBj5xCQL/
5aR4gH+GmlzjI5X6WrUMe2Su+M0leA/CI4AqaeL77Vs9Q7PGmOaN4eTVU2J/oy2rru3/Eg+ujZSw
PNbVY97NwFS+psLcNrCN2+PJJJgbiyUFKm5jjv/PmUBTlh31s1elQvxNDVeT3uvXSsndOxDFEbmX
xDRiLPIMKJB6ybwPMDXYbb9YNX/BrxIIdq9sWntWTpgVw2KS6n+nDC7p9HZav0dP3xt5wog5G46U
ywhp5W4GkfhNlAmxVPZKHwgRUzvhzmiue3IzV0jWABoitY8H5NMtRg30SJ8J4SLsTr3MilCflldE
vyC0NiotdK7I2I/f16UQo/1F7iZjwzIH0WF7uQA0jN1MIUdmMc624Dpej32jB59H2o2p8iX7N/wi
Vu0SCTncMyUcHRi1lLcVgIZqt34Nqy984YaaNvfQzIz/zd2Dvs7c16wbmpXL/Lcc50C/S10miZR1
ivM9fbO6g4iXz9iiP4+NfE947kO/lQbYXpJhUI3B9/cVrq/2KsVpL9kHQhMkjVsRG1Kn9EKrDvr6
Z2HH3BGelxRp1/o9wIHZdAPFMU4QhcvozFtFCSFTJDDunemAtTgTHsAc4NSfMNylEHEs+SlACOmQ
elrPxTD7RDO1Fnwg5Vtf2qiHA3WnhiO43gTbypnwALVT9CJNWkx3qR2ldS8j+ewcUMzyqoPVqFSa
c0khlbmX/pAlxyZuakmB8yr6OrXqUT66jhm88Y49YuIJGZZU4vGHNVU3jrY1Y+7wF2dvXwLU4s61
CySNkEbMaI743GnSRF4SCJRrN2LQb1PU+VeNAm2bD0Q0JKy6zqMoJajKE+UPKPExv7FhU4gBp3xn
brCmgn42JBHYgnGbcIMdPsJbczXWMQMyiBnV5Y/93L5eAMpcuaDb+XI+R2mDPgzgWC/grzvGnsP/
1ZPzoQGtWZyx7QJsINNp5gUSlCG4MPOIgsmZIH5Ok7EHXw1+4naZH7/3o0TGEk18rMgHKYjCki4J
LZzEOLeB9t3P3dXvpqISc+N0U+gOTXGR2f38DcglDxPZZ9DtwOuyHszyhEotTH+6c+F3DAFpryGN
oNBSlzSQYDxBPqnKmUoRl0oV9RNIKq0bLwtYIjaOLV8M83tgjxh7n12v0PJt9T84QaCYwnR3hp5W
ON1+3+yKCc0/o/KQZDSgW2dAXc6Xq2NhWutAtG8rXI9XqlzqZvBjFbCd7bAGdHIs8KbWxzgyj1no
j7NPtovoKrUWqfuypIZARjDqb38WLGMa7a62W/YJBAwagql5cCFyXTp2DnsaRQjr/Cjpug3zYM3u
TR0N4sTETfmeJSEJodvopSFS3jK8z55CxOVNKBQHDAxxeX1+lemn5Otj50uEnEJgXDQsNFkouq6v
8LEGUTJbm1/gUYQ3z8M9IwGgrVfEUrxsArURp4TprE+eGPHi7KfUf1FUAaGCtCxDS5gO8UKRWwsP
/pRyk8VGX88EdYdIWgSEPfkMDXo09n5CvR/FvghnAEaQwTyJx1zmvtX9A2BD8F5xpxQCr5KQEFcE
DzBZTCi2H2esL+kdMAX60QGP5yFoEwccrGSwsP6KimbezhRZ511qGP/fkQCfpZIixElm12x+J99D
ld42A8N0LcyWYOztXJBxD8qOAb1kAzn3hH73KIDMFgJA+H5uK4WzwEJKYZdUxDZ1tkm6Xqa4/ObS
CUldvABNkTqw2hE3E8FyjylymnMkr60HqLOrh71PPiI4DDxPnQ/O/bTcVk+figiLy+E+oCAb6u4X
NsyU0mY1u9cQTrX4ncFCOe4D/ixPou1BfQPCBBydBXGly3f/qLedZ7YchrTMV1gjAbZqzReSUf8Y
d0l5beKjJCuRMAOSABn5eAQ0K+9lQn8vUOrrcVY/QbWVJTeqbuKJgfXF952mCWX6i/E0diRjEcN+
kd2T4Zjuaw20kBV5v0pl4lFEv5IPSRCbR/hI09XjGirb6Cv5t0gkxDu58ycKitnn1lPJr/aQztjX
AAnNBzT2gyYTTtWRFuzd3XrGNUFa3ZSVNbf9H92UaDvjMa4xvHfJydrPD+uVT6/hGFpL4gXRQ0XE
EIVaNraXzeEilChv6xJIvZEq8KROC4rLoGFMHyA0VGNxbu38ZixeGs4o620KncwcSmiCHp69gmfC
/QVUckXwUdR2dH1c1LgmmX/iHWhWmWe4O3SCbuiE7WffjfEE2rl92HD/cKMRPyF09SE/q+nH1O94
+DdYLF1uiR6GTE6iW4/PxqR02b/uFpjhQ1AIck6F6BQIiRR2RmZyW0SYJmZmrsKfbLVIH8LvkdFr
xmz04U2XM8U1nMee6Qos0mTa/tZZaB3uTNfHNfVLYJRbFKZ/qoXROk069pIRHyTc2anCu6VdApXE
L+iDnUrSO5GEE24T4g1mOaYLeuYrEs00CngB4czJ15oXjxhXJpyXdn7bhpbTjS+1j8Ear/u0czvz
qzSEuL4uKmGzE0T5032VO0jFQVxwWomB1XYDnE+3AistQshhnvxOLrcHKjRckLNCvTM0J6eCia+0
nKn57IZfY2DacjSV3ylMBNCULt9hgYxAyMqbziKjf+dyUq6IRcfvDjSUUOzLQwiKk3dA4P2Hgcxt
YQhDWY1mEYozLL/hTWakqSRc6/H2FNh3957dlodVFsWkG7HzpTfkiXJEJcVG9G4z1qIOMs6/eVN2
syv0kZoyAgCIK7aWsC9NWEEGroDtgk8LFgD7J08procWCXbNAY/psCzIikfxrgPRvVjWAFTfdNHp
OTIK2rOB/0P0M0mEYme/hmnoNoim94lCfMMPLAHicCpMa7xhA6ACceAvXHUjWXWl5QJF99GiBCqF
lVHQbwmzREr+5b8U4DRGdqD+swJSSE4ze2wHXLwDy3hW6GOVwQJqStwTUuQBX3kPuTVQk4FCIUxA
ij5DQsCkBTC6I4ST5lnbMab0566SsjYoaXYrV5lTUkXo5ZatRmEUoiX7FysQ9p/nXUqSWySiHOp2
1Ix8KmvSz7eSkiA7rmslkLBdanDyzksLKZRHYCPlc5Bd9IGNxrdOIkxQ/oZaZQyyZPggRGiZrPKe
JHCoyMgpB1Q1lI3ZyyK3BlgZivsvpPRLbgLfNV//AXkN17llh2RBvrkrDInl4wk3NmriW7zgCgoW
1yd4bzYqjHLZyrBCYXn5AVnctoqcPmp7C17SBPT0C9uAgzkDI28WZRAO+4P6ZtZ6Vv3m0IFg/QIp
XgheKAoVKcq4nC8OkKMfpOoYRKjC6cTy7pfN219B2MX/uPFVOt3zdla9WY92oMm6G3cVek3+NQ6C
m1fMvJ90zfUHQdexSfb+ZP7VQg+nS6cKWGTM0SDd0TuzKonYBHIcmmAe6Hhj7bz9yAHM8ZG28J8w
BUSFktAjOeA1O2eg4OuNdy+Of8THF3EEkv4+CsWxPi3AxvXPM4f5Jk9lgx/zdsjCOIRGWv6Hdkov
Nu1P+9+KWPBVaiTdt9e34pNUy1xXYXepYJ6hqzZLUD2tFNjGksJwGmhJfDM6uCegSPFU/x1TJIaA
iQA4t8QyPI/iCEe27a6+UAgYgFC6JzUfQfgqjugDxCQ1wowxQ7zud1DzICb8dBn6t3OUbB1lVey8
uZS1yzZIgluqFGjRRNLz4orYigyJJ2qaA+w6mvB6ZvtJHlZSG30xP3tOalJkUpEax0JiKU0gPlKD
EW+f/ALYjLnnYjsVQOc0b4zLce3SEcuc2kTw+eJn/qmauQwOBLJhm+qii8raQvxYOfRUORWBXHDc
nWsU7p0sEnFw8ckUfmwUocAKPI35ziDZ4PrhH4qNnHrZNQq0wpl7TrkCuXMyS9DBUZUmfWmFH3N8
cOvZck15bE6VSr71QmwkdUPRQmrDRtnDSzQFSXT7aw6vZny/Q1aEW8ALu7Jpn1yVa6Qd51IL+ICY
/9IKqO/IxgLUGjgswt84DVWh37fM6XU/1p9tNkcCECJF2g8VwaepsldUbDk4a1okOjAEeBpdAIG+
J927kxSklSFplV/jRnDVs+iTSSHCzZaDeq7/TBOa9y5jI+V8LFtmp5HYzD/2LSUcwgLreOr976ln
+5RYxf1P+1Q0p2kZ+js1PSJ73i8JKPjSB36ubmdfF9oHkHQOh4RMvHuCKbp6cQFxKOShNWUzhvG+
tF4ioFEDaXSsYKZBqirWIU1vRs9MtylEbWAPiT0iyfoYQ53e4eeaaFsLSGbzgrspdBU/aIMdGVaF
JMzAp7q8vQG2r79gNR5Dag1yL4Yl1mS9fvFcHHPQv21bv5lPnZYW7aM87xv3d2a4xFZT8a95S1wT
xQrv/UREtvA1o4CDnhSS3Nnmccin15bjJX1RTAT+pp4fSsn7YF7qFlwMyMlhHBsswxuIuQT8JzVp
CiCzaXdO3XMpaxJSTM7SkrIEfMawvoFpk0ZEZSZbI+FfVpeZPfcH08iVKoZAm1QMBytvuBLR/dcu
7rP/K7mspA1TXw89py6TvAKE4AHdUa5vPf5MufcEW1GUpmd6eJdi2/XLY5OIKNJGssWEiZUFhA89
sQLRPh0+KBli+nrX2YH/dFLIngsI4d0qgPh9feOdNMIOjqLdoP0IXYFMXv8Qm/q6LMJ5YimYnDk7
7XB5qT55YZ2k54jhvvC56jbMSRaneucFTn8qangYUF4RkVPiTQKpvtPuVBp4hk2DGnV3WTOIHVVo
ryKwy9s+TQ5AUOhFR1HULeWBSDLYrDTdoTUwGMdJj+Ly1jeOeodzGc05bLpw4IXEyeZgLtqKe5vn
FiEjJqt0UZqJWhcDjofiVKliaZfX9cidMxi0zDwSAKWoWg4Y/vxi++MFOzPdscl/kNeVbuOVceVd
C1f8QnqH1e8TPuvHxS9NsJyW3lznZzZf3MJjaVDOFjuMZLOdIFYqPn6jMC5t3bMvE9lxmBaPpe9E
pkUJcYT41VItxFPY1KZcooU0VfKoQKejix0g9lNnjQAKCaf3l56YTNKx3oVPj7lLETrP6SHSZC/K
sCRhdH61eub5CNAWzGW6jud/ILm01C22Rvh/lN/wOX4fDBOof+0cA8kDW6qRhfTJ0P/yDf4ZMZLc
B5oA4nz0vZbhAkElWseoP1vBMEwkQupW19jJT5rSQaHPvRp5Mw4qE1CKM+EWKs50dTqfvYqTmpL7
M9dEu1d0QHk/IF3uc9aDFK/CcH+cMsSVSh+85VT7ywUd4UCGVXy6ls1Y7sCfcJSgbapWV2VnDWwj
YaDjSK1CNMRvvF1dx1jGLpkpOiYvnUQY1Yg7TgXsiJH4NFVRNvzaeafueY9zDRtJ+T4tTcWuA2Kc
KDWD5bNf1Dbz5A2LwAFPl7SlkJZzSOi8+rJ/TH3Znx1iZfqaDRF+Dfw20T4FEAjTO9IeKRL/5cLa
aesty4MeckZACbwuweMGf9hmL5obPdKA26AalRF2tvaN9/lSyRf7T9QQRzuN+D737hkGEXI+scfd
iIR9yJhlQDOfpAS7NDvAXWAY9L80LcVl8i8iraDwfYrTGHD/+5HpepqZVzZgbSIC6vufscfAhBwy
tD/qZLzBNb6rzw6PtIXhyF9JCiAPe44qQz7E/A57M/xRiWSWuSmUjrAtgy4+Nb16/bQ1313ofY8x
N5vZLXU9nMgzhRw5Y2THn3nyFrclsnvkS6ZE8PZUzlcwqsyyXB1U0uqBtpivVagcmrMXde3s5ft4
+CzWmnJPWJiE+vUbLa5mzLqX1QbEt3/OCs2vZJkqEH8sCtouTC8vLA+pohbMMV8QkaahPr1lB2qk
kiX7VJjTktCJPSpvyJwtsiCKUncPm6tNgvsBmy9aGMYt8azuXuxpoJAG6PIqTrfyTWqPEHdkce7m
a3j3tSRw5XO0kMnE0Dn6oEhfMFor7jLRtcV/9u2Yi8OE+jcBWBuSQBdiyY50FDUrjfeYkyagVxMS
QeVkw4mGBJx2BrqKLo2+RDMV5LizuPHtuc1WGE9MBC/8boHYiY8iTvo7DtoVMvtzRc9QjOYY7RCH
A4pgyQrJQbyJUc5oBniJ8Eg4kqH84+88zcr5ICs+TSqjwDHhUV34vvSktTpZzkB56JaA+57hRuxE
KAjKfmVEFSf/D9ob0TKxXjqVxKFQhFL1IDtUySLp2izD3U8DvSzZurXkZ3zSeIS2xGJxIN8wNfye
TNNx4RW/WkLvNdfER5AgkMcYuyozhxicEWvScFek/sSfLJDQxT9F172edq2t7WU3F07sh/F5JQeV
e9fS0giY0vuzQhAmu6Q7lJ1ovBVdzKoWWozWCTndzb0wmanNyAmEm1QVhsAIgJNezMP9s9Jk7abv
lJNLmb7Z93On0THv6Y2LtQJxY3LKulHO6MeGecBoPUhidnHODkeB7KGTci7dKM7Bn/sqxTzBbphC
iv1H06VnoERQg3SSBhJWD+tDme4JrQfB1C0EQNxcgb11y1DLHF551ZzW7KT+ZOvH0CGSIxjE1FZO
Y4Mk3Aj3aW4lsJp+8kO2BDv9DuwGBJe1VrbeQS64SyTz0cnOXo56REcmSYUAHGUN1+icxYgcY0WZ
ON5RVbNHVz2fGl8r1K/NAwkqVinPaYY4Fm6F63VjYqFdVq068NZg5ZFA4mJEWUubk4eom6TJH7xx
4RLw/OpiRvMy3hpYI3q3T1e+LgC/GEStnGhRuhrdO98+p5QpaoEXRUM+M6BMCXhYt7BAzkwG4ayL
iNZ+Z6Ly1ZWQgsZCU0OSihgrr46SZtPWnGRKMAstldkZucl90ya4SP+CooZHwTHRTyKq6PGRhpIL
OjTmPPFxDCD1UI+chWM/QKTf3Y5FDPVJETOCIN3LwimQg1hfFmUS2zNulI5mplAlFEuLra6aDD+K
n/aM/dIAPcGBLnoWH+AF/GthrVvdocqnVvjH49Ic1eDoH1qqchYKbB3rkt/tsG3+afY/NqP30hp9
hJb3acHLXK9RuNmCWLvY9MRuodqaxXVUsZTetATfje6hcBziCRIgWCpmnor2gtykBEd9pXjY5ULf
milErFIMFNJ0fAbgZx/NSMoZpJJV6D5luKRGZ0X8V1bwLqkWRH0G3UxcnnZ3bDbfSE4iJRhRBjrS
i0s+FixLl+66xp93yD5O/zz208aSE7WPYaesdivLL6lZGjb79N1MYdiC/Cr9mohxYV1SsNoZTxHB
YdaH/n1eSR9NvPr9MFtHDOBSzG3zw8j8AMreYFuJrPkou0AlDqeUqgPhNOAHkQbGa/wj18QvHern
NH1JTHDlg0KLLmybWkzTiIuQcs6mcHjtUKcuus6x8afI3EL3OQmeR0Tgdb5PlhKYjl7p2Eam8085
Q1UF3HtwnlZPLwISi+FUm2iJ0Wshrohw4ZR6CeMuBXS2duOPz9rTorb6Zz8KiwcqTJZzzHqQDHM+
x92VsPTIS15kLYKMJ2TdHDpx7RpLfRg0DumYc/c0n9nkDtlrtZTBxRX2iyRijMJ0F5QosTl9ySf7
CdgBqYdMFjgAMdIE0mK+Vvef2N2VWlMA2K+sAUOT4+Va8sNN0VLb8jsouKMy1hyuuZk0MyFJ39BG
A48idPweBU4+vzDV1O2qtphxgKC3SC9yFHC816HFhX4L3/LPkwoCtm0BeDR0wh9Ge9lP3t/Wk1HS
T82VwWFPgt/BqeAFt+bvabrV33JtY171ShsLvfhD54lGvALpH19MOBRvmnjg+ZyD+zt+52dahFao
B/1VirpON6TwDS/qtHt9KIDM/dCLrLBn57h3c0HxOO/mtOyk2VUhqkbe/4XHgRctEFKbZwXZKBzx
9gRyf0ZUurq+9v9spjrVPaDJJdjyRuMGDro3CO+F6AKHC7bTAp0FWv8rsTB35oRnsBqVEme3UYSA
Xai3M2mvOdfg8+5YoaHXnwUhyvTw5tjJKYFVZmYB7/rWslvkTEIRyUq4Jg2YggdGOwu7JWvUHi0m
YVaIeQiOcz0ftnfu3VEYBOOuWIIukzB2ghXE1x8lBo2/rcmFyf60jaOc2QeWjbCJGlJ/Rn5a4fO+
xyTuFpV7P/LlDSq9LiOCcnHT/wjmGiSkT9DvMBLq/D2Ld6PBjb4uSR0uxUj/9m99vLSmPmuZYA36
HX3DV503Kg21DXxXqASUwuVH+tdW9VmeZSfJ8ZCRCv4cyv4JzoWRwWn4xMT+Br/pLzpbXp4HbVbT
XVyc/BPpYbv75f4S+7xRaA7dldraeduBPngKdiGGWmSrypqqW/A3jwPHuPpnpdnCBwhtyAKELn06
033UuVLMPWokZFKaHvaDDc3Lfbz3UU3hziSrBgf3WDzJStckoVzSrZ4ym7MGuT7zzztSzoG79qXm
dZKszwjoeuH673KTLPnim7bILzFl0DCABxCjj0cVLDdM33TBUUH3g0dGdp1PchXBb8iBFtCGkkUz
YF7U+OlNUZXq6s3+4X9//gaROidTX18mOkSUQUS5oZEr38ppi6fo/FS0WQKJneToUmUNPSYB9jMF
wvvC80FoALuMCKOxDrX+aoe6HRU/alpHOp6B3rKtukkEVIgmje+XlRSAigfYh5YNy+RUSxk+zr80
YsodH/X6ish319a9wBIy1zC4ML6iYMoS4w+o2fDhNTkStd/q6HDBxBgRuxBnA39rXbcfp4RuEqpJ
U+0fq4pUnq3J+k2Mly1CKWOqjl4BDyi+3+Akvo6XJSVyACU33GjCHfT24D8KUF5RpbK7IJfTAE7A
T7JrLn6U/x24RCPoRfNcskxijgJUj1ScxVC38l+4vT+gv9sRvVCsHrEBeA0+CexkWMIA6ZPVFMYC
DhGVzjhP1i1aeYkktmQ9jow4XHpF/VP+E8I0A/IZJ2DPmL19sLJEWdSlQqGkLnyY4zpp5xzc9ND6
3c17udwcAYYxc3AH5G3W8XDNBPt6GwsEM4FzqFn+VLVO/TcNlnlt0uIGC4SyE3Y2s3xF10epTYpJ
ZplvpeZU3qZDIR2fNq8y797Mxj3Na9aD+ZHEIiJjBv9az71uYy6QoPXV+8C8acJ+CAN9oBEerVTq
vcYb7Ttunnon2MZtvLTGcBR5FFA96uDmYvqYPin79KxHYANpvhcqPmkbkyqULNfHTYx8y0sxvhKQ
5CCdz9iXeVYNoRElYBRv++7Ffvd0DPK7T8A/Yj+2MhEdnLvT3FJDceqAIkUZzZYr/aVftTK5ANMw
6gyb7Qu0SP2PzzBnRVl3wqjrmayB8Ota0sTW8odytA0e2/CNt28NJDnyWty0jr00DQYofELywRMy
R+TG48948xWcQWLwA8vWyTMACK8iAXrjJefUoOzPr2sbwuhmBzGNKltM6VPfKseEiZK+gMta8DZC
G8ThKSQAB2kHsV2J2DYq9VadAuulr7psVlr6luMrwXQMgIUDlx+paoiPq69sasJJ1MRQncSNZYgk
V66P6oKa1+vQgKUhgfGTDQtGkxZSR3ub1fMaSvLLEIKWVXjAY2JbMpcqvA401B+IQkY2m2gyXugX
nfFmvP6Zj6qbNKLH1uQRGUlG3kN9CAW66PrJOcemgY0e47TV8TLQM4TuQxtAp0bmDvN8v5JO9OjE
3VIxqNa/QGjgLawC2oPc0G5WYmJQPa/cB/ZqhVPwc+WBBJVEAkJ4WOn106fNgiMrhigLlfB4JiVz
2nvCrWGG10E8n9ot/eQYzMFrdF8pPD4YoYiVXwMDiqrcF6o/oSIak/nl6mAPl78lEdMc1jK2caqT
WO2VZD+zS2rDMCG4IKrtzOg7vpQ10uJkG0QskDhupvYwtUOWCK+TnZQFBw1FgYkplG0n5KBkIAVg
rlObk3BSR6I2gX090E8brYE2ciWTL3SwU57/mSJQJloZhNtNlVX91L8CFQ/SnSlHZP/ggvyn0RJq
RK0QIgK4B9Gs/12GZoRN6dll/p6F5o0ZyGYwJlGVhRh2hCeK1WzPH2ztUvsoT8MCw0seYOw/iKk4
UX3I8VRyZQVDsZBekc63Oj3k+O6NnJn5XjY1mpjAO36L5wWQfyylwelSLBgmxBYlVkr565XC7gFB
tFKSA7LRoJrovPY/gQZ/tSyLLc3ch521DgquKUikc5kofZJSxF4U4/tH1VFbaPumQySCKtQre5xM
8dfbQbp0frmMn4u8zzh59M+F3AWeDhLv2rYoHTAyACofFv+SE2N8F2alEzrMBTNLA3k34NCR0IJh
NFua9Pdrm6GRorvjrnTt6g7NHnDWSBzy/wBgCZWj6SCz/7xWno7XlqVI+xEtlqDwWWOyaM1JbbD2
W5oWn9EwEpcxcWsHZQr/LvmSXrcaCny2LLla0jz7tgFOgFS54+jOfRZVolWTyrc66CXUN+/lJBgc
z1C7ZpR0Qu7GjXsKSicUX1k6UP0HWksduTDFlJMGYAFy2yTADs7zAs0LlcgmehOQZrCu51T0N5fF
rphUcxCML2GKIrBXZS7a1+KCpgXP9XprpvoBG6YA2wmg5BeuhWEIS3IoQmRD/l5A4RB3aCLuiwPf
bZrxAgbppZqVrTv2LM1GSNdtOtujMegjl9T60OjWlJ1qGEMIDRLQqol9256jv8vl4YRzse0H7433
+ogHGjdkB9XZRwrbFYvjUBd3FNVARpW8cJ4TTQLW2p4B6K0XxmEe5GLZ8hmATO+3bUGCowpC+aF9
itymGg5bR1UFrFww9NddqbnbMwranma6BpYpDUdUghUR24Z31kv4OFFLfvgAwz7XbJvmD/fAh+L+
SOwWkSDXEOuVZteYNA7l1iWJQNvup9yV9YJQo/CUIIIdg+rZU8Rbh2V5q5fmYQUMP4nEE2Cf/EXy
ChVQBHTwg3e4w9ogVyK8w68n0QP9/8duA2OiiGM4SatWT5lG8Mnna+1GYbqz72vcf9n4+gVa5DNj
JcClbRama7QyVDk23+GulwtLA/dImRdc8yeqoAx9efvO22HwNNuOo3jy3rUfr0C7mmC4OliMG/o5
ncSSl64MacZQ36rlj/vTcU9JoJpWwWvVqMaXjkvnnzW0BG34N4PfOUeT5gfNRCf1TMvoeEvIB8if
JJtv6WI9PEhKg45r7mL1FUaqFCHKOZxeUBCz7z4wD+E0sKkCAfyoNFP8pPF8M03vcNBOUXda9PCI
500R0nVrAo4C3vTi5Ke3+wPyjRjiXhmg49wsI97UEqLKrl9wqSXYxcrrVTWEAxcRpY7jN56rPV0Z
SbzGzPV6m01Bmj00Y8FtKvtDgR271CRX7lJag3BKDYtqepGcvdTP7Q5XUaQb4o1Up/N/CZkHTVOl
nEG0eCPoGgkgZbrziXbntzTUWKyra7Wc4nqoPT1N4AXZ9OMkDvBQ2g5mqXYJ4h5l+ERFe8O7en1h
VqXYsMv1GgAkN3ttPGu5nisIPDHRu6z0PVQ/ZsEBQ2wBoke4vFs5kHvskhji+XCmOLQnW/OUexqH
klz9jg5iAPC5RplqKtgyFahR8VTEsl7kCYbL6WgOByG25+nckxotoPwd0GennGjAKbjHRV989E4a
hkVuFKR6U3XWJit2bSGLiNRtc2vGM4O5piCIi1WsEkvlEu2iyNitajv/3INJMb8QuZ7NDwPPEMre
sqgm0/fJB9gqfV/gLnUU2xPsPa3Xjz/7xJS95otQWc1OpL7ryzhM/klZFydE3DOtdMzLbXkpEcMh
A7rZVH5jWJRPXQ/jAwfKdbZigBJxqb/XU1R0nTMjEBuUMCNbjCR4IMeIZxuAGK2nvrdfUu/EvUe5
WZSBBqpBxmvj/h+jQ3CNnNOXnknWIiVotU+8j9J6jR+8kq3S1TNKeTMu5oFGz8BHozHJ58jX2Wc7
xHvMxARo5EeKcTuoBIqoYfzJAEkCh8jFkvJmMckPInbgRBGXND9ztQZ6peQai60MzV/FUJArAs10
Dij7q2VEyLv4DDLRLFs1hGwd+6naGwzZPGJmf8alLWr0r/xzUWWNS0yUX1gJ6AcC8oZnS/qAVPmp
dl3bzbwrf5IjfQ+YYkqGwQIpLU3yb1jNcb7+dPQ2pCj9y6liAump+xq2a+rCcMh4yHxAbR+6MGf2
YPGklKh6WyK5cz6jKblBKjpOTf2tJIrQ4uoTt9ZgviAEpgMlvGWw9Bt8sgsL84fRDl0MUTBCDjyz
SXoo33V2KNozJojGZXb6emUrJ4vnKM50FbyfNv1IXxQ2RJP/GHulwU+eATp3PG4lc2n1/AL9eIaN
Ow0VSqRxi+QVKX2cd1vjzD4hZEwOMFM1YdRjowL1HbelpX1C7709PlfVnDdI3htn3KObx+Ow6Xi2
3FpHQV7KEhHwGEwuyqh7PRXWwe+haGYxzOm2MXDmTUfM+WCUy21O9pKJbmrvRxl89WOAGDpveSeJ
IGpxZtLpcfIjksI696FvB2JTQqKgvZfxf+N2CURP8T6Ukog+sjADoMFKOKeA5TbpZ2GbcQ3nAYsZ
Xd0E8c1GVpI6Cz1S7ZJvxFhxBBf4zA5Ylti2qWVgwZOczbVQtmPwnCG0xTejKBH6s0uvvLLdOyhU
LW42jWEnfwH+ZKZHADlzmuc5sHePAgkPJQY4lCo9OCTzmgVq4CUnGXp/rByqRxh1SGJahkLFmbTS
jfPBHwDKuRjDcpgilsMYRAZuYTrRjAi5tiVJ2m2IIpyGxKHaMwEr8ZJyIcsugdmijcYNoCfQs0qY
jZeTPjcNNPCs+TxnpQxhkU/CpYcmSzsxOYaY6d0m2PUWcg015TBZpf/1KQ4Id/UfM7LRW7OZqYnZ
dMnQAUmPrv0hC1Dig1kj12TNkZ7dIKgfdpMLgnpBoz2YTVwpN+ycFuoN9ueBu25Vj3pWncSaq575
nO1ie5paPDkTtupW6OKyed6L8sEQMgbBM6peWrApyKPakOszHFQyXHz2BrifV5NG6m3mIjWp0gGK
mvlPapwy4G+rIKXfsAbGzuEsSk9EqQczJhB3kw6dM71RCl18oLQlE5b9e5TaJ6IBB1rZU6gsH8tk
InNUkgcqjvHqaccblG9Di84UbXruvzPmz+zbHM9c6BaBIWDGLnz0uEHoanLWylWmHlfOcqPq8kYv
5uBD/i7jLjVN3ND9sfLu70EnPlvYEZBQDQjgqDUMSjLw79FzF4Nd0e1tumwcHYZBBCjbIDMCBzKy
SvYhtMpBKz0cXa9hM0/kMByIHcdRYPXtPVfM0vm9HUHflW36zQxU+0LdJgOEBXGmxJgKVuCnp3/f
5s/pCL85yeNzE2qKnJdSFbaTq9FqLi2Hu9yGZqU7OYTWfxJMZXdoCPaKvlSuKtwVwrgLnmwVDAy1
HOGYzZpd/jA4vVgoTwNZ4Lno7IEb1XqUwqIPrr3w38+Vhu20G7hN0DbpItGVpL0vi9mcyzNbm8Mx
JUPOsPYJWm1VnDXOifm4IECbkMVi1qqlPWzL2p4tuliuOHJhpOJISkac1Xn7wCWB/C7e59iKpZDW
4Y8h/cTZXJy2XhDvDwpxFW1hnXHloTJkgBJXFPpYNRsGbC7tyVWhwXWzcAaKyqbJKrqYMUHUXDKP
AQKIRLpEicPf0BYj2Q9C3/pJequ2ipsGDGKKKA13ofd/lDXy/htPypvh05woxpyCX5ybwzJAO56h
vHkmxuYz1Y2A/HAQ3pyZiqktLNJur9v8CixNZb48iBjZXWRS6y8LPsF7zyjC5iqgjiOkNTsV/1Mi
BKWObc5v/jxPc1u+je1NCONWtgymOBHwSLI39H1rBb9BJ9bcHVFc7BTO7WgmomNbi3yaF51OScGO
LAXZA7jBivloDVDAk8USV1fE+RRnBv3N3fvyP3RmHrsjm2Xldyk+dKNXhgnyDrJgblXYvbe4YslT
22GJxvgoStjWXd4MZE1EhoAIWoaUxRM9Q623YQ3QtiIQuW0x+sE4lFO2s1kwaTR2XKLFYEl8utmj
tOan4XJi1tdwzI/nFIGQfsUBvmMZqEOqtCUWsrmMjTsQHSbunisA4ITdOCxjLXBIAFHsD/BYwUlF
fmK7WaUTU/XzDLB75UobAl+CfJNtY4d+Wlb6CbWQQ74r0Kpy9HfoMWgzex57SqOhbdg37Sl3CKY6
h/nfYFCgvrwcoIflD1AmJMXkYS1Ff/pRT44gBcjqe67bobsO3AwxleqyMY4hBU6ggJkOTJ5+OWKK
6kUsKWEi+/AO4o5AnA44CwmwuDcoC2jX5rR7sIP6xObr+dAf62h89V7PE8+M04X6YJX131tRE1wj
duc+KUswGXxX/tsvobk1nbuFGbEJgel4cf1qF/g2UlgXR1H+0r6eL8nC0Jly7pll3vDwh7CzKqMo
ZYHiVw/QOw+vjDtSRm+tY8QRF6GE4/ZoAOb2qapEmg/blLFSFjW7Sm9/zfjjC4meQHbPRYPnt8YJ
tG60e6B4azdd3YqD/1rkV+d1rxJR/8LtLW0hsLWtX6WwgCoStTxrK7LIZaPhugmgHPKz7C88/KOY
4b2n4O8r40Weye4K6i2ENkwF+Q2LXL99enorj8maHYPEorSYLci94Pjf+It1o76rkPcqDJakFTw/
n0jmRyPbaKw+Ooxu9E3E5Lc6OuHga8m5rgk+3isv5OVXgJpVX5gpG0VusxkcstoFkjMeDUuyv7Ir
8qSzgp3owIE40J759Euzkb0OpvmTlCaK5OgYw5ZTYEtcdsJqJPG7xhFTPd1SdgBDq0wOxCzyCbuL
riH7mutf5XHapRK4eIsNTLJ3ujSFsWm+miMREF/9Y28+c89qvk9PYpUCWJ2+ckdaDnMB/XBZQTg2
gg+K4iVmbx7F9j1rc8aj9loXovCwM/j55WuvgFmEosDcql3P2nFTnyudBsdMrrf1vyhtg/hJ5ZnM
VjaNN7qYrXfTlcORzP3WEX4qWobfdDyN611hi1uZe8vqtXKHhTwH5MjdNvKn9HNEzMqYZ7HoRoNP
s641WZTblpQRc0E9wL1uAavUMqXHLKA9f6dPjOVcUMShnPLlvF6v4ET3AZyk3PlFFAaFJF+PW6bz
R5nlrqrqCDvTfXPQebhiNWXrKA5PO9a28mz/5h8tMsKRA9PO2KTbvsC8sbPIQRjUaHm4qj1QU04o
bQVYDX2a65mopyVXB44k7s+SqLedmIb6vvWZ4wf2aN3URNATVbBduVhi2urQFrQ0uthcJctiEJxo
uk2+Tpf4CAwbjE/Ke+t3aVc7GGX9KvsbEW83kVDQ69fUa5JaBqBIp6TPT34L1onQMUXSsJKF2TME
3SLzfFDFSsmQszupidvuxc0m47Ns0Vd5Q3zng4Z6SX7hvtE8aN15DRTt1vrvDgdzzNNx20L82mzy
hKK2s/wv5JofGsbtjCYhGI73WP7cxbRVJG7JlMXhP/XRRZ91Km/gwehF6mlUwahPIsIoTy8eIoQS
szgfiQygGieVnxBUR2YRFMlav3wKU9Cb9wMuowAcp/m+RX3I12s0uBBwMPuHAttZZ0goUTmnUdKz
IUP/Hbkf761MwwRzz6pH51uIVsoabp830ZXscvzfADEmIHr7zt+ozSOUpkcsVIuu1ndAkGt1rpnP
6msuD7zFSLR+rnJfUdvWdRmDrrSvU1HdTPMwKj8sEF9fuiDpBzkCE4lD1AiXXvtYsR5QlbDd4qMV
CeU6W4vCE8gZ0tuewraMtDyaBhhyOC1DU2ll9ARnWNPaAypSrE19kj1oouc8+yv0VlIhi6rm1vMj
qHqMS9jb6Ur9coINVG2O8ILvFScfjcCXpeNS/tRgShj9BETVjOKdo/fdfR0RDptR0A0fe5r4fGG5
co2BqaZLBNhEg7v8eo/QGFercbp2kozGB/Trqd4r71rWZ2LsviQkP90gm/mddGj2YoSzn1gw8ui/
e4hr4FKa85elZrNjJZMVNaczyc8F5Q50LlOx81NcHrjelw6lIj8lCIiuadojqioMFByg8LIh+2jJ
ZXaCMu8ny9ZUMRworQE9RWX9OthrD5svus8iBvpIjTtX3gYkIxZm9inSf1cYYxG7zPWvZqEN9ncb
uv9pTNI2wYLyvyk4+LgAM0ps7W+YjSo8IgMgvvgsfM0NHGJpLFzj3txKfTG8NIHG3PsJ2Ww+MPwY
zvPVf1C6AQYn8rfAHlfNUZXsMxOKU5QeNXCLDh41btjYnjbJk7m8whhoGz55XdB8ivY2pG5mQQD1
EoDSi07qL6Xl3nGHApBExIzgpRQiW9bjHT7nJhlpnKJKUhNmUvpSkel0Cnkc1Q5oLkUBfAAIEGf5
wTGZRL1TIdMt8LsutCoHqWYCGESiclzYYtJuoGLfqovgJMocyp4W2E3FdY3+WiQCDnsRrK2a9xuP
YWFIKwHtvhdP5DRz5x9n9ytKUnBDEJuo0nygKmn9xr5skXGyoCzuT0vE+hJyk6eDS6sw5tpUYs2p
IPNNK/tDXjBEUbh3frqVs39g39iAfu61rrgkgxmiciETCd15o+8GYTb3jj81ya8Rzz8JaP3M5lrM
nppEI1pa82aYfb7LtuVfWLiHxp6QD3rQxeq6e3ikdfs4OnqDVbRtcRbd8U7ASUUqOFdvNLApeV3M
MQrxSGNo8CmK6QgKzNzfQEKZOLwF+6VXR8VMPC5SmAUeGsyYQh3/t5WYd0zosGaRMuu4ui1BZib7
kPeBSCl+U8NZqDBRobA8K61JZJAQSaX9mzeGcTS151S3bLaTWfvRSUFmdtDTmoMOl7L3AFh/5tqK
d+Y38DTJOYclJUnKoRTXxUT10imREZxCYx/dZ72HO6q39H4CuSL1VUALX5xuCg62igG9xkCQmV9j
AkIdSmxvbQ4EFkR6AsfEXvbuNF9IU0DYToHnrLWkMJlyGD/g8dQQNzxjE4kqcao6bonUE5IBmoKE
uKWesqp1359XI4hAWN5ZcqVuVeW5xJuYSxWA0xSgVDhkTx8dA9meuzDeV9lCG+fV1hYQOtVuh6cS
WJaTbEma4p6t7tsQana23rFcUfc73sPtm+ASJ81jR95R70F2me+Kq9Em2PDdYu9c60sr8ke1w9uK
W4/Wk7SfKDBRUlMLEI43Oo8eBrvzOveZekSp9L2YAZJ0tEDg0MC1vN0RFLNsWvRoLCzQRklXYIfU
hU6F+qZXdh9w+q/MnQjLK5/RNoqjeJa6fG3JZnckSb0HTnVXmNF89yylEtd6Y+3wZ2xn+aV0oev3
9AeqTJ4lATsEL8zK89S4WVhOYxi54OXVfWMJdBFZ6GsKwKuH2TSR0zQ0FeV2uQIszvD2XPYbOhBl
I7vbGe0k93zSuyniFkBCEOaPS8I5P00xbqZWa9N7pz3g4AcUQC8JaJY0g5avLog/7wl1ipgfCFMZ
f66oy71gvUly7TKj9Iwqlg+IjNnNP1tyY/r1tCqvPXoY14QtdK/j6YZzZCNTWdI7BfwUKCDFP+qL
ci99DzQT5dzhDoz5vdVdi+w0GbilN4MmSn54ABxAQ9AxDQP/ImYpZE5QVlVCuTc6uA+iwSnlLgpl
sHHTB/pAKLn6Z8UXKpJzVdAZ+k24S4UYHRdMTo3qwx3F3Fvlni6GthbKrndJM7tD6itkgRuihhI5
eXMhu4nH2wr0dUa+gEk1g9RVSukjETLGDAS4q5HKtnzD25R2afaemBXD7wno3F3TBf6nqzSxAmXX
a4ip2xCqU5fXFlFQqkdkVtSTiE9D4EdYUQiWnzDptsOe3Ycx41H2cBulJYVJ49i9BuOEB4XxtRTO
vZO9bU2b+IoFsdMaPXRYW5fBwqqqgTPjqntEyChtGS0SKVneFqY9XeqtB6ls7Wdc/5RK1SWK7kz1
81KY7XWP98Zi3Fv06d++DJgbdF7RxJ7YAIPb6CDBva8s0qL5QYSy3NSHxB3vM0VEesUsGMuDAttv
jFp6S+6fqbQMPqnx4P8lsuZ50ITGH02oLQEUwlbKs5alr1kMigzZr6m6zRtv3WzSp25dvo+uodpx
zedyZuBvBxxRCp9SCUbWW4W9EK3PHZ8yRnvDeUSDck6bMdbcmnY06enMSuyh5OuoODP/gyDuVaI7
h15kmewPeyaIdaaroRdk2BB5jxVahw91ISm84Jnq2UxVLbWjUQ4VZxa1R6aK5SduYM3ZUIbqVMm3
ozxKk1ZcPLGAsdNYMk6HQpu7smIEeSJv+t2q8KJpXUFDR5QEGHQPvGXUlyAnrJY842e/GLPJAoo/
nezUvSpPpIN6dqbO159JZVhJQ6trJsQFqkv4blncGmuECWQseO9l03JgHIEMZjVBoZcKXepkeA3Z
PVTtW3nC+/hLa6ODbyfr0rymzRpKJS++mxYXpTHfco4axlrRWleC7R2zdErF7XD1zu5W3TSitMOZ
/IunCtzqdCVsy9A3uWhdeM8lPvHwq0kPzh2f0Flp8x9CscPCd/aWw77ywIkqh0jszoExGYHfes9a
wFL5lUCsKkqNQKPAJhesp97ohe/isncGFf9kZCPO15xZHAMyI8v9YgZrnjWCqR8ah3bmqua60xV2
leuQTeMwTk00PPl/3ZcrZe0DYLkq8oq4THRT7jjwlXWP5JPCORAzO3q8bcGpn4VY1y9YRR70gavW
NEpeo59aUXKH/kTiA+Mm4uriJoPAKvqXqxHXwSug8I0ayyCMtGHWlOiwarmCCkaQ639Coba9zcYa
cpqLr/mJJTfRLJVyNldhKQY7W+LULHJKesqyZXbfN8ChONoaVo9v8qzB6xuFopvDTLtx9dTNMmsQ
AW7IDsuA/EMjuF/c4UxDTdULxezScjo5pmxx369JCFE1yxL30r7+DotMlXubbumSA/qEx0Y4tyFr
G+AWva/k4sAfcMZ4U/MlxDBsY1/FaGNAP66ka38O7obYoQGPPtHRMPDi3+Iav5kDix92U48w82m4
0e/1S46YVdpvudiljkG3A1RB3+zr6pgQYIF5JkAmBcAo1mYHjk59i7q3kms+k5S/B844o34O7l0o
wJJ0PdBVsdgEgyZ7JtxZmKOHyE9Mg6bDhdCHguaD4ozVHhAMfivW6XZazIcu2Rryrv/P3OLPZrWK
USNuQEtDtertcK6MlLXPMe1nDHi52ZC30cw4j5kDkhXmGigue0f1/qIsUISe3cJIEFl4pTHmxvIh
2WLUYIQAS7eZ5wbrsJLwlRuqJ/GVkMaaXsjQGgQZzPP5ASexgqZRvV29Ih6JAlhilLgL1povz3B6
jJzc+hEb+PgiB+gSuFzDKDiP+ACWCj+P232kznnKDue/N3v473D3pv8wUDfVr1NKMYRTqqzL3tea
Q1TnC2pjuadRPHuqQEIt2hrbl1otzn5GJQkPpMBOE/UXjHqs+uP9nZ+0HhIG9uB8lFQs20J1Ipzb
84ROdK8b7qXjVYj3zHT2o2+MN9WhvWuo1yTgYinlzOcJgzrMOl4hZfWqWZwMLm70MH37U7l8PRJs
utAqRGeJM9U2P2Lnjh6PL4UyYVkva5yLOAYEdsaQyhwBUJESOJKx6Zjkyw2g5xsTqP6yF/4p41mH
Gpu6FKcWXbOWMfBqV4dZg9nErtzDaOwsunba4iSbPLvM5kp7e+sUYAD14BhuB0kx/URJgcjueVaU
hIDxoTeyIWEFV03ncRgOg0eIZzSCjyZzq9A6ckaIb5fAcshP5KEiSxUMDjet/0ByWGMfz+qTznbT
bsmc1gIlIK6BilvpEf5eBV1moiy+MvsQg3gbCGW4jnGLw53pj2qzDh/J2kDJCy0HSM06TTjyEi7t
nA2FyRRQoTWrutL1VvJfSqxVt84inMHC5S2A+G7MWH1+5+G0NCNkBeo8fglLJKnnLlS1bRIpwZ5u
TGcXXIGBEDshqu+DpZ5csXU/Cf/zf761hTdVIxOLjlAEmM+4RA8DeNcX7FgT/nL90BgjlzEtk/tc
o6bqf+toxbN9geOVnxZWjs2mttHu+Qp2CjknsQg0SjInJqgXHmjv30mtet4ofJof2WudYv8Z6Z/3
JFIAPRo6eu532mWRQeksF96UDLkd6+lNfGifVw+p7FLo9vI9xVjZs3045atuHqHXJ985xoe36f9L
rv08MN+FIPcrn8zIxCzltATyHSO+/WyVviuqjcgK+m44qvyOreXMRznobDGaTnr21r82VSUqft+E
8XKQRFireXEXsRzoOxudnNBSbEvH3+9FnZ5xn5Sh0Za0F1FWZ3paBIsObbFRuFK/Zyjysf+FFnaY
ebcAUtVWZ874F6Wsu+hh5zIIeYz379d543F18dtp7Y6DDXvn5jCtqj2dERQ1t/N36uqDHHbM1pkY
4g1EMDLmdSqX0JDszeH8+MFt8vjUq39EhQcoIyL1usiwPI4yDt8mkaO7Mtc/k4sYuT+91EXKFWsJ
bcWh7+z4CkK/MrATFCPlbPd5zQWzhmYSBFdCrkeQ2UhJ4AdPhpw+Fk6oWqynPMzfckMDgFWoo9Hl
lgzqfecn6pJgxv+3l4h8UUFQEtW7a7oBZCHPv84vNSVzdnIFFIJhP2IVBu5593A9MdDgs9DE1L0u
s0TBcJFsREUr3f1ZAGohZ5mzc1zO6msHeOFIOjd1EKxo4zLcenCmBvscZPOQ/lEs20OPlcTfAkDL
ZX9gxvEP4+YV+JDmgR64ZjJJHMdb0E+TSY0gxvtUE+qL5a/mGHgtaen3bs9j9ve/qw/GQMu0rFFn
LuNWODX2mZX6dNU8Nh8AeXCu/oBLy3JbpBcngkfsw6IPIQE5esgbO89fjjWP/OI3mihCVEb1dgOA
62/NFAT7j2IPRj3uoANrYs53IYt/BCP7akOonIu5C/0cTC1RAeNzuzyPVvEZktBRZETjtgL579T1
pX98QgE5EzBALO/VpBVzhs9s1fTy4wP36GXY6S+PXhOsjrO7ZC7AuEURsbQC/I3Uibg1qim8+dCX
h7laAfu1YVUMu4nx6+8t3qZpcfFcy4y4RAP7qxfomCYxW+BodZ4Gbe7AOJwn2IsjHMwHQjf7s5M/
uiLyHnBKw+foIJp5+Ljxt+FgE2XqmTg5hbYFZRPt+1V17VGf3UcG/W9nkLOGIkqnT7GDG/UeMWP7
LgKAq5V68A2iXbZfY0uZZSwMlWtCbWbKd2e5n2ZnsXYuGaC/s2AwzeoOr84Eg7TDE/6F+hCoSAPB
s8S+M8GPKzPtay9XuSnmVTpFSsdwOAyAELCbPgAQFh1yZc/epmWeCcbEA1Rtl9pMl1FSiNrGmjiW
AQoleLYLuo5lbXNAkwcuXDrw7G+ZmQhpbnOUTFbDfhE7W5BxKVaOQhstLtX5BCE19xj0vTyjiwHg
O8YqtecGM8YHLaqSYYGSINM+k7vtvCukboZyEaPsmidrTdQgH/g+pZqgNmBTdfqOmACIJXijnLgH
ODq2NRUDRK6buReNtPQRVtAmDhH+Ad0mtISHhIsnYf64R6l791l9R6pm2iw8Ab8N99pA0sqjCj99
HGkNtN/8fXhFgbBipS2c+YGfqfC4ypp/rB0giWJ/wPCs5M77Y6DzxBO6ltfYH6ZTTewyw63Ir6V2
ke7NpuImUCcC26KKBllNV7KUW7GtMh0Venm258ICYQc3apknBuNHiQRY3XMYLczuemphaB6eJXGo
LCfZFAHZ2r+zrUOVjpucEZxhpcVqNhoaQDsi6Y3hUMBnx1PF2tVrVp0CeTiYICF1EcnSTs6rXZ6L
JxchlnU0jR5d+WClr+TIfVK6N86dW+9zaQtIKFMyhPRGvIXAILziFGeJsXnXZiFB4FhD4SGnVIXz
4VUzwL1A+9yjwh3AfEbkJ5W4bxVmYFK96GVlr6VJNHghKts0kKqVdEAhDayXcdjunrBV9kDXbFGo
3eLGKv4mZpfwjCYu+7a9TDSODDx1ptT6a+zHf7ulBkAQjRD4G2rJPhdWcAcNbLldgGYONR8ilI0X
jUq77COOUICfMyITIdMdYeq9Hj3cFBPiovd8+6JuyqfepfAbCTvqNNtIcEMq7+lCg7SkI8nKaqIk
QssjeIyP8B7ikrny+RU6d2vVqxJkYh5eCx+8JqiG1sG7EePla10jUDvT8FUsRsDja0TF0u2kzkd8
wcJlyqZZueSvGR4gQF6DGDdRsyWj/pjEjXj6P6U15am4OVQvEEgsVTy0iBTH0fhiFVcQyWuW62Li
L3BzNMozRoiGo1tDzmqVfS6HI6ppN1iFrokF4FBpHO0Iu3C0MKe34qT7/007x7YPBzzjvtmWZVYr
sCg2cnkUav2tzlJ+eNJxq0h2vC2sSl3Q4JyJWzWCcXI1JKU44zrjtN4Ja0cPf2nA3RYzmuNZi/zo
f2blK3ZNE+/KxzBrjCHfGX9iihm9PEmOR0vzI52UKXF4+LXLsmNsxDHRN7VigReiy6ytchx7fnmD
vPEK9dJkprqF+S9Yu6EpZzwvX6pnPDN32p7wQ5s8zz2fAvq90NuhJcxvCfBINy0PBjLeMZOBQaN5
/EwB2IlQYD5ne5D+KDe0K9fTMKQlIj4EChiW5pdUPhG0lmpd/ScpgC8sWQI4lQp0kwdHjV6mefA1
SzGcprKX5qKd8K7LTb4Zgs+JRW3VD0+n/fs8OCKBTOlUBG1PhzRzAVRr6HLL2wM577xp0aoV8pTQ
6kZyeOrKCcK+ub2fOguULIMTTqWVFHLenzh9GVDjpUkxQJe1hX9NNCbEu6bOzQgM9Fm/N8oxiyTd
SSZTYahTIchSDR1kZOeNtrT2C6/lSx9sZkyRITllef4JfBCfN3wCsdZRmX9yh4LQuDOyF616qNlV
gVBkWroOY228Sz8WEaH3H5X3mBv3ICEhd5KUrOwDZDnxTb7Xysvy6Bp0fEADlXZvYg7N8tSQ9wxS
L3ddswCY++yFxTvWWyKKyJhGyfdbCp7pW9/ryqLJ6xmKRMY7AFEtzmf+tGNTINel90OrnT0nSeWB
9JbKZ79zfjHFWUk6fJe37ngi4NbIM0MUK6cI5QbMmU3izI3BekA/3wfMkw9oxUtsSNOVsrTXq85a
yYl9Ft/Y05Sp1Am0I/+dKsMoSCT4YdgkSL31fqorQHbu+miJM6Xkt1rvAD/a4BLCTegMrSsx2jpL
bGuzC/yiYXI7WeHlruK7S05myQdK95hoELk8u7KRt5oJ5nNtKYdYiH2oaCfBaS3UUD3i9zLa1dZe
jrUvoM4hrs2WgPXfXYjb8HfJhQ9QUjoO1mWKJxp30XFNMbq5kXzYXVQgfrP1EDnhydsGXabboTms
5lZQEBPeugmGxWPwkt9Vfz8pbwgIZpsprAldG5vAp5hCHzAczAl+e3NZQfeI8LTfFO6Mw9TnwkpF
l5rHit8KmyHmwT4RwtHFqv1VH8UauU3TeMUXVKH7u3ban9VE72FP+kFatu6hTZE9EZ8dY95Ux6j0
5QPzH2AFOTmXhyxzBg/BF+mW12T8r7qMMW0QtE0Vw/TBVw6KEBeg6F3yWoQYFTaqO4YJycxFjaoG
0auM6ieI/Cqg1bULF2grf1JFs6x9OA5C/18AEXy569XigWN1ElSV7hrEsh1gZh7dtFzVxwFtjULc
+DJVPvR0A87I59Lg9ae1cbC7ksS3YW7Z4PVpypFZuRQOiHf41qAZMOSuDa5TDTjfL3D3bgzvvxyh
NAf/rz8B7rXRiI9mI2X8k+QI03btXx1HlXzLlWKluil5+3ag6VcDK3Ec1zaE8+TPBW4tUhSWp9DG
JX9iMdGcIP3+UN/lhoVjD/yZQSORYR0ifOc7DDWU2EsT+/PPrYRnU2vW/jWJATvSZlMsUVY3ni2D
azEf2lt+TO7UW2WzX1rmx4Ok5dZalwSqikweI1oTUPWWtrdq6n22YQVbV3kwEj4dJp6esZWzkQAi
aXUcWoZRZcc4+VgXz/gUUiu28A/XAf0fCLlyEFHOraVajTE7eDoND/l9butKHV7r0NGM/jM3edo3
V3ddRKQ95pCh6I49QJLWRGToEaZguMfgY/jASsFhJiUy6EUaBlNGHv67aQSlBgrQxjj0fyEiH9yn
L7CNUKV42RiJkoECYNyfF7Kcx86gitJHGSoGW0CMn/M+y9GSWml/cgG6gIZylEYkjhraAlpJfk54
byY5cJZ1uE2IU4n7Bmk5RR7aYQMLP/GrEaN+0b1QKtToHl/C5SQmbWnnmQPP4sbCwEVKKe8nQq7V
vOBSMJYgkMrZEQArpZAp0pg9YPKUEEO0g+m1DTPgLW4Ff7ARivH93tnIolIPDFz5tWL34v6wIo6n
px6KpWqXkjA8KMwv3b3aLmYWlZdhPeVbLLe56M8sN7w1mMS4JZqvjN8EqdMJDOoKFeSCUw1v/zzL
0d8ws/v0UhB8w128gVmo8FWzaqtQj45iZCJ7E0zLamj5677SYexx0cZvyAfeF/cTQDZsxrI0KTin
L1WfFUdF/L/ueE9uf3RzH5TcGrxEctb8vvAe01AqGrPhMhbfKLxpCgr+xjPKbP/Hv00uYulUivij
p8S880C7sGKFSE3J5GmFE7AvkpCGpLPca9IgiIV8Czr+Iq2zi+GX3r1OULzdET3wBfBUwloX6Qv+
29fyciOLdq/TIhuORcC2Cd+C4Iu9Ci+9Z1HskcF+2qNLmZVSQOuJLaZ55hvxHb4Q5ekOsdb8PI4T
k2K9hYtHgcz7l4jL6dGSzK+WD5jMEfIuyl3btOipF1JMJ9PV1ajmexIrVnfJyS2rdTB9JwWWJ51k
ntzVWXT2yBICMBJrrMtRgRJzzdfYDj4IPceZD1gbddBjmAlCNHqELiVczN8f14ojn7fIqvMVe4AP
A/6uH2Kj5aFLGlJcHlYqXhUGmrGwZgZEw9SUgGV1d1HRbt65kS0BS6c71u0EqLa7cOhLMQyumBf5
U925sc+WnEs4w7y453NXhdnpk8HJ/9QGcgXvDhHH3WI0cm2DZ7zZVOl/x5C3CKD9E1ul5UkLRK9u
+WGHqMmW/rYBv2fWrROjZ8N9aWjL6Hd0KooiWPEBdaRhgaVN3yjpbBTDxQ9z/vPRqDvDQ1Te145K
JR41U8ZQVtEDa4TiLx/C0RGQRcWp6TQVWvHQJxXJYrd6Am1IDW9bWa2WjoCoNNbW96F0Dt4QvV0I
tkMD8+9pf+Q434PKVNSdZe87S9DS5DWDtuF6PwXlXFCE1Jmp5xGfVK6jLNces35kLTpAkI2ZAkzb
o6+wE7ONUnCT9PHMwli0wj4fc2qDMNWoZAZ4VzUj8kZGIIl+1JG0WCKSGKbooVdGTs7P4ExC87oL
dTBRH0CCTYNeH9+Zz+lsrESY9L7XEaT+CCBSl98MJI63qPH0Qs0WGzW85xwhp2Q8rEGWo95DZrph
45pOCwrDwTdA/YUr5FSsgRqHj3e8thZk1ZdcSF/7edry3Lo1Rf8SiUgmYfPTQRYTQ/U+omm967vz
3X8oKDBPHDHVbUS5lUmGBNAy7nHJtlEYjQZFS42MX49smGJTCjNPe1GeWuejfsd/J4ina+1VssJW
icvnGuWIaF7amWWghOsUT3zVORL0fBqhWjZFYuV9UGOcK1cltM1D5bBUfSBLEK2CVerJnn9CGD2j
3p1r0wGrAzqsZLNcUgwWsMPZYi+tswsNneIiEYzR1+VTHfP5VGB2mLN125tQL2ApbaUwjN+R2PLJ
8aHAwYV5j76JEMLtQBGUQjdIVm7s8ErS0Xc+abj8Fsx9GOf32rnM+99Lvw8wqgttn+OgTagUIJvW
rKFc5yoa3gHsj7QMI2yfjNVmb5LP7pr7ZU75boEGjnaMLk54+7GY/SJnKochmNijLsSSL5cProRZ
eFwUD1sLzTECelfnNK3DW3efuQ39qZ6IukqZx0GRtM43DnFyCAfPGXhv4lZw7FYOXNP/lnbV77XX
N4sci6TDYbh0OXyu3Y1HN4EqHrvEoXrB6oY/FmOGrR+j7PkbSp0lvUTV7w1lZyTkzYKv4U/LTgWj
L7PmLHuLjUnPIUUqy4oJNunKUR2N8WZ/j5Vh4AFmWxcjBDx+JmyarWaqVeSYksAyk+zNkCLQjqYb
sPPAzVUlC7u6L4aUO0ha44Ta48vOkzQ97fQ/MGsuVCBP8GjD6KXb+CzRlQx/drjdyojQODk4RE0Z
BMeqoaCQ3PzRrV56vnSPTXdeiEOLVpLJOaLm2nCBPpibRmAmtvSmlAtBOaNJweTHfO9u0K6fvZp4
6YchqiFsqiL9s3K4ikyLyrwPU8FT4i9tcrhLT75uamySvm7zGZOEEkwqXd3wdfT2gmC+WFKWT6aK
JpzuFxdvg8acVus+1QT3YxjINMVYHblX3o5FGexAocw/JRiuz4ujByYs2wm/M8A16Cd5qeTXEscA
4M8yRCdy6M8XeW2gVx/KvvSEYRbbF0vjKQ7eASZmlXHQ6FX5+WkepIdYSAFBXVv8ghAOzTZ9UqBv
rxg2IOpsjMs9dzcx5qGIdjLM0aBtA8lAYDg9TeCmNSnWbv/h7TGsuTqtrfLFaF0A0/Qi7ttFLA2V
YOb/RO8F+9egpmQcYhw6wbfIbYwczIaHmKaG8LchL23L3LPwjWd1Lkg2XzftsuzFLAJqjfYZGY3K
5tFrV5HEjPvhzkgOiSv6mjGazsYwquOFh2WGSt7CGj5vdI44+uumscWvxKQGdac+7g0dOAsHiroY
WmRwREiW4v5Ou6oui1cjVxE6zf/1htQvmrqhqpFLGCqv9ZIxE8oeuMQxlBv8LJbotEwnDLLgsnfI
3T+3XD2zjEr7i6gFsw0Os6aRHUbpWSb27l5dj0F0sQ6hWdNT33auIUfQTSl+P5g+YwuI3Vyvh7Pq
RIaIRJrxIRN3madbEYkDPyzCKUlbF1qWT0Svf3mNV+1BpTKfptsK+lYFYoidOFsUiehWhOsBtNHl
wZZlGwYCYnmLHClbBeNqaWsdLTPm7MqygCdTMr0CGyvUtMc2A11UMIPABlVnPigl0N8O4uDw6/cJ
ew0ycEWyNQ96/lSOWrVapoWAqAQZysomnn50QjWJjSQrpGbIuCdJAKY7VGyUNqNI6zP84DTot8zz
4AFRw2A62LrHp+8q+qTK0hEaznMqnRhEJKCujRGiroGmfJNfHZ6LcVq19HbgVPqfviGGZrDUMD//
0FrYWGwxIlsF9RXTnZRW4s8OLhgnuXeWfmE+VIqgTD9USzhr4nGfApyXRKwk7YH2FNDA6TDINRWz
3aMpjyud5zjXIe1oAEyP3hQRA9RcnCc0vvWYpI+FO9LxwepoWtwpnOzvV/HlTpMclQJOSkcY2uT9
ZBxfzvlRZFz/mAxdSL6K+soFBJY1xG3K0DeIKZiDUXFROiuv9sCfRRBUNlH26SGFA4S54XHQ8doO
A2H0/tr0BOs8VPyGiBs47vt5cxz3Q0pnerM0Ptq6nULNdq1rh2WaAYIHVseBU63atWjlgMC1nAux
sWfwQWhoZw991c+aAcSbMyPTWgm+LyVmy9Sqw93cajbpeDYjT4tlNZHpvvx7NORR0YxvNP1ekPDF
pQNryQfhhxqrilAQaAebFRSY1XJYSd7cNLcRqYY6K0tFPzKgOIqtPTKUG8xAeRfIfyeSEnPwaT3x
6rGz6Wtyu5ahVuqMxEFdqiOi1696KFLWR4tytp/QpSUrjml7P8jP69qU1Gl6w0C3/wG6UnxHkQmb
YzDuMdSeholz8japAcYz1qmkRZbXcnAuVPLaOCRP3x1/xyo3bizok4kd0rdxi1BHySnxLHyFJkab
JMIL795i/ILT6U1Y27Qu03eZ9eRjHwbc7GvO9Cqy/srOlWDRbAf9fTvGiTm8m6HhEvbOk7wOfs6t
2XUfWj/NDVyvmXm/u2YB29W9EmUgPBVxp36dHmPIpgMZcLm6D9me383pd3Hd81/e9Qw3FOdGgYtp
bD+lPpDs3BToyoH5BPq7Mib/O/z5jLfhZT/9ozqM0pIg4PY6E/ftASNEgV0DamHZR9C9QZitLm4G
XYCkKL6Ar+WWLrJUB2tRVsNZ99vzz+SLLXsM2/I6GktyKJ6+UOCaijUkkKGSSCukrDtGZRdtB6tb
gkH/enyllWXqUJBKYWKQfwDUk/LNPJiPILIx7MdYQwDD3DnC6uv0pE5RYlkBTY96tH6jBM7IIqDY
ObRUV3/JYhjmICeG7oUT8Uwtna6Sx0krIbb5zIzq2TRwmGT1ZZ6Dgi7v4HfRUCwb/8OBthqv4luU
FjqbdtpuWE+0ceTMnrOs4+PBSJ0Xt2HMms7NjjA3aWrXcuk4uYdgDydFPjdKcSkd7K1JgxGfAt0l
l3/ZUzHvijwL6/V2sTejq89MHURvxa2tSorEuFpupR1K5KDHqkj2NhLu7kOpo5//oHeJLM8iAvi9
vyeiE6AOkwYWmt976VByjj/JdZ00gjAIP08jnhiU7yioPEojgRkzQLEfw5yUHyQaSA0ahpbtCCsb
RDvJbW+CfaPWbn0yFa+7f09NbykNV7pZg8ayiA4D6gMQBvrWljM5upq3dDr5QUobWu4zfw4JtUWS
s2+Qo2HN+/sY/MtOjaBmPtSCqujq/d30EUSDEkalXupGYEaUuN7QDbEHvNtdBNe5NBgUlwu3yebW
TCN9YzwgOS3KKFvpzJSd+G7oYQTZQ2sfW3BUBY4rzO68BT9vZuTGc6jmN28JkoIkXunw5ysuxk6M
UJm6uspzmk37V5bHbl08H++KZRgsB4YDOdeupm+zqo1IKCmONARA7FheUcAitX0crp71vRhPFDIb
M4KHdIxfawrddM5OqrGTGvTrvypyWGnfOxYGuOiGRUC+kK6CiX8j3i51Fm2J1xMFXcj9fcLekmNq
IIbKFQnSZOyE4t8grz9hvxcDI6s8XX4dVGaJXMdVOD1e7wFrQPHlf0NeILDonjOo5Iq0XhwmvxLt
FmN7CNSmt5FFJsHTYj+5mDAN5/vcZdXYVvaiQK6dioptdHxb6Vud/HUi/9r7qGhCJ1q+JPNpD7B+
xLGjzMAQjlT9Gb+lxoQRuCZr2fIsuUip0rWBGP7h8xhn99Pi0yD4LS7FDXmMAqJyncl0Ut5YGOp+
zWMpLKVMOCBUlP6V9rC86bKKKm/mQnkaCLiCX6FBfpt2Pdeee7frUdD1BHpZaYPxenwARvvlG6fF
fuOpCFpNcLoo7npgXgsOX+TzadKUx3XgmBxRHjZPTxhcDpKAXQm2/aWJgXLByDpaUN8gZ8EeJPyy
FgZYzVhLA115DsDak6Aec6xg1VKP+0IQMtjTaqmrYz80OPemuV1Mgb9VRvyxfR44LiafyxU+aMCo
W6oAdN891haymFt4IFCSqj9zsvVEP3F4dpMSdiK530cyx2YviCXUd6TVZ2GH6IqQN7l3VuQFW4Xg
PRGQ9pJ0POc6oWvi/sz/ejCuiks5NGx4xx+G3EJDaKU7GQgE+MyRRPSYoAuNcrn2RGKUNVYukuDd
zlll3r02iUJJ3blkWRkKlZMZIIarys2kRjmATLugJJBTnA8d+Flb62zPE7CAAVB38UY11bjxzMEN
jqyuDoujorXs95qmYUOR55UxmIal/zOVFrzTSU9ZjvsEq+YnS7zrOpjEcs23/mqyBfgLXvGcfYXo
kT9epR6ntPkxNNiLMQNqgFNFDg/LLbmk4iWeFnyVenU6ytaBhdn81BhvhmmLZzdP+Xyw0kdOU3Wu
KXCTBSoGe3vM9UjzPEM6vXffAImrJeb/vVTxJbbSZzvVsCOP5yjDTwYvTXFT0EHwzTVV2A0XNwZz
o7VdZxPluhBHIwL8aH77V3H9Qi+6Wu8lJM8g16FSCXc+DV96IqwezJdmySBRgWbuqLQ7vQr4u5gh
ap4r79BqDNi1y3k3KrWvn8rQA3ab87jmA13zZ4naPX1GoXs+mGp3PjvdVx8cZs6IdPuzsXPdeuwa
AcObnLH3EDt19KtXLlbkboI2BCKqVsaePrLImLpsHm6vzZORS3c+IpY7eF5ESIIQpp1yFucgxQq0
7398//dI4DJlRyBNZYUBwre2xFTAejwOi652qc+FW061gj4I/qYjSnu8E8yVrt/8werwrCL2Uw+2
uba0lZL2NxbxhefcL/DyRCTzFWroYAunFfiKuwKLjpajiCwD3tD+3ATbcXzxSHQzV/6NF5RH7+sp
mWIbKBmwHeic117SyhtA+apsaQTD/QzvHaIQjS+UpaUBFKX4TzmFdEFPE1GhZe+tWMDVDyeidUxO
IVUG73A8j+CJlIspujttrngytTt9ng46+zybyS1dN0EpuArRt+aLJ5HQCf6T3moIAenHKPMIzECB
gEjFJ/ZvwXcbgLHgpl6QPcsnSShN9YNMJeR3mFVDykLZI4vw1tHfHBU9ofu/25xU2nugvv64Vh1F
LvulNecPrx7UROWqwzid0JLyEdlX8c2fJcB8UBYFGDJiNbUtHM5O3Wd+XTkpbJbeU8Z2WuL5Xakq
JKaIz8kY9+gymoOIq8MmXFUkAXIH1EV7Fc0jBnsUX7dBScmui/Lv0J9DVePDIa8ucbfX9+fJMCF+
R7ouyxHrlz7IUXAjNVsjZLd59HI8ssbUoCfv2zSU11TmHJLXNW4Pl4PCyNjvHyL+wyJtJmYdn04b
C8zdoCynTL8mas/DS1duDbQ5AVJKgzXMkm06RKnPQ5gA99GOObLc93oWjhwEiwbc918ZzbLN1GNI
2DCU6hcUB+HmZ4aF8h8/qGqWu9FL2OmLRyoJEMUKZXjYeAODoBKenXfZ+x/tyVEJqtb2+nHYTBV3
Sl+ofFLD0ksBqQ22+yvEzJOvLnE9F6L/9W72L49ayc1R9uKMo+bMt5WNZHBDPMTsQhNX4iL+wyZP
Gc/2H6qKra6LyUojaQBKSM+Il+bcW8WjX14p0d/WhkP1RfOex7k9jK6Vj3TNY3UKi2B0GjgwG49a
b47pN3P6ft797fhmPVNtllJAIyFxVPJ509/hwS5gxYLb2hFeukF9knIr4LQZKwyeVEQjVJ+zeqZp
8s4q3JwU+KNucWsHMGqeWPZG3tL54xgRUOphbuWzgvspyaUW/YvkUYPAx9zXaUZEomD+DDvxxAVL
wNgLB1fTJ5lkBu7fc8Xz31r5eYI5UPth9zDvQOTxBZH0hgZBstWN5sIxMTQo9o2WGpne58/FVZ7n
8L1I+/c1gYhzaoemhT54d1Su5KvfICYIsPOIeX+zTnSjjpnRjHHqSsYpIN32CVAJHQOEn0JPzZOq
CFvDNzgI0zfMzzp3vtJrEqqQwMPXthvZzC+U3MK2uejKIGv7SUQlc0tpoUipUJRrX40M8G1O9r+e
tLwDkgfrs4L91GMpCKSBDfsIFkkFovttgP4FSJ4aJmaR3tvuy6XB9O85vJsXSGEQ7Q4nBDFKVINt
yfnUf705d//qYVI6R1chQaou0mp5GBhWmd6mUylkDPP7QDYCIxHZIEMImDCkdSmgSsjd5/uwLKFC
b7QBJkdl/Tso/1PcMYNjV2NrVBIgYzDemKMLu/nXiOdMtennryCE5waShnqs72uZNpeh8qmPoT5Q
0cQ+2Ie6sFB8nfH/Q/NpQAO43FY3T182bML8dQ1P5xfK/bz8haw4XMlmVUv+spJxys6w8lC/7yhc
fn8okbYUIlgxF50LQkyAv7BMjZLQPszBLQ79oSgDOCxKkTwVPQWU9nSUT5ZnC7uP050FiJqntLia
PVpwzvKo/jRGjD/vRXNvgZg1DfNXtfYoPS891CdqEtyQ+3niMA3AvGK2eHCIZngxBMtOe3rJbTVv
Y96QMTNLX8xiHbLYKWj6SQ0XhUjFSNh7rDXiy0wsSQhWiWVbjLHYd0yJ597FT5l6AD2/YGNIaxsP
r8GBFpD0vByX30qyZLyK4yJZs9vpoq1E/c3w19CM4FS7EEXk539NcF8gAt1CZ6dqeZV58+IAZnJZ
6Psqq9pJvO33UkzX6xdL2O117907l0T295yXAIo4elrHF8ZdZx448kIKoa9cJpKEbDOZSSrzqiry
iQQ8DTj19/oxl2FSc7svY8le7ti83r5sdDBpcV6srFQzPkNwLRyXbRCG7rv5lb6fVf51fJ0hXwaE
BR9FxTSr32Bi9PneFtoLvnKVhdgmmQWJ8OBOAkHgbn4iba3z5aP4xZHlL9eGNwD9Z2z2LaY1Xbne
NJSMF0NbZCmmJpes5CGzWONk/c0ZYbZgPcGQHZUCNtZWORicuHZqqiz/R0rO9BSoCjYPUt6Wj8zh
QByQLjKYkvJslkf4kQ0wNvYUdvls86ZER4OQEpMAz88XMlgP5BU8JbvB/IMyOALJ6mvvwyRQsHD7
ZZPEbRlEgK/GFZ5ZLTrzoxJMEeyQiOiQtR2kmlk98G+jMNS+9xtBmFC2Y2rSefB6CyliO0SqtFog
UVQFGSTDL14ZwZCkavnkiD1/72VbdjCPTfxX6muQQrjC5aMdzmhFdQl7wwvhSvzcEMjvVNlvH22w
eXElT+mfXeRXzyJc4ihSThx3zbWQag5Zm/5VcXUxKtiDCUqQfl6l7hNSvd+lRLlDMaTn6+NmtNhN
ACaz9XCsCCn7nr2kRywmQ81OoIonVcbIsnOjRjky8DhChH0hew2Qr6MRrhQKkLrMxfpRIf/B/ASX
lmu3OmOdTpN2/1dyAwQTt7JAist31GqymeQI26U2m3AsRuvs3ofa50k+PetZAIltxcjgz9OSVh9Z
WrJHSVfPNbtHH3qSeP2K96sDvLIXIWAdyofB1Xb73xoptGPBFTYA9dUQgicPDd4L4thvx1k4ISeq
510jFKk6hQ2qKKkNjd7Wl114wcG2dTR2d3HpYkZq8W8m+Y2p7UZRaDvX9yjjqiCebrpoh61eB1Gt
Co9g6XD6SDrP/VRnkjBtemkTMzrHQiSz6UeH84iCm/o9IAqsvoN2HMnDiiZlpWgw/snt3kbb2UoP
K151Zd6XruXF9P9ZaX6jxB5qFmCQbzN8CIEjOV62T0+hjL+KpC2hS5AEphgO7AHcAHRZPXTPt+rB
8rsU+awwRXTQz64pl4+sx0xXFSpkBzJq6XImAGMZQQXVsf88ZoO4SujSeI9jzYzOy+vgdVUDTgqT
1xOqNcTONSdIUHwCXQnHQ8KXE5avnag2VOb8RutahI6KUzZU9OcYRG2wNUxGO0FpCLKJ1qm9ZuM1
MB3XlRbkN24c0i+bG7kXzRjS4NeC3BH3Kgwx/ijc8AfdGwSOqAUaPuJ9pUg2VhyJgEHW9q+wfkqy
MQlccij5hYxDArFGiMZ+TuZ1DRbXGSwhB4gm7Bqu3zuso0k1EKaPXv6/CarcCYZAERZGgjeXvkpQ
UDaWjpPTK1W6b2SaplgP8sM6oe6z0FPt9O/H18Ou/TcMsZkbXyoW0QxAVanJGR9v3n4HbzwjHSJ3
gNdtMc6DQwcOorkYdoNa0flxs/Mx26mU/AB215b3n7eN1yASLOf/+EItGEf2WtPf+JsNogeb9WYf
Ws7d7WuiW/a+7VY4rS3mToPZx6NvrrVpbUycVZPqYuXx46te/jrYPqb6JBFV8lGqsTq/c9nq/pGP
zTAiGNT91IuFZxNl/FDXIV3O+LpAPTCuz55BH/5B0r5WS9sWYBqtVlThnJAPOU1mBVk9CFKDivY2
3GQ6iKDzDmGOUJ2j0Ythb9/m4dr4mXynRAk/kKU0O7iCy/8D4ADFitxqEznR3627jijWAntX8J4m
T8HO9Dj8QM4M1sxA5T9qlGsST6aqXY7jDG8ecN4lbc2yYOFCSupb1V95m68dwa6DTke3QbzR2gZg
X/VrifUCLva9i2swR2j7XwmPvm2LqLUS+kl0MQ7W/69eHDfW9IUDGiemJdEDEcsvZUWqmq05iD1h
GAH7CeGPYr0sE78aw5R14bXUPqD4IFB4fRVZ2GihJWPgNbwVzElxRZHUtMU778HDDxzvzCxFZ2iN
luh8ztYxm4ChBLrM9gUsRoXfrhYCyq0lymypNwekEQbQ/ANu+rgwGJg8MiRI+r54fMvhYVhIjS+b
P9bpj1nfcF6fswZaMDSc7K/L0WIzI/sryWdqjtJvYHZTRyB2b6qBHIXZsy5nThs5xLCVhtosib/b
VlQPpGg2Zn2ivsGoDNiD5RL90tvx8Ib6ublhIROX2fn2fPoj0ZakIDSPtV5DZlmx0sxTbGJJKaHW
GRmrBrHrMG+k9qUhC3UHOLmZ405iP87NH8IOD2XGLIcXMWI/w4LFukVdEkCgvoosEYueOuFgtr53
Zmy4tac7nC5l2uHF/fISd/6JK6L9t9LmsNf18xNoGe2sKVQ2fDtQOrDOIZYXl+HJV8XFFO75Q5KN
KuV9oTp0q89mQsGYuYMM6ABGw0ZkJGLobTZ7rQgL19fU9SIoQgXO6hxTUTMc9PwfWkHslWxmXRF6
jX86mGh+cIQwPfEgPy2Q42CuQ0dnUYs6rJ1NqkLZmRsUcVTb40bnljuVkJxL4iYmWmV67mVjgJ9E
i3E4P+UZl/qpR0uSVYmD257li3BwnBZKGXeMIH/scSz44rrcn+3jm3ucDLwlOGMRcHUk8NrJDY6P
U5TPW40HNYMVkqG1ngTjtaApn+2GQirayj/chArLcREEl05CKUs4JZRVvoOrdF0zffN2gnK6rMab
co380y8WQPQ2AVyYUyVZvVGjmpUy0HYf0V0dEBLFkwfF+5hyVdd/XmfDAsJhMyEsB5csCXZL3lnk
/27YlXxfCu+FACMYEWj07CR6BDp0xfj6kDoJQeug0vm3BBzBJ38eMLzIGzw6i6lpwjVRNrVmf7yx
t4rH2TqiTD1rBLMO/eZNqIwB87Zv2v5LbPVjTfafMldTHOzseyVly7g/fghnYfOJEqyy57Fh1W88
IscTy6muRjgAd9ipisTjBchuMji1RXImQplSooo9Ub4kSu3G5rW/94ZjneeTpBM9kLkIF6eoX3pz
d8yMVp2pec3HLQ131Os6w1zlYexKOB6JGlzUV0gmdRqix4Bc+5ixchOcFZEk9PXxiWnUHascmaTX
v/eJQsn/Sv8Ep9ZjzRRNt9sPXognA9YZaUbU4Ok7XcfZKWvlWAjXStFJCkrIKmxoFlZHl2yQXxoK
z0gvOHAHZCFxK0i2P9Hxq6AuJx9YGJG27hfBXhCjxmvrJzWEehoX5u8gX7LHRHxWXZNl70Dx7Dj2
LBASPDRSmV4u6GsFfXRANIuChkKslbD7ox2HFStGfmqfc28NjhEC4VueNlBt/ybcqds3Udb7nnaU
aqLBnfe/KnIPoIykKVQgnXijyiiTtffx+nzV4hNQZh0IzSUcz5oFjI8RUlA+f5fU2dPMQ/TdzMm9
JHHpqUKTieJUe71KHSd8qKNj1lepsrmVWceNGGRFtfLMCB+6z44XaMuz3rqt7an/YhlmILyZ3/RK
jYGg9/L2DDv9/bjfPEvT+/GQgWIv5KQNfJMDFxjiFQH8X2+Tx+FJEP/ihO0BW8+QSGlPnCGtSHv2
uuyMnjuZ+25Eyhrr0syQl0kvCJL4+xlwyx5F/hTR9jvvJunDn7TgG1xmGl0ADr9EdtXeywdEt8Bv
q9jkx+MUmclc8ERH157CPQM54kyl38d8wQh/l9o0xe5DBvLl0xT74vndF6u2FcU/Ubukh7hr9o/G
404DXHtOhDZz2qPkJuSibck+DqtfeVPIwzp6z5QSrY2fC5W2NePqaLe7a6IhIpCI5WS2eLS9rsPH
POyW2BQa+VN8p5sJ33dfLCc8ZxQQe20ivsPxPukmTEIO86/7Xy2nvmhrv1DP/PZ+yDa2Q2WlRU4w
gPW3GNIYNd/rAX6UdSg5FzmF1/e0Mri5X9Ga/P6GzJsk8G01jXy2Bzq4v4ynDmSH7Bq4mIJX3wvZ
aDTpSjXHMUHkAggySUeUXXglt4MGMRsX94a59QsYx14wEqGDTD4rGgCApQPCHUF+e7mvdSggCRrW
pTzjj6/vRtUuKmVIokDGMIaFfu20yEF4XgcpA898fzVimoQBzTIHgwyed3x421LpUtpha8FWGb89
jloh9350C+I7/L8H78KDEx7kJJsRaOomSJ977hEJJbd/0Sl46szORnPakYoR2QyRcCscIUV2hujS
9gdkJ13aGfiQAiuZD4Zt2F+ZgBdOAekO54y35p5vY5NYlhk52yBsC9VbpIhM8Vg2lYAY7jygSbN7
vgy0rKsSGcJyV3D3ovw5WVb5hR7JF4sAVbm37ko7nwjH0rC3O9ktapoB7tgiAQv4/+p5abYnALYx
4HFCnQRVlF59GQsedcV0gnHRxn38aVo5QFuIWkSxVpaj8gkM5VDKiqntCbGhtCQsTNiGmePoMZDA
NfaUyJxMq7UfPgVV6u2gkaGTJ0+QtER7sRh8WWb10q8sZt7DE14w5H1dHyF20fkgKhPxf0x0/XmE
AR3JR0fZ8+SUFFUFo8focoYgjdiDDKKyhyRt3OYJANQGR8keVLxhilSXapwc/A97jg8Uj/ySHwO7
0OJ4FtB+TLA+TOb8G6ZF/WU4NaGzND8qhmSkvd5ImXruIb9dDvW1h6bSl4G/9KeJ+ea3moC5UmmR
rgqzUEdjokGSjRUVGImu2B2DYfGpPaoBPpXY/6FmSuA5W60mhrO0diythZGag3GvVVMNovCpyvow
r9iswtNO7SGFSNN48b75dD9c+TuIZumIvzpHbL6f8NaZCgbKBz0cPlL1IRcOtnJkGp6I/50W78lY
wRrOrynyYzAGkc9UMhKAYuN7yjgi66dhXvVIxOMuqFrA1qlQcLD5VExTldZ2oqTxTyrd04odHe5Z
zvTctGfJzhNVxRusSj4AF7nv5nWHnCQDpI/7lnoXdCYlHkM5yYChzMiLdgZyCFZnCItQCIpWVyM1
IY9ByS3SJlrs+MEdborj9TRaZCBiR2dTkmGtzMQMyyjocUZY2KchfYMqQW20SHqjlBqqb57zLb+L
RVlPSx/AC5/8Ni+uaXqW9Umc5lviuaxi1rd5yalJStDHXw4TQKkMvirb/WDhWnJ+gJvdb4z121yE
U3tmYCgPCVE2UKkYEo5+RoVhuqcsJKrn/+6s8jlxXDS9LM6+yoUCZMUawxaTv2ztU3OYR1rlodSw
0cvCYuk6HENVvnxjfOFWBJsmNYE2d+k2FHCWC+5fGFIjxIRcaQfaX/2hUxFOIpLCU44fKyF0b0UQ
RFf2gVcXVnhAqS2c3gyJkMf2VGGVFdSBO28hYU1+jsM45a2S+ACMyJAY1uoGr3weY3vzi3cneTOz
kOzXIX3oY0q+ZfjWSXgYkB2O5X4HOkYqCkEmb7NEeEOvETJWmzKllBiqfCUCTYHQH6bakmkCmuQQ
s1zawYuKgkcmc2P8iRoIvgOmD8D7R4a+5LrEQWzhSH5ePV1npdJhw3SuVmRSWTOE8s4LOgu4eaap
Fjf6nQEZdeLSSba3b2H1uWYchN/EWHw4MDh5ZhOytTTnemhMkyKhno9MvqAQfzgFx/6GfWjFv5AQ
P6mWthQtylLd2pVejh8h+eGAQFg7a72daINUMtAa47uVx7R3fWiMTNDwrZB4Cdyj2yOTctXuGQSj
I20P7Vw2IsJHJra4CHrJ1h7xtttbDl+pjRF/0LAQuOLKu0eUpEXMg3uP2ybTPJ5o+s7isXSBvzhX
agbjv5EK9ZEQ0Wmifdd6X0ubmiHBdOxWsZ9npSeT5a3TS64neCIYEufZmg/H60rsNnD5xmXEsZuH
k64MlCTNeO3mBSV3kHgtn7zmJLHKMQR3LskGUaKeTKLcNFALXjb/5EhMi8sR0QUBUJdYn/MOU6zr
gQgI1VdxJ+9FsJANoDk396vTcm+guaVPtD5mns49OkcImE68IZxEkqast6MyYldZD/9+Ep08tY2T
YhW9R2pprP7k+O0Th4SLL2Zg3xKD/sDQDaOFMVovMROpe07IIR6D2u8tNNLkc3S1B786/Ri4n08y
QA6GIl09L0QAQg6etyHOehT0ZjotuDKo1HiouCxxDP8d/5cOVsIE3YZuaeKA21JM6A18LJvK5T0o
iEPIbZsMkNM9AbPdRxBb6l3UfBDejoh1G5qphBEXAQuTtJhV0crGuWc9ocXhHV3rxfGXn43ALeVq
3AQjXMoUY9m+vWNDjBcnfrsj8/YBSw08z5q+BTPQ7Gqpo3Vwyey1qSLXkuRP05erB8l8wJz2d00M
QE0/ED0Ijea155Lu/DNCW+n6SHa+hdbfsb56IsyAyLo6MCWEENaajx2vYlpy7D7vk+iYk0n9KYUL
Gqh6Rpwdxf9ekIcyq0MiOxnnR0GSxU3MNOYy5vA+/G+D63nZE1C1bqIIOPo84YwVhiLWPXcE2HDU
L0P6gCkSNMR4FfvN/5yt1iyPVe2BBmnZSIpvka362sLykK3ibWX2xd1vtjC3W51z2+fuqJe1H9Od
aI0tMdeGwWnS6GP+UuiwB6ylBTHnsT23bUnkB7um2Sgrk1zbX+hz6xymxYWyWNsIEJ+Ep2C50grE
4wHRdmp/Zgr/R5qgmrDGf6fKA0MHqacoUOXj1JrYL1uVCbXGufaBmEW2lCc01/wTA+e64TmbVTLz
Q+Crag0ahHz9V3PFIdQYZoR+2m1uAwhAzBGctJaepc4Dh0I9mZfKFnNZH/j87HRHX1p3rcfL4ISo
PsE+zDCT9LftMRkjLwBwP7QXvnG1gjWCIKF5SLURPPnUjvcd4peIuL8Nd47ZtwOH2KoUqITUb3uV
IPBEBUxK3LUHWmUvIcxnO/jTnjArClCrQMeRVppM+HRBLTic/+V+LdZiNV/+3+M2VTAi8FMqsASs
J666LVQy6KbiG0VkRTUmd2mRrzNGA0Uxs+8JLXqX/pPYUlmMHtCePpm3FYLTgxf2BYc4hQshV7rX
8d5feIXw1iyVCxvs/wkXA2Xqv3knHWjISVrdfLLKXcIQoWqh6XrTqwZ/rolJqodycaKzQUo3zLkK
OmKcagRpNX8QURprRk6OKjxPubhKWE5zi5sEcpn+GZukPtdUyLiRxM7viH5t2eU7Vj9f2/IEC30x
wRu+D3DQgyhug89Zo3UPZQ8bQEaNXUNQ698mXQr3kyarWTTaaReaOdUtIQaxlgEM/rvIlyvZQdzT
kZMa6oaatDqMftVRKP3/XrtLv7oUosTT/VS+/sjQxR9GjWtdvujYW9e+Pc+Hi7f8kKglSCrJrr2c
zQlKIVxjr2UuwpG77lDffrARB5w2G/nbuC3yZZD6yLnn3OyFSWmIbzH+5kLEHwl6fsWf113n6PRK
vEAbVOZ5W4z5YUyYyXE9d9aK3sy/jYGsosLYPDAZtjLq02Nv/2lk6FNMYu4MjOTUTffpZCswAkwS
FfkxgrQ3KYIgYuNoSKcblQ/ooMmFRygvQ/3uzmU9t70mA/qT+9hG3hGVM1+Fn5dUuiBQDwAmbsxz
uWBbnPgDdobvssptaVl0Xhip03PDG47E6vGp2VBW4U+05boeRNR3RDQjX9+DgFqNWLB6Rf3ld7sQ
puD9XPryzLwgFFzF6nqgDAh9Esbn9wYBkEqIzJy+vivB0P4nZX/JeWkTJ4HoGJRw34tjfW4+GCs4
mweg3TI1lhyzqjIrDzCYTOOZM6eIi+qHttWBbRhg0VBxFl3cuUB7WB47tYPJDXf7t3JxwvLBN7fm
qW6+v3gOeCwfFO8xvNdGwE0Eh449zq5KfuV7KOoN9EHFVwoadpN5g1zN477q0z66dgqy7ETJZAGz
hmuBM/mwrGxURsOO1h6sWW/JJhpvpA4ooBKDJ7RxdoFk2SUAcjQLKlZT5+TngGPuHX4Mo6sitJh/
ATdscKatvAahT/yQLCN7OFvNbtwZMo4eyAFiinbnjtnYXFCfGRhokCtfo+oK+6t6nF+omiz8KvXx
HHhyGDdo23GmQ0oVOMSCmKQtwofTYV66EMWeU1szr4vwNidKPqmlzUbL5os5O9kZ29WlZ1QwtT1v
2aSQ5UJJqmneqtbO+Gpic2E4l1O4GlfUnv287C6AUK8Cq1kXx2IAd3QJg5QxadzE+t5c33VgeH5G
fmmklloQ8f+7twbQQQuRyiKG4EgZ1S62wSyDBt4CqisOioyUCuaaoGdvZSLIddRqDANvnH7v5tk3
LABkwFcjkh7XWXc2xJzW2kVrFtgy6PwHYfoc2+U1Y8P14IV9KrgbtkngARr3wus0vriGbpD5XFqz
nOEMSxkCe84mZJ0OU16VoP1sZPz93tHTvvQZXtN0K5fJ5S8d+6AymdKJQ2JFKNASVY+Hfvf5LGiH
G9fVUOrrq2yYOdXj8XTLMGU0RQopKSJMadd9iYVBXr+tjKzrGOmRFyeHQsZK6qMR6fNtRVe/XnJv
hk2ES+2UVmdyieTcLpBVT1Av9Xvyb26G1rXdX3w/MxTGMRuX2Xqz3e1ifOGgR8PydjYnuQeFxdoh
t2F38+a5TzsPVfSh6e8rwLIi06vYCfiOK9AoV1It59bxEwhEYENjWstO6Mn7wnE1Q52SfXQcMZql
L3Z4H1L2T5G434qoQqyFvzf0gVj1mXUo50EGKGHOzAj6rGg5pJA6hDjLBx3sjuiTk4XsNW28nQzc
ndzkVnT26LeANXAIpNX03oT526/fDV3DpAUINNuwY0Q7mX0sAUzEsa9A7ARM3eo3VZ0HTbjwJSJ7
QegsmQ0fc1gbFyCiJMksGpmi5+tuEmrlDgv7czh0TGaZq84Z4kRAzR/Oxaapsuw9NmAFtLjdMSC5
DngwQOEO5UInvTpTCEj2ekE3O5feZjDl4ZYYb2pQ+aPVyIIt0VNJ8o8rH3zVIYeD/2GUBlGKsLyS
WNY3gjZdCDSHKMXoLv0pnYKzAEa8Q0XBj43Tl23aJlMOKye44fQMNwcx67UAx5MntWVHMCzn7/hy
Y3jLxQdgWgUNfUwmjIJpcKhu+9q7O1sJvMaz/LCdcPpsi3O5JiN0uPJsBnl5tHTG6qNX1TLVNryH
6DZidvDXn8m7r8IE3Y1elqGFD1pbz9gPiWSDRrLWyopHAATcq6gGeoPHod0XnstH4nlaOU57/VFQ
NUErGFA2PBoYzmwrMV/u888hHQDBRpaguOkO0u2XCBkbfdTYtosbcJxatd3HJG0OkH/wm5ojcZe2
B40wnM27/SZUk9Ku9tsJ83LjHDyye0DNJxqs9GglHcnBF4VkVjWLIZRtdWcJW74UILIv85VdX242
njYkwnR5Rj/JTwwvaKMEvcPRbAMi2f6tyIV5ER770wjfVMO29k0xqBBmmXHswdVWCMlINfKkc2u+
72YMvbZQXeiiVGCXu3lpvdb5GqiOpJ9DYDua4lsoN1xQaCMgitO5pbeCgx5kn8WUUSsOkvWsmuU5
amRihkZZP4bWtaI68Eg8Bz/DM6rA9B0CAQXLYI39pV7amg1BK30FrjBRv3JxjtsrG3wq/Hm3fQMu
Ylfm0p7GVKI4aXrRPVibURgh3jT7AG5Th6zlKOHzNx5o9HQ2HX+PBRNK2B2+kz5gu0XmSCEgKMue
gRZvVMCMdJJUHkOyb2oHBa+ELCYqOfG/8Tiq51BImcTZkFN8f8hZtUM9QrZH9BzD5ViRq/ac0t/R
xU41Yy0QJvGweMeYUQJHkUpPxunBKudlT2BC2icjtKTDRJ1VY25gALPLpDlAc4CwehBUzrVLPZmO
//5D6bE3W2gI473V0YZtjCv8GAF0sa1SeTP3OJZQWtHoaBOvlLqCYOFqDSAmtjXlroryCtUT6EW8
kFVbhl0Uhs4Y9Mxe5ggRuWdxhxjKx5jLrp6S62QcV7m8CbmNKbf4FPze4D50O4oxxXGsRBeJXPvC
CCpqAdFQIF5DcrCXdmbp2zjMwNDmQ3F7vVl0HRjz9DnujWUsdOZOjy2hUNB93MMyDINClPeQlu7w
RIbh9C2Wpng7IQpyF46kfxXtLxWd6h9onFVbSEF+FD5zLYzYurXN4H5LJN8TZUP/MhmbJzzhpU+s
yuad+qlnwmPdl+m5yM2fMNdkNG5VMem/C2bst+4vpFrs6GCY55yQmCOjR6uNd9bQdK6LDpuyIJjG
qL4x4cgRNI/Muqj2LdSEXAnkwPInvCQSkVRRhrsZtKOjKLNNH4tBeSToBJ+Z/u4DJdRDMRGbOwnV
dwVfsyHvjDDacUU64LJi/txbm6yefD7knRIzVvNapIGoiyG4lzhK57QcjkaK2TTj+Cnpq27r5x8Y
X3NsbLQx7ABNAe4WFV7w16wPTqpFj36/0uKoPrMmtAwZ+FuetPuvBGPXC50AlPqicX+x3KVhFAvq
RU0f03P3wpZavahOwgYDc97/kzDShnu58jW2XqwzjHvwdVUUSjioFPMLq7De9u9ODiN69oKyimS8
YNxTye6AhlLHp+fHClEJsHc8Iva2wsX0F9Swzo8x35FZPSnHzJ2WxGDsQWCHy/pMwIFJT/yRfE5k
ovePuDKCE8DZHsrd/TIQ4piJkCLOqxbn/H0ORNAz0YwMDzwX/QrNOlrMibmwh/t41vt8rSy4ln+n
5DajgbVGxbAHxAkWqjlboxRpErNa1fxpDTe8xOI01rVai8+WUAQHRMFa/6aKHBbyYW81s35YmN9r
tMEdFXPXfaEAfxsNEN7KfM4Gv5jOWclVHFbJ042frsyOVRwuuphipjUfykD3m4SLyruzBM6215Dy
hNBu0jFW1s/QcU9tNuBLS7avJUa253iyhCxjcuDWZAMyxqAvqpnx2viBcwRI4D99iX0QjolWcSpe
oL+Z1YkpFSEHzuCKOi/v6nc5TcNUK9Pb/wSsjJANZXOOliQ8kJOZ7bCXqmOk0efUip5GO8eL54k5
9Ra0UQJM63bKrVixS0U3Y+oOxSrXlLssHBX7AcxT2h9y5PJgbNiO4saVjlnhA1CzMJrxvpxSvNpl
Vk9XGOG8t1NF1oe6tX07yqOYT6bSKp26fy/6RnYubpgZ70MlxKZsrMItW5PLLCkM7YZ3+KpY9587
nVZaocT0jkkZaE2U7zDkwhhJWa0nfMSexuAiFggUamGsuhmat9hFTii/B6wh05+BuwTR06sy7WYY
oXX+TYILmdxxxdO/G/Mm/J5nHWqR8hsn4xljApdofUGI9Z9TIf1sGnmoEY7mzKdjqOLjAvhPZ22R
FHomOZxbNyyONIc0Caw11DME2BaQ7uRmgdgKtvAvJ2fZI7b+EEcvQlVtYCUG4tE258qnDhOoL9GY
ysxD+qtwxuf1XOQdSfDzZVyj4fBES6h68PwoZ2ZgYgE13y0rqiEeaIB0heo/CqraxD+WphYc2I/d
7mE15BMQ/e9Zos1FcR493LO4xZPTVSItBbm0RPhgOv0A92bonEybkulnT1M38io/JXddcLzZvAcx
SAD5/lwkEFhtyBuRhK88JDVByc5XVulJUqm0JHEvsTGcUDv07P/I0JNcwW/ztqlz8/4KS5witF2z
XImIVXdi3nhFpTnQ2p5MWf5BXBojVrUlpjYT+wUQtv+PDHBZuAwh1yOwUX4P/TUYTRDExolrIYx9
H/crlJYKFDqeSYHxrKI15TPcUj18SSmd0G1VJXSdrcEPVfqLyQtWkyFJNQnPveomziTeTKlrSUu9
/ABZDozNW42drCPTi18L0PZM7G4z3aj7nYXo/OJ6uqxzTQTHhw8LA/LZ9PzMiX5AQUEb8o7AViK8
utHSey8xTVr5gS+QTQFaPMNkevof9eZpvWhS0koWM0jAd8P0wTtVPtHwsj5/+bdZhIYW0BXZX5wE
pgx8sRALaXvDP9TYsygCJv1ZVhAKucqIb4mn65qapDkE+3U9MWJvuabveqI3C/yD3e1H5v1I4Hun
TIPF4LWXVlUlIP4xsqvZlRiH8tUbGr2BeUrm267P6H1W9sWO3ufdwR7Zv3/D7Of4mPQ3fqsEp80I
YxhXyPm92uxjIrUOxqAcnRQnHMD9VY2K+6ETjyPrTpe8PJQMXLPRBVD7GVcVwH1m/O+hr1JPPPs3
EQWeaw4RRiPTi83pglBbxemb3P01RL7CtfEuEnAge86tRAGI1G4znYNc8s3FxCclmqKAoXz86djA
lnnsDGX5fFV6H8NNS6+1AmI/sBPyqm+OVbV6NZWCvYGmcpsyElWM7xol4r0I82bjJmEl1PcV/7P1
lHOcKgXtxX57JPF7bD3UrzFdo9He9LEokfriWKi4302lKnz/hfU/KEa5hdIyT3b3Nh2UXB2fGVlp
8kPXW3quwJI4zApQyFd+TmcjOTgs/gcPoG/eDPqgcdZXiAvI7R/yAznhHL74IYgVSTCtH276mY/V
BIi1gKTnzWZ2NDdzrcxbDcjbjbDaBItUBVgvQu+yTuLD7SVhV5ZlWPK3HohxWTQSdvGovs9d/QRN
SShiJKTU4SYs9oXmlLg0zclQkJvvHY/kPlUaX4mVparDvTu7yo8mJQydDD8Y8KYqDiCw+m4FzRt5
11r4RNvD4MDpFEJ9NplEKhwr+NPYuJt1TgXAIWRCji96kj6LyEPTJ49XCBl/wsoxqmJ0vtU5jpYn
P2SU6W1fiUoZ2C9W1OUAVfw2Xu/pirCE3epl+V2OdeIsM+EiUx9km+puagj/oFuWeWrNagXnQ1Ub
1ibmXWbZYJifAHCklo4dDWsP4m76r8Pk5XYQ8JVgr9FTbkVAzEoiOtDw5rwYD3KWgk2Z+AdeFtsr
qHSkyLZrHSsVAU1yVATkdDYxEiuUNwOfM0eLFBXzMtqe9azcQuoR0am0xQFbcxVL3Kn2wo/eOIzL
xu3UrYD9JL+Y8z9R/AvyqkXMGHhhoMNUSPL9KRUfD61V8sBO0o2f7iZVQWH5A7k4Mg/ladVqZwLT
cnz/f3OBbapFY6oWM3+HlR1t7R2ND6qZ9WEFU1FHoXz8yNXcOyQCPAZjkeh0HEpQqCxk/NXbboGD
qr63XmD9vfmLYo1xvjOr4/cRXfP2bdsVxy6k5vjchG5fgkABUkkt8JFhsLzn/f8mXdBWi7vhVqZw
jXOEITqKRvLhH9gD2is+ii4ah4cIj1hvdBCIXEAG2UCsEQGl+a6+YgOI+drJVexAeYpWyv6S1fXX
317PZd3WTAP+N4/L8hrT5SPvNobBy6UxJdg4GF/mOoKmWZRcYYXVQaTX1/hROLEGxEXaCxvGvfpV
WOu/VM3T6SAzUBjks0sLWBRfMRdzWlWXod9WENbJqQjAcGzojxG2apz4r3zVvA8zU56Y6Sh9HhUh
2asPhcY10YrW+zdqybBsYpsVF+6tpmDkA/zNdQKQVAUiERkVY8lGaghyasYEebxCKIcJey1QN7A6
RplkTw1RZmVWNVFUIM0pHvG5z/NcuoMlh9im2ceteApkuqzYWiBvz9osD0iQuD+VfZ4LGVVvN+1A
HrmWdBLd3jBAEAlp8oenDo/Ck56VHtRP2ZFc9gzSqVCMZGBL12xuLNjEqxAUNybIEwQQVg3Gl2q0
M0NVlHHTuMooxG5BtkvoiwfEVe0QwHwgRuiAGkmGrqszhbnomZWnzlaIyoq5fiByfvUfZ5RiqRSc
0qQitjuE/Jqzhw/8zpLSfEKtGx0xpAEeReo8Lh0ZFTBej/5HVsOEFuuH/HUHDPz5VSm1rx0aYs7V
KJE9P3W09CObx9YERypsURalrztOLbT0suTDL689+MJxh24eh6RNGEYO0Skyeh3En7FZuZtIYpgn
5XDhi1KcAwl6d/73q3z6BwB+7B+v0TmENSmZ0XGIBQ==
`protect end_protected
