`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
huhkCp1xAa19GTD/MrQ7700+xBmcHqKyTDC43CnERbyBfXNAzAU9CUqfNPDxhJFOirIWv0yQz8fY
cpC2z2ueew==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
K0Vb7HEDNytHh1AcmV0XqdBEo1myp0RAQCKEngK4UJEJ74z/2Wob0uh0z0K/+fxYCvEzodPxdjX4
C20ARTbXqXdEsRyxMb0WazQCOYKyx9sfganvQESYcC3awPPMaSSxGj6hMhx7KiWA2bJ0WVgoFeay
u1HXBKRu1vbxXEMHXbY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
K0ijBIM2uPO9l3rfd7jb7Ich9JFhv7WRcXZiw8JlAsDWRmKO7v7kdQEmDZiNnbQig8n4mYZKS+3D
mliSQA846aZ2THNkvMWn/K1TeT3tNuOkaF+0SmWdEQ9CTT7gnfL9x7C9RuvvERDmCeohU0zC9Ncn
H0QF+lgho/0+cA/sR3rLvuBS9MREgRtLLhXRzh4dvnIpeSMQt/HwiFVzYkwC2dm3RrU3FQn6QhxC
zlVTJSaCNOp0QRA0nWcJmQKzXx57exuuJIV4JiE/qV0tAq14toF2+kyMhh5WZv2wDTC5qhjwZgTI
pzBtgTnpiE22bERTHruJ+/YjIRoz2zgz7SIHgw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
1zCXIUP2czn5r2yOSzCiY5mHzR1PDiAtrLqvoLZf/Ssy+3CH1wUf2tME7aGhZ065dKcui4jteByZ
GCoYfDV/l9VwJr6EyQ1F9Hvi2iLet5Ieo9Pw/vMNkNL8X2w/ikVkmAKdNfAHJA+U4hgo+Y3uQkp3
gx+JZOBuAqk1yLwVppQ=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mTbfMzkG+sfin88PoH2kYiZi0JQ7pPZ/DI5s6isAMevnLfCePc92Fsof6SEGLTfTvVp7A1uXRwHi
vMMF0Ks/aAM+QOdFwl4qm7+sVTrE7UAAMP2BnuV859OYPNRRsWpQ5iDm3YSRBh224I0vN5QnyS/A
pPA+zGiRXMIiYiTezUgSfPtbBzz/zpOcVNsomEvkDQzWwT1I5TL/5QGRRdr1/nK8DHNt0e4IAfJL
wPjnBnMedy0cbzNKNkelckGmLvKKRUJMr+slajjssXXtRtiKqD/2CMGgrzBMEIAGI8mxRn1IqtYB
V3HR+3I9oMeIVzlBQwnJ9tIH/CK20+/MTNUegA==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
PLuU6qjTDiPB6Cs7c0HqWqtCN4uO3BI0ZvmET/bLOpJGPbVwRPb4YiMW6X5dthC2TMnTaeZ7NCyg
vYORdyZmpsmS3pI4XF4IH9gkbZ4dqyhad89nDr2Ubt5do7C9dKeHW9UyZUC/0Js5XQBIKxAU43x/
OTfXGaYe5afmhsL/UATZtaujZ4ORCV8r1aEsSWqmV6ZvK/Z5sE73XevWFLcpADLBRpJwBuWXhr5v
KpobX/Nnr1ntsAiwu0xjB21Gn2mXLuQkKD3YD2vwv30r2IlEVOxN1QiGxMvNP2+YPMI9QZfqLVmR
aPtg5yHTMZ2Jn4G0fPyXFN69e3lvfzwdGhPvqw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4960)
`protect data_block
FdiBo3TnN0Bt9Hkm5Zy9uJDnGOzevT96BnjE0bwVotWoyRdLA5W319Zwhsv6axrcsNcViddwIKp1
fawYnNpz8YZZK5qOAC0Q6yhTFGYdLQXbKxM9o/wDwXqnp6F1IMhWxjZW4EVXyBpMqLa8hamfQr9y
mcyJRilPp6+li82Z+ZaHPsVaMugH+ZM4eqgeX2MXERHOg/wPhUQ6o4NmaD94c9ts7cmzl/K7b91W
PRZ8qGbvH1T7z5yV18m29KtsyVDKLzssV92e/BEluTfC09Q24oo3X2iDUoW00kYOTF0+A1yDiMyD
pBZ8Gr4P/8OkJbKD1gNKGQMhlKoZvLZx09oX+C/Sh0dr0SvTBoBogkCI/Z10Jk6ol+p9AghdfEE1
Tr8WilWoE2UNDuLjOMB8blehjluD/X9r8bgllo+9guwmrY/7NISOaOqKNwyvCDpXgTViZbb3LuP3
mscNkEjWTWfQTad9jvmU+33XuJ3vttbR5zzIGvjgYfN9uB3GMfJq66O9BDOeS7QMYVGsh4HEdDXH
3fKTgHdABwXv+h9AxI16TBYPI6C3PJmLQR+ABzpddt1l0LTkNS6XPHv85fdmhjJyP03l0pfcqO5j
mb9lpLOTfrghhzSfuwxyhxWCT4KsPafpo4zBkNcNMxn0rU+qEOSyUF7GMCD3dB24fIY0FrCLLFtk
cFVH65zclKs8JVT0g/t0c8snP9931NVcFfDfWv1YC5htpRtkm1GEq6AJ1nhELcpfNhoMLX8NK1oJ
XHKJjckhdpAYgH8sFKm3Ch91KQ7orNXJv7MzBwSGmV8mF2OsR0k86ntncs2R0uv4z6hnQrSR/Ja6
IqS0UV/j0hVWdvMiPxnZIyCnkfDv5rEVLKxpZ2YM4hZDq/6AWjCon669bLbI0GzoXcwhOe5WaU4X
0oU5PvJKT5b2Da2w+sAWSw7I3GQ/xBO13/JDgeY7o7+GOBSRaIADHFHvIS0FkASjoywH3iZYehht
qhbyl4BLajaJpyojJbSXVrUe/mQJQcn6X/X5xPIma7eVbvD905FhQ55+4TxaFNu/qmV/MapzZeJt
vHCH8dcsd5d4eQuNWiQDl4zgE7jcMiJ6fIEmzV3PBIhVe/TCbZOBMah+Kl+nYFdfROt5c9wDlLVn
e7ih6l9R8YWLWBWXliEZ8PICOklsOYyGOL2hts1kJdFIJ1OrFiWHfwMiOcuFVszSRBS2XI1Xzb5o
pmF5Fp8F5w/rVXBfOu03p0Gps+mC5b5l+Pq0ubnTbepSLTBdP4gVKwKFpdyLb6WCVY5sC574EPCq
tPznkoy7q0ruPA0kkPDkocMbDdpnS8BntN+hpFsZx6q5hvPoshB9EjzV3UmBVebP3YwA2+eo1R3Q
gXMpTWEXoVh+ikDAIOm7JvghOUHMaub8rmR6twQSyMAHQMbdSWMiSAYcLVji58Tx1E+cb3kytGiN
BOeqwxEMV6LFMKkW3UMH7HyBd2EmbbPNcaOLEhN6GMsPEMi0z40YOtD4Z0gljDjlICmRawOULWPj
rtdHiNqsrdjvVLkn0twlutVd1ql9eHr3ecV5wyJWBCk7b7DASSdfnLeslK8aR/YTE6NsareYCIKl
P4W9sz5EL07ell6eGoyxgWSyzF67oFG7KzeuO4iETjV5h3fS1kTD0yNr8IYRg2ofCfPoyOQmcy/O
P5eWdzGC5id3eplfVY8ykrluOAt5RjoLaSO+G/vmXx26liNRVH1QQLhjaKuebVI5R8xW0kEu1FC5
Ydn5aUjtfCwdnxLmvsptq2/JysAEgA87p8+mB+NFFEzEblHxPLMplb82Kpu4jo822B7uMChcf8nY
PvkJRfL6d6gSGLPczuxHnTbuO3jJN7QE+MfkR5ckBGHDFaJW+IjCSwvjKvXo9dQRtocK7eXZsHKH
fBu1Tpe49SWWaSJiXY/RVyscSc42RWzEEP7chDKujZj66fKvaUmptB6sWnX8T4QlwYjX8LPFu2Gf
+zPzjV1xOcwWGzpuTBbfeUju2oAv4stfrWwhMyYM2IAqzasTNY+6DvMlEu5PFuwQZFMOE2MdQNQS
B23Z3JsVN/KJWpNHH9IoZ8nF0KvnckRyTKziO/mCic//9qjYsLr+uLzI3asl/OR2Vyr7E1Uek8sh
Zm+yJlRsxcCfSuF/OLW4jblDQ/6yj7wpkyWGv5N3s6EMcdOdWF8gZq+26QfYfhDTjyBwuFIyX881
FD9NZmQGgwpfwLyNM92PsgPOmk7wkhf3pknzfPcYABbG/l6e4CzeNPTqEmH4VMfmLOYi03A1e0A2
i0WLcfmGcTWSJZ9FMaGCKxyQP7qH7UojqrXsoKI0T+IKzPcVHIJ1vhC3vG/O36QNAx6q7C/Ohibo
Usxcz+BTp74VZzJ1zRisVvjQW4oyFnvUh4Q5WjATKRiQalXrina8kmQHSGoJOKIBZ2EmFrXLNbQ/
BxqbTpz85edAEq19pVcsEem5wp/CW2K2XHX7yjFdFZkFZiPt+AC1N1NgnZMtjIr9n+9QHgDfJmRC
GmIKYgbTh9VnWCpipT86LZqA1+FN6kRyL6cmY7+x+I5PvaTuLkWs9ZzFMGGB4lYgZ30v2QBW1k9I
6VErOHS9LOvqf2gfgdtvrCfx6rmmpbRdfnZLymTCS+AipcwJydKkSesjgAowZZaVytrS09ycLBle
I6D+b9hMq2hhMZIPs4s3APZEkr8MCyMFcxwq5r89clLNGy0tF17AMNHSzCTj6zlotIhbLODO0hDo
XvnobQyu2+0gVjaKVNC04K+49LUJ3WvA4KegdamdfbDFr9zgL/TuZWJ1esTqaFi20LkusfXCVV+e
DyCjLMNA+O/U2ORhzjWO3qcIJYHhePtsvynwKUtXqSJlKksYs4j053YN1ct1vZT9oEudCC2rGbxt
5DohYTjuxASoLVzxxjJV4EPaFzvtFswE9TjOntwdNfVUiGB/Gbv84ntDo0wLrB0NXVYHMhBwctmN
jKOCXprvh1EMfh9dOq/dYFHUFUPmAxlIdJ/RkxR+3DoqSbvDdJKjdBYeZUqzU16sZGB4HaSSAWrm
qNv9YGuuwnKP3ZUdw53TkLGlIw4gtNZpsZWxzbsyB3u5oPQzqDt/0DgJ+7C/NQN+RA8mMmOp/nrA
YwlM6c5cLr9wZfz6XjTsbYFoOFWd+hbhywg0v1D8S9AbEgV4hefC94MNQE4jln6QnuHbP3X+L4Ht
lLJsRpB0QA6Q3qYcrLrSrIr1chnCFjxQlGpKrCpVTf3rYufDd9iNpuxZSLMPWWvVaZYylicCXiaI
hPDwT+j3T6Z3k5khn/hnOTop//j0Z+xs5BABhBOjdPOEeiIJBxKqYgQ9q6z6tn6woZE545oGa0Ha
htld2mSfAoJTGtHjhYzQGjpjgX3ZqOj989OdMa6myp/2vfL3bl4+5UxeAU2Mkhkpe9LzHFEWNI/R
t5LEGcRjcw3x5dBgymML9tI0trkD62TTvVh3gY3v/ncK9bG5jc2F8kWqcnMQbl4KYAPFvdterXge
uGK6j6I8zZeIl4IfmA4BMhty6BRRu2zEG5iXORxmHN2+cLtX/m9DBPzo7RPgkCcj7QTYAXmZvEer
HjIjL6Mnzvdc4+cSU4WZu0otE/u81v5K6PuMcnej16XIil3JWUNcD5MseXyl0W7RZJSv78nqwaS4
4myKLeele9TZzKdy6/ukEp/vdmw3FQktO/q3K8fCPstQ6Q3QLb1/6bKhAmUl0vgt/LDhXrykVQ4v
oSvuK0FSo4ergi05ap5i5VAdgUfeESft1QqQobi0cg0OIvA3VnMFGjz9PmDicivI6yJ0KF5nXc7h
54rUv1VOPy5jpnd5r7hSCEVB3CZn3yPc0EEmGcnfsgQ7+J5SJ+bST+/0BSQt8UpG51Y3a2N5IOH0
wECSKKOI3W6T2mfEe7UkMuZPmF0FonUU/21mb66JxMj76lhNvGgwh/Ernq2zrVRI7Q4dELRgVX7T
oaeneDPV0cVSG8TxH5sfU2/BZH8Q9LPNC+yMpB/9ObSkTM0h7bzerWjOJC5rb/ZjdmwavnSRh1k9
vGY9raprrAC7BCEy9G97l6/2pR5ezAy1aogCaF2qMUZTxrmDrxIkusry3sGkJVY3HGCaDNNNkYju
egIxzwfCnrVAMBoKoWYvC8J7fAnMRjLFTV7gc6z8FojEG/7ZgdhPRY7Yk+6L2gFEZfXLHcpfbWtM
yKMXKHSgYT3f7r6FPs3JP4DMvZEWiqS2+27I0QnPtvRGf6wCH74P7HtW9Y8QnDRIO00TpHoNm+L0
6pKwwTO/uzoracDYEYAwr7jMRFpVFaQed2KIJb0rsa1VcBzjMPFuNuUDQHBjWFfY1RbRILuxpWai
5f/a6XxhvjnVbcaLi3uygRVP/OgKHXi8wPTmrttzuIhyxN6xzE7RWbykBVGTq8NSDfi39AnbcoKC
V4ix+Ke/17zmKzKNstiaCWUxnk3RD9dwcYnOTSspCSTBDeEWTJGCZeUe2dKuA3Z1O7wQcuw8osxq
TaZgsTvEfceVZEJYzGmTZcYKOZ2t2CYGuG9EdFC6SXpHbXaQiWG8X40BUzmVCaT6H/RZQIH+VXBP
nukg2ynC6Ct2HC7t5a9z7sN0HYJCGnW4GGCxRpKn5WiwvcZU1YVMeOY5hgWX3c86aSgV8d50MZk0
s1kgV8uLWFW+uSm7C0+VC1J5XKHiUHRYppcBzKJ0YZ0mKGUYATdEUDO8/I8UQFToXPS5EZpiXVvF
PhDNkFJTW1wmpJVdlPuuGJfhD7AfHSMSXk4kkx0fwL7ROztYNpYUIeDL2+ZWpedDOSPHrhRzrPV9
2g2ZeTeFUYyuQX795GE70uAS4S4SpPMI9yHe1xGRbRJ3VP6TpbwgHQQrSK4ZsoMrG7NltdGXEJIj
qK43wehIALudo5amnkWeobd2z8K7Cd1xkaR5IS1FX6flmVgC9pTcmxOZWkTMnj+W9Bp6M56+o59t
9TMTIRws6ggtcDSJdvimnZo38EDFFpHp4Lxzkg4RvP8NwHRGlNZodbVJmL5x6rc4FuVOMieM0FsH
ophyuuRF9p9q6iDowkwqJKPbVIjUs+dNSWPkcaqpx236AAQxFunDhUj/qt1PFiNgiCfs2yAJxkDY
2yIlGZw8Aw3cq3JFJ72M2jsfscFYNp/9cFgNMoEM8AU2lR+an/mv6d2xNf8YEiUtElCLvhPErY8x
6wME4pEJWveJXv8qKJsy9i1e6YWAq3uvhFYyIvL5AnDFt1zYpLV+EllmobJVvYp69hsm1nckvE/6
g8/jGgNiybflM7oXxtwk1m/KhgKRndJkj40vglnlqS0jYaLhK7HmWJtd1IROpuIK5O0LfyvQt0sf
o1bU6RYeOwQZKkyYKrfRQqY+2uEFu9Rxlpg0oAK4oxAnZ3DsYRLw4+3kkFWFV9nTRmo7pmdrlKPS
MzVVCFBZaDHfIDbxKvuUOCyMZ0xQtUFlkKNIj/NPdCRtH+o0EWit0714ekLG74ETcHJILwZojBtn
CPGaz2Iva2YndMLe0xVKCZgZBoj2uAQ8uryAY2dVk6bKoFb7LAKy+7Tej/p0WioaiUrdgk3M9+pd
jnQDx60GKSfKbg55N8kIlqkHHhn2aDQPZlAnvZcQv0kKxX6Lpvl6lVvXJy2so98e1lzSXm0W+SAy
gDhpkUGPjplhq6bpLThZVFI40JumqZz4hW9Uv5vA39pdshCyZQ5r0ckEZJ17Ktg1qOyCxYa7fTwd
KMW7HLHCXsefXId02one/w7IYrWTAXwKcpYN3/v/NshN18+FU5j4Gt8jUkO8yedDQTgViBarpnV6
oB4Tnc9dz/AdwxJwi7b/uo76I8whaIPg9ZNSdFHFC4Q3PdjMWoVP3e6PjsdARpRqRQh9riLvUvsM
2/7Iw42zPvP+T3QwnoxUp+8wIwetUtdTVg8tVjmzkhJVUqaiAZBjqJXiJvoR+L2H0Y3Jg5Xq8Goc
DMZWB25jgvmZZbcW99em3B2tnoR52wSmFWXRlbf1a/9/Q466/SRS0NBnmIS7uZuD1CKPGlYi8fHa
EEXYwxTL8gkNfo3jKGo92LsokQDhjOGhsxSvRWv3XjbTvNQI4WA7WkkOykBP8h55NOe4LTd2qZE3
IVTo9JkKStZIdAj2iqhtrlyTd/0Rn9dmigz8ObLAAeEglw8qnapzsU1LSlJpavQN2whAW6akL9/y
iAZwD5xC6ZQerGCgsAl/7PdguNxnN7ehRt+lnSmQhx9b2by+jvftapY4uXNC7pVHUJJny/4nSfFz
E//smqxNBQIpkLcAUJYRzKYAPDh7LkZOeSQXKEWhpBjgacToEfVU5mUw4GGtQcdqS3hbJc/5JOPu
n9NGedJIyAhAq3l8KdG0w8Af96o/CNCVpzgsQwrNsryaxIYpjfUxkpIxfRj0pJ/bT9VO7mzJ4Hju
z8A0PFGphOLVvLn+2Nupla4DxsP6PHO8if8Dt7AtfhHoTtATmuWFdxTCRegIH5Hv0ILTW/pA8bwD
pLiXTtZteRO/dXZOaYnfxRSZQtpL46t2OlvLSJeioANrwddcRkRROJXD0RoDBYhaUH59FOQJJpMC
KhkhubbwTsO/655LrPkfcAK3X6wlPxnyGlsh+NKxWrC9hRlQmuhtNe9C316LPMiGIMKEhnuW/Qpi
2w==
`protect end_protected
