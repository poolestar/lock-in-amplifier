`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mnyeBxGkesbdpoJ5mnPm9lGgRzZLbO1lpP/OB3LNddzG5vV8hs1ZR02JYnll/fMJv9W/BijeD/Ds
GRXpIWkMEA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TGCFvcPRdDBG0YEmp1lTZ+ezzVZ/UkhwEsQGokdyCZG3IDz64Cx9wgQNj25QFT2Nsqb2/Tlx3909
hPC7+eYxWPPmzAOK57FWLZd8Ms+LWRMgYYCHtbsHrGgkRKH4YT82AibyUDyfb1M/bK5db6sZBHGd
hl2rw66FSGPXEj5erZ0=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jqOeHaDOLDH7cGFZSAVWs3mVcUILaaQVu78WnvoFYiUKJgKiDYyoW1eAEHguaxGb8M1XF4t7qRPt
NGG36i6Vk1R6QYRlZqtUbynbvJI831veZoWCb9macE0fvQbbVJKxlwq304/E5Jv5z06ZAJ/pwrWn
G2KJBwmKeVs2x6uRzYX5qysZubirMvgoUUpZAEUz+c0OCHBVPNHn4Y+hiEjO7ngCafzIzKBPhXsO
ii1vVw5KDVl5cfWS6FBwwFrVkShnxUnY1Vu+JlVDoXYRr5koTOplFWAhRTz1BRPiRC7qqVrNDWfJ
9Rr39R8mxAS59Hx57XJTa+Zfd34ysAGkAJGUXA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
y/1zm83TfzBPWMCSRNXjBAKSwilBF3rdY5k4zaq7joxxhF1fcHVx7y2aOijaIyOqeKgkNY+dgkAS
n847VJdj6U8i5yYwi2Wj4sDjdps7GIDc9YJdo8LOkt7Roc10qHJ9Gp9DnyQ5orrj7MC2Ruqjpo6H
4RB0BUUgP1Dua2WVIII=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
M/P5pWHqNuaIkrBGjLLlFOWYbCA926EoNggnRaALnS8BTslbDIXEJLsFtw/wsEAGcgMse39BUYtA
K6aHty2dxAdyTozi2q8c5wDHzVFwPIi8S93Lermf5SOKQnB1eVg+hFB7NKDimJ5N5pXlAKj4LTcD
GBVqV7Lqw661xgoYoZ6vS1h5HZKSDJvyMcYGHVauqKkgtar0cZ7KbD4nd6nDKcHC5ypPtuSyoDEI
YJ2eFmxmVhY25qtfS02tC/ol9OKX0TEeqz2Z1T0t/eJ1TvecYCN2GqRbDsS2hE9atLKf0ezqZtmP
1fIXKeLVJYsyLSbEnY3dH02TLBiCbXeNxBUvFQ==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bgdwJHCp15hQb9R2TdDSAtjWfcCnbiVGxjOg4DHYJthTyLtKhW0dcHpafwYJwdjA4a9jfnll+BUt
VR+TjB6+cVLVB/vJSzCdK7pqbG0zZsInd/PtgUd6FwgUT4rVhxvJ1eYbISlGNfp5Ls2CxOwZ8Sq4
zaGHq15Z9vt1EBxHxVwSs0SHnOtuCg8S+iIArkvy5VR7j+9XukbgG9hsScDPWZaNNBSQ3FPZb+pi
4csjWx6LDnla+7rwF50OQQv4GyB4h9WlGYuZhTx/GKTJ+fdrpUpLA1TBnX/qz/xNqF9QZGSXOJkL
8a9AI8wBSCsWhvPdgFdjRI5b80brauOkGVrFkA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22080)
`protect data_block
p93TERkFAfEQNkalI96DZIdkz6lMIi2m3z8yvN6dDpKGafRmir8UPbCEjVwLTome4NTHMjd1v/mY
obk40x7Iid39BYTAfntBcLkvAf5S36yPTQoDRjTvnsBbB6NB5phb86OnU91QXRMn++2XXmwN9DY3
kObmOoHudPec+Uk2+4hCmDsq+JS+eURR7Szv2j4ESJ+ErOH1gffL3Gj6AC1xf7oqI4qy/aAxfxQB
qc8HcTP4o98Hs5m0Z1J/QZZsyTCt9w+duob2eVqQOmY9+Yq0+/L6/W5xLF/jvjfitZr9gfi8bm4h
B7f6fLmNG4ExmNW8hJkEKBgHfscet7WcvHOlTb2uILlztbByAGaQuIwP4yI0ApAerNBK545kGLNf
v1zfEG3WmgBbYG6iQjKBefC2P5qgVlgbQs/r4RbChWlWJgAiUovg7tKX+hk4Xn8DDEvPImdxkGUH
3+kd6pnjddAlV1JGTUIAXb3I1Kb0VHjxxrsEviiE8sJq8RHZ+hTSBBDaBp2lnw4j1BCxy60pKYVN
E8QrFWmQx5sVLsD9kO4ewc1HwtJYAkEQ4LvVe8qrH06U8061WWwFDw7ktRDykCkJNF/KLcG+PGfw
AT/mbGWCUWH9wTqP3zvcbWaT8hVcGVOeJUDn5lLUBtzxy+ivT49fKXctnQ5i2avipJiiJXFfmSoa
hNIUgd1bdEzGDcPZ1ji6C2wNMWbIWJF36BGki7ftonv35m2I6osCbw2orIK0KaMd21sZtRQU3qt2
Xq9JV+6uFuZqWX6shZIPXnnodH/QVnaylTdLxwPkjAWfof6fDawCvXQcBmnufdkMo/mu4SBQtbfI
rqyIACGF1thJ1l/7/GRDB3ikaAIIOlAVfNBjjHmkxMGdNQwCMHrzvbgEtn58WW95cEf+vt5A73Wy
MeGOsIJajpmGnBfZV8KPLtWaGUQO1txSkZL0zFA2AGy5bDcyVvIm9wG+3VgpXdBlIgjEoWt13W3U
m6SN2/vTc4byPqwAKWTOvJdH96SWaZraw3rvl8bcX1hKexT/W4m226LmrYdKxaynchLwkLEGh6Z/
FDOFjxdrHNzOyliTQPFEh2Je+E+1UkehbL7VuT4uXjH75DfHpWTU4YMLdGqTqMbAO7LOT87BLYxY
NkiEhCvInhE1d/StsyUalAYL9ysVrUbqBgVMOeF4z3DTUqr8Tj2ttcc/1gVSG89QH4xvk08gVit4
zbN3lGY8senUCJQczx94v94CernsLS6NT2DUJFmU4C9MS2zl0ugraySMOPR8SU2DI6ZPmaOPA8xa
6Yf6VmQc0NNp0u9gh+WX8DkvowJbXnO3h/ZGZlroJQAvbtJsKSFHvLc0xsPTWiump/gkrad8xy+B
/mBJUG69lbf1IZ5d7Upehphvbz9QsbD4NQlTVprg/R+RGPHAuU3CGThAtTf7BU/WwJV6RsZuU7Xp
Dn+fdU17Q2Y+we8X01pmfIeQ6IjAzjIGR9xQ9YNKRHS5NwUeAxaKorb3+jzEK9MKyHbCPbdn+JQd
BekbC9/qhFv+c8FY+bj7eH+v16BZuN6Th+649Lqv+dGik5fN2a+jxQiTWr+1rbIoAhG3/AbDljCZ
ozbht7l1Oz7eQ+bPVHKLR6VjYyzyPEatIkNBV8kUCHJFeJ3bS8WQQ9j4YrjuXOH8yKg7yHevb4wK
BPVc7nWwuyGkpRvs/UugMvwUC/fzHuRSGkuZVoxNDIP5zug55ItgCZX7u/2X8hxJsP01srImKlXC
WtcWvZrIPqYxRK5Th6XxePgR3VxUNODHx7UEssOwNwqWmiE5CJtpM4KCbtvY+9Lq1KAzAe0mQDYW
JwIjnsgtsLsLZG30LjXs8ZyQTMvZS9/Sj9Pz8QOAks0FFP1f2bbews2Q7j2CX2dMlwC3V2guTz3m
RMqY1v4Hjy/tbENPQwQuIdHuanMLDe7LWg3v8Z5qxPvJYFK4W9iafC5uf9ZpJk0FXvjMpjiyXs0s
Gf1wYXcdXRFkV6DLl2mvBPI2AEzyhMrVhlxtIxn5AaDoogF/G9pP45tmZzyAvxqFGFN+kg4qS4qe
TwQLXnY7NgYeNZgGaaLWTDnpMJY6SprU+o/x5qvMQAebCqdByjHTrEP/Cg4512rSTGnImmrzSF4b
I4Wpz9iDIBONW5XuS58fQSLtLBb/H1DTTWyExxE3UoEkIMVQLmcwjfG8s1Uypp4lf/oXYeKlrDKF
3ovjWl0K/MiMWTg1uT+UEkH+xZhyAMEOSTBIAihrGO/DW6tBWUN1/FQkiYmHV8iMJwziauJ7Ilcm
UMWjMHR06A/hfStMDKYC4wItsNAUxSpCL4mGkw7x5lKz/5Y5LYy+MqCaPQNI5qPg6hvsS22j3pRv
rqlxr7c4gGULyD5Q599/5zMDy8qVP8yFsnLnpY1dw6lN0gEoOMaYU0W2rvPW6pkY/EZIKP101FxT
HWJKESHvkCrmNr/wbg7b5pX3gkFvoFV6rH/sdIn5M8xOC6C+atKS24l+nV97jjVZ2URIDABc57oG
JdF962mbiYffrTTo62pH4emVPbc+objJJnFQKposNmkSvl1hCtTQgEp5Lybs5AjBkrAS9mcCq3d8
8wXcZ5jK7bB1bNFWyBQdxqn588QySSOpJpYMu+Yw32FX1ziFRMqbdwqujPwVQmEsN/YW01wsYAEm
KfwVCrPzaiE/r5AWXhsLGfrfp2cluda0ddYD6MfSRMteeMlswahlzTctuZuFMfTCunjkPwaMXfLK
O+3i8bf/+LmlOxfPCU9n7DuOj74LLlTtAGQPaYDrZ5SXhlbyQZgQ5jMCNNDql/2Omy8sfuOIlyUJ
svi9Z/Dae3k4ZtIWKlmRD1Gs28n/715Kd4YDEyXlsil8Kun3qRioznPzeIA2pxoVrMTwW2SHG0DZ
9LZxJS9RJUUjucFJZu8JyAfBMLe9PftaOe81oExpNuW1rbr09m6r1HxILKY+JUeQ+kz+7aH2cYqD
TlW/zkQkIGrZyx+dMd/6rkv81lFlRGCBT8uv1P/rCUFPH60UFYH3kAZ8t8pmMMDu+zA9qRLhSyqI
X6q1VpC202cyclPrCZPvNC00Pe5RyIHa6V+6iurUOD/duCFWzGCvcriMPSVbh9/NDllbOzdYAMDj
2z5DAiLmJnjnVoSrOdFX4rTJBpX0dto8xi+dpkNuL970NaCzYxJLr12l3nwWeO50p4OdQTJDxBMi
NQXM9mqny/g0+frm3tVglJ12GuceXfBdfQld63dwgsBC2tvGZrrf6NdCs1u5KCxBAvwCXl8Qqp1L
BkjYGuB5/h6RVYzwzJJ3Ie1nEcRRs4+nLCZ8bRA2CqECxHtWLHcX4hwLzft6wd063axPrrw1cG2v
wwPsf3aFqRf1NyPrfKHHOc3KMb+D6b/v2qMp+1Aj6uQtTi+n9hHzzGVp67NBrV1bqXXtGxXqtQRJ
4g2Gqkfjls9xYTtZuvQjW4rD7mwK5rnoIHRhM0oY+ItZaMIgZTnAFUNYD6Dv/k3MItuSRu+SYwV9
fY1zDvY6JLhAtDmZ6Xsg6uCFXT7OdpMvOZWeCqPKxPM6zGDySf6yvCLpBFgAUIEyGbeg1REJwu5f
wumCy9/yVutd93/tyKeS/1OoTe/efrqT5W49uBvmoW6psRorZTGyFT/Tv9K1cywT02LDBl+FlzLA
oqJSXAOKmwxc9cZJCGrCoaVFXKN2RfdtvcV6L4PutDdTzddxrQpG2HOSAIsRcuhNDgxdvPxVSJON
/zlVxy4Mpo1jA4o3LDOHjYEt1M1n/GnrpCHiTRdEA52K7YTn9BqaMMfVr8LtuyqkLhhwiHNpI2pS
9QGBgFxprlpvYL6VHm4GxmLOIwK+TTqRqinuyJSNGKsjRkMHONk7/kQmu1bXTeZKLOThLADI9FPJ
wart+ke7dFr4PJpVK1inxz86cOiyNDYnTAjP61Okby/fucs4ykptAVe6R8cWnEDQ4z85Trn0JkCA
/kEWOVJisBii8TRMBXQPNBRmOin2e3aoZoY3HKJQ0ztAQL+syoDyLm1CMfcg6bf/oW1Y8ZGBZvAR
iSdwEGVa6wKOMYHqGEOapVVpiJpsKXztt5jjfETVrGij+qN4+gzzXeEMBarClivRwBM6h/OFQ0vp
Hl5So1hj5w+DtpgdZBO4EGZB4L9yyhgFrFslrRIQzT9fT1U4Ac56RAGQFal2BsvcoxZxvmbXWXYJ
ZorTWB7M/zZi4bR7EsyDlpX2G6xalEQj7y7Sz9VJyNbBucWPB/oaOy8BIPSHb7H4WTBvRrSRUfTA
AIjX1hpCMLbpS5tbG1pxRccRmRX/y2UdcC/vWN4bXoKCGXLsVIZLKGgLrkKXXaDf6vHFG7kT8Nlp
8gsTUeUj+Egs+fVb7HMNfb57YMKNgpKsWMuqVfWooGkJWFZ40RrpKnRTysDfFlA6Uo1mY19GiFox
DVyUUXTcEzlB2u5VK9MJsy87X4uPqYHPQ/L/ywuQEQzbhNhuoH5mO005OzGR+z3Ofn6J9kr+nnZa
HLpbEJfSTLxpwebTa7vL2OwOwlByUwdmogFR1lwJKqIgq9tWCzV8aPFP+yuheW5XFRbQxvKK6D90
f+Yurq5CVAWJlV7oR6i4mY6ydgB4jfU6epPpZjpbotdgKw1Mls0Yj4NHsDrcBaHMpIWgg+pHVsuj
ntZVrBEcfxF07nT2WCoCzhCdp584gUpoh4/ZClzGTv86bAtopO20UJQl0ew0k0FTANpJgopMYX+C
f4+RCwzOAI5Ag5hkwyQJmM2lPbHOq0b3NN4nKpROtAzxpz8+9unotRZNVD0iKdS2E384570mBkIY
j7YG3pb6QHybJB6AgZHQE4LvG9ba/wVHlGFn1FtqSRbaengDS1h/0dqUDLbGNI3TqcS4lFTjd7AA
8ggqBElKFj5RY751Al1zpVfyA6h2JkURBIaBjxSHmuiiKrRE+qzLYZ/aKRENSiNQD1a7Yxy5a7tT
8deFc9GiR+5hopab8yOUkeg5YeLo/d4Fpj5dnpnbALBcHbG9swcsEoLP5uPcCSTNIHTurZOBIb2M
AZenjm8EozgbSrb3IxdkokTAh29ntbv4PlxduefJeNTT+ijKV6z+Z89OR9ll1QXxrBQNDP1euoDV
Kpr4CLHLz4lTerR/vJ7lXYyFGjdig8gZ6N/UxCo63R0mzhcacHYRchJfw+oGWMJnBc5RF2PO7QfY
ie9NEsS5mciM3qvwLrHmoFWif+qZ5eAOSO7Rmaxx+6r8ZcR2oqKUvfihUHNTzYvMcZUE9ZOeVJuS
yUaYynhXGaFM7X4lCnAojlAhvKdInmn2QYi9CTTGCKEiDMxzB5RIy74mQIIMBLFVAykrYN8lI4Kl
IJfJsbL20uR2wY6f2wazOVF8jer3vFveu+SsGeq8LCw2acyd+a9ygDCPVf0kpyf8NPif+GtirEAO
jsc3QorIYjiHEMoGeK6BsG30Lqjchy2VdoAL391+6OepPbzllZSw4GehO27Ml4J23FWIGpPS3MpW
FSQwr3r3fPi1RwE32us50q+lIiNgkJICUoEJm7pTSnZHYUWnCkBjA+7vNyTfxifbXy17spMJ37ec
S7dO0mE3GruzUuGAJaikPsnGAKZyrsCEq37E+d40idNIZW9YZ2G7MIMGFZPPpmDw5PKwWN4QRgcA
5euVi/HE0vJpjTQn8zF/1dWDNE99EAGJQHwfVV0JjjARw8XRyZ5x6P1a6ILRlo50/E9S4WjK36Jg
8lILIp5kUmyr3UzqaoJ7Rp+woiwWVj3OAabTugNLlWmkDAicO4v64MnHhWO4qDQfNJOZeRooregW
9lSXjUDB37Fa0ODKgym6mo7OKZpSKQvpX7px8+g+/UhCB4AGMYWPEJs/Xo5nNYJf6RgLmu36ol59
AhF4KKM5Pze2TOr5T2I4AqWhsz3y9Exgc+/svcpAPqlzKn/86D/PIEpIHMtBzsWS6o6J5TL4vhEg
wYmxu+7rseZ3FcnDO4JdfGz13PyM9VCR9ddIxib0zMuhqse+8XGgbDChTWGezeXCcLpxo9PC4nQL
TUtw3POzYebz74IDlptbH86L26fkRWYpm4+5CWo3Qh/WfVY9ilhDdidQHInYg/9fSFXg4T8W442S
R2MVzb3hq6psEKxwwaPhw35RbZlroQMiAi8Cb1zM66VWGd8CMDEeN+Ony6/3694qNfZN1WoDyDe0
qQSN5NqXG+XCl2R4tqpkOu18e4QCUfF3FZZE+LzEYfezSMKCcQQhV/IZ4YiDeiD4Jms9fQ6nbRxw
6jK4uhQrcWKTbiCmF5ACtdWfpVRIEY9WLpwGNvu/bXUl4TjLlSDBKbaoNPe7AxFrpDS6Bfxgmnbj
8y1YRHjOPBJT1L35RvRPqGi5bnygk44/NLt2qlVPC9RbF9JTgeCiiObVwvOAvqTVVSi5ny22suef
J1mSQacoSXhtIOB98uPTQm7ac8PQTuw2DaWgJDh+ogWIv83xxDME49+pYaVMxWCNL6rXctuUzn6j
yPb/qQhwxFxXsLm6qQNVCUINcLthGcwCeq5PcHBwsF2mMvP2W6UZENm279EdVOyOsKsNBqAtBSq+
g5Ne3DIBeZkMwxTOUZhPC95GJkyi5MLn/cwIRoPaQGBDUlOWN1HcRO4G0zTd7sqjyeJ2cKLyqlED
rj8cgwYXjG3LTv8JnB/Jm0ghrAcmorAPRG5K4vIEgdP5LN+AsxKMCCEH9OaROTd7OF5V/MctfHmW
FMDw+DO8fBzhtBJaHL8LpJrBZykewLbOg31JWOG8S7l8q3OWNtDPmFINeJ+JD7G34QgqCCtA6mWi
4RWhhiPmXwY2NiL3kIDKY+vp2h8+uVhJXUW0VqjcF9obHVJP7/CjUMKkX9SGSGMta88v4W/Y+TJu
tHL7jxYsj8mKyeQdvQ9cKaIcrfhouiUqbCPSLDdzmV2Qwt8CpinBkGNr1gxAcmZzr1exwMkd85tP
yBgar17TpGVc0MUwV4tT98jiFh/gmVT3j+QP/uCKqv1OYVwg3TWG/ztIhYUPJFrMLLC9mcDN0uqG
1RB6hs+O3GASqW7+ShgGPNo1r9Ye6+MXL5vfH4gnrU6AalLp7PdIcW67kVNrqEKVveV4hJRSunmk
gKGDDd49UB7v0WE4YHgsYbxDys4QFB/m/tQfvO3TdT9M9Atx2aojQc5he1QZoKm+d1r974dx4MWK
HldQGvZSK/SEiWqfqlZj7lejem8uuhv5dlm1PJs6YAlRT202q1afcSmFqCjvj3no/QTnBUzneJ7s
8t3oiENI/xqAXchY5i6egp1V8EsXPAdoOiKdzutv3hgKKFYPBv151IF+rio5YI4TmbzeWw1Wqoef
dHfbGfBdAswbDPA+1wMxLD7ySszyLxqu2Ev1qen9Gq/ZobhqTSM67cYJmXuE4hDFY0h4/TfwMl8h
612ixdm6z9HoloyKwk7paoR8zDMHRgvDGUcGh6xXujBMbzNVXCmIb5yNh/xW5BTnfijN3M2pQe/h
OrCVgMffHQl+sXy/nkuLsIyzOGkqlUEoMXIbwfwWuYExeK+/5xuWHOmoJlSBu8XwW2VrmEtE0Sok
VrmxdQIP8ycicSZSKTDdbZxHuRu1CY6lthsDLTPCV/aUwThhgpkiazS1FrR79wR2ubQaLQqyk814
gk3mvOw4/99Z2c7i5RNwp5Ip1TCVmnaBpseUETVyhlKr3jHHw8UFf2cUGAM6fwJiMV+UTIPhAbR6
BIpOjH5X1wM/phb99gRYU8v0Rvb//jFeQdoxk6fhU89+mLEii86KAJ80UH2RqyrIAaouCIMF9zNs
sA8mZ530D2AB6epAGZ/cNmrrem0YPbESyzi0UIOiPFwFSO22j9MRqS5ZKZstU0efGv4ztfLgN6Qq
Qj5ozVragwo4SbluX7kv2D1QRMYNmhzWA3TQ1e5pZnzVqlqNcHVL1GF0A6bB0ubKcKSxr5E+q2Ne
rAQQ5qgcSaQV5tJpCEU0iYENZWcXWTbmEkqa8UUDHGafeHK8gDqvIuOG2hfD2AVTwJqwJMiZH9G4
lLoFxlKt18h2KWTERPhAIvk7PoG3JY8rpkqgcc16Q1fL0qhUWKlt2/nxkKcSYwZzJX7Nj38Fxzgw
n9ZbsZXWJQcQ8RITvqBtZyHQvz3VG+FbOZrDFM/7+M2fPSE4oLJ+nJDofsvEbzT2Unwkkk9PIbeI
NYYxwmPeI8rDDycU/IoZCqT73vUgEz8SbpxaOav9T5N/2LVvrwo9m1lZByx3cbBs2dO3966pu+ue
Vr5KOjonuCUirFrSNM9fSfZFKbw3At2NGky+LbHBFSTI9Y/OTpJbEiursC2TdtE3grd6YA+rh1SG
YgS6/7T1qwEflkAFbfPz1aTC3G2/oKVEa/Mui4Qybs0eBz436vcsMDheomCXLzVTEdJ1gfLqWk9s
KrwQ3YS2wibRrkrdED83Yk+z157RSf2tx6AsbTuyh/XjjmepxmspUVUrSwQoEgqZwTGsdrRn90gL
uAKQ9PBTgIIx8H+pR5Bb5YfEosJvQYUaUHg0BrCHBsHzETB7o1k24SZxTgwPm+sxOJJDLMeDDDvA
OtosT6dNg9XKjVzhmG5ObIMccFtL2swAp5YXRE0OZOK0s/cczlNeHYtbyLe8xF91YUeEHl1kh8xv
6LPo6gCa5oPJ9OqGj77zrx4Lc+aCNA2hXIjOzM8GeFcQP6xVYp3VF1O5aF6SKIXHCr0LNJEF4ol7
webvQ7mfCw7O074kI5oaHHB3JI7wPK3V9WHsGDOgnsfgf9vIKslZhdNK/4C0jAV4lLHy1O50ON+8
bcwkUtJ+QgPdhMXTjGIxW0R68BvrjMio2NoXTcfrNq29spHTNFCQmwoWkM3WWUO9gm3E/rTcPNiL
VKajJaFE9JrLrWMGQLL6nQjdwR6iXtLN+gjWS2Qvz4bg6eTPkmHERUBomY1L4B9XjoFWG+8VRrs5
jDqkUyRMaUw7n1hh/Wa+zFBrf7UHSyHlIHfFwrgZDS8AGx+8IZ7muWfWUIR2iLCIm4xg9VmPDsmn
9b8D/ZALio0DaS1apWd+McY45Zl4VrHb2kFYNrZL5AFpTEVhMog5EIZlB//0O6ZeNE53lSVtVQ8n
bFmwVdBL+683H+f7HjaysxSsn/GpznzEc87nT1sazjLA9nofqIIt6e/o0cvoHU1Ir96YwKyK9wOG
hCKAGZp2EKsZdWjS+tnUoKf+ZEkz26QO1IOAqiGI3aa8yEyaWQ42sBsa6HQ/cGspKy7WyUnXiVOJ
5mVdnph3YiI1uQTLQa0FGOmQ5gKyv6kQM+NHLkkdq5FZFFCDNroSLrpVL0Kf/pr0Q6rCW+Z2Fxv0
gN5DA8sUgQvZ9JvGGfdntxkUnVepZBB9d/Op/w5NPsLJ9jhOVvYzlbGeQeCbNktg+MmqdJOIqOvV
orRNQ5LXVXZjPjoAzn9HBPS24NNZHzcx6aW/6F3/3drgIMeAWsppOVAtTyOWv9miFfOQI9fO3y2U
XXMHPODP+0XxhlhN+/eaCAWB/DhdNqAcDAariIHxCjQHKgMW2qxWk2NDKf0tNHU07hN2xAX1SZmb
fBiGDoR3GhLCFOtG8DS6Qr4/O7qX/bILoju9fLU8frusGZR0laKu9cpPbyipDeKVO0tgGs9kYemo
K2FUIokILgienc4n/cUggDExVmDnaobrs4OEohqfrD8gnKak8sZqcCmRKzKwtTkNkuAgghvYZ6wR
U4kvFC7X3Yi8QnqXFUwJ3CeBl984VHjyGo2qldoEq0CdZBUecgPdAh0q+grSSm4yBy7b+P8nfkpB
8wJ2hzvlBg43br1hIubZawe59zdAQ6PKG70N149MXtpMMFId3Udp8U8Dq0ev6yKpHPOSFLIhCPFV
E3cvvvnt+2beE2loU9k+i1aVU50kSuv9jjQ8bTaEDQJ9XF+nXrBeH+Tt11uTB4ms/ZxAa5sv+LkV
SB08knrJVJww3G5O3G/2g3qyM5NfGnOJGLvIouwmWh1UxBSHwkfU3JbrPWCkiib5R//K/ypFDB+m
qfwxkq+NxNDx+GqqK7MzwlGyF9Monnti1gk0c+8MI8l88QDhl2rn7t0aY9JIzQ4hj1VZAb6zjgzx
h8T5I7j0twN8syGc5bMzWU1QIloX5ZY9sWmV/HVj/ojvR1EAS36f059WF4J+uffb9h5PC/304Bjq
7a1rdWd7vW0ue/PY/VElVHkqCpzn6UYopuCC2R8/BOir16JSuScSejv7hzX6uvO079kp8AufAWv2
GW7T8/a1RPCows459iNrGJOdu3ppveIg2v4IIgtxqk1QMp2mr2v0xqmjYnFX1SFibwA5sQtKr94H
KnvwAecOrt5CL4ok3y1tZgzg8K8aVTLwPs6GLop10mbDq0Ins04tLP0S95m8KwqVyQ4R6neW0lDG
yWdMiuVyjNtLYiw3k99cdWhaJNeBYVQdCenBvQzPaABAeG4YswfSNBxFaH1hED3CwXx7VXeHYtgy
mtMX6zantgpKvcmLIxf+RTmu75eRlUzZt95+ZKgWFYm0YJh885VsnXt0j/Lg4wXymlKxc0Nlq7O0
JrpwrDL9rSEyi352Jkg/wRZ1wBzKUGGng/wdKXKNw4sB+1vmeeYoarTFKrLjUXYAUWTKeJveSzRb
xQ3ZaoaX83NQKjgnssaWQ43+ZWqJLPOdsnLURM0uRvClHxaw2LGxN+3/LGlnjvt1Z0myscOTv/ZS
NnQZIv64fpRC78en3tf///ar4saiqlE0HSsmY066BqB1E62/Kt8XNiIVYDPQBUHtRqxmxYamRjDA
2ApEJPMNH8OResLHgKeN8cK1L7iagLkwxj6qRhE03qGx43D61IPNth4QOBswewFRzr0rVTAn+12T
zheAtEPlhUz6xAB8qja44yj9g35A9jkQPrhcnBbAEIT6wgDoDCDbIy8oLdLn1S+XiDegUmA5MRUa
Eora9jnq7MSK70pg+h1fI6swQfQ8q/WW5R9+dYRyjHbP4UE1KU0gyb7Ro9QbGEshMIZ/mmgSpO6T
iVCYYJ7vQvzTMjl3UhtdbQ7UzzanlFAQMpa/LTpfrlixDRnzXhm8P+eT1pn01xAudeGJZXgrJ3f6
VEtNSyVL9dyuGd9CBms8bcN8uRI14qLg/nKQDOVasvXXxnKtHekX3d7dzOAJSWGA7aDwn2wNafkl
satfnXIEdDtKRWYH+xeGa5XQUhReoVMZ4wPJwu0DfHHqTRSCgLKFavAyjOazXLyHWD79ShKYCRiV
XUV94KDn3uCoqeasoCx9NgPmZI2M2DTS10jXefPSqXOHx/uBfdiNoPHufb3GrGBG7HoJy8+ma828
h7TBt/fgKOcwH2O9krXSQxb2nMY7pil5+Ko6W12/20F0bVp3yI+9pfScXa/8dbFJ5IQBsPLT4Ixj
TKkonwSGE90tgTFBCiuiz6dKi9RvQ9Atoyy4RDRFGatQLuJ82QI60JQvoFIhVIwWagUnogsT/Q/2
vVmB5d3Ojb6Q1SQW7w8fmvyMj9aKd0G1KspLFBhrOnxfH19np6k8EkzsaQPNuTLSZSuUjhKWYjfa
crM/md22CSgkUi98ZyNQRwqnfKw6zKqSDXDHPFYeFz/5U0whwNfYimm13nEzvewAm/KPpKGg9jTP
LDvuQyiMYIUiDedjW1sCgKoULKGYy9+mvsRRTij7PKtzfZIxx8WKh86Lqhg4xSN+5sC7etek0nyr
nv/chgzM7WuObXy329I69IxHLXYGIilztlmOiz51YI2nBPeirBPtqSmDsdMj0NgnVfRpFpyYdD2u
JRMI65D3d88E8yixO8tVo4D7TtN6ldzWOfKZ0rdytg9zsSmVsd/xnQ1b61m+x5X0RYRM1UcTLw+K
od8ZDZAdR1Fz54sCBZWioycDp+XgJEwoM02GTAkM9zDibls1ivdS98Ci7jWw3H839J7rrBdFxEaw
PsXojllJk/+Mj9K6LEBq0bE5ZAp0w3foQKo+gQIGDLkS0HU95cLEPI2/D1rRsA83OIp2JNj2A0cJ
wdfnWC59gHHFNMJ1rgEZ96cpY/KiefwsMpqQXx/L9LqahmpH/BiSyXTIqkGLtGFsRIxsIPksR12Y
lIxcQimWpalm6uk4qofsgr9Nge+pLnkQ1NZFPE95lgXpiswc88hB/BT65TlYeftSFKhnLp3l/wc7
nU+IRmJst7tasajkY3E1G+THdM4QHawd9Nsob0XYTFX2ENw/dP4XI47D4Ygb+m9dbXAkiruxinMb
EfIVFzut0tr9r/z+lNRFdsC8A/pkp6V5FGG1CE4WTCNZzR0Np7E0M/jvoY1kdJVhnDXbA/k2rQm2
gZ22eySMGPEna/KFGU4w1u75dXdpN7n7sMEsHprNkJamkMUJ0CYa6KX+bbIA/7PtEwsSqlId/xh5
u49ltnXm23msHaqaK12rxNDI8Pum5tQbNI6pcd5ebfdCdEr6w2qf0bE7lUgukyS7dJTlenT3aWm2
PfFfTw5+0p7axl6SmRIl0buMNtdzARtiiDcCZLdXg1iaLU+0LdSnWd4SFzgFHN3n30mgWW4Q6+EC
KMW0/7EEA79XhevI9/+eEIkVG267/czMuss3w39wj7w2hg0m5mYmjfWnnrkiTVKPcYixbpzCUSvJ
APt2pVUbB4GchZ5bH6eE0sJPC/qMKI3GzBCAHFXzhXnTaPuRd0JCKn8JsRnYGmM0g3YoU01C8wdH
aRckCDBMmqxiBlV/ZFTW/sJAIwC7c7rR9C/icZ6gims0/7xLg3cbvfm2I16bPlrEfUfqA84/7lVF
tCZ4dHBpOUwVK4+laTwjze1+2luPQQU9PLF8vM1HvbbFwegUKufaJX1p3+mNtcfTl3Y98ZUUHngc
jely6Unv9DGoinNzDxPGQ3m2eoI2mlYQ5w45cjZGBWrLv4SN42Lnh5rOxeRqb90LRP+Di/JOXfMB
COanxcJ51JYleB+u3I0ILHpemGrt13xjRZDHKh3UK0+CQ1PX3EtC6fW59l1JEo3y4iGwHO0SQuZD
qgoWxAcBQ59qnXDLRFngBZ7k3CDHJXwPKTC2PUS1kkIXbUUGHntPG1enezV5vmB2qTtdy+A5aeFU
+GRrpxkE43bLFjTgGIuV7wbaRXvJI8uUEFK1Lc5LGbtJX8aN6472rUhEczq8GeazLBkcunQ9cYvY
9IIrLtdtZijOj0iYZZ9Mti02j0DKuKQ3ZnUf95AadsxkUUR/nRJQJCI2HN4YgiiIZzGMpVvu1gkj
Tindvxc9ITc4yK+YEO/bZ9rsppDXA0jxjHQpTZ8Rk3jk3kS0Y9ihwPdVkXEMDX7cMVDU5AO2qRRs
cHVv1SZ0kxH/JcXwwyaS/aJzBmp/Fzv1Qhbnu723kRsRV0HxI7/uEqo22mF2Y3G8KE8UKKCYcwzK
xvDXaKfktC5GrwFZhKxj4izDRdoz/uf9eoNzsz5zpaSQP/cMVDX3T4VI5l1bO2tVk0y7iVlhwGom
jtKEvDhPd4jRWPo6GTYH9lIkwIfk259F0fHGTDfJe6vo4uB777yn8vn8bmskBkChW3tOD8ce0noO
arjoNqa4sFJ33Ry0wT4tIKqafAHZhc/LCvPURihxwDLlQdYCK1aZmWzE+RaybzAfpy6aBl/wSiZK
bmeuN7y3MvCOTou5s3vxCgn7KF/0/n5v7bi1I4HvXbXgKS/kdBj/mDYzh1GfzaMS/tuUgJh66ST6
qEkv6t00xbLLZ3Ew9FVdxJpcqA1kpgyd26HO3/cheku0RAWwAVAkFyeuaeN1+fQ5DT6otJE0HXQK
bTvMpvtVMBE8wMoO9lyRN9MYeTmX/uKSCJWHhDe+s0G64LYkmBoGfkymYvPwzqYjl6a2VmbCtbm7
lS92ZfjeNqHdhxAC3UL8pDz+OCrDqkfPa3n4+mZzgza47cl9cJ8J3m5COaGChLQ2ZuDksf4AdUR1
yGEc9c/62RVpBppKTs2j30WPSyFUWPFUxkEyYsFQNTrYK4Zo4F7Csa/1SnwRpkqrp91gIW/sBKGB
lL28qDLTgAXsCpnGvCmQ6zS7FkCQj5kbTvaF+ejiA2giDDY9vBJmJ15UEdh3I4wjg+5yV7F+xsHi
lk+bYfTMo82Rs+X6wkHyLRl0wRvcrnv+Hoo0yHvAYMWbLG/5TUpnRHTqh0yPou66WfTPZuyu1PEN
HRuBqroX1uGpRHU7BtNz8/Yiqxxpl8SrmBIqK7/Xsh03KOmmdiifbO3yUtkmAW3HFipr+JRaE3JF
ZJo1umVHdZFMHxzQTUh+EfDhdCCyRXIWt0tT+3I/rSDxc0hj3nEZihhziGSoMq43kqIhc4iwIVNL
ImAhP72Qdh8na2+uVezaUbyGnSiZ0R0YTijkCuG1CePsXf7bIXIaCdBBlu/jRM17KqPjHC3924AF
T4yWQ3SqN2cCU9cBO3Nw5q+yxTjLIiTp7MsYFTWle3kpSxFD29W+JWM+qKdcW4++YMOfo1Y+nJAB
inWK6rxCzuwfQUpDzU99HMMZl96YVr6gAth23azHHmqvpBb5Adbgs5Qc/dCt4l43zNjoaK7ayw9f
ZpSvSww+YuYX/AmQDJX6ho1kDvu1yhGuy+ce83JGVfN4AsR3qMZyNLw9Y/sG2jA2gNKQxQQJs2ME
wcXRVd5fAV1QnrwVEG0KGMtrcv/ShkbiRtOTm+obfhF2yNtAzZ8qCLL6c1db1U1AJrbhBvRuOYP5
JMM0ELOxsf8ep22tBAKrttvVadkP55WcWIeBoOXlxVjMAQByEWzmV97np3ieMgKryPO+uFcsoRI4
CUFmRPKn6vbeXZ3CYs7P/kCnKtUzGcTRRkQUIihKIhCYhtzbApD6wQiC118RB8LAKOlN81fnvbtE
nrQcu4ChiEUnRz4xwwAuR5+RM0/2j63BOaoPRTqg1jehqTbDlteFQ6Z7YOzR21Ie7rfeAlWOfxsu
0gPYmuewpi00OnJxlcFkEaRIaPCITjT20/QjZbgBH30iP8mRH4k415gSj3bKW+h8KYzfeZmh/pu+
JvrOj/lOBRJyrUBNzhiiTOqLvumDW/ns4Z6KGZzfJv5p2J5QYLWp0nnzi4tu0EkrIs+86MI1LCQx
plBvcd3WivZDb40t/DAXiYMGsB7k9AglTIMaLNRDdTMPVneQH9BCfqnwXPoQQQS5BOX0dP9NzLZE
DLwE7v8B9pcm+e0qUQDis+M7Zp7/IBbX25HIu5jhXUTb6I3jUjFrninCek12D42BDc8aQ0wscMd3
wobfugPVnUNFamxd3hjE7CR3FUNO8Ok8DNRSxHi2k56yukPDfuCAtanQAKqz6M+apmDfTxwOcoMu
UnykD6eLjz9KwkjT2lNlM3C5rVaQasydltz5/3EiPRnBpAAzPyhnWTYlb+sTeDSeTpP25/CyuXGN
D6EHKCioAqiix5PCCzAtoMcuQCfzrtJYPJXpadwekLIrWFNExi6TK59X5g6H4ykEOUYUIB6P2cDm
6uKLJuBZwePTxwwUL6Z145nWdK9lRKNzQxY+HbgVg2vP6v6FfmJP0dU2oBKQkDhYNvIpiS5CTjn1
dFaMy5EyO+8OU13MFUdCUAjxbj8vdG6e97Mjud6EHU8wFgElulyhzG7GYcqaoyYesIS32uiFi+bg
MDGIwaNnLfp+1oSzb5n0iGv5hqMOhfOf0hZumL3Un/GeYKDertgpjGGMLjYFl9qdBiGanaNkBju0
coHg7ZndHVQu0Sjsg9DsIbBJSZXj7lXknRf5HHrfUzcLwV6JjG0tYDPi8lSjmyRTynpI3lfmoGjF
dG8E5r5PxjjJZt8Uwq+8Mt/TmPFjpYfdPR2ShS8rVFeWs7dbt/p0aTGWUQi8TULeILP0oRvNb3Nr
x017NvRHTtgXDtZj9s4TlyT5cRD5lzjlZI1q7tj7TYvPudWDs+Lss4ml96liONU39nW4z5ZW9Smo
6rZo5TBExGHwsRknFQgQiPA15/J97Gsh4zqjU8+YT85YFtD1vDFIEn6tQlYfp6ZaqcAsb26ZW15G
5SZxnD8Lx39F7VPkCDHBAbrAVAoGi/NbTtXoYZG7VEPXbzOL7MtlIicHyYqZGc7eFXXA0MPfuFws
GL9oaYWGYYryAtVXww+gfLBtNIRl3M2wA3KzsOu4TZYbXfch2MnGKQJDskvyGYMnVBdC5bcwZeFg
t04dE63LBZ6CwZUX7htQmwEE/rcsongoP9MelS8knn6tY61o4ib5I5oXuGJgGpsT86zBiEUEH9b4
Et08SLs4Qa0vxKND1xiK1FhqZVWzkIR34/k9agU7iIjYd1MTZ5cRyvXgVBRADn+cGuG56nc7jwRH
vChmqeOLaYKHxC8k6+OzqeivkHci/E1bNLNzwtikxre7ql4+BCNSXs5fBpSVHMZCnHuX1NTpfMqD
HEjwMCGjahpfGqcuIRBdxg0/QIpHlXvAQKP2/IEnq8yZpoKdqTWGIfAbmIZ2JKY7eEn92TyTBaHm
bbbAvySVYC7Bth7XyxJthSsw+LnxjcmLmvwlsb5UuVLyWAV4wGTdE/5GjKi0/F5pIidsVZ9iXzeO
6nRNDuqlJUZRPRBpZehmxEIebzWTJ5H3DxIalqfUYLhgrkj78HLzI6BvbqCJAV9kgnjv+B0Vuf5q
4I8IitzaL73PhwE3RckjXvfG8xpxQ9bgZX5wQbbI0nnTulUuyAxIaKa98osaCvEwQwG8KIa0xM3Y
4vjHd7B8fnFDb53u0qMBL899dRftn3zAM1cR6oe7gUnabuVyYKna3rGRhVEJMfmyeVDN0lF7EMny
wzG81eV0518PD4F9MigWBu2BHSFzpgGLhSliY0UfigttjrUh15JcnhR/mINoDaMLmkoUZK61yEyW
+UcDBpbSoX62CktbOfEX48jl/P/UL9ZWUd/fIymZjZY+WWTb+BH9ejw7EN4TXnEpvdEM2QGzb7b4
TwWX5KXn8iO5HCYUjPjDpCKjNr/03KNXm0uV6/K/via7DCctUMb9/fNF7b11ZtDjYanaALcAjoAR
J3NBjE21F5pQNgfIi8f31i/tAL5cMXm+Imnlm+976vlhpAlwiAU79eow5xIvi7xSbSoNLjqJvoVh
uWh9FMpF8r9pF1bcllLzR7FEW1T2LZt+j0d/gWAByOGYkpDo6s7OznUpV8l8vwJ3wdoy7RL/Enke
864Phg+Bm6OCQF9tXnuq7iQLBxd7YiprYJrLqfx3RYr2rRDNpjMLCxMYz/pMoL+uLnJbTjWWT9pA
TBv1dfIMlW+I8LygRn2qaF5DTwyvn+86u0LpNkhZUqf8KyN6Hq2YmP6r9Ut7iRD80JJokQcG9gys
sHKhwE6GQ+SS1sBYAP7aNlxyxG3jd4tB26FKTs30xQXEpl1KSFeEIsMOBz7P/N68QhQS4AB8vfoe
EnfUf0GXhQEbkZPdyK3rvzsl70T8mQRxCexmANKbj6oCL4ID/rhxySG2keDT+FMecXT7ESO76uWf
F1mbtviMv5bvr3WSEaO+PSCIt/4V86KUBIVRgoVJJJuTPujf/Ga9OZ2OaSnpWQPVcUOiXvK7FwTa
xKRUmEB99Eke8M6/lxD9Ynxny6vB4caL0zQ6GQDjma1D0y/odcAQMsws1cSMy0EE/kMPPUUuaNGy
7Uf5Jeqy8s2jEJ4XPBDZ6HixXMPvHNVr7lXSajS/z8cKaK0kVoXmkub8Vlaj/hzU7zDHK26kCWuy
f3yY7VrLy2cISsp/Dzas152uue8lkbodu4Nepmj2hfGJ4r+PUj51MibqqFYhnACituecFLCkAnEy
0qU/2tgi2WKVrM9wWH5cgvhUKB0wOCFyuZpdJ4YUMKhnaymqXBiMTZQ8IWFERtokdk5f2Q17mewH
dA19TxOCSpikhLXyos7tPsIpwTacRMpozZduanCnjpkfyMnCGPGXcYyMVAhnTEeh+MAKWBKqtTil
HV9hxVWOlPruyibTBevHeg+Od0mGKeevfZJqVxodIGlZl7sy4oVW/fNxT98UmQKDVY/RtyyULPtm
akQBDIxSfX6sTMCJF2rqfNShXtDS05LOalnpOeZBJ0U8rQAV9jcc/HtZ+T37ryNi7OO0aMC7/NaO
oDBw+Fn/adQ08icJoV0m2OZ/zDM0RNCOknXjv2fjJloH40h1OcTeK5CRGdcUoUljumes/A0RoeSK
H6k3DLcEe9kElsJa1nQqjGAd313eooGYSFLRmANmowgk0uyXXo0mfEXcITrhqRHUekiPgKHQiShI
EHQcvWxte3oHMnBUIuAR9zf2aHNWRq8jYgXqnpp/hIZPE6ofbJFHiT0Fkwv3HmxShgqx7zladFAQ
JU0Q0f5f/NfgyMUS9UMmzAsBxAEbXsxGubIsfvFjCBzBk7vpVp+fV7RWOkygsCcRdPZMPdXtwArZ
0wep8xqroXpRWtHDJBXWIHkbeS/BcSYn/7buTdxja2rKhM0I8sPjqmnv++fIdaw2x4mDoiiZdvUu
3UmZlnC4qh2wOMtzHvc/aLUi6vbeVxAloM+s7UqlCY/FrNpXTeBRJnuK8Gv6C5xaJiyPc+aEXSNV
PMLHAUR48K7YYL/WdG0EuEF6I44ado6E7kkARkBNrTqxDnFnoUzXIMqzBs54hFlAnlSaLob0Iflk
391/o9d3V/giZ45EW0Kqd81c6EvVyHpacP5Blsp8zc3LynfKqE81z5jtKZPNE+c1mBXA7Epr7dOZ
5z8599KF8vCgrKtfVvsG+L1ZUK1nga11D3CL1Hr2AUg7lqYhy41kvJFr05v9rnUyC2+GLjvOEVNY
bC6plPa98oSgyACiCQk7wF8ngaEauRpTMtsEIRMyDMF3f+K6tMMHuBCFNf/TPizt4kzBhdfNtkwO
us3SzJ3rXaBp6Tt5TM/SfIL1a+IGlPcXBzwoUxlIAgg/stmafBITC4pLOC3CdlmWpyeZ0rEkpeCe
MWlfAYnECBOYMa9E6OZwoeGDwQbXxTb0lXd7VQ/3zX4Qu9t1Lc/CvXHoo7BXzbCxNgGO4Et2vGi4
7KjI+Q6AL6ycN6sAd6TKWWNI1oiEmtoYvtDUFcQVvrk8s5v68YOZCgxQYsp9S1EVOP4Xt38ESp8U
HwJUTSfBIz5qre4GPiJI24b857UwwzYeUC/5l2lR1Wu77ZkJ9KNfBuF3220ieSyFrc32AJpCJGfS
VQAA4Jwdb6AjXGKyOHpht+kYWdzq2Y2vi5M5TKfEEeP4kPKw/ej4py6o6jKTmxmclhdDb4HBhNVU
usDdKoEjutE12h7oUmKv+0FyHEHvxJ4d71XBm7qEkoQo6qLvoc9knOXtNgvB1X+2YstGWLlkkNmG
t61FegfFIattMH8AJzk6DpjEniVZB+dWHV9898zPH/EhUoDGg36wevfk0vHDDtOiT7VJoVYMkuny
vVlEpa4KsDxWOE4d8i+fRJuX83BI2uX7Pl8SBSPE7QtgaXeD7cOqCuQvqCAWT1861i5CIF4rsGHY
lU9Yt/29tXG0aIIUfxxIVDBrel+oGfvwBAd3foQ1ySYDulqeA8TEn/GoC5ci2FQn0UEyk/y3Dryg
2RZNlI3rmoK0ZE7GUlBHq+DXBXu7PCjm9Wwx7PaLaBqpNEpDQpkfj34hOYivW/Nbpt9AMog5MS0U
LAOlPkThxObDOQTcxHJk8J6N3EoG3HADDRej67hU/qxzIDydXJBjkWbxSq1stjTjFQGA8X5eQkGw
fq0eRcsf0RR7icCA+8R7n7ON7ajaBCqQ+i5d/krwxOMpA+L1Kz/gyYpeQ6Pqb+um+nJt+GQWnlRJ
vqBpV1FpKuzAw7+Y1idxtRQSMqixyc1r43jla0kLM2g4Navymwa1CABisesEB1wFN8Dhvqp9ZxdE
PYlNLOCvAm6/p8mzKreJo82/eN0xpU/qHSZUXoBG0leA3FG7zOHVnqbzlMmo8EkJvx+vg4Q1Dd0r
N5EMXqt2M8+o5d6R61ItMzr+cyNWL/K5SBXf4o/5KML82KBArBmRrROtwsmktgIHRqr0vQfwff3a
VuIa+Ugpt2XACj+2GJkr+HwS5uq9tNpHO3eZfsAqk1Z2RAVoOaVjf20Dm+nUSr4aYRrmPEhZ0eFz
FnmekzDdGdm8ek0yOiPbMnadpxU0Nr+e/rUUGVYPDoE6YCgqfhphyIUNDwDOFisNkZhOJMldfCTn
BMcmNyXcz7F+zQ3aFRfCCa4U3L30o6u7coED8ezxBYAxuX7TqXpj9TNPCvAThSVxLnPWa0mjI55w
0c2EgqhxgUuKvjhkJDvUl+pgNBbv6z1P/SCubpme27SMHBsjeHuh58Pvv8CZI4zn3MorqHh4eawk
3oP+vrPrcxe5yaQJBLFmDUQ3jfG9Ho2F5t2tvGUErm5M7D5uMcySkwl0e7Pb6x1QnU0FT7ien5k2
/E1zpS3mmf1mBogdiK5FA8wOYaGjj+dQRP5EQSx6M9smU2qW6PbT482emuskDFMs6I4A37NdOPin
+Jdc/xWscesg+ldsiVBQEB2jTWujvD8BhgPHvI1ZULE/TzlfvbOMpOhb1JN/36i6uQIcu6mCCf5l
VlmARwOkqV7QrgjaNWrX41/C/f+E7SkXW1cLFKOyA1+dNL+2Ot+hjiBgMilFQjgov65hmR2Ifxqw
dIQw+janraxShOWZgxdxAhgO96GnYoEN9CCZf2tfI4cxwUCYbGYuaZ39ABxGmrIBEbZbBG/Kfdkp
LSww8tjYUjehOdl13u02YTs4AeqSEd2XVYFJG2mmd2/7Td/gLlhdR2gSnwQehDy+SIJOiAySQB63
/jfknRbOCaFY0kOsijMVAjefjJ/DBQuGsWS3plO4ylTWje/QaSoxhFSddM0IWjwCHMMfwNviw/7A
+qaHaOkabKUz//3SMM16bOU+x18W9dSn0MtcEkBkuHGppU+mwk5WUcx6PSb6ttFPer6VFJlfxVV8
A37EDHJ4nuEMY9b7+yMlVF/JhTqEwnZhZdJXPWKlBm6H+Li3kdOjgFAuBaF2wMaBiQ9amUZtCZ/q
LWaIP4WaMDJvwEUFvSlKPhH2KxhoFRsGycT/i4pT7TmkYRyI+/bdXqM29uKWcCGj4zz56qqYUqmY
WsjkjA3gFtQgZTLjURN9lf0vy9bK2cpR+Q7X5NVYQBpVOziyYm3byDGTkq4yHVSD1gV0yBpowq2B
zh9KCsm207UtOtrZYYmzKjmL1hilJ2trkZhwGjF3pJnsGzOjLTPNVLcptGACfUV4pzxAN2jf8yjF
glxuR5IsZyyLr08PxXks7Y3qb3lC5HTP3opU4ojBvXAmc1IJ8t06cBTIfHyn7J/RfnqFcwPiiFd8
6wm/GI9Z5xBJUPqlZe+mRbTRrlTYjk3vXUg/Iw8NwxsXNJ8C3u1GF1JnWF5l90eZ9yXkSs7xx2J4
R0adj3EYev/uo/IVL5Kp+Zq0QOM2H8rBY5GQglRjb7NojtSfsd2o7nEmpoV3GCXcaASZ1w3lauK/
24BNaYdeiQSvqh+Hk1tGy+hNsx0gMF5XE6uANfJzGHuG2PBBP5QixQGItFBRhCLX0B0kB5eS1e74
p8zDpTg6yI8MBeHPK4gIlTxwUMcyejJL+UBY0Jti3npE2PkQqWOMO7zzh22d5Vq+kVuePpaR9lO+
u8OdvWOpIEwwV08z4xJd+fUpc0wiSRhI8DAuiX+0aIyPOhaVdE9DBgFS/yx5w0jG6MJjv1DKsiqD
MLr14E4DzPyc23l9W5cf4UMsGPv6OStLr5neUMh/Lxq1vGzqS8ycq7zpZTPu2GtUDCz6+RATnSnL
dF6v7TQyWku1/SNDW7bLvEfwRpEwI6P384pbhuEBw7yQqGqbR02QlCvSZPjoM+gBn/h4DH4FWGnw
+D+PxKDhUMneyIz7bB6wQMVd/Mz5XuJontw451p5YRMpHsB9+qNytoXghlBJ8hg4MTPXrzM/9/Zj
PGwFVLx77+mREGstalNpLpHh2vKlfPPmFsDz6kyXsIqMHeAi+tX7et7Jrg+AsvN579GmEF+v1zva
EghEPKh0x7ff9QSbg1u+qdlYyzr1B4kXZw/3r4yVXLuIsyGQtdVzqke2A5fCR8hyOWxyYd4Vd6yk
RZPD5Q0m3HhIhtvfS+yJNjcVT2kGNd5bzhRe6kX3+pVySVuz3txK1GTeVQ2dvyqzzeREztTdwTwd
V4lPI1xRkNyMw5CVonBkwXoduM85NkEuBhCvWys1+MHO3YIOfdL5jVjb+lSE0ntcqkZuNEXoHHDM
tlZynD+1EDAOlKxEWllslfaVpbMa0VkqbhMZ0pDZkafdR6yzq2/S6Faz/rsytS77WMLz2NVoJUgg
pTXHMqzSbhexi2VclKt22/v+WqtG1o0L7voJFAND8Nrj6e8rPCNBWHRaHTzFJGuNmWMNj82BtE5n
Afs6hGLApC8xaJSW3eTw1ATHmmAZ+fnrDA0yxEE4wPHEJxWzG5z0ysoKddpUFPD8LnYiGBOJ6fZM
wqPbzDV4bIzzNu7CZb4nwIVNp9voQemjrbl37E3pBg4M7jskPxZwYmxUDJuDqE9EM/oM/cVjYXGT
ThC9rm8w9ULT1Q2AmLqDZ3ApFRHBP5Etlfnex60b39Z5ptEl63RzVFhMcCnNPKVGyjB1kskohNii
wqs503ncz3W4NJj6ZAmQ4p+DdRP/AdIVjtCQVD3OQBPAFF9OBZ0Vh69Y9YL9guTuDDhhwL9XjYRO
sHBXMk5BqsDNguxEsOVMfYpvKdqcFOioSrLi/wuPKzy4XES7t2IJ2f8Y9z+tijo30+Wsu/bukJm7
R1ZgVbvv6L5SYbbNOyiG0j8JqluIkdLiyyUYxLuu/UXcTTVef4JbdrBOJ5nYWjFlu0SQWmd48QCZ
1eW18P6WhPJOQJ9V4RljAMSIevoYfoqZOPQmgrLNDKVTuuKQk5dteRk3EppfKIv3ptGliaqrV+R6
tA74iz1ZPpsPIzd8PF+h39XhRoeQDas++EomSnh4yjyekeRA9rrSmS62PdN7YEfLG4Mh130UUnTS
rJc4jNQxHp7gQMLZQan4Lnhhq4FXfGxjz3iGD2qWxlHRm7QOXh/vAWixs8o1laEnoIgtzHxzmBy6
AW6jtYghF1IkVAMI1jPOPENsq8pZpKeJFTBYBXRL0FfUYx/sjVhht6UpaX77ZHCDZyW3twJbdseu
RFHxSGN9+Ungmq8AvdgrmTZK12azlE32gl90lQ8GGjoWO+ELjBj2wZyLPyUJlR+4RxcAVIWIHta3
oZ6fwPrAkzlahVHsiMLachD/vMOA+xbQ4Hq5gxzlfJm/fpafU7KlFOf/gskhn5+2pQW0EoLWVsd9
Zu0lJ6hc2RMYCx6CfTVQSFfi7hjbCnLpAMm1J5+SEn0JiZXpoemEb5wgwCz0NFtID9NouaD+iz/s
NftilCPyHolPZ99T6ZiIR/04+nr7qCl8rP4JAAUvtwVMiHqurHJUhrAEjD3Efua1zM8CPWYmzOtp
j2w0rJv/Pah5xCc7VXDo6ILJ4DHvnOoSOOTx3tqdWIkmh2VL4r7x5tjAfvyDpqKvoDDzYutB0rva
E83AedK6y9Y1Gj5KgmAp3Z/imw0Tc+XfNnlolJ+2n0hSyFWHbnVx7VXYMXMAeLVqYOkddDbs9n2t
PyeIEudstbv3Chey349q8MdyEEbwOBNlAmPoLrRFIAngIESFchY53w9+2wqzjHdRs4B3uLrhehlX
eAVEDiveFwOuKIRsvC2CrMskhhB7K2rZW6L4ggrycpzPVAf78sApkvM2pff0nbGXbuV3C14o3WFu
w2Wzh0Fg8khGEqzlf5fYu6mm558imMf7qV1+bn3D2JevoCV/Hc0IBBNZMSmu8HiAhbfZYNZokuTF
/eZIOJGP/SDLms+bGSzpgAT5L9d6FQFJnRFT/iA90XX2wvld3tgII/q0HdZaZqgQemflAE4K0hUp
DnNPzSdbpiX+a8PsHNxquawWFI+r+2c/tsd2jwXvDp9eKlI96eayeX2UnaZ2LXD7NOxOgxVuPkQA
772EjviPoYWn9WkEBqrPehx8ZlY2u2O4XR7a3sJM2t7saPfEI/2E7QX2YQ+okDz5eaLz8uVM2ZyD
sngr71v5FR2yH6DBoC5H4q2ABBo6UZcll1ozwXwTKvsB/NY9LwDMFfrKV/LLm4WCXqkJOOe7V7h5
bWbvNO62lF6QXxeHrRZnel4sGDwwi9IWC2kTi/cpoPPx8HVfgnzDfQ0k4cm2sPTwzS0brxQ4FaIm
ZACejMNDKPGwnKdy+4ooyNPGv6+pfob/RvSDXwc9F94FtRp1/M4kV/fjF+8o5kd70GmWc/NnmfT4
g1qC2I9B8FTwfgy6V3xQSexGbsm98oHO6qIDox9Lh64vgK+xBVPh2KO0VFhDr0Y6Wqi5USsZaxok
M0EB0lfY5L/+xJEG868+zv97NOxIKtMz2V4IYMBrgRlNV4T6yVwQEx+xe5jG0srmdGxukU4IJ0J7
8FyK8ZOUVy5tWZfTy/bD1lhoVEyS+7Q4q5Zs6nQgsmSJSd66WWhp8iaf4RMS1X5SFKLTgFPx4K9h
UIROW9e2TLTJlalO6oGiGKEYgzBAwQcH+NWy3+PuXw44uPMwK2eW+FXCD2Bh8UCPlwhfywYYIQ9v
YBRnwrvcZRT3n548YmNtMA1QaayxI9mXEVivJVaJ49dsLL0AGzzbxPbhPacY+j+DW6kk0YN8z1Ab
QAVclRYFXIqQ/xTJecwyaPSoyyuwUAhjfL/raF/VxHK34B1Yhwk/yOgm3+TpHgaIXvlnJqKw1PxU
4zSnNhGM2fzpIc4XT6o3VGdait9OK1hc/S0hwn0vjx8hamWNDLnuXksXtrmbdVtc02LIm/MEfufR
hZ5fk8s2/RuKDVbkjmet1AsBTcdUVAjdQD+MmfnEQ3SAqPBLBuq0YZYotr11KiRGMbfxx8fpZM+1
BnNsQuSbvsBSVHGHRxmzMEECzl6xxsEYDWg6BOcJUB8P91xnuwKAiBOspNeNd887xWD7G5Bc5x0V
tC62wE69DALFKEJEkqKdk/D92suN937AEhuOyZzVh1y6zd3v2Ikot/1zJ6sLJiCiDRFp8vSgB6bL
NcW6+W4uRS44evK98HkmOo96kCzB10scdmjpFUKZQLSCKUuH6CIkIRL1D7uRo6RuRQWJ+Wwmnrr/
oeGoUIo0iwV4TG2zPTQK2YCQdUZ+8hU6R6e1NpWhDEtdWR/fYfRvXmidh9tHCrYYNE40SEO0OcqD
crupr/aUb7jlCY27yb8pZqcJNFXKpyrw6SQzxnqwHOD7UOnm2XLGFvm4ZKegaz9tcYkRLcWNyP/Q
NSV8YR85ID6gwF9Jr6cKWp9IeeZBE3rPDA3ffnnh8nKjQIIiLApLHxSufbdrfz2pXY2WjSkFlDeR
DU0j+ub2z+8ARwwS3ksnPFIMDHJJfU41o4pfsJ8LeBvmx9GOkmYVGrH9SxP6CECFnejwmDXW38Qn
pbwQckgoVHLEQxd4UAZeHQZCyQ2V0O1dF5opQIXXrps8GFZg8N/ne4afp0qaeYofqWTKthJuyx8h
uDecYu6c2mQucz2P/R/blS13Npo+VMwAxM18RcYHvslyuBuaPEllfEHRmQ5wNgjnkza0oJO9hQpW
BYwDQEuVoCRK98owGdWM3JjihG4hwctcWAw8YyL3qtuvLvPNVvDq5e9qoC1O91+g7g+FEyKnbp9M
5HCiybRLJYh/8jjjKExjzxtSVqjTNUYXp4mSNb8oDrK3YqVkLEE5TkrwPSRp/kqThMrqbv17uYpH
FP0xvm8BxkB4MzCeLdlbwaDWRiavyO3OarSX1//9Cw/fv+uksMKdzjrXdF0Mk7JMwG09/aUbjgZz
Sg6JZ4+fQ1x1r37/sKqecPo3PdueES0/vQJstWQ5wOoO351pv7A/LXQQTP44RHhuEVKRAoTNwLHi
c0Qxu1GIUbzJfyRR/sjnfM4Pw9lUdWDnhQhfREqaLQVCCiR+Asx/pk2T7nJ1Sfys12FhtbJ6K5w7
w/2w5nMLB4lFxQlh5IJ63zVMJoKRZpUgYfl5Mol7lYbW+zfhlu2KAgqIrHqjPr65Dgrns/CBptd/
TKt/rrLcWevQBp/0UIGAG20fhg61t+7iALwPCoItaM+HaR3Y2/ji4D3ehNfEF7ZazZ92T26vVx+6
6PYnWfzqix/qOyU9HAuB++SHxdeSy1ZQhx+h4rI00IRHMrn3vZBihuidkEUihgZMkSPvZHUiqkru
kX7dXHgGrmxhz90jbkzsRJwtKAtEP+QPETq9QwOZIn7NB91D18nhK33tQw3pypMygX0mTf54SbrK
UxhEaefxuUFxhQCOvHAmFzM9si7B+2CmKj/xTAbY/VuKw8JFRTp3Bd/NiN/hsRvS4O01yXxKMR6W
5JnJka/QeYc2H1+jtwGkrxt/xhImq87W2wCMxA0xgY2gPgyDR805kjcbDNTYBRBvPtb35rOsQV6a
85fq/t8Uf6MRRJYDblVS0ShVyQAVpbVC04Zzrf6MxEJSxP5OaSlFldpj64OaFLtuTPHZ7kDdBmRX
F069xUTp6hTmI4NJLeJ518imPFdeDhlzfkJBDsggv7g5pTH4q8OGaKYDWgftVwecDZ1ZzYpKBi38
YoGXEs4EftX6rIVrhPHOoR+nNCCqdPsUkCW1iZLeljStifTPj8lL7tQCTFSpktGEWrboNDrV3tzf
x0oRyk50YRAr9uK4M6u+hjp2DAVveE4J9rJcW+clBCabZVmJeOTgY3zQkU2Cjs9gTOKH1Zey1ERI
kuox87iQD854VELt80AAJ1S4WYQQXBSSU8Zo4crXKKgifGHgUVbtbm56yoSf62SNXDvihTje+c2R
jTgGQ47upkdSeufztdBNLS1eb+YBSk1lhSNQoBJ9JK1BqWZi0I00gcv69WYEAmtIENa4oh+gSYt5
JhFeVHPrYizi0UZ7E205d9JLMtg65Km+sJAJ6NXRNv90gZeO4ukYuC2s/PMCYmjDy//6YkmaX/Rw
QbdsNO5SQPNGkXK8IXynlaS2gwE+9NcH/RM6soe7rnyMODCuUDQWHW60/Kak1nl+q+lvNUweYrh/
jgvyuX++pjSDEnQQzf+oaTk872QrRttNmJi/JhnRtBhbX/UUIGRbQgHQM5thOfWKKB/iA5zH91lA
tUmQ+UzBPYC5RfPoZvZmcI2i/KluVW0pJH9lJzUaYkhvt1kiHuBosLKCfC/GInSL5sjXCoz5qxQB
9aN4S0HiUFyhoHCr/7bRlgOIlu/fAXbF+G5veB+vh/EhBJVkTvXnA/W/RduFak/D1iqgjoppxRPE
kFKqaEDrAcnGDE3lRLPnS6gJoGI6eJSXOo0j/aWVV9wScTJwAair+zKIskqXsao1yrP8RWhoPpWo
6VuNp7r7B/KfYSxHBipLbp5xfMSDrtjc4wDsYkO/2pLR0LFe+Q2SBMnkODtYe3gSafv4j7EVHPZI
dyKOGXL189SnR/DHFeA39Qwn32v9qvTElfRAjETNggkevzONWKGVeaX4riktNtPJ1HNqipKOWXud
QR35MO0gqc7YQreleLi80QJe+xEJu7Uc5ixF3YaIqhnRsRQUFSqdRuhlWVxTJhVQt4Yd6nWalL3S
qquLfnRQswgo9md/2gUJdKgp5SdWRb/VBXWJwgDfN03cVZTJTqK37PBdtFkPu4mja0yes/OGevaE
4mhrildXRfswlodDlgmr6SX3r95xKjasExIE38CdwdEOFWfr5kGoY8aOzVcsABo6LAJcv3IqaUKZ
gow/HZotexTAo+D3A2Ekh0tG5hnqMsXk0GjwTQ++ZjzWnDBy+lPnNjBKfKxKLg2BFpB0ot0nFA0S
4JfwG7J+pnnTDNTbSwgMIQB2cSK6hO58Yrpnik+dEbWGIopBJ4FPUXj/SH3IhorM+SU0ruucHjZ8
Krn06kXkpkfjzF2KnGjSje3pov51x8Zucj4nowPLnecG4n10WWDVVCDNZ1T4T4hgHMsOtpBnoFpK
QkgLQPugkUyHiaZXlVZzCijl1VvrYKsZJXEaqndyHF6NPQol/un8CLjCdrcEOxn83sGbJ87aoeHo
o0Oqd3kWlxqXD5QM/LortEZdxYXkA/vLeurnDemJZ6wjcLJMp4LIeOsJtJeRlQdPTCEOLEr4/tiU
vJodwifcpzZ+G6rX3coX22y3Gu1yyE+f92XY7riOSECRtHgNZZ4jf8ZiDJnpPLEQWchaKIxY/loJ
o1FbwH/TuISZt4cSVF9Ds9rQZ0Y6ROM7BgsX++cC8Uv7PuAGOWIrG6fgNgoUlO6hr1nNZijiTU53
7VzsyZMr3ODjNbtuDbdun6xQWmqtYv8SNxjjlJXN3TEujDHu3M5eGgVq5bPZuclXG8u2Dm4Gc6jL
8mad1IGUpkz0BHL8LzOLknPKTT2PW1UcyV9TqamWAQMkjJlEQiN7HUu2Pln/SIe/qzHpUTXkSF6t
6xEQxbxFiIhqm134ARHWW5r72I4xhoU70BBpZshwJC07FrcauQ31zGfIGIgfIT1JYqlvlZgC53pV
1eA5HqzGuVL6hkN7eJIOy9OUI8O74awq7R5Lc0gllF9genaBqeX78Q+jDfSEnj5EyuYZKhSu4PRB
+0Bvs8txJlGc5GjtKt6R3TdDPlei9IbfCTRvROMhAOQijfFyDM2LeIGbYJbczcLlmIpEUr4mbq6H
3rkoYTq0QKXRqO6fiWz9fqr/0FZJ1W/S49nr0oDf8YfYiyxl5sH66lWI1NmykkflJCWU0KXfwPy6
BjZI2PdddLxoDwAFp+P3lVk3RCcJv9B48mKZ5VAyFywW24iH0cAErIgJnWCYrUbUnwLdAc0LUBvu
uy7fNakzIR6Y/tylrov9s9FhJ+KxVshSBLPrAkH4XMFaD6BVlz6RuCClSypZGzoZDnoLjjFt6+hr
5a3uoIQfPXpK0pRKRd+R76k5gR8yXvHWhLGbu5fpNFLeKYB2+sxH8Zb0uoVzinRSKDqv71fW1FYM
XSX0VdSiWujz3D9QMvMHXvLBXICCJ/AO7mcQP3LNzgQJimiphUvRDmPXlBdxvHaqcYRfByu+oWhF
cNAa9mHCiUiIvw5egKNRcAPlOOqTXEQ166wjGjZZXy0RAg7enrM9kZjjZBpFzng3MJnYi74kXdLL
j6IWv0oTFW/YqqRVgChK2IYJp1N6rn4XrRaQSUI//Ob+hBVh2Yov+RGDapfDbADQl4OVHTQfxAmL
2zaYUFIBX0MLs6PUBZfp5EEwQDGBl5iAXfV8QnwAmeP7AxSqxZOoHEsMta7tW1Ugojl4m4P6yQf2
HquohAuMs23vU7/bJVi4Ke5ztx2yzsTkA36N+c+5CwKMcSBdLX0wkguQU+UwHuQUyLUAk+iPcY5l
5UGzPjBaVYNUTbr+cKkOpsRWuk9UHPff0tULZOI/FcCc9V3zeDTBxim8KYT7Bvn3E47P8r0L6qK1
vVNnYC1j2eR81oGr92UqXEMS287SgtRhT1YWby0dSgcvM69t9KAhw4A0PgScDTJSDeL7tcD225PG
bjf5TAzqQalA1R4R2TqPVg9j3FiAeiZZLqk+yrHa92dbrVkcHq4pxL6vMJMVUlFJiUjlyo1dzBGL
dUYMAyVVUs5MAmM55YOI/ItOLJAVaYnfP/awdmITzbVQOA2iOPb6db+Z/m2c0FCmAV8JOvJrQxKb
XJR0V9GfKXmZpkIJnxfSuVxi6rYQ
`protect end_protected
