`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
IH1F5cif1Pp+GNkJ2YzUUpyT4qtMj1bWmPw5b3/1i9OlITTDNsBA2eqKNG4Nd0qRdEhkRuAQfLS7
cYlNyJFImQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QSQsA/v2ZqhmQWnpnBd1ViAfOagz5g22BwcO2IqBH7LBFWF2zGkLl/o2mmuMHNMARxHHdLe1Tz6s
HE/PqUZD+WmmDXuseymBsO5/5LW9GV1xNz4D2pvw8TKzeUQfhfKvpfW9FtGUm79vVDIUa424nzOM
OtORVYO1TYBNaONeqsU=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
S+xvC1scVcMwrEaSnSGG3Puf/c8VMJBLsc3RrO9ksHQOccpAnBolsYcICrHfOy4vgQAc2Qj61XSR
eUNXANj58ozkixs/ohs5HdyBgX5XCeuIY0HDls8xKkwQDtisBkzQyQl/J0ZmkqQv3cg4oZO4fg8N
JGJ6LAc0ZLAQVTkr8NA=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QBhICjDm3dj4GwQyyS6R1ne7LZ4yoATbZJzcSdERhQEeKddIssgU6NfoRRMPtQxbL8w00wQ07svu
2jU4ACj2d8IqfyZBwZjeUXsaF2Fu90HD0qzNHfp0SMgxUYH3IgX0uvbmlVB8wDKg+/Xk4jKK9+V9
fLgeRkBHzy2vpLR7Hh8FfaKciq8kCPfjAs8/Mn31WlEku0ZhtgmwaIgyNGcbVyyUIhup09MH7DTW
Y3T++zEQoz22L8Q/2xsRZpHm8x6tztaYx2TaR0RHv5OD17kiiia2WyRYS3Xlk17fIBPG3rwpi0FD
Zz6BZlMH9CMTUPLIxWL8dY7TW5Fb8AQcLOqV5A==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JBNEjetAq3iKH52609figUunHzlzSseS4T4OC/MQl6TvkTJDi36sHW+aYpVbfzgEIuoLOlkw7YFm
xp+V7fFTLftU+pQ29+B6IUBzLdoscpHtMuZqjyDqhJByD8B43kKubYMYELVoqm6oX0DYj7M/ilhl
S0eTkrz4uhA6E/yqig6/UbsBegr2Fpy0GSpiNi+VkCcK8KTSUardVxmmjz+frvsjhhjrUwSzPJJ+
Mz/obUn7k+eWCxaaIYlmh66KyavmeOWS8RDEdjhTdr1qkDgXIxWG/YNkOMKUq4u0ziWMXL1iXehQ
VrZ/g+w89ZYN1ROx9+S8e9735Mjq+ZWY2Xpaaw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Kpr2QPClbWnB86r9b4qBHKtyy12DsjtkMaU/1Dh3uesNEl6sHAmj9yO6zOIGFv45GS+XI98Ny0Hw
TKPwhE1ED2KpO3WLs8JG7vdTxZIMS1tqJJctHliH25cJ5ZeqRJNi2QCtL+1ztgcu2wDo1Rt/n7hc
c+3GhDyiyyTb8x/T16DmlMRak5vwpTUkrpjl6emHKEFcFXo7VRao+kTqHNaRdLqedjj+h6wBXmIq
Rwm9sq/A2BaDizRk22ngtlDiKhrzSiRy3StUOqJlrpmih0p2OdkBUP7y4IuCQbK3M1omovdu7dql
0FcOszo6cpuZ8NEa4d/p1Oz7m/BchT25zzMX/A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74224)
`protect data_block
7AYMS++uwa0ZELq5C+C3trLKCtxzAonJSTQhmY3f3TBuF2YXMVhMeMZgcNcyh8fKrD0JTFOXC6iR
hBvDSJQ4ElLFfe2tPeVIv6Dqsfyl3aapH0cucncXRo7agBv7uzQYw0dSzrm89O1dopMfPHKHnqRX
QsZ2C1E4/xs3SwLxpUt6gpu7ypufAF3+uLH0yBkZuzoaNmNel8vLNXQNsQWV1RK/2JCiDj2HPcKf
v0h6Cuw61g/IISZHonE6kjUYIt3cC8AgcwiWVNhSt2f3rIRoDyQSmUv9engXzcTDXoujneh6gIe1
90xI7f7tHHAF05Rvj31yv9l6IeZODBoOF/dFRIuud9/F9fBDrmfsptIuxRII4bUT0CnnSln/eih5
bpxc/TSINcNg+Q7UoF7xmUDjcbTQuimFvynkc8JnDzG5uidZ30f7TMr8BLfqqJEI60wblFNgRtzf
Nl0Ei1053K2Y7HIwZFncQRh/VGFf4cVo2n4glLxGL6K8Cykt//ZMGmB2c8qAtKOINHrtnxqVmeLK
+8d62C8o/MVmDfvqpZOL0M7FuDbcdrMOJ+TOBrZZH5h6booFErXimenQTrdfnbLr3XBueBKoNYI4
/v7x8P79P6zUQjrqhCin6hzX7jacYHSsHiB9BKgIaOrYDepEDspglGy70WfpjGGjhPm7LuqBp0gM
iM8xWaRE4QHiQB2xg6ohLnUMuCW4SCO/k9m4zq9SXQkJfA9SRAO/DHjBEEg/9yzm9tzzTFDNcCaK
qUw8eFYbcgLGZZQyQB4TpEw8YGj7rLug8BiBRJenpm1VbeXZVkyoPQNnSNjXr3nFeRx1szowB3qn
ouqBrphTUiazC3wh4Kg80aO/YDbIJmBUW2D8iPLOS5EZndKY6pu5ITvFNDc1F38GdHHRmp31LXhU
8sw2sV9pKd20uQiCJfE5S42fCZgiWL24zVSF3Qsx3sLDXO2HQBRgMs/RDwSCPKAAKUvIfsytpKuL
sMJs7A8Ve7vuW2+N/lknk1EfP3xcXM3L0ZJNpFXpEuJY80yAwERIASao2l23Az/e5XRd4GkqN+kE
0m2l6bSjc4vkrqDRSEbwHDJEqgNabbyllvIzXkBbuJuPz0/0Xmm5TIvVDqP0eKHhi7wN93F79o1j
SSG1qY4tGdhvHuwDX8fNLXFEZ7L5lJSmzunki7a26bI2OMU32u8KZ4TDdSopjKl6q8Hg2KbuV/KN
DeRHjsFMU3v3S622zchG1nbTAI6hrmepxSTrK5siHxosBiyVm6OkUfVyEzFd4VlZ/wtyX6i2tWYj
r+CDCjlj1kJ3xgjWWX3Php/JtWzYbMaP9XgLtyHBkcdWiVyLJOOZdXPbvxxP2I2ulSCUUHfER5Ew
wmaIP1DBVzUiUj4nKLOU53GYzb6e3qTWF7hygpi0pzC+NzDdTNnnEoILhTO8zz2wOaEm9q+jnx3v
5ZVOthaK/hXDNQ15I1J+PDM6pM6zJ2SbGog9phNCXQANiArOBpuVH5HV42/YQ6fSu9btzESkahWG
/u/U0oEP2ZsQROhqjgbGPNpFxaKu8siMqn2/ZEP3w8j0W4KpW7p6r+NB0E3evYRdFCIhT7KZjbuh
sKs71UFyLXSUPJln+3iyRWK4FFiI1N8Re89hRcIJQozuxa5eKYTqQ7Qf+v3TQ2DZWaRw1+vxhtk6
Ok9oNaSy1m3oCtNoTrHYaBLjn9KwCBRriCiAeuRDeHvxO4zTIf1AQYXyuB/lRlJU9fWjdPlTnUkq
b5sE4ojSYFyAVYDL/Vue5Me6tgrjv7zX52TMinbz9dGaAzvwMlBswQwODcSLn8EHR8g/JjoFKHAC
HWOhjoFTTkU4cUGZE3++G5WU9Ko0Swbyi2pbSLydloXMwTgHxFssjgaiPD8gK275j8dl3Fu8DGEw
dEji88429x1IKH6qQYT3VBGf+FG7EJdyKsyExejTrH7Z5HSCueX7UvtfId1c8qmAYuQfQbH6TYsG
Lj0L/MydYNgPGxkWe0rOyutWYZqMWhZuwPJouSJCrPD/N64CpnD6JHaGM12m/Q0RlFWC6RcSLH5L
fNv9QVZwl7jE/GnOhD76Tyn7egdbAueVjevZTr3DIVlia9HWdN6UxHn9vslksGCzlq4uhEmiCoDZ
Ai37vLkv8jtYHhbo2njd/fuN+xMj90d1GnhAyA+sIqDjdHGDnvv6dZpbWz5zn5paPDr+jvhqdW7l
/xIdq0HlADwYi+eHN3SrjGU2mjC0OIkEFEOBAx+VCNrprmnlNqelynQL6+WEAqMR8/Bp1EzIl4NZ
jHfvMM3ZfdHY6cvmHqWOa2ppZyMPpcC/t+yq3ngIY/Q3uk0a/BF4DFUZskjGBjwCFA6YMflWv0GJ
H/ksJHOD+oEfD5eNG/kBnx7X8HD9+k9uyEChIplr27OYqaScSFlclduaA/u+L6QS+aAbQBjD+mXs
Fk0CFGl+Dqjl1HqIk/QzsZtaFD1hq1v8MPvNNbhpQBwFHW+8F2KBflAeHVjAGA3B7HRFjqBARQKq
RVhhTyjxdvBVvyHKFWJF6bjWb27SE/QYh382a7e4LsApu3UFJ2wyHhthzslzJ6P6Xp6qY6vOcL5D
S6+vLG8VmmwKUGiu8/YfI4xgieHBuarDPF/Tj5NdipbGQLkCTY20Uu5kvZSpjYYYbG4gbdrWyBwV
pGghMSwoIEWl7L9shj9eAduhkxnFokNw+GzDVr9sGdYNAM2OYgLj9UJHljQnWZ+ujlX3HMbe0pvm
O0B6ATyZn6jY+po2m/hs/I+D35fRmz01bgnum4t/G/HqkVp9F1gHvs17w6DILrQA4XaKIKUks/DS
eF8fOs2ZEdfHSiWYGhqT6GHBr8x6///ucMfaOLVgmsIJ3n0WRqKV70WKUiOJ5cbCsP9uy55QHIL0
CHrH9TzfPqeOIbuqBOJD4qHy9GMuaMvE29cBISmwOTi7bkRo/cuaGcpfq8VHzxR0ECjm1ToBCKuC
umRx4eOSAY2e/hrSCX+r46+OuYVpqY07gzHavDOD8ufeHvqG1ajzfrHmBC+/x23n0K28Vm7w9DA4
ni+krcnYdc5FZkSIndn/3h1b3LiDvncJ1dwK6DfxmjgBInHefI2v71d7Jnw1ebh7KlYfj6/i+1hs
OBMBmOmyYLUUpHObztoWqqFBUYHuxNPyjbbV6Gw2RarIIbD/vpdJEd9q/NJk9xpQYE6oKwjr+2BE
fSdjX6nRCkGKw7VEUfeha4ljq1CYWRQ+I6KtqRXVcyWNV8FKKaKRh6auyi0AJDoc0/m2BfZ65UlF
mABwzv32D8rZ9ZIfMajZQFRVdF5pkOHaC84c5JMUHTgryZonvm6Le7i6XQH0UX6jo8v47qUv9c/s
txkr14KxOkgkyGE0QyfZWvSEhO8ncf7/PFMIJnTbZIEJgOQ29xmAix4o6N5kuEOC0z9HbFhngER7
QI019Sz3GsZDOT/SK/bD3mwCUULbJzBrOKckd2qgaK5v/FJRwFBIVSkERavqIFmnT/SO+MwXigD8
mQR+mADEfohdMdFNZvqGVYd9JmaMrxSML6GbtagrV+AtkygvOTGPK8HuHw/dWlvkJhx8mZfIpfiR
0fMpzdL+2RC7/BuDQrSrG7tqtIHFfSAjR9k5rbbNqdEBhIMVjZCQl3j16SHPXjQhxc0UFUyhCcfY
ZIaq+k9E/MoXx88hXatbNG+4K2+iOR2AKcIra7XZLSy8r/w6heMQFlX4fHu9ym0B660GnkjAkuVy
l7lDkQ2Eac9ITFi1Tu8VucM9dXschfVjiSXaScky75HzNOWvZtbKJZgivLEdCOdIfwasVfe+auBy
ESUmczrCPeBp0ytRYC4+lT9tPkngbgkQMGDTStfylQ4qo4JMFbG7c0CaxdbId3rJFeP1x2ucro9Z
rslSjyxVsM5m8UjlAB8KROhSqPbGAFik6FxvpEv6QjELKVGdpp7jLnkm75SJtezR0vY1bi1sBZCq
WVzJ0Yn5ulDuD2fUs6nqF/GKyCmVn1M9PNMFKE+z2GiuEOHWrYq8sUyapOOvrGweDeeP9tNSGLwf
vpJgyY7UHbYlagy9S2UIkinVsPpddmUw+SfxoWLfhriHjAyuQyXEp6ndkZ5ZhPi9VQPCjODZtbHG
ypOXXMDrxFpcRIVftVeIXf1sFn8CelYYHCWGCsh5Gjwb2P+sypTq2v8Rx5nh6tQ9dmaUwXRE1dCl
9gxQxH5wMPp29jCumUcE178YV/L8O4FkQyrqTiIiuNqVbiut06wYy2pdXR9XEaY+jzGk2a6hHVw5
cYnrY61imdydaJJUR628s/juIh9/MTnWztFBPYEuU8pvOGqveGd9hymjobAiXRUbksbFSIqo8CS8
d1gX0jKwqnCrdZ+lWbjZrdh4vzzvejl5WmSjX/ENas81iyxgt/IUNUf6gp1EJ7yjp0aQRmPS4y84
io3hZH2rjX7oOJROZoFV6w5DT0ncDenLrRy8u2EdnmRLW+Ghkaz//5K8NxfO9QmGu35Ra0Utfeko
c1gmUeabg50Co9c8R5eA8t7Dhg7OwoRGhgmyRl6puqtRxOUmJ7rlaCJrngajsqJ7EG/N6ksLN8uT
yCkGbI7kyLQfQ/gfSSMD66c2FXhDP/aSFCQK+gIeU+1u8iQiV1pbVGasOFECeR3DJHunZj199K/7
aRagGjcWDRtIF0JncT8FI3yIZ0bE3+Gv7NuPpiSRcMA68ItxApbuVNk3TNFYv4XPBRXBAkIbPLUE
+jQRcVuhprI1LK7DZg6UDEev+ZdDal1PC5GfGUnIUyE8oQbgKKGsxBc6+JZoPYS6VVu8OFNZveEj
wjjpLtOr6BlzZ3Q9Rg+P2ZJRRc2TRDWC4p6jhcp8DnlIoMKVLAkcV9cecQw06kmiaxThDnMbX70X
P8m+oMa/ZJxiJMg2iquT+Y6Pth3+qKLvAE7JYrq05gGN9+jYl/u+a/XRvtQYQD+Mt67O7AnApjkY
NvpFBTBX7v9MmMfNAIO3jGS6CzOT1jS9SIdpnwCa9rJ6sdD2/T7KfXv9ZXnEL/cp10ckHXoZ7n4T
kC7PCD0Elzocw7rHQL/YGt65pH8FwsehlL5QiwBjweXbRrI3BrcHgui59gIgx9G5b/Nu759ZQzE/
T4GiFmOj5LLhezwjCZU+IkrDt3u7mAJDBvx7v40uwK5j8qE/Q4nhZ2K5yLUXlRqrM1Ef6duBJx5R
af7ODEo6fbq02vwiVFW46wYtFVJpJSL2W5NVhDsaPd/pXopo7iejspoy+yLneeGGduTD49AIqZKy
DvJQptleRspeGTLMK8JeTAdIjJ6J75S2zR8mGAUXy+plB4IqTgzz4/x5Q7mBhc0AJs8C2HyR7BWt
nqg+vv5+aYvkaufaVjQX63WyAmhVg3xhLDW5BzZHGt0X6CDJpThwrXp7Jqzg9yqag72aaZ4Qo3HC
XxiY+/LK5yxq77+7soJ9VpsKa4nr6CbMfmAHEKKjEPRVgg8Nb5vxv2PmlVIbovuJviP1XLcxHXZ4
Z3B4gHJtO2s1b4sVhHn7r6A33q/dnWPD2FemxS0OQEqf0zWizlWG+wcJip1QyJnklJbX155VyedG
Oa9rGdpRxpngyfmu24ZXW1OUsRjgp81mtu0+BNqvcp+qVeCarE3ZrZgaUM+1R/FCiWilOoL7lj3u
vb75bdMbLEb0D/G+1zy8b/9NY41dTYnwpsKnx1NDVC5X7RcKAtA2XbPaO2ixBSzcMuobyvKUV83b
dMEmMbPJyqpLDC54dWOMufTy4yrEnh495l21MEPEIhwteC7q6cYvWTQMLae8lUP/Lv6N3w0cfaU3
hK1RNm9lRc7WQrgpIMxO4OQAFhZ/biM6VbK8I1iGTwMiLlBO5Iy300gnSC3KbaM8I8aaKiNSACky
GcEorT8c8v5FzyuxS3n1pvguMHf4J4SLP0sDWInaLALxddHjZYcP4g2qBgQbPdrSOtjdS8Zc+cuC
u1lxtHQXT/BHpJyvL6CCpFGTrryTAzJklRDwwHRLHqYji+GIfn0VfYvd8JInHdkpQtSmp1gcXY+Z
FYr+op31G1xG4sBWvzGBk8wP52ClERhJ6L3by2iB9pMGpjJgNULZOMu8EEJKCQGSqcPH5N2jphXR
UQOLpTsKhOYbuXOtHFvxfOKZzk2KYyO6hBm5VQyIQ2TAvGFzHSl0v6jGmaLM9AuWOgz5x7LGxAgb
3hF56QAYUncofx1lhLHTbXcqMaI+AeJwKe4sU9Vsdn7/elsN1ZaZ83iuXHeZOK9VLxYBii06JRTS
8vvqKgiky8rj4aZ9ql3lQ6nElrf2emeF/hVn/Sl4j7aMmMog7kkT0mU5C7cpHpgwKcFxgfw6fKYM
vwCU7Y5/fmdVZ141klrB7y1vkdPP970/Q2A1DsGXXnpX31fUdwOI5J8UCfUyC/kQA81IXVRFr4d9
3KCwuaxEaxdTGesgP1y4UcmIAO5hIRPV3xMdwqfpu1BY/0hsVa6erU3qBfACaIElT1ENxDg8nmU4
oyRfpGot3xYOp4jVxExuNv3HmayV6dhl9A/IPgFGsBEwOIVWuc7np5bpsKmMZLjlqY9xnBLIVHVj
rIzdI2q7lCT0Lwf0jWNbQVk7RdbePqpGsHBEgugidT4mQSTwT86bjqa9h3YKGxN29ihAZL6CK1j7
aGo3XA2PMLmGnQ5zEQ948fdN71WFBNj3egKqnum+sqR2isxLohAxKQpAIJX87X569AwPGF5siepW
nO3Dj0Sa4IQJBSO6YGDOL1MWXI959s4OwdBQ86/QEmJ51b1Mh79yT34cT7aTpxH+2PmvTrYtKd/g
0Yg7Bc2xThLy7bd5bHQujtxg13tW9C6k9xTz5oNJkFul4ilTxiLqsjoB3cyxsoJru3SmRtjhThZm
tzuRdShVykoVX3TXlxJXFe1z2EnYms4bCw4JAFQd/tiVujDcMltBLvqrNCs+VPTlOcwB0Xdu6ND4
7Q8LQ/YQgC1OChf/qxERFK/jKloVkiDP3BFaLmiBfCbd7xKbEh9HDKC64gYCzHy8wrDQxvccvSvJ
Kj/1T5rnp++zRyFlXLhySpxnIGm0i3gln3lLKZ39l5sw0wgRtppAVp+3RaHiknDuuiOCJBak/31j
4mc4Icxu5T3Kcwrotqg4iBL+jSwOVfZyvIwjvylMoRDgLDa0076JQqfHo4hx1Vhv99niOep7npK6
8xTbkGwgI1DqIeMsUnQSkv7ncb3VTaIR06rC1QwOLkh89WYvQ2mlYoIHWlPIDPtIUZJOOAm764no
kiaMqsDwfKJ55U1BpvsfirOWsZe94rfcXML2zalbU+Z2I7Ej71slXOSoVWlBAtE3GaYt2X805dRu
DmWOFpjg2/HcnVZ4D+A2tH9+g3xKHEKvgSx57ic74cC7KMg7h01p8lcGkwxxYJRBHjTM2srea5qW
3ZBBXczwytEfBybARHhsjyPbbfUi18AHiwqNdu16rz4sJFo5GpsN+9E6H1zzHKFQtGU+VZXQy4wg
q3O1PTnzRlhwDW0pBSyVEovydzw0oHJnVjRKeIbEiOzRI/eN4fYYtcDJ7dG4PDT9kAByfi+IAkq+
a9D7jBhNZGtf9H8J6RZTiJZhKAsfn6xRHdZ/0NEgQj7zhg5FsklxCZcDOQncEZmveHV1oZndZMRz
r6qw304LYvXYOit8iV4yJc7UPW47AKkp7g8VjNmIh8HiZzYsKYZ53JaKL/Ouih208vScKKr0kRqz
wtEgwiPDOf/mJyUcPETwbEJ8tYtHa4UnFEC5rJKcXB7MpdDSmkWU9OmAiyUv4B9suYIpvfXmDGFQ
Tp7T4AmQgHjUC5I4675d+nYw7s8nE7MsSamq3NC38CT9KZFL1s1VGMWAAlg607Ipjcy9IWFrb9dX
3rqnlAZRtLxCXm6b/qbTzkUqqH/gJgk5M8KI/Y8HU8VHetqvHYqgfzF473mfbpqh3PRbSnIdbSlx
nAk4jPhEnAsnFZymv3C6mNcnzcrKAr+JAtb7VHMk4dNxEDEHtPEy4+nEh+YG+Wqufoin3nS4gf0I
qk7PCszaSj2p4A80GaQC4vBGRp5VvEINmOoaKJAA5NRuF3dnNfxL3ukHDR+np5Wlhpvqft+TtcjN
BRyT2BX8UpSTBUhjDTsTgbP5mZ4p1GqS4dUz9afF8MeHAxC0Za9FzrjTEZPr52KXYN/Ii/sZcF3V
i4KpU96ulA/MOw3S05WvCeXx3g52864MBitOrkZZb9CamjSMZfQBD9gbeQZvOp36i3E26fhUe/Z4
JPOwSlQPsGTnrjXsZfPCiAlcQv43f4HZ+xSDH9l01hlcQVof3FVF+EAmmbYJ8htCZoU5I06GteqN
i70oMl6adPLcUrxwBjFZddAYAgX2Sips2mh0A+biCUJMaTEjKWH3McLrsd9SsWUsMPodzp8vhVmn
oOMRskeCu7D8jUrlpYMQwD49gTN15G45/Jmc8tspAkcUTeKDxnnimnDIZtFr9ZBZdZnDi2tsbyhw
hXCvL8/5uaeCRf8nOMaisgjvF/Jq48El/55KaX2DpvmfGCA+eaV5bCvMD5DB1+rv3A7WpxalxWT+
FtuQbLSMoRCbiJqKF/DoSSaT3coCNVBQwS7Cl3rxT9UzR3vesO5anSY9x/2YYJhmyyNeqxnsp7w8
AmgPV9/CDIYHrrXS4RitAYaB7C8C+djcfKdWgMvGrtE2+H7ahdaemxs82Bg92pdHvxxeJ6nSGqS1
4W+e83h1PbiXzqx2UA5ep43VjG0E9D3XvjxDPAVC3s835PJzSZtDnwMNkWryXCmWL8QXM4bflM32
/e8k44XND7rbIHhVNUEEy9NuN3gckmbPgOaf3JiHVcims00p03e1k4xi6EDYRVx1XysiFQJ0PFCf
yZ+pwe+HYa/eU+B4sO//aXzISr+Fg823C5bBdGPe8o8Wga2l+x0Mc+CjDwUDZ6RhydNiw9jOcw7m
rZF9MNzwXgWdtuyvjQ0QWK6da1H57uNmrbuJQJyVs5ac2cgmmuYsik6eY8l4iABKdrfV8D7SUQuV
E/s1jWmfapowutcNwkMWamVGBHbi4WTYQJ9MhPm9FQgQnddjblGjNTkJIIBD+f4E5zVP6MDtRpo4
oytivXKWeSom4psNGzt/+5B82dpTOhaeNtg73/WHVq2KmFKzbs6YOVmJOjL7vBeO5M0RZA4ZU4UU
17D/Gm2Dq4LA4VALpH8Z/YpFvN4okqr/SwwC/UO9R9+RmA1FexJ1Kl9xWVji+5ih95do8UN+Rb72
6akozjjK2uKuUCjzlGL62WRZICiaTRdOPp6OCFCFGxQTnHi6egvtbnbg3BRISOK20hW1UD39lyCx
dE2h4BGFoJwrkjq42h2nL6bJDYf2LZXr31gidl2ePfPUNJoOX0whX9rR404PHv7BFdZ8JWjuCqc3
dR5gEPhdKKVluBtB0Q/SIZl0+5I8LYe0vocnkFOmGR0j/Kney4k0JlgurpJ/03/urAchSJpxLF0Z
FXtI/h0dTC57gtjXga80CKLJr+YlIreMvMgNW0LCR9koFPpWFSuSSFW3yeDy3c5t7cEjGNLAHImx
kWRmC9YHWqeqs26vWcTDkFBWdi/yJT1WBsKRXtVh575HINgVm/K5xb09LT5OMeCDpz/l4J+hXH8R
PfFjDlIpHUiFXuP1xR1va81/q3VhRJBKh2cB73AFfqiwEEaDxqVJzOkvrVnrAYUw5CLoVeTjoiib
zhVzcGfqj1M7kvi5iHyAktNmTntSfmrY7JgPnNXpIP2FE4tFygyhJQs9cslP8xZ9T/X0nxfu3kvU
dvZ6NIbK7Ud1e6Jkg3Ot7+rpAAm5/j46+Nm/uCcuPCsqnPiKp+I0bN4rknRb35aVBWEWDRdhrwiA
iysJKy85fMdgLqY0HsxysKmcsFL46E72qfXlRTpmwnbxclvqgRCbsIuLFJx2UQQl/39R1OkM/Mq5
a61ZUwV7ZekTVcxxMkS4hoKUHu+uXGltQXNjw0eEsUX6OfEAiMKd/LD4lAvd9aMXBAo56irCxwf7
vKTr/uUn8DxfDPlR8YCxa56Q+X/7Xsq83c1jB3tBc8NhmkvAGG0Omr6xiLOuI182o8zoXnXuaJyD
o+yvZqhQ5qugk3GNXqmiIhoeh8ZZYzutn/R99sagl41lZ0OWjqtaRUSd8NzoilAg0a2PiJqa8cE5
FvGJGybClNditFjf4ZIUpG/DztZM1iA8DzjT6CJZnfYDuhCflVmJY9qkmCmX96Cf3xRqMPdTgl1o
iQjTRPaK/ZHMGJ0bSeAMvBDVeP+XoTiIq8gadoS55ZovxI0Lz5kWl19Rd+lAyrHjUr/+bq/nIF3G
TcHwUCazd5vNo26bbY18O2FRr7mbyXI6H28ody1iPkSsz4uujpHbNHu/MWfsGCaRoxjnbb3ptX0l
dzIDnRSf0PrjodLCt1LrrcdaS7rOSp47Buy2kg8PN7KXZ4kIFF0MCGmpUH5WKIYlUC5snNvul332
VU8KAng6Xziuu2+h/oZ2iiOyjMby0YbEseY7FBHp++23UypnxTynvfJqVtFm8B+g1CLCD59o6vQ0
jMgrxxX9+rtxWgLfu+bXRI44CRefkZ76NJC8dL2+Qn4aI5GOfNFUn2QgMIJDtIwCwWQSBeQRYJph
CTWBJ1hXaCGJsQNU9Yf8q7qDfKnKh8DNYvMVP3kiZ1UFq0LK8ikR4+o+99CkxC2gQzYpJxVsdz8v
CAjCW5zimhq+y+LT2KG0M41A2+9zbiUXPNh70JswGLW9a8uTklYzRqVpLYd3G6BG9EiCPi79h6Tc
Qewp69U/7PhWQD5n0QvA11ON3SskU9ZY9/AMHwyx9rfLCCCYg7i24pLvT/AbJmviDJSjIx/x23Zy
GEcdmiEEpgyaq/dB44yBAsb4JEkrYKt8q9xTc7PLtw6PYJD+Y5do6ZyJvjPA94paStvpZ2+NantP
xLGYoCBKt+JEvbKdr2+oSZ1q3wTCXSqYhi2mCbSIcbB3/AwgT+hYNMjpci+aVPt0iZfpRnBs0KSB
tbX/8GXEd4DHjS4XoLaWuV3w20rBfwh1GGPM8u2b3x8QuFykhyzvAiSMmqxr0SWLxRBbODq6HdKO
PUadnJxNQKvQsKLTxDiWvOrAZmdSVeii+WmO2X5uwq5jQL03qki369ugzcs+tzUli5Ll0iOOFB+q
jMNBHP6ULKtHvVfNYN3SNYawvRPKdsWZK0DXueJJ7r94Y1RHyLIF+qj/zY1n5xUqvF36SCihNtQA
uwWH7QJBJDO+aoXvFclQcUSyqgFvRUaMm7NTbIHw9wh2LQGxXrHGIZyRlehSGN6OiGAEMdzxehBn
Yvwgu1WO0UJCjjMppyvUDpTvviOVqg9PLyjsc3C01/OZfFtMMEXN1+gJ32/Zitqyg5BoTAHbqgP1
0vL2unHiAwyyhiQ7tva62kG7GE9PnmrAt8u7dx2ooE1DeXY7cEjRRrX8UTHq1IjhcSvs1JtWHzdm
NuPPuvHXjrSIUZ839esx+g6EijSwgP2t2sqYHSRoxd814hg5vDXYRrdbBZ93A60SYaDekCgdnD31
3lc5/38JDUY0zucNaOJcp2Ejc0s626Gd+Mk+yuhBBqh0gPPHv+1HQi5cV3ZQzkngE4l9VGQ2YYzM
/Sr0T9JYSiBaqcjlALFaoG/JTEgBx9MnNZGNZ6dv4Fsbu5SIEm98Mfobhl8ERCkT3AV9Xxo6AcGf
dpSuLzkb7z05jFFoVZDPA3F3U3XvAhS9Pex92sKftmgsHGX9ICCFUIOhUwGDnjtr3/gkYBC/0ypw
pG11qZ+8w8tgsm6bRwDhK44UzuycoXjR5www4i2b13JOCGv4pRoOU1vE9Wix3NqG8UCUTfJcHCCr
TdXqf8jd6vZeBMmdoO94yuet/5jIa8gLkWlrr/mIOF+4umoCkeWZHI3KLXcVSRovDHy0GD8C35ox
sx6PWCFqVMHigdtk/ogR3frMAIm9DMF8MB9ENmiA4NxUjiOAFnpA2nNCiiuhYcFfRDGyaN73BO2d
9FnLYMI+wlv0mTi7dRXHl7ft74YH+uHi0kF3Nh/4gIIv+OcsFgNhW+7h23X87VhfKXSzNFPMXgBG
5A2oc4ad8WonnbsWNM++f6CfXPVHallBGm+Sqe3uqmMVzueldRklBxLml/5obpAwZ2HKnNJpKmbz
T/zHLeftRNbYxAD7duO94k+7ZnpjeAlLkYgPCRmj4scAwmEFNFmEKx0vFM+Bw5vVc/YQvjk0jFlu
NvCllqXvldze4U6cmLBkuXszPxZyIpAhpB+p6VRodwc9sj2hxYQ7dlVJzsCmGd/UcI659TCRxMuR
uvCAn2fUQW6pwV3aWiXck+RZkJJYIJcV9PcFDYDPXysVlqgQTzO+F3IERBjBUE8KtUqtmL8w7533
NQnOXvudl1xH4RDm5Ch/9IvTX1Eq1zK15lXsutXXR+0ZeJSmAzTuX6rBtMji3HMOH9mp0UrOJADK
dPSgu92QglgRgJmZkmWCy2vhWtTdZ0n9pKwj8+HY7FB8O8NOIBOHErqnQYKjQIOZAtV4Es8+cMEq
93p/nlGM/SxkCt13itwK4GAyXBbQ6rPjVLBiW4tlelfZwdq668dz4BRU7io5lO4yzNhZ+BfYQbKN
eB4a7MFMpipe34KcRGvGyaV7kmfQvjuDQA00h/40qRI1E82EVR5cahq+eA77TsvSuzXdJfLrgpnH
nNakurvbeDGdWG2dtvAfZb9GKgjm0rGR4d1W9tPm8ErfjIYe4LpWbAw0Tj1q6xms+WAB1PRxhdsh
K4tWV31CgUHO0g0Krf5EeNW/4wEBmdU951HzOsLvzHVtiXoZnrxZknc1aHHpW/CbfKRREHljoAu8
/u562u/xfGPE4DGGy6ZQDo4e0D5qmHVRrFbid5WSelcIxjKZwgwY51aPK+ZTt0DRC8SVqus65bBG
LdYW82UTwrHtX1ZmlI1W+97oTRrXAIiIy1+T4orZbcQTXgqWOE8RQ9UdGyaZOz9qQEMYzdytDmAg
ysrG2qRZVgGm2qsf6pSBuX7ZcIXWZJSLmM3yUx3jkDapwwMx0w6zYLgLAYIEF6mPfsZgp5kxB46N
usLtCwMz0ypXL9Ao28l1Jjq/kLhgwEuRbaUBq3YGbDPpixkruvSXLJTARPo3oZhBF8UisqZbdeVE
4KoQg2J5CtgekdYR6B3INY85mk0s+d5nKtpJmScK0aEKYiNCvdCvVMOGX98HzJa5Msfpo03F5xkG
+Y5+wbbVHemKHhaAE7DjK8FkLeYZ4LR96UHpKbxdSh2wSrML2ouNq3U2IdkRKy9e6GfD7Fv3h9Fw
GuSItTby214MpKrki0TJYYWjNfyBLCFP9vGtxzMkl/TXZ81lI9ePY88/upb2mCSzfz3MtDJ9s/kL
fye+y1Monx1mkp+GrYnninT9hihaFlM12oNbMQu4kkovgNs1cFNJ+3dGl2fwh9f5HL0jMl0mp8r4
7YZ0WG2Wj5dffoisFcHk6g/eNCV5hl2g4UFkV2VwQt9CbrNwBmwKkjiv2uYyUpnhVIcIyui7gGdO
QG+xyvNeAZrRpIAPfrfuELSpGPkqQGo6SgnbqENBAxe/QR16u1as5xgvj79bYsC/Zt44RL0ElaNl
NP16RtMKe3SQcV/T7JoXTh2fAe80M5ZIpSM1tqXsEMcXHKt1RRoR9+HXoz96tOrO61AxMwnvuBCj
dJy/twNlsfapWyx3YhLsbMEh9qgjak7WKS1BvHlul+DLuhl4VHM1FP1s6zEwEt5ciySKeYW3U4yw
6r3blxGgToIHBPsMjLQlNJyf3B8njkLz5iy7IN4jcGzMX1Gm2fknFca1W5YtHwa7aiEce7XVWkiB
alAxp+k01tjQQ5N0y7E4PGMt/wJ7r0Z0zdUPXKCv9wDo72esgGOQ0aMvLAz6aQONwovrX+G+zcTc
WooJtpTsYUY41iuZixjN+EA491TJm15AiSbuRNbHGfAgZA/Jhb7s2M8oN0vzD3hYijU2miQa9xZh
aIxpG+LazaDyXO0rtF4NvUrSYXSijKhEyJN0HVLnE9VoPVVD+52Fps+/OhyuusFr2cZzjQ44ElJ+
i03Zjw9bzFQUSLo776eZXsl6odoZG2nNieV0mZRCvrgKzZZCfzQDidb6pCTC5AwE3GF7HvSqScz0
uaBSnPIWTOS0KfECcD0zs8X8qKM5XhcvAE53a3U5gJLa+jaGi+q+Y3i3Ap1NY6NwdJ8dqqmK23ZD
A5qAXwPhcItuKghWPCW+CXj/oSIfO88WphGevAvzkzi7eu73N6QvYs9NeqFBk5CYCLX8oUnTvwPF
D5/xjo9qShPdctNUKHGK+6M0G5OsPHqlsuxlnxKHripuCUkqbxEM9n/n9xFULoRn/Yur1oCkMpvS
Ulbdv+shpErx0vGdDURbDVGUbOo3/P4XrkcKcvLEXcoG8cO0c49aP+F6ohCFSMFR1cwlebqlf9sD
S9poiEDgygODPShOVDUQ4aV9Be/egUEs3Nr9m71a5H6hD02BEcPLhi8yqYsBYB/kTzw8WZ4qNJTp
u51mljQsqj8NEud0ROkv4/HGZou3aldRx+fItsjgUFchttlIni7kt+MmWEXr9jya1BVNr1TRIpke
xBffidaJyRbHyUjeX1xm4oYpb995+kCuiu3dIX4WaV/qxC+UdwmHCjLLfQWoynMvUCN4IwfjWgAt
fCS2eE/zkbPFTvleRiM8WonLQ4weGnRXxy154Xy9bHydhd4JfKAasWTWpwhNoI7CulzlDrO3wpp3
Ti8KjTa4w8khZhD2S30q2HfDU0km32XbgIHy+GdGJSnBs7Usy4jdKTTdHQjr83Amdr5yKNS4nXru
fVwfkdaWOAtli6poTcMqVIebiWYU9jxU1nf7riPzwhXm+LxRMCTF4KodqfK9VPDlSSuEWp0j47iZ
8apja/wcJeFV3D/eCX9Z0yzWQX4sosETJuUZ3F0cZ08PBRaKOfxo3rwoYkdY62oH2BvTYh9zotwQ
hGQJjMZx9cpW/755DKyZ3bGkizzXYL3+EGzrkNACwgowQj1P+8MuPMz5rL+kbEkpMlLpuwIPp/Mv
Q6PB0wdbRQtVYD0YXdg0aO1Dhd/luLktFtCeBWO7nr15LFK6SiWI0VgomJwauMzdiPVWNlar9Mad
J94j5L0BYg9ObtVsNbwmAzfIZ+MtTCQU3aDEL+OUUO+TyYmRuge1UjRNQ+R+KQca/RMvSkYYe/0g
d6+YgFk65rABHfGSrLbYMEGrvBJsW+oYdWT4rmnwLlcpTPKi8gHRhp5pbJJ+6LZZL+woEm4SzeGI
nATZYQ5sHYL5h0bYTow8VuxM8G4kWDI4bipJHY8tIyaneR9PZ3wnWfxvEIGUozGq7aJsK3xkBabP
ETb8kW4zbzrQpaxsFFYBlFAmDR3hrUBtzA3yBL3KpNwYJEOjvwWK8HJiu6+E5LtKN2Oal2EXbtLk
aXwkLLHELlWskkbbSNE8r2m1yHgWLDlOXpEs2HMaEcsdEQb2mgiNAFjXoeu2AR1weWu7TA2HoD3y
Tae0MXFXiIONk2UBv2jsnZ456PprAv9Syl1sHyQM8ufilmbVzntRGK17gGGa5T1OMe7kCpDQ4zpD
yYmhak5otJuPh8CnZZ2phhek939eaRep3cYn2u7huyoUoH2LvrScvWmRIAkhk/Q6UZyhuyvdH29k
FLskGPmvLTuUAzP8J8RebVcx0xQswEKwINYFPo/r5uKpjF6ledmi8MGxs5m6SnxMDqrWdqb4TAN3
fBfrtHQLBajBi2VyMZOeunlg6lyBYTfcjcuNzc47T1tU/NcrmGuzTi/pMYiFU7EEOwW642R+Bm2o
NDk39Oitwfq86kZ2Cxr1Oc8eO04Wl367Gade7Fch29zhSL2PLgQXF0wlV/LuzEQsE5JHx6BTZHqp
uK6wmJeqMolp1sIdhKPb26++CfulCaB8RUQmqTtznEDkmnURdChVqdijN2GcAk3aP7zJuJP/P057
d4KZ0yPl8CD0sRhC+nuonYoZp80RrXOJW9FKK71DLpl5fB7vFPKxdkzH9u+JhQzVq9FvRJJpdsuG
/Qi0EJVA/nFlE/xuWIAbyi0te97qiriPo3hRhX5lezIjGdCuml5OrBOUO4Y1e3FSAO6yoayksb87
UOmESc+ZNIWjcXJOY62/gfZMr+bvfptaDlTwvfvOdsy8I9Fu0n3LMc4Kwhr7/UuOgY6a4Pw5sEZ9
oq61xeU59TIdMO5kP+ZpXuAkb6bLxkFYHi3qCtj8HE2kL6fHasOTDCED6ZwwJOPw/T+K3AvBRNTZ
GOKDtR+ICZF/Hi6S1GxKzAlahpuAvUCbOEjJqq1jpd4Dx3A063DYTawVAq+xlqWVpwoZpxd4YJLN
YvDyi03RHyiWSW/QUT38N/BXUui+qXnmCAlAgrVR4dQAlWcOwb6Elln+bxPGAZ/aWDhgJCZ2YvYd
Au435o5XOcl6Cj3Qggu5RHBPeHFWlkHFSs7YMZ2iU/wqpookXMHHvWqRmvHbbqLa+F8uoSEB5Qis
I3uuA94CCQJ3GT6ea6OvgshSbyV3BSlTQVZrKQ949+FkpWqpTotzP2zMbasYgpongSNPTQS/E0L4
4ayHsdIsDtJRNFh+kFpMoj7rAAGIR/t5HRe8gOT6h1HbkKnL6Ls1NCPPAilaGq82nBFqcFjc8RQs
Z+otMn1p6fuJL3oKe92M8ohw+hDG+1fsQ8j1503iSCibyDnStQF9gwbk1hnZdOHU7R/RG5KkspGq
2Avs3vnXN9316T3Fg2hZ9vJxf7nF/muyFP0Uv0F1mSkTDnmmgALoCIPzXGXEbNRuWbCOFtnKxfI2
6Jx7MzkjxXte5w6PM1rOmBAdzPNMGT5wVXZ1lbW9njm+YiqpfghoTbVF91unYQum7JpLDYGht40O
51jKsuJwRuCI3Q7kCZnPnKs++VfTwo0j7mYCr709PaBUkBRAtr6LXrfR0JEmVXyYR1a8vZKhoRIc
qyvrMrg62peFwvLJAVi/Lp17Dc79sTwyZCWj2qGLal1VjqrHyvFR46dLJ108ii4WfX8/QbeU7ttD
20NyeiMvalYBqkMfKRvrzOtCiDEBSlFotpIMW2wYwXDhFRFdm+yEn3oIDczH7f+VLxBh6FwNTggr
+gSjeTUJwNH14YYkmR5zQ/YINRwLQXLq+042bmajaO98bvbDBa6zvK80q9ScbeSl/OFGiO0JxJgU
FgSkImSiNbQzNNc0cBi0Nr1iauSW8aj9PLIuBNki/ybxU/q4p5pNy9UrvN+gmCq5Q3h8on2VJ1DQ
FRPIqG3/C8yS21KPd5x6a37kbFHjTRzxC1aGoFFqwpehuEbDxxgJfUiXvUJceoIzt5sfmS6H4W9G
fpnbO1dCHneFabf3p0kG4Tk90bmpR1pbo4uWYOMgLV7LSF8Bod7+0+8SRCd8w7+NJ7wtUxArltsT
nmT1FTM5RDPMljEJ35hi7lgPIwPGzeP8QSCicV6OZtOLQHxdfj7nxkjzxQTm2BaLH2cfPLrwV8tn
uK16gMGaEapeATbVEtytn4BG1/bN5vf96dg7BTPhT5gg/RQRRSMykV0aqFT9LVz/ShH7z6/VDLu/
btUqB+3Yo0ygqzQMbdGW4oT+isoE4Kk2SxS92MiTKT1rv6/USbuCQdFjQROOHp+PtW5VtvXAo36c
zzpdGZzt4OzVzr1qbZ/EPU3J2H0/ep/96Z8FKxcNit/j0cYG5k3nKq9rSO0xyN/c1KKx8aA4F+wi
/hCOfUps0Og8m/2lRtGZiHoLg4OjnRwrsEn9smUt8UtDljel5FWEsioBRVrfxJZ8EcX5+x///KYQ
U24rBnRUDfrPL7N/q9AQ/6kMUoQ5U31g/pSt27b5FQAZIW8CgDVnsDUK2fck3jZIGmx+obyTnKSg
DNk9NfEIWN7VQlp5vqvSPPGULScd+TGeC5LgVh+lyuqekmCr83u7GkPBW8NStO37QoCE9S6oUr2t
v46tp0bXcKq7rrSm2hoCjyUSRHlYIOB+8dgHy6TQkNhmCxKIWOmk1cu1xR91rpIMBRhHDryFcuND
WCrVPCk2FOd9wgFfqfuQT4jCCTFUE2fbBOQLpdONT3ekT7QjtLgpQqzhaw8oy+azLDrj7AKoT3O4
N0N04r7s2anE4kdV17alzldH4z9mPOnSmc2Hpxj2DXK7x5u/KsLwGjZaE04EGnFhbZwuYjyR1IQM
yDHnZkCBeHFMEvIVNCbdJ4E7ECdTpT4S7iiPXXz76Of7uWr4z/kmNdE2GleJh7lEIM4rqNAuKTik
I5Iy1X9kzKckPJ2hgGjEdyW6D5LTdg5ekK/0r458eEeDVqZnUFgxRZzJKevegKoWQo60K2LhOsRR
pi1NOkpKkC91SFBbhtUH9GBZJpd31tTDST1OdtAh/q6bZLasxP9rEBLm8zAMxp3BvqJ3YRjj+T1j
QMZ210bpq3pjokaBgQmeWVi0yPYSg2xTlwJOgWitNeUeiQHp/zAeCEXOS+ecscDMBTXI9/UbgGFW
AsQiUYVjT6v9Yznf8sqcJGPzJ6g9LAKfa5wnE3wCWjwjSiqk3Z2WalqWYMLofSTFvz/vrHWp7ZlT
qHSUpU/neoh4JXdhBic+c1RtXVHNyEVtWgrNZYyp6wywbeFDrzW9IhKj0NC6iEE865qE8wlvpUyM
29exsHcwH059RfXub178UNA56l+BH8FhRQ+r7TZFcKa3b6YkELrsBDmV9rORDgTgLOKO61ZVdWYO
uqRiMCnaqMQBcQmYYIo5QX7LJDwHb9nbFoHh1J3CciQXZrwtfwqfNVsg2G4DipiKoz3vjeNm55GE
xFekNQ8LhZHjwFhsrot7MLh8eg0sMT7o9wqzgMOnoTRevOZNTkn+rNWSI56R/Wg6eK5uIaa8pxZ7
1yhiSWXdt+6TClCXUDx6QXSDl4Sj0dRTI2vRxGEQnYD2DZRLbYPNMCk2rDQIbgZ1bx5N5Ik1gnCe
q27flhu3+m3fiLReSHKnwRtZuF7OUmGiwHVTySR5CXlA/1eNnv5AskwtHNakmwhPdKeeKgclZdFY
HtXq341jUm8oVuGg6OtpBwJPNReatleYGi6vTWsMY1j+d6Y8HhyERSijjogdJ2mcN4j8uH0+WevW
VyxTG2Hve0ceH92zxx06Rom4VMJ9e0fbLqaTKvddEkalikZuOIbEE2wQLol8SjnhfEAhgIlomg2o
0nr3zqOjxsPaPnQMIoj72kVVWO+7++9oSTouNN6x8uD9tsb0BEfaYpiS230Y1hUr0v/A3bK4uvqy
GV2B2XAcRcaZR9w1ySSrGyi7iPyITZFSw2ODck2qSBxlrT2cjM1u7lnJys97D4rhH07rG9M8FHQ+
3qPhTjyjY39XrF0jhNuS2vKGF8MPMbiYAwiENBC14zeksaLqkOBs21QCAM7OCRTErEZKh9peOCGg
X7+fbRqmVu+ZhWRWKSND9QB9zYEE3A+d7RNceHO9nspDNiu03og2xlSb3i+gCTV6zI5ghTq5Upq5
Vs+lAKuViR8s0IfCQ8q1DyMlm7ZaJ/mWM8oJ/ceItdBomrWkSUPNn9Gjo/KN5lXSUToPf2jJ9+Uh
0GPqsObv5cWtPgH59jVJk7/XRQaGOX/A+LpJOrzl+dDp1rRtF1SdoqyZfhfap07Jg1yFB0nz50sI
xy+ofYLJErP9o+KDMnAHqBpmCLm4zw8X3dDRgqvzG2hZ9FatNhOMIBfkaNv5nbO1Kmmd+m3tjfSw
qHbA0+UVxLxXscs0UXw0qW6uwAqPm1+uJr3baKJCEc5fB7+2EKsv9qeWUYinitg0w5/hH2NFPEPm
TmQ20BoBf+00csV8bsBlqmlrXaS64M23XobD7ZVqLSO72d0oRweIpRzgH0pEhcMguih3uqi8PprS
MxJsU+fT0cfbKLlG9QTHCuHqYGX3u8O7mBNY/9wDXKlxDQ4D1lKr/YNZgQj/Vu3WC173hFkTbk5J
3vOeLsylSZZnt3CPpae4MaKIEg485VKwafRMOBdI/8V4q16BmIRgeEQq435H3uEoNNpzlwLu7x1+
5/gIsermPlZ6wHzsr5TtwFHhkf1r3fCbDxqXX7QJZin3rlcQeHNPJFMA7M/oV1L/weDq/hlzCxPc
kKmqR615SD6qklX0VZYlaH8G7h2SYOOfJTAYen4Uo67c1Wp6OtohDImbC6C9s5suBO9lTxQv52Th
vHhyjQvgtobCWLm48hpCP1AfV58hdc/muiyIZMglVX27bUvadBLLGa8ogElx3+qBCFCAty2BxjbV
UX41dMup491+lpLl3EuB95v+ekylypAby0Ps+dRxMsmsv3suvVivGVmauT6zCE2w9BxOzCme/pGF
HKOWhv/7Traxb6/L1G0SsrXaYOrEuKXuBCsQ8aSv66u1NRcqbSSs1bgXZ9vqU3MILoPxl373PRdF
pJC4wM/KvylVfA3roitFWgLyX4miiV8ZjkP6lC1DKt2wUNtN0MJAxBN1k7kdl5Kbuj5mxRBZcbaa
rC2lhG3Ta4kbK+tPq51xxiu64itcTPAbjKLBCFGaTTkeFY9WOXeFR12g+HcSsDrH0OVtR3MjrFlb
BFXv5V+CKo1rHKP/YdTQ/ap6NDhs9LpzSJvXwzws2iJecyB8SvYrxmdlJ/VAT4CLo27qNBoqPY/i
CFqGw9C6BJbmLATm5VKVly0QKdq7NbWf4WAFdoWFVvEeJyut3jLgtE9wS0MVGPQdSfTdKed/dBjo
cCdtSJCnIVRnICKBllxtrFTABDgOneCPbeYCx5ysmykQw8fevYOgTujjhPw236e23TOtZ39wdutI
K7TdMgRaSYlC4esYKwODW9F4idaB/H1f9/Gmm1/DLUOxdwQn/Vl23FwnYjyKqYltzSyo3tKneCNu
xG4EnV1ziELI9sIw4GeWz8dYiSo2k1KRX4C0bDS6rY+wPS4f/9vDHn4fl2+eJKbe+TH4Hp1Icy35
GNt5+VSVopaYEZqyH8MlekVx4zIji6lbxIlCq144Vkk4YK5mj9NPOuKkr2zqqeCGHDJcsBi1U1UL
YbbXpLHloZAA+uevuo9WgFXsCg2ViEidyJhpWC5XogXop1ANuMgT5X4e6vwHNQ94YiinGvnrPz7v
hhYLKKAekxNdMBmZ+hiso7Auja/WCbJjJzJmLn2cy0wdAoU9f+HYsnkpS3dbYperwgDW9Xc2M56V
UWK2JWh2syHzCOhSD75r/oTH7SBDgGoSJd6LcfQo/h02Phbq2i5IwBuWSiMmssYwrbTYPfm/S0sW
4BEfw3iyiK2PWiJEYkhGy801azt+/ejvnu6Voc6Nqz3skB1ncE1+kKFDFf0V8MtgIyah6JxwmbgP
styp1B8Q2UASevxOQWa7g6u3mbqVaFm+Axxw2i9z13IHm3fBLzHweqepORdKmipo6adOsr+4PyvW
cn0yyUn4VFdIGeLVOEA+NRwzM6YNQoLeph3wALsWwPq6bswz1/IvxxwrDllGsMdAvkPKVbbHRZje
N+ewv9FycOQ+t33Fx8gD8MGYOadb/MRk3qTeKx7HPjKBIJnGp8Q3hjIru84Wycyh0UBBZkY6VBcw
WufepyZOcpOJtiDyXMATGneepabXsG3Z95JSQxeyDkku4VWZqTBC9vQh1OCLzU76v3bShQbcm3wH
r2OKodm4w1pzOGKwX4fJsJKDvWIFt3Tx8Xn0zrSYQGpF8ktlzZi5NgrA/zkMH1SCOrCZr7O64cyO
UMA7qHjZ/VAXed2WNVxFtuKeGlT3D6Rke3H6y+fO5CBDU1wyxukjW189L4Sf4YCwc0IXNALL6C5t
JZFlyK+OOIblKnivigQs2OM7hcdmVpTgc1dOF+NSyBewJzShUya3CsQkxoCpkEj3toLyO0qUPVeI
sa6Mcys4Stn8lOVsuQne0NgCNeCdxU0sy9mpnCjeFJLNfJpvk+U6MgIhjWO8zVXWspsVCj9L0XAO
Tev2PzNYp00ehWxFMwLUWElz872nlVkAeQGSoefwSHbRS3MBU+/xaxh48XI2f1GuQJL0ppHQHECi
V1bheJTAwboMGjpkIVO9xAgHGGsfOIskhNh17/llbfb24cyJy+n5/ei8ZwKcM3qBthS0JhdEo117
Nv18jpbZ77AldoPUMDFxjsA84AE1+4hcouUW7hvaUMqwW2DpwWQgmh9Fm4DADedylh8Gi0qDZD+s
V5XgnCfWmsvWSwz9/UN3r6AZSf4XDSlDAiBPhKApIcBDCXnPVpEWvpUZan53rZlQFvnYncJilHCM
e8PNZzGP2P+yEahbG9RZ1+tKCxIxsa6TfLxNY343NlIj51EKqgvP/lywsbCi0kEfIPdy73xNC3Hn
JuK1SQ2Xl5AkbulDjmtV8L11l05H8Tc8HZCpJJS5eemgs6CUWJBANFuz7hvBzoRMo9IFO7brgdeF
ogkNULWiFsKoW2UPIaHrkSZlkg4g8MZCNUlRIDv7BT9kEVT/BSAAkkloR23wWEcBIAtaLlLkxnHj
MWrdpeBwfwHkJuXZeS2uL8Z9FqiN358kOeLDLGtrisMlJkVj7sOFJP/zehFossbAYlIN1hIznP81
icNfHikt/Z19rzfcZWwQ+Ip+iH8JupmOp6axQXAtWloMemlsBrymi14fCLOkrNtU+F5OD94yCmci
9FzGzgnzsT3d/gr8RSlxOSdAKT31e7KjDOwggisHsdzegLsMVVM/QnPCVAkfeHKqCEqThCePBazU
tuFlLVH9i5LJLLJhb6ioZXIh8gImpGwv3SJNEUxlp8/gUCVWGNIYWEICJA63lrdKVLSrluTqC/hs
t9unZmT5Z5S0Y4lmjLtMro8lLugvuwF4tcjZMG7wX3WpAtOHt4JOVFG4wn4wx4S/z7zElmOlMzVk
LNQJktrRYQBv2b+8torxvmCf77jWWkhDCtjSjAAe3fB67BFthKCLOqb5sJNvy7SY8214PWdTFTVg
/WGThB5Dc5D74dKFnDBg1Fy7j7br5RYk9mZEUkXZyZk1C9Aqz3EVBG9dSCRGaeFtjQVc0oTlvA0b
3lSWPAHmDuV9X/+S2buq2KNgtq/vewjV9b9GGnz2HNbsyjrRMMIM0YTTJRKhfS28r+IuMgoi3qMx
9CWzVOOCKdeub+Wg8dn1I/RMUVNZm2QkvYwWwov5fEIBYDKJaKysMX1K777Yq38xW7coPFKktaqU
eGVF9z1R5UGvFiy13Jcb+wg5sOTZV6kyxlidWjEMSAno0spZW2D8L1oUnEKba8jeS2jeBNfdZvMV
lGO0fYkvHbvs0Doo5Gh3KwlJhlilcPJzOKGN0sXpqQwEOkkBSvKtfUO8VJvVgy0H9y0buGWkosyy
TLoP0w9T/fj+MywyHtyR1cF7izeeuCWV5UUO4Ye3JsVWRdQzDQ1KWDxB1zf+6FKrbzO+z90Mdruo
uzHQmx5VCEn3/iC4YD0706jj93aL1A3aLM0JLoSr0cRyh+yvaiYp7LKSMHal63QuIsXEPO813IkO
ojPv7avxw+mS4IK/uDNL+0TN/1X/79haJCMtd/Cp62rOkKUDDnNAaZHU2dyGusKYVNAg2Cc3H+1k
lk5snxgNVlN4UcX+q8tbDrJArONsMqVUgsuKE9UxF6NH8YozzKr4Mdv7TfIBme7aAebmv2dz3+uU
Qsxo2TV1MfmMrTRErwyvd5uJag2B0j5/HCF3IlJbuCI5BQSfyMHN0hs8JbKkWonr62tsDkLN+K7o
980CT6b987ABHcvCf/jm/a/N7JdlPMADqn0LbSoA74/ZshYqRLavw+xFkqZhwqTg16uzPDgw9+rh
/5WH2bdcYKo1RJbwgGIe1EKTkKxO3pSwrcgJjThgCLLAdxfO+OOYuevWuz+/Vnl/pHLDIKmPJiia
Fr7V4GBWpJEmAD6H7DKbcU0yRwy43CLP/TxYi9jofOaTlwetz0/hvfpCkef6CWtx4MInXH6eFGPJ
c+jmjEBoT2zkEwxmPA+xzudjnpTgbSSMEJRhIO6sSEIwYghRXNP/C6jhqLhiPKgIP8+OVSN/ckS3
R5ngNF0wvLm2QNoVcfTyRso6gGCnToaZwbWwZaEsw9OZGqEk0VSneNVpF7T9kM5lqvnSFei5Um0c
hKOJPoSlj0oOdTazBW/kc9cYx7C1uy8XOSyRQUH86XcpyiEh8AjgfibLbzESGAHxBRGjbW/37YWs
zIKm8KE7tf+3As4VJhKHc6o/1d7sJByYxTiFGMZLwyIjLlR7WmrE0UE+n3fXcz4JR6cl8+okCJy3
msGMhiAQDCintKhqKQdqzvW+VG+cpTv/tXHaKYM/3ZWKeVVcrh24iOrNRKCXedD7ijxsfdkk+CKU
rWmC3tAPzeG+HJjAz8y5ffpXc/CKl9QI1jJJf1Eq5KFSNnUeGhPNAGm4s5zADsQ0H0G/k5IHFqLv
Wg9+KLiznm6G4VPLB8FMx4gkKifweM8uYrCPvh27KdB1i1DaX/hfsaIyf8Z9cbeagnpzhwpg0SWH
RBX8RewOeQW+G8mpTAGw1brDDE1jK8Oy6P1Hd3tANtt1OXElS9T8y/4zfy6/taL+fmXaXzax5nBG
Vy/do9VdG/bJpSkzw98CnyF9xkoMjmyC/3UiIT058PmmKMPDBiRtsIgvrMR4PhkZ2ChTPiHHH1VS
bKCHSdbsiKpug+QpocflDT3zNZ3sm0duSIzOO5fW7DccMzxYnUNi5j3tRjhGpRkK3Old++gGT0fo
8lXS5PGrM2DWijqRs4yW/5EWlZ8yumYAEORGlUyj8ErLN3JHcClp7pxzQYLaZSeNJVOK4PdrReO6
GowX7HzdvsF2yhhcxvF31Rsiw56yJq5L2pr1PIEXxF221LoO5aLtk4tekQ4lUECRnquBsviWa1PS
+pdruTa+Wc6evKEmSC813X0CDSIDyPgkO7pPus2JLPD+nzLBG5L0xMGq93/NBh6KaDd2Hmeq3vRu
TgMWYCeEOJJT9mUF3uKPz+nedaIZb9pb8xUSviHyjElLyguFq3XdkdWDjwVcnu/zcawC2RJs6dTm
nKLLddhYZhedAJ5hdKapKNRiPEzIAYPBqhj/yz6snzlJbX0hWr6+bUjaPmLmgfKC/VIiUXvKRq2U
myt396m1KkLSZXOgZ0kwNmKuxvJ2bxMjKcDoF1VkuJAz9bqi04P1hWM2OAhcVxYiZgwj0+DtxP73
X9Wq6rkSuNceXKv471BKv1Lv1LhS0oxCX3xRV2I78TQVoi+NKyBXA4gMNNiqym5lZXMviGPqj/Cg
sLkQD2Uw0B3XVlyUX5lEfWZs8AEy0Nk7doZeGwn9yeL2dsFFis5wwIf1HF0KlfpAMjIHxIBTOxRw
//hAQO1vKV6szWRtO8oghtmLSdIZ8BDxV5RH+pjz5KpwlcG99ynad75Nsdta4aP3EkCIZ1OLLD+/
1f+ZmPIa+XY8S4DKKmknNoX3sUlhiMTm3Cv7bxkRsoX8jS2xff3lCeHJ6A0YIidA4A7iWeq6ZYUY
/uzBiLKd824GqdY8Fc054UHNVcosImd1hBkYphNUa/i5+znmSWAQcl1pQKTaIXLHg5RJwrjYgHhg
MLy5AlxxTVZfCRYZq2vQhThnEOXAvqDiSsICxpXVXlCe0lz+mdUFhwz1IX+kJ5FHwazEXU578uJq
owXr4vtd23ltLKuNkdAqWzDFNqH6qRYxecp3wr9pM0ClF/ZTkuCZKNF+XYd91ssw+eJvWZAvC67u
wBe8sQ9lcOqIajTPTR6BJZCqtDmlJS8MzRn0hMlDtdzaKIo9gYGAG6sTXTflr+reDFMbX+MwKyl6
BaE8HUffsdpJpeGxS5WclRInrN87O6Y/mftPSVYqUTNU65xqmSNx4cSPcNO0SNZrfFwUYQWakpbk
01R4snKlGf0BJZEybLe/GOX0NMPAl1GBO4K7y2aJhOf8utNtxBexbcKVebQl6VrzEFvCZ6gwfCzR
qQ5DRVYk8s+uw08ZzM0YmdLQPOJIlS4+Pwft+KuvD+9dZyrOdE2PeK8A0FhhDDf3lbp0UnV5Yfcj
R5ngt28fl9iV8Kky7/1ebSUkWibxBOwBECTQ1ypcVFfC7XCOEdIdW83b7Fd1NJSkCAs0ukfzkE61
oNwziA5G+aIDVs9J8GHpdveNb4R+oG61J5+BUwCQ3zev0zhnKln2KvuVmfNXqloFg+XG6u54grYL
PPRaoCtE9PXmEuvS51/TkTtbCtcpZ+3djYx+p4SmuarTlXY7rkwXGmIFiVFGyC7JWxvLTL0GmCbM
iR9i6ZCbePagPkbWVKsKYy1wl+tvj8Jgvy7gGhPeLD6dtvzI0+ZNVniXDX0fkTZQbyyHPogZsk5n
UMHLTrLdQwjyUjUBYQdwOGNhejexmzDsl3adxkbvZF0d6lIet2ezIBxFf3XSBCT9chitpNMji73v
8vAdg+4FWeRjbkwSW4idfJ/CNWYHdADg4LL5hys3/Sc0vOlPO6JSeXVrDq9JBM8kcVUeOIWGI3Qy
iO+VYMSYyc/uP9PDwKmom8e4UQ18X7SOmvHz5aUEarSlllAD1VQIFGbeqR0E1cn6CvcEqWyp4cze
og6AICy44i+f6ZTbjBMuKlXtzsqRV5bGRmun7CzVbvoI0HRUk4DAJJsPHRdKieFp3dG4bQDWyLcA
v2UqGzfGJtyVJyKG0UeAT6qYahQFJE/JE2s+tZLXiTE5ER3Vd45FsrfMDreE/cJYFW9KJpucuA15
Mf52kQk/CbLOmyfV9pIa99cjM7aqGBMOXPdb+km7lwTA3ShMpdYBXPY+fg4O4TtZc8036UNrXYt5
HYN5V02gDULwCIyHQQosoWpw1BKxMsXA5G3TpjAVp+mgoDT6oVp+barX+XBDghpxN/Q9DRt53odz
ASudq01PlLqva20OaXp1tUupDxI7M3cKFdlxJk9FEL0Rg2FNs3CcjMDiTcODsKDlK/+6xmDOJ0wF
rSnh4qnG/wHlcQCmHFIhBf7kyaXvwE827HJr5wpp92j6MA9PYqA145ypZ2QuP+knAVWl34lcU3cj
vP5qGA2sEYJt6K8glRr2I58gLK7FIlRDdKalM33qLdL8gxaGBsm2CQQN7RGDevjpmFbdgZFtd5oV
U1EJm7zHW0lJC0pkx9HF3xny76lkMI68xahu4g69JJryLh7UG8khFa06YDAaPxTKWC4AIoCi0S2K
K8o+iqC4HNuqztsYRjiIAIWkrAxvAWyQdkpcQ/eQPYeKjgC9ztmY122+5rfOi6pLNt4VL6lt5CIx
ZZ3W68nxek42dl/uISUQcYxedppS1I6hHz7ucl6Zh1LX6+bTA3d2x+1MwQ1zVu2ndoapEatuyBWo
0d0UeQzPkD7U5uaJAvRt9ERJZ+Dc3oeOjoDJYY2zbLbvtHbIIJpKpzoZg8KP/DK84g6v4ZmsAJgZ
zrMvAd6wKgqvaFvKP1DV5+naWMgO2F5/v2dBxxIabU1+UteU5WCQ94byOkmZ/UhqNxiU1LOh7DgF
LjjnnmqBT4CwKIqpGJRrUSnGnl32/f0WCIeVofQARsKwSeCILc+BIJGfcvhinMLGyriuZNoUlxuH
wIwHi/2UALEYrEvO5JlJpBjANZQTR1iPSMSl9lUEKV46U1etcCvUvmi3kFu+F1Aryw3xoUXLv/oG
n7o+xcZ7RGfZEDZscZiAr4DcEc57+BWtjc/UBQgQNkngH19Na8AEL7QaebmNdCEtZsaT2Nj+8lEv
5LRIgmDdS9a7oFFJN3sgXiwthRiZJ7j7In5zdcwBh3kMiXrDt6kS1aDp4PmiPdEVjaKo311BAvhb
Ic6347G7l6gxK4UXZug/Awetx5DrGAFFq5d2utp6O10Vv61SNh5u94b7t9eYLxuMClE2T46fXHiP
nGE6B68DZVQpg/eZwlhbQbe01QMzlHQiXtDLhaBwss6f+zaoP9M7tfauyWw21dC74j93wtr0KYWi
bHlNLebDcZOLqLQ3BTFcHC0hrFffC3P0RXtjQJnGM+WCD30+UCi5yZG5Olv6EvrKStwov7i5KWyy
IBz5Zn1VR1XTE0m2kBJRcEdsRyYwkYreKTUf4Y4bhSo6cNQPExzQaiNLWG9IpQdRCwPgRiUUeTKF
rsICFzPnF2Pdxy1mZBGeh6Zca+NM76DpHu5C6RzfzgYi1uL5w+hQjqucFWymvsh/4KFKq9G3LxMv
XF0x1ZAL5Jua9IIWzX0hH+fxJA6hsFmbQ9UL6MGriGouQNeamhmceu1F/CEChvjiWTtl4TFrJIE1
XuQiaU2FTwFLjJ5fPmA+wJ0DaPbRfGMhPWgTSJoFOsjspDAwt4kk1HFwlas0kEuEV2bBa5M4yv0e
+kTN6o9uNl1megpVSHsOXIrdiDvdP/sbfliTbu8xRxkRcIbU6SPfS/y+kPRGk3dhljQW8eio/9Wa
XrNc59Pp8sGp/Z3oV4XVjLuRxmF2qdmcU9xbQ36CYzsiCbyX5JhqtSdjTf/SvRRSd470rACI5rc7
5H0g8e9lqfDmkiZoxepkiQx0lkWt6bMRSctXXlYEPlmv/LYTPALRl+FHOiLDQRjkJ/q3xuGr36Wi
DB+VhdrAkCqUS32Q4Tl7sc8Gapr0ZsVZ9ALhRsiJj/8f5UnvKbP/7a6RClb/PBWQoa+3H0uL6Iwj
mURthzu89AMk8ahgLuP9UGcHy21rWztou/7uZtIoqFWwO5ML8lFX2173aURNy2dSq5v7yx63Js/n
YB6ASjqIv3a6hvMvoCIPu6GWGq7lPlsfG7IsxRc3rCpKKXAVQ+i0fl3ZIajbvF4LDgz69O/fEu1E
h/QV7waN0A79pGhmclU/iUA8OCt24U6zroDT8J+rs5E62v0Y4I4CYKKK2t2WVyemma0Ajrv/nOW0
fPbF/zFFDA7icusZs6zKVcaYnmidbTK9WJITyXGH8pDwyLinO0+YEK51pYgVLZx4zAsn/63iKFsa
xQn+O7hPOmQuRb3poX2BY0+B01nZ1MxXTO3PjbyeQ7to8a+Rdj8H3Y+KR6/jLOvXfrSECKKJGZMN
SPY9A2yE2bZHOxlfV2Xqlbfsb0BGbltN6l/ZJ/+V1GK0aPTjf3NyUPS3yvAA+Qkkh7NEjLn1NHKQ
OAMpCoipLwGBOP+LoLlNufEtey2DTr2rHgRNO838f38+gcOW4eNiP0eRsrOe5r4KXW6+Zqk2Cmsz
IQGbO4uMUwf+scCfrikmRSM6XlAdXUmsUSpPWSkwg+dlp+LJZxwKpr5PmhLYdxOpS+KJ9uAvA9rX
mh9a6uvT9zODUdoFIF6CLDZdy0QxHyWPggazKS834Ngyt3iF3obcGjJuRTkk5YDeVfsdmjl7AcnF
gpeoix1zi+/FmGI6PS9a4AAH1sRy/uUIFGOXIN0se8Onc65UwjjYTH4pGnY3ePxs8c5/oOgYOZjF
3cYq/2D7hxQvdos/g6k1J836PpO0/NlOyLNMjG8D1kZR2Oe5RNi7EbKBJUc4hfW2lGWSH9X4RGnN
WK9sZ75Kms094k2oyWCYH1ToIZbBfiuFD5qUfASUSoZIwEDZsftwdJxigiGMh6WmU9LbKbxNwxwr
QQmwDUzdfiicydnUuG2JWGHREo5UERQJs4dFtlBUmEHboEQS9xX2s1cYSnGE1odAHaOeAxRKEL+p
I2JoUJrvjnssP0ju0+gVkesq95WEnBD2NA9lMm8kef8wg+zaXIw/6rnRdibhb/StG13HqJd3PXEy
oKVWicoSXBQanHW8b/pQIyc6rV44YKWbqNME1G9iipSwOgSF3ZuJtZ5lUOJcrzQW6axh8gUuuyX7
JNyFWekwsFOHfsmt+n0lGHfm2Ez0vieoozUPcIhajZEo547ThD8ONP9honc4Syu16Jlh5EY2B7x9
FE/jV8bxZ+n9sayZvf/Ontl0ymu+9E4hgv7LFbSmjKidiQ7Uag4WFLB9ca5mybU8jItK+33XLf2f
Vq8MfPjj9Hc3Etern8Q37lmhLfCnvAEwkNGOQUMjQ81qocm9TjNdcUjm2K3f/9gxIRBz6BCf2+E2
A2hGX0HbMUioUJcuA9miLOKx/PNqOPudXUTX5LhaQCL9t84W2NVPQmxRsme5rRsfCVaFniLgeLcB
UWwSlXocJzGrlCbuOrv62p9fbOHjZj4zyBlsCoG+yWFjbnlyuN6s2F9MOqwRFHitBkSteKvICM2a
3r3DzXTs1SJs8mnVUlXUO0xi4A6kzMLU2icHqPah6AeOrAnAdC9nWi6KvYnd1kNlCBhBgbqllgLs
vMwTehA1klAaMHKW+r5chKwpBuHh6SoD57XYt9Rp/v4kq+Q3K7cNxxkWA9cZTi1M7As32REDlESt
1h0YU1I458mxzWhaCu2SPiQuyZeJc57ufEQAlL5ng73uYyb13/lvrnlQ62W6qol5P4qqWe5yuqzS
miACypEb71ZLNCjvYnOPNHRmgjZfnViBTV6XgPCzTbMbu7MMBwm9qWh4k30yLKsCcBaLEqE1BxRF
/K79BqqXsnx/mQ0e31mLHpuUqFaHJzUP291lvkW17eh5qYXHIlLE1E/YGu8NAYmXKBtbbiUsUdEh
DAR57oVbuLE4txTVA+2y7l2PVNUWwSEeLrDJTNcxZ0fVhD4+WV/icpkphQvxhATNVsOsNHD7JICc
1mORW3QvJWxQ0GYhZ8exlaARAkoRyn6WnRpiuRo9qObISWCIP+Bhy6w6XQQLiG0ltArZkDEg+7j+
ajtbhlCwFctyyqZfXi6qtQzfq0tL//chhcCgB9+3eEYR+GkLQvJ9vFVs7yewohlbHzXHzDDY3VLt
G98DQsLmC4lyHVcJiEgvZrDPlTOSpCoCc3TSWL/oiQbx3LDOfFaLi0hna7cRXVCzGYxHDaEOTPYF
FhvjJqe4bx08dNYAoGessEslrWdmp9zpq/nM5d67tfDWDK2rqChs5GWHShUja38GL+EO8z2CMe/p
nAI0F1eBond9iEVV+3SuhLbYe726yEPgdQSQs8HQ99twZFVshTXkA8Jbg1Tn0mt9quUjFI2BT5f9
FRV5Nquuf96yPRbzFkBA0I9kZkCCO295L0SNd+XxidSxIRNzHsnVQi0Y4HMCFvk1wndqvZx+M2Pb
VQ8awl0pJJGJcGkZ/4hBnGKSuskXrSNzJP+HDyUTOvT6FWzYxlYAZWKgEVQFzPdJykSkHqbaPMD6
2Jivq2zLmlCFUoIOSuKh0tMrGVU6PakIWBqEP2Pb3lAxzrBOysfuyTDewIXLkQgNCKzeH+DpoUNq
d6uSr+aW8faH1OIZpcVSUSCDw8+b89dIrDg/oX+HmhXFTdk9HTa8RXBGX+Orq3IVU0PGVxhfmgf8
bg/oTUCAlmM0zgpz1hJA3fWioIBFVzGe1t+P+eyczi67S5+7fP47nyk4s3yH965LLVqBLvCcq6+p
O0XKoL3o+NEY4YioIj2Zvbb2UhB7HGI6IY/6cEPecO2oewRgJI3OCPhd65OYlkrKvQW5Gn96IpuB
V0IehNR4x57CjAgmrOiqBBDzOb1YEjk2dCvGzQo04jDlEUlgkb+GnuzHdwEXMwdOE2oczYEO1xJg
JgIie8hks5Q3Ey1y2/HNl1aye0j3U0k3dpeDFCLz+WJuX05VtazWm4lLt17lTuc2HdXr8b7HE58E
Q+013NpyUca4tftL8C8ZeoeZvmoJOPCYglBZc80a6fr0OxXPhJBKM5VrIolqnqu30XTI5mugTlmZ
OgzFI3On5k8WIJXYIwUvj8HCr4MfiG7EJOsMv2eLS6nIIaZdEhhYKSspBFIk4MLeXUmMymo2qfWT
UP4AkObwEnwQEbl9BwggrEs5jot7RevFfrEY4k5ZbzGGz+rH0LqtaABF6fWfHj/lAwfJi0BMTlQx
+dNxGoWx9e5J9gzMA9XyWDaxTAuUMcic97hBN2HQ5Bg83kElu05OOiBH868E6uBotyY1xEA9QLbv
ltgRrV81rU6NSKyLfxHMRScCTylH7IV6IEo772NuP4DJ9bcQFSbQW+iKJfE+GTPnz4hJ1OPekfi3
9ASdvNdM0C7qYgYq6s1oVFZ4Y/xdMJVXo+Mi3c1NTnoBmLOet599sahRgBTZPrLh3LnxeYTtuPMH
hUuN6x4yOHIT+FIVabb2zNR60Bi8hcppMogMpgKM1Q44gcIVCk17rBIVcbdbAH+QYfW+7MLHTHRQ
W6qnPJk0f58wLvJiqOv77YKVWo6G+d0RhtyuKC0mLt2+PaYgcsPCychHKtGtiRuYRtC1gGM/6RH3
h04AU7953JNSxysySPejwGmJYClpGgaqQCMka9Hk0qq92WGRfhTYETFYl6KPsjotoYSUF5WD/cdU
gpmAe9TgHwd7eC4olW29J9JJftjjMheH33d3nUyPWHspu6lDYIyYoPQbth9qlTJBmcsaWPmH/Ke2
FXJWYG7FB7UoIhkkP08dMjz5+EAQHKr9O4Jl0WGyEMPfVtNywId9lMo6K+qar/yL/VDfwyaaS+47
CdO3K2Z/L4rkw6yHUGV8k18Upsd6wuKA4bfg0cdQ6MkmmqQNvlYWKIT2HJKzkQk2y2TLGbVWHYDZ
iKVcSH2LoTObu5AvifRGfYFbhP528HXvaFpMmPnpT/CCI8B1V+nQPghdR60xjd90onCGEB8atH8L
Y3ETty45mt4f8D6Z1AtG+fOyH5Lp2s0SNRvdxhIsneXUBntUYr2Foh3mvfduHD7xxRN+vmGmzBYw
J3j77LQcpmNp3mzfaRT/K16mwOFe0X7Mhx79KN6JZveKt7VTYlY/L5uzQ0H1v4b1BRhc9hJItolp
jNM3b3qxnsi3W+eXIY1tK5tuRB3GCI1fS9O6a8EEM3RpJ7groohdA/CThBRE4+qdV0gu/FhtNB4M
AooReSP/pedqOAxa9OzLs9aDXkiSAMp9C3Uo0wVwbNyDtneF1hPuoCGJNfOCHxmtEPnSFd9CQ5ex
u/V2g9ZYkImd7FqVgerAA43ipJjjFeX9VzQ3TXV+kbgrNwJcQ4x4YNgOc3/nI6a/9tNZHcVmmoYT
d3jkX9vBwzohdPYxerRJLxA57c/gw+jwG34ChutO4GR0bAVQBCNceKtXj6ZBdrfvuLurECvZjWWn
rtzSX13eLlsrpTV2lpPBA82wUBZiYL28LWfluyDjukmhH7knCBeFf4HoN1ZGL7tj9L+mt+KClG+L
+Dufo19iLJUmOL5hvjkpkr0CnNvS/WIISzMGHOqnaiA3T+j7LO4o57eeXkWhFp9RqXh+Rxfty/px
Dh7m470T3+/rA1gQ6J1dOc1n+/KY2gTxqlvG8Hj7cSTEEXkeFavbVwqKm7RJ0MtUi2mqPCmK5db1
tgKk9EK1dIpaT44ICou3/7EkCgGSV7KuZMiFpyMQd7dLFUXgM3FqA+R9RPEg/2Vo/+MmtxnbnrAS
Hoh+raF1tlcVZ9qEaBEoe7PVG67dK8k1GD6p5PgtgnmLCznGT7/Kr1zJq1Taht98lavk7pBZBylX
UqlJnws6Qu9LMbNxKYRkOBzcR5sBcdO+TjT9voZ4PhjwmwnI2JsEOizoiHEUsGc+Tr6Bjd5uSynp
45rrAPbKOcWTx3jdakaO+aB9DQqy5IVOI9YVAr8ozV5T7jdZ/Bm2fmXx1fChJkSek31h4Jaw11XX
GuywO3eBXtfKPnMJTvbxnQa6goBB/Hd0E803CA5mlRgDCd82/ppdco+hI6EfvdTPXdDuJHZGB7Vq
9HecvgjMDev02dlihwiYIYWJDv/5dDuigrC7R96lvYkX42ZoQL4W1HzvLQGmY5l86GbIYBYgWsDk
hEEJY8pkDxMASsTXf/lhO0g/V8YColed3/OHZ5gbzTte4dFVa8ojgSa/5DXTfyS0Yx5TnGK8SWbV
q1p6YR+VWhza3Ew4JLVJcBqyRcC7Jj1PQ4hdYSWODRpRTG8Yj18kTKMhtwCNnsD1/3xSbipxKeU0
u1gqZGldntB5JaAWltjL/P7UlXeQ2jcoN9muMnPSMTLxc0zT0p1wIPMnZW5U1eEvWuxdIz68rRZY
8lYls254CN66XkpgaNO2gssTRWznnmLW4zIJ6cM2A2Uhl3H67DuAR+aHpyZTsYyG0D+gCnThYTau
x1SwxfcmmAIg//LYjxozOoryH47WOqOR8kQjXR45gI4cVbwFIlSCDbc/qwuxd6wOTTTw/yZOG8OE
NM5nOQ60nDti9mPA+86w7G2cNqUPS7uVjkwpDjI0fgPcf08IuQfB0zJD2xgBsI6hAWqI3l1TQv3R
1yYnYlqMSb2DfHwV9cwMnyfElmcxt/AuMWfha7wrF9JqyaNEQDIPdrazsZ8Hsnb9Q5PutX1xHChD
dte2nqJz8w/j5elkBybuyVqmZA9pkwZYGhqIWR+xOZc6RgU8fQBnxUT+aacphSdY5V/EvYGbN1nQ
YrHBTRwIyKT0UGbq+oQin9lVH5N7b+1TbXVyIMEUPvgpoPwk3qTMgp+2bvbmpb1lVVUuKuWrdRDR
8fxWWC8kHnyfYLUe36hOHFL1jRHDN1WjAZmOAP9cPXzsIpmwNsXotH4hcS85u6ivLrfkWAnHCB8G
4GxEmfvy2Uvjaj/9hwWoHRpkTDDuO6KzUsmnCswbYeLkykFIBNdaZZX+WIJaA+TDOEtILQY+JBKI
Ywn2J5Ict9KFaM8xjR3Zh0TXUaHt5efBhBeU8D2z4ozV5oFcpj0yj3rcczmQUk8zrYxfzCftraBo
l/fPVYRnvyHK2lkeWVoNhBJAu4djp19jqB2nnh/VvjPjx7R23nUU5c0kevancjfQVGXSzrKm+inp
/sGRXvfvwNRMLYMCyFqwDVZy41SHG3aPTgiXj8oix7SGcxKLy3GT4f80MTCyuB1YR8IPpQZfHkRD
1QXvQrYW1jlQABVZrSYC4urFkyZ8F9sWIH1Y7ByG9RbsMh0mR+1v7N8sDIR9Ti/8mVN+OPAD2XS8
5+AmLzDRrSuuOH4Or219SQefueo0q83swwf3z3KENLm1R4coKVKtftUl03yV2t5gDU6rnGS5CPfK
0ehLRnXUpoaXDPYWUabO9mY8Te372Cdw2jYVr65yejgPRuLxYuYfZzQpAmLUtM1toLBVu76YaQrI
ZBAuXzM0Wcsih0aDjhjC4AxxScW6awBBttDskBAAqF2pvaXwSPi9VcPBvFuH8xiKSLAlWAzzpR9S
0zs8o6gnv7Y7EDdFM/pEOvU39gFN9KrVOyIVE0CN9tlvbmXQYcGNMA7a78GJJEDnzJbafjGK3zSt
EDAijWq8pZlIC5q2ILih5bZ2mYeEFU5Xt60kNz0Zxv9dxi9zfo0mf+/9c1ho8pfrYxyjoJuJY7gv
f2XKFpaOgr5m9r4iFdHVPbaR6XvvJ1oU44/R683Jnu43ymZZqpt/8WjgBmiBTq7JH06+kN9NpFo4
1klBl9YK1fHmZpObZtATITHZEPf2Iffny2abPBREYvBobBLfuN6aRrBN2tgpEgLnry2CfSvodTE6
JzDJpSKKOhPM+PpUVfe6GNKZOoJSonyLWDKXti5yVENlIWYT7obr6ER6aJZtEhvxB6VHDCe2ynPm
Pd5yNlbXH0O4DWx3dR6DiJG4IDWmEb0mAnVOZczqqD2s3NrAcphLRVZwTdP4zGRV2t9GEtsRPGAw
8yIkBtYG9cSqiUxEaVCx+MX8l6I6J7WDkKGFdGIqJ7QuBh3DPeQzLrRF4uBirZrOlY8vFs6TefG3
4msOJv2tsCXrnfn/dEn4Up9hwNgrY6feUABGNeAAvoWdlvhRTuZOjjJpO3M8x61DVFsp0Fgt8BkI
eAZYeElSS4b0yNYXiKKJfnGsIe96KLEHVBBo2u/uITbpZN4TfETdTYMMMkEnd14GWcv49EZ9yQEc
iYmTASdzI9Q8ogjLiw/XorZf/P0ad9pt/rzLyPGrZvYlqxHuS7BoDzyHTBjEWM1I5PSxlw6Aq6wg
lWaHc4sHr/DNZhK6YUKGLu4vSryF+nvs9srafhX5eh+H4+bIcFcVg4IRA62sCdaz71PkvpJ+RT+J
UM14hYhbbh6B/YX0x1cganL0kWKqZi+GGOYfa9qdO0Ouvyhc49rcnpYKf08ddxEP3YTQ+3LyMaF1
Je21IM1KUAtyarIdSJjNtEBEIBZfzUnOOo0ej9ZDiJhfePUuM9Zqn/ZJjnfPP4polTW4Zk9u/2uM
NujcQXcs/g27+FKOd8vrSwliyBrofKSh7fEbb/qorYA6IYkhacjUDW4Usj0VXMlkj6AE1+6G7Swm
ntpCc4fW1lyeu3EKC7hjz+LhrztzaFo7fl5RqgnYO/6IAAenzJIiwKim6NL/cKA749ylkzRyVJCu
QVgslv5nFJTalQ8Yv5iz7h1jTgEWSPjod8MSiB4fIZJ5Z3GL+ZypyYpCvumT6NxLE99I2xjt46L9
ZSQEpvmnBOyPa8nDfdB/bvKjTov4TivkQbT8nykiuGB56tnwuUDh0+w7GkCqWlW5tt1sfqMWVv8p
tqi+awoR9OTxP+/o1XO88ldurUcmz/C/9ROsv2iSoG8UuUUA9IddiOvWJbk7yX6ZpDIGSf13NZFb
Q2yNKU6BVZhh/yxdcGC4gkiAUeC7zoFouqopZ67ryFlmFy7gOzlgbC0VK+PgBSbrjziAZXBtm5T1
W5LnpLFztUiEmbKabfanOcsZ3KCUzY8D9rmx+7/6EG5m1hEthSzXdT75LOJhrrvgFloe+9/laJ3C
0e+y26+3Nw2AbEcaRfjm2JJQCEpd6gyz+J7cB7tTKo04PtsdZFnOjbxyDqcroFP79b7TnqhHhxtv
m+UlsNwv53xjzeql9H7nm8jYZeyCZ1TB71nC2zAKLLazvXzAUJOMGV+HN1D/Zrfpd4ipbBd8nbFU
Tv5pMUvXNXoNXs0t5E2c6kVnRQTuGvgEvgnHEB2DPWtJSwTy2Eeg1FJfD9UusUeE1QBTNSvYqW4i
SCErZuydvcXo6+Tvszbj4yyLcrQQhRBQPAjpMGLagWG9HUz9/kZliq8C1fH5Rn+MBR/55gwLpkvb
DdyoZSqfTBggbexnhnThEzeHAZuOSyjTErWUOTxOeXT3+qTAHLJ+FsZawRDVjCiOO4ql3kxZG5/f
moG6AA/6grEGzuGa47OZI+ANVyXsi25ylz1asLgR5taxkVD7ialp2yxZwF+0q/Hse4X8XAYXirVs
v7aWL///8oO86DffgZxtbLbOHTXHRaYxPr5TWZN9jLWAxKjR2Q9Kuht8n88kzA7YDvcccq1eT1m1
AAqw/LwMT4P64q6ZtVphle0YBIPH8eK9JZpcAQa8Mc73AzwVqzKLbvj+T0gRrXAfyFiE9IX8rrk0
AWRiyMz9bjoieDnVjCT9/KSP8Iwbe90VoReMCW61Q9Uaabf3z7cPqGhAshiYqweoeP7bFYDDCHVV
KPBGVtSxlpbVSz6OS6ClydwLkoKwEqOQZ2YyWeaRScQIa89zYRW9ujh/nlJv36CjnTCqN1/uk4Y1
Nx3H6iN5WMdOiSvtzMm8pTLOTBBfikUaEhCTaRCsL2WVUyrI8j1O2O6mjsJnvnX3m3knplD6YAYJ
b2Awq+FpjxeQydHzUakoxN9QT0VWkLRPbP5ISyGfOPJfYsD93MkS6yvoJrLspTIt+oMo9uVXSev6
1ckGS92wNoEl9SrYAthOfip2d3u59f3xQYnWXIE6saqGMVvAKyV8CYfwj7Dj9ibpBCABbsaJdgOF
QdDek3xZ3HxQJfv7Rf8w93rtyzGl+LXsUNABHFOxq19ojpfE8Lut55uyzUksy3LsQ0NMiLNCJm21
3BA7YAQ+2xDxWvk2+hE9LwH6yJv1+EygqLM4b8l9xqUYjMqI4O+6hZfqHI0tWs058VVNCzJTSiYy
8J2uTeFo1BDJzTCNZGEiSGUnsa84ScGGtsSp43F5+mZTREyw1LNWC3k8YXeLLADu4siEOmP7/ciS
m8ts/QEQXRLqzNrKzViUi7f43pqeFB+Knsm+Sy+gbtkJY2HeTdX4SCagshqZALoDJuO2ZDpgVGmP
Wo1qXKVzxp2n8EU6T4wo4EB7aicGgSATDLDU3SxsCzseJljoc7hHOmDlcIZOgw970q6FNgUOnU8r
ItZkINr7GOvl3s3faf97irInLDYIazOdJGi3cVIP/mMu12tvHJyYTLpcC+0xkCknb0HMAkE11PJW
wi3jMqkfiIc2CSe2og1+PjbdkC4Sj7rNH6L2916Gx21nfBBhexxp5h2yLjeyNJG6YHhrRdbWDwVV
vo15YfBweal0ZKB+M47kViBMz8bKuD8x06iwZapJAz9sGHJpXBFCgwsevuXGJtulrDWqUsYlrZix
ad1OgzBHkLfQ7Aa3/EquIBB+PO9EkF5KRW9xEIy1DJHLyC3f+yLLRxstBydRYVV9UFIsCMJsoCmN
rgN+WsPf0dp23W9BMW43JLbIKKMRiQUzOvvnQHblaaOyjlHN3O4T4kZ+gStee6Pvo/JY3mXQ//Go
0oPKNwfo54GmLybW08eO3Y3KFiIqUn3/1Psa+da9P5sEzurZNHewLxi5deVUO5XVE+aUiAj2BJS9
dpYoMuo/HJmayJTrlMqGKsTs5iHXIFSKxq7M9+Yvn8y+1i2FOj5KmrRgsR4dHlcVrtRzNmhJn/hl
F9UI+gz6huhHblii9h3eLNRKB5MEgWyZ+ce78AvTf4kMo4t2D7Ehf+SdBbOASe44CYh9U1MOd+un
Imj2pSYAs0g5BfE9d7yd1ZF2KYCmTM4nXiMDbu9gyfR+ysha6EMz/RNhh3LI+2T78W2hpUmAPYCa
Q9Ka4qzbWmBGbk7HYwg2U1vNbZDvNVgChb9kF1fsaQ924/EQosptSzsF7iWcqCatfxdcY4MBNzaa
lQoshHAvOgxUiefL+3qjAWVgc0PWvia44+Gum0NXH6EdgfNsXgzC3edNCupDftxQ42VMHkzsgg6P
UaTpMszNHu7z54JPkyJLwMU+pw2g0JGZQrt/rD0QxP6QHNn93Wx09d7nQntjtck6nul8OcJYN4CI
9uEgtTaqxg7EhysX3eUr2sst/X4FGQC4FrgqA7fuenZK+91dvGDseSz3gQOvhiye6EGVDYeAZ1dy
Y4BK+Y22kY3fQDeCQqVcpMRhwztJy9vPxkCx/LVpUMPTFGRv3ZBAktAksSGb+f+6m0c93iCzsoDf
uNE/ifa9rrqjzRol5wJexqwrbd5KQ/AhvWds1JZ7M5ma7xB1KWNcDYgPsA75I0i1DLcZ2ZjMqOqK
aKkIixxu8oEmT6tmJGghs9FRvzpntrSGpwS3579ZMDbPaJwN25dQNgw5THmJEF0y9Vh9nkS2hb0Q
oKOEz7fzy6xD6tl+UGAAPxTfiTLmfw+DmNKzbEJ22h6m6SqNjUS1ohAlaBap9bwTNdPoGr4qXqIN
pXdkeZX2CdQ7X8uTuXfU3tHMZFGfUkOHcCrqyaR6IK6LfZ2Im/eERDH8+cQPUuAsWYoemb3An45f
DILlPuQ18LIj/W/EVZw2/x83kDmHjtf39Je54ukdmuKv35n05N+G6DIdX1qhx59TrjIAV2vzZt3F
LqM4eq+c1/V1q+/LbmN/sV8yUolI8Ma74aswrQVjEXb8pyIaHPBbmlHqthj2UL+76N3xY4b3cJAT
AoiBCb7FKem//ilxZn5vK1tlY/GcSs8REZdv+v14CkdkKmBQhVCGkbJgXsKPUmnagqCZjr67BYtk
X8eEfaWZDm30gPf9szrTpkJnCOdzmpYEa2rTsHqLDCd8TL5OWbanbO93xxOIxwycKbfyID36bJ0b
glhocP2m5g9MZ8xnRF7JK+fp55/8XQ+VuGJFyi/X2GPNgSqlAdl31TUTlGpqPfh6aY/3tUEV0S3O
TGPu74j/HhxpGtFBar+QIX4SDK5+qVZlTkr/mt6sy0RQSrbPot1TTx+IR6tsvLYQTGr3g3BFduxv
NV7XpiDXZbOWVf0o7uesNzRMPf50Jw2qJF57fjJ57cOSMudcgzhV3mRvoZE5xFNOcDOo6hiumYGS
qo1YnmvsA7tcoyNK4T3E+njZ9w+3hxqLk5qBfY+6YPKZ7dLMSnkw4rRZP+zFYRVLr50jKCrT1Hwm
PpEp9xMXpA6oGEQFvvtIxd8IuRXq6P83u5eU5Wo/MDhJXIDdl+mtsOMy0kQhCUpebli/bt7H8q1D
D3jwY/EhXQG9rf0LyPMQBpP9i5NVDJGCmTO0w+Wh8rsxOclQs1dkzakJN9pG3z0+BW1ftvzRiH/0
0LAkmpXMtx9SFac+yqsrNkF408KfYCq5JGqI/LWEZ858yLgs5Kxwce62vtcj+SawteItNNmHN1n+
V5hZV5QoEUV7xCEbQRxZdieA+XsKePtuUYJLguecFP/4dIOdSDxYi9aoVqOPtwvaScou3GZkvpjh
9kfBva2ZkCAHgeT2mIrrXUsGaTmlkS6BKceM90BSNLw4kRYZktK2EX80kxr9T6i5ZW4xFwlOMvXP
D8aZqiFLkwlAU8W8OdTSFZVFBJXjGeEatsGdV2HozBJ/Sev9tm65TT942hXOzezRMESpToMph3jX
tU/nkPIr40wTakDy+HoUdkHH4aloyKDzy91UB5HuV2PTJKh+sYRkbGO2273cHPXeNqA8LsC+0RQ2
kQJcssZr4yRv5O+9BG3VnJfumU5PfuxA4VIIYjUzAlc4IX00k1NCL1i7o4kaGXc4bD725u90gcGc
wgGSc7B/U8KYxaPX+OlGEfectzJtYEcUECZIhBE1mda6Yo/tO/D8vh4vCPNNswC+MPx6xqZnjmWd
Y/i8rjgvimoo3Zu89J4HZjMU4umcK/cWiNuBhEruel1J0eDKltje1qg6ajlft3CfZYUAmpivf0ru
zcxBlXG+wpiOZnBt09xCtMjpkWpFdZxoVjwGatsTvCigKFTvyZ9/LiQRgxSpcgoDi4fHJOG/TZ9J
RGj69e557AAJmsGifs+MnIOZiOMUYW9ni6HcJm+DsHx187w6W1Yoch+Ib8eNxZ/MrHACR/BorJIK
RSe6Yu0AK2acE2M+8q0GK9vl4gAOL5y7UkXHnDJTak5P8u+thf8yvjzXD2kkYO28YTwhO7uWMjJk
KyvGwLmVZJMI1MOQ2ltOUmmSXcLAeKAj3IabqorrS/Bt/ihqqMG1WWd4S8o8uI7IRjNLItEfd8oq
1FzhmRKXQAkBLlb3QzSw8v1E+gyFuYpCDKihhN4kHQj4a6uq6LXJ54jGz7uOXRlGyCDc0WANfpg1
lZ16w/+cs9xGS0haAOMwHRwfSxznaseULLPNQITfKrCEzBTiYkSlzBfp9slUe0sVTDoRQm/7SvBm
X7AEHMvAHKgi4dbFw6k3oCSJ0uam6Kh6jpzLGNxCphaysfCOUju/lQ65BJODeLhYaaSpjt5RKRIZ
QFqcqeUQR22NhEG/MVvJd4jKWBCyOrfLdh0/oipyXTjWwDD+jXRtoelWiTG1Hck4HSiEEu4oAD6A
bLSXJaVWOhspCs40InJI9q88etkwvUE9dJss6YkR8bw1PeHzF4xmGTb3kObiREzf0SFHBI67PbLd
spkO0qDoaqpZfxjd3im+K+d71WojgxXCCopaYl2yufgU2TuoGw3BY1ZxpneSToOy0ZOrKmgGyhSP
zn5IRlEkLLIOr2zqCB/AsKNgmAsiE6Dgb52Auxsdrh+3FadElkh7m+2JBMaLYhirQQ1nQTAq7XRg
i3ztG2V/8bBUWq50h5A9/WeUjBjPaARCGibowPuyU9pPNqMMBrqt0MIjeJ8wagGTLdKVAeWNRCsf
Gdt4tSsPJd/ggG6VRgxUHM5aL2qzdwvudNekSvbUzDCpbQZf6l12VFOWHA8HWJ4vnPfDyypDH9UQ
2pQW+yEJ1yom2SViGjQSqJahtrhtFF8ANba7FRKermqIQH/nFopkyfT2sNnWF38A/sASNuECHIpH
ewbKIMcQRf7hQqP92hURBXohWVcKdAMJ8HdNFt6FnNK3ENADCKF592I1jOY2IoBTu2kJe87/3B1R
OZvO1mLri/k+rjiRBu7ru0qf2GmGTX2XZjD+lMmmEn0Cilb4GdLj8yp79QY5vufXbqwlI4EvK5+D
yrISAAfW37wyNqUuOXtjiequdmAOmNWkaSpO7jTsNx29dhZSxH57cUowrodzZT3CsTqxtnmsF/HH
Ptmns4kaX6KLTSvQehgcSSwDc+zhuaXUw6ftRsi/wc3MZI4Fqp+cf57eGX6GUqd7z9gD9Qv7b9Tl
T31RqaxTk1rKrom7Zw8Ini3F1Px87tMdDlH3kU5ym+Bx9OBKenRRfeM1OJEKbC9Pzx+r1jAfBkkG
brb8pT9RFNnHYnFpQvP0HBCMqtTpX3vrE2+yRPt+pYvzBy1OmMdUhkCKQ7bsGquHnrNB64TgWK13
XTyzcaE0Yq7LVE/frdMQxYtaXPRBW3PpAWojmsCqYKb2rNwkq8zAIyKaUjPu7AeKN8jQaE7/D5UX
OKun+dXOUdL+F2oDB2W2anbeQxCo3PgE4FMv3+dosiJNz3OQGTt3x+3ohgqJS6bcHgFELYJ29JKD
1OjYzqu7idUsm6KmpVwHlOYgIqqbmI/xGaWE0KJJtSBJZ0R8QZWnxOGkBSnKjinKBH9AyoOd4Ft9
P6ZB7VSgaIG5Dwl8sMTaaaUxhUbeDLm3w8MlOI+BIcLIP99zvINWEXaK1A04/PtItY3xgir1kdNP
VLg+RTYUvu1DY+1XW076QATJrBf8INi9enmqGdY8/Za/mTxZtBeSjeRhwpQVMDlQc/Nh/FH+e35i
Np296kjiJK6481IubAChncN8yn7P+P70jnuy0/xbwwNrvwlTk/PzcSEbBuOEWCUQXXpMususORCP
3h02tbXhJ6BbQGYleR/SNKKYN8khh0KRIwILS+NSZvWODz7mRn8ScNb2SHhzTFwUh/I/cqtPDXB/
dLKYVaUUAC70+SY6r7Uo7oLDjfoIVU6t7gkUrrAHQ455NtuPQZgMNBEuK1piNtXAyeUE6H4z9Fkz
M4aN7H5XVclM9/Ci1sq5f2kD+Pts6BfBMWDHBKSSPEGZ63XVag2jRnYcGjMoX2oOdofc/14T5cPH
GykmaDaX2W0Pf79S9Nethc3npqAlirRfYws4WQfGY/y4a82y1z5scgOE05Y+RUdjbXEtn3KkS4RO
k7sLTcXKKMH0424BKMzx6nI4Efbff621gEx08hFbs/Ji5tl+GtSLToJRRf6LuXWLpgQ7yW2akHmW
sZuzYunUJ79D1WCws37d8gjoClm+v0ot119Ti477Bmh34zRgQYZV37v/aSRpLKgh6XEEa97BK40T
uLv4OiCJbgZOwEdr0feeat401VcKZYas4a67WxUmA6hm8spaj1E1ZQL3Q5DrQzvlPL+pjqXD/c9q
KgbuXe2eRk3o+1TlMf3wdJU+m3B/hs8XfmHInq32zdza9jkcE+3y7/Z7itdxD8CPYYyyExp9O22Q
dCL+9Hc3M0k/o2MXQiECQORHtpIHdLXpuenE+hRYSPeisGNtGiCo9P1ET5EUOp12VjQPlPh8oMJr
svdPWR8m61alXmOnmnTYg8/WxnsNo5kKxd2iPlXa2sSS79+8sTYLUFzMCe0ZXgDBt9nybodu8kgQ
lrT3Vdk1VLbLLUujJGBQpDhFCSzoO2ol+jPSLIPmvnbX3ttAgPp70t1wrpv2zgodvtegBMGl044C
w3FFj3T2QmAWjxUQT/tRCBo4oVLJysB21hITUzExkBGhYORVmkI6Ar29qi9OqKbE6xMtvcOkNEsV
FaeFDrbPxXUl0ecd50k3OprCGFCWvYcU4VuJ9L/oEHQ2RtGtiwRjW1lOsWosi697wb4IB9JUBbIm
jR+e9VGeou4m6NpfO1pn/PqUHYa0K65FGKh9VYafYPgFaZ6xPHmAbrhme+ZIrFpvr8MBiOAW04KB
Tt5Tjlv6pIvHUE0zGsg1kpa4nIJzyuQKm1Dr7UX1TmUckZFRqZRIcMTQv/467QhznvOaVvWIlGL+
dNfHU7jJiQ3lFuQE+TM9U+Kf/WkEaFDIn0II7RCb8V8wRUQR9MdLB8NglNX1RiIaO0kdpo+kkiU1
frsMET/tIFcFwdsy1e07/QE/4EpwVPJg96EiRvwzzliE5CK5p9nBiQ9qy04KzN1fIYUnT8dwJxLI
NVcDvjsBuQhWqH1rvM2cF4rfd6GJ3y5RODj+aPOxteZDQwnCxdSXmA16QKcD0GDYvvv8UyA54Pd8
judzeT/s0TOp7589wCcC8SyhXdHeGPxywx5ND99QPT58P+jeAPmERMIJ4gUWTVtpSw65iAQLXr7o
8TOEppSCiPKarvWclIw2AtYuzKrxuTNMWa6YiCongjPpKqs29Z08iE/q5NFqxcL+mqhDdoptCle1
70YWtBJHffUViI7hiTH1O7W+V482bgI8IU4NOGde9fvNH6DaSW3OQhBQXMXnhBdAOBTOEW8DShnV
Cyeuw4KGI4L4zX+JCNDdAC2acbGVZJnXNPpF+mSsTzXotToub/EYxj2n9pRXOCznnXsLS3v121qc
akq+a8ruB4B4ixi39e6/aRLtfZYQbeIZJR6AME+0F9n7LTUCHX1NKtijAiSax5TPnR0zPmcNX9Y3
LeSnwqV175nYeIIQYHEcptRFuO/oxSD++lEMDEZjpvMl7bD/qmi4SjjT7WU2O1t1UdidS6rTI3F5
I1h6fAdr3iNFa9Ftca9BraFet/pPmS/OAGdCXqZeQYVrK1jdpfhBRH7N0MCXf/tmU23WCu92VWFz
KTGqSWo5fZoVKjekyjnK8gX6PnmIy7xw6P6KdsYnA6o5/rbOD9XGsaimJ68jntPhD4r2/i8aX/oH
jBckhBgSXwVyR3gW2rF8rkMt6U6Bt5YXOeWYXTablrrMhtzDxaSLnxyLFfagUriFFzcOyYz6V9R2
CVNCDe4kPYDN9+J+x/LzG+1OCN+Ug28dcvHWQvNQUze/txV5umNrCAUp1nPWcyZ19Jqo6eMm464J
IW6s1c2lSIsjToYG3zqd+AfuShoTW3s4uVBw9ymVKWO+u+f/W/8v38Wc6sR3EEBYPgVgoDlPlYiT
q9RHxLL4JrXfy/RaIRowHLEwKAMX9xRc29Ni5NVPvsQuszsB7Y4HtYtdZ6Hr2mxlEJYFNiocLcks
HVD6hhx0l2CN13HXj3nBqMLDqvO55S46hwLd74149WUSDe/T+O/qSMVAPf0a70vUlENJfYfL4wMl
ajG/TJFd4y0DES5YmQW5AhxDyOo3CPdw2yBe4IPZ43lUZYboxkXo+UfZ9lrFEFW8xT7zntdHpKZw
xg+bmjjdnzen7Wn40IkpovfPJtIDFWOnxmjtsGKhWIGGjMMTBHppRbDfA7+3DB9KNNIg3WxAzouU
ZXOxRH3ToQQuGgffLjiEdsEc7rCBGkNTe20vrDD5eG03KxOH/w1dCBdkFY1VQlJr7jFsPkI6QCTx
feflZKNt8GHjFBZ6lkYDmX3dDLokFicsqF7S8dpop0ZZFJQf6amRX5MT7fiT7FS5bDH1PSBC+H+6
lOJKDmscLfMbW3oZev8LVrrOb91jVXyjCdirh5kgyjD5rubNUv5bwz64FY6TAeZuWQus/tVpmjXv
uDFqazgo9HRxTJ1Ym8Jem4TAReUVEfOVFFSh4blzIGuf3Lw4Rb95FL2oklv9YBUTfgFNyBF+NsF7
UrUM0nCCV8WX6ad95G/LWzpOR1O+JhdTUKUm5RpSha541/BA6mdTIvC2mg6mTug+3c6lGG5QjY38
CtrBzBCvj6L5IMRys4mUtcJlLSOPrV1WxT87bEVSZaX/NL3gPMLkRBso5WHQbSJ1hq7RTamhQZ1k
01i6FClt3kADAqzooLAkqnmv8zJ5F81Nxs29TY6IffmfRHyJ2ocpcrokugVrVXvbbIwzDJ+qmGsn
CcbGyljhgl4GAp44oLmUGPKAOI3r5i5HTmO1aDCSqfoHuivmiVnOFmVd2bNS0U0yy5PYyPivkwVc
fH3s6VrOvjN1ouNcGxwlLKEPWegOfaxOxRkionM/aeT2OrvpHMVQfXuhOfiztZafjMPf/JF1D3zj
WpSPOsNvIiqBKt5CUwFSlExZeXgTPm31diAP9aYNgGhULEGaBx+uJUi7XQ2mmUkDqMFRzlUkJkv6
dgKX7h22RqSIv5KgCYfdycTXgJIcP5lnrLZH1hYWyUKIuTPPGGqnpNYAhWe3z9WdhYCWOXZz93Xo
S9HlnnJTZWfFfctueaTxcmuPuAhuUaqt6ohjNK10i2hRt2RS5qgfbhQPF4BAm+akkoa9lPFCktx3
RecVpDmyG5NV5sXKv+IM6whVL3eT/EKA3ZIthivJjYJMkSByq0JsgnwWMj04DSZvQ+zCeUmslIJv
lgs39X+cHnAnD5ewu6VMeQMBtVCHduE1axPSRD3j51kXIL2pNWaZnEbnko07OmkQyZQANdWW4bs7
+skhShmA8V61rMU35r5YUJO/rpoA6XsTK+MfBoU6TFK2FyEz+lAcVFaR8OFC1uuYULGalmcBcYmw
tr9PHR2LbCWRSiAa0Gcxx4YDWpo6OtWKpS1UmmBSenEwukOZDTGCBXMPrNPV/Zv8QhMbaXM2A0JE
ZUMRzn3ZAkP99FpPouHFhthTit3s8sddTS6HDknsPWzhiyuNBWm2DjrEne9WdDOKLQHFzhIpta5J
h1QfBk5Ki5czv312ELesRf6U6YWT3WybMFOpP4B+5IXaS6qQxWkpWUz6e5OqW8+9Bi5GT2l9CH/U
qqfWUIHS0SKxsFYeNVRSG+PrEGEYU31K8DBHvL7MS3gMb4EVSjv7CDRA6CT6ofdVB4LOxBXDfc7O
G44rS0uhJcu7Ris0Z2XlSdErc47Q/n4rOzYu/pbjl4e35kvt2DPDRr1P8K6eTkzSlTbzNROeYOdP
bJtHmnjrrK877OpKL6FNVNzaOEuTQmPrlB5z4vOKbBdXcx5cOjmrfP+k1Po/jnKn7DtDGPhgzFtx
boV2EUD42RUJNy7R+5LRzBWZSyZ/TwIUvhcNTYwo3xxhng+BkB5EmmaDMPvPBOzCI2ZfszdAKnUx
HI43TRpkLbUPSw4vmXYNiflnyOklITTuBVmnMbo+QGLEJzUQklzAk5by/2IWTqOnOxMgBEl9u14O
NbWFDYTalC0YJbhPvDKiFA/p+V72ZPSx7rPvYoIpUJPvDCWvOUBuFmQ5+7jtzQEYOnurPijbZGkc
W7Zd9NRTIZ7Li+avg7wtr/IazFRKnYijtJ7F2V+Mo1R8vNGg/7Kj7sxWthc131/AKw+PKqBBTe9p
vqgXoOp4Kzjuo4bdq5sZEwYLi7NmyPeZ23fFS6hRgl+2n1G/eXzM4ypqWxw7AtAAmIIOUGjkYA0i
C63jm1B57GFexBJDDCA1oAWG1OmTlx1hcuFpDbENqXpp7qn87o7CiPKegqmgs6/nCQnwO6xgLyug
9GLF2iBKWpEgY40QLk3d8znbm5fHk3VnaKUAOMg3Oha9UFBfPUbvyrmQUDWXIcK5BEN5ZkhD+tOz
yyp/tGRisLmgwGP6VopLqJTB1reHQQgedMnghYrvhGbx5Wn8bMBJl+WySeVofA2TjCnUyVQVXEq+
g86skejF4Qkw4EpYO+fHOIsXdrGRIuA1e8ZXl/wwzUlP2FTU9ygPaIIqZGDFW+aPXzSYOKqLS+I9
pt3ZsH6mSEx+sX5L8we6wIsM/shzJYlP3o9Kn0Ti7J/zNivYs5C9o6NqBwFxUR3yoe1llbe5BSEz
5YGGWKN39Q/ZIdrkRvYENuL3sLrrVJHGXcwqY5m74RJZC4O0fa+5ptScpjpGMnvMy5jardFzJFki
cpYbdcnf56BmL0QO8fflkdQyb33lIsfrkG3aLxNFWRyiXekOQT5OjAaspf92zkVRNPauO0ENBijo
YNuKluFmWzBHajl6gBsSJtU+JO3f95k4CW48+Zl0CbdGZnP+F+x4JbwByMxyskP32Y4psXrhIy+y
eBmWHtwGRbWfUnZoiRw+QBumWlBy4Kj/Q1ePn6aIuQv4DnNb5yVwKf+EiQwERb/xIx0nGYQP7gCb
+zygyBtMqiNUO9q3fLTDYNUPq6OtLIgry6dQjYCDp0ERNIr4wFkhddreTGL/CpAQguNidrm5Fhea
0UV4gHb0PovbxOcxH7Ao3rsIXkQ1EXtULypceqBliA/Yyfn2dt0+6+wB5JfFtYz/wab5Shvz0NFj
GDJ/SD/xicpflEz7C73oElOmz/Plbk0w/yEXRwGMrsiARlTRtAye7fDOkYY89METW666VbphQjau
3NUCDJciH0vtTOliEIQ6DBCnwCTL8nDqYgjBsNI9NxzzE62QoPxIG1ptYzYLxSc9p4KYRarP+OFL
nnvQyjYP/i73tWcp2gzZTeC7pTeBbLvD2cMj6yhleeNapGw1O6ufNq5CPTXnUKArl6xq9Z1dBsPk
qLxNEihMX02tHX84JXPkKz6ssRy53tZGm7RHfZeXvGA08ROaNml2aQlUXtbOZMF/BJmC1TUTZKw2
dwe803InPa++b+5wYqyAoP9dkQdNjx7r6a3aRvCfUjz1cnZ2M6OZLtZCqYASxzKw+wk7s5Tf9d20
hLt6OOaZ9CDhKzQB0EfYRqSVeeuh4fhuDItxHyEwL7SdyH+biPdwjitkFexjMBnVQN55OMEOOtTP
Zp2x8LTuzrgRwjbeHKq7Kd9J6MziKyGkPM1NYZKkIdcmlwvf/UkT2jhPsN2Buc2WI8QlyFTqpNgt
pLuu+DtPR99y4j+0OV9a+/eX1BaXPEdNkbjsO2JD4aEF03M90lZ9IBl3BnZLIUu6HHyDS+hpThIS
uFUiBOMPGfjWcLgySkqUOIgG1OY8TK+LgbIbVllxflC5txI/nAn7UDJQ3HbUf6cfRYtN8gVBoBpz
qvisEPq4y0lPBs+fnItxWew97oVRukMR+VhYNM7EvkoMzGsh14kB/Yldpso5Eg5oA69dczb37AMy
3CPqLDOpixFoe/s/isFjeQ0vSpTtiS4HiTeeyuVJoOadQf4bVvb509Prfw+Non3/5EZXmctCFkZo
IrhHG4PWtHOwIo4GpaLRRwyP/x9KvqQqOxkQooOVSRyq4v85HmAtUr+BLjbWL9HGAaKRUsHToNoU
MhQyryjx8506BG4ZnuSPFQjoivH+hqyY/RgnSzKJFvNGvwiblwpo6Bs0CWjLwdfwZ2o+Rz4VmqCY
4TiRBiOvFPFdMAtEAH+qCuHvGFOcbd0LuDBbyaZcdaKkZgvBx4STzALJXUzbuFkEivB+HEV25vsM
s1u30y4rNrqH371f65I4coD6aml6CF0iwaYbUCRLli5DdQDfj8X1WjnmImfb/4+HMIfA/ik/BEum
6hbD6d/EwECCHr4MJ/+TxcJ8JbBAiCYYB2nM7f4SatBaohGWYVJmIjm9M78inK0IXFau8TqytdfV
zE3g7XWJZzbq9l3H5N8K4+CYDinAUBkkZLcZKVbQp6zh+L5ysCy3dTQZhImc94AU1tOR0Uaf8d/u
aYK+m25vxutPTFPZ8vMxWFxOIfjje1eNxdbjJM90hJ2XVzuMOfIMEXM6TxGRVj2lDuYT+mY318g4
0lNfV/pebUYOBcpAGY87J6v4gI3Zwq0Ddb9HiXpZDssdwpCUNAb1evvMlGGzptZfLJcx0xIDWiZr
1bt6wW3xQXHqQJ8UGgIoqgANnHQeRGBxdR/5XJVpDll/mMVYZRg5Brh+1Ta5SJmLo1fcLcXAbnSR
1uG+t02mh9lpXJP8qrjkxdxdhnhpHdZ91ahbBJCDfh4AX99H9JZnAOBRSeE9X7RvUU7WwCWWgtc1
r0jZlg6zWgp/opAMGq4L9tMSKd9+JfKJ3nqz2RxQgmZGls1SQqpc6CwcD2gt4+v+Q1L+eto/rYJH
8fzevdBSSFHqMdD2B6yFT4Ly9yF+Ij8ViNpPeCa/DwP7xuFIY/4BmJtKynMSn6ddwP6QiDxNobYp
UJCI+uyhnDfkvn8wD3LWVLzmzLv/UbEyGrLgjBd6pO8mKjXxDsc+jzGRLYJjxZPQoVpevd1Xu8rh
52da1vnVkcKXzJAyRZk3tWiNqUa7Fa2gaAsiZXgDd0NBajBQtrh3Ekmagxjzyhl0w+vWEyGRbhdA
XYjSVu2OXJWf4YvwUqWhSiIDu/spHuW1cHIYgKEQv6lGMl2sqmG5gqOT3mFE2FQjdd+RYwqSqEtd
mgeFtNNWr9Da8OMPUZtPn+EoUnxG6JmRoghYzKdj8h0fB//JmziaW8BxRjHMv6Txz9sqDrrSI0y6
Vy5Y+/ICYnUm2Ur9oZqgZhpJJUXD1khht+UKJTafP5Scqimd+RgprWauyUnoVEx9fli5c3FjIVtI
RC2EZaXQK14e4dzygTiWPqWRoNjBPIo0kMJ4TaccNeWzxEgqVJaZfk/frZS19IAKBUq8Eto/dzWd
G0VlLwIrgS1INZzjQAWLgIWM7+YfM/wZcQ9XoTZigAr2YPrKZrTDvAxDG4WQO3tR3GJaC/ICeup4
idZCnO8Cz2bsiNPR2gWc/o8iJ9iTSQm/72Cuf//3Zq/egWbRNbrW+FY9hDF9oJNQuxh7cMb0WLrV
OQwf68Ogah26eZ/rGk9qOW9haIjyXQLnwho4d9J/vJ1aaaQ0N4NvT4sIlUztMRhv8LNr/YISQYeU
9P9KRRNW1AB0mdFaySp9lixKzFr3/utpT6hUlR39z6WvkTTTKyFeMZPNJr3zkXzfTmnRSQ7U2J0L
S5zD+QyhMJKv1mMSB7H8CGqORb0kfiARF4LuB5WadO9L3Wutyw+xaUstMiZaGi1oP6oSZgJZu/x8
NVdJCcBU3owVyiqd8uGYNkEUWVfcMs2lpE4R0k38yFwZDsX693Gp2wcqCYmF8J0he+2bKnrtDn+a
oup/lPi0mv1ml9D3Rfx3QECZzGqIQKLOnJqpHHEwDv2FEO290WATai/Sray75odypJPmYKF/EqrZ
3DMb0V9OWFuwEKZbdF5AWACoCRYt8fmTTWuxu4p2gF4mz8U/0prbVj5eNQ0FQHA24NaWQ1MDYboL
JeOPzWlIHDMT/mxOxF7+QV/vKRJoYyPr/Ajb4qjrNZeGBcUIaN8T6twi7yMCoze6wELhlBCzuEEP
LmOyz1zMgK19C9c/O/4zPaVSPcu33ZtNw89rCH39/n/XiQi3f9ovlaxTXNwUveMN1jWJ2ex5KS6X
NQF2yAOMeJQwbKFicOeE2/AAtuxMHhBQ1mWyycQZovcDoGv9BuUPx9g7ktDQ0blfWMZI5K0aW8h+
Aiv/oOKKbC0HXWcaBiuAgJrXyQqakKLB3GS60UvNsJg8AA2vo4obZD32KwW2tU9FzDZuE1S3nltA
3ZGyK5E5ABYd/2IrMj3ERx5gt1gVtB7Q6gvEQaU65PM9SSTcm0nZHfO64C3HDcAO7HIb7/nB6rFh
9pSRj2ck10v751OvvhwuHg69XuidqlLa5yEdB8lDLqwzSATI2rcRFaI/3YsYpfbWHc/fEDDZ7B5n
akuKVX9rULfAOxtDun2tkJusIMhhDOQmlJK1RV3EPq2BF9XoAj9AKbYiownAIDoVPCEHf4jLJq71
2ZXWydkrd6w+1pPT7pXz7xoxzQqfMc7RVg6H5ckFhVWo7OHb1ACMa1Yi0RQ+MyMNpJxWjExF7m65
61R1x0QhPGoyZuxKVLJdwS3GaEQ6ib8Y2BjEHaar3YGU5+FCP9YTx7SW7tEA2IFOeVTqrqFHe3Qj
6VKHCfKijmPuVrOQSLbdPoxPG/v9TYcCIwcYPpsQ6zAtTETjLWpskqB1LFAferykzoUtkoICB7Xc
NECMqF7N3jAl6EYa43C0gaPKS2ZcXkA4cv9/COsl+v7Sbx5kgMRej/DcRfHfS5yVjeWKOsH52rCS
RLg5Q0fb7UQFL/NfeDxQSMvGAcmeaIfYKvGTdauRaahfs3OqKgvF6j06Bm1dwmlwHbFAw9FCstJX
fqccrluC1V5JmP31IhhVLBEWTxrWiZe7e45LsEE3vAcyT0OHwu9PfhKvqPYP54O+ubmbUPs2S8u/
bYOyE6NLkpR08mNGf9vohsp+YrS6Hcl6JFENjiO+/aUomId1VkrRY0/iPNHBhxIUacIk8eB2Q2gM
T+0LQu8HBfv2Sefkmhug5V3Kd9SRsk5lIAJIvr9j7j2i8jFQq0oDnAmv74aDspr7LJb0fa0ogbxo
EvRlbl2mjylq+ivjMf8bmcVgeO+P8E21UxUtrrv1wavFvwVBux12JlhtKklvXd0/oYNMPdSTmB83
0Z7dQWbXbvyznVohMoG6f3WS3PMTPoCw5slIL+nHw6cV4YUj45bQPlzjDkfbkpG3vooWMgWM0VyC
T9iW5vXtcdwzWRtZd4P57YLU2H2ap2NgTNaDG/+vchNIxdNv+x2ZhlN+86rQwxcCALLBjtZ7rB/1
ltrK+9MkbpzQxYhJNOMZ9T77f/LvwaGiJRN08smzwzb0NyF4XHEbwsFArDE+yJ0ngpCusxeHXou1
zo1hJnaP5QRTDPkvq2RUagtf/rbzlPOiiDrscuKOli7PuvTU5hvy8knddndopU6CSIE4DKkI2pqh
pu0xl1TZhqizBtVQOx3pZ0Ed2Re6bKECfrS+mw4rvuhNpl1nC1qXtv0WBgRcdiNH3XTSvGDzX8PA
a0TKoRSLDYv+0jiEnPATizzNxv6UxVVexuW/v+w+wL3+xftT5B1d/Inp5DZN4ydScc8ZGo2+sEF8
oMab8RtX3U3FCm6R5+25LcFblYm8ulgs4u85Uqp0vnieN9Zw7Z8X01fm8rPhYUvvkbFsEUeLgpwN
GjbJsDLLm2Sgspg1TrTX4vzx/64udVAs0e/G95K7tq6ejlOSkmW7SJFm+65bKEd+nzRLO648aLwS
2BIsiySdJcpe61DnpR9hMJzIUpcBwizUOq4aMzC2mL7Ofige5ouROSTVYiFPdK83X/TRymw3uvmW
01X1uMbIk0JKin7gcU5RNpemEZ1DQCoAGaMHhHGr7aPDqW42tLz3CoQfkl/cVpoPYZ5V8ktL2XmX
5I6P3waGePLCDM1OQR0JHIzeyrJCVLCWevY6S4R7ekujN3TLInzZPpIMGPHiXewX3BpQLgAzxJMo
1rArVk570ZBiRx3O1yCHV8vLV6Mm8mdKFtNqrL+PEn/n1fZM8Jc9PfQ46k318cvKZEuKsRz55b4j
oFNGNa3Kl5rsq3rTdvJAufbdR3fNlBq2tq0smZlWs/m5S/OnTkALZxNDGAohnE1GZoOd+2xaaZUN
PSAQi/mO+1mmrAFsdiz8GxVoer5QVAt+m1d7gHHXLPnwgkyO/LJOWLUFs0g7PD7Z2PFHB/R4Nu8/
rGFIiLkAkNvpQy5n94y+B91VzwYTYbkI8XZCARGDku8ca6DQkaTFgULyLIvddBr+SCbdmFKaNC4+
xE0YkuulHZC3kmRZ1Z3qwoAZCJNgaDsDCknE0gP/1+VX0t3ESdeyLX1ab8WgL18iEOTvIUqDYNeO
GiTVMLUahCQvrzXXcqMpJg03iLDk1MTgOQtPVSN/BtP+sXfjQ18tstusalQJPJ1RoFDIoofUhf3c
v/6cWAl7SbomTwyrxFGzHaKb11CLhC9t2SLKAxLi7lrzIQkOHJ4ULdqN5u1K6OEYUDRCzcsL0gio
t9WOYNxBzDsqjIhY6kCEpKlWwisRmpcDqE3CqxayR9tH12xAf+zbAIWi/0+9K0ABPgJlN2SvHthR
8eMh/NwIqlxK9zVHcIPf98YR/B73qM2LCCfOInIe5T+vUbHmMhW0Tpdy3mk/dOOSfW30KJ0HMQNk
3gNMAnLOrh/SEP03DezR+5chn2xTtLR1KyRs4kThw0YCKbqIXrD9zA4vLjQZjG6/WNXmvzDrBKtK
8qMjGO7ik8KiNgq0fElV+EwK9a3aKvQNbR6AhNWusXOe5699U/fu+qx3+2wo5F67p2O6LXE7IPX9
2tG4EMUv+wipHBbMy1iL0ECDoljloppLh7sGWie8NdDPwNSei2I8h4GDey0IDXs5ndY5eyLCDo/r
l6P6w3MTx3SfJGoLYaGSL+AoTHwaCwaQR8eKYnzzQJaxKB0UQn7u0+a06YSdAVerkJ2AAoKgig6a
3+j0ITIf9aD/Ny7IM+X2T++Au2+f/0EKMxOmfSNw28QpyGjtsl43uNydhIwJpuTJ7Z3sOWmM4dRR
LgPdg4pXS/PUAiY58dtiG34HjE9OYyz/T52gpapWt1momV4RjRdlk4lrbO7ZpJsMly+ZjYs7VhaY
7CcZQoT7xMOAPQXbjMzm+rMABeBPaK3Cji83fiBx71a7pRuCN5WyVhrB5VhlNFr0kHJKERE/pY8O
XLGj91ros4+6H1bSL/d2jab3KAisKpuyMdMGP2sKS2gEqv27dxG0MH85SqPVvuwStj7VGs6fnf4G
pcz22dRFmq9itnXxmSt9hVXl7WO9XgV3jBe9UldnA2RdwuEiVxYlfBZYhlxvcAnCwPbUK/SOE6L3
kaPu/LYivoUBNr2geWtUSgoua0J+z0CKJjnMHDItUpO74j1pudNOHJ/cZk0NbNOUhocXalA0GUiB
aCK98fYDl6jp7hh+tj2IcjSRT10vl7xYB51uJn0rHXTew3Q3uewFwb8KO5TcKrfuvF4ev+0T1vh+
AhvGlEZP0/TKAfxQ1op28+KtyQD85C9c9kfxY+Q2Yu+Rpk+bJ8UYcbKq+FQrqiEdyR5RbGNW+Coc
o9k6+uR4ljJYXNPhg0eZyHwUAufKWb1Ka6M68zl7Xb6dUTLwyP6Bk3G1gLliKuphGvsRA2LIaRv3
k54UXoM3pPmxVRpAr3NMfysbhP/8ZOeHl0/oYs0QA7Bjpa8baQNgwSrGWYbZwmNdFJqFTf9+nk5H
VYclRyCPITNTJtACJPTi2rKH7gj1MZp51fYeEsAfnDf7CeD046yhT8J4Y5/rInhUMbUxC3oUAb6D
qZetjhjMoC0EJsiF7k3YD/lyNAez+hMG3vqdYu1udNsBOvWIqpidNND/+hjogvY8Zuq4IQseM9O8
meEar+B8S7KEK8DIj1Ywz6DqOjao+38eyUOqpskJzEPbPStQ51zA6SbJD/Gv7Vw5OZby4BmO6QmV
MD6hC3OVGBlKtLGWjIBNaZWu9xN95zCPpgZ/phF1MpiYza8yhL6vMmfG7ZucaQo7+Tj12Ioj86b6
k+Os0Hb7NsOMMV8bNZ2tAksnj38SAtWzz6ldQTt4zrhuzLIRXQiHxJt7Z17PWypvt2x1n6u3aY6X
CM19fZmLfzoU0FmqaVa5godswqJUCs/skulOm8nPTotBJie7GmyqUXuG0qe+Qc/gLjKhNSGECzAp
Bt8MPb9f8z+m8GiRVdBAFXk32uLjm53JKaP10WxYWWjT/QfAKa9HCKr7gRC6RJI5RCgmkepiTkAx
qi0X/h6NFkKhmzm6O5aZ1VE1Z78WrgTRt1PERBJ2/T9e69m7UJ+/+8VSe7RmCmw4FzQxqIDQx2fI
cNQ55KpUM/U9bOL+ORUtCHxVydiHY25cAmDCImBmLlzjtAnUJgGBz/YixU7MQiF2kRiQW71rqy+T
DvcqudKzvcA0TrQl6mB9iaRRiamGLfehY70D+1DFNuTtPJb7CW8Pdq5SLNGEw1InEpkuY3u7AkHd
urQRKn/mIZqKntAh1lXPHLRWxsEomHhmT7FKuVgxbIycoinWNjMsyIHjjjQ8VUN3uvEZDGjfzevv
tG/psVJkLwvBv4gNdLDJwsGNFN3vQiobBd31uGX8n8R08WBXwDwd7cRVXnC+YYTMnRGJnT1Vdzjh
YUlHXThLFczwgCducR1pfnTjSP8CBCM59+IFGx4WPy4avJAHS6mE0LGel6StKh2jf60dGvQolT1h
dIqhvje4MHeqPLSzMS8t5xNxYtOwVyC/eTnR6m5r9s0mIyOd+0GquxenSsSxfCfvYfQxt6U8PyZD
d4QXLzjVVCR9OlvmM18C4ZIqFvlogc3ulKmqNn3GNZv6PkD+cPglrTszciOSfx1eRQAk8V21e7B7
4rqnU78pQafrUdv1aTwHX7EeTT1J45YdDfEr3Q9HpWCmxD13bgAg/Pu/Vq30MKhx9yuE36E36lgP
zfnGuA5LQDRl4TFBgToPrK6fsomMdElRuzU5SRxzI3ljvrQ6q8O5lysyUKNnoUsFswBZH7e6jr68
GOCT/y4QSEEKLgPQSMyZ5TtqD/xcrN2faXcHa/1G/4EB/pFeBmCA6e7sx9ecCJS8O6WWfrlddu8T
o4QWQH/FlRnu89Xwm+GVHq9wXUmKCppwnPicCWMhSZSu+MATSLln7ilVcroQ454RoOejyJ1ZySwV
CHHxwqRgRDDsQ8+sebd1mdNHJwOSua6yoLX/kPFjMjWlxHowHuqh5Ipr9YZxyVDQ67pS7s4fHxuG
/ID444F+YFtNWnjQVRtQ7fPfkXCkOGkbmhrLpxWQkUIjbUipfzvvqYXxDNHb4+eOVJRwCXDHfosS
TuD3DUuYrMUIfTDz9uN+gYOGABO9fsgahw9nkm32a7j/409Am6mmBAKAGstikXoHRAXa649OlHMz
Cf+siuws5W3AXZEAO3qcAxPql5BvmXtqivhyJEylHaH/PHuHRMvnv2+kF+GBXsi0nY0h5p82pcID
TKHTXuWAw9pdxdGRDVNVDo9VeVbXL3TbEDaab1AMvkjLIjoeFnRwZ4MHEaH103BYy7FWLM1Egcky
rBvxfWdSGHlsaRDUcOXytmvEEXBhay8pL8mYYgKS7UAzks5OaAcdrvTGzPk96+zN71CMzmnFwb+x
jQFVAUsn6wcGvaI48A7Bjq/kURV0UWXLNhnyrutBa0g78HXww4HSl34u6fkD5YfYsu4ohW/xylrJ
k2JkF/NPz3FYvojT85t001AVIWHv3hRPSulG3fU83Oa5eocxwvBPID9wtvhvL3ue5Yl16N+iNBJ5
eFZpzukL4sSuXZ4m9GzslU/+HywdY1vfRx0E7Lp/pspJ1NTiO/+wwWhDsSk23SrA7ljQcchUeNlk
9QFU1kgT0VXbL/3yLaiWnoTeUeVsOnJ9/C7scac7+m9s3yuM7907Xpi9WzDAZkcVGGCOlcIm4dX+
yvHyFpm5e9MKJAZ5p7+mybWljKldPUONcNW1A9LJBxm+xQrH9YHpsYMLuoY7SaRDRF8qx3Rp+Hfm
U7w89DatF7h8S3pWbaBsOMycKfpbsRpDRY0T2lQQwQwB7mYP/BnFxY7h21UGcHBLPzQxyn1oHxJk
6j4WhsIddPHJ11nyc2dku0RkgimnlexubY7oVdJsFisHtQdY18gtTqeFxvSie0ALtmxXFOPjk8Ca
g7XUlPDXyMlIZgVhhqzmRWkKiQI6vsI3kiRpUWZ4wN/Rw3v31RJR/1GuABAnrFAU579uJlfqyxJ8
FXMcKyXft32vgxuHkjRolm8/c6om5cY3E4pFVuWeCiNb5hmoFXb6PdKiZov5JKW9BmPjZP4AtM98
jsmiEJt77NQG9MNYjKKRWBtGoZ6PmLoOnerF5oGwJw8gxqkg5AByVeKM3QbBa7gxGq0VEblMnJwl
gON5JK9h/R+yw6S+6mRa9WJBkpphMXRmN86QvMwDy+oRG3QVYxE4DHdiFCFBQZUZmm+eoTEd+AkF
xuX+IdntOS1SgZ1hoKyX3PGTkCrnGqbXi0IsqH7d0J1+j+IMoskk/dylhEwpZkszxaXPx0nkDRZG
+31EznJ8/jIyB2Y4KkqgnGdxltIJCxk21tlv4vTpC+UadMQS4SEwerBNmJvEdo9YJ6Ux90Dh9L37
9fDzRQvr8miRBPA9hwpbL3UNEL3imqgCAqBGzBvVVFBKaIu6Z+pqMONrdxz2Ch/lmIQ1YWhaxcpM
8qNN2mK1sZKIV5jYLWdmivWhZ4vcM2jsaAb6XIDL3Y2AIDSu3oE+oa48e2p2cFtAtl0kdyTqi0+8
edcPFDn7cvWYsXauvUf+pibZFTkjGBze1vDLIoWLF4mxrpcjAg0S/TzXvZsDhOnzVHqZXvkB2q2m
vAahEEu7DtczA+o4SRFJq1koK69G+F/yt++uLoYnRySBeALum6m6weR0lUQyLFsDgQrCtcX+XRSB
xOakWi9bSB/kQ261Ahh26se+n9P0WwizCuOic/Bh9Fy8HYi7FxEFnSNMetSe+cr4pDrlogyLU9Ux
pOIBDrn8vOuyeX8vftbsVSx91P7Vd0qBD+n9lF2dJQ5z6gv2torGIs5If+2ZGrWr3w9U6sgjAHZQ
hY2EeOIN+nBMQn1MjT/O/DjyNafVXr+pMcUQ5nFl9LUdvB6A9byw3eZVD3Gw9sVX8SDTcLDwuBqX
cANVGIS/jy7YdbO//S1jLQqDAF0HeWsFi01SduCDd1cmj/ww4vE350XaVtbKEIy8bV6/A+BQKl+L
vaYQ2D4FcwVAMV6VIJMvV+jFuvhZ96NCRsyoMOAS1bk92655MFxrt/6lUSV/kcLT2cKQ/463JOwi
DP5RTmSOQxeWeF4obNP/IT/S8s/eE2LKAyDe6160RF+71h6zdeSBg+dGVFmvnqXxiw8lTAzdJ5HJ
RejjlBT5nlyUGBil2BFMZ+5s0p7hoz99JjVSfjFIfUiMzsDWePumLqfnDZ+HmGlCoter9DTWTSMG
3LV2NnQ58q0RR1OfarR/XAEM2Ya7ZLN3nEdYFX3zcUcP029QoX/SUlx6Drfkezk0ykKkuJ4eI9NN
/I3jKIYrgyDVY4/uGJHUlp+IAAGNX3cEiZJXAoEQ/3rwp/v64rpCbLkBpc2qfiHBgCUGO5LUb8is
M/egePU0OBVd23nJMagmklr+2CgFqbmm0Ngx8iV5hJOxq39tGtF8Eo845Oki/xN4B1owG7oLK/Re
W3jmW7hbXxneKXHODizasDHS133ppjitlvINCL1u2wWUjN0NpElPsXtcodITASHZ7BFU8GytnXS7
jlpjJY661fivcQT3hDxLSvkU9NNslF0V2MukWTc82YAvkyyKqZhcT+v3FNPcZGd7DkSIrt4Xr/8j
NDbFAQD+rCOg6EAuQIxthMba7DR8CuKVmiYq2GnX7c2H6+XWDwot0DQVEoAvEQsM7+MfzR2BQ7WD
rX/Jn/eLqf76qSwF9y/Lytwb815bKduOjfv9V+jzAK9HtdrKr1A7k/+5kyCnjRRIa0oCYuylccWO
miGbrzQzxW8DLYtck7GEXcCzYpunEcXSouAHdg80pDkODKyxR4+wpzm4Q1gThG7QmeMKwH7yzc9N
wEa5wZyKYkCkv0FppV+0LJ/iu2R2QUSuYcDqych3+DgYH1gIyjRWsUNhdCbvSpaEX421XUPUwDhp
UhpoSHMlb7u1JM5+pxUwacU6FWi/pc9OWURTUOj6rkYHNruv/N+7WVrWSzDXnRa4dc1uSh9aaEAH
YM7XLO/im2YZDigtqR/psagTNWFrluI95PCiCM6Li43WPgtNWMphhD+ZZoY7Zed+SYeqTo5KZZiL
gzBdrClVZgD4Spt6UzH/wFkVTHJg8YjJwb/hIeS2D4zrxhuGOONgZGPfPXm82NL2Lao7c/DfngzI
jRiZ9DntNu7jpE3TjZR6L68J49oaVFSx1Ad+ZyH9Im2/vbNzJjntwzpp2pBxESGHZrTtaEf4BowP
KPzY13+byGbtk6PUfWfYlTnh+y5XHFXDkfEpzsRoELYYrTw12D5sZyJrnHZ8BAWJGMquyFZSbWE6
yfsPXnDe8Y1wxJ1mRnZ5PDNFxwnsR5BEJX33NNuSAbbgKdZ6hPGj100eYW3uu0l/3S7KKWboFSxR
DVVAyDVIj2EjO2Gq8uHFR0+p0oc9tJFW7hnD8wDl5HhRUPJ1rHBLQ5sDgEQ/kFUOUVWW0JVKnoT2
Fb5pPF3PPyu1Urz8XB4tshTdYjH58dwPYH+kH/f2xDho8eOkplwJzlnzWj6D85X1gjONkApyt2ml
y6ZVCjmX8AS9dCMeF7hp3fQExeShy6m60QusRddfnD/AY8KqcRJFgljULcRl8SgidvLrdhOGGANW
vIHvOpygaTnjmNJMMl+Q2QWf/h+4muUqqEqDQ/7Q4J4MnMpb/5UeTGUUuvGTpOjt0HDbEOv1ObO6
N1mBDJeGHB4RvN2v7AWRgqShG82sXpAJEGO8/yi5rTjCDMl5K2KO7xEfkPlax/uHOPMN/jwX7RHe
S7C0ngVhx2ML4KbSt2P5og3els9syiyCmtLmiRrY51q7D653HgAvD0cksUHzZI8Cns7U3PXcuf5k
O9E6GUkbyG9FMMy12gx7cjNSXYJGso4Az3gWuVxkFo/XYa6RG+IYZ0Y9d85ODsmtOhiE6jQFc9KP
9KyeHtSscadQV2MmwOQCBGYMWMWOA+mFESiUrc8Mg1LmButJiSL4Q1x3z3/p9vr5bBdYOfrE7ZZx
dc+X1SNPF4PptBc+Dtu9X52utZgl0j5wfze35wPPo6wtR3JTR2eiHaxctC8x6lWOQ2yJnXqs+8X+
VJlgfqBaGbM1g9Zb90ytc2+897kNglguIMtajHTuGRst4U+84zK6hCeSy/qeG/5ZPGZtHLpJaQ6W
h2M3Flzs/QMUmmUBamHnCYtrdoBiHKfC5Z3jj9H/tDi8zl+UhMbRYl754wGVlayUs5tGw3MQ9FM/
kcI2FyuQrrs2D8nQa5vRG6rHI5Xo8eFBzlzpEffRw3PER97usfLb9rX0ZG18R4LgFWp9zWgweVtw
H/hUx3f431JF8/TBphaweSJk3hsbvC8BkL4cBLenIwLI4cn25GdulEV0gWrjDa6NSTN9mosycceD
GHCu2dcweD2skI2kTJRhfMO5Z3rVlUnlRYt8G38EMPqP+Lg+xbyKlZiZ6pAXv0Op6SQQUU2sEH3P
ETRWlnKyjB6ZNx9B10BWKXMsnddiE7i3aXMJ1jOR2kdC3ryGkt+AwUaiWL1H+acOgtf0wtGwZN6T
0FXbMJrPw8vKmZe0XFXyJmSRoom5yEQj0ZI8Yzn9N1cy4mEzXz5pRDjVcC6CIUESIqWrgnrro9I8
6QfeHKebPQMmO4Yt5p70oeCim/E9mddlB6CUeE/jppK1Ug9NUqIFvuRssUdnDqvn0WJi6qmQs74b
yk940qLm8+JMUKn8pPshXqjnndLpVOmjpDHlRjVrsHOzHGn8XZd3mTMVOEwdSjxnuGhdPTR4A85n
QII6j16TJB5PIei+ysJXN9MKhGHMduwOgK0cflXoqFPL9UxV27izUzWBeMOeG3dfTsl/61rh9gXJ
Jt0fGR4QHCTRf0Ded3gdLMrYcxegBlQwBCwDnbxJsVWGsbmpd2XvHGxulR9q9aB7YyiftfOtqGUv
fUI6SGpGj+nI49OaSix9tyvfngrldRFK3cbL6F9x79aWbeLBDjZPfrSrmzi3kFMcDI6w1ypAgGTj
N6CGnUSkqe5oym6mZMkCl+Xb0T2EO5jYd+zicbTGTBjX/4+NpexzrS53xs/VCZ4VegHwYkykwTMN
N7x7IJLBhTqoYO8ag3FDHpwmKvj6TQAfGb4Fi77aI/hVYxqN2xwMTtBK8Wg7QZ3jRaq9YdCqg2Ov
2z0y87SGVOmUwAMcqulM/uNxaIO5DdcmYmla1rMz4rDO94tHRWdhMPLeh9Z3avlskHeMKSQP8jzZ
WGDm3KX0QB5CdTwVo8WFn6P7llMIzUmWK0hjQL7aUstuXsJvkXRj8ImkkVAJ5F38nwd34ftKtWXE
lBVbCi5tfmJkhcsZxP8ACyY0fUG9xnRB/VXLIfGHPCWELF05OBUcZjZ8y+66QCfCeFh4cHV2FRTM
hG8jCNj2770apfJOFUZtXYvQEYBq6Ncf9/y/fH80rt/YgCzSRf1EnIv+2EGrf+JThLwEIHrTz7kE
285lxR0iPc/+NI0OSwDYVBPTShFj1jMTG2Mce9bG2ar4gRr3j6Hku5Tt1WfwhKYOXpzcsemmyfCl
g/igTAjexF3AA+z8oFmegwq6zFRy7dYpPVX6X55eOt2FnWO0L8ZjhMweo8o35J5AeLLU7Ff20Wo4
fG0RO1Uv8UG+96SxeLZ/PmcH3fgMkjeWuhjR8DMGY+FyGkC+yE7fWpJYBeQIOiZIulygKGWhVJGn
lFu8Snh6bWdsKbqmi3L1PLpVkk8t8+tDP7bGJJxQJcE77QJL0c4YrGyJtxNPYND0Kdxs6c2zCX3M
OJ44M/qCm6eTXOor6WGhwsgZ40GJ/iZLembu9xrq0sY2Xu4+qG1BP7YCv5dKWdzM5yB34dyfb1Ld
aXZe8a3MAplU0G8It4aeW0zOGqvVz/yvu1s+PPP6hVJUaoUJDCD5QaUjl1HeJRB5+0y6SGN8SEy2
pPlE68hHYnqTOuUUa7xWxRU5YsftyL97ApFXg3YLMUGsT3t2/blnv7O3AK0sC/bxmWGAD0ckFRjS
A5L22ffjk7esAjrz15rHH+lTXf65n66lf5pFFP0ZuCEU3OybmPvE5EDr/dzUB9rJKhSEjyPzDQcT
KoCQxvLAwyhDuEmK0MQ++eWxc2wepbQbgFRLvbfSimhKn4rX/JVxPfHPHWn7obRzMN65ykjBG5G+
JJbGPUhu7oKkKD3C6Msg2MTJnxuc1HdEhts0tiB5OkafQPvqggD69Sqgyic0SwNt6zTLgojepTvO
/Jb9lOFyovJH6Un/gHkkeBIHzNX1uwuxsbk2Jzhzn53+We00DB5zsv888k8Fqq4mpVZshB1JDA++
ki5svuJhGWB1wvQQyBQWK2iB81EhSlRca+9OwYyvO87Rf6Ok8XGBLODlouoBIp8REVoNIQBp0mAX
KyZOr1KgyOMIQrBR4vThPUBT2APjGeJBRfgQZT++XD7vG1GtxxXfMNlnWKSj66QZ7BNuFmR3yqsb
zVDZ23QhqyFEmidTASDiaKyouo5Yh+gOUFZKbc0B0LqUO7JQ5uh/DO/MKWL3HYOzfjX9HIQzasNQ
Mo7l3dfDMk/eBgYjzmRk72Z5W6fmfl3pBAcWrux7y9dS1C12FfjtvPk0/Pdc8imWGJp6QIIB6Q5R
Gt3UpNfl5/3Y+SG0k8pLTqEJ/l9fZZ/miC2j7QxeD0aTxhg9odoQBijDtLSOOKcLBTj2Aqojly5a
qJW+Wv6ys3kqrlvN2F1AYKQBOrhgjjwo4YyAACnynrnTINJJdykqacZfyyHrDBVf+wL8ffgLShcD
nQEkOf+pClzvd4o7JppQ5MvoJiJP+nNiIJ2HY3wbn9HVBjhKftD7ePe9HnsDOWQkIzMz6M7ysu4h
utf+7noBYu2CtI1bQZ7xp8KaVb7/VvsVqC5PegaOtM+dfRDm3kKDXt+7EhAIMANYqA263F9wC+nP
V5N6F3e2Wkk+tveEVq29dheJ91Bp2OXEBX+V7rEoRABw+d/JHqoFkHlX919QsfDz4NpxnRPvWXHR
HmJthOpdLXCXMN8GLweFFIgUxeoRieBLWFik13G9L7g2rP7Px47gVXDP2683pTLej2j92IvdxZ4L
V9rlSszulajC2lo4aKfBlSKHKLlzV7bHWN006MDIRjLwhGlXN5FIqq3ngOZDxNjR1vhtZpGclcbT
ARz3IvqSM8TPmNZZf40HzhhXLs8pb4/dLTiwmj8NFtLVe3Dk0g0r042YxR9EflT1U1fNG2W/N70e
OqPLBQ+Mkhj2AyCFsrOddC7LcG9zWrmpMmS+4OrE8iLWzKK4wVWvs6B9GEYMDHn0EnGXRCC8mNDz
Y4Qzg0f7Uquc3H627cldkEfB1yHdxa+x9Wmk5CkRcSgmjX448BxYJNYuakLpEF7tdzu63JtE5wTt
Q4pEXORuc8cUuDhrebaGctsuNVKXTJMxGaONqK0pDU+wnpsnsLDgbkpxQWUOuCZhaNxavz3SF1hA
9PPfnCRi87wuYNcjSjvCA+2LYbKZlQA7T6lAob/R+0lZujSDoco88h3xAYgjjlDWnzwfd5oZgVpk
pMEecKXMBJGiV8KgYxt5uYMJxSdNJeG7yPJhZl/mI2qKxY7DEqmN1dAQWRlofkOu9bKh3eBrvPXS
aI4mDa1h724IlQzysSt1bW2l9fx8P6UEtvUqnn+wsoXmfAnkqkhdsaJ+F0NWCwwVcTi9QcjLyM6A
4kDW26Q+4OlnqJmyjxNvhQjOTjB6jI2oMpUtJUCT17BJlKBABIGXpuW5Rd2RUIOOjkIgogEGXk5g
5dPY7Sp+7pV1+vqZD1+EtAza3M9L6GtC/dPYEXEmhOHWqOkqSwj+1IKdkfnT+YgYj9U5x9Dfh0jH
YePrrA3AyssnpQbrqWM1vtQ4EGo9fV2mm+30Yh+RjkxDtr3O7Ia79rMcF+IVMQlNWPoYKTk9uvkP
IR3Y53WDHIX2WNzb/kxvmNJmTxv/b29bZaVSPXh/PShDa/oqhiknflARpUcA/HcOEysgh6L9jyX+
gPxV7SJepBCwXT7KWiD1ssTu3Lci9NeMQGL6s/vtc4jClOLKBZRJhs2atNDGpeEBDluXcriEG2cf
RYwEKm6z1MkSiGuIuOIp8NYxBKzOQUKqCoU0oe46QKG0YtpvK0DnYB3AlAq8oZGBhM1f5ExnPQm+
9tYyjfFPau2XG0PuVv5BgWJg1W5rSZKlNA9NeiBv+lFejLxjNEcrNsPeq14Jih3xH4RmDO5lnP7c
IyuAasvkBuvTPfVzvc5PFw9ROIle6+zBbGggk+4d3Gc3mxIQUtWxh0/t1svyFhcgRxEc7RfTiMTD
Nh69ILNQ9+xU28hniUPYXpjleeqeJatIrbhQZLJHAbLTPsH0PiTSxZ9jU7TC1gQJoppR+veuiznr
aXYkl3YpRWPVlMhlYRXSjPnO8M941GosIMfGxDwQdMt36YqqJTbzOP7H1jrUofHlOUGAcOvVWgQE
7AARRobnGECS4fyuglCp5sIjfwcwDYY0kDtTU6KYvBOFoAPdYMeD6U2sPbzKVm5biAyMoTb0rZBC
XSVXndmrXlhh0Lv65MIntlWrI8VsOsU18+/zy6jX2+J+OqeSSsc5Ba6Ng/JhVB9wsqe8FmRC7Skd
ZRh8cRqSJ5ERzbXE1DqlQWp/4aNIi883LHAQVQVdrQigE5yX+y9lv7y9Lsz3R78hCD/SdzPDFHbK
0J06c2K7FeGRRFj0DfSrB+aLacu8EAjvBXBZn4dKOfVfVb2J95MeQYpiL5krGBw/muZLYrV4gucU
BXNKeuVHoLoziKo1xQI9Qq/4JcFJMz3ztJfoPLiqOZ6AD8VuOFO9MYSZLF0goXlS1ZNZmuZrRPPZ
J5eRLsAuvt4oPbUvke0orRtsmopkG7ZbZY+tiJxgf/LQhqx/Rj2tq+kICC/ajSalO6NoE7JXrxmd
JI7pJQBz8Z5VGUL4huDnmXlFn3OXbtcsxikoUCUcpRvQ6PUX6cY0clhVrt3XEdtGBIjJly2fHwJU
TURZcN2iG/jU1VDKZtqR7sLgJyFLb2EAmEPijm5Yh4bLIMc/7/Bu8I/Kxht58SeKqoTMq/NVk7ou
hbsEmVr7KQIOQIQnVEcpJVLN1D378ErCNEW3n6HmmBuV0xtVUvEsILP8efrGq3mpw73WPHp8Ib9/
QfN64virEX5LynWZnKlS7TEYuKoK+am816XTN1ULszmfbo+W6pAN0XcbfVfwZO578bSfwsVK8nJ+
fYTifO9bxlywFYOGDVtSCX1Y/n2bEm32bSS4dNDnertasTMjGvihwyt3MsoEkqoqlxXmUid+750N
jYgTXeVCwmEGjMYXdrBYfVJfTcq5mY8xojKzoUr5l7XTX2ku/1HVUZi1nOok1UXce23zXpoGVfxc
YAexobuLHBqHglAc8lzorqF9L5DnW+r2sfhhrhw/HZ/Q5Y5cd5lhbOodv5QMk2RGKZ12Nx5JGGYt
vTKilMioGC+t/WXlj5b4yac7lfrC/oZXr1PnxrzC2bmeKzAwABQlFzkzoG4fQiPOnFOKoIJVC5Yb
sefRPQxfO4SfUyMYWZK4QMFAuOrHxOH5u42uulqatGb//uqJwvRpWZupTuCAX5Z+SbJzrA+k/fV6
INNrQD9xUfy61Sy3whs3dx0jUjbW4iQhAsHKeDR/OSSoDe5VcgGN6mx7ESnopXmUXAcKnJOOfOqC
Hlyy++8hmCa5h44WATrnSzxizuu2rQcEeqCMcHwGimLU+jUjswCBYgJqY1RHXSLSgAZxPcZRvQ/D
OqSj0fqrfCzqpIKHPzapqr6kscpE5QixapcU1cQxngSmJwF3c49uNgFw4iAO8y53/hvUuAX38tpl
o9tLYvstx91pjqDcGFA2SwjEMatSeHy9lP9VKUvK5/GlC+njzeERN2U3WIYc4aJ9EVbWSaJQoBfw
m4yFH5rjz89iF6g2gOc9dS3MglSzxelXfLESqcaNfiH9oq+PUvH0LwwhvIFuPBxgf+be4smg4ELP
OyfrR6DsH4Xp9R9yEVnW4O0L8jxP4bR+ygEnOJZ48WTcHum9BLzG/Thctl6k1ZW4wKHG432vrAT4
G0UXkulGIk8jMmjnb/9RY9QeQ3Lvgz45txUlscbYju6T9fK/b9r4c8vzINKAD7UOpzAFyyIynPh3
QMnyx7Kzu914+/36CQ5A64ZeGuusuhpSkYy0tN+Ist17BfzbvimdmcpPUbEfGtIgovaPCuh2Oi5W
rHLCpy7IF9xKYneslQ5wQcPBWCVL2smjyPZKXBhSIi1fMKmT54aFQeUxZZNMUdPlqoYvozxNLewz
J9D0oJps3vSUVgWdVhtaHyCe4Mezt73vBi/zJiSunrwnKJRbIxeZnRRhgB2qZt+y5gqj+eKG0PA9
HKb6T/CZ9I/A3a1sldcRXlDc4e9dsvN2yEpQYbNPoT6duVc7susrKY/1trmy/KV0WKAidJzUiQDS
nTh1X1Z8vt07ekYhXsLjwddv5wFC1+QjyTcqt02VQBOFB0nvPFoTVOtd0A8WCkjSTRotKyUiooeG
JudWgHlgDx+opLstDfqb0s7Fp4eHwFHrUuSks5eUn78vmwVEt4l6dOjuCAFlyDbwEOtqj8r10fOd
LwOY0wYpIDJ2wLi6fAYnDr+KHMyFd3riOjc21U0K5iRDIbyhf0ob9EQJD1Mjc8CqBkFLH1a//DPv
1zUVlPSgwGFF0zjfyAIm7xUlpWUHNqi8HI0l5yboFS8H5Qe61wwmskc1Vc7d7D5tNFGYHzsVuThD
f8D1rYEmxVlOHjc0rsIokjst8wSU4bFLKMec963qwQzAwfDJz92aMIBNW7ykNubPXw2sqt+hPujX
446QPaWlOH5szKIcrFghlD7u6uNi0HccDkeQWeXYpisaNv1bj5EcST/MUrlmAvU6VhAMavlFeZwr
Diu4dae/3zKL8FY60BNcxy2aLCzoZrFiOCKdmDD9qVpnhMirmTojiBJddhr4nmS2ahBQ4H4T5zH5
j+ZFRkCuM677GTek2KVpdJPx9+PZh/nV4g2XwzCsADMynnjmSo3geeLBvwz/WAeBkOvlsm0kSa5i
lA6txr7hnqEkSUq+JIdWblziIeh/O6/lNVbg3iN6dbB8FHriuXzQbDigVmBhrwZEneqLoD2gqxIi
EIFnTRRyf7pSBrmKuOINsoMS6LMgamj+dZm4SR6cYqgZ2TnjUfERU4Udwzo560o2h4GEGfGSH1w9
dp8HcuCmTA2KjFL+5H8cOWVmgLG/5/bnRJBdGDv6Lte0/7+uH9a2o5qsdSXKsRYcfqbOZmYzc504
8A6eSPR++x9Ih0QKmA5VB3DyFc8OyPDQ5tf3TGBNXLYSKZ2Z0VSHCZlZin316l3fU6ZLl2vV9l30
+bW9w2WNkcsX7tch9Cm48+Pho++fygJdeRbOg/3r3AchEhdefdk6cOtQPAZQ4sPEE4eTiknplmah
7TyViWN0Um9gK9PhbThn+fAh2e1oXmmY8RRePsiiBTWeEHJ0GOL30vx7PixPbRHONHaTwrZ9O1lz
8TgkMM7elyh0QvhSnbAr+StKMNuGrgyJFQSK2c7GAMztzw9aUZ7C7IT4YJiioSPQ+4YtyPUZCnb/
RxVaWsE7LkRfhk0aSCrRTDw92wwLJYo/h5HZh3C7Ob/6kNd4eF1Zr4hZrHb25Q8XFLGK+Jr2hfpo
tXHSnFrDRy0z6Z3xzUM12BsmRTteC3XGKF4wIrAFiK+OwcFosxouWZgRDFlWKdkrwr8plaR0hj5V
SQk79jcFSIrAQlvhWrn5OxNxPNw2IBEL6AyHgol4bnjpt4nlYgto+zVWR1hxbttwRYlC8mXyOdmv
6lmCDkHh95HliHgrUwipWhnaPUcbz91sQdcc7aM/c6JDoBCHQco8KXw5VR9xADlkO1xn6RFniEOU
A4M89q1RMlRzR9IR3DAtBiGZLeAzxI6bzfvP+l5nA7oL/KOfg2oaBt9DnKAIyeApkNDF7fST3PyI
3ryQnXvOvmsZrLkror8EkKbPl+bmm3eZXFMWwpKIDaHtjrrFb2cvjF+LHfPs/7XnN8b2E5IZe/c0
FoEYtpPDx/nE/vgDq0EuI9Zua8/6y6CYs/qvvuEEjGi4yupY6zeliP9RrPMLM0qvUjipnXF6M1p9
rI6LoC8duQvvpBc0eAZsXfpXgs4usanlr5Cp3p7EAqM6SsaACSoqiIWAvOxeX+/Qo2mrIEfYTW39
TcToYIyjcJA5jcWIQNUeB4y3E1VduCSlCU/One2Pm4coPVqBfuAN/1Fax0ZawfQZNHoPb0/LZiHh
4m1WvCowKywChE9+ezsN2HwS063KOXuNKc9A1Xw9pDUpeOt5E7N4TlL5lzADy6I9/TXmk/5u0RW4
L4+6ULlg433fkbF8hULcB9FEdCKqsMLn5SZ1HZaDzdQm8FlNWOviHRTCu/3veoxyqqp7fm4Ga+d4
E9rBhPvyYJF94c8EUKI0pU6rphPDCr+LzAFozBDxp75mGBdO26wjX/jdcQY/NZWE1P6WowVjiAzg
DjHyQNdZQulXJMTg3RW6BGCOzG3jhZ7ChkfsZZ0KMqOP5vFUrT2GRR8sFSkJppHWOAzv7k0WAB79
1vOnkE4nXkVo7p4sqBUB2Eiou6L1SvCUuRV7fhejuHn7oUrysNuIz9UWUPX1MBsUYwSOTSkpf/Dy
5F6iU7K5C0idE7wl+wmWGIWPwiMnVhLdTvo0svAYbj4AANekcD0f3VK0L+XIjZJl/jYckcqr7VBM
JXFA9C7aFXaKxiZC0F4FoeGBcc8gXAkItvC83tWKnwjh+D0Y7J3OqxxBEaWAQayCPs+9aZUYgQle
2q2rmtomiH9V8iPELIMIhRhKfXkDenuBaEXCw57X84WgvKUAVzD1761S97+6vzjwAsCDw43Yh+zd
1Bb1L9vWhYN+Y/vDoZ72ptcefOO80rdyFJjgIQ9WdNiTe//X5EsDVGRdD8EBSkpIW6dkdI5M1b+T
958PCsWBqBU0PtZj9FrereF5R0mptXOG3TGnLfro9rFKUeDE5CL/SDOG3/B9JFclgpVWzSSgWwlJ
C47/qlbJJoZXc+Ne/hGe/cUDLTog6Mi1YxjLMsMwUuASEyMDRBI3sX3y9wAXBznkJ53M7dSYWmJF
LkuiIpRzTh0h1J+WIuIvi4qOULk07uY5F/Faq5mYm7zFPjK6jTY6kh13GwkjDXdKz9FAVw91LJj4
5xJZNFyoJc6dhx4+glBTC+FCw23sk4OQ2ebV19oiTAInGU42POJuWLLIMdqhZayPL7ILx782dNwM
HIESobG98zbN/xBnGW2QljmVET78l0+VWkFT109oLoKIU2BRIBS4BRJHBsosu+YkUSo35pSCVOYB
/4I6YtXZrA1f/LhjtGRaUqMm1nj//DCqZppB9/wYs5FzHJUwsyPSqz7IiCNmKmb2mhWJC6a065dB
oT2+fg04x2g8CByKrQ7MfJ4I8Y9NkRWzEt1AxOfBpxFr2u84GAIEEbwQwMXq0NmC6NrtL9DUvOzZ
4qkqp2w+dZANiGQXtGHR/KBqvEHGYHlyxC26LdOudG9FQG4z1aLLwqlhJD9gsokVDlSDeuSLzo8R
Wy2LmcYe77WV46HB0E3wuEUixYPfwwsIfvu+zJCYjdqWk+ec7StHI40/V2Yenx1VYwN+JcVoCg0u
7EI3eHKmHC2HFckxcZmTWSPe3CMDtUUahk5AQ3o2o/SbqnykgyG/NJ1o6dwRlul3wE/WQ8jJsIfR
/Bp3gpL8WjmQ8siW4R1Lde+DpFsJDQG4BUp1HJaHPd72QAmhBuaXGl6oPzrzhV7CWr/Byju14kUn
muBlFZeIWgPrIAAJfwYZiEfEDO6wFpsjbFKGOSrPSnDTNin5nJhfFjO/LM+j3ZUgM4UnFxeIDLaR
AsQpGR6WOJOAn7BBbAQw/qw9ZT0pFE6K7OLJtr80bV2yYe54bt+cLtO4CXcorZwy8kZq7r1xg7MI
wEepwDfVChzCSEMrWgEpOYunccIvfjIsgpuT0ABbExsQ/OSxRMx6J4qOxVde+s7hsuLTrGFSJo/Z
2zPL54F4LDELlEbpHNC4HWma6Uk/I6G+SgXgvqR8eV3T0ueQXlENly9rM7B/pEnxE6gUY1qZxwJf
XCMpYWaXSor1OBgGCC0vR7fZBMgMo00d9k/pJwfrhAK+40ngYfi6AmwFDAn0ZYc9tiS+5YU0AEn9
BZjrDzktYDhbUhPa0Ol6cFcpcaj6uUpJ2cTmsUdkYh41yqd6dfknanF+qmUxQw7O9hXkdTyY+JsY
B8w98JPE7kJir9XrsSj+Wmn+/eF69jsTypDhwx+Wn+BbSzis2zhDPwht4vc9w1sY8HRYFRYZQfBN
vydQ2RdUficbsWCk2LkVeFg49bLDqd1+o9e/AVMhqql1db4cDF2sLL49ZdlJNmsDcquUfhhJDPY0
3eSZftUQj7CABf8c2O+SuS3cbnJtspMyA4Wb9qAN+1wVBiThvP891vflrr7PJw3pf1Qb5C7ekK0b
o7LhrNGLCFKhNM9cPzc/0dRFopZsV4uKa2nhClbS3ila+JzTHnKHkE1FqBOVXfyBtqN8N//2zwif
3rzhv5Ao9UajJMkveokpnpw3FkRYCzBY4sx0GnD4Jno6XN6v7/ONk/iNM9zsfWiHUkLRJKI1xvqM
t7/IwX4YvI33N60ROi/BxPsu38nTu/c2KR6tzjBD9xLgNwaJhdrMZieWhwt4qidRTmh8U2AMa/sr
b2qkC7Q4mCugVoGUWyDgPdxMgqtg9AdfPLflxfTRvBi9iV+iha0affLVhAD6nc6PuQN8rWRXezsV
vbY1vsQbgSiFWdAaiFDs36dKEJyrU07F3xWZHZ59DGpH5G7ygO5l4xVAqexhUB+lze1UeG9Se7Ar
Khq600BOah9DjZJSATENSAMjXPBUBFdmJ0LBxVOP5MLXS/sy2iv88TZMFY3ZaliSJT3/aUG79dmF
trvnot1blzVHx6YNN4B5DHZgrL3Z0YWjkLxq+iEwZAJ4dLvkOzca1ffR+vpLTNDUfJ4tleRbB3vk
lSugOIEqDvDZEr72q6tBfTkYkHCf1CvJ/VDRpMufD1ipmL5wCzE2izmmTYbG8kbBHUVqcDwY+Tty
9sosMm72x9FeFsaaUOAoQR76omhJSCtdkd+jaglp9bllva19SPW3b9+z/n8V3j9PfGIAo9tBFRWr
aUJriFJlX6pCcbnZhnKt8/9DmOTizqeYtr5oXHqsVrfwhhxA4oZi5/u46SaJhf9cy7WyVCA1ynID
S1PkZTAJ/k4952xYC5MiEhqCOUSuMaC/eg68Zm4vF7kj+dEPuTMRT2cJ8HSJow5dw3O+3zsDipwt
upPKAM6Ah3CNCiZgwpYEX62SuNaXMpwl9kL9bs4m5ZcEjEIPZpNLkX28/eqLEpbILyE4k/D6D0ek
umdziqcyvPHGnywQnlN+/dACRq/UuL8W+UUK84m8ZL9Uw2zxOaCHJjC18Grch0SmkYKSvP4VHFsi
omA3V9MvYD45pctCl4lol9dBLAlmAGd2Fh+fu0ewCEhbG43k8LQSeyNEa5gKYLi77GXYzr2m5c+O
Y6DmF/EhANRzzpJsfr4Pdagy5ekzR4AriceaXdPJfeyinFML+6wtxqtrfJ/uQOokrXGBY/rucQwK
Tt9//9hpKdJ9TGCsEP8bY+9yJuHqStrMG8wCVvbKoNAm/PkGnCwb5ESVAtPtoZTSu8c+tm5gsB+d
+S+Ag0hbVYzeiAIPBePjcawYWbcf1U4FkZ1qQTdmp9FkQn69QXmmygQh6ao4NDh+tObywhB2fAui
ihStPQLRZt268XNU4ptjtEIe+WAxeiLM/6yecgJKkXBZADUn0D4eOx/kBKkwXHhrfvXi10s5Z7LE
vc+4zsxIam+sVSgaBSNfUewQFG/sAd/dWE381GQhhc8bNn48ud0WAxkCRkJe9D3LJ7AeqpfS+wpN
BquORWmkWe84RByVyjlyMgmaHMuW7h0qP1PczxT8RgF2Ll8XfseORcmjUIgK0qN3ZFq981OGpTtT
xbz0cHFjcyW/mEMBDRjfuX0NdBZP+LFRBwuMY1s3Tj/3FSkhVsUfshzVGmkp4uBXEUPG5bsTO9Qs
9C9xosj7fDUTvjsz6z59KzRWzCUit46nHmTlDyj0VbWTzmhRcGbWvTXrVIFKhZCTqGH5PDhOOU6R
qV5wRt0JZONHGSDlwHLCrKLdUslhKowhqL94AXrEyCygdNzsFg0Gxy1e9OpxWCZVrohqSDPZv2Sj
fnoR/5gLEFysb2ETbq+yu8qFJXsXywjLVEmKu7WpF0BvQF6hBkbZk9gWXcBr3b4iMVIXvmBy1Kc4
nlqDq0KP40vzdlioRkP4p4Aldiso16JKBzUbRJiYhVFNcCS76UC7d7+oYC5xuvU7XPGRoQQS1Hlh
RNF0lvxvaLlSTprgYEtZvas1YrqDNZVtoa2G8LYopRy2K++JYBynkCb1tN6BkLxXqf0Jve4jp1a7
AhVApW+Zl6Az6fSPoTv2gvMOjiomf8PGmJRpi4MMLaYZBKPRtwJbzGNR1vRVV7bi71mRmj0GLe6g
wj8g5tlqDnXXcXrgna6gd6yw2QEtv5A/PFW3fFG3Zhy1MNP5LV3bdb5hK4Iq0+IX4ORHiwEcEBuD
irZp2ApQ9rkAd1kPsaXvmEXq06mgPbWVSjqLVnoX6ch3ToFyEKUTZ0sh9GfUMZ3ABliQf4Md4c2K
P0aUzAjDSUTD613Bz5P4b6RJbB9xKsqBRmmz5Q781ZcNZBx6fDMYdxShVzmPZUBr6vKf/bIuYXJv
CtvTljzV/Y2HriD3srSXqh92g5lx7zO6Iur5F1RIrLDqefamRydQYUoCV5SEbX88yw8KQoO+xyUz
GH2AhceE4bYMb3fDpPUcotPXG63iZXSbF51UECmKT2ZrJ/xDGEdOGtxv8ApOp0lMorrZdvsdmz4q
vhuWOHgf4/bwzs6OD8CavjZd5eSfbaU5H4CvP7bi7AJV67BdZMNiz939XBiRXO2S26JAL1Ewy46O
5c1uNlI1Vl44S6Fhdonp161Nj2Rsurd4w3+fCv8zgPbrB0hs/iqw4WSetYfCvcOSax5h/3zXZIrH
ayfIzdMke363lBnHSvkVx3LfKqNW8IsfcpeUQIK2MSUORtifwLPb2ag5qFe9cDERCyXy0Mquso6X
2VjAswrZTRf4ihOPlXlHslDujbvEOipTVMn3N7YqzmtztWoKE6UgVmc5Lt/FRVjqJo3qDFIlfeNi
7JUabHZMGfB+EG1LlGiTi3WHrQ39Xo/DV8gBoK5xByX+giKHrKi34wvinFModE8knxFH2Z9vpYgH
GW1kJBgh1QXlR/ALlKH7i45eekkjvPeDFtjZbqpFKS9eD03jlUbwIYK8XNWcNF2z7S72br1+t3rQ
tVXhADfxbkIDY4HUCtpp6Ra40YUzt/MWbAvYJP8Ih634rx2lGZXzS3KdYpV229dcZQQq96v7wt3s
3cqhRNWvHq0FvS6SyMtK23r37sNSudXee3RodcHhSij+tkEIzXDACQQzlr3QzQi7xqOC7XxJgroi
PpEWMF6RX/OAxq2ViJK/4LzY589ZRaPVyzBXj88N2fjizfHHqGidImhlhMrUH/MD4aQVGf6ixu7I
Zf+LPuGH4rokiAKdch4YrSyjUOnXkugq4hoBUwNm8cH+8Io26bloBQQRH69yPSnlfgZn02bpPn2/
0GUUcSt4gOqbbcj3+e8jJLZ5BnbRO/2eYwJ1/kPODUjWGF29hsim2AoTapAyiumLKtlRwL1/LpGP
Hwlh8rgnD1mrIUXSqvsWBbwE7f0b4tgCqwepptZpXujQi4WwqpkFD0EGtiCSxv/kKT04yTJnm233
fvxHsQ5pjqpkzVctt4pRcAeqnzQGGaVItfOR8o7IBXj/Njz6OmAw7TndfKiV8KvkdjArtd5mLBX4
Z3NjSniHGQIuDVgcO4pOnlzcHAjafHz7vv6XitWP789z7KFzEq1857zKUKLwKjFb8h2SUWnFoRrh
CpswknFiFOXXJfPbMpbj8ua/sbwpKf5oxd9wGNh9lBa18VRTIN4sTe9ZFJywY0tUftO1cfgc+OTZ
QA4SSiVoTRXBh0gXqsR4ggemk+m0DH2JOejJEUjpce+8W0+6Y0qVExezwsbImYvQao/gRT73p+NG
z7O1gyL2CwoMpuTP9NqF3iPHNox8Q3Ti01WPzM3cDykvbHjE2ls2VYKmhPPsYzy3/r6GdeBa/UwN
/FjA7p2s708QsHtB/EL/WuR0jFjl6hb9nyRnIY2EjpMpdmwS3SOC7Tk6GPJxj80V9EyYNJXydh9r
jYc5hBNPW80VUGsOixceYGsKCsGytrMrdrJTOAawf8XfNoRQ4/rjUqmoSVaR2h4pYWGy/p3cymJi
1YfKe8vPzZywlxyYtwnYM+jmC6QxjGsLe8xv+LNm646doKs9//l40hTJkW0LclYac/8Zvfgrgv6+
8yb0ngrYd4+2WTDc86wlsa5+Wj58Rvs5AayHwnErj4XNVoOUJs1WwRuyDyUR0G+ppM8ooP+4JrOi
i8uzeItMgjsrGMSOtNRc9pTn3XUSVPgQ9O451DuFjkqddGMg4FcIEPPMob01a4n+1eCf25grPY3V
djKikUudyAOX2pphf7gcEuh8lKqRMkwZJayWq3Z+F1EggiNC+AwiOYNY2h0uS5d4YQaI6Rm0Kq8a
7zAB0GHKMhainCBG0y9US3jTHTTXGOkfChAvojx+ZJJV7H1VeKV5fLsybyFs3u9cjAPJ5MAqCCz7
ICovanVIENfL6SSAv+MvrW/wD85k9XHIwNVQfEUm0wNPrFpneI86MFkyimirwXSkYL1m09rtyoSU
Zds/A1kQCpgR8+I2WRUkisHTtsRal2U8Gf0dp2cyz+4aAhQ9jwtfSxYkSOtfTv+umDpzE0xEhyiG
3ekTIe16vIMj1uKYqj78qruRFpppmzvxexOqZvirK/E+c3Cjge6pPbkufsNK79oT+WQZ6OgVSTmj
JvbyHw/s3ZeDIGW5Ntv5zMOhc8W9HwMNhSCBK9Ip4YNG2vXYHZtepZdutBidLS9giDTGPmgwKfDU
EZUgTnSF3FwW0mMkHQnX6J25lZiNQGbN8ec4lzZDE26DPc+JjcmXvW4xbYuhxRuVwt2LY+yM7b6F
lBPWhquRZGO7ZUo0DD2DVko6y1C8mi4APwbvm94y8+aHfsAxYYb7FN1Ej3b8x2BwerY8qtoPLElO
FBvnvgosiiF1mhdfK5B6rO8L5QFRra94JB1DvqEtImA00tDOlSWB9h3i3prjb2zs9UA5rFw+Z5Vt
DzhuZaGwPa31l934jmgAUPEnAdIO2Ap0Aq/TpHM4vCHbBXaMTeAFrmzCREslOOe/nPycIX2RsB8G
Te3GtRgFfLhd9t7e6A0WAbIqseGlCHzRAB8j35NqfnCFVvursYmzEr17RIAMRjR5/9bvZ0hdDqy/
JLX28S/XPrX8oGGes0hDu0gWU6Fsd5OE5N4dju6JjOuF+Mj8OF3eVKqoOV6qzKhbDzGwFLlBGoFx
6neEaua1/00vVO+YYtUNU5XqvONg3YiCf5ZxNHYAAoRLSsAtIXGKMisByAWKgkouOMbAL5v2y7Dn
qPylkwx7SEqv03CVsaKCj5x/9/Zp/17Ua59/Q6ay7il165KOI+tL1Wj/veqLo1Hy3Xc5eWB3UNeT
iEpiVvJ6a1GyXAOx1q3whH+H27qneNaXOxka1W3wMfaTAXDRbqiasFYYqZJZZ8yksNflUfKNRReM
Uxo4eTzKk2REBo00OhH/TEeYfikVHfI5F4A7SkqrSI9NptMfIz6pKrAN5KVYOfnsA5qbkxVbV9Nj
zBpisLPo6tghmvTCXzXK+B+V37O3ZzgxUe9ZjSAHUQjGkqmyBx/pfqDDnQqHxcJ/GFvB6LB94+Gj
1GDDkCRZ38QMF8OgAgqCZTMaC/lk1QI3ez3BVcMr/WA0MvAEO0cga2mJJY/cW1YXIGvrNt3lRdpm
WYDluvj5PfDArVcDK9Kd/Jtkq/BPSp8eTAAndeFHLCfpCI9uXojP1zyhcDtKILYTRmvXogz9NOnk
9691Mk2PAjf4ZFFvS3S8CbFMG7E7FlniaNyqDfoH/yI8Rxvsb9wqW966lKijcT+XcIEHf2JCzM2T
IuebSLaewToAqfDF+vjVKb623uizBOEQOB/CvKzQhtJpWsHSrPlq5ASbjPplJzM2RxLYE6dEqVl/
CqsiE+/JUHkzTv53OR28hT2UyYl6GsKkcigjd++RpVnCfNw88njSmBr2IRhE9qPnyL0gxOFTcaIV
BIq0KdCHeAPdXZO+Q+/NA8XaRxkivxWDEmd9KCBEjVBg62q/18TuFrxt/tfczgORt+gLIdbo5kKM
5R0wzVWMcvkSA6YmFPCdl+66BRlerL4RH2rKJrShmh0HZtD2rDZ6NwhN4n6KeovsmaWX67G/RnYG
A5vFbd36OjrABOQpJT1qmDAprjMqm6UAovIhU8iuy5Qz5LYzli3r2b2K9zA5C3MhMipVv98akAow
/l6OwoaG04QsmTdq+I/aDuzHe23cu2Jub3yMbObqU+OCFQGJCyQt/4J/GF3kvTnUhzECcOn4rTMz
calvOBXpmcvGr0IhDO+JsEcpq2vBNu7YaP3SJMcZ3EFhvlfBLUwtArP47jepeaYn+zAWif/n1x2H
/72lAG30CGqpDAbDa4Jp9ij6FCXcHaJWjSm6PtjLkDoYt+kXWPY77m6LGebAZdyLoXAjKQrrvgVS
yZK8ZeMAmqbazncMjinlWmy4UR9jfDFutAdH7s4JoCG8HMtdivSO9PSKishAO0c9FmL5aZDxp30v
Ux8jcp/HMFl0Qtrb+reqrEaTaC/THEJngE4mgEpjJcza26suJFBz54RRvxQ9QPRwmrcjMv14JEUu
Dy2AjclDEzhvdApyumeAMCCsr1CMWS8q4LrEkYHQ0EiysZAl5XNy7fJCVu357lcZ+17QYAzDtb+X
0jx9gZPtGD/xymXU1CVlo3PMt1PRvfRQCtGq6SHtVoWYCxiKIHP081F57f/J+SWr3O0/dY95fbV+
OQT+dqmANrg9UK7QrRN1ZbHkoDi8TmH2esm0JCKbEDpzPa8NWa9PRZ9RjJEoWW6S1xJY7t/uK2uT
HTTzL0qJZWnqci9Np4ZJPlXb2YXw2MXB8J/oZ23SbnmkKPFJpTIRfbCJoHdRN5gKrxAiYeFSMlRf
c27MrlpApQWJD9VcbLNDO0vRT7MunItn0uPK0Q6Q8Qtr1DZiuTfbgTTxqHUzmeJ2IHsysJYIrRVu
l86wpPIhhgb6wmLrIesxoxTlgwTlUIi4FY467ufru9zEF8sD0eqSyiB/nZaHKHfo+NW9ZaAcQDSA
X4fRGVPeleMENa+Q85B5tFdBm/d2O0exrIP5rd/zR+l22YTE4e0hI0N0zQpSAHlXJqvz1+4QTgDk
MzVhQdtc+1j6wMUSIIOYMgj9O278p28GWKAsNnf2NRpoBVRa1grDOi7lpwIIK+EpgGzRJ092OZLJ
cfOkxMk4Q425SUd9tbAKmdf8UhuF07kb3y32DRfEU/Y0LyZwS38b5nz9dO4kN11G+nnSQySTr5Zn
bcOCCWjXzvWo5yO3lUuOcf1Gb6FdSQqyFvKL/XV8FKfbLuLbl+N7I0+zRcewcP/U8PZuw6wKxwJP
4cX1luEP4k4ZmCf+VMr27ly7i5K7wct560Y6tIVsEq7ypa+IZsCpfcaWItM12H0B/9I4nxKWJwHh
GNKOIlm5GjR5ljK0eEuklOK0D9HlmwGUBhdzrv7OA+Db7xBX+zi146mVcEmKalNDkAof4MrkI7XT
maY7DrqUswjVJIqbQQJWKyNog4R/WYNtM9XC8SrpMFmU5Co1CW1SfdQaf+bR52MPS2pFEvkAeXx2
NZTIAHq3tvFRkTCvaHbSzyZUC9yyu6t+09TqNyqRD/iV2XFdIN/WrmOJQJvh76TZtL9Zti9w0Xau
rH7uTr2bhu6+kwVtxPDy5z4tkNhua73HHF9ELi1F2xyrj6wVL3bo/5Wy/1174dnUJUBD2tF0WiZ8
An0JOz7NXA5Tk09jhWDeM8al8lo4HGGKFOJUZQvZTH0ENQSDiVvN7xeqPMa7VY97/aViQkJsKhIr
6quzibUYrhP4VC3798tJrBrPu6Lc0isJRyp/fInP/KE5WsEhlcw2B0dmcMRBs7Hf//PdheJCDbmf
ynB+Fx3ofLq3whFqoB+Lp7pU5NnizxUt7AmgSK4XecmRB0iUfeHWDuggkRc/nZQwjccaaK8qmbYw
rgyAWg3HGzAuiV6NyZNFM9z6Az/bi+qNeqfDZg+V00YcP9xEC7YnCBkLLEaqn7P0wEFJszRz59Pz
xCuyKOeluCsZTG3RSnWeIJcx7PoAPD7XWVyA0enEQUcPRyjmmMVi95Z0soG5kgdv8N8uEtfA3Qt2
Qz/qsAVmc7SODgEB61dpkLF2zd2K6o9e4GZtH2Hsj4PSLoY1kKK3MYcjk7o90x4dYCPSXXJ/9Wgt
PF0Jt3NT3+/XaECcOsPsEPGriPEkaKGJWidc9doofLSeWPtubYV5vSN3EChpKrSZ8Euf+UPGE2MT
gQ8Cebh4p3n6+P2JFIjboq5zKOwr2CnMfkysRqazaCUFLbr54/gPXNQewrYKD1ZrxiFD5+lIXlAO
wr/Hj/4ZqgjTpcvQYHqDGCC/GmngcVi3tzmUPVRjkBjqPszpZ6FtF0PKWEBqbzDRG8YCeX2aQb24
rEpePI7tj5Vdw60QX5IgbUL2H+IWQpzVIgJJvWupZ9U+Lj7c3BpX44jzQKjaiZWjul8/eODoyrKh
Vxea69MbYiAS20ks4SZ1vRNnvCZ5rc1/y/FC55/n9fziTSrOh1EMi3YcDFgSZA4yEp1mwt6rRBv5
Od82C4J7tyBlMrpw1dVdgcFb/dyAUCVX1JoSglvQ52hMPQ90UF6AuilN5cqhKVI5yGRJRRFAHZhD
sMyYl15lgU9AWzMt33vgjCKRJ1pM1im4s+KeMXsglWpe8nDooENxIkynr3eYnra/G4Nuh+wu431l
CK/XLERPRqndr5KOiknX072EWRGMSf8EyAiwP/U11cSvNLptt9EmN6nrerQXlV66ij19McKBCFOq
FWtWgPyE6AWIcWd1vYOO4LF3bo1TpcNjvjq9KZXJkRSqWF/lpRZuYxKYHICMIN1PUKgyvcIEw3yC
+Fk862r8i/ZXChVsOcUTpUHAx5icX89dFi0z0iBGj8oke4r4K1/ATahdMffDILYoT5CXcKQpM6Bx
VwIbeePOyg/l9ruChnQohcZEtx0s8XpHKD6bcRtz8+0wL0E85RteB7K+lWhfw/3zzoE4XX51IkLh
ONFcs/RqvV4Vr23rfGr2acOD4Im8v9tYeTC+l/2rSLeWN6yNZdul0McbZi51t0OQ3fh2aReH/nKW
bElbeGqR2oOanF5IYOcQDdZaSQugXCy+YXLcX6RBNNwZY5ozcIFQBV+RtW3/fdXv61HcXi0O4jA4
wg2rMaHNR1gnx2QPLAYE3HMOutDdU2/zPug20eYQyuBLC/ysjRfuLPOz0bkAfhlVZLgRbFEUNXCK
Yyx3A/+BQjlh4EOLJm4n9G/Y7qSYO3pyeyetemRmETpl4j2ybwfGu0QQSUCuY3qZHASvWe56Xqg3
pgNztW7KXQbR47I/QvdSogxpJr70Pj+AIJ+RGNdagRVTsmz21RCMvBzNstZJEImtmmqOcZlltqCD
/WeLdxUJs5TDjWqxSOR3w9P+0ESLO6QXWlCTpx+pPzu++8JhGaTSLv96npEye7wmE+30uLNQPoiu
+PQ6aaa44YKqkri4PtOapYxpyAqdAz2W1xkU20cY9QQEkJrMleeU4MPH3iuF4tp5wQByjA7eABq1
kwNLYGf2hUJe0QQvaXgN/Rew8zn8/Pvph8mP5/wxXVX/XG7hjF0jmmHVD3Xg0lvk59W7BRQZFGzl
7gnSJUVrGclTjx+WoRsU1+34dU55FIFX92vK2wVOok1N2lcjqMCOh47VWGNJmshwLbJLKif9rw9p
9R3dUI+ptO81g7s+fHwIidqBYppR77Efo62hx/hUkohmGXIfUIOtXB0xwuxsZxCdesAxsPM8d/Jt
v+7nbkOH7RVsGBOC0JXTLRe2ZMdKFMN9OjTe5srQPPca03kggb8HymVH8t6FiT81wD0+W4d6zOPr
PUXVb12BkFt3POyS+D6+o8uUfYFsR7DIAR36BcJgI661HV+/j1pK5zUFkO0TwSimVOylbQgNOfBO
5GeVQyqXgoxT1PqhwO87LK+2aTK7F/gUv9hLD3fQgkSwrYvUNgLptJK8jD9+Ate20MQPSSPz0lje
LiU9v5aqs9/2h7JoBjT9Jqkd1oJqiWyM0u0dq8JublN0ZfGe2qRsICDwgzSOlnJuFtnNnrrooLIG
Ubz2BeqSdSSbooa3zAEFT2vEvCNt/3Qh+85xh0aPu4XBbsUdC+YB94vt9fGOhf0FPcdSCggKK/PT
7th4TeFLYn5TllxaTXYDRG+7bpCM79bjhVNk3TYtEyC03EmaTjU2moJJtj6JbjgyCz5pHQfJMDc8
lLAxEwN/RJMMchcmN3BefWweGp6s6hX+gEswwMptlF9s8VcXft19giR91z25to6a5UZBFtVBR1+O
xRuoozJAmNmumTI6qJrUu6LVGXxIBX3UsRihs6ixT1szumHCxo0ZK9VyaXwgMiEESXJcxCo5WoN8
75zy4TbobG7Wm5N9eXr+t4sxQy9kqKYryreg4XshyqQasuN3qfw8q9WsnWJ5os1Sqv7TUjCf8L6k
s9xJFZqVM49TtQfP6I+WuNYrFAA28srPs9xhixdkMTxMVR8nVdHuZXdsMLW5Ojqs6ESyROL5xFG7
nvW4PaM4EXo85YFtVEolBfKbReYq6Do24cCwDqWIcqYE5ge1hHU0kVdXObKSr9wLJsrVsfLNiinx
7vkiQgwvKMbZEcvfvhk1dnHyGmz21QJIFyovVeqRD4d6S0iUCoaUy9g4aU3deJLO6RSix8lW2tEp
heP2XwzWl3NJXU+SItQktRNIxfqgrsr/0YHOaQJH/oKKhrzAgk2nkCRL+4i2oKnygySpkOIuqPv3
n4jdNOXoSRvJgPy7PG5XQrurpX3KbkD95k2JxsMotbBgK5IsyKIULxgAlskShuN8OxAceq2fdoZ2
AaOitfzU+aicZ6tXD+NQJmpB0DMePHUZ1++IpUXXDheVgvHBgR9ojoqFGurpvupnq8Dz5hMbuknG
ptmaPoMlMMXzjWMuExJjUuB0thgbIOv+eDo8LopGxdU+SWLXSi++9s3aP1IwW/E0zTSiaOMlfjQ2
CBuuWb8C6I+KCM3kv1UIOSAH2RRbYVbWpJoblzNC/a4c2pl9d8qmekSGYw14J0fJsydPvdsRlMB8
ljNrQmStoxjNm1roG4mlUTWyDyuZYA6wQPINW+DHwrVSO3hooWizHfxMW90NsF89NnxmYy27k+oc
1G0F2d7ZzbDmRepV1TavCHk0ZCdYM82enveGji+K+PWhOiKQEbmooK+1aJQfYWG+EKPUUqBB0jfA
1LR/eT38InmGoqqQ9kdqygKiqiLROiov2RUCZws/skVjjvCqqnsC0psdsO9DSKB6oRfvU+2rlR+D
mC9kaPlXuBB1wpKfGMnW9LfHAOnF5UZcMrorD937uJERQQbtGiWt8zJGRZtr1XxGKi6y9Udaj7JH
9qHd1yJWYjzUXSCqMerq3vkSSVOj42EdLI+ZnszpVipVddQxZslRQK6Y3Aijfba3mzHv9NrfZn5D
Gx3zCp0mmNS2Sv0QUZpr7jLYolu85jUXql5c4WG7YAgiQbArgsbPEuuhoo5VTjtEPQKEIWPg4AYS
4oOkT7rQTJ0LcZmKi7vFBf8dAN6PxnKcYUbFRlyZCR+LjKjIntyjyGm6grndufdjnf8XAQb00n2M
bvASgM9sfgNwVm2VLXP7SkRgyWZ020PZzDaeEylZT13MxOFSxvGulsEaTkvZEMTWBNDb5UNDjHc/
sLCk1k5NrqN2cvroUFTaIprYwdDVTiLvQJOPGWH9pwGq/rMMN0/0Nk+cjjgiE8GaQtkGPIYvYMuN
byIwlOwaEOXqD1vgLR8/x6Ulk2e9OS73XXTOZCgZAWYC3gtVJnBdqNMip+qILMYNcu98UDKKcXZJ
CUy5SQVJ+MgSPiyPr0YgPGxCKx5+26qOck7g89U1MzC3LDN2ww+9ugclZN+nTBnG8ryNnPGHAb2R
tm/VXB+h8sgcWOVxC35S7JdcqA4GckAIJ/RhuqsmiGXaEzujg7gFQQPmWEr2JPDMiiK5oitNzIqG
Kkt2PYz9ZA4LV/7F8vYyNaHHdAYH1ecyv6PI6lfLauV97L2iQZ8DuwnoEvzS9uopIeCClNddN278
8RbUg9eLTCEjyUIqd2oKcjFhhHy0agt6LmBXpJYIGWivIvmmKQKkg4CpxrJLOfDfcZtiWwq+chsR
I6O1pUg7PWEuE/YYbJtqO/LBriGfuAnmZtFQjrl2E0hJIVJAbMzBJw/UN/4eRGFRv5OBGI5WpDbA
cZOm84u7cz3VVDmD7koSnoUt2vtXN9VruLSw22mStUz7Lu85soxo6wV93rFdR8UE1wD2AvSAF3Vx
kNTkKbDhiLMM5YnQjlR8ENVIe51ZcES/XS5Res96g/sAgkS6zjd5GqaFPwL/Xcw67pHnm/KhrMki
JkdjCtdPmknw5i6Wb16maWvSAW8LhmBzeJY7y5wU8R1idhZg46heoTfpZcrQij2SgA+IBB5COd16
COwu1cV60GC5+M5Q41JjaXh4/O0G/OsimWmln6oCJO4TGpxB89YvBCdjf0admyJR0YB/nYWX+iL2
LEjIClsAvtqL+ar0oHCXkCy1jj4IpukE7vz/1V/66QnUJIsdivUdYsoRiwPG4gWcnm/UQEvhfhGS
rnI9a3ow8emWHKKYduUdfh7eEK1hiBa/lzYvPSSFGkj3ftGhRyU08qNrkOB3PrPT4sR1OvKAWnwM
HFJEBSXaemrmGeOFDoZtVee6X6lwPHi3dQ7geNuS7xiha0MpuhMpb+eyzSo/tlJEUhKjcUe30+3S
G+EO6nsmeVEeF1Wmh4bSd5C3AqV8CQlAoMpJb9M3LAC1HMFDjXmfZbV7uTJj+DXes2962TuftdqS
fh8vlGC6BrT8gqL3nZKL0k4r5tVn6U/iBUilHUTPXGYpJKzrl7AYjKGSe8HL/QvVkTLfNzXpRuJQ
QBCEK9MaNxAkX64fKYKVVtxDofT7PjjTMmtNR1e92Mvck1fHWe6+8qJ43OtYXFltMF7xF3NKCQP0
5oJRBI8l3ivm0sUVO78YmJ2/2kZLFaWr+UfJBjrQaY09HtWM8zyycpML64iThhBCif5cbdOs9WAr
yWU57QQ50BOptXVe4XAN8ek2Cqv38aH2WKwRhRGQ1WGljlYbZNGIIu5AstXWw4+U8BZC5S11TRTf
yOWBp8s28StOBCdJ2RE61kY16AUh8fK6FyPX299cU2EXgxqVI5jtbUqmgOB9fXQTOBsbJHNIB7QB
K5PnQA0XAGNeEpU0MjQIiXSXt7XXM73FQIJVJCcrcqkONO15nJuv5rNVlvRIIwYspVVc6TLYp6Kr
VkFyvzLd51pw+VKIMxPL1bKBM1TcMc15D4c1O7EfM5aGH58bsBnBPQkGJEeasSfwWmONUG/CZxs4
gcTP5P4HQeaBg3W/068gEZSQDu7ObQCqjDzYecUYyaRBqnVw+1xsWYTtKQakF3BoXD1imjhsYCHs
6/Yg7iax3l+2OX7QKhuEhdQIBJlZ5H3HHtosiZodUc2BJaCB4wM05AQsHmF4flSBSoks/XBI421B
T0QIByJfF4SKP20MPbBFnJgMWZrzfjTZryc/0zl2QqUJYMwNlPQVZetm0AwRpZuyN5rucR94v+FY
N16gtUSqavO3+gkFBWFjKnUjM6dGLChFVh6WVtNDJ7+sgt4pT+wSBh/wVB3GWH9fvwp0hgCU56eE
VIdpZ5wJ/Secn4EyIe2dId6RRRxRHms7+Evm+jQaxvvRX41+l/WkfABGgYqByNYwTT403C1ySoOS
jscoPWQ5fBQJ+zv/3xQ1nFIapHoPjeNkj2Zc2Ds2w2+yntbBEFTXFDcL8/zUBHtVTfZcQyN/Bnu5
Y2yzOkVkvZgkEgezbJR8DhWMIRG4IrFv4LORXPhQHItaNRAxWv0gfCUwbaNMzySS/ODSYGDx+gDi
tBgdE4/ENNCInVWC5h5AAv6OyFOS9wN6DdRH9Njx5ZcU4sY0KTq5VGCal+9iaRAAdxBdH7w8UXtO
s1T8NEcxbJI+x1DWH1WvpWvVOX2izJccDmJqE8kwjJSEkWBj5mEFbReW2lXM9/PkPcdqqO4Um94m
yczOSIHHsjfHSZg0toH2nqJlYHIqHqRwOwwLQuP2s/3jhE0O/YTFFFy2GH1kVEFaQKysdxck0d6y
zA2kqJWzmiW56ecF0MkSXFiT+zgsPZ7Oy1PNot80TLyomZuRhDGZ5GRd+FoeM6AqtqUAlNE48UtV
pEhkvk8X4XCT6q1/tLgJsUF76sGY7aWLPTJsMVzBpo51TFFaWylh5RR25gOHoDfsEDeurRkW/2YT
9/f6I665/TSdig9hBv0SS3y37v1WZD991yOV1WNfwlUcQBNU3fPdhcLU2OgW8IsFW0ZD1fOhF9Wg
BrVl+bQ4hSjLcgKEQaTfwHWZkg/yeYPYokhrhfSgbWmlehHv5WJ1l/bIbNCIGQaRNH/kOJZQ95jX
taGpBSM+WsejDR9HZWn1pFBC8epKRGhkCuLt5yhqcbn977NaLYN4oWxTc+/fbESvU7Dg2DqWJsYn
4Kj/d5JmkDKvqVez7seIejdUCR3zrqg/zFGPPp0i7UMYIAIBijNJySaabJv+ex/XpbnXNFRVJvv8
vQwZW1OH6f5+ALrpgxUlP3DajO/FlV/JOdEjG2Ec7SvUYlCPqHnxduKGd9XAa0+vWAtKy0FX9ye0
kREPtuZSYqHxT/ps1VVZhflWhF+AF5zIxjdTmo8otqh2WvyYvgLLUmssSfDrsaGvpH/poS0SNY7/
Erds2LPuPceyK28xUSmgEdxGfT8OLMsHu6z0nhIOw1TBhQavut5g3pe8zeeHoh56gwcG5xLszNTP
Yb6Nzt5F2LtBYU2feyFAAQITPYx1TlgWfPGIbkfdSotbzmO87JYGHXAq11TdbJDmaduCSnwKpN8I
aBMalySDjWy2M7kp84UnAelkTiKschTP7sELE0Hdxt+hJc5Rh5egDXFTUBPEzWbqrh3+cnmRB8WV
lLiNZAp5PuCFf+d/IkoxRh7iq+UfBE5KIEHcMbjY10OLINuUjotZuKKWUA0Bp+WX96HedPLj/4yR
h4MSnKk0myDacqDGV8h+wa4wErI/a35qo8bjjuXCi9boK/4utBWhEJM8mKXLU4A3IwwELtET5Fta
l7sPT+jv35g6StH3W3R1y1ipzmCLzvbpLHDVk2hLbbNG43Q8wQgVZIyei9Zkkl6bSS2QuAv02xd5
lSTbLwR1kD0PYirq+4Enqc63ljvvkRfMkAFK+gyXfYt+9Aj6R6k0zXfAZu9SAq9ltpetd5nrUCXb
ZRI7fO+QohTNWBROubYvVZ/PNqqj+fqbeo9meFAAc9h9SyB7WWZ8SE0b09WOWuxPt0uQKLUxm75O
vUfDt22X6vHuxEUnuZ2IyHsX9RA4X6HV3aIpw1zyeEcuCP0bAr7T49YFtYlc6ac0iWvce/jFblPE
CqUToCp7DSdhxpMqv1GsOcO0KHBTJNNa4z3jRlv6CsYIVqmkT4XLyR9TE47TGos8n/ASteOMjH7B
IamwK6WQgjnnNYrY2I5EmTus1x/6Wmf0tEUmwH/LGPdORnQtVe84+pm7Y79vZVDFNi3IVMfkM7/j
pxVcT3CocXu5ppdhbVelss/JXILhO1M4dtanubCjuXNMBI6vbyZu04nIz8EQ/dSBvlanTQnZIQLz
8aHLIPn6itErthiyQS2au9ScPdvaUnan2Kjy2mifC/l6l0x8xWZIXYZ2M+duX5Js9J54YnowWygE
cNg4useXB9JI/qQq85+Rh0pJi1EUEGE/F3X0C6uDhjHAgnnpdZQIpDLd+bUvHXGHUWDB3kl5Vliq
JWjdP+L7IGanaW6/mxM3kSvQSY8FdbTvcEohGMJqyd7hrl3Vm97o66A4rNe7F4V8isPJzHllDFn6
jEbFF2KxfGE+NNZ4HlUE451uJVdlSdoEpfm37DbyjR5iAw0hd4rv9axAMx2lde1gPjsMZ1ay8CNY
VCbmphBJFBOPnzlEkY0tp8e0coKshWLYVSQEDDowLPkE93k+poXXRhjtb0zrZaNZ7W10eQy81zbq
bMre7+vd/FM0qs+C8CDjJed1BnCHxx5BeL+Pw8sDBQWrY9tCyeNeLbJmWuTZJ7S/RdUJYkfvPDVy
PLtsili9wTqBfli2K8A2Ep1rCMJubFn86RuvYzZVsVoQc2k9GTJmvoPfGTZZU9E3Kk+QjXb0ro4t
2G9d69fvcNjtzI9RbnHfz/1hH1I5eNpbIOmZSN3cLNlAMujDb0KY+k2W0SmxxBJUbSQG/FtVqO/K
sitxethaEDWHKK6KwtFJ97wwPwN4dK/s5DOX/uyjlTgJZrW+f6d2rOOPVYWkAadF85z0c3Z8/nva
8E6BFPCWcUI/I806+Q/4/0uEegv6fv3N4pKjzIpLJeRz/lX4qaWYmMeSV5d4X+Up6VhiKTxDKuA/
awHyJqAEL2jMhWiYbRMMuINUhV013yb+NcLEWhMLxRYvXryaVNTtuOqdkSvFAMBFXQ/C9Yz9tSnR
0et03U72exAA1/feyZIH3B8nbVurNbkKrJx9Bi/3p9LsF14nx45TBq5Y77fttfS0TS3NuEWi4jlF
AWSb7YFwFd0ygNdTLP5JZm4bBxaweIe0TjQ8SO1mzvuyE/7jbBrEbi5vxNbc/U/GA1597QlXkUKC
4R0IGow3s/+821RBUR/iFoKVxu57iEyB8h5rrZHACDsu1sbuFVO5ifRv1X6iEaclW3huPc8Qkv2W
AahL9ZzS++KlM7oWSgKaYLiZp4KZcP7JS0G4gpkch0YOX9hQH2ihP9TExo47pISMV22baSrAycFy
64M4vDG21FT/BCz53K1eI/Ck8R9pGd6201bpuJUQZ1jGc3RY7fn1sSWCPqvKDj0sTdUkr8uOA3Jr
b6nw9eHWF6emigdJtJWnx7VcH1Z+uWTgy6S1vCXNquEHRCRx4rYH0NX8wTrOKd2VtRyYfdcs/VL7
2wAejTasdGHL0qdpHBaYw/d86bafDfpxwUxCcIlHmpWB54Jvkc7pJBIzAqWVn7slmWVx0uEpZWs+
XFGdGr7Xny/vR5mWCX7v00vaLK0DoYXJRHUaumdKMfK3WYvFmQR/vK9wR37sUKmELGkgo1HJ8+1U
s4LjEWk1H50+GX1bfPKa4e9ud4biR30D8H2I20Ghwy1cYCB91iCYvuC0RSxzo3XJkVJ9yi7tzuDw
/lXUMv7d3reQTWSS3iqg8v2HHKTNnvbgglphQ/GpqLdlxFYH9u/4Y1ndF+j6Lv2wy+5iF1HQPER9
3lDcFpKIKqZqqeBZJLfxA1rRGCDYvi7Wbt5q4+GMxN6IwQoGdOgXqCnDupE5HDKGE2mMxTxW/yw3
EyKBgmHxiMcnWO4TxLMgyNxXfGFBapgDy5kfJqKjYXU5b/lHDtzo63bUcUhpxHLij3FVwHynDYel
Y0ryYah2K1sUYlPs37Xz6lP3MrFxtjMCU9rkUbmUJChYmhqfi3SLw3aD8OHg2vwMEIP6onZ5skUF
gbNtKpvo2p3KX2kPDxE0MSXW0biZOXJJxa9VbwoZOIZMOJrVSszZkrtjLUmM1Rlq5pXOBP29wiCS
hHZZtHm3E6FruNQ0UEw05ny3Jal2OXi3KVm2cfC7Bh/K/FcMXj2AuofsnD3I1ZE9Sx9Bvrj0XYV7
+jkmBAEayFh7owqZnxz5s07ioiVtddb9E7U6sx40GBuY5wLouoNsz0bQbxAgikuw1nDOgLfPujUz
E0JjT6DcZ85mh4R/fLM4RWs4135m4odD8tmxZ1zj3+jXgzsgqXJqNOJb7IfEx2cNUh7SfZ/HWy1Q
WWgjo9kjNj1i75c8iwaxAQocXMghLg7S7jheRluns7uigkIm6OZ12Fe2XRjSOvLE/USt4My8lIcl
K+53EU3jwrtBh96Aur3CvHdpdMN/5JPNaIMkeawONSZ4RtClPqPSUYkRYOvKx1DI3zMCSv+XyLss
GL4rTBD9h9qvdmRkpSQy8pCM81Lgs1hgSppmlmOAYdgWwePfnLxLwGkJ5r5LqVBjgvCxFMiCP4IB
TzSisKt/VvcaMjEW3vmfPKGvvcxKYYkS4Pek7JchA3EYD0bHiIBC8dhM8RgrReTJNsE8z+FUypEu
iFZj/tGjgc91vfmJZzZ6icJHPLB+QYP+d5iHlJbQ3Q85wD8aznBePVyiPAuhBbhjOizKUzvSltoJ
EdM8uYsNZ+0rxT1gdIeLBxf9G2W4GEN8lRGa0D0O6e+ixWkK4Q8IPEmSYBEs29fzWEC61fvWad4A
rEbso/OraP7e/7U00hPoHT6XnWohzBz6WYw8rB/Javfhs+n1oroHMGSw/WCAXspecUu/clQNwAwR
+2o8L8oBdu/tQukJOOGniqrtCMaZD6S8CIyq6koK/Af2wDPgg/8d4dK1iMnuno0VP0LEowBLpwPl
ED1Pdy2d7hhehs7O90jqZ4tQlwnyGsIGyo+APAEJaE5GO6RLVaZ14/H200lWifRbbAxe7WhLMocH
vMMJkFcktCbQEZ4vsf/Mp8OBW8YUvE7vyOuKBTHXWUfVIdS1sqJmeab1lv7oJptSHROTMZ6lruF2
CuitR5UVLqwfKUyA12Ysju+7q+PDncsnDnK3JU6oC14MeHAlSOoZRIuVrCMQ6pCGjqzKuiDBTzLF
P9BAw0kxbf9Ou0vxMG0+aDPwBIa1Klfo5wrgtl6dZ9jghw4FJlF/7qlZew7d0voGJ3CNsQEOi2Lw
Qb3OtqgDrCWobz3zp6JPgo0Tt40c21S2w9Nf27LhWcPQt7KfUDVhl1/mh99MEk5B6ywBoFnnXS50
l7N9j548PNGhbPYQo7yZatFZ9aRIwx7VQCrXrDPF5vTID5Z1W5DF6pwmqiS8+nM6k2HAb55CFG63
x05VUs0m452DIDXJrV1m0nZhKs3GYPJ8098DiJpUS4MglBvgaNWYIhpiHRJN/PEKzy/IrNiSW2kh
ZbGtZ7z0srtHRupxvqSAb6BVlhZylPESzBmU5bxv7cJ1tTrHCzyDPu219azUDUiHhf/jB2zP1Crw
EbfuDN4YoWnvUKt+JGpyJo9whkhV8qP1mFLArWZCD6ioNfgMdzVwpoPNuOL0aGARjZwQv5cYQ9CH
AXKPWZkkGUOcQxU/IYNmPfMD8877L66rDu9irK1i1DIrzl5x2CcR3ZQzbX4xZeUI905KkYgac4Ip
eypB+WTlUDGujBz1iPPHxe9XmYpasT8HCHqi+voJIECeVlKW4GlZDw0BFSfgq5WwEHt3Rnz1G7pS
YNdAd/sHxtDIbuyYCPq+sPC+Sf6/ttcT41N6L4Lwpb+wvVmMhyvaCCNDl66nGdLJO6nLZzNxu8J7
10AW+uxTIDjEaOyqO/AtbTfvoOEnjfFuuikAHQN9HR5mTwdV9cSr3wBUfZCOGg9Zni8mqe83JMbJ
eMtzUnb0/00AmW19Z+nEHSBTdeLDgnfbFrcIriOYCiGyaM/7M5WwgFffVEXfwmsoOLv7uhz0HmdO
L3kvArwJ3C2e8F68vYNplpJuznonzmRWhi3WldOSZio/0YAgVZRwBxY1z4HrTDER9k86svf3wMQd
6nOZJnBNIh4Yv0mjQfzzCnUFopIaYcwGyzTNk1zpvEsQqhWLSYMqEplE7rHx9lWXta/2jjPcPgBj
eXP5tDzx0k+7AQNvHEb4doPYCfIJGoGc0cdP2XnBg7NxaFsAPlrKwJI2gnMclgByQHTJ4ztPR2Ii
2TUqS4qFlhNdmYhhPc+PvLDtxBPf8dynjNJ7ACu9ygevkCQZ3Ml20Q726q2NdOYW9TKTNCReTZZK
Orkntc8fQARgIygOHAtO85P3N14uRebv7gpycIm0XnEzJiIKwOcCMAW4ZlhP/NgAFglFrouLnSU7
xPEEyTaRtSvvsV/0oNpxtIAlvzmK5DJ7m45Ui0pasCJcNeYUOPiXlKTqLNKDNOV+wcEnQzGA/D1T
ki37w4L0r/HOdAbp7k8BSATrS1qMFIXCkfOeKLujCX+m7VZ5TWT7EQWBUYeQKpqjHLqvX/rjXtEe
7sSmZW+MoufeVDuPzPUN/s1KF0dA0v8JQIFzDRfGNnkMlS5AsPmkkjvyaNDBikC+kSf0iPzuveKn
pGUWfnZL2aXISnKKrkjRw9kyEoqaEkZ9hlPkxnI5qz0RkaMU2poxDswlPo5zZUafVNJ7iQFlfMAW
xQ61pgbrZxM02XAkslx6l8bh9v7rn9fRfg173XTPX0iprc0Q499os2TPPeUlZri7Y47c10+VtVvr
uRiGD6ailBuJzqyLMUEC9FGwKyGkNAyZjw4DuO075Q4ekv/CPaoq3aHeNDA2KeIRnINHgAw5VDoB
7jqJKCusxr83G9W5kXn1yW3ttgCbvxHhx5ypKUROfLCoSNHTb4IbC5Duaa+uOhYiU61ls2Cdo+7v
O8w7JgxY61cNqFNdio4ENySD0TwRsie9eLVrruwIUHor16tZNVX8TOoYZ76tZ57zOmZambDstNT/
Vw3UcCMtf9PNwl/Cxni2Y3SHRsRobTs6sU1weZuFmZ3d8F9VyuVzcmxMpSc8akqaQdpNgU2Q6M/x
2W3ke+2Gb/qfjGH1IHHqjnlaErGD8XTlQkxqAyiiCkATbvT6Wm0cmIqqBTdodzLlE0NFeYd4WEHR
vp2Sio5ck/5vJGLhPDcNhwH/3MUhQuT84xabSIuEzbLq1pZEw7OXTCziQK53dtT+Z0NzrzmGUecd
UdpN2UiMLaHb3VNtZj6nA2s7nforB6zdY2Rv6h7gjT3DjogQJzoGB4B8Z/wOMSJchFwTUxNmAVFl
hauK28B88Fym9Qm0ByHLDinyPtxHCC+yN/IexIR0f6Ky4cLVk0RS+82CMhv53IgoQdwEg/MdnROs
HS7txTlmboTryZCYYUnjTGBnlYk4FC2/EN2KE8RZyuozrYBI38uMf+5+K1kogWmlBt1oJqltiRZ2
sYRo1aX7HNXX0Uh2WncZSlmyop4zpjP9K/xajdadiC6op1JlDC6NaHUDGX2WYXOHS+9wO2NTTjrL
If0YOpUTzSCJdvcebCs+5biOGaSB5TdjXmWYATvcZbPZ9S/yeC6rN7VwPmNZQqw88M4eJ0CUzUj4
ryU6EFfuFUStG2+oTvMfv9pP/M1SiLFI/HbMpsBxBS0xHKav9DUHUcEDn74bJ4Xu+r7DGFKXVNNa
xlyT8KIdLPmlieQTm9Q38aISp65upvXGe+KaON7DuO3Uel9N1weSbAbGbTnnxxmwDAAYmnNtxFmN
IF9ptt4wCWMXLOt+eFXINt1FpYuxomIke9AIMeExhAj1GIejBaKhfu0t8MnKTlOA7fhwx64uG1Kl
7bQcPF1t+tjIUBe72mgF/W2SCcLfYO59unpc8z0x07UxQZpdNd0U2odd/rS/1yUsN39nFLEdD1g3
oiYALE8HwsDGdDYAsg/bw2+Wpw6djQ4hqgTXp0zCrTOppsJylXl8ffmJzCI2O419LQdh41hpuE4+
oi8eUJ6Qi90n7O4Fm7+SFNVYRsUWYzjYB6GH+xDFWdHQpiR61OEsl5SU8+/7iNrGPi4gnHBpM+K7
NdSpYAlUZoJlm0FCoapWPa7qySNBNWFkl8biW6pwdzCJ3VCsrJa0MfUGZgAomWM2n4E3dzVA1jv7
Xr4qi9JNKt60q5iLv4oFJnd0RwJqE2IL3qNOxMn+Nnhwj61CAy9ErGL+QntbaWPlyl08jhu57C/T
TDKSPCpYDD/k1OEEs9NOgIIP+G7rmos0QsmEjliy9vH0E7pb3XnCbqowwvpwkB64qeCoZb2z11+u
8wCNzUjcAW6c1SzKnUEMUmCytz54E3Tr5P7IUPg5D5JDy4SiOBXnqMf/jBVhEoJyRph5tAVNLg4a
N7eVbBYfTitGSw0wSUvUNJrWdzCISOmuZe8fDjUou4Jjd71zISwyRoHJ0EDdiwsJH3IfBUl5i55d
VwmTKCTJaj5nMbadlykUyDBm/ApsowT/nbUbGihIIqprCm3Y5zDEaSTd9ws3b6u731ECHDYXRkX2
lgHnm0g4X1ZFxMn84ftRETEyfdpBgwLjChMElHVDDHfkGpZQeMc0kWupPPolL9uj6Dxmf91pp8+u
ETyV34wLeFrY1KMpy23UhSxV4mCP4HIVY7CadylVY6DVQqhTlMI7BY4VOZL7/L1ZXl0w39dYHsmi
8ggMJEyR58udOiZFXtP2jDpjEylyUEc/CeTIQWipMOFhu/QuvhhusfVPO2m9IrI3JLdJlu/g+CPI
52mx0tdIDtxdGUALHnf+UWPEsUs4m/USg8nReiIp0RkwEuV0J/UFfQm209FeiJakkhLF8lyJF/Yw
CdgAarMpW7saGh3go/k0l70QsuzWTScRJyH9mZJ+GoBUEaKboItZiiAnYPbhgm2rRUKOmdyQA/6x
9YU6fhqpjfl4G75pYukxMdBaQwCuRJbMD/ZBXR6+bNtIKHGuDELIMpwZAwOLYut3WpGF/hgxhDvh
g4uT1iRTMMHgVSoMrYWNFO/Jvt82v3AuZ+QssXCs7zceNQbSiMKzpYyA+4iEPqkPnN3NT3X9z2RP
p784rxN0X5d9qgde++Bz7ADGtvCUOttHislj0U0o+35rtT7DgVNXNpO/kcOqNmRT0/DzoBT6MLaU
B4wCz795sXsJwKMSm7r+ZmUx5pokoaPLVoWfVvRB5KA5M/iHG0ckcQxbiRGOXi0fE42iiw3SNgkl
Byk/fgAmmLnFFovlGc94M+ElwPlxhvn3jc7vjisU5FoRhQgkea26+8yYWtx1D32W2qOdPIepzbK9
fcG/mucrFElpsx45+fBs1gSps+Mcwpkjuc9TdjSXWZ7ax/gGG1uTALrbmXBXToHEihhyrxEpyXNm
YEELLsUda5IWGu3bzdieU94ntZq8gNLmLM6I9a+JH5BRoukcgffyMy5k7f3VU6U/JDoJPw1TATvF
Hk7db2XjuNLydknqQViQWOm+CtBPWNis4z25rocth4evGCU7XS6gaU2RUGYYnT8uGfwzS3J3zw5P
QnN5cjrBSMUBk4cbczPqCVfm6X2sD8A+WuNQzXKti0oklV8TTmx7nLbW+AuzMvvkWMticb+gDVms
AmiAWi4yzH4Bj++Zf0EBTziGslZFk+sjS2ujjc7irL3uAKyg3x9jbRqL4pjuuKnk0Cq6ry2zi8TU
09shYqObIw4NNbyki/B4kIiRNyrGI6VdIa1WqwfSyr8wJ+qS5+rhvK8N70C/ydpnN5AD1s77VC/z
dARLbqWQN+01g1cT2Hdi0DlrlH64mDl8MNxkM9TtRDi5hjlc6hWGoUy+eHqGcGdJ75bIzOXjJcxP
QLVoo9RkwfBeXbQibbZGkVEYI+5/FaQ8ctrscZBa9xApmWMorjws8BcMYR3IpMTpIhKcP6SaLjnU
MVVmusMrC995fCfomXB5UIBQiK49PJP/gsqmFmca2jN+AjJ6K37Wy2yDFzzSMzdwHJuQo3TRR8vw
CLCdR1eQlSx6zkPqFuVBoFJ1MReZASN9FnRA0/ta7rFuX5xjDgzoMFxLxXh4TtF3EKp0QHiuEAQu
OWY6f7J3y23h2SruRfhqspXF1Wini8cjBrvq89pQ7CrAp1Y6euFMQ54UTsGYPTxnJxmIIvuZyXk5
hBLSra5NNvW9cY/UlaP1qH5UcCt1zLA3duFU36Dwt66uNZyDytuiu19ABOp3LNej7FMZg/eQ2r95
sxBhp7aedovaR9Wkh+hzCxQCMS2w53U+4GBlhBGExPjpqNqxLw6CBHvJamS0ONgWPxvFVIhpH3HE
oWQHZmCnl8pgMh1vCqlLCY4t7z7o1J2Uc0CH92eO7MMAT4sDV45sxaHNpBgWrMDw0DdJDkGOzfPo
arzD58nT4k/lbEi6m6kt9y4/2/Nl31Rwlbt35+TWHG4H7MkA7dkYwpTYYHeWAABkPMpu0s9RuM4F
oJU2ZaPtR76pfIQE/zuQoyC04ZLh2E9yw7bhzdXkq8nmPMrk8Y2+MflVptaEPBhPSgshRaIh7Fpp
6jEWW6FaWE4vVd+oAPsZbaBoQSLk8jBhK6yua4YFb/bKopT6SKxSFIEpu/scAdss8gPMlK5h5MRV
6SxfIezruNNBFQEgZbiRFJndWV2pwlmCEa6ZnaNkHcLvei27mJF3X5U3WmCVNXdTeDzXt+nvJiYA
W0CXPnZGn6F5WrvuprXi3L1Q4E/+oTZc195yxGCE7Vssr6qHoiT95JiLJUgzqdGjoWmRt+ODoLkz
HWQY5dTg9sMeVE3sCG7eizbcSGe3W/wAGjPsQSaclXTdgJXelV/6sAKjYPMndWM1fXmnDqRIrEeg
4NT5wrHhpANPrSM8VWTrspEyqBKJso5KuA6AoqVW0A/OP/0kHlkjmOY4Nq9ZTKyaekEH8/2kLRbo
MsachMOwakrTxFLOIzSdG96A6vJpX/ojE0inunHIChuiVTQqUqtWI9is2EvMImWWhg7fDpnlsCSD
dzeCWCeiHHD7nb+hfQqSG0PuTwDcCjSRqR1TwBqFxs9urMlNLS68nlU3ws00gHSyVPdUk4dMCsRj
KxCiW9dlfN9pRzEARmLhiOTbIbjbLwnp7Q1rjvm5PiNo7MQrV83UkN967m3PSXkdSy9fR5uKEnK1
cs6oN+zcett2kTm3abX5UcaHaoP+7KHBCIXSDWFIqGLC9y/Gxnlm6RidZJpGKNAfP1PbwXUWKsm4
+yZAIsnED00pecOp7oSeY3v9iVSfLWRfXZpqI2GYYC8VBaUdYhFssmrA80GQaBOXZ9fiJZ/axPBT
CmG2nKqaqJS55kzklYo38KSY2U3Hw3urgtKYYwtyhQwDRHpFknffFFDHHJzq3NSMPGW6bABifE51
IPNWO/egcd1EuxnLxCB13TRr9Kox1XJA6agYsebBKxBKnErEpV1xnYjzdJyr61JeLULLiQoFemYj
KmQm+5IozWfR17D5k1p3GslB4QZE8BSSgiBfap09kCVL3qFgfWMGdRmpuL1oUX4mXU4CW9G2RffS
HYstgV8U8FKF1BToSALgbVtAr2ZyQ1IMskAWfWuuYjOj4nSs4y9BWf+AYZ4XCfENps5eo+xmKl4U
tAK7Sas8VygoerrzIlZAD6q2qK4I+DAFQdHPdrjYGj+VzdsdHIJtUBl+I3sLoyCEKtdtJm6R6Gz7
a2G+txj9BwFnUgSL0bttn6K6ZAxo9bhwlTqyy6kg3Ahy9c7RDXDzTXzh3M6hNS3n7SYSBDswepaZ
ggRbetqKiZ9FnVFOdy0/l+JcKQgqWbpWzrTsrw6JX3Y3to4dhEFXFCLvxAAFqcjykTCmv9MZRM91
rlfDkYu2o6k3cnGw8sbfSwzBggr9ni9pzOhvPlCx0DHMZtRWoR68grMxxCpCTGE77mdB2PhLNqdI
S+eUsXIm0gyYpmcH9nhcWPCCBrP1qj2KmxSixwMj5+iz+pS+lKj6eyx3VXrIayOBZZs/aXTKHbRS
8vTvpxTqScHgQPLOWZ2O4LgY2Sh8ta7JxDGJAJlsSCU4vuUlXu47PWh4OWgSzoD2MSQmtFtGYdvD
nXuF6KQRli8JAB88GdCXgm0fwLxb7zL3vBSepMtyRqVnaYU8Tcw7gZx+uGfA/XbZ4C+JAJ8LMQs3
7v3dMWHx47CqcBX30Y1CuOeAgyocZ/tgkmL/VM7zM1Dz9O7ejamWXQLSvBU3D71gZ16xsiHnfWCh
ciYOTAksWFxO2cesyn2PUuoN9kZYxLVf+gAJv3zCHa5myym3F+KSIxpa7tzrtquqFbm3CS/oCfro
6zoW743W/8/KIVQh7xURxoiY5yK2i6raskwYhRVXLWq8oCtKBJ9QHxFQkuS2AmTleNQ9vpCRjU8D
gVU5s47doPn2Am1mKP09/5j4Ho86yrTJLW1laxytxv++TrS6P+5ojVcxMXt9rD1DoF5wvLiab3Ec
4l2F7ZrXDNvSVnTpREUInb7H1ENFt23KbgnLSBOI3S7qKV3nMuV/hfCQx5DZj00v152xcJSoXV04
uXBTnGvmHK08LMOX9dBlnQmb50BS0uq6YSHCpaJvGCI4vP/BLBzg90ev89v+UxcgekeyXWnOVvk7
mOLKXnLdEyrkwJrzzxq7DDa2qHbqbPcFj+IJdTskb7Xx8NTfkAUJ/90uwqtcJN/+E28rhBuS4cCI
sICufOwI+8U5/gv/Zl+GITzmh7SNXorSZdm/8rDAzalMGmBwp6vpkgXfu+iTwvXyv97h16FNe2xM
+MCV0A34S/W371n7uQIpFZFiV0axoTVRu+5X/ELfZ7kRTLnQsqJPRQ3kaJjEzM6ycmpuSa3bC6Xw
o72+bIP7VpsTuNQXnjgz/4/G5jex/sCeAYqEAHvlWUwCnbcTLl5TztVG2AsEpoaTmELXog6E72YX
QlhwVWG3RXOlwn6mPilQG4sapDLSZj+TPf8LUCkLKOwLeyvxOGUIfyuhRI87vCdRuoWN3L1M1R1c
0EV1bxVmP5p0Xhb0K69d1+Tqnbjx4FIVp2i3DuTJorIWyrZ19eo6pckimWYYo/TNXsxxV3+3jacP
FyjK1cePU2czjSD9rMncCtpkrv9mtvfTnNT1JNXL77gp7aMuZhOvY9GlNbKXwoZDWVxFWvXN8t9C
gwWg4Dd6NIXrQCxjX8srV8ln9c7/Uv+twU+XSp938v7GSnrFPy5loxO435FBpKsT562pAQO8a0rR
VFg5LkrjZJSLuT/1UInrY/Realqf1bM6M9fqR7RoDzSuwx96dHeZjUnGzfT506NtYChE8rpFi3yA
HP16C/rdBnBFSnx0hCvERXLJdh+Fsjdltl5ZnMIvq7q69gx9YmQWe97qYhgT8rfP0225H34t1NOh
E+yYyOvH9DwyegvCbK8jz8qyXnaVHTkPd4fmsFe21LdDEoMkwxWUGzwgynp7W0UEzdrHNKM/1WHR
zzyftgQ5F7ymmfnDbBa9ifl2xfnUkVBqoyNmaQbuUyz2uiyqe5sgi6Vgj7WJ1qyhhp87erWAnVVN
pwjK6JV13O7B+7GsajifTcwADSEeJsGqTiOinZbr3W3KjIXojyl5phmJWIkZ255lyo/Hp9IRO4Tq
c9i+/2kCoj/noRT2oYhmh0AKgxL2UsLJdoiU/Y1/Xer8cxEug3U5cRiq92U/DuiRygTBzTeWIzs3
Le7r7ZmVIvrp8+QF/g3awu1ahoJoWNbqIbJokMzLGsElvQ83uZ6+y0riPmndQj/e04K/4pNSqxOT
hCo/etZa2VUt9QhzKHGdblUijD5sgvFdF2xVnzZ3MZvprByu+ttmYA7GfK00g27+6MYMcPvHGN+R
WyUY+6JkbC0GR/RnmjfeibC8pM7a0dnYnp5HyBRLcIsTKQ8hRb5xsTT8JZLJJaDOpMlDHCGlWR2H
wH8/nv1SVEoFPqn52ykwOpdw1yeTxmwgrohRdj/1GoeSG17FKpxvYVEhSWmuf05JcKtvHAxYFFby
xwlnsLM1kjjmt05p8KsRFXO/1DflJWGzVgF6mPSEUvirq2yd2459GAXn9qeQRNk96NM7GBxx80Ir
IlPPgU1IXJ36BZl1gFXNA4AomoNjSqvGr0YBnUXBUiaDr1gM07ZHMALlP9hi/c8Zo/10pJi+HUYR
xM3jEBhj61y8YItv1HqAIP4eVWmogPabHCjiEGua3UDItefE50Sh9UfWIe6DrMekKaAkFORBTaui
y3oc43h9Efm+ZAdl+ikoVmB4fLX+ktyiZWccW9eefmOFqPndyceNegLI1jVJE8Tp7r9eGrM4BlSe
VdmDV9/s9DF7WzNboaC7t46uCamIaB+4HwoYgGEWY0be4QTUKkOFIRVQvvtjKeiBLv1xA9C9TrCN
iG3sOQHhFjNtMjemH2D6chgHHQP4rsSLKtDYMzk1ZHV3M0EZQqZ2Ze5yNMbdJm+ACmT2MFRkZvec
Ph+NCayT6v+8v2ogmktc8wU9iTVmA190Pk3DEQPPIPVnPSvCIuOlG9NTEqQYRzVJHf/QvNWFk8AM
uUojlBY2hg0Ps32xCJi7R2o67GbSVn/Es680uaPLRk+JE7dTMDAZWl9CJFCYTiusH8QTnGVVgq4e
BGBY1OZh+vmGuGGPFzqR8CzQzpBgqxfr9c4taFRpOjve7sPHlsQgIKeuLIciM31op0hbK/BDp+/g
d2TRs83lrTjg7sTY8zbDy5dg+/O1ErIdMCsrZsNclym7EAmnXkSu92+uRQcbREEVk9ziXLFm1FIP
+iDbI6fJhL6qROsku4AQ2cA+iAMDbvyaBBjGFXUZhFV62mtmIxu0mBOZKmqJ+aCFg/nRporeBsfZ
9yM+FdsjJowUI5IgnpTFkZdVCJM4FFUHvBhoP1j2QPQi5QLjw+5voNkCaB5IAWCAVwKjPUYQDsfT
MkNcbdqliERdEWRk3T+ArKclE38/WoLAdgPAq2a0rgT/SLG/vL5BacCXpV3m2GPUQFHHYxXvNmrg
7S+J3bBhAP/gPbEnHF7Ff1X0Kekweh+5uI8L8lIYBXNfoDEBwqK29cSqq3sLVl3uqVVInPCyl0zS
Y6/hvHwz9gviV0LbJk+8u2nq+DXL5RNyu6wVReAg+zlLOgMn9jWx/SPnF3i5V8Lum8A77hFVqlmm
Yrmgjn4elEBfqWuD4J4q7aBvS6c3neF6gcyrzzMsgpXFS2RWdej+LMdwKnvFPNo5f4A2SKMx2pAW
kx2ybagl84E9I9mJQFXD8xbVF2ntHxG/Stri8EzwG3y7MAdwYb3JKLYGg+Zb2oQKOBzQ0DSHAWkQ
avyuChDhUkQAHeG15DX39BkBJZCRU6mrFRQJnCv+ninSGvdCEx8CZyc49Xh/LWduCNLIVtuECkUR
jbn9UFGtSquZgiztMWPEOX7/EXrDRK6Paf0MjgRHiPJSJxL3KxkpRBMFpMilhNyOQmArqOiG3M10
vrYJQcn2Cg8Oog2RrskrZF4MBumvGqKK+XuCqn6Z2FyOoeBMm+WUDEBqPu8M4f0ADkpNiK5Le81u
lZd6zGMNq6g6pQ==
`protect end_protected
