`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
VuMqHrS/xayS0NiRMUADTngebRTMa20uGoJ2x568TTodUM+4Xj8dbIVBgaFt8zKLsbW/KzVw2dDN
8gRsioW1Ug==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UmttAWTAeIeyI2E4omE2H1fojD7i1LJuxYxoqrIenLDK7GrToBE9ZQbyxGOOSm6o0st5sDPZoMV+
H9VT5ab1PhXyxpglLSScoQgMQpYHZ0RT/bqtWYI9S33rXKErdm17MfnWTSdBRAu7Ix7eBp6GxHI5
rH4otpYVFqXtk8wk8+M=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hyvJ5Mo++nomOEV79YebXV6OeFhphscP30m3xI6gx5/d9CnNbGTNCcm1TqO309b9bbk8iiZzgacC
6S52jtPn3KfhWRj9AibzeCSCYXoohsiOJ23FkaCk+mwEkKlJ3mDjcZy26GLjwcjbScJNTsm/UHWK
PfIh8HPiCUpa3bg23lV5ulKM4YGRj2sBTa3W3JHs9lKcUGiQk9bOc/u28OTs135SpVlqZdnYASTc
tFBfJN2JCW/4L17BBDrKeCBGTYwLhUnmFIdUzMWbvQ+mjBjMFto9Rb5EwjveEvWs87csNxKyyZuU
4BylbByYGAIJOeAfXEyNVDuYfcxYVsz83GQjVg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
apAayz/ZFVHW8QiTkiDBE53TYOOUM27cyrpNlZPLylxG4talg9Gs1bWtQMhuv92kudZyfmMDM5E+
uVJJL9tgf7BUEr1+4j+Bs5mj/5T30ttdVw7NZtOBJlm+hnyis7VgW4moDk40uVRcWGvW2grm95C2
yN1pqt0YyFxA5XTvaQk=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
T3f2toNxNbI/z4gSmTtpZtoPSBtD1LYAig8ZJobiZAfaKcWJhPBPy0uESvxqT1tSULTyfOYXy71/
VHSw/hyQjbeWrnnypABG1W2vNN59SDdPFmNmIFh9Rasz7Gx3MAGlOml71nz0dK+sRawYp7dZ1/vg
irvlz57fdoEcM7tFi/NkE33tR52W8KfEwJz0lzGQ04cPC+ZwPWiro+BHMU7qo4tuCuwfFx93rrVB
uKWgxmZH7z85MxGlI28jxFE/WYFBcSr3yneidiPyAV7MwfJzHAARt7LcOsFb6vQ/mpIu/r8ImUmi
vu0EWLSfp4vLOhHmrc+hpFewJYHknRAcDik5FQ==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
obcug/Z4bGoLdEFnwbW2QJ9Ih1MzA12XZ+BHpOFzikBdXImU2p6kx/taVMG8aKD0fb9peqKJkrfl
+78bTc016wuX4T2h0OeVEOKMNfDZxJ3sXpS1Rk8YFBIk1Z06HvCCospfy8NSG2wnZIXaB2JHOSAl
tliuIAfzuoMjmeW8+tGymXm/tGg4TJX7PJjXFGALfRYEPd063CVaTkxVCG+3y5pm2OjjWlvsdebP
syQUjBCH4s+4D6dFlMH+C9gj+3lClfX9TaajeeXZgA295mNzShkA/e+hiwdPFRhACK6efYDTvX/H
UCY78gKh+fLozqDExWHfwXLODd4LMyNvc25qgQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 423440)
`protect data_block
9sP0Vazx6v/wYVI7D/hLnJnp2A+ZLql17WcUhKXmB4+HZQYo+YG+NqZSvQTowaX1th5kcDD0QCuE
8CoOLzhHWnxWOgAsIbRICo/nOoaHxtXaCna2ceqeal/9wdoNo2iNVx+a7jJfqp4COEw2K60agIcE
DTGO0FDLiOl77AN6uClCo7Vqs2j1JmrYqLkBTgxtYXXDiZ2TYbAfhef1A7vh6WPsZdrj/8K2G3K5
PRMNJ6uhWfdPZbIZcLqbq3uzb88VfkxiFHK90EWqZc1t5mzbuPV3ncXEzsP0+IbSHOYkhH3BcBPn
OBznuxWiIcv42AbW19fb9NnLKme3CJbZltplxaF1mXUA0tcEkERThIsuqcpxN8iRNNosRirPe8W5
XMIB2sKgFeasPAOOPBt/U65TQ706Gss43nbIvf3aX1DFUIIK2tinRNX0yuAEWHzU+5QPoLQnTzaN
gpJe8K/2abiAnPH4wvDojj+/TIRfzmpMvnRzfitFqHxTSzWJ4iVhyN/UbtsJiwVquqaV3XdC+6J0
9z+EnFj8/KCi5n2aKK/2qFWqBADR6lWc3VRV0TQwydbPyUt2jBEfLy3fTOLV6Rrvul3vWDQopQ7F
DQ9w/EAkPh6krJ6DK8Wx19n/B0dcP19uJBxDvFUM/y4FQy44JP+znr5o9AO+0XqKh//TrDG2uKxV
QqRK4KjovmzZGo7MBIFXPxsT4L+YxIqbFdpTGxSEd3tcoJrJ2kwIZsrBDGSLp5EwFnuV+llhGcfQ
U3lGANoTVrl4OVej+nKj4bZ0jkWo0ULHbX5rCBI3xP78UfnbL+S7wjk8fuXGSw69vJLGHR4wNBSa
5x9WuDkRGiOmBcfMm4OlcTclHqOdwHXotKKpWez3ML1j8q7fKz1YmfHPZrPwCTv/QEWATuQQAj0k
ilmZRHPbqC/+zOLXBzsHje4AQOPbPovK068pjIwY7kl3vcwCOV0YnV3UIyYSvdKTw5duWM9ltLmt
6Q9bQ8Qd5WCRVYOKbdbO4kkTkyNSvUb6oucYQqTBOa1pHvYoKssVXeBD7ZfM3oXA1i6N0p/2Qg1B
3TsRVAm2OrfscIrxc5K8NZNKrPyccgrlDU3rND81Cp8FDcarPRt1ix8eBWvNgPyJv5z+c4Tyje8u
WOOW+MSUPqvCSwgqMZYDmt1Hj+UzE0/Wc/tykQNfZQ5hd+FYlsbpenneCsIZXkJ1CQeWzR8lCTH4
6+5l/psVz3QefjNNx28YQ+KkWbP0ocRD+AEkzAU+TVWJo/mjJ+7cyvtMFvXgLObW5gpzc2aoAVt9
TPlRjrMY12Ec7twE0yeceiVBSI9QObY8fP+RZAotRTuil7w59bD3Pj9TfyL6bvVzVdlV3L0R/QEh
9zwbujWrkrGO7gJiWI41QYie4UQeOuJ+pGd/BHkHj7gfViWJ+ilTGok0tEXvnyflA9VdPuAA5DOw
4QmTLIGHl+GEfQxXIF2tdd4FyIoi5MYJBKNtsPPwnoPrMtfdux33bPIq9GZV/26KgykoHEhqa/v/
Gtkk4ULvSpLoz7Jbd1hU+k/BYvuRepkcy1GDNEkfv+evGyousbiiZjmwnAQ2cLNLHntZW66QbCK9
cVSq0fStaAv0oAZaUzUzhfHMNFZpliQuZUf1YNwCccTCkyJluCL5azpApuct26/bRnR9jP2pNzf6
vYOOQvrqRjtCY0lar3A6CXTm4dgG64uQUmrit9Zld2eejGSIlXrGxzxbfy82hBgHfZCPrQXYW+yi
IAWnkboonVsemnwU4NC/P0LIchC5t331cCNsOCTHN2HgOBsxwgytZ0nT4tD9TGc7clDPg3HIzw/E
UnE+unFrlwi+bnlesVSluKb21qBrZJ3U5YeCna66rrsQdRn5VpiVl9zdaA2L7dmBfALpIuGMEQS3
avrjRRiFdDELEndV2m2WR9icacO560czZV96ySO8y2X3aVNjwkWm9+yMoQ9+21bYoGliqM1pA2oz
biYRXidEXxyXupJQhBPyw5Rm+dep8KYtsh8+u5BnLpvookrxMWTmEOJonCmYs9cdxJydItIPkvBm
H2TssF8+cH/+ONZZBHuWVtn3E1YuADihaa8cWTh7bZAosE4qawCAAesYVgK04OAvDJqep64YFlaa
3werA5+23c7CUA3618qXWPNR85bTDse64XZ/QBspassCexCrG/z6sXkDxO7t50aHqDHS+T888nH9
nzHqbpLkLVjEOuOB+issEuruANLTYTy1OAetTZX56cWFllqgt/ZurDtAvxmdh58xJkZiGyXOkhno
uSK8AU1guZLSFEh/i13ltGhKwYI7fuiobVOjOo65HpZ5m5AV/fT5t6ovC74nmN0EveQuIgLosWiJ
tSNQOMDPLXFDgcjGaIz5PTDYhnSar3ZTrYjRWMQ/OzJ0DunASxFUohQsVqVyAauAiVHz1CmbID1L
7mu04MWCxsdYuhcGoE5I7YnbrPNMyM5ySsxy0QiR2bDz/DVlsEW3VsNp4mObkZKRw1Q9fePBxFLv
sad5F8XnPhUZPi/70+CzsluBoX5rOZteaopqnv1BhF9+YcZvPnLWQga5keEXUMz+60A0tii19ujq
36/H8+Gz+Zn6t5ukMhc7EnHC3keIIlxYfKSdMpPn1tp+0fBOGN453KMEfHGZTcBs+j2oXYwWiWSE
F/wgfrKnhxtmQeKWTSu9gTj0RO9IUTMWF33Gghim+qni30p5ZBfiP9kAOcHHtbZlz3pJis2V50SY
x2/y9ZhJ2b3o1uyZg7k+YJAAIWMOVruv7p2ZL+hilBhbECNJEhQSm9QTZQuL8/LrJlBwChw2/orD
3AgsNaZD0PF5Rm49Oi7o81DxOitrPje98l9FLhiE2oOhMl/A3wRpxYYQ7ta195SBi403ET1pv0Iy
4XkQrU6J5U+Lpg6GipGQYgC3v5cvHdoTEw0NFcAO08XzvjJO8CfwkXJsPgsz2NcMdFPCuBxr7pu4
fxe/atsaj9Vp/4GZipWn35L6LzLLLIHoxkObV94gcDR0QCi8dXZPEILJTYo7YCU98dNOzbHN+OVZ
9QsrahsRak/nCG+PgyOY0Kijrm21c07TAeMKhmNhZz4iYwsvv3mzhEwsifXjyNIS52PBKXcZ5/na
kXSNp+OI+i9eOQvCiMjm7KETFp6oyDIX6Oltxhe4Usm1EQtQ0lhi4IXi9cqrN5l6QB+bEYG2/84I
m/Ehee5exm1tIi036UBzhpmbWrUGhiiN2vN1BcfazqgFtM8C2WAxFTs+NTpuHjRAQn4oew+R/12u
XsbAR3uY8iXPPhbE18wY4aOhg+Q/B85Y4Q6lkzzcIw2a7U0NJ0ej8U6UY940KWtILxvZqcE3maUZ
1D5vIyo7mY2JlfQDNgXspTj2hBq69atve17vf22oigbD/XeMG5g5NrcE/Iqfb2LlvyLmKsF8Z8lN
HeyALJbeT+LGgQrGulxQ5fa6h1vlR3Gtn3+gUKiQFj57B/4dwEotWre/YA71FWM94SpoRjR+Y13K
gA0QmPwEQ2+o29fRMjvty9P3EJw95RHDlkUwvAY8lTYX6zTavQFdAAOAMWKNzRGTx16NMPP9h/+/
AE/6UdqSbQdK0mlIy3GS/RBGMONuXBBhFVvjd+20c952Ag8OkwYM5zJRVWWomS0DK4YyWCH2u4xd
MgWMzgcxor0NvDtoYRbnj57F7ws9/tDqEgpup1IIGPBmtDvos+xWI7AzMXa2QrayNw3ygdifATb1
l/hNbeiKeHTM7qorogFIrDdeWo+C3Ux6Y7lbCdjSP4qBPsvidXJ/rXm7xDiW0oQHOlW++SVRo48L
cyvI+h1PNyrizNRod4ZdAOynNQrd43ebrWFUvCN3TFDVKgRBm2dR/M6yotcRS/qp57347Nc6KyOK
rg/jpMfDtoEzwASphXQSHh8zn4YVB+wJMmXSP3zPxxFSFCTFwE4I3fZhB63uGDmempLqS4ZGd2xo
8yraIg5Vo26+bJXDnOmqXTu9YhniCjaKV6K7dme03F+Sov0vPd1Demo5AQ7jL5/EFFhruh8zUD4r
pR3TZpT+gs2Reg/wLz4eIW5hl72fquT0r+f4hXOAgOS6imo/wyi9uAp5J4B/DWBqURcDuKpdB2sX
cbrOWp8QaxVF2vpHGq2Xhg5dFjKlYtBUzto4PT7Ja2A8xG0dsdAwvxmoZWrPccQDr6eTJPa898bT
X8URvCZFaydL1X+mQZkN4iUz6v35uGu3J+qTXEYs3DtAmDBFzUXsrxZ4A6RYaqQYMKfpU7y2Xdoj
YrWKK3/M7B1YV/rPEiGvGvEIPu4Al9Z/FSXlegQQNr3XlR1vDsY6nMym5tmrxPX3GbmK6qXoyeQ+
PSpAh6EbhNWUtvHQuCTVny0GJZyE8J05vIN4bkVVU3SMWBZ4XQ6qHRrZ0l3sp4e2TC+YKdPUvd8q
mstA7i/vGEbW4F+KSQxJisFOOy41ORDVGXyombPZ9aA6hrbgUoU6IBTWEn+t7QVhT5cHzeqAW4Od
xcama4PZCSUwps7oFSIRs/0EgS+Dw+Ta87nHdLXWM4czfaGTprzawRf57pzQCSlapn3+zxfmSJf8
bpqghaEunPzr+ZhFn/e5esvbNAInXyZb38H7yNkBlRplaVzws9iUUDV/pfOQxfcHTtldvwJD95Hk
jBz+dLgNJWx+ADzr1/1KiK93W5w62IDY71cTrvjuJ+dj1N2zFmBFMlv7ExRndZcnQCRmkH/2dQqX
d5HpdocQ860u8ZXwOvmOj4vkAelVTQoj9VvQgJY3YINquYUFJuKp4+cf/2BdyEVEgOf4aY/5zzIG
fcxmgxdjncWgexK1lYPAPewPfzXL1gmHcpHppMveTU2shKa/8oljhFRZua7crfBzwTsoATKSaa7/
QFmmBnBMXbKn2qjm57s9iot7yPgAU58JaROyoBltNsMAQNU2oey48yaQhBSlnLCFFzurtCRptoVS
6cpQsorldLuO5Tw+T4ggBt1rLlPJPq5PxxQa04m7xQ2q/6kkxFcxT9lhiRN4xjRZTB/MJ0tp66QH
U1KaBYgUqwuNSkPvZhqbeBulUeOxnXbzESwzLL43fIrJPS6wCk+YQZrMUt+jGQ8QNWzXXhR53nOv
ZPIGT4fa5gLoUoAQItk+qo8GqJofo0UM1Oi2tGNE97ywEYyyen3TyjBZBsSai1JfBwVYHVA/O99K
saZk5AASzAmcF7Dl6NFOMrk46/hyymIccGTSp75XdiFyEPNzY2skDQ9ECBqHLbU42a3i3XkOQi3t
lnv4IYOEhLrOIHxx3LVZCQM8JhlvnYcSxH5yQg7bQgsL5ZLUMJvjSvMhNkeKZ3oKtr6hWvYL+GPQ
t/msO4eG5kMZu0y/dknJRQZE5mg7QKZ1doOB0IBbCRYz0jdxMPxL0LOJAr955H4cDetCmiJHfrZJ
vFuEXxY679TiBji+Fl4AXDQV/kNqNhyxxW5Bz0fAADJNTxz7I86XE7CtAcO7AoqKkBE3J5ErpaGG
319yY64Jo4VnUmtZ0C8joav+x7FQrX0cIe2wIoWknZwn2uHLy2jP2juplGRca8Anrs0Fylp4eA47
cgvmbEGG8hZVTbDxx2BXxifBQNfG7PujV61eV/N3sGhHYuQlyge44G0ia0D+Ixd2hR4sYtEJIi8L
IT9LAILphDG0hxaEoo/aj+pHxM1vAslKkwYEcAwFSkLAx3U2RcDvCzx1T5P0dmyJurMH3oPsqeO2
mpSDImwELguGiLvLp4kPAcvxbuKPmEtK0iNpvDInlIdNqC5n/knG2KbVJxj7qmeJimBWJJ/Ag7yS
pPngHVsU0HrrLuYP3E8oEV9HQqlLZ5AU58pYVkFrK6qU75c+ioSmsqxSd7vXyufDyvvdgOkoOvEH
3MX0KzPcKFi/fZEz21YMif4O/OGwjJI56N4gD5DTUsWD5uuR6W2GomXWJQkDglV96lnCrrgzjprn
ExL8PTjlWoyxfiIboGvaEur5+sKnYmy6gE2YpAkTYeXRMp0sjkw2TsV1QblpO6qnqpDsXKYp/rDo
ttg3ij3bE+dJDKYYP4cyMxi8qsG0RpuBtqdTwggbJcPZfkag8LW/+BJqTOyE0sqh2AadGaNeGghh
4S+oXfKRd1yN9+hn1UYxNFhf1mtrSIhc8DpM0SvtGKNJPM8xqGX7DXbDunpVW4pNlmIwyP0UqZOb
zkvjErh5ZmSD/Tb3/Zx/UQNae+CCasFhxbuNAhDwjWFXKTPZh5BgOF9wXRzO63uif+c7GcbZGjMM
4s2eLD9qNMf48BvyLSPBM/PC0hTH32nvmj8Bo9m8jg6+DJJMYFjsknMVbvCs45H1NSxdzl61BIWT
MdJdmSLiLQOC71+zeTINRBDgez3NEyQa6LuMhgxv8gyFEqoXNpHJ3nb+qpih0Ea2nyLyzitklr5j
iQfUxHpI+xZllVoR/dv/VdPnz9ymnWIPvc6BD9n6CIpNZ+OOJWcMnhChrVEUf/SRBkMyp+mWKHA9
o73BZMcr4E5Sr7er7tOI2t2ImT5az25Y+h/StXRXhwXvRl9Ifq59zurysqgwYJIlzk7bRLyHAscX
dpauLXFCqxWv25zGWNqYXuKt85iXWgMVIK+AO90dFJEFTcjfQVi5MDmxTz3Dn/DygqbjYE5g6A0r
0muypYs3ksZctCoiQRApx8QEQ1Q1xHOr7Mt8HqvEHHtcymEF67051IgWpQPnjvtu/jl3rNaeycvz
SmIkPUu88g1v2oVi8bo29uzM6anErBKyQooK10MoEgx+fWGxACak9tirTE+t68rVqwzNRPEGIFwx
iQDJFRKaGi4P4QcCd8kIalexDhVJjmsIHMm5nYFIgRfG9aOFxxMnNUfXD6nO91Rif3B1Td5lRJGB
xw887k+9OhJrtEHwFiX7S4OHiHlVX08DApBz/cuNqa8OOGxvu2aYOdXYowwqaQtJQJbm+q5SR7zF
+BcfoutNw6KRDYgdjdRnwXgvhfCH5kdKdl5A5lczd82w+wXu3dVyItUimlWapVrVLgse98rtiuBS
/6iPbc7V9+wLNiJGxnJWYKtHSKaAxwcIfQIb/D/z7roJ53lRqQVgQ/FYwogbfrU9DGnWreFU2syN
idfMno8vl9hdbNXcWLKSMyVvBgXYlRl1MjUkKTFF7Tt1q5OUX4zZSF3DnpyrPVuevnmR3qoXnK2Z
qZPqhlirAX19ObRVcBnNgh625k4q2di51VK8rhARFX1rPmlZP86HzpFTBh7Au9wnpGegeClm6eVG
H0XODArEkAjUZhmsv5CXUqsw/oiRVVlaAzRs8P4WpiS8KEv3xzy5Ibtehs3sH1i8TAwXco1twEzq
xKUcUYr9EKr/+7Lq3fQqkljxB4exZhaOcXCsFDfcGpGuETCj6FhxPKdB+e0sAqPOJTjKUqy2IJ6n
ITYDktLGVjoEAq0RVWo5CyGXGGLyPYJbw2hzxrPpRVuTzL3+hTdnBEhu8D9aycsU72OQ99l7bmpr
eSGae9kibdUGuIGsljPBmpsUBsQcVgUnqPeCW0mAzAm3c79yLM1rj51x4/9gVKn3eLrvO0HOoljR
dNZwmcIMDu64aSlIadVVwYOPpb7ST6b3qj1DZsDyktSyxAHdm3eT4yh8c+MeryYXE/ptk2Xun7Bl
VBvkWHJbZYhRRl0EZvk2+Vvp0lViw1KKCtfh4Tu+/201m3y0VVal4KOWSy3DNInTYf2K1Jqdt3ym
YtrTbkoFpzndrZxTr7/52AgIsayYSWZftEzrU2ynCxnL1wEpp+SWPu67JrXEWpQFRkxwRPteGHeN
UTBEqK3uIy6JyFpYYGKXub0hVh+IuxkAHOHBbkw20z+WiUeyHlm8FhI6AzekNHzqJf6vPavRl8ke
1+ydsbmU183kfjA9NduRxats4DmI6LkFbWbc3aVt6kQv6s7vqk2ARmnun9uVNbjikCEUZn4JR6lQ
qikGRq4MSts2sDjSuZDFgsS1D5j+mpC8imNxKNtpH/G5DZOMV6mF/AyYtKx84B7+NLWnAuUBAAOf
9i22oE5mCJVuVOwlJWADRC8rNOrbQt4tkWTqQTgrFqSiTYOoYCBwmVoRsWLQBXLkaVGtwEq+5D2V
eZztQkdbwobKb0ZpPHss7NSEMx5Xu5fyb0+AtFgosZ5Ak4UMYizx2ZrE2BQpysZlzhOXFePitBaF
7drLE/Nm0NaxZCRyudU+eXlOBX3LOzlGxMQg7BZ4gUfnDTugsuR+5IvRxYAF9pNZofSxSIgUngHG
gKz8iJ77l+TiiJNo1lT15kfBp//MQIU6fkagqSPtx+yccdLSbwefcYS1OZZ7KqcGPSjVYOFeVcd9
UVrEXzHycx96QmPHkGILGuLdeGWrxGKtAOCH8Gu4H7p6O6FnMUoI3FzZG/ed2U46E21RFpimZlE1
cxK+V+gMF4D0OIv2yhDkZxk2XMrdNPPF/VsEXQoo3t4Ieuhyr0CzbpMkENSd7k3TwDFP1oNK3fSz
xcshklqsKtTrZG2a5j792nZmTmLCDssIucGGrKAmZGJIufty6uRQNjnOZGHMU1l0QgubeINujjZq
eXL3AImULnhZDSG7HTeQJgFxeWnEExHDrBCTTgTcqTroB52+X0gBuCOaRIEwEyWaoIEtcUZkwvN6
KPMlD/x6V18vHphcVDONYo7NZ+a2k8bCBzkZL8QkshLi5jwReB5VgZMmdNDk+1a2eKyceBbvnFkn
qWv+mA4kfNW4BLvVgswvsA9RH2tRDASAzc7RrKIiKJWfL6p8dyi4AdgL+L2924BVtl9bT+yvOaq/
XbULAp1u7ECUReyKRjUiLVQ9GsMNSyeVA20+zoqOttJgjt5IM7Q+RZmDMrQl/iz10ytvXDIIwk4i
SBmJBB5HLohX/ILJ7wzysBA1w5YDkTXSkoKalwpaH35UD38xSOsOozFVm+KLb7I2xW/X0J6VxdF1
uE80N/KJc8DFN6hJKkOQOFDjh0WKJs7Gzh6a3JY46xZ+dRciRU/alRldOsHMQEHnoc+L3j6sU5t1
q4LT046tFOKlt7gzt72JmjysJjSHozuC/oE4UoELPYKwlZICoT/cJ6ll9EXDhSu4LxzQwxZ3aqOk
SWVNSxv/SIvMbooRZ+rqCd/xGcDZZkofz/ZNqs+wIWED6dq0/Ajnz3brkGpTErImw4yLhoK7svkS
4wNOI9KUIZ3a/s78nie/OSC5No21ZP/1fp17OilQNl1TWMvMTPsPXuokuR1jxzl9kJDhSemeQ0Gd
G8+MxKKYJEEfQujiEkMva2gM2m+xfyfUzGWXOs1PwvMnhV1a4BU0ho5jumtH/Jf9sOGE95tRIj/m
aSsnOaiOP0yvE1uqvLGi4CpUuIc1wB2IcornTn3cMSlF8KoQDXASpY+9mwAvu1RHttmOcE/8fL0y
L8UmwmEoE9MdE8bjciSrQaCH4HnId2OCppGq6b1DOTrF1CzNNGnBUsp8UXI2BdvxoQFnld7ouII9
PGZlFwCDMHV1XDK8YmRF8Dy7AB3TlFrffs/KWKgp3+EP7KeJOJ09HWB+xfG4Om1gbvj9C7RK5PFt
dstU7yaZ1YUQnh2rsOju+FQCd/EEyzqJdlt95/K/OpEdI3e0jBWgWaxr1VX7qg9LO0QvwgpA4Jt+
RVV5Mgjja+8ucn1iv7PXWxFYxZiXQ+G+eYwCd31//GVNdAFt0/RdGFR7Tz75Gb2Kjf5476nf45s0
aP6h64oNYPIWyffEm9G1lNFhuhkjEibroRr/OYJY1WeDlVx2PGya4TxPStmQsMf72oCPYKIOH34V
TI1XKrslnu0ot5nEB8avCMFmRejDakZb793se45F/Zoka0lcQDnRJ8nf2ICG93Ga9iItpbCWPWRQ
ap9O82E6cXs5pTAuCuM5v9lG+Nauz0j2Oq2K+LYbCdaY4JXlU4pgGF0MnHMomoQLOzBIhNY7QrT7
bRhzieOM3mkvnz1SQkuSkN/a7c+GlFg/kdXcoxLl49yP0MOm2OJce6IxMzT3pT6btIrMqWEQ0EBo
x34JOR+J/dR8u34AyghohWn3c2mfKzDO5OS4dSpvrMmbTM2juG+FehKUEZ+bg7l+6+VXBO6K/fZV
h8CdoHKpeyTVuKHWpNoTz7cqGd026ZanaCTPxlzlVAC3sY8QjdO6tklZ/vhCTdYh+yykzm8VX5se
1CvhCEYDTX8ysAhINzWpgsyVXdQJAKeTHkWLopLy+uoNy1XSJzdo3aLDV67YnASJtyFA69FFz/GW
RAbjMuy5Ug+Wmmtzs+AoGePG0sKrE1s7mp0pUAsR/+cETGCPgwhJGpVhfq2k7KdurgtxgiCQaAT1
XcM8mgc8rsPmA5fRd7jblZybwDVbgtOF0CIqE56XGGqZozFFFn94UN4/I0QDdl35Bx+LTC/cd0I7
Y44l91Hq/QPcW9gKNirZhCK+XO/EdY7sDOf8FI1UCDsyDiuUNP1pWZ0udBCGfgLjuO4G0Xd7wEYi
cT3QB4xZauLNrAkFfcVHKUFwXeSUTukYdZaofwZtJqX3Hs7bZDzHhvjkRtEp2n2SSX61ktNtGQ9t
FtUKSmhQyTNGiUJtPcbS/nmQbesuObnDdSpZoKH3XOA/pFDHbHASknSzdNp+vUDH47ZZmYQGtd96
xeYnYse6vlOaGzcPCxY9WyEk+UDWFqo/y+7AWWEMuRyGQKQnhCIxkcykw4Pgd/K4u/aP9K4ARmLZ
wzcAm4BZX0x/YnUgqfs3EHpVcFM8emWweBSvDt5f5++SOmIizsIK/AyhtrCPcOuOd8OEYzWcn02Q
U2ZMSM7a5KH7rOI9fZnTlQzaey+UtyRlRrYYzZQ32udx1zpTH87UUhcX372cgpp3e2dDzoAs1YkL
k1zPDLdDZy1S/VDvEFgAUkNYFPC/C+/gbcfkCMrFA8l4oa/M/fRzuI9tkOj8x6uQn0nH6y4XocHW
08E+a3CaniGFmF8yhz1AVsVAT7PFj7ZfDqCdrhubLn0A4/K04Z1GQcARqfFv/uTlHlVAeQxMFIpw
0/gqF+3mom6FW+J4kywMzJ/2RmRUbz4kY8g1YDuzs7HtAskSms4Tr8jxfETpVc3An+iJNI9d51sG
hJd56pOHNGbwgN0wMYM7LTRIFBOwmN6TpxdeOf+5N3cx2/mq1WGzfQJm+geb7D3ebN2kTh/dOsWY
ucLnuhE5hbY3JoAaePSFz9Bfv6OCWG8Ohu/DSOyYqQkl/c6Jt5j/qUan3Eg/cQJKGRAI474ew2sy
G1iQcF7OjKxN75Dw0JZz3DdrNhS0LkwsgAH9XaqW+tuAV0FDqlWn4Zkm5q7afLSCyycuoHNPeqsz
GdZ9KdA1eqy9Mjfm74A/rVDjwDaHH1007Y/Lp7B1E1Sx6gl8VhIbRiz0NCTQkdvquHwb/fHwRECv
2kC9J6fB2hRMBjpHR24gFY1+VUcntkMQDswVTOmWccUMf9stXKPQD75fXsEh61xbA6fqE9CBjMRU
jrlbbiPqiMc+ynFcOq4b+vMCP2eTj+bfIt/gnW15JNpRx7MGYgY9ao90HscIOa2JMvFdonTBHpfG
m3cH4lfkmDMw5yRIiA32GZk8hZ9qGIpU9z78zSJT5dPZ5ve6nTn0Widdsj47TyS7bH/H4AQ/5tHt
I0OqAcJopnROqX28o8okNH6rnXYd1pbeHqURssex1i3c6EaLSgwXN5cIKSRY7Dn9YX5P8CukLAa+
KaX4RNzzq/5yz2dQ4aLsjKcx+WDQne+WXQ+O30Nzsos34sqdntS3ibbuFiKEXCdhRPg9DHugnlef
OY1jFGiFodaxpTSoyOBL8zdhutCnS0TnkMeYs4u3OKnEmnMtwXSmkCrtMaxUR0ZPLfyTXJAmFdMU
77QNs2yGG5ugYm0pG3zO6iWfPtNQKKQnqyHiJYh33og7c+gTcg9ok/5aATxUFoon0cQ/cNDo5neP
fLVpvRgrFpI2biAI7qa2+o4g8+nadx2vKt3G0YgBLK3zODHIhlbgPRbFhYQndUC2Q6igTOuV4cfj
yXS9e68tS7JL1DhJQFiu62G2GsQGKKfsDJhs6rc9JcCaFJlS05aWtLkrh6u5IvFTI2TM5oaZZUSK
Hkgtxqxb2PUsRdaB/T/gLMk1S3SsSi1wkv13fvEl/ksQ5XgLh4wV6FMPasV6qbyr7h1G8sEn4TLu
V1V8Z7dIV/PEenPgwgzLlKDcjfP8W3IeWAfb1J1xCKRG6hBm5tT6ivmKVsW4qbzQN9wM8N0MdT7Y
XVkYgBGO4Rfu8FolCvtMG6I4jbtftxUUuhX+J++TraAgQ55vJaVecwZJTs1M0ngipanHUK3tcfGK
qoL4Z3BqOdFjloK/MJscbSJ8b2paXtBFajSa8mj7Aw+N/QTKYBi3OIASIcdEgqmJrba9T8MIgNHi
NbiX7kg630fAaoClM/M05kIJAUvcaDHUQmXL1tAadRAAyFj4QZDEwQ4UyZR2xOPnO6neEtMPZm0r
AoxbWjncxWI0k9U68MeE5VkNQiSidB6XVu0NsBWQxEboWrTkPeMWf7hbVo6uusdFp9pfwHPLXt8F
lnD0iGvPe0fV/nU63lneMIMBDugoz8g110KClT3FSfa0yr4BVYVAycd8dVUjdnLh9JB+iwp3GV3e
Z9C3J6tnuX5ZzQuPx/eMGM812XDQQEEdK3dS3W4sBncgjWh9srV5dqB5cg/FtPXxh7P0yK8LHcEN
gE0ON8pSkV7s6rqwTuSr4x3PCi6HVp1Rdazc9a/YYs+OzRNgqdkCiXtmOx/9xThlQuwosdskdAFH
jb/l/2PjI1M6WXAUcXndUdAEoiJV+cbsqXOG8IWIj0YLX5gGIqw6cgRYYufz8YXpA6683mlBlXkW
/M1KkUISLC4xT85s5oaW2PRA8A8v05D9iYt42sHgdX0eZBqjVJCdKqiaAcvvHWVSGZQCiOjD7LHP
9ziex34o+PliOoKIPO3OEheFBlZ+sMzXI//LczUns20ItKMq4+FFvYrEiQVlcYFolUwEVHYKiNNL
i0TTadD//tEAfiX3PHyT7gxRZH4oss9yV77XGka2Wa21MAXTQ7ka++Rgb8Gttp7S5ZApEsjIeZeE
u1nYl8JgFEjQ5CldknuNVxHlLyFwmQvanIAySKZJzxbbfAlYuuihKG8EtyBmonfblyDlGbCJr2bn
NfpgjmjLAnR8n2qQDJCJDYVOKc/wQHl5MbJmS3rcGKWIxYgO6ZT37EWpg2iKtb4qGKj2P8n3tBC/
sRNLEjHCLxLavGbDVdUJfu+8e/gHBypkF7Uzvm9W3KSjZ3iWPZJruGadvD35yeESMM1xXNR5YsNK
iQslR4RqlquBf13cGlBzpMfwnCWc/m1Zt5IB7ffCkEgIBaX+e0tsvK1VGNukZpG8rTaWmk2iXse9
kmcrwgbD6LbVMQzBycZDEpJ1Pgsq4zGkKSezgvZI3pT49r5s+1PfUW4K6l9VlPRrGjG7IYkHXljD
k4BokmoymUDA0qzVHLTQrWPqHFEFzJy5UVA5CduztLfWvc2S7Bvi6ODOtCfFuN29G0g/5chxWGEw
X2Q8CnJFiLXqV79EPBHMjn0t71tGRj7CwkiKOdrQZMOaz3oNnfScPh6BBMu3uYyCP4K4DWdvS+PI
wtI+FJmtBXvZrAeAbevmYhZyx3XX4fdAh6iPOV21BJaBf9TWtj+iLFzqm0qNjCtM8vaMmJaq2IaL
Y3gUCnYuTTgXalPvQ0TosYYq6INrFVLb7RPaInvE0DfPMgT/Klf/3JV/P1isrGRxZN5L4OoD5yV3
aM20jAy6ZCcQrCGBe2YAAJlIMqhf3jyq6Zz4lN88pjnwqYvl9jQIkFFSNE81fvHLslfdNujGiuzw
ovdOlCgGdVj330I8krDzOzLeuEDObXpR08zl0N4/huj6la1/Jz+yPl1TJa93ryFvn51nyUbsYrdM
gAHtoV1PkBOgZhnrVEY8WhIq0IzTn2VsdAkm+wO/3VffiAnkTPmRwQwR6OU4+nZQOCKFf1mktAK5
JlKc6H96NoyW14HwfxQKwTmdnMX4CSMDuzeUUx6EmezT/u+0An0H3rtIWV3lQOMQQUcaIGJOybzh
4LusqbofQAHHMDp5T2PZo4XWOKiVrnFslNx2sdfBgpbByN1eCfSUTZEGiTVCm4Azu/ZbB4/RUEpu
xkjPOmUuInt+L6S155lYKFaGMK2F/CgbzgN/8o2/e5WY/9q/9EpBSQjJOwnEfdYQpoQX7r2VoxFO
T08S7DEA6XJQBo7Cnq4h86MvO7NAvQ6wfA/Q6bxE/+OzvaNBd2A6iwsHVLdWQgWFFeXdBMlsjYiJ
p7rqz76p7qi31+OBRIREcvzlaLGw7xdRHdqRhaw4gV92HhrD2z2KrvQR04aSkWiXwN4tZkShwppM
3hPQnunLvj6E6KRt6cTOWE1n029+uyJhvA1stHOYzQCFRTsgSJHzRsXceFbu4M2eDdtToy19XEDI
KZQTYkiC3wvvJTZQQZBmnR9qJPZkanzvHQQ1Wn0++WtY9PlHRORnqvhsmcU8ubMNgjA26r+4mlPF
Exl5Oh9zh/B0RRPn30am6LLm9IZjVwNk2Tl/55a5B3db471YqD6T9k0honzrzhNUrK3V+7ejHh7O
9FnieI6TWFz3YHhBhnr46DcnvIQDE2XBAhqJANXKrxxGsnvtzWZFbwdIgZ8b+8tkdBx9UWeXmrHh
5FD+D21QJY49//Lr0qj1HvX+98GGdv0LzRqoFt/osnjZU/PYNjCM9Istyur14nEO2wnt4r51bNUR
5jBVy2TzaXTS4LwwDyyYoJMLC3hYQvtLERbnzhxpiIu1WMf7h2LmR1ACyAzvj2TSSYeH/fq8B45D
XPRctEw+3CT+64OxyeAkvTzmplkZeIaRQ955AaW8Zmu+00v3OS7hNPfHU2HnQSY26PpYsQDIQKjh
dIDLCgaatGImujMvsPz6njn9wxqHT6+0HUL3BzvBna6dq2STpv9aczpgn6sJE9sNpesFtYT8nDmI
IiTEugVys+2fUI/dnXYixuUG2UnpZ6wD4WFkJdURYKMNb1KGLeX9rwhjiE1ymF0GVaqUs4GyMQcI
ZCTYb2UZzImmLIOVKRd1EuIIwq6dqCRZH0ZIiRajOSb5c5n2+8012U2QFg9R1Vl/dLbn5Ku1zMyg
Y4CK552ND2ys+5x2+8kRQ2l4AmdiNp1Lo104zjEtNvFJVEwbOS1b5viP9ATPNJ8xwARky4YCVtQA
uoulifXtVjtd44dkSHNhIB2+3I6VMaVwbzKEPimnDT3vCyjTGv6Ol1YSnB8ctLCXIm1hB6c92WHO
xCvc6Pwz9oWBB5jG3mqlTQd+9HhoukTMWVLkrqlr+s2rEpXv2ZEbnp6ud61I6sCKkZzxQYojw3Uc
YvjRm42puzh0skbPAk7avp3hjE4lEOM7s1LnaOzY7/MtJ8de57MtiMcWQUcaFjtSmYO2hEsdrCp6
8ifvty96RiP9B2dRy5AZyRzPaJ4JnuGCku+p5ihtYyKSQeR+synvz1qVebIoXFFts7c9Ym1301IE
Q744S2voN7B92xnCsqgzEavnuUR4tXaMfWrxWmv9Tg5H89MzUOFI4i7BME+EF1gkc9EqLLpHbwzX
AASPANW/ZjhxTXTpPo+wIolQ879tWJ+Cr55xP1BuZKMay9ErZ7WOjxAkDMV9vVjoDAuD2mbbUSdS
RoqCTMOWfj4ld8K8bq67EwuseHS0sJA+TkMaYy3V889NAnlvPCCBwf32PUwbQhn8+iOSNXOJCnob
Qqa4yYiI8TKRDj+ub2iXgAe7hsXgzYLI4wpNxP7G2thXKfgeGz6u1LOXodRK6PMSnHIsEOTcZz01
oS6+vL/6VG+7a27FzjF1Yxc2YuE2RTf+JGhSN5hcI0YzHpmi7KyPCsVN1+fYh5tbLl2HKmFNnjUr
/gobk0dsTzHYEufJE2dm1J/FhLgSyq2OfLRxISEgIuWUTApro3sw354z+BUMTB5Aht3pqXe5vK7C
qH421zy7w5SM1z9DfWRpabS3g1ItaJWlCgJBzvkZEMCa86ymuNAfrQydhEwoyxqJuWBgCaLRaP5e
UwOsHEqSzMY3Vpj1iEr8zIuC08K2H0PfBVB7Ug8YIDPx8vX1IEjMmEtKR3L0T+xUtwg75XnafZA2
d2HWO6u6fwIsElV+++MincYT2tRNLco3yHugrJfHewRqI2sUL8CynWeQRBPxSygP2cmUn6UqEodT
LrwVxuhRamb6zr/VcRqMJRiRcFR0ulcjDlJ9Calcs7ADaZ1lyMhVtJNHVMjr01nqxpfoxMsWGIe4
Q+RanW9T3khdm6hV46y2ZDWKIHDTBi/DEtywQ++SG9Ujdc01O34u7H+u/XgyHYGkAlveReftFoHg
83fCsVJBEWvSOnN1tT+sYkZTsfqUANzzt7p5Dl6Odjx3k5JIJRHbqEwALRXRpwjguaasZ+5lyaMF
fxUXzMOWgEs4OBKjnwfEE0rlPFBsx1nMUdTuL4msLp8NHwFkLxwFrP8b++u5Q0pUij1rjoz91tfp
yiZW42W5nTtU9MgSB8ikwxp4odRtyeEJBZmIn7m+85/Zieg4Vo5195zsjxoP5XqnuztlVyr9VB4s
skzbCr6gyzeGP3BJy9abtA9g8G8ETEq6XI1XdG/x1FLpir43SRFrTFGjK9+wsoVIdLwl9NhrHMjM
aaDRmMqP51twrvbZvgL1zvZJz+va0jMxnCx0NghYlwXk31smsx20zY0Bz+AQdMnUNc9o9m/Jx4sk
O5lIZBFTgPCssGFR1SkSzZ/KEPdir6byY2xWCNefDSuCFe7VoLc1/2p5x4W4CU3d+Rkq33n8ftOO
t3EqTkqKUSTpH3OEB6oL802cnKvkHZ8ubjC+ToSCLQdraU3Fz2qQuuSnqxgMtiyH4SVcJ4ZT+4uT
H4yh6jCZkPV2UGP7tEq2BllC2RNl4QVyfulQ6VE+ZrxbZ2rgmbxQCZNIuoA3exiS1Xlxh8CDRXrl
HIUszlpVauyq9E/Nn4ViG3O2g94AY2mCGgRtX8s662pCKqdcQTouBANcGN3ibWxN2d8qXc7Yei6m
KHTNJo9ez7DHsIMVeeYC0YkvoY+etYt5fimHFvlNqE1Ru/u7+w2GDE2SthNgzMLvvSLFBgzgQ98r
XJ83EReMiOYw8Z3GfoYm2KQqa0D657TsUtz9wUHErOsBmCe6/sXZk+nZS4TCQFWKZJaVvHTTxqi8
TZPaAUEedWPB38y63tHNBIM+MCfywnrZDI9x+0Bqu9aw2W5/v6fGKy8HrDmXRAhR53E7X8g6Hnjy
pZWtcdff/7uGHLD3YfRhnyE+RdF3IfsrkLIwCn7uy5NYeAYVo4VbPgCr7ydpDbXt9Q96aSXi+938
niciB+mcobOIX3uUZNBx0G3cRYoPk29h3jwTeKIg2NSZrXZaFek/szq5IzMNkYpcMDHXFceOJ5ou
YEeRFZ8GgaFnYDu+RY7Ro6Ijy4arCdcJJn3Ryksbhhc7TCPsz3wq42YDYbEpRc7IV/qOcqGQLszZ
EyGzZl4xYCArKQGcweZi3uoJyieREVXADaeFeiVlS6BHgom3PvQtODMAKIHIsKVymKpmZPoNkhD+
BuFfXXrcyQGO/iSnl8vrjmCiiQcndQ2gCd9cP/p52DMXFfWWQuhVdYrmI6fKqqotObFXH+J+TWFP
02QWyfYXcvGpP+4zQX38YeIxexxb+2p/mvb6V969qGyMBOLUIsKkmdag0oRPw3ko/8O8O0uf6jTy
OQrcuY7qk6S1W2XwOlyo+HQcUlNiV9eoNVjPA4lUzQDGpFCVqcUbCU4L5eJA+8WXpZIFbsxdbDx0
TubWsJYgzd37bRLC/Nri+o4+/JMxrTJsW6V/zGzF3hEYZWw64Hou5ZTZg2VSNJmWxZNJWcC0Dc57
5WuxPDmEEJDAZi3mu8WEGhWZgUinNHWnei8ypghD1+tzIQCT9gA6+kauXzX/FWD3uQVxFsf0HP6Y
/kLzUa80L07i1YLazmPjCVzXzbiHseFubKQ8DvRgxVM0wmiSQSLFc9CasXFHYYprHn2xaMaLCfF6
UeVUfXAQEE25dumk5nB29crHdkCeVwnkvlLtwb3jHFfJsgPTZe0vss6J95iCeRlkiCafQRLYUn91
KQoTNYxpK8+APq7N9e/4VYWUWRjhjdf/4Y0yZBsxBo0DT4JdI1DtffsrgNtRt8f3ejfe1opp4aup
7JjCrQXWoI9/OMHYOKDgwZt9xGSmktzJQkfHnpxEmGetv5EkFw15zmTVh9slSCgoVvopwSJ06Z38
B0cOHArdomNKNlCgssP8JAltG2YIImnyYpqrS5yw3PtsypPT5DOoswJyRmyW/LCbagdhzDkS+9Dv
s15co3cg961/v3V6MgiL7j2pR2VefEfZLBnmrqkyeL0u1pzXO62/S5WwTLGjz2Qu8AgEUnHHIyK8
/v2hpYrPED7kEkykR3h7iVX02/DcdQoASxE9mWzT9jls+DwfgBoPk9bXmM1PgUH1dOvFsI2mRayl
n5G93llzr27IN4QA3Ma6N7X6LxpuyI3CH75km2zUN7MgxyKbQlgaUAEjxyNZ77Z8Oi0yrBta8KBZ
pc8UYrjv6gqQFZA74zbXbSJ9DYU5/Xc3sR9a0ReqUv8CBLJ6j6D5u04vk9K8EZWIOLEoAlL1oLph
J8Fdy+nG+pqp28J6TnYqpoknaCdtX8IrchX9bXJ+v/X0awfME3drtJRCZQb+mhN6gj9LK2RMuMIU
3b8fHZUlIx6ivxGsyDZYoUUmSVwtr+fsgLTOmzPbPbsqXspIpIXwYrOJNrCeOHBRDzJGLAhpwoRN
ze/WdyqwLUqZ8bV8cishPMEQs3XrPZbAkKVI1NO2bOw9G1rPCvV/WtVDyYYtzXKllQyx/0zrx/k3
d6xZyslteD3T49JbdwJzBzIZsR2ThW72kfr4YlOEZJQ6SJlclt9nCt3YJ236eLJne+DB/B+D/Cda
62sduxkAT1AQd2UP5Ho/omGtOB+C5wEgTPcSV9uzU6gDPBJb+xBzgAJ6mApdn9bdB0xLjIHygZnW
0RjawcD2pSF2yr28e+eM3BcFw9AGthBqXt4nm5Ew8q1rXXHXrVadQC9WTDpp+d+bbn3kXyA68Thf
TPqHdLnucAfXAzSCBuaLjemuFI0g2kgkzU71imXKudS19Qcajxc04FJllt7658C0Z5mYTxG/GvKB
Go6L1ryq9tk02av3AC9gTLeBIQSxxBJZzvbLenoBPeb5llG8KiLDQiwyAnIwfu/GuPcAAG4gIc4+
GFKgfN/qMk9IzOoX8AizN5/h/eRkHDU9tL4DVqQbUMWdueSN1teX+wmDtmWIt3Xs0MQQCbKwbPVP
m2Ze/F/EKeQqTSIuaVvmkdNJFWrZzl8d3hE0eEC+d4N9t5TiwLt6Q+XOAedbN7f41r12I5y9ByrO
5m9GM4oXEogEo8gk+YbJOPWIFHGERGOzB047nhcgMM5XtbA/x5qEXpNCd8t5H4Dze+5HWEx3ORh1
k+S0y4TINUumtguUnFPq2yffoulZOEJdUO7YhfEBUZt4R6jdF+JD2IkVNKDLoP5rmuDz775QUuDc
W1rcOZmhogodDUJ4Qqz79unUhkLPoAc24Ho3RU0A/bpCAVXHXOzNLoFJlrUINPD6T5l0sc1dobyp
OuKa/D+4hutzqnp8+CW31D7ycaEbtfQhjbfAIWVTXrSZFc5AW0W7pwDUxzcbsY5SSvd6bJ3F1p66
s0/Zwr/MSxKgcIsvvzFMeTIYd54+YcUG3PqWpnoiwUdZ9ioCRyamGpduqrw+v7eQe9Dajp3imAkv
n97OexdjxMl16RFTNY7g4QW0vvLcajRde4PpU0CciUHfUwTugEW6vhTFl1n5d28As0FYFJyEBIdX
US73g/NCKYmArTVBK+wA0Yeg/xpqr8wnGxPRo6enUUPYyHTwnd+xnL/wxGJzTzzgIYVcz0iA4gaI
a52MOEtC7Z5Ve1a6Qps+GOLYesAeVxDKqhptTvOn8tqOfTboKaZhqzX8AqqAF7YO1vDHG459IOXT
yD0BlIL36se49v6QBqhhkhNElGn1F3mYlNhS1MfcixSN7yUQVi8Y0uejao/Mync2HNkkgVvNz1Sa
Kan57smA0CMC+PFjmN/tJCCBeuZ3pKW7AIWlNt0qvJTBvgp12UfdGL1krVDlKY45cS4Nok23u05C
1vFCwZ18Ksr1jMa+5u5miR9giDO0ZOtNh63ZU4ANzNE8iWbVlphOoBex2feqMnlkJGJ3ylRXw1ov
q6FJi3f48lCpxMSTUXAZvD7vHwysY+X1nEUy2qqIXnLUHexW8hXrHBnuXC6uvepAg8Ycft0qTJtY
6fTQwMPnblRjI6F63IBaQcoBAAjL1FX7UsnZUEujWvCve7ha4s/e0bl8w2EsWfF8/c5j2Mnzu7v7
5jqIjuvmbcdpiz6uZjCiczZcIGv+119G9J2Ph6TlYNimf+hhJJn6CLZQjbr5By5Gfi1TdF8FwrDP
7bM3kIqiFsyBoSOtqCy4CsJBiqOyLcSzXCbuA8CBiyed3Gj6Dnsiy1o/Ok2leVBHXfMsVJZZo++4
MTyU7RM1irLBfWsP1v2YnGbQxPxx7oit35Y7UmqsNNN4rpavH83dGnR7MP2cU0BuWzCz3jTsK1qs
/rSJIyzULsar5Ld2ImF80a/cJER6H+lE89F5iyp5iwfnRBCZZ+2lWSL2ZleCs0+giA6U7Sfw6Ib3
4rOhH7vX3sjZW/N6uiXt33ntcxAreYc2OvvvJLW//JGP0wUKPPzWKFJjxEooBKtQJOiTrAksnO2e
Awu6LPBILd70Ru0QFBqtUM67Bj0LjdBcCL9+5334jWT4pqbrXIKhcq7PhnyHl9cL2cQ9vMGa2/n3
RI1QygvwiHnFo/htkxgYxVkG2uBqKd4f1z+2tcb9KcIWSbW5KrHtWeoav7iDAHDs3z43sIbuY3XZ
lgBVmxk5c3RgIqp7wAlU0Efzlw0JRM2O+oFVg5pfuG5jB4jvOmlssSzclyu9tlmj+5IMrGBiPmyF
Bz6O6tC1gy+Wf8Tdx9Ir2yhbTgWQdsmXHlvECeZC0HdrzZbsudHQP55HYxC7DgZFU9nugy5wARc7
wYlDfDIJSDn+52ypd6g3OSaFzWqjZd1WnW7K+t4WyYDYQgKCnLHh+X/FmP+p6IHDrKvqcve+Uvb7
bg7oTu2fmE9+/VIHyitVZAxk37rNzh3ROvzEpV/u79cmFQUdfEdHZ/3Ca2eqTtouVjat+jdAk7NJ
vOPbI9uVe8fjYwPC6K+kJlaaOcJ9MQg1ezdYOcHZ51TYfMExyEGomAlV8EdPVYohlpuHJlqObGud
CqGbzkXxGGaHWhFMRNe7EBpntC8LWNWIt58jZpFs6NlezvxDu1wZG7P1oKSNTdTgSzoLlNQ+olgm
NTxnsjipG/RbEXVwQLAJwNnD4OSpwhh1L7WSOLm4zFIyHMLeQlKJwZcBA04Uibd+TuWg65j3mGCJ
SGKeQGdGdKaIYeJ1klFqShLvo3wuckW+hovNR6nhcw5psuLB3ki0mWejfxse6IIqkvZbY7LGI9ob
qktUVKUHDsaozu1/U+U0e8KH51u7euMyGj+4yKo8PMl5HgMnq3FcY5f356AFJX3ZJcVY6EJHz8ip
udIwa26tG8YUX+oaBUgE4rId8UFBb0IvDqM/sqkKubKw0/m/rBOu+FWecbBVl/uPyzPMDD+36P8w
pyka0fl/iOKVlW3pTqpWe7BGVqzn3XgIi/sGSKD816QZPB4jcvZ1//GbLcfqDgdnkW1uy8QNGnw1
6KKuMiRWuU2SPYos/hiEMnq9FB0aWoVnsoJ/5IMG7BZOkpbE8f7xOH30Q5C6Is9A/gkEQC+kJg6H
+f98dPAWvGx/q4BKU+AXB7hLRlpUPvvivXQYe0lAaVyGh6LoCJWm7ESdvE7m9Iy7jwhoRH3auqVP
fYqD7KHATPASAoo+G+4urAErhywGmaYzZudMfgN9Gb0t4omRU7xFywHwDzM2gnDQsCocVny6jjQ8
LVyFMvaHYr2kfApR8x84nP/Bf2o5trc+WxyFiyGI3U0m2/fEUkp2aFfY0nUNBAa2e1vLrfn+ydFd
U0FS+r8trUAsQrQ3kzUAQtPX+89M0CTcQx0UDTgRM+d/uRe5OXWdfTjS01dNba0LyJB4ZvF+sk/d
1Zx2A/aw0Ghu1aNQUvypnOi65LbwoxlSdSHS12E1oxVcKQDgTIN6XmSjRxL8h1gV1wGHPmVQTVOX
pUZPiRBnOEJ2UcRWVV/3CFnBYTFE4dVy6m/mOASB/YfhZyabAMAQVLScyv9SrUDZR4G4s0mtouHw
3TbD8jaKTjfxCRerEC1gLxBw5UyRleD3zV+hLwEwiWQFYbIDC+MKj0p9AZLJSB4BEhVTJfBleGNg
5ovkSPYgjNCuguZAiBMx0KXR5xkyovz2ARr4LiHfidZJZqqpsJ92A15Ic4jJl7jFC/P8WDS1JZsU
u4OIBbH84zMshD2AELlAXMHJXXM1iaQH4YjOCWZ8qvIg/Ujvy3EZFZIKHawQs0HXVSOXJTthlVBc
Ul/x/SOAg3q1lfhsTKAhCV997Js4nI/HgK3bpknHziCBj5oKifbGautxVQL28AV2piJYBjcCG4f+
+X7tzave4hWiyI5i+nN3R+09ZcXP1DI7Vh7U/SHvxskzp/j7gfpi1Ms7x5hrQo59Bnm0V5GmpmhU
6ERAvX6WRF/+1rrSfB+55uCk1F+PmDvChDdzXIf581WOYjBNSfqTWxDS7XsaMKVuLavRLd3o/cEh
9vLj5cSLy/TbMS47QVzhTyVPdKSANUuCMtjNsBW+g+2iAhYM/harq6jqiTQ+XnlbbUB4JLk34AUi
8QNL5QWGtlryhyWPhFIgLEQJJJuWFl5C7CnWRWGmMLqaAt5uRXDkce3eJi9DjRIBjodAY3entkCl
OoPwfZNC+NcvvX6KjcxWB2XSP6ljWuoR6JJ3iIpc02Vf63wLr0XvLjqRUwrVJP2tbTlEGieJ1BzA
DZO4bsDV28GxvfV/h06DguxKYHbfBvTm6rq4+LvfUPq12KItpQqI707MW9fNNIPI7soQvH8BhKEI
3iF+ukJw50M/8ymD7sTPhyS7NRNuo5iEkVFKL5JZEDMharKNtIdUQNTwbuP17CKD2tDKWo+1uoJd
FpNengKVcKWM3XMc4jN1CuAbTMcgRa7vXX9lzOj0Vc/R0Vf4uZArX3gUmmURMNYYnhbS7Lz5t8K9
DVfkH4cnRF49bvOgAqWdLWorbUrRDSZNXhoUBfPvjPAiE17wvmykIbF2yCS790s1OcVyPxSTIe1g
m1a4FLEBrR0n7kj6gs3zlDBC/oXAmw/7O/aXrp4FE8g+6+B7yE9xDJOPpTu5kmzH56lu0Hdn3ACI
qX9DIKogiuohIPoHmaXFo5eJKnX0Ba15uUwBs8zhuHx3+Zdwfb0CYmwefN0EjMPa1D4EVOt/5A/4
7VNHWyaA+EH/S1m1UipWm8ZJp7qzoH7xNIKhRkssnIjsmqjbojGWbA2L4dJ6dSmiUHHFFhvQRCWk
HxsyxykLp1sohNzyBswxf8mZxyDgePS26OXADHtnQlBuTMzKuMUqHmcR8BHmUpSa+4L1uYWIRGse
erWuSOPDiVD5Mi8W5BvRgQzsf5l1xQH78fj1f77il0m6OfZz8tv3inB+qL2SHZvjfnJWe9/Ubzfv
5GnoRzAgubLBBCotso9kC5cMFEbpIz0c9zbIbzLMce1qnJHDgKiQKz357EOlETIldnM00J6rIGcr
JWmLbhK59+LYHHZvIqU66HnStLLk8PnrDke0s3Z0frNnaHcs37dEI/DQW4lFoTtFZSTkyzSryRNx
oICTZcSXvwHKUMNfk7muquc44CAldSN9l4sf2Dp+XvsBsQdDnZUXaj57jk93dF05+3XrFK1CM+7g
Cw4PfhmrTXU5oqdDzACichGqlJk727sNh5SlPs6wW0QVd7ej0mvWxS/41WhT/ogVE27HM/2au+cC
PZ/v9k//Hjb1+mTDCQKkPstN6eVPy2csxRivbyti8+65f6SnzNvZV6129Cg3cyDEMldHSCrqi1U8
RJbQ+cRWU0hGtS+7FC2pTi+hvpWt0ZbBjhZI1J/ffu09zBF+OJT9WWlZyh9QRqQ8KEO1pAwjS+Jl
LhrUhXkURiZ1uqr2k590chkjbOAo1CcKyv4LRU47MU5lejXJEt7iRcP8fyloNFjbBQbsH2S4IirB
K2sa69qSreWEHL+F1PPLy9y9R1Aa9w4nCG4Le5eQFpselTolp+iVpsARa4od/l8nDjdqYiFrrW1o
56LEB3163sQ5HrA3P0cEWXtG3CirRbKptSsnyLteNMzuoyUN/HLsBdWHD0GDFVyQESSoazuzRTWG
DyDcMp+bDkgSVGvoqwxCQgP16x1shjyyZiaa9LLspi1G2SwQbo59fYklNxyH7cwRmybKbVV2eBwx
q8LU+i/LqkVD7OCXAK1ZvRCRSnVU55FS/cTk+aEfO+UCfPctOuo55ab8xUbEod9rTU0jKclOcHtb
wl5E2WpnH1ofZHGJTwadhGA18iqSNSPhrcFc2oZCxkQ5AAb6bkuL+xMZpTHhKgS3WT+VpIYqpF/N
SCv4fxRuf5F2Q25PBtPBnvEQkAmfmi8Ph9Li6lojRsk4tE9BlfDT0zmSOmUm8Wff78qFOPY6s3r3
D124WYsf/0VuvKm2TuatrWK7eEYhjrnJqvpKgYY+y2PrTpSEBpRjrWJpuRlomCbFpDtSnRfyuGw5
x/mveqDnLzSoafY1c+4TwY8wsGOBskcUgA/9+zUGuL3oPQi/xuGYE04ZoQcnndoMjXw5piICaOrs
S/62EKsh2jswXyTOg2+h3j2iFls0T7MoFRoTLBmG76K6mmGudP1ZizDXqtOdZzfpH/p2e1pRyIaW
4nqKA1CQxL2n+bf+5jroJQNIhA7SHflhY+RMHkFG1tJ7cqJYFxWwKp2uLCfR1RdZRsbr+8hgJ602
4n9bDlOBjDciz04SDvLp2OCeCqH6Ew4pna5nBhWaemQcfyncKWgVnvqHctN1WqBBhAxtvCa4Bi4z
zDeq+hnjvFY6lrSS01AaVYQWISBUsKKk/QbLzGjYWa+ppjeBMlGt1LrzGAfT+fxN0suorS4v/eDh
VFtRFSWOENOM3gkcgTx8wDXD48zp468F4yT64kQznSoOmsixSa613qcl4Y2cIWM9G69uoLfT5NhZ
jNI+RSOTliNWMOmrUkkx2r3NsxFArx6t+v3yTXdaaPNYJ3TJXoTD857Cll23LG2iArq44NWqd6zx
YgVX8socr5py4qMsbSi1iS6MwboGPkSYh7dlrxE9I/BkcBr9rZw1qoBqDau37DHvrcNNMQhjdadQ
fB5WzUPp/Tk1YfwExoh4LjyVDFuqgpYRkoSXE1ZvB1P6fHISIl13cHriCtVSx2YFkHHXUBFpg6Y0
t2rP7nynxSburhP7fJh/8aNpXX1jNcoHGbyLGDC8AM5aq/IKXK5eWKODrfHonNxa+wpv1B4IqMCa
OWTLNQQ/9ftsc2Mv8Po6nJjQfTitq1DmGHbpzOVjPjN2QBsYSJjTUv1b5vVsy2aFa2EW0cxueh+1
m8l8vBcdjEtMFJ+Oh3n2gjKGKB0hklOt0BnMHHCxRCWj+ZhDrKfmWKUhWvGYRL72pW4AB1N+asJg
tu7W8UUzCDA8DnLFEQbXjjocHdcUm8MA0794Dc/5iuMoTGUSFANpLixsoZxGVo284nKArpxxP+tU
mUz5KBBQZDbpD7nOkU6c8Q9pO+cldPJBfVRPxjJTXPk/CAlB/Xrazf3VJj1Kz3U5n3gavsM5ATxY
6LD0SH/fRGwnjRDo8MtvjtbL5knBR2ck8d+PSbAsWNvu2cMTFw1DAX1ugXb9OnBu4liAh/XCkYn9
kcljKNJjb1OOB8wxfxlJuaNy/htxTFYx8eP15lN4SnjKehk3d5F5EF/n1KBV3VbYkOEe7dkE2Zgh
JLizBpuQdBFcgnVEEoE7g7HHVzrO79lVhxk4/YUNtRtr+QCd2VgkNcVMJC/j1DJg1SBisDY2aiTl
2VMEVfKfPLUgNrtTPGfQWsB1Kv/dqsPMOSFzUVymACfqH219Us0uF//6Y8moxBzRBWG/i4LYyrIL
dAP/YksWF8NpbnR8BGN1s/fA+gV+eRyImW5SCTffPkAX9Z8oxjMwq5JXi4UsSKU0PKmpKHxEX5y9
VBA0ZbyJj+eY4CGX87R5RyGZsoDGW5VmNBuAEmMpLbv+YBfsxzphR/uk05w2DA4WYZlrikDTvEOj
wHzLt/v+k49uaWsyAlyVilBO4eHqErfQ01g5EGHhfYQylWs+BbM/3d73DVGspAdGqGVRiQTFQSgW
ZvjEPMDuTkdIms/rKZfD5taRU0leDSd6QWzMDCx0Vc/mcMi5MBV1suM4dmiqmnETvHfFrH8uBocY
elOqk8RzYwnhg6cqgUKCojBsj8jUMPE/mdldafnEACbqgnTMqE+NLUg0m3NXzRxbYIykS5WOds+p
de68baOWyq7mTFcZscDDeKg+Qp4RQKZjlSs4xl5U09B/a+CCqGpvZvlwgWgTKCo6UrAapgS+35W5
u1ATXypu4nP/ZgDoMznhcE2AePgbuUgGnStHjvi9DfksW19mVT3ma5V3YLSudQC6f/pRQYhLDhwa
zYCLcp5+C5GU/S2kYCakU5/yYpjGyx9OK+52fNLERDoIYK0U5R8ys9/UQcs3vRLR+mKJ1UrC78GR
noV8Jaxlbhr3fRKyDTjzwWE70Nm5Cs5eH74mRzlLJsmazAtoF4LPzs5K6ZzAUOVKoMlIZPU4ylrR
1X4562o8wYwxfkwkOGjhwo02l19gqGvxLzUvBoPws69uex2cVx0bjFbDUPxHp0PrjtKyDth/3bqh
5Bh4ZZye3tMdVlZBVk3akKtLvpydcXDPJeMzuXkodX8bS/zCMOUquJpqPHxYsVM2mGIFR6Exdz1M
M78FQ31XWfB4Nytl06Vy7qQJs0+l7NDts2b+lNRhJ7unP40RyinAe07qa57QY8vFoeR1aMtXWmnP
jszjA7lI9KL4+0U/rAiSSMIpXWDFGxW82z8i3TG3k536N9pNVJh26lNyjBg/RPTH8KJF8LuxT1RO
qC38nH7bSn3bQ9B/NQMJR2yUOdtQApPiiM+FVLTkMxZy7OY3/IpskFd8jVxaL6fkE4L1ppD+LPha
0/hYaSaUa9p6CxKjxkTxIrTMuKhY9+UrgwRN3d1I9E3jXu48jpkJJYm+v6/vMsqXuUaFUoPq9C0b
JmKBMDtyB87tU2L91tmcIyd0XATceygEbqgBHzxkgrq9/JKwstZ7RwhwD/sUb5rp0HNmNtPYvq91
KUSWP9ieJEVTAUDtffVY+EBq/sXMuVbD55NmMjjUszZZ+XAAevwrnmE4dLqZ3iYWjlB4zJEHBk6Q
2vviLk2pQ3tYrTt2n2q4LapJBVT+XdsH1mY3Lh2y6OmSHGZ86BFN/fsLSKDKqaZ/RSKSOcFrOEQn
5biVItkbXMtXcmlI/NG5hYmWfR+D4gMkf0oZishg/M8JYxcfINdgq8o1iG16NF+aV8NXfmf6dmXX
esaUwK+WZ/PaZNnbNYtUQ82TB02XTGZ6HJ40foTPhjbXpuj6JV9upCndCJTDsrxj4UF7YQ263Xn/
n9a5TPC4HMV68/W7yt8jsZm3EIHC9WpqqjatuIcfIR38h10kh08GDZpYuT4Cju/EEOqUaH3L8Ujp
h/ndMlnLekEs1tjnq11vVinQ+dEFpzpboC06BtCJ6P0UfMcx+QvhAzhBurLx8Zbd+b6beOx7irhN
dveXNmBdUbGt8PHD+VXaxJOkquZyb5zgHAt5Qo9BxgDlnqANxr/Ghc9kM6MMj1ZjrxVzXsI8TclO
KPQ3HY6LS5D8BhELpkIX1NjS1O+thz23oJn8XXG6b+GO1pSTx8u3dN7ognde4fu4pFJ3bR6zkY3D
C2ScaAFkrxVbHXCVDVZwANsXRGTay2rInJgNan3jxNENKBqRPtLFcZc9Gn/EfmRnHt4xa9asHc7h
XJrTk3cUjMYoUEm89W5hK/2IUZFPCzWR687apd/K3Bi4QdGjZ34/Bendm+DR0u8bS+/rf6ULebpp
GJiqwyDLIXbD4ecYkwElTU2u1HDUI4q64mW8VPQFtQQ59J6BxsIuIivzXrVKqvoCJvwLQTa8sg1N
Uvx9s8qU6JXgSDyBklCl0dd03tYIB9iiE5AMrVvuM4gzVdCTVWK7YfX1TSTLEu2a2iAibBbxxDhM
1sgeQM4TYQuaiYw7+52bvtGKRHrnxMHYVP/7XxfBNSWgWSJshDy0i93GgCjXkdGxuE5sbPl1XM+O
k6ATtlfMHoOHlbF6la+5BLW5q3BSuXk8Iac+QScHNDAPDfbDVCOC/dYtMocEsUQq2sDFb3m3Itqx
gn4WYTjW6spWj/EkgPG+TYvvu2IFfPmj44xGH3PUmt2ruLIeq/JbSk7MSvkGr0+VJUn3HLRNdiIv
FCuKqhHG2BR/WdnJlV3iynofiefTNNbx9wwWOIQsHw7Vdjctd6PELZTpRJpVxRlbd68yVt7IQ7A0
astFjVynjbIWo0Y2uPJk3oLwaxc3u2P1OyOfAOiq6lWQYOFNBbuhMEtQC0mOuR23h/MtmBtpoo9D
rvtQr3Ii6ooJQPtmy3YXkvHyXjwcRzsi/PY8FdJ0hgxft/oSdOMfmG4JTFAi9Z0XXJexrnzfcRQK
xAHiSwjqdAX2a9yPFml9x91TmRpgyJOs9WsK3hVwQk7OTLW47Qo69S2E7VML0CRrCXulpXhuDwkz
ZZOSUskOTuNw8o28Ydl/HQvyLftT/ANlGm2D02BOo6XeU/S1WqB45jP0Pymu5CSTXkSwCgQYjGQT
Zfvy+q8sxS+Guif4Ylvsbfr3SqNgy9naXP0Smw+eMg85HN6vyb+CQmwoCk1s2ENPjhU6w6zYOPLh
clowuhlpbwdYtYr4fdr0MwUTSn7Z21JZcWZHen/vjjR1K3ZBYzw40hr3k3I6B/KsmsWbZZEzxvjQ
3phMbXoSNPHIM+GQ4qham5DIkdtR4zFlhE4q3GdmeIdkFiBcVrAE6ryTzr3nSzF5wqvjq8ZxwLuY
4OvPKcmCpts+1avA0mHPrBayG023D+DgWk9Kyfyo9EBzMalzpyLhb1ogzQoxmpXk9ssdzZRD1gFu
pKQe+oR3VmaDegD0lkPnkTcmoUcZLQEQlJ6OmJBeAXSUxwjPnhp1gjgSAH3pi1geTuAQMUjnDmYQ
zJqmyn/QHgf+TWrCsWPug69O06iMc79SsGcLO/UOGoGEpXs7bsILpSazqevZ6NFz3vBh8JbcSIaI
J4vhp9LGiR4TpuaiyCoI5CumAOD2+2qbxrsPRcfdpNJIv7CWBAOOOgUHJ8dtHb2togKtvoHrtzLM
QhUqgHB869vdYHEyA4mM/APGgPv79jeqhJ3+LApN/vUhZrmg4Pf8Gwdz1UQLArJHKoKA7My1hels
qUUnvq6OxDAkTfh9VyJWEg6OlLxL0HWVT+O67wXSfJq0tczAMvYPCbypjgaceOYNtQQAi9VNF062
q97DPMj9d3msxFwjaH77WjEScrGw+Iwp1SOhB0WocJAj574MhthAutezSiWEg/KNjS3OAi01IgkR
eQozhTZ1lfRYGOP3XfZjjCWAQS1e1kUELKaLzg+mgzmFF7i9y8Njgm3keYbQFCEJLRIu1JNZ4jBQ
1z+SDNRNwZpJcd9kbh70IelOsHmXzm3ZDmyYLxMa/sJP2xcbJ03c/ckGatGBUWUsRqLWOoNaXPwA
VTmj+/3o7UgsvbqcsmxmPNgZRh/j3Z9m4CzpkKlTlU+kB4+U4UhRgMaUa2bNrKXLv0rAa9ZoX+HB
M8AVTXJc0SPhS1pgJRDMUdqcqhXnrppLAoAIBij1bHkA7hyOJpcUP5cTt2z7cflD4wXpRpkhrdUv
AdEoBKJG9qa94pyScLhsSTjdF7AwRidSoVX540Xdg+IHEnCmxyZ/uBHAP3XvSjwCYkrKJ6NoCLFw
4qC4tNKwMscBBbptpGKckqx+cVzNdalPM6TKAtNSouNmtj0Y2BGiD6u2U46QwgEGcGnTlFjavK/H
Xyz6T1M4xi3H2HdiYxuVKXPR9P2WH48C9kGZAlm6rc8ecOVVJwBr02PowW0lEg+6v3JUF5UySpyu
I9i98V8s8gCvxirqOSo7uiex777nQxJmalIT8nt7hfCGyrpcp6X8gMEJRp9mDAFfOAfKrmhXGVUU
fCiO1iIpLo/FnJ7I27joY76ZzW/E6uP7dLU6tTMO8lDUtjZRcDr9J7+JnMuzwErJFI1x+IXFuAxO
GQjJN+SdwmcHSKqjztgwEJqWvIU4B5xkPPMn7HhQonNzzMmsGo70aoFZXRSqDYlvPFbWYZ2yXBFa
CB3N69KoCWIsmbhD2nWKtjLUOZkJAW+ujbvqAuYNHdmkeehS5eXPRNE55u2O4Tl/wiyYFQv50ZJy
uvK1Fj5Zei70EMSysCFyo1h8iYDf5kAchEet2DBb/3ak9TUzIe+FX43GXOVYNpt1t3W0DV7edo8A
ctZgKw36jD+rjqA+QjbAfUM1Htx7BH+8TKwEDCnKXIh3gL6axJdO82z7G6uhgDg5XLXPaulnUk0q
ir2AERG81vbe+BVDV95p+qf8HhkL9VyAdSq528XeiNsdiBrFA3WoZAW3QiKDz9poYRo1aLKozg1+
adk/44YMdyMK0cGe/CSEO83u0PeOSZCWmVcdfftjv7LWFS8ZFxsLvrqA+/KBnuNGgnluQQOKUF8Z
jFkfbsSeccQvnlmcmMkTNJUYRUt0VlJYDNSeC/RJn3DLeg9toRi+FKvp1UMnAAaKbZHLcTcx7xaL
Wffn70Cmnag6LQNvuJ94ipliPvieW34wPnSvuRi0HouHlljdLdLdCkSThcJSL3j/2sADjVB1ujtn
27AHAELCJQE8IrD87U7p1XAz5lUyGIc38g9zTmLTtM8mLYJt3WcTSFWcN6fZ2+A8aCxMSr513fRr
qqRkhAk2SvPFP+BYcY4bOT2yXzc+9GILD6s68Vlzlfm3rs2qIQNh7+9dDkZB0BiZNmXzzGFnPl6b
rNKH7TOaj07vRIfZfaZG2UiL5SMfBO3seJD9RA0vhhHo8JrU01t1CpTBMyQ6bgLVVKRBs86sGCa0
NFFZhyPG1mDKbdhnuCgwB4axl9+wtSWeXWilPdxK7HExbqljJD8HoJvi1Ypwlr4qEmNDDaxKLO3I
sOkgwh/Cl/TjxnRntWlrtLtrsoSfQAsSTTVWWtn/J9niW5s7Uay2s0lJNALMBo5FJlKV/z/JWGZt
1pobv8IOz70oCBUZUbBwpCQzRbJ4j/1aXbO9mn4lbbLmOH6tc6RwXwpAeJt+l+oGuy99ZLSVRHEM
nx/SpsThALOtp/CxDtGIKxf2OoTNZKdnVMUaq/qiVqIvFIeKHbXZTA3/DMiObE3uSg2VW/dnE8TK
7Xae3ukJ71bf1xK6viZicTLZ2MnIEwTc0UW3dHTdHYKlVuoYIMdhBwHssqlsSE7KfEMoKo8QSi48
qe1zNCC8sFisWCE4PHNwIVM7gfSK71DH0oEJzQiQfHHhbKHnI3Q52NSPqhDHzVt/pv6isVOfNhJs
ohaE0BzUddzGXFk5mIcdbfBnKVNW/DLUQ825i0gMZGLFQdsn/PpmxccwiCTvGofgE61shsPIPFOr
dXwEIkzUb/yH+q+UFMaEW5YHj7PrPF0rtGGeC2JKKA9d7EceALo8nddq5XsVSvnAbzwQdu/TGNwK
hXPs6jXbK9lLjgAXQ6wEhCnQUTliMUWJCGmFT8K0A0eCKUMj1xmwjhrbE7EarbCo4NFeVBlNysir
I+mEQKLw1pwAnh5VUUu8cCY+OmIkDPzspICkM7e7ICiOo2mNigeoVedbOLcTiULRplQ/Kj5NR7ot
+FG8G5WWWzg7YHxCjaw/BAGC/q14+JOHgbruF+tr15Dz4AV8Cb5w6KcUSVMJmM/F7adc37tJCf5x
R+XQKBRk7mTr7sx74dj3YSAElfnxMjakRbT20E5gIU8Fh+oEdNxO4nMvCd/ONXJw9vqUUG/2jmIe
Dr8pdCYpaI+y7Ffx+SbWJPd38cNgnFhbO+2gVTztk3nm8Y1ZrmI6gShK/bkhKQ3ecwxaBjzwux2A
EF0fJ9DJD4ecawOwUkz+QKSEamaonY7cItC1TOzHV0Ji4iHI+XylS1WLxAtdZ3esAefTQCGICzZ1
BYYIGuINiqZyqWOWj58ZQCalgZxIzMsFkjRderzCK6XwN1f2zTtQ/evHgB62tCOkAekGp3AbQczE
aAMxRPAhZkUQgzimbgHYYaI+x7KCd5aD9wUHBkGjN/tZb9A6Zl8ubq9A9JKNlLRpe0uV3lfGkHZI
VzMi8Qj+C4a4Vopk592Zw5zZk2Fbg6pI3vx0xbFdgQiwsotBbeH9SlioGEdRYQKbm7VhcounGOxo
Awo/UPw6Z3OSgXvQ06e07xrsZsN4+hNj+9K2DuqUpnzOHuj0fLtkCSqyXLoOYvMUGaq5i14EUYeL
A389dGFh1DfA85yE/4uOvxiWy0RZbmiUOfDUfFLPQlkgdBDo01h9sBg/QuABu+l0q6nIlx491QHT
pBTPVaANc73ZfncL7GisatW4euM287lK/UgPlp3X1WE3EvOYGCTH7c1f9p6tM/EB12fjwAcvu6j6
aA/NtRAaZzhv1y3AZQApHvYAqeuu80rNi13b68Y4vtlB65FhhPUxG1DY3jRSn4aMMtwq330AOZqX
JkxEhidmoN9BfMvX1yBQ45pps3qAs7NqkA2krxrc7szHwWML1+o5RC/7m5mwh6OFdzhR9f/l4btF
N900QHf/ZSb3Dc8sBpeOUCzYOZ2uD5a0Y7TVbH+TrRc7MdDoWHJR7l4UUaJR/Pi+xe/UXhYuJHds
XyHR2Cptpvhf/xTcd5++CF3xK2M+9WtLyh0l9YL0Uu0AKJLCt0k04O323NwspmGOVjcIkG29cogR
PYqiOfznt1DsNVySvEbwlqg/YV0K5bHfPMvkc5mnNsMeKX/wjyZQfyV41nT3WBLU0LwCnfOH3/wJ
hdGyOEMpXGESTxicxdlP+lOmpFQMTma/hAJLfe7CkbC9BkBxopYQruU8ake6IqXIOz6ZZVWrtSxp
d1oJ3iQ/rlr3uV1ezPyoMhZyIU2KGPzVcF8MWxsJZGyUfIO6L/MMOb0YosgmWS1ranjqVa/ukmxD
PWtMozA2DB2Ftkcq3Iahbi8yb3aonvbtHnjQR8sdudNFsgElIzbgfqaY6vXX5gGnfAboKwJjweU4
Et0FRBZHB2/Lt4PudvRNosZmrcbUlsnWiTQicQmBxdmpLlYl5NkFsRnbRoGfbyk7i84Ku9Qr9d7Z
z/+Ku4wjyX+OeuZK0RDkY0m0wximFkFWL1Bq+DuZrDVxH1QMI4xRE7himq0GFmZhbHRhH7FkRvLw
bcXNujAkwZMvnbHqr31ydLDccx9VUSiZH75mm8FSVnELb8HJBuLAgHpZjfOLAdzSi0vNAQuQO2k+
77WMXYpi20YONGoF9ahOe5cwGbwV1XJIyyHypyay9QMAzwk4s3beyuC86mib4HOWDvRnUB2vHBBQ
TH66ylFHlGuf4OUtv1uffOHNel8byJJ53z502QaS3ags0B1QYrrqKnk+2RsDMgAHM2f2ZWk7/3bI
2Qnu7s9WYLZ1MfrzOgogzBLgXLGFRT9vmcDE38NJxvGXNbmDTdtrwAPZ/vRKbFhYoONQHs7tZFbQ
z/KSAdOCQc8Y2iWZPPFrj059TP8y0oWI3+2foRqCK2b9IBV0A3DYR5cf2r07b8Zuk/y68aos8Tkf
Sm4fbgIRYSlCROO5JBhrNe6ABhzOkKwg6eiq0Raqa90nfk1y7nUMf2fD1QjE45gX6/7M5QCVTTKo
0ucaLNZEcT8kcPLgTxWHxSULnapcyouyaTtPo2IDMVYraY3haNO+I5P35an5Y3L1t3D5szWSp7hW
5XQOsvNwxOWs+akDpnkyvrH04bQ7DuleCU0RzYzPaNe7U/VKuhxmeeoYAU8ym1PP/koKzzA5VtjC
ZONSaum7bTc4Cv7+L3I3mPq5P1KlvDfBwAOKBzrzl/AH/JUx0TNGBgKM6IVScJXi9/r9/mrtTceM
dnbE4VJAJsuK1uVaKp+ZOB7+5VQBJjTjkGlIMRg/Nqnch74YPfNJkfo4XtVkiQC5kz8WOB6r9959
p6ZSd0N5kluokQaGXB20+E5QWUUG4Ey5Vmx+lO7PyWJ9Vuy38rv6n+ZsBDTqMapgJOS8FcNAXx+7
LyAtZRtFoWizshlI/YQDe4wp8+iWEUQNj/vuyfeXX27zP/ux25dzBzmOD5PyIED/cbvXcKzHJsOd
2tmW0b/hMwzQ0m3mNZ3EbBuV/1t5Tz0XESIAdwDnHNNedLDvNHtQqhHhlSjV/NK3xO0IOoh1TWP1
6Rrgx8Di4aFo/nUQPv0PzGo40Acq2w/j6ke25029RaT53beOXkSljZK+q9JjgxyutjsPQPFExLQU
evCxmJwAfpSJXAIrT/UycU9bWLxJLcp6+R613ERwlMKWYT9Xmnbl+uyJpn8cB5cACasPO11L5Lcb
oDMvlebl429Z/TK+3KMgXNnNcSpzLcAQb63s20bW5YxiEUMQC6zEWUGxzxNYUDA6AE6or9IgpiFD
osNXl5FS7W7eb3X9ciYd7iN9BEcFCPhNEmct2LxiyZ/406bSTyuqF7mdRqQWmJikoUzUSpUaeCzE
VBYOjFHhf5GgCemiRezKfYbr5XGvxgtl0owUBwGItiK7EUdAkXN7ACioAn4obsxbvsSz6Fq42nWa
Pa0K6gQW7QOIH501gdzZGkmuP1zNM4NqdHgDUu5Ry+065+6WSrizX2LhjqyB+aBfimD5UBJyL8iJ
gshlqyBAD8CMQ18zYjHH1DnP4rfEkTBkiySTtuLhdUKQJCWiqR3mFCQYl2/ldS7kX2iNKDPL0ig/
s8iP6mIL+/0By0GKLpWkMUbPiqQxLLshZ9jSWgC7uHcUPEVwz0u8E3lXH4GB+vxziUEIzEhzLYza
cfL9ZnEV4gVhndStOoTx6iwGHCxlCd7IzUfbMofpFAcKF3lQ/aulCIqRa6reyJ9NigdFqShj9zPd
sEAaJAevkxuQ5cHPYDwNXHmGAJ28oeMeYRpt4hqw0cxWLnMVtqX18g1blhHY2Ug+gphwFzpTqYAQ
5MViAuR9xmM+pmTen+odenmlmOxLDRN4pttDXgmeTmlXaAnTsXrUHYyq5DvnRKXTxsOSfsGXe1IC
lPO7M7iA94ez85eNPXn/HU8EPtiiize+G4hnqvNzk30Q9V1toMd644rtE+tsyh7QnUqEgRVECB0d
rizz4RQfkZLFX0Sa1vOXQoeYh/0dyR8m7uDNhaJu90WUmFhjGQz76xDdlO/1RgBDBPz1ksebbI+r
vO6KonyYhhJtIAjVvPTtw+deqfW6fdtIVwedVZbtNsV8oE+h6i62XPBcMQwHsL7IVT68YTfZ1/7l
dIMAbC5aykELkK1waiJeh9HOQrwVPrzFiDk7luszqk55x5+X/BXQq0QmeIK1sjACdabuNiVFEcVf
X0aA2UucVHZVO/8z41LiPjHB2XXNb6numLG3y7k6oraUW3gujZRkYSqedYSRFK6hXE5YaRaRB2l9
23kFpIQTYokhwjjI8/bs+6Oun1IHULWcq2kuJwy1yxdwO5Tsp807wG08p9bZWYSsajYBtWEWzid9
+TWuKkoJ1IMD63So5KbuwnTawHDpgwdIj6XcenwFVtQZ56tkFEi+cEtD0zFpz6XC0/uUdmzyzQ/K
0uYQ0kHQKK8ZiLEc9kifANT1xuyHyPnuVOePd5Z1aG2QG48qpH7n9BauK48pCU1dnpO/7z1b8PC4
juyHCqBS1ppnmdKde0lsMygMt5+iPobO2vF2pXfCgKd0VNUvGJlOS0WuLG8DbaAZlJo+TigyNCrI
jhGcixg2Nz7JLHQGuDzDiwkqK26X1cgqU9zbM3RR1ydpdKmtv7/Bqzg/0HYE79HEeyMyXTEU5s7L
5+bO51JaobScujh1y2/LYKeAoLYPzugo7tCNADOcCGtfcqrdAvThMz0arnsrDsdtDr4S61eu2BsA
zh2SpludA64MNuUqKh9lVPtJZWHWknN3CMWHMWhJhPo+oETjMWt0NuEeIOmCE/eC/6PVXcr2xGvb
809lj73I7XIk6M7u/i0NFb0RfJWe8Q6XyaGZQAoZAXZDVYpuDQNbldg3AgjktADnPVZ3YGmrBwMn
hnU2Y0P/Wg/BOp+l8CCgfxQX7eY9De0+qcJhrwYOwWl87TQIhMnczLG8HQtexr0Uoba6UrTJrNDY
FyuRYypeRxUeo5OWfrufPcB2o1gFiCzyAAgwCfqi8ls3P8heTUaP8WdA0UZBoi+jkh+Ga+7BkA2M
J0AXM+aMj/km/TRtZrCDr+Si1CPnrqN6OLuuy1BoialRHIcHk8nXGeK1c358lOr0VcwIlIjiFmoI
8aQoZzdwMCs9OA/bA9tPcjeSqyC2a2VTQERJSRXYnWPmT2eJojjRiTNIoP3/eTRRbzpFiKAVhLX/
HVscmtFheeAnMKh2DB8Js1vx8rasUv1vJ1Ec8hnSh3+Cr3wPosvsAgF0H9S+kQmGyAfcNn9x0bt0
bjb4hruFCOdcnXMVTDRejnpm68R6bpwg2CbniNhQmuPpvItRuQ/TD1RRO3HL7yV8bj3n9Ors7Czr
Q+iBhw8ffqy8JTtWRItjmL+ouYr1f4av7W6ztXPaXNnG3fMVgGmkpsitYi3Sp/1h4YoHXHJhISkd
0LjfABzCH6WTNY1xVAzf9wGJYp87j5guoHttTaWBqlJN46j0ixiiUTc6TbwgzP6bdRvgGRYiqmxt
H0Uo91phaU3QQPCZY5Q13ePIBHbmGOPK+x5Rx+zfu16P5U+nnFgoOJGzjLZ6zRwwrBhsIkY60jIn
Vdq4lC+ER5Kgdh5Sujf/0U023qLmwRRHEvdTf1WYYHb6kn7oHezZCex5Rf4nz5EXBD9IAqEoUX5D
6tqmF9mPGJEhjZzKPOTp5QWf7cplNCs8+aHRtARRiQSLvIH6co7w6tKyVxwGO+LZv18I7Q73odzz
l7x7x8IVO9NcJ+YgSI29Ip6VQ9Z1OQpjMO1uCuT2GUtBZlPWhPJNo4QbLvwiMFUi7W/NILBEGsQ5
V4jCYiNw6IgTRX6K2N6mH8rlXC+kTOd1SW4sh/MMMctQ88YxB0CrgifNqXKe+iZP0AzGJnErlv3P
CpAiGhca9dvgFGjTzcOacu3+BOuDJI66xSxFP5Fh/udJKtoly3XE+/j+PQBNcaPQ7skC0HenlBe4
+jJyHr2QNbc2nS2aTNBvlIfDMNZnxFOviiGJ7esEW6yjIBChZTTWXOX2L66XsQm7A8ZzoKJ/fMj2
18rP8MeRZS8nFuuUVCCZmsEc3k9zjshaHhEzSYQAH5yyKrRsGV0L2qaLLdMUNcFDsabvd7dMaMGR
WGG/8KGlJefbxUZWj7QWvXBIO0IzVnRaaXblvefstBmNZ1AXC/MrApMUobqLy5uRP9x+L/xBaFI2
VXuDJ/2HAV0zkCLNJo8976dfpWvnTJbnkxW8o3DFF4IcnvS47VDjc20g8m6rGqsQa0zw9HU+R6ZE
NfIDFvprYC7/VRBwy3e15eLKSPoE5FBFijsCqOmvwAajv2BmnQ4I7NPa5Cz/EUScX1pJszs7W10Y
A5uiOQKvY3LW5mxZWUdVzwyJMUhsdZHg86VwNpH00P4N7pAuifdoSK1MHrS4PtKhHNnJNPyRunrc
RnvZpUAi11vDkx3kNlL5zcT7m91eRUO/vqKWpp9hDS1MWHgZHINDqinQ6LWn1by5ymR+zoWi6JDR
7VaePJm6IZM8YhJvTI15RqfvylbErBfD01m8aAVad9MlBYPNAm2TtM0No6PFqu+FXY4DhqChVl0t
Zv1368nPocEdOXocUzE3c4Nw6ahgBS5aiZagCdEuP7H+3mcJgb0x8/py0K0pEZud4GcPx1Fgio0v
yGlDRnCTGzONQMXhXSPweHQrenyG9dwZSq5DZ+RYYeS7BbcML3ueovp9TLIK65+qEl6G5k1QL5bq
a/oimtAMjMH9NedZV1X/CEBZ5Qg/EK0j7C6Mq+m9jJHmWT5/uKx5+8BcUl1p3V6zbo9JxOKY1Z54
SGlU4ESSAzsadI3ynM0eKp4hU/rC8vO7o75tzxL2cIBWtlaQDu1x8t7X+qlLlOuwEqj6ZUiUPtw0
CNZZRCoaMv0bRhUBGG5D7HKrAgrwg9r3kYUZL6ITSLA1qLPbGHSeB9TA3Dpvbnviw4hpM0tnWrFC
BMHyPMliWQ4jCSlRsDszz2zQIOTVlPKGsbe/1h6ZvLKnY3ZC9mSc2GpHusT+/E7oTh230EpfKPSB
hvQWxTWuDyDgR0JFIItNIgLP3PU6inzv70Eg8M98BML5BQMjXooGEXKbPyM+aQAXxsORva6imkUo
Qb/7xA8mjnKJZcxDMveeDiPMBHXZUPnzvxv+m2Hybhf5cVkQ+dmCepNnditoirhj6QzlP6+9qG1W
cCublcDTEvvpSObpSBUAVjY7fi7eB8taQYi0qnuPnEQq7g3Qd4GP6YYA50aJ3u1/aRQPbxloFNXX
Oewdz0sd+dD/XhvDL3p7QEYBVFZ4FoGKW+9w2q1FJremCkRwrOM87XZREJpspXipby48R/ul6QJ+
keAP4jFTT3gq+ehMFCYvTVjdHoQaOQqQhE2rayWdK+AptqJntEqcp8VPoqi/ZvbfCwv665WyXWVI
qgGcp80zo9vIEBGJMlknJlbBgLSZJADSPKrq1jM1d9U3+56t2XT70x+0qU5kI1iiJjZ/WYAs/e5T
JUNjcvuPrJw6hsaK8urcoJI1JQMMhv28YIB+Qip1Kr0+6t9vZiqSEBArej0AiVEpDBLKOjuEFGwY
ocCHzznZ/SADCLYQsLceemIGBfi1pF08rghbY3tsrNlP0RFms8aJD+znDKogSVWd5o4dWpTETfHJ
OpX2nP2YS/89Q97fLMujgD9jmdLvavQnfSDpFOHrZ4pdwHnq2m69UQOYMBno+nLWcSABsGgJs+RD
29J7HIg1IZqY+KrCa7ZyRKiLNtVDjAHR+n2YTKseNZ3yBs6v73RlLXRMpyqUbqJYNxqmhrNrYgPI
JUkcRrykYz7ZZKBJ+rYqZj+4bayENP1R1VTmMOi7ai+FdIcJlyKVZFr4XVNTNTLasV+Tu+0eIqlI
ogU3vpFiLFmZHJvY5FavEeReLD4O+xGm0TBFMTpfQwzdNtdbOOGbpT0s8JumG/1QeSQO9MVUEd3B
gBGPiGQyLUYCp2mSNJSRZwQ/LQ68s5GZknTbnVLqax1BsuvU2pI8MqzjNILnP5wsihQBRjT8renK
RROd/CBifb6Iv3hc5Bl/bx1l0C2M4UdxJmMlgHKXT4mDc/kF+oSSaDO0H8MlKfwHPaxThztvu6Sn
cMt3YUC5BVz5Kb3oP4m0vZ1lwVkopqNUKIDkx3IgBT4TlFuPb3FXc+Gp+IIXKmYLkDbl3A9fOgan
hviW6vXC1+LfI/JteAY2kN8SeZZKLmPqYAKftNrhusOA3CzkokQDf+QCDwd+W6bbBMGsht59ORmX
Ne+ke2edbamm2pQPvReHvnvWKmbd30vW8bSs9cnEv/Y4J09I6UwST0aIMeM+GUM+16zmObAo/f1g
OLMkq3aWVZS/reoM5IcK0S8iLH7rmy83Q/tuKi5w3OYb6DSp6LY2rs38IWtTz2V8yB8md+9myabJ
ue/pwtEQfDaGqON/GdHTjVk3VtQWijnpX9/X7rpGU4IJc7aMlXQ1VYYhTj5YPLDoC531Z+Efs/6G
B7tKdRf9e8Am4GF4irNDWzzR1LBxHD9jX+Nfo3EDzBJ7PFvzVWAtKQLrmJgWCG8ue1IDtnwjY6yX
lZ/GgrJFT1n9M5BNV6bodaTZID3aba7MLZCapucjqxITByFIU9XwCDjg+MX5F4i/dBFnHVW/q7Qn
dHOZ4Wmw0w1lmsPpZOh7T3EEecGcRY0P0C4YJIpDaDwKYvEVSCSQYqdhkPTNJ2KDdJDKiAiVQ3g1
ShefBU3MdYxLLI/iUNJ1Z5uaI5/IlymAlSaCe6T/b5K2Higg1c9yVyjlCK/97rRcuAjDPRu+nuh5
TSh7c37wHziKtBn5atig8jyjbPt9jrDc2BI0l1vBBkUK6m8Q1+mHS9ipfobMJ1S+toGm/REHzfHW
tWfGfzZLZ1J2aL/spSPIvp/I6vBNouPvkvThAWqe5U/lAdjZ3S6QQ4RdiE4uYtrR9NIAhu83IE5x
StTnC47iEh5lBrGqzZl4I59wwz4VAzbfcmgVJ8XRu/T2u8KIdSlFLZ8D2UGBJ3F8FwctbkKIsaxd
EEEob/5u3vySKnPOT8V5RFZ7RaTcD1GxYs5bvUVXFAhAsSSS/BYaKGmLqp1XRypXjKqFVK0Efrqn
wSgB/+OckIe7Pjg+wVT9uBNw/cWfC1tTSDR5oPnjxynW4vas4OFpaLJIe5VFq2xrQkjRmm6XWQ++
s8bxlcmJEjD0rhRJyj48RbEdQPaM1KnSzCTVvPlkAEOBdf3blZqhcmKYGMJlGLhGQry/543OU7KS
WRQluhZuNHhO8aTqB/mx8jvz5nOkjZw0oop6bVVorimh1+2L2sMmB/CxUnLM3gPTM0SjW0GEcu8c
LCz85x4fgHvJfMd1JkvcsxbsXinkSXoO4OYHBJbzpFklPA+eC85nnIkwqwSToDc9Tw0NN7u4qzdJ
h9DkVA6i3lzpJMomBqC5HmzF0GTpmkd/geF34Jfed8Rw5zqho3DTEF9cV3LnZSGrK5DeKlokTMIM
ylpE5BPH9HsWiJ2irdRQiEkd1fMTVExjAPoXdG51072hLVnGVCu/fh90m6sINZNx3zYKSJkki9sB
j6Y2znr5XBQStVrNhbIg8fRcHz+YgAIZjjjM/5tH7h9iHUsbzaj5KBgELs7gduyDoVDNqpHo2wj3
M1Avss+ur+0gzkQDQwEvwR85X6Hm8RZT10UgxTM0+LHQIoNREZHi+9zO+Dg3ai4583nugf7i0wLf
3vRLoncCMZcOsRw0Mc7qcl7ZIIew05G1T4BZmCbrc7ZtaFhziNMxT8gh6TKJP3HshhwnJP7eDTbw
MruZaU4PPNV0PYPtH2a3/wbPXxnLTh7OHTTYke5JyO9vyWzbg3nrmOd1zg9YS4hVRYUoghklE/I8
lPLpiwFG5oXCXIGSu4/NkcUtlEOPdklNccaWeVk3A5+vQMDQVHvl+NBSVNPjpHjid75I9Zv9BlWZ
xUUQF0EDNHpfhBfeyBMidVKZUvjBWzdI4WmbNzaZ5LQgpWSu3bhVU/F3McEgCpWWySZ3C0v4V6eq
0rgZqBSW4VhdBx6gWKd8A2mDLtBrk6w3wwEuQRadi2AprcuAjm9lbUnEE6JqVPTsOhR+7r2TSshL
wp9rUtcB5QwCPz3o7PGcs5CPpD1bxD0E/iLyKE6EL19ROzVmCckiJEYCbqF+LHvLyOWffWqfoers
xt6Cf7lvUx7V8fgmuZx4hzxfRvAdoEy9cx6kaJ4JOh+YcQvyAafhtMY0FoRXSHe8w4g5Vdw95b0I
dLs/iHE1aKZ3T7EKvqzDd4uvsXSWMvmcB5JRX1HGEbHcHuhfdfrBwTOshnTLS+nFzXBZnr2crPBG
t2+7HAgbuG0uV0p/4vGq99HzqXdJazL4xM7UqiRTczz6715qBz/5X77TuIafnxjs6b3w0PytauG1
j10LBx6OJSn6yn/mq4eC4BfqFYvtlWU4c39SsPup9FmB40SPluTseuxHYH/X4OhTqHEg4wnvMHsM
1F/weQIsM+B3M44vE0fCHdx6w+3zew5jiMWTqng0LhrhAZxeavyjmknaG8WkVRwjZaxyT/t8om4y
5gDhysS+Oe5foFiPQfchfCegA9GNczheB8H6g5Z+nddvVyzhKwT2gjfoGOF9sx+6x73m7TTeiJmr
dN3LcJ/ndQxEVuGjBmTlVE+xwWw+HzqAvMtmoYwPWxXMXBM/njf8qYv01HrJ3AowmrCg88OjRiEX
zIJ3xI1UoYgl6rNIlVTYeG8qfc2vxiTleBDb+YWVm4E4dorXOAGTJ8m8m4iGk1uxqhRRIlE96rfs
S1MKPKXSBL4ou+VlJTb2Nu+QvNeYEHpzf3405VAFbGEKqScnSQfgZoDVeZURyhBBpdbsXN5NiTg9
GSMutm2QM3NN8ASzoYy4Xj6SHWEfIB9zuy99Z5nrcVK5hHqiwzpMqpTNz3L2zxOkCab+GPowJ3bO
3QhkMv4D3BxPLcAZVKBnSAvtssG4RP+WrrhZXjatrrWyxPk1AJKLwcUdwoKJ3PhWGyt3KBuPlBSy
9COHdnThsR7XaD8Asty3U6pPX8eQgr7h6J/YOSvs1Rs2f5KHvg2qMHVKtultHdD3H6W7f/ROAUWX
ug5/h52LloZJcfyVMMRSdJDi7uyJr1xrhSFs/Bn00t+i3/dErYPArhFGY7YiYNM5DGNBIvyFNH3V
WdoXctW8u+y1U3ez6TKV7K7a3TcJ6cOfHcy1GytOFf+2fiOcnJmv1NpHDi6gWfEC70XRqN1JgavU
03wX5ih3ST8v7VDfiIpE49pGcH1Ccl1JmnkpMt+7//y9/Kt0M/e6ticiqLWEblJfEyHdUUx1vE4p
3oP1QfyeyIpgB2mBNYm+VDu934qKXGXhAnsBII1r368Nc0kXwL2cn+DlVJB0AFEd0Ba674+F86DX
ajJzeXOKJvDk+5s5xOCE0U+aTiP1KzN1XVlbCgq0cVrIFS2gMCMTfR2GMYfg3XWSU/b8mQgxwfdm
G+clzUfWZX/q38X2w6m2EO4c9dxoAJCz8uRBWwEfejz0IAyaGfzWKMduKR/0yZU3Edsi/rXnfSV4
UTMN2JqK4BdF+Rn9HXwPHULQp+O16+MH0wZa6SrQPu7KfQnSNBju2ueyny6r9WHHSyJcFNSkMsRP
k+0nOhQPt8ZuXIovvb83tKFn1NzIkAvSjt0ZvdJ+hSdG3oZGwNKw+vz75eHUcC+Xny0xvAz0Lzxb
Nw6iKL1R+vYl7BIix5JCL7//ZoQ0cQ4Ow7RyB7XwUaX9H7q4tPSPUqI24haMxILgc2pJIlymRq0m
uUqdkQigUp8oRxD4tH7eA7jq9+hPPLdyeEsOCcW7F2bQ0Dvesb0W1hiI/eU2Jqy0k7BGGm6N6bZH
GWEgNIcv7cL+qmb853m8aAcrx5yxvjJTNEYJY7nbtD9kX1/1csq8ovrNdDqPgeZzmsjteyJZXs69
h/+CQNCPL0ULSA4YEo/IqvjZtixq1ZL59V/hhkmSu0vaOB0VwWs+8JuCFz3kf4h9ayhtaMx8RMku
qLtWseCQz+qNzR6MxUKwn4WKtvvWfwZrMEbwxBjLupYqOq8RbdHUotocu50ZAEO5QcWhHhKhVYDD
o+6bs7dGtGhFkG0naYjeFgPjCuEwN4MdzuksjAo57F0PItXRvrQ2+iEcc8z74P+dAk4J6BfDRhk1
xWaacJCXeKA37d0Z+TkK8fBBzAIzQeUvI6fmRYuj/F1g2xqFpDy//nck3Ua+PlMy6diEW8u1qto5
/Oq3FbPIknfLwT0u+o1AuznQJbgijBd9puOwhd1hSr5yJtRUrGLzAAOJhLjTCqb/3Ff42PIB67z6
WqCa1q91ErukCTn7wyqolSNnMaqKiBtL+7IdLMwnUmMJOogZpjEXFECLmGoLRwzFgJ/Ymrhvma5e
jiyeCJWIg8xS0UDLFBGtOT7xmVNXGS+tUm4W5H5Gji0zR08/ad4UqDOaQGFTbr45lYDqE3ZBJaMX
YKWr1pNpGe3scPvcap1W8uu5VgzNOLY6H0FwGaQLq8YlIs2NoVJK+kNIH9uX7yZbklTplYR4LysJ
KEMQb+EvHoqeuNubJI6x5aqXxUTTpXUr8bEDezn+KU9CuJTQdSvKpd+lH/5nMBT1xdN54AQQVBFM
0xfNIQyCpjiapdoJYrNbdRPtbuyF4hhFimQEnfyyH5Amu1nSHQSgFhsWUIlWuITLEmn/gr9sTI4s
Oc7fuDLXU/AGwc6QEtwbDyxpyL1yC93lLmiZVRF+WN/6cQxYm8zqJmnSRKTpVfN9+dQcQnFpyCLL
EKR1swYSgj8i0JkZH6bLt9dGOqXNCaPY1uDOYH9lZgXYaGcS3dUyn67oQUfXJ6efB/o4kZUQkuEj
+Ozgdf9kJwesbMUUeqpKQTvT2dFRsGiXx0gzJ90XlW+kXtWitqOoCH3GKNfocS1RqRgAHqmIsMyt
rFKPsZc6kyZUrhjqVK5V55kE1nxhG0HGyBTZFxc6Pw+0ohxKwi4Zrfoif6i6WcKIaV00maUqEPoH
udu7ATHVapCDHwIEssqBSfZy2YGt06nj/1oVqKTNG125eTMjchRLv2VyeyOfRuzjfjRuAZxzQcEK
4y/KZVD6MCaAl8BMf8Wq2nQLYAOyUlHruQtum2NWHCzJvF5lty0jakvJSdwAm2r6bnbMGQfh/hWC
wgviHkvSGjs9FsFDfnvrzr+fLgkq/Cpv3wKJDtuwclewxaOmnKYAwO2G6CCcWm/ScuOHzdWu813o
jjwe6nTKYvZ43cFHeQzhsHTOGqpes6if8RIAYeYJVtkQiZ/FuScaM/mYx64HDIYrDVTcePkrH4Ja
vg60sG2JTYsGCqmP0YMtomnka4SNM0FIS/CMk56AnwNGq/aMfWYLhmmsMMMsWxWKecWHAEJ+bYGe
Db3ohHTYZPB9pjmpo4OkzEahfo2jpmJ+gB3A7Rw0P4DKO1kUJZYHyLOf9elaIE8vqKPNu5OVmBJI
jNKQNgVAuyc0wP8QGps+CtbnCjQnA+s5TtucXfZGB57YhcmUAvkD/77uwTJ5v8+PLrigr5LAv9xa
1HczHBEcJlVogNHLOsiohMxHrQukcCVBQKgNtaZ4Vo7uDnFtEvPiEbg1F+1i2a+ZBZE7EnUM8Qv1
MRKP9Ovk3QnIl2ZD+UhPL7Hxa2ze/cafMfK8oVXVvbi6no0Z4QUcYS8d0XxMNF7dIotDphI5Eygz
vCNiUcLIWjyIK9ySkeJjS95rE50CLFWIBSfIkBNI1O7LoHxaqTyFsKqmSw180Ob4W4dm1OS/DlxX
AVqzMv2kejwV+o55wykskaMXx5tzd8S9HDa/h0QcfIa5LpOKK2YVxv11KtyQGE4of27KS8gIbm8X
4qHT1bqhnAUCnGn6WfzgVuS/h9T1ffa9/BBp6ZAfMuLqyNnx3Qem1e3Nq0DtY/pDUCGFPXyWYcrq
HDMXFH6PLUeMadAzkzhp21B2MW2vsz4yD6fpiPk5X9gMVUeEsa6BIa7GWhRnYyz8498Mz16vbhgj
r9Q05IGxkCjfh09GNwrIJD57+tf+gyM9EUGMe6aDqeNfyBplfyoMFwj7SRc5aitPP5znKbhbMWST
4eySHDEi/Ft8tsND5U9SrcBnvf2EJJeAmnT7cC3hXViMKrBERljRVl9TmbgksAn/ZyCc12mYrCfk
ZhP3LrayicoEx5WBGixYmSXiBpXWzUyQbWAHRS5w62NLWzJ5UYkLD7UCEai0l9zKuXIYPkIqUe4z
A4Otc2WgL9pZkwvCGGJyeteEukwB9dv0EVDDI6QzHu81pqBSH/HstEcmtabHgkfL37oEZp1nhK0a
fM8xnpBWY9P9ZJRbDVPYQki3t8y5UMjwFURmlvnPRwSQvVf5SasF5SxGxy4YczX6pxZwYi/VQdRX
Ia6+gr0sBwnVOYXZlBFMTJV3aiJSeKGzC/SEtmvWuXUZKW+KZS1rXZA9Cc7os1rmjbxNelIpwCOu
BPmJ7nAK5TsrifKbHSJg4V1q65gOmMNYwGYOHomH0gizuaUfZaNi+Smj5kWIhp6U6NRtnJ2qzpCi
vNQ0KKgNeaVwJEK6Dq2hfPn+DUnt9KetDqZC1GSassOoAm3YytawM3jRHSRySGRIJjIeVqLWNEDA
kkvuTkUY8dahbAiEkbtIVFRp4K2RgM37W25Tp1ZqX3bj/JIbGCYY1B27NUFKYfpMg6g0ub3qFqXr
yOAKcy5wGwLUB0RoD1lFj2zYggye3xo8TDiyyeMoq3Yw3EpzrCX45J/bSaTlTp47V/0ytXHUyZEj
c6rFMy9oqvVsS+g+AAHaBVZGp0qgN/HeLnELETneNzgK9tBeCG5ykGle8o0V/qVe+LGZ0YhFRDi2
psopk0MZ2aQIKZVkJvV9ZyxImUVu+wM3aEPkgRcoT20UzB9mhiWnOgBLApZ7PaHtlhps5pGQRz3F
ck1qpP7m2nA7upMwXVKLZJ8rFhkTWxir5TND1SjmhJRKkrmmpK7kq2VrZhl6jrcWmXJ2EDD5F69p
NQ8Rk5HoEDVjANdtZu1cmkqNozqyhKB6tnEsI51weWPU8HBB1usP42zVtoz8mha686hV/eXz0W4r
ff4y8ltpYMDbr9V5PnR8wMPQHHaYFZqJ83eZaUOlvZhuLKl26ZdUeJVGEwUUB0K6ix/DdqdJ1Aj2
Ax6mCdHFFS6nqZ/BL9nYhUaS2Qo4DuaQOOmccBUSavpyZcBP7BIUAqPvPZAaaJxbQ+QgrP4JdAIR
UFBbdPhJ9VYOXFd4P8VUh/axtcBXmKxG949JCt9AgWA2AeWnYBKoX6OY3uItJ5604d9pfsfA8Yxp
w/D3gKt0lcb94e3gy8uQDct+3W9QVSZ/a0nQTijZ7bPH1w44m91wkygPzS8IoWd90Gnd0Q77s9s4
Enl5bJcYOta9C9QYIC3Lv12oiKTtMbh429vhDMgzlx8o4zIaPT9niBkd423t1ejs03b/B5RXzyX9
cWJ7lh60twqXdNcmAH0sPkJVr1gVw2X+X/2ldAtcf6HL15Hqx/sGxzXFZ162WWVRIeeaS2udMkKq
oinmVRQoGPUt//XZgocdiuo5kIncbXANtAy5UEor6aYWmZLjkdaPUm+L2b6vD9ISglrgjRS7prAl
41BdgTkILm7L1Rvq4ZgCv0X7VmS3asRi9BX2LiKZBERIZ1eEZf26s4/EQsmAOm/t2sQkd6vFEyQe
EmV0ZNz3804f353VCWafvGFHyTonXQNABy31FrrlWpF+QprX3IGCEwsNnlY/ISqs+LwzrGzKoahv
Bkh5qo3Amehv8WHZVgYFgrFyfiE/DzZytDLc3tueU5Ocz+pALIUxmUU+Ozs9GgWV33ugTnSkLJwI
NTiFmKT/39BAYJdxYmIYbbnLuHcJx30ggLKx10W56xua+lmpqz3Lkm4qNbaDXzMJlhYQoV4fMInr
/dtDJlHXwDkJ8cI7cmA8MxrXBiE47RKQmhJjSybFSs3HW+0/nTCnVDLNcBbFXfLMVpY0LYfPHILY
ZJBktdeuOzxL8QugytPE1VzembCJKUicjX6IFbGtYrOYSgqgklIwjNZZxrl+vYkqPwJ1Qk2kEZII
x6HrA10odtzNsG844ZX84bdjRRrHatlg4FLP9k/ynIvZ3oHyW5Kf4J7IQTTkat7LqbDMC9V5z6hk
NbWeAB4hy737j/4ZRL2s0D7zH2f2cbWIzZjl0Yg8RlOWn2xruea/vQtXBo0rER69lckjSNn7pI++
BEXFH+LAmbAFt0ODcDAHdIcUscOre43orCRW1vlZf3MHIyYiHstU0Z4XUeQ8006TS2BxvWxrhWv5
tS52+iXPe54n4I2crVUvx1R7diindI9tpADij+Z8S7MdQHWvcQBWvb+BNoNYsMMmueA8EIZFKT74
CKatJ8OrNukinT9aUzCo4+M5jzPgLPWTp5yXDVF9o1x+bsi/0cNHrt0wZvWUuOn+HYuaoALeK4E7
6ZAD7656ghEC00A0h853wSpkCMX27n0YF40GA24mBWndr0/tqQ0VDffsItsFzN+aCdhG317hqIHw
ENPCPH3For5b1J3hvB333HAON+PTsGTRsFgNmPOd5JRPYt3rRkvIBwT5/EXANLdkeuuVKE3KIdtE
oMqTRCOlouRXgHjFLyi3pu6cAnEqYr8ben7bIQ4SvXeL8mZMPQ1XdBKNop6Va4qWiR7T1lwYDN0V
+vbrg9T0cMRN4uTtO9CpUFFLtJXc9Vs39wuyMs/tZHiOQNa3PInYg3VNoh5wZqnq9nSGw8hx+bGc
paT2X9rxmr4afaj2h5KNxUOVdHBxNVFBxrCHkWij4yn+oapEbGztXzDjqiubn/P/MzDMOTwufliU
XM2u9HUTD4kXElkQ2+UcjcZtQtNmCZ4JJUFm1BM12Xg1E6Uk/n7Dzd5v7SvsCg/m7g4dhxivtmGf
qd56ktIjiCWxstKTG1CuqGiK2juoHEKDr4Rc1WzytKxVSF11lYqy4D2le37eMqgp56z4Dzxbykn8
0+4KTIAd4LTPu41Am803jPeZjM8ZdB2UcBr15h1PhHlw9uk7TAnKv8RQwHv5/ogtFZJpUpgNoUwe
Fhwzk9Hp1Ouo/sGuYTx5tLw2pSznQInWhtFaQBu8V5cSC8TFnC/QSrI0gNuoYrZENf9/oUOovSGf
oAh792fZb9UKHq5YXOVg8+erLggfxoLXCn9b5DSww8XIzb6Bo4PM3RmXlGETHPU7wENcRKaKJXkS
8mOM5gqnmeeHEaslO/pIt5l21+4wyjHESK1TW/pCZbvdcBJeaB1GACfCOv36R9ARVWaHiKQu4Elp
kKO+UvvYIHtenXsTS5sBJSpJZpAPXcyewPLKXpHdWebUcb2iYiRb4JyhSk0f3FxKIip9P+2B4obg
9+IaN3JXKM1FQxmgSrHnUy91shUYobcd2IMehalusKXVXmYzW+A8dR63xYGX4WsVHTTnLp2g+B+U
LzJ6VRRcKk9A590Cm8pj3gmt+z7g5hZ3n6f4TsKzeCa+QRtXKgYyfv7Xr45gtN5m0zG23fMs0vAi
TPmMIVNNzooDW/m+S3p9gtMheaLpfmZ3m/hgY/wbAjZkJQkAQvqC+TXjoCe3bF3OGwD6QgLACTRy
YN1+FyNeaVdBTPJ/Eu+NU6/c/thCmw+WUuSLmYQHXHv2tMP0Dn8LRMN0nyp78EMnjYs93UYW0YAR
DK9VQSjlnNfn4L0AawYiJ1mYIgFrjlntx+/Ad+pln4IO/PFDXh9klopAb3P8aXwDQf4A4g/M37Ai
R6USOt71dsboxDGen/4sEe+t7RxpOHjLgQWiLklWyZvt0L3dprvScIdvRVvLt4QOzXbQMsSmJ4+o
9PZcuOSG5Q3YENhMB1zzX1wEzCroTBsk6LPRdV7FijXL6wJF2hJpHhUf6QlKivYeuP5guSxjKOFf
9j4m6rACMw1G/Awli+Ia+UURdOOLC+7qLoX659IrVTPu0QRxaD4drTorGelqEKjarivI/eufRMsy
Y2lY/Mw+MIvW6nXy8PUPe0jqJMmO4jotIbDsdcIKZPGMpsgCXj5N76TVrgaUMB6Et5K2jHQIi0ZH
wWuZL3dlSg1nw7go7l9Hm75ovuDLZsCTOLXLoUJQClw1p/SBwxeQPOWex5eX0S4d5zSH/Kg80ll5
7ebwXH6wMDNQd8GEdK6RH/9PZf/GZWzfXnzz9fN1xhVJyMImCCUs47V19UzYrgOk73RTWu8e8ABj
O4vCdDTzLuEDKdnhPpdLN8lkhpecune9io1xzEEjKJbhsWcWz+FK6ximCmeD9QfQYrgujPgy8G9b
ii+n7Hi72dIgX9Y2e4nIYFZOTa69XL6WHvFqewOSiBQg2qb9cBv0JBwFwcXJQ0N7oIxb2YqIC8Ta
5lFaa37jeAamRqNEyBULtAxBJPPfb6DNeqM441cxw8BfrPqAOEtK4lwDA0TyBqwqm+PDt6Q5iVhM
6BMW+duGGbMoIQ18Sp+L5vD1qAvN7xgCW89AtTI32CdGkN2mOKZOO6NBeG1hRe6KfW9K2BSjpRz6
plDH797uByVcBmM69fA4AB3wPzE+KTbas4Ubcxlhnvm09IYXSp4Q77VrKZF8jN8HXmM3/zxXLleN
X0gzzX+puhz8XYWMfjHEMk0MUYVWY6U0KHmctYmUPta80cPd/N1H0+8ky943nMNac0z3JxEcC1ru
FKoNeWyOdRtf8QWq2RQnv80YWlmiaMYnWeQ2V7ZhZDLqSe5ioUH41xueb7rden6n/t8JftObtfNx
/QmA67UgHKfyy2yhh6dhIePizKCNxSjiVJY+IQL2vqX9hrBYl089PeyJSMu1M3Sa6gOzcGyxn93Q
yaiLTfQqSa90Yc8KMrhlVj4n3HiZZ9gZbMP2FlkWqcgJOE16nZagTxLgcS4vgSFUe1yFOvo9XSlO
AqS6y27V/0Y34GIAE+46IVNKnpA0uj9PXdt57Cs7+Fqbcgt9ynnAnUHoUni2Ol/DOXTk0DMs/BAh
zzuz7ToxRoTAcXKPJPYnsYj+NgWUFva0pnv6YJLHGmnHoEJ/xHjNIKGwt7vJzN8FAxRP9Gw4g6DX
fYJoC8rr1KXP+OnUCdNVeCugIB9t7zg4ZtLw25LSMWVkGWtk1tDi7I7y7py1cYqVVlr7sH05MM0E
kmm8XiICVcJ1n8kyezKSkc/kAaksQlgXV55D3Yw0kbyFumjhoeceFShEl6ePjV1bTNtW5Z+Gd0V0
zRE7uMsLbDQWGdIKh7iSM3tsnqot0uL2/UKN3yEzDqVIjl2gPnpUTObcNsod8bec3+1Q9H1P5iNa
bh9ICL7LpzixNrVupuxLvxhMOIe8vkWNd+NM1w7OxMGgGJvC9KeFgiP0kMMA+BDt37El3EwdBO0G
ZluFxeaSCTP2W1Gyy7Fa8y+E1tXE1Y0JyFhPakOggkK9c3XwiXKXGBgokS2lYmo7R0l8eWXH9KP+
QsZG6Wvvgo1wfJiDeFohZymHRbuyVUG1syn4jUllZjE2GYpYR2DPTItmwoFNmxFZkeORxyf65xB+
ofjwZs8qv0t6klhsttW9byFbnS5iXNY8BG/tc1tSIk5zhPftQryL68/6loNhuEkB5aNPws4iqmJL
H1MNZDFEZdNmLsI+lGC72CihQGhOYMAJwPRfAKelcLtYPYB1RZTAtzoCZRbiK5AD4Nv4snCAGCC+
UEi18TYmBdWwuZejjQnW9iQXrcPSROsDO3SzhJOZ1QXbLjmptSyV1N7/5/Wj3x6RocCkxPFTL81B
FDsLgdOTt2FykpqeIGCB+9N3JjtSNnP12tt4RQyiopbavoeWXdOttROI7pnte5rBBYNPw8yQy74z
aVl31yKHMnwhD4APQ+uBaZVYE/joNHu6NnJ5tEYmV9D2MWIDGyZurxFEHygNFpfqmPDjoddYOKd/
Ara8Cp1k4sTpviGr8vdVc5u6LVl+53wG9Y3G0NLi5Q7xgUeaXqxKKdb4tsDuvPuxM+VxJ/3j4t0E
f8BZptRiy2vo0eIqPej2dhF/MH1xHcTN2aCELDplzF9Sx0ImWozI9eNIk9gwKONNK9dowhfvGYO3
fGL0xDMMdqeMsPAEhdcPGZo6F8w5WN9ogmoq3+QHk3eT/dKH0PeZT89owmGto2GlK+oBw9EhXsgC
Pdvg3uT5aHo+01BUWBx5PLC2AbR3Gz5/DNFy+wKlwybaDLBaqrhhW8ATfvXKOdb6YXc3Sd/MN3OZ
Ca4jBBMgsJNrAyMIeqbhq2Ofj3WUyhv8RsA1QKk+kG7mgg9V++LW2i1z4OZXcErM3Yk5Z46dAKrV
OVwL5BSgrfT1kbJ3EovfP9gMUbpaSmM8JgmYrpCrFIYZaqxV76FF+MOaa8OR5E5HzFSq+Txvv5+/
czpgo6P2IA31iGx5AcMveSXkiBGq3F1j74CPpfj1kGy8BzyX3z/uveKCFjJH291B/LfFaLiOmqVY
8LJKqJdCe3+Z53fi38YwcD78BBt4AvmqF0pDTXTRe6UHQlljaeGJa0BVCrUmceuprNja6rYB/0gt
W6mJWESFhTnGDlnGGN2itYXO+gkQgsrG3DQPXTYNXZSYYWigVBdAjIuI2IYBcxITr1p4I5RsYiLD
2oN+8aQ2Bwr6nWdubMfStF4+LBRp84AA3an/EA0Ld1bMmGpNCmJpoggqoK/vlutirOHGr9D6DBIB
akBiKaKBg1AImihFDjuIfwNgsG5LcQiy1gfdbpj8R5CaOwnRjzYsiZa5BgYYEg3XDtsjA6JKmiGH
8Rj+Eq4/Nv7XSw38ZC+XFKLvRI2wn3IhmeP5UAmP0I839pkCkR3ZZkmJE/OYXkmAqse8vV7ySlRg
eARFcE9DAV0H3S7fEwqulPfZ+7WyINFpgZhCF7OlyxVDcNVOJqZxiXCBB3RALe0/GmRlZR8Lnm/4
a0mQMAKIm+43qSNw1bmK9/FTp6DNRmhTyQDba2WF8fZ7HT5WCmbsD3Ck6SoXu6ZzphFt9X4YGpa4
VX/1l6HFKWnDSSOqJhlCWMzM3cR8Zj1WYCCbPuW9ulxb7Qo3pZ7S+ETmiRhoPbWGCqAJiegFfXy1
DWuH1qWyhdJ/109YRt+loDrnYlp5pc6BxaSySnR22A/eebu/Hptn3z5e7kf8CHEzimjIPHcwcWE3
P+eTb+BDnZBM4D/OHbbiocfA8yrQ7winrSWnwxHJUvJp3hioOeIH4K3l0OGo+pUlxttB4OB4KaJY
OFL212SavteqYDPYk50fUOiuQ5qf4rEvsC7BhirWPA6mpeThBiWrRHpYuHLtbX8zA32Z1WZzl7wN
dW/0Gy3Z1GXRR810FmwCdsYKKR+3nu3YFkkCEsOi8KRi4vGHKrLzwdbnGBR6acSSqTuoruDArBvL
RJ80nH/6azkRuVaN2lJ0K2m8IR2P15W2ITgS9cJ5AFrxVgOt4n34yryqN9lg8tjhqAZ83iUwLvJN
PyV2Kkzr4ogz6q/9VWutHA9n/NT+h5bRxpHYTZC6ZQygvytYobAXCZDFNClT6LppOCYS2mbmT4wQ
KCIze7HGk1kLoUb2z/iUo6z1NP6w1jrpEgrc1exj+2MNzq22RMbsK0W6I1bx6bJ4DWF8CrEDqgvM
FYOg3XDl9kVrjXeqFDW3dXTmdSSDavgbYUmrB+h8MHOfCCy9duzYsW4LkYWXSEDVzKLlU6C+DcwG
cxSs6oC3NHdRmPLzfm3W9NdVq7pkT7yDFVxFZLD1KceddsDUKdrdKDTrU4dj0FqIw6AvKNcaoNJE
dWzVliOAk2Ha521zH7OLIzm25suun1w97/QTf1JycjRDPMRodQemxA40cwqXR99I9vj3hOF7jkd/
FwOT0PoobMpLdzWVsOt5RO9HT1ifDmnouAbJEUhCbmQ26FAGK5S6ZElo7dgXyFkuDN9B8gaYq7HK
5g5oUbkjzSjIxf6zyCgJtFgXUm5vX5FVwjgL3mrVymZ0XCHKNTWP2IOwktW5GIP05WyPPi3TkOaP
pdHM4aXJiYAlDo8gNEQolewnx/9Xt5krzM7L/VY6o5TOnnJ8b1TEVL1C71vboNj9zZhQfTOZWD5t
l4b1C7IOSa6cAQB5Bvf4x1sqlqsjER/G0VYOyb5oHPoIiLFUnACvm+qITGOx8utddkxWgAjAOBDM
bOhtInnsE1TYh8v3pw/At9RYvaZforpoXEqhSfKYIc4w4xCZxetE4HXPTmorP3Hk+NoN0O7QknD/
t45cSGoeB+DTKUsOf5LS/KiBU5SXc19ahY69VjEBlSihvdWKeKXlg0M3Ot+rO9pIA09pgCs1mlES
09UfaO+wc1tnGKjk89svGXs4KXta7D9oTcoL9iQh3k4wrbZxoh/RPYN7fscnTRd5KuyjgCi4HF3f
JvzD80Z16190ejRpFzKrwdjC9IbgPARS7p5Pzv2AAV2U4SCep8lWPzCsKWEIa4auCuew3cIJFAxT
HsQZJ6Ksy+Mjx15m6ExpYOFXDdg3dMd3f1klNMij4RDgk37L4hnOtHLG2Z2iCoQ+EsNXRrt4C4c7
shM27O5HXCXL7XW+Wm6jVBjh9nUQ8i5IYGcRUh9PCoWymwjmcSNF5ShTzCFLLmZJrAkbY9z7tGom
nkfXk//Zc3SlaUjI9e/RDci9icjbMWqr29SMsZGur1mc0XGKUS0xSwfKTy5z3ugyWnTnU4oq7F7k
GgvskksTscm/9I3D/d8aFa5x4jHQ/OiT/iXCT+eBBrCvSPRxOuEAetA94WNRDKWhUwIs8rgPxvGq
QbgZrhYXi6P4SuU8q0CHVvawNbgNPNeeVP7ltwoJRXBeIIbDMkT1YByWoz5KiZLSwBoyC46WE4Ja
GhLL1DDskR1c2dq0RwNWaRcK9uHg6rgUQxR/PUphFUVIaQhvNlYAVJ74tfSlV5gHRUQg8YKeDmJ3
JYQpUtCReInMxn+Yhp/E9ffe6GPWCuXRDgiPPqadNtxOTOVQgb8hQLPswS3GZCHYHc4msYtHUG0+
0F41v7hvbmvRuYP5oXvrW+RdfwL2n0QiV0T3bm3uutxTUvfpNjVzoekvrHeaaKpo76vexEPMzmSs
lEm5iMWVIq060Ck+wwlJhlBDXnFoFIWFB96k0xjJvIRtWb/HRYV5DzogLVjN1lYILj+xuccY86xF
r4TC5Wkm1YCGJF//KfdkFwBtO0Q3+J68ksAhPBmhbfNQ3lWS6++AHmbTlj1lSYnbdM8sw8ZaZrX0
Ha7OrTZ+1rDoaWW8NgWrNE9oQTJDQ81YSZUPFIQEmR9Af9qVN/Jq9pz8eiKVBQJEHQmfCPTSAoqz
1MXVKrfabAjlB0qL0V1EWU175eZPmhWaDQ9wzNeFSl3+E42avO2YQRvz11c7bVxHw6jal8lzJW+N
eswTtnRcMJ9gd5c+9IEbR/9FdboHw8wfi8FS1cXhl/sEX/+smMT5AByochpR+UXpbojPVu/am2fk
AprT2dfn/03DgImDD3TxWNd44sQvjjkm7e/1y39iQnRDJXn9dIVgKyy3fYcb57x/UKsLW61ial8A
jyB8htBEhO547Sp1qBEf3dxGFvvnH1+u7xCt7FuEvLVrD1kBXQE0X3gwRMsIFAZjYZwBq0AYZ5Bb
y2KMHFggA77Dvkk3rCtp3ZNulJCuu0y393PUUIrTZbbEOSo5N1IckUzJL5LAnPvQ+6nQyx6nyXJx
8fGucM9SnzJzeJtDWvlDJ9VRR3rUHXO+RaN0in7jCCJZJLeig5Q9Z3JIuoUJUAQvD9nEYRu/Su7Y
upu4OnickmLL328jBoMh5ZHBis51Uvo5UvL8gHwcC8K9La4z/ZbKOVvt0EKy/DbvvU6RVRukzLYP
USl4zc/iR4PCOO68qdboRsl8WPGUd6qbSuKCwY4owm3yckC64Jyf5vjQogB7MjGx+7Yeb6d2gvci
dHWToBky+Xrmke94VFoQ8JkIp8BGlkszHZw8fjcWCdtwujbVKVa0b3r+bN3xkJ8I/Nf9h4A4ZuWi
la4CwdhmR10t9Wm0Nj40KwjmdIG2O9Kj75ibTYbAb4OC4zYqLOUD7+bqvEWYPfB8gc9P2A8gRiv9
GJdAVzYY35kdH59PDuHw7tQEpZhnQNi+ibrRQRnVye30FBbfxQJUp1kyFRFbr1c3m/dQ6fw0BS4D
W6Bgcrc0BXmuHiTJUIrsxirlVi+vRi+/oOqfY/ayOI96/VvdfJxxOQk7yrB21IqxZL7ZXAGNmJvc
/KALKz9yzkXDx09Av1T+IhGkYsydtmT9rQD0oImF4O2uRmXCnw7SlDXufF5eCL5MQ3JQ1tnScaDL
YG/20RVvgLq+gfp5QatiD69yGsbsCZayMi3B//ntJNgkAenEsjm2r7CuH9PQ28d/TrlGr0Da1E77
V6omKv/gUVeXudEI6WLF+4r3atUe8jD+po7AeBDnajcRYLjjYr3ij/j4zhgQ1m53GmuLhuWfEVh+
1ABrS/9s2T/bT42elE5mhmYk1siiuralMCojoJjEZkkdOVcj90xxvmozbPGOgCjK6z75aQg0yVYi
hEE/nLAVj/zgvA5GrliJj/OPEzVeCkemrtBH5jFkoS9z5h5PW7l9a5Uv2EHyYw2Q20Dv7bQsGPJa
f9MyiEXqVANzL0nlzdxCHSYBy5n4D8TIub+PfSWcqPEF8/VdhXGmoSI++jhLL/vL0+DihpZ3KSF2
v1MmwPbYmPIzfmycRB73nW9VcL4GE+1aYkLHbAj3kZ5KNCR/QOJq0OuAmdgKDUrn+Sy67BDmYWCZ
iKkb0Ou4CjlEQyWrBX8W5wPs1OrWFlRyEdsDuEwzPi7i8ukCUPA4IrlK5Fi6aVuBkAxr/d1ZLQRf
NeRkZeS3VUCltmIQ8W0I+2tSIa3tY8NHJFgO740dDgxfELNdljVq61Zz/Lh9W94fLHAsRu6YaL5b
/14AbuXmSqhF7j01SdKvG7t9y1UPqE1LePL3MT6Ajbi7v7Ko0Pud6xVao+GLQpvO4Y1K8yWntvaq
amM0NiIzxsB8o2ewLVSf0RCGVeAswyh5saITNteu7m2wqLVF2f5lvCqngKmIx+kYBTwoCoK5d+Rb
ZhTOTxQAhbfpYP0rema/9ftjXSvOAPRZTU5r9S5zKTXddlxdt4+EEpaTMeULwbjhu+RM1kKdFp13
zLTD/kHc5FL58fEniosB44K7CfryhcHFYgVZzS8LzkOw1bj5vBKuisMCmQ17IFpQAk3egcE0RQ/E
+nEY/UNUNeTewsNbGbgJbdhkf85Z9hnbwHfmrk8gRr99SedyhZTs8jEjYaCNzAEGw4TpoTYxLPW+
6lLnB2pygBeRqywdmJ1eGRsZnFLCLXlF1nIH6rQzM5NxVNcjSCljDO1nYLcov07k7sv400dSbXUE
az0PGiuzFM0ETNuISBCRh6B0nQrq4AA2dAceQvcU+JRUPwALGJQFjkb1+oQ1wZSagiwF5YYb9k4c
14i6nWHLtszr7yUcLGSTsOfuCYMk36ePMv8qB4+zPk6WPdOECO9MqvMhoRMmuGYfjLcNZFxYOqgN
Kti13bAwZKK+YYeseZIGOC4DVqqcPgce20mWc70iXuEEAmSYc5Zh5xzJ+5zK3Ji26PWHqfDMjWSh
jQzuwwvmH3/hZVgXJVYtsGJTU+vowcAWD1SVU/uyZqpbrRooKJTBH2Z033ZUVxL/4SUl86Yj5Ed4
H+saoIq8IihR7YvzuLztOngiq/pnw7BfQ2o6nVr7bAkRHkMpvAS26cpuXn0pYW2WR5noVSDADkMF
P1I+/oY7n9EWTuHv+PVHfy8m+TvOnmBVYeCuxi/qpbiIKXn2i212t9G0m471VOmTf7MHVbfRsPsf
8lF5E89ODad/IcgIHXJKhp0RBGyQtw/hiGOJzgJ131V2FvNla6IDQvmucodN8RUVhldSe6uIeUWL
dQsi7w/rrhWeOBhFqYEBb4CCeYPZqspJGBVtzT23LlIRWfKACxEosyUtLAM3+L7EV7TaV97nDTb0
EONeRX/fhJ7tiqAcXRw4HXlZfzZJEySSHf3IT6p8+vrtTRqhZRu8tc6VgJMyp3xNUtG5bQ/GoliZ
prgCPLqZKEU9lYhydyUaU/B1C57/lU2gZSymNX7GLCZ3PaGtaHEeFOWQJNPK+IzpOzoqsr0m0v2d
EejRWone74D+dxt9n1rBY2bc0SNi7GkXGcXWhLjjV36+enmOw50FOpeInEs49VSQZ2wkEhfObOF3
ErzGGbg28CjC8pDzkNP5bqSJ2tziXcZ62cOzf76nk+aGKpsOpUPn/+Bf7wN+MvoCtg47z4+int55
a8+ovFWFUD5iuf2qSwCQx0ZZJUwhUtgUCfskpTqkjJAxULJjLV1zgkl9K07eNgne+mFEoeK1Fogc
1M3WLptqSlp2TPNgsxz2PYhBW850Fr5Am2qvKkpj1YGnc7PDSGil8YGh5LLadMz4LHYhUM/Dtb8r
ivPmNmKqSEWWbywJ165xiQhpD03oNoHYP2z0OGOMzD5Gqq1TBhgvs6wc5WvcA9BdjaEPk1+q1bA4
axpeb2Hc+yAbSDTPqKq/4tXYm6cAw425HwsCak2PGdjlk0/rUfbxDOGIZaVzgMd5vqtIS7F+q41V
rCvdbP1YdXdsQN1u1Qe50Ic0FixsR4rXrc37xogYV87igD7j9uyxuFSljuZaoOXF1ZNRK8W2cGzg
Vd+2RR/XfueGzroUGqCojVTqZIkzxslo9AVHegFnDzuDaUmtphu6AVatSRwfVwqqgDQQczi+xziq
sKNN4tSQj99sQLtvK7zwpb4cA/Tjt3+Y6kVMKSP6uWz5qSTmO2fNQEXau2tcONxtaiCRW2WaCkfo
8vfSOYEHiOVi82GfbiHjLPG4xf7rUbUCxkF/T8SzyIRluaqqeV52Qmvi3WfOwH1gf1q3vcmGwX0Y
cg7Mfvh6k3er1djSu6UEJIHZNwY8g8SJQjDzLW32hohIy7+4IZj2Z3cqn/EA/+2hZvm3yMsY4YXD
hP56k4kR3MRJX1kpiauqKwahysUl3WtGZcVa9MtiHh0piXTD2lFUXo4iH4SVGzAP7STV9Swl2WrA
6rm/JuI0KxmHXOY/UZ5bR+8XOGQZSZxLr22DpWF9oVKS7TK/mP/QZKaCAsGYi65t4ykvsOWlwbJF
qfVTCtlObRsWVys/bUSp+j+Q6jlUavUsh78Jm9ziOUJmp0TEsHEkWavQbg2XU0l2BuEB8VafrcgS
un4XAATKt/ziEviENBq1Tw2stWKG2DRzeU/t0p45glDJfqNdRixBaUbJRqhmW4wjPEKedR9bRLyH
WdB83IJAmfJU31H1qdaFpg6S6JFR6ZwuDLV6aSQP992mF/yNd5WjokTfJur6G0PVXINFKX1qb09f
rNPz5AOmj9gyCmIeIa6rI8FH4/kAjqmmfm1PDrDMiUZC8/Q5OkTmNpUE2F5o7w8hW8LmlKFhWkzZ
TmP8api56EhU215/iwBJfSFy4IB2l0omTuCZQH4hhsrhcKiRhIC3Zabcpa/CV/EEJy/FdtBWxy6l
shcyOA3jzN2LJHmL8RNHBdHdSW6rBkfhGnmMPccXTiyBQ3iiNr2gDDRd6+1LEouC79DGCOqpiBYS
Yy7ddfO1OZGXwNZvEJeNrS5W2lFEkslETBlw46iEMDuPbzO1wCmhNn7dbgiJej4vbxzguaW9rg4e
8JewKl+ZxIJCloOEi4CkUxDvT08PowKfsDrTTdz/q4kxs9c4qwcY2MpwUkdXcsbWB/0abOhD33ds
x8ZyI4+X6ZCvdunyBLUX87SiYRo3q092QJdqrUxacy4ID0yDBQFguZNybLOQLnPhIeY/NgU2UD8w
4wRLovWNPS00KPCENSiLuwGCOSXPsDuhZoti1q/XsZr5tSQVG14pSkk5ev2NYT5kNZUkPEE3E82J
O/83RT0mRrJIx/+8UIhjV2gkkbZysylfCsaCdaM5d6YeOUWrzDcQhsAxAB3VIRti/MHOEARfXuuE
17BV2CyyShnBIuaJC7DT4hdd+pCLL/vp00NkfiabSnYUGr0z72pplsVMR/DHb3+SeqIuGlFuSibr
Ij59GkBWQSrpnhadmhtrtRpSom1Goth6zZAfC1RJSUB43NfKyzLM8ALM6UEQMcpL/VddVFauEduR
10Es9ziHrizMXz3X6K8FhroV1cV5Mk+hdxShAVLakecllI2qmbXxB9FRu/2h5b34xXDq5ZqddLe3
b20ZvJGh6xfdiKlWSTL1ashRCRyKKmsUYE09QRpKH1aJojXO58pmrBbBO3PbKqrEfvYLK+S1B9Hn
sWN6Hr3JAM1vH7lDAJBoFOf6Wecn9/6AmThNN26IxsynhjptfVEy0Nym1WyWBfHtLDvXbeTWqq26
+YNrvhizUYc0SDkHG/EyAA+Seibn4QUROL8OEgEnuIJbJ9/SOV2qNnDP1C4lKbZiqWqgV8t4IuUN
I+G2lk+zv1GSbNA9PAGUna+EU5rorFEmkVAJqIWDKBr0EjfmxvAfnts0jbz/IIWEG1TF8A6v0F8+
UuubjdunP+vbP1PRRDOsLMUUHMzGodITDsYKRWYxPxHq/K4SKDM9Cfp+aIbh77kNkvYvMxixP4Jh
Oa64+fmW2XmN+LaDbQwUpjfFNtUSwpnwNteH+M11nmNrmF6rNcTIhfVsdoQrvRZSCkZAqEP5+PZx
u2vSA0nhJ71t3bcWuiLxVetWKIWmPZ5nx5/vtBDW1mHnlAGrA4cloN5IbejeyMYFllxWAv+ktmpl
Ba+GnPYqkamI2u/oD8R2rkr9IRtksU4XzykyUNkUHibML84KFiCeRp3zbgTjzRxxzfRfqSjR07L/
rPOwKKS/ToPERlIYzOzn3tM9gW0d2PwR6N+QXDitvuxJnt5qS7PYWgEgRvt9ajTuVFanfBiviSJY
ZKc5F+MbuGbLZ5RZLpyRtY82O9UmPRwDe7C8mQnkPXgG++ILb6V3u4mQAKydFxOvRwwtQw/elain
TMsHbuFExW175jMvOiAs/Xsm3il84eey5tqbTQTBPtbcR0pQ6JlLsasOR9R1VQsdT8nG0UGA0jba
xvMCW1lQE+UQRYa3+Bxn8oaX10bPqOf8Vm1e5rVqcBcaasgJE+MKmExkvLhz/SEQ4SnmAYVzW1Vm
AFCiZMHfZrCWQnkjLvi0+uB4A9/oknb5Fi8iEBrJIRY5ZalmQM6bM8B0OzFzn09JtjfyKExIeCA/
M9DvVnNND1YrWxPbf+sQ/ipuXGxVENOLiBo0AiVXYKyBDveVkWNQcpPtMO8S89y5BWMKHK/si/Lg
Q0qtbSZEz5ZuGiIclBqhM7/GORW8aZwXmz/NJXyshkszdkcn1MpuD7hKxj12ggWehHT6Ncux/626
e83TY5otvQQZ4mwUuc+jnxLWL0UDWFilkI3ms/ByiUT8N/NZq1/DyNbxkoAo4RTX31EgQH+8xwFH
XbsIDemyRUBa8L5LmCyJUAq/OGDhSU8m5ZdMSAFsJXahhNnZInq358NAdMFfDYJKJ2OVFppgDVOo
MQ9vD8VziL3jukVr6ZQeC5qCjrmU9c7KUYDYvPhzTR05l9slW61D9mBiFKX9tWga13mkEITI+la8
vf0/1n0QCMZlqEE9GBlH5Z79+CrIUV+mcJY1Sk7ENBtReMGOl901hmLUY/+t387wniEIPaV5+rA1
TQCd+/H6vR91UpR/Qkj0bSjpjjgRyGOETuFu4fYQ+DzBw1FVI0Q82CAK9W41KpdzKs02yHRcB8Sj
+vIzpLlDn8A2a58xe3H7X3tp2PjpslMQqaWIjyhfIklMidIzqFC+gxNNNmRIHFyUms3AGhUz6B7p
DEj9OPQVqFneIJO+nOm0NunpJgfG5TB07MOWnrerXljE1dC5dmaPOypWls2TIs9jo9UZVL01vbSo
X0QwH5SznkKA8umJGcYwGfjFUDpEQCJyCmNiPKDhSQpzOLmXQ5VRsRwk7eTcUm1RZC1L7CyVwB6X
oCn2n9u1DI28/BCLPC7EFISJNwMpnBEeJWyVf+JdHKdzkJd+mBScLUjG7D7LSEFMeP1PFU+NoYco
rFjlDtLWqp2dglVA9Yehvw4q1Pbn4SPyGbLauD77M5XR3bryQSOwxLemb8BtQyKLjCNBmeBaJmCR
1gqH8Av70PsqBJ6tbuOS2hDgFlR92wTxLVeCQlG7SqjTckMPriT7Xoj/JKzdr75rlWQoZyXCc9PF
36NthhTCFNtZzq/i1pok6Cx0G+XH1T4ZySjd9UyPvvfHoJaaHAF6VAEROsagW9ln6Ovc2bPIU/Dw
/WgGQCAJPtnSbbU+m4qSRX7UwKCIN2f/IzaxDaOZ9tydJ3zLJP1FPgdjnG/KFviz+x8rGvZPOunW
/XKnl6XQh8zY5eFyrYclgQcAI/8cKlUVwuIyjPGshdrzeF2nQ/nd2q5PuxITcfLR3dX7H/JIhQ2P
xUnla1m8j19mgOhPG6t9S4MQlED5Ynlx5ALVLCZ80e2BOa6tUfrFDTQy0R9T67C8IM6JsvRQi6/q
F3wuug3nMr58I6M+AMUdMQG/O7DLgzqIH6MF4LZhUJUexPEewNppcBb/oRgQc61Q88f3Mi2qXa8X
wPw2ariDQ20xvEsU6CeX5WfQQ+cIq0P6P+wZX3VZMoJYPW4nkJxxuc3sVnmRp1phRai36zVYGzZ9
tXbKMrOeRQzFONRNNc8IXWj6nBGu+QFkECfWmsGtOnKOJwUeXtlE0gMf0OW6YFwyFGwagjmhCzqM
vY5a7mh0ZfmBeiMLSYJ22pjWxZS6de4+mUzOTASG+q5Ig+xgwbZnmBsYC4fEhL2rlEMBkvQQ9Udt
W0nOniDltC0MT5z7eTB3BKd86JhLKD/v8yy2o/C055r4CcQUL61v78Zo1rOoKQ/CvZfqOshf1E9k
eaLzefm7bmJFqx+823U+etEyrdE6JTC0xyT5WThZ7hHMRCCf6VeeSdy4UH4H71csABBkS8PPQ9PF
/rJtIThWmXJt6q2CW/p7PDVwaHVxYAAKRheO2KOCOdoZCN3iPECiI+e6gdr9q6QoP6mDnpX84A12
Ib28HDCu5f9NL/5ggvLl/TzM1/w3alj8YAokYVCs5fdQlF3KIDcbwjBqHQ5Cc0Po4RdOvq7sH588
OymrzVhqdJYrOciZv/8Usr0j8m2ayDNOrzuxvLlgJcKMkfFlNE/51ytjXzJatM//lozTiab4Oluw
LV7JbRqnj9skBx3BkCw5j2TnWBKJhBGvN5p0BIOGBI90QNz9U+L2HnSNSgohUkycCrpW6f0WhW2X
F7W+h1tHJJoDvo1/8tfFny4uc0Yc818JrV4ZmZlXP2ZGxsaCwugXf3DqgM5iireYgW5mTdI0lDE/
Lsx9mKoQ5QTUBkcJPlQIENgbdhYXcc7f9u3ScTik91gNDWFk3hkVDNTs4ItPWv8ZKB5KOcmE0TNJ
3GdH33ufm511Uy4jJQ9bC698YA/OdXRIYRL6fiQzuhRVgaMh2p7S6XokX7UUOm/yxMsvZiv3km8b
4Ib0YJ6W3mkbjZrvgcr6ozLPB8DNdfe/8xVs64WSQO0Gd0sE6n3X7q0D7drWfRdNdonUIDD1fucg
3+VurrOm6PWduFA3v6Kqcxn2R2iUM9sY848dLi/H16fIH1bUNcoCS6us8AF6sCgHPV6VW7bkva54
3SG0TFlzNeGscquShCL5CrtImq59pRfbHlnmz5IlnbycY+RAa33vxMS+rT7LztJwjSybwgsjrwzx
LS9DMSbkYhd4DWSG/yAqBrHqZ5OPF+mlsnY1CTVc+TmsozJFZqKH1ozeK9EeyyvLUA3ifSqx/bZH
N3xwQhjhtpNjphED9PJyR8KWzAIrgKX/O9Ggr10xfsD5S8ibvbiHcBlPETovaWIZUGZ3FXMjowh/
hNVyIb/RAKqvhmKg8rcfkG62N6ozp0ln0EgJjJq84D20Q4MaixXtRx3cOoe9EASBPt/5lbypQV7n
ZBQzHHAHZJ/Jo+dMnvTssPiear+G+4AT2wTXieLwFhGLluac64mtmjqRdOavKA+NBGQnFRYM02PL
DFZOQJ3EgzYXStmq51TNSFof8+HdizQyxDjDAogL5uIa3AG5lJpGrJXhILHC50eFinB5fvEaw1Dn
djC3GvIoHvjPC0CL+ZqFjCBZnx3V1bUXuWhqRDYFbJUV44OZlH6JNzH/rkf/NPPMzHi6xOArZhDn
HVisHW4fMZYk8slRFwqSNL0tZF3uJxs/1oFMZVnYhbu3Z/h+33XJT3ASsQpdn3QJgYcyWM7ixn+Q
b65iLIeDv7vGgdVvCLRMRN2hhYGsKus1dnpwlpYrOL1F36mSALplpCJcMEwvR2KDkgJiWi0HEZVu
azW+c3XE+EbeWf0MmtWNfF1cXeOJOYliFm/guIHWfd48C/W9awAM2UQDZF5sUlgo7Z396o7U7RpZ
wsCt05m9TPtIrkc187cMr4HimbLJOqixRb5G9yPV8mb3EN0Lq4nk2EH7u5PCNP4gHO1oD7Hu7aw9
FKQCNSeh5CW17UXkGZZYjuUKdyy/MHW6wfQm6B1NyRJwEE5Ao0QGm4uqD+x3L9/LzFLu0RM6dKFl
cWzNE/ghEd/9fgRIfyyfTgwapQ5aMBElOI0ygzceWnLxgnJXHhVFaHJpPtZtWwZOK4Cej0x4NOxH
y2Xa71No94uaR0UtgSq9OoxmvYEMIr7z3wnkZrPm8Pnc/sy6u93ZxGD9jlrI91v3/Rd06i8yTMYc
IFJW+No81jrYlM+gI5/rCFZ6EtDF6FYAP+rQEMI38quhQhW497m61sLaN3mmNcVAP5EXSpC2VlX+
/LRtT2DO6ALDSjFZJV3HXJtQjEeVF0z9vHEcJnRy2adKTG/yC7z5pIpgDliRQ6FFjLKE44lmOy+G
LpOb+Jd9wIyhOJxSZ+uS/iKhcP0d5rxTE4Lic+qHzHw8yrAsCWn1p83ILR/+XBesxG10DKVKaMzZ
FrnMr9/vUd+sBc9NPi31HpRMrzMS8l2HHsvjIzdvNYI/jhw9wjptPwBMT+XD8ipKHfk+YYQBiQ4z
if/u0dgdOQ8QiI/CNZCesXLwNgNrCmmCTf0Eer3gTzHl0Cb7Ia2rztVLZOnbGwi84Qjww/DKNlsv
M1pNOuamfT9fsnhcUnFxqjXEcnnfzhbIMmPFeco7JsziN/N2iscICpdl7ZXTg8+tTL7lO/iMZU3R
/CGTx0/cnIfhLMpK25fXHWF3FLLMRxvQMR8CKNaHFlv7CEfvi6ORtrQXFe8Hx/Fhuu8978H5Jk1j
jT3Pm/gK1rr7lMrObX4ocTMVXwZW7T9EcS50bEwdr/CHgAB6C7UzPph+sHVmeXp0Jjg2pJGR2tcJ
p+hi+B9+qEMyUXIDp86+Ky364Bf7RbgN1asvnvKD8VYu/ijm8uHMqzwoRRmLAvz+QIu+7LWQ8Tch
02xLRkBL7mbu/ZxFv2IYC/8TO8sVDfEKsJKYVQZ/ngryq36adRJyLtwjpufjZPyq4pl5IPMW43Xs
fjJT5cY2+1iDQURcT9o1+5W4T8XZjKmiDAhSf/W2r/UNelerzihxzWa9kz0qUJ2PCjkzaQzNGdIJ
1IWybMEHCmFR8ej/VsoN5C85JDkci6kCx7OeCggBFkU9EUjId9hWUr+G0gCqsh6H1h2vc8zSrxxy
ipRTqU7wFBT8y7jiU6rmNHs6Xo7y9SRRuiPQpvEZeRMSaeaB9NDSlNO5I8M4k6hzPgje7h+gJzfO
4JMhrZciq8kBvoRp5zyCihXrKWiltPui6Nii98QOuE0N3gFbJfTDCZJ4jm4gAwoGuLK8JuTW+7+d
tqCuVu0XWV20SYNsZzC4VILBG/zg3dJpO/Ku7eiEgy4d5pGzUxN833C7bc4r/MRJmjnZlShxkCow
2WnGFhPbNI8AnO9kdc/9dQIb/JwxmJke7ojVV7SDwS6bBUuFFiqaydJFNQI8IgwUjcRcsgJ8eZ+B
w7CVmQbo3HfyO52c3vJVTsezVj0OP4lk9BdHLbtjkFYQ1as587tjO4XoavRb2buv6AENeXBUFTfT
yq4Iy8fd+6Uuss40fXagKBlfeyGpNODLSRA2JUKEaRRAP5nugMJdpme9wWocZE0ScVMpjR28n2Wu
Z8dBAuwE9j4KNFGqKq4gXsWuu+lTkk9wJ8eLq3aPjk6Xftj1taWnBZWScIOAf8KUFwPulbG8dHqd
F7+liA0fLIZuza3DeVt34d9AM7a6bSCnyOoxfmJLbdWKEcrier8K3oswVK3PRdX52pE61z2yxFNI
XUT2yiR056SbudNl6r8rmL5UdIxCiQS2KqDJ3vEK2UQhC/3sNnFa0IUVUH+2kMb6PFzezY4ZvcpO
KDX3X01sq6OiJcaW6NwwrHYojhWEt/kv2V+/zSZkAuxYAnD4fCJNCv1eR4C2NYKTa8ajzv0V0gs5
Apyb/Rd4Rzxx1+DAYVR+bwdFxG2Zr0t+pCv5p2ai5W0u2lH8YDlLvrPoXIDX4eJVIukFQs0z7iDg
1IhhfxwImwAtg9v01B004qIsA8qPR9UBvpgbE9sDWPxy3NoLUfqUvDyWyfHdf2kI21UDqr4W/CPL
0GhL/uvqaS5ZC7/fnAd4rUdUFFDgFBV0mMuuLMKmGd+vbY41ajucUyOy4b1ntEyUzqXA4/yLdsH1
kUfq2sty+Wr4Lw3vFLxiCJHJKSdzr1Wqo1Q+nHjQYwVGTx8i7g1N+Qdvgl+kr0yRKSzjGILzqDOH
zNbunlTFSVJtcqkOsbBj6XsvYrk4VEQuwlpjYi2JWWnsRnBfydHehEANvP5cZ1w2PMH9QfxtISCb
dPhh4a/TSGQFTtlUS8nK2sDuTsc9MlXqmEHpr9crjx6JAB7EjqPo+69Za0vHfRi4LRauT2wmzdxH
DvjB08Zgdaw1+mzazzP+YlN1VjPm8KfT0ByilopoDjUIOhZUVM+j7smlAljXQuQgzeQlV1o8L3x0
njOYtyxp2CR2C6Iwmqbhwytay3uLsCVFV9oI35XhH/9MgnT/StSmAdhccpWM30QrGLvM2yS29lxB
xLC5hjTzGtOfZDd1pfly/1uaMhTPiIg/NkQuUwO5wyHnbz7IejGptK+HtjGNTqqH75CI2XZOUW/N
yuOIbGY2OIBo+iozRCu1NDjBSyePWnbaYUbZwxyOBif1hIZmvSBFm9CCFp6ldR3DtbnfpVlfJSsR
UrLiNzbpY3NfmW3Pmjv+gWAo6W8FWRI2zZEdUeXFUnvL4ecu3GhYdXxb4zbUSKWr6WdRhXgJJj+z
MsF2INzYyEzeuhtJf/NvtvQt7SzDL+PC7rKS17I2gGdBomO3w+6QOtnteAGF3ofTER/Zf0xpo2ER
VewH+fgtidZ/S406Obx7wR4ElBfoJF5J9RHkDaJpb8sMJPmL2LTLvsNiJZMKw2cm9gJe3Kox7FnI
eEjtXW+1XwVsmDpCj/xZvvKywHf4xF+zdgvBqcnXp0HqiSD5EqM3z+M/CnKOATw03eZppHuaLVvo
8L3NdQtGo6fmgBmtlvFa7a8g1JPHnCZd9qNsN8SDthREA9iDjQ6d0ATL0Q7BtmcxBDtQIkHE8WoW
kTq2GcOgdAZ9oCFHKq+ofW7leqfgPKygUsq507VMO2cGB4uBgr7xLRCb+PRNTwAxXbAJ2bI1nLsE
IIdGtdECOz1klot49a52H5khZDV9qpz7wEMH+GBcziOWCjbPqBwG1fl94yL97rj4pMcSbA/AKSTM
Bt8oYTsTUjWjzxXvePWJb4GOr8bUdaF47hTE+5IKFXy2mBwTlxiHavEQZz3KRPdkzcQYHoYVnaHW
XNFTYKopAq3dF5WjFxyetS3xgksbK11bp0paqoYcILFZEiN+l5kdt27lTCJcF9juNkw+6JaWl+79
T22R4apmvObnB1YZwcxottcXqI9uCN+nTZFsQv4pZP8KoIXoW4qI//J76tEnCeHdexBgXKA+++MK
yMbnSIYukMvqLSVUebk+hayCY6aCInGtkyoGUdnoyaEgkMPfJKPUUBtRMiDYbmrMs7+PGHLW8J3+
slzfx03opFHwYjuMLbgtK8qFra7ltJn26dmc4DhB1b24N53tCd9fpqFT9XTwu0CySshF2E9x1iY6
jS2Aimekg36QA+7j9SJpmGSsfosB2XoiJmvBrdc2JoPeXjz8F6NGdrB7hkSE6LDLKamDYYO+PnmU
nUhQQIBmgOPWlZ+2bLcbyby8kl6KiVQOjBgfc7XU+sn2RBEO7U0r4BDIieSiJj9tQKQHn3SJbTSe
CDMo7hAgmSU++2q5jvNtKtljQRrviIVOVEW/7lJoOsu5aXX7p8mhFsYg7yu3qGIVsvkNUwKJTzh3
dTjPlP3P3mA3ftyuiU2ztBKFmZXdDg2/xGmT5edja0nXW2HbMJ7KBqNme9FM4cLFELAmDz20rHV2
/StSXNVa5aEXO5xa8ljFAYTF1c9R+ERBvMk7BbmfRROVWBg3jJhRgX53ho1GTpcbve1v1xQpDAR9
kAm36ja79hOC8RFjqVuZ7X9bZ4s7S66UHuP1UcWpW9FCGH1ctx+Wj8BYWxh9IujrYXsCZetTyCS4
mv9ozQFYJZYcHP3Ni+wZQN48tLz+vsAlEa2LFExLJVn9sYba1+JxVNUR2MHzNh1QDjvS+LAo57lA
bEKu9rBP7iCsFsk/HbbcluwJfwSyU55IQcxH6CEBZSBbR3z4LwiTHmpGbW0B0QZw9MPzGIq9SkLX
1/4Xs+OdJfiRTPbbRRDzGip0QI7rpmQA9uE5WJEEh74zQ5mGu1tW8OLwGvmD98QdvQcuNvyp6sVg
fEu3ZI9naERtvzvjDJuqDVhZ+cHXl3RPBlBrIqnZZLhQvNHVnzQOBwB4EH2QdtL8tZgf9Pt5GRLQ
k4Ic7zPIjg4SaDrgYRdRREUmbqtavZz0djsubgik9egsGj6P8p2X7ddC/5LVa0gr5y8H6IiRZmMC
EMLXtg3P5NbhOTJMaWDZGp4Ww8pHChe+GlLn+vX9iLhqsC3sXXu4iXuMH8ksjM+Wp4WQJ1q6E/A9
N4JpMlQwD1Z+bVsrBxNkINTxbHR1Zv+BLSgAKABWrp/0u6vvDbVRm9NP8jCjrCxTapOefAL18Q8U
V/Ydko8taOP0dTNsMbjJN8MKcc98jmsJQQC0n1qxKzXUNXJa1EigvO9XXh+XerEHhSNbOHdK/YZP
gM9JZD7/z1yyxpDcyRQ4QlWrT+VqX5UY+L5n6IsoSHfoALfbfRAYYEIQ26h9DSp0D3yJlfChlWQ9
kRPajf5io7ZTZGajWPwDV2O2piS0tt8B3aPO85Uv9zweYOVQY0IBmrldjk8uWy96jPW4AqtqQRjR
UrqRWA89V5LZL7lg5hC8nZiRmLovCdavrqQfO6PUgQ4wkVGgHwgewnZARmqsJJf9lGF7/9OC/y5s
jvHj52LSG7rg0rK0v9DHgRha7/CK9zb7T8F/J6s/ZkjxkA7PvRijURghjTKmWgnxMfHj+uITpTS0
XadeVSUjtlQk2+6kiWwux6zb/AVBvYHBD2lmJkh5BsQD/2tu1fj698WJhbqDwYjLGYKJ67OHBpeA
JDNro3lGAoOhMhOjC+xlHoHFDCSB1TLdTuM9Nj/ZclDXRBn6q0S+Ll4S6vjWRY/qSxLJ9dSPqcoo
imWC/JZ14/M7Pgc7yQGohq9JhdiTIn1p1yDinCyB/k4ohftLO11vl3Z++ftZuZ9ZxvWiTMK+bBHW
CNuokWJ4sdL50cKOs26xeUz5kCjGwRi21TD7CNe15DaebAgaYCi5Ciyu1fHUHm5eZUGbBsmd2wBD
Te1bZJOdy5wRANFTuBQ5HYj29SK1hcPx0yG7Y5+eVoACu7SVH75q7kJ4tTX5xP5NISbWwpqjQsWl
CKJ8XpdgiPGFSGf+9wdIMtxWw82WKH51YnV1iHN/sEv8KoV8yBdcobEqP/sOuj6fNG31fCjznhhF
aDJdoQPM+b7v+imkDoWCuNP5yUdq/VQSRGrXS2QHlambRxZBibJOjV622NdYbcJ5P8QYCe0QP++4
C/zO9XPr869uuwgH7GAit7lU1/SiaGK75MEsVXkosNOo7M4zj0zRLRASD3+i1B9mhSoRiNhjOQNd
DHs3JAoAQxXyNDQF0i82rY32QtXfJkAKEintiaqjvllRil8R0GAQfCr2wREAmzZntJqmJtEdJHGt
2g6IWS7tu9z8ZTmyZP97LHGnkvvkOgcCo3+mRQblzdTi2fRzPfcCWi8KpDK1Eumun22qwbTF/gpa
cUnNSmPUh/mTvXNNjlNCMfxXsDCIg3g+F9Jx57vj20eYEx7lREWS+e9763qaIMt+ot+Wt9NFkge8
UxWt82VaG+6i0z6NwZHr4OaTgiWslEC2b1jTIAfjOaHZ/JL5x2vjBMrRDefaswdfMxkyPe5dImgw
2E7ImbJ2X0AI80UJq47NouT4MIOfZWvOJtviA3TsGCCw7IXl8xVsmgXyg7P1vvHPW4xw/16419eY
h7ZYgs//RiKLAh5JC/dnpKajFwPT2mjFvHSbya9WSIeRGe6ZsYkpTSwd7AGf8qSMiew2Klbea0yk
JWlyEim5sAqGvqTUj1d6TlUhV1XC1BFeDbjwE1M1cVp9vj4UZVdH1kbAICQH5rYohECCd6+SmkoP
8AO19IeoVL6fzTuaW1TRc5MZR5RCATQHZ1WaLfcfGUDVmCOdkn9ADnWoZyDb0X/3SeZxdeTH5rmR
QYhmquUgdA6wxazkWRs1IdiiVU0Effl199SQJf0CzVn7zQc74+HGQUwKMbq3immlBzy9sTidwYwh
tK7vequIRnvjLGn64EHGFUaKzIz5IeTr1aK/fx/NTshfY6PJmNeCINGRuQII0s/xuD+goJUttaoQ
8reXkIRiIptOEUdT3IRcFrO1tZa70kKBTnw3+CcSC9+YmTxKgs6ayQQD4pnQk0a8ODPyv4GpzoHx
mcF+XCKqsDLGn6A22fnKSh9WthiF+e3XEOg+aUPZELd0LJQM5nBZWLhMQs5qzykhfcbuj9+do7kN
b0kSQh95sqd0nHzirVZ4GtPCssfw5rClfuuRA8nU+P2xDfSKtgG8o8xGNAzPYEbkEumzWAw/jlsm
dO37/I7rJzd4BMV36FDmam5NLkkN24q5Wt3up/iR0YjedZM7LzceXMkKCJLnjxMhYBgVhYm2Yudw
3xeLQZBLnB5cSPSSk3A2B/kOA180BRfAgywfZiCqmdZ5CdZIeFtyLkWxU7x7bzj2jgR7VNZLp7Lj
M2lQnpcRoeXdihP3aHVz5V5CY0i3QvrCqVFCI+y3yfVGaj7cBFilIPddQgVhdU6L2PaFwnT8veLv
RXuGbvHplYXgXuoPdTq6PMGk2bBtQzJV6qP2k9gAH7pqBzuT5TQuQ2o62sHS4U9BbMJE8e5XXccA
AdvdUAF6nyBQaLU2FfizqSNad/mQDSas10inY7j8ka9IuQPYjEh8iJbYnt/oFYNP8cBjdLInzrxF
OA9ba/6Z6ygUc2r9OF2siEdh3qSQSXQJimNIo023s+IJaXtGnuu5QP0tCx46QY3gtPXk+QT2sXME
PcXv1ANHR3egZ7trn73pAl/hnIbAh0oUUF7Z6nLSaxGT9wl5CEciUjwMMYGkOe238fZaVilODUK2
0fNVnOPe+iEGhqRG6VFVXbAq+yFgtoxzSXoBSRTA5S6s1a2DmPlgavfq5dalhOhVyTBGfPhXXkxj
1/4k+ekbaI+/p4/F+hUQdYuqKIWvTKp0aNWCe2167JtGhu0pRH66l0JDih0M2XojmxBc3jOgWPkF
7R74m8uXXNj+Mwmhu7/9rTn5IPJdzFLiurFrlMKPWPWcc2XRkas5cB8JcFpOqqnNsAETqgVc7aGU
hVDq8Kr8cTmbZ87n++QHFFgMrIg50HUkMGMeZ9zKvmCQkooW9limYdEa/fW7djm4ECmRvyoktahv
QaWV1oliZLN3gTK3Pq60eD0LvWvkM6ipuA/3m47M5Kz+Z64mfyunKh+/DnyI2WlUoMNXJJL0yLSV
yrprMRfqJaXgml4V642wK7ZFeTL94fiUBxIJ2Lx+RtidD0zrBE50BaaYiuK9aDB7qg5Zr7oiZOE1
+LFv7gF7rr9FHuT459yc4p6uK8dzXkNvUyLaIattiE/Qvf6tHI/AumtT6GXhOJ3Ajz95q46NIkKn
IKzSORW7s0dPSqc6Ov0ppPDvGaW/e50YmA9LrJszxDf+6qqhBW8x33+Tbzstc4/NUF1FRohLjxqJ
w9zqZi2s9xwQahEOI9XbfvHRzmyCQSHqWY8qGnSfX8ejMWTDPe4C9oECOS3AgFTo6MAoKHstRJCY
tyqT/0A9XP2oUEGnUsugsEN79S0CSykdh37xFkYupzZb0I8h7HwdOdN6r7MM9TKbzLVL6XYlRswF
RXx+g7rXI1d5Rv/6EG19Nzqk2/JFWyRtqV2HxthYm0QfUTfrJ1qMdmFLDl6kud94VESZbSGArXW8
EdY4AwovUYl2qRMKvk631AWWu22lGEBt5B+itGhsjPQbAfYqn6q7B/kx+r6/IOold8W847OO60+G
WGLQ8etOus+i4ZfvTgrDS3BmWLZDrN2F8qW1nV5Pxq+RM3uuPCVEkESCYe5gHA89hYv1hDu4sLsP
6hZawXsVAoao1hQQqcZQa8M80nKaW/91iFGobPLtseP9D/cfhdrZxSQFZ0vP7YOo19rFbe/Kjj4u
9oEtKetkAc7OWnNuIYyh0pW58umRNgTktxbYHDHdpPNjIPW8FgTvcQKECvJSXGMaKjylfII6o8kQ
oc48aeB5Cuu9z6h3Wzo3XnMZh8R216WsUrP89FLi8Rie+cwUX4XNKulTM5l8D9uf1Qvj5FVR/ZBX
3kr2j1tkA858iB0Fj0XMax/l0kn+gx9J7+gr1OvxQ/FtnfD/rjQLHzJF/Pb9P1/yICiUMe/E9jcU
KZSL5hllaQ4uEPMRhvwmJXfSogfpm4P2SSTFJzN+uWb5kaJ525ZUhPRpj6YY0YejiPnxg/FbXlDh
/tAr2dk5zLSlnU3pUCBtIjWyxW80kfJ5AwJYlRCPBaBSK+y1159NyaEy859hGlomLMBSooxtxd1R
ER66+cEBZhbIz7rUETgkzVqq4d8pYBQ8MdhCHkxNlOH35U/U5xFIu+z0lGBqYP7CUXkHzIBAtFN0
Ls4xlgb+fLvKeEXTGJvjPzg/rtzf4RjeZ4bpht/VII71nOs6rJllZlZx1rvN/qghA192hOUtJ9gY
a9OVdr2fDihbKbSklB2TySjE3PlTGwlo4tGotBMyRtLRLOBqz+RlBFH6bABR7Pyf0+uqzaMR1Npm
tXZVm7hQhMJ5Kg3CigcMKoku6JAWrFzIMIEDWTM7RBr7QbBQUEpY7r9zdUcw1OlnF8PUjKhn9Y2e
ZE/lrSieBB6Bg4T88euxPNn3ijutVvpZE47GqBajNgwIUKN9oknOBTnBMVHReJ+Wy4Mre9Uy0rie
0vxp3NMzU1lcFWZ+yDcD/loORaT5+ibCXvL7Vh4GIX7Ic0ng+gY1Wa+k6CGXSfq/xhRH7FZ0Mz0i
if29AWs8O+wLvEm+zOG0idLgOZo6p8QegK2P5Rs5Q0fWh4QG7RuV7C18TF3746d48fSBNgT1WAcb
oUzGLq2JFSw9VDwz0qjY7iNJE2gbNuQQnGsFnRFcxr1JPwWxPBtGOJmU/+CDBUsQ4GW6u520lA8u
zpvuqZBlNI/5ylytS4s7z0FY2dpj9pjmXRk++JZ1Sb6K6Q0awmZBxXOMDfCYoOd+FvsmoERp4a5L
AtRr69GJOLzZlOvoquPSv/jmU3/G5LNuqR6cSGt4cKpJVnwhu9FOK43I34EcZBAaOW9n+iwxYrnP
4ZzXy0PoE+xahJ+qnVxkE3VQDhVjBeo/NxEp+yp+A8wGq6JVVaMSD7uO/TpvmUtpa4wLjtIa8JE9
wS9Rut9ZRWcYFj6ciosD4fcyOvz//L0qA2svDGXSNUorgBsX82Wh1MX/8JGGoa37Dcj/UNNyl43O
gu0m//t+b5LrsnLxeXDcDL8MMFrlpuKsOHkKXExvDOmCn20jse8oBpnq+qTCdocAKFT5/F0sGBVZ
1ZMUhv8VCB1dHg+onW1pjljkuUM+shhnXYt4SWAVh9FA0zH44E0zLFP8pbxMem8W5+Sbj1pDCl7K
RjISJsuqZgVPw0B6H451MQ5yOeA8VC9ADXLrXsZTPIwMtdZjo3jysk8WJN3V144hh/oZ+UaOMnXI
GSKy/s6x8QjCke0sy2V+YAB/oTp66e2rzV0GCVTDH5v57m/27VY0fvyqqSoXvtM1tDTMQngxm9co
w8hMu4dnsaVk8WDGvBlFOhbubU/kV1rz/gsIhU9TmBbEMVpTSVKnMl0567FvDxOkuCNnF6JwvbHI
zQ6q3lDg4zYfWNR29ZO6DGm1DiRVtcm9271MrY2oBiekm8ykJiba9Zng7PUGJmOXj7H+aBEEFTbU
ux+HPBFvhqKsiGbCAD0gYZzfn6Xprggy5fuE6d0LODLRPXgFQNiYeIqaV64VnpfGlZFCNhcLhVnh
9q3w654CLllr8gnZn7qEYt1qji6dAT/1d5DfbW+JCTRepTRPgBjf/xXRCR44lTqIriiF306GMLMt
MScQbXsJ4Tdo2UCas2jVTxgvKH400AWdIFChwbyqOR1NidHdFq+TM/5z9WSR5iMMebO4aECcy/ps
RLDF6DemJ0KLhTacgqydX9Nqb19IG4GG6h0n3k0TCxM6k9/k+3/+KqNmpqM9eTBhR9WC43g9oWy+
M08A8IPM+tlSpQZyTe2bqBaUMeKfWeK+P/y+lvztreoTyy3r3Zn69exGfJ8sc1rKeCc5dMLhWNnZ
uQ3bTaSVw7seDLeie6EAjC/ICLBQA7E++IVondk+IK5CPEK10KRIAF7P9q0ivddE3eqqaLjTKcWg
nzo8wyL7cOk91yMQHJwjeJdogVgOQ/y3pIEVmA3lidJid/z8qWU6V89g841sWPcIZw6ofnFrxp4E
5s6q7G4B6xz64vc28GxuyqgARHOekXKZu9FhaTgELBQ877V1lhRXbkNfYtQBH+ZmY8NHEqWdqV0B
zIKE+ewagcvYV06Dfx2NOzj5tYBNptUGDSNcV+Zn0/KpLm1pISaDK425uJfUIkHAnGTeToL/t/um
+mxYY+BNpgyfI0wdtrpnpNvVJLWHMZcdmbbUDi3JABDvAm7Lo3YHWUR5IPo9f2cXRKxt1T8skOKB
Y42bJQ722pigP77EniRWedW4JHOZd0JnICVckI6N9OFTl55HFEcYg7edSXzZ9uNmUjhdwUrlj39M
j8bNgV4iK9js3OpoHsYnnqt3x4QZpgGLPqwqFR0WjmwFjCUGJi9L3W0mvyp0D0OlLpakuomM6YNQ
DYRG/FWZ8h1Pi3i4nI1z/LBqwMsy5C+HVUhWBYbKE5+aRnhVqtQZyy+L0fz7AgjTktDu9KUegfej
Zuuf3scYOVwfPxz1eR+lN2L7jwG2k/7TgdorJrdFpnxUUhfpYbYS7gDWP5ars8sKTfL34mJF1OIo
O7D5OLtpgOpW2ekpYIHSyuwnVAxjzvH4pmKDvp/KQkmNIGvRmT5962CIAzJ4fM1/35j6D0IDgRoY
WzDMtKAbErWG7TyOLO/vMY69w9cNwALgtdaVF1UA5SXJrEikmyLNph6tiyUiTG/hcgqJFZBSDUR2
wYzCg/sUvk7cMTvJhEENoF8IcsiVY+S96cU++9h5WBOYnMisrMs3OMqGLYjIUNBO7rm/uW+37kZm
rtdLa87lMmDQjilbNJZzc7GB7jrS7mUt0XLKXYyxqVbN3SIkZRJHDuEhLNqHohoPqeGrOdPRapjp
G95fQScovCuQDh41V8/bS1PBJqTcmBSS4GVMe5k2SaKhak75k4kKynl1se6y6PKQLZnMuP0Uh4oe
BMM3NSY4gdKTa6KTL4XOQmRROBJUAsMoctgRCcNAX2U7iJHUUGq6OFnBfsSFi5gXRRch6a+yl6Ig
4C3o54Z+lnf1vXDy/Rvlarn6UKTXszWPX0NDKCfqQL5spYOnVyqLPHyxfEVtTZuWfR3cqfR/e8So
as9UMuAi4/pSXqdB9RVV6g21n6iiAfZb8R4OBUwaJfQUlKyMheW/dg1+pMC9317Q44fJ9XlV6/EU
K9bkzDMImclVTX2lNpLwwmfj4KIJMtjhr6XVuEt6U7fAw8yhNuJnhPJ68Ly5kBPp+YRFL4AhwPIb
cyCpEXtyeScKRMUoc74hVmmNl5hHeTmjClYJlJx5Tw5a5g9aJBdhkGPx01KqG0lNpYLKY9DmOqL1
4Y87n3khFyrFQI3R2aAb7dCgqvKWFeXgSB67zldRQfvkIxlBmAQ4PJdnBSBFmcY2KlAuakLlvfXH
oMl8u1Py0giEoCqb6ztUPgkRl25Q7zoNnDi1PMBzsm5kwlbbuXiQxMMUr/CA5XaHYgsfw6Xvpw1S
unWPV4VO0bvikZJiE75SnHIpUOF+gkTetQm8NNGAFivnjBJoid1r3IzZ9XN2bgPgy2RZOlshdb8c
fL7oGe1wfAS8f644iKD83jsbXuUxC4JfKNIf3tweAN2SuBGY0iAY8/ynlrDpXpOzAlXuqzqSW7bo
RPHi068c8PnY/5wBInW7xoP4ym6oWl2W8qdH55xOoqff2YxltcjzUyYK7bGX/bPbkWGwOQNqbXsb
YZ+DJOCDFQmIB5Vffsc4DCin4YBTuCorUK41R3bxannIGl+iRTYJXHS450w3QmfQHmfRxemMr74m
1tUYtzgBkG5WX+gHvAn4TlhVTCI9mj5zXWsoQ+rDBzruKYvfmNOwRqrjzoukIbQ0r/N87KDRUOuH
uB3iz3xuv4V4dSseh9HxmO5BAS9i19V3MlxZp0UwmlX3vIezAJ7TLQJTpczSln4dFLeTJXSbAxav
Zoslbel7dUccM3z3brozwb9hda8evgBHj85oOCbxHAGdctMIRW/MwY8hQYZlgS87wYNBcwxFeaQb
lAddHZM5rBmfoHMtywaTVzVrDRLJLDInwjK0qEZGxu/3sqQSqL8lLwFlH4aoLOgBFUuftODblyXN
WqFz+07PwfDOyRRDyWu5zMuaD1/Zzr6h9CS2pnaERW6TEWpK5JwF3PRGsqNeD4jj4tzEsTO+q40y
h8OAXdcb10J1iZ28OlIqSi7M3Nmzkvfn0pxtRq4fuhaB+booTRFTY2/7eekW65OOnWPbQYBzdPUc
mhFp3kXlLlxc37/TKbpGZ5DsLeOzTWAyOwu1PkfNxwQwzBaaI97BnVHkjXJJkUakMFus93XviUpH
KQcBe2SjSgNDY7JtN5aBEME9JieudTwVEF+PYd5dvhsS26Hkr7lfJTIDbad7wYP0r/ddu+xvFhWp
eQc+oMAHQLUr13+mAqrSiHaMUQ2+Jopk9jh/0sQr1Rjz0tLkA/eFOhnPsT8Py+SrnqHUydEkHxSM
KW+7GLtJC4lsq9c0Q0aaJZYnf7Fq9cC75EHQwCoYRC4u8bF7x6nFmf9gfvW6QhD2TRnEvHpgiHc2
jCZDIRm8yd3+vrjy2lBbj7ibchlb8DS7aWOiaTwKKd0YVk74dfj8kYmaLGZVlOSqeqWin4h2LLVY
Z+iswvxnARuARt+kKRZWYkJ3R1U8PCOb2TojEcNRfJ0DlFlFQ4SwY9+4s+5shJknqdyUGqW5KZzs
MqpZZB7juZ8AVQhdhMUe9y+HmMaApqUMQ8BZQ8epZA8pb/CzLwaJb/3vpbgZVuTO8lsQ4lPpFXG3
i0btSPwIgyUc6pzyaKMCOGqdZEUdTHrkaMdEE9eotSlHBTY5c1C/uzzM8kAIJ+dvRm1SXfv6ToS3
DEvBSvGRKjQxP5rjAkKhVcz55n/cI+2SaEdeA7fnQpjkZoYAeODjg/7/ZJ/4j4QF3MwhXCHaD/Bp
B4e+V2Vec4BGAFIf4+Cu/Ziv4EQMCZWpUUOzbKN3h0AiqIwzDoIzlxwFuQZs9mpCgTg13XQfjyiq
ubKR+IZtIo9KwsJkHtZy1sxxJ8SwL1fSCygZBvjlrUm40ubNWRdxPws2CCZWYA4ElJU27fuPtS5r
JWqFVCPoqEblcEevQn8av+MKBnoOgWqJa7l6JJhXn1rWBiJtGFt23uNA+Y+wuNKPesy9fJOcbuq6
twc1xeoMa9ulnpOKG5CjQ3+OWHLaF/fAVpefXx7CrLqDtRE8ebDOB0/0v7DdcXi+G4Z4o8pHxw13
AnJIc4C/Jd2ZHcMzagNfU7aXUq6KRIG/3/j2xqZos+HJw2Hn9+pEXv3uySTIoeOzDuIpgQhRfCni
dt7y74OO1BhKyKW6Q48zPwm86QWbUNTQX7+lN4Y44ybybh0fWH1nRBLnjd9gxwj7eUSm3ogSqgK2
2ZP+1AukCQNF/qJNRM+70wiSMiGo8DEuG3ala+AMnCBgv3YHicmo5PfzgKMPdTaReT9BofqWDM4P
2DxUEE9UJeEcglaBBnEHYERZsX2nzWcjqdvSMtFzV1QFEqWlPpa6H75e+kWfshZZgOCDhTEDkUXZ
PxxNf7WmPlEUdY9soyf2MT9kO4/o6VsluHfR+mq8XkVSSYg3QPWYzRZoihJl0H5UXoKcOBJ6vtDL
w2ZiSoeRlU4osht+CGbYE/081W8EGlNTWWgSvpX7sR1A4bBXH3wS9cxd+Rr0uE3sAZ2LhLWRQz8Y
hSpVP7y3wwJO5Vl4RPOEam/K5XKnZqmfmJ5p8ii+Qea/SzFXX0aAXrmefKTrLOJRRouys+kXnMR0
3tN/W2gXO09jWRK2yXuGGVb9MOTXkoDK2/VSrk3Vx6Sn5kQAFeelPENZRL6PKcoOQxC4Jt6CtfPP
B+NQ13ig2G03gvUPigxUJ2mT5kXMCvx/9i/0x9E4AySImJ5iP7CTfHBusLSoAHD+4zytXNxXWc/p
KrnaWweptJrYHCoXzS/rmeBkyBNEBN4HvS3gTvJC7P9Vs+b82EsIiUWSKzDKwG28SVpBPq1AJCw5
NjZb5N4Gi+xNjFmeqg95H3rBy8o3n4zHUrtanBirX1sg85XFhdDE+LGmxJAujt2p7TlW9QiI9cQq
Gaws9BEyiwwic+NYn4M9/L7mFXjNbpJ8GVLWnUdp0ZHDxMQtaDvGE0xpUG3OUySE0ujJFbf5LHdL
tlgoMMciElSglXDuFmzZ4x3dzISiKNAMz1cEEr+A9I4l+DNo84l+ITw+F/NdR652dU8erYlAADjX
p8Vgmyf5KnOIa8dJyvzPOulR3pc+3uhXzCXWY6hmb9YOIUq6H/c2ifxLzqnJqlqHNEmwwoEfM6aP
tWlbOjXC03ahAYJOh0ble8Brq9hBrGtU4TLYIH5qFvKkk4hASjBKJ8KmOGynAioQaB6bkLzvrPAR
1tnhfH+cogzQbNG3w6L3SyEbdQMm4PVJwO2EZLkYMRdev8I33oAiQQflDplBGwvVlrr6OiVvEns8
L7/fNMobKKf+cWRryJJCWxrNage8kPTgGfYM+/YZfD+tPItszXvY88aEMZI2kfxsQj38jrjn88LG
5JsrOKnfmNbmhzsSwmmsv6ippZviC4I2Vk83KmQnNcQUF890FswXzMVip8LuddrszepjR25Uf8Ao
lNcdoO0L6Mak2Dux0qrIDY2bXOtSPxB0Y9F5eelK0KMRRmAIdPZ0qXqArTyvHdKZfuiMAwbYLBtI
f6jBnQ8m9IYXfhzdAcOe6Lh75dgQfvbnk8iagcMkUgZTSVuYxPQFhxHuKNvRVQWTCuD6qG+Jtt9V
HKtVH+JTXksK3kUL+96yZ8SM5EMbsBafFy26pXu5rRw5yNNyDhFP6SsxEG1qPIL2dmr1XRnSdb9A
h6svHIdjAxf/RVfWYIRzjzQ3kFNdbiQkgD9Wr+txdGaqQTf70g85C3hUTGYhEz79kx2vSwSZDht4
eLsxwVhf+4Rs4ejrJKCjirevC34P6i6gd2LgT0MZEOY38ILBFHXNdd6aqY+FRoWgErql5/+jicAr
x6Qif9aP0YHg5KI7kdzq5ITGhhWtGeBusVbzpvrN+FSH9N0RMLFMPs+IX/sh4Y44d4HjhIvwN2Wh
q77zMbOCKkBi58lfWHShOpwXyzrRTHLrnfcfOy03tWnZY/qwIgvj11jxiYjAhX2DBzBNdb6rdifq
tJZ3jzG19dvp4oQp363Bv8EC5EmmHO7Ze9NqGRne5PzYiOOR5kPEzg108dtV+WmfYl/Vnv38VzJc
0f683UqrRsxXmVgnwODgEfi0sIvWLdN+PGt1yVGfx/EgUkSsivyF+ZCuM2YvxXMlb2WVa0xhjvMz
hiME/n9Idriy+pI03KF9SdqsIyc7UeWJzg7UuLdK5ZQfSokdtxoOXMqIRPGrcJHNdnHpX5PeG/vQ
91C8QdsqIYZ+7NBpra+HtZKYShUVNWtLnvH/YSpS0Qupg5iw2zkVQTER6M2NVxNdXGEjIS28Xpk6
mmxkZoboPs4xddQ7G+5E6iSrPP1xqhbNTSl887q9evP5Ee85jfUOFfHcKsJzfuTyJoBT3ZWMJ1Se
ejW7PhcJaxeTJp6sEcSU97PRiV6XmUJjcXkJvwATsf9BYIm/Au9dlGOqhnd2TcPWf4IXVt+mTk4r
MbaPv1j6ih4grbaW7fL22uD6CbzihO/k/2x3fcmGtWPgnxCilQURnnvOCDst8jB2XQxHfRl8t/TE
mUmhEdgSeyhYxTPUKhm78J8LM4SpoxCbFHzoBQY7oD9aDdg+o0pKOFyOc3L0Q0UzaQgrg8cxjKAc
hEJKvEj8SjThf/JSibS9KFIN8rjOpq9wjYCDsZhtvXhuI2hfdQf1X22JLC2sODIkCgLbBoUzb/wv
hwspBkRhNd8hg07Th1tg6RKzBcITdGozDabmf/BCzFH9j7p1Q7YYZJCV6jQTr17SkyDWV75n/J84
fCGmyDMUyrV8P6T0xqsV+t+si6dPMK0/JPMwUZk3CYJxUc+e5dReoIPbPFe5brJSnEb0kaIAu6JL
lZRFqZmDGboQFNAqN2DE6mEBy72AmIqV8euYavPsM3dnu2IQ0j34GVuCXm/cKecgKEzqT1k7Jcui
xY1IUFicCXO3SsNJY99RUvEiwj4zww/D2VdIq8cx038rDAcA17s83DlIQsxUVBfQbKinRiwetFGn
vpy9Ck/xSLYqfUWM6I7qQzPBz7PLsFhHpYVHSFj+GVHrEY6cgZOzEBgv126BcWHuXrIVbmFjhpB1
m01YrsVcEP/k99nH/nNNO2pk+VqdS8M4sOPQ1KvLSbMMDWr0M7Nk8xfY9884JkBxNWalI2Mbbf8y
N3hWiMdSz8r07qPUtfhlBhRwLj2ZbzF3Elp91LiH3BkvrrLg4eHif8mIVD7GcY9qrsMFOzC/ugIC
7dLypMD/28E6aEfY3QOeHwg+pd00D6XVYf/GgzRHPfKktxW+C1ytNBEH8AdrUMxTeLUuFLhNWC0Q
JjxKS/dtzGCiWCjpSGvCH1moLyNHyp9774wFCgl1luo4HO/O2w7LMstqsNt47I7aRbwYCfMo4qfa
kkH7ZrlEzpfDtkJEsFnvPkk4o2GdqadVafOIapqNMDYXmZ53M0zpOQ0aGKCZvYrpF71r+vZ/J4pe
zu1JQ25ToXtVUfKz5A3P5AFoMef3QnjCcsver3sXhMoNlp+9qSiLaVTP3fp1Ascq4J9jsMW4/BYx
BHNUAnhrqqQ7fblu26YlFOmtImQEhFnLnkiftUCj+wGQpnWloXMUmS91RMme+TLrvLRZsFQvl9hd
IB5VAxopAjtie4yTDccIuXAt6mJxXJ7bWbicOY7WqUnCvJs46Lux+PT13MQxR478pGKpWK229tgp
NfdO/vdzPEWJZFT4zLYGoucqFB1F/yYMgB82BZM/mHdWX+bly+VSTQzuYqilDYG1VGIq3+GkLUA2
+aBtXhFFhCIn8MlhLPzZwGPVpaPwXrqiFRA+8Hz9R7fHByoEWd0ETS+d/wjP3KDxiQGzc3Yw6BCT
TMsg2Bpl8O5YSHIJZXY6t2RiE7MUcZU7g4Svz14D7rBGyU7OFMMO6VEZqZ+zTojAq+8gCi4/oL3l
T5Cft44ilDO9MHIYbrSV3T+1KmyaAabt0L3fsWwiK4I/KWP3w4u8JJJTh5iPHxGLUQ718Jdv6NXQ
IaCaDlPxIRYx8E3nHzmoPmqcU15ZzsK6apaPpOBtcuhnE0xYiRFXS87+XZO3S/rFM1TfBdLczbry
y6wybMns2MlYskVIZf66d4WMAdosxXXmbXoPGZmhq09nQCl0iqU9x71tJbhDIVhyJiFHVmghtERn
TRC2AZ71Hb7FxV1sl4qQWWIZ5WtQdQG9MEGNcdBRoy/ktnQoYtC0fnYOZK6HkdwBCrrGNa3otTCR
jnb6+kyWajnolgHj1hMJa9orj+GL50GVLbm9PwmVCsR0sZPva0j6IzZlFAQgWLiERgIjHXIgHnC+
ZdAD636QjB1/6NGP1EHT6VQ5fjg80eRruAVo64LnpRgEXDCfa3WpLRXFvHge0/m5vk89/2lyJo0J
IL8awe+MA77OP42c85+ivQw2vu2A2WyezPXq9Qt59dYj+XSBMJsZzgJkggL/s+7la8DEb6kgfW4g
xhJAbnzYY8eay3cwJ3e+A8to0VT0oJyViCpYCbaC/RfOX73FK5DvexrCWubkLqWW0ISfCp0VvoGD
KBeatf0ZVqJvMCq3yVSDJ/ijVvi748sogn1FLcrBk7HQU7rdI1IGYPzoAbKw3E5ubjXt+Ge/Y1e7
4sUNgmqFOJp7Y70hmbbS/YfGnVJ+4/wTSstaSXL5SOlYgFT7wUOyLno9qHoZI4bqdea9qxZnimFL
+B7eRr311vdQdqh45x3aCC8eueDg4r6eKAJ/Ybu7YJo1ymkoQhiamJMUAv9dybFGWi1oy+dLFoSi
FrurTahuAM5bIrJweSiSSdRcgj2GNgAKBUwF0i5aTMRSp2twLQCcsZCgGLr2q24hBuR5SQxQAxGR
S2w+lBPX9sQmorOFsMpPBF97bb/+ZmzjC6kJaPUj36JstLq/O5TAC++T/zEpv/tr86LT1rMBCR26
ZUXeNfdiOhSqCc18pz4BfAGcaCG3RffY3TrWYt11e+AxLS62tSbY3AqY/LVb/6aKa9M2nAEmKF7B
Pd9P55WVg0rMYjkk+95RMV+k63RYcAH+O6Mgd1AQC8XfvZHJOMzOAXqn4LnPvmdDQoT62iDQzWAz
YjQvSI9XrX89zbMxZU6FL7Q1z3n2GFcs84ue9AQMsL8S67RfWKx2chXYQc/LtcYFpwOd+XGic42/
61B6sWq70Pz10oW1AZ5Eihboy5qHI9dAYwURtzzU27h1+EJGt/1mYb14mdn0hHotafUiPiDcbFPb
QpCn821KoipwEfMU65yoa39YRKaU74KamuqVcW3n947Gq+biMsZb+9lPf9Mhb0qOI8yWfp6TcA4x
t0iZuGG3+CJfQpA+LNAgpCSAMWg/QzHmFyBKdMQDTOicfJEyxWDa6GS2OgxoHw/j+xpZq5OIzILS
bWL8m1WrZu8P6a8ZosIIgkppp3pk+f53XU5TkA1p9bFMPPTLnD1ZpC0Doezz89h3NZwZWMee1IGE
x/wwNoXGO5isWdZlFEwo0IVDJKT7G+7EJ4m9wl2CA+BrA84PQ2nxQ+/LlQSdRQjffWB5tXiAvl73
o2tEqoiSQou37/lZTCvNVYKvJ/zyNV9cmunmPSIdSy3jirGHW9wQRAy/YtBAU+APOEpyLTsVMnkB
iHMPBiFC122+ZG0s2isDioa1riqH7RFbSP3212FBGGMiuu2maCiuFbuRJjDxo1ZApaKg4J/0SOXn
9BmE34oL8Xo92wKUZ94Qr6VEvz5boYSKFxlBf0R7xnvMS5w1MKEil4BVhjxU6V4LIMaW+Jrw23E5
q/wbJNZRdX9VlEUSRVc7bYI89h1DcGgNd1+0kxcSwi9a9kcEbDdX2t7SNjNVPvScEPKQ0lgu7EXv
+DWIWeqtwpVZsoi2FM+i38I7X9Wm3Cxs491gVaDLyd3LN2saR15bAVMUGHubnLBo8/3Xn1bj8UmO
t9vUQ7uc4hIaHdyu6hMc9/w3/0qQQ086wkWi+A43t5C8duG9tFQBr/r13GyzEMvZToj4904FOoLc
EayoQ/1ajpxMSaJOjjkfRwoXjWFA9Dm66nU3Uz1ihp6+GALkDO5im3pW9EpF2opeLsprYuBjfAVR
Z9/y7x3FcDERJGwVnsPa7FXi+EEco7sJN4S/7wEUN7zuXNZpnmN1KbMoczoIwgonYiLls+N1sb3c
KSpeo3TyaPl/9fI2KNQuuFX7/ifP2jLqOk9fyQADXSRCWF6VdKPCtGodygqEc6m1IDtYlzbdadqp
yjDDC8KpR3XLns8vFuj4gBd6VWem02LY3dkMgdR0IXT62G/M71X4ajrDeBLzETQs00t7ubhMYK67
fdIebK2xC46EZukJWKPP6bpQBIi8tsKUYDdOua0Xy/YOjJZDaQB27UgnqqeJNu1MUCuOSAQFyMjx
Ne8I5mr+RS9U0nExWadM6wvNkNs8x+S2f7AoBgcAc5nUEPMoJqb5LTxi/fjPIBQn1SAScRN/DvwH
g3iUAhv3wk9YFRyiBl+Tco3WLxcLdyST8yxhCUVbkqJuMHibqemXhy/YPKA1ntpbLbbevhMyZfLM
XPiW8nMdUjrcRtvBjpS85oSfKoPDk/i7ZUhJJXl4YnKdZ7ZfDY13D5KxYakGYzsuSuZxAAXqgL83
VbvVQ04Vlxl362wW0QXzuvqiWnh0wJ/+FAXj+xIizylpRyo9qDoN8acnFZvXentxXcQztt8bo7HY
ZP6k6D5eVXJwd4PQ4AY2SZKN2uoEbrCA+ilNKKsw3MUZwso4KymyefmO4/guHpU9Xa15D2PK7IA/
ZKOzl5URLG+kBWK79hHbszKdvPntJHM/YkN89hJ5m1KSTcUVtkU2ZnWFFxJyPwQaSBW8dISrXX8v
6mrFoSmR6zpJDu0jqo11SVETwB5nITQ5hLB75CQaclKE1Ym3bANoP4HryY32D2sdvVpw+iTnZ64x
X3jXm8S+LDS0FK0Ix8of0Zusce6h2+XjUyowRLB4T9F2JWNkFi4SeP+VY3CMv98dLSSdo4anNWLi
w+9DrE0/3V0k72IWxqMN52ueeTReYGEIQsiSRKjkLRN5pc6/DxUNBqKR0Dm2b6bSAuKcnYeO3AE1
1WgUDMHDR74TMsRecfp30jlqNBXKi3iTEOoJPgGbw6NDmtAfgAghaXGH3ZQNuc9Qv6tBfiNP2V8a
tmcWudzVGLYqXoN5XT0GLGIyQCpkz3f7bqmgyp6QYdzeNzOU1ZL9a5564VV4P9S42LBZKkUAj7ZZ
tINHBpd7qhyb91Ln4boWT24mXe53xdyv9L1x+F5H6aKzvx92wOLCiPnQUKfTKu2cCjUH/AlLJebe
lgTPahxch9Vw5r7Ol2HjZOuRqcwM7PwwBwUUKmZgWKwF+xvcb1FXaPYhO2PgFLCwL6JzxEjYyWX8
f/u/AfDnuJv/M+JQnLhx6hkzLpUZugzPBlaJjiUTjmfEny9zSSUEAg9veEZKIjqULrzQw9T8isV4
aQ0HEWf6OzQ6iMSyEGPR9+4QsW2Ek/QHsuGLiBsV0JwsHVvO/z5w3ZwCxB12ETmsuB4rSAoPuS/K
jTVZUeZ6SbS16JfggXF1eUs8J0MxOLyl78FDmqLYjT+Tmmaz75vQuE/frCP5miwxIuI/Y/usu3ta
tBTIe2ev8SsKygluYvrorH1CIsJxFKI6PPc9Qa5sBp3IwhchLRT6L76hbn0yPmryknH+k4V49yCO
VBWpbBjXxc9QtY6yNbGXRttZ0GwSsmRjXskVnx9NSRkbcImFouPrXMU1ffiCyLPNNChwpEzWE7KK
OWqG009Az4U6eQyEV1IOiSiEr/yCof9uLAdC+HUT0h3xGkKKKPLJISziZMxnrF+HkDAn8VqUmvWt
y60Y74zitBsUKm4YkYu2ijVcR9H3UeVP8aNAqDj8vuaDbzjwIe3bH9eMPUNq0lkEmowaZuU65JHL
GjQna2qPElO5OsbrA/q9pzm/5ccn66O1ZRJ/GNzgkk7R40Yslc/nkPfexui5dB+nN06DyhzW9JjV
t/S5n1xbYMcjWaUJQJNYL389vOV7CgzfesCuqc+GZbAWXlUEQ55VBLVP+Z6mYOyxj29rHg1x8d3w
EwrRDGTinpeiidi2YQTJ0SHQtoodymo1Gp6oWx+jf5IqPoU+6M9qBEl85OFiS0NxAzBuUzzFmWOd
fDAf4uvBJJZMa4M9J41fGoAeM/Vkm6l/mf0L2N98UFWl6OT/phV0dgOC7BrT7ayaeIh//pU+Jd/v
RQY2lCZqBMTXApcDhU1ecANVIZ3dTQC+EKWd0ITg3sQsLl3IIYmySNWjDkntmfUnxfianmBldFo7
akI+Wpc/zHyGzr1fSe7eHhI1pF2U5uynm0PsgA0bNyJGROqHTAwtx1RbU2zY72NN6rFhM8qmh68r
PHLLcRUXx3emr7D9CbB73O3sYisi4W5V1HSe2NU8RXRV8djtZufGNS9MTjo3YFlQXqmwg5zv11Mb
hqm1ptCppYBnRMK40alq18RtDsENfjbLlhe1j9KIKtlKS/dRCrer0NeR6eK8qOx/mz21gKbe1U86
uzuPlue05mg11ffCYLpo4wcCyY3XxfAKEHIf6Q+Qf4fC9UjehNVQidou0pNno0aFw5hSIY4jDHzZ
aG2ezbm1u1VkvfJLQm50ruwPsPu6rY4cozweJZXs1RrRnP9aFyd+kTll5XqNAKlSsIqntaKf6lWz
X/WnOC2IUNcTq0ZTZm8Q5mddG4ttrnxWQroamZjwO9fzWnejRMU31SLelCeG+aX6IrTo588cq2md
5dwcvs8awqexcKRqQD160uwP1LdHoQ/Z/XRiHNfDeIaa7GHrZQzUFmbpq3jLh5H/KmOBGK2KjZAM
XFthKptm6anCcSGkFueOXBcB5nIl81MZw9bi+1f/u525uMH0m9q38XIrgnMij7vBT1IsBhBVBnSs
RC0pBUs2U2LrOlVa1sepcastid+9sEpIiEAR9BVf8ob8ob0DegJ7Xd6eqhyDy6+MZ6wnDO8GLBJ+
4YY0pybkZOYqcHK9riiogMgtnvO6LJULfnSA0ZeHujFCRF/2WS39WxtwBwqazT/i3QAwktDtP3Oe
E7EztfNSvj2MR0jSggCrkDPqxTx6srwE0Q5/cehULOZfQGtx3dPC2AQ1+GdhDsWIJZbYl7H/9tM5
Wd5c6UQqBvFUiLNFWRXynBrCo8n8lLb+Zz3I79xjys9EXVAJPUKUq3c7XQ3HBSug1+YYOG6E5B3b
l4jXeL6ve174/oVxi+UL7m1FMCjNpwbs3DZrMg89+Zt7HG+agWVp4sTYyEvtHwU5xibAm2nVWoce
28q50fRY2okiekR1W3EP6IBQZfcom4zJ9DjJkpbXKJM9hbKXfcQVeCoSkDKQD+KTCEB5mTFIxITt
hWtnTUoxHabILLh/KavQFFcaNo8fkNpdEa8i78+Y1sRsRWw4BEdyPgMYw6wNiBYI0C1PI5in0Gsr
XXpxfnuZCF9Ou0PuTr+NPkGOSKu/GPC/rJUgI/bzAJnRtesYhqrj1bIPXtukS14PZOFpjNRLBAy9
T3jLMXsX4PJRRVJAMZVRZw/9iBayDtsINMRs7/hPo/bpGJsZ05xXmQJENtZhNx/lQF1EWkmDETGy
P19ylEovYtSZ4eppzWF4cFF5gYmsyFbq/dYo59CRMMctE6JLGsnKYyBP7q7qdegVmvvx6JqAzVsg
OfqI1yJBAQovSiiXTLz7QPLD/edKQPlz0ziDMDWYFey7dTvyc0dN2/pu71suKm3sVXSaUPOHk1wY
w97bHSqB9vFaFvkA+m6j9VVD09cMY6j7daHcWA6CZO8+t6layU/8oVAQruz00qN6Fc7cuFx2LniA
B88h+Fl5YfjnpK8YSNWCa2E+ULsNBo96/JrHJKdVZjR7HNeos3w0svfN49OYPaCj67jNN6SxWX3q
RKBAuKnMxDnBxI11U3LsR7yAnw4R69fP4IfH8cSKTRULVq32hL9ocICEx8QXGmI+2be0QsLIGTkZ
ZFUvVo6I4CjpgJWjEiD2tBgucZTR0pyOMbBTrlFPwIqHoWx9ZSYLsCtfmWD312SSg7MOS36ikeDk
NVyLIgymOQQXIjFREYOjWZ0GM5QfRDBRJSJsfUqerjnYD+3D4SzFSztMnVhxdgReQF+WA3eCJZmi
2OowMIE6D7Y4ctNHLdATCQ4JXDbDlOnPiqWTxBNFEHI5lfpo6DzG9kBFL0XE1emeW5jrVfO4lKOQ
FDXf7rXyE9v1xDQrxxf7uUZ3ROLoQC6djDHjnoFbGX2+TvzEAZ8RYYIaD4HXwwjkZ3g9aw6lo79t
xwzeBoVmAksvwJFMm9lW+aEgtWPM8DZUd9EOIfL/zqbYnXaPAbafYnq0aERILUeGlweU/ATYoQfu
jBml2jVO5n8ynJRrruYv57nG3NCobJLKUPleMTHJHdr1QX7zatQ1X2TgxYRaBC6wywYDk2ULhfsS
+UmOBJvw+2Rph7sJm+R4Vh3Nd0A/XB1G3uTJIaGM2WdDPs34NnUhce2kN0tiePrwbTBI6dU8QuzL
ievPQ4bfQFZjC14g4jX7pQZ37EjDL68HFPjRRQyJDxkEp53qWtP23P/9yr1pLOoYZ7uCgZzjSuTo
ytIAUnd4e+ILDOaVIptX/Pt+DQQFDxHvVLva5UHi7KTFFQjoWKKLct59ikjqcG72qrGRVRH53Gy6
jmRDjtfeJCCU4HA22U0bOG8b3c0NIZH2XDAV50WhtA1BNIYPXyGLhTjSpPO4lIdLRunzoeHIU1+A
AfJ0WvFDYsJeqK5gcBdg+hbbgbAQCkCkVpmbtGzMThvK6zZEaXHV2wRSkLicSHQmYf5A6eYIyxN+
t53IXyJ4ZIjEVr5QIYbs+che9qZMXy5mXMUc9eB7yOctO5EB//0ebpQd1DgCa7PLxV+bv/haHQS2
wwHF6BcYw8k/CgMF5mk9OJEf67lqKBTiEERcVf/8p5CYFfB8XBacnvUttK/JDgTh3kFoOdDUBuZu
wjB63XmMgwLnRiz6bHc92QaxcSlwKu7+vqCJZFlelebpyp1Q4rXjwubonV68JODtSySVlqNeE53h
/BlVBEYnYMwm25lL4RQe1kjHBkvuWsxyfnd6Vo84HUhoul5hC8MGzHcy+/x9CFnI6v2Qi2XpiBA+
dRB8rlm47UltTD69/xnYBm/SXZYg6C8RUiumhFK+Ki/oR3m1PzSQgmvQ7PllSHFzyF2SOPB9NWiL
L4b31mohYXFDt/k1KoNmALJoDd+RD2oeYPCT2caqhN58KLMRsIcOfJnvsPGuB7tQuJB92w9daJsg
8N3dfiCIVs6zktD26dUcxd3fBNbUS139SctZlaLdpWZKTRtUEYKr01S9gdyHEzjMqSd/wl/Fmlss
sUye6u0kP0GrhF408e6Ycna5txoEIE0s5nBbVp4XCS+BOMjlhknZmcyUi5fgKWOUI+zqSr7i7xLQ
RqoQv/TqgIgDnqIIo/Gk+i7sMb4ogcc5X4Cjv4YKxK+ySLG7iaJlT2kiszKMh6aH/DQXZ0IZ+4nX
ggQkbgXfEQ+aGolxOvkw6qS6GL95LAbOvwREsIXv2TLmdp8U6f2xt2QSzzT0h8rV2B4BsCj2VKaL
iRPazfh42TfENfETx309L4T0P41/DQK1EZ8s/JZlmsbvBg1xhGQGHkachqOOs+wYdcmB75VRjnBk
2ObCBRB5EHofJmpll/GMeg4yODxSVL2VPPnCP8HV1ezixlgNhHsVpemM9xuWEu2w8VruzEBkgRA8
1ufMw+qAt+TNSpKHpUvglL8Wjl/C9ia0k87Nn+ZGYP8hQyWh9IisUA1Ch0ml2gjHgFcBFPSsiMRP
MKi74qHLSIEfw9XewfBqosrcM7CKL8gc+NYTBuXeUPeTvJDGVLZDr2MjEtbdzc1I8oBxpJPB8WgM
1C989yY2GP1q0mewBFoUmfm6gmZi05c0HqtVHKxllheU7NQ3qjrXOD0cym2Olm0C51JiXlAP2m7p
UM6y4UGEl6JMX+cLsHNZtWu82sLztlEmBiJFYS/+k+ivs0Eq/3AD+FoOdMqurG0JKKoX0N0yFGSW
VC9exYEXXZolUtsKbbVnqhWgYAfAJ383pwWrF5cppM0Z0uLVDabUseTP3uoiZs8BvT4wF1JSEz4z
TCse1oXoEMIDjIpLGJzqI2QuXDuUP+i00uvLZdd4/Vz6eX256kVUsGIV1x6HVut0D8N1xa9C4Njw
PzVkIx1OoAcWsAHsSe/2620JDDc25A9KtDFUeQOapwK+MS0g5TbCTYu3x7j+wY2R7X9Cwx8gCMRn
xz0R3j9Yiu6DOnHbwEFjRM2xjjpCbQlpvnnbzRhR+wigmWw/jTbOw7PatIAUtM/9aZKMLGRUu3HL
2DjjLr3ULN3L9nCBvlBr/DzMlkjVu/tFNzPV88idOV/91SZStMtZgMZo3HcySseDX0hy32FXeOEl
kNOa48O+27fGDaVV/3VLY1VksggAQe19MFSUX73n+hHdHuOpTaS/hQDh1wBSqIe3mbmjgtAYxSr6
cdZvZ8bD5zxJFJcrQVRUML53Tv0IM2h0NO+XXPI6lOrulp7eXveedHK4+BkrsRquEYB6s6cv8cXq
jwlpxH7MpaCuZ4ytj2TIuUs/g8ujEH6NrdrEBStSwl7BtITW0U7S1Nj1tfG2x57/MX2UIxApaaMw
X8Qarhr2p7n7eNgND3dDX746YUaah1Yi+fk0mmkE92EAmHPd2uHhpasXx/cqsC+39M7Bp/QvkvbY
c68brzSPs9N8YX+1qvju7hs7j9ciRNw2l02L8ux6SenovAxm6oEyOgh7DIM7iW5A2Jb1nQZ1b5Ql
gHfW075aaj+AN+d11/dDoXJ0ObqgfkwnnBlIVh09yE2998ZDERqoEVIaFxwtoaTf4AxkSEchxEeL
zJx8SKjR8NQpzITfJ2ZHpLRBZCZw2FgIFpdIWHh7toH7ZTXqfQdIbQFikXD6N6JXqIrVgFSor90c
Mvpli6hco+fVSDx3hdWwrAeOmum587MwefY1RhDIzk+1M4LBIB3bqRVclVtik0gafEYB21HXI/sX
KxOWXDnEKekJfPyhNrTTJaJCgxYj3qXoO1BY+0bR4z+HAlO6IREkId3P386a/rweQX0IjDE41FV3
qOHeB7zYzkIgWwkXivJBM2Rcn445CuFuLnm6FzHrt4LxbL6jla4IOvVy9Pjjz8kJ3VdEjc5ETNF6
9tuLUFIdoUmR5hy2IMt8YXErfCxuEzQsak9bFjtAwzgVXcWc/Sokv6xbg9roj4Oly37JHAda1YSB
NteZ0lmIwBSsZ+L5FX4hy9JPPfh3BCWEWzNkXuW/Uzck9mKK8ijQWM/VBIC3oI2twl8JyfLissUB
l41be6VmMh3XlIFyvVJKNtkplP0oaIF1Onb51V5bi6Q+cKqxYRPFWju5107CkgceYNfxQq//b6YS
IsvOuLqO1QIsSSaiqh3pr8RtX3vGAOw2BrpMmJZ7NiyHMwz5gcyJPIM62V5z0Ciaa3kYgtfJ6hpg
HxyzzPPbBR+VvaLz9lLixB0nHd2m182y/O9rGqRuNpoo1aOPO/KwtJomSP+8BdqVDPV60Ug/Etjo
NpiFLLs7puyzg6ISyZ4tGy/TL3fIdmqhYvkL46AVDfWIbPWvta5u+R5Vjy7GIqwMkv9YPyNxPMwk
HZcd23DiefEGMXvmfgrFjWJY947dG0jIG9QG1xLGPVovsGQRN4Z28yKn3nQykdjwQ1cfuvkpVLrp
q46i3hV0OtEm7KxZmV0Y744r2Jayh6I9R+P8FKKtZEu92jPOWeZxUf/jNWuQkSIEbexCBuik/KXV
2IJy4Lj54iawo1ZiQliWBhWdVS9PgnB4c8UT8wBUwJe36eo7KgRTS1HmY4vnQFpi7a7IYjmM4cz1
61t+nOrmavA0ckVKtIE+wa3CE0L1x4gnMSgXgEtMR9X+0Stkb1+FWzrTAQRN9hpdyCCDiA5fBhFR
g8ZQqiuqnm3ntUJRLwERTsQNe0b4pKaBE3OmMYzwwHQph3OnSRH0Vz2w4melFySTDT8NLVfkMTmR
e2YdJ9BxNvSgyyYXzlO5AKipMXc4OQ3IOsMRakFnIdNQXh0Wzp64PYkyw6yejKam+QgNFVSJXcgp
K1HiBVDw+CHQgCWJ0ciidKzJrl6tQ6cx0U8gu20N+QHmzct6yUhR060MNeZtJ4hLM+68BaBUMVwg
+IKfkrfJG9X8cTjTkix5YJv1EUrq73klrdojbs/XamwjsRwOLBxQFzdFS6KnncLkxRKpApyX4ZCU
FThMWMWUrIg27SXufenMPsqYstcvtxTri2XkbzZt9DdNk6lbnV+1WsHQK66sHeSYW86Zxk+q8nTZ
YHYILMSRaeeUCKsTwU5hmbaPdhFJ0Cz16Ds0TZuKeZmSVwQLnrViqP738RuEQ6YUFeatrv1TMPvb
19rLnkFTAU1oxlUdql1v6X39WqTebYsdG++l/F8vVPut6EgIdBBxqn5ilFLc6KGPpiCd1/R27rIR
FS+vJHp3G2ZoCoumnd6D6IY3GjQSdYUtfqGFt9fK36swrDW0x1hTqt+cZK7I3dy7VOWAmf7ujAh5
htODk6S0Vvzpb/pJLPGk+bptQV4ffrpSQzVGk9JAXUV8GPxmLZy503XMA6OIXuGJtqOxV9P7/iVh
BMJ0mLOpcM3bkPdygcA2L/BlNJrI+E0+2oq6hUR+ul6urc9BBeWXsOKWrNIxN8HvAQCTkn4sK0HJ
0lELX8N5YvtjVdAtD5tSDCw3J+Okhj+H5YzSetkSTzrGUxWdAb7TkZeX+CxPLXFvTL/VWHeWjIhW
YftVk3DctmuJjxj+OeAFgrbNMMAXKaUrYslsCvbnO7D8M2kLCJ8P2UspBuiwEmzP6Hgntd75Qi7n
aFSZKQKs1+gLwFzbIQlhwJJKRU8gXb31t2OK6PyiJG7wHAeDq9I0sv4FnWae+coCdNcNimArWOhC
NiZh9aSkbHGC/+uRJaqEPD9Olzy3zh8sgGDhS+9gbHVTy4SWAm+5JxByUGf/SGJp+YF+gDymbAgq
uW/3x0oqXhOjQz5jq+svoUQ1JDoibJbCp9r2IeKt7594WCtGfx9e+tgh2LyzdTWJaT2CIMNGqjoW
CBdJMH7susc1NPzdi5xoGtOVh7czZXqWeJ3khbp5o9E/cXkUV+itoi/NsyHtmEii9xKV69/SdO+N
mr6dFGUdO6xXWiTsqxz2NtAPz/TujQLCDz4PDeBOG/ee+wTPrjfJvMNrpR3PXOGJqsPw7P97FStU
hEoKPx3dOvKL77aFY3mZ3mExQlbPmaOfozBRXw8i/nn4S602KpHsu+AM/HAbSss2t4RIP/0+RWcO
A8TFg9wO9wB13rs371r9zJ4kQNBwJ7aHUAxL6BRjWRAt9rhelhttanK+SHOD7OmmVz9PpF8eQi8T
YQJCZGMtoU1jFuN9sKRdZOVo48taglmdPjhrVymiLY54mGoFGK9zygmtW1kidGxUXR3mLzAKEwgT
AxsIdlKXM4E+HO2afa/h5yfLYaLbH/1bdIVgrt9BDgh8N7KpGKdqlLfttIaE0zMFbfUA+gNZZZtw
FJ5OcebcA7gS/35BEkD/VV58QsHUMKJPYGES9WP2hn0koHHcE+2Vv8S+PdZSH7hDhK/4hNeLXZjr
sap/SrsTMtgh6gKLUCxN0J9ACojj/dmOz1HpaJFWJKZN3gMFljM0W3uIdl1pgxqpGcGQSHqUzJAo
CQLgSgGsyT/80aDcuk3pReSSO4UYA9msNdQ1FumEGA2rkKrew1vcHg63DP+rgrPRqOuSi0NlhBqC
dOBNNEbDpyAcIo5KMtQjybC/+4Li/K19ea5Onf1OgHFiCsmmNoV2l0y84XBxzQax81IB1qAJtKnL
UNgsRQxZ30sq0Elo2mkh3IpoWAVD7SPmFqcBhO07WoBTfh1fca84pM3AnVxRbX8296tPc5ISVSvr
fMPiIB1b86VdYXe1xbqAMj4h6Zh8so768/YY92cAP9IpUKBy9szPtTogGhR5dVfad1yEvqabOMJf
yRfUBHBF44gX0j4AqBvlq1o3HfKEe3S7iNpqi0GPPF48n2oHi6HVpWVvvQihKtDpvSx1iM7rq7AT
4WksjfxRJ2YRZVuSTctD+eTu5SJHNyod9yXkAyCa+cIrzD+BT4kjvMzIDHVplEj67a/G26HesMXJ
rRa4xiNgYYbB/Rc3QVCL/L4iqDASnhBdt1Dkq0gMnJLxPgWC59PDBbUTGHEgZYp2P/hjc0o/FXd4
1BE4Giz+BiQnwsHCnObs0BdFfhzKmoNHH6Dz6oOmMNsQu1gjEc0qMwp1yhYPAeix0trtlRnUlfsD
t28eTTZyUbRfOnPafqehIyTe15pzzDg/raaMbgyA/ueqZEWwPyOalgyFnn4GmTFmQY4jP+KTieo3
XYf25f+SQUKdmqN5rDbTbKcac/VTM/32Fgyp5DS5obG9tCQFpyAXHvL3O//TOByXCWofz1KcsAKS
7D6OST9FzCePsGsgIDFZJi7fRNteQZYhJJhQkuyQtutvk9KaVaaY7B2LnGNWLioybFusdYstvo5r
n4UUnkrN8NTjgFPMARm0tK7daRemXhNxoDxR/JJw0kVZq39UXsoXT2+WQjazy76ll1bhUcNmPSiP
BjLwZedEMSIjG+prVConO+biNn2yiatZsQzTtx5OJ9TyEqfdqPlgGIE1+D966Tia7BOv0YOD2zeu
EYJ4FIFtjrl1D+RiY/fyM09io1xN/eqkpj4w60odu4aoYfKMd1TtIaYvn9OSTpe40dW9MOoTmrIX
TSZrqMsbf8Aaom5ClP4Z/JsWr+xGfV+l7iPNXzGSScypQdfdfQnoEXa3D7XjgzOdKk5FgYYqZuye
Q22VFSmky4CT5b3xCg2Th7V4b76fY5KOoAsTvlA1sHjCrcr3WGGTcVwd8FfgZErHFTIkvv6RzDtM
Y9ZZnnDhf9kcqyk0MCd6MbbGBeFPq0we/VcQtJv3wjnDJ70wbH2jSE/MQKpCYCLj5h+HyRpJ+sJd
zXoAw/cWIqe9/YhZYk7JHTWEAQ+aMRwuauNUL5YK3cXRM/YFXnAf1tjtDJQbNN5U0Cbv2c41iEn6
N3QyP2deltfJjjQ0PcAPbZ4OWMvTKrDut6lr2Im4fPjaEXnwR7zgtlOrzaiADdVgZPEbu/U9rlCx
ehRALeOrTMbnJAxwvHbfbsTYp6a1ZrYSVofz/FYPfF8Ku908b/vkqAca+XubihDNDJsoRqZr9kh9
MNUGRfvg9adEB9APHugAFXr9MladWM/wD5vyhIwamgXX+RJR1k5SFdrqXFzJvLcLT/PHDACckJB1
CbF+Q4S+EGlc6bUB23Vt49XMirwqCYLzAo4JGQ5LjlNH75P93obOYYTIKZSSL1s0kzKWzXFdFNOl
HPg52O/6G1MIKETUwL99jzSeObFZhm+iIzvIjCtLgJDfgZ4HGEEe6TEDhfkf6V6z4wXZKeaCszi9
I/OxlG9v7F2dKC/4K/xDGieYEAc+lSSPqecuucrYlt+q+TTGj6iCRk8gCZn6ZAvtZ8uvBe6awBjZ
jpEBO/ajysA5fZVfpG4Q/l/vLC6YZZu8CQfpt6d/3krUB6jkGDLSyEoqm3t8CXj5LSov2YRX3Ihs
jatvu9ilWhMqY884e+er1gXRWnQeeghhCbtswtPQBSnhVMDrQY+dZqM0HJe47S4daoLdiftfnzVf
Z+UrqMTZ6TuxrV5oEbgd3woNcyHj/jEmF3ZlXJ0Yk4UQVs5Pe9CxK4TasJ6qwPImAmll9gGKesrn
/sNPQ9L4Hbrs7InEPV/tTm8xbQv0qC2E81+YmQAcZSiFKjaDvowUlDvRlfbAXc4BAIPv5Yk1huFs
JoeZ0rMs2eDbalGu1Su1WAR2V4AwUwSGU7pRGoBz0fr5wp3EGtjNU2DD9PzsfItNYV0g8dknuzsP
zIjTI09WGYUHRVjt/rC1bCwthTEDhrwQuN2v66pJiDYCB1UT9SsU3Z6qUYarkmqe2TIFMSqSC6Ry
UdsPRu4Lj+7UL6dt3J1qbi6hBRCxG2ePFN+CI50/u4fMAZ4gD6mBQsXbQl7oOhjYSWxRn6+QUwXm
6h6NTtWucdzm7DeGKxd+gMFzr1qZ8pq5jKQ4N8SGWdHLeEhNVKFOMvifGssv2zgLLoT9SJh4HeOA
R0yBnVguX/VEomscWebTqgpkD9wCuoGGxND8DKJ4Ehink9Re4FiQ5H2thkk/EVQ32D0ggfqIfagB
O0WLqFvigO4vQ13mGqGDronArwsaR4h5c/bXao4njxskoJ4MowTbVRdVEDqOZeqJTr9P0ezU78Wl
XM34HovVV0+hps82o9HMfSaNG4dDX9Y83cV70ZnxaCrOr843rpQaqER6ahlVBwaOp3c6SZYJVazo
oZk+Z5+m7ionLmrN/HCKx0fnYirDKpaHIr9Ei86ekUbfyc8kIEv8j9rlMePAyiqxok37vSsNiejb
CT1z8WQn7o85uRNJOAxofQXLRkwhBjiHDxM4oyW2bFKHybUURowmU/Qn19ELKPg/Ycpeb/3UsNeV
uQ6B463c+cIuTD4VxPonO4xeCbqgSpFuys3TJGWJIZ5a49Rj6DL4JvcSTsEl+FqV+4PTjfl01eSi
oZTHrm1Ew4LZIsu/ei7b0g3iWwipFr3psgpy4xGEDuRz9TIv/UscV+9HHymef5bIvQ+t04Sokg0G
CHiGbixTUUPaCVnpV5Nh7bthVfTZcvM5Rmd2P3FGsnNDk9glu8ylEWmSr7iBAT2OJcgjyOUohigI
SIbAvVWlUwlswOH39yoyEjkl2V3T5MfyBYbkwwJKamZWImVaQFa+lhGYehx6up49ldBB8X+dY7z8
gvoZFEZFEnNqLaOl1ORu3yvJDj/cAfD4JQK9U5EqshyxD5wef9e6ZMln7nfsoL3vHvNl9HvMPMfw
hYE4/+0JS6nrnCG6bfTD9LVKaFivh3uY6XnHLOCyH2THy/w+KHBcnlCUdC4me6Gh92/GnAdYOjsT
pRTbqnEagpJC8kxk7HC0t5TXCxcM3X/h6bTM+B7cD5q7AQh0f2PysTGhq6Depa+HtD87JkrpcYU6
5UEqL567CUvL04l56e8ZMSNO/Dd2yv+aTStULfcBDv7ffwjsbp3oFH415nTD+Ps+gMkI3HEhbxjD
agQfj7PGm9f5YhiJUriOwTInSo9l5rCrzwelvn+ROttm2M4V+l1tIFnNpJFWwKy4eJXZ46PzP+cF
GWRCCB2mHiOCsHJwctTex0tpuSzmZAC1s7P1WMNoafbbrT1nkVM1SGHMF+QgTPIj22NuAgN2e0bY
PY3X11y4T5D1iKH1qA3hnSQGroTs1WY5QCRpZG3OThh1Nj57Yhb3aIryvc4j0MI6/bwO6SadDl8B
aAMg/NKpwV0Tpmf0PblvcmErisOPOGpD9/guJ+sHhpWEDaUSjT+mchADOkesmxpnxIn0TMYH5icb
2stnpHN4mdCPH4xU3AhfAJoJfwxUDvB8QBAuX/mSjk4hVXCFMFleIVmyntU7wi/5NhPioipAkuky
cpcHxfVLCgt9iWPEID8sjGMolfsNDufErcIV/GUCD8TPedCgUpmBl10AtaXltoh2N5lvknEKQwaz
pKYKT0p9Vi81X+FMTnaH1ovGuDq9Zo9ulQ8I19wE9JxwWivRVgX6THlXtibloE3+6YhNUDHC71gn
fHkvEIqfIOJbiBvjGvBMCGBlC0b8XqukzPLsFV038HRpDF9DzW+WPfWvzcqaip3GHwXcinS2PNgn
67E/0CIAIFKfVhQqejL7hUzMrECl35YOf3dhxLYqIgCa8pIqkDjxADBCViM6R9u5LdljMijgiqSP
N7HGQ8mjDcC4N44C+F7m3FOSKscBBRf5bOyILXluYdWiYq0cEMbV78pnvDGPEFCWEhU+6/LtCsz0
Ifj82GOwYB2QtZ9lq0fvioMKA0XLqn3X+R/WN70Tg5j9ZnsK0tEEWCUjEfQiYtLdEfRYwo0r8sZx
DmKg+Ajx+erePVVFofw0/joGaiCMe4F5+2Lmu1sxdSocXT3+a4Rw2Zo7buSpvYzHLrmOsfy6hhKz
Ni1SfIPoZd8qoGoSq86phdBpqWCKIAALqmOTBZn5IQf6w7wuWqc6Crdl17pOGIvTblkaxppdIAKS
XkYlZi7qfEqLpls2KXhjeSczyfiQy3SkBzRmZd14k0He8Vq+BOea+FupVkKx2A72N2rvbl9cfna2
NTRyby7r4cugbekNSXV29m4zA4LnvNQYmVJeVmXWcXHOg0JpTz9sz//Q6QYJDjsdIrwngV6ob7KK
ctc/xmYOOEk0o9moKc1VvduDadNlapzTnz0TgSncHHZowyeJ5eZO8TR7wdEJJnIUKkwxHruJ/0hH
Pd2Fo2Ve9aySiMBR+A7FL5ZUwAwxPE4UXsZssL+q5e6E+AkJaQ6GdN95a+qTBIs0Oo/BR5gL2IMd
QR/GkkFItxnhByTqeLDwQDHOND4Jet5yevBouaB7S9+FkUQWNyEXddvLBdvYDeuUjrAOPpodTdfm
/RJsoInXqLSxIq2jNpLNF49+lIlAZlTM/D54xLdnvzSjTsPV0RaH1Ohycqt0lcjTtY+V15UCjvjd
iyc27R+KP/4oKtSK/j4PITjmL+EnsrhZFL5diN7Vx6paeRDTfuQOkYio10Bp/AUT4sOEYY8ii9M9
7ogtUSjucNu/LVQIkC9umcbmVG7B7h8CkFioCbm8hx2YAe8wjO2gUuXdgVkiCkbf3SqMjjVZZx7b
zDLDgwJK25vkLXLHHlwW+cOdYBAx0wkUQiZe6+3dkG2Q6qf4FidjjW+QNH2HKtJrWSbs8Gfrh9fc
SsDPAaWBc+Ss2pPpSz1JzeXROZuoC+3hVgSdJ3IRSR1Nary3r+WygHTuiS1utAaaZOyy8MFOapv+
miUP8NQEty6Y8NiSl1oqCu34FjmP+vPnqTmMs5jy4DBG3cvt8BL2L5czDgHGd/fvD9R4rtTPHi/s
pgb1Lp3lUnulfPjecZh6QxFscg1XeVuDP0Dm5RYVezpRXff0z0rQWiypBJk29N6M0hHG3ymOrcee
u63qu+iZttluuAqpFFIdvx8V0oUvEcJ3uYYcwt5NAPAMuRPGOB0Tw0DuGJT0nshoiQTIrn0fRrjn
SL9pI8TQO6MMvzuLO/+jCQj/lyh4IZEM+HTHJ2H4hfdPucidsb//vHdiZIy7g/mpJ0UnoAVftslS
hzsvXfLxPvlmVfJfO+Wgyut8zMyQTu9y5Y9sNVa9Uc8oBbiA9ustzpGcfPQ3Ibc823HeKkkOz13K
i4Ri788Q2jtEFXIMcm3+58FeSoAlzV/M7ULzidyeFWgdiVkRgwy1s2Njw13PVnmcz4bOjFnJ/M7S
jR9GGlwdKC6HTOWenkbMUn8hepjWFs4G+GxgNYZD9FA6ZDWAe/1O9azNnXQFnfCt7/40DpMp8gfz
UGlgEIs0AH6V2erW09B9bna4KvXf1rhv5YI2lgDOnJDXhJkJiZh/ihidRazlnXvLwCSsVBRXXJ6q
E2Vf/cC5MQY4jp4G2/fOgaU+HJ7FSuFHd7WA6sVZpOeZcUZDSe5HAlTwdwNcp2YFUhgaR1xLS8LI
kVtfewxWViUHft/mnzIhvxNnX3oPsGpqoDPjOlL/KYBfmEnZflulECB7SKneB0Y/KAkdrllyKVvh
vcc/k+lf4E6BiiTCegJKBWcMPP8XtnWDaeaVNBY42/UX+hrej9anUkEstrR9YNPm0tgjohpqor+j
fRXnEndSiP13h7tw3b5xiySA8ikfUcqI3onOyGN0l5zTNfXwhBZRDqKxHVAJE9v5cVUs3u7G5n3D
BZa6tB3JjC13Z2dExPR0RNdhIgbFB0vZFbKPsQ2c+LgXCgxcNobjWmaXTfWlN3mqVC0HYcOeVmpW
DgrvkeM1q8s6+jFQWJrGBtkUDqA+FC34i8Kkko7LEmXGswAStP/Of2lzIr+zp9qifh2g5iX73C0a
bPY5cnAi3q4W8mhl+tOPSy1xQjQKh3tNSmtL3cxfiieEfXWgKcz2iXII+Y4Vmnb4xZ0jbABP4zZr
F7oppiQkFqwHJLvVr2C4Tztr1dk25k4g7VxflYHD+3BJp0jfh/g0Vni6nBXw2soWMG737lMWwe3j
9n3rJ1bAPHz/CBJd7S7jllRAhjYTbVZwtuv1GCBiRLvyxxJCwlIiimfcXx5pIntV9ZsNwpBuzu5f
N80K8EiXGlLpKYMVvmj/v4j7wf1FBiy52qJYy68kgNsDu1BVQvO+0NuicukkqZ5Z9MlO6jmzewZV
T6UAmCo1rel+7p2iXmK/gnvNz1D0etDSYg3PJ03fhn/1NLGepx0FuPXMThwU/xCb5r+vJ3HsfCuM
MYl358mNeBl9HyqJ5HzxmNE254RDkaPHpkExj5YfVIyUJkBt8mvTOBX/GBKapgagRbmsTlbi6KNb
cpb5d0XJv80FWcDrDCU8qZNl1ogWxwr8acRgrIxBenJg0b61fQxoEG1UiASpoV9qll7+25mAuYz+
ujPrLzMJwfBx/dJlzqSsvINI9k9MeC0HFPZXf+Ghwc0lUl8VaS/409Lpx+IyaTatgTWA46sOAldY
P645W/p1LeByVy+plmRcgGSCGM4JnzvgM/TdFYauDkkC5+apxV1j3/Zg/XBgB8RTnzoiYuEtMmuA
i09YgmP3JD00a2SECP7c0RBd83GNLr1Cr6B2/m0SvD27sWiR96JkzftCsX2UJsy7wkTi9Vxd7rd1
hAyNpBcVQaf7ircIOmW6AsqweW80ScSEvryz2qkFZiComeAN/xybVLrjYGfpE2dH6wj0uOMFl8yY
Lp8DLpN/8ihYvl1s3b5GB0B+lMoteh+PlnzOpB0J6r0vd9x+dqAupOc+F7WZaVYW2Soo7wlum14G
TuwSf25O5r0Dycc4LzFHRiKmwPoO1e6LcHUFqti/aasVDfc1zhKpTd5kJ8JGtri4kgl7oL3d5lFK
9gdi/y3umu2igYAgt4FtBEb1G2gaGrCkWiCGXhDLJpRFlXlTtIEi22d/ZKXwAPY+DP26CC5Q/IzH
WUiiJT7XtZc6/XOu/3dbfj5FWbWDmRml9LxPQWYgMabaRo++v6s9Dzaa0EM6zY2deEf2eUyaO16B
Eqd3CoMSclntHa+Xd7zPF1msfxIzBWfC6fExSboyYbNnHZ6iAl6y7XxAP8mPGX0L3YNK343s0B3a
57uSgSg52Dv5bDWedmFO+AX89uPU2x/SoiZyBP5mfSy6liU2kTWfpu2rO5LzsbDXDd+WuVxmCKk+
AG/F5jsvQtVtfSKrupfRGU0sWD7VNrnlDY1E/e9ehZnjJO+KNHiIjMXgnu0XSfabopZvsckjbXiP
bDaHVW6puCadqVdi9kRX36+tYLyeiqvhqibWT6qakotL99LuoS4v6cn+1hkGldPpNVZj12Ste1hc
z4hFKGp4yzp7p0p0YVSbumJZUPWgU0K4fWi8DN6QmHysPnaQjArAZtRw8bUcEdHng0Z6OCAdQJbQ
mrv92nF2Mt1AOwE3kz10tcfjqJUsx5A6xD9cAIVfgsRSXFRfN9CiT1qvnge11DACyRYtYMqIiaDe
UZUocFDpZy1N8fyxomS8ugUmdlRzF7I45E0JFoCgiwLFvyXLyH1FwkmXC4VzaSCTmXt/O/klTGj4
Q9ngLSZ634/0QNQoBvyv+QyrkHR+NVdTrLqXftZf2/IQO3maluJ4/VZY3L7UR4tE9OZR/Ou9ro+H
iiz3Ffo0kK31IgObr9KDsfr9ilMI74M07g7FDZGUQoj0jC1ZhFy4aORoFEVcHAzcHvq0+/fWwXeA
z/igzvmz56zmKYuMHN1oqC6F8I8a8kQtWjx0WQnP3bJHi+9TE0KyqOdPhgiASdaxogMbchVF8Ajt
H0S5SU2GD/q+eBG7ULCpts7A3ZNLWr4NBf5ikPxZNJsm4tdA9HW7u7a8SzL2pix2br9Fr+vfFWNI
nLt/JN1IDO53jUdOidGFPON9LMHUttRN5fK+l2Oyo7ITHOHXkwiUHgF7bF7+zIa90mWHdARSftUR
zSUJN4Xn7kTHQqGP+Ui/QIjqKBAxWIuYsbrV/z4K5PvDGZg5FEbqkGrilEl+zAjw2rAwoCHXQIQs
gVl4hLkwbqKqexQSkk4wzJaZWdlZGxTejgavifpS4akg5Q2MwvZjhaAtEnf7JuryG/SSGrQCTdzI
tlRGoll3o4brppl8Iiw+UL28uPT+de5kbTNkz0lSPY51GtIwLFflYydQ2rMM1Xvo1BlB4CbM3M0y
RZOOtfuitmMegX2P0JsJR6TrLMRy8PoOR4w/EifYmoz7YiZfm+xxVVpb7euRmLGzNfPBVD9hiNC2
v2c5FgxqZZS5rJXp4glfFdOeK1o+cnCj2KIcRiZ6xjDf8AvtT53rTXuqaw/sGOgAJ2CqErVspPRH
+CpbqQKOLf6vACTIbVjesHziyHs8KMIOqlexHpYPgKTfVx6I9VsKoRJdYY65HRuanNByleUPQ1H5
i9udJnFErHwj/dIzPC83HAM/lFL2T7kuVSW1z5y3E+3O/UIdPPVLjRjxrGfyFVwljTcZOl2O/9ad
tkHg6kAwcIZCCj8OzQtQqgANjPKI++MRAuSwVhI52thHxEgbLIUrDcEtPwJI7bDzYz1lXiM+ncVF
z25uA74i7SGY3P0ljhQpSiFj7+M87cZVz4BQuzH5P0XoIPWx/6WZr3plclKTaqmLy/QmcTCd87Cz
i/enyUoqSl/F1PCdZr09bxVBgpEMslPWjFBef+6ApOvVquaDKNOSu8q09k9dggTiuRNNaP3i3NSe
SddAcHW+7qyRCUMmJnj/M08SKzNdQ+XEyCZ6kXD1m8g+1VIMOagN3a6KEZsbKUJA8c9aCza/ciZQ
vUepBxFvMpQ9vl0sPppoppU5zdkR5mmmn3Pxh9neYM2AZYJhu0wnCkXr0/A/cGLWsiasXI+ihnfq
fsh0EUN3GjaH+gofp7cT3OFNmg4ZLSAA5LeQoPggYaNYfS71MXAAqmVOzsClZaSao5Pn0zV4E8V3
IgHEr+tESp0x2WXJPMRAdXo6PFLB2e8tBTPuyjGSSPE8gr2RBBUe+aHAsxU0Ieyor8/0IVuKlIhe
GA7EL9KlrSHm1Qc/n95NoeFPYg1CWVRG1vbGICVPxaKtrH49FRtTm0GhCWPV6mHaDZ1I4kVMXFeJ
vR1dCl2InDd7g2H6YUy9chJg8N4/bz3cNT9u/L5fNNOACTYea4E2bFKiN9ODAN9SDe2SP3DgJQYq
CDHWcEeQTpOlDbCprqPsYvbGPOhnpT/xRWrSn7okLwKHnO8uKZ+oh+vUnlmy/gJQayksCzvM2ysj
Qavh0MoDZFooHtNJ1fAsfx4PbBuFNobD2r/SBQLnWuGoz+VvTxpSs0Wki9eyngVHMG0FylgTuLnP
f0rCmrVBpl04VPBapd+OG91bGdfHBkL9XVzX03iGD9FIx6R+MATTs4i/jKCwEMpI3nH7EENNaubu
ztV4IZ1hKE6W5/Bivn+B+8EE8Ob5Q0LxWOyVr7tGlXO9RytHn5zqBay5vvzJOgvdjdinN3h12EDH
jjS+XLr4Sjyl1JvQ1zkRL65fDFuel4V4cNgKEH69tYBoF4zvvhZpore8oQa6vuVO++pUrVqb7rq6
gBlHaT0Kbn3DSFMfSOFeqjEm40Vfo+Q+hnHL0Z9K8I1HTf4hRPHBQtV40Q2+K5qWkQ9vIByay9L8
SzepSLCjt1BLnyU7shc6zL9hPDFm4SfAufNY4XR0SI0uRbtA0RqhZLH0kze6SWV02a59s//NNRmE
7pwBg2pQ6BOuW89J9Q6lauLrGS8P1NgHa/AV5MmyuMgHAV/dgRmB5dOBmJCShrhqanpExx7TV66/
fWXBTHx+5jxNujWO+oi7xN9UDhqy65op1pbmRM10rERLBFBf8slxFoT0R3mZcgBy37ORb7fTRS9z
XjaeSFlZEARi2Nb4sSXTBYDLUAhwRIE/cxC8CmAoYEwxHMZka8er86zNMOwioyUfiW82C5YM6JD1
g/mqhCU74bG3TTmVT9TRlfRTDtwj/SAMyxThm0Epo49iANDO0/Q9xVdk9poGa74k5GpIDyJNa1XR
lapcXxdl9L2bmK/V17dKIpTA50Drev6j+ls5AH/0Rk+qJB2KVfUpDkkJUMSD6eQ3DdIHS2B6pz1I
zwJq1Xz5AgWmQwjcl0UL5ha5o/Z1KButgo4B0H98ZUSfmVKHjgQqS49FB2jI42eSkqR7cVDF6BH9
51ZtZUOSj8mR8Mwfrhm4YkecconX+pWMW/hUSOP5XBvhzIp2P0ZytfZjTUWOQ62lfdUjhxUveos9
Kt8IG7svmMdeGMhKdhwCGyXdXqspVVD97NdPUJyNh1Mpjvw9VMCOGcnar8NC+3XQ12HE/0pP/mLK
tsjK27ZyNj0g8T4RvLIR6Y7EZoO0CGsz5ezPIgXgSD3AyYBX1Q9uWTCPh7+lgJqIt8QxM6j1QrhJ
J+HKGPeuFFMc7XVE6rGdpLuNfBMPgxVb676KgkyMQhwFFMJdQ9cC5RjaBE+MYFYD2Y4FQVqTbCN/
gzG0hhDSGDkBCFhzSol12HuYf92OqUeTgXzrl7UXKwX3GulA6Drk2MxxBIhZrBRtTwTeyR75YlZt
VckSCZZM3ErValAsh6V/U5KSbJZo8pwUCkd83ZVl7rzwGj91kKNp1+iK4NT+OLb2N3DqBCrwCcE9
7hQ3K/eDSfn6OwQ42LuZ+7uecY2ZVaBiZAWdedhULL1PHk5/InDhTc6X7QLUgi7YJ+VH5MDx5m9c
27lvNeRa0UjG2qfVDkRGoTNx5M40ByyPhORI0xr0F7kB/tKMcnK671uWa605XjNvxThps/YljnMC
x9sO66P+PmArh9DQQao74a9y8oyy6F6lXIn6NSy99+LnWxwJ8lER9Ko5+PhvYQSDPhYz/N0RWIwC
htRVqm5lBBNikMHVvVCY+s1Al6lmTr0d0dRU9E1kFsioQCbjGvd+KSjgwhn1ureQB6h7k5yFXKi2
7t1Dvh0iwBojQbV9BInlh9/0GjIw1TEpYoCoeZHdYPOZfMr9Bba/qdZ8g3FhGec95EfhweqBlmHM
fe/9d86GarBvicRU5g6GGO8pqAYQyiqks2IPIsiKsaRhK4/h+U62f3hG+6qJvl7QKvU8TB1AKrP9
OuMChFKX41LgDwi2xrWxtfoPWYPAsVTFnDuH6DfY8UtRPCFzrMEUMXRbL2i6oYW0DeNwd7YyLBX2
PIA2GabduJ5RbzBMYXOZhxJExHxAiedWG8w9B/GO2hmyQ3SwW+RDoMjp2ZbElN+AydJyUyRyGF3+
kTn/76QD8XXECi63J9p4VTMtVuqTM76NvJ2qi4h2V5arNIr+/5mNsGyWU0WyWWeA3te083sEPY9u
gIBkkVThJgAXeRyH6fye/KzasmvNUtgXcatjnxZit/4z0Kk5r6zMpl2zlUMLV2eSHdog70yO3PDh
mHB6sgEMRfszxnT8cPWXCT/TZTUY1w8TW/A4R0FXUVMsxikQlRY3fnvJm00QmBAn5I8JvI1YWc2+
kS+hIOXYSGCvc4YqS5OUUSiXv7Xm+Lw0JaUjK2M5zFnHde+V/NZCtGrfxDUFuYuApoVOKJnCd/t4
RwcD0o/eGYy+IegZequKOhtRBXMTr1pc2u4FJEdsyjwG7uemXtaRmI0Cm9ToKFuEztoR6eSOgy72
HvxYPhO+wmMoCNIpKb5cVawxasLcYGe4mnZ5u3s/lzdbUXuMt1W9DXSA4RuzZeL5HcQ0CahrtvZ9
OHrdXt//bYAsn+N063WjuaWW049JNe/h00kSCKNGVYXmzjNeQ67J7+bWdd1i3ph5Oix2FPRb3lIj
WcSDm9pcS3dFrSVoVFWHTQVR5MgbOqMgoC7Ktg2O4luYQf0/g/PnrBknRgcHooYmhrHz0hyBcKGn
Erv+WP/SHTzRnbyULKyF8jz3FLsMDHWubFvoJ0q++h+Uwtf94tyYlnhy05ucZLUMMlKrzk0O35Lo
5xOK3x96qMifzrSFop0bikG4qdYS7ot+Jhuhb5Z1U3BS8b/sRADM2w5x3YDOoIWbb29+0czBfr33
iAmoHcejYPZiXZF+bfA8gc08TLuAQPghJGgrHuQYA8NVc0UgR1GLuJjp47DrvLcz9nm1RjgZ6qk4
E+kql7QsnhYWoYihkrodSDqPpzZOIdWkgFUa9ieV0UBDtIm7RX85e050AucgQZ9qOl1LZuGnfatZ
oT+HpZYMItRMFm++TJVFSSG7g8xI/hcsvR92ErNf6jOzJZYiQ+lHzB2WqjQxZt8dP7TLKAID0daL
YAy6WWruEq8+aeFXcDzCkXU68taAJLh2LB1k+mSb2PSAV8mRddqURwcqwnKsOJSUu0l5TdNZy1+Y
j8FVgh8ScOi2pWZBLd3fSYZvc2yN8y347rslQX/YqrU/IcErTuW5aSxOqjShRolKPN2wqUh6a+an
lzR4nyT0gVlhMIW5DAKFEgfTh9dMzNEPdkr4SqXamhaPx0RZg7KA0rDz0CqLVbZD6gwWw81d4WBp
kz1Dol6AdZfd6w6cQaf1GrUWShtpKNIFbWVeQP30s1JpuAyrQMAO/+g50UxQx5I+kIE5lYhlYP7m
ID/NtyeXfu4zNJwp4M0cC03dyZrfBzqmVt6f/knIdWiPTBDJg7dgttC5sMXU6UIhdbRkmGrEDU0n
segHnUsgKb6Evka3D4fp1qYJYoRPvX7xzc9k/r+CXgQT+otVInDZI4hsXylU0DqdWV4CUxx1KGTp
98uCyKVy4+fO7bhgylWOHAtrHMfXZ2Bqg4Wcb+udx7aXfoCo9rGHBc2j9xxWLBpI9HRA9UX/vj1R
6FHnOEMmnYvDd7/BNo0rufYkkswUjbY+D/ZukltihCK+j5iDvXLTa+19IdF8MqXmEM+p0fl5m/U+
jbFSy6G5jbqGy/pq066m3nVN3xVRD6fkygFjG8+qLVMa2VGJeH1Ip2hF5KuaxSwwsGI870XJ9efC
ATlPCWaEMMirPQkc4rm7CQSG5LEuHTZg95VI4XGI5czbGfNN9mvJGq/Q2iozkj8mUPl2qYO3RzU1
9ddgOADw51c+gFsDUDtXBf+UC+4UAiXkD311zvr/pQsO6HPg30esl3lCCWJjDMB/tQI4GwoZkL2a
1LEoG8mVG/5Go9BteWZQLFJn0MFk4FReHYf0JUdPKrYkZuJ0EoLTDB3VLgQr1TU3pR8nf6L6ceJ4
WOJ1AZTVM2Lq+9UgnIwNbH9gbLgUXy/uKAwnZEY7WnZLGQI9BYa4xu/pAt/zqJQ66ax/AcFn1sfM
NOOi5CSiRH4OPe8ACbECQejBoCXc3ecHJhBcUqejmxc+8abY3y17Mj/bjjT1win7WDKGONOVDXGz
8oEwL7yklQPZpbidblqJXUPNXtLRIup+p7i7BzPYmMSbDdLywh6upXf0BsBPNHwZqQ3W3TRN2DxA
jkZmkDTyH4cPUs4U+t82C/yZNMsE6aOgyqoh6vP5gnHB7QrywZGu5SyPaIl0y3ASg0pCll4iXfEG
SoULRmJetY4qm48avWb7nIMDQDGaIt0xjUPTHxUte3Ph55hL0M0EQylAxIw6wQ1YobWiwbOAFYwm
qhn4EKQYJR6vAsoaXKF1VjnHEf8llXqYtuQt6WDlsbTb51p5/6+F2i5FNLXkQnMEvv6MYnbGMKWX
rHOZ6ScCm5kI5azSNu+xNjZgH+Odcegl7briiMstZQPECxjEij6fHMB5zCYyII2pfmzkAcSDEWM7
yU8hDuHgRsbJabqJO3dUr3grtK8P6S+FVomIjNRcBvenO1atdYEmo8q8HkcHuup8fZCdBu5uVvMa
JB9f7JUA8GG1Lk1XzJAq//nsrHkV4R6v9A1Rj3v9QFuYZxfma0jav5uPUWo0iN9Je4z6iHTJ8WWp
X1zxGRCLCCTXLkrdHvsZ7ZMDVgMDMWUXI4FWFMZDW/YE+3PNRgwq28UGGCW6XUjNzqOpQo3zvD4m
zKg61o+I8cB1DLzMQdMydQFmEUzDkK8lFOrpSTGLfAVa4ENJcgoKqyimZ0Z6VRGgjUa8crmhoJj1
/rnjmHfbMJAqs5oa7SzkgdiokFcp2CtPaJMd2KkM/XRIwdlBVOpAi3wL5x/H2b7ng995mZRATLWo
5DvnnXn2KqKRBkFqAhhF7b6CrnBpO52AOpv+o16HEnqTPFeCyVwV6Dz5va5mJzy3NK9ROo9jWw/O
qSlr4uqAjo5ET4rzyWgty/G2VHMgpp5x72XxE7l9o77p0/bm7JQaOUcn2Kt8Qiei1QpFhy7Zhoy4
kWMux//3WOW5uhoWqeXpVrHOfLZ798si+Eg8TWmzwlEslXP3EGpkV0lesBPEDcSCYZum4CrFjhuE
RQQ5HGls5mc4XaTbTp4Wt8PRhdvYJUcdwVhN1vbNVqhZZ1dljnRgwH7J3JKwBKSoLT29gb7eIKVP
a4q4DskHl8ZPfqE+hitrUmpC5/+sNPluxDswIBnXlQbsjMPrtWqC4evdK4UziQWbefZQr9i7EaR7
Ax5sC1OiSJT86F7euiqeZA9HHuQK/hJadJ/IBE5cBaTPY/TvZMfcBadzkCy2upszwmFF9Ou+GUKh
UOc+e66et/CsqRUmkkn+L6fJP4wtZKy4meARc2mPTBIbMHF9dSfJ4xLXmFTZvIeB8ucKMocPtH0d
Ps0ssHHJsje70nl3FI7L5U0ypMrCYyrKmyvWWbzU9FcG8s6wSSQCcLygKknTFczuT8/HOkyk4nxg
XP8DbfV66rE8helQdzbpoNFI3tk9GM2BrbSuk8Nv2Tu6EuJIQU4QQQBKI3/3vW7oMG6XWXHagwm7
2r0iPaQk1DXA1MFJpt7xxjkTVos02xPyUJtfPskLvtZ0tyyOOD1R2WuTbH8UxOsNGK42DbeL3EBw
6clOSd/QLU3qZWe+rAzAVrYE/RBPGGgd/LGsnrvgG+RFnylf88Q5LQdNgCTi9Isdvt36qmbtPJqN
WCvjP3DuP7Z2h7mevnjFCPTOZsHMK8B0AK1h8jkGTj+j9UnxawMs+CdRX23wARqBvJ0D7RKHMQNR
frqr+CDfD4q2XZyoA1jxgXO9txs0YUUStgsxftjqp8bOuqeMFtvsMg/wAQThuxL7UPFiBp3e+pj/
jj026xYhtbcbAGjPkSv8zeLUzD8obGaGDGE6A8uaWCmd+XH1e/wAWp/xaNLNF1DdNU7sQUwYBTEL
hQqlncTNq2nVZtW9jfUzYWQ2+YpAMcDlvr+MF5gluXO8dfU/+NecW4mnv1h6vSI13UTZH/NGeBpR
k+fPJM3Z+yxPaDmMCZre7n39Hl2lYBWfkPUuozpeeLAcg8nM/M0bUN2R33UQhUBrDAzweJGdNeWU
CpLHtGLv1gM4ZOkDjtSb+LfL2qEMg5u2OYjtggGeGAXOjJPPKoISq+2CrNn+5HF0qWb6WeTATfbV
ztp5CcDoYFfw1xs7gAtgLCdv0cs9SKt9SBeQ8L2cCijAwlJvt2v0qTKsXo8ZnvbslklOVdYFxESu
JO1xInVxzO65+edzjzmb5/h9An9HC1FOQeP4qXoGD09DZLNCtLN81lJ/QIuKwND+5Zskqgfibglg
/07ZtR5SC0xEvrJ3EkOUTe5IshdqMlweC1AyfPDd2FaCE6pTWjigSxUYh/e2GbPkdQ2XL09cZGgg
U2KSUD1lANSZdnBz7Gi2tOgxaWwN0r3QnzJFGo1wCvLWJkg6/sOsDzW6Li4F13vWzUojf5HIxUJS
yqezmku9z9lFzd7V4GkumjUUqwFtAFaiLE1daWGGeBIUohG8wlF3Ejkl7o1uPKrrAhFxmYmxdb/g
TXUPu9bkPW5+FH0Hdg8XGzHmTB1KOa9NRsD5Hx+rKB88iFOU2oksyWNFgCd7yfKfojqLrflhvU4R
7ngMBzKk2ZQ3UodIi36czDdErhGHFkiebxFG+kgGTRtwpb8dfhZcvLCAD6lIfzx7rd6Bj6VcYrrg
UXsATnNbzWFckgI2ftih7LNIMU0aDsi3JsceKN8Y4kVN8pcZuqSmgZk39xJdgbkpmdNzW1D9QPJb
vTF4YpIiNJsAAL0v9LZcT16DDbhcbGskIyV4vb3Pnf7Df2ym0CRzvbCQGEnh60+bKJ8gFIc8Z+HF
oBaYxoHX9bEnfBQ8Y+H8rHZFwGVsZNqC1wsE/H6tpWEqgL2pMSoVJJwpoPtSHZnevR3ODdkgFBKi
m13emhToOJDBiKmqT/uki1nEMgT4k7S+i8FmOfpwO5FPc81Ohp7k3Kcja8VbzCou9YSroAN2JNyX
dVjhKtiNG8TY0lYSCeBtVOuIc5rTySae2VlBlAmVaC9nFJvKoOm3OKE4Nehid8y/z8tLW5sdyGju
CN9nM/pd4gzYuI693yKX9ItNUN7pyGwN/rRZxJYDNxOgKYAdmh5KlSISu0YVSJJHY3HB49WQqYAW
fR5HATRH+0KFmBVb/fIzCD/uyH/T5xZmrOn9m5QpI7enP8YLLPliZpSg1czRwiwuTb10hYgyVWAO
kf8qwbQYmnrk8SuhSdknfz4qAOSCmKoYzrxzT2BNjqSer9Du/c+daXf22fad9hiflXaW6l7BEEFS
JHk8JukHXVIiRDZqBeXQv/JZUyiP6WgnRGdNzf5WulLkVn+7s6p4yDlycL44Rzx8cgt9oh7u+ldz
oCU8FBiFfQb7Kepece7ia6c7a+GpAFdGRPzq/cF94wSGvy3qsYTGeNWtsq4n0zlND54Z9Vu2PmFU
Mvmz0jzG+hRKq7WfsmZfFePw5RKfa4grqAMdr2kS20v5QcMWZUysYWxkS7J6naE45J7F8lwYG3ag
ruxRsaVFZR0Ps9hYbwfyCcrofKI3AB3/KTLEd8OYJwxSSrPTGVj7DYSRw3MUC4QY7A/e6K4y4RM7
gp+81gpnzUFavK+49JRHJDVLJMOCx3WcS39w+a6g00fFGNmbKePRbQxpbyjTFmQwXP9pAXi8uK2g
BPjSSfa42YWuzfp5V8RSgc1he9wMkDJd+QhVzFSSbAw044S/4LP0TPq4St93+8My7Yuefu4EAqSG
iq3mcoFEPxBqRFRNofGDEdjqxwXQJvOST60GQ3VdAc2QphcY9r+YJ/OdxeBtkYtUqKiC3gW04crY
RdKipDWmoPhBJkY5rf2VHtWiZpc0iSb+6cEw66Ps4vtfEFIMXnSnfC3Yjy1nBExQBXBeAEIylAfT
dbdK+ya7czyWMMAO8E99nxkNtE/Q2TRLgk8yXVdh/pBi4Y9skfe1M9k+O4aT2SmqyF192h1VoKlM
gSc4zmuFNZqq4S2MCa9c6u4q7ehUJrtmbuGJ7i300iZdoL1yvkv/HpF07T9unT5MMgTqGSbGN/Nt
kwYQgHn7gSwBARgfdl5S6LxjuUFPE43lgW0Nk/XtwhfQmjJPglEq9trG+upvAaZSGeKsfKh7b2ZG
IZjYDoYKfTgSg3pC1SoCTqtm6dKaZDrFXoUD8FJgWr8usAgvCBcPWFWIzfIyVyT7yEd3w2UvQCNE
ZYzHTzoSJZD0nPL8ctdDItQRDUaFu3ffegdMacaiaE9MVuwpcPcgLajaNqEiyA877clYLkz7oSRj
v6f4bClTSb24ODpnDrGZ61VCtp8ugbk0Cj64qj/gjdhpl1kNQPALZih2kyGrgZKMYFO/YN3vyF9y
mGpRrx5UAUowF5+hpVdJ67xSAlwTeVAsMQMNLCHkptMpGTpZ8dou65BcNm7lMR2OrurJdIREeurT
nTycaZtaVJQWjyFQkOXamXiTntcBWsBGQ0LYP2Y4cyzgAnmDPrmK55JkHKScSsCQnqW3UAE3kWoG
rP5lDZA2BFCAjwmvjZ9qbSwjVp6kMSqWB52xVW2wqyclMPS//VA6E8Rgj6cAQOFRet/sm6Ka82Rm
ulUHDzNdt8fFlYUnjjO+fcTOfi3uEQUmnv16YvVTMBfMEQWuCCABwIxy+mCH7Zbyaym5Y3mYQTOU
s4TPFa77/HeYHtXoqV2hJHqC7j6OTWhMmkXiBMSfvgToN29Ie9T3ALF9gFG4IKs4LhjfdfdUrj0R
5pcYFX2zxDXrBkVrOYSviDfaZK0rZ7At8CtQMpzssY6F5YLcMms+4OnEwgeWZxSf8TxE0jZ1zdRF
cxGSMlKyiwchavo5aBKDJlAaLPhcqHhi+TfB0rcSdXYhRywcGs+pLPPLPxNK/dwZLRXjbepppZwC
bxCSXhmXVKYXNR6Y9oa7YmoPqYkH2KuHe+EcrqebCDkj7aIcJYVo6hOr1q2//E166zZ8rHKhBQJ6
j6avALeJTtFZbbB7qiR6xnGwnBuFAL08HqA72iyFyDsW4JS3dKHubr1WRAeuiF4xTSMEExlPLjJt
qTeVYr8n/vSfF7S1Guj58XfISTK5piS3/bfNmCkS9qNg8J0clIJj8f+6qrzRhihHecXMFBR+Plte
1FR3N8Q6M2T42Gjv1owo+U33dsO5k1OK1w7/+0AuPgH0iY7Oc5huPgdeQGPbFb0zmidCK7eAo08V
42IuXm3Kn2i60fajrWQiECF9/k3jqrd3h3HNgSplzhWO2rwiU1jruSYY9EHCe7o3tVvZAPrkus4G
KKtU1QNh0ZUOiM/eYpNPamL07mOEjnarimddonZqs0BdhHrupCOGP/c5rgQCn694dEZmgupGRXO/
Hj7ip6LaIqTHWVi88K+eFhk9M2E57ZZyWUQvjuTb9sZew8JKKcC2/eozPI0m/mzLV95J+LZvmlgV
khlRbx5jtGJmcU36HBQOVXziF1HFnjsz7ZVnwIvYn3uRe7fhagJ1BBGt+oLGaLVx4s8GLRxGtRzc
eD5th1uEYbLNlqECsulH29mxekQ+4fNVf7+MfVkQXqxzNx6vsn+tghoI7+w22vYzjLa3HyrV1bB7
knhl0ZeYRAYMT1Dao0o6TvRJOuDxmH73QqIJJSo1id/+qB+Y7kD3IM1mpD6QvJ/F2mmZNz7lGYuE
RR3JZ0K8C61K/ymVpk89pdTmRpfrFZ4sKwU1eaqY9SuDaiR9r/cGSXNfMwEmd5OmstqM5QyjJOBM
aPPmBwJIxdNTFj55sc0HmDQ27HDt4QWDkDyeIqZKMW84xuHsA9wAcM4j7mPXyRxYBDtI48HL/Aik
TRc2ntTX8FQKa6CAV0P5K1Ukdk4vE10BSQGyrQeSZsJ5i4KcGswHcoSwzMCr1p8znkJgVeD19W5k
ccA3MPEsbPVllRkbtD4bIaYPygrkjEQhkqZlxxzpIETAnGYPdG/wXeQyNqH0vlSPea/GoDzG2tsx
SrzUubQ1KT1NsMEE6EW92w94drx5TTlAaHQAGJCb05GFhOtNAmQIvH1Q2S1mc9ZEcrxXFZry9btt
S0NgOE4M80D7wOaKWwb3v0w064lAGPgnG1PzzJms+aLZbdS2EBa01ZV9S6wsfOeUuEwYLg+O1Yzh
oJHdsP2JGknN8rBKU0tSB5RgCPOaf8hSp+6960K/c3T64RoQINOSKaSMX/9PYrZBViYuCiCqPHOQ
Lux+uf6p0YYS/99vD6s3KK9vbrcb45Ezo6mBi093s+UkUdQS3fJhL9faZ5C6WAikzo/1oFWOwskx
IyWc3m3Px9rHKfTtVOMAh03WO09QuPSMzqfg2W2gtkVMZr0ZXkTwj8ZqnNTZ5J5WQQ1hqF8TK1Y6
PupFm4SRhO0RHAO4Hodo8K7L/B9kmU62H7xvVvfcq9AnmXiT/oQJdLRU0MmisVeb6S9j5mMrYO56
U9XYmrgBWWen/ur4dZyBOIK+6yXMdm7S+udE4iYllj0dVK9AgwTGnIYiqvs9QXQgxkg6xfbIuHDl
NJBfdcGEoZaXpF6gJ/5zaS+o3JRjZisjHH59/3IVT6kLzyMtqsB1o+13ADfD2FEtRF4Cjv2EVxWe
ySUshXivQwaeO65B0QP5SS/iLFcZ5TzSddXXKK7dfE22xAm+Bh3oG/fVVoXfsSxCsrXpF9b4ReTv
ahO0ve/6a5MCchlh3/Bd8CiqApUGnngfYpIdsxYIG0VpdJCPOM5VTLEAo9evlxwXYfOEgTUFhwIM
z13xm5B5ez7YoMIhuguT6whrWIg4hjQhytDgRaCLIUgU+aDfBUoJgTfBNHaLmMkYdcxZkDyQ0HkN
SBmiThlIzqwjqVi31tbywfV3Mkqva0YmtjRe0g9DacsXlOXThNVo8pPcRKhAntRIA8pMG3UwcTUK
wuls2yTZBgywvHzQKk53CmNGWDVpFS5JfE0tKAWxXFOyEmYKU4O2AjyssNICdkSuJsNqPMsvz+6F
uHyhaPKKMxGGfOGNxL6ENz3Zbc9beIpJesJFY3j5TT8tSGnh0G3ruanXBOGnwzAGv56ZHIlSPnnD
q1kdmdPx8365c0i7grrYRWPlsy8OsnF8kNdbrq6w4RWEtLiY+cfJgMZFIvEhY+nwbxsVfSbWTR+c
lkOa5/gWG01302cEQrMo4He/QoGUiwNHuYKv2Hrde0XOH6xhTQkzBAPENEkHNHht1AprJWDDRNSr
406Q8LcFnXs2t7wbrurennqA74cTkhnPMYQLmUzssTyFaJSIZTaXuToJJGfkL8kZY1PievnrfuY3
Ecjy2W4xJ/Cyh4JIDDQz4uNDqx26yKf3pXEC+XfAYquylhqxRmY6NUSI2pVV9b3eBjUjJGXlzizf
ltNRwGgmACitCyzgizWGoXw0sL2lul9HKXYMbaLN86mb2Yd3DzOGGzqNSpVfO/gdlExV8zFmApGe
ikfxMcl9GZcZDjGKvsSgGcu0nE/4ODGjyMePcA4BspfnGURWnTHpVdOx207y+P/zBtg6fsL0QZzv
+oZJKlBkpKSzorgEhpu8H37YF5Ql0Eelhu8oeZsxxXVOFJiaNZQGSAskGQO9XG07/l7GZNEWrkUv
gHoWlq9qE9miV7RKbmEKdaEnfvUf+qraCxvTTGQGca9t1eZCXBJV51PXkvlC1k4wmdLaLsWJ/ZKk
W/mJMPf84X39rIYp1P2nXdTT34f3HXetJgxLpPMBXTwcSPu2c9QvUz1Xb4HA/VExVtR6VZ7XWfoP
/N6+Z6960m3Wzfcw+vupzWyvXACVa4taBtnVjRwGdAIqrxBzv3iG+o6M+xrkwIXIPLs/ujZT7lb1
vKd3lvF3h7/6GHxe4zqyJPAejhUkMZ3VXFGWMoxcZ4fb3uiQfMXrJthgR0s7/oIO/LqvMsUmZKYi
GfTVcwz1sunYAhkpwFpuLpkRYOgVu4Udt3vF1YWHvI1OPiG/7e5/wjB8XRCl2s/0/mENTtu4CMzo
anWRB/p9YOiebzxSmeGtMM+WZ7XtfODBriG+sABdUAcshGoTtCNTy+h8Ub8i3XETCUFINkpEQPuJ
sSmnxlFj2Ikp97ZBatSHAkeGevtqMQzy9mja8xBJ/ZssVa/x/PfC+KtheY+ZXB+nakbTtxG1RtHZ
PFMOsEIFxpRbj4pX2iEF1jP/iG6ZeZuDK9ISXIFb8ihYM9eborOFpG46qnOczeuECBSsPb7okPfy
fumrmx+3+8sS5uQYckCCJtecmzspU1m78yIGVy/Uu/rd7E2esDWrOmbbzkq2TWR/BkSoRKRFR3T+
uuaRu8UMNpuvd8y64u6SPpqD5EeYigvsF2Mh1APdlKP5A3hWZeIiPx2+7fofbHUt091TeLHw+OmG
SDK0k4w+zFNM+buHsOllQbIackr34TCx6Gcq1bc62Of4Fgj52p0lTKnm7BABAOrMpQbJ91aivcNk
Z5p1RhPUYtC+O9UW3vqpFVe3jEFC4EkOxzQngAEFJEI06qB+uVSnpjivXcyIT2RBPPrGPVwUSRrq
0pV34tm4TJEXZ8Le5ezOAy+YIL+WUQxxinhklYW6pznCuv7W5PIOIeZ8hRumesVW6rpr2buFWVHF
nN7pewCBQcdmzYxKhQrrMCVvV9o9y3T9n+O1jaCN8XhHXVNbRpSqb66EhdA01aQn9B0FvHTdVx8u
ka+1ACj40lw/JRvl7hRb6AXdfoCRkhNMvKU9HkBpLaaa9inu4iOS7jMrxVfYZUVRGY8mIXmLspVW
QPAQkMPw6PIWqaajsYONg+jSOP29m+TtTFy50UqbJWEB3rV8lmTnoPDoL6KU8CYlw7sQ3pKC61gh
wfzpKNBVtZcY2nWPRLmTaC5ojuMj/Hc5fvfN1qPivW5kB88xRl+X9g75PFlqSKJQVJ60kdxHyNi8
/12vv+6rx8UEL+L3QYT7hO8TWp713A4bYXEO3R3c7Htpa7tbyJuEjmAkAFqlZHXZYJubcAm6cXPi
bdAjOL0BrEY6F4UkJhWwnUZJUddneTQZdZyJKBUog1W8dwRUrBtjZ4ODEoNu791D6xdiFmyfKgf6
+Or1sFUq1w5XSTKf3MCuwqs6Sr7tZKRirLQe57qAupdBZLo7z+6lS9t6zIzlqJVRMwOCWXQ0i0hx
EMpXSsCgeqorPS84fgmB3mehXvlRqvVGSRUQfMxkukbbZo1F3ighnNXlNuRd8gBvh1AzQ35FHuCs
1OX1TlYTWFzo8bPQ5x5LuFeDVai484hWqgap2S4BCvjGqpI8zj6zvS8l1TmmwfvEEKNtXp/DwZ2p
WrHGUca+fT3pU9dUscnuoiF3uc4+pKUtt5SoA9Scutmu9e8ks7bfa+Aqq2l9lUHGOQD0FtBsaL57
Fb0hmArTbdHDlr7zSxuLBMm9OGzTr9zk9Te0/ILUqlOaLwMYNAYdzhkh3Uk2uKq6HN68R2y0dQ0z
fXGhpFnyw4Bqk4B1PGUdpawrz0Kkid1X3NTm/P/M5UmaZq/ahh5ql9Ul/C2TJjXQ7OXDVVAA44mx
LFgypJiyhI7Fb8nriKUgDLNni2rIOI6uaobZm6NbNPWoaK6EgO3iwp/eKA2tnzkAkn9RILg3mNha
Nrrh+j619iYtS4XarzyGh2+I4H6VPbKJFERZrQxYy0m5EkQtHIlv8mHAupPuTemd2525maOuyT4B
eQCtEmDIZ2TKnQUU+rrCQoBzR37esEWDQgkoqlS/+FR04bZcCiW3z44757QRQrI+/1vNlQp7ega5
U2iFdOxL1xk87U5kTtGGmK64DrUDwI+BboLwO6R+SWPkXbwez1we7Hgig9gXsSqWX8jWn/HNCx0B
x3T3nO3nX9+xWrDYe8VSs/qYASz7UdeXp1P2R1KkUnConCL9msLt0STYf95X3YD+LhS+XWZoGh5/
+tfbahni6u19516CGbu8h+/xu59CZ/ISQ8YVHykTnBVPTzdvKA7NhhWkNZOe6yIvzUOI/jNvm8va
IERRVEQN/dvNt02gUu7/rSF9tDFdJaWAbD+0b2S8L0QKoskrSrIISvEYLIIWmcmgOcZJNA/0S5es
qjPGbzSJy7c58G5JadB4V/7G3FOQAJyuLzB3ChTfjDkcuy3WJeMxRRPYxeid1gteyvNWYau7rYID
/jqeS5TARv0wPPXh+WO4JkYjbqy7CSc65g9cvX2buRM1xkhWKijeUSgmRq7CGISsAUDUwWIgNFdL
GxXcPaoQ+P2K5MKnhksrbc0YgDiL4cuQRS/CJDT4acJbNo4G510ToMXFRbX8x7B7Or1AQs5o8TuV
AiLMaZlV9PJ6DEUzgrB46aSea3q9dDBn7razS2ZoxpKXT34+m+uIg/HYurwRJaR/jg6N/+wKcZPI
2JnfysYvAzjNyC9ddM6tV8Fcr3wJWfTaPu/eqvKA6qMJENT7+L6MyyrgMPTmiaJ6VXliWIju5+MZ
QlxxeC5+oBbeRGc56MVp5ngHD90tRvU3qFhZYfg+P/cc5/GBPec7YvkLsn5TnqsNk/INqJgvp57l
4i4a4Qbb8s4mQFI2cMLzP0TqIxnoxYPztEltqcZvWimiViHOgSbDvdqgw+yINXPw6AJqOOvqfIxX
RidHaXC4miOAB8vQ0J6kDDRgOdfOvvBvlAL/RXcEWgsoZgk5mZtFPGfKl1VfUcW2ak+FbtQWzx/h
N6RxwerEnYdxWazDenA1qQwQw4tHcJOq9qWlWNDEgeSvS1HItWNbOssYO6SZGVTUc52zmEMpwRgL
7LyoeypZKgQX8t8N009L07pQekgy38s2FoZ2cxaZhZJYyubinTu+EKQanM1Xa4mL7vrThfz0Cc0N
3qnDppVftm6q1ppI9x/Xr6sRn/6YTRkQNhpqBoY0qyX9ps6WDJBxCDePpjsaEmQQjrDuG+9lwzgB
M4gniqXZoTeP65EvN2+n8RrTK33Du1DKdxdxB5XArw9O0fCJ0F+uo1f3V6XJYYMvaPNv1xyRre6+
44sDQ5Z4E2Z147n2SP+T2SKfXBxE4RUlPmG2nqRzQCnHkJNtvWPX7Y0gUprhc10NKrUPI5nQI0Wb
ulavvBc6ct1/dHmP6x4te3zsUzbfma7tRDykzMZWn89L22TRiULh4N8NwuF4TEx7iDZ9gdowiGNl
H+V+jIP9TWy2Og4oMF4T+aFFSVsOlGyPOh88pNFM7vFuKRHqtLN+1aEhnQgo0BpOf3vFKfwf1nCo
uIG0Wnn/lKIUHSrNPQTQbS9qIAW8/90SdSDiqIxzzJLCULEX3md1ozMm7MqRzhSQgiHXYFu0YOqO
BvE1SyhecWBSwwTlw11WF3GqrnOSRJ8xatWxJsZ2zfzwtIYMndoVrGggsnVNtZlbQZIQ8mRfgoyb
ETJoYFouA4/qhW1EVPpdLjwNOqs2QXf/SSYjXauzkt8pyDNHCcPWreiZ8IIqbOQ7QITMdx0q2uyD
QohRQeM47iG7VXvfTMasizOiea+F6+TLrBTNZamCJFHPVdRXo28vSX7tfjJC8uIVv/fEzxt8tdrv
XR+/lZuoTkh3elYH2HIdUmgGJ91MtojOhteiwXd25KISGAFGXw+nBtaRgATCQOhcVZD+W9eAKb64
098XpwivPFU4Pdq7PdIgGqU0JgvGv4IDnuejBs25HZpAcuDVi/oQSdyzpRSUEY3CYmmoX1ttQHjb
nvYwHyR9DivlJ9L1QvlIEjum4LnOoazAM5R2MJJj0nUnN1YbN9bb+hqWA+5kAgaaLTzMZWzOIIPQ
aXF34IiSX9QHX1hJbYZzIIowUZa8PfmSQK58ws010a81rCBz7+mfPzYs8oPA0Ux5MkPOq/eJZtRS
OxKx4OCuBK6b7yPjrPRPRiezDW34iAQDW/G5BnCthBEPQ6oRH7b/bYp8JZfF9bZXBdhU57hBk/fB
UeFCVuz3PhPv55RkIHjjPexJRjAXsvRKWsuVzfGbBHDH9mMEx3KAzjAIsljas4yBVhqkfQ1ai8EJ
3m9z4cQSI/A5ZlnIiTh602LkFD7MdXWpSiiTtiihURgqESw0nxctqZlF973pwmQJT/O854y0lcKv
1sBghryxQEzbvXdS8cUPO6iSvW5YGQFzO410x0VSrlRuvYg/kSjnQkfQFW1ychqWkUDDJdb2YztK
B+DWM1+/bBG8+gNI9v9VBXmeyNc7bES3LW5Byx0WW6FNkUeZKm8EZDUlXiqJ4MjVz4t03vd5PLwd
vS5Be7QMyuRpFyDRNPqbaGnj7Fn+WPm5JArsc32H+3Vc0X9Eh2OJJMfYE+MkCl16a2iCOFv/GRon
PCJsdOUYVGGTL8H6jM08rWOnlA+0tD7q5rBADQdG5piBupNewMBQQ9AUxITA8xFkxsxVFoxPhO4h
VQSpLjqzyu+3VsaydrHtPqlLjAWpdrhYS84aaWrwxmGZvoIN6WKfn47Uocf+2eyK+Fp0h5JETwot
VJQYl8Dmh92PeapT1iWD3RSFNoxZ277waeje2ogjK8Ww+w2PaQah6LnuYwlENBsKCt7BoZouyw7A
GCzfldBJCcP8EWx5ovDQRD8gnedRH13zCWUAz5B+6Nz7ZnKoSi43Y7dDBWl+HPVogY06KUQk7TLs
hmD1O7FQNOGYyvCCt1AHDp+IOGFwKWFWlcUP2f9lYb5kf1vlJdXp9jhqMQsIhy9oksC8+1tz3+Cr
aEKgp8k/09X2qedxKXQvBi9Q8HIS4G/aa6vWAm57zi1PLtCr+RQlUWRGvO8Pm4cmGmEmLrLI7el1
+GC8F6ttf4fclmBdOAOccyVBbbdNFY8i2kbA+WvsBZNKrJnddnMiM0+xvoo6eVIjxS6GdX7pK/Ps
zXCGiNBZPeMoko9aR2r+QwnjituOxq05OAeyfeWBVtkizTfmZ9dr+dXh0zSNthvKw4M/iIVzjDJD
JII8U5g3qQ6fS6+k4R7cufNhPjSig3QFu2bldUg0Mpv2SyZdO8zNZckEIgz2cmSJWhDCmO2w8Zo5
S5FbPNBQrZpWCDdvgfr5Tbd2DqlbirzoyiX6gusIwXq6Adf+I5FgzaN+RPXTzayP6ZO1xbT09jwW
lcs95o/KZJ3cJN6ifXePr7Bk0prtI7N6sTDAgfQuPOr1qux8QdLqfny/97DUzXIChQU0he8kzLfy
nKlyf5sOF4wUiRGPxvkJ+62Fd64SsqC9G6thfdwyqBvwiWcc8LV8wiDp5owVcttUG35ezo4xmnm8
p9TpnJDSreuRy1PLxZDiWontz6HeBZuoZWBm0a5nbWdm7XSNj+cdHnGzgnSpmuOAKYDO7VuFopdZ
3yi572rg8JAodvW9v/yaX9Dk/O/AAOAlAJ8yfukw4/hTffJBtB0u+vRCP4nyfjNbMzneXmK8qRt7
okWqhu9SL4pl2FehVTpOEnese00F5pkpWryvDrwSBib4Wu9LpdbLzWKevD4sFNSTLAwPSns+/IRd
8Wfvo2PPDnv1Iq6ERnIN68qhfcqZHPbc4sqy8UR+0Y55Ckv6EpjKIhhnNGWcsJRlXAYymGj6SJd1
uWnSXgsOAsDVznGIAm/QKQ/Q8RVFoScFPS7QME+GD176L9QqGlAHBTIAhXtfW5EHkKmQJbXL6VbV
zid/ko6EMQHTW55svaEoJ5SJ8ChyTmpW+UGHn/fI7aJfGWjv/iOUGu55uoYZ9kSNJN1bJQbNfEvA
1uqeNb/prL04k3a0bNbc2qs7AH8r7ARLtENiMOwBoBLGRA9Az0ZB36eRF1BZiydnnNNtbTn5KrhI
cVG4dLChS+aDfBuxNqLQ1q+859+cuqA48MpEeqX15Fe2brg0mO+r0PF2fG7vIn62AfsrC4OhD/mz
V0wu9XkYU6hzZEHOqPY3kCHkGSqZA2bJgLVZU6KKOF0wjPmb4BPp4Ib1ooLnoF8VKGYs8rN3gu03
qiVUF8cIMtRqDAX291mghKbvkZt9gtJY3ORtEEojgwQBj1cJzzOnujaQW3pa9W8T+pOIWz5K/3Hy
VIpohRrYi0XIgyyWYVhZNTiM+w9Ig9g4EiO4esoNZabB7crnglHGmGcXDkj0nZR2qZnI2nu+fpdJ
HgTXJjA1TbUAuqyjpEYh3v+vRYD8QgL8SPUJP9eRoIFUuG7itN2/vKXloVq+OiPYEHIjL/19ypsn
muF6vE6f2BVbk1X2KsE6ZwnXJY0eXVQqTgMCBnJBtumSN+t0git5s0HKgiP3T8n3RbeOEWvxotxm
fyOTvbWm53ZBNLU6Uafe3QCfAcvbg8iZiODpa4Ud25JY+lVpu4pqmWkwTIrQCLeycQpNh0FImPxE
sqJKva5u342/MCgvDfIc/15ILUpn4m9zoymLPpMHbKrnArTegOdHlQwppFUrlnmeoK5gNOI3PlvL
/+3qLdkK9IinYSi4R+/PGmEbuM2xqn7Jlr8xjIcMe5fx2z4PDjkquyCAVsU3Gv1LEq8fXKMoHVvq
miWJNliYfeRB0fRwRcsuMRgBd339wFiYAt1AQV6Fnx/jG8aV8qpwKaMZ55XqMxvlI/q9A9NbD1AT
QE/bKJZjzZ2oEFC/AflhUANEzMj7oMQugRItu2UsV+p4sRQjLFX0dW71zDP2AU0EggCKkAHvRe3k
/Zl+fp/McDWjFadmbQF9/76b136RZ2B6vIGqcpYi+tEzfnFNdzUBYQLuy9iI02YbcHX754DWV4MN
mnks+tSdr3vQelL7OQZC/SCLvnz0tx3LR2PiG4dVTOgdUSPb2fepooTz3peau2dZ77K8e/k+DPBZ
dd8yA2TUt18h+ulffcNJNAQiy+XuDbLcOhm/XqPKXy9s8b4q9sB8vzyBCL7TKj8cDJ2tebv0mw82
f78xHypR+DFo65ykVESLtgc1L0fspukXPwn7eKjb3AaigkkRZ6CA0tgnRQ/VPKctTRJr0bke3LSA
eTlQJPFdWjnOMLO0ke0HpeQa5IO2Rc+Jljviv/X6RWc41/eqYLRK/yr6kCJEkCBsPv85M6cS6PH9
h6yPQZ3BvhWz2FEsHiOOXxSq8EQHOyyhBo0r/oQZ0GpYZBAYChXeg7FxReOoyPjwo5GZC+XnqPXi
kCBuT48364ICBj7qAIxCYQMrV6uzDHhNSYI2XjwcKfN+Dz2q1kdbniCQM5/D2SdIDbBN1mKjo7Mu
jpB5ycMLlDA9wT6MSokLJt1gPFQo4CZG+7IvWy8c49UbnQ4HyONUUyWIQ3Hws4xuMf94thnWZaIU
Q/vvv3a6h4PyM0D0cwqC/nAeBzUdbz9KC8vMN42MOv+YGn0i6s12oF6dDNKn0E+9/HvHh8ncvqgk
ypeJ6/UQloiUa9lKdBc3zx7TSKh5fXu+W3w69yVWJOefZ3qMkyynn2UfP/uRRHxqq7BYj6OPq3hL
lhmIKbgHjckyc8V6XzZwcW5JeBW4YuAmiwlOYZnYUHFWZ8z0n2HDA5sbWXfvR46VK7mh8raH8Kz/
DQzxZaXi2SweyxVFnGPomJPRFxZpnUablLcv7Gg60yqQtO22awG7BActB4mKy8MvkvUkDHVn+AJA
0aF/520IbvZTUDZbSlPLd77QI8RHf1tF21FljHoS/bDD685v9OPcoB68jzRGk0BTt5zuMtIJVkk7
W53zwoQOTIHLb0VjbUuKHt44+7bPHot8SAmdZBrHy3azEFZQjMLhmGAPC6HwCa29fRCSak461nFa
KCDwa09Ru567ePkM0XL2Y0U9kswufHbuyR+HdwWiu1q5Xsgad8blaz5xmAhGbjP23dKHTrXyzyVw
f2F/UMNbD3DYZN+UKlAVdCcMS5RFkDMCtEZAFGwurXxwfBvMOtCvpsAeZfTxkxNL/rWVCzkynyuC
BlJvHnXieQpGLw6qoLXMFJzuPNMqmTUm44sJEmvQe82pv6v41uuxgMCZyBF+RetwXqPGLA8LOAkN
6GcpRyD+xcWNXdxEdnHuivbHlSyN5q/2uFGmzfy5ff32JQerxy4Qa2seE676UBv9TGf/YAKJdbnG
POF90kD6pxrT+XiwsWjHXmQJnnC+ak+UhXQbWmtCaLuBW9TPX79sjrucr9ij/CWZ10E/yZUgsGni
eh776hlTeRYicCrWRpjCHiZNIMC+yjf2G4Se3rl0Rr2XxNXxQC4lyMWC5sjYrEpWBP7NrSn5wmfz
4AUdFfQ0czFH7/Y58Mn4VempDEiWv6SF9ra3e7jxEqc7/T3NUHky1M/rxfh7tf/yPNG76q3LwjYW
BhPvrugUCwYWPaMMUzaYCxe8IRWTO4gKIEbT2LZ6huqAxF6yudLNogbTSRpIm/BmappjkrMtTetW
oA3wHHi5bFePXvH6ZAqZ/BXP4zhv/QCooYMD8M6XRm1OwJDbz3haHAR2l3pRqK7mCbikyilwX7mx
3E7ecmXmBy/KPEJchWz7FZaA9x3hzTZXJ3XYaqxWd5n8VWslVagkMxEMsEHCGrQvAOxA5zZSYaHe
xTvdZj3+c9bc0RZRmEJJ/+NXqEZjJDn5DYJXcXpomkWuWGea/w2i5lyU5hVAVoxineH22xxiSvC5
Wg5O49DcxKLAd1JpZoDjqcJ1sY8yyh2wQ3Rz8MKtqkoYECBDRymd0F0xR2P+zqz3ef9F47T1MaH5
IwzYM7WkbhnkTh3DwQ5IaA8oFlHT6desoLRp5dvEEngQefbma/gwfh502wA94ZWVdmL+9HSheWco
KRADyQAtp123juOTqhhAXO3ZHuzqT2Lc+WAH61ocIEiIcwZjSiruqyBk5eh6qkKbLTMU3NyjOinH
VBwtlPUr4eUf8ukrhdedw8Rrm9iF6wvBqmRw3TvlHMabVUANQ7KoLNuRUbO73N5jZWMjR/wiDGCM
9fGp5RltujiD9V+9FQqSdvJTk7Isxzk5EFjl26aYoXx+jAeHeIX0QllmjxjayTEgT0iva2/26WqX
RFJefxXm3dh2swQ9ub3JCqL/KkqLWSPMszpwfea9USryp9BtdQbzsqwDJOw4pFzEbKMyDEfYgmF8
lcBfBClNfp1xwQodhlBY3+Ov3fyvDzWgvfC8cOveX28OWrGZQGb4Y+6CbZY5QAgN1nMyFCoGku1L
ild5zFaKzMl41zUcu76zchpIXr58fJK6+n6WDf3qzfzztnpSL4HPuRlscFwxKalMzoPt5Q3Jw4dj
dXd2BVDXRORcGPXUeA+3uUxJOSUje6hNbJiNvpgPKJSjiGTdcZsng6U9m9anuWVXuQ0waVxU4jZv
H3ljE1ttatL1SruIEdBqmvD0r6MOYC6g5icAcdpPngf7TvZ6C1Fvibe9cM6lW1SmNbtP/Yc8Mkxa
5HkyssiBHbstEKmSz2nF0zTV3PeTH81yWUf4XTIVVJnA6ZqPk+vAwKVxFwmYDlNBROm+g2qWZRf5
TZ8hDV8ys+a16m271Ed5NJRznzTyS2i4nONpiDRLh9O3k+fogEFluKE2amySpxC7v3sySPt6oQXi
T1mLrSJHLm6SZsx63M4j5tDAqn0B90fGMBwW3KwxETR/ZM/pw3aWl3ZuGjCd+ETV6x+IMusarFIf
ILGyamWOpumyHxVW53Mt0xlM8BESCn6UAuVSGb+lAk2JzYVM5ZFfIzOush6DEi7EY+fDWZcYMRte
G4Vb3AWoQbYNbmvRi1NGmf8OoOPRpRcXRxiBOQavvD4kTukSKo2mB8VeEnvkEoC7wW8q4IDa0bZ5
ivLquMxiGAk1vS4K+KEytoH4xdfuqCTuyQIBhc0oov3icP2+F7yg/5RD3ObBnb8x8jV+GWYjUD4d
Z8JZ8UsuzgMmzvpTsQkU1gXKxk5Uymnn2wT4Z2Xtjhw6tfkr2KqCoieNZMjkwd3/7sZvQQZc8uXt
QAltBCX4eWtul905JrrulgS0oBK8O5pSQ3zRCGMCT/CFKK/6fI6Nbgzq5o8VKrstF0GUHUyDDaZH
RHoDRI57tPMaR2I3qT2v9WSJmnqevdZbsyZk+ZdJEmNmuRsoEDOeCTem2PgqzOFZ+AF418QxV/dU
eM3hSorO5CwXqi/j/I7rEU0eJWvi1uQPJLrm1u1nnnnf6c9P1cXefZ7Em9xReQbG3Xbm2V4NUPuR
2Yv2/4UrykdYRUQKLIGitWhWVQSRsTFDrUV6iBlQKDow8cOyucJanL2fKxgcvumKlSV6+4vLM1Ac
bQ0KgyH5GoLL0mw4XWVY3zDOHSu/JBt1VXxJ0dMvLr725xyturmLkDJSAu1F5IeUpKTb8gPx7md1
4WQgIbz3FhU5UPAlfZiu+PEyoSiCoIDNiJ8oPe8BX3g85GqhJWlic99EuP+30Uu20TEcK3NyBE+D
RnsNRroa1n3ZcR1toSMWmOiWYmZ7Y92qj6VPgaaWYBI5/0mtSGwYNNz6bTDVsKgacCq4/mQ5t10X
DF31PE+cjZ2o2xPdZTrtHhAo9o3ORiD7aWQI/PGGd/pEzva6Fb0vHMtE+1BdQQosKCTNVrS0YDcy
1gmJxAdHYmoVCVaacyB310ZoYIqjxIorieyZv3PlBk1375krAV7UuWSrAcKwMOK7Ks0oNT6uaSuR
jqbwBtsT1+XW7kKXBVW16GOu1jZ7RQ+2THQiQF9cCkdS21ZmXo4Rw3BYyeY6RvQtLicJvnuTaFCY
R8NLUpvUSfrS/R/SRlrw+NCVaxVotMLUQawMj9k3Qol6EbedPpCfv29gUdEpz3sad7thDcCpMxSW
5LLP0hxasWPsxcJyrdHg08hfs0mm1TbBM8tO/6FGHxgRm+jC62mOSop3P/XxDAxuxbUiNG3zP9uc
jApHr6+duPogkJE6np0KpWFyvU1xBTgX3Act7/sVFh8V5PaE+xZysLUGzN9cSvyFf032X0YvuqNY
2Q/lBwhg8UhJ2ygig5YwVY7srjvZwD7PH/Ybk1jOZSvncwsM94ESdFNEG6C6nLByLVH65ohkQcdf
uU7HmcitazAJMb/2mcY9g+cmy5WTsPRWVHDUOPCy3Xp0ecjFp6vgTVdTBO9//8CifoI2MoC9rCdU
kt5Odr0W5HzWQ1WJaPWpEXXyMOg52d5FaH91ORLYLj4MxKh1huVW2M7rlmuaoRMl3gC2mH6NMlou
Ctbzpc76ssD4KRUcquoAn/TqwIrhoKxdeey4Ta9VOEhWhLzZ8b7OuZKfYp6b4G29CRvj8HM4xKrz
NP6cgrbJ45onOMAc9d84aYIBZ7ONV9gWUKTbPeYiGBQPR/sjrEEjQPrHbLXoSPMqYP1OhGDDu4dO
WdDQglVvWZjPvev+8A5DL+UNBIGjjm+zcpUVItnB7Gj7M+EJFpejHwTaXquDyq8SsQKtMmgONPTA
9PUFJicEgjJSNT9Ch+eJmC3uEyJbOGgzhujDs6rBLisfwcGTve4h/iqSD/n8MON04qJnNZSsQNSV
IhOCms4YaSPJxazGTau8wi2IqhEU3CRQiq2OUvP9Gqg8R0KscbSh2D3hu1egEQQ6jemhfD4q/h80
wR1enClx+DyCMgKcg/Yknj7JI+26yiXFrSknp00qA4BH18UxJJgjfR+8CyBAd1DWumLVaJuetlTP
DEOQhZBGTUEKnwFRtCODONUYJZDN40HkoevO/AB92/8CswPJMph60rtVNwPom5v5Z/3HDmAh5gEJ
Qqj/9z9B6sGJOzHh5y2fdtUVbyCSIHwZIu0fNW/G+AqrEHZUcdTlry+M/NpkZs1FgSk1BTOGMvgE
aeND+Ey239Uu64wftC0pDiV+P/xv/6O4IIFbIHWCger+HtXxS08D6cKucH4hTOxvQ1Gtsn6wy1YD
Jt/JHjcKAJ0uGULNKv2E+3UfPSvsXorOMHi1KwQ+D6Yt+i9jMGlZhnlDGGpjBm48tgGAxPmWJpHp
HjRsOVZta80Ak263uJPpXArRut8wIyDhJ6Z/h+R9GDGPeqfgY4grrqIt0A5gInLXeSeNMtJw/QNu
xTTtxGPv7GG5hFuIVQEz/OWZrmnFc91dpsX0gXSCh7oakxn3kTtJlf3Jkoy/gYxHsaMLJzqRtaIZ
Qi9YLQTP4qOdmZ/mmOc42VRk81MlSdOySAAvS40PHJrfmnOf7NhtSqX2kQKFwe205aK+/s/LnSyU
ML0BnkN5HIVh/psEZSclITrYoyTZDqiAnUKISED4zER3JnRSmaANZm7upGgsOFmMgJPMmzm+QFMP
DgvASzvyeM6+7pNepHI8W7nwZyrBCWK2vjklwbniR4Kx3eGNxlttTX0yX+C2QfVNJpzug4L0nQzy
BT0fsrsGh2AJGG3l6GxQvL3foWAdOaQZwWq6fZJOOAFEYl3MgDTheXwmD3W5jKdVlzs35NHiblw9
cqfaMBJHwhPfADuu/TF/XK5I/d75yBnWWAcec0ylY8G6P7aQ1N/6jww8nG3C/fGfVpGmvE2jubg9
IFE9Puqikbvwqg+9Von8NPFuzDh7oDMFO1775stoQSxYY35vqznbI3EBTFdaZpo6bHBh3GYGu8nD
eT4QxcdSx4ibY9zak4hPSDmm9CSda9kRzjVmmokVZUDmtj9AEYGtMgZ27tuSOLVm9EiKGK73UHdM
psScWu+jhr19oirfsQtYQF41UWobAjbZf8I3WjmCUcBJqAu60w6lGOokaAkheQ4rj+XyF6s+Yhrk
7bffbjmxRTlt10JW23dhOIkdF8VdRbedO48LczUCfSeh6S6iFKUWKGz8+Q56ulMALXzNytD/KDHV
VibOftbIW29xsA6bPbV2GYpribgUNrrw/AI0zutooDMvwKB//xUco7vR3eA0WHxKF+50CCHXUQ0F
6omU7+CDGxp3QScv7xvI7yhe+jrGEvxvACjhh401wr8Nm8LsuFujr17NMjt8yJCDKBBtcBDppUvN
66neajdPtpWCHfzjCVxPUCGlOqbUqi1AIpScjrfB+AGu6hiFML96d1pKzaS635qSM9nmliOaIgeg
vbQwGFy+FglIniuQ8A7J5v7E2BxxfGa36D7+XWmZSbZ5swgFtDBwA3NZiU3mXue4wj2VGWIsOrbB
oH2dYQ4m1Gmai5aC1KC9vLM8GgTpxVsIVIdjY6lW63WxGGmSI5hUT081w8vZOz4u71rI/8dRYQxZ
JNgIJ8DlYUGXmqVGuSxk/UoXxQsWCQZOEOdjiNaFFjeNUiR4bDAMEAILAM54NRkdJ1og21am9xio
FIJyGKETPBYMGvFUtTmNWXpyGUd10HNz6WBCmekaXvQoTpg9Twx3jBW/rGinYSaSF5RCBvuo98dB
oCR9Pu2u16qcrqA5/gphy7g+i2vPcoOI4nJiijHkh4+HkB9tgGPZ6p+kbZpUfxnTvs40lFefZBs6
PAtamBujKs9fqPDnbX11fTKOMNfEev9voRbWs3TvsWG2EzdgObbiIw/RKu2ilA/UMa6cKy+f79Ae
DDdjx8LbeWTz9PiDwUYMvUrIheYu8yFmw6whcaJiJuSLbvYjOOitr98FicC/K4KjqRSL01eCcg/4
Tq5/tjaW51y2GClhTlQMaK626V8vfiRSQgJlaz+7TOl1V2iEL+CyG2suFZU4HpC2mRRMr7IOOOCp
lwHNQn/10C8ETLz7CM6wYfBGdyKmOdE8hTw/c9jA1o5qOYT+L5mrp14y6QmrWsLy1mWxOFDczBv3
d0n855g3csRdjzUhpp+RGL5O3LqxvbufcEmxhPHd9V2btrgj9hEIY4pCXndxgJoYLJQT6xkTW+Bl
35Rzv2tOeozYkrcIyu+/CbW9NzZm59UruOj8BeltqHAbzJnzdqrMepylnn+YWCIzQvlwXylJfgNp
PFTwLGMa9eS8E/TbKERot5BISKfVfykIbdwsoGnKiMvc6qhifF2obtgaUfyMncTAJZh3arI3z0wt
AOG2A4sCJBkOXL4tPRr+ldg0+3WJIfxpAL4pvNDPMlYiImoV/HcPXV81DFOPQq/dSAic5byhuWKl
ruIaO/0LV07ZZqWGGyss9y1gqH4RLZ/dEaVFBkGFX+yAVCz2+H2BCzoE3ACSz7B5g9+wWJ8G6zln
hGj6v/DuFss2ICecmeqJ3lbgZSDMJgWFxG5t3RATr9v22uOyFEQdtclsnE0PIVbewFt+Tz6FeSN6
O5b1jR/3r1UWK90HmfYpxAypcjkJb3NS8V5n8Pcy6JnhIGgYgo+WYmst1peKC6dvVG5i7BNjrgPj
jdYgVzaPhmKzV9UrwVel4tABxzDKYaCSTlPJSV45JpxdfEOSaQ8InHcRStFdwkPE+GYj4THhep30
OQ8aepnhNpt7iBXnIgGKeRRQbcIeCDSI7VDSw99Zw1mmqcVf82HiAs7IXUGEPYIefExEnWhxnCyg
21P3JyA35xYzU099b0VDRoaad2+DiKQ+t5mNi+zGhmIBTdPBQcbYdK8rb5ZyFYaGdciquC0Ivj6D
BnC36xEDTT/ELROq/wU5ohsPLm4VCI4Hfr57DD1/U39sBpIl9Di+/0kQZMjb8sTvBs8KMnpDENDV
Ho4ioO94b8Wswh6htHuWtw5CQi5tPffjye1xK5CKW/UkxB7tuACBrjZ4ILbrhik9kLHBbk12Tx6K
7hkHzMP9aq7NOD5uI3ZQZCpPB3/XSICBpvUm75yo3NaqT/9I7aAaOZFPhfPFxKeOPi9ARa5zl8he
lKRqzSffUUrenLMyjJu+g0HscViA8mi6tqtHhW/sQNfihaThrPjgzTulBMggpDvF7lr63CprvWnL
UVwIKsNZPcSXrALxpyfaeM7w7rQl2h84ACORy+LXC4mLfeoffo3O/dKlWPqx2K61X3rF7fnKOSFs
U33vHyf4pfazZDmIMWafE9fROH7FaZAuAzzGXUGANOHRfJ1/ERK/hLwn5fCwkE6o7uWEXgD+b9RX
JMGX84jCCrzBNoP3xKka8VVbuPMqH3lD1hUU/EVL37YRBnUOfUJ/OCj1aqF96/ASw5O/Z8caiyoe
qr7Po5R0gzT8Moq7TVZQkhJeyXEKQSerQVGp9XUXlnmZzOFZyM7DB/tN/dGe7u0UkOKExXPX4Y3g
350QrUcOHEd/UqEctZZGxL0JdPrZNLV4l4lGdGP/W+Plk27JbW7lEZC+2fSQkoHFkTamFICscbQp
chu0aIKOHfMLKgdn1pSspna36a3pP0M9Lacs+tg98NL8OEVb90sf+HkwvNSF9AHb1H51mTbpUZ9n
d+v6hCuCZ/QuFlUxnCIEBQZGLzfgokxqDUVjHH3mwOsL1lyyY+lW32iERYx4Dw9XoeJSUTd1880h
scrxNQ61dhIb4Z1DixC6vRZwWBwnNzj5smKf861fGvu1C+/wrkFYIFdzRY6BeCfFTsygiRH6l+lz
RBpjUeFCZvHYKRtB0yx1dGcjMIvtkOOlmVEctXxaijFE2sdPLl/gcqOHddvwWkmLKJEowjK5pYzp
ULu4TwCCsXefxeqP3waUFuQ4+NHZGantx5eB4UIShpbbdGrG/gHKY/73ToRJNrtlCU1ibl24O3vi
sUzui0EbDONIEsa88zPpYhBM03xnd7TRdECW7TF2/7g+bVYuzGftzqskRfwj7JDnYjeW7ji3pYxv
pgVif4U6PTR9vfQ4J8TegJu+dZZBNJ4a0Xb2FJ8RMdIsJ1K7dqFrSg5jLdRIsjuW3nuEopVxBcGs
ie94Hd+RwWzvRCFmPcBy08v7L42nZcmloTWxNvDCFsoAYFzsiVUR9/7pdV5i9Km/nI6Q5eaKN8zy
RfWMP7dZpUcUZfrFee1k35dTyRFAavQYU49665OUPoCNIZ/991G3V7RD4ocxYV6zMQJ+euE5UA8k
qZOGYCiRiMMJcpDpoNUr6R+lQqEuUXU0sokka9cgeS7mvN3gaSuzEOeYow8rcrb7PkeE6MT+5pV7
ywqOmTUWPhm6mwrXmwO3eQhlPcVZtFxu0rr8GS/+Z2vK16AMwFeBXuqIkD6SZyLPjeBbC9KnHbcL
zFIcNUwAHsHN0dDoS4MlNoGc0c/lRyBTmE3c9VEKeDaetzr8Kk0BU5hVpcNUvkoMv5rF4znT+X12
W7F8ZU7h5vtzBlHzAAHZaVxUJhgn8H3ub7eumoejb+fC9KXfY2VpnanKUGCxX40oWluZkCG5nGdq
nn/3ITDCACHkGTmFE8H9+pICW77+A1t874VfsGLAIQODKWXdkqxA2OJfmNKajvVK8kk4+BpZhwVN
lr5sV3LMu9ZsHG41FNOuVTmDypi3fx16H/b8jmWDg5JlcP7TqEugUT4NQ5lLYUM6q018ABifT1+f
LgGBZa6l2fCe2Sby7Sd4+8nsxdaT0sFcyyAXUnVsBdPVLToBS0gNne+7tHfyUOWseCRbA9m9jBYY
klpHydMDNRkvEglGwzhEceFNdg7TXjN9B/8qp1lqPnxFvBaDhh/iw0ovE3tnyTzjcPX94kYRs/hA
RzXjV8m4pKPaBq3q+R1HmqtQSt9wVz1qVwfGhq7ABRU5hzcnQ4/0SoPyHBs+86B7yZReLDm+AY6S
v3C8keTV9yUE7YPBOigwuZp4kkmlsp6XcboSsUlnGVMQRVJSn8h0E4oemsoqHPnevjVXuBreG2up
5UZ3ZWU/xCDG2TbOEYiGX0Zanb/nxGarmr1thci3x96u/KlfBDQ7wrfnRyyJsA/Xb1urlZjR7l9z
wsIPpuaS8fGlf4Eoq7unef3a90f8D9UbLezWRTHeg31UNazjZ94yg/HAqsLlkwRqN7C9NYtnoTsc
ncU6KhXM+iPXI+lR72RkPpNphHO8dasKJDT3mzpjD4bGW06Y4B0trlHtigf58AO/cT/EYzd36Yd5
ZD/76hv366aqHSQ6UpkG3rYJIQ4zN+pjqqqBGq7FVIDCDeUF0wbCc7T3jztKRI5nA+kMQAoZRgXj
8PEqSO7SaDvmpWnjz9iaGrbZFD0BqIRZNzH8jD28M+9pFaaUYxn0VMuK1LZjeeDZCbSyJpVG2tvm
ijEfnbErOkD2PTUIekR6NSUx5bKEdlIyMo/wFXr6t093jkXrpXfY3YCwfMFssfytNDLf7sCMusWh
/20m8GPCmoI3PZT6xxwu1Q+ocCwQDeICLlDBY5WK4OCqDEr07tOu8iOaQ7QkxT8VyM7BT86dLgeJ
aPUh0uoshOn382OLlRkg0mQtwBfqjwg4GiSiZydcs/l1Kv5yK2Z8W+j6K6c4HAL6vktWRZYiX5Wf
Gc4VoK5uiVl10YvOX+Npu1YWgkUkHV2rSuSPIoxce+ltMa868W/cE99oB8j13FG5Ss1yI91titJh
ZMNWmgR3bjv+YyrL6pkqLRZo8EnJzsjeBDODFCKsaEvIIuMhunwbLs4oUjA0lI1Tassax4VXsY4v
x4f0eLmvIDFwHcR7ywtvFKix+nGnvpVOSpUy6SjV240JPc7XWYLb8UuRLTYuBgrxs25DdKHhhswr
Y1XJnqQ4kLcIH9jN6ElhZQ7rLTlleCehT7NYiVHlWvy3nZcqmBq860wmE4PCkHgLEVv+DdUDpGOk
WCkWWiZGJ4sY7tjQ6r4V7Spe8YMkv59UcYGOo9bClZTV6JxqmY8Yu1Je+1guT+Uspan7afN50X0A
Mj1hMDtqyFr143uoGMaXFsObYV4TBoVZID3PhuEs9TxabCuPRdjiieqrgvhetlzOcFzKFV5Hpe26
PFxgo8u1+9bMElzT3fjTrC0P+3yBGpwiCiGFy13ZusIsoPtyEsKSGQz/ky154FJ77P1Sy6wwLFht
Gqyd9NTGSbdm3tNX/IA2vPOyaYaQirXJRE2WboYf77GBxhDguoufMmVjBhrLTIUmIJ+5wZM6bpvP
Kcpi8WICnjQQk+Laye0p+IQ6sBPwW2nzW8kq1/7VSlGi0ncZl16CZ7MsXKY3wc/tanOT3o73Fjny
C6Ch4u2x4D3wf2aLRPtvoD0b956TCP8xPLuICuL4/qlU+XSR6fHu778cUWX5ztuf6TO6gHny7pFr
sYl65gpqvCg13OcXK39ysIbVvvE1VaR72UGKGcLgDtHQfyxSVNcJsk8hwGGa0SWPZN1cJRhxkX4S
AqIKWwhetxjE6lS7U2a7vzz+BGE5tAuOk3oe6AVpmECOCQMd77/3gkqDbyI5h2Wksj996f1fIl/M
6gsKageZyuDUK9DPEfQ2IG1ESWut1l6MZW7SoQnhBdlZzmdVApBuKcAVhzR3aOd8L+e/QLuPa9Vy
1kf9FPaeUXzh1KgkHQuM2RH7hlDPkHA8fiLHykD6rh4/PrbHnImUIBnnxB+3H6vjAHPnIyAHfSWG
9mM35RGXnS5IWvjyz88uBbPluA8RDANaCc6Scrqt4jf1RBM1NK/opi8DJvssgm6WXsw2sUst6t/1
AOu1n6ibFqLDBxQWzOebOzst0y0UdjvQmBuSLKNcmtO3kOzgkLe54o3IFIddYjHxOCXv+6G8PcFt
OWKYEXWSHgTqZ7mR4h/+iXo+tqjfFJF02n/96zck8gXi1v7oD5HYXSMSniX5bPabvnQB56BeMBCL
jq3ZnpVhI0MzHy7WGpkJtaGVNRRTC87HUXUjGJpNRxUFhACscy+Bm38kPgggW+kkvfx7hwJ1nYpb
C0Q/kca8vnl+8+ah2mNIt8GIPtNh1FjwAsND3unaVum4uFByOnUNhDV1snTlki4b+VHlZceX2Ll7
CxtJKxHbwj4+SWsfB5xRVww12twFfGEGVdYT57rauC25I+UsZQNtDOKsXfDM0I1CvLr8g/XX+L/V
OqK53NGR6YFeYK+vQCl4BE61gklG7gqUT1E1tC+gyTGxDlj8NrFaYbcznqdAtUiii8XPN02Vshy3
SMyHUZD0aDGESL1pjdGf6/sTF9FQu5wAg0PLxVllwkOSiytEY2ckbUz5PFN+aSlDbrREzrJVzy0J
V+YHz1Jefgz0oeGEhwt9RZGNQ9h1W9xQqHD1R+TdCnxbXErEVzY4RnYrInhYK0gLc3vCmG5k7KWc
REtC4wRjRSRF8bZEhjNvOdQmTEpC1QOzd2dL+ZC043yjbFDHHwaL2Av4+EglTC6ZmzVDIzBE+Dpg
HyjGYM9YJ+tvfuOfbI0Yg20R9n5+4mNgyAkXS7iLHV98KLOfXlUoajveYWJwk1PKqFHTcmc4bI7G
WIweuCswgenKtpftGUxXbm2TlX/JXjY9kMHIAlWzjtw53E2zPDKYPe2uQ8b8wxtG14HT4VTOF/nE
pKn6qf9Ifi4xYY+kbN9sMQAoCFX21s3254frvFha+cVm4kaIkxx6JKOzqXYqCIBKR+X1O8ZofzLp
MWHMVSasv1IKjcah5dKPjd5GfaQRJhahM2/XGNLKSyXBIlKlN5SmR0i0a3Ql3NehEa037qRocW5z
ewSiCWF5JVXTZWPQyqz7FUErZYPMutqBOduVa0nKkbXWn9wFnVyTcGFpskYKLJcC1EzitnCQsT7S
HqILeaUGFXfZRsbFI6/c/5f40ASe6ZS/MBNkQ2ltsch3CSiUZnRXZPptnY/ez9pf8XBawv8sXcSr
2E+oxXn0CJKTlKoJK6vERxVkFn8YtNpPAkzYgJQsulF7noRVWkDoloMciZVX2a3SDd87RdlIYnHE
2KJi1zL9WYPmDmvl8Lelr0lxzNiHS3ere2xJ6WozzyC7wmATF2NDMXaQiIleBL3MqM0Yg44kD01T
S6HpneqZ5FU6o90JfYn1rknHzjqofa2mT99YEQvptazXrIqKRCxnPDC7sKO8dj+fYm3Ux2nstAHO
d8Ovhl/ZmQW8iOidcVmEYTIK+EE268Ga1OetE3fs+Av2ox45PdE8Y1Q/UDiyfUF6TDNhmw9HkWxN
XOMtbuvOFxnP/UHEyuBbj99Y7kyI6vUuNq3DfJo4jS1ivSXepodSlpp0UcpqLJW9cwX4k1WzxmeW
GV15fhvFSIblsLt+WzLROk7cuq65lWhRo6R8PzRpxrqfcnycSbod97w9P58kSrAs54t2oZfM0AVE
BeZ4Q8UA8OmsRGzX7wOeggISUiZEjhiHbzLqna5Dyxdu5S88JRNd/t+rodMqLMzlGz+vTL7eFvKy
Jx/JWQPdf+i/ly+4W44SJ3wn7p19EcoUBkJRfEwAyDfZKaMPz1iNcjH8gksOmqjlAh1wdyK9TxOh
9Kp4YjBTm3rjYgV37KFf1WmKE1F08PvNy/mlEbH4Jb3OhJ9RwAu8Nymfw2ARVmEulsrdA51viql6
OKZ6zRli2Jdy5Mo6IUpHegvSfBuYX1gX8A+9iIizb3ZnRB4kuHIIXtOuRZMicsDkFhA/Hl1GnKIH
eLR+NeAU67uS7bGjel3lwEa2iQTS4hVIXfNNF1+sizOFltMeKsnxWcPbBXZWQLYOG1Gto+ohkm9a
8rvIf1mPaR67kkNVol9E5HD5Zp7Y7rYk7z/WhjCgTJHpqtS4c3zR+9hvIhRMiBaUwvLPTznTPep4
1SUwoEfCglgNKM8RZ83T40SYETnW9CTPJTVnEB3SFjv0vrGvcHquS6xsRYOWUbwkJzgmvbJd7MA1
kh9kHl9H/XsaQbkE2gOx+1wqpXp/uEZwudTEhs2NkU2j7Zu7UcgyjCrWd7PZXTRA500V6cKkq3PU
sgv2s2uGGChGknctavctlVBBKScR4Rbct76WuJYgwbjgstclgzKXF/DoNYKTkM443aQJYNo+8NZP
5GlDyJsiPUbm7vd7SatBTYV0g/2eImm0REhBaCTD/SKmaQ6WyR6Xd5J5U6XB93N2o5+XZI1FpVRI
haTCutIAFdaNcRISnDB9X9yqoM9lHet40u1UudgDhB72A02oCWf2pcBZP3t/th8MxBCKmvOefGLU
C3XExHaPmYn+U9xhdF96sqL6qZ2PiYu5Uzoeu/Oqi52aO3OJ6ua1jqWUDUvZkHARK6g2rNMyn7R+
VPJpgsvgGSjVBUeGcHuYJqwMJZrT/fT5HaZMYF7XXe6rQGj3aZqpYYaJOvYkAi5m+It+XwaQXlsD
pigN8YJbEm3XF2EP2kLbwjH7PotIP3Gnqad3W3a0afNIczoGgVfKgjO0ZnGXsz4TJ03N/2+jj4bv
gvlzSe8+kOxL+4AdZyVBd6vxCqyafWDSZ9bEQm0QTGWZ3iS1ZlQ7huET0wRMgQWShRnlSJ93baZM
NFac1cu9hNCUkIqTA7E8YW8FzJFNNtm+d/T13p6A9Su6Fu43Bmc7Z9ef0kCPthjBqTH/L3odBeMd
Xh4mii+c7d4XAUrM2k5pek8Eeq/NG2fvWlkclhOFcCgGC05DA3/xbNaEBCstvXh4L6PzUP18HwKt
3ErHa9aAFRSjTR7HiHBpA4ram8oJf0fptVpDc37mUMo7IaNR4LWLs2Ctrt11zK5sy5rdl5h+8I98
1ulHAfT5EsOTF9gmRsIVEKBZH61ouGt4X61bczFjcg40MjWeQkKLPwNuHKIFfugWAGYeFLKFizGW
0woWbErgZJ+5sDam9abyNiipI0RUIPlEAar+cXzYTLI2V2SzdhWP20XovtBsnP2+h/tmIuYe6VuH
Bp/EyqzsLVtG07gjeWGJuoq1xbNfP/qirVWtGUoHWhtLsmbSrg0YKmVWgyU3tuUOoiTtzZCLXo/U
oCRoPPKnEol51JSnfbPQwdPW/NUO/a9BZoV9ObNFpq1Ee8PYEMWl6ZSy4CWnfQu4/pso/SZj8MTv
juxd/a0OpG0EzTU7AAFJExZpPXkdrDt9WKTpEgN2ALZMbiuaYe1DI/iO6ZBsLvJKiXJBjzR3iru2
bvbgbbwLJMfq03DbBO7GqihgPNiZCvxdftaM1aF3eCae+KMCLmOQsxZEuCcUKD4gJFBNhjwAKkL3
t/e4vIc2Pgde3jtyzlX/6pQybNi9ghr9u61xuj85oEXj6jiHzE9Yq7y+2cvEWE5Yfv0qnZB5ESad
Y0lBeYKxhMoJx9UWKay5LjZ8ZnMxeSXGtWWawaMTHYRzkea4ZG3rYKJYHUZLe9A1e0D8RLsiOCon
fxgyrypNjPJqSLbx+b5ENsLhhWbfgyymeje8qpRGlNBQl7df6PFkmEDZSRkk01tVBZL+XzN4g8i9
4MB+L45StaF3hTcgSHz3gORxpqNFOQc2N+n/KUiHo2q23OUOgUE9GbpYPVF1rYCv3CyTrULNGVyh
hswQD4WtOAEn4h0Yj+pDTQZW8N8XZf2IOaRFmrcnnoRTtmoxzLp3sAUo3Clpin536tZmgu0qAVsV
ct9dhcZmr18zAf+YO3t14MvqGPHBP3pbz8r8/3VqMBmkELKd3MpKPm/IIglzN4nwxINFkDRx+ySc
lXibg1dl29vnNtqIBCatxES6pcLRlR7ZmvNQf7qVeYj1B87ABdjOacXDImvwCVP3T7brGbpiKTFx
YOOnLxHs4Kr74ioxceTHDg+MUzAECIbwPkuYWu3ChYIjyV92x/WiRVtQvssvVy3P0S/DpCgxlAcZ
ahMMz/57IwIYGbtXVkKHzsZHcVj4K4qafbmTmaUnxbXyRXoFAt2Wan7R/7XwdDjbU5+L4Chpj2Yg
1QqfmlRxzCay5TGoTpAs0glGceoq311RISlb7wy/3vLHZFTdyou21vaETfInS/uJsIrblzac3abx
LmGS77s1OuIpe1m7RwRxyjWOUr2QqIpmWGoiIg0WWjV0kOwMbsNLlK+pXyNB9RiXJ5DZL3vKhO5v
0vNfK/0pAaSgqDOJK7ThMPsAx71f12ehAR/kdn8+0Alqim/9qYueTNOhYPzQgpqgzzY1n7OAv4Xa
KaLEUj+3Q+HuozD4RE5A4wbis96pbEgsVVZarFDO6QLGQw/BnPRgPCLs5QDDcoGiifi81H38I5/L
WQbzbW39SzfBNM6X6F8EHZHfUn6GFRzW+i+SuKOXTVAiYOFUqPftNlhY3YsN0j/C9bO1Ve0VHxZT
/9//TBti1rCVNpoZqkIjgyBGd0oHre6M2mEc5i8xcYiSn0nEE2zpT+4I7bA1QLMS/z5fsKPo8gPp
3jo7idZhOwd/0Cb1e1J4c+uRsmFxrgN3K9lLoTFYNm3b1RbIkPwvkD3M7WZxIDFyMJBrFRlleUzU
KoZ1ejryWJZJtaoVpQGEJBL5LFTVwgwE5liQ03fePj6wdOPrF2EXNiSquIm6bXTO24TA9xp9oNSa
fQvSL13WoAm9zNml92n8QkkfjSs2RXS5zoEp7WsfrUwS8HaYmMSyG3fXmp6kLfwbOdJsUEXqrjB8
GHSkKT2sNFGLHPc0dB0n8+CovcvkKjwX+f72hYtH6OqeJttFZY/J/NYVqaIwbTM0Ir4qWTsfqZkF
myV8JhJ1QFsREhCZ8YPep9AizLqikkucM6Lyut3wMAlVm1fS4bZmPKfO9kG8ea3tqXiTneeP7c5l
DuqtVTsUhbAEq+CzsQzpugYOwwb3YO6Wg/gEesca6VqOtIDfzJNqJGuDoDHbpLsEagpkJaepwL7B
3HFcNYPaSLw+uIj1ZZrmXo7Ne4mgw9mcxIQSTQtoeH5VZbqdFM0ZPrNBIATcrJDwRrEewZMgBKet
rg4NrYbaVoB5IOhWzF/q+Vtga4/kn5QG7HwoLAP3rPoalVSnVJ2K6qKXGuL0VqZy/v8S8rlE2nWy
lwFnGyS6HfzBs/Jc11m6jbZdAlVhk3VmYBeEtTpcqjVq7K5ORx9bG8M2FxPTTuMa3hY/HfFXHVuE
r9ox/441YZmVWdMEDckVporK0nMBsdOv21+5WjD0hdHCdR6JgBq3F6qC8jyuy40FL/IK0aDZjk+p
HtLpmXfNAOXmILXsdbeVOPNeFFHv5A2JN4uzXeLSYSA1O4OVddL0oRwzSJawSYI9/OcWBKirWt41
O8wuI+cvpAzbhMVH7rw+Og7FWRn3p5HUavXjkmPMhidaFnmgAsAhd7ZcOYeT8j5DOke3aeJujXbs
S1zEPgKI3aDt+6s5YerZM9lYZVn6k1HqcdRf3GWE2tx+gmFt9L4n4a3ccGlqqQPZ/DsfUVUpRtlM
L9NR7+VQAoXUhHuZ3y53aozdRmylXPBuip96InzpahBZG7ZV3lCWL/CGZmBWg/oeKmmJrgIgIuso
yp6SlTq+m8H1ckLgzw7p0Zb+01DnMtNSVGBwsCRxflikM0vnR9J8cWOJg7eWsPlhrrFSn0ZgTfBf
NfqCMAqI1+KfYrGJwF81Ekz6EOFnVOlZBeHGr5eKGXhoIwemtUcroqeWyUmPbxOVLdbzGUhcXiPR
BGu6P6gw1bpL7krOO6wBPowOBque+zBv4tvTrVQHxJcSylcLlyqEbu4zXt6Gdz4dWZEy+ZPg7/Ya
ADDDp0ctJET0dEQibWtmQy2N3ylrJFFWmgrEZ/ftLd6Y34k/j5n3Wq4X72QSalq6T6kAR+jWur8/
Up0bOtxnAyTZoc51O0BgazxcuPnEKUA5qqBXy9TCWM3HeZQXbYKbB+mdUUljiNziGm3EmNZZBKz+
pSIlEv80iXKbE4nuZY6FYGljVPGrBAe7REvLibAnIpCo4jmlVe2NWapknI/wBm/uL4mecJRmKM1M
f7JBGUjWPSppPJFBgAKJ3mF6nXMiPPO45tF+cCrnNrdrhIbAGwPoPYKM2+jKkrJ2QPFoDSgW3IFY
aICCXSdcwtwcx7T9/ZfVZlDOoSsmbKfYQxAR1yfUvNsanV0r8Bg26ynua0LUmvUlSDbengsbAQ81
sYIrzUyG+VWvnSWK6sixSEL1OIJ98/RI2KNYRpr8y7sOoXZfu880CcrRjUhP7Bw70rbrZs3/ENL4
E3h0rfh/0sZtIDl+eWqBFqosih06VLF6MN973ADgfwM4FH6/V/U0G1cp10nnZNRZEUjxzQM7mpBH
q4V/rn8kU+eB/h2rjkflct8JJtYhiS2uf6italF+MYwVRt6Y07OdjQBhU5+eeuppnDRvPKI0V2VK
8l817DRNRRAi6GcUiI2V2/Qy2LgHxrxFkGS90NfMGKuj+sU2X2Cacs+mn211L0Zaqpd7kwLPboPN
ENBZZqIqI6g7Dtn0p0ON00TpWM/ksN1VdKOy5YK5f2mCWmHfOTIXWnihOg+l2fv90GZszYZ/PB2E
/CuRT/EvLt0rU25IOQRWq3LJRe81DgVXO5f6kYMRQVpPgdXTFx59o9BO3IdytRhD8n/47qKFlQTw
DPpLYk2HkfETmtKY2C4cmUDabjabUyXZhV4g+wscyfSGsqZ7CdAHXDBpwvWLzDVvkCUCjvKXLN8t
0IS8k2X9uX5GW3DroY2Owp5s/D/rpgP6JUEgdJSDYe8WpHpr8rgTzOkaJTTvlXvHCETfSwum3lGu
J+BBAkogdABaM0c1Aur0mXSlUqKc9hteHwBRqHT1n6Ivu8orkFGshU86y4Q9RcoAXr8oAUduKiX0
wqZfW9TRuHgXvlAuXYDpc48yVM/iyPzG/lnfIeTBg6Tu3FgFe3tW8qbCIZiWBw7zMXZAI10jjPTw
yfZwDe8BfnN5UBBZNcJQAzqpi+Iwok30a/2TgzNjSABzs9Ua86P4+MN4um5hIynL9/9yVSieiGLG
CIn1G8V6Z9TtnuUi5amtzCAGaLjELteFUNo8faY3L/o1+Vys3hVSpI4JRRfi8nLLJpHrvyNiGQzZ
bx/Z+xn2rF+8OHiZj0hMSj9IKEvOhyU2Wo1fkUWdCFoH/Uqfyxz7p54s0tXn8K0XEWlTEHvXGNjF
D3s3X6FOvl5Nb+bGaMw+fUkfe2kA7VIQT0MIntKxE9K+athHAQUjAXgSxwRaGmW7tGiHf55FjmL6
TAI3yUDur6yDcJl0G/DrotYUZ0aq9Cw7o+NEhIVmwfkRe+zPtl9S11fropmLYya6Bm8py4MY0OAl
6dE2cS30kvrPmLtzYrX0QnxlXOBGwc9K4oIlp8r9rgD6EFTekpFec92YenKZLLKRfaW/OwwG02Ut
OsbTEIGPpRl6TAbME6CBDEnSWdx8V0RN8BqYkc4mi5pWT/pTazU4YSuOR5QpBUAGUZPIwAB5bv2s
bqsghAj3xC9vdVFPziliAVE19UI+GhsfdSHWyLHe+EZbsiftENsgCUdNu8mABWeW1WCtg5DGiwcu
zMI0jeN7DC+bIxi5pA2UV74mh8khRgj/sxnuSGk9qqOexvN63Qn9A0DmCHZEq01fRv2hLxwzdi0n
CuLeBgVwsr4i7erDITGhDNCNT+S9reZoTFtE/sjYrd6Wu3x1wEBerIOFBTvCtSCfwgK4tYUmZset
7YlQRRGz+buD5lggDgeHqQPaLyphcpu8DEni9ul/yUY7YxJZ3NAMDXcg0hq+IBF6H0B+P0E7U3+V
sNaYoDdvSj/tvfDAX0tlc/bOmkpnRf3jlQ9SJNDBytqlLn1P+TlFiG4W+lkliIXUYFpHd5xlVglu
2wpF3HUrJ3HFcmFrvO6k7Qtm0YOx4zCeQhNS5dy+J5AH/zs1OLyIpnkN3Gsgo+fnzPIJZXesnXxH
8MateCrivbEXVEXb5Puve5IEHakNaPNHf7cUAC7aS59jZwzWgl5tpdU+KPk8BqurGUXfAjRzJofH
8mi5lDlJ+8vYDLDjeiHX1YkVcNlsGDCNUqnMEgtE1PuGWstTsRSil9dNNwlUabun6TBX6ghxHsWd
j7LZg9D8S7UKk5wOfaYHiPipK06frZXNSdJEW6FE5iE5Rgit2DLmWhcJFvYzMCPBFkTJenF4pk3w
aN9Tz0tfifJ5LehYpQrqf4p75Iq9zpMhyvIaCqcJbt0uJ+fTlKoK79ABDWiUaCpvxycZfU8AV/CF
M8zmnKBT4E9dWZ8ndIji8EaKuvRM/2dz0goH0wQnHiKNN8FxQC7+Key1FWCHfxBtfU1NrvIdgXT1
lRNRDO8NuvEC6XjMz4NLBIPF6gRJbxUZdw8kxWbvCEYl1CsSJcKkVuHlEYtFVhtH/MC83+A96eMr
U2a4xMQMLp3CtEDn+hUQdszlyHYE4i0SJAcpYyMDY/2x/UxFUXuw7rrJ+zUT6iXbT1siGCjcvOvb
a4+257Xaq55toYpDlLDTSKIAE5XZ3hv7WRaMREOQfz7woUGTgw3gWXB6wSGkmX/+yaEabU13iUpC
0qPksEqSqd/pA4JVHbWoSRe5gP6GQBh2LPSFoPWVMzCaXR1fokko1FXkY1oBTBlRnNH12Xbszb8T
a55KjpeI+tZbgm8lm3R6h+ZOvkhIcUaZcgxdtgFVwST7PRWaxJkuRM6l00o17RJql53RCG2Fx+ZB
udqU8uwB2U0W0hwdsq6vYJ6uGW8i6NAfC2uexZLwc+s0wuPdCk3+zhmtZoU1eYW2r3V1Z4ZN+siv
zBOxUcYwBNxcK8Hsd/1fb6UAjPUQaGS6suz6BYR2iv6TciZFv9qWvHkfaYEWqHPRW2xF3BIrG4Du
64qJosoS5OXvD8Q5o+22ahZXJkG+Gs5JTjGG84EmEPo0bfRsuaeJEqrTgNoLNVDDp7HbyyO5DHCz
th0fTMbNp2gPZxkFEO+0QW//yDuj8FoX7+klqQk9m8kjj0p2walolUML0Oub5hATzFxWI+4Xfi81
939B3qmZv6PQibE5NERC6gH+mJaSUZieSBzuq2OZOOs7ZhTSo8eZ5lodFbcoR3nRzxhkWTaAvLsI
TYu1oIngqQaiEXTfS/ciKZaQGjTwWAEYT6ZVvMO+ApQFl/DaehxOfc/buMSU1bxGvCC81SNhJ1i7
8TZkLz5sycXSiOp/vvhdXxIGacL8d/9CUxWrgQgMr/qE8Bt10juPub8vFtuq0UrQcjhx+Y0cvqsh
wDZKIlhCaRpxIXXc0LtcNoQZDhXzyZSoIK/cwGQIEL43QR6LE0twsn6SG+4fQOlFOPRiD3QN8s95
g782GhodX5FRICxAZSx9ua5i9sCfCUndzp8dMRflbDczugd7wQ8JSbjiIJLZNeur9IWfzVC5hu+f
tjT2oaT7cVpRdu0cUQblPM1X4wCq5joLCdTydEsfkXAWZba42/CSr9Vr7dE570+/P4uvtxofWW5R
F4gR+LMimW+LtRjBUvV3zYAk3+Xepr+axTtu4wfw2QnyNNt6sqXEi+rN/U6RuoDy4gGi2zGWWphU
hsUFEtguChU3Pcg7xEBBk5RaBoh0ZDkNqOkSvQg6Nb5Lbh7wyHrZgQNBV0/lhBlDtAYAQD5Fa1yO
py1870LRGM820MzR+NwaDiwqXuw6qR87/y3Osx+gSCcn7YSv3/GRgZ4UQ2i5KGzKOITdNkvYRbrE
7zikZFvkBiDwe0SYvwwlO7Sy5CGSpNydWCeenOu+3QcZpLZNhu2qFJ7p0LOYRtQ5r9QsuC41dV/J
9P0Ri0Oi1Q9HaVQ+ecAIBqltLerLaT6iIcoXugbXFRakmGsXe9B6tT5AosJo1rz8HZx1pnzHZXOC
jGnipntRRu7qlvLy46askirkIv8xFswUFLAOW9n0/jVNzis0wc3kvtPQPVlkMznboA/LheUGFTz9
zvQp+qhD3PRYEjzs7VpB27/SrVkVdCM42G0SOz+5HdQUlSuAlUe+ngB1en4BS9tUVAldTzROurDx
+6VscoQsJMuBp3AiKnWQ6qhqSXjFZKJyNeqAPE1FR7HlNvb5cn6aoL1SxnhV4AcaPgdwm2SGB7qh
X6JBDcbInOpRU/XKXfzH9rTsOditCPNE0B0k73yTh2Mjn+QnBfL1LnXu6ibUrZwlff/WdZlR77Gp
zPgdt4js0fgs+XeHoHHKuwx6SYxxwQMDKLZmu+ttK0gKsVGxRCuWzG2zm+lpS+yqTm7P3B7Z3Zui
IR2OilDhymkcRGFAKvgAXfzm9CTIgDbj15Z5I/BnhOvm+5YQWPdEwBHMQsAz02cSkdRYARWQkqYj
5q+6RAaSDM5P9XeP/9iCIPDzjKI5+rmIduxAvUXfxDr6PN8XzFR4UIndTSyVXwHaZhymiX1CXxrj
GbWLk69kfMbAge9qj1PpsS9QErw9K0kZSEOILLv/4MSVXui2fFJIxmFwQUDxhcLAhkiDSdjzVekm
Kv+Q1/oHXUG3L8uUn8kwiuUAjywCB+C6paIGWPDRrc7gmRTiH7fWGxBLWiSBsYtr0TjpxBzakerm
vP7Lke0XiP0qTBPzqoyNly2SswwVxMKN1gnn5utxN8hK/7PGJ2a+TlBleVkqCBOW3xra+3VD5C5Q
fIuDaf/RpDXc0oJlC9tReQgy7VPCWu8yVBN0fBBQ4lD/0A+BNpTbbS3jQ3zfUjckh8dMoP3Q7BXL
iDNI0i/YvEejIf7hgTAr1WEehF+k8aKTASRUDR6KgTZjjr8jCqzUISBsz8Cw7ZFhlPKyM2R9Js3E
dLQFdK+cNdfmrAVf5XhGkS7Og8Bi4qeawL2gNnu09F7DEgvqmDsc9eGEoMCgNAMdLGxqsrAVKk8I
mB2pggvdNVrVOnicUUwrrcx5noFHriqjHZkQbHrA/4WVtEgQN4u2DNMZEg9v0JjduBCoK8+bgCBG
mmO0Fub5JfuF/a++HdH7JlWEFjAq2aAr9Jx4n6pmfS14ZMgtSTGa50IHcRdZPqa+Ty9upBg8qZrF
kzB3s/nZDH+Ga6bYcntqYPdGinytNwZrA5hNfNXFkejkkiEOiwnDao+enkhh5tk93za7lQnkr3QO
0B+UTBYQXolM9jWzQ9aRkS/MQ9dSXNZUngJDy+BGs/CawcP2bIGEQg/A7tVP+Qi9ODQv2assw1PF
4XP70gJT6826gNWT9fNqZeiBu30TzSojI/tbfEq/XVOSWosYAbVfBPLHKwyJixdLGrO/EYguVyt1
luJIodKG4hbXcjreN6857ZEffXFVkTvN4mfjFkwGcffP3QLAiPvt/VO8LFb/UoKhz4lXyJ54IOp4
dhujj5gLGd8vvdX5OaBZPptBFsJuaNoiElAtlVaF5yVLOfCG/9rJ/NZpnksF1n+RQOI5IIXXxrSL
Q7+KbK3iyGJFe2MLZWBRP/Y18n+7gE5f68aiaWbCvAt3cGshdhK7hEmq8jwvkL6UpbqV5HG5nG9w
EHF8Up6SYX0ZbOO0hdH1VrOliL6abBLGvkEx3Tl33rphNfZ0VqtgXRt+x5aCtIgluvaLqN/KBWdw
Zebz6VnNWoEjsTUsO9H4xw905MhFVSg6d9vSbN4ca3Rk5QPljSlRoLgNmmbGA61mm+MMY4TlqLMp
QrWqiRKjlk/zkWM//h8tQHGTCK4khFVUyLub/OaboiPZsGa6x0hRwVCMAW89m/BPKGKa2MmX4M2/
o7W4ZNvHn6QaheOj9pyGGDSgzTqhJYhFBYDoriPILN0yjOBjkwk1IGlgOoh2YRUi0ZvDrSiT4NK3
I5x79259ZuSGnnMF9jINWf6T6TMCvsJ0byBQ9mLOPTwhfDstJQ1QhBiDWVGZvMO3bycE9+Bets8v
RkDdblEDQytK+1ldTP+KEMC1leKQ7bXmyWckzN0H1/F45/+F+LXAk7MYSj3KTAieKmAut07JZ1MN
DNvcuMJD9E1zH1Vkm1QWSN0hnAJZpAsR/kMgDhi4ZvWcRVPzd6TQqJFAxy0U8vPYLACCWqnTiZVo
KVcQ8+m4/RIx6FcIlGHI2Anw5WPsqa4yJWUCqpFhWEz4cXRqUvtJ0i1KH7W6yQXBeY2EhjUEK9TL
AHcu29eESfaB5b+VN9uFq7r+mfHCj7xwBx92RsPXkbTGNYb0vyeu97YbVuuwjmoR8f7HWtYJ57W+
Cuu4JiXLV0JXngUyVqIYwAe+2EmLrh9Uoz73gGodOcZn9iNXWV1/leXsl2o8LDhpF5j4QHqOCkgC
PF/M6N55QyNXT7FTljwVIYYaBJA0vzf74mcik7gLGCXMQMpYdfRB4drSeSqoVRsABkxTfxex9ZrP
ut+Na4exz3O5iy3nI2YQMhBAnnZtYM6fv5yOE/2hCgqKEXyGNZUz5arSA7xMXtxnvgvMlqdLuKNH
J7NSyeZGewZ9qrpo3pSkQWHP1E0jpin/b8TFIj09MxZJHL7TUG4bAKGqQxpGWN8fFAUVel+ozwHE
tLKOibEJSYrJqLiaTlJZay7ap2ekjoDmMuhGfzXkR3+cUVEto1kN1z+0KBy8IL3Mi+ZjnB3PSCv2
pAVDxYH2ZPiCDKpVDlH/ST75z3LzOKYBtwO4DKpVOTPezz5wMif98JS5yeDeXzbtIi6tTXFWsC0Q
LIBw8iuO+v3lngouVA7OkwzqH5yRaTd60lzLXKt8zoX5mlddWYdYtoC24bXoAO7ouRGuIU8XCWkq
ctTmqzf3CGKWQY/izc2a2qQ1x5tpkWD2c1mWja09HRpvFg6/WsEj+dpD6UwRFJxboEECk0mgD6q+
VFQIBsWCtCHK0rRqhDJ6nbhB2dpOqm4PLvvINdmwQy1JjeGeZlEI7Idh64oDUK9wHF6z8MONaksL
h17Q+YXc4Wq3GvUBOAj8cbggScsUyPV6T4w6a+Zqd792i/VU94nnk2ZpiHCL0t3rD98XN7AKKFPV
YfAC1Hi3ufgzMvjBCUjB/+qgbQ1zktG4OtFQditbbO7FCFjl3RIbG2LHuS3pw1w9dO7v9zoDaDyV
RdA9TdGA+IOU7DxN4bKZUexIryR9AG07Mq5WYKynhY3mkGTy87CEV5glC2fQ5T2VwMlxO6op2tv+
IPSXoYxcW7UXzAyOGSZeqstAsgvR4HEphE4Wxj9kN2MIFWh0URqz2D9FcWv6Zzl9TsyuydbOYDYY
c8zVt11NClsEKFIpu+zrM9NKh7oK0xtWO88IvqnO9OobgJBw9srWv0iX6xIk55hwbpIZ1LIfuqkR
I42JHh75qDqfLgXC1sekg822+23y90Wn3+yJWQ45RzwqjD9Jy0Zx4nsbqOr6Lb5z770dVuFb9XV+
FvpBX+iqg4i/R5z84CnVREjqkwPxs4e8cMLllfK/RkZ6gmn3S8aj1NXILS1PN0tUAgdrBy6ms3E/
Qunb2wMbCyBylQFWEKc/JoyWnNVucNtZFebs3f+rWLvys+I+ZlQQaGYyXTN8ay1x074aUeL/I42j
OHUq8bB3AZ9+6AwqTdquzDKhmKIQ5d98ICySWPnu4FMTIKh7SM7GlScGtbyXkDGwaZ36T5wU+glK
EorV/M1br4i3sn8UYgBMDK0aiB0KP5B6tD4Bl1Fe16NLKX1jE4IzGS/ydFDBjSbcUXJnnU8Ka7RH
SbPBbtxBvXQVDqVGuubwM7WE7zlXR7Np+DJ+9WXrcfVsH59rd1kVwZDcl2usVYioOACFRZF+JS31
dp781UlLKj7q4nc2/aVFEMcKLkRSJXjXLpBE2iDZNMtR2iW80iIC+t7j9HayJ0+oRyPJ4Au787co
RJedpRGmJo4HlBgqU3ZPFtgvS9JJFD5pon2346vTEvuFu5BsQp8xIJN6AIhqPWSQMaFcSfU5ONE5
UQcZgiV0CzZBn6itLQokGOnwr5f53HTQ+aESKRPmhN3IA/VjPfxWWSick/lrGqaq7Z2JkaZzgG66
OPqWg7BcrVsC2Yim0bF7hgzrv6mXGq0kH57TF/wyVhRN1l3dPvYD57CYKYZuUidTaRC2dhQqNg+X
Ze1l+IkL2JaCnvbKCvaTD1qsASadb4nmQbeoz8Gpb0UnGMwMjoCGeYhahE+YEpjbeMrhs0Jrnj6I
OS0a1haE50g5vlKPiSRx1SJ2LkuBC3ErDg6ut7xxuwgMnT6aMNPsp5lVl1uN1OUtIG9q5RXGIZY1
EBv+80LoqfTMfnSl9naf34Nay8MlhGTfw8iQUjXBTvJixfAkxhdNjMxAtqhCgdE3OvOgGRMzBMeV
WB4dsTxqi44OnWFeXOo+FJpY5MgxRZReHrA31wtKPrtBXwjV9coTb2ogLh/kXvCAzezu7iVW8CJb
fbeQHqFwJJ4HG0eJrsUqzjlErTvvN5w3FUNaCngBEFtWqP14lQxHeCEqRKSppUVVtyXoLU60CMsu
/524DufVuH/DqUKA5wyssBwFCteOwYrFUrKzPCgC+paxesqlhmClj3nnPs3XkbWiHG1P2htaF4Ds
jp0onGSN4eNIHACIDVxK03i9agld2xyx6XhUhsVeBzyX9rrli/OZew1qIsvwcxaWv/4Wbqnsno0O
z9bCYMnEmCcGw6CgKP3OLrZBqNnCvkzWLOnn+pqJGVF8HwgzfsQq3iR+UqIWShqcN5ZADSxiPgnj
HsJVwG2X7AWslSjkiY94AUIT3fP8rxL53kVkq7gY0JxaWVkIJ5VptQM23RbDKyZLNvGrdCqcGmc+
iewKy0vAbd0N4FSFcWooGwplG2OhfKSJ/xHx6MkK+qBEwGEhDbjlHJnV1krOeeXWGfiHcnW2RTJm
47sTMo44PdKxLEpts0AsnsIyo/bzcHyAvnvtID2R2PDCkSQlzNVmFLvWswKTbMGoXV9kBgSaArQx
9ATmjaF5//XkTRnlFsL+V6qkNVNBaCfjX9vC/MIl5DkmuxAgnYCSltFrwhw3UIjACyhrttEUgaY9
SJ1sEJpNFPHPFSCeSOYOxquDEwCxHjXkZnpOVNMHiKjatzAQEJ8rSBiz1naKqPMOZgooTskHiSzt
KBfKUJxpeoqvx8lin3m7yKlhp5WzCudz7wb8nprEXICIxzcvgRL4n3YY89iVDOl0YWspbxJU3xRq
TsvV0GfSQYKFCTlcV9H/0KzxV1XcNqSPQMN27+nnBk2M3rfEt4MzZ0gnMEov4ojVqZozdt1HbmvL
cVtLbTrya7Op7VFLPXfNS93wfapxi6FZXL9d82vSJUZcY4ZelpzYHJUCbshLYB1hm0yTQP4S2Ypv
wvYTlZYDA3ONmghqjQ+ZKzwOTUeMhkPWOFcAZHWOdfSlTTAkcEHs2SdoyOOZmvzw62uSpQmoH0I2
jT2YUghWbVZt/ZgHf9EVwB2xApSMO4l3is0G9LRSp4/y+MXYCf3pjapVMT5jvj08j/jiewxNqUiK
dUguHAvjdvvsPQjjjL3doPnVrwO4R5o+mgQf4EKhRYD1qXleEseAWZvoU8fkXINYh+jwilZ4esK8
/7aI6/JedyyBluyRf76XfmDdi/EEs8GleHNEsn4O5t5pNn4K6zeju0C+xWeloJm0M/ZaanP4RirC
NPRPXUini/biIomokQQvoYZGG0wMRSFcab6mQKnCYuDbflplyPYF7evNMvrl5CFifXW/SQktJPsO
UxXlW+GM9a0BlIvCe8nlvLNIDIayP9hpfIE0ZfGbp7djS6JEwLqig1tojn7qDC7dS2YFVp9UDBI4
Q5AkRPAtzLvd1C+EYmpoc44jk1sM/jw39aER7Nii3i0M09ilR75YUP0d/rexk54NPgiPJNsZRXw+
jcB3IS6Bos2y4ebnk+ZFNGVzu34cWJbTD9+5+AjJtEfRAbgUOo6MJyGaliJJczZfQtd5FhXliNPM
X9TaHOkyGd2kF+zLT4PNLs82CqPChxcrkuQzKYDf/Nxy11mrgQeCabn92CXKuXnbHBYI6nZv61RM
zicqmYayVkNbONbzuyAMw9OnhnmVcE2lFloGF4+KtvUPM8TYG/dQ8NL3JrGBK9RE0HOp6NRRhEsQ
r7CBlvy83rIQ7InGpt/v4odsEoGDTFqbVfn6+kfsGISWR8G5AmUw5QDaMIenhfqgS2ika6uhAUqc
hH5xnal/qBBJ3MBgfURBvv3U+pXvnrM3GexOKcUPZ6DnzNNGCFjaHWB4FrDmEezv1zpaz7wLrNSw
f1EOX1BoXK1K8PZX3XI4yoEGifIBlD7EAcBPmqDlr2BOaol2wBkYLTII+8qbEnSrDb5BxT00xrv2
wPThThrlOt1yv6i1xQdJHlrVLsau6zOnImi6cNIGTCi1Z1yO7phzUwWz3jKMSMdGMhRTcG9rkx/3
kHKvz914zet2f53QUpDjoJgw2D8RGF9E+3jv3iwIpsUFTZUtksxltzURpg1N/3SdHuCtAWUQwJu9
vUx4R2pJAZN0Ja3Yfpk91OHbJpa+klc3dsljnNU1OXuqWuGol7IAw4vDHvL8NePdaZ8FECyyDMgT
Sg3TK4ovyO0SSCwEV3Ahbo7GvKoyRUYayJlHHVVqZaljJ2MwQ0YrEGhB4zzUdvquJIeL78lIq/Xx
HTT+Fhboks26GMZMNs2tEsKe+Hu7cDpYWhDx9VNtUE9e114zIA60CSz8Q7Koyr+SNXDzOaKtArA0
YKt+ZjIO/baeIg0dPsMepcjS6ZiyxV4EEfnNZlh7IKLO5pQZoN1z9Gpz0pqI0DthlEZn63/7/mby
NAiJuQDvnwz9NH6dojjwquSBsJaiBsNeK21rCaBJEROBIqMD6URnWJKlpzuOzIlYQSxs1hqNwe91
HProJcW4FrFGle7N0nSfJDWzCHHMSjf/fkSLOGWcuxnf3nxuDKJjnuxpi7SF6qhKzgLTXBmqkwPX
nTK37as0j2l031qIr03TdsM6vIAoFIJkI0bzsYkeWY8bBWVKMoBwclFGc1+IWQTIp53R3dSUwOp2
V4btUOzFcs0eLzeTjuSXhfwSz+dypZYWBT3xzQgVugeJbGV7u4BlsjFC1eYejPxl8R06L6BQr+nR
U1CLABFpAsbNKYrnNYLfUFof5NPpeiDJ5Ds/th78Eo+4HU2ePFCIuPdsF7JDRlOg/49QP05pHSzi
htRYGDKIe/HOtrNFUNGM7rXnUMrLXjGn6eSWZd6OiHa26prl0i5WakXlRBYwdSW30HNczETul/CJ
hq/FaC7pMrzQ+2R8aYRhyv0zWVS2s4gcVYSg/LC516H5Sie3RKH546jH8bVDJRL9BhWe1oM+B/7l
HwWfhWMV5J9znIp5IGnsg3zw/+dhbdKjxyLysrGQdgw8jmopC+nXSEz0126LeQRoXv4+lJde2jDu
316AOJ6kS3340uG7vwsnNqlrtC4sLy6CZ38WX23SqP/MOBGc9bcBsRQL5SnlHKC6gHzlVaF2S1dI
GIs7bsJA/HGZtWeRyorw/ZeU3AmrDTKE/18zTPYd2eOK4SJmhNG6TiHVutUe2zN4NZHnZbrM+vov
2jlVq8wDvHQvwR/3j57no4SMrxGMX6dREPhNrzEFUl2c6dcTMMMjdkzCbaUEpKPFdAOEvZRPKEBb
NU3IxjsseXVPKVFkKRq0ttEYDlPca7eqj5RJk39f9/29PfN+mQg+HCN23OgokS4+a9f8WEYaAgGa
i+qOvusEPKcqt9SHr3AOOKVOsezX7iRO/0it+tyye8C9jhcc0CtSn6syegxdomJSPGnArQ6452FI
N/LituXzCaepwwwSiE+x4MuOPnm7DbThVSLefjeUX2VEO5godx4lr2gu042Ez6MhAq7UX/843AOS
JcGnogNf+WQsp376VwE0cWrdVurx0EV7aAZZ94vtOS06Ypb73z0eudXQu29zLByBOp9Y/+xYd8/F
a5tAVnJ/l/2m4Fv4xs4fcQyXwJ9KCjq6CFyMhRBclJ5TM2+vXfQ+nmzCwdlklyUnoLe2PR3SxRXL
2tP8geDYjvYLty/lguU6EqaNS86pSLIGFKXCo3Gh4jLEBZ+lx4Dkyy1+7lZjxfjXQMLCB/HBFHgr
xBRNh8F80SGYGTxmzYVKyKbmvk+7JIv5MVGGfCihMAe0JJRe/OQXfZfaIXUvPKHhtR8Po27Rw8Oc
7QeaSdLfF8Y+BLfdwkHDW11n+DiTK7RaBiR42PGE0As5pmVpmtEysX3A5+lf5ZtkOeWE+XbAPTnC
E0SJF8NP+lVXZM/keNxEhrumYmS06Mxzm050Hq9kQQZJNe0fOmpPe/JhalL/CBJigJIbnyfLBiNU
dErKBxseEHxhbj1anW2Ozl/VhglN4DdHAP/2MWYTiaTVuJl2qGr6uFSPdlgh9IctWzbhM7gYqdaL
VSWzs0gBnGnI+wsP6OguPag/Xlb8EtBTqcahChbeZJ+ew0bA1BFZsveAGaeIgrPGTS1cOH28lE77
DjXMS9BxxqMtrLfPSWWlz6ZNer6HC2ID9F48I7RSx05/RcUC+jLhDr8lpGAVCWBSeCKk+BWpnjXl
UHo+3ma4tq1yn7jZGGPpxblmNkE9R30lIiMEdL5rEci4qkUkn7oxQopmtxCDV2c5+BeQsXA2tbPe
Xt7j8VOcThnrIzBpqKILrQryhOtVnloOgu70N47FgEC3vrUKgLep/nncNUSsR4Z8KNbQI1xoKi36
JO1btknPelhT5I0GA1m7gU85AagUZTkptPlOVc7Ar/NXz3cHs5nWyDr9IhYXaxQ/O2zkhtTP0NQR
CrW4OtELESRBioUf9h50tM7LCOMcJWO2qm/Ec9YL7GBX0QoRa+04ee7k3db8hKtIa8YKVTx7K37d
y27XUlR3fnPY5k5l+fgkpQbqsyZQoavpYZUUYA8TLGxwusI+WcOJBqWTndblP244s1pp6TOmD2TZ
CetPBjthCGGQAjRn7e87t94v1upaeYOEph0acbHomzlxZ9h2E5PeDI3/nSsKVPMj5jcY5kQKzvd7
dc1Dno9AQsbM2/6kpbr+vTmgww0lSkzzjAgAgGEB7n2qI1EuVu+4gXBS1iQEmKcPopiYpyvYk4ba
CwB4p5nAZL5OhukObEzq/m7leWUdkVpqEtCiL5uxQee07q0WkPc2FUZRfAVIV1JDI8xo7Ks+tHQX
4JNPOlBi/V6yo+v4YSTmdqMpfCxs6a9r7em5B89VE6hRImFtTU/0Wsfk7wJjkmN4P/fmC6pasNW3
5DwSXeI+jtwauMcWFfjutr/I0XBP4bPK3utvYKxE//+BoNC4Rwske9/eR/GJOvgPwoGhUebiEp6A
jIlEQt/wfGbfUJgUutRUAsiIAcZHXyNHe6plkFVhE/1AYTrXhuO6Q1nrD2aaFvZLDTgc3XpC7mGk
ZCj4b3TOwfbcgu02uiCyhfiRZT4/nQ7dQA21npyTaI0BIjYRSPZ9kESJY6csuL+KJZpvqJzRYjBZ
0E2Pe5BrCmj0BiZXS+5suKYKMDk8VfDR/k8bQ/i94AJI95TaPpfSmXLKOgsM0rJeoF1GIKwnBl/e
zgE/tjq6cndO1kSrZWoT+zRFOA6wB9teGr7a0F6vB2YQcV0uKfLNPyR8SqUbV3Wr6RfJAB1itrTQ
O2bdJPk6XI82Hd3xnGW2LVygXPuzT3x9HCrFQbI7jamUy02iW+jgmc5kw365Gw1Y9XXUROTdMyX4
jb9QTWsPKYdvHYcbwHHL7TIiR1vgcgvYKleJu9AmuNZxP3WkqMpR7gZu8/5Q2GmiZwKOH+015Wva
XgzEjULPPcMuwy/mv4Bcd+GlFK4L77O/kinshPr0oRhH9Rt6i3Sm6qn2jxwCvPq3ZeMIT6oAMjok
sU/JAEQWtl+qEKxiq8XqGXLnPc3960dmMNTJx2C3LrhzdyC4aMAVxmowb3U9p6MgJglG6fdlGtrR
EI+yh2M6g8GpfhdXoAQ8yHtRdtFZVug782JnVCaPN/zPnV04xXZ7pdvSlZNQddU67HtHrk5rsmlN
62+OcUNOcnn/JHk+3pxVKvFc7SfBiO95OESZ495dD4ZjSInWikiNJ4heMWWc4m2wR62Spj/0AnEJ
nvb717dJ9yToR2oBBY92bBffBdzRj77Ma/+gL/qpzFhxabRj+hU4IkCixL350IBynW1vx8TMsF7Y
7tYq5UsQujeCs5SbDUkLQ184CNWKKOshqgc/TP8LsaoeTPhx82C4gLK5wMs+5/RyiVgkcsOxz3Vk
w8oTS7iR9XgGHXwf4qe4aXG6jl35m0fmfxbkPi1h6z2NoXij4TY6RbiOcMSEvqKs2TwcGqpVfdEw
NQmyiMSQhpfjvmakeimiY72IfGlEqu6ONyeXlUGcVq7wtVHmvfcz82ZpssIxDTjRDUNvnT5gwmLv
MYrxEVENE7NTsHiSjXrq8oIyH2hPO5CTtlW1aXNA6hjwuK5eoqCVMWmOGVvq8mQ0z0McOaDQ/ykO
fFG9tDTJ3rIwDJAJotN+asadsGFRGvB1aDHx14XtxzYmyxy+hCCoK6frQ8+/0NJ7UDxT0R1KMMlG
/Ga5cDM9G22d348nuxsv8tW+FiGjvkDAD3b0zL9oN4MuooqiR+B99yst2Hq/UUQ1ivepieG7Y/u7
gRf5c7vWyWhRiT/O3EAoK9fB/0XXkoFK/k69xJPGTeQ99tonyEV2Dkp6CfaRI+yKwawg8oTWHGNU
6hOaJ27Hd7SH6X87QqrVDmGTTkOmxCBPl7Xtxsiw27U0qIdgnRu3d3Xyc9a/0BWxjeUCDXKPLaB8
Y4bixhk2YjD+P4GFXwIePwisQ9WTL9XOgkqFTiPXGWusv+XglyhwGowqj8Tj4r6vW2ix/H+Z+II7
/ORpj6+cKMc4oBsIMxX1OAa7eLeojNKs2v3wzzi4x5bizp01lqjg1n9MMUPSlwEFVeRD8Z5WoGkO
YxNE9mxf7fkUMT6Sqyx4vqcMPzhRaRo6n3ZcdaY1pkGFYZu8ZneBfi4+rk+Af72K92q3uhTnvasQ
3436Q5sXNe3hAVXJbmci6XLawECDKf2g3I9rmBKrNztHdk8fTmI8KWeC/CiBuHoXVkNQwmUIrd7E
JpBomjjFlN7aEV2YdF+1Ft0GDTLo2tQIGaVYSJDDX3cAcq0dLxEQiqbEGeDgStDnQDLNeTLi4Bfy
V7SvX9lJCb1YKooPYN1U8LLLeXDTXFjd/P/DlnF4JeTnruziQFuRdmZrCAfvyrL9+TmjQ4RtJ7h/
dahEkSYkE3HN8FvPwg/GVXqKBCvhuOiH1UAFHfOCSom1Ua5rwrYsj1Bm7QzQDHNAPGRHK7+1gy29
D4JG1w6+8EwAaTPo7d5m8Cb6cIDtvcaObnR8KEvfPUh7nJb9F/DNg4fOH/YOwbebWnmZ+RDK9V3d
nc7FtEhMwLVHaIYvK7neb+VU1bsERU4kobIh4HBx7klzpflki21wdTwzNw0z9R8Rc8N/46svawEm
oN8T6GYsk3PROrB3ZwG+gDRFDXPi/L9tmMO7aiulu11L/aOOkVllufNO+40gQySE02pKd6JFyrui
k7WGnFkzanbCmGTM59Tyk5NB8nK+Lm+xZhH4MIV/yLCnkHHH4TAxVCBFPGzPIvmGqrNvWZVyz/Gz
H3kaOdKzeH0vkTKwaTbKPnIda63g4wzarkq1kGZY8YF1hmB0ib0djPKVLtDc+VugLhbHkyyLAx6v
LLBgb5e9/m1pVhAWzi4Qfc3Sw2GoY/wCaeXauvOgj1z4nCOhpw7lg2+BO0u5EJc4T1nfBcUPMVrs
OgXP/iaSc17DPpVSYn3nv5BkR4QBObGWv3BS61HO+ZYgSfNyZZ31QQdeQNvKG1D3rQu7c7V7Psk/
XPcFvn+/jVobPAtVHAlPCibe/75beMMwMY8YABaXD1QecsQz/P494FzDOXEvs9H28fpiyHJCgIS4
fM8+HoWlOPF5urPBc4LH4a7QCktSjhc/USFGyDv+F01NzcQN1LixXRF4O2TDbvRzvvtLbKvnFNf0
wCTcO9dx65k7sY00KIC4GbSKKPaxjtcn3Utu74AVun8kzUrZGf9SBo2zN54c6mZrrFKkwsM1GqtP
BiEqaztX1WcrJCSipWMbToMzeFME99xFBkr1NrF7KCD/btpRn6Dl8FEKwfrXnKaGkkBF3NhrPyWA
TpO2dPPNTmn8axr3ydeXl0gJuQ3FywBjcXp6wbBbLgj1fNMVCAlvtVc7GGEZzvEjwGFN4yhHJzBX
OmS7OS7pFMW2Zc60/P9sFrJdhlhECtDxAdsIlsPkrnBbaHJSaeNvjuF0U2XsMibV9f4hT6P+jhm0
2CUK5LnDHXMh1A+DnYZmJxDV3NNog0hvOkpuHVSoT0YgU44o9l0QrHYvF+kgdN0GEnMSeP9IMkKk
JSb9m6H8tkJjl9PxKBOd5eL7CZgPqw1i2UdQJxoUHX60udJMzeiKrteLDvlw0kCND6IeCoOX1y0p
dO9i9WisGCjrZ3X986pHO8Pu7KLGMh8R5qhqz24s+i1ZJYEQ2FTkIK7M5hwU3Sz6Zerm5Liz8Y5i
3neMg7+SPdnul0V/Wd3yX58858gml8tLWeiiHQe2PoSVRqW0Szq+50l01pwVbpQ6Fz5Cq8EHMaPk
4NLVn1mRGhwaEHZXR+TwBpCMNb8mPoCNWbWYVByDDy0oRss+kaekQOL6cWN1rw4cO2RVzqlSSojv
cx498a7flei1VFkvJUFASW7tEsZQX7JuyYFCisPr26GaDnjIkk0IiP6BmVvoahBuG+h2Wlg2uV3y
FCHAJTDHOChs6jwBYpQrxmJV05O0GA0+j8qDKObrhfgoK/2Hsbnolb1rWq2d+9qyAONNeCttRzV/
RhoO7evfWWJave1wj/Blu9Re5/aaQ5OTBUQapIOJ7yT+kUMzXR97mB7FyatpHUoA/A5kzqSHd2fi
lPBDfxgyObenEP9kIJtkzDai/GiSCdkk1yk5kEX3x/gzciUyUz6MMUG5A6ttdQOPONX/3Wn8tdh/
GBBZyVkKT6EMPfcRFy1iMxdZ9YSZGN9ZJ3r2rCaVUe34rc332vN1bQCxsWUNxqkabR/g4DSNO1yE
P/1Ep6KiiVGw4Ow3S0E6uhBA/MuFQGdQR0sJlhI5VIB79yz2eBLaJ2Ae0ykt0r99bQgN40gE0Q0L
9/1Ju7SgBiSOL3IebIaKuKWLq7F1Eo2TuL7U4PWszUQCrk0z78v8FVr42OI9K5obhOOcB9L9aUFO
rGdkqjME4NaCajB3Zl6PRooqy7+OZ9hKbbjST0GxETkCy0Ke4iDwhfrD7jc84q7CXF8cJ6Rqfp1s
CRWdD3PD24wD1x/9Cr4bnbmkRhRoFUnUD6zdoUsM+lTCMGtAKkIlcjfOr2GwIStH7ldKElu/5X10
t9Pbzhwx8/aDDUeOBZ+Wu/3blZaCZlZYOcTfMzJhnK6WyeNSx/MEVKHg/QeXJPfWZEuggNsICQ0c
5w5CioW1XDuwy30MHUUJXE1YsSwCqo5IEA2126YmOc1ytF0TZ/vpG/ollnoH7q9kIxFxU0vCNh8K
DBWvmlDyWk9Wrjq2wqkdlHn7s+QtVoiWiLwT7bqAVLexp2IoIxNRPWtg5EkCVncPZbRje8it85e6
wIbkieqH6520Idg5VVsPgDlRkMXbga1czUA1ndpEHKLq31vhxtAaH0vqU1XfaTwcZexMxvkBLlD1
3JGI/T6NUuLUtcWutFEYqmkBe3CpISBumJyHiIAansQVJYOWl2/Vs+L98QBvYkvftAeK8qYqap+Y
WQ/i9gsXTmEI6bkFPaBt2bXm3FyGMvXoVjrsB1y7UHRI9zZF89iFF5rBNZWWPnUqou5XGFn7LvT2
Xtb2h8GsTLk1MpDsuwcVJ/YZyaZeaUVe4pv2BwloMq0KqTidjrPTFUH1U/8E6wQDjqNIhuWppHRH
dJpF6Ix7E2LIjhpSS5xiio2cOvIBEe+K4bK4/L48odjGZWzkyMKRK9pdKHvIxLOUWfVKu05ISind
v6DJ9ROG6C6P4CkIr5qZ3hc4RFRSUMg/ls/YEFEu9xd/8BPqKyEu1cbEm9FeaRNHzx4yqWQjcLoH
YPM6c2k2+nRAY9V/bm3eaq8RB0BM94l47qnpPTpJ34taio+ybRi1fTkP7bAekMWfNK7RxewDE/NS
46r99+UrVT6xsdCycZh2LyN/EW2l3kWvscfDgTANkNjrqWBQ3UNY4vSCGxSb4X9jy/W+oBmd9C+1
sUg/UkPUUfDWj01lvVnVknOaPK9HWRegSGP86vFnrNtRkoZXyk6E//eXU/rBgItCGKYtwTAWZ0QJ
79TEUU5DQOHkQJ0BA2Fz6uu0ln3CKYAHcYCBsSgXN8I5us9KFqtSRyvb3m7pPn6QWshMDW6f7jcm
xojm0nD6Ex1so4v23uWtd0CHUmSsx8mxgNtk6FIHSOarNZt9O4UCZVcQ6sCvH8IPmLTPBjDjGiDJ
UR2tCl1Pp3F5hAshFg5dIIuM/wfOcxYkxf9qetycu8kjhMY7NcGhdR7YAmbPjfsAxogRLthBnMpa
a8DqlTsXTFsYOsmp181ImB5c/hhQX3wgfymX+Nbvs1az4N+qbQZIvfUGgDzF36V2sHKg1bHQT0kb
Yivw37NR9t+q/Y0nWVjNj/+MkL18HBOt3ZKC8gl+agv1yEfW8so3B7AV7icZavZYCpWgfSSUM/5l
nDcDMxKoVqnU/5wXztMgmujBtdNISNKXr9FX9zbY/274RdVOq5iS1zdfJXtwW7hc9RV0foVCYpe7
rBRTVqpPfsVG05s0QvgXkj50NrrAPwDOXVQGr03qFDMLp7tibSHWrUuIXPE89xbLaSYGLJxH7fKS
unnE3ZCOsiFPAietAo/Ylcl34NfPVos5STf9X2wjJFDM2qohJLsOmQfWOxAGipW0/kxx8+xTu48/
vDQcpOKmba3W15o/DKgI5dFDnZQr+yEPH3bcflxEsxaLXEJ423WnQelyS5LJ4707/uBT/ngjv9JX
LR81+zd/CdDuewlm1to9GRHU3Qrfdr3MOZb6JwR3WWtL7uI4+YmcAtAQIp1eJrhyiZHRoTvrhJLZ
BtmhA+TfUclo4y3lFcw7YyKU8WBbML5dphG4T0PTZjiFZsRBe4JPCr76O/s17nMfYFLnMmEHPOtt
yNifR4K26H1clSbExFBljf1A0TNKiRwRoBu2tHqmHJpZWtf/m2GGLF2fgb1KNydWKTv21Hg7lyPu
vIm4VQJL1QTQgstt87nOv4hWnMtVZcYY9Sdz9oU1b8exBqDkPDC1MYsEb1kAYbzd0CR0RmgloipX
Ory2u5yZ072eC8mkciXHmXOIi9BsWH6em6ZhBOwQnIiinDEXAHoyspYYx4Tsa1x7SYnU1gCr3J2G
WCOBMlnxumcr0cw1mhA0np6CQJQPVDAdlzS6xCvN99HiIlpou+DKYew4vsev6/mXi7Wm9hxaaRvG
EUIDFcYhc2V4JnhhKwFNfsmJ6tYy4cmiLFruOlIDR+uCnyTO8Sap4Hf26PFAaDZdWG4ou3XCT4Nv
pXMIpaO5WTV8E6+77E5yvLTplpC4Y2kHjletvtOowm7OG2LWh56nHy9q4MzcEVnXIj1FT7TA2JSx
0xSRZK4h1H6n/hWokQV/d3gqmWmGJLskTxZHGFSnmt7l1oopnrJxUzOlhY0kr+F30HbEtDBV+nGL
piPaf/nvh8Gl/J63hXMQ0OoCNuHUjZr1ERhBUUqbi6O2QM+/rwC45FkeL75jNkbBsv9gM0LGnzSo
e191pUKbeqZ6hbd9t+/tUWestBg56JCidQTsVjjfg4egGsPIjrYP1GVklErGDLLowXNEmRRZi+nf
uJ/RVrBv/njzK/g1vHnJCLL6vUFQ5H6Xk3l+RpKyl3H+d5w/L92yednqhOw4DxwxLG/q9GEBpVI8
E+oQMPliem61+YgV7uhyphfH18ARZDwwwy4JJdE7x37T5/yQ0Nh6+n5412CFPNiI8fCNPHJZkk7p
3CjRawI24uJW+9XSEhd53op29Cl7T4RD4UbFGb2WBPEjOURiTatmfyvyYYv551ULrXjNfZulN7kD
Tr4gP+xd7UhaJ3oAc+s/D48QusJXf4B6grHIwMgMntxRsfJRWsIZJpCdSO1Scbss1IbAUh4D87gj
9q3dlO/ZhtCigdXb3Mn7VQemEcuS+JGuGXSoeNs+8fEAUGmZLDHh1ar2caEzzrV/zSixeMVHaXAT
ffGN69fOBkIbrbRxUAfmSd4LreSZBb2xDAVbdB78WOsdcikGpURiwExupPdF1duR1lNB2zPdRaEk
k9cFKkdC6TRX+qfLRRZwE7/aXvKIuvmt+btNx+H6LzoKdZ/v0GV9oFK5RMAHi/5ixa39HZOROZK9
Vu/ET90hpy417IZZMFRNPP6v0g/G7z0Su45xWggD/lDL511SM/xsbIdomWjvrx7Sv8BMuPvi/ru5
gaC7lK4SiOa9o3PRxCFt4ey4dKE+sUpALVUHvPY6SrEGyqKvfsdZD9nleHnLlTeMj5FJ7mfDuN7G
aBo6XRfOuikQOlN3amPfTH/8MMQ7b2dracHInJL24b8YXXwxAEI5AqQ3T/i2VMW2IPISpx3wREBo
b13m/fmpApYXLlpjTZOZsh6YkBldYPJbixRk4/zxNUwnd+/aSwdfK1gA/rTZRsDXAm6vDYfz/ZPR
6WykUUqCkWBs8R64PGauFd7bmNFVg4O5Pv95WyROdjaIP/d44F/1r8U20+2rhwag8vp5SmEIgT6h
JqxozuPXKba71JzeJ69TPo/P5WIRhcLZvRwTCWFBeSjX/9W7QY+Q2JMqnU45DbNM8+43WUdLUgjP
QjivyZGkyMz7hAQdesnvSRK8wMKw24R5n4TuQLQ3ZzLoDOPzyyj2r/zwz5MscXIpM0yYKeY5fm2Y
tubzjUvyTCtIB8Nimu/dP9jICPgpGCGd99yr/Ex3HiOPVWuKyu0ZUxOEVo4ryC2Vid8QXv8wfSIr
LT9X7Q/mrM/oWgilzTo4y6cLJzcSxYLyTO4Dj5jld2qHDyfdPKWtGnUCCMLTxHnb+cpMpKBcJfKJ
RtNzEOF3vuJw5gv5O2QV947z50o2xnH0e0R6QGelth7dH4c/xAtyNFrKwfDCcltXicvR2snAhl6t
SkZ0RGaSdCpEchXT8E6Qsf52yEFLDYl3UCnDYudfhilImk8II+5SBtNqqGln1dOuJiG9ePNkrE86
TtryQ+Xl96U6pLHOE8qSWNZ4800wg4jzA9zix0M/MGwiyAUioqqb8gtgX1qAE+gDhEPDmo8GnI/+
Fo07OBgStnQaZC89fVBU6l/3o1eq6hvLoZXp4TkUl6uZ0W2vAXANZwfzcU0WFis4KfMbVQwaKKr2
fvP8DhIRWXfvk6y+LncVrNhqMFCIYL0uGDXNMLJVAgBstECqtBpXIHJ3pu1US2t29xS8H3EyQsI+
dxlrDuDfkUerl2sB4QqubDBjMa7SNcNiJ2213qy+5dv/HaV6EgB/85rLJwOR7b64QT+QTFeVkDGs
qJ5qn1odu4LmecIk0k8IUawKahdX93/MMYYvIPdWtrCZWa/xhqmZGIJx1+CYunvd4FPllWiGqgw4
r37G12bBDjs5LyO/wIM0iYtzIISco8VNFvKRtD02SG9fn2t5LF+m16MPJRFiMZRRdnLe/Ckpb5RO
iXt2MJExb5UjScp+/ybtjyc+2I5t3kTmHzmW5p6rRhZaT5pu+9jEhc1U6LqFgXJgoo1Lhif8bhil
mB+s1tIV2A87S+OhoYxaxEY9PPp+6xEhdpeh+8BuVFDzRoITAtDyocH9kuawL3PcPvxYMi64mS72
qqdQ2cNhFAn5770pSYvm/VMb+5+tvnnGX9p57ynjDWUV9fZLYffRyMTFkiuTnDSwAhEEthDfBk3L
YuTdql6rmTuyyXg6A6nzf/S/NTCLBX2M5OZWPuT+wBvaB/ETqrXp0nPolZFt6G6vvButj5bbkPgW
bfegm9MzIVH8vL51s130Hpxi5X9HfuXNduQWLYPq+Ft6sLfbZdVVSO7y2KUE8UwGNseM8gHtUkbw
TfFjVtUsRzp1AjVt21+nIdraAObujzo7KqLEPjGX4x2Cbe88kfNx0yNrTHFxxR17ol78ExlzVc9h
bwZCmiBLemJd806SU/XJeFhvt3VXAYERpt540dk5nLxnaS/qoJEZbGq/l+ZbUD2jQQmzD+HHGZ/M
ee4C9CGuPIVwGQqvXza70WzN5akIYZWgFq8YJIS5BkcGxKt3Iyc1AG+k4JoQcAuRDiWIedewn031
HyKzD27AsR/1qCItAQh/vkmx2+o3ns5AU3MTP3OT0APhUHnm+1a/lsW42cw4ZkL8Wb0f8EwmVQVr
NKhjdpJreICYkdHgSd8XsIZpehrdzkC8/wYduqkU8aXZRaE126TU1Vpa7Z0lOg5zOgenbxTul7K6
3D990B/8kBonwfGT5j3YcZNTSf+432FV6nBLTkLB+COYJ8m1ePCkjMuQOYdZoAA33LT1rIMpI2RU
kFJkRzfSk5FstvpuZn+dR2xcrnrmeNfgxyndpsU4mZhLGP79nPVjiPwVaqz3Q4hg9Qj3c79t1SB1
uEL/R7hf67wSZ8svwYFrgdl4OfpGbfTh3VVoyd6EBVa4A06b90w6D8p2Fk0UUzPHajd5aBjfVeri
YkQ/TUuJ41CZK6aRQyxgubniH8Wv38l/m77k2MrcHXvpKsVryYOe54Bi/6Vt3hY+KiQFypKWXnTs
OlTwUU1dw5ruE2nZ7+ua0+gGV1JSGiDtWjKRke+0764+3JJFT4VKUncq/A0SGb2eBYwCAg2wZN0f
acGfw4G1ogwOXK+XVLZGlfA2QJGRYjhY869zQZc8r6xj5fT3vb/ig0QoBZ4U0oqw9hqMr3YXmrJ8
WKCPLqLYf8vl+TTeWbfLIgcmP0TLa1Tq36ekF7F8XeCZNAdDAzeJX0Kh8228iyyLm6x59JPhw887
E0VnbvHn+pK9GK5bv4V/b40kijOz5M32IF2w7JnQ7/qh7dn44EF9ZgPj11+yVZM1h42yP7IMNv5r
1PnRLnWq99JBbTBeN54I/eQ9NGRGOd4V+dP6/m20Nopj7AFP/EkaBg/B2ZC2Ri2QaGo2WxMEhO2f
lRYu6QChzgKLA2CoVl30ahaeEBfHfGwqko/gmboBMyGWKhP8V+qTLRJ04bE5TibLrtVXnwH6xX6h
LnIlfaC2q/y0lfVMt2knwDwi2f4hIVVSKOuEwsltp5o0xOzw0fGgE6bOIBG0xfp1I+zpP6kLXkEM
2bi0wighVzbDKbdhS4ia0ef9QINA0I8mkXiVij4RBeGOp6fujNpq+I0c0gD+dRSxah+qXzWXWenX
dgsuIfWAgsHIv6GRDuLyOuMix83GhMk3FHGTO9eaMWagLAvfUZH3NFbz645+0HV0OvtxQMpSM1vA
+JFL4KA/GiWNldIl8+1Z3G0VABvHfsuu+9HMn7DVMIn3Wg29Jy92pDe7IuJ4JxkfMy5b0U33IOpN
PJW9+udJBI637MHicRq6A+ln22BVkPil3omqeH6L5QE0FhK9b5u45oR13eKcBlEpTcZ4ZAyUetRt
SCk4ujtaz3pEmguEOX+aMi8B9Vv62B5/BiozrdZWKIlRw8+88qgDtu4RmmmQUk/Kw5VHq5IOnC3e
s8zAGJ4yA9P5QkZE3mDdnvvkzTE4N0nca4fB1gqWXjOPAhAES+hisKO9tlCNV9FCGjuXxKOcUtzn
K9HkTlSp4XANY8Vf8SkLiLLEV9AeYMvtNA6ul37kLUpNeVQksyAU+Qa+GIaNqxCO9CV/0bL2IjFt
6aM7wI5pQ9xnQcAFt965RvOYRmTZlVUhrzdN9eJB5+D+oYeQ0hxwvhprLduDTK+8km7KYtW54Mdt
TVpmHfLw9R0VNo1J2eYdBGBZl28cxErR6nlMu7qT0yUvS90Rn3BaUzO8zAEwpo+JS2X+CLcMIlgN
cGO+24q9oHnOEv0RNBdbgBq5FNNC9fRJWExZBPA6OBFGMj0imFTWW9bbk9lUqfDCvW4NKydkUbVa
X2lBudtU5+wmNodsIapt+nHhGWhggRcpHM/yxGyheOj8jDltaNBKZ9zq6j4x5cSROxF45pAWZKhn
G2aBCAz+wrk62/v2/fValHH91hzzJwojCi0m3e3R4t4bNBmkii3iW2NxvrDgKp13wu+Ki5tDnWmc
rvqymqkIHAX5K+Ffp8blj6cCyltrWD42WCVGNG1F1b/WOXeyx+ijokZHy5tKY+DvcNDmem0codjf
rMWyPfGj4DqPJycLhAYMJ3ke+TTAbY0YFhEWU/rYEhr5dxZE23wmLSwE7KEI5Wx9fN2pY1UJvQnp
xUeG2M08iEr7HOh1TJo52ecUF4JdSQCYTyTKA7LsCDAHA0Q2tR4MP2X73O8rLsMiwVxCeK3X/eHL
0TVVwcca/nv2Eg/Go0V7xvfwIZORxlGos+D8pRgUtbg3I2lrW2TTXFSb40kYQzd+Q3xrlB44u6o0
MCviv8duBqXf8XWeKRly3G/+6ulWfj9R/17w0v4FXLHAx4IIcfuDYMtZe3GhvHSOdiWyVvgk/jcQ
cEXShNpkxb8W20IuVcRjJmq3I4q2NUs9C56/pkOO9NIkm1PAWBnLuERIasDNn8EUpBwa5+E8YWFD
Tx4a0LUxZwvDUCLyOiJBR0DYgpb9Ak39ZtdOxi9hS9aBmszZgUREQfSmkVgP7kmofNDDsmi95tBQ
LxNHELBZyKiRk7lGk16Wqa2bCLlgvd0+0mFzl6QcwX4AoKphLu2C9gaBe7XpUVIvsCtKVcy/Tolk
K6GQEKjkMlzcq+IIP0GTOxDTHbKg5K1FwuA5jqLPZsuQ90LubXS02ZFBCthDkdcpjBd5+Ybz/awo
W/gkFkUwrtkK2VjIU9TCDdhtKFEkj0KnhzWLME+/YPpG8jjH0fvXRdm0zKLlxC/37pVYt6f/shpW
V76YODTByZbojntzy2QR6QwJmhLh2tlz8PwR2kbJbFDrReqND4r7B5JKVWRmHzePIKz3mT/j0Eg5
6eFD+uVgej0o2/o0R4xJU3qdY/uE2LeUlLIJ7z6DDr9YSD1JjAJf2cxVtnj8yFSn9g5dtwcruXc5
MMkK0oPR5ZHu1UdhPt6NFi5f8kNv1TZ4SBoEtXaStuq/ZHO5sVDiAlKu9HW7j5RjVVI9m+YJ8WGq
D5juKWhUga666Sp3ljSZ5IoX8N69qsXUkrcG1SQ97kPmq99khIO2JRiUzASomkSp2zlXphRThUQh
2uAhVNObQN1g1GOBwOaeLrT/yd/zpD+sEVb8t+8P2Vllk5q9VqgrEW9F8Og7SUm4ghkrBeIt4LXF
2U54mj0FTQdFGwvF3jix5vAKUu6kpq+/+X0bTpgK/53NEvK19UAg2lLp/9qT9Nqd3FrJzOBAGZR1
vtFH3qBrPZAcy7gZ47FuwwEVggk0IAX2/3hCZ3bgtRJtqaOZkG7+lT20SCFMAZouX4DBQkgPEmF5
xHdF5cKD7Xmh5+nbgOOqWzkz0D43ulPy2jYX9JkMUj0RHtHSpext1EzrAGyucIUr4kX0IDgCbe3j
2cbM1+eUdNcDdfyY+VPYBBSQuuoefNQEIOQV4BsZWgSKRpKhJlqKhS8A9ELjDbKMjgSw7D8XBi+Q
kCYTPnVOeivQQEBcNWRdKwxMICmePIoy7Z04z1Tty6SDqhAFgWBpc+1lz4vW8J++rIlK0UWEnKhL
pI3D9FncXQUSDkeFgdwgVADxnQCvFojZDRhVmQhqqGBp1DsTzNqAk2NY2K7bIjeOvBhktNEk1o5y
LBeHyOp2qHqVIytzaW+bxn+OxFtZaU9NdOfnt6SU70gGYnsv+vm7X0ttOSKH11lwCbf4FU59Aasg
WsPDosjHDfyTwfgA5NTyfxqs8U7F7wLg8Mz3XrUAr3SoO43Id7MbvOtGspWTzcHDU8v6Nqcmrnka
COaJ5hUNnQSDE2VWiaW/zbG14RyeJ2dSxBgewUxKmT+8AiVEa0zo2yMJiDdF3/HEaCAcFqcSw9fT
ktWlU8vn6PJIiDg9UNI7phldjnEmuryIzJ4AZJNSN5iQ5A+e3Ljyifti9gvwfaabKLZJQN4LZPm9
TXR0G/rObEsUYSeeAW070ztqCwZya4OTECgc85GaM/Z/bwg/StzfTDhDcGwgIQgXDpaXSBMb21c0
+eTVGxwokIRJkaoNITbY22XcDnbuUjbv8ZQHdj4qGdUc/Y88gF9x67CRrEvOyvgygvyfpjrnqaGo
YUwQVqUeOKIM+Oy29/bY53Z3NU7dPMSQDQGCNZM9vNdk/FIyXIVUcQPx5jAIXsU5dd1XkAL0CUXZ
kFFkYtCC7EbbhtP5PO1VQQIW5VoqOSSQYBdwInzDd1/FugY0FjCgKYmD5xqdzegUKRFHdBF4+rvD
BF4YdI1HYPiHx2UiZ+IusSJFsPeKj4B5jYaC363s8OoXH+ZU6CDVrEowxL32nLbrLCezENZNDOQu
JTxDZ+wqgYC78h9I6yy3mgmZ81uBVgKdGgYkUi9yyoZsuQZJpQNquTIc3W21CcjskPwpfrB/pHcD
AoKMcrD/bebz3P2O1VH3vpUj2Fa/XI6s8bsnBjoo/dXsty5B7TuaLY47+3LaarcLRy3mAVJV471g
ZZCRzXz5QtVvX/j3rKGHmBOXC6SDXA3ubQ9HjwHffnoKiY/dPVp3b9UhiVCIF/K3jJP9oROXC5XD
TyxIeLnFhhrwVwlQ1K1rcFVEgnDu4MuUjrJcrzOvlcnU5+9FNquYl4+gJrPXlMwVqgeaOk2Zwgdo
BvMu7UDfM8T13dkNK6J72jX6XFRmZnD7pYm1Yuausifp131L+OxdPrdg0/Qkx1UcZSN8UHxeeqQ+
AvjUnjLrGnMFkY9aFW3EkDnMI30BLrcRQFjo4BPCWHOah3OC40TEozXO0F4LaKVVFNd1mmTNDIgm
gH9nxE2+dxMoRJWMAB4/VEgAT9pVLh/YJUKB6AtbK2RWW/JuzAqY9T5AmSgO/D7fdtsufNkbUcAI
582y01zI917xL6WzjiFjcA80tgkc7kBct/v4W/jBrfqCWcUw6IGhN5mIJ0bh+fiLiIvEwFIm6ihi
mEyrfI6PlWqT5gZtdUiZjOWqX58AH5L7pxOfP8gwv4TttDtBZvbV3aWLcmOIiNzZXQI3okZ+MOkI
264xSJY+zvNlPuFpZsYa88k8KJvU/ra7WLMUo5WF6hguaePGZyKPJ820+Oq9om2oab0IwacMAgtE
J59tBNv/JOcCQXWFjimqaz0UwqUexj06tqHAsSbDJ8H3fiys0YwPN1ql/QKHGVxHgDDX4X/88clL
/VShm+saVnvW6glNbuOszxI5Pn1/Whgt4sxrxW6DwjSCsAmmGL6jz6uw+IrPfOgM00dMw9DWh+57
+Dnc43f07YcDUR6C2EzZJ3DolJznlw/PaYNmnPGsKt4Pu8GQSjD8lpbu0vt4AJgZivVVbfPOTvcf
VW5XxMUpmMOtKhYSonlCAnLo9Aib8/nmSbzx2uviGjbBAJRhv2mTj/c2bCUPn4cLixAMjWmNK9s+
5IWOlq4sdlIi3U+PCKiwLYUzztU+FiZ9/cS2IooXeQlu0ooKCCLiU3jC7carfobTcam5Pi09rRhE
X3Iv6R+RbZBRK2nE8W7/n+ZWFVNJ2OM5j6WgphMHXjRWwkODa0PqPTGNpQ9GIb9RFcjbvP+PPBhO
X99SZPYvnNnr46/QEQCuY2ICRaqAgZ9aKG3Ou1FrEnGcLe3DmRpFv9jn4cfXbSIvRX5kiNSWHux+
vIK5IqqGhTEHh6HXvqQGQTh/CyX2hXd9sElaSFv+myzXRANJhbEVqZayJ2uEzJfBOWVPPZpPR3js
3cBcz95yapxs6+v/dixX3zvPRd60SiFViSAbwFHkSOiZkrypKVAo9q2Ur0Kn7ziiEVw4trj5q4/s
4HIP/TTxUzYQ7YS54AJCsZObSTRnJi6x5mQUepBwDG4lpFYxuIxrixK47Ev5QosTUooctNuLIbwz
ROZ3YYbdbm49bbHcX3jljcTmgZ0NsfONfcZgDSbvpro8YAFD9qD30L9XFLoCJ/IV9IidJ2UxN5W1
X1B2I1NijOR8KO3Xr74+eB2QAr8iwQ+9W3bVBpiDGtLLCMYv7pjDqJktbCxmzgq9T0Rcx5/9Ta4D
9TGbOY6S8svoC6RQtfKRu7/KqxtoWtv8EzHYzY9oyQaeZLYvAcYjFE0BKEXBabfm8ZdXiVQid9cF
L6kAvlEQ3jkid4epVcfU0OTBn/epI96vRyDTroPdtziBGO1aPJL39cseUUG1YiRPxagfkN/v5YcN
HOXYyWUCDiYV68Lq78fo+Dg0t+mUqkJ6YIXZOO6T4Cm3lgbgXBKuLLz2TZnIXkEQbDlvmmG33nQJ
JSM2/c4moiZmcWbKdu3G9spO/JncZ6ndo+E5mVnz9rxCq+aFjw4uI0Tw/5TrTiFd5xO/rNg0OHLS
ioy+eXOwi+vcY6ijPLCxpW2IKDCx3w8Ikxwyc7wma6CHIyofONgnXmfq+bTphR+JjjzqjWCyhEoF
lomoJDz/njBCNQbNzk4Ro1CyMFCmXa60sM3bSxXsGTHuc9Sop/8bRkPgiS8dJTLTDpaEGCOp1ZyF
gLriejCLJzpCB87KW0mn/RWy86HO5aOIlTkszUPZe6jlt6Djo/Lxi+yItSPLYWYoKfbqD0i7spc/
7VJp04wRN4CzahWz5f448x/At6sLCkrWF7PqLpdFBRx/8HhN9nXc2g59vTvuxodaR7s0YcR7ZFs4
58lrIewfo5WDbFOxsaDG2l04sseCuWKXbyAs+v3H4Z9VQpTelVfvS3RkcTzlaN5XLX/Lk1RA6tL/
cdcvh+fE41aNVHoK+4/oGQ83Y77OozV0DkpN8jsOT8kJamDxIiAjz1xUNBlE6Sk4AoPgZpMScVw4
v1SnK3CGRSjtmh/SjOt9qKxukBrKJiFWzPZxwzIUovRw0DXY2gcZyWIIMjY1dOCVWHIR9JuWBTbI
srAIHLbbb1/w2mJ88wKPy6t6wf1OZ/WBg4kmqfC410i+HtJZIsFj4+7tWUM858YVlz4koGqxWSBx
FucYLNs80BogwbsuIWnTCbK99ve3FvoHNUhMNm7s64XDLmHVYaoUq268AMNTCVM9M/ifwU0Pn45w
044W2nGWs1difov4dGhO5XwIIFc7I3kAgphK6wcVPP4r9yGcC2ON+L44I4sRxi9QnC4rINW4TB4I
xKPFKMgIN9AhT0zrWUwyUyYrnZM4yjC8FqACvrvz2PUIRe+u6sieQrma6uaB79s2DzMTSW6FIui3
hjrGQEA2VQXYunPS8bdvMF3EayaylVpuM0f9Qx2vp67LbdXNB5Pnon9x/ksZCjYJJn9olA9CN8Qh
u9qX6PUDmyO8yiU/ynKEigMryUi6Nzc+miCcjD1aGKTSRYlqxx+uUyChlaa10U19s6FmhCJRa0Tg
xFde/IYgMvPVOIwsU6n1gD6rvUEKtLcv/YHm827bnNzY2hirvN6YP/nHnGMILq3lLqwwn9DeloHF
9KUfHhYCp1C0/9NLdqGiP6pzeyrEnB5NyYrGHbPu/x5zRAKtAzvlYOsa71ZgiOQJD1WT2o9ODjjC
LmPzIHfehPzRCa4w9CKtDhZOAxtTIs/02+DbG4kleWZzpgPOcxvOY584aM6Egmu9lGBvs+Lv2gzn
nsYLAgY5nOMtoBr0HDGf3kEMMr5QTEpmKCzQ1uJ3OZP5PG2KZ7HpGeXdo+TWqWgZwwOcHuzdxg25
uG295gPrSca53fvL34XJ/8QyEQHoflub9W64mobilOPyH48Na0xYTXQDshDZ5BzdW69D2PmFRw+f
uWaURb01mV8JrFM62PUnlxvYuyvvwPCG4oEBdQIRI8XrgWZ9xS0N/Jboe6YXiKx7keSQGUl1nSgl
MrG0x1j2h0bWDWzusyg0s2lgaqe5Gbia0NQHeGKNv9WVXDunvm0RVcAzScKPubxcM2uq8hlvFxz2
Sg8OCpqTSdIur57yvqg1CdjPF/QRnMJYV0vO/ybdAxBiBQvgQhn/8wpQKLnLq8g8+Nak3BX3mSYq
cbMTMpBu4HeFN1O935XFuBMTCsTlHol3h2IIXaxvHFAwAmfVssqWeIUaLsA7JUB+7DWPonL8Y/F6
NPHhROA4uhiTUKZkD3flt+K+k/jApJRvjSc65y/KQJVBOjXobRhmZ998T0/vsCKAQssiyf8gQFoZ
T7DK0djr+eM3o6jl5I4hlOx3ZaDgm/IMnxMibpJQ5MaBm+yBh5KomnQQJiF2HoXxDMfuGPbiqVkj
o2xZS9ztmBsstAKycyxhvGE0BfdyUB10VFDW0SfSnG96NzEct6XBUPTJNdeI9+aXzDkZ2TfRBEwi
I3em86seUKjzRmHcWedVP+5eT++9xedqYj3ZqsdlFulgHD/3vYlEWdr/dQ7shIA+pTgz0DVbe20a
3Djp9TK8yeWtRkANsqwuthe3ydv4ftWl/JNEvk/ydd4/99syIevjwEcOpe3AnRf6tXbpASZjvYkW
mST0A83RBSQYev1hbu/hOmc0CPbDEjqsSfXTNljv9v7BMT/XECxt1ka9LjkPN2agaKioWTgNFIjt
leLptzmVnCLEsxU7xMP2eAOl2fVB+y6xdCqtKcaYE4CfSG4X5fjU7YZ0YwpoN88sPC4BPSuQG/O0
zoYy5QYn+AMekOYIC2FPHu3Z87P9r4T4ojYxoWen09XzmkNllBShoNZluyccXETXKjqYfCVjD7Nd
BMTy8A7bBhOACsNiRlQ1OXbexqXBOkG2A8k3gDoTRFOzWBBuYryjffsxai29TzfdB6R8hRU6x8Cl
bitUT8degyRS4/uHGx/YdV537OzgptKCrbjGFg3mIQSfUmSV7Z5KbPX1M9O5choPlm5amFkjTkSk
UU/iHix2eq5xGyeddyx3V4rQDXmNfu+IxMfTqUx/MvB1Fm7oNKFKpbb4qn3NxXSY3iE8CPpI8Gde
yAU60iA1ldLdMdn3ijMLz2p7lC2UY/UQ+DmcAQDhWbxkjIhizrg1WCQoRnQJmM8Ynew33fc5VrWj
xlB8rHhBwewAhs8uQ1JDyp6+fBJTmTpe5lWAaa2anD5x5ojlCYaK+ERvq20AHc4Ir5nXpE5hxjSB
1CPMEaDyaw6gqt4t6pDQOHiferXFGf8E1nfZ47ckg6zMzEzzHEMOBeMjSFKyJqlX5orbxHjZCwyk
9khrXL7fhpJ9wH1rEstAI5IbdJL+hhmauqg1gXRikPb6eH8chBCMELsNEtwCe775AYAbupjxS4Q6
aFLzBpV/c7fCqqrAsxcphrhNYXzuTTFuNnbDoWgjMW3BcnKHEitpk+i4hMMxpXgSEIFFeucO820v
Ww0HX8ttQTBRhxHTLR3hX6r2BhqGLYT7tHkpJrgOanhvqMGUFtLyuetmeXtMgTABj/vm9mjQR21P
BXaZWKRJ46C+H05lD53sin6NT0xshqtKax3+SEc1DLJwAiefDf93b282NseCuwiygoBlxqfAsJSv
zrN8AYWW9hT7XLvAQWXEMFMU3Q6Dinyz5Q2EGaqyYz1nhktFL28VT+IOCp2nYnAe93m2+PZ/3p5C
S4UlGJBHi0s2J6ImUz7ljy+F+WUEmBovMhz98a6D+FLrnObX7JIRhv/m+mxnWDHk2SpzsiXFrMZu
MG7aOHIkltH3zJoRSXB8/ag0AV4oyn3DJDxcatGrMGRi5NxBq6A9eIa6UpRbEeS/dQ2WAco/oXGn
oMfQYZ1crJ3jA6Sy7YuWJvnvsdUUt1aeJXvgpUPI7GOVWK8RRShFRFiLEqXVKfq1tHdY5lNqq2LP
tGvJtEzj97uwHTRaIswgqVRB1ZF0ZCPCvIFMASWJK87MgIPrdZF3dcab3VmNVMk6dCce/ao0mPcR
p6sYivMfOp17qchT3ZgOYbTVac9qmwkugkujcfEKjSchuPv21DEC4PKuI7NgyH3XkMbG7W5Sl/hO
z2cS9no/rWcOxHnsZUZs1KuKphTTxsgj+4siMD2mcoYJt4NYzL7s3QpsYGC7fJacSY3Vsols13Fg
N6SGRYvCivqdLUl0lQLYxmvcg5xkNzgCEj70XM+b90ZMN9JJxLtBQ50TQSn9CaMo9CgMseS+7sp5
+u9lmBZk2cJJxRaL5vVaK7LgxIQW6eDBHcM2IFPsTZ7Ka+MnjYweuILPa3puezHbQCKm145CdxZG
N9003M/4d4iIBI0RtCpvhLbPmoD2o7XCvlYJZQKaRhO4mNwQK1ecbTK1qZg0TXQR1Zr2C7IgGRz4
xhlBX5C/Zh2xTd0EQjQKHl+XhAy/KxxVUBWqL0uPL+kalxnShfuYnrOL5vDRylAqXKSjEJKCBdbm
zoppb3MzKXjhp3M8/TojTkXhrD1M59imnNqNbTjUCandg6xftwjI+AFR6cX7aSKLqvi6Y8G4FDMx
GKSx9lrcrOV6v0ddPA3W5/arNA6apkHmP+cTF2YFBNgXRFSrZ5CfdGQEnAk/T5N91od3jLthxnX1
SRdawLCnBPSMGJCmb5guLJC51cEdTonVrJdMneiXbS8s+21ATsoljyseAMJmvFeSbDFtk6N8ZssY
8WTgzxlbWxVpQDodEJyq+FTDiovUaZoynUk3M6DsjPDwXaiqcF1d2pPBYk+0x34WDm5IiRKZWhVC
HJHr0+H+vfxjxpWglkgkBtUUxDJzCBRzy8tlSgLLYm2QbNevh1tj/zb+510u3pRLeNKCZ7ZW4/jH
QorxV0FLnlmTPNdjWYC6U875oMEqaxy2JDSCMBIKPTGf4U8cy+BCZQ89xYG3yhcRMn9q/NYl0gxB
WdxxTZNONenS+QJKbVxxV6rG+G3mzGKTW46NE4LkEXUym/6DTDhQybTkD+EEpu6oJOeaBiTx4hi+
8C8xIFMIPWEvAM1qw78ym83fSKc5xHfKlfzZDCSpZrNVLvRJNawSqeY/8304zKlDmChGffBDHx7c
riMW0AMJSZseb6/9aC6KZ48cdhWHVMSXYnapS0I0SaSbvzaCO4JhUZT+17wN67BW09VpOHeotid6
20cfWELvJySC6ko+c4Rb/Mx/Sw2xpUGjkncpuEcsJgH1XM247Lq4KGlf8ANXnG/7WxFBHHN8wy+T
nvimPzjuoqCnTEpuGl7QYchElZIAYZ4wmLWp/fx3bkwpMwSyrQOfNUuw7541kPjGsPIWdiQJpALa
KybP0Enll/tkI6kaW9BydZEEYxHlr66J8OEA0BcmBOqiHB5pGNWWaeAbJDCs9ekj15M6biqMk77d
pHrDovHjtmT33fvHN0K4ClMbJ4B3Nc2rXm6OJIL3aBV9ZfFB0lC2FUImykrlN/uY6Iq4xz78Jc4G
SZV9VkRRy8qy0ty7oGlXrDDJxIQ6gc+VtxZrwTfqjM2hqSagQ6a8lDMRYyxP81e2sE6p/tvwzaRD
H2ZWIeihlEt2zidwkJAqXGdQ2t0+s7Hu8U9YN8L8y3DJEbs+FuYjpqgvdD2J7bMGw/JjKDc5e9dY
mzrp3deUP+wCaDmi50HQB82pWCNwV/E0PysALWiJw4hvrjiyNG7RcM7gVflvrQ+QakozCNUPbw1i
xPPghTo/1XZNVfB4QKoQXXHBxx2XQAeFL2qphcL0Vh5yFbvln+Fnuu8gudZPWaE5FCDg8gyP65t2
+J/ZWe65exl5zOHvfJId1LFthjDDWdgpkvgH6uPQt0aOG0k0GQoF1SzKpwcnVNZ7Y0l3UEXJLl/t
AmReUjPbSdVwkWkXMEAO/S9QHje44bbl8/FAtLuLJ53G4Kx8b+5SF3v3N/TwkoMWTZilgxfQlF/h
rItEPyxsZ2E4jPgEVAxY/N/CD3OrZz6YxJswaPEkpk/F68xWz06McWN5p3CfP6J+jxFa2p/JOjjo
0xJYnwRSPMzcAJxjLEyk7Q5yW3h/IkxMLzLSdTJpJEnSc/rdfNJz/fwbElFMpaEsfN/eD0cJmaQq
xc4PMD/+BIqrz8xGXLWVfQbRtTkPTXrfv534rKnq/9FVB2Z47xcFQ/U+z2YNqf2UV0yYrv+2fi9m
Bvf4DoT+zNxFXxGEW9NBM/kMXhhJg8beBCLG0cfW5aP82G5glMx7zlUT6TQvdpLSHimbhocJhyYJ
MdGnCZ2GxwWHxGumTAM8epLiK+rueSfo3lfOTaYgjWafxDfbnn042oBtxoGRRmDwPyxv2WNhmjOR
nFLkLNSL0FH85CvyGI51WMpOr9A1+r572i7gzzm4PblOkKUh4hrHGaTtN53vTLug8E7YFIetLUXr
5RY3e4vveYUFn0LKsT1cqvcVdnsF4MZduYaG4nHuGohs285RGbjfnqmL2daRM7gU1mT01zH85IIG
3Eu57JWxwCs/xrNGycID2NYI6R+1AWjJcnxbdLA/hUIrOiVYUyn/vNdJCiFcMUjhZuGdHeoZc13I
wj2ZjK9taYA3sG6cVwc+ruQGS+gvKKgstT92TMTmRSKwCF+HwIo1yIDKKX1vRjUQvs9NNgLZT+jP
t+MN19wS/qZGqOiQTG5Poxq+b0ipFxcynqf0n8jyY3Op1+b07VN8/XnSjVlbX254XCllU3Yp4bm0
weLwGAqnGyPfFb5WRcYCcJreaIbh2s8Igv0+09P5u1jCxkYKTwZr+XEzTH4YxSXqhrUUyvxx7/fL
vsdZ3Q3C9+2ADMfL+YEg5+0MtBhwovzZwZmqzRiXYy6CvIhoPmIEUTB3ofich3xEFeqw3LVqxkrE
0wUnfww+8t6BCNwk7F852qTVdVGDxs271i3Oy3SSd3SGvbvn5rKxbFQT4DWyk7X4uurxOxF5Jo4C
n4ZPtifzpGrFAiTse1kHdYen5OaMa3hdBzjAVbZouVwdQ5UXbIgSqjdDoWnL1x17N2DsxkyULKcG
ZmF7/wjE8fEcUKaLHj1IEhvL6su+fpq7sc/NKYpiJY20TrHY+IyJPCy18zduZ7vhkAjrPFhl6FD2
zfsoh6MNk9uSIHWnV5z1dns3YCqTLDlThU/j2cvc7l87zXtq/HUBv5RPDApzHhdeJkiETGOXw0c3
aGUqF/985Rd48cQZimSGsTgWzUiTnfqXK7GEX4eW8kSQFgMMQzFTGjGPNeEVMeBxkgDjHTciNBJZ
UNpoNs5HRd1rZ9akfdDLC2WP3aYINAJ90zEd0A5M3EFx3f8MC2FKkwQqDRY1nrVnFRWuT/XUP4kt
cQBQ7AvZrE1o+weiqrHBRG3mik36OtweVYnIbGycFMu4+pMrrwcweexbt5UaIJy1jfBwp/WHwavS
P/Wuy7Uod/wtr3OP0stdgaMT2ITIzlD0n7LleIc7hB5CTsi8r7TO8LXPtZGJraqw6Qp7LF41PNHQ
53ymi61kffaq9ZTzFerlk5cTGWPg2REJvjek702vTI9b0HY6ttvbePGL/eAdoqtbGaKAeelPc9n4
pIvs999IYdhZSyWuBv+hF/9VRi8lvQ4f413/jEdKH2JmbUQFFKqeljnVlLGIUU0xZQf3P84heFCC
yY2UdFUtBafUbr16N7Pi8Nk/PGOTg6WrkxDtE6+xbtgMipPnxPLXtp60vZ9LXcau4rUnKxsaRh90
frpy453FKhOBm+AktgIaSdRX+jl2Oagzua4k++h+YTukq0KNajf5TFjhyjdCqqBEHxX3W/eBAsSG
FyvuJZxTGmBnPWAyeHVH4rA+3jVfJJQ/Kc467pzZs8zeDJzpmeFDkM1z81htgBeA3Khb9PeguBL1
txW3SwrNNIAhn78MTvAGPu0qCG/6Hr4aTDIlQgoYTXJzS5gSbVHMPa0zpKWsjnDYXLsZIgudzUNn
QjvgWa1KiLxb3POJZ4XenX7wkV6mDJ/qhXO3yYKO7SzTODaq4Ill99slTP4R2Gak/bm3eBChJfpN
FZ55q71Ga9kF6RVoCtNLfc25r6l+3lgmqC2v8pssvqzRDZU2e5oMNIoYnqsbVAq2uTixI+q73H/R
XzxjlWHLRKXGpMzDQu1GUugTMJN9IE/C+Wrqb9HzBD3Y2ox4c6vfVhwfcLmJr1giwtVOBWDAblte
99VcMswf0hl57HJ4j4XQUoQSy94NHcqyV3qTSnnneUB2HBuB7ltQfrlThE2QMrHuuA1RvFOtRqRB
fcEGXoE+RYnwQnPegHVoOBjtgs++C4dfkZYCeGJfoLinkDWETA27/CJ8AZpiPgc3N44GxltZ/Lk0
h5LaKGOj85sylZdLUJC9wjXrQAbsCqlJ188NfxiS4Yt/kY03wbNW8ItiW9xGwh0p7oASilen8AwO
DceHJIQtBJCj9VLZMDU/vSpm3dCg7FxLM08hl62a+whoAgXRYZNbGr5OgNl8TPwEdoFLTzwDT8bu
n+6i1354Cv1ur4aDR37wAxKL1o7LYAIsWqiF1xAni8d0ygDDrowrB85Uqqwnk4dp8IFqSXOq/AIe
YQJF/DMnpcxkEf9j3l4cNVVJ3sgN94SJ5pGrLp6WRgL+E+QDDWVdfLa8U+34njbA7BeRZ4aIur83
rg2PMa1LXthQYB/ZBL60C7Ko17xXelvsk0Im337E9TnIs8Odq40f7nBNuvnTfSA829ELRCuwggQ4
HzTiDvUVQNRAk4751X91p8DjZPOrIi+JHYsyeEW8AIemkKCwvBZCHlvCpTAFrPp3HvUv1Oo9LySy
xPAw0oMXVzMV0gJM1+WbV+qcuibHfBQfl73ZicDpMZ87RcIBpdG0i6eB2ObMRYt5cW+bfzKfYJJO
PVOFWzYhHFNpJ1zgETpIRU7YKS6FxsckQMhGKv/YzT1Ix87KH4onplBsvLW3mWwpFy7t+jDyecXF
hd2ebSmQnfpoGzmKIcFDdTiWOZ+9GqGJwLqJjUAtAJCUNiT8WpO1uhNlx1PTJhHNhSHyZdrPBWjk
i5lRKEn5JitPPmMyH3Cv0sJ2J+knZbTMMZjrXyLLYJCWiC1dIZNDxBQHKwGsjSoKuGT/pXDSoDxd
3AE3uTxIFHHPluH22OrzlharP9Ke/fnVJkMmyLNtu0WbVNYWb8HxSHGogAAB2650qL7ZLtl4BRAv
ACvyPfO36FGTvcjycxWGoaFvMdRf2aiapO1Pq6lt2zWcxn3bmgfftmwrBLRbxbj1BGYltguk6cX0
zCMNpPJRiGb9up/0dzORjjetlYCoehxzQQ9q36arLFdfs1qfHIL2IuireaKxIMs4x2XNu/Gjv438
VZr0qdbRw30Hz2zhBOtjbbf5qRsHZRDH8jTTez1ReS0OEJKiFz32F8huApRMSN937ETcWqEvfVkG
6+2pn96olTib+7CGaUFtmSWUhcr7KQXI83FFddx6RiQXNW4q8mgH9NUD9ctqEnR3eBMFhwvR44lQ
d+Zo7m2LLPFroGOMIdhn3l6wXfL7emShiz3/fNcCqhBZA4xBMQOmIXxMM2dUzdFsSRpn8pbzjmrq
WaUNlidmCyNrYke/FlAGAY/BaIHpo6UoxGPygfXQ4AXoGG8HuSolkzlHo7iHphC1t6CsQbab5zkf
7LHSzE2DrwV7fT9mWmjb2M8BRfHpeBmRyFQHQaJDNFyoqgNxyFg56qW2552V34qcYCvNPtgnDFmL
JlyIVV/bq02h/QXHzYvF8CCy1tyDKQpV8VZaSWLp+cK8C46w7aKCNMG26epWBOp4/c+i/EmX+Huv
OlLE22iAXmi2vuSNAUTDUeOshGo4JgkjwjVhj/9KVz+zvKD7Gvxs6fbfRuMRiMJbjGfMVFI9Slil
/jF5VZo0Z8etzY1E3faai8R5oNhJ1qgOrErWLNnyav5GFUapgBO8BOgLbRQuVlTj8dRRvV+bh/pt
juDeCZM8EhCAtbR3B2mZ8SBDRK5TT3pPVgAlk/e7/Hjj7cpFlY9eFdczIo+yDRCfwl1XzjRRrD5/
1F4jcM10jK+iteLs3BlcxNxpeO+gkupenAEbtd54VKSG+rBncGCL08vo7tn0HOX3AzqSbJvH5bw9
3tauiq8h/weNXUBM5MEqRGydLBA3EQ9CD+8cRK7/7F7NW/du2qBeogHt6uCrXCqSUaagxmHu2Zr8
t5RqWywgYMZSTeX37FFBy2B5oISIT9cs3WApBiVrQTNFlpNQid2ZOqsLUsJIF5d8SWFCZmDcE9CB
0rOfEBY4LOv3FwVnlkx9ymuv0CzzG33p5CJDlsNrWDVvOoh47c6T+MbCV/c4NeAeazwoNoJsV/tS
+UtJZ7JFhQ2TDFjQEGVnQe6kFvOqUHUvOT9rPZyUxF4G1nvQoTFGmfbbU/Zo8atIuE8DC+yHgquI
5APEo1of8+C4xcXBJwujRk9PhadV9NU7yVvcLlUb0DaxCA/Q++OPgbb7nU0FBWlAcXKoUcZlGWqN
OOzd0VM1oPWGPyLE34EfPej3n2sCc8ZDc/Htzwz1kou3aSvXmEXnMFB9dScMl9pLDNrfx6yc6+OL
NFbzIwZJNe/efEDrFSwQn7YTzq3Orx+jRlf/3GL2BLM2Fyij02NfbAKw3jys5aATvSB8Vbd8R+Do
x0ep5/rCRXvfvQqq3cNpEVebJ13VGkokkcyv7MR4uTmgeMVT/w9YKMMb1QAyWMdvU6gTj+gYrXr2
/aCLI2HQrty7t2wEKqWpgyUqhEkf1ZammCU+699gWoEC7+rLAoolKEFda1FwC+hiU0e8d/nvyax7
AfB94sHEq3iAV8dHiurAJFDVzh9y55LzuPzugsKvogp9uv4V6Fe10vLecDWM/uS5ZT8vWKTp16jW
uAyPaMSS1oGPmZ0FVq/Royt5B1FkVn3qFtabAAFjnjk95mwF3cbQNd6R3tmzrMlDR9eAAjxm3br3
GFyeE5aUHuLV0SZFyvqHW4jB0XHZWq0yxOPW9I3EOdVcG/N106+LNVQYZIzU+5t/YTEUfPGM/k0x
HHvNIMcnRIBqTpkrXh/MGe054GqjXx69HJSmIVAo+b7Y4Ohx8n09FRjJJHUfb/G2ipihlDcvVVXm
JzTzNlcqNGInzHLuHEDl+DAG8kQPjQ5scJYNc3meTG0eGlPR6NR3wsTwLbChoL5KnGgvkCgQsn1J
qNDfFsvW9eV4wmM+U7BiQ3e+rWzvgzcx+3viWvpCixvCXdayPBYe0OnGTDrTot5BY3vuD1p1fhzB
/Oa2j/nnBMB2kHjaWQkB67IHaD73Frj7kPcG6WVqLEU01VWiej/VXKOr5yI9n3TIbuweoNvlEiQj
I62XZorvQCCgnXFtv2ciCB2cGBSR7HyJm9vAYSGBP1ZvUkJgvT6pTwxaclPIMr9UYGO/mEag1Y2i
br/X8hZ0ksNmSgwih1B+rqKGUeqpK1f7TqAoijURhFvYgtyIhJsWGV8FjH5tj4Q7W3mdJFmXc55O
kjGdj31UXPfMwZDRMGmA645+9cBDnge+qzP41mk8XxdN7fkeTECXMgCv/iqPzZ2bOVDTOWesrqhN
UN61INLIU2x/GS3cWe3NzJZBk7IL9ZG3OZX+pBrDVFj1oe35bF2smURo/kkfhzCStozOT4rKlTB5
1E9tRHRk68fCAbPzuOXpzhJ8JEgcQVmuDJBOvz6+QicDVnQYg7NOJZrfd1WWNW3yDjU+y3s7nN5I
2mVYgE/X5/dvzyWfOmXN0AfGTOCtU50MuuqEiEghKGExNVnl6vW9fDqN6rmbru5Ah/1XaxIl8VOr
b4cjr4Zg4Qu3lMxSQgjhbXJVMkxwWI4l8BprfOiBHZ431qLAy7W+a0O+0UJqBr3WBfj6yK8SCZsS
/jg0ohbY2Jxh6ESA/OtV1vTkoQNrHH+IHvzPAFAqDgJgbzerAzFE7yfhpiBzMNG3fFIzinFvYUKX
UlaQ8qkIwrf2pcc/TmQTa7IecscftQk5nagP2VIZ+TQRK2MtfATPW0OGE2VfCmkdabsSWKtkUuIm
Muof7846Msj2bAToedAb0xRk8HN6wkE+llMrF/qrotJ8fWwcT/GjufuJpQaoEZfKtttF2z+8kHb0
aacmonT4SdXf1KNrtUow5BlB+sbMRkC+JN73A1FRMk/ERM+URvdRFf1J+YWDf0eonc0YORquNIpf
/p6UobcT7eea6g412eOPs/46Ooq9iwI9Tf4EdDtXtkD9ilmUMdmzJuTA7tEQEUahQz5bypHRvEfD
e/8WBenuikCaUP290roEo6kvArsB5coFWCkXXB3ivZn5mwzIPIRPpkpJOM40WuWwt/2sCNSeWaa1
MXqd8xKkjOjqp7zpOw2wDbvAwZrit6vs7143T/IfA2rDTjAnF+ynh0JqWucCpVAdgwL6mSJF3EYi
RmOX6dsQQ0NvnAZ8IRNTU3w2AAv3iVjenRbnBZwobnULKEpGUIBXm7bYlavILZJGeY+KfirJYq/6
yPyCbJm7vD3Ekk17/BP/dcYWNZEJrNDvgdLcSGYmtR6b6UiPsHKYDvVxFxh4kQy7eAVxvWFumTEL
h6yla6wVlSk7HWwg8Dn6k5M7QD/+I6Pvpjc/0HABP4bHf9Bx5VttiyU1gS6Bugfjg+3L5GMbImBP
AXavEyITPl9dgzlq26F/VBy5TOuH0KgKqOyFMjCCY8ZeB8DZsUPZubDO57OvWnetUYgGqAHM0GyN
Ajl255dImGllK3MxoZivy/YbDrptkcNBksQWUxQOj4v9ac7iw0FMqgCsFcV7eSG3sd3qE+vRJVyo
wwU8L+8wUhR8l+m7Y4f8adLjXDGmsM49zwqCLDWBBlXYcdpYZAmx0qiFo7OFlZkn2El20mABFM5V
Jg5P3w0/eHjv8bgzcATl6sosotE/+lrP1FfgExJwZ9RWvgjRoa659oSf8jnsnQAIGjyNjRRjQV8F
PHjIQwvc2tW+buorlq2+IqLhBhnRKC+M/J9/mAnh3JhtAfFBjrDYdjYvDYgnpo1T061LWJkWIbqW
yyp9xb3B4fqxTFPptOdd0BTTxd/HHSzfsbQBkrBUD3evNTsWsXjewfwwyX0BNVFSgDL+FwwWu4rM
/dvsjWWslR2S82SOCYnbQCIe8tSS5NZoJ/xo5vpZGHeVezb5VfYfh/MoHhsVdEnxCbbXIWcR3FGT
SXdV05SXCvPSpou6ACTMzuVkk89pReT8BnxNkTQ1dSICHVg48UxgcQ/TXYlm3uVxk3bimEgVqaMu
cVDWDUwUkI23eCmBqwey2g7G4aJZeIcvkjD336C0LpnYucZjS3Jq67eBd4tKv2KY3k3Md5Z4MgTh
gRI1VzfW1hyK7JQksZRI0r5KCMz5CGRyvvCgmTmMjsOWqkd/BUNeaZAv3XOG/v+ioCgo6soDP9BK
SKhFmihwDzx0BHEvNv6y1ulhVGb6Tr4pLighn7+WGxxdgp3ucByUdAGNYvqdFwgoNTqEnkZ39UmL
P9nGkTFwfxnOUUA3Wg3CU1x8HCrz8MraZy7tstiM/RPHPgSK1SqzvTIIeu1oFgGwBTFk2SPggm7j
qAgtpJ/j1q3MT5H/D3RykLu6xOVjLU1r3pviDRaYqooqMI6uVIHPm+K8/Dqgx2gUZumAueHlwEdP
NpAVkz8fLxFAaY21h0cjrIs0aqEvi/Yupe/gdgmcJLcBLzI/29rWJjgEJZpibUivNbswLsFXNJo1
zfAH4gKjP46WXXXUsNCfl6zMZj7K4BaDlHsRJzGGj52aRv2LDECBl1VdPlZyYbH+ub23IY/l2j3o
EMkb5FCFkEUXkYD/OKD8uGKDROjR+w16PmOBqvatactsFUlJ4BG5GXbXzYaFv67/GBi4am6JU2DU
qng0XF2BEmBG7Idt2gzNs6mJzBy+4QcsCkBru13uIlO4jOjwUhNWCHpZePRTszt1RwdQIAu1M2gD
U6HBGO6x9Pcvw7be4/bRjyVG/uiDrMdkfJ8Z9fGYPMgpQFKwV2uleuybsTY7VMsUZWkiZV84vl4G
1bH+/GBbgwo+WuJ6Pou9eDEzIBZy+X52vKbUFm9BalvtFOfTGWoyL7ACXqunEYfps2PbHvRuCxFV
5jAE1sQ4OoQUxlGbfdKuS/4uGljVwWPAEBR/+JQlx176dxGyVrBlJSXbPmK22CxKaWvUXBZGM5dh
Qv8ISq1XyRvgQ6Jly6wPxKd3nRo53UfG3fB3avEipfzaA7xQMfDlFl1j/LMRKQNlWwaipVBaw+WJ
vjwRwm6VIGz2Ix0W96HA255/grdNr+BzXHkhXD/UoWALxzW/4bN5djQDIW+dfWNbVQ9PrKJ1x0WM
LYaMB1Zju/zSx5sUmgUqDHGVa8ZS43WbCvcuiX6tpDWJ9m7dgxF0VBp4vtK3OwO7F+s6MLKz3AVA
r6qoIZX7En1w/YTsgFJZyQYK6X2QjdDm6fbSe6edk/EiwkkUC3Ewrc6IAu7C6Jh5eNxbG7VVwO5R
SQheNwHP6fd9bGejL/Av+bsc+xPUxewGLTknnpQ0bQpQ+A5O+6PLAD1EV3Q7MoiJHeiM9y6WsxAm
ubOtHAxEcs3DODfc9Brwfn69cxPBC0H8H2yl3MYViXDDikKpLbN/DRAKUGr+Bh7HzHQ66VoBs1Uu
cY1z6Rvi+F4sJTrcFljfx33zm5KSw/M+Kyl16lcaHaxy2PeESIoz6QG83wj3/++70g3j+0lXuHIr
1S6N8VK4sC1IZ8RSqwLOCBK767ktEZn3Gt8Dzt0JJ28EGpc+yshq0ykybQ3cpMSJINO7eMWKwqvf
DF2AAPiD3hxOvzcaeThxOuDsul88O0YFA0GVvAWb66XpFj5iR/z2C3codmp8ChYlasnG6A8YEq84
HfmD6obi3BbI+M7vlBcl8fj9cn0Y2+EmwPWA0TfaTLkSAmAZd9fkvyMUgSHHoq5+OTIOSfrrFkV2
xFbDUQf3uf1fz1db67TTCV1ZxVjjK8q6PcAM187Gv2uDx0zFK7HiQBJqq3gLhYaNs3vtMRG16vao
fvnS8sEc47yJHi2jg4jaJLwHmq4Y72mlgfFHLBX+gBsrhpR4GLK/Vle5uwlV2GIUZKACTlsQ8HKx
UlXX7PDiF1Qkj3F5bk5lCscSR6ffvRCnmXZFGLxSISbgaD2WxLoRZliyoyKuv/VLHJaQbQd9gu47
TpbgsmF0GDKwhtSuNQHnD8l8GGvD4L45e2hZiJIBIy6bWn0S9yEIiBsrXKosJXGzteBu1/PpvTN3
7id4RxgkPYNNLfLnr18fVrT/sUqGWWLJWgJ016aG4UHrZPJjMAW9IUXZ3pZnZ66CRRrs4mj0ylKT
7tZVwInrHnnMksokbV5a83QkoWLZe3a8Hvt+BWge8Sl278/mkbv4sq8aer917xLXjmtql6Nt2NF1
PDTuJaLXCni4kkJE4otjEzvQVMo26+2ibbYssthlaJpAh6qYA9CaR1icFV2rupCw+wPEaDl6r/Pc
/F6SDO1TU+GChdx+aG5EdMiG2Xp/wMlCJn2zBev49iuwBPyn2T/sQwP/9X9u2+jhROcALLEOjx8w
ObYRPo0CJ6iy57drN9twu5Tj9DUUfpLdkkYcNVmPuPpy+NhnSvLqnpW+Es/tvwheXQQbo9nQn+26
cm1G5P1sERLU4pAB82QYVPMXdp3SBAeWQO4odCgg3YQf7L6Iwp6khnc71P+fJnQD5mwqqrqy32n5
9pe09z0k9SE9X8/+e+m0d4/88n9j4BroagzriS0KA+QrPAZQrI1N1OU9Tk+L8nxFKmTyFE1cSf3h
9hEuXCACF6lYmrMdmUawocWQz4GlT5y1Kmoq+ESO8+Ao++eL08Fs4kuqQAy+tgzC+Al+1v2y3v2Q
PfGiU2UBOzJNmgwGvx21qaARnNyTLcZHFDIaB2wjJy2EuybU5wRyAVO9zHdx3v/tN7vf6dkMpmz1
8kfrnWl3BNtb9UBLWGXNfU3zOO6OYs+fbYfk6psJfzev5PG5qpaFIkHFfyvdALPKvYuKET16vNlI
Md8qA6M50oiSiCWfpd9q96nOgLk49/U1iOjGQi6H8fjFRpzd4+iRfub7/593sePfe4v1+PvgqKag
QYKHl+oW6JJq0KgDFzI5m7zsxwlW5zemNgREESaBK670Qc0nrDIC7OrEzx/xq1nPNHG9tXymrTAp
RwwdOKiL16rQQJ09pnJoHzSWIL7x9eo8FsSPBEG0I8PjUKb6Z7uzVgba7JAbDOaiHlHbLHM+T8vC
LlFU+8m70aM5EV0F+e0o05XrMrIE7gdcfuxeeeHpbww3MXE7u5N9nIACQP/964Uf8oce4+uBCGK0
a3spnVrOIjUcgYFOPTiBb7ruyeonYI2NT9eINohIhiPSv+6WyQP53kgy/MTS8Y1MP3UsM+1t0ytk
GcD84wHOI9BmA6wJ48en/tbcYqxQfEApEH/LznzzvEZK0gZE0Qfaks1fOvQkTkeRAoNykBXs8a3n
tmiDgZYENQCRzQ8/deqcTx0WD00sxrxlMwhN09Bm4nk1mF2ybFkSHnxncUuiw+EWn9nH6pkGBg2k
E/vX+3cUZlmb+BPFoz6PEPoWtcQ17bxgJs9MNdUdOUqL7DPdISVOlR8RQiS0QWAQZ4dPElbNOzOb
7edyQfRzeus8g4Mhy3JwmOZsEae8GT4n4zCFehZgTu84HPjq02NViFF2AcjRluDHGuBaMjc/AEfu
NzwSrU6qohoK3n4kEIEBahKt13BLzc16yzdPopHrr5X71BXSNtm29/k3vFFkiTHYQnQsHOVQENjY
46Wn7XnR+tc+8UKxH3TnMWVUxt5/sa/oD6RugSERK/elmHZrg3zc04o2O1Mc1EkXByDoFCU3cvCV
KUHu/BNjFPR2xFOr1s2QgvS0xbEW8lKvzoxH1jvCtSWguqksyh9EAk8PuVfjUmUeRRebB0w/gZYx
njJK0SaXlppNFcpZigrPlzumUnKdfdzkoXkd/7TQv1lzgnRHUmmDxTMqWOSRZ0V3gUujP5k73SCs
iQWQ9ZeCdNgb17Ut2TTWSL9+Cwm3lJpZQNwMhgf8NuDER04ixU9qiibjyItbkakRLAvSN//D91nm
PsbPTkj9BKQkyB4nfntP8Iy2MEwUwSDCJGiYWtf4gqB2Px4KoAfaCIetIqQfz/bKPv/KaybJzraK
yS2rBcJ4VYIceoecTaCaph4c6cZoOKstLgN0Nj36XLc6rP/iasp6f7mB9shRUVvOQRdkMDos+iRs
Lx2es4TateOScOgtDW7pKGigysGTuEqwSBXLSAiHoA7DHJZ330EA0RFpVOGuWdPXaN5VDrWD37i9
2RS9tfrLsbFEyVwmCdC5TRMDn6piZQAFS0B0L4qrzDFsOIpaXcYe399XEKDjyHn7RuvbkwlcL8/g
Dz4JVkI6GJqrX42pdSfBi0PcvP/UImr45KOxuXt4s5MPAu+pLAse3UrRwWLENyheBEiP8rFQVBa6
WN2kNiLEEyZYpCFDCq2qCYkR0faXTNYyo3feXXQ9mqTnRPYdPij9e/Rf6N3E2t2Iy6ky1ZpOzuFk
ViiN9MltZ1SNFOPpjNeoWHKAOKoDpRND4wWRLmXFdRTgjtAR0AdvRoV3okF2IQNC8D9ehJAUS88o
0mUgeCXHSSVXG7ZlF7K/Ktg+0Jh8kSaJ86Mu58k2NKdPViHvwWHt+imwrBNPnYsC1In/lukyfw2W
Hf8iexxFa+E4FU9zVU4YyMw1FO1aPXA/JpJcqopypOtcqM2Ttoz6ZhsbwW+alUP/lxNsgKxN4k7F
swtDhn8RU9Pt1tMD6JGdTvyqD5Ik/s3zUGVt0xah6npDXQsU3ziZyiGpWR7fnAh17LwEFfyCKfdA
EgUBi+HcaBhTaMAlWlDsC1+riVtpw/VVD2arYNhAV19WSkdXutBIGkjAAFWKcvrAnq6rIonLWcuV
AINTXmDqn9KdjFPeYo6+vDGylr/TLCK0omQ+4DrCmjQBfcRGDbYwgGYc54147xYBJtTadQql/P2P
0tORsygLfUJSuVivC7lvpaQIySNEZ1pyHzf/Y2cbH53kYiqRNeAqH9h9+SOHbIbe7WFZ2WH7r/hP
37RhpSD/5l0TlXS3tZCNMyBsXeTI7YVgT3Zyj2/9rI3OoyFBn5+vaZ32OXIjBFMs1zg9IS+R6DS+
L88CNZKd8oV7wLrUE2a3SqcjvnZbSnx5vJKBh5TuJLwWev51sP3F/DNij/Q/KOzorHPmJ//M8QGo
EOztE/HkNFFxL5Y4JpOgrRGkZ5T5s2hyV60yjbGNCfWtO1782qa6iSEfNdvR2oryKOuvQ0EBJLb2
9B0u9dthiJXWWenxDecWsBTe1ex23UPQ8CteTmcHpJBrJAyO3WPE10zsK1Fkn0sGT/yXMkgIZu5H
03WOnuR6POzUyjYFg5NuMX57hSdx4hrDfHJugqUnBeyiTPpwi/dRiumTtCZiryq0/9it1xFkNXxl
/4iL3D43qwsmRzGcApR5XkbCpUUzBamRfUmu7uXq4vEGdrrCR8x4x5fNkOQ+UWWTAmEcYapjN+u3
A5xaKFsgDb60qUdwj04KCAEGjvuPs+66xIQ2AknmmSx5p3tHgGgunLFU2Mnzk2TlfS0YKa89NcwO
cg8l+rqXwMY3dx3w1xTDUtZHqkcpgOmZaU8D3+GI0K0sps3CUZh9Bzz6kWDrGlRfD7J2pX0Ct7YR
VVAilnkDchFCzT0wiJqzaxdPQSxiwnUJX82v7UJJsObtKM8Gt9TMXooKPv6GDB/wYcEGyNRzN++B
G4zvHz/Nvscuy9oPPqOouiuSqrVP/p8uFftOiYZcZyjz6StycRsoMTX32creWyW7h5OD+PLPxM1C
9lstHWHvANA4uKIZD5LtfrTmDIw99ets0DCPZX3ISs30r87gJe8Pg5jrxccjhyWzw6s9B5hLh/eg
GEytejshOsmpkfd3kwWY9BWtfqUdy7A9z8egpYdoNGwTIpyZ1TjEi+bALwWcKYogz28V4+ZEy+fA
gU8fm4m0yOWF3R1WzhyiQcriXByx714l7Nj5hUPgEA13TSRcOrkLqqgbWDvoYI4v/lvqx3U1y6LN
Zq4sYA9jtBoC3oaS0PYaU2N+4lgmT4Xxw9sHJ+i9qWILM5RbhDX1kWADPrVRhXYSFP4RQFhviUCa
z/jrW62gWXIOjjrOFUh4KOvcGCE1P2s51dWa2vL2Bnx7Ekwz3Nj78i6WX1l6nXhVdIpGfmYbN/PZ
k3OkhhNQu5Lf0KnIHXAIn1FG9HzRNYeYlcsx3EMpwbCNwGHoJxUvEhvxaul723VMDwu23kEShIVq
rwOsD+p+nZI81fspr/apeOOwzza+BOlqQHX1tkaXaA8xFUplviCy0IDxqSxGKn8fQCpoZ3BmGE7z
JpKBPWXzUweMzyxI9Sv+rWpF+nnCOTvJIti1nLXkDNYPtI7zm7znRqiMeuUwG97unvBBbAS/6uy6
zlK84XcxYNPNOL0MjPYWi8rj85sP+Lq44tkvsUf5a798BWP3CTzV/L1fThqEtvZ4Q+RI7t/mosJD
PAFmVGolWq1C4mTnKosKKqUxOOx/iQiOJ70Qdc4/NluhosMz9iS6kyMOw2g1B5YNjoBW5ReFKjAm
SZ7qZ9afAyxF62DrVzA4KUEUct1KaFaFUNdJO7splwHnpnTVohE/Ln9AGhrbSVWZokF5wvZ6q9di
dpLBSTK81wS4oEa/ypiB/xZf3F6zHIZBkv48UmQBTpobZvAKUy3I6X2SX/jV+PX8Myilz3tSfoA6
jRtYbQxTmZpTS5AGgR74u4T1k/b1F/sPCH7WaoUyO22TMNJeQ8hOnR68xhuhCc/MhEmFPJLv0Mii
Xa2fKzENzO+EeH1+qu+r/S5okoRO9qkps/euw8d6ZNL9mMuxis2ey9AvHiJyVcr+cjKExwOB5NXb
+Azwwvn7Vu9muicIgw9H/QucSyNXG4MBiPi9dieAvInJRhdlMSUeEh9hH3cKVR+www14bgupNe5I
KwovAvFVaK5kgFb5rNL3jga0Q7b8Uck6f/khypae6/Y/5vHiBg22xRA4TrY0D7shq+5NObIjmULS
8fbHmDeFNxdbnYf7TPTwmvjuope/R96aR0E4GbDwBxAsU4kUQRTjzsQ8z0mEmptlziCRAF7fQQFy
D9ZlKBop8y/RQHX00leXArrezbOJXbvAfsV6ceXGKo5Znj902KgnlD9EOoDDKPgKKOtNegyPsL34
0Rs8t9MQJtJRnEMI8nvF9ciBIt61S3lUXMIGdYYUznNSC/kkHTijrWypp2uVm07G/eRRIHjxlGr4
Ktzqp5DEQJVpTvJ3bLqpin1QKd8h+TqXKfb2fI8uV2tBWZ7QWAOgyU1uOJ+0ZyU1LpjowqKJ0btV
Fp/9BMEiPU9nNC/cRN0NNU9HbiTMa1QigXNxgaQwCeOnr8bPWp+ZhZmszS4Z1ydGzf8un4aj/+fD
5br2fAIj7VbnQrUY+a1cn+pcQLYhXTVsSmi23BpzKPDvJ28zLQV7AnR+ocb+edMJW/+G27cbiSF4
GFPLCTQlv5w7vEP0FrcmEoosB1Jcmen7I+HuTwXe5fH/DbRMG3MdcZSABCkY2Ve3bflUfESkYvko
50h/iEOAzu5KWuVl35z3mYJWb2bYc0Cpv9dmjzSFcbzVrmWHzguVo8oEEaER2/FnNMiHyfxl7CWn
XzwIZt81eRrHJ4UeSVYnmkWhhP/6LCsGfKLzFn7rlmE11qEc2W1o2J8ufR098A8hf6rAOsqyb6aO
SmB5Aq5HAM/8Lq83F4fpmofjmeYuxlCwjRfyJdGpwpKOovdvF419KDRgjh/TqzljRdgQZCjJwPc9
iZqnvxZpKViPZ3OsMtdzd3/awHDhEv2WA8rjg9Pme8k/mffQCIfW6V4fPmwAaay6YRRCs98pDlhf
6Q7YjfdVcE9svVr0Mo1YIuMiJyz3Hr0TT7DDNMnHJtKP1je94T4rUrnAim5GVT2Ug6HteQsG8V/g
eZ1GNVrnZP6gz7c9ZktjUIseum7Bi6OE385zhCjsLrWRyzSkdX0GG2952/Tuw/WUGGYYBuu1fwI+
lp3C43btwSOl6Tmpu7FRNgVDoMJYhigv7p4BHM4a69GUwIt422treU+VB3/ILEPdFA8FANjpLT0e
tzH19mI4F0J8jKojr+mdvQf/hlBBjP1pgQPcGg0CxxFUdioOoEGBhWAxBHrtkl/dZITDZ4s7dJzQ
cxzb7yRrQN1M8Pn7kGnSFX28MisROyOGfFU10KdCpJh5Qq4xYcPLI6eXBNvnwsdD8XNt/67L9X8U
OVkQvlpS2KcLRqyPjPWrd9AxI2uXHE/xaogT1X8t+mqCjM8WqH6HvLOHuxzjXTIC8f83HLp/JT7J
oq/sNW7qzjO36kidpc593oQT2xPZhu8zKy5iLMNl0WsGDPV83E8teFBM+S6u3NsT7ZpGzR1gMpgn
HVXANJwREOKYeP/oD9JqhrBz2lNOTSQzaBznySiRmtb1fv4f/gYCk1Y1dRUc0ciWILZ7G/7AB1Vf
LZRHNR6Dh6DoK+AErPMV3L2sGjTHAkAqRjufrG0bBwCQoF1uFMo5sj8fGqXshQ4vCB4rpHLC8k4I
c1aLUxzujY47cLMFgEWILSjyeVlcPXvhWSSYJaFwUlECHjaSqMH6LwJReQKqWJ2abXb+r9D0OakX
JB5DV36x/ot1ZihvoF7vt/sCfqKvDrxV0V4PRteDjTHFYaJzVsbCXnU1HbWgx1vq14+kSsxQfWlJ
+o1Rt62kwWFSdl+uDVBRimTneOg6fAhalu9E2K1/sRTZu/cyZmSiFzWAB9USAqyB3josLxkcwA3b
HteUxfjGeLhB5mhMpUmMQSj06GZ3OGy4fqLasnRgcnZpe+lkNKUGKhUo6uw+6PEOoysnDDfPg5py
ue3pKbnOF+BplYxas//bMG8PIwBXSbERSCCXwHxZXBMmFBIrnxofk5TSq45/Hq8lK1w9Gxw/+Pzk
AJ5KVa4H3+PId/drTm+odF2tnzhoYK6p/bnBWF0nGRrs+ylxeQtQny2zh2p2mZzy8+1AMtWsKCTU
j0MxsuKHzMvhs5nYwHvCc6C3LcKoRLll71uuTZHlZVHlddE8X4abTd/kYgwWxANhC0u0Cmt5aOxO
5ZBMefO/PQUqAAVOX5vmWN1nP5BM+C9wUSeJk0kXOTFHyvfC7n6g5z6s5H3tMKD9PaABKgVGPo3t
Ib5Xfo1l7+6zd+r/hw0hZ5drnml7ZFOiIy0l3X0fu6itCjm0HUwu9HEwsVtx1xkyGeA53NycZAoU
QhAjQS5awWBpjdOo+up4m3a/fi0KGmD7E/156C0tJPkMUAP8tneeoBDffXA+b6ngT5E0qYt0mQvl
qPVZlVL9mk2pZI1IS16jXm6tA6RixpwiLu1ERN4nuocKmFBsQ/SsB4b7EfFXwUP9ni8mdyoWgcrG
pkQwP5CbVbsYqTklFX6I+kiWapD7R9vdqtzERBOapdkoClRKw9OvBtapmXiy3SR+GnQF2TOeyhPd
kMcRQ6KgqRaOJFyj21fzsRpY23OZAfvdgr49qj5Le/GZGv4eqML2gnVwCkFruCR0z8spLGYosXl1
NNl78rWWLE3l4XidsOg1CbQLDsk/dpzgQRNdj4yhhKL0orqP24OO5AbRbF8iOHSmKfMbQbfo1srD
dw8PyZe7RByBnkR2KOYvISDpXGvkRns0jkxOq+gJyHaByL72Y++R+FB4U1lNF+t3Ycv6Pv5xpiT2
ZwNKBmb5gcJlVeP/dodZYGwbALP6rrzifjC1wxl098VyL399gRn6tCX7Bz9e776Gnq3LTRnnXKJS
V3gK30ROeZC/rI4Yf9Kz0PBeIt5Xw+Dg5wE9f78Gn8usm+RbhCQIHf2rUBViOLpZGWSQqE/BptRp
s5ePvdY63llmqD7kJ5uMGz5E2IJNXXb+QgaJuyRImG9YDu1fQaqDjE7m0osXFVrG49hMi8fP28q/
j7/LhhpgXuoIxZrc2Tnzgxjd5Ux3JlXPURlizAH9VsSrH5uWb7dcztWQMyleIxxVfX3HXyH+A7Oz
4UBssyZTpJlBOa45sjzyKp1dHskNKZ9YTJWa+YgU0zR/Krll6r8pb0sG0f0s3sOXyH1z0A//PaAI
Iy1QZLbglQdCTMBZi+IMowFiPeH4IXexDYw0qcXAUXZRkblOPc8uW18sfS4AyaX9J372ngt/GGBO
/efuDqEOmSHvpwpK4sjENkPr7V9HLINmMcAvLX7dHAMqyiwM/1cu3xX+SzJGGk1GFhv8mTZroXZW
vQ4g6ykBTvJV4rdfZ8X+zF8abJWqgrv+WOHr31eZWD8Hj9xyCXT+BnIyL39REiIyHR5gzbZyzGJA
FE6tjwrDhgkOnYZO0yh8V6NzqFWMA5UZk5k96eAR76l3CrYOZfEdpfTVdDw4Gq7HEvgvx9F+D8P2
vWtXz+Lge+v0kX0pRhd16ETo3y0VdwSL7tJUNmSSISF6OyqCgqvX51xPA/6nOxoeTYsSPsoWlk7p
/Kf+VrnMbnbipOfMWqpMqxLjOyLWGDRlQJfIqYfhBEgkQhNaqrNhbUDL038Fvdr7ssDIK95E7Gr1
dEAd/2O9bCKePqz7NlAqPlOjJw//CI/yIrBxq1YhTqq3zf1+wbcVhjV//GPZb9JTFneUb/9Md3BQ
ggAWY0BbhZQo86+7UjUhephe7gAn02jnZ56/3Q/lI2R4mF3C+Z0SP20SCguVUN4hhfXydZkLDdGc
OwTC0mXt26cnLS9e4JM6OU09tpQXwS+DNdHRoFQjUo4w2j+jeIa46moZhYQPx3WN7eamxzIim6mu
l4V7IPZt3d+bR+lOv5goT3d5Q4yvcyosCSyA5cOrjQ8Ooaudut9MW1SrsoxJhyO1HqwA7Y01+dvH
iEypmaduTX4HAqd+uynC2AUhXUZfrGpwNc0MBm2Df2Hx7dmk7FJXMhoQF79QYd+W/c3Q/42iuoqP
CVyQn2HVpJXVQawU169JPyRlxIvy8epY0PrQzvuyg6I5wETpUQvGbbY5eWSsmCgWJdQRwPBhJGu9
d8enI1HlmBY6CtTqgapVcHQ7Gm+6cq5dBDQPhSBBUx+ZrECC0BOen1TgvlUMjNlACopDk9qbuo+2
2YN2Zwehu0A6LmdY6w1UJylm2RczHztuxBgSpJeiULSoFwvGiaGFTPrv6trxCHEA2D2Nu+V/2EHT
9lCYqUaTonnj2+m/VPer8rkp2YaAwRkPtihJwxlw75WoU4AEAjiUsEma1Nun9r278c6lN3We0Feo
ihRPvYKMwmqD9PdOdwmswpzd7GhqHjcVTmHD4cWbp5ea8tSYJiJUeLKmdeOHjnUylleMzVaRw0+a
aWn5nxOCBtIA9VfxwCQx3dH6dXmA/sUq9jdAiT9GR3GZhMUlnswkFycKPkCLDXMAkQcj2NwKillx
gIdsSF7/y1C10oomAQ2JkwsgFXedqwnPpERxuNEh0WLnmztdz2uW4+Osa4KUyBNDhqeypuSwULn0
tsQ/BCkyhK4x5/Ea+hBmdvYdQ4nQmgTJ17b6kX7ebWbIzpiC3HWW/5XhWKes3ZM26U/VMwk712CT
jCQwHyRtOBeK/WuluBB2hc2dJGJ9GucwfICWsRVS9+H1USoRe1+/IqrDIiI0rwDmwNtuW7nuYE/4
qlCLegiH45GUcchRcYM7eXhaIG0izAmwX/tUuPpT+N2VxH1cqGtgyyzuaCDosQLEBohhzpoxULCg
3ClTj8AkBuglJx0wHjw4udGpuF13TYixmB2zYBGCEF/sYyIONr3w3VcU/3BcpL3MKNuZCT/bL0F4
JBteOmE2Yb3hf8RW7UgI6ViadYGH8LytIBnfujPLsAik+nnd2WpTcqyK5pTAgR+NbkC4IPL3/CYB
BkEq8Oi8ZB3jrg4O4W4bm+COYfLN3ygqj1/0iwDVyixME2clbU9Ec1YKGz/2ZjTfW3eZxIHCE476
Oy1F6pQ/0onm5BLDX0vMJEMlAG1CJzheKQrOvBD+BupzJPBzxYW5wcdIx8kE3IajBGyjtiX4wQD6
e9RukRsUcV3kkuVakGpftkQ/nE/XJZsY8zFhth7nlTj65XPoQFq+vk4Pfg6MnPyEaS2oY2i0Ck9z
cUJor0krkJhZqBh5rUEC8T3kLsPRoNijVXbk3ZwA6/Jc2VRjIk7CwpDAgVVxHF03pYs0OQXUq9Fx
GLxl/4b8sAUoSiDrw9BvPSVwWK9H+j8w1oAIrVbwyZUKA4NyQLdYVArckhNvPSLHeIOEgMT/EX71
Ak4gJRGBsoiqrlXOVbyx3TZt2iYdEAxjoEw7UglB09/oKbqnjY9EqhRpjcWZH0VTipr26oIKy7Tk
eRlMfyJ+EhNgIHbZkTn2EIO4hORsA9xSaw6+ZP4qgr2YQe1K1Ec88K0g5PHtfM4cPuXYa6u5ZDY+
ZjZecWMrW+wnGchb/blzYQ6eBK1nk80xDGJ5fDWEU8MDCWcuQv8ngsYJMkemx1D3lEl7c6GIiv+X
T1gCy2EDdAzDF+sIwLYjWtkFrPfN2ah6YluY0HZEhDCVuUBFOER4Wh+5G8vdUhhdBa+7sa4/Y2k7
ff2eCKn+EjYpsj7WFmY39xt43Cc0X6JxJJLO/pTfDh4G9AXurBf39Qh2lEhROVgB71ePSRSozcIv
cBkxDrdbEqoEult5KH+BRmPkQpawYNO+FjRrYj10isOOVJrFWjuKx/2/DbGf/mVvQH5dtv6QZmSi
iv73awEm6kLom1SUpJHuvZFaaZyiwfP9tElnJyrlSrHg+Yvf1eZxzH8DBMR2/U19L90BDrLyA0ri
qJ9C53o57Qhac1+L9OdQNdNhKnMnk+6cvYM6IFEv3oleC9qdcB3NPaNZJTJFqYGNbzZsHOq0bvLh
X5+JScmnVguYOCgLaICLzEYkPgTAUDRy8Z6NeIyXp9gC0dM2A87WTVtkmc6JzKI83LiAO3NGPDy6
/1GHp/lAZJ+8Su73Qsx7XimiXxcct96VevbFgxaaPDCXafVvLOTREzC+L5dQwguAo3VT0FUs5Ter
Vkvd3ZTX9t2GhJpdJD6JYlLaS44KdPbspNKWXcm3OGNtxTk9N8r4mpM6A5vxAOTNkCfJ/h/QADJl
HBl+LR6FhQPoKIaoM7rU1Z3dEQ6tXE43D1qecQObsfbKTj8G5nNLMqAFrdiouOqQtql0fFl5CCCx
gvTx9t6bNgIAjz2yOiFRhhXR4NcIdmcy15oSAVwB0Rj9O41a1Pp6OqjjLtA7lQzhmkLzp0gj60Nv
h2wvYYxMaRDfgB2cIFC0PEQTimubNOEynb67selLFH+EBSmH/EuRoHzLyniMwD749hoYpzjwS9+Q
z0Zmwfa30qvMG+W5lGoz1uoBOlZsuopGSF4/zFjbnaCHTOkeIWP3Ra3jRyiwu/3k2KSkeInrNqCD
ZEqzlPS8agZr0ew+ERO6Tgfg3oBn4mENMGqCRCKGd2TGa+n2NRun7EZfGRPqSDnfV561+3McSd4g
AsbowvaA0xYUpDrbXaUMyd5ni32j4bvgcb56QWEVKeB/rITSqA6bnzXhimgEyFPq58Ntc3vBkXNh
YxETu+5zWR+Pf1biIvZEW8dkHHkgslmqujalCbGEaZYeZLd9nXDH69tyRWTuCIc8avUCbGE2ZOcU
nU+ZpT0qPDDAmHeu1E6ktQCKESbmczpGwuC+LNRLazTwhvPg9lzHRtlupLLHhi0+hlGY9rk3XJgI
7Go1stPHXJlvdJtCGQAHR8/sQtA2G4+9zS/m/AWKyS9cZuusJzjgg/SMbWbWOENOih4fetKDMhSR
ffLkiHwsxAipnfb4qtGhn63Mf8XhQFvd70NpnB9DIm6B1a3wFvje8usRkADZNE9xXD/ksGihs0Lq
voWdoH8VAuFfkCccazoBY+aiWMHUWdx9rSN4GtM7nWHVG/SznR85azi1S2Vb20USPrTDdwBuy2Xy
5Puj/xuOZ+0SMiHN+6WSADUayNTLOaKgXAPkj0aOkim4Nhj4SK7+QGe4i9sF0ltLwbueBMQ3oSSd
JzjRgSFhHQmFHDW97t+BBAa9AGwrrH3h5sinwKQAmKD1eEbuZFTBjLxmetM/qw5S0bN3nAMhI5UE
ypSjhmLYrKBPPrZwKWuSIYIuZNzfHtOM2nMX7b7sNTClabZZAQfmPjWtcIdydEtctz75RIQi6Q9L
qROdx7/7D5CL5fCUQpxPJoDDfZHuujY9LvJ/PZPAjT+Lxnoe24cumK+9jd7LdS+gcssisUYCS8te
8gLGrN24QDXVRulPuTwYfC+dXRU703J/8v4RlsBoS6M1S0Vg3mdLAUuI5QQAu7C7HKAgcSHx+Jl4
NtUC7HQWcmLM8YaW/gmOfoK2CMeUlB8Mgqov1fR3z8UZiJdeRcDsqNZUqwQ6/qllhVgFUaITIsJb
SGPgLTkfoz3vsXEw6MuM9lZxOn0he7BwOdA/SCzVE8EfFbOrvd6u1hE4lj9KbelmY0cXSkLRCTjG
X/6lpEx54ZCccSVvPUnGObJB0Nn/ZS7L0bFwePX8bUZNgg+gTVQ+daB39hFKJ2cQZDsMNWFk4CFy
fMuIfobTjEmKnevDbFfjDEwRI6Ng81I1I9F+htnyNp8FL1bgfCMAwsj5qm8cm2E5gJ7GoTn2sZlY
HzI0RSYM/6ZpdWZnWqhXIiw7VUSfGrp6AP3DmuM3YJIin8aFd3rW+X3pwG1Uo6y11/ctOt5h7GC8
UD3Lzrx0Q7VHPx1YChQ0Zg5KwvQiYWNcFUHA7babSdeGAt2vTTE91GgyBb2SJGa++FgWedFPmyXV
T4L0ekhcu0bO5V7a9CWZiBpw2x8T7w5aLQfECavWt6FCuG9sjQfpbBvdWlvofBOHd3aqol/zKJLC
TJPoRqBguN/ungrntaKbht+x83MddTTI2YiGR9OGWIM8QpjNQl2ZYutGzk4NOFDHK0ozaitACsHV
TQsKbzBVECWx2P5AErgM2iW2ywYFmFG/1hpecL8AJjqSDyc+nGKCq1r60PezsckfdHBWhfY1S4eN
+SBd76b06jFmKZ8Rwx8OE/lY858ydJ+ZfCYG5CSq2YiNrbeH5ecdu6NCvDjnWiGgLgqsyhTYgwrQ
VroSEcmWAch3bv40fTKmuB74Ep4Isnk2Q+ZJp045tvgbvwoOrKMhp8ZiTdqipoopAKJDC13geak4
vJJIaIGhcjpFWJPv6+lKjGyxtlVCShggn/ODZNZOaUTYz0mLTdp2+uHkc82JR0rfcKKTXM9FvGm7
Z/vq9g12/PL2QLDE2DIZxRUt9AqDFt6T7oxtMA6WVpLU7Jrl3WgaaC90uTBOOWDBF3qcIdlUZqTE
s7y3t94/RNB0EpRHm1lKodgTP2WgN88ra0AcA4iV8iuDDFW1co3YNCs32XMldtyQFkylCPmSvaBM
LhX3vUsoIBtsKZIKq4ccf6+UiC/IAsBQpcGcE2Mdmkf/0g9zFhfvT48AjxndpPtEKsmLCbJFe5Mm
P4eksEpvZdHNyvS5P4tynxzDODlRYqs2n3sDttkVMHbAFtnbP+KhujYLZCJuY8jJIQ1z01WZ8q/A
soEoTW7MINnu1PBT200Nm2X9JH1raMVCXn6QQEvibqv39fpx4Z27Mk9aC+aTluRUXagBJRRAp0QY
1nG0JYWRefg9nUXJNfSstrruOn9+EkOJtWoEtvXWldkTGZoDBu1koAKmYDvL5pb2Pt3sNt/dZQCO
zvBjyGw2SzepmvGYctnv37QxTIFv2VYYKA02U9qb/D0I8ZrU2L3PFm+lAFWep39pqv1e5uqcmsEf
5P6bC2QSJVmWFGLcZ+DWxLJi6HJELlgcswYf0MK1yg3YqwbWVV0ZYpZUHExh3krJ5GaWxgJlcLej
LaNH3JlQyIx8tIFAQq77MvNcBvrUp+A6OH6Z3tJEGtV/5eCj7Br6YUwPW4wzQ0mDhsiSWH36VP/x
g1/xLNOgb3W/eB5gW78Lp+qLODD62IcYo5Bgdya6RErZE4aEoHpcN20qtqK6ICTANsjDxecaHnCK
94kwKcp9mECb/74e+hgfomvVNNeup1BcBt9AyvXuWz3wA/kmvjSlfT5Gkll7WYMlmOjO6T/VJTvg
w20F3mBdlBRBb5tXj/w5hOgk9/QaHvBNpXd7HH8Cr1AM4GLsydPXkyxAHG+AoPAa2mur1yzfla8x
V6l9wBz5alUn0kllKyBnKWV8KCEOA0QUXM8SYnh2WwVaUGbBfeCkCOEBAFmLYw9R+YnUwX4dpw/4
o7081PMFKlyB3bUEvfzmHKiDR9zTz9incBDGeOfaQWPdIELUSYygccwcYtUGkDxnXNj3MJ2pDKfs
+H3PEqjGgg1qvWFv7gCcOnIScvnXBC8E6TzO+/MDyXo2BzCScJfGrg8IXUGTJUktxho5sg2Q7r/+
9uQ6y4RuwSnunRNY580dlQ+tqT7dYpCvCykYitTEQm7+zfX9taPx2P7tFezC7NlOiI/AqrqZZzkY
ekv3c1aONn1t910ndz4yoIlzEsTkWoCcQWdcj4LL9P5Q5ad/TRJ/IvqPzAb9Ext3t3OLDb5mbFbO
ej9Wz579zS4JIJfWqyItxZwFh1rmxn3FZlCbUo5IMHpz978Z/KN48jvvakkkKSuAiVXuSY4IgO2A
tISNn87gwgm8cRPdOzLp6aDVVwRi9MTC5ND7OUgxI/dxbo10RUrMq+penM+RqSt5CCEPlq1tYeMs
LBiVp1d+IEGlDfpe3kJhtudC1FnnIq64T/5ud3PkNbVaEi7mgS1In3e9QliKw3K1/p/18QvIXMgP
hSND5rJDE5NzMA0drxR7AJOXU3rTLnsiO6iT8l7lm+ur+bIj9dKeYPdhOjKC6MWM7tz6TwQ/tr+W
Vi8DHYOHAHkffeCGezsYQfbpohpnkOvGKo9Yq61ksEuDMMS49U/3ARP2iKNlkj4U7kkhHZ+rJKSM
gzKsf+Lfae2KDpHXcJ2Z0GRywfoTklowBDjFJ6nKD88bhNFfdcB1PDsX+ymE3La4tI6O9748CClN
7OYmkEn2Yb++0gfDdZX6shZvhKxd26LZq/u+Dw6CiOdvz48NnarfB3CCLuiWGVtZxesHLCJZ2/5t
QNr+rXT5GF6tXkU38s/Cq/VKUmEHsvteMwbM0qar2iRtr2a+RhWtjzU9GRvOTL7BhKLL7h217iO3
DAnAeR3XYSB9sqC1feeolV2eILZvBQ5OKZtqKmq1JMeO6lLkDlgh2DlvIhV0zt7fpJX1iZO4/Hvk
MPqerVEShEWm40D2v3k8J3eA2HpuHZti/OS3y4zKtoSsnh6RkRXWPdd6YG3bUuRXXliC3gNRevaC
R1JS2Oqr4OTxqo0cwiJBFnSQ3AGAuC41OoL3PynD8t4SFCmjgBkiq2WT990wLc7ioh7qjz6PRgsF
E3x4KpSgpGmklAkzxoQuUTCpfo+ZNV7ql8pu+0u3oj+FouYGq++D4/5ROR8mS2rW95Lv4UmikzLq
OfPxx/HL3JiIkCXiVujv7nNJyuZ3lDa7E50J8UYF7YDo4gWuBsr2YJzZeT7+rM52gOzJf6eqA6Rc
u7h2KtAHk1RgJhYHk0bpmHU2uQwt6c+EDnQKrJYRdTVa7ACsnRw1BnpbT6wcT9XdSxl/PGZez4Lp
KR25GEV8qHHuRfhEzZY5fX/yAFP5LyVs0ZUN0D8iO3U29c/l9IxVdc6vd6uVVRPIbcg9gCkdZYHQ
MZL2HYhVhpaL8ss3gbODK24mIre00r++LooRt3hCzJjKl4k1sogyn2jI3kciiSmSRdD1WPNqDN9z
anB5yn+Ft6MACeEP/Xt5Tvn9HdvpzC1XTQ+08mOgQPObSCoLRBhQ8KipMJCwtJzE4AYwRA5HXfWz
/jYj1R64x4SaXEhpYiulmxMDIwexfL9ZnLQrTO8TEao6jmux+2i7D2jevE9yRiTZ9dv+6/YKZDX/
bbjvpI5aYtnNUz5yRbR/mXubE8ebhYWDmf4nyw1LemTZBSylyc4VBKzNErlKgVQiFSiN42Zj1N4Q
8X3Ig+ffpXVA5HYm8brPO4RQG8Yj/hoI1dwEZ09lrsN/s/IwNIpl8EoKKEh2Avq65c4JrfwAgGef
3of1Rh+hUa86vD+mZ4ovjy8/Fuf5nMJ5EHPVCn01Ejy4N75WdD0aYl7nyhl/dqpBLt08uDN1NCNd
vaJTn9dh8JrtdfgMmsU0fbJ8SKDv27WzNC/Z1AiFquBKomK9o8H5cgEzQ75dTPs9aR7ISt+Tk5Kk
xRGd/b4Edp26x0ygbvjKvupB+SQLn71s8O7nQfzxo41IyAKGqKuFCSNi6LUTPNFjoU5XHqsadDG9
gBIzIKjDk4u8lsib82pj7OjpkqpFyiNwZsdXSc/ScWq3bXOgmbmNVfCdxIPtq1TR1Jyu3tnGI/EK
lN46/NhOirK73T6j0ijqPdiN7EBCwKuA7Xi2zUV4J2kCWoGDtjib8rWgyZmBVOSSkCslWeEkkbD5
5Y5hBwABwkT4vIwYvElF+caPmMJWQkHobVNVK/O9Y4OIYLbh1RyusW0vH2ISYvOpHhvYRBCqT1jU
+JiQdtPTYegxOo3Gmq2QF07KgcJ3oaysCftU+8ZFujbo+OqOI2nTj/JiAXjppMsvWCRp1w/ZJLVf
DVZ9qlCrN6k3itavyQybtASX2qUiTa9zhhUu8rP7yvC9FI1xWXgeZG7mO4ZOJa6VpCDX6Dn4mXjA
V6L8qbv2prtkjEYh5OUHwwE2fOeuL+40juGg+0TzRqp37V2Rcf+ouHBWhZMREj2OpaTiZ12Lre6p
5xnOlU0ewAkzYgiyzECO6dtEnFt0KNzcAf0SgIGOU3VSkLlO6+3o83uy87L7viaeOiEYfOxu+SRw
YZXSFPOSFKwAOpi9uDXnflZPzZzY4VkIU0Oi5V0qQyOntSJ2BkEM8xO8M1NhIuRaOG2CXTE//83/
CN9C7P9zcsNdA9Ay/LZ7mWUTMw/2pecKr8OfX+b62d1he/0781hItZgJ2FBUJ04HhwwjcbtzEIsL
Srl7grONtVhnEjWUYFE06qqNWBSyA1TICsSP3VYtnFrYsdhGnIHuom6UaDKa/wpeFdmxFNsK5NKn
MusLrqkM8XHf5/xVKHLZioZcwniK7Fa6WdphmCA3jhUdbdNJR/7Wlq5/+vaZk+xBd5IBaxaBT3DU
c6HdhSUR+SFysFKJZMVTDnvgID6QGctZfcsw0FTHWrNngIdzGIqR05F0e6Tq6NW7df6sVU5yq4EP
A2kGwvqq9T00FKolKS1lgHZMHXlYW1H/AMRM6IRBik1mdzkIo6CTOeifnfjhJUDmGd7F3Xk2tWeE
+btn9GFhw5hOoQAresxBBPD7QEy5F1j0FLUsdfBqg0kCwFLE7BA9L5lvVOiAdFOhps8xhQJ9LmSM
xvvnmSZiv9R9M0Z0eMgoZpESIC+tIIxMrz/uutW+3xLA8dSbNqV+uq6Q5WxekmNP4qhhog8aLZ+6
yBM27OZX5/WABFTLX9PSW7CY4s9+NH5A8oZ8Gj+WWfq5+RE9KskUFfUSw01qsD3tbNOKIeEuOwVH
A8dQzHhhiG/fZqSXKPO3DTQYzV2hfW1FabUNP7ynV0iClpEHjdLJm5E8Hhh2oW63qQZ8jemuDQV6
nRs/t3dM1iZkhjO1/oAkGcoYVtKDFHGe8t0WsQM1vU4QL9N+3o77RRTfiKMGNlF7Efp2YmJTR1Xv
0dAaHB98F8nO5i0VG4+UEXH5zNa6MdNCWfDhWtSEh5VI4kWNYU8uSlEHyYRj6RWzfux/fvCGa7X+
YgydXYuM5ylU/wODrGaPssL0dxXbmKXR20I7NZeqDABRaAM86UZ3xiRla6MtVXrrZk98tP5iEeiP
mxnx25r+fdAs5AgQ20aH65ajEmzoBge4XM9+hkTXCN+iBTLR3Q0uVZ9c8z6QDaCjOESN/+xQ2xzk
ajhzxG9xcAmZylCCqSY1nYYzC8SgXD811HYvpxkSfXdEB0eHnqfMWkQzizI0thaHrBHXWliFY4zY
kAs1ykKFLetYySsrRSrTr94wns//LT+3SEJwlS3QJDjks/+vSTgDjXBgaWZvE5M4lwpCGTRj0DbK
lfDp3J/rcYbYe67yxxif0y5zmP0GHa4LOJscEMP6HeTAUbvwCgU50kSmlextiZ3UwSrZYECBqN6B
A034yX6ivavM/eaY5bJZYBiHkK3cZSxmYHbPUjpynD47WqtwgcO38KCQv0s1XOWWpq3mvuSmaCXR
+KwHXQMKct2YMeYnvaPmY1OMM6p8y+zPaeI6Pm3DRWI40vJtaQEwO1fHnRdM+s5F5MAnrcKReFey
wWtJz+4K545K28AwduypkYPKwqY0nNds+Pdt+HwjR/e7G7jgZRCU74RONmtvKB/kuyREQHPaqz6A
pzQU1conUYsVSeapOtQ38yypGzRUAgNsdtQ6TBT/G7dzTK83spjI9HV/Gv2zAn5phnlRxpxb4vr+
0IU37+CPxB1oCtEjOb2kg4uJcjBZSiaLv/wWU8cM3mUaF4fsQIsqyK0zxLw3WnH+R5fbLXLXHn+P
Rssjd3ZgRsOcCera5e5Y+zX25MY5ofk5Rg4yXPurdebqA3srEwAf7xtpGwPd6/PS5qV1c86WHJM+
kY/ePfGRc056BtybrcEyW4tsFI31ckbDjZUG5I4E/JDipV3GLmElD7nzraea/uAZl5pGpBLc0dA7
mdIo4ms7suPf/QZ7RwGGI++lFb3/+1uwxDQMlgBfo6JL6C8KnjjPL6O/hBZdOBvpEFnRL+9zxZck
dr+wKP6DBL9/cFEuNZIOR5E898e0a1dqgC67ANZrN97cLLzPriUW4Dwaa3Gu0nNkcs15eMPb+LZr
fzDeIcr/WweCpl5WzQ6eiyTHEDabsrXVBY/AYywBbG8RamRbEz9y3YbK3sqHzHh8JWdDNeoE3rjz
NpRV4Hzs6YddyaXMxUFPlofGUF0OpqKKZ1lAoaWPDxybr1jTriLPdGEy4PZgDGlHVw5pDV+ZWw2p
Q2VtqxxeIN5PSr2crX39x4zK+TPJRXeJFYdgpHP4Pa5zoqAGOtrln4x6/jhAgHJ7E6anIlQu1Fkk
x9heaX6UnZqLwIZ8LTj/So5acYTBFApUnthZdQJNIY4DTqpAQH9FuSbxFxxIN+fa7G6kkZq9axtM
TfQJjJPZCgzahy6jDMn3VlyzJeVuefFBpgOoUPBiAmgUb+PTqtKDPEnkSC+P7T83EygGPFUIkGP1
zsEfXlu07eXXeozoCjumNl6pMcS20N6oJYKYsQbnT4Q0XJcl11jjafCH6v98fyUesL8JE+UcxaZ7
NNFiVZFcqIbdQG7GbxUe9y5dc55A93lISk5vct2groVlVFS7Q0TtM2ThqVV9C+C3Gb59aJ91P2bm
z62lmLFC2Dn/B7DGyFOP2/d7A2I2Tr2g3x4F8ktpwBfxStrfDdnkNAIPhg4pQKQKrP9+nfCO5Yn5
FPTQyzbhKOTsrk96O/F9vMETNZKelGrGI/6G1GaIL6jre9GhhhaMnBJpACU2KUq1VxuVUsAxL7Qu
89jlJ2pMBvUeEgIn7FTcj4zPEe5yfcCmx+NARwtK5yn73ouyKl6xkG1QPrgQ2geBhw7vx4sAfj1l
KvdvluNcqiNc3XKT7e6Eu+hC0tBpFbD7X0r+imS6tfMzI8nJxofpaBC7E19qR9c/HzbYIAMK9R1n
gSf8QFB61X/KriIS1RPpxnG45ZDYj41JizC7ueHvNwIbU+Kz5QmAiK2mvfPDpkA88VmAiw4eHd7x
AU9KZYYnnxZQSXd9rc8Tbv0TSX1Lc3Okd1odXst274bEz9I4j/I0lAJZbDjDSjo9Rxj5b4ZQ95SU
SFnPec1xpVXd//SPVuMi3ORjJqGjEl20mk5ZVlp9wXgFLLo13BcccBoKOngM6KIvPAn5A3BbYJ9T
Shfk+rfGiEvwHk8kDAaFxw6akrV4CIlny7gRRFvoVDPftpiz7mKnVZaKFzLaLxB7gpASONaQuvAH
sHQHqnwckmSzCaCNOztVqjpVQLRvOuk7BXKrqsvmizfKSF8Cfopn6DaJltxxr4VuY3TnVNNWtME0
woAcSOODBHTaPLb+qgDl/1IhhR1pYTh4QOYA1G/cIRdU3Xzq/j0UGkMU3yvEljciUONup/U6sOVI
XiYHuapLz/4YC5MoNvMPPm+sCCEKsXM9P5pQZPVNOleSuUeauKAkztWcpZ7px7+gX1tPItibA53N
UwaWJWvo9xp7HxQR2qnWQXOK7hCEEREHbjSafl4FfsiUB+MjwomCrGRnNp3QDylNADZxfg0clgCf
MZfRJKbXoZNPxsoEAKfJjDTtB5pkuAEHUdVSSxs8eYA9aps8MsagS7PrLvhFf8tP/yI0ySeHUMwf
bRPIUCIhkIQX7mt/UFyifUjHmZW4q5k9g4rXLi93XlCNl2TlVY3Fl7LimEoPa+jYFDZLUAjf9FXr
PVfdD/qUkXITiqEJ0mzPSIPeIHmDPgzuayHxYQFgS/n6rF8SKrb9U2ykY1bRjB6m+bF4J6spj6mt
oUW/RKiUaPgGSJ9VlyQhLYnwrkVnfFGg73AJ8/93UsnXYkKCkEr9+092GXTAmjVMls6Pse557ePU
VK3Ft2dqZdkVYRRwzCsn+CYzpqN/8p4Rlw5CU+KqkfYT2Smdo1aK3taGcuzflAi0nvs4uKy+K3Ho
sfkvz7OENNCOqN0VnmviGjK3tjT7jcgVBRMOtoihJ8AELt5TJUj/oP01BVxDwZAe/3CPYkG2to2i
Na8SKn65RtdR/bCAyw4ef+HtPrX1TVlLg6f94uaoy3IJ9ES0GGoG5pyqcG+hkKZP+OVqWxQ7MtdP
QNRyYIfcfES6S9j+MeJxNBOpTAvdyBYaeTOxsMiylB3MbQh6q0ozAP1ii42ppfItaSR1KDtN4Ale
wrd4D2hQZY89B3siSkDKELRLbTqqPFqjRpxeFqvpXPZ+Ex0k/PRrBQVopL7uPBuBZJn426d++4nJ
npEYRa5nk5VZ68vYG3D6gLl/Nv0/2ubIYZAVpZ3cJN0BzpRcf7BEfHaj7h9xQyq8an9MNuA9yrx0
/4cU2gxUfs1AY1olusqJ29UIIIsXPFO0AToMN7PwCeGVUQBTid7Vki+roX+aSTypF7nmdvvWy/FT
nGgDZEywcP4f0L7Np2UKEXoeRDgCFt7E79TmJP9RbrWSWscD5z42zApdu3SIBC2qei0wmGB1ptJ8
17PveqDIoee5r1n9nF7IVEN3YSnjDZHTycEQuaaHtrVVkwFLOZCP89GseyWHzdnERIr+oIROqL6+
CP3ZGHlcQLfcqfZkg332sxi/CuqmVgdv9Glxa0vzvppiE7Lp15R9GFFfNtyRPem4TVR/E5dvU6Hc
F1G+5KspCkHTVeYfWiCG3sZ+iyInrnmmnBcLzjHLJ/O8wicWThb3keup/GocPYqJ2bQtN5QR+b0+
p+fnpD+SYo//T2VaKJeM+rD9WMZ1tJDGNfAnHj1uUlsXPirUVZmVrXMPQJmxhwsninsNrbxJAMLD
/uGIGaTSHACc/5eJGrK176nVugUHj9dh8GgTtb/du94DTHOTXxOOryZgdD4hpEqxLm+V1KFRWgLQ
2Zzthp3VuZpN7qaVZzqlim2Gn5X9wetKO1wR+pYjVPqgrPsD6PVrTkfF4/4Hh8z8rA6jb0EIxEjm
znO1EfQ9GRxFoNzs0JM/z9EbVFQUbl3H8cv5BKvKHZ8AsT2cxKHZ5tDeOrNiVWRH/4jnRsS3pLKm
89EnV4dVQX0Vbt+Wz0iYZsjC6UU+NP0lJFk7Y7ZHIBgOl2RPBWjIh5YJDjTfH9p59wSN0imGmT0B
mtrV0bXnHuykoi/LahIf+AiFJWIQUbXgO3802vhgX3pngBvm+ozmXGRP9WahD4sN/rNMbsrtzoG5
m4heZALhHN/AvTsPShf0r+mrbh2J1mERcSP+3oynlwUJkP7G3S3uN09USD+W+IfNtKCVEB8sTV56
TiOfxvwvyMfBFOMYhYwk51tasAI1P4DZl8fT+tKqH25h5/QnEluN4V9nkjNPiaT7YiuQxJ5MqapO
olkG9bvSmOdCIV5zZAbRML8nYb+7SCFO2uxKwOakaVXfBnjIPBGsfQ+Pa7ETFr6vYX75t5Snibti
b3qtt7JLzl5enOWO5C2R6/5CdHDc5Rj9Ot+h2o9l0OGV/FxkKlm7Eno/hRifw82Gljiw2MHwYZZY
5ZtyXAdUrpRaF79+Mg5oNBE9U7iz8ez9b1aVqy4y9XU0526RYcv01GZZAr8SgPQU/eq5v3EJ+1Km
Hij7cSc9EJ7TPahXI5Y6ikWF40DBNKTWGZbxBJdtC2d+T8kIzYOsO3zVN+AjZeI7HQO4omu/GydC
Ssgad41pi7wzn3u2n6XN5nRg6GAgo7bM0AFe+YHSVhC33YWngjXesFrc1essmAg2k0XBdTrcU0la
6wjLn5GQCWVR/mTFpkaclbmoMnVZqGBjIvFQhtcN20qzYC2sqvKYbtEUlGB2Gujc05foz9OZnfat
GV8P/jf9Nk+RCHzX7vBcmkLB6LDxeFmZ+nHnJO0F0EXH1gYzWmw5ygqPqQ64x95Db5VrVUID1LUG
TthGhBaPl70wPI4klZjC81zIJJzHeb7YYOpYu4wXrzsB79Qjt0zeo6jEl5VSlbYio+7AKphF1tQ4
0qRFwGVpkSI8hOn0OOiOVgMPtl4gsX1KldwNcp2OGeV5KVGApS7kyA6QItelpeM72Vb0vMV8IGDN
45WPJov8As3eo92lFU8kWJFcZu1Vn93R0DBziUrn6CCYvWdTRt5F2HBUrMIKIl6kVzmQl29czClF
o35kjrScWBDK5FqDOWhnkmjTzRV1/ZuhZ7kGgmm9FZ7k3B3o+HOuBSiA7F1NskF4xBYGMwedqCHb
24PryXZWPc/eCqgDpwusLzPrNuXBbVK1Yls5x1xxeJ6mh7XmCf/cNQY4Cy3LucARLhXlHFCNrWt/
HOSw5baCpIJgq/elAQD7y0YPW5wMEC7DNK4PbZ/QCyF0hpbUz91p6yjMBOyaZe2hyYf4MVt9QOK1
RItBYV/5teMqmKPFzmppNJFA+RYxGuRAnIejb5SCsUjwj/RIWsNFibO4HHLW+UNMLm08jsa+UzDc
hV95txAWPvXCnIPor+/Xmeny2jND3ckXyA/RK0apRjnOv+RLI6AkTKMbSjSZcJJcZkzVijX9qLxz
ZGgAzHYzGOdjGYBcgT3TkxV1poup0Ux+7JOUgopsFenahLq9oh5tm9E0lBFbwixIBeDIOToJ5a5l
ilNAJdvKUQZ7qpzRvO+Ud3TgD082fAo1QvEqh8L3aVUGX3SaGzO5xlartnmQ1uf6XMeBwRaEJBb6
DBqq/4Fb7R3PI7Cn6tDqSxzbCLhxUmFFjYMlqM5Qtfh/zsHFk0kS6S99GY1PfZuAYTWrjF+GyhK3
YHxwdaewiuDs8Gp5360JRxW/2DpD5wnRZa7oA5zRd1qtISHCgYqOo+Av7nTCaFZY8/AOuGmpsZOh
q+Pq4fyjx31XU4oyQ1hWej50Azp1FnW54nCLeQs273whyMWO8Z5/mnfzjW8jTxQl3oOEN5c9+SmZ
ka20gg/9wYN8tEuti6wndhFV67sl/ByDudD0dmGn3ffcjEOZ1G/ClfOwdTkudH0dYiwLZouJeGbL
3leTvuAahrjPwa0Y6k3NDuTtFeMbo9Gpo0TqGlY5I2LUP+v8EVZ8LmAX/NYrqQXi1Za3gH5SY1JG
8Djyknt7IepaqGNyETVm7IFyNFQwC9G32WAlq7X0JdBi+nuIzrEljBPJEbLIf1CjzO9lfQ8f9QyZ
B8KElTxKvjTFFKW8c8DgWbqeUFHoAw6MHh4Olr7Br3JUwWKrVKdFeXift/wYVzcKcH51Mwtprf91
5H03B6JF7TD7oK74E+P06b2jYXla6kRtR/jTQg0BNs7oq+AY0+MTdmxXiVM0imFOC0Dak5bnJl1k
T8ibuXtFbvHY82J5wgXmEBgcEV31KpqJ6sqFL7uzYra/Ads4gPRKRUUfQjxf8dr+AcMoKnv/bh4I
4uryh8LEF+AlM+2TWzlsPMmlvUsd/0/3A12Jh/aQOdfpdR13eUC23m/Lim2h3DO83Ro09Y2caUBu
3fv/D77/9WsQpslKhZknHhH/Oa1LU0MUIjdOOy07QBGfSLjE0/nbdLBihRzItZjORAnTMTbd4WwZ
stMIRc5ljaigW/Tf8zuzSrZBNnEeFHps4bwYiedyTQezvLgR96nK2NcDD6LK8FTCK+aB7yNpg0xz
5Ad1U8it+cm/MyZ+Kv6HSe+6U8V7LTm95iTq8OR0/F9lgpgcqDpk2+C80PJDgTivPjhNgHkjnsAN
f/8IckVKzLSFYHzNLAURaR/XkB3jR6suSxGtbHNgUwq86/pG9DdENT0XIGcqmRFyBtUMCF8Myefv
UAK421uQMYfxo0y4umuwj8Orm3Jo8WB+Upe0Fxd4Wj2jHQDwJhFnCh2T+OxHDW2ukqMN/inmhq3M
7LsTwc0hB1Flc/Gnd8MZdAFafEXkC9kY3WRPCJR0ErhtuqRDSD0AntqXnmgQ9t4NcqLoOjPpg3F5
DVksoxBy5tQMeBiaSL/h12aT56Ppsuxp67hXh19BprygCfxKTtJlyJ9gRyh+P4ZSmOVQZGajOlmK
KgrP6nnkn0/iTHDnSN1jcUfOyiKESx24opUQRRLZHY6b4sBiBbZOG/wFeRQqB+b9I10D6ERtz4Ms
Qgw9+14Q2eRSdSW72c5NJ9d98ww1EfvCFLVMBCEahBdcNKeogfDRNC+evzieLciRrcSadtnBIl6f
r+t8ZMGEvdemqS2gO1pn8xDq9ThJT8vsJGdHn2LZ8a8JZA9wCvtX2OwQ+BPRQ2SlK02udoBkE/zn
3yuFzR+oTltXdKWxdR6h+sV0B9yCW+HlEEZd607lvrSrNC9+TJ+fqKU+bZpUpsUVCCFRdoxp9bOW
OTcN2AQFjO+vyw2hp9spYGwFHpefZTcOu4gSntnaHt6zS/EvbMZQT7kn+rpRM12RNHyuWENyuxyT
EyFIVWCbisuFyBKr0YhVYKqRHUQSDqaWqlj0ZDPxb6+gJ3U+BwSOANw1sw07rJRvn7zmW0r9feLZ
7t2jzzfJpC21C3Hx/yg7Y2oaqh8+CScuRUvWzkZQ+228fGyhKt9bv9BYJvhPxxIKt5/lPct0WmOa
7AxCxY51G8DRD2Rucm2I0Xk/1rj/c6eQ8OkDbjXGC8+w5Mf/oQ4wS/TQjB+ATggdirFHALweQgI/
Xas1XNyf1eVd9ukLpA119J6jscDCTvCesnWiFXPWIYqc0hgR0TWPEcACUXy7jw2hfs3K/FJgPY/a
FsyiAjTcJHZvzdCtg5Dp/XAYxOI3AuDDDyhFNqPJPborBgAr4CeBIL1WJAfzTvk4bSGhoC4DlgSk
4L5SutauTH83dzBl7ZCfcGqWD6UsxAWu3xhggcOBtGhd6NtRKs3rHycunP0IXNLpiPzr+XldZ4gZ
IWpwLvbL28G0XOPa2hVMKGc9hgUMQD1wQGOYEbkctbSAmtBq2oMB0Q4RQ8qS7UN0SvbjTqcv65fg
CdQx27fTb4X+So/sOrn8q5VcDt9JoTrNJo9j/aw3DEHTB92XH/ZbUnfiSqwjHhgG9tHI5Vv93cw1
8b7V38bokTSXcIH44TniUyXsHQgnVruYlZrmrkGGs6/oCPq6irg9OW3+magg00XMALx9KJdQNxow
A5iQp0Rk3YQHnLvCvQJO1yEvK8gM25Q/tHCndQeaZ1I16moaAXNDL7VhzN9aWiRdPWEHC5ic2/aL
Pe5u5TTRtvNoWlYIpz8kkB078JVCIcWBlXKRjCBYv3pBBuwUfRJ1cbhZ5QdImzut5357Cv+kKaeE
g7WYuU1P2iR+5Iek+o/Bjh8Q/UVdIHJEJr3/+BWh6wk2fwFqMO4jg1OrkJgfIRnfcFs/U8phKOPN
wkBNsu0JKpBrDBFQPq8N5QJvcWSsQcqgkodq5fCt50qE/pkIhOvuwoSsQKct7TEkGQA8P6Ii/IS2
NlbNEKHKt0SFZmreWlN8Izj4RJZihezKjM6MfIhQVRkhWP+SUrCzR5cdbza2YTypXymh6MNoydUw
OPVvC8ausxWK5C+bDjgFX5ED3sp11M3CvOZhYpm1APTJuxeUJqU6zMxOojXokPvsszA8o4Z7zGMo
qxgehxkRB3ekjJC/q3MclJEg01UzTUU1ad2V5rc6opxc5jKigodVHNZuvUwhbogVPeQ3e89zh/6p
r3CqYFzUwqvHy3b290FCnEtr1YRIQjB080dYUis+DwNwpPBVevAu14FxbRwQVYHZGyxM5wxZ6ldV
IdgqsiamtYhq7WwlY9ptMM2rQA1f/Cx4RWTxBCd7dNuysGP0+DCelnGbQPwxKse3fUEUrxM1wHED
R68v8iKMAqVSUTAsVKY3/TpNSQ3tz2SHh+JETOj2b+iuCmKHI4d56Bm57Gz6XgrDcGr3Ymdpqui+
baOZkJMRYCiR3uVNheUlUnokNRZhRiDzTE9nxfSrxcpDy5tg/kOW5GeCCAu3/vaNik0RWPtwC2P4
qQ8wQlyU/LlymCfbQ0Dw9osdFuoNRaCylhWBcBoADyuKPOcwTWLB7ZEGjtzNIAjJhC77qGrcrLMZ
6N8EwvmSymiv32TBTKKAPKwudFXz9SB45wcQkpMqXnKCp39b2k7yo+ksbT158Yidns8GWxvzsMR/
RE60N0h1lz4eUeQVa5EfGPD7FLU81Z1GyLFmwdKGyfKS9ap0U3pZ0eMt6sAuSVVR5Udd3lryAw57
GbUyqoJHwTwMzyblAiuMNy52KMAeHnKBOUQoGipYNU/wZcYD07YVSoX4dRINAyoAvJwjqK29tZVx
8prZlv2c+goDlPT+Nsay0l2YnXsjSiQytgRXsNUeJn5W/WkdBFtIThhBqCHzEJCOMUFp09T39BqX
4MkW08AUi7evL+4uIxsplEZ4yGeyGVUT9GX+uK8QbTeuHk7Ul/rql2R6txKOoztpBR6e3r/UJlFQ
AcLuEuzZUJQ6RpzSs5Bx1h2PAKfCrKJaQxvSypt306JS0Xx1dpNnnDl6jIIgIW68TAFX3U/v3D9d
zBqT8liHnb5Z2dOzOqS2+PBte3cWfk44Lp9dnN6sbo1Acodl8uFJphHzH3VCObpO8CvpMVekxr5J
gNbZlP6Ih6qFpkQu0OunriJdU15nVXmW86slSmroRtvlgKqFyw1M72zTb3e5sMSJc0QJUXZm8A1C
F6wY5lEb1B996DGJdYCJjjUpizkVRbgoncnkZFxjr49RCy0diCvowgTeRGsqu5j1kI8nSRpSu/4L
wdNceIoMlLtbb7bF4ZoC1YpmjkPHj7GqkPK9yW6Un6Q0KVz8aMluqVFpwhxFAuRidRkuy4KQRqVa
QjmlVD1SjcXA4rSRWXnHJUAWUcRVQ+WTiUgbaQ/NsyYr4oXKQ+CxT4F2vdW7QOkRuaKvG4pbl+x/
PiTjxn1ROhrDqeCAnnIhGP5Tm0gQuoGHtWUyl6PYcfWbUjCDfWP0EeVCyTYBWT4Md0WZA/qpEor1
Z02UXjfemocBepj9cLenenSjwceHpew79iZqXQcQ8m03RcLQvV4Aj1ip/UgEFAx+5OvQNt+93eC0
7RAnfN2cvABBRoQvSeWx3kbQ63XI4cEGANCI/+24I/fyFrsv2mCTv5q2FXX4DPBMQ3LTkn3KeCJE
g23yai6e+9J+k1zk0sUckqz1n/EcnKHf5qiT68ox+60c/AL+M5SrywowXO99Eqqx7gDHoBGkJXFB
WadNuwxH/PtCK4UXJ1rZ1NfanrFREE9ORLV6KxvtjVAYxlsaz/ZExr5FGAYViQII+xcenqKJB/t1
YEb4deOAd826P4Uo1ftBiU7CaNQooHV7hn2Ksx1exHvlP7xLV1/+Vw634ODTq0TrGPO1XrICr0kb
0qe/FUG63fGP6ue9CfqR0+kfBLCFgYe0nQf5F4z6tI+lVd7r2/HE3fyc02z2wRTUCGmZ0BttraiR
Rh+oyufzNJWhAK3jO46XIJMzOqQLSewQ3+v4QYVPFc2V/x7p9wMfwHIink0uZYJ8Ye6tpuTWetmt
Po3r853YXTfc+lVL2rW64rPPFZ/MJ3fnNNTJHJJ07XitBjzlopl4sZPttEn90PH/1tclYM7heGuQ
/nisG3U/XFsBVmoNBVqquhVeea/9ubsMTmEHDdylgIEM4mRa3cDarnMFCqorVnoHfpPfKLJPEVZL
ZF7BTygPVMaLAZfUd9epHQjNk5Loorp4WKshga2yjRLCI/chZrieAPCDE0adBM6WvynicOmYQhx8
w7WOEs6EnW4ka1kTprSO1BSmgWaNEfzTfsLXLcmfcKbrlBXaHmT7TwpncYbxzjalKRxEAiAcE62l
gV33UP9c4SnrP3a1eXiYtZKdERYyXG3JYmp+6WbHU7/HIU2hXDOfBRboK7N30FJGitZ/sG6X/Eqi
HA6/fsmTfCmdGVtkXyzMqO9zGAZRo8Lb/+LHzBVQ8WT0klVkaf8p2wGtBZfAcq27t9VjPPT6rDKw
/N9uVEfIvBP/8Mkx5e6OyRH/aP6+QZ3XyC1TTU/wFy7dd6YL69An5nP4ktGQw4OXgbdWhXv9uOto
10abzojSrPmzCsNhZg4k8CQ8m71JrJ1DmPaH1/RsOQ+u1NYo6GHku3Lyn7OOb6tDvWzlAC/NB9Xc
BDoO4p9Tp4AL+P0B9SgBNCwgVecIeDeCMhVLP5A/s+Ar6GqsIZN7KDeoParm337QsUErI5kZs+qo
WE/JOug+mdVnG/AVKj0dcPSGmvZMVsz41JHychsXEvhuClVVPwd1lHj04n80GCWqE/T+gBe9AZfp
v++ddSI1uw42eZZ2o2pOMQmUNydKElr217/SfqtJPiaisSVJrpfr0/ZadD2L9yUH/7r3IL3nhhAH
ez1ElMzwrZ5SpWqlUCcPfZSCw8AbouGEgD3sh/ReM7J8lMz/ZmmdvADaxpsEPEpf/3ksvhc9VIMx
QKlBvaJp3a0LfwJfAmcePiKv98eGGppPdFkoK55Q+oE5jhpYOqDoSTyhaS7UTmODyxMQKNzRZ96Y
rPSAeAYFYdk6xDeBtxUbHjwgY3Wn61L2GTB1QER2B6tgqkS5algp/UDd/Sdy77/gusmCoGsaXaat
FHMypm9jGftDM4V3XWHmr58wTOHkk+USN+ggn+sabH51kKBvt3ytErWM1xNCG9ynpk8NEsL3VWSh
5/UGemgTqpwKh9GvQ/4wQQpkdp/lBW+mDmX9L3BSjewyam9iyHcDTUjyYjUeqiPJxliNII0RbHgY
VMHDWTb+92BeITbPRvTLkOUXqwWYc+ORkpcE1NePG905gnuZyiHqf8E2SFG+HJGVHTbHd1/dUjKM
+YG0/1ZxvRELbRRiaHcWMIWAu8aqdqTphchRQ8C77VkSrADJnhHCI6AQDEW1qSmJb0AJugMTwILM
T1dPcSg3bUkQGqBRHiWmNhYj+ax1Om7PMWvmiRoncmi4MWhOoNInHoDG34JUjmzicsfAj1Sq7VXv
NqWJsMYYS0XmWzY8m2334qqYN1QXbH0Rd3cwVgIrlxLluRigb0WjGZDMFrumB2qSHCxeW9JJnlsG
CHvci5Sogvl1gYWePxKZYxNVScsJwIueENs6DSOJzWUVo1M1LWhI++KsoVa/Oag15yEuRUF1//iz
+i0syCpa5ZDp1fhH3tQrErI+ww0Vz3ULoUThYCoRBR2OYqhC+pRNElvaG9JvBgwcFSc2Nr4AnUe/
tK88swkii6F0Jkux8/eJI/E9wdkRN0R3pXzLECqFd3yt6xcRFzhjU5nzO1u98QYyt1idQOWuJwK5
Xj1hI+bn2KjRoGZWSK4Px3jPzf0Uyepup68sX3dyqPAPfxzn4UQEYSEc8b1rbqUGj9yqOKhCNPsk
1n4N+DfkRIasJFE2MlcYbmKBpLnjsd9rLZhNBsgAI3/l33kDAM5djt0S9UWvrLMSIhV56gdU6Mpx
0Kr1zAu6oC6Mk4QCX3Ei9YzbPpnl1dX7ZLR1+jXPc0nowzmsQp0mKULd4HkP0z9VFsD7h0vWzDm6
o20v4EA938XbQAJ+NbnWLU7dfJ7LeQuf1WerctVqifohN/a19PGFUOjvOnQFk/6wpf7UA4qrwWlC
MefB8l7p4naSODtmtCevU8RX8jq16YY/iwZNrI+R24XbB+jMrj7IxC8XJMtr8o9Fg2jMmIpaYMda
wBS2hydhGoDfUH+xBJZpzZAIwbUwkNFBw2qdH3H85vqfMor4Us2W/3iw/+2K0KwFnFVukTsu6ff1
hl8XFPGmqnoQB1WZyTlcPeDxUtg1KjG0Qs+QqcqtBE5Vc9GyYTA0s6JnKho+Jd7sdK3/P/OsVIns
AKJswA15m4wej0yg33CHtrtHM9Dm9PI2QZkfXDHt0zucWmp0YSn1rpTN/zW6ZHFiBWvTSD/k/cwZ
WMLugFZNxr252NyO6OT89dY7RLaRTxjGwX/Jjd6/q54vi9Wm+EXCoVMSbimTo48y944GW6CF0JbM
FOFAp0gGdD5bepWCO0zMzvE4hhTnkfMRKR7rPFl3LVw72xA3AUqarAmtpWQbe+Xj/UF/pLVr7MG0
T4xEJxLyak3u8ukK0vM+k9PoSINq2jCsDu+pK9Gt/7TLZomyHwtYCjSf2CSy6BpN86jN04obiW0G
PxEyGVevpiMz1x0Fxfi+h/p3Fzs/ELLa0iVm4eYy25W6wBYH3+YY8lvxMRaDJoAIbP0nncPIdDyU
+LxP8RqaAPIok60obeZo6quRbgAunBe4mP1dkqv1EVPmM8mFXynwrcUgfiz84V0evG1c5KzMLHyT
GvxI0/cLtKv01DzD1k97tqN/nVqYe59NNyRCPl3Dcd1AqGzc34sjp0mfcxdCiDovEJrBPValcKXi
krsMd7alx9omRdJ015YfAowy/c16iMruPyTRU1lgZyMUqlOtNyZkYW1E0YcWsUMHcm/sMXdUkeWX
6nUWJpx5i0PJBUuUMuKddzEIMPYxPJStOt5Hri6IvVGHsPWFQC5Y50hjY8VE266GFCouF7nHq/vm
ikaD2SJmcCJQlaCwmHwuYZr3jhqoHAfXRjCiGpCa0JYN4WZJWRBF5w0uDgKHnVtzmegiuUiSI96P
0X91/JLifcG+ssX4zaCkHpopGPK+GOgAMI1x/U/rLT5jUJrOdtQi4Uf79ZD62ctE7Cc0r/dH7/UG
LUZVfkTaGiRw9We52L5DJU7GJJVcmBeC1NMIkTM7isguJXHchz3Q5srmP5qFAaNCZ31gpk1ygBJI
ijVSvtWn4k4d1H7ERIjats9h28BF5PeLrCT8FSmclgb28+tjLM/eTSoQk/DHzAkNtWn0xAiTMBcN
G+t6DmDeW/hWPMWMmpubE4ad7F3KQq3O5jFGvEn3wTDA5tbGxkhfyTieU8vtroe76eiC+EeI94tp
IagZLHTb4gTlypjizgjiq6c0PzegpWT1rCHZJ+pEWSybPG3/m1uMsZtGre7MQRm6PS5A4Y5NQCuw
0gcMlbza8+k01t/vqPOo5LgGTVWFlcuLxa9hriU1A5eZokyz3hU05FYWmRFbfSurYBGv9jSyDYaE
pYIkJLX2JSNk8F/cTVjJKpEX866HkcP8ZIHNcvhKF5TAZuoZq4yWOGC20/8F/rUuvEWFCxcCE6/K
H4xXlW+ZRTgvzYfpChmxXCDK2tjfz0/wpbhlNWYvhDPCTjNEfN+CVFq3ezIwVf23ikQZlnOAl1Jc
F62ArpjhBnboSL3gXeizAtxHhHdyX0cMBMr7373vgFXUUzREohEmlIfFSTa/+NVHWR4BbSEBtfp0
4XnR/cx/0weOUZLXD1OMsSCJwJQEYw8OFrPwGCx2JG48o2uxQk2I7l/LPNnZJ7DrSApRMP9h72XP
wCvvQAg3aGKLGe7xYf/LUzgWFrhaJqB/k3SsuMdZu2IZuxmAP9zd9KbFvzvjGWV4QM2P1BAH0ZHW
RqnKvYeRwMKYpkCLkLlRJnjSzj/bm9XmstuqOBcgZOq7lVaxI5STG6f8koDGdb4YK53wzupVlGts
C3CF4rrucFrT7fdM+rUTdu1Ina4VDUAxRW5LpCeVWBpKq32/WytfhhLLb27ZFfj4xfaQWblswKjn
E+kn9ZdsMFEb+Zgx/5rrwoPy4FkaZfZNwk9LK0Wxus0kItQdoJYGhiXahC8hpQSp2/LW9iMdcTKr
Iwqb4V6uYCnDgENCUDai+S4B5lI2rsBHIAAhJZvgsSiZq9aa5t5/oCBGPWlzossYMau7USOyT7Bd
XAuNeHvECALd/4ZPxD58qdAMyx9LdriyAiUfqhejK2nnW2UzknuUThj5D/PPzzg2uzkxjTEWNj03
DAjz/laSGBruxvnTg8Uuhot7mUREOW3u7NA1hMz76aVJeQfbtSkpScFVfuyKtQ1cSEdpbI39FIFt
RoQRQSnyQtlwVzoQ1Ii2WTQaAXtVIGtjiA+877kzhOX6xSaI3idqv/Yi3mnjCrviOohdC7mu/f3u
3Wx8XPaatg0Xl8tMb8ggu76+2qD1fiIv/s99kzGyOX4bTxdYhM+OmmkcVmWrUWqBF8qIk8eRSVyw
iLoexMs3ATmRyWTnNN0kFurQJWRIHVd21o/7rEZv8Ek/bMi2NcjLF2gDUYo0oWPqaYkToVprqhG4
Fu7wOJzTO2iJBHJW0O3E4xijlkq5CHViNXMDLr1A6N0XP+9+nCjsVMDMDWvbzkHHQWHs4loa42J9
vH7jJQc8Pc+fGgzFj6dWRBJjJXE8jHSTE4+OIDUICB5vM3IT1DJost4Jz9mdOYYxutu6ULXg7uqo
Bks6eCRoCLlhrin4teHmc9L7F0pVVltfRbXBhllYdFBbTGXN/a7vH0BNqWs3kB7jTgwHlC2OJMSQ
k6ElFJfALDqw9I1GvBECeJJFqGhUsXbp6f4ZzkgERJ0591Sk6A9itMMrV0zgOTp9j7u94zW5DVUD
b2vJsU3+I8IHtTBCSSHgxImY6WYN3hw3kKQhTns/7nXjXI+OGAjqzvowHgfYOJ4vQXJ2RVcqVBmG
KNPSHdldac2AZ++Sxmc6MlgMIqBLOR26YZ6vJ7AhUt/a4J1m+fdv8ONcXD7OmKVuoj1lvvQjVVve
VhDsplSPiX1ug60WhxK3JXB14WapkW0foQOXbZ400srjSeTb2kx06id3o52ZqTDtEMJ6a8g7fG6L
d4r+Zm1QyDNwaCwLOi60nYSSriONTv5jM+AGE09t2WDr67bTKZE6BenRB2xhNLG/DTPMEGs8cv45
al1VUKrErvexPTdSnzU5sz/nvN34Qj+gaOLTyf5ZzxaLUSGgKVtk2pTAdNs0Ypcr1Fh1SLXbf5F2
c9yUyf/YBvJmF6SRMc01PskveTo+nlmNWBEAQPQJ/bmkSBG7P8bwuJSP90E1h6zuw++V27S1Yxmx
FVF78AuuaurTQ5Cjmb6+FEtJ/8ZqQ1mbW2LtRpZIIfBObM5AnV2v3PLG73/tR4TABfMFsO0Iucu/
d2XkKq8gqY0i9xNn1aSsPTxP4E1jXgYRbEHBhbcoJ0uOKcYqW2WMaAq3mj2QeFLZ4ba3R85xDpvt
ueUHmckz9TAG16EEQVJ3Am9VOYa2kEOkfAZsHGDs58ToXSEUncrtSsHz5YzrD0eoYBANGFZKBUiL
wq6Ey3hYY3yhfr5TeMKRe4Losi91APwuw0K9bI4VMQ3mDH/pcyPSDRiLwowLKfSWtOKYoxpi+vRM
cS9fUIYp90TpQ238Amx4IvfbhtLlK05QFYWXFV37cc0Zrxbykn3ssd9BeBYZ2ORPsFQIJ/NEgObV
jzs1agiBxmCykIvNBEihPDhW1Z8zdey4wUMzQrujFxWhimH8Ca2Ko5z1wI6Jl7ptDfRh/8LBJOub
pqgrInh0eY7b44YkOTZT0ADuq07aTdDs/P+NBn01K6Q0U42osQn03xtWAbIBLZHsoLHUsbhM1dD2
FBuH3ucXA5PY80HG/+g4IBoowQL7F3EbN0NDl3Che0UKUiQxNFOPN2SG70BgVLungHHgxAvYrse2
WObmjR6wCJ6TmkP74zYYpQEwAFcV9zbVVxh8zu9NpyQThh+pH2Grqcrr6xKrcrvhQah3Q/2ymh25
c9Ch6uqtmhZ1TuUs7reWlQW/ef/TCYyl+HkFSfczcPgZnySuFzlFCCehfnS82vUveNl4VcbVljRN
+4+8OFPIHwfNlAHPjx0KN+Q6TRWyppZjtEkqe6KW0b8FoN0U7GbARRNb4fQFwJI+Ygrw6wM2V4Ec
szxaeWPIsPDoHopNxcWNpMMaJ4GGpQr0BKVcFTEbKcE3K9EcNOgSDTLdjjOpEAdGnrSNQYblt3DG
dPINot/PgWAQq1GlUyeDQCJjogJSG0H27+XW4gIJou+lwYgmhzir6edqTaRdl/0WkOJUmoZ/3oSt
9ZMxGnaJoJ3/IWl1VvRJyfT1X0R63BeCmnB/2S+tcpruZh4OC9KGXqh/WVjsJht+R46rK8vD5VQz
9tyr8ZxULYmNf6OLdCSaCMSI1bk0cIt0ToTRp7p3O5uK/gwG+lQ0EMfO3AfmenhcLB+C7qBpy+xN
/UjtOnkzwqjvrBQr1oy4Ak9hSosAyR7eW+WMBcgypANjW2HXaL6GBlVUnPi7K3rlAzeN3eBx/6BZ
wreBoJ+XPtWVYxmXUjZBxLF6aFgceVF7s2H0426VB3fDR8/AxnMmTfSWWT9Brdw9+xWhWIzFfM7/
Oti4mEngmbHyLbbY0GSPPhby6f7yCfmyNt2ybH7xBh9cC5taD9t/5YEEyMFStyibRMhecmfP5vji
RS6UclO+zDss1OuL/y74ulXJiD8ZMgvo58BvSVcR7ApKRRAQFfyTGl6DgemsmiKfoAzuxumYkh+F
LWFq9s/lNLGmCwQpwRpmsFB45ys8ArsJkp2YJAJWuzLxhXiO2vNQXpW5s89jH2PmpM5Oi2h1+Zrd
GyVWMEOGpSts00Z4OlVweEs0iEkS4P2wNVDqkEb11cRE9n25FlN2YUIP79loZCZ2mVUdDekDEUTL
xvEs4mWKbZoavWeKtTXMdBfO0ktk5QyAg8+Ptc2lD7s480l0N6XxGpOrC+geP6rT7j3Hx2Jahl/a
Dwx9ygg5ZreZ5jDDOvd8WJyOpmblN2IQGCf5tAhqveOyD6RmnVFuFxUXvWHL2EM5B25Rrpt/BtK+
2orZ7Ih+KErZjHGlWaoniHurpe76373DLR2B4EknQMV/EsE0vlnmyW5ZL7xbyujQ6Js+V4dMQL+B
zfy28J3WgzsY82Gyu7/6LmXCMkJx5HHErLM2qBR1UXi2956EKV0nUJYnNGVVjo33/clkw3MvAMRX
PBaWt6qvdAr7X9Jiup41LJAxLvrMd3AJoF3qoTm2OXu3U4yKtL3GYOQ2nUNCkdEYsCyfIj3ZVK6a
yojF+y1MBfA7hl2IVplTEXNw61+uMCl5I1pRPoltP+8tV7HGlDbDjxv1+JYpPS+Bc5ub8Kh3QyAB
c0wxCdJrDvWaWE8qLOE7jELNWJw+QiqeggAXBNZaMA89IDbm8GmWYYIpaLJevkMWiVFqsgOHEnwE
lzNoI0z5Spi2T0XmQKdknEm9/LfyIW6gR8Linw7r+4QWIFIMwgKWCgzSd+GEgBJDRSOveg+56vqh
gdXgFIZJyj9ZVYjRMTbwkZe0c18OLrooXypUgj3+Txc2wiw9n1YOe+r+5oC19295zMqrGkThLeRH
kqRfIyOOfydgx9k2JxfxA7DP+LMTS85+GQjpPQOdkqwIh+VQmLOHlPpUBLSyuvA5ljhNaZtchc+b
PmzZqcSa5CyDwejPg7QK7WkzG/Hi58uGZzTXHyhdKdn+KfyQn0yZviK4pAm7VMmh80OjRDVB23tX
ZG0G5+SOkSxGqDT7KB+r42MUuj+Da/2iKpOnai1T1jE8VDOQU481zyq9fpY2Zyo3YVJvgBuQd7Gg
YFnKRWKtSEvKOXIHWfaLi2FHtKEIINbZYwRQah5LfnPKahUGU3LZkFy7oh+kfnLjxnuVDpWWll0C
AagAjmmL5QxDLzjLHAXnwLeD6FMDJr55YO3UtrY6sdOKZO4HfWKBNXcKYUv5W6XBdYZIpeBpItkk
uwOYIQifBapt2Rs4M5uQ5+AJl7cCruUNtp8Mlcvkc2BKSlQNZN7JsaJBIEKk3JA61LwckScvQA6L
UgOWHAkVQe/W143K/XqmthSsa/zBr8oYol3/AAZq1bIzKYbYtVwRJYV4edsRrv9+1eekcykMVPOB
lIW9cBP8GWXoc++VUC+Fq7MUb2y4AqqgqkKydtDHbdgusAqFdjdV2YDo2lYRCO/FtBohVfoLqc0k
PmXg5rvvFxK6Rf48qbcth8dOKxhkE1Kv7Hr5nwWm/y/8CoRTGUX9+bizwitd8jpU6lJobFh87uL2
gWTFhMbG5ncm5B+dBUJlDR1QwlQqh391vZe+ZDaKiXvwl1oMugr0limN0cuLPma8bq9bB8U5aQbD
RnkuYIJepGqoGyHzWRSGxVpBHFgyCpBy8R7EdanbGHNHChqBN0rRTNXIXhctkREGhtiDDDr/e6fZ
MGar7ds6M5QO3bDS1eo34hDONgPgkwHLRsnxSx8eUP2zZOuDZyAjjqvewLgNNd5ZFeIhMexYec6G
RtTtggu2KOnRLIIPxyZauOiTNhLqNef1tdU7HW3NJmSQ86fS3qQcNtJKDnj0ohPuctKvueAiZCkO
oWGCnIU0Z9HDbOW3yjAAofO4EkKpfdbeDRVk9hrcfSJqXGI/ZAlD2GTkxjiIr5zFZMjf48frx2mX
k0jgtqhy9MZGfu26x1dzOYsjk3arzIydaPUdh+XTf3bKKLDePybOeMKjLfjf74PTXRb6mZFxNOP4
TV0o4h5C6MN8DFGWmCWgNv3Ep5QeYujeWguyefBeTt7P2e4ReSHLTuFocP5ffQWQ52Qtlsa2R+yM
IsqHlrzCQHNVqZESJEjPeqedYBQA/pC5UhAMBPw9Q4LN71XCtAcaoJDbtV/b4hYrcrlLf2+T5yWf
sVXBVy8HkLBnaHeuLkftxA6tqNq0Sg9Yo7wPwjWrB8N1MeGo5Gr+sw1qe1Z5cIgMQpyOofQyJ2FB
Jv+CgRZRWMZiyhL2bpDCjvVBIY41zYXTASx8GoRd/FRqonJeuqrr90STpjOZgTOaGvjPc9EQ4xcr
6mlqKo25bKCnQqGiS8jpxzE9WpuvNTzExF4aF4Qq2prttBpwjYvMTCkNjWSCbZI0pOZogDFH9Uyo
0zcgtYy6b//y97hjm8kYurYRZrfuEG1aluti9FjM0PST1Eavr82PvkM/QXQsqXk8iJfQfvnwTEjK
s3Bumawgd8APmF8XuCJJiZ13aWsQsijbPVKCpxU5pf036lJ2gwari1LgruIUJOyW0DQ+4tNz8Xrg
sHqeOiq8a/vOaJbIRPG8N8ACltfyhoB/oI4OAgdSmFqUdRPMVv2rL9+SOl4eZHs/KEN8VsxeE3sI
xYpMLFRPIGhOEKkiNaTbZ1C/r0Qy+9xPPTCr0numXdPSqdlkI2/hCD2WKbhXdmZwUzyFmHVR2pc9
ifswGecnm9Tf1p9sefswduOpSe/QANjF5c7+6MOy5z6NUCv20rIVvkziHGClusi6otU3+JTXd0Ts
g52VjXtW41qjCsf3sABo8/o/LUnKHRj8VWLMOAGJyPzPQt6VKcKh7Mj6WDVkicH1+i+oiNZIkzm3
WHCgxtWl3a7Gcpb7XSzsKKa12OkEi8EOIUEFgKyKz2ziLHyYd4nBnWj/1kaTI2sGrm7AfuPZbKJl
sy6aboxwZQDBv7c+SPVBD4klB084QMyjq2oG0zHb+jK/Mxca3+8v6D9+qiUklA4L8MAgJEgZpCSa
rkAGKXpBQc9gyqY9Vis65zdCDfGfnhmypI0uc49V6ZmduL4VStsgQxeS6gQ0uxtYj6/3WbX3rpuw
7sRBB4ajoBWqKzZkNwd3zND4rwq3U7vcd221TN6XIl4ox3A+B8kYDnhjDKOw1v2wA0FDRpOg0q4u
4Wx0V7o4Uq5BlQrwVXarzUdDYIhQYlWMBFXmu0Px2l4PbZEBeDmfIPTolXtxJhxg2l65YMxSAUVN
olMF87u6GMahE+OPbLnvjnY7rYJk3OeWsHTYelFvfAnfE09JmTcSfaB6W45tTF+T+DWIj5tzKqZi
wqXQ10HfJRg8o00tYqOD6Ao774RnbFi3HgfI8SUAZdDO/rVUShMd8Yqw7cTsUYVMP6Tt6emMXq63
QY7viEt7vGeSI0VJgw1lT7ng8fjieldwYK0JdmzNeta0oy0N9KG/0FI8YpUGcA/oYaYFaO9mW+J6
F+YcaZ1nLLIQY6jwBtk5fcl0ymeqlsNLwMpPHIx3V5Ky4TyOaSbtTZO3bRgHTGItqpJnMtn+wjPA
UgEPMs5SQExccUL4moB7XviTsonMi5xpFoqsTC4meTmoZ2IpEIAlm9sW93T7lH85yCocAsC5QT4t
Ukor9W6N3qomEHsmNx4Oqkh0TWg7PBbakxTIBZ4SFccl1YJdWzbG5A1sOqAiPqU9GVAyAHjEq2np
i1/U+OiSbAD7hyS91gOwqG599q4Z/qdUixcacopnZbQdKf6gUpXbdkb4rAAQbCZVvnCnqD1iVVwm
KFGEi1lGEK31bfIxR1pCV8Y+9GiWIvwcKX9aCjmjSkOf6ZRq9EG/X+Y+hd2toU7g8pRrj1KnxWrO
t5Wm+KhaG+gIvsuNojxVH6lmewu+ta5aEwxUc9TjZXWJXSQ4dhiIiw//iniHQIaTH1kkKd2f6Ssu
R3Yzfo99KZHglur02swJhy2e+x57/noXQDbV33RVAXCMC1s+rLKTTPsrbjK7EIHi1xv4G6UYypGg
Ge4OWEgkel9LWFiGHinkV9nqiYPl6UvU7/nKO6LiUVzFahTI/sEOtYvPvJiQoI8Vm5deatet4h0z
j9Cg92GBMHdaXWkG0PpsKOg0bxX3xTagPY+SDolD6paTeq8FOeqATtO12i0Z8gfb8kaRB68PJsDJ
hUBIZgW+rzvNHlwx2zRxQ1jWHDP3ZJs8hf+UqXsOBA6qEVzLsvKm9JX7G0KJWjqJkHlAc5uhNlHO
sy9wf+QFIlq7MNetAnAVIdajECXzflPJNbPeATmNntSIiK4uGVF355f25si/boRMxzoff+c+S53y
tCscoxguEruUiw7UWQ1TinCL6zUCQ9is9WYaVMZMVIF+a8GKT9vVMBblKBhjaw5orqkL0XD7FNJO
TizePfY9M1WgO8TjC53QpppmT1eSCkTpnI8BSmO0pCrpZ1nR/Smu0ForW8lwIVx7OKK09pwiO81+
GahESWaqnXHI1/+ZS5tnHi719Ujy5aWUjcqCP0KBAASekWiqHRa/N7GrHO/msUNZIjIt+u2ztTEU
WTCn02hsGNeB+EqTBdzj7/HQmVtqecntrU4XE1Bra1iNq7PryV3LlJY00lbt3VTkfQA7jfchc9SD
ODZPFbGNGljv3bgdTvzixy68I1Lz66/CkS4qIjMnS5eIrr7Y7/fr3TFXmP35Yj+YohdKNFEnQROY
VTbM2U+m8hfUMx0Pqjw8Wm4ZRgSPIr2kQT4heck20L3/o98tbloJZavULrhBRXbEUBM3vFUYoszF
4PMfk9KGtDkOZQpzHSAJnhu0HFCzQBNWxdeT8fLFl2zYkXBAh5wpp+I/5nFkcFyKA5LsVvQax+Mi
VPNpbTqjlCBbc2AgfXQ5Z5dvsuhYzL9yX7NgFob3QZl9jMMGbsFsVeLJ58DZ5bxg14wuyrnaCiSf
txBuxSH7H3Lnt99r4/fg1YnRAUhs6+uMV+LJ4J2lfUBtAdRV3cZJGyepiLhCqP+q5g2OoiwGvsTk
BcJH00ucffTofRBgvoEj096xRFqkYg5o3y7vygTYqbQkgBruxWLLnJbmQW6kYSBTts1TEOdj+XwN
9G7u05m/LwowLpyyDNDGBexlGGV92jA4/DlayZEJSIrgSSsui4B1yW1FqDo1GpkBKOs+yDGNJwoG
21pQU9t5KqpW1CK8YFnyvTt/g4ICbFPY7OuekxwHkWsA8FK20eg+QPf8jFzf1LybvIeGXgXfuIbQ
WJaT6VAbrqWBq7MElzbcjjTqZlpEu7Pw37PlMf74RUD5NkDX0vM9uGy/N0bSzRSqEFVrJnuZJ+Ho
BJ6JY2vXfrmCu9fiaESL6KgnmB0n5hyNs7Y/3f08Qby6hKu9xY8Jl2EMHO3cZQ1evUUVnH9WOAqA
//3L4phZhvhB3G72QJAWRFFxXDXCp6yhcdt3DmkwU0A60jeQlAorU+CPBQy2X5xOyLE8OD1dnM6j
omqEZNL5ErvY4zL7wfJ9n1S9S3PVDrNhuWPYc0ReUNmHp9jbojCqo9HDGZ2N6hgoTFpOt/nxy+zC
s2NgHSQrLs2NVTHM/f584bodjLp9hPEeonBDO49KOLLRVJA6dBysMI6QK/kD9Py0wbRPhDkVgEub
EPAmcrhvaKA/DvLIDU85AIRoDOPw3ZUwrcpI9kVMTy2TNstEaCA9rTSm0mx8mQpFB1MfraGlCFdp
0Qc8ernJ/ZLty7bL44ynOzI1yavhlQlTmLuZIf7Yzbt60VibakSDdXojbSsoQne4LjUcMeqSUzWv
diIOUROHuchgINrUYB67u9TLEbwdcwMnnykR93ckVlifD4oXCq/ACSzav1b+2wwvnAEfYN5TRQkI
hUWgkyWJEKIhc/kQj8ERlZ6rBmj08vAt/Rk3W163iQuhUhg8rsl0sJKPms7f5uz6eQq0+m2nzRGf
Ca5+53auQnBM/CwYc2ojCqQYjJf/edqcHkP6n7mmXWWBplwWizZDfedfUUNIUtQIWaFdURrxcDkv
X60hTumwsxzb3bWaM1h5dco4iHGyV+0LsQ5vE2O8CAku3ZwL/NIf1sSHCQqnRhA/TBaotukclWRx
xEbVt9ymcRJM7CCddLAb9lhOOHR41a54aS5kZCzI7txGULD61Q9kA0NGaRaxGznFnzO5V7/lBQzE
dd8Mn2d729WydRriY+hJ7vlZ41f+3L+cmDbkDhLF3c6LxruPSf0++UlqqOSwjLPfxVKv6WYbXlDg
EaaGyKQBwyIgssYX9VgrKKO+uS0cvpLQgBSwHiPmzt8qC0J6WzzuwBJTUbdGuV64jxBo3tr2H0RC
GiPmMUQFc6lB78xb2nQuZ8KIobOfbcMYJNNZrEnU4o5u0CtjpS/VcLDhoef4pBc/x/QP6+O7MhCA
I5cpTgFr3vxe6E2wS5WFwq5ibPyEqSqOYusrRN28oPmDBoE+PUFSyY4MC5oheIQROQeJmYpDL/PV
xu2H/XaNX5HQNz7g1hdLhqOX7ZXVWswganQccQnLvWK0OcbATKkeQdREXir2cYEQtGpFWE+q5GQl
6EUWLX4y+du+ytZ40f/j2E1+93Xm2zCSuY9i1VmpE7QbbBnWWXDSoveeP1RxbGOM+l5+N+7nvR+U
czknTMpe86cvRqLUM7at+UDqaXzlEJzmrV7nu0JsHfvMDx26esyorHCe8D6DQYvJ4YmFoFkl40wz
lL0g1Jy8tYDrtdiD+n+FifqP1GUiiWy5L5lMrO9siFYbHW5zU8NeTEt/eXHs7L5GhcI2v53shmhJ
MoP8VT4jYWP52Mx2u6V9v4DA1SCSV30T9Xavr7CaejEahxJcYl/CEwp7Wr03MZlsPRjqJpJCRNSk
7aVJ070VkT6scdoU5jefv+P9BC0qcRYJq4tnogOplU0FTnSmtnWirndzQmaUg68T1/fZJiCVbsMA
y1W/yDrhI8/w5UAM/zpuUnPWaIZOTWXWL/1CvkfxcxoZylDbWHdAdlgWEoSbxgBm1eQIjkjB5Meu
Rtm2nnxpJVdu1SjLUU8RfUkPjvLxnWjX2S1m4nU/s+nsTWejgBce/LKsGaOK0TEgmbOsHzD7GEAd
LtwiFPWDUuTKFRxICZQD7LwkKGkPxDzrbP08SdIEuMKliKXSpIa8zJUudnsxJIwpmR4QSla6FKU+
opNb+HIGTy9/J4H54U6/pAh6fHSPi991uHmb+tjgOSFRDSkDYLzGk3FuFw4hWP4J4A388vvxuJCs
2ImH9IE5MnMpughoMhfrcECsbABEMR0/dkXYOfjbPlvkE/4FbcZwgAtrUEhgKvEnIDCsZIx0L/TV
3pHemTcrEC7zeufX7HsG8GDj5aHmnx8n0bhTiGePHbkl1Ld+VI0CiocptHK9DQZm+E+al4/KtlzR
7Px3Ph+sn4wm/3EcMXNbtWwFj6MnysoAjR3WIMRWgaF2ZKMNra9+PAyyNdiqy/QGQSX1wGB5QNg9
HPEppIHLacfzL4y2BSZd/Se74VsE9w8qH8/YgCm9/G1mROQzTL3zZYIiNNbFOJYnLwkPVFTD8qty
UT9Icw1MLJDBl2Kn+4ixMO/SuMfBss2uMJYu+5yU7nEp5fUcJfH6H9fE1dk8Uwqpc9x/zlw95jZI
AhFWCmx1dW28qeCmRTzD7EIbBzhAicHp/S7G2BbyklQknCH/DYpJzv5ruJEzOi3/r3abtBXnDDdp
A31l65FKJRcepz0MNX0wlWVu2D+JZllIm0S/9ks8HXrq19Vwllq728vgz5t93IUYJjteW6VeMTcz
vv/KtMo9gINNLKLK5UYH3fQcqVToUg3CPmi1p01WZ7n04Zg6W00cUp1UHNxBUsLtEQRWa5+MSoBw
u2zd++4OHtNEOfqRibq7mFRQVj1C/MN29QcGlC/3oeCZmgmhVHZXAdrHHhHWRZs49sPGXQl/wZYA
ewwSOshlfDhH7uaLpo7MYhfTerRvErXi83sLeRxQC6gCX6AIrLuVk5DvKILakB2yFSw5Dyh+MxDu
07/21enwrOxaMStF06jI4/dukKrxixBrKXlu0EKk1sgqiNyRnJMWLgKciWLypBocem5PIbVH1RUr
R/P7459HuewgKRqgO0Bs/+LAcEK2trl8K8zDlzuVyfpRQQrWRZslvjVC05ZihRGiTTH1G1iRs+4G
04bGraSTcSy8CAnpFk+9d0dsf7FppG0c47vy3EYC1OXcz/XbgYvWkuqj6EaX64IDA/TBMnmnBvAk
DzjU3fvHxD8Bx8bWTofw/y7zoNEnYdfNc7pGQ5KbXE+tF6WTvBAI4R5nR8g+y9w9ueeCTovq6FWF
erSSJ2sHPLxymrpcCO7jOvvFDn96GVyhUH+wIUGhq4xv6X6sXu8h+Ick1cjpBojgX4KcPvPReo5C
Df9kSlAePHs4YNychQxofQwB/w5ScLakk6ZzA99OTOOG19bczt8XKk1UiU2rzUmEcH3mI+DTXU+3
xQPnJMLTF37ZYI5gxWz4HmPniXundlEqw0YTRvndnqqPAp8SRaObXDu0UEZ7DCeJsPrEO9wLQLkw
qhezhNueXNfYblPma9EnDZ+VSnEAv5IgE8iYkcdSvRn7F3Q2BbNp6ziIztb1OEQ2udhDRrDvI3xq
2DMCBchrvdMaQG/RV9Vd2ZMgD1XIHte5KCkrQbLbPISsVpNITEDAk3Z2BeveIafQwWMEuDsG1k2F
HEjDM18KLJbGP6gOMTcIRy6kT7d39KNWqEQ4dWX0VLPfx+iVIQdfHbmf3Ck+LpJUx/HL2i7QITKg
peRFn70Fn2kKjYv84TZJAjKtAtP10gNihf57HRDGWT4T3QELu9UQYFXqn3qCIwBAv6w+zygTcfD5
DFQU686JAXxSRTrlX2px6mkRMbTjlgtwYA+F9fRov2ZVQ6nB/W5tY5x2UvlJ9ozR8Fec3SAx6Y/0
DRguUOYlbIM972pPygk369603tbeqWyBaud0RuPzpHEF+lolQK4uDbR7UpDqg4bACP8zlE+gNkF4
ZLJbtERD9VlgZNZf+KSTvNRZa2LXZyGLYkFS0hLQjogIQe7F+jFWzfLCvH1TjHu8Y7VhGJ/dLJ8n
GhZWDmPGLObfsay0a0TOJ20UU3UepoRDPq9Ur/DJUoGPcATZ9MdzI7RuuTwxx+CrWiwD7j2uXzh0
yfzzv78qGAjruzJLnM8gOkYVEfLds78QZCl5dyL/qiPO3hD2uwQJlMFHUzk2ac7NLPxe609X72C3
VtL4uaYeTyEYmW0BA+cmgM5SaAlc0QkpKQ3cnCApG3im+mTJ1Eq4Z3eLfxeiXUxkE8pLHO48eyco
XjXbfC3kdbjnGZBUXS72Ox3yJ7/CgcuwByTzDK5yKRj7S84pQfzhN+skmL3F2pzuSQOuqKArIF0J
H3JgL/MjjLd871d9nOicOKIdPqRT2DNCSu8jn3pLx34cRGHCMy1cXE6g0le31i3647EEFBIuzP4V
r3UhHn5VgHnhnT6gHvDKVMQkJbE/+ZfMipJJYFWG7s9Y9s26CbVZhpLghfi1dn9JgCUF5U2h/FcA
vG0bbwagqhblHvse4WSMbGY/YtXf0K/KX3b5ikE8uH4xUjnyeo6XDWTRqn60OQHX22tymPoDAFoF
WOhv4zJIXdRiwoJBilFela7vLv+4cuR6pa6kjGO/VezSg/Nx5UVOmy5jRIsLuliF/VaI0B2dgpZS
Od+Rfj+TnyWXr0gNxFK4L8O30fdEppfa/uJpFW7pvMYAGtbhPDqcKQQoF7t6XgQDMRteIoybzrWh
O9ncJHJNuTdgFtADIyI/qC2XOt6JD0IALxRZ9Z8Dd83kjQKb6had1crocnjBlAKCMgQJHhVBHFW6
W1lbOnbxzTCwC/6x493r1IPL9zAul4I8M4g/Wz4cuc6Mc52GShk6gaVZGa17ObN+yzXs0OxHoQfB
XkEmvs7yhdze5m1L/aOGS/v8HJOFdIiN7VPowod2zTCtG9EbPXzI19xy59LluWnxqD8fNUuuXM1p
GXkjC71nKdLQguoV8pmsye6JJcuQUHHIOgRBlQYbINj2e82YJQZm4bNm5RQPvkvofW4qtdpyCKUD
8QPFuIp/vRKVGngmZ3Ceyhawssrhb1ghb14sWCYj5SM63AMJBi08z3jki9D4YhHKxjyb+r47dV5b
f0HppOGrh7B+4gl+YuDqaVZOEuhXwJ7DkWn7nxwbEk61sqIdaihM/MOlDYdLvAp5zmrpoaUa9S0v
T93/Hs4smJxqcF2Cd9HXEYeFWVikXFjXruSDFjVBBCSjXPGCZS5LBz+Moas9bQ1PmcNLm8kY82jv
C0rdkWusTPOAle7Wp1oqbXW6qYCwvbvLURZ5+hLKzbHNdWXFbHI6bDR7ciSOjPpvjfi3U3R+6nX/
lGPtqGXDZpWVcMvCINBj+gSs+2KESukBsiY2myRG05C3LsDrclT6WmaMz+hvaa/QU3Pxz07CMzU1
u7vLIhs5COslip4wzk4MIqCk/vjYTglt/HbsQ8cO2ootmBshK5b7TsjyQTiVwt1HhM9rFqNCBiRp
WFVUoXmhugjGxDCF4w++jQkDWqdQ8SJQxSbHA32SPQFUqNF6emwDS9Q6IV3Bs51x2+iMCSp1+FOy
1tya93kkHbz+/9OO0BsVYkSfxohMxr5weQMnamxWooTLWSvSgxVLWg9DIEcU1KG7RbgddBdrpZ2i
9TgUFV6Da48THb03EhcYYgIzzjyqN8kqsMvynGdotHBI5v5aVj8iOGeIsesnDFJJKm4mu2NN72a/
CLBSFPYO7B11KmjRH6/LGy1qiMvPDa9q1aRX4lWYb3u3pjN4+v4IBCFgjt/jKzGKXq6XsZX8/tOn
Jwjf/w/qOj9U2R4Iqeh3UL+M7KeT9R7j1bazNxvtm8qWmbyEzKWgr/YEGO1v1fDibKfkYupqI+Ew
s/u0Pt3rIEjU5VL1AmK6RKZ4Tg2XFk5RT9uEvfqvtFyCxe+SvXTEiNouocXvLbvwTF4yqCNsBG/+
vl93tyL1F4XhXYtmMEL58EEita1ON2v0ks8SgVWE/pP7Af6oxVNPK0SirdZF9nL7vX4wwDfJOhN6
4JS8rZUTZxwnASZRgwP2ch1h8X/S6oDRFF4IfAETb0KHCDyMLBPBjXhrsND2MJTQPQ0ozNCZnckx
NP9xn8j4F8yromTIO2MKrd8pTpBCrFcoU2XwXd8/oCdvKTq7dAO7jmMEDaW9e5fiOoAolqOWm/DI
YOiZ0mBTh1JfK810iYpN4VnIwuCm/EHrFYGyT9w91yrTCrA6tF3mk9ZxNd5y9maRHnMyC6bjOgil
OBdZJ5U5mw8+76Xts7jB1VcZx1uE1u5bnhXDneTLy+ARtVkL5Ij5iz7UQAjkW+ST578YGgQ9R2QD
tQd4rkSMUY9a+4IZoIdRAcvyz6q+qjbxH/jr4NTj+TE4bHYm5bWEa56ki/Nd4gA5qpNn/Bs/TEt7
qy93lWB2WAvLh0GY4nfOaNWeesLzFWv//hA7VELu5TpyozaG71rG0Qe+a4HZVNzkx85LIMqXineK
pEjk2SpSvVwC4EdkQIyEG9tLmP4bgDRsMVEPbnMXr1cotQU2T2BzZgn1kp1aVVrTwnA3AAQhqeNI
91EzUaq03HFSpzoYsdPUNI1/F0/oHfcalCIfD54ipKT2KwaAtdZfbIgWvpFg0owatKKMsvIHG7ke
rcAzTJHEemOaxcXI5Y1kuXMqq+N3zJZAyTrcSFsjwlU1UB5yhb+5uRUCw86t9BMcX/zBLhKNaaxO
6H7BsDQX/8POnQxZ6pkUi7viKBYYrORJ2owUd1zSGNMpKe5JNzC/2ukfwh/VHHjl5WGVnVarSwFc
oI+M9kVsGVMEhC5dXH5aexL+DCwsyyn3DZex9uG6wkkR/+0Gw/iR2dX5LMAZgCl13lbnqEZ+Us4l
JEC3y4r1IahF2Wv0WBlTPQkmmZzf5xFVt9Va7oBYJDwtG1Ec3SoC6kD5br4Pcc9+ka9qe8g5gzXf
YTU56yqNuHFqrjB/Vq4JvVZl5XtbxkiXlNLifUjOmKx+77or8UgvQ+QRiTaHqoen6EniakXvs+WZ
dNQ95DRHpx4SUNEsoXdIMnRtoa15KegTqHNJV5rkRC2oze88+zgtujcBgNB2BmMQ5cm48dKsSJjU
oeWdz2/BlSyTSjqXlrx9DGEG/ipguXqQTaB1N+VTH9BX7lL+LqtaRtqBMli2z6BNp1k2LYzpp8Jg
sflOJqq0TpJ0Vt9tn+e8dZMd0h8Vq/1K+DXManfUS+N1XY9UoSLXn+EiGkvY3kgLUSk1asg+rQcM
XieT3DHzd2pgH1BcaBt8KRo/p3g3800pMEtSTvwTxWHMa8VOlPhHHo7JBE7JzQZ5d2Nt/qAkX9kG
nb6W931kG/cFF+gA/56H8SchozHwBH2dGXkV29SCUQGuTNIC0qcTBpA7A+vFGrE/ogfp2FlcYQf+
MCsU9Xp1GgP3WfDWqnRlDBRqk+WLwS+ncZ2iqeNXS1C+4jNAViFcr4R+tAb49fpCP0UhrM/OhPUX
y5BmUd3pAMriBOKBnzo4YdCr5/MzFqJg7ExkEoEiyKdfGp86bGdEC9XEM1/54S1C67HXE1unUiw0
JJBJpsOtmfccuMqiQFBiqY9Los10mara8eBWB+7WoDex15mVWJVEXute6lAR2CbDxKuk9vwldm6T
T9DaU8I+xFn6rkkd/kgCEHKOn3Y1HfkE1tI416Nbk5vTrNhVJwh+gEwq1BRXjZp83PGEisEaMjIr
mxJN62/fxnxevR/ZDUl6SqHePo4YPlOdTld4bQXVeaRxLZohZ7GsBv5hrkt9usoGRfPMfa3j3R1Q
GvGHtQ7dbzHX0ajK9dGOCJouPseyPlp6CBTIQzO3NkilXqJh7uegKPsif7+Yxf6sVPOfr0Tp8/dZ
WM5rrPQFjiTpPj9UnLUA1gsQqbggVenIu2n4/IvQu8/yX0Oc0hLidS/PnII1ZEPcPFnexsLMrUJ4
2v+d6t6TkJGZNv4i/D/9M3+fLSJB2as2KrsLwxAtqGamVrKFGBuf8ihj95uWJ85R5EUfxiaCPr+6
mIxthTCDUclnImbAf9yzXN0gKbH+HR0L94uVb3X1zFyKxj31P9zxQiWMOZKRwgyXk5zbYEt0M3Dc
wV8pJoqOuThFxLxl0LGZ7W5yloJSHfOLuJS1Jq+61+aw4o4m4sgeLfmFB3KMWE7otz9UnRu/bWAE
UgGCA4pqhwNUulF5UGOt0pn89WM7lHlNuvNXrXMS75YFnvwDhMmUSNL6SDf9EcuxqXzQgRDSvDI8
QcfzljJV0MCANmeuJxJFlO9Fv8tdJRhibzmAb6EWDlJULk2JhWfONQtKq+eKM5pTKTYQ9/qv18qP
n8ORxpB3HaJTmVJo4xQU9W9hbnVQPeKZQDrJjPFoi8mmvsKDdQ4nT62EneADKjaNBevedMXNnkcC
lWMsoFsr3kSf9Ck4XGFlivJT9Dj9vXFAJt1LzDDICKoAMy40szBjWExXszOywyZJiznBR9RNVWrC
/dGs9Tx472RfWvOLZ2M9aruW/geI04uhTmQJAgqsisbF2zOE/lEZLuyJVsdNV4UwJts3WlFcp+40
mmhJZ+VwGMxN722tW2m4QPsOkukn1C2mw6C+Zt2OUglRlB7kZkXJEbJ7fT/CWlmr7/fqMvVP3x+x
ExAYNuLZrCeAIKaCw12ix/0iXBShV9pSHd7Cxi2pBJrg6GV+ZZoaMEfgRSjEX9TkCAR1TE64/A03
uBMob9QAUMps2eQh2vCKu39nhUvU8oof6861E5nVVPNgP9Cczp404aJOmwRCjqDV9qnoKNuN3CCH
RWBhpHSAgHUl6OpdB0Ehxs/K9+tVikrdLPjGSJRNMOOsKBwKCshe38Qx0NazOoazq13ejd/EstD6
aKvfZTDj/X2NpP3q18Wwjt9PNr2IWY0xUdzyXNczXUwzqahL0SQGwKRbQI304jpRvc1AWLhScw4W
fugnBt4vNIiiTKvQjh//imHQvDg5ZEG0IjEOqxhYZr6TZuQAH/6c3uYQsU91Tp+pqDAFqZFjsJEg
g7hgD3BomoRnfjETKMf04D7YLiaJ2rAkvUgZ0gvW0MfdpIeG+hB9VPiEDPUsI2Fx9tU05oKhnagp
a2tEZdpxBdOrj5WcB0+14zLK5h6Pwr8lFpZ15ANvl3H8keNvPj3GyGpm6NPZbwpjcV8slpAt/Nq8
SVjUTA6w6QP0J3DmlTQbMdxQMzjEhzzZNcjHNdYYtQmZHBuzaEWVnxQ5RsXsuNubWOYnGwrIU0YJ
AtpW5fXX+2lsGi8z3AvP0r6HjwkmdjbVHu6rzvJQbQOZbeaknL7K0PLlA1F3W7KKT+GH9tDYQdNw
/R9gIP/u8LdNsMf+f9eL9lUYNaUZNe27OYyJ3KfzjPUc2w2ZFz1xGfvyp7J+70nrRTpXgsVYvK3N
WzrSZca7BsAofNpittA1O/NmFyqr2+x83NleS0oqJN1zBe7n8aTNIlZGp6yXl1SO1va+5w9u457u
yZDC8M4EnPN77Zky+SsRpM94//Suae6pVStjRCWVKxIqX7xtqKaxwu07FqEj1aEMTigNJ6ftVmVr
zRV65aPI0mUpxsb97jBQA67+04LooMAXiHJk1IHjBgEFgVrub9ZHvcN7tDs3wuE92qAT1NsVwgi/
MnMfntv6Ua9iSLb3mKIPCOCZOmdzPvwDeAZrYl+O+jHkl8b8aG8Z7pHCH4FpEMcgzSO++EE1gtLG
wOD+7M7XgspOpQ/TnZqF5kYyVjl6QOxurhbgFtT7FsfNoYlf+nvFXlHooEgC/9jgU77DNnxTdX9K
avqK/CwUZtU1spfmBwsuNy1iSQGP8NNqtAeqN2wwQIIuWTo9BJZGGYKBOGnukc3Psuf0xGm5iux7
Fz2J0TVrCVsTVGoEkjHnOAhQ6KbV0b3WbX5klVpvjuZWQKTGLnSI00md7QplR0t7jY4zFTKEUyXu
1WLBTtOqO9S4mqZVAqXLJT4xSZf3VMY9IrgZoQupTtojBtFu+9AfjZXkQCgT6e05QWi4NlSaX20p
ZzL4o7BLyJvdkoZ9jUzv+iIBcNUH5dcZYu1N9njbJjA3868fNdOoVnctjahuZFCx2lKEUYnTV6GC
RSe6zljmhvaq0N7tFuJ2YMk1+2yr0y9OS6TUj2zOkvykNG52rHgiftXHC7zCDsiy6vIHgbZuE5Hr
tcmfLqTTBhdlF1skwJMv682luewrBS0Gsoq2gQ+llMYeuYZk8k2UYsRtIz6FMWQefi05aKwsRUxD
er2PYlhnWByWFAcuTn23OzW5Bx0/IV2/8d0vucl34L/+akGbWKJQcgh2wARzQGLdfxdoi/Ne++kQ
7faEs5kBTcLVhhMFVn+RpxzLbrpqSKyxyowsdvxIYS9zr+n80dg5QVHicadSNW5/EH+YEdkLWZoS
LYZH8sNhV91BMBMwALPGcMXmigRTLKRsw1CeectgtO2Li4C0lxcKZYlqyLb+UOOpI8Onky3I0XiW
WyuYnJG93EM68NTmQy+tqOV+0RJ/XuArEVjLjvds/xb0QeRoTjg9VGDkOya2JYZeoFVo7crg030q
5EtsXyJFIH+V9V2Hshh+Xkqmw+n5hzQ5UvA04LvAtzT8Q47qEucKd2ee9Yd21vLAPSp36UIVNDje
uJzM1R5ppLh5V0GUoxMJIyyikygpRPGsjZtWcaVdfaXyKcLHIQLdDbAFv1hRJidUJYMcRYDripWE
/Tun3kLztgI//IcktYkahChMqsvHwfKgBXekOasz1sT1EIWw8YEuAGGTgixtVlirXKjk23F9Qul7
yfasiMLxRWqqWVqI4UpbCrO9Tpjy5bNprc/RGBte5o9ccKmOt9d6gJXV/5s54RCysGoHYjF6LnOz
nDgRWagqpg16HoRhthUnfS5Xlx2YooknFHaEY1+Qh6DM9BZVVRxT/KotwHGvoPQ6mcRJCWX9JdWD
3bg2KwhHSLfrLU/L9wsHo41O42EFMHq2aYSsph2gankfoKZ7xdmqboZb+cmuoC3RhnG3iUWDaJGy
qQdtff//x+lw8xAJn6tLqD0lDWLD1RinEk+GP6rqopou7cR7iJh7o88v0Eo1MqB/Itr90UXpOxC9
tEaKRzeYUcCz12Q6I1uiOKXXz4m6U+/YeM3b5CJxaLD1XherLuBq8rTUfPQSvmJFeIxH0bzl7g/B
gzEwdGRU9rKy4qpifhIqWQlRyfXG2xiJ4wzLS0kIuAkCN36BtYXTlfIgRzi0Po9HwY6euiBP+DNF
Mlr4OgYqbftDE8iUq4IeY9UyiGMGGDDyNyE7IDzq7jo0i/dwYj4kNNGgLWMhhBeU65R3HGsVVC1Q
J8A1QRnSfET3eOi/4a29AoRTyfWDX+rbxdipsXDl1ZzC8TXqWzE8jnuQpxNxiE9pxli5gVOlyKDl
/2IZlmlcVMTR/clfxPtMCh1HFim2BBbplU6CGq4L84rpoZRsFHW//cz0Rh42SLQQ+Ua5B3Xtp0d9
4z5cu2l9gJIZPLJYIkumF6k6xbdIAAUQmDh12l1ZSjBNF2cnMmTVQTzU8up7DuQPXokYXbnAFejr
GmBNrONr4XmvoAoGwBc38FpkFv7UgAsKl5xlTHac4HvH4F1Ta+o7kEz2gF3jqv+PierJqjREKDEA
IUmmshNr07sYTrPC/TBo4r/homv5ckERzJcIFIN925h1SIXLA4rmk8Itndftp22raaGyZADCNRIT
TNNVtlNKJLlQ5+pZ5aMyI3S7Ya4LJ9YPfVGZVrjeMq0eUUMrjiKzBzT32O7UonltxJZ/TwKuYlLy
PGSZ+gBHn0YRkghfqUK9B8yEMILmlwiKZPdiDM23QRmTuhXKfepLy6CpaTan0XXr+jjVpAaBjqmg
kz8c/acngByAAxFya/Z6aWRelf3p9s/L+Xuv6di4fkXDd8ZxgjeaiaDDOJHuKa6Ud6ZCpI7T1ppF
zZFLapfKrZoXvbE/ePgkg+nDR6B6Xw0pdPw0BwIno2+GGmdJ+ZRjEJwE+QPUkn4QrdAhDADw24/6
9wdfWr1Q5rdfhYviSQ2ErBuRTj1118OgHWAMdc1BvUAeE1WZmwlyIcH5ot8tc5LBOyRS89HwbYRO
njMK50UjvWbcY7EwxcMUH7KVWmg5GZU8JF5KloJSEM9GH7f21T5rr89UTdSGYg9qFDSnwiD+WSxU
swwWCktqm8mYVRtY9DmMyTkG9lYuFIPWVoVmjtlkAhB/rCeg47Cm0fBplZ7Q6EDes3vgSieuCoOg
8dGt3xRNJKy/UrEx5CD2f47GhCIylib2tclXtbSu40OI+f/NrSfMRVHug6oP9YsOKHd6PO82vzO1
leuG3wg+3lk1/2wnNf+bMgTpws1IY5+cxRWjbg0i5/p+1SmWw9/PiCvEFk8Mxo0EQUli0At5KxHf
SZ/Adzsl51pMAVoq5P7CoiV3+NefaZ5pbiold9vxB4jDAYUmYm5rOyOLjcy1L1vox2HQpS9ZhRpz
++cRcXH04ruQyBcEUQnbvUcQE3d5HZeBD3frBEZU6TWyhX+eALxV9KdAfcXlmXELeU21Dm31Deto
5nMtudlEw8sTEDeBD91uaVWCFVwgOY/mcVg/OrWPoVW3D26lEZOutp3I1nHvECSo+zJ+QnFxf8o8
9hglN0ktm0HxGHHO1oEa6aAnk3mMmAMS3zqDNuGFVYCdGOMb9Mw2M5noxyctnqxQeQkKU5WSuU0o
+x6C4DqDf+qYtNLT6aNDOKkRnCadTeGe1gO7SavihFgyz6Tj7s/rmuUMHvof43noxxKLcuj1DrSe
TE4zNP0FLu6HPfjkzDpjXs1OuNLfVvHUrYSp6sJcTyA25ldb/Fxtnu2aX11FS9sSg9d1iRLiF6uT
N5e3ySHgbxSJAxDCYMXa/5z7ymlQAXnmpqNmvKCBIwknolU5VR9tCXknI0AasuSr0Jrnba37lgja
VXvfO/vK6K4sx4EFG4msZ0BWQa4ZDePal8so22F8fPuqGTQJbFTgRploBiBUysMRkO2sbBSsVul5
BhtftMrs/xi/G5Roseu18wOnqm2D2FPu0ABQ+ag6uPVtKXzjaeNQzhawjGfZp+dmZESYyRZMrdDq
ttNLx8zMlj3tsz3dLwroo0KIXxnTrlz1eqlx0ov7X7jfaM2Yzg+bnUz56y4z3kTNASoELl9lh3h2
Fjo+Z25Bjr7gEtnTgASRozZ9G5GzvI1+F7eKEYs9vRP8IP9Z1nqh9JUzk7oGSVOSMJ4OINEppXyp
49NQoUGgC5UWcpyPgYAjdJGJ+IKqQgtbnSH32SPleBYoeI0Hsz2B2+JbUKN7lSizVwOBB1AB3IXE
uVSMfOB3KqIOSq6+K+ucHGInKW8J0hIBDIGLXwBo5Cs/q2j1vO0A4bxLrkOpN5UzdFlDLsxNGVJL
rgoYpzIv8qQyOep4HGZE3qKg3DfzcvisFC9ou4cUQzijd6J47awoTEhrZZBoHHbqe8PW7q5lFjBL
eCkUv3rRMawT11gxa+DTnXDNiuFFfZWMd5JzBPSOAFApvjojdYI6cX1PLa4bOUsMRv/hGe6pClZS
jPGgE78muFDR6M+lzDp7WyAmVtduDRBospxC+twiRqi4R4oLc8xgne6XvCj3RGfpCT8eGUhK1SBS
k1sZfyh7Wp6J/s8VI+D5Yt8PyZmPlkUHT/1WVjnl6O/iPxWuUnGVpqC4Yo3jibX79PgslCNoV6d+
EaocVzX+9NBzx4fZ1/xhI46SE7i0kRiY5+fq32UnUkZD+Q+mCFUuIeK9pkPZI91UPGIk1+SIoW+T
/oOE38/ANCeZ7foYkyMbwnwQCTkXvkR9+Jb24w9kwyH0iCtUupu1yinly60+1HENkZg0GLfwqxip
wi+z+YBGpvX/2cdHb8pAUfErXcbohQNPUJrpd0RrHaqYGJQySrE9zJtDb9Hq4WNsYUzbO53XC3gL
LG+dbdHaM+D8BxnMUfuvUPBtNeKRmHmh+ypo0uj5+IB0EgDKga2Jkv/I1uXSEkRLDXQOggiZTbz8
/hc1BDEYVTQu/6pmXz73jXJLA5MYUXk345TXnyxLZR4mQExZdlsqEFYId9jjxMyqPalq6GYtP34M
bIiqnRT2xHbzrtQ4IuLqyaKeRZLj96+RWumOz7VAk5e894LJLXK5A1aG8I23OXYoe/qy4Rpi6Jsf
OBjh9Mv8EQ1lJTU5VHTTO/E0XkadNE5/yigfEJzInrASSBymofheMW7QuFwaMuk/NDXkla87ChrY
d0ZBTwxUpb1JmegwbAwENhF/YT/R3aF5ojJ7xxNTq2Khc41FjIzvTAjwSfPcdrmxiKoIiRxszzHn
UedImVPxhbX1GeGRiiIheJLjMatZ2miVQCYzTInG20v4C4u5Gv7uTWujdrkj0bI102Dx3Dg82zbL
9qcGDGRFESTidzU3B+r/4euIv1cCqHoshEe3hsiUNBIT/9PkTfZhX/N3y8CJjuJ7ukSnvHtykLAE
SfWnpdXx1Aotd+wS+U6JUJbADnejTqA2HATfuamAfv3+FF3zp9+YCf/uVi3zo/pLcOGw4HS/1qvr
v+lzYONUnnxnr/210O4ZFlJ2fl2MsuhUGE4oZ4l7QFR3ob3/u0Hosj1C8oe92n9QgbxqlGsg5oRL
kMZExVInwa2Seow8HTCtV4TrCtSh7s2OtctuiQKQhco1O63Jrz+x8f3Og9mHGN/rBztzrcDfETMT
sICVkqywaQUG7akaH7xb2DTf2EsYjQXcQdod2GHIYBlHXUyHVRJVD+5mByhh1sbrQsmEP5NXAc4p
cS7+3o6HXd87B11wwiElEcOj5k2A9TDptMsEaEfNHbFtVzgOdIOfFVR26cpFaQ77AlsH0MmutE2N
Vshp3DAQWwMZZzCYXooHauE+muG7DYfUuVC5MPRTv3rCfiTcCxkAnF8OCA0/5Bl+FuPf6CEfStgE
kfr21lGqQGMgSiSoi/B7ZQqPI6DQEly6lAG7Q7Ou9F51Qshe71Oy3P9TL1Wvv4+RtKtxlFeT3dEd
YuFk3UYIeDo3QH+PXXol665cvO89uyE/g61wyo/p/RGkYdTU/fsFYiNFf/JdFzISTe6FHu8woYQq
goRiaMRwU1XmEP7UNyObfUItrdMOEZExrmmbJa1S7Y1j6UNP3J1QHQOBeh7m/2ybUlyKX33yhSda
39kWqfNajhGt/4beT8JZ4++1jq2Pq8VSQUrLpThoTQSTeYQ8GO3liXc4t2n/RJle4O345/LIlV74
UbIlrf7WyIo/JqUeY7EHSKpjQXgcI4nyVqC0QwSzVMZCjhcbjEuFMDziwKjfZiiITC8M/8goZcNz
BP72vosVQe4H/BKwbmI8+tlXE34KWGAwOI3L2d5PqcslMUw3UWE1QrVnAxsRNdDHB7jyAS+g68ss
yCr8H4TPOL7n7Jw/m3n2JZcnK5YDlwyOH8a9lIDWQI1bVquexHvmSWfWByADk/BMoAchRIm2vnXp
EEmTszEaiftlecmd25/YjDMns8DP6hSuCWLuP+nqZ+r6qXT8l/VjvRJulFfb3R9M8xjt9zUIvwic
4sy7G0KXUNWU3I9pBIvB2K3IU9h+J7RrrDHKKcfVZAxXoFouUs5CFCVZ0yOGTWepVZZJ4Rb74VcP
qx7XfUTvV31B6xvZF219VUiXu2bBn3sOBAKIm9XM3aLFQ8ZKn4Qxv7hYU/OntLxKDJ5i+popaHF8
ksePgXYm/48UJ1d+IPiYNA2cpwAYqEf7JxUH1Xs7fShVw0lYz+9p6/BCn3FWk6QDJdHrTflVuFIP
97AajvRVlGkqqmVgIcAws17XaRcl1VJuZ/5zejT93zz72rErI5Ygv4CXJ4yYdBq9RDiLcwGRBwyo
ljH5PK+We7FcVDSG2LVtCFFWJVCd8z6qrdDD0S9Dk2vtI6qtdg37u9tgNdy46Eab4EV/NA7xSiVs
WxlSzi7nBXK8ixEs/0ezGsO2aN5uB5lkzexnkAW8JKDGrwLbe8WOfB9HjkoLpZI6MnPMqiOGp16g
sseXYTwnUi10EdV7HTaTkFPlLHDBqYUn6d6M8ZOR538Fid1m5SC4XNiW76MFThGdv4iDW3+pxBe9
GRgYcdx3CSnF9sngMbfkIsyOUb2HxTMxIoNICTtJJT2AG3x6DJodv3GmQhrmhK+Hojrc4ZPHhcHq
sxDDIkkKWmUc5hHOqRmRqMlYiHsnetELWH9ejlKra6UqnuqGb3oiZgmEGKo7tjtX5aq0n+106N7x
tWT2++XyjV6GGZDwKfWDxmr6I7z7bht2h+mw1HAU+ainYkrAdqLixgBBODSOtToOQjDjIVbjfVVv
ng8BF3mtCKWA1tahfDZy1XdFiaydr9OaBwhYHTeo27s6PW43jDx5RbZ+M1r9enwatb6OWuQjSIKq
Fo54n+iLJYqrAL/La6vPzJR/5Nxd6WBUTXHyityBZzPForW3cD5XfMpfpkeCrhT3tDVlLQBOk8vQ
lTHdLU7HCv1vhWSHaF64Qv5hRx6aKRwvJ09n6ZbIVQE4TqNSf9Bf14FmYZK3bZkYoFFsIpDh5lrD
j6CXcsznJzdKQeJ9e5zAsrclO2VpEreC1EZHFcYmx9yv4IdZcWJVtPXVuZ62APT6Rx1+EjVNPRYo
62pzRHoHuuFLw3N5Pn4UeTq8/5Vplx/B8lk5w7DNYtvAK/+if/apNzzg9YDDmiDyITYgSKT9tDKB
XAuZ7eeVkSf/jQJyLI0T/P12arvGVn7IW/TZ9t+SjCaSQL4RDQGayHO0I+KWhftTp5GpegH0I+tH
uPNq2toeXIgS3nw5N3b1oaH9MDHga/yv4sDS7MgcIhyUXYMILTHpcAk26AMm4wd6Z+lSihXsbB4I
2q3iQfiPvx4Zx/0bl6LigD0h/QuBQoquRBx1PHc17mS0elhwePr8LKlNwcF0PzoooywhrppzvYlT
JyTjOjhdLl5QEJC6nMBd1kq1IY1zo0J/sQcqBDejO0QcHfcGA4Hjg08IulA5Xc6RHA89vMJOWeUu
IPWN6NtAciEg7S1JHS9uTtRZfgSXkY3qLGcxhoKknIiBefqDOK4A/vTRvdaXD41VVMPFJ5Z+ZKzp
MXLBCOdCcWUkNaYN2D4rBeRYN5lH9cHXOCkPnitvCnGMNTIWuk5DP9gFnAoBPWOJZdpfOeXp1xdt
kVopSlL34YrcrTkZKFbIIXzACq5E+gdFsmO2+LLKyIDwxH+iN9lwickMaXl4JVrSbjx1e6zm+I6i
eXutTGjGEtpJhynS/+VAe6k9W9OI8CvCOtY5czuW6vExDSTX02jpRGBDZ5gwy/ZeYl1+KHQZzoC6
6VsaVBhlhKxPyJRH2yN9ADrRKvh4bO9+p7zx/29qRPAPeMNkuyIhV+a+su85aM6tPW9dQyS+XMAA
sBI3bfcab1yUo3LIeQLmyP2XVhgpM2k/Gr2A87l1eEDwSoHaH0Ln1VUSwL0msYX7B8MyeqdZOU8H
2h6XQ2e3vzrJAEuElrmp5dDRaT/ROHwCm8GEi5RnHnt/Hm3nOWbf9t/KGrP/4enAxKnBsG35er9v
5lIfcyi1bwAPGAINHbVWRafWsm4TaA8Psj473GQKZFY4AhWpV5Hs2gI9wSCnzu7Y4wV9wPwELKts
9k9puy3hKAPW0+15f7OHknpMZ2NZcyTGrY+k4BGIhcm0jR2L2g+0E8me0JN+hsS4iOKQdQl26KTD
PkFoKJjpiUm+fTAWi6kfg/EHjcpPmzrhnedefiFvzl8aBVinLDFnknxgxbGwwbwIMQyCzZDVLjRn
AT8l+insgLIRN9u2bW6Q+Y5/ZPoRLr9otKk8Ww2UL71LMMpvJ93vsU+3m+gTDdAgaqTTgPqn1HEV
6f1puUcim+anFnxjxlW+rBH9SXEGP2bDd0mob/ZgEVsU4DgmWBnwRxJXibyeFNXDgoy0Zj4oQoH2
xNuY2tOsu7U7iGT87eoHIkd9kGKRvkUWAwvjqPGsaY0teyWVQVTHoHJSK+WCrfQ5YJyHD+ZcBNxc
neFZ10Fm2IXgCgAYoWYwo6x07e8GunxLf+R4xAs9o37HGc+yelEzDVfjNIkg4X3NBwBq6lgoe4U5
8jAVLqNsWU7ts4GpFRWj1iCWmpifGTJG3of96HfK2EExSWgHikvD+QWBeZQAaxbqWAqka2IU4jdQ
TOlj8V+xL9j+h73s5VIaMbb++PgzQR0U2mRNl61QLbrF5a4Ny2pSNOSwxBvwiWlA6pXLT36KT4AW
kintZYrTyaKdTQslHpQKU5pnWblFe8cIkiCFmudv7oynqo0c03UOGRjcpuectGgFR6PRKkK3KuzX
qwrOBUpclHneHH2J1tivIEiO6Jlbvog2xbnbvbRq1P7c2FAwiXsUKDCckxz+m+N2yzn5GREfEj+E
1KfTX5EnVx3GRi3VLzKXJSHmMhhVeMzOteXWnsMZCg2u+/2Q/QZPy0t8m7Dxtik8b0yXsnzVedm+
is7jLRbNssZOezGetTda6vPXrTwDac8sgZvudsIAM4yF8vBvjzcrSDxLd5Sda3aFSoingPHRGlJ9
b/CMk2R/WJpjBQKDzWatLp1eJULsHAIPKcu8OfGI+/ax7sUKIcc/2VB9cbUPOu2fRd3WAgMFIgCW
4Ga1AQ9mtn59CKes9eK7ONdbH8z4Env9mVFA/dw8pIQoIHMrdaR9Rbt+0MUtRsGdiuqeZzmIMnHn
XYymPCMtdFSi6UkaRv43MpQKc1Wvv4iDnHFK2PRJ0bdwBtGnE887x/EpMpozIjpfDjAVfN5zEQ2L
usgYBZJdqez3PGFajewvc73oPfrgXW4cpN/5vEGOSr1CtBS/A0/GcpJtQ07Y5OC1rZPKyrXDhr2Y
54sp/JXNOMcb4pQefk6vXxsbyz9e944Vo0esH6fvVijYLTHNX5OoNvWbel+Gc9WJQtRyZN7fHXBk
dDgggIY0dKT04wxg8toxRpchc5VJp57C/1rS5qEGi8B2DCYHW5fqoVtRiUcTDhi03CrLmSgLoeZL
vHmYiMpHORYlQ+l5++ZDO3xcaYPZId7kF9uKstvW2zgKdzGDRRBB9xy7Hu2gOalCHevh6M1sfSpE
BGKqOo1FX/H/xJtRB/aRdz5yC/rP40COt2eRk5UWL182mWzuInOwCkW/YP/GXFIuVtWeLIFadhGm
lVvvnZXzCpYZWPvA0VJ/bQbx/HI+UReUaYX9P6SjFQkgkTwFP1SoPQJM+xymJ+KIrfCqSc/MfIal
6aHBMtM14dmtM4ssKGLkwf0Q1qKR3D/MC28didFpHYol0qWr43eRf+isMhy3NlXCzD2LE8PRG64e
IIRjkpE5AAqLrNcUUZTB9/tIB6VvBW6CrjUOmJ7Dsn81L8RAaCfxT8HboXgqKQjdscKRz3ynSR+I
wZVulNM3Lpvo700NWZ9NLVEDl1Umq+8Isf+wA+7MxjJBiWpk2DlSWsZfl3Ee3MOyRZCvONxx47he
1lT+eHYo5U+KDHJxzD9beXVmpcEeD5pyuc7bSNCmDakxEAwvQIWJ/oBFdF+Gtm6UhUoFV1SEFenf
KMdukSSPDwwwSZkwfmPB3QAKZu8G0Y45gtNnnucc80Ei6gzmb723reyHBHbkVU0sYuipBXQ/6CuU
Hjoyph3dljOvakcpxnNTmKtShUA3jp/abiYZUcoJCnq15RoJE2XHrRzuc7nTetEWMtxqDZ/smYnU
3iJ+nsmD6sEnje8+8JzF+RXfwSdwenA4GV82Usaq/A4DQzfBk7V6rfh8fkZK4o9+i1tQOQrWxDln
mMjqSoBCkwYNAIz8BiIbpVHewz47VjXzQ5szXhWNdg+XKw4JvQ5rJ4R+f/Tl+id+pXPOKU4X2HH2
Z2HaVujZWGurJ5zSlB/ZmbHADgoET0oBQjrGsm/Dg1hgxU/aO07gjPSEmkhpo2MjNz8Ups+H1xsb
B258Ncm5gFXKMn/kyXrwSZsufyRyKlzuGNelZ9zP8/fMfdq2hteSBL10KD/5cSpt7TWBJdzozg0W
L37tsabrQNXT4AjAMtNDHJP15cdqLsPsJDINTcGX1mDHo5HELjIX9A6t6Hu4szNx0ANgAXlcC+91
oMeWrsrGqUSvNKMo3RcyRztFFt+tSaF3+7VoV5v28b+wnJnAUFKtf5HvNOM7q0Hy25gLXRowf1Bw
pGgEbhLcEPYGt3/pEEQDB6pzKBYpuFRPYr6ulXWNbDSoA4zcc9e/j5ZaLckhC+KxOlbiAbLWo8/l
8Z3KkTZjoiXhqDEdf4EY2JgID/QHHV7u+TGKdOvUHatXWUkaPTWS3N9M2YcbzfNvsTnJ4V+gYfx0
ChW9o+FX0xTDGLgp0rOoGB1iDVlGByt3IUIz/37AipQt6oznDiZmE4jRvThRZkQ6ulnXOOq/98yH
UiKsRxZxRdVjLS7/VkEMhrkPasHJOvnajrU64aC3zdQFYjiYWnF6YvmkQqDMpE/c/3K0+v/52MBv
zhc84qcB0h8JMNZSk2aIoIPuhceCZThNYVIrlkHNWcQTfHX5B6lC6faPC4uKV4CbZokoxu7qYcNT
60dgb9HU4MDtTvUAWvOtbykvY7ie73V9K7e4OiY6Rttlk2K/KBzGNEUhX9fi9uQBrH1CJ2iedCdK
aD+JMl1Eu2Xnd/9DbYC+CwikII/Y+zmjIqiCaiuEY1lmAA3tsEj2ee/mcvqews9+DjJJR3hEjP8B
BzBAd/c3Up2Fpl+a8YsZ0uo008TcyVWuVPTQDOrBJ0TzU8TrnzLMHOtHqZhAtMeLuAXQkp1dBP8L
EDatwnZ9eBewdHu4WmewU/ygUpQpgukC5RfbqUEGfccIpI6skSK0dH1qs5/ip3qDKOPnTyYA3wae
9Sld/mSGa+KMNSXSI21CBeGQowGSc8bXcMzDu/IuPymmS/4qnAFNI98I8OCPFfD7+/TNtdA/UNOR
9NkQtu+DxAxQMoWhLDv2WrumKcFtG/8HY6NWnVsZSlAGj4IvD+1Nt1OtUxdDqG67j24HyRj+remd
hsSSz3nppmbBBccl1mDXrRqm8VuCow2mKXdKlBijFEBY3ZzzFeBfOQN80TVqgCxI4qO3n9YGJRs3
8ihu8ljuO3Svc536fLQhHXnXWopBdX1N5BrEAW3zxh3hEOK94Cj5irlP4ANEYD8G9deWoUZWrrZK
g9wCrgmw3zmUOKYPx4x/6KidWIStEKG8y+W1MO95thqWGo63zm3zhFs452hdqeafHtlf7RZ1zy8H
mmTr7dvp8PCe2+V4B71eltWC3ZUgVciYMfOjqfPgqpcqvbYEi3EIPYvZ32p5Kl8f5tdaSqnJJZ+H
wUNsy/HefEohhtaouz+M7Ces/dIX+Dsfcrlqv+MzLcnDpyZQkB2jkzUP5z8+uNAKhPJBjrl4GOi6
gBHht8WMRvxm3rSHUP7x5ZQcMjgPQ5Wwy1FpNq6uRH4QbMizxFLLbSykG3RykPaiQnlrJ29vjfhN
vnFrYQrCij1ewBt0N5rf2ZFrH6XUNcmP9pA/os7Be2CtszQTyYfK9EpbjGhAf6SlffadZ5w9odXd
rC67eH73ZMKfX60XeBFC9KHsTBa9qlNQ36M42WpRgbx9+TlbAAKsNFZj0UmmeW5tCe/V+e2bBbky
CnCvhuTkKi7jXpISCwkEt41C4NaR7+sYB2JKXMWPVxAcgIBistNAKgwOPWC45hYE8CBGyibPu3Pt
i6BDN9t0WueyPUlc/xOsvt/43lc3ZRuGqkD6mEJOYqZS7D8fQnR3eKEdWGsvR7hJvAqBJgdnuwqu
sXTkFLc+WLtt4ghfa31UCLMJzWtH0NsIV2/KJoFSujlzL9DxFvUa1p6TTxJgI2CufdXMDOplkE29
7uubYkafbTcnyUKrqUT6X0SMeBdYDPfFH/Kxqm1/8Ykkz60RviW4Gd+pf7RSRnNmXAPr7EElUyUg
nEbLYUvCHCA1UHqDJvqpFJLgL/P7JDiQmYZIe+HDP3QZyW/YMT0TOEH6/QikBuislauwze5D5ntW
fGmJMgftZVnHsQQ4+GOWZy+H8EROdblJTi2eqlSzrtN/EtMnWJiIJjuJtHvb8cvOjEvSsLk5AvTL
u9wiqsLaAAAv/DPTANwPKu1jtbDX/5hfmDb3Y12FSgWuNogFKy2jVVpCepgZXD4hZ0HGApvY7Czc
Po5qoFYjIQ4DXaAIlaQWk0f3qKljubKq2VR5cpWcmBQVkum5/ZKStBD+NkVaJ3T15DZnZ7F8lywZ
hOIz/pkgc7aQDkb4AyVvJZ+7z5Z75etT8tO3JVovjThcaGvDWedWl/PNL2CvoT4z633jkoI1miYn
KpiuQBUMRd60I1T7A75EIqeT065quVDZ/4YszEI50dysogZXXsc34bVXagdBDhq47SLR4JkyGJ9t
vxu/C0v9Avithha0F5vfwFRRBdVvxtSsz8XdlH6J5igpmb1ikns7dSSuvc49e8YJWbhwuwhu2Nlt
39KpDrDP/k6s93wH77EvIFcqWnsevvte3fphN4qCIOHv/8PHJRIdrC2wn9WJZzaWSnFhPMf18h5i
y/3gsiyjNI+PI6MOZ0RQ0XpqdNOMr4Da3dcufzpwrxGrQJGO3PNZAXd9/xVPupTe31lN+g4DGvJw
EAdLh1kXJqmUBdO+3nvk5+sWNDhx8bL/QPoZWdHrLP2X/2ymYnEeuxnLWI8iF5Y06jTN+9UEm1Bw
JFIKH9nIiEm/hjrMna1u8CaqEqn6Qq76RJjO83vU7eZYJ3Go7OEE+20FA+dhb4lc/M0Ptr+bPIDP
ArW3basdTpZcmt2aZU0vLsOAMq6MOqXq1kS8LLujzhLLVJ9SjyOAhlpkn4dSwfqUN+0XNhOUdWim
Oww3yoI5SQj2HLXfSor2dQ4KPswZkj0cTaqmVeEqrEhlMCwckyCz5+9FtIm0hCx5ZDujtVhYcD2K
xL58AB48NaxeG1y6A7e2cJo74sSQDQF4faCBms6kRH+VeONNKpZdSDDPsMzI5ChT8dIjSktlg/1R
HvukqpdUCZ2YecHgc3wwrVeD+Bqmcf4wM6DhwEMLIuDJp5Plxu4RLO9t1gwphe18HEtn0ThnZfZ7
dHeiX2/Jq6997o1ht2AJUiG0EXV2POn9ULawH2K9+YHtfOMZJobBVQAb1h3jvqTIiJUh9WgQV+o1
aTuyLRaxg2y1ItlUqPH608FSczdcdBFU0KSSCNYv/LL8bJNCpDCxezZgTfoFs3dOLuCzFD+NdNYo
PcRcaX2E4UO49yiJ1Ge6gs3UK/EucDQOzcIBHbR/pLf85kWtu2YMcr3FRjvca0o7X8PJqc/3RYf4
EbWKZNHXhPYY1szmU8bt2TnMcKp96YmM/gxWiJLhE6PLwc/8DJPHmJUiuZeUIR4ivCgPitsjxTR0
UgnNbsf/9uWM9yRtk/rYbLLWlmORs2BoYrHz6ThuaGC2o3+vK7RBEj5LRqy4pL9qMEhZNXeWZViP
ffAUv42RrE6utLvI9VnOEZdpdSzXLMBWTQFKjn7Xiuxs/JKRe7UOZ21kVIH35xo0XrSa+8sgLpBs
aLj9YQcEP73stSGUvoEf38HpPZT//mRWvLcFCNekheAO+qYyzptsswYUxaafqd+a4uPEZFyI6Y1E
jUfaDs9riccSGHylBhjR716QydqsrnZa3SI1ONxu6z3bD9m4ua/+S3cu4TNQEIIz81REKbDonYzW
CUeFikJgeV9D5UJQVGktrBIx6MtB0qLDZ0NzqZ5+tOcksGcQLaIW78SpGUYFOFixWJnEKyZ3tOy/
U54c9hn7EkqsQJSFnqMDCf6r+Ytp3sj/DJ63/tKHlzg8rLERimqwHk36RvKFYP+vzQo2GGRfyQ2K
paYxts6d9MfwWbZcsy586yiPBM53018x5hStqK9ZOtlhg8WNxase+xFhfEoNVAnsC6zWs0KJgo1v
7VYIhbn1g/nfgYgFI71lBFv9qAtLhhTN1DJv8iQBVU2IBWGVaTGq7AizCsef8XaMEo0xOZCirLXk
s9Jh9Z2h6XlmprbwV8GlQatm7zvP2ePZXHugCifRXg2riOmCIE4qUQnJB7GO0NrY3fMz5qMfbkAX
H9+RS6FLVc3mz2rhRxyhzjH90DyudMYWJN2QInfZ2anucwcZyzpcVsKF9kKiJt/vXKn7Ubyl2HOp
l0N2LQuK2HUYEs04tf2Ldrpk1DgIdykw0tm3rkh7jfWuU6tIeZv6sdROTrHzaGfMjtXPdSNgXKX6
gJmLU4r1oLiA1buhG/PI9+Fy9q/XaET7BUljQC4/cf1yD9Ba/yfe2GpE+8CXC3KH4gaY6BHi0UFD
hWu/ow8otCNG8bdKVrE8rxbY3WZPnqoqqZ2xwFkaTDt5XeWvHMslgIYTqvNRE5BVHpPA2W3seohS
g3l3Ti13Hjltixdx4TJOvLK2+y4qOe0KQWc73os18jepFyE1pLUiXvstjE02WLXA2CreBtrZlWQt
BrgSmeRRObufJC9CaR7DKAdH3Q6UlBVK2Ut1x/mGorajKXM3wCdNQjzI367S2ZlV+vvyRHEE9xUM
27XWiG1HhSJIpT8U13qIV5e3WE6x8SCgqFlkSgF3+cDlTtEB+SFsgYge+xqpvBKIm+6TUnxOND/4
iUz7VEmiPPSi9CzIdgnMsESgU9RfQHToy9NW0grxwPb634co54rNjiW1YUogL2otF0UBT7b+WICs
D7fRTmAnN9l3hBTvgfwwJwabdH8XHiCicrQAl1eleDM44uMb0QoO5v1enh1YwucmOzBZ+knwN0yG
d6VTFAmTyvqGulglc5Bn5jggyPsDlUZEdeG/Z3gH7GfWav+NG16IlyN4wR/AOVfe/aeVKb9UpdMg
f64+yd5b9Uxd/J6fwTgd/psou8FeUZGjMAIuTLN97JVZOLhmPMn9pvPfI2iPm8SWx+WWgoWrq5lD
W3ZuA5MgYfIdxcXjvc8MR3MPOL0FDscfMdNVOEB5peEApT+F6cu1KGH2TXZzu8McNmAV7lAtc3kl
dnO4IxAVc8u1f7M+VjMjAt61b6otsYCb2HlZuAcwH8mjFqKIbIQ2+CalSOnhTni38M/uLDu+7oYY
h+F+Cb9v50stxNiU57wgj5+0FzPW1dWZjvDGu9PENmtIekkngZiDRl5vAla1bvD4V69jfoOIXHbp
ZWG/DlZixB3HwoWVx86ZjzveUPdDtrq3/CwdKCW2+b2YohzfVfCToDstqTC0xphTuTb6c2koeyBR
1RySY8DeagfONBvNizKFjg3D3+PW5Y5Am7plm0Is275RdhHbzCn0V80pQprnMfpxfPA4E+jAN3X3
XU9kS/fo5WHRcPvMusRqn7Kg59Zf+ApeWOj27iniFA4tz8xUL7bdkcW19i0Ro9dPhSjLl+v0AFgj
cZl1FVLhs3FmhMXglKO41rFROX/0R1KYvGkqGIvGaB29g89ebA4PTL6w+Lw15i1icGPS6BYqI59G
6A6WYUhjDPvy9ifM/9DI3/0l3p45xjsKyeBggBXcey6d5s1y51/m+KL0RPd8oRx3eB03vt4Y6ad+
SPEkHGTSPkQrnRz38FFYmP04fXNVOXKP0+Or+/KutASfnAFk1pA9uM9YtZ9ZOdFPgWRUNFKdK3tc
M82795yiUFiQYP8nBi2eq14Yn+gBx/ra8KrBwr/+FWyDs9FH8NqiSlnRZXyCagcB8JeK+6sFrngD
hQ1VomEKEWlqN4zmQPbOwAGgsVlqSc4bHscFtpSGNHm98/RFaLXhSytjKQWZmrQ6ppIamSU+Y/0W
eqRKAlFpYDzw981PnrmzPBzTk88bFyOgtXfV4xacBOfDtbTHIkger0skJ9HD/neIOFGtTGbV6wRC
kK5KrnNLTEuMbgs0iT9KbOJIjvgaIwaf3i+PujdEwPnS4Rrz1zj+8VLPlzGnE8G3L1IS/nZNU4KV
LEJiam0wyvbielXh5v5KfSEFtLKcIyXPZ1eEPrb45GYD8qw7FEGgNXOgqpfD3rGT8njsi4rWRRgi
eLUw1PbPTn48QJQY+HGvUZrQC5VEMCR9YJhp/4dRdZOyTmYDhAD9uO2hDP6Tn93wEBk5qde6FZ1A
Jl8wR7xEOh6uTouO5p4jnc1nlk7HnFRGNCT3XQ1tZf0q1VligBAB6rHofTBhnKmcKumljpWPFBQV
SzmTVuceZJymXZxDPzXspOPUQlO1HD+BFrT91ycldsiU0u0otVqDUhsNu8r0LL6CHWrDwmakp7ua
iS96lvfmQd6qMNsXV0x9j9lAeyzRBsAh5ZmN4mVOKBp0QGOeAJJyxUbJGwc1yDzuka0R9hSBEFOk
xD2tuy7pBeJ+Xc7vDuYa+tRnQL40JOntk0FcJrtsQWTA/gvIx7BBgvt1JmsyBFWul4Yg3VDBzv8v
GsHVOP1aKngoQSN+OlIyMSQMSnJOMoa+A9Hw+e9BjslSNwmp6g9T5Eyi8kjwi/nskt+g3D/N9Rbo
GmLIZvVId66Z2u9C0tmleYH955JR21ORMfcDA8+MoWkLDo3IavBs/4coI/he5FbPP8scnu5gAjx6
lvUDwBgcwFeXtPp5EuMoWsOgWtQTacYheuPkr95+hI5fj+QE78oralEkXj/bVq588qrSPQmXD7nN
KPxEv6V4ctWz3185/JSjBuzSCGWF2E1XXnFP6ESrCMAJxD0IHv+yMeIMfmq3A/yt9YAK7/3Q8WCg
MMBOzXvsVuXTVNjZxvRkCHLhDXAUVX/nJyUCGq2ErzlS5hTYQ98RD7TljqqBEr+6GcIfnB98i3WB
twsTu5c7JA127RxMKaQ9gxjGO6Lv/slYl1vL/zKC66Cn7Bgko4/7LyXF6Ir4NvN/pNU1Fxqs0RHq
Dgauc0C/Evvgi72uH/8GC46nw2f0oC2lY4ONWTUOn2VLC8prD3FO62MocVWanX1zW8CpZcyO48h/
gTDLp79REoiE6tybY/zxvig6lr07480tv/lql227vwzUQx2VtLQiLQ9V2RM75kVbh22FPE87ri42
/h9ZPGquOGAR44RvMIKaY0c8yx/WxLWW3gAr1jWkAOpQGs8EwSbCQHFkMbSX/P9oQqs3Tk1twCYl
1bLPgummPJmqb1x0Y63bY3TJ8gWWpuGycOaIny4ak50L3t0+vtl+98lt19E3C9mEDQjjVzKdDYlB
yfqSAP4QlyvrKLI6xN4FSkQaDj96IyeyY3wqneiR9WHKFG9RaeNnSXgD7KddoGdTTEqRm6l7WJ3M
MJWAbJRkdA+Mlt9tkqSVGYEQfVqgfpUvIxFDDx+8Zoby1g1MLu2WP96ByaSd/adYZur9DrsAHcA2
3CtfUZL5XZ3ZuA2F4gW52uLMwTdKgNc7twyAbkZyFniJhLVqC+DEb05SxkZudhhV+7rXGuU3RLHL
ou6QOGYEkXPRyAyKTcnFueUVu6jFvxbxHi36fOA7pdMnTEbTyzDmSaji3QpkaYfv3ucmLB+qJasn
xKYdgzV+HFugS2LQXsg5APj28F6GxET1rFNmrC7653+OfFuc2hCQcdvPPFRCqZEe87c8gwh427vc
MLr5Zhx4p7rJJf2FfY152and5gcowvlnUZVHt0qaTAbf7FbPxGr3mw22EIHBlDcyafpDSN8NbcYe
WWwtWKhLAXrRSi98Nde8IW5kdaQdPhWJF3ZnUKK7UM/EUf9YUPVoO68p6+yw3hbkVO7765NuIAWQ
1nnSo6u6SJ9TsrY/qvWgY+qF8TXF19TdrMJc/6yRN6xPzmZ8JBz8abK+MDcv9C4IG3AFOywPe+OP
IwyY8isvubxZEvDakT+kgGBW8I94fi72yQ9pbhBbozgtPoQXh0DboLJ3/NsIIedsy1xfQ5O6Wptf
FqZucAIHLhVIeqZjcptVBoUSHfMYQX3uLtVm8Sn/nvxImK6AmVXQEyywtJzCGZpGLFqm6SJY7U8H
A7n+j+rZH1mA3d8oKGajcMAFmzE2Yc5M82je2V1u3fPY/0bJqcwXH7+v5gXtVQk1jzIhMdvae1W0
i+/9EEOh/D2sDYVzTqcs0oQZFiulkeTgg3mUvyvudIove9FuuSWgfYCHhl9lUDmHoig3NNyWvdfY
wv6iek2vHScyh5VwDBCUmXJCSAyMn5jMcAoU3vGXb3OhTG23En/DwjPrxCds0fedVTTUfaKIl4S/
av3NvrfqRJZw8Rc6qgQovANQtaqTQGpMBImCXpzrANgvPcdY8VOLvIg4O6DVBOdbrqyHin6Jj5Nu
FWGA410OrK22MhufzKPc6pSnR5WN1MXcVypI63IoYfCwdsX3Brt1qLLujPD4F7YYnRfvsGPEYrIh
ezEfyu1EGKTugEZD8qts46MD2otRi0gWI+GSyNTiPhWnb/vPDHw3jf3btfCIQBHm3A2eOPEYPERW
OrCEgDr0f6mURWaYpfKD31vuyZ1N8yJZKsx+HkwvM24rUuLNiIZM/xcl6DwFJy5rjAylSFChHptr
D0+0pYyz8tcol6iGsBjLEHZAHNxQ+TbkjWKYXi3CuWY8SfaHvL9a/DO2/L060yFnqckZJizMif1X
OZCmT81G+Bv4M3nEmt846H+a6Wqbwbk0nbKRDVKOT8x06cWaq36kk7vB1vK6MQupQRw6kyR1Rb5l
qgV2MMXB3G3EXiqouYi4esuRmmmMlCwf+lji4+vZjoWZYhaf9AxTPSlEnHEEvIbDAtG0KgT1oul8
IfKMSQP5AjHzNuEmImHRjAsL4EJf42VJdntNWXYb+b5a6ZL0uOgU57pCMZ8/1VlXdwzR1ZQ136xb
7aSiS6UZTuAKumfAMpNb7NCcfAJSHaSIVkaS89ZwM+1gC5zh4TJ/AQ80LUYNU8IF8ZIqnwU+Ztyo
Yyp2R2hunKgY0/MSxco4VCMTB4+thYk3RSLOtlf8ID8mnz93nIMVzHJXNwRrzrCStnpK/rDXJfkK
SGphmoERlYMDCZKhVkG8rxj8DjzAf21YgZPXDXGbrfzbJl9aB/HToXMu/xfUEdmrKgl+AErmkK05
miin+f0wZYDrBuyO3MCA24k5867sB7zHGFDd9wLiTfdbTGtGnp7TINPGR7iIZMJmYH6x2FBuCAh3
0OceS6hkiPd178MZiokklucnBPvTjDGDj1V+Ieuzzxzz8Uhc0NQveoOSF6QbBgsjTqtUX6WOO/Ox
uj6hdYHE+qzoOHbSqIcj9lA+b+aY52bGWYyb/FNZs/HNOYFSDFc0TQ5qhXjORg0mZS3viC355Fd7
Vb2YrAOpKRAvD5EgUdanpKKjTRFA1ARPy52gluvHT/CuS58WuzgPC1gbT95aS+3zt+mE4T9f67uf
cJze2e4KAIbFCrEWHHK7TgpNr7726cVKUZyU4HBOxeLdMDwjAHQRKO7pjIFzvm6bvcQ2mlo8dM9i
+XGJCXwiaUAxpX8iuvx3GdlLzGfinGItmCum9m+IYyGeD6GUH5mt4YOBg+mUmSdsfUcQxtCeRlLH
l16Vk4TZDp7Glwv7nfjLDLvzv3HBrsGt10U02cv6G+6WRLen1boSvHwLrSBxBNP+kbUNm0w/Vwx5
snmQdHvmae3wipjFpYI7ROe56CwQbPaRY+qH8ebudZgp45WtKdKPc7MzLt0XAFyG61D382yy0Wd4
2fzQCx/PxfCIxPDNLx5lZwIWxEl+sfXFFKIb76djl9QGVPW6Xj1IxgzNH0/WpLSAXWfgvWcYIXH/
Ex3QBT5WFlx3GwqjCQZcgxY3Hj4EiusPntlwxvocMCUXKB391Ee/E2JZsdTSNCHgd/ndI1Nf3RYG
HgZd9SjW+siuevCvD5TB5936FacmqDoqTHFNc0oAZD+NMtCGwdGnRntNPUXi+ibD8dbgxod12tIi
QfERjsBZs5bRy7HZULpTjoSvIqZbkVbjp7fL6OwVGiKxI3aX7zciG5qkA+yFtLNlzx1a+6QCTDio
fJDErMsOz6oZ9Gp17yXCchsvgrskRXvKAVRZFTtWh085/W8GIsePBYQlPBZchYyuhEUHvDerlg5n
AC+rsNx6Uuy5zRkiAbxA1SKd4rD7zrdRMbGOnGHO1MHbcP6zJdd5fW2fmufSSli4k0qFjeLDGWY2
0gQzWXUCVKv93MpYT8DQKYFChIj/qmkRiZdc/+YAKKeXefuTkdx42UNumdUqVFsf+b+WPPhtCw5U
OCJgVgTkvKqgQBBNaw8MXnnm277TJ3YGDe6AFJ/lgQ0riMcLH7MuOim4ZpMo4asUsVfE93ZQB6jg
C2K9Gg9mAMnJ5rI/l/+clF8O2uqyytzhnkDy0YVAc3ado1RIZFrAXlUMe/nWscxJesRcg5yNv41Y
9UhGZnbWSTYvGyvKenKQ17Magot9aUotszc+8mZQUcklxkZ0X3D8CTCAQvqmRYbqoVQO1lGQz55k
2siAEr9bz5CglvaCgixMNH1N85ljfSI9vZ7GE8Q1vPdQtCIuvW7SqHqpJUWOPSgnlQgZnokGF+HE
MrELtaqQf/5VH1at6UiK3bwQtu7PDBzVZKEY04XIgr8sVXjp9tQmE8MELt/GpK/bXDrtYiiWbdzs
R6l9ZALyiWCCBxgb0tlnTLqrdNZtrvFv/+whmD9VyOo69NHQwc2ZdlY9UWergugnBAZ0Sce1Yu4m
aTzyW73TSzfBpe1VqWDlpNKIEFvMGkKMTZjlB3Gn+hMxLQnnVMrN1BseU+WDw6OCycz4rNl/Xdjy
DJ8K1SKLYY3xiV2jbkSAswKqjuOF9Zt3fL8Ptae/F/YTzY+jz7pkUnEfvIKwKn3fnQVLkpSJdMKr
HC86NbCNA5uW1u/1jc8ka9nXjv4QKwtzxKpu18GzXDGqcVsAQGlKcEpvsUl+3u89gG1ZHCm7jxSk
0lP1KHwSiw08TKhbAKqWfOxa37v+yMeWoSczxGOj9rO+PQhE9tJH30X7IMqV7hmDGlprBMX29/uJ
RgWXrImKhABJ68f/QXq6QTUpR8Fv3k7oJCbfj0SgZp7sVQCaOcwo+CqsmuoDfijqg5IfO31rQrRV
09WfKe8rjnKhx4LndbUVZapQdkntL+ErOwZfnIC2B72Fy/X+6KqoKxrmUtHzNqqp5hme6UCBCvuk
37D7wAtJAhRdQ7OARU1Dy4BTqxYjJOo2PeX7GqJ8LgFgVGm16XzcFWugiTDPIgvtCl39o7wInBaH
5HdtEDWF9zTb7a0O7bb5Ta/Z4YliUyD0uj/yrc/Vq/ePU4Q76oJ8SqhSVjvt+96ZE30NGAV7q4jk
hOBHiEU8sJpwGpQkzZWHhFREc2VRAvxq2RKY5dGpEDiXqRDR1VrGaFV7bQ7USEd/0coCpO9WAD/D
cjkEBuQv+0ZuqK4YKVXZqdVbHIMgg8IyOsKPNWFEMdOnWSX3T2wLWJFApuehCu3/n2cH2Jm7IaT1
4NjLs6FnWPesZ+UEgSYfmD5GYeCP+oByPdARbQYj/kMD+5liW4aVl6UyBCquz4CT41qaHERXb4Il
jvbHQilz8zk5sGlPbPcRT/UjQf2IIFHKXwqC0Ndu+dTW5uzJDPP4GtrDLTTQjAmM2IUdV5mU5BAz
qkxkHx5slbF/SuRYmA5A7aDKsGPNA9LO09t7RGQ+ApqnV8brscE5HFeiJPvhJjiBR8gpArt048YJ
8Djgcx0E/3pKC01WE85Ky05YXNamHRuKuv76TDgN0vgb7fxqssxtrUQErDF/3QF1YSVShWb8u0+7
MU/ay5czIj5oWgvYUCpNCA0jLaHTyEZgwE2x2PWgTnMzUg3JnmGbaTSktmbl8JksOrfrB0RZx94z
GpQFWQjw+9CO/5fTKmShgSSJEKsb21v7kFR2heesLGb9YgZXaVF4KPqQbxpTVLMEHDuyfCoduVe2
mlZ49qy+6Kauo9Zrht2NVt6VIjAdOZGGPIh3XKFzB8+ZdX/mQpSTYyZ2FdLKTkiK98huQ5fT7ESQ
u768gzri4sPncPrl9mdfYzupdSphjZw30SrnrOQ2nnUA7iCsVOOJQMrttEFbEEj45j5Im/n3EeNf
BzmkwNOlh7wJqVZjMhdHa4Vjvin11oQYf7/uCI7epVG/3ZErPsiG9Z1kfx7qLpaJ1rXvzPx0aftv
xWkruXJKDfO75BwOSpyEokR3fmezlGiUyVkdABurAVZKxk+ZCLYXLNBYhtxbTrCMlOiu5XE94YMB
2S0OvkZyzyA2huLjm5u8PoIoK7mD6QO45rtqPj+w4EM2QotncZWm9+atfPTHQDQA64/sXG6jRO5s
H9oFtDZ4/fjShsVR5j5E/d/Xq5100P7CHnMSgLui7qzqXGSiTmlcdWhNmWBIvWVt8qWoOO2rqu8h
cEuL7blF8Xhc+dzHywR1O+DqGMhkEHVJhPETfWpuOG+MYysx83LOmY4Ufgf24SGX2vYIPUxfDYZs
P2mrLPNTcTLRyJKJVk3irHsRWnRcTBPd+v25qGiBrzXTdfeSwZwAdz1dvtnNdGMnKF7Y/UGlNSwM
OYOGv9v+qZLvKQmNrvd7uNWi50IRrJYRNLlf5/1SPgMKjmaiFal1DxqB42JexgxNV7RMGCV0aBOi
1aN0bvYjChmTnOqQSCLgfLFvXGMeDKnJREC0VjbC7b0iQZnASw5Qg2/SHAn146b1OgbEk9IxtGja
PAcJ2cLJ+Z5rWSP40vBIzG57rblu4oMQw1WpycoXqmpmEvYJszZQAt05iXA2oiBkh8XAHDESEGpA
hBTZA8B9feHCAYfx+xNc7Iq4kPuL+urT3i+IEOV95LjOGEoYSU4n2HzMpo2kk3qo9tlxqcgpQ382
RJIzKJKTLG1fIyfawUUr0l+ToydXVEdI/8zWF/0lHLV86u4PvcMTSl5H6jCArcBxlmmuOdVz3qUw
DxPgHuhgKR10Cr/jreMpucqTZdP5aHsBIpQMs5ywaU8FupRnnSYR1/uzm4Z/xy03YX4bFDXG7z80
3qpu9Uaq1nxf1QlpRSqJZ9mTGUWayGp2yi35YP42SqWiUqcTbHvMMPiyAAZpVtGX+5yN1O3O2w8i
3hAw8lbyBPfc0btc+mNQUHLhQ9F6T2KS8NqIcOETF7bi3SMlBX8oWzSE1IUenclolyIvA6wapzIE
ffFpBiwQuQDh0+8Zr6yc6tlEckWFnfnqbNMQWP+b2ZfhsNc3JK5uManXtzuV5GIf0KvHZE9Yrm5X
DV7UxRD6Ap1/jN7Ze9KMxRCfyZSuGwxRQV0OHPZqKGAS9+jY6ekLfbdXItptp5+YV8EQleigO8H9
2RYQAgVmj6NFx2Ox0C4kKGhJM57JZ15h+vyl6f3hEhWqk2xQRon/r9jhjP2z9HiXKaUgVF93TAa4
SGlg1gAfmsVZf/sLD6RHdnY8hrAickoICgNoWVbjvmxOI1MiQDsasFOmmxDMGOaHASHuJOLARKB5
lwgwjiE+ws8PVUdknuHQtsxOUm6d+nhLHGW3N5qtjfVtpyMutKYGtjgA91IVVDuBP4Nqn1pNVY5/
P0Cu6HFAFCBFTzkNErii7a9MjuBHP/0fH+Lkie+Kb61fyOM/HO0yRHq85uN+9LC8TUY9j1NAOxkv
tyL/USyIdvqQ+Tuomo9JzTG4uptyRtglw3GgLjTqACU3aYlP1yiNQVArDoYECp0E1fw71vgXSx9d
tkNxb0sl4IzAPsDmcF11bAdI1OYZilGAWF/y3tLRX+rA2tkpzGA63avTQtTs00XJn4/0WxHaWcWC
Q4lNVpVZQKuO1z7G4+geIOCS6LmVorcbeeI6Dx4lZ/xxHwEfzEoJlZk3AMun98/PIeFdj7YSY3JA
p5Za0/WW/7VVAxwc4hudlEgUX5FkQVSTFtiuTPaSFSG4pEfp/rj6x/nflhS0riojLgQN1IuGWmJm
MOSeXX5w+melm38+i0d9htcnjHHLwT/s+VQsGrOXkZFkerLSzKF1npnXIgwGNeCdHucItdTqOhdq
mGnZYMGNcwq8KEnYMSxJ8//iAZIY41pa9/EZ3T7b2yz1atU/KQqoQDr7aO2YZUNy9LjukW+p8089
c43eN/JZaoqQikVid6ubJrMQOg2pY6i30IktNc7Ok9zHZKikYjXDjreNmQs+/0TtTHOQpfS92jBw
bPmTgNa2PQXFoadLOxnVjrQBLuuEP97jNNLKMs/pX9EEdBCslmZ/zlak8NaCaeEpTE924UZCZqs7
9wkqatFj+0YzNY2ScGeENYdftz6mOtxYnXBTu8snqV/GiDJl2lvlyTOSD3oLRuRNLG3fAwhByA3G
/XVsBT4T1h89cDZC8TZ7cGujpt5Pnc3bG8w14y6seZ6325jvYTh4g8Fx+a1QVodlzLvkk8D3u6Iw
ePFDJfhCDfodh74oGly+gCpyqrivhNJFCT1vIEhOQB3BxZUS+PvVFgXyxzntvLvJfpg21Nsc5Btg
dpv+UHs3A4T2XG7F2dKQBbZ0bOzO0i71P4FoJn9lo65CAqYOsYgF8P2tqkJl3iWj0UhWlS3+TsgE
PG+hQ6so6VofUiBIsjjRfDoyJumsiBBfFZ9S7xROLWfj/4gCZTFVAvL7T2Z3I0ImBMJ0Q4EQejb/
cUtAjEcBTZd+3xdy6zVxwjz6tU+QZ02uk3KkJwVncXiMOTQnab9be/veR17tI+FdcJd7GHtaCY27
dvf0+zm3KWz0+6s4sAhx+brn2k2OGh2mDyY0P7qTOVMxN/xC9LBs1HbH82GjY38wC8mvZ/E7gV5M
XO46hn4nOi+gcGtlDQD23y/CO7+XnMJop+4rbCVj23Vtqi/QN/VJo9fldiLlFGPSbeXNICh+VGC2
kk6PA3EJrsKviF3KFPgSlZvYvQvXMTEk71aEh4ZI+2jqfhJZfbLQ9jQ4/Q9GX2wBdeTKaCZtqbRM
OKEFecnxevn/8+lRi+3w2rXnSeXaTbcReBL27YGNBpX/KiUMyuGn6iiD6EOrV7251oU62iVZzWCI
zrMDPfQ/wjQjUlurXT2bdVaeE9JLa0jrLtHu5c3WQw++wRUD7b5SsqNk0AyIpuinnArgLDbiQ9Sn
qxDw9jsCkJzJFaka+T2/4wrhPFKbVlBiLQUZ6dSbHZF7Dhpt6+9rGV2cC1OuQRSzQJAGQACb2u5G
r37KSammk7taicKaiufM/+/dU8skt9oxIDam72Vw+iyD2+m3yRr0K9fdg0zR/U+hWTdeZzlgxhqZ
glTA2af0GJMxPX27HbTnzI6I49q6k7cEb+vGVAOZPhgD6mjW7Hu8N2ScxcumkDv3/hV1n2JQpwW3
q2WY2a5fnLf+ZFUYmd3mGOxT9JFRBTWGlZQlun7RybH5kjyV+MXEgnhPXDcBXaNyEfQnNGCgVYHA
hkN3Ar1vYWb09Un+k+6kb2PjynhLkmRBe/wYIJ1rAkT6OnOVm4iikFWmoYZ4AltBddZDFHlh9a6r
boN6v+R44UmMhURbFQZcRDGaf0iW4eu2vM8aTdL1RFlsYCYHeIENJ7IWQcH9Fasp2XBgL2kJ3Kv6
2JXb975rFW6iSLTowN0XZF4snuIPc8b59Eb6XKO2rObxC5L2KzCpTeSGQTD8jIhUAYY2X6R0v4WA
e8rrYbbcBpGRVYyF4vmVHpmVkCZkg/foOVQxpa+sbnHTjJLRD5KTqcfI64oQNx9/y1o5t2wNmpYr
JtXinoGvD9uENNmW+WKcBM9eU76GHEIz5Uym4zhaxWsAQpaDYgUNM4QAQRnGLJ0gjfyDZPcQ2bGG
GnbioZ7C/t7mvWOnlVA8UUq50az+8FEM1Gm1tO4xKVoQ5nUI7xPw0nbONaFNo7aCeC4ervrEsZhj
xhwIndTEoNzC0btqtiED/qj6QGvrjV8WQISe0H+D63Cpezh95EE8QXoV8tI22Mqb+ZZHOgpj9d41
i8ZlW2madbfYO+gMu9QkazNqf1Ad89v3LUCiTLwMmTvQ4s5aMWmj/AMRKnntO1uHZvvOPs4q9CEB
E76OldaT0U1AlIxAqI/7vtOsQtxHhj8B8adoVR9podfRBN+BKmjmFcIeuL6e+3soUGKHPUbhwqCg
zSd6HlNVci+I2b8dYlX5BzhlL2Ar6dycymqE6jHM/rci6wK2LllF1lARQdhdoaEENTKLcOAtBHis
0NQphEP6XHwjWBM2Gda1LiwXDlrKWJrSqnTpXLUl+0KgNSoOzfeBBDkazzRmnbRB76LGQDNUN7kl
XOO+YzGEoCJbhvGMXeyx5RdD7U5BeW+7rzw52h07kEyzr7z+LN2wN9fc+lhtGW9QNIb0lbRTsWRx
6d3b5TpQGymtkhAJv0pVw4WzmH0Y8mAVUK8zaztcDsL85Qcy2udIeWMVdwmJL12AtbYIgl/CqsyR
RBxut/mTbkW4IepBtXhlFh010AAK50dYQ748fr2vNi5cEb4s1va5zJkkOE4yBhpnDf+DuRa+C48T
08itvw/jDBw3EoiIreellEhbInYeZgdm1vJbewhPjOS1j/DZ9Dek+G270rUKZI4YwdmpfIMRvWvc
e+3UteF8glURuwDuG2DGDb3R1oWfKT26GmSW0EXt4QTYnp4V98m1NL9jy7EyMSlpZGz+iMO/UXIn
83YzVEtQaPubzGurf3eD6Md4gZfFdl6BYyxdS7WAkza2ByloGzHOkz2w2pUiFvW29Yu/p3z0ZOGk
HeJDtkAzkJiuXMFH811I04xmzL9MvAXjYE4MA3QhpJzn3AgM0xvwekArBgR1SmmaUru3IFvNMxFy
TtaBNhLgS8rJau4aAD08w8uckq4Y9x54SrHJPeXOnVv6QYvfDiQOH08amkNWn+rrXRp8EXf5c4GD
YJETOonhf9yvS/5NzHUUZJmb/IWBxqS5UASDhmjtOWSP74NewbFPuFopn928F4e4pIkOQjKcgywT
CJJOJfEr1taOojKOZPROAMAz+UHKinEMbOgq61YuOhLCijZmGEvlKK4TPlhEMotDRf3DQ6gmBr5F
n2zd+sv+vhRSWHzILtwh2owDsIUss5x+ytIF0MIG+PyWlOpuh10r9jmfIsmM4Nc7zhScITNAW3gz
jZX2H1Wab/OoiZS9wba6uwJwqimUGQEot5dSgWw3aWwTj39UhJv+XrLuIDXm+jPZHfubu74m71oW
xUGdTh9iWxJuPDX4DGTqBQMdmV2X8Kk7OSxT4Z8snmMWZLI+2jepZF4w6EGqHGab9sbCRkClg8mC
7RulVoZQnc3MV5VLqEBFDKjIT3tlISHKTjDxUjpiZesD4cyi/5YQn/CGxmCIgUnGCIFXVwxHLk0y
qxt1/tmvrPZ0Mx2tzWO0elMXJZnP5DAzg8RYM8Ogw7jGBu/52RD1HBgRYjXo5/bRP/2LDCkevj0u
oXFqzZjcah8RBVV8h9VZFcvNncfYBqEchGfRYHrZtUrgW9AkAesR2zgexkOaQLjAGQT/zBx6B2yi
IHO1My0rABsY1/U8rjL1mFoSeIICRfxWEQRRvzLXjfIrMrYKzYpdGBpLv5li/NRNZiKgBQVYdjMH
MioU+bLJ/HDN+7WZqy7V66f8IrfVg2Jr5mXw3bhJM8Xb/i3U5X+iZa6HOoZnBCWxKMCvHZvPmB/u
eUXuhynh3BrrUlAmWXIgcWBjgh7gvtkUlmKpgIJy2rGNxnu93t0RWPaTSap6MZMK/8AcHBGSiRRd
N2MdoxJaxK0rr2998gXi7dl/xuackjPilpI41XTstGLFpPlZl/MDyhxdFtxFLmqmsEtyL4U7XftT
Nl53jX5ewkQxfJSXRinzSaANiO1WILT9jrtwakuQjXGhzbUZ36hZ5pBmXWS3HRrfjvI8nNl34qy9
1vC1LQMzK57X2nQqVfjS0eHQo89gHNOSpiiL1jBBUQ0JSGWswfLKr6S0PONfXCHL/oVbGYmfoYI2
bwJGg87Ovq6pcB1xBMO7z3/rHo7gIfRWPew/gWCeUGI63lxIITr2+A9aH5zohPhUkiCfAovm8Hxc
lswLNF8UD/9/9FuUK4y4ALzHfNfdQ3l0EQxx/S4vn9gugQZ1RrWeVpSjcSarUjbgN/ZJdfNJkGmt
0naQ5nQ5vc26Sqcdb28Azv0ltafhTDMBlEwy6oBHg9rAhhV2Q/7CMcdbbey7PkwzGUO88GntGC+6
BMUJUci/Ub2ZhzfojE3ZoC/RkX9CMgNlUVd8mDVD45QI8VgCt3yDC3ZmT+uqWCWjTCXI9jPV521+
dcDwnmJY74EgjUdirkkODzg7eOEkRax9gfanOju8fQ7DMY2zN4yatzilkMinzFD239niAxoTQAz6
OUPPZsGaztjZqumQ5RF2hL30FETZ/6MWIJzgQ5ghFUmGPKZ6orWj5BE2vBxXZuetDQxouf83wxX2
WAOSepDeBtktfc+XXHAv2LG17AQvrz6kKKKSYE7wETdtJAEhknrF2YLwUkGuVdTDG0eGqmS7j858
scp9phAiQsRfuy8uUY4PqjvvVwy81ifEAuubbqTm/czIVQpO/+EiQb6S2TwM+fZXCCXLwQDtT01A
t2zPuiOsUzbyKtr6a5zr5jobVuVLMru/dsYpbgLm75x74dn+/E12gs6wSgx6oqUXFrEIXt9EG7Rb
z1S3jjlUJCtIJjXCTMxwVTV59vWcU9fY1eNKJXaGOLZw5Nbd0j56bPUn5titAuNp4LwQ2a6zpQRL
vjoyA6giyxiUWWKKYjHok2TVw82CsJXF9IXgFlhAfSDr8jDOcKGh8q7fpksN79w1g8wfyAPb9dln
Mw2dr4NSzpk4y+EAAffDgbfV9I4NW/NMKtbDYbcTKLTbhPQA8ksXN6I1KA7R8BPLgKoYFcSTOXp8
XecuDb6rGRV3hqCH2E0RyxnBVS3aMLpD2HMM2gY5jyKZ/DF7joFz3YTaaNE0V1IRjyc1inl6/N+3
RlRLZiNNxgcWsTQOPFQxD/7QYp/uNhwC27sGTKCSxhD9Z07k8GM+lcjLEHR4SMnhh2081MLPvrzg
/me0/uBk5NeYr1ICMvedC3H2ttxUWiFWTjy59+S5wBM8uwSPZ4rZ6/TRceaQtUexlfJv2wXva7H4
bkwgkWbn/TEjW/laWm0EYktVosBkbgXYkGH33vbpWzaw86w+objRTwLjdZnsNwAlp3VcaT1nO3el
UuU/XI/MkBoPTiIIjjSmAs9k9A/F4ZiCON9GHtXxx3poRIFvQW5JHMNeLdaQodTMYzYQ3wSz1pqM
BIlYV+MBjkeNVRBc/En5g7lXwU6es1lQg7dl4n1wJ8gXpW03oFg/lZazK9aYdhNwW2nHDIl4Rvb5
vsOyV+KuPSPRO00nIcDwsBXqg5omn5BR50d6JfyoNogH+tDulv8AloX/XCGCxKnSmg7d8V91YvSM
iaS+YKIuYWRzI0BKDdN0vP9PxcevFTW1U8ybIVZtmcZUoPV/GUCqg15TY1RD7XzrkbZ+ra3MJRhN
OuL24HxGhihsmcy+HN0WY+6ODa13dNjWHn49vMTo3dL+caqQP2rAR5wS4rJzMB6fwIzyCDn5sGTx
gePzERbM2SmbTvlCoT+Ce5bZqXvd+24w3cxHJAefHJeiCLtfpurCq07vrWBADEJLSdiZzqPPEHCg
2bpGeNX8UxyfCUiw7W8axTLwoZHb++tSvGJCPeVvTOORCKlzSV+oRI01Fmen6M9ICy9F42Lmdr/U
vRjDedVL1ZPVolGBB5kFA55kxprTDsYCfRG7CwR7wkFn8xNVpUjrHFf3bhCKRmJ2ariVQ6FRto0e
J9APyjMOqvAVcAjP97t46EZP4BTVxNwzHoxV0ibYgB2Zx/oK8EAGuBX+IYbo4p6KFQC0pfM9Sain
Y6WXChuEK6lEC7PaXI9gRMiTP9Eru0NerY8BoNp4Iufuc95MPNprwR4mc/9wz/XT50vzi5traxb7
Gck1jdz5UpeBH1miOphrnjFWJyl5wcgf3F2rdeyRnc9hYGA4oBxzkrDa9aZL22RZJndzwq9ss4sU
4q7d4fzk+REYDmVv4MVwoHo8/bybCWdm2VasldXKnbUkNLoVftx1jAP7RThdzJobcxx3G72dTU2s
oGM376mZUpTlb2/8UX/Ag1MBswG9z6VYC28DZ6ds3FtcLp2rfmS3tUHI5Rho0ukI6JVjm15VWKx7
xzLKVOl2dWUn30q0BaoRBwBpgtwCVtE3V+429hGnsfUUYC8c5sfnLmI15jQ/tzuVM6HYBAqeUMzr
ZLvr5fbs4gm6Hz92162m2QolSepibN/KvLQ1ZRqqCdBzvfsxDlwZDVMHNUCUeUcwPIuYhDlYwDij
r7CWSMiaFb5HLTkdVn92F2MTpGQtRVyAydpkKxshpCi652Bd/LNu4vrb2K5eoTREivfAL3C5OAsj
6vSuvLD/G9sQF5qpxoUfvgLtnZRRb9eXQ34ib14ooKb0A46vstpbOYZc9zGV5NZBABjYUSwYVmyQ
2Jb8xBauXPDDh4QpHDsB5WUx8LBo4EBEHf/ydGuNk2ja0dxvF7YJin3QD62BNRhBPSJpTDx88Ll9
BJhS/Z60aptlXw3iUC1XoIkpIRe5c+hCoDOpN5m2hY8+fsdJTMj1MmaPO3O3FnVMueh4FZPt1O1M
S+WxXMqHMeVCI8vSKHiY7Qwh61up/3NCNCn0zL54c648xBhT0+zrjF0ACtFZQDcZcKEDC9CN3vAS
FvxwDYJLmVjxHrQhKs0vc39LtPY2N2HAiT4KAOAXFAI4/FJP0U17jtYh2uwXbPUp2rCQpGzRa+Y+
g9GcrK9Vu4lkdpcqKGXmlYu9EFBSbFLVi/os9f72uAmO2InMlOUbAFxkbNHvQZKPm1OPT2dGvBoy
J44MjLlzTYaeZw2yrZo7T0Nwk2vBIBdhiEjBuRR3rv9XyyHQ6ftI/9iJh9cA5fqis3rHdQ0cHyRq
wxXOvayl/QCE36Nhts529doOixf/Q+nyLi+J/MQHM7qndqI3Y6w4FVrYC1twIlrP12KXI0RPp3Pa
NP5jJsllMGApLID9gkbFdyyE5pcM4hmWDB66vqFO9vPz0d/jw26SauUNsmGJLKXBznk+pXSM0Szh
dOytSYV0GV5KPZDuggXkEaxwZQLYHjdQhOp/OXVMbjCiVnRR9SijX5ODIMOSPBd96IDJm1lxVxld
BIJZax6TjiuCx/MVv0gPxUmUSE43lyqcMQxjEpC/huvix0HWde/HXQqFifAccJaiqOqUaHuFVd0f
ARGGlBbpMpqAOvPKAEhUZrSb5/mtbLvF/gr4A/n0YtP7i1ajrqshQ4Bolu8py/AdZ6SzOhXQHB52
K8GhSv9u6sWkJk8XjQaCahJrZcyFqz7/TM+ahm46zSfoCv43G9UeRRaksPs34fbbr4+9RI6tj5iH
zHTcs5AFAFY30fqc6u6+j/sn21QIrBG4b5XH1/S5iltvIY2JrIKu/tmY/6yelCW0VX0blo86sQ6m
J1H28GA33exIfN7/QKWAifVducUC7ruw6qk/V6xuENjqR7io6FwxUVHEGAMNUjZoBcNula0I3g66
c/l4cZUp0HD2EapsowaeypJmjhLGeVjX6HGLawrKFLiizX1zhIjRpaANkDhvYkIZ7801xAN4gJlW
LSEJx3nAS7yt1ZsmSQWyXVqW1Mf7oOxUdDnhDh9ccmNf5aOp4TvMF81hZ3NS0M1CqRfkPN6ZwXa6
VW2aBTxcO0+VDgdbB+Z+RF0jk1REjXfvIV2SBUpA4WKCwfj1c9iV3Gw/QEp4NwdB5aSdGjqR2fYN
FqKcgVcBz+rxUBZHzuesVGB7wzPdcxtQPKukZvOVE98c4/0y/6Y44vIXOggTc4ESUxi3iBeDYhrd
bg5vE6Bmp5fjKEqKUio58hj2uRcsEdgcVQFiZU9ec57hmGo20brQIaeYs4FDj8HjGKNxO2+JZDbZ
Xp74pThBMzcE/YuBeaXPM3loXZdf5qfcfVyYnIC/dTJAhF9HMU4ptLquMgDfl8bfF5cTCoJSPY4M
yI8KVIMkabonux32PljeHu8DyJn7D+VtuikI51eAA992CoBPBEY6aBsDLIfiA3h3uf3h2RTWTaLJ
NCGsTfLjzcvW33h11/fhNM7i1FzY15tD7LIYT67tSdnI9dlQs1X2UFYYMgaTwJwECCHctyBh2rjJ
2RxBHPFBN/7hfwM0Qxp56Epa6u21M7bfac3W2w+lWVV8M82LQnM3x1j4QzdySY+B+yj7iAkciUE/
/Uyr6fw7bTJwKnb63FjW7opYsgP082jO+cIbqEDYg7Z0wd0t3edJvE1DQ29iqAF7LSxYs/XEjDP4
NxoxWqUK33s+gqJ7Tlwuxs7kDGHl0BTeForewSHWUwPcy+hY15xXnLg1JyI6bP5j9NhFdNeg3ddZ
9rQC77+I1shMFsuw2bqfC1Og25dx8iWXYG/27p/DKTN/kkHKjmRMHaWnAmjG7QA9K1u16xUEFMcj
+pQDsHef+/zZjyPlsBN1lFmffkXfxdCkgwzAl6PJBfk0c1r6MUDzpEopkDNFQ0xH1hudRvsvhumL
817Zg8QSudBJgVyBipQXdz5ZwDKn4fkPXlz4/a7C3FtkkbT754/sPl2mgDdcIeMhiZUTdwHosCua
7YTFrTU+9oAXqAr4l+kCM5Tn3pKZzKXRxrrgQQqsv3zDIHZaWaoDdk3JRzfzj9mQWE/NhIQzMAfG
QV/k/0frFcexjMsC6yr375vvSGrRwg6JFCBPCzl50KUaiCglLCo5w4E3kluexR+f/rsSYD64qRhX
yFEahSS6E/O31e7UzF7MIAJVsAr4f1MXoAHqqqnse347Xl3I6sWHxvFiHABWo+f2fqyKuBNb8XyG
TdATKqRcaoW13S3yUyA1/7b3cOXKVGK8L1qH6vyelXwCO+PmwqL5o11Lzt37dhskgwk8O5QJJCjw
QJNYUTi5TzlpFk19MFt3nQadYFObCK0OfP6zxffS9JvXN3hOaE8WBopMtjrsIefZqAoDASxam+iW
5MhUXUO49dc5Gi/vA/vKdliVtKrTQyzRz5Lgy+KmdR7cXz3d/qzqxqd9/HQrdNc2v+PavVUS45GK
GykzxtC3wBl35v7pHeaa8elGKaQBItR1nY14N2C935/yhIEVkSyWri3qiLctdsSkB7gsFlbO5WDb
MQCZM1qxhIUVxVzlWgHt2As8IYADiPqc8ffd2JIOxg/S3LH7kvIl7hB6hIYyVeVju4gJ2J3Cnlv4
6Pd8Y/2edo82VgAYqY9zNOiT5hvvhWycd6zRkfyzKntRpGehptegBGf/UueTjAPVUSzjEcPQlt7J
Y4EHW6ZF3p4CGVtXWzQGJCDHJYy8fQs2iem4QQGOhDcDMrnu0G0sCDm3pF6McCAPmgwRAXe6h716
mHUOO3Pe3RdKcdVOZonFSKBg7vzasJ5K0qYZO0WEqPYMrMnB8qLBHrrXFOieb6hpE5noQBRCuF8e
q49ENnk8r4TxN2i6jNkXkKE9LbAfil91WkHOKYuhhWy+VMBKWXNomxq+Nq0Q64m7Tc+Q+sWSbJBv
5nmMkb522qyM3MPRizgw4zZdmjnGPP0Kzs+h3LACVTHH+q0SArsn9AF1tgHESapPpc0AVdyGGGWE
oSwRfBO/l2aeZPzCQAwtL5CXbzreoYabqwv+tQNK6RLUPq8r5JJ+JKfHWce6oEOKRoSpMV3ThkAt
mhYN65b0oJc5rKKfis0ofrrr5vOPNEVIHedH0d73ujo/axrIAI8WM7mgId6RFw+ulaDW5t5di/2t
NmOGFgmU+VteSNVrrK7QiPKZdILAZuCtmL9Y5Rq1QNrGPXO8KTK4626D6O3pyjfLqmdluvCl/8zP
q8y20UCO1dmg94FowkqOEVav6psVC9CAX8A8OdkD0qxcxY2dS4MnjkFUN5M64REKcsnDbCAyxIS6
l0hsneZDVK3cZ2R3AY+IqBbjcrmJc7Ull1ayEavumkoW3erLGfPyaLlcwONzShW8pwLsq0vtyqDa
zN8tzeDv6ClCvrydDfRQxPSBtCJ6yRvGuYDLbFA1FbQypejsrCrUd0SoKGlWojESaWUkZJtWxsbY
ODTInYDLVxc6kz5FdcgKQRPPDFWWJCisbX7/aPZQ6ZfzTJWrSTdUXRiAMT+FZWqYEMa8D2Xj2VZC
LJ3nbXIEU+cQG57c+UPxLMZeNKBUVe/A9Q0o0KS1vClVt/i+68TiXoBpAZmVqbmdc+0baj0uFYnJ
cPAT81uSdruu5C4ar3fHyAPc2h7HUcys1zOp6p1ZxRArgSxscwM0Ob0yleax28F8KpTWxT4RGdD3
P55qLEue7Mv7Jz7q6e+LKCw92qfuf7biQKDMUDb/ujRn2OAAuRJH5P02CyIh24mBBL2F4yTiVGru
/p2E4F5q69bJJbvbplmxWz31cFoTzdeZsjV6yDh/ZJ4wxf6IWiyQAT827RyPu+g7npkqE/fHZa7a
GkElntsIqlzZ3kOAaRSYgjCcLXVwh+x4hfFAN0ms7uvQJHb5jf6yXNx1/YyvWHiIE+mMxR4oK2Wf
uC7/Wf0bsmGaAvF1Ewo8BHQsIM96qs/ulZhFzZZMAV2k6v966GNqlsibnjEd4KA/Cv89jjbyRi6j
y+3JFchkTfjT6SZxNd4j5SMs0MzwE0XqUMRmKm8MlHJQ3lsdfBKHpA55w9e4q93k9Sq20+q4zhka
bK2PC+LjuJTrCFOYCBOe/XspoDNWbn5Trrj9s9Bcra5uGwBvnffmwz3mr819qSkM1E78NiNVa3Rj
LaOJ1rJkX5k+Dcp6IPSitY49LIuzgF8DUEznyJm67pn3X88X7+6k1MPMeUvo9yC7Gqh1CZ8WKpt3
0inWp0J98layvFuToa5q9yxeMidCbQ/0gyj87BqNH6BwLURPBfQa4VK4OZA2mZKZ0k62TmVDPrv3
FOz9y29ddKdR/H57sfQHS39fktjJt4YLod6yS6VTEJEWMDoK+V7Dt2Puw8KwvtbahVd6EZx9pMm3
Lo/8quyP53GGCmSlR4MvGclEUDVlg6vgbSgpJfwBcOnzOXoJbOBTaP3qDcxR5jhrCUKZYpwNDrVw
Etfj6kALT6GE00iu/Pvy7VqDcsFHrLFR3oq/cfL7/phppOxmYxhVIGqn81C/adOlvCY0yaIXP/tb
79jd8GoMpHwcNH08bPqMOM47HCeYGj+BZkh/givluD6bRKr850A5dHlFrH1rFCHsul40dU3SVTEX
yer9Qsng3b3b+/8/a3vxcGCpGt5LRv4DAadfYwe8Uv753hdtS2RLApux2YXw29xTvIMHqGDn1vxV
J+uS9CG4s5DWK0PpgJgmkmm4q7Rn5T5H/ZrM/lcSpga17ayS4U9I7LtKRVGyxGALg2xQ5+WTZGTA
lMH8vJPwJU2ufud5AfdV3qDRXaS0hUzNbE7TTgp0MljrfXNdNM99DaYlh2A87gVPfql8KpHEzI6U
+te7QgJElZjfhL0CtY6JAytMyEpZEsVO1Jo1i2BHDJ4TajcGt57XrvoEAAYldb7af+dm2ZZybYrM
bkYcej4zLyQDM8v2gDtG2in9PSpL3NixPbNX44C4Bi4UZQqYZRKLTtL1HJUWtr3Wn5WTVtdU6Kir
boZL9li96E3YufKAct18Lf1zcwOCnjg7pEJskCn/hpB5Bf+xMbq2k794JgAQLz4f6abq3L4ldgyl
iYJZeiqYb2HrV3Ln88Et6IYBP3B+OPF6cpSAdOyfzyGxs5oNxe/91Jqxhq5ADugA5qi04v0gWIgx
jz76pPZZW8XjpGsY11nsNHxQaVY1GfRQOEyN23yWSMEXIn/CiYsVSzT0Zwfr9YrnLY+sEVmj+6gB
W8WX3prM0mgF7hQ1Wz9K1/V9QfgwNw2aqbOQ8pL6tMDewHpSPMLVbzhYN4DuKPYgKsiN7VAKTR0w
T6XjY/mAf5Oivi1zuYBRilueYn/roSzlueSt5/gG9rBt1AdbqaUWQO52uIYr5HnW7gIyAxTle8Vq
b/FG3jHACr92cgdhHRjjBtTV609b8oSfv/524OhydhsdoVSn7zRxwSFIccDbozh10Dpl5G+c+iDY
JlP+XVfdW8ADh/xP/lfWnrKEO21ao/FBSQ7pPka63KII4Mai9CT3PTOF1ynZGS7+CUUO8GVq97+c
6/k+iImfvEoo/AtjMkeB9BtzODddbftNM+Hr1R4HrsIa0uj3S3cUkcjsB7+JFtnT2SGPM/FEdyLm
Iw2klTu/tH+ITaiZ7gDQN9lxBAQ3RjEihJNYUlT+D/seMga5Sk1rV+ceMgL+bVWYf/iqYxaUs/cW
wnyTevFmhnXm2IkiEQjbgKPmwmqZSxJaG/LQN04LH6ApWiFJaur4cC5WJM+YRDO0/yxPlLMS7zzQ
aI/vsduMZhFdidbXl6NgOShzIXQtBPdfl/Cm9A4fxDty8f/gau2UhTS9GbT2BhaNjN6ULgW831c9
/wOKjU0jioV9uRSrz2AThAkd2/DwnwOrrDL2DxQYToISgVr+0tFTjT5sScfx71C4TIA3gCATl7Ss
6OdhDgGH1PIVvezYjd6gGFCJX1i/sumLHebEnLG19rn/vQlmgBXj5Xwd4HevcFPPNp5ldOh4lKWf
axV63H3RxekIXNza6rjw27TKWTFu8s4E1KVB1gpXBBqhSFbrH/3No420zgyEl1Nlb1CV3Tcvq2NH
m/aXVtsOONwUoFlVNYvyCl+CCHYMbGsqRZl+gN/zXg2YFT5ssYs5Wq7FlS87qz0HcI0sklOATeBA
Op4tJCv1SqWI7HD3NSdu1sjttpAhYk172iouy6Huqk6VfbRVJMX+RdChnjn3hCz8Yr0eB9sCiYhF
+HZIcbk9kM4s+0tNpGtnhbvGUoByvz/S+xotNMrhrvTqxEV3IUoXZGd075tGfQGxXNfV/uth7otj
Z9KXwiPx+GMl+s4NMquzNIR+z3OCd8DCfao6Kf67dxpLM9+eN00UmTJN8oPFxb3wtFPcx4q1fIlu
hL5d7SlZE+ub/YV48hm8eVWGgJ+e67ayWWMizP0mJvnPAfF+OtPnO1kHZPOBDewa2qmxipmfIogt
V6k2m2P+ZFYduKRe4IW0VICyBCkeNAfm5A9OZmDJ7hNjsE1H2MPW32mMMNkhKR1mS52f8CYP/Fc8
H26KYcrbF8KyaGBb3Iq/hvkCRZqWYspCffz3NTOpAV327EDgwH2ju9VeD+oHYm2rTlaU6keyt3Vg
ecPUtDN+xzbmbjCFgzXWLpl4D6SEUgRPJHrg9KUCUk+MQSpAoEAWmNpnVooiIq36kUM5gCveqjeU
8Odf8mfgbB6cWC77dhGvM+Ygn+WLkdJ7iLzmQCIAtcXBEF9ZRatVA5I68A+srz69Nfu/lZns21Im
26oY6IejsHrZTye+yjdU50fx8GhBslUm/eoNxaitsddmxUXZV9B7df0UuFzSyB7AY+RnA5mrjvJW
L6Z5n9SbG8fB4IEbONbUazqpt6iF1TdhULMT21Q5gGSb+z36Ido3akRa59qXv7ZicDRGSZ7tYXOh
Zzw7mp/K5HTITdiCuLAWR1Yep4SYRKlZdCjTB2yYSCZOckwcj9EPaJZ+TaOt5vcKSWJVEDyqWona
OT3XCO3Rx4fN1wYeR8DieOvdwrZyel3C1zUhJTkbqjM+Fp5UoKkgk5ycg28bWKaDy3mF4mJV3AUV
lorLnA70RoVVxevzMQbyRhCl9yxIS+vbpQj86Dh2Xfglv/4Ht3A19eYyALbOGTJTkUhb3v0k8WDe
NZTihM9caRvnt4Q0ho24mKy6nfwxOV4eJ6vZB9gYUMvuvnzJvVqtiIfbSMZjZH7nziz7iVvYkm8B
XphWHoLlmwVeklg1/+JLKG/qaPgq7kkLL1Znm+lvejh7KbXpPKDEIulju2toU3i60KZaCVoZmv3S
ch0mNUpSuosm5SQN/xmkRm9nSkBQ/Wv3qoJIiu97hVdceAOg1dURgfgkBQHzhOn+vKWTxb3mHRn0
QhoXQqtY6zzb5l2/JIgJ6Y1EUpIvF9QgVtBWp7H/YqjpKKa4SyrCti0fbbUOWu1UWuDU6B6huWHy
kRBX1qig1VQWgC1eASFGov3+K7a89yaN6ekQNMFKdAkcg2xw/mlVz11xaaSDa34PKCDLvVYLmBQR
v5xLnmE2zSu42XR4OVR3rDkASADKNFzYev3xWOMS3EAmQsWSBqOXNTDIwVEQkGZSTyAWhbA3gaFE
dYQLCb0/NhZ6TpgTAXtOq3/c7yFmkKcKouWU4o/w/xQ8IKSZL9ZFPOcl+wChpQGyyNz/sFSZyxjq
bC/ZaUVAuWrtqID6AXaH3lYrDcdvNIQpfTleMG5n4ce8pNbhAlXQgMrOEK2vuKXyfc2jtaVbAzkq
yl3GhUhNhH5TfVhxfkaX3t9T1FaQspf4NKsgj1BgVIoyZtVUqXyp/ty8/SU6WAh3tbQScXUi7mGL
fxvBj/PmKQlwogFJGIPqLYf4LCulAHKnyOphKBg5MJNtZf1/Rg2upgYTMNF6Qo5dLmLxaQsnbXAM
gO1tBPIWup85GoO6/a542VzVC8LEafMbu/qmOyOlMkmWTw9+TabZU8SJqyTctWzLiHgolnapilqK
+wRez7UW5Khr0Lz92AN48CMgnEJPki8cmmQe8BYeN6QsL87eI5CR4T34qiSG82CuTgYxfOwMG/S5
xY74n9lKrGteXj/KaoAv35Z77G6zr2ZUyDLjdWBIMenVFrs9YF3TRBjvqctI/0ybN2bQtstG3+XH
wszsXuf8SiBJovgXk6adwEF1FyPOIpJU2OJg6Z21FUBTnOZUUY/HPyWZSLnJIv6NndDc7Z6zgZiY
axag2rSZXgd+Jsoa/A7NaGLBqR0nWvJUC4zRzcU8WntqriMhUKi8RzvVkxFralXzoY7M7FnnWiBy
mMeEACSXwUKJvG9Trd56LLMjLsFQNyU087wWVosTR13bUaKJ1Vc6kdyT9IbJudFah7r2y4r73IuG
3Wt2qLQW7hpYCFwiStfcLJo8JR8QMLkRLWK54OemL2wVHP8KM9KblP/in+gNNySJOrH+5w4ycHva
+HJURZi4gb7I/CiALapXeRjtkOzF0hr07jD2yGV0NAHSB3CybZC0miMAZR91AN5hAVewDNZMscrJ
opmFAQNhvswIb5l7lhuYa9L4usa2bEbU4v6njq/ZIowv/I2ub86Swsk3V3otKfo3feMxBLxY2MkC
jZ5vdI9uO+I6ZKMEeEJxcE/0eX1VoSqkkILyAwaSV0c2ZS7pPzOF0LT2tpzef+Hwc+tivRVy0uCj
ssan3iLu8HSrR7uxYiwx9dXO05vddsCdRMRbPx3bLyqJ2ox/s6tNWfwvSeehtq7TBRHuaASNhkEp
V9FelNwZdHO9V2tl8c/19QbttdTQ7N6ZB6gAlCgTXuV+0MAAnwAr0B37ZYwjzNGFSPagfiSJz5RJ
tzZxiog6k1h+Kq79YqF5J8AoDvdTesv/ceIiYLgr9hVLzDIhRINo9hBuro+v1PrB9cGDrM+aAHma
fH7Ny3mQWYHktrw4JdUbVSDA6yS+fjdEd/taIzuSUMLasu8SdCWJa4Il1PmQKIOZszH9JXTvAwBt
xVb74sKYhl13JkMi6yu5/V0RkM65YBF1E0woWMIjv38kTCEiES5u17/wVotVFjlwCXViIu0/cFMp
Nlk8tYDI06228NxYlbIVsoI8rs3q5B3n5R+b7+uzCAHhONBVZmHdsXHbplnxO2TlPizhKe3ncf8X
ViEwUZBu4qm/jFxnEpBCMR86XjJUKuVxyzRsS7d/tvRFkoHung+enK20CFE8TitalrB+n0oS7YcN
BpOJ5scyvxRDSYu/ZHwA3/pd0Ycp3QqmUTV/aQuAFFGm67eTlO+wklqgE7TGHKqR0BDqfTR9a1NW
iTveU8QAfHD8muejhqOKgwIx3OzYG7VX0fLFsLLzVDnYigaJmn27EzcU5MqScR4r1Z4QAXqCyMUd
CR9SplZZvzybf1H9ho/jlrDCWRl4X5aEeqrTo1PeJP7Z+RbT8TS2VMmEb/YRzG+ZDY/IRtk6EhQY
7oCJ3gbM5Llb5x8jfdV7HCjNbJRvv8By5sRO5OCrklTAO7+0FWfzldIb+1QqvgF44RC0mD6uFDfP
w9yBZYxmEOzJc9Lr8gV5qIdreSkkGbihO3KBvtplXux5sIErV39qnfcyF+84w2+kTdPqLMlGWRUG
dso01vC27qJD/pZBSA+DIaLATfwJ2/A+KSZa2Nq9SOhYiahea4vmvxqjsJfVZ7MbBEvjCpJtrIZ7
MD/yvs/vSg1rO335YYWJUYew7E9ZntOgMjArpg3c8mNSOOlQkWmJGlWpCDwz1rDdIizG5q22KXOd
i+VnUjhws2FlG3MX1LnLrYzd6oyM6FLVEC1sO+Re0CvjWn3C2eTTozMp9AerFlgUrz98B+nVitv9
mcRuS5zAmffbSRkntAtYEqNbUp8uvGYgfX8QK6KMlp81C6K5D0DE/lw92C/2/bmuYUXPLQYoluYv
W2gijVBAhFGfajcfxWIENJqgAwUbyYP6yytqZy7AhyyGaKRtzBz4Ep7UbjWw6Skw5iV4X62jNwgn
SZ6jhUp0iRsWVG1XtEjIVfkAPfpR09k6H3lS+4Wx/OtxNXk3LVXnkRL9O4eEgFoMGuyBQ7mOA1TW
Odnalpm633gyVASz+dvK/Q3dGN9uplf5Y/Y9F4XdtzC1VjWEekDpp/y/yl6YatAGLxaoFMhco9rN
IhBrq6Shgy+2Py9WkT0ozN1VepV182M94nMcYUVhYqXOqLevlFuvUeYH+F6PXFbQxwye9CggbO5+
Z8/HIhz1a6UQISd39qUip3IiQjFpKJ4DIKOqJIuq2j9CbYTPO6r2YAaxZ1oS8tvl+ZiuPew88KRJ
a32xJ4aEloCfQwByooKstBWFYoch1xqr4J0wH/xoBnFlRgti86egHG3Iuotc5ySvlEgsw4nB+xr6
oRfMh093Orm50ackrnvJORLAHdpztwgc+VlRUhowKYBN4oWnbAdeOHGs3vd9NdsxUphsRpAmBY/S
34WFy3W4PMDbMG+GYlIzquFCUgHD+6T9dVIBqid6SUf/E1BqjHkHisVDp4te0i0Cb92HKRjzbWjg
lPYHfIbdoW5RC+2ASwbfYgBcyTXFVQXZCqqE0avb6I/jFeSYPx51tVtlR65mn3rVxeDYPFUkAc5X
Bm1i8dXGMx4wjQJnJljrxAAvYl3N+Zsxkw4OK5s4PQGYoEh4Td5jjbPjVZ7sroF+e8xRONu8aeTm
WuyhC5L7kS8FTQ6XgbrFCT0cHO71zrlnYLcdhmfFuIkmvb3lsnuoct6YyIS0lnp9BLglwgCsSVyb
62FKlQbLLtm/f5CnbJwoKkbQbw1oFoDFvRZ9Gec7RRPgnBrBVVo5riYB9lwqFdZYmTCQ7tlC9eZN
etFfLpMarRDzh1lJGX55kBRIlOJH4lMqFWZJoSlOLy6FaNatnV860OpkhuzbSquYibw2vBcnvb3K
+E6Gp8P0utSsK8zq/Z7SsDnxRa+cLkSf5O3jV8XYNZyYxNpSjdUd16xxdb7/Kwykb9FSoF2tm/H8
aSoIPmZ1UexS6u0hcG3qsYht+pogC0FilDvKdobMyTlNSIm3KGdcyFQO48+dXgGG7GMgdc70tvXD
VGnBHt6wpREvmGSpvXUJU9+z1UzkrVNbuhJzDgUh7wOQgdFiVquRkTC3W1qf/DcFANhRyBo9maT3
dBdBFNNJvdhU7x2ogGDEGZ6uVp6pNyHiaj12ezY0IYZ1d/vBR/UIqOuoAGzQ9CX+h1qbvymoY8Mh
/r+YKxz3Igo600Rl/4P17Cq2PzYJ0CilT4Bbloa+s1YGOJnWyxPirpp6dW5/P/g2+4WZGxlXfoH3
RQUEcb56T7r0pq07y2dVIRgMe7BWtQBWbjM8fQrQ+dHO0NunNWJhRMAMRiD+5Jj7Rsp8FdIKGRga
v5KQ3CH7BMUbhV8BvcgYDaYByJP8K22XbqSoPxru0US8R7tqV8SqApGI3U0bbxu/94EFxHjy6O79
NkcL7IKYzZbpnBB3lbrH0n7k/NYRdgsqOrgeROK+6aLePArQWk2wJxYEKhiJbDe6UcCgBpo2fMOO
xoiTcSd8ZsfVo8ogiF+D/umdbkdRwrs2SRY12vXptCnKKUefGtc5uK7pA8+KxN6/xw4zVM09iIWV
2SJDrR8cMcl7XyNVp5xxc4Clur46p2gj62O968GYeJc3o7C+n1EzKDnyCFaTX5yiuD51dRMYxcnf
d1/C+kn9pbXf8l69p5cXSW3CJWnwB2eJo6WU/U/7cngyFUBGDMvp+tevdDriA7z16cEZyYwthmvb
7OGO65kfZSz8d0TVXLoiSSXc+2YvZcMQsd3jKQ0iGIGRngHVZpv7yiP45sN3qys2/V6G8awPj3HV
OxmXmn/rQ4URszmSF8wVM7gsPry7vGNFOiGlXVEgTNaZ8+F2FqTq8tW2D/9R1v+TIKKb3W9fiIQm
F58V5qUO+Yu1nBM6d4/gINeUmF0oawAVtfvI+rW6WToVK7cBuNeW6O0L1CFkjNEyL9fvRHvXZCy+
A1sIN8Df67vc9hCD5Hy/xdl+ky2DLdc5HW3/IOvC3GJadVqILSBmvZRN5nuc2On+ojFjH+GdOm8/
K/ApyuF89dRtCeWDtZNUUnX1Q18umePbUCPIbttBaF/sME5Ll7+h2C53JTePQFYLpISx0TO2Yexw
J8OQDcswe0L51sojUKidTxWOiFrSan/V496ShtXlX2Bra+I6VBFSxWY2YXWH1KNJ2cqZ4EEfMJHa
1Q4Y2VvRTovvkO1AoqLOPbXzyYl3zZNyzqI1WmMgAB94pWzlXnTGMf9oDJ86FoZQ9YcDYCoizAlg
UQwMxC/58oBi66iQlzdPFYUSS3nrujrWifNETOhVKKLsABXwgAbti+MQjaTi9eN+SnAqJxlmAnkW
TeGApSdJdCyvA/rZGTEQwVJAV82AepCAsO2av7wbHb1SRqMi4SQg5SCleYIrgq9EGvXEG/rM6fCi
PMkMazyzaGBtJhxdT8wtcEYE/FZmbcthznsihaeiU0elRRro3LPIvpqJDEljn18aYnrDUw+d6Blw
8a/IMUm+V/p9AeGcup6UpN7yqsc9YACPcNKTjendCQ1sXAthYIUrwbRNbYScHqH5E0p5igthKdwc
PzG/Mpmq8NKgeRPc/f5xa8Vx9yQazF8oMAepIPSQo8U0axBRhxLPSF6Y/chisxj+ZmeRk0lv+bOQ
plLkguKuBmfc/IWfflaEr/Nz0t7Dx4aIAknQIvnAkfRyC8+nu0DLFFnZcZ+TuUj2yx2njDGoQicO
/m+O4goOO4RFmrXv+jpXO4beDyyFCOwL+P9JQLAH0vO0i2QT0/3otJtQ4zvFFO+WijE/FxH/lWgW
4hBCVf3J65H4tLddjrSL6lVr8BeGaiKj3/yzGAJLqRxaDMoaDXniGpVLA99GeS+IJdsM/N5LxiHV
sD/UT5X2PEIcY6jf7nzZnHmmupqN5uyXjHdxPMrhHUtvkYiaQtXubr7NJsa0O4+ZxxQR/q5sBZY9
NZf4y+cTwDM39C1gOxVVmBtdaT0w4FfW+a/KwbwxdTvJjyVzzuhJoqXgB30yRnBknVLseRjUERkJ
zBVkw6o4V4epZ60eKlMvAK+28hs0BARED0vu/ETmuOWA61oG4uhzABPXwfl73BBPLhnxSsLkjXdW
ae+O55FPv/vkcCA6N8UxWYH8GMBeqIZzJrqZsthD21WXRzZdgqfBMEGIGjxwSvvis5eixDj0pgKp
ZG/rkYBO/C7B8emqCU4p8YKFFT09JhX09n0+/ih9wkkURbcP738sfWfB1Ug3qel5s5C2yJL8F4wz
oELE0Np8q72SsGcYCsBwufmmBixk0kZZU2kEPfEgJmxaJivG0R/ywzTI45LawXrDeTSdncByvD37
njmiZ2ISvpdiOsh0/upntvcorTa7Vw/FfrVsJy48yRgFmGvoFoZwNn5r03mKf0mZpqEPb3td6hBK
h8Rzs/NlFyLxqiXmiVUkcs8aFZe6YBJ2wKpGuxmco7pKTrry53VC0IhQWVIJ79P/qtQWP/hqELT8
wuAAeq8WGB2d/fmKxHlgYYOrebtKdn61jhsT+IL1+XADz7b9CbjnAyM6zgKnnNyV8vIfv3nfQMKs
KVi882TEKiaeTfZg/V6ldxNEsOgJtANk2/sJsOUlz3O6jolbAo26NQ9t7od/sZru381LyiIYJ2D1
Rh7ZitLqGv7y2z4X+agkweP+SySq2Hu7yAYPX6BpFkilhj3A/oRlBNr+RsaXqQcCY+G5Bf5dKMf+
XwZhw4ca3ATl7NtyFSczs0qMgI4tHMSPx/9ciPKYVqfxj4cLZhVmnP11J+4t2ACwg7gxfGGky97M
2buUSTqGJJR6BWO4X8UKid4iK/WFK5IZV6upQ3iIdPk9hpNzsh6Q4ckFDeNJo/v5Puft5kVBG9FP
zp9XkfA+H4kGf0ykJuTgA7sFfqTpA/wkqVicivEy5z/rOiAHbAnBkvr360F3NsRs/L8RbEtwoZO/
P8+fgN5hg0eL8zEofzYXM1iiG0Pbzl7buzMvkt4Qjq/reHP4zK065hzjju/NiP/UA1BOHafgWwOT
oQAftV7pznU/1zIWu3gNnIXUnzDz4SzooAvHcQneYSBjkJe59PwsHrpT9w1dU/ejtG2V9tH9Ob3O
yh1q1pA1qGOk6sSComojTmmU1DW1lts4mTuyaZISWoY1b0ZhWZvzWzPZwX82koGACS8/m8jHT9+8
hPyUuhqyk18leMIHAtsc9VagSEhTLBHMa7yWorXhS12tvDKbMluhGSrBdBYrr0dVFy4BcgtKssmA
S7crKTSEOvcxZ7Nxa6Rc/1zdEKJv4fY/UD4GuGs/jrSqLOX5qvVysyFUiE8n0B+Lt/FU8/bWUDer
0mk7a8n3Lcy6WzTSz8RLHWHpAwUAy2UaG3HzGCKbHaA08On5H0xsGg4Y/msq9R88TvAR91G865FO
cYn5wx67nCiQxf7YGsS0Olzc6wTc3ctS++/EQ6/eQB+ylGepgQQepteiDDsfCndKNxTGOC9xO+WY
CMeyZP1WEjsAay+rV3UTBqCHtJSb237MhSzXMqzyFgieGHFEs9UHKAMSm2Q47oJXV49VQshOgFit
Q1e2AueygpUBMgbg/D5vvJ0MaJ4XBGR/ZiX/0GBYeTxYjMosGLtXV4g00pkbFzvjk8tlia6hU3gM
9rycbptdTehpAdjxd7LJsE0dyywltNbIjeaD0WQJkPID9TbLt42SeIc9/2A4sgSh1DobCu3/s6HG
TKv5gTTHU6eK5KhT8E/lsNa9q2Ab6+MlxSzKhnLeYS+OPgdImpiwaM7M4yk94I8iZm7p9S378ug1
CcROWJRqqdpqIBcLzXrffJNo/xnrISmuKpBIFc7hj2gjQIjl9E2COAv9UM1mnQZN8et8ynGgd/XF
2iG5qShk6P5ru64xGvFqaMm4zSxlQ5e8VMyQvfAjDZmTfk9pmXXWtX728bsdmkFLDGd4kbHN1nVQ
R1/z+lFPAYCvwEuKGE9P3H4+TAj5b/GLJI9z5GQsY2h7+cvO1Io5l9oao/912u+uIkLj4Pwt3qIa
2pSI23vH5g/kjHWZUySCKak7I09u4o9b5xRwpecuwhyoJUSWmlbnxqiOTxqWA8LbCN7Uiu3ae9Zq
kXkE+GDXQ4/yfei4keA2ptcq+NVW6JV8Xion9kyva5ww6DTMRtl03gbgO6kSV9PMfyZhs1l3i4/S
kRwRF0yPQrGeM7p2t6Yfd20PTvDatIsqaXv6Zw2GVf8RGKJBJiD7utetMpAaPsw7AyzB6WsfST9k
e+k28506P45xHlCNslBWLZs45BO8MI8RdJXZWZSqhrr7KAxrDMlG70Pf09w5NPZBv2eiePl6Hp5E
jlfbVsFhnBQu/HHU7eBTbZY6cm7yZCQ66C3eG9qdzmzlfw+ESk/ZGtj0fU0NNQmOKlaixsjKq1zV
l89IE+BoRBWTQp6VRE7r5GmugrH5u1Wi9zvsyDOqcJl4p7FWFhLJAceumwOVmFvqXIzSUP6KLWWI
3k3bJlvvf2RKHaRJxapCLNFZzwJbVSEUTpNwKXbQclrDLtX2usUm5SsM0/as17WYaRiyQfjN63ff
wp8AK/MX1FXMggiiAAprdX2CZ0HFr1nAMzHWcZXiCQQWLkR0XCNbhE47eR9a58bNJFODVYMDXlWr
hNveEYdEBozIrK0vjcBkhLH7+M4vN59Lmx1/Smz/pRgoM3LYVhk11iZYMR0fEjK3xzuIwugxKN6N
N5i47XoBMpugZ436OlWhZP9wogCJJI/uYbfTgc7ED7X3op+Y8OZFgt3Olrh2KfJh9YCAVhqe0YoZ
up/15z7pHH7/4BMdsqKFj1SLwI+WyVBeWIfbaHS/16NO8WMGeRPuSQiUg0fT6Hk6FoP/M4samSAy
S+f8mQvfkLNmLCP66TtC+neGKu7yqFyE8jetKDYsnCHJ/x6eQetGlFjwjaFIajbpzbahg0DrGx5Z
1gRxLZHH8T5YrLnzgvul+w7T6I10Gnpu8/3QuehqS508DDpQY5NX9/rD0jxRerK7AaS8Rrt+kiFN
RzTuQVkv78A7NhBtHDQU0PrhBMudtXWnkjzbSXdHu9Gyw6I1osZlrXBnqxPkl4ebefYybrmaB4V9
TA5og3qU2mKxMDEpXUAxeBwSZg4sofEGlkGcn6e/8Z7H75ITReLoAukOGxY9m0ziZVj8dDz6G3P0
UwSpyjlwbR8XEx137n7qi4L/xPOcbKUL2OnxC/kxdVb8Ssj54rUn2rBEmoU8HiZCSBpDxgr5ueEu
9OSbZjIP7HSwv1TGO6ZFp4y5MKoHK0CaGMfLwpHifUXN5Ut1F6k/AZ3u1fd5G/Z/sWQfUJeByAT2
jcoffvDYMnAcjyQkSV3XKtHgGMwT3R6N3izDcQUWvsNqz0RfpQVvyQF0CnjHw7BQIIgQTomep/G+
XQ481fMVgpYCO0lQNnyYFiJ0QDA84SWM+MxoGrwKKDSuDASVhWWY8PZWkHXTbPJOJ7tVPRvwHlhf
KnwmnMnppkma4xtmf9DyDpqb5Yz1Kb6ozJ4IFPPmstGJr8DVKYkQvqtOI8OUn/UYucrqFFoYihrO
uhtWfI/U9gUxiNVCYtIGyTFrKCyqQmW7wJdb4qkslXvSOXufiEftwbC/XPEj7PoiXDgqwbs741ZQ
v4Fo/HXEOkRm5sMK8wJZhna+11gxI8EaWvZoIyAXWVLz+vJPftT///hyoGO2z4bf3EC0ahPJpDYN
VHvyvJWXxZXdgiUQeJQNU8Z56qhx02BtU2zuZY5LleLhZ5Tu7EYX7+pjvEfYEY5YjLUWdmhHbiGD
RXK79dS7yFtWGrpaHl2Q868T9GyGjB6wi4WCeyaAoDCBFN+pHhwmRrFph/GLZp/FP9nhreZSg3dZ
nnMDlSadBNX2odNFlPYU+/S7CX9Zac+AGCNplrpDeqSIhqJv4aLrOY0fU6cktQ0UbWchxUA7d1KM
NX1tWrJRuGPYjlYtRuMTPXASI6s8O+LPgnpcjuE004wxe4kyNrQq6jiIALZiWS2ZX5js62/+UtMP
8KxaZeZ03XoA3C8KY4S08+Kbv6UTU2Wh0FLXEueA3PnRkyU/GGGIk+HKy1uGVQUUxhGDTcT0cAR9
DswF96eBdc3LygAadaB1k8dahOTd8Srnwkd2OfhHbpiHoFbabuXn9rXJRqB92gAEoDes88NCdUc1
HQIqJVlFS0y+V4s1TQTeGtndLrOcAQ+yYBkgYW/+b/wfEcJv3xnxE3qYhZWo1iXjwCjO8OKNCwwp
9KGA2TdEgVVl7WeVsbBJ9bASA4/URxEPAQTkkv6XQAe0iJ2mTK5jesRUQAxW/OwMOxmRzfCdmdGl
q30d8cSzWw8wsGuTIEYAHJaXpg5Re2tgM3Q8EOnaAC/14BRG3NpLYLZvyIRgbJHuY9ul773u5+ar
ad1NUSUK5TRF8pYLdHC/aRnXpS0KaDtO4gTKD/Be1PmoQmax/ztlwmzRJXfz3Z14Fp0h3W8StkaP
w5aK7/zD8EaGU3Txbjq+VViI1C6Xz9kdwSQPxp0AOoR9KYbbdhMOoy2PyKA0FFVFD4wM3DTQ/i+Y
TjoWX0nNMfVPh8M77YcTRU/qzv6LX5NiRTtjj54nX6PAtbo88Vg3cIMl4l4yh9Cd18lgIvnLl9At
yLZjbIHK+0S06KOfq0YiY88I6K28YNRrtUUsIv7k0shfpojBS7p+EyrT4vU/IoNBmWeZpbNmg8jS
RMDR/y0cYf09qDyD9+77ojdW5q1LvEvF8+Xqp6Vn2hKwOf4r9eYJ4C7ROznH8szLeQy87LavmRQg
kAL3QUWcHaXIF4Xk955t5LohRZ3v+CzpL8swgyFpflTJCfve9QAcBFaPv2h31hSJ56zCj1G86MlA
pXg+bjOFy+ol9TDoqUh0hD/K85EltXxyl56FcMKvkQl21nGp6pNCXEU2FsCsWXgRam3zrivFV9yi
jjRdXUQG8fQv9F1BGm+po6J/TN8sImZJXQI0YV+5gqYBSCET2NtZY0L/1C8E6unCIe5nNtiDaAOy
gce/BMTa4FHp5MbDhalSlQGwaIifzds85CE0wzBkT3uo0g4DUZzqBhKmF+MBa8MZ+0Y5SqdhVi9q
hCWRUl1/3Lnw0YdpilwbVPAhXrVZOxgDTapE1crSK06y8Sg8AitZODoDcthhL/liwY5Cu2x2L+In
Rcx3GyvZQm7ytusDi5PXSG8H7C4qFnEhbzwDqxSpgm9F4zR77tKKL/3HMNTjvBpaL7S+q3Ak6IcY
D8qfzwHgPkauz5Hd852jCszdE/bUxs/+BfPyrXAV66fbw7MKao7FSAchnljv9T1Kp3rodJe9ohI/
cWWKtrX2yTSVq/8tfDsnI2GxmB7XpVjAq0naotYsWBoTV6S0PBbjBQlbN+6n5XmEKod15RncvOAT
IdGFDzgRlqYodz+YZifPnf0ql2NUKdgg/+NV7WF8ivRhVsaxUWtFbySB6EdgncymMpNu9u/YpwG0
+73p7q2GMCzc3yJww+vZus8LppLXrRQtb7ic62wHWbH1X55g8dN4zk8xyiry4JtDZzX4g7nQVyUj
NJHpDouazEkXGl0mNg93etoDq79X2HYmh5j/1b4l5nwjb+RE54z/PkQ21/qM1sw000/BHux7cZ3e
TNZhH2W2Z61U73EHfbqXSU3da6Lg2nh1KnimlVaPdnb2ZJEIDdC3pyorhFAur+9mh9FWs4Sskhtl
8hA155AIi6CqnbigmIr9hl80OWTrNlt7zkNKrxZtrlPsPeQv0T0fDG8CukVgjnh6RXMQzzIqsopT
rCnOJ8X1cPHovL+n5B6F97O2pZAMknT8TeTrQL9xy2K/P84KJ7/3AYy9epDuebeMXZmrxGu3OxmH
9i+fmIubI2QwXuW4YZh+8w1LerVDTxxjnZEY5vvG0m2sgdubBR7x1HzXmvC2aSDa5OnrhvVu2QYx
YPgMo4vi66id6oqPXrIjB8l/PdFgav9PmYP6Zn5DYFmaXBRT+4oNUGwQCyqfq/eOyCa2XS5mot/k
LD9dl0D9sO7XQj6bAYHWizthfeflIHfXnEDKmm+wJ9ZEBbCYm15DnhV3fMIGaakws57asfpkWLUZ
zL6E5e1PfydE+GU7FGtnso+EerK1E5H1MehOmywGFytPmmDJmHuAR7y7gRvaqrYGiV4Z6+O4P8FR
1TiM71Pyagh3QuU1X/dfyHQcm5T5BZYXlx+loSl1YSW4i8wielI0ioCgCrjPAPmRkqJDgfNTODeG
dQTyqSmwDLwi2cTRCvok3S2h5zVhp+LZzMW9ben4Sw4Lfi17igqobj+kn0ZESgsqzZmLjfiT9vhJ
v4Hxwobb9vXfhiC/ZSKqJmD59WNsKAYQNjuwDlV5UJB3DRZSvsjSfCB5Jwe/k3HN9LiaOg43bhNk
uWYKR4u0Mg9dEBkDqLlHwQ2tgKja7jOs1lh3c8rjAHiznxwxjT20WwoCrdKOI0yPnPkw/gaJIS4P
356GzJJMrY2iRI41v0dI4MHRuPqLY1mjJRzLiNyqeAUfVaOX136238vfvwN5NuVjan7M2u7cr4IP
JbjA8cJQuz+AmyKPk3Nip8VBHAFC/RbFYMFS8biQyjl2C3WDZNzUTCIYQ//8LVD/z7VUQi74zkPe
l47NjZy1flt+GB1r8DZfx9Wbua/noCwHARejNWD0PTVr+DfPHEtz5KZlVlIgjLiMi8ODAwNfnr8i
03WezK1wj4qSJ3KH9P5XNhI7vSuJ3aIifnlk93B51p42HzSOKz3LrAbfUtC6nL9bWF6+AzYmdrAX
S0TfNG4XNmagKJzTRzp4XO2pqk7QPb8wEddZR8dYiRfNtuMnynR8vW4hXNPlZ5GwtXJ5ZAA9yaaK
L3INvRG6m3cgE+QmBQwc9IEE87XcPlazzhL50shwEtObuqaE2/bGPs+LXH63UW1xtSGVZyPk6Nxd
irJHm2NikRY8V+BiNlHBP08+cMnAnBE+PCN9TzkYHp4fjd9SHbMlqwlBcJyLCiiyCXj+69afYNgt
Vs1SWjchAeji6XReDL2zvJd8KpxiANF+Y+yO4Flga6jPlC6mnLcVzR0FkvRxGRn+5fTe4y7W/AD2
ZN91vvIlVTu2vGSL7krJgjpuzbyIiqtjogqv6gGhRkbH+m3PMMeHTtC/oRvMQ12aTQcpqW/SZokW
nC/1nYh80l+T1qO8tnkT+AZWWCHKDorkxvQNA+XWpo6vAjTrNutIxcEO2iLwn2OmUXkO6BhHx2ey
Nbqpica1ZNc8Jx2+KnpmHn/m1SMKlX60lZD9nejq8OgbLEWJYfqcgkqKe4ZRCd4gardlPTXFJreJ
xrB8zJd979pioW/pZ9B6kwImvoa1HaEFgR7uLmicWrE6y7Dg6NVCTJVP3tVQA87ZivR+dtWUu2Hs
W0TGECBLG0RBwEoX+61Mzh62gP6qDTpOc7bVFUJY+NPseYSlgwLH0k5RYg6Z/XmKW7Frj9vfoRAZ
DJ8KI3pHw6li6dXYDrIURlC4MOlhiLgSSWGN7rNWfpslgQlsqsNcZuUriMzAQhlMJ5Lf8kn51omH
jPO3hJ23NfQMnpY5QsJLISYfQa7Enim1WZH2tPq4OGx4AiprScIw+pw5C0qMRuiGXUnWWk5EBWJx
ezwRsUCawNxKqhF6uJCefhTOT9zWBxk4BOY5BBnwuAfhEUSuLOhAY7ul52eYu48Mvvy5xPzk2YAf
uOa+6HPwQvIAbAgQdroDHSuPovj70othh56+kPFKOT5RgKLhJHlKQQmD2xSj2Ny0SAhYdLh/UZzI
6jELU6ROZNtOneZzFYVI2g+SDdP66XqnUK49h9qi6qTCAzBqL3jw2vZ8Z3ZX2A6Q6IvRS9axZmAq
goVDIL708EpuGEtnQp+3n7LB9GxOigZcAR6M/Q/VNyVtKWaYy+8oud+2k7cIrYVTXi7+I9lfuzaz
M6K7SyzpUrVukxzQGm6m2C/GHa2wPVjv0oHReiRGlk5BW+lfxC/LswQIVegHnZEQ3d/lIW1cZpsi
FlwVUe4Zt4XcrBqI8L9fZqDLu5mih66Xdtn/4Z70ghU/w0oY3WDL16K1eL4l/a/bk/ELVmYpyRv+
5YJn9XGCFz68vLXNEQ82cXOReTCeQQehAYE+LQt0al96GdS26Wt1wIuMSrEZnNdTdpL81bG3qstP
3vTecA7RbwzlWtkEzyRDywY9uM+gQCoWOTvA6hR8906N92MoWqC/h4mRXAQR1mT/Eb8gLRE3QEIz
y1fEuZ4ZrTtGnfjrkkoauR3vo4IryjNAR6I4re9N3V0Fg8BYtTvPLqnwiGvvIURb5O/5JRuyOCln
Jqj3Uv1nQldrUDEXxbtUSRm/n0ggU+SZPlaaEtJfj39tIVdYKo4XqLZPfD1Tsa4dsU79DbuFQDeh
+r/RBqOE5YJflrj/QgUgGb0ZD0KBKv/DyX7oMUYyOnZL1xymTYMGP6VMWYurSxw+Tc/GLYtdEqDU
0LM0Oy+VgkX6pAHVLaeJVnmXGsclJL7uWzG7NJO0D1Qf1jayVwtgjIil1JjBDVt4GxPDt5rChCEv
0kOg6/ixDY8CYFZ/iBKAVQArLwnBANcb1jsspi8m0v2eH+spL6mZ7qOx10gXJqpsvvBQF7twQh+f
+3jXk0iaUlna8mox3GTzMbFX1m122hmhR76XcJ0MWT1CFfy2H93VuZJ3uYXuYiv32igYn4kapVR7
SSLsXGWt4xcReYhNlSsd1mCfmJOl9cSshfVJ2F0oMFYyU5KCrfEP4WpDW9vZ5HrX5kyJenrmEIMl
phDiEQvHvhUPU6u/W8Cvx4JC7NWJ0eRenRuHViAcYGh2TT2nSKPKNi1rlRvW2Mj7tHcjaSWYNlfR
fk9cwqXCH7kOizAYRwF82U3Mu1tuM+ew9n9ztsxkxx1AO4l+bUfvbkVvFdW6t08r9EQKxvUTa+hj
XVqfj/L+7LT+GHvPnMZSkR2oSZMDl6xOSRInj7/qeMS+p6du6mOuAJG8Xvf5xJiVq5I0uovEm1B5
A5zZivoux9oNu7jqKnymIfPTconJ//IZf5peZGk9m8wzK7dYE88ukahDYpub59VCOcCPi6SIQCSd
qn+iWFeBE4RUcoiP4SK++lkhvKIJ8CACVGo8HebGeq11iIoZe+0RO4nEey8dNeYu5wlxjFrvyzPl
/eNZ6eg6pwR5RqMgpx3nd7b2aj59aADfCB8QMo6DAE/VZIMMTirNV1FAXvihpV4pxOIgXfuf4eH1
y121eMNiQiCXmz4vn/qXtZVqo8BST45f2OxkmS/KIKrUlt409RREbk+EoujqIG2/2gwzH1qttdcD
chqSKblwjINHy2q6edbIULefWlSMWoHrePwlBVIXMlgaEu4pOErSoyPeev3xl73HWsal9WjB1jRT
AwboHgoeUWc6gbmOu3l37qczvCeNpPjPxT+kZpUG73gS/9lGir0JgyZZciamzxvP4XuE6c4IKY6D
PrSQikhQV4gsFuo8nEeuTMHC/PCcvs+ZKHnR270ufYagDniC//nVef+6HqBwmo3zcp1tVd49i5mJ
M6dF3pukXQFQ6whoRqKfRnSLHK7K8cFWf9n7sTqKRuHB2ha2f1bP5PfEYHaioQVWvRgMaDVXd3ED
OWAVRDGJZi7+1DmSEWgFM5L250QyTaCUYf7wHvhlbQbEZjGj8fepL60mvbT0NiXXAFlcYge4sAfR
xaLAeG7+OuCaNWw8oK9eqiQfDKIbeeWAOCHYJ1FdnCJXeBiLYVFnoLqtVpv/yRb7jHIEwMdUxN3l
hx/vvKJ4rL2Ehg2e+uMfQNasNO+olg5rXJCR2QUPgKg9av00kJ+5vgzSIlfdR+VGGITwLboBZmdW
gldErTLa3molxQmaNBrjVw2OUHuphYR9fofUxI8wgOVJ5PcPYx/C5pZRQvGEphebAV4ipzW9m93a
NVN9MROcbFAkX36HhYaZwfE8aYd115RATKKomuBYT7i4lLeJuvjAjedgfBo/aPk9Mc5e2HOhyaM8
iaJzxRtM1hhHiwj7Yp+VJcGo0jS3VmN+4Aljf7xUSi/MGOS1/k0O06wwvU2QL4XEXIl2NogZmk7n
DM9d8qpe0tu7UqNfliQ0360VMHMj7MVF9CAqHGeINPSP/h5akn5TIK9luvtyVoP56Q4R7cx/MaCe
2FRwq2M7bhqwNbWq5Q3EBfJaZONZtO2BUO4kBD2GW5zzqLRFCgxp+UH6VoDECYvOTBIrxoUS+pPj
luZRqcrS+HBB++WOj883WwAhbMltzfLSq1ZyFLxzYtdClcuIouM3i57KoTxod+3nVHvk7yy75EBc
43jfzSxyGj3e80TqNbNhV2F1IPoh3HnsUgBJgWQI8FcZBuC5DLsPNHD5OeyvA1w6uZUhNVVv/7JJ
/q//o3dSfb7bLVsSr4zvj1SjLe+rlEbph98Cv7fSOlroxNvsqWH7bV/vM2qi2SSVptsyNQ6QkRSc
7wIW7Bec2qGCSTAgZ3FLkQfOBV70yGtGfKDiKLCrnx2QW7GOJb/BNSsfK8CdYzgAVcVNaT2f8jQi
3jmN9FrPHnc7U3mNit38bZ+SOJTeFtCbhdrmuwBs4z2jLzJP+/PW/u/c7iPkY4s7yjWwnXKDCVt9
XlDlHRBVIX4sfrltEF3Op8Sphgv+SctrL5A2So7zu/yCyFEdQLVeuzGK4kYmzP30kb13igW7+mPO
kl8zjj+q2v1+kQQA6WFvzOrOAITLU/NhdLAKoMALjCof1Gp1Mkui80xLPL5QroFQNYvMH6IF6z7w
B2tVaFfWul0Nod3nUefC22sqgniaMOXZgmoi2PC706w7UK06qhyxf6IeEoaojRPUnXGu7wygE2h0
XisSHFV1Tz8IsWOOyLorxLyE+w6FIPPkjnqnH1iZ7c55Ooc3Idkq79fB8OuBmmm16dmD6355gJ8E
KEspXic5f8uFlI2jU8S5fhd8nMQ1MEKmaniZnPP4eszftbR34AHUtrPgNC1MUfxbYBDvLLHNbL5d
Oh72oqoY/QvusU9feLQbRY2S5X9uWSx1jeHlcMfpMHHlipyKjBlaCtMQx6dtaOBF5vYTFoYiXc1w
zkxsXtX6nmaX/cO/+WDkaO1TtHlfNV3UoZl5SIkbnJcAPEX6utsI/mx2jIrbofywEFSJX5QF+UCJ
xI90fPBvlscWZDsnBagtQNyFLPrcosxV0dGYKGQiZcOudCBabzVWN+hbZy2aGfaEJraJ3pA6AiKn
7/G00gEuKG/kHisWm7HUCLDJbY0QBvWpnYtyUdH4zema6yne3tVh1475747ygDqaB3UPrAtzNqXb
h5SJDVDH3e+Pp+bxiCFpDljUJmgjBBu2F0+D+9JURRf03un5jTkXFYBZkiA9K4tuax2SshTpMicD
Ty06tVeBLFoStaQgUf9g80ViPcH729fsWNarhyQbxIUBE6FzgWR/t/w2w9BdeJ+NJ8Gzmg97M5v3
YVutZOUqZ20zyI+pgvc1TZmGQozn/LoU89QR86Ao9jKasIh1ZFQls6dRNiSXKzZYfLJybG71/vj1
9nOkJBX5zcl3Q/DAMAsWfl52vbUUC4Zl9o5zXEe+NcIEyOC1NpA4Eo8JU5uWRAEMYe9aI/cqZ4fO
z1hD3dE55rdrZN2Ypw9pWyYQbaD+ObmYBjvGhV1RfMq7vOYbCoIRoE61ZnmeVpfMMFKS0wMGjs2a
k01NFTUm50gMZlyZNCAD53c26JxucJ/Dk5LbRNSh4Blvaq+HKjZxkACA2zpOkZimRucWmdrAiUXm
AjxRZA5WyvcMYmRLo7yQRwEth3ksyoFXQq7UuAjVPwcMuMrVDRNuuyhnxefYmGzcDyLqDD1j3Y1K
CObq0qoGlmuKQM8cEyHhmisq5j80T1CORwf8jmhaMjVNS9oqKoxdJcUNCkx6sc9PDrp0o07wM+Ov
eOM1GHIP3gbD8pQoFQ6lho60a1C4ohGGDAmDb9n3+Ty3qmw1o1x1Y8wRFvOZLWHSOgvvq4AOwjKi
sJ+jCMzrlydwF9kC6JL/gpnSdUYEq1dt0MiiiNI5R2Z7x8yaToVyFC6NpGJX5Er7+VvPi6KbkuPg
LuBnlSjyucr5UXZQuH/nNzYBk8wQ9mZ/L72wcEOKKaL198QTH48zNSfIVKQaw/QOGEpfMqr7s0lX
1Qtw/AhrnBohl28irxw6VyiaMO9o/rWQPiJrSQo+nnOSussJFWLWnGNTj2dNEGXrsQP3/iQgsMV8
S3XBIn1si2MylHY1AnQaG+S4117o733NF42nke4dla/W6Wbm/2iD0BBC1C71OP6+LaBs10j8cn1S
Y0Cv4mgRksY7++wLQvvKZNpl8PrnUTD8yYVVFcEuTKYqxkaQ6m4nif7PzG+qU+QjcoDCcKgu9tV1
Supv4VAdxD0P7ZRSAfvAEPLlG9a/1Jxdb/N3cEdHqsu/7kJ3E0tpYI1HzIU6Hko5py+hVcTzCJwN
mMri8TR+5VacT5DzwZOQ5IpZt3UL6FUFfamo61JpxYy90dxlO8drcFDHpJ7dYYbHSJum3tGfqyij
JaCCkU9vCH39KhFFBiRR4A5xrL4Pb87r/fNhyUwpP2Kpo6M5DA9PG0/IACxw94Vox7N2iGleq7dX
4h1kpz1q0PTxQS4R8ThphkJJ4j0MuUsW/pDS7dtWfV/C1pkcmF0NRzoUqyytekU8WiJKwVE+7sCX
kINKsRUO0YC87PkOp+y36U+J+4ySYw+idIM2vmNiYqc2v4VhiQDw1dw46SYnDPkVJLydpwnzMyRI
boI1eoVAhpa54GyHRlmoRV87z6TDdwuWZUhGVE74uaEeEXohFBsojwKcASzuZ6KwnaLj//idw47P
3SDPB4s5Xl04ns+qPjqS6GS/E6Y84scVZBlr/dhfMCUgAMFHXOMmFornZimAKNJDTenihqQ0xUbd
wuCsueIRtSHwtN+OG5f7KVG675EITyrCarOk3Vi7iYXnrEX+oioGZevkb6jR0Ogu23Jqnw0urS/j
5K+MGFqOeCJyz2L1xvOwtPrmf2q8sSKAIHcK/fYa1yOPmRO6q+pSstM11m08K5IfHACMuRVKXiG1
EbUtsv7wuu4QzStOVRe0hASu9gAC9q3dlfZpFRqPTFlwTyf7hsIuzbzS0B3BIilVVWq7wP1DMCl5
NYh1l+uyDoHiHir7ZmWnQ3RyaIXGGi8OJ8twMgv0R2h5tWn1d2u88DFQwF1bAMnYbXKBycj+GYch
ThRb3yKd1MjV6YQB8cQH4bblWPdpPDwJS8yzB3v7+RaKO0FiJldMNwMxtLULrDqf9X0tC96b1nCL
QVH/LLMvDXZ4tcx9TUl72EDQa72a58x1YXkovJ2njhP17BO8r1GSmml/jwcc7iVlMH03i/Qd1lvl
5ZGm1+pe1/R85XoeyUJtQYJkY14Mf0CAduXw8WlFJ5sMfMFIv5/LZaLu+y5m/fuShLHHwZZUgSty
k3OIGZ3/hoES5dZAujUnt1o42eQj77LO0ibaJuojGeXwZad06qNKNSLjc1V1ZqzrQGkNJkBAWMUg
6jbXE/YgFqO3G6k8UVucHWVTyQk7GPkwSpbSVzNLuku/igjFkjBtPtWKJF+66y5YJ74n+I22s1lE
QWzMVnLNMUqK3ZTQbnoIbwNoqpXi5JPOpgNWvk6v9TRrVKBzmgKButMmrX9gTZYiLu+z3T+0ExEQ
CXcBmZgD2VFLZr0S12rysxcl0QsXwqhZhtHNEtsjzWVksVvdszJagmNHWWeynl0pON/4bb4GB29V
rAKTfG9nsQAjx6ZitXTuC9/xoo7k4ccz60YOou5EReSFX0Z31FIS7Wwz+KhV749BU4izvnzC0UV/
mAgCZ2pyyTRNjRenx2jE//y29TmGcrQSTxcOGP2qwgRcdtuGZ4l6g3f6P2OoXXiS7glQVz1ugOEV
rKErg2D1f442aAJGfsr9VSSVWhWlxRkRupCsH29MzMluPe4Wj9gmkpr7b/2GZhOHLbmxCqY5cPv6
fYo8Sdo68mmU4MCYO0ugmdgVwv6TRuBvCq7V/11hAPHYbq68jUEbm5LdPQbqd2CfJippceEa6T9E
EoqYJj5aJdXIK9IYCqhP1RUPbxCah9S2BRK6jy5me+T8dDt9kzLYZTORDyP03/T67ROvYyvzhA3l
FoqOo256mtd2HG9IrMnEmj2/PYD+sxBeHfry36eC5k+cYih0zTpE5vCmBDPr5xkC3AXl6l1raT2O
aUNJfDXvYyQc9Z+XVZU8Znzfb/GsPE4M1ulj5qwfOGCP/4XQjb5jxXMo64fH6xgyYoKlX9GxfIAW
kO/KK1EGnPD6DUI1nHLJzHWcAReWX7DrVO290Xh5sEQaEqo+PTAEYp7Km9ZlBwuaal6ViXc5/sgc
2ChjMp8qQd8cxippkdvCJrYB4GsmbfBqkDuI5uYQ5jmI3f+Cv0hZAgQ3FMp8YhG4WdiHYozjUeNe
7rmtow7icCu2JgsRVoLESuHbsYkuNAfppCCCS6VDUBfNDUzWhLX9d1oQvtmZZY9dNaFFfLx1R63W
MLnFhOQTCkdaA4irfahs7tER+eSc4FpKHEZT646Hxx4T6ClI6EoklIKxeBfp8m1FZAZ7fGMX5k66
J80iMDXvNpjzhgefrnmHIn1Ybr22q/AoMIdkzJpqbObqew6Dwz3ChwkqNj7IwAg75pOXWzJM1uaI
yqVKDOhCeRTj8elavKKxTkHBoMP67wntt6JJD3GG/c8/5OdqrkirqDThmEajU/7WmePq4NdipYi9
lJ5CV0UTTH1FjmEv8AHKE8XLwjKv+lkpwFKOIFtdND5ej0JTuGxtO7mGfHOpKPGVBiiaZ1+y9Pra
mToq9XI0XUSX7Ui8sjEeyPsy9wYme+1t05dDjc+Odbtdg58W6DRV9oFzlTLq9elfqeO1KuqYwX8L
Eq3TwEHB+wbNakjy2MO9aXD2UoVAXlDzj7iqOw6RsvbCunhCUHyLXbdkSVz8yE5kl8m5+n3TEEJE
Nw4I/pWj+arw87RXf4dR8P/tgtA9WOA3MbEMqceCbj6BmcOBDzZ7x+AeHKJ5O97+isIvVpToqbKD
yov1QIPZ7bUYd08iUH4e0EmsqmsPfXb8ShQLk19CoGNTcuGovf+sAAFg63V8BdryMumWEpeCzi/d
9aRmgfvsKLA1+3k7in6t2F8W6l7zBAKL3sBfor7bZ5aFI3vk3QTat6kkjQLf8aSHreGGn/tRwRrm
oIF7qSeZ5+g8z3z0sRZhIcjBu2DVjw1GlQlss9gC4wh6zZWmI4ozMuQHR143uB8zf4HYcDM8fA8U
CFmTMNOar72JnwZoZfv3SeP2md2LTwsNyW+HFGFFoFfmUYIGulZo7y8IGFD2AwCjwi8f1Ovr++R3
xkzV4LqI6dH/jBaNHihp+yCb1KqTL8Jcqs4irRT3EhdIKT05195uacjEylgvxYZ3lWLMLaqVwWG2
gbFe5WEaIoMSHtN6r483wec3PtCD+tc0J4UNBI83iPSxROeHWs6aSzOOGUu+ZD0HLVUB1QViRMae
gO3271DYMgwMUC5zZD+zqQ2F22pPbfQDrz7jnDeCO3xsxGiaF5thcy+d42c1jbwEaZyLyvubgajR
Bg+hLmO30TTmG8MfAnlE07jGKs4+gAL5Gv+sWRT70EVXebm+WZnTtRZv9xvI/HRZzRzxxmztsRmf
tiiN1QO51b0aQHWgKejBV9yBC+pW5oYAdZVGGqHWxuuIY+ReLofqwQQ22P7ITfQXQH1RHtE84KPy
yMYy4RL9iz8Vfh5UsIDSLgN6amI58RsWG8CPyQ7bPro9th45JqEabFcaeLyyOcBmT2QUENPNDs1h
PG+k2nELhynQ+eaMf5aQa33CUcZ43jnDohQuhMChfUX2JefhhsjjhfUrfflV1T/TvIncqCSCniWc
iMTjU6UJdcjFuApTgWm60zo3uCwB4Qx94fv7MujJZlUymKQyEfoRYAJL+x48Tz2jR0h6ZyJcB+s8
6rUPHEJu6GbdAmZV9hTYAq8mrLdLNwGTJlU+n05CMkDZKRdLCht5WsDojg8xY35FZFAc4Km0Sxcc
DrCzKBGmeVGDDBtfgg+ySoh4FK/l9WVLJU2cwPNoFxiiv1iJiy2AjqAXO/EEHnPraWiaK5hn94MN
jPXVKR323VwF3CuO0DT1qstgFZSDW2T7DqeNZv43hgB2hMuE60ThfXAJySlfzmNEyNzaOC9RGLvf
CU+XFFcdF/uy5K1EJIxZTctpDd0BgmmWNO53+2snIbhDdgUsrkqTYusBw4iyPX3pK4BpV/jN5Qj3
ej+x+GfTgIXjiBuNfSRcLqsPL6AJtuT0KEIFqfSo69ohsowJyWdHVm6mFX60MZY6Fbf9iWiZb1o5
hHLrvCmwIL+NyoJkgNoejmB6k6cnIRKHPQMgGX5j0GgPD90wdRLwVNBXfhrQUrP8dplhuuvR1np/
5XQQVICj4juLqMMtzDHPoSuv3GKBMpG3J39K/D14JPFK76ypknM3ToRxaGfcueEkAkTJr+zxbhXE
MExDxTJli5uUtQLdhtnN0NyOh+JNgEoAiXS0Yh3ofi1Z53rwCt4s3wM0N1kSfs7z+Hk03RE6rwci
WwMPDQvKqvaM+ufBhiB/0cfxgU30JjUHHWtGNmKwlp+XPE8JVKeSrTsUrIJfHomNYyOz9MviM8Y1
VyFZgQwsOTj0Y0Ug1jj3c+2SzkfxjNwJcVlluAcawA5hTUVCXuri8ToXTAwmM1V7zJExg7/BIrHK
mwoK+6gPl386zvRhCpOTm8QuEdvi+PGefQ5l3hrWWjIXiDTW9ZTFONJZFsTvr68IGXWXsheH4Mce
AL7G8P4x2rsDsdUn+zGsv619Wty0SQd0vHrxbrqUTpe6xuq7Wt6A/Id6oDPLzgUiSmaMXZZu5W2Q
Vl5h2wvGEu87S1sKcx/ldeA7u5afd23CLvr3JcVK0ChOYO89Uj/VCrMmOUVddx3JuxRH+y7Qq6zK
yZgpkuAopx3L9x9urq7SrC92PMxNFDP5RF7yinwJrlNxx2w+4b130rUcQf+in3NuW91UwFUJ61OT
wTcJqfad/VKuaqfhfYxyNEXLPbvsUcHbOi41wWcY/GxnAzQVpZ68tFQGdXMHjH3pg+34pmax9jC5
+1kwx+5xggzG9wEz7EcAAPZPjaAlDROOJW92W8SBGBk4sVNhs9LjCFDjN0K5qMR1O8JXRllaoU1/
guBxm6ma3xQW9nSctx9P0Sf0fpcFaqVV/BsOo1pgtbYGDDWOwmc9oqmxrTDukwrvcfDA9KBC2/bA
dMO4Wic762WR/eCsQFIXW/6z/M9n8YYMQDFLZ2QsBTpOYR5P+cIeFZLlg/5UX4vLQgFw1/dc+gTt
ga+Zu0+sb5zgU5G8MoaTjWPk476zpzW3+hNnSEYwHlGES1IIgvdZ/RqTlLNlnS8zaXahFUDpj0hw
m75D0FmaRrLOz6SiPzytoqavu/KoFJ8OHTsmGwRt7+QbFtntelCbjI1ZbbLi8alqTyvx6OSrEDIe
wPrH2McRoE3rqeNb0uq3ewdK/JqDiM+nM3nALKUmCbG9zOdpIAaesRi1PwSg5xvy5cj2/lkMKDAa
d4Ug871KUqi8xpy+2pPOhtEC2gGOnnb7EcFvB7v2IlJSBkY+yOywKrkmcrGitZ7neuSo7o44Ym0Z
wKjwq4sNbEPP6ZombC4peCBh2N5MmAtAYtc5D5ThN9ZD6f2F8VnIL76nct/uF3ReQfgMCDfaNl8i
Al6e2IPDxDXG4ONn4UztXVdjExRqYdwwox3fHzdsRSq5PDNSRiaS4CduSLZGfoNOeOvHI3MHx9ar
cEajiHxZePF8+6u4FcQYVdWUNcuVB2UYZsYZ3v576m6yVbwbhb/fa5m1OWWfBRboNxe6/pCVwhGT
FLnck0mvk3mWaNYc39qLsBvU9KemqkrPdregOaIczqQPRbcrHopviQgK2aDYIq08OozucTLm3iza
2q51PJlxjfmSAM/SleyyRQw0/rzNOLEpFXK2Xjt8Occ0pXyB7HU2pIlJ4ifpvvjo6/skCyDNaKnj
bZavOJTCpKxavVrAUCWn2/qTMlEjx9V0AshHK6hNwTSI9tva4xPHtZxPhpUCmyV6O5vIE7mZ93s6
bpIzK8AdRn07UrehpW82SKwZ6RT1AqCCFQ15xCqynKac08MhDXI+OhcRDzY8orI5lHd9X+fnBBpE
L39vH8PBJeXOm4rF1DLgTzM3My8TEeQPQKYBi6/sb/8AQDwROSSEIbeK5ht2ERydJHZZuJE59PSi
TJmX30RB03WfHFy/pPTVXDsIbBd+pkZz0JbAXzhT4n41YJ7faoMPdhj5J/fYOVNiMysVxsq0SN6V
Abo9DBncgbtNxy3w2rK8mxF4vYUwQQZ5Xcs7TZOBjGIIhf/XHKO/OppjSEYrH7fHoefKaFCZWlIP
jt7LVdQtBS2CAsKFjSrJ2jeZIVO47ftwH4/mQUuCH40x0vRdOD5Lj/29dyWL0D1Kgrpi/0rpFZoM
g0wDUobtUC8LdtM4XYsQ7Pc6pi9vO01XETZF+fImO66TKT90YjRR3Fx2YydINS737gbMjgfal4vD
Rp09Tc09l2DEOU+FXrEwiYndsPs02bk55L2xiKAK5/RAlFKIaI+LW9kuS7iOGLvrbrHDqG4ZG3eX
P696pU2KN9z/awpSYhj2hRZq5Nw+nKWjpxlMDKigdSpvXp/irWNOkWTM0xQgLwP5rmuF1iWdHm3X
EH1Mc/WuuWvxesgLh7vxWFKir2QoT27BYDN24jo5nR2A4xm/jOiaSVqB3XM70UrE/fgHbvZAGB5N
wQanbdYSWfvPiRkfe5h1R4P/7mWCUlH64H2byykLNxaeqIFa8CrsAYLQd/kwj1G1joaa9pKtffcU
S7mhB2WMphawmLkhU4v23JCt5LCa/eP0jyHleuLJCZxBcQC6ZJZmDH+XLZa1+5wD+uEr60gt95Wf
NLWkfJNguudraSgpYxKUYxMbBtoRecd1iZB+L6/a+ZbPhSKbgG3A3wnMRUxtb+LNxhDKtF3znojL
iRPBTb//0Ag1dxGO/YSHlhUXqHURdXXAHeh6YNBCkYc6MFwvHMgwktR3cfE4A4ZMU7iHqV9uJODL
7bzYCZYI9YjoHShtAWPhYPRB8UDRfo+yWlAnhD65XUapV5t04BWnPxxiPWT44Y2r1zAn+CiQmlNv
70Ptl7CEMgxkBuVJ7mhgZ8ggwbRcttBchXrSSS/rqPkk0NSfCDU7ic7c8l3EFKawNkdKvIi8cJuA
s3cApmVb4IRqOnK6djCd+oKzB9zYDV5vcvWasny1vLrwXqLHchCVQdMIUXBfFzfZyIM+hKiga+GU
pQdN4wy99Zkok9MFngh5u0o/Z1tco75lisZwdoVrzrljvkUPT6rFHWliIlp82PfBMNf4hXtm6cd7
GarUzYjgke9ZMUk77i65WXsv98j+3qe0C2yXNGehRwoNEvvid1a19OWhSaMwHDeNGv0vcjk4pkbV
OGawl4RkcRGxiBObHyR+wKVFIZdjAHNwRu5OrNonaH99FOij0QsUP244RE2M2LVjPyPMF6vUb0ON
mEBuLqrDjQSCiN9xqP6Hkq3W5wmlnshebFgjAPigFzboygeO+MgJ92+nhD34+XtcKLCQMeSaJCAM
sFvPx1QMG4Awzjo4H6WoSPZIZEanf9J7Z5fXD0VMi8RYUbWhrhwX/mJay4Z9Q6IOeZURVrSxfIOT
49VRCh+/2u+HXUKW3vgxEfxkrhP8FjwuO8TU9Jh7vXB0cDQlfFqn4QC5bHLBZ/5xOHseS8DfUztt
+r6d+I3JcKY6Pi7cX2ICYRH/gjxlyoeZLahk+jwGkjnIy9JQSdPiXE/qPzvywkD5qRNKvJ21WGQ+
WYmFdMHJ0QyqUnT2wwQS252BXD0p+he6vf1+cgHKBbxnqCB+d27THQJCVcZmU+JMegcFGH99XG88
Nj0FSsZHxzoJwafZP3mTz8VyI27JSw54bAyGD50KwGGTCXR34CPcanB9qQgWvXgsBeTW9uE2VVwT
6iq5zq+2Buu4biisNptypmNoPmOm5ZgIfYhLnVBCkRINsWsbf4HZGeOWzLjWr75Bu9MgVZjfhhp/
pr/J1BVRBNZyi6Rc98mBvCI3wyRBiZNrZSq3pn4uYX6kJ1r4hyQhE2NaE1BdIHz+FwsgFjc8+Dne
Nq6mnTS0twzzVWMssijf1UHe7ruOZyZY3F06gcUNJZgSnHnJJIXr0UGx9tXBPwe3UPAqJuqwbL9Z
FZhrB9MHp+e9Gu6nPKsdoH3hGG2DhqZWhkAx4K/d9+drspki1BmVWWYi+G50a9muGfDxRQ3O/X8Y
dxpugpGhEXUNREzhpARZG4Y24qKdW4k5xNJPSFDEDwZNfXpXsJwosIpaBECzP5jDoVPjQWgGEEqu
izkAAouFJPxBULm+lYB9z0Evu02Sm0mLkJ7BA7q2bxxgbxl3FI4nWXaMpbe6fbdm2PONW1w4tw1j
aGCsOBehIQw2UiuL/XWE8V5aICOrBO3HwXP2cvvjlYKHD68LxsBxs6pRa3gSp59nV8lnwXpAzC+e
7Zn/hBqFb2NIgPdYWxkBQG3i8Ra/vQ9nfp35OBuMnzOXH+3tyfztGbNljNv+P+12XDuUUuRz/xZi
shxRvAetZSRvNktQK+6VmP3auRz0a4HHpojCdIXtVYOekwWu7bCZfXe3yASu6BBphlBHAcWd6zvJ
VdA5iebAK2WeqwID6AcVmmqhNKfzLjHUkfDBTPh7FiHZcVVkzxNSUdhJT6rjrvyPtF2pCU6ZeIMo
TGwuqGBsE7MQzReD+Z+kfQxoKPwuIsO5nV3FKHrDgHS0lg2SILJe+jJV9oYrWVxp+EPWHmj92GUN
VBsOtmEoRgLEBGsg3iLj1ueQPCbKhvj2h9pjgkYE8isDWRgcVHUvBICOrvbPJhiVje9tljoKGLut
8Ak1XfOpmSzSfbWH5a4QTiVDETv/SYPSwnHQYBLKKi3ZkuUROAG8xEjol8hKJuOuCBB1xSyfIO+W
imLllvJ2+jONZrP7AeXvCrcloCqEunAq0caHusNXWKM+n/VKbHMc2//cClsYDUd7VNLGwz/sQaPk
tM5MJmHKQd6gvkCzgxnDEkWzpbqp0+1UQeOB0oXT/MzmIsz0yqgHJ0I1CyZLEWsYGS7YSWJJOPUs
0nHW70o2PKDubVuCAcldsRy8YTlLLZ5jcjonSx85U0rPY2UTDNbuBYGDJLXyEY9edkbYG3r02A5C
Moi9dGh+I0izpNxanKdtf8V0WrZ7gCehSfll2602cTXHC3QWuETG/B8o8A/30KwMeF4DjcWKxaC2
kTXIV43lRNIXfdIPXXEaa1I4351qs3rCzuNb+H5sF1K1L5Fu43lYw09tkmyAbkoY7pmUwteXN6Yx
bj9QizbkRPltEOJMmMUQp4HhykaX9P5brXQuRLnz2HQCohKEejbHfA3FrUVimUgqwZq9l77Uw7Ti
s9QP8RQmZg5xMmU3HzalE2LK800kii9YJscWVL9XwNg7H3fPqX28ipHiY8tlSTgR6eZo3TBFgSbi
rte01MFOuGTurwg5wIaJcPWvxcm/+DL5vJ+anpJuUBFdFWibY1hOGuOA2CyX7EGgCmsJ2AjIj93/
O4DLa3srDeJPVBedOOw7Go0kNUjcFe9gdgulz110xXaQvRA4XnHaDqe/olyv73XcDMnsjCpfZq5J
bGWhtwknutQAmvPg5g5J2DbvZPztr4cnx0TunVtUpggcvUjeyfJ2JgU8YrkWIZgCiFYfsUUDBxH2
sZJxfgSDMWl1zefuyTMtuJ8suQsHaYS1zsBLItH6T6gOzj9xa2zBYix0HuPFEkX6Yj5Z1vanLHzB
ilEw3Bs78ODpx0FRJX0f2IyQ0WeMum2WJiaSnlzk46wp1xaQCRtL/nHyGYqxrT1d2+XtOxwfH2uy
6HfkAgoS26pBERapzZ3Z9OCaS+5hZbOZgBGjhpnG2UW0z0fYGrolKyUXsOJbVNc5mVFQUHtLDZYu
VEI69erUVMn50iWFvJG85wJVM4EpV5gyrCop2gq5dMPH7m5HKB4G+y0o3HFQqBQYLslMVvJe0YKT
zvRyxmYViyvH9D3YlizLJeAT4QQFN5bFkQLZrjdvY7biJnXpR5R1xFiTTQbmkhvGzYb165l7YUQ1
Yr8RmTV/9myXDiJSZjmKdva6Xn3wig8VxsB9AuZ2kvElx/Fm26jKADwgt3kh5JDjZNbN6fAne95z
0j2fWUwTA4+E8aXPodnegITmfhSSJ56ric1W3zGNeMIgooXbfVyxaE80EsjCo6pboi3QihJyiPsP
DuIyRUZFHpCTIo5C5KIOHVErUWHHwXCItCUaLkJkf91W96dHn+P49sBNnEPrrCsR4DUsrfBTgEVF
rVJeHEiQ2L063fWlaxYh/nT5Xf4mFY3MHaRJ5+bc5Y+XHh47CXabtNFK68GqTMZE649QT/xMBp5W
XFtPHhhZOUTu38pbYYwL8lH3fjrxiSKvTkobBFbyumVr6TreG9Xld5mEzA2jczvdU07m7Bi0n7bb
2Wh9K0P4GE8As3Crp3t3UJ+MAaeBSaHPm65HRQawaiZ25FI7IXwpyGW+2uhqrhnYLY8XJCor+MFT
MAJAj/TtPVTcrQ1OfE8BsK8TjRDIZIy9DF5NG3Pxih8BFANTspmLwPLlCUaPxtuJBEBaTFHTysb6
HP5nWcr1hsuCXRCtjRcvCO0kMDOIh7ijC2+CtBOPeFLgaBJtaZ5YVJaGxT2S4GOeX7OfELkwPmGz
aNkq5Z9GzSuuBZA6En3z//ttfveesI+OKboPDArziuFStcnMDtwRIAfIL5kkT0s9JJInqRnbghVz
aBS7pFOrh1H6JVKG4K77Bh8jMTRocoEZ72D14gKCpmrZ5fU8Ulv8s2WEO1QtzjBOY7km9uTo8eNM
O/E15W4oHXuoLuZcQNHRfOegQeE477tKbSODrwqCNcKAFpsb2Z4Nb5LvX1L92T6EvvD771kPiSD7
V6BA2eZmAVXfAuh7+cUIxsRjspWOcSqPyKqhLtxxs6Yjtv6GfjicafVpzl6wArjP5dO797fiTag7
7WY/1cwvnxBSYhTgzGiy3D/LJSUQrcwjQLLphpsIOKqA/ux6rDhrjMCvnm5AmM6UZskhLR23UMKr
TTs8CFcMIqWqsL0XrfgPLt6r+x8Oc0rGYSW28zKJZSwuNgGpV/0g6BOLXkmEAdJct4WHRKkOk4IG
SvyBWJx3KkonXunBIqvf0dKQ6dcR88opmIUkkCaDpYkJqcuQTHN1qnHbkb9LQiT6Xoocz2QrCMg1
37BmNiOgZ1BjZxEfSk9Fw9kOoEgImZVZtDfdkD1I0BXKDvvfBdhxUeYpwBGUYU2PGytcc1pUQ2Pk
One46xWf04b7VLoOLmwgiUwnx+JuVGHt3LKwrbFXCOIxIdDfrONVxaP0uCtFwxDXi44336mTfwx9
fugX5UQ33AfN9San1v8iNR6/TLiUZGXCMI1uDSsuRuH8sip+vHahrfaR/LXRSadel+jm7OLyNGBb
Xc4GE/4y6e+FiQuzP7RixsawJcSUdPF6YmncFDvkQZ+imZE1L06vfMN0DEY7LkwH8hO+eLEq/gRV
MxOYfJFrcVRT0pe+OasIyr9k+LNLzXhlIIylJltIjr8grsnLp1RQTNi46v+nMVgqBWgxoaO0wiNh
zXkLrwqgrwFuiJWsxgPZPluabxP4K5W2dbjgJ252XvJOzWwluhW3LEctHyfImRQgEPdmMyLJ7HK1
yuAI1Pnui2Hn3+mT25cMGYnlriMIu8Dv/UM1roIKQxmQjo7XleVdAYvm7evGdRbcoh1yZymii7Xm
IA4+IZ3CCB/p5PWkNApJXfhu0xuk6n1IGGC8u8l75l6uEGhz/xWoA4WUGzLTfgcxd16mNIydRK86
NhcHdG49eMI/Fd6GCYqYA3S1XGyQpB8+yx4Fr0tkclljEsHm+IxRdPn2grP7ZDIHxTIKSZsERSxH
CUthuiV4RzgGpHN2SoHJD7jB5ETU6lx8a8ifysbUlp+Eo4YzVLluEvvUNycCJuFJMTxD7PaNjiHG
Xl5TSBXfat+ETnJM65XqctlwNuB7mUdnwntKD6AkmrSxOK7HYSeyGHTdNoUHKVx0ar7DYvEE1ins
ZdiESuX+fpDuwkNa8Mc4al+ldH6NSmdf2fHSLOfKPDDuSLU4F5Er4kdI+77LUsleaLPqzn4xOvTd
VLR4wPURkN/A/g/jrdgFqyvTE8q/gQAJhklVbxCkw5ECWmT+KhWsuRZrxTgvpZpN4dzrs6ohL7ff
VqAgHF8HLx5O6V5BrV8DUqDL81sXT12bkQ9jZUdAAqF86616MhQglCTDzQt4LCV5vg7Bx+h6dKFp
alrD3m3/YmOkyqyLnmnRf4ejqrJejnJ0B8LLtBPM/ascYXN1MHQ0Xylm8DmIsXCQ/DijSGGSl33U
22pyGYnajaXNo3wUI1Wa9Xw6TuOzUVFVoEm+/kxX4Yvy9XWuwdQW9/CygIm6Z60FADMgyc909pFs
hYrgTKJR4sCxoDGiMP5+dNauflm+9EQUUXktAIMiTmhrON61F3kVJdTSnGWkIct36Z4vPXUpM2IJ
36/O2Wyo526cKoWSNrXVsOxd48Zs5eAasZ9W1uawEq0vFT6p6RmYduL3W7m0j+MXKdRlDpQfYHUu
wkS1cNSX/Z/1xP2pNdiF8g5OG6lV0T6Hnah8D2r2KU721asBka409CRGG6UWID0cASjuS1uyBwGJ
tVIgaRUwBWbeGDifH7IfolV0pgKyJyMAni+cCJRCoNYJpTiszPAYV52o4Bm1XbB/xHjmWyTt59QN
a+JbTdXq2De3rQT1twj6dNeij9FWtqM3Ia3PT/LLySzrGcVDfYeftA+hnGpketNYWIb1toOkP8wn
gqOByzpmOpdzgIejyEihqw3qVKZpGwEd5tNRkNJhLp6qqOIH8fJoDd+6V9x14jKryp3eiHbQJ9/2
g8vj62g0d/jm18PIgATb58Nqqc4jqRPsw57wu14PoCUClmsyiHplxU72qbJTh4PsXZ5g2VxrA2bM
tvaupla76xJg+AwBO7RpgBgincurHbwlHUzeLw+BpnSkq8+MdN5+EmXA2q2A2dZ1x4CS6g21+6J/
ZrsAdB6Od8jl436ACkx/aFZ06Ep414ArEvX1ckRYU6Lq0n4jOijjup3hy8GvUHFfBJD7d7jpTARf
81quV5vtUXNW1OZWecz0dcZKkMLl0yrHbky+koSKt55Q46zqN1a/bSLwcJDXkHf4nwj7reHK6I29
/S4eVdqwUAzD7HV+BWxHOdGjOgYQL70w2a6EjBiMnKsGW4C3S4IV91Ao2Giemupb3gMeADX2hjQ1
5IUKtNNID3vkYnVXxWJ3MLroD+2KRc0jdgWEHyUEo+LfYcKWtGJzQQPXkX2Ldf9VYeoNTnutEVhG
iiWTVbyUxyFxjJ0/RQ/cPiK9QiSb+WcifoXQXR7erSIZ9ULYYdZrkFKC/4PNF4dFNnlPXYV1W8Ig
cM7K7nSMrmjNGBCynsVRkXSkB7o6eETzAruR0Y1F5vIFKh6JROQsp4J8cGM47Y7xfYwy8UmXGlG1
fN+2BW8uLGDiAnFDWHJ8DDUBMDFOrPBezRM/NENJCU3xvrArxSqM5TXsMZG2TsSnqp5Ju5DocgQk
+1SH58bHR8C1HimndonNPtFVCnW9EFXcuLVe95voabVQxc9kdv45RcN/8jKHDdj7hMr12YdzgGFS
2Yk3oyD5MIvPJTQ3EOh+lOBHzp1k9uMNcmEoLwHBu4ZiohmRn9SrW690WwQ1C3c623N5ijAVAzpH
C4J6f1DhGwbHntDFwxfecOpnpWlMHoh5B3VQMgzlDTELsuDuySA7qxjQDGiAYeOF4s0LlDXFYybd
bywbrNUcYdnzL884lfjBpv81XVBfLtrpZkPJuzUA5TDynw3+dmE4HdvoYO+JZ2aqTLIHiTwIN/pO
Xs8kj8r+9BFH5qr5gTnZkpY5uOkdONuKFK/7IrqhA+jbxzeYcrzxHiNXh9jhUdw6f4j6xwZR4VwN
Ag4N5uWFWTZQftOsOJ6hRuOuM7FT+h49/tbAVWI//AgcjrHCBFxLLFL97LYqWw6XaDpnrhSkQx67
8K3NR+DKCUYIHv9bvGe9EL1ICbU6hw/69TeCwL0AsIszlZo90jm1a4nVVrOWO5UT+il+2Au/9cgY
T7V3GKYZVnW6ZDqr56Ffp63UWV1qTZcU6oZtb7Sir9d7oAjaos6euCKzx2HT5eqQyDFmYP9h4DMY
SH2AHAeiVc+WmW82e4mn6kSkWarHidfZlfF+g0DqsNkBu/mtAjM0pN+VlvVmtLVUKjTL7mSMgspi
NcDfQbRS5yHgGodhC9dFqB7CM/xbRiK5L1hqKg3LX80C7QalHsH4MZqaB5GU6MwuNgVwowEwG8pW
VU4gh+IuozbRm3i3mpD5EvIdttGFCvCr8kyAQXVnpN/lpL8dFKgHxRcKwmhvgasrQLBusPlCGI4r
CioPkFdC7I3yxa5SdKD0qvhFGS2xAnYHZ6mwe/mFuRKPgNasRZMVMr/x9qAHryrOVSVCLDQeiy85
8A/7O0uPos7XOPOrgPZ7Ls5wDE2YJM0w367i7go3BRVlsBVVvFIIdrVKQs8kzb2v8/OWwVEsqWWv
8r5wsMmrpDkW0kPtFOxtP286/Fs0hQvdpcZQSQLQbuaCfVQvfyuPdEgYaaZdXtyYqinqV1QbOSAy
jSImiSBp74mAjn5SxC5Um2mjZitEJ1nzBVTKPwnpAdxiw6VPrAupwrfpJ2r0cZbKEdpjADwMPinW
lLH7Ty2QvJ/5nfPd7ObaKw+TVD/2UXXYgqNGlpwWrlxr2zbrhcaTBo+vq3HyxGGFlbm8eE25rTTY
BRjxXcliN9N9RajC6uiGgrl68V1xEtAlbrUm0Mc8fXcp0rCnja2ElGNFhEX86iLfJAdd9YsPMcUx
9EczB0Vpwo1geIysC8GDDXhEjOMFpse9TeaTrCVNK22vheCo+OF+QTSmxag7js2b9y5mIiunFvpQ
SIqnNnYsT6qijYorVmHfH6Yk4Vo1XxoTWncgL6fPQOQGFr5yCFnliNM5xGBkVDTtRcUko4kkOY33
HobMZ/+U9cuncyfqCd1boPF5/wJ30GwJnjAumNPhZolZ5hsXBuAlnpcRbeaXNKVIGuAmmNuzjgnm
3zh5uysof7Wn/XOV9djU96nT0TCBhuuNaXIErrYY/1of1deozCrGoIlF1zpVjsO3908pmNuoczxF
gsNbNbswW6gcd3P9Tsg0y0SYOwEBL7aLYX9i6a88ic/DZ7L7YiwiC33+PRR3b2jcGYOOAQrP4CmW
YrRSZdFZvtWyZ/V6v3We+rId8blSOmX8QZq8V6CiOB734ofk+hRL+mISEGXyqIBxAyAwsojtWQPc
qSd93mZvITwFADWHKFCL9kzrr8potYKmHQN98JUZrDObbkuQqM2D7z2NPwLYM412WF9VpvCzaXEV
mYF24pXKSYDHm5/+v5QGYRljOsxu3GJu0e9AwjFukUO3PuJ6bMTDHs57FgiTNWMjIdvgLaDscJ38
PqD8l8ffG9QSpfLZhd2EuvEpMjLQCrNg6WTBS8S09oO5RbtK+gguXc8BFPluW6FBURtvUXYEBMlD
kM8hCo2nrcoc8L5f4aomJE31VDosziDDsZqwvov5ygBvsphkpAeJeHqzHs1f8guUi0iEOUGmeHLv
TbjPygFadYk8pA8wh8bEK/YFrADE2f7Wn2jxFItR56lsyBDx2X9F029qPPXctMGsc9Pp27Ywa8xi
lZh+O6TtSsvqY3edS7oxUZf97qZe09hofoXMykq2fKj71EkYcJ24HlPqXs+xCwPqKeV4FF6qg8U2
PqGboWOIyrPmZpKpAOEhdeQfTY9QE1OELD0Ff/SG/baLavwrBvXBzb+6VRUhiru8mGjmJObJtFOB
wExadIgVMafy68uMOWVZCSD8tbmjpqnNXaNtbaTjE4efOMIxEb67jMdJ09ciugNOgSJRz+ubxRQ5
52qeFOuL+jO3+BOe3RV1moNzX102DBq4KOKy+txTjO8Wmt9yWVXQ3xgFmaPCfC26QbNZgm5V6wJC
ywxqcqrxm/pIXxcPkKbpIXhY7Ai0JsATQPuAmTXiVp5DxnLHdlxYfm5wNS6BtESsNu29jYRbFOvR
pBGIvGJ+KZ74bDHJ+ngTStmY7c4G3MgkciJbErOUfZVdXzPqCYRNCKPlZfH3sZEv5FHFJSR2eJo7
9O7Sakyl+DwHcE7lDmJwAFxN8l4XmZtq4SKdQkPQYwRiN/aQVqIUAUrPAGdeWSdPGd15vbv9JWUf
i5v6T2Bpz2fb3Pud4JI7yN6c7vcd+blYXTNQX2fMoCaZ1nv0g2wgGXpQJLCeQnsDOw/5kmnBSsG9
DZ8wWbNyJCi00LRA6Io3Ymx1nv7T1LWe7wFyaaFX3pWyoqRiqMIHgkS+0Cli92KMIQjaUnHdiHnU
ICnHoXmOW6oGO3EVblAmOi63if5I5ajbr9ledK2dwUYJ13sJCXJYTEGuP8VxHfBTJRFilhJXmetP
7dfks5gG+H2qv9iAmfCgsoYjs74/uX7ti2u2071yNzRi/5HhipdgQDkX2BawO5VP7iZrcPCUAGqv
/GGryyKQCoUnoAozibP6kxPafoDMVJ3EqOYBl4EuYW0mqV8dz4OFY40xMSaH5qUz40Set7VSGr7o
F3imm2ELP58kXHffHzIrBJ10lRRbTQqUqwfN5cV+GKdxDoMzVYZoYKodBThfpuanpLCHPNWUNjJU
I4MG9bNNwYPwsEmG5ba4QM+Z20mhWjlvh1X+/Np0GJ2BU5IXxttMfma/IBbAMmOXM5xm8/lrfc3X
MzU9YfiWP3kvSKZlzorYJ1/lXqcCKt6NF87i9GEX3mIAwScJ49T6aXlZXd5vN2JW+seY6jrv0aAk
UsIZQSt2bBdYxAwIQ/Xx6HkOuW+DGDnjPSHd1WjOEDjCtZfZa1xh0gWK0a0NAR0KQZrvNqFZqK1F
sa586i8sqzd0BdPSoWp0dUwDQ6VeuotVwUmUSQD9GZc2PrKFAUHCLdXNyfItxCqP+tmo/q9R1qIM
pZGi3rgToGDaLbVjdcL9G5qzmAujLx0z/5rTScEncAtAd+uEvU8Y4+svkBVAFPfsWoJ1hEykOfgE
iLmxhNa1vt0wzAJPPaD7wdfhOJirSf3LryCvyc5ZoldQlP+DSPpq9gdudXYpIm4jHXdR5w8CtmWP
VcE7/Jinyr92hqIfpBLLeS0TlG9YrBwG8NLgq1ZfIWvk1zmlmQQPF7sqO0jnceXf/+sIxrjnXyth
FEOfZIuqULdfoFamFYp8O6PxZhEt3vOCy0NrOaGj+mwe3n81qiuhW01uUL2L/nhC2v6cPHwlX4Pv
TkUtSyA3cRTUtvZ7qZvrOySr1igY28WtTOYct+QNqhwM8mURgm9XmgDDiMGqRZJliceAlhvc0Pcc
ClzGC19JxwA+P7dBiF0/1lKPzKfgGkPxNrcbUP1piYHVlDh+Da/TfY39MBqqMtPskGmd9T6aXKzG
aYEStYF56qcfjlyIR3WRE6WNdeFvhiRkrbpjUwkx/3TUerutz/osN+qZ1G+WfUZmyvk9mqVP8xqw
C0rrqEloTneAS1fvn1VBjOeLPLazIxuzblXGEWuK/uliNBwn1nXHsGNTBXkmeLQXB9w2OslR2oHJ
gvqKTuIYyzZfmCw3pL+9EU4ySy28BBkUgJAWE9umZkKmXlPkA8y9UiWm28chd8ZSVrOhebuHAUW/
qXAbrXoAl3/XWtrAf9KIs3bmSV5q8VK3zStxrQSZPmX176YQWoccB6AtNKjktdoNXPjJcWofiREv
0MdobmpwfQ6iBYhQ2uwSntBJtqpt4lPuhTspNMz60FlcBZloV6xbELdKo7HT0mW+rhuX4W864sFj
w9o+TnvMfG6ED21LVnw3Z9ovV6WwMrpnNYWlMunfCXd9+uRaw7vSF2hU4RhoTc2mLVVCkVduJnQf
X/P9FdfJTQXil1O0qpB5Q122bWY8e1fDiCkjOd2XGe++W7TWoH0QSg8K903TxnTLnYw0ljxUcp//
d/IO+uIWYUg9HWdowgxkC3wwYrI9qDOg+k0PuuYS4HGxyyeYFv4AVkIDK5gsPo10rEOOt9mIWAWq
pm0cui4f3AdMQ/K0aRVJHzOt6UfHzyqGJdYyt/65rloPAULKHH+/sSedJkzidjue6wZn1nxclcy/
hJ8I7xRdrDzTZy/9FwV+6HuyKq8fg8iRbdEnGRwsscDO74We1uYBoB0ys7f+IxtbYu8EeDXn0L4q
Y41feFhyyyfbMLGHLxH6uLCOlBCU9A7DyWaBERvQS+eon689CdfKlEz0LJfAo12hYlFverDIUaHt
HnKj/C2jDkSot6zL6FwUO5vSmz1bAMhamT/w05GxuaVi9Ii608DFBVDfjGM7AJnkrWgqUH14AZBf
KC8d93pdGeK+E8VwHViDXf1KPaC6pUQsbYErLMFA0WZ/NEaX/EVZflTe0v/rBYKsJkFVDE7clThi
62Zi2nCLqoN4NONKy/kQk34ZjACCL4X+qckE3HPZOz1E32l+Qpcm8Wpl9a9Diud0D7JNmAPkWEeo
+ZrC/lsvW+WLKBTK6FfqZqzlJr/5+J45uzVWxH2Nn5A7V66to6uLYlFurAICJp/FSUnxeLp9+wRG
Alj4RltjUWfQkxI+ocUZgFUe/PJdQqeZ8XvYE5sIxMsHRcsUUWMUBWVYiOZUl8Vb2K+gvmlRua6F
ZprubeqWg5z6zxW7N7ov39CGR8s2sznNLnUufqqzZn9g/ud6u6UlTVER/PyfVe5iVlUOpjy2ECOQ
PU3CLrcJA4hYD2v7ybem2jKXiIsUjPNfFS8pCaSK7IO8hz44yTU6KGNBDyNmVB6g7JAxqD5VmR6v
CVI1Vc/RvSpKfhllSlJByPIIrQhKe+LraTTS7tSwUG02bNF9ocyxUi+q70wdc4VnQva6/02n/CKn
itnHSiWDc6z9ObmmF/CudDkiplQxCWh9br1ygtZ4TrdgNczxK2siRi9in/s/nCyJi/d6tfzy0H4s
ugkebzZkF132OxeARXEg7ONFZSX6b5qcmbQINynoA8IyTUnZKgHqPlJJ1fTFpyqYdGnAbgUJ7xhI
eZ6tZyHRBWr6hLMCapfTb3Ltgf0opsBE51yqZQVMl6ahqcfCFT+c81cj52AGnqnp1WHdZyQ+vtkh
r/fZIboFx1VeGfOZy+QhIzlvV9X6fo0V5eMhB7nJ2IZaGfE/BY0ooSlib0k5EH2rGJg9pAOHiIwT
+sNCnP1JGQsCIKM6gvQXZ/nsy6gX1b7aZ/e32KIRhxm3LmyLPjoaiyj4KXe1RZpVpUBXx/hXRIJQ
ss9xubvqWu+RoBhrdE2pl0I6wy/5e3643KmS0lHu12KIE+PTnIEqWAt9GayLElqcbMC64j9UlpX3
ULZAKQlWrns499JuRVJBj7hJCyfnODR5P60K3JnCC9VJStMEgmGrTiRXFdBIkUDdjptQAkONjUfp
PH3KBlPlgE0d63omNUJB0BgcS0mH71xpLlLD3/SXqgFCJKQxEH2khigFo5nUmWCmADm7K/1VNGep
HZnoO1pt9UE9oYWnVMxuuqV8bKFXvZauKEFRtpZ3KTDOYalFOipAodGJ/RMaUbUGpxaZq8hx4s26
SZ6nT6eWTPq3TDRybnjHxTq5DwWAxiabqDxmp5JdAFSvPsb2EMRpcekNaK8rMxVCmQsiJkyEo2MB
TK6ktXMRGVXFo6tGIEBt/yrcorwX9RK/nPD1q89/fSBxiAoWWSPmBsmyWfm7VCX5p+CfQLaphHi0
yb3ccsUYmUStCQeIKajjlPLGHeZYIMMfdecensFlWcmjOVobZow06yjPmEoGYl2naDs4pydVuL0u
V42EBwEX0KoTLYVZdZs0LdZ4FKN+RjxWLFXVvFx4pwzCwZhz5nEHZNFGQMOIifZhz6DQ0cWEnxEZ
Fx/O/ADUn0oA4p8PZ5zvA57S5uvaWH/azpgr66qq4bLFX+ppbk/qlcfDHSGNkW4JjlGSoUi6mSU7
SQs+tCz8ZbewBMUcU6MQhyKnLggimSm1pVRds8w8oavhTDHds03Mu3a07kxnFzOIhle73HoaWmZv
OP8WQhA85+50iHc4tUyb9W76H9SMi42YXIDJda5DWEe80hyIlnOvLQI2o5/OToL0+ELc4rx4tdzF
3XWqfhTcDEBlHUSqDSLehs23jWwhzAqYRj7TU3PFTv8bvN6CxrKtwKzojfTveZPTSmYkWa74NBrP
KcMSox7JAMzG1XGc5Q4F8kIHuxpLBXONCh0JiFzXdTWiV3nO8wrb/vluRa534WXYK5kjLrPOpMDA
1vSi1gQogi1Jtuz1uxTkoVNZfGOX9FcxisssBBvr4u5ydVGSlu78yBAkiih5jWYgw7+iEE8QF9/P
xprWeCWfoS9/L5EoZAbU4GjdTvCcUiaOUQqqjsj8foMbHQFwql1o9MVYzxMKyxvZC4LPgI1+2ZSN
39Zax6/YyDQRlboDhIbyziVsx2ydzt9SBNAIm1PnbTnSSIM0Gq4BMj6u/uSAVTFjDpQXTIZjR7dU
hpQZ51iWW/5dvHVRx8FUs/wsb6WDzSYVS0jCdhHrNgC307RJuxW3s6O385Z4U0zsTqq60WWGfW/E
CrwP0uQgjypP2Mr/z0JEGR2SFDJR7yIM58yrds1eSen8POEQJ1o+53Q5IoK1B+du/oI/8bp8yOgZ
ePFHesNhaqvHbE5MlkUPH3e1NV8NMiVIEcsUNbICXnBtx+egywfhgOiCMZ1kdk0c/6LTTMyGUMXc
jQzhBhR3KNN5ZCYVpRMJIWBT1NWSplwGg9r+qeDC/jJCWUO8qQKkkDIsTLuWioIh9Fbiy4WOAl9a
1Bld+zGFNKJ3LkuzXQEojNyVgSrt38RYcmFWbfcPgGq2AiVe6WxqnTUTY0WgPcIjMKy/YvxNRuBJ
zj5KN+dllu3pbScJ156r+5Y47RsISe45cyFsQAOxrUqD1BTOhRXY/DhYlzguFnW2molHxHsMKq/t
tNSHN2kbb7oKK+/FUCdDISt67QYHUUJt/k1vsO0KRkVH54N2tEIjydvwEu9z/HHXmaiI0dhfXn4F
bZUYc7M2+pFhFCUr2U5/TZ5+hL63Q7YtpugO/9wOUbRTyQQDq5sNr7v25TL0Gd3oVJIv+gh8WjPn
e3Xk3psZ/e8oEsC1neP+lmROJFdnbvHMljxLR/zVDar/RGtotoPfdmIFDxIH3aFumZVXnz3OciH4
ELX81KkG8MGh1JoB3rgmR3Ai6KQdiUT7j8vB8ihxpHh0ku8zUxo24tSOKItYZ5VRzZO3Z2ZHBNy1
gzCKyZGL0Z0xxNP7pGsfTrNAw72WsyNoGNM7lhN92emmaPAOQxCWvNdWpiyDIs9r2x3NxwqNeQFq
+k4hVQJ3NGztMNyAEmHvwGxhpaCIaUgf2vQgzleLHG+Mtceyyd1RNvmgX/7H/JoYRgTH7kXcbk+t
cHzNE591GkQB/g3MwMtK82S5IJSCCCr7scDAX2ztb628drdK6JfUEpJSUr9WyzX4J8H858qQo/hb
pWvAlomSIt2VzBumsKxPIIwqLf7PBLb5K909hTCdDeHnp0LQ7jToC2Ritry350iw6nOdARNM+vcc
C5hSM/dbOELul33uYA6YNU4VQWv/YsQXE1nKvU67jKjGEbUvF/IWTDSqxeGFAChbD5NUzMf5cek8
P/QUVN8LQDtNBwP5Kkz2v8gpigyvdiWd1J+YeYtmQT+MgmjyYqderUpvbiGho6AYIhqJQHbOPTKa
b9CanrF9NttCJqmy7kkCfuzGO04sHdtXrihgz2dR7on0HW7QHz2ONQGbIHVRfJkFIkaIZW32AuGP
JGn/t/fuif+619aOMicUk9330OsQ6/37c3eYTgT0O8oHrE8zWjIDwrmBtm4PbkgMEF5D/FGMRjkz
Ldei6XqNc4MZdAhORBVqD4NUZ4w5DWVzxKHyy/9eKbvMsNEPu5uwdJECjIydMlWXpjyXIR3AmcGr
nKPn2Q3niJS49O4TEQKZH7rc5eg+CqP2spFDJnV6UNW7wotAb11SaROsobyc23db5FM+6LL6jHTb
GTiRJZ5CWxxjgTw82kcl5Tc8/7i2QwIIplJN+whXq9J75408I7xSXrrJYtOcTKs4FarhmCbKmtrP
gzN6SpHLyUogziE98KwbBwmd1g6S50A59FwGlPOL5xOKLPJB9A4Jw5xbGT6RNEyQQ75JAPveVgfF
ofc5ofLnZ/Vei6Qb/wK6Mz6d5Jo7+zwU8XXaxadxlipVYiqKi3ER7QwPikwK/yO/RspcLi0lS2Jo
9TwIUHVYTaaYsK8pvnWcbNp32Qs9hxzvtMR+gmNPatlN2AYwHKJGuLoU3ANnQESbiCJq0F0563/4
Tb96NazjC46DlIe/phAl0oRrEgft1ycLEOAxHi6jOi63PIxxZoWf+Vx3rKhCNahchuPVVQFSwNlo
PTDA7XvnPNTtPqaX3LOT7fDCSq4a5btAwY0zKSqQdbkyi9net5W1TWmq4MiM1LPg8I+GekmPs2zP
mM42Swu881NViBIpokkT4b7k5hccHzPGelyXEcUzNOWsJOD4stMnMCo69QSg8eDIIiIOf7aSRTB2
2Uy8g8KwfrcEaq5lSHRxIvp1aTp+s6aq0BX4lA+2mfwLn2zuayKn51t0Bv2FNdubHICuGmCrj6Gn
lMfwiKZT3ZFcxzV8lnTTmZxBAsuvbCECULQGSxLPp2HcOuKenSAUpLAoH/SxmcRXHCJAU9g13xba
VOosXPa1NCprsPRl3KfTqhTZffVOibZ7Unqa97VcCRIDCvIVfcqNi6DpObhdkVsxk71L9KZW3YQ4
3J+MpWAwuJnOe3s0XeClWPJdFTC7fK1shMbJlWsPjN2QDi79GoVj+hNLMtsyy2ixjM/r0fT58V0G
htk2cOt9r/A3jGRDJ5CsYeiYoXfCJHx/K1WdDDp6S6pNgMMLunj6IpupZpjpaIilWIghfU+26Otm
Ww1AXuxJQMbKGLoRagdvkMbboPVxkk9lDC4I9hdhk0h+j8W1EFfliuiQgA67mc+3UDC4RHtbYuoU
G1NpDyfQNPpHlAJg7b+P7Nq2omH/uaAu8fFCMLa4g2Rn87l8JH456Mp0CgAAb0aTWddBpLWz0Yuf
wrTUFMRjMQCmv/2JO2yQb/zAHoddDOYGf4RAOfBEjBKiYgN2WVxaaRFwyCF7n11reiNm5lpK+yWo
HbPIppc/f4cCBjTEGKLoonmPkiV+kT0GiASq75Dvjbq3SPtT+O85mu6H7fVkl8eCBPQnXnbuyUsL
iF+Rprhl5xrsutImknJcD7f4SE75/z7TUTLYPYy26d4vDK9c7cnmjzyHbUJ+gJVGzFKmedZfrtpB
0fLZalBAt0UXR5RlH8pSrJi84iuv0cJC/xuCw39SL02IlRen51MWPh3iKZelwFTtEGPwGbiV4N9T
79FMAj5dUJpFTl4L8Awph87rZPhgyW+pl7rXy8eunIDpws69e6337E3RL9gW+Lyzw0MAaDPIljUq
rciQP2ufxEkqRw/uBHtbWz88+nPFH5BbNaOk/r28VcAdMye5CVxbK1u41hoVn8ncRf6NUQMafRGo
N8uyIllGTZP809uFEkf57d7vIsrQJiZtv3+Z3781tMbQJq37Z67vqfznnPeRtAOUYPAB6jeKBerA
Rmv+de3l+5c5vw+nWQ/EoCUs12H2LxTCNggzJEi8SapSj+lTOVKurvvHIvLX6hdHRnlkP5gpgz/X
Dx1o8IFLI+ycXrMZMju82KEw+9AxikD0nzhoPy7F6jV7DI8PuBOhEIknSLdm5vhX7D7tXdXWzmkR
0qE2MGDY71H1FwZ/rU7aBHFHt6Cz/flsf3WyY7xPKiliSFWWjVaRJUXT56XY1EFfpHHXCH+DksxG
NnMKis0lnYS7PQZ2bULYXFI7yFF9S01FkvSW58cSLnVtwIwpjycyOfVO2QQvfyyDW5gjLSMCPqN7
TVCZxQJUx7J47lsH5XkJuegydrRfKhzCosFioJMzZT5cxQVczH5ggmYQCDaeCgye8+FO3B+gd9FT
QqY27Dx+bESoQF1Hn4tfQFFEBuMDF6MaT0C2Y58WDP2P+YlHK7MviOGFbLKTZMzxNw/iXrP50Twn
UcwOTRbiCQ0sziPZCfim/hfksXHbmqKbBZ/5yLH+S8A64OzHTAxscAJ5YI01sOQlx1847k/+Ql8H
y6aAcjBaAFWYs6l8se78767Z9MjeHgyEhfzpczXTXNvkyuk/jq1B8isnm4bLcytERuGDzEi4aMWC
cr0criM3jLnKJAKBRUHQ4lFdXv9ydsR42DQEGF8TBjz0LTRDEXBKgWH/dtnq66ZqjfHPwLWMsUzK
71jAtF8rGM9kRbYQ8BjvczHD1Nk+nAOzNaYi81RfeRMJn34ADTPCu0ZaeTPMnPfnZXjHK4dlD1+t
hh2PmreKuMz6WBOfjH9WpLG45rR1+lcLZZzdeHxk2FXOSNEMkHlIBkFbP0bcFnZRcmEms3l8PYlV
/N1cmd/WRxYxu3W3g+fiTEE0TKc1p1evxIQpz7jLlD3OHlkbe01qkGfVMC29xE2IEGPRmche4Xnm
FfEnEVYwaOnYK1SXiE2HTdJYmrUKq9Y+i//lVSJ0M79EGN9g7zhZKmgfjJaL6GBYymm9UpY83YgE
1i7pJ6LeZdoyIm6VcGX9M4P128sW17c1TvUHm8H5IZN3U49savyihk0P0yHqvQH1l5Cz4xaqX9fU
pXlDcc3mbmxlfWZ2SR4jSbi2TvpTTymIba9SMOmm0tqmf/Bv+IHdcuf0lvr5aV7DxfR6lv6WS+sY
BTYxV1ltujI6tbHG/lwvKEv0yoxSTSQP3rGgyUgXOwGWcrEIt9QyiyCC9dzACuBbIx2AYYRQalWm
7papswd6kCOcR7LPLc+elT0tc9AyBvi/AwzJcId7FkqTC4lgzbibAS0sbuN6zwwAWyzMByL/r+5M
NBhKUNa0K9mBfQFz727WhuMKAjqMB3n27cFOBLfUwAWTmE4qsi0rgn+hQQb3Qpn1r/uqzJWaPciv
/iubSaGw3LYRAJWE+ZOnfAP8TVUUhqsEsg7VPz04qwK0C7Th9KRGCX0KLq0eHGk68WKy0o4mrCgG
k/Fa6+R/ooPV2myf7TvJysQK7gBs6w3BVv5bSebjypdJ5fw0qi3yUGVBmNMAOyja08XZQbddcYe+
4/Um4YYeAV05CbgzsEAuJNcl4Ae+bnB26OPsHqd9iCyk+xWzOgkEF93QYoDlgAJUO4UoxP41nYpx
l2B9Xibv6ibcgk4gYzSpa9R1rCtocDsZxXd6OWbayZqTlCXyOYeu+BfdCuKjPqpswNruSGFanDl2
47qWz/W51a1Zv3UbaS5RHQpEco1kpAN9p7mHSCMc2vVRCHHaa4PIcGhNrcnuiJfMP2EpHp4Nuh4M
nCKEBy9dleU01OMPemUkaTRV4bFTh2QiuJjf8wRaz4ueq67mSJHzBb4EfyjJsQ4EBhENLiuhRism
fOP9Hre77eyFg+50xZjf0oShFIftBkMjjVJJwLtSbOtcvfeAi9vkd+6XOI51Bo9bA4YyJH5yRC+6
bOizrkqt9GJHo70ywaaNz8mA6hDv5yAdB3cPMZesMuo13+amyvg09qkj5OzzMmUj4iId6zAWSXQk
o6rulsdfP+yLbdnZYyl2xnh3nm6dKYeINzxwGqWwFcCbshJNLLkFdCMHZbz1AAOAIR7onykmqVEA
+Y7xxHrtCA1iyDCGpoXSAYOTwCKO2hDf2Bnm1R0xAth93TVjPE1HbjZJQEoO6BkQVCwwMCgIMvpt
uLklEIjFElSkgUPZi4vHX1l0FQjkeYTJZkeFm2WnouD5bV59tdANBjUYcJjivKV6xWlrIizSV1Qf
G4ysomOnOpNH7C02dRp+GyttOy1eLxUfqtPwkZjqjkvpK9FPZChHGwb5GAJRGJQywHalxanw3JFq
J7t7OJ+YisEVzluexReyScHI6UB3mwdf7tRsTFqEB/IeLZQsGKBjLpignJPEh163RZZdf2SqIsue
3i6cydJlXNRYRUkMGPr1AZzOjipDr0sYyAr7MguEdEDAgCRzQciCvKUxVRmNqav/dNM8dRaVr43C
fFVofjIRwCQ6I/sqrY54AOWy9Z5w7ieNg31HOmhh287QU5MQ8v13tU671zwCGwnZn5hiBaNoyaJ+
Y7gLdiI1IrPNhdBaTT0jeM+xn3EE1DLYU8xfQdMU0ThOJMC6TQWutKU5zOYGwd6HUiz6prSOIYww
fsvCjWWQqhdZCOySl0/y7s0E4iYkThDeoaTSymVvixSSmoZ5FzM3kltGwFugoHySF/0EnXh2pEfi
oE9MNH9WM8RyY5T6lHw4CNxGkn6PDizKuFAybb8ELuBsZ5oS/xJ526yVlf+iLv0UDG8tuqcds3AP
HGjJG4ntokPRsEcjOoICftg8svseR5SJOi1UTNVz76xhpqPbi3tp+F3s7ScD6ML0L2aZzvgO1psJ
wCwzDWSA1ADgz+tE3fdduN/wrOi8qOkJy9oQlec9wzRkhZcuQKpKxVlQv9/dn4ReFtz5i+ZFrEXR
4UI7plyIRUIgIJ/rNEuYUwU6X8TVspT2/7E84ZzyuG/a5Xmns8kEbd7I5mdpDjvOCLldTvyidnik
IBghPM8UlcSfpgqntshji21eQkzKH/hMQptn8Tq2bqriz5ps0xo0d6iAsK/M8Hr69Pm5DP99webV
fYUJHKJWoeWBBj3pjimG+jt5BLzMUDXiJ/0UexXdboxN2qeC4sM/AbxMa1CjNRxzK5bjpBSKcg9i
nPGTeQ0oHiAHVtsawZmShVyPlMebAGkXKaTaxy9E/h87HqQRO1XMSEOiq/L3ZQ1J2A0txv/Bt/Wx
68rmEEgYfeZNc7ea3rwQ6ryYs0h0bL0D4DOKISEDh0aI0UgOMbVMPZmxAWLvGHUjczyBeKQm+h+z
BaVHjprOSGi0FY47pJdDKzsFjxCNiP7+O0cTMitUNEBoiZ7RHMzwhbXr5mKGVg6LXVed9ewAmCSq
pLNZeioKthKVwyavJ1mirBgAcOW3xvTYsBDUZ7pGZYoXgmSQ9vuouyC/zHM2qhObxp2QiX1xSh5T
9m47ytG0w+pvbAr0KKqHPDfcAJU90amtiIvWLY+1QyuYM3ao+KSnufQ6ZMiExjGM5EtPPFAiQkaQ
8CQHLBzCphfNPX1GrtAvsqLOp/vRepSsLG5onjqxFWZRAbWx1OXU+g1QuJtuxqNF8JkZs6KtylAo
WVNvsitxCNSBOpb3hTqu9k8vT/pWGsAMXTuqSK949adNgUWipfAFe8BCKljcnNx9PLs3ahctmZWl
mfdhQUlTo7lv64yADieZhlOX5APwXesua0Ko+V6cICO0Klr2hkG9MDy1ds7ZYPsIWCei7tiopyve
hD6OTw+0SOAtg3i4LyfCRrgeeXKDypkOJlpfD7dxPHUA60Ftj04S2eW57LvCi5mIzinwSTyFNwJe
zHGQ/hWJ0anqhPAVE9m2xhLAgVKjQ77nlcY4/F6jPwOGACqSmATbTBC6fVq0BgVJpOXQtJCUBKTI
9NrxL3I6IP1tqoIHcNJ2f4ZX2kIK0XQrOTT+yMDMmkUNcouC2x4w0GoBjnUH2eLGIrH9ELd1KHCB
WMlmSEKK074VJTQ8BschgbVrmFOX0sDauWmHLp47KwyUw9dnysxvnA1KoX0JUnaGYFv88J1uWdfE
vwIhjurILRdoVg8+ttCFUPPg1yMgYULKayTZ1ql38h/nZK2fIjlNajwUVidoogqw0WkRkeyDO5QH
suvOgXXtQ6cGwxYs8xXWEMAkCscCQ8022rVA4A+guke5cuknyftS9W/mIF7FID4DWJXYJHkZ7KkT
Ys6Qx8dQJzO3hsfyU+UvLLV4SkiNcx2Z9TCn45uYdFjCgLacfxOFY7c25IGsYmhlfUSTuiufthLU
OlKePZmwwiWsxrbqYmIThMwPV2zw3QvgUmIKqtPAZD9W+nFsMWckoST9n4SfSfMlYtnaL0JQRdrx
k8lzMVOoW7GaIG3Wd7de6VUZ1pVGFRHKnV2EF3IRf/nnCLGaEewDoNeR1iSBeuCjak0RMZXBOYAi
U2UJe9K7LtxngYuq40zb0qYkHLQUXUJJ/zo0ckVlGBmxKd2CuxXTLxkPADK1nfmxzrFomJsyj/S+
5+mMK3NSJo9tksuc0pInvY0Gm1Nd1uWKArgAcLHkt5E5+dY0BqzgtoI+WLtVIwfICrwPBx8+bwCw
Bww/zzZnwSSOrK0+ktcdceinC/APxnmgn86wrthE6p9a68cpadyNr48lbteiuWokpFQvSycOWLRi
dPetsb92mrYuMzMXHUWIhXI5a/7SY7RAfULWeyFk6n/oZaN3f5COgNyEprdfqCvKNxPUm6bEiosS
32lAnftyZL7x2a3pXerIJm/bGQGtAvOpBoGOpy4lZVn+QH/aiDWp3VjRIJbBCXH3VOO6bX/UCkkc
Dd/34kPYckO/kdXhPkQt59MrolgnqqunHw7QUVAWG13KHBZAMaRCwY0JJRw95I2jkhVD/bDRceWO
OMCj7C+k99XCRjDhLUMb5ykfHsBkl9KsMQaBojWTDHA+tU6SM9WbhPMUT5Jj19ZSXpmxc+BYJcxW
Ji9votlnM4u6SWn9e6NQLzSrJdAPJjJQOnesI2w0rh3IkfQ9wc7ViGm0/gn9LwkSzwMh50VjoPil
mccFD7l4OrixqBoFFyL1H+N0wAMWqrlKbK7a5CuccoIOc/5edq518QDPHVbbscs8iTyyQRuS7GFo
9OaMG3lXGr0b0SDmqI4WTwkYRQYMikAY4ML+AlJdGLop9Rhhi/75KDajKOfE30m6FZiaFpkvi745
WGOIWC/mNXJ/K19v/sRUwhKoOzECZDvSMKQ3bLye5acvMbulV7uWitgQa7vXQR8J/MhmQI1pBnBZ
31oM40XcoCoeAv2lMpulERUks1uBOG/N5z0RBa4/2rqhfPFqAV/MUEnhx3irInq0WEY7IydC0EJ+
88tsRhENWCAQegIhI0/0VcDdjv1g7ePYTN+DassVOm0DFaejWEhpACVx++btc6NfyKOa0m703B+Z
yMhR9YzyF8fw2zWO6+xkG+bQgd80f4yxQLgYOF/7qwHhCKAFf7BqgpxSlQ4Wzg6TomO/AlszJBOw
plhaV7/tErFopBIx0i5319tvnmnGfnvj3Zk5HT+q2GWuyKRVwagLDMZl6jaPizrdJfviSAqfqFnN
57g5F4P4/GHD7T6AgnnO9DuSqG2bqy5zTzZy5hnZ/LafPcldPor77N1n6bTy2lA69G8fRGCRk34C
+Uyn+d+ghbpe06E6gwN35ueKbLuq4TlIk7eMMJxdX3Fu+lnCio6jvvQj9EbGuPvSSdePCaG92wo7
7VD8qC7fAcJpF81U1XQdb/n8hOuI6wb1uMWTDkVstQuwJnBBAJhIZhWXQ4OzwGR+mj3vFwfxxuUn
J99Xqnsz09diyHlX3UBZ8YW6ZAqizFdQ3iRu1aQAqgpIV9z/UL9Wa8XoA5+YNAnGpS6NQzkAfNaL
mtFutpl27H/c8VebvQjO5oFnGew4gDsT1h5UarKrub93EslH3JozUV3IzkAChQYwwoutnHWy1Ge3
ZP+cYSU6u4jLCjQredRRMf3w4uDO3YTSSkZweUbC4Qg3kGJsgjYAhSyg6j37XNAt/fPN1Qv/vBNB
c85n6u9Y1Dhck3gWP3flSVjcztjeXMTemEQ3t4Hv69iXDr/qJ0/KtM8d8zenYqfGkOVK8g4tvDvh
a8wqahJavmwgKJpgTid5rJx/vLEcoMzkRHqNzSoAvQjNBj/nI3ldiEBTbjb0Fcg0nMkDsa3jUPE3
WlYcMcrUY3OyViNtZksQd+1zMVPYnOlSwqtM+EWBKwQtGNwbj0t3oQLbr7PKJT8jjog4mye7mwRA
080bSSJLOBcyWrzLgGYhy/FkPkHb748BlImTz6yaWyf3IHnR11xjyUjfYyRt8anhtFw1NyDRK3qd
tKT4+DupmpJXlMtL9V2hTGQkDgCPNQEtuAa4aiks2hjvHP8CE/pqUC+VK4LQZkbnAw2YPoGmNPxF
cxNOnZdSlwRIcmSuuzOpt5Vu3sYewN2EtzUwWYV3hiNKqLwcxnwTZ/eiAuGfeTKOFdEse4jcZsb9
9BryPpXmd5hVk2lWcOgkuMpCdmKDiPfSit8IcyYrXN2nXO5zpFdsYhMtF9SJG8Cz0Q5G5SYFY4I6
MarnHCSn//5hN4SgwKCbsLMUEFgzXL0UlR5SE/sCrhw+2oqjj9z2gbk1Ih/RaPmc6FOHkS+QLM5e
ZPrQCuETKY+32KEF05k+nzwiL4O0VXfwKtlLeBIFtTE7VT7iloxxn8wDICFA6AajUtX0cIU6FX1n
OyyRX/CiIZRVDlMK99ujsC0riUZ9CO6j3C2xd8iLpFpqe+PLzlXNS0+JpFYjlJqHnV4AsxACuHMM
8ICBazy1/6K584thN+edjj7bibcvVOsw9rhZVzVWBdRV1pm4H9o7YFkgcAIfrRC/buemhbT3Iryp
RsmQcexiKZOliEoHZxoMJuOQoi3LfDztZNR3zvUKE6dkMDEq28IRIbM34zFMt9ZpdjcCrYnxsyRL
TkH45dV5Hptx4/fzjcORzRpjmmHA7uak/3jQ+oSjx6b7iwd0oVQ3+WjlPHKD9OdRDxvT0UsCViFx
I70FiZHtIuBVEULRuiLi9N5AagLk6Ef4D3OJ20VmUP+e8TY4A/ag6em3ZEmk/sZHNaD60EwZAYqK
3mPuw715UnN5p9OaYsWkM2MGchZAwkVHdH86lp2CXjebN1UQfcNcxsY15R6pBnuoL6tHLqmKj7Jc
pLfmLT6zZyhs7i4L3/Y3UEzSiUU2XIM8M8vH+ZcPq+VJaaLETtzUphRuHYa9F5kBgzxekq2E0YRO
69tnatUN9b68XqUadeK5A8ZzWQYSUKBj5Je8S54VxKHF5efm9JwYCWYKShDmTFf5GDXPn9gNsGGG
lSdrdhVXCj2bpK9LFKCtjGtEWhJxGFP3CEE7Yl/ihbYYDL+krsdAL5urmjSq0qeaqCdZ7Yi2FW0+
k3ZSh+gU7UU7AsYfImAcRws5TZ+eYrudtbkdJ0aTI4VpcnqujTu5o1JFyczWc75vtQSmWWr7uxNQ
71Hp9o2Rvas0tAJBqAPAlsaN04bc1qdWBpZrXeQN+XHq68v2jAEWHaQmukYR5RiYfGo3Gvg8wUA9
p8Tu8gbuvepr59ab4bZSdj7G1fXAi4VrEIt+7VkKu8pA9jxolbl+ALpLVUlJJzxSdpElXk9FglcE
r7p2LNPMuoR92JaXZ9dfJrgZHF7B0m9CjMt0KEAfN23IRWxhIAe4yOyApxLNNlHq4XMXPRkBoKy0
hMJxqta2dMPpChgFTTphfvk3hRUUJqVRI7/xXmIr45SEmmyleqsqk6wngKAwbMRz5ENybfLs0HAB
db0ltvAHyBt9eC+2RgUDRmJfH/1k6hBbaI7j3LFQHI0Tme43AiArfRTLEdFNmtD3i1GbihjXWOZh
RN83fsEJb9ttZqIVHUBW1iLGnVEtem5ZIA0fqbN+zw27H05aNTTFZkPSdCl9Bd1YIudmM4UUV7lt
mslkD/ECumAhGlxYczwkQxz7n0UlKAD61DeDBRA9RKnIptfFrHvW4XUiI8gzt6Eg/aYPxAzc5Ph4
zHQHP3JcWrM2LIsrI9cPl5s83kTwTq9Rm1e6jNHid/iQcDG6/iYF16/DfUGwYkJKlqCYYuDWDGVG
+MgWoDHMOg5Bhw0uHf3QQkQlQl8203Ok2Q/nO4pZVN68HMmGuOYOoZPLnwOSJcBsOvruLlwfmMP7
6lEX1RH3ldKdyAygMO2Qrh6Xt0rXalLY1xZ7gFec82VobJMaxCZVJQLs/xBJqpsnSmMYPxp6P6bI
GCFe2Wqk6dMluwSUXkQi1pF5BL2TYFeIwiWx04KpdP/3nad0xsKl8hmwXjFWJMv4uhmHFWqpn0UU
ZWrvQ1vt4icwf9OHUpypUlYsJdCfB/A/cp5nmHrWLaYa+aWpF1tOM0YdQlu7FTXmisIYaQJRp0kE
UAbELIjDOGanNIL0NLaZStU3jWysOau/NAhYZo+sG6N63aS3ybGzbRFe2TTCi6wufq/oaMuuWUej
8mZW8i+rhhfg+wlKbirH0bwQ2UXp3nMyHxZM6A6yqDOwdBzoaSj5srYQyxWC0PGabGfqgleI8Xvo
4Om8izqXSlXIxIuw3G8Z5akJd+gcS73Oc3FdJp60/fL6IP1cpjm3rY6ycF5z+WokRviioZxFmxSS
eUfMlLqVhywB5dQs71uLcx+KsbyUqI6MNT1bq6D5NQj3RuwS/B1XcYEcQ9EPzcLbHhSFD5gdR4SL
qvoBRZ1p7oKfRIVQmMQUAhzOJJIvOEHbcUHLPelBhaBP0AEU3dP8aru29f5bPmyytAACPbxW3kM9
Ov8IXLl2dHib55VZ2RuRwT7Tl3a7tkNy1V0qolk8uE83kT8WQ9x6ZytsHZrr+BPkIzx1FO6Vl1gc
EXa3OD6sGWtSSjaxq8hnl5ZKeqHoNIFAfs9Sp71BQNqOOgEklqaOgdbjzSm0xP38n2UHmIMGNv3V
xEcx2f3kY6BzAXD8gJivgH3UdfaFtAN9Vt7ngrzjbVlkk6WhOHrLq0/RwEmSW87zoMR9PCuveX4c
x56pf2FbF8c3xjhfGvLKemjQ4qSyBxKfINBLsfUvTGMAv+rgY7PNegEkLR/epQLmJkt3qEdOdOTy
0CKSVQvRFsdxw7KvERDxW8FOIb/9pUtam0qH/elOdsqJOQhuXuyALuurN+xYEyPsS4fvcFkJyPG5
0TLDeallag238lyNE9ZISF/2N21DixAwlIe1pVcFKy6Q833ozGdJFhfNgChgF0wAcvsvoLjxMYFj
0VcsZf5eJRH+rzyuVL+8xjCgQms83JxBzaNnRF6u8tNwx9eaLceLI5Y28kHFtqLBjll3Jg4+xuOz
M4zg3dGvfanu9uZzHLAZQa5sXvF4iS902L9kFISG3cex8BaXUItvKR+TE3D7BaH8PAkTAT3kAxNr
EcvBEu07wrF32EHqYIM0VxbS5VsAvw7Y6V6EvZAoDR8w8NlMO6W+rjj3hCJEci1Ar8TFbT51PHx+
UqD4J/1Mdb7P8dHZiQTllkp9QKKCFUihe6YXch8FNdinCU5Eyb34wxMNUhK78AZOTAFqz7gtOoRL
U5JT5Pi8PtKiIGYvBhNV9kRnG6CYpQna68lyZDQYiu4H1wdMBOtjYh5JbTwXp4MNB5ma2kFRE5Qx
loIdEGgOL9HuQq8NrTn2bSWrBXPFP3vW/6m1cfJW53dQV0a4557MiHVyhBG0XW2BP1C5E//2WUas
D6fOjIqRVnU69kYw8Mw054LQnGG2Yb7gIMZ3PYmk/FI8ei/bJbSl1kvWvICF/OTCtI/Jl7G40ZnY
R78Nor36h+HBbOIA4biMywCDZSNAI54gPKtfSWcEPiJyTXqDsNnHfb+OWv+HJZ2tZxo5cJBF4pf7
WCzLDNyrJHGLJgOB9f0OdjCDn/cSmogYTlhGnK1abWaa3Twg3GKAXDZgUFz1SwxpoljC2UG++Zqp
d32XFsHguRP71leavpIlNfrisNMMZE2uQ6iekQBmDYoNq+cRhpxmPAKo09crf5vTOo2J4VoNJTUC
1xgYg/+XG/M/GsoaisSCzf29vER3Ui0IeuNIedD0Gcnof389RaMxjmDf1i8g2rOf7uTt0M9JO4sa
HTYOUXrPbG7ht/hkZIP571UJ1ehwtcG8klMgcIsujXKYma5EJi3aT9JtGjSC1tcUzupeAot3XCXQ
KfGfueYmEOGdiA1cp/tVdWlVyThKvTt0oZsvkyqs12XdUL+48w9OtkJ1iQi3wzAHVsvzQbhjRbbU
oh125pPf5sl0MFKV1pt8P02hrktWz760fkTGTeL3ZB+8jh+NnKkYuzbkBPj9ab7nXKIqik4WWrS6
NAfuBWSN3GAEghphpf5F9qOkKtnroGR4a/2HSt7Mb8aRTrO8PVUt28GdBCYquUFaHqFSCFGEO1NR
fJsdo5O5ocf/zf4Y5hK2nOh04+h9Giaoa/QmmeJVfuoLbPHQ4XO45LtRARl/sXfR8cAcGj/kjCCQ
45Ek3bqnNdLVp9IYEbtjDm65syGHvfbyhD171Xlj2k2nhgMhLwCvr+0G+oaJ8BkM6Plwohgryjrd
ju5IS4LEgX+NgRKJYvMkT2++ODn5sREWRO0jQV06TwYsi4XB7EL5593PZQUvwcI/IM7rTu3SdHmi
p/v8yiRWp9Ttsx4g6/jjcfIUUQWKzhH+RAGkFitpBjwoxwUDAFiI8h5FobJUUe5RDQUuR7K/8e48
Ng7WmfuvaAUJeK4Uhr8iGTJD00qQ4aHDyrNkrz4sjwYRmScUI8gTdr8ULdkJONa58HE8cnfHvPHB
BW/TmmuNy0NYAWkDvmI33vSGopYDW9PUq8f+mB2KSdKSpzGel+0PeVJhBKDdVjKom0JTBNOppBjb
C+QtEHNj6l/FVnSnOhjXgcfiyo0Gun1b5v/GO7uSo/bN/8BEuOxvgloNNLHtaTBwi6EoHOC3CB9Q
xjjZyLvsbt+etg1if7yVzsYCS/c7blb7S07B03HUE9xCxXNNjmLP2s74R+a9xEjjVHrEKZ5xMVEE
qzvPkthhOvoE6tDfxLu+ijHh3/abwSs/iME/dkaRHHOhdaOe42Yo/SBVFZvzFgF5qFDCJWiRy4Tq
vxZTNIGgMZcbZUeAjjOYcZ0zpXwnY8pagPHzOuka6NGrmW1wlFrO0AnaqeVBYikDQXrvKRw+qeEm
NO4EKv4iAf/JdUuf5760kTDeeffudnfxqrzlwj938F6lBH+DIQXD2nFOa/L6+ibO/X4mNNydt6tO
gYbgNh0kIWGqPzHiteZ/Da0Qp7AGsTL5SjqBzgki2V2fdIgp3cC53fNU9AUTtdlGmWKT875li4rq
MdvmXbvJMTsQjdu/ULHz0Ujd1AWv1PjzoQW/F9fX1uvBQiFdt84XYPj8Udby6JCc1FHRFT5Rx4t5
4va1Dqn7GITScyQtoT5KH+hgAmPShyDhndbHjjA9aLUkrcf560mgTehLb5vQPgi39T5J+E+Eouw9
TRK/5v546msbehcOebEev0+MuBGFra03iCtp+8+EALKno9gQ8FXwxq7fEmbVnZRqPLtNhvZnSCJB
dUwRlyAzOO4hbrFiiYvX3In80aX9PrtrG92bUPr/df2R5qBLxl5MgLmPJMG5iHUqR2uEdt2PWkFD
x6L+3hfEljFdN4EfLSikYw0ZDNdAFVkDE5muWQbT4ZpvA1LZOWRHiojc13Ct1Ao2BK0aZwkwy+r/
/z9c2Txu+raAS1PdJKdphMjRONlQ5gf9dLvLLTQxU+o18sOahj4xbM6vDsMRaNadSwSaiuClhfjg
v8KB6osbSSrzwrqiT21Y5sF2ZoNDB6dCORQQaU472gk4lNbRkngT6mdcNc4dVxAk8aaUCHZ0XzR1
cqp7sh+xbZLjU5t57H7pwIZ7vtlrVI9LGmR0T/CXM2x8tIZDiqAXFTdKvd17lkB91jgDRYVI7fZi
Z0gX9AtSY4rJPpukkJheTqCCwJaJeNdz1/pYfpmq06F7/Sx5uCdgruiYwqBowZUgKGNG0bYWPtq4
Ydrm00NkjBMOXYUr49OEs6RKkq6koRYkYB8qx3Et/9dsCc0SmpJ2ykotr1MHV7YNvrykeWUDoawS
QwJoyGhDViBGDGdyfPf7RrsB0V+CNFrPVxB5UZqkLKQwyY2iGsJ9x8Fubi/5xmMsg11sDZx5R08Y
fsda+RnpIxN/MKq776Q4qHc6Jq3ikAd4sA0es/nJX7bXlkuH4THwhL8QxImtFIKfcUqjmgyaEYRX
SVntbnS7CNUy4MFqo8W3q/U3H1wiVKmVUZGUEWb4Nq78J6jshoPA6Qz7g4ac/mTlamJcxvBaSXnG
l6FoFATPBdRxN8VlNkz2806KZ6ZUHowt9Czh//30sAo3WpHnFCuANOJhQfWIbTBN73NKJLS1VK0e
euhNPU9e2F16DIgrsmVd/GqFnw7i2dXPL9GKa214b79antO1uij2QQxll/cDdtJEC/lw2061o4Dj
sfIGXubA283FVjA68fy8VXarfJPld03TEpgkmIrbG1vB7qQfzXfyTajgO8PISVl7l78FeEUcRujq
/Ls+CmsEwFXBC68lvuwF7Z8jFD8dBtwh9wF1gLlkSviNkBSiR3+eGdEBcQZJ/LzHVcliAseezeNQ
JoO/zl7iFCCSaC/UqT8KPsQjrV6UY0/1F2vkBX0FX2+0psXSBHVsmmiGzqztNiYBqpmwU/pobEFh
9mxITIisOn5aTv3fFY6T4PqyjOzd+mpghxl/wnSZ7y4tZN2f95QlWUCDRuVb1/jB/MQGKBPaSBaC
qpE6EP5GXfYp0g7qJrmqgbwKIdXxoAbg3EPcemm4YU66je5Q5+Tjs/W8iMwdilai4Z9rmC7kveEl
O29ONbQ+8xHbfxQ+KN77Xs2ganBsNuOPS23rDBQ/WM+RWJdL/eQsC4gVsZ7piWizYIgNETQUegDH
SHlOCGBPxxyXnpjQSjgOFMcM9h1+ebMWDcvn4Dlz9HQUxSBYb4WrVKKLVADvc6DzQ5gNC088WXPO
kdAt6/75VKN/hy0nFtMhvWWKW7uJfG5kuCXIEhMQg0Frq3XdqJ+c1sX9roTNWkcp0XQwmzru/uZN
R0fLz/smoz9H0F5EI3L51JrBw/bLuT3XUnlcfaEWKri64Wg9vnaDdsOv0CHwOfqrtV7ZcxtVZrFF
MYyf0eRTGqFsvg/fCmKKdQziz1TPv6LwyGlBknfGXTE+7m+7GpjD6tXi1dme0ISbSJTsFNcyOElf
/KPq18f/da+XhkxMS31TMg8Kp8B9YZ/RS/jSf/IOI1tZGObzln+CwPC4N8h+QSBQLpAA2W92Hi2p
3ng0dvA4jMJtqHmpeKE5U82eMnG+HMLZQHOGGDHK3l0/+t2O2T0X+nKX2FL7jghrZvDgK0k2TgHd
t5hflM1ZrAKt66bvPDJXU6fAWVOaIdmvgEWBZMZhve2itBuqseW5wgfcOQxAd5o8DSy6J8vWXCEh
Pt2vRM+aH5JjbPy4d+BR6ccdRw0plVUwY8v2Qv4ZYE72EChDlGa0qurhwlWCE3K/f7MO6eY53Xe2
fk9FflvGOW1AtbFi37NyAVDf3zvNyQWrRkfGGkjBfOeuV8iIARThfDB+87aDb6o+VpiWi6Xx1wLP
IVQqVcFLsw5x4mNjECz0o1tCe+PPAnGsOBdYjS0hh8l9zSRYGa97OFodcfsFnwRrov5qhPv3Ug3u
oFzC1s0bRAn0nCA3/yKIStVIHvzAXdNecrnUGcLtfI5NIo1f88fjKk1qXoKMFSmS1ieDm6dDdq9Y
uQOTJl4qC6MXNQBq2Trvr3QAzak1dIZl2B9ZghkUWHrB91nR6PGEQoKrCp1GxS97BjFnTtPUCUkf
bCQysayiF3GO9BegVu8tQ5oknPgwP3/g2B+IeBN7ijQyZFDApSzz4oqJTjWGINstMCCrtBego74i
OS1nhRLDi0Gzlba3i/kH8nOB+5KWcikXE23ssLU5d52gooC1dXYB35+6vP3pR/tarlZx8D5F2vhz
ZOVus4lMuMRVSJnfFe79ooO8FfSynuQKxKeF7bqVHLqtIOcIos9Au/j1rA+hbOEIKN5oVPXKdRby
kQILXuiZn/sUtqiL4vl5XyGB4wlZ0gXAPiG8UTLUFj2kimsMO0gkiCVJAjZ85kesm3+hsjwJAAn9
hwHoCOC2avw+svFmn2Hu7ZPY8lhi64Wab1q78rfRG+28idKOr3YVo/Ji6vCkw2bcpVaR6GCE82Vz
klmDARdLXuj8vHIlojxh6vVpLnrHtVN5xdGFBB1ZoLogmmq1+mUEXohd6PpgpREyLRZSBqG4vR6P
ypXt5CqM9SQOSbI2B3SgTivUjaoPdsHEvfRxqZvw3LBiDhnJ+RmGwhfkws5fCdC+sXFlB+SvkkVy
uyhrL2ycxwg/ROY9jeku665hPwsUji7TvVv+z6MC0i8xZKWUDnWfK95yWdpZYMhAYi3vzDxuDK1G
Nm9pm8T78lP5y4ReyoYGamtR0YU6khavSF5TO5WfVunivmX4AUzqh2W0KaU1NophdFq+jJHUOKPR
4pI+1SDiBzwHWm0AbLtYUKvgYLAkzj789cmwtm4tP/ZdaBJMloTjwHW6l9SDgCzVTLPWbKCWLgvr
rsrfY9CuaGp8U6Zl58gGdVEJSoA+/XE28z0K2ctRKoMlRE+VqTeZuzW/beLxAm4xI3uZr2PIPcMa
N1R73J9AH0er3zpexrP1ZY1UXesqasn1fdXidoRQqtyFFG3UqnIOvNEAJmCF1vp9p2GvUFT9fNM2
UouZgkvNDzZmaqUQy7gAvtJTr7i5yMUw4DIEgxcnpJQqP3wzzyn57g348qZi97M2Xzg9fyyVuHml
Qe+NlKHuYssbEtukFUYgc/D3uWWlq2Z2NVgUr5/ZEOx1SmKs908um1+ufF0DS+WdbHVPc2vg09SS
VszoQHcAYLh14JY6rNITu9irATzsmQ/jiKeDN6rCkKENY7eDYG3+cvGUNlFbmlriayTqWtJURjhS
JAFCFKeIVEv8bH4qfB2sCUI7+ZJHrKNmSzEIPR50g2d/kTwYcrJZsU7A6L8KvzlyD5BdPXqyvl7+
WwYzX+Wn4ZxRCfR0NsshoF2WG1bBPsBMSrXrwwwEcXnHYvlUAVpIwXxCnqqqcpH75Ldxq13TFE7c
59sPckanQq55XV7NNar5e+fM2m8+/+mUFDk7Va2EYUhIoRJdeECJ9JsNi+BKiBTvQ2NmTfBqjmou
jqJpd20VqBnbu3kOXfNfPMSvX9k8ruyBp4ufsOrSQRP5VFHH7il+jMWrhwkgvmdUYtgdALapE5Ry
Q2MJ2UwyHr3NPWD/UFJH5hnAKJ3z9d7C6DTvy5I9YUiOO8wP3Q0zH/ZQZD9vK4yNu/XyhYY07Axy
NFuTBCYLoRN1Qhs/Ezk4+Ta7qyGYKKY/mK2sJ2YtUCbJ88+CNKpBIqYHI/OeRytpki44jRP860Cl
HzgqVy00FkcUvvUxHu1d3F6gFE0+lE0IPmYraqw84iq152E51e3vAx89FUV5sXXeeczkoAClhXmZ
pzOKlA651Weblipkx4uuE/4xM8plPlBW/Cfwa1tPTCXnNOldqv8hThdJUtcKbIaisVY6CgTK2nNF
dh+Bno2PYs9gnlDar38geR4fxM+M3ZaNDCbLzLLL0OwhSKXOzr0vbqByx3SHfWVCjmoaTOmBK6s1
6KxdffE8FOpDoOjKyXYimF6axpcECWweZcfxjOBFEPkpCwZrBDd1PMH6ZbsttLPAnrnEf5B4Nvba
BlluQ2YHdnAakaBw/NLfPSWhZ9DRuX9GyYVO5Cb1Y4mFMlp+AwEC0zXO4Tlu/p4PjEvlHiZPjze/
/Dsh3J4XZ6pC0r6R6iLM72l/S8Ao2dwir+U+6jriQnXoQJr1esAd7INeSDevJlfAtaWntPgyHeaD
VaEIUconPR5euSwb/YqAKQ7wmGksExGZDRqooDTGJQWD9o7i10NA4qEupRZ+RZq8A+dZu6kUBwKn
YyfjS9pGXKM67Ac7df7khI2NqirDTbbZGdlZflEgf89rAKUPc46Tcg53UW0bJiApe4zxPxOqPVYk
JllbbKLzsvNCoxnZ4GGzR1dvNhAaxuM7J7g0Kp0Vq/ml4c3Ad+uPzdMpIVGpMkxa2o3DQD+TAyBm
2szDGvfhOHPW9g1kN38RpeukHni0vYeIiZXkx4Ghf9x84fEbM76xNFTbq3x6THKVOgZLMwpW7ULF
tt25ID6W1VEsiJWSW5vthbj/Zvjjnfjki9pBACBhSoREu3JtTNmmTf+A25BXM3Ajz0dN7ebEv525
FI+n6sS3xf4CVH2ZwksUZIUWkxvmkJxcjICJhkOGk5lctzuzM7BhL3Xb4kZMSkx05PWKe94F8BOW
fc9BDUbU7+KTFgX5TOBDA6lb9J9yXQiBOwKXl9cqhOxoVIP5XOJPLKvLXv/GAUDda0U1ISLVpMin
zc8F3Zm+KDCnr5oG+aZFk8Lopcq4Osff9qnrMyf+eDjrzCvP6lMSErKGKzohPOHBXxvkcGsCz9fF
qC+kq6XZWAEoMwkTugTXWDvwSYruDv+GFThe1BWD/cvJ/1GqeDrAIh65ia6R5b9Q1ajmk8bcFbJ7
iiHtMy/K5rK3V45JQOpdlFDWt54LXyLbNkdK79S4m5KOmGFupm13x/mWV1d6FlhUpecQrJ/BL/Jw
iVG6hsaADs55U1j+HkqP0YDZ4y2AAa5mzGlPlsze67E+MDvyfT4UlcwN8uglBQOVscOzPiNt+Y/q
nybPzPN5FmcmmNdbi9UZASgC60eJXpv+qEJWCIv/aXkbq9xi1nAJUt451W83Gmpoky3b7bMNUNya
0u2dlHDPGi2ku48tQM+kSpzKWJmEtXTZ4waasOTsO689qbEBE6jvcnnSFwEkaUKZjQdncNESUkdl
rcQwAbR3kKlqRnaL4DyXrBUPm7BvpF4Ungj0ugBwNsGqOl7d1qPKFg3ndj8Zz/mi5gGwkGU+PmGM
wjbtJ8KzaRhbBSgfYEUQJGR4qlv1nRahou4L1N40zCDvZg3Kx137J98nJYsRLTF3uB5g68NwxPfB
ZUYLXtnEuRg1zlRc0STfzjgk+DLT2DLAiQ0DBGjqU8tGPLdkG5XcXuyw6DE/3RTAwtQdyv1P/KOg
BuR8CRrve3uJntycGje2lSg56qo/6EdGWup0ntMOuERe8rOYnx57tcogSLUBBFUdskId8d4Z/PIY
lCjKevZ3NepcpBRmndK9PatlsWFDDKYhjtrSDWvIURV7hfbMWTb7dhEqa0dWDYm1ELu9Hxx4L4/L
12bj5vFV2uqDETsPKKXEIeRYQv4DRvkuMjbQ0a8lPPLSMR2IYjpUou/sotES4JMlDUKyxPNP7N/8
tsfJhsSYiGHu0MBLWVQt06bZ0j4Ob6RoGTGogL8wdPUz8eilR935vXsW5VFwgwvK1hDr7qp0c0Z1
wT8DBj4Ovfse8j75inQHGlqIBDVop50gEDXH2FA5loyzaHXo5gtwKyXVmNo+NLgFElbmKUba9YgS
WkKQKYlfY6w0j3z8uAAf2XeoRLlZ4csZ7hvHH2KuP3LV+ZKrrac2U6RVkT2KxEGKgM2MydZgrLfh
gyvNFMmS0hAe8TsOJtbsdclUPaP7brNjuWl0cagWSD6f+/8Xi+2drL+OhIIU+d1GEQYgF2HLzkgT
TFFpiwpqUrhejVGtWl4ZjX7tR8j2lwzJsgTlBeSuiXQGEaFaQpvB9eIO0TQgnaSCgVyg6JDTIfPk
5nXyf4HyWh0ZGT6MzVavT6S1v3X88GQ9wt8QSaBOvsfkvulEDzwSEN8b4Dy+09UQLfRf5n8MD+SS
jE3hMKUzI2KlPi9rAptfy0pvl/JVNp0+KGHJtU4Sn48S/Lh0bCoUZiexKmoAHix4ijLEgpZOPXbO
1ZH9l6K2hz3HATtPZT+SnAhrZkcJ8ehulBIS6ALjZpMYRrnn1SqV2kpZeEAgOGSS2fMjMOdiAdcx
b7H6xCfYU6A8RRDN1i8hDDc2zLeIvYYA6cUeMn3EdRUxRRFOQkbn47QFLb8NwzSeSBvRfcE5kab2
ceS7vWmgmQRrmHrB4mfOemqXRQD+wQ3wM9C8Z6a88u/2hwHPPf+K0lUoUHBO9BhheOyaIvXj4zJj
YrFnp4MhN+irxdeeeTNjVxF9ur6C4lbs2I5ERsTJOYFtP3ypFrBrgJPoTpYjIjcLtc9vz/BInbOc
mGxzHjXdtP+qXh8H9PvOGRj3/rHNDCTtVIjmLhnMIgWrzE3awjPpMDdvQMb80gOG3JIJU1fiTfRA
LTeEeZBfUOYykYddz1eU2F7bLrg+UK4NpAHEe9s61G0YVoG0KLi5P+8Lts0nD1uzpcFxPtUx5L3t
YL4gFnFB9nNQwQ112lbwZ1qTjIMNTOasSdC2pVfc5/pbOG4YgVbtSc5sO80hP4hQ1xCpqZqZMzzK
XhYP4ukHq2ruK8I+zLlq74VP9wjamzmci4vqN9SOd7lIwK2qOlwE4O21cFLPVoQn4hMBge5ro0AL
Dtdep6B6LR4r5Iqk9kaJifQ3lK7T8hbhjgcGgYVmOVdosDqgo9U1kNfzP9IOu+fHcimf1XmItSAs
jemlq0s8+p6Fom9idoB3X80W4wRaxlLWCvAhQa4u9anLhQvupo4UUvqJWV+LIXFMZCoIwR/gnBIt
lOQNhELHWosvtNKFxDyaPf/VD9aGOb04THpxSYQohx7UBsSDxo77WVa3l3T0WLIWbCw+FLhMz2E1
6PFKI+mNiP0v9OXC3dI2J3QMpTShD8ESWq92yUay+z4fhSEHEe7VLTXEX++CxqfLMCLmPHAiUZOC
Pjp9XTqAvVPxUsUU2Mbstk1GTans+0pfgXhOnV0xzvbbGPyo2ldAoA1JuBOHKJREnUQu2CPJcVcQ
lOCKuPVShV8H0ny0/5N1aTt7R9Hvhi8PVbErKMgTtOcIIW/IiWgZeeWT2BU8F9CGP5porktlG3xE
2CSRn9z08jukCKZbd0ggGnkGwecelOaYnPPBNmUwulkIxN2wmaPTPCbkVbkB9YD3rIGUdQnCi3SC
7Ls7AG1HAP/Fgl3yqUN+6EJ+DKDrLpii1hOfRf5fGYVrHGKYHuJE6yHFFNxFSwFKLIYrjV8D/63B
KgsmEYCQCbu8qTC2P32+7gwGulcWZ9BNs/YaKRXRtxq0bFGeG/ySJ69O8eRzDT1rGzA5rYhHJ4LO
G8Zva8gKaAHsluWdt4aYpB0nArnoYPJ81VzvvSl1ouDUvjDoJJVEs4J8SmoNBxFyA1f1SH4blfAi
RltZNNYC3VSDHNBU1XJHcmiv8hQXzFK+mwGV8Y0R413pab9FdPPjff5gR9dKmGd1Noz9Iceu20Uc
PUn80Wbq6fj4CDRJpO4QbRa7Hp7VZZ8zHaBCP6jpqsFoqYO1j7IeUlHpYxJbuhm9qtJf5JsanHkP
N3i/uiWOmGsfVxIzkUAZNcX8iCU3quCe0do9g8vk1IpM5sLCxa9P7/CUNrZ6o6cm53Owp4R0fNhB
/Pz2uKqM4N9aLnYu0f47DBBs9EtqoYCpxir77CfYWyyn+Yb/pqJYReEuzs6BhfA+CubjsPuAl6Cz
/gwRLCCtAHLdVwWzqWd2L/A1qfwoIjX4aUX2QrS9+acBYAV8h7kxSYwSi8EPaI4yAHq8ERINZL1V
lOXBUGSW2r3+gk6Y6bT++ZQ3v7KdXE8Ad6T7CLDP8XNR0pneyoRN8j3U68GUE2YdpeBpm03Km15S
EgClwTzUne6a78FXj3JaM7TiZyNuP7orsmQBHrWqDaavpz2NxqpkZ4syww/7mViSvKoIObdXJMwN
kdZ2vy1N/zN/jjMlRXAC2LJ8wR1EpsiryQKg4ZO22EXsqQ8PT30Or6cPjNQidq3hHBZbOB+tDlxR
GTN5ogldAwIgac2zIwFcjmM0an7OD6TOAeyPy2osBnxFNw9Ft3ZoiBMtBV75iBFfMOLWX0Dj3EZK
e79SEFzl2vS1Al6z/Z1yJWj46F1pV8NdF3jOk52twQtK5kDqfRFne6tfrqZTxWHrxfc5HXEvi9aU
shHyg4y+9n6yLx1ndi95FvF+nb4qkUXQ8EOhatqGZFnq+FLUthGFuIMASfToXNu+8qRncaZxmgyd
WePfvWBvmvwksAx8DQQ7Xl5TbegbSwRNI4CiKZYGQ/Gs7/TduvBbWr33hDHYe4SzSzfrr7UOnhYT
Bl7gArUreDIn4EmSL627Wu0Rqn8AoIGDVKqi+va2Rbi1zfXpiBuJ5MfhacE0DJdSpaOqVV2TwBKb
3VTFlqmWF6AOvwnCUmrf2D9XorXIADSYFIYz6Rfcht7X6I9mvidixh887OqHKlE/KudWhERe2vOf
iUb6Gu8+Lbxz5z8JGhcs4xkXx1+EYUKr962Z3CGTeHdv8LsTL0wHt8wRr3e6/yqcc/HRWhPRQF4O
hPeWif721ao30XE5IOM6Kj3W+Wj58JtJk4PD2UBaoXaP3IWjwr27A1AsqbISCEfQbZqFHBp2fNrA
XDt9/uYqIcRN5L3N7dk9rdUsQFr5rdQFcaO2zqCQtVQZf22TRNJaCk6T70Gxdo+sy1bUa+7NG5DD
7oTuVsXUJwfxLDkrW5OiIm/lyNBzggPdlrJtbllYvacA3oOXstcCZdiXAqgv1h13euJTD4vGge0w
hO5I9RN1gVPeY1we54Q7IkTPMws2HkwYrybaFgg60XPm2Et+gnSgpLzreP4C/I/asxI9fu41N0ui
Vwbb0MJ75NT4dYaL2FAmLchTeAU/vp3RVS9sA1aQdTuHlDeUN3NatJC08lPFRmk99Do4MYdIroWm
1eAhutOWLVJz7IQnrIMnqOr86JpB96tkKUXMpk7wp9QwvNLq3laVsHsJQoSgJoiVBzQ+nQotFA1h
59QUbnoVTWk++49/9oWVb+V5zEx0r2zwhXGceEDUoCDibTonQbWHXgADKtGMT/UZbNxyNwcJ8p3M
+MfJ1OgHzWX/mEefHpnElMNtNAPzd7fVXSjhoM/sHe3M47os74R7vy8plS4kKc44KNW8+CNl9VZs
FkMVLwkmmYVdhHWS6iS/5zygzVXQoADQWpiM3qB5aJDmwRTmPZv9H+3XI/sfpQPW4tTsjWL2f6ek
ChBPXmpKmyXleo3ZwgzPMkSTlzhAnjqc9MdwQUWjyFaOC1S2f9oT7wF17CZm5UhH0xGpe9MnIC4d
ioHaRCGsY2KZSfIgcnRbpEw+06vZIHfTXCfYF9DN2Fm7AX+3mocjQtZ0Z3uPcWoG9hPbqZpM+/Sj
06+dfmK+0aX46QZcbSCYmOfE8SfacuIYTW0BH168r0SlCLyOnoEdBlThv0lYNzOS+NsEKHdJPdfb
T7Vpr/PfXfbWjFM7sf6Gk2XdboX1V4EDVckvVqM5dZKASo96VrffH/yWOGv+kzkJR3RZvUmnlDIa
I20rF1byIDiXi2XJpWQqoYzzExU6B/nI6mGi/bRyUWmb8NvS0BEhIk9xAf9bRyD2DqSvkB+CzLbt
LcSdho6Z/yOPKZpvmJ9Aw0c3i0m1nzH5FtKRYww7BBbOCC3cgvQh1aO2/GIsq/LjYpsXXl1QSz4L
Kh41cNkNVkfkNHEzDDW1lcyOv6+veqSvrb+/WY/yF1/aNVLu4h95juFHT5KTK0moB9OBJBxuvpvB
XO9dvAdhUUfudNqSWtFPX+P/s6Ye3Mj7rmvRt6J8Uo5v3e5cSV0SM9krm8KJ8leglQsUg9MbkSWu
Q4Zk9LobLpVzUdUJa6s2m5xJTcwb4R+49BtQpjN6UHQxyEcAfyeLPNx6ZPtUM1IKEsP9TLifadh9
qJGGCEmJgNSQqljcVuWblCVDVaUzURHKlYZxuRVIzRlXiRjghDoQ7vXm3WtR3b1r86+wx1KaRgGK
+sRn9prdKsHPelJKoJiUakY2STmuAj+OqNKEJIQQrfDZhQnck8VfBWFHpd/XkgyQDG7AxwrEi+a+
K5NjEaYiydt3N+mEKsUVT9/1S49womV3Kwg88Vo/22EbKBTMZKEquIqdI3jxamQZ69gdMfeszSps
rZVek1KT5fUigDhDBH8D0JNIv4EObTr7uqV4vV9EPSz3rVPyxJkP3yBRvLAyUe8x5QrOJZNqcwjN
o7gdoMvU62W0DHsohcpAwFcXRCVFFHo77BaFoMrZ3UnOFKWw6hDPFJwDlUaFlUEDR3SUh9VUsAmR
k5SF64I3BYOagK1cE8FomyWfQW1/bL7oSxBtz1kuNZgDtPjquA0ik7A1VanNQM6ktirVmoubkZuh
wDeFqGaJ8rB+3Va+bgLjN5SOaF20TPWG2ESvs7RDrsMOO5f3EBu7tmWD28W/LGEzBK6HawCCZ4dr
jxN1Gibk8rFxYlfQvgNFZ7NPc/MX68eTu/TZ6TemtYhNSGAQV5cZt/hby14nOkkuXYasLRFq4IaF
zu3IMf/LHXQa4VgG37935j8wOhS00i1RlDwjj105qaSvNuNNtUY89D8ZmiLofYvf5DLz3YZcitHV
+2xEepAuxbJk7CVqHcskl50TWcfv93sbYnvGDI1JU8oZlG5Za7YlRxURhxhvlff2JF/0GNB7JHNw
HBWsocqGsMAbXQBTmX1DemNcdYYxJArMUaPxUdqq/+VmViasEUofTKzOgpn1KldFXowUEC2t/g3I
TJtr6WCKEwdjn6mmAOBHa3jlc8OY76rLEcB6zMdYOzJxHr0GZ6m3nYuNeSxNvaXPEmLoF5j50HHt
GRfumsxjEKq4yaJu58+rkLmG32r1lDGyMukuDBBAzfHMypAGZn3x39R4TOOBf0bFb6NXAZgcdWm9
I6Prg8cVHmNcsnT/WrX/qdy07dHfRzLvaa6rJP/I6ygxSdxW3gleyndvj+VOnXZWpTBFgeC3hVpt
CCUFUAh565FQJevagUAYPpnrD/8SEYdp03EPqexEbRx0e/a6K60lek0Zk6KQj4hyrC+BBKmb4mOe
ISZwtcvP5DEkR67mie0phDbWC7pvxMoc24YQvxBcZAiyWxSF7AfilNAH1Q/7sNbi0WcRwVT5kHA3
n+qOv9/ACT2xj0lbmutclJcuwpuqsXWPZrnipFIvTps4IuTwfmSp4stcuTKSOn+cT6zWluF52L6V
f0ublxti7lpxPO9RMlhIL9Ym72VeT1qDSJmWQdyTZM+oiViHE3UiSEslmvtZweg47I7RePqIs5rd
mkoszDPufsSxjkW9P/fjr/9lLrFalVnfmAs5VqtHU5VvnegvdrHdhyHOSXtVRxwLWwZ0zQm6gZQG
OLHWwHL8Edvl3wRf2rrUiRgQ3DCtwhDDq4tylghCq8YEwLTUCgNC6VF4l4g5kzU5wbvj4fRkfbgs
v9BaPtn+ylnevwFKOHAJXNmvsa5s7eaZw6GkercYpsSYqWJGoAg7eYoITCkgFjhfQv1aeUsQDW6u
exa8irDn6XK9V/hShBpIDfWf/9psmngdOkeY5OaU3zLi4NYu2VIA+zzyZ5XZFv6fcEQlh+4azcty
ciVCGtC4AyZKPN3m+2E9lLbdHyXwiGrfLj2EDQc5Tnj9dECrouyZcYO5dEu9YqjqCVM57f294cCi
LTUVwOl84ex4bj5A9pUmHyWfJbE5kSZeOppXatEYjx0VOBdFzfF2XgJzgYGZis61U/zkPpLXQML7
PxsrQeLRIzsco+Q9BunOcmIjrrR9W5btLNXBF0iW6RF4xinWbAdcHgidsTUsBQ1v8hoNBtMYH9fG
Z28kStS3DGpULOYhdwxQU+hsFOm8Y5g4QOrssJWNf9DPWrSjZg6PJ1YQL2Y1Vvw+jNeBltSauofx
loC320q6VeaYuamzTv9Zfl/7TqxAgsoHv3b4HgYsLbqGuk4n+Yb/EiRNYXpHky/j+DT4iA5r47g9
aliZItzWSsOETJXZyA81z4lShjvB9nCqpiBzXdwfTo5SAxdBs84KsVAFVEONwtble4Z5uC7RQpuT
MEy0abN8uZzArON+D+Mx71G8MPDLvaqeNg4dUuYjpoRocJhb2WgOkT6LrYh710a9VmSq9fpWFDQ3
hleoiVnKinctZbo0MoYyqZuBf0iCiOJfwoVkOa/jHmmRWawUXL8ILLu8b3Mnlk6VSaggnuOCttKB
p3I9Ta28G1CK7UQdqqcF6nn2t7BU0az9Uw8f4pFNnKy1AnYKn/uBcgTTSRF+ddnAyGC6cVDB9SfY
CHCbNMyRSBt/XxpQbBanZKnLkifvuLwgAO7i0juqKNNaGLIzHj/GWYhHrDvRsAxK6nNwvc+qtiB7
bQ+jPP0l6IAdf7YUoYFUVLfyXQgNJVKUc1alA7Wa+AhOYXdJVkVl5Eo8BiQA+e5ZCiGE+kRADL7+
xV6esBAfhEzNQGSwltBrxCVIu8CRTA2ZpH3QoZm3c99YWc45ImTvl0PEmaurCKEmsJ5mAZfgEeiO
KyXxtpmkuDMl5ZJRN2WlbYpYLcFFkvH2vpivLxOvSQAZvBTjYHmU3oERiS3G/URutu/LjIel5As1
y8+kIByyXSszv+5iGTlDXFzzsYUTk/4vnkg2CDDeQtCR2/vABvLXPiy5tEHJk0IN2ELqz/iX51gE
LBBP/wiGS3AUViNjUGKvX7Lg1RRn6si0TNuAIEwUcjXVKgcQDjMwHp/lZs+LCo8y1a0XE17MdeLT
SNWRnByY7JlCQMaU7TLOyFGKfji/sYE/YQG04UMvbgJ6AFw3pTlmTzVvqapknd6V38seLVVQpdYG
ANiRMN8Jzq6gxMm5eByqOZpkCM0Wc0MRh4ceK3EUBHPFgNCXWuyZEcELYVuU4NjFQpIKha8u/2NT
koOtCdCApR2T2Gfl5TYT4o1aUvIbL2woLxxWLM62Yt8lJZkd2tjxrKdq2s4P7OolcFPa/gsDcAUk
HPWvB02ibsomZRf2FzJ6p+nFlKT9Vv6/N2yPGgQNBoRtOc3e8JG+m4EEEyz9uxQh/5YJjEiHSta0
r4QbYPqXLzOtH6dtdTmvBZfnrYnJOj37hDEOBtRWHOZ2/u6aMtSkpxqnhF0UN1mwPVIzwc9bUINa
tJVHnaFD+MbtakvCu3CZfluB4lq6KRGF04ow42C6I/otEfTm6Zv1eRNeqgUWZtwC7pTqSpGLSCtW
F6YgCwlphNIH43o4c63XGC+dlYXQBmcP1b76ptoWsIkgz3peZa9SerWccr3BLLrkFFd+nZkCgnEy
ihsljbPAKNgIZRMm+m74+IOh3IiPfyRCXrl6FlAMO6jQDKNnwyg3ESaKV0V3U1budw3Q1946TpmC
ep40ihQrL47PXUKKgeunZU+6CAYeQITUTeT9hHeKfn9RiDntZ0sBa/Jne1AhPV96juyam6CySA0q
FiFqsnMDDGQ3sgf53Bv+6Xy5mqJP+GltL+aSW+VN/tnhqsIh0MG6SaxmzFPOYk1Np6nJBeAzDa+y
W3UUwVTAW+cQzgtqVhd5Nq5sCmWjdo3E7nfbSAVdd3sBOG0Au+pWHyDZh4ZfxBV2JINnGcoCqGRT
i6+7lNFV8UAk98j31KF+j6Jruj2W6TvCZGTLTLptyV+H7AdvGyIKdO/UzIco551tRxXohFn+0aQz
fOIjBb87kE/cdKkd6T9fJ82AZb2LJGGqCaDikdSaxd/u4WOQVNhmbR61w415wdR80nH7Dd3Dqde0
alpStr74p/DxlnDdXo/cMic29v+xunnplhy3AaVCvjEPanJDk6/LesaJZreBFoqksVKjZ2neyypX
E/2a9egoUTJqVL/IWAcGRi/kjn3BuQT70XBERBlU0FwH5vSQRwlOWQCu2wpBJ3iwFbaa6eingP4t
yTe0xFpjOW3ac+f1cswo/SulVigpveAkwGXLZspbuYanagUbobqMauxgBTucT/JOcqRXqjh1cDYu
cyBCJIAejDYokZbB0uilo7noc5hk4eMvLiSz2Mb/900Ozali8AbbD4OXL7u5WcCYRSgXcAId/vZO
z3StnJkD/71LfAQinNci1gJ0wgdv6jS1difptpdna/OAaEQFdPHXDE4WDW2hpNGv7gy7MsG2XF14
3WbZOQh1g6+mS2cbCF8lkcfeRjtncD+oq1wyXqw0uMu4r36gfByHm9GvCBQ5FLfCfa3c1eZBZM/1
CemMEvlxSaA4mPMyJ2LobRY7KAfU6+0jzspK1dnHA5qJRMdMDd2aOeO+AcVKmorwprsHlzLbM+lR
85qY1C2iCZaOB6mHtY1w1jj8pxrM7FTJiu04jYDkyHdKHEdNtyMCUYYL6kA2hQfs/T22nM5r7tYu
16t7JotbbDrr5Hkg88Q+1DGMbsogkJO3NdY4gXUfa8nJILeCGQYD1OfFOZhwm64alA2T5P2ZD9P6
iC6Mlws8C9CwdSb7d1mVZ6qAgygrAd7AXyJYGRXNyMU1WiWyEfOq20dF0quFMFxQZ8JsEbJIWY6u
tPERULTKoy5eDsSdjF5XDFIkCbbHlEUjJPp9Wenn2PvwlJJNv7Jv5oFRWCS5XDc0OnpB2eeAhqCz
LBWd/XNWvUCfKNfhQhcqAX3m9WrKMRpmveKt4eAC9ZHk3mVwTHZdQofbXIgR0axfFw1F2Hv/m05C
5pKleWPeNRwfvqFIwEhBQY57wbWxK2znuIvIQ1utmCtS8BMr4neoazDUxIUsC9ohy48MsDvoR3rl
xwnF6+g20NSAy7MZnTM5rpqe1EXuITDaJMbpq8vIG+1xfeH1wUWCID1aOVtsDoRqEtOvxd96yJKA
0MZPEczXlP+wahzcNG+XvvjbKqNghpBlFiMlherTCLdHDqjMglaay2VYoFa0wNqzTt1bJFwFxUHB
hB61rT9ze74pz9nE8m2n3CSJ8iWMk0ydDgsoSlsCGFMrkhFblHTM4wkDE23mO0z+kUf+Tn6XtO+S
O3NYjpSQqUG2IgKipV4bVkUkPjc0BI49VP9O1OVfOAJ5jAqNVP5F/6V01QI7HzxsVZjYtfJESLad
FKkj1zLuq3CKAOIa/6+UbkKiDUEd9vYp6EWbGk0JckLhjXJ+AJPBECSWGN88LbveMRuDf1g44Rvw
jMZJKCjmIVZqh/yTpJOlVIe81wdMM3MnZLHcPNCgZE/9EzBzsGuqbHvybM3aRb0CpZQbLYjoivvI
xpL9osYY4OrFHaPybbFdcbCNUa9yVRmBiLx+BFGxK4kOvxWbjD5nYD51UXUQThafWAqQyrHWn8ri
n/KAxUtAJPaRACaXb8v6yQF/Zk51xJlVki2F/x7tclsIeJuPSqShL6830lBsDBWwfg6iHG1YMG6D
g+t+EC/BQdHXeFZ/142xzAszgC3amN/s9z3Z7S6VTVYrTzrE1fh/eMlk2Wl1QMldXDlg1erXVVGu
4vqL46YP0KY3vO/3fkO7n45LdIkgVhhIjCg9tDTDtSmEdfpx6IqLVVvrZe8IbzMHEA0F+nF625yM
A0mXgC5vugDcc+JtK2YCGE+ffZ7SvUqAG+W8lcYTPpoIF5DauOG8IpFR0FP3U1NB++UC2COQTHq7
19CNpQDzKXng3wllLaILT7wVf/ZVsm9mAj9BiaapFMAIMnrkhGbS4IvwmESO/x/4E2e5pNeq+ClY
t/5hdMWnBbXGdJ6egp93ud3PKYBJjfK6XyZiWDyjG7bv/Vp1sxxWE4ArfoL9QyCGExz9Z0sSAlvU
W9ZU6eFRMTHYS0FKcA6+hHdr+FsbQRQvq7mJDYOQDY+IDWYnE26LvH1ADnSAmrgISVorzUtpSZPZ
sGeP4VvWmIa/Fzdi59txRFgg3rKMSvsQqc/y3DyTe7QjTDINGBGWqaD0lcLyhpgXGqaa/XjjdsjB
LxW2Ngi8ffw7oezTo2M2Y1oyQPo0r0pPQWeGkh2bZbq4A35KpELLGnnrDr/hTkkmbg/DrK8jz3Hj
Ol8Re34fbQNuIXJ113JWZyQ0S9ooL29OjHOnrBvpcSxP2axU5NLiYqPnpOcM1eTnq2DvxEWAt4VH
UniJnNdsHDU8djv7lHGhfH7a/yaK30dMtbDA9+0f+FMYmcwAwNlGfhZMPhIpomzrZ/AGxMxvMa/w
wQjG7kG8XhDFckied0vvevNoAOMIwask9gVwJkaRwMjTWJ8c+8ImJ+PPn0njF0AWGAY2ehCusrx9
dRWRlOvMk2j6V7fDiBdE/NsLzP2HT8Fes7dtWpp5kkVZiMuziuC8t42xtiSOfX9MKGjodbH8HVby
lUu+/WnZBZrvL6r7IvM0jZQ1nMDdEJ3YOZCXWu+JiljjO22XqG6e6H1hp5WFqXStJ0p1DClOIKyH
EbaQ9uO+e5Vp6Uw3/A8RD4tGqKxh84xiM6dELELHO8MioTW+hO65GABU3vAYV9OAfhhCzXUq+XrU
rGIovVddmfFgi2aPM7w2XDatL/RPCoirZRBZ7cbNo+1I/wHfDraYK+h6C575Q5fyo27I3aiMlnWi
RNUo8l1vvxJtSQfO42hR/8A/fd0QauLJ2IpPd6WV722R8fHTR3iVlyFNUtaDDv11XQb2W7tSfPJk
SlhAhkPZTpHJwh3X29eApkdKpGaUEbf1A4v7TJuxf6EASH9sAq779YXoa6pMiZ34+A33Wtl9S6hF
iviyMin/vA9YcYzYK8M3mYG1q/oUSlgAK4xhAjrz17dY4SjdrUpeFrJAmrw7mhsXtRKilqj+C1ZD
2z5P5yY64fAwuvv3W2e5l8HxZ8b2Qpd1rYY+2zbT1IiACfpOeNAUTGKviFZip/fc43RWIIvGIg05
6T6QCSvTstRXPWPncRtuPZ6JDpZbaIShVhJF+6qe9Ej47Z95eS7rBPJQD3IxVzgGetsgv2PDc4Df
mibECMhH87hRY9LI536p/VBnETCkWt6EXW/9M1iyZ0O0rDKsVloXqmjIvsDRjtQ1Esi1oDusC1AV
rbmvw5MzRg4/24UYdlSMMJBypK1hn8W8mr3Qs+2C6Vkry0iWHbSt00z5mcat2jnr3MC6dDBmPtvg
1b+oo/bNrsupLGo+Nfs+YZ+C4qmfpZlBaEewH5Cvm0MiPSoygTmrUplIUwCeRk2oF2VkRdLjVxDq
aW3TxnJpRQlrcBlIrtMpa/ZCeAp+7IUWtfca5VeMH0HWV2sMPiHpIIgh7in20TSv9PvxqJgSJR7D
cX6ct0Zt/Aprk6Xav7WSA5A/y0CiafGm62tfSZcZWwnSCcjTBT5MZQIpr7vzAhsjq+f5bKkbCCWO
VdSRlaukn7VwmPvl8H1Y+9ZoWh6XMhSJ4CZLEVnzFrWggXJiBXJUe5EdvQ4Gqo8aNsVC4SWyRfXO
2sCBILIOQ5woCa/18f80813blbgtkONK6r971E7GoAnO6/nd8mvpsSGCsdhn6EAFebAr4nmZk6FH
0SBa2al7lC+woLzUX2R7cENMUrkW+CUOygtaBKDbYPTIrRmDhtremOywDXY3xexr/8wEduxlHMgh
ZINR/1Rswuz3GXqEpjcpyPvQix9rrL2qE30q/OLZ/KKoRmAjtoVeqDk82CmoDhpexnr+FZ85BMFl
YY1m6tFzS5rGb/wDZUGygjfdSE1tz95OiF+GVvjaTrrKbTtMBKp9wefflKf6+jVUEvAH/ZEff9iC
Z4KUDTG7G3OdzEmvhwSs0DXJLWwxcO6E3IYJNhykNujRKYkhNY7JNVdv01anoRECU9RGEUW3g4u7
FKnmgUM8s5B1yO8yDV/EeqTOPPDPuneQOYmmk4kI9pTXDGjlyvuM8gZ5ZIhxiv9oN0jGJeBgRSe+
wNUFZ9jwfaxhtSDTB7tbyX2RQFG+oWsx34xOM1g0aDYQ1fYTT49jeqomheoh6xMAuv1QA6mocT/h
oxumdw/VojOiQllhMj/X/HIvXe4XufxD07k3mJ4tmYtdxAcgcaw/r2+UawtFeNJVW4qhow0O4IsD
aQB+xS3hTofmu0tjQq3PwTcoQx3G4OcqHhmoje5dZ1Jn1ZaQnIPe0D8WwYW67XsVVjUMhkR6HbIz
H2hfckaS8er3XqdUqCrtQU5QSZmpb/jbNaffcm8DOnq+9HRdz1U3/Qt3gEE9OrWpz81Dclehhi4X
RT9D1U59lFQ+wxU1eiBB09rkvydZuUViTw3z9/Q5qo8nuuMa/ubIWvpsTIlH+AQ8WDC8F3VBeL5Y
IRJsIphr7/VlAyBeAghr9vJvNhhuxXI528FJc4v/yV6x5z12nJe8N1YL25OLDJnX11aFxrjjZF91
kpJF8t0P4O9R+8eHX8o36FG2waYHK8MLBnKyJgaA2sqoHVBYiRW2aKcQdLvQWcwDLsb3vIB5/m8F
X8AYQEHmQ56rfsR0uX29gUpRtqcfo2moPEo6ck4QkMlxjiNL9GnlGwg4Wh/Vffz/Q0f+9Sovuk32
5Q80VJ5/kaw/bsDdcdMdg5QNYfhBLdk/wcd/EGvCfk2AAZI9mKOmt2+owIn7rwx55/diOxyqrkbf
th/Peh87Gd+eBTzwZklohZ+nF06pKJh7yHEiQ3zen9vKAkNZuZFsr55D5O6yQOscBRfOThjWLBq+
1YBzxO7yljV8Q+NwzwESpwwHZkqs5sfh10PFKgM6K7nE2AO/e6RKujCcE4w+CT5XxChKNC81ORow
1m4QaPK3lN0yD0gt7ReoCqL3VcJgphhQ4IdrUIQC+72T6UaxAa0D+cN00DxfoNWdEei7ty3j4CpU
D5Xqk6ex7xlgn9xUu36rLYdpUJhZLYep2vmnsdsLR+lWC/aviv1nsty4pikqG74p3/mJfiDMfoDr
l32B7S7OhYVcE80o1ASY2CF1fsQftJbgvwl0/KKrP7DS+/LR2P87mb1UOZVFBLigw8l4BAIwOJna
lGbea6poT5kksj7nFyzhxSpw75DChrbJy0pgsHWySCd/HyJvihJc2tzMA5DQmQUX0kLbrsvwXCNw
NlUiAPO18UYQmZPWIYMjZAdnT5RDQumaONTsZ+twBY4YRKdGXfGupEfpSOnjcnc0AQ+3IIBh5hbf
ZTE/Ye7Isaxi55QDqry9GfFoPUxJEzaKD8lmP4T1YiMicVQQ/AFv5YDyJvKiO+UkDevcl46Naz0c
L0MtupgcZn5ABikvzaRvka89QRYPiI7AgmBpsVrgckJY5b5/YmcY+w9OxHqJZsvVetyL7E7sQVpz
uMQk9wtupKeRjzhXTZ3G+o04iJhtC8vN+KK+YiCDabOxv/YpAiQPLZd+19k2OP7ql6zgPAXCATCM
cHzqt1DaCOgBmYO2koXbKf15zbcljTzzZHQ2RzskCB/ecpj3Qdz4geGxJiKQ6iGFnjlmxKzz6kmu
NBFkGeCmCcLzJNmFBIVhd4X1cH9F6vmnJDJ+jsj3/GJtP1x/gGtxChP8MrBMb1NKg9drQHC7vgs5
iQg+UnjWlx2q7mp1teT6U75DXkvwgspvXtySkAC2X9iC0VfM38iLLS7QUWspSYk76X2sMTohpikz
bGexzY24BT5bFJssvlp3PbkcIYpKQ3r7nn+6b2CjxwZOsgzyO1eVudmOV8kvnzQeYKaNXTKzcGg3
9cmG9uvtjMRCKFEgDldoRaagAE8gSCztHQNLbmcWnnDKkszF/qMfp8RzcuHOPNQH2nMJbfxoj+Ez
17h8sPRc1JOEmStdMHECPbfVZbmnZ9nnpdbI2Y59GnswK3hJrXmYLxKzWn9PptA/rvmQnxtrvw+Q
A/plYfts5BSOQzs8pS/1g8cJvzPG4umQ/NqR3j+s39jK/53ijoEtj4s/TZqlt6JNkXURDk5ZDT3e
0SUk5wQ3MWttjH9CJhIgXD95L1FVDImxi57eYspuBkuOTCQvllBX64qle/hf55hAArDwxTaUAlcP
n6GJObL4jbt1wB2J+xuvdEXgnZvGsy+XTyEOkOqjFBF7h7DaobUUcQ/KzHsSJUSjSLY687ZyUhIq
W2b8WgIJEuRqs9f621Elw2H9QfRqV1cdymJkZvop7XxhxW/lyvQG9m62gHZCp1hudrdBQKGEltva
wDyD5PUJXI4mzeKEnbuKHYZFgugSaZSW191aD8+U/GosQiP2Q0U2NwvYI9KDm+V537cby+FarODX
PSGd6ngU9PLxyDhSY7hegsX+/yBHPPz2uCmg8xikOAWk7YdSRme4/BXNjvIY/j662sEcfHN1+h4t
7mNl3TDuqS+jd1fSv4jNyKcvypv17/IlaWIK8Jv/2mvs+vlJREqojATN23rk0Cho+7N0FtW7GazO
P2fMVbANEWwxE/2FWZS6Z3B2p13J1g43xAIBNSHdmNAMhmpCoLdB6kD31yz6OhpsEnC094G/QAQz
YaoJRyzfnb3pas7EiVn6Ea7OAu4+xDb/GV5JVO0ReOtVOCRN51o2kDFX24KkNzZJoTPZG71JeFSf
2Ixce5XNhp6UpSgKEBWXv7VKGB2LtquNGVyY7qh/OPNQfEqi8c4sAScilRBJ39PQLfbFIAMRVyV0
SI/pcaEN2+3QfjTdzd68LdaCOtSgNWdC63Qp8jFL8eqstwvNN99Xu2LgZJGZPe51DjbHWyFjdxHJ
T2OgXasdaa5Hxqfc9HjjNTw2VoCRlntLD9OLXaYZjnGu2kShKRn1XlqpM4eQueM3mFi6kr6ZNebz
RFMPYg1a+a+1NhYgI0TwqNHU/vWKLhdZfo1KUIvfXW4u7eHMXRvqihEE9t6ljPtVJAwV2BulMg3Z
9MEHYOx/vXJI8NCmWzzQOp8sKclkkwaEzbVfSBrIJONO3HKe8W8v/XlaLZnkx4Txb3UePxwytzlV
VpuRR9lf6HAAtHy2rrcqj8V0FbHr4vqji7OHH/w8brrsekhrargsZttSMtjd7pcXMroKDeFaBaS6
j4xYHBPdgOmGuiYaEGaAv7rYfWZ5NxV4qniDRjyIaxScmTdTV+4RTPu57g3r5kWMvlh5nBQ+NIL+
QaHojkkSn+WohwpZ6tMT6CyDGS7jHWoamh05+K5I2RbVUZZ3XkhbtAUc3SbFEdHmoub7CZ0N80ve
IAtt+6/+W1lD0k5MB39aNuR4kyktVvolKNYsK/orJoGWGghKxxdCiS7xkNhYexdADdIGKqZoPKBl
8GCmVh6M64uQ403gENYDYdXtQC4t3/CGhk2EC1m/Y82MKn+aqOpAFGyvE+3U7MIhhWsOYLCFIRo5
naNX/ENM0OGoM5yWzKzW8EfTTyM8WT+KQubB/h0L1KE4NxmJctmpKPLeKyG9diov5/+a5K/PASNc
TyWSrG7pjXq/b7hdh51sLxyff1CnRTamDxblb/OGXjbRQSdMB3VGET20mWOt7h7IjfhTCjmDL5SX
ugVF04ADunrulgHdF0u7lbTKsrgLNccOMFmh8RPdGGuXx2jJbNRj/OBMziF7XL9yNSqwxNqJq2oz
QNhYQjBmiRzy5zOeoZOFxKsJocwYW6RAFgZtQmA7FsAQrZ18snu4gATTk3dQ6U2xJsomaNUjrbij
pURYMy9An3ZBV5pdbZCvDZVAMGmJsm+mgsGobXzFXwVZOdjFtKN6AuW9CIiIurm/dvbbp7S7oQrO
miN3LrdkqZ2pVEU2LUgGcHyk5zkW311usDKCOpkEw+4nmwqqht9E9NGcnB7BvE9on7gsEVn0ZGLL
Eet/8QYXRnZrRH2ZhZwHVrDxmJihpMdVjoZ4JBH6KSnuGio8upsWAUt/0JLc6UlHVysRqA0s9ixA
J6FKbA9gfYntOgCOED+YgXihcNIGoq5NkW+xxUxzv9yt/QrjWpzwSs8yusA+XgLGfprwBd4F+Q82
kkd1Oln6UgTL3KVsIQZ8ihGxkjVj+ycgenTS/4Wl/zyAxyuzYNDeswmRKyiXCeZwRAqE8d7LiCjh
y+kQpco7cyVAFl1XLlVEm0ngi6Y27kJoAApaCJyJDLX9l9jEV7OsGMZ20qPKZ1d+CKllntGKenSP
FUqIoC4ZwNJ+sKwz4jZ3eVF9w9JNGcYqkaTd4PpAyXAycj6NSenEOze/KJOYhFyX0Lp78dMJDT+H
FOF/mcs+IeYCSM7CVgAm4XIex8WPaRQ/H3UmCWZQhi9Z5L2Kt0rHCJQnKdBludKETV8P429+vc4T
jPw1naSApBCulmWrpDVacpkM5FYw0nBKzeu8diOVdeeuTUnyz9ltQQaHmXPHisFOr5ZEZhpo49PM
i2lVHC7chAOyKBD/bKhvY2pip1GxEc/jfowPnsesBXFVv5gzbNU/ePoYs0/rG8b2/WEQHJ+XXrWo
nDmH58HgyRDrdgWGOyci4g9pCbFf2hBWLzXDPAejhoP3DzU5t97Q+7UYtCeCR0JgfNbz+SVdN22z
wmfW1pXwolwR9qhKOWE7d73SocvR7nkcpGil4Sc7KB+D0R7S9omvoCvf9ercCRMNdUgTnJhfmxJj
I1HvyzrgtZk9IvXdE44WRY+BA9vhFKWV3ikLOYZaPqySK9FYOUO+Es+hd8C7yoeFbWarOxQCdaGz
CXO1yHvEP7iPmCscNKcbUrHZBo0MEGmI8D813LsYSQ1ZCmAxTyM/JzFvR9P8ebaZ/ydi35Qaq+rI
PcnY94LdOMMkyR50XXE+WHT8Ywx6x4KG3G6aqW/Y/QtRXJfTiLs4Nt62eXWCm7xJfnWzMYcqPUD2
kY3UKQOahhM5ahiBe2N0k+cmOkRjwQ7GurfN0AtZlY/gGjdAsVMnivqGp58Hp7qXEmyui1LdXoXi
NrLFot2KVxWq29cDEMlqifLQpct2y903Jusyv2eigZ73bgoUIGMOMAV5YMRAGKYSQjiGYzOAHrlF
ezfr7aCblffek6hlqa81vfO42dEhiAjE4zGuaS5HVVi3vTdQhe5T6cPryiRA+RADso4Svr94wgkG
3USWGTpHAyVOgQfQZoHY5o3d/PVplwjKZ8y4Ug/OfmX0cSR4Yx7dVx2oPhOp35evKvCgI0FBdzWj
jUh2yxJqUq2178Ymw/IalOoCrdkJHsTTdMYEVLiOYYc50ufOdAKObySw/wN7f5/JgtbZcTgw5sn9
QgRMJDx4PKSmyubpBXGqzAwt4BTnG24VZkvko7izw7hTPgGR/9sVsOYSHF7TpOA7X8j4WZIBn+pd
/BO+LCOcjCkxDtFSbIUVmcXz3Fu9+ViPodSNSe76yWRPwEt6S9rSw7fM3+1KiAwUV8Nxb0UN/pFE
mjuF9eaB+TuskysjD40hWqLIKqaqkDizH11+9xziNIJO6slF47Na/nKtfvFbpQwKXwZgoE78nRlj
J2ryFuM8t6b+WJ56MMtixsRlHK1/3iPB0YXJUcfPFmykhkSJKVeBanWx9jynE7PdBeb5u1LFyiBo
8MT6qCTxXROXig/n9SGlombyLpcQU+F/n628J4gLT9Fuli4zEjkECtO+Q3iWaWmSlYAn43j2aEcn
sIBsGnaqnKx4Zy1C2QpnNfIO7MVR0XuWfhdzu34DBAqWJPkJOCiXLxK4yLQQW1gWMDW38pqCGAH3
CifxrbOJ+rJEzrofYR1ZT9zLqFbT/y010X6+78+VgvDmij/T5Yv3d5ow1ES2puOXQAIrOCzhAGW0
vpu4iifal2CobGHV14i0LLptLOOqA5bIj9Y2R2osotsDZ7T7yuhNwmFAP3yWlPvuIc/T+LCSn22b
vBrydLrACe0zIfvKC1jPBjqJixuWPT/RXrY+7EGq9wS0RkngUIT8Ecc1Y7/F1mr3z/sUSSwiSKj4
Ui0YtUB+enTtfJK3iD/xyLdJL0TDhTozU3jkKKaDF7tmFfWKQuDT4KkIPLdfU2QIlzo848z9+mvZ
0mhFkShhg3ZmOkcXjdBYJFhoSB18kBlpFihGmH7vV+idpiKv6M8HWFcrchnl9Jy9tkkQyLhp3apQ
S9yUWfe1Wweq4YrYOGiA5lWs+I1Sd+DttQWCjjOEncna4AWi4OAbTIQ2KxLaL3SKsJbaevHF7qlM
K65kap4Nlm7maOyP1CBM1bfGizClpeHsizRJidI9FOUpWMvxd9jkjQ7/SEFpHK9FgDHTcE/uOdDN
TG1eUtdSy9Gk2+ir/wFrvfxKob0VonobT8wAFJ6sCxvT6zKqCD6uuJnmap1vbTjrrTt0EeGs43VS
CTe/H3Ph7A1cDnpPKoijQv2KVN8yI9LR5I3PcJQmAIo6NLD5bNbjlhWnAz6bk5JrvffPGR4mxHdF
+nSIZ0deaZsFbvatsmqAm1wJopieR/1vmNLmK1yGw4e2617TCHEOUIme1meKL2RCUB/19weM9PwP
8zLDe7Ewp1FEuggzjVT+gUWyBka+p2gDeNQ+Zto7xKMOrWwDLkF0vhDBVrAC/WONKj+Q1I+gwysI
FtRCpfIciG9bTmRDaQaE703S1JDvRkRBfzNdIHd1ZBd2L4ADW4iw9MojGJjEqCqPhjmH1oN4ZSt8
4LJBx9/Jdig7PPbU850H7h6XRRa9w96Wzszl/WivXgRSJtTqIkmaELvUOE0ZODyEH3p58eGXA/QF
B4qiaIo56jirh1HIXPnrPtnarrbZZYCJVxFdzwR2Pnu2i+4yPPdf57OLbdMLC9wPoRiHu+UWeUF7
ouEJ1Fj/+pw8+BoanFd9pdob/WnrNOXK5rP4Fz1EyciELYYjT7mduh9MmPRbBcugibUG3M9MXVq+
Bb6n5aG1o2Xe87sl0mjalsT+8msHBG/2IN0h7dCkSnoNR9VqdvZW2nF3GvzGcEFd5QRhdd+WtlAB
rK5UR13BiycQSPBVG+/aHcJ1ctfr6PgYSD9obdFcW5JHpmGyVNws/7ah+UXHmMVAjE9zCgvt/63F
YKks7lsLNTv4PP4AT3xumhbzYuPziIOOgvrL895oRHHM8339uRmMhPw8Y8tg6NgyKPx8mHzCLmVS
wc2hi1QgBIYVlbSFuxD1uIYAVulsQD8fJ6GjeFTaV0Ar3FkTXrtxP0IoeLsqW2w6IUT4mVUsg12g
8sObqlb1WN1o4rvMSTIb1sUO9Qh7UBkwA2kE6X86D/RkM/OCbUSylQ3O8S9/Z7cB7LIKIy3ZZ0sw
5YHYCMZWAsGSrgfY1TSjkATeOvwPUKtV3Q1plPAjLtAVRj6OOEvbFhB9FsCXoU6SCrSHbkPFhEij
+ccwOnJvm0MIR4N/GieB9DZQwfMert6XmuC/4heDH7uoqOGc/2/e48iIZQZcnJ4GIyMfMqUwWCBc
QQ5ZBxe8vD8Mvz2O0y7z08WNj/kAWFiAV10jnvScKlgtTeBHDxVNaOihX97Xigg9i3uPo7klFWLp
Tj3kC/oz9NMBoMs3FDQEMJVk2nFFb48BtRwEEVOkOlP5cCF0Iia9xUxreuwkzGls9OwoQoxlxIWU
VHKPDbPvM/fQP7F7Eejc1REstvrYZfRtB0GSE7IZ7hYU1cB/CbUGVXmb8qXSY1M/QyU7Sq16bBj1
TwzhY+wcH+v8keCS+7jCtSQp2ASjWtY2t1yKpX/Gha8+cmfR4hKTK9jpVJVQUOsDYpPWi/XMRdSp
o72xzT/1Cl4zLmTLvxqq39erbWrw7tppLHlivrLoCqk3jrAV4TnVQphsu0SD9qFXVGPByHaHsilk
zGNxjqZR2za5APhtHzzT9ZADL49jRPzHDe2Buaq+y56Pis75IPHnbXTf9Hegz8IFU3cm4nRqsPHK
+Ci+U95/8/iZr0R88WiyHgvWv0hAYEFpyQv36Sze1pJQjk5eelKObECxVvfQ28LJEc8HIhS8j5JU
b0XZmxCu11auDwuLuGvuGzNmFXCWHJZX0cIHd8xO66KFh2Q4XQouQur0gkRG+zXTlXaaCxUHXnmm
mJvZhEQcUXxJTwvM9VlvQhTNI7kViyIsJfXq2DuaGHzobFs/eA9zzaaFbH63J8fBlWix+r2LCkqF
YGKVWVanJZMCUbVKQFxF0QEw62Bqs0PdUFmmlxW4gJnIJ7oDBKF2qTVBkJgzN+qPt2n6eqNVMEO9
oeiaH2+fdwqySSu04PtBBL5P9nN7rkVnHTB3vZdBmxIBfOxcjj87hYku1muUrT8CUXbMxP9tDTdu
+zhVZn0++2y1YmeeaJEdhQMnKmJjZjFrQSgxY4rgXbaxsyx3lz5quXtW/v12XC/VCbOcY4cdAOYT
KZ2hmoKgYPh4c5aBf3/mnIRgR+frFDZh8B6n4xyGTqM0jdbUb1aGWfNNM2W/ExRuM3nzpYsfNUCV
yHOK+Kxefb3ZsgX6xIwkNPDf9rpIxUZPhtL1I/sxmJaZLGXaganaXNBCwLgrZYOcK2qiyqzbx3FR
TIsmTQ4+dUu4w7YfL3KnkTlDU1bymvLbFJ+Ld1n1U6M1qwnYexPZbY1jeusUX9gpCvsGfXWyT5Wg
1g3e/tkRbe47pz+J/2D8jpJylFrWjFQqITtwEYJfSFv5sqlzb3cSADgq14URr6gREo/J5SLsuVqJ
CRKkD1L0ZTBBZnxvU8n9/W3lJnVKk84vzdWA5khhlPXHx7O1KBh+Y1d1GaeQU6cwyEsRDibPDZXm
W5l/tT4UWpoxoKhcyjO5AvhHdbKKsT/bfNf2ToDwNJFDKx+N63k1YJLrhvj1TpZQNlcRXXExEE0A
e7rs9ccS+PzlO2edoZTMu42ndDqD9e38+rcKPtKVGvQpPoxfYsqGwkeoYKy2C3v4Zbe3px4WZ8N4
GYmpS6c1wexSUugfHSdBVz9wj0i8JJ3x9m2Law6hDroxDfqpFgGa9b0Te5NPnRcheWfi3wbBllOE
MjVV/I1FUoUK+RAxebNRFC0ECTizc3Qt0HYjYENK5xmHsKX21vcRhi93HXVHnosPL9deOAzV0pfH
jgfSApDVOlkeclrLKNobmdBgDIljezqtYv0M0a5FEvTnswigwTkkH6j+uSwRwvLB9Md15tJsf7yq
mf9KBrTUW1jNoplN4pZgRd1YV+1jM9Xpe+2VpfXnR1z9kgfP6zkHpRlNlXwyedA8L+LFhKOqNZBZ
BPXDDereqyPSKh+oGdR6JVmod33ZqMoz9muwDPvvZl54STouKjnKlhcA7k8HUhAPtOdbzKEaQ7EP
1QW+9/Rg8JJYU8vCvSHf+K/ody6Gr8qSOkeqymPw4GDqs+26OsPVvP59b9tuW3ziDyGQGclU2dbG
oTSkQvNi8vBCds3x2idSc1LbizFVagrgzyoKe9c2HAplo9y7t40XWNCYxg1ZP7bbq32ZYQfx9DPb
0zChLBdv8C8zabKYqVxD5uTc+AN4R8ZVKjtYZCDJsEQQy5pLuZdu1E1zYn/49c4y6yV3z2gBsvF6
fTzaRP2yrQrdHkyaQiPh/aDoY+As61raj7EyYSwIB16t2MpFNF/zymSdn70+i18UkewJh8m5F008
IscBhpYXicj1KYrxRoS/7Sa5gelTCAp4SA6B5/Pal487LxEabc2HcpIj9rQL/nNE8kLTo60aBSYQ
NRwzpXNmQYlF7z4YXOUxxGOCh9v64DP5Wx9AGuGZGTFPU6u6JAVGROM7g1N6CMvV1U7XLmi+V0/U
fRFkJnBNdrQ0x2GZfUhPpRYzJiOQeAt9ksSEU3VnQ5hbCttO6MHBD4963V5SrCRIyjkqHc8NhRhM
fXcrsyRj6aYwN57trlx6UbfSO2hNVO5xhPFMjkiUU4kfSEFYc/2GyCfMAkQA+HkaeYMMK5TRwhm7
CpNpIGwUTvUAYZ5ogzzW5b7HiHG3N21iyQiclHaWXV+1a+AibVsnEKsBzNtlot8XOhKfyK3hfHIn
bD733jHZR7ZdATbAirtUWp4vd+gIiNspa6gaJgVj1yFe/1hXB0kOKcf6TFW5AfcswZU+U5AL6Znd
HH/4epAW32SIMdI7kfLXS1Yt1gIHeejBXplNGCspcj5fRrz8Q6w8N74rnO6VCK0Af9FVxR8NRyeG
9nmSFCpBbGQIrJYc9qYVqIeirRsVuLLvaXNXdNfSGSc1KAZ90DCpzk/IM2N7+kQI/aqhGoXP+91W
Tb8HWEHsWlsgBPSy/JqUHzoguOKtdYvJlT8cb3HBOpEBMlNFIdswSJ0wKtL3GFrsxcscWBymUhgQ
ViaZrsaloZMswCGDF6WMx9jpeXZCw03vol2PVcQsUYxbYRS92+HRlfq9zAtHyuyjV53rwvkjoGdE
/dc5EnnUpuNAxglo694wMbXGxKbv9AflsnFadoL5oSXw2Q6Wfv/2KB+CKCqqi5ppzltynFYdT7Ov
RnUXLM2KnoISI5S4OVtf2rF48FewGUBryXo/9EnC76ZWARV+KecDLVB/rk74ckIevf4kk8hjQ18m
P/2W5njUpaNjLTv5j2uLHR/zPyhiEXmJdh270Kaw5vQT7IiZeSiXekpJewF5e4aLASQ2M9UlMBiB
UAYU51okWuxDFJAt7E8YnIdQENon8WX4wmFR3Y0UsC4B4d8LF+oeN7pDsz6Khy3m+tYncEy/Iak7
ySosC+cEh0j4NG1t4HWoBJEJjEUBu+GTU0FGOsrGkNJPG3Yw4Aw1KdaXzBGD7QvfpOVPTLRyE3bl
FcwQ5bdMZpcl+AVOLjZRb0+jo5/PIVcU/f2Y6smTbL1GY1IZ9VLT7D3A9abiRJQqyHGljH5+2jze
YHivG0y9Jy+dlfP7Z6wCFmM3QE0CpBdvHb0wn1R22xf4VwOB7pqmgR3LKR1OIs4rBxtjLTPVuaQ0
ZJ0x5L3Uw/7tI8IePfqf+6jBpmOrxo6OlqrDhm1t71jT6SiFQ/K4uhyIlvDsYX+ihd7uD7eDvTWm
tQeq0EZD+NYESG9dpdR+bL5NABgE4sXjz+g5EVXR2gsyt/jM6rF4E5J/zZsK+NBXXd/Hqh2UrioI
sV6MfsEwPCd/MQdghuU9ERe0sveyAFM48NsQ2gFn2397xI5aorSaFuTG1LV/PK1vw03ti2f5+R/u
qWMPnnyLrN/GSZ/bEN8HfnwBT1WpJtP0gOx+LycunNPB46s1RuuabZCUUILvyl/3I0dQ5kCHR1aT
2+HHERjZI+W9cTQQeAYWKifc08jY19r0PFpiqWwlecaal9WJHahHvQL2VE+54bIRZv/LiJI0eNUF
p/SVOTIXycF09OglSVl6vDAoob8l+pj1DvdWgxNCVIR9Zim8YtLmTgFp/7i+owV4bnbAZHjOGOer
jNtYmXAtqkZjn4tEcU/LVFeLU0ASi30QNnaPZ9v0q2vafqmOkvDOhqQ+pN+gw+4BvwrejNwApj/e
DW523LAy/+AitG/fo26pmjuYr1xaRbfugkK20QFarPZiDMpwVHEYvfDBiXTTeTIWF/j+K3QXWN+b
Cppr21rxkEAJvRJOHkJz80OStGY2FRLQW5HCiKcOq/MBQbvY5p8/VhtFqgedDWtEoCKLVqKcX1jM
tIYskN1njg+2R1+WMmt28d6R5skpOM7TTpfL3P5PQ1qGYmSDKZ1a7IJyZhGl+AFf9tHEyte207uh
bg++DF0XHcYGDf+mVnB6x28GC5XkAQKbGy/A2BYzrz7PCTMNkow7y0fRnkO74eDk/lQtptPbw2G7
XopP+KpL7q4nlFTXTIRW9y0B8oD2NQy2Xfm9laDKemeUk9co9XyBgo0mikV3PQdBz94mGXLy0AZ3
79oLhECb9/peSlNbU1TaK0iFmTNVSMgSfOPLQnPNcTSCqJkEiGR0LI/x+x0LJGYLn8ASIYMG2CrY
e+9eY4FevD1Eui+io/jvxwkV3u36RrYB45uogiqHOGIaTpif6w7M5aBAfIl5M27N8f6cLNy1Afsz
Nt/Gry5JAIwD1GHOz6Gl4tRc57wKgFVotAcMQWZoIW5Vt6Q0nbFqEY05xpztijygCmfBGi/xO1ia
W1rKXZ3707l+dzVAxRv00QFxmE6knfJB+zvVYXuE1Mbl/eU52HCs+qJGCKJ/wSCkQc9fGG45400m
o54rj8x/Zbrt18aB0tbpq/hYucjjRbmbN0TpJ4JC8yzkHCtRds0UbFKtD1gi6hAKwpdwHX2Nl1px
7bQN/U5VjIXS+XZ5m0U/M2m9hh8BgYyW4F+mbIfmRkbtssYlc3leeAiDhmIsmhKQjd2d90kNWeH2
2rrfPY/wGjHAZCmZMpjx8NC200gYdxmbuMQRVQ8YoL7mvpPcFe4AkNgQnrvFzdXmej7JXpz2ugPw
2XpC49KTM2TfcIIsQ+sJVWc/RVfJp5ECTGVw8164K4vaPPWme90B4k7zVNvBaYVXVa0oQx762afQ
uxkUDvWph7GCMVloqoce/hB1s71qnYmgYd7U6Id8AOlILVgIsh2Ya12N/GsBQOuEzaI8tht4C0y9
D1P7TBF98Cc6bqYYTh48cXdGVnVIboGUz+S3NI8c593oobN/AoGsj48VjcNHhZRGiiiQ9+qxQ42f
6X/YKXEiqaj/UOtkZ5ZCPMU4JCziXCZFAl5QrE9/Mn4p/PBvH3kSNRMyzuRLzYHvoehsOxVWe26h
JQuJMxYtQcN1QfXc8VK/oYfJLCfBHh8kXXfSG7TDgWHexp2zc4j/S7nhzWULinBRCyK1BC19dt1Y
5upA1GcgvpV7wdRdiJA3A0ruRgw/uLnHFcKHUb3XeJwjVTAl/7MSsQx07+nGxvICdmAqQbz8EbBE
09+88spfOF3CM+54llX/vKAkszW3FcJcRLxqAQedU8ov6sUULx/TD7SriOwpadje8LYKCU5H7wrI
qwNmHrXbqFuAkAbgPgCYKIogkgz6vQxJ5ng6sMFfsc4bGwW92bKkysx6Bewpjl4/xD0OtxiP7AQT
i77xD5QeIB8XN6Rhwaf6gzQJArF4s2l08rYwG/cF9+8OAs+L9rnPTSazGWiSk6G802I3um4CtpVQ
iXWH5VEos781ScGhd8cwdREdHcP2lc2UaVEU+pbOCqCEtPAnK0yRNwuN0AFFpajjHo/1PkhroIu7
mPj80oHxvpL5wFCfWTgz0S0B9ZM92nO/YkD8NMbualdadhMDdbVtbjc7nN89hQxT+G/S25zaSqia
y2qWl9jJtdyj1YQfJlbsZ6DgF2Ahfja+cwul8rvfg8d2u2cu9SMQLZvKCspdfSmp+XpfDDA582fF
2ZwlMqtELPicylsH+srcuJ2JUKdFvXa/89taBI2g78qW9MLyMp9C51ejoVgU7vk3z3gh1+Tb9P6V
ZAgkhEnSIBUe/7kYwzJ77dZOJjxMT0cIRXFZu6YlVUL1ENepd8pn98mafdgd1J6LwL+5BGSlz5lX
fXgmDavNVhA9x13ymIzAKnStA/9+2OVft2sNApFC5ZQ9AJbY6czauy5X5ZLEMwWnSQDcWP+4ft7V
j4JyANqDhKu4liMOnIvQfauguC/gy9erWbDMP0q9+nD1LyXufrsxc1383QBUKCoAwjMtU1VOn/+J
+sk23Dv6kV46Gora9F0UFIe/VBL4GkN4joDrunAGL1ZTAdxeRJmFVdrzkYc/q1QIrYb67IkQuvPB
bDuzYCGow72hr11TOoTGuMtIbrwmhbUAn1HMHoQXgxP/Hcrpj2yZcXP/O0lhMhkZgnVg3YBkeMii
kWjugyzFsc7ckqcA4hxyuIA9sdlH4OpO24cdMe9vl22NgfQ2uyOVowd3qFEYCPwMSeVbayBqdx5u
fWY720+Nxc5o/B7z0zhkpELv9PC641Ae5JmHFzxwS7V0rC7rQBwiVGO4U9XWOoFxO2iK9DIeudLp
Lw0jkSHNwA1tarvMESDWkjnt8Qo5EgCFgUNAPbd+Y0f1rHrbgEVG6jzr8TH08KJSH24oiO6bV5rg
oWPsrVKSetGCf6e++HtI+nrz820Lh7SIwvEyrVgQkF57ZYq5tXOu7E6rolHCeoDBkE8wSwJkzdnf
Rt0jW7IX6j3NL3Yc5fFtlKqtrd3I6fs2Y2bxsYUI7IPw0DwyB+OyFR2vKs6+vuRO2qVlXkAcHGoW
L2YOc4dy4Qcw1CnSqhVY8LuWTCZ47pCA3jjJ5WUSX4j3rCXd2UdiikLgXP1aC05Dvrk1BQ4sZKz2
f45MrK81UAhil8w9LfziRo+TDEiHpC50sJXclqU00MuIzNvH2RyAUor3e8yr2BeH9Qr6116hx8Lp
1e9T80vYFUvJBF/x8ZI16lW7mgmksYdMhwwKVPo4zDXWL9i1s9nGEEz5OLdrX8lslt4dmlo01GFk
nht2ix+91kwbtnMQ3YZSox7jW5mctAwvfcYKriL97RrwPvFQXjc/94k1bc/m6b454XsVLfce72lt
+Gl6QWTr/RWijfzJbVZZd6cTgKOy9DAhFBpva2ifrLMxta/auIW5axmVGIL4t+SAvGlNrFWM3XU6
dxnDJ1AWkw9Gt8JGXpYKInlziOXWgkKgfYDVW9bXjeVbh+InGzxiotzZ8FWh8t0KHDHr/EWS+APi
QjrbkR9eMwF4/W0bWpLIUUvo0L1bWzXzLcNsTxdii7mI+vDa4gWgdIb7zXcDUeFU+VlgQokxdUsQ
3dj+YawhwJ2OSgnfTOltQm6q8OesiU4efuQ0l6muciQNDbhaJKzP2AzjglQ+sYY2ZmLMkW7qkOIE
FUgl6kxTBY1Jl911MfKXLZSOr1Qllv2oqS8hLV7ShYdX1XdZVaTsXoAwU6MEnD74lQXeLweIv75V
x2kHDEOObyCBceN2sr/STF4XWlbxRtkbADXKCybDVyry1bNZcvHYwPKrr3Qs/tnQUiPglpzVMACU
hZ7dkCptCxgfUhyVUfR2sFZe0bZFJViJ86maLTTlAn1GphQUCTBqvcOg3v/WWhkfzblIaukCJvSu
gmxd0hTMT9x3E4cdUJ19Rx6ho29vjIIlvEvR6Iw3hnbSbOjGUX6tzb5TVRSDMAQDYt12BxxrAIB5
Zvq6z0LVIyEzlOvCmc6VuwY5RXYuuNMlpHIl+4X55S9NjEkhxBAAqYrGONYhLXemyPfM/vkMD5hB
7vp+Tp3WrUv5LRopW4heZ2mddDE2BZrAq2MEelg2KE48Hur8MWDQcZw23FwR1QQkeABAUT/HjYOR
3Wxc+ADUoEjR16YAlnc3dxC6ASmtyMJv3v6wZI4FgLtfRH2V2MnqSwAVVEuJ2c+l90B5RpApXbJv
fuMZtAg9H/1VJNBi+bbvB5MXSZSHnkIOc7XKGq+7xFB2y/Ra9xQ7t/LqIcwh0C8C+UZ8/PFIfHLM
0oPra1KNzykivZ6N/NFIfVQYypA7yoenBmBn1wlpXqITHk/narJljgFMJHK4NbjlcmhbMVgJd0GQ
EY237kPN2JwyuzCFvBOHTUjoBnFCoI5wk+zuH1BbhHISjedKJsp9/w/0TGpZVyNf+RBqm6rfJibv
X0TiyKfIBItbhgwHzLpGnFUeNHyMy1uxpkqKFAV7jhtnxmP/lCnrnVolwcMSEi9LsPXAp6t5mJaw
sJB0LK13XeymdVDQepYRzAJeZD08hnugAwiMXJU7uEpsfv/8rV0bWEZfwTHcQ865yc413QdafrtE
xNumLQrAwmtIRcblV0GKGqojnGFzDyyJBz8b20ACzh4flzz2Pw+I9pMrWuL4z14XrwSX7chZ7otH
fD71tiWa9uJ0pqtWbZBY/iLPPYZ/qFkVlBaKPUXvgikY5Roffpd9NRp0fNAdfeG5kG4vRvGhG6cj
qK5yVHYrBqahsFAtPEUpmRHbBTJdY4HIOzi9zesOJUAP6oUM5/jAZfEECuOgwunwMzhkymgKAHlS
Kue2j5ldPz0fS9Jk+MgjuvnM1kzgwHbj6zUU/ewWUKpqTJeJ/OUV2mWftEiy63rT9DsZjmtn7fC/
u+x9OKQsj+4XwEdqGyU7NGUfGCgI/MKW0bIAr3Llb042ntT2jrjMSn154HIZzLdo2H0QUz3sLlrV
BC+lkgjfglcVvzCTyfajFi27obkF8I9rdx4+zxCAj53RZ8Q3/Jnn/ITB8Fc0sJlb5YOIRniB3dAd
7aRgu/jin75dI8Z1MyzoY0NKpGg/+VS0aX6dUP2jHFYHAZ2tVCMI7svPtTyunDvFU72GPoyS1lpe
NhIZbYNNmeMNutcfqcx30u4/XgCFUZBhIpHX7amGl93XEp7dqxg7AYFQf+OySwbc9KNAktMI+oUn
EWgF5s/b8hf0vkweYH8gOFcY49lHXmSa/IP0TL/W/5lIUlTqtTTCsDLoRKul5Q7BBNJcaup1ZmiD
fqShuzd0aq4cUo5jhmt95b8lzja1F96q4YDBRLz1qVXG1oicEEI+xVwLUCf5Lo+TSEPmDviw3wmT
7VhHiS4xUVwYXo4d2F2mVP6rwujCq4XO1qHTTMlEgf8hz8vGUqBCocCpjXZTxn5/aqSXffBAMFPU
bImp3NxSXWWM53oVm1DnuFYGipBf56nwtl1ID2Yf4sSulcBW/dSMR/Y/q6M7/KDejW7dUywbLnb9
TcSohf6sQSs+2lgcuo50Of3RhXTZJCA0shnODjHADtkJ+7MmTuv9AsXibusOvsPtuObL+WpfsdIX
k2Zm0Fdbbl/qu+iDT9hrD/8FsOc85gL4hioJrEn7QJ0ed96qbV1wIi2dooLkyg9HyU7Voqy/OFOV
ii+Av3NWrl8B4/e1QhgGYjlWYivl1DXzZ6FOiu+qLeb//2ArPto5/bXjqkPDOKOw64xeErdFqjn5
ireM6cJTJKtFtn2AHh7WlEo/wweZTPYD0+mLTk1XC3wy+c2+Zh5ZlQVsA+M0I3zKkRfCfCZjhT70
RbinPctYK0nkAe5Jzf2uWj2uP4H7fkbA4zeLvvJ1b+CIc4jaiiGCka3rmCeJdrnvQVQwHbB9Yh8O
3c9sqgxJAK3aKF+4bSoRv3aZhl9SWPKkW+4RIQzYaAYb2igCNtb/RJVSNF9j79At96p1FSFqLtSV
I6eALemM6UqPahIbli+Q0t1b4/7wuMKFlJcxuv7bpVoH5gtkYDv7Qer587jVwOHShdoU/N0IXKfO
5RrWVUJ4T+tYxXxPvchwhEjmgvF2pgEXhvVcX0GA/HYRiyj1/8is8a8e6W/9Ag5tPZuUUNx1Nzu7
pGSmd50eJa0Aex5pOiOUpjSBC652TwHj44wy1Vxh/1Rhv78JnLtOLcQ+G5GXzgROpLk0bM5gcQcZ
9qlRHCHvRX3OX1jiEVqx8k83za/PSMGZ8wElD9/jvE/gF1auWnIzV+I/T9MoCWi921ZS3dGBUuJF
PoC/AliGvPDwkEix385OfLGDsfZtHV1Bj1r0bdaS2vLag0hYVQaI1QRo4ao98b0zTOOZQJK+mQQs
/jaTJO/gxzsb0pZ+p4Ocf7QsHqkKLrGcOu2uomkCQrx6hYoKxpYB8+5myQO16TTmM4sinR3U6FZL
UpQ1g8Cu0KFkhZ0y5fQpBoqqR62Hxi40KAXK3CTMd/UX0E1daTF/9Oh2q7/Xvad98xssFRYhwBga
ZE8odvoHTFzWje3nLiXb1Z5sjUJW8ROer3Ilhvskcg8JINf7GACRXjWnRZ2ci/x5s+g+CU+ZjJ3k
U6zeQToASFomtpJ11mYNxGc7nKN+L7UMbHBtUX4dw8q0WCospGnfqEvt0ERktB53rt3fLB1BKGOl
KwTzHkOtBOtgLs2Q/qPaEXLmslNGNrVhgwhQHqsaeBJgGhoVJBSuh499tIhB7AcjPMpeQfaDNkpq
utJwX8vcUYLbFTjf2yMnGeK8z9RkPgXZTKy/eVtD1D+PVmCW0ArovrCY1Zs3bahtd8ooEY+fO/Sv
OJ9VMZ24/wosVv9uoMhxm3rAMtkRfmswB3naJ9o2ptAtyqSfQBzcJbCTp9OSEcJHcNTmdOHXeVWc
mCgaOb2GE89KrfQTO6OEwf/deDL7Ms+1DHOYBRytEUH92nrOSGnoOvWzgFDbVK7KmQG/TqUCgfy+
kIHHW7QqQJhYUKvxb1gOhXo10CmFAnqdxCqkgh5ED8wgDDyv8YW3TDGibJ3K9qAMrlIr3eFG8jci
r2j3FI+Fuj9iLQgwAYLDUznqAwfFUAoh0NQmdLljJsk/YjBu8Tl+YxYnDxPhcROX+hCZhj2jCGM2
gBE2pkSfhT1QoJID4tx0VXLToj0RZohjF3WR7TDU4D12C+Ju/jp5CtoHvQ4G8BqCPB2AManMA7Gv
NJhlMgViV9e5gI4Gv/dF7xBpVHLMSZqws7swCnjYnGcTWtNI5ZicjedfUvby7Ud03J3lhXoiZQxY
IE1g012naSXcV3nTXJwASKFo3UvOoXxLCyc6i4xO2oSBpp9ioKb3rsATrOIDcxZ5fkKlCq/J9WzP
DT+XVFE0L+4/k4U4EA/3gf05q34CivNxtnqg9sNGcK1rQYAdCJT0w1suKIXh7Snfes/BuqajIqbJ
eGaOUCrKZuFMOe3/cClKNx5eP0j+ddUwtxawg5Q+xX+NilLaGwCh+zYLEu3rxlTqLOmrcQYCV0qF
sZVXA8dwoiMRxNe4hPyU8JN0YVdnm8MZOa2O0gIENhtpxxTx6hl/+ZNDR6+jgtl6VgjZ/+4XpKoz
8NxA8zVsP5cPM0sHx58QnbDsLzAHJAUVqp2djYp5Zo9eze3qBBCO33e9iK1O/ZtxTNrSwT2J1Wz8
XHwNDDxT4XKe1X4dmuNu7uQdGgcnus7KWoXSQdMmRj9hqxOWRM1TbFcdzokEa8Pncnzi9osWBYg+
YD3JUX7FODpIy+nbQbyksrh8Cdq86AhvcZDyFAHZqsFQuBotzSDdjjR9A8Q57wTmdTwXJx52wFvr
byOv0VZltfaD8JtlF3uUwZFbgnPqfmo1Ayk66+DUkMIIFeqlLtnl4swd8LMuZ1ypf3RIXNQM4PzZ
asJOimnB/xiNEvLeord/EgMPq2r/Uiismzj0be7z0GzS1dF3f7lKFuxJHAVY1c/rBWhDsat/dfGx
XbF63RR7T3Fa3uWlyMbG8mjnBu2W2zVpus2wp1K0tbVo5c+2FqHV50tGfYWTIn+/JoA0YJ7I4phA
SmQ6dcHM1ym+9OZ5nYaXZ+y45UzlltKHLeP9EyPNYpAa+G96oymvr5DpZMF+ob9yzFoghB3Ao6EN
IJVLi3GbtBZ0z/pVYCqHYsuJaqbg4Duf7VocOs287ahaGYmbEWdQZjdQc1KRREvMq9UfdAsRhtEq
niSisdijmLV63rEvvl7H6xzFnMOB4ZAG4mrmccaOsjTK2dXqqnbqWKuhzIVsQUJrY6NuOvbdUD9K
Ndq9wchy9+q3g2J2cnTfCHZO+DavuVpGLoHsOLi8zzEfO544AjRQzKu4ApRZ13ZPzTo9EOnaklau
69x44eHICjR4WwjqS7n+M1mxsX6nekSGKAZDTxKBxgS483XqgNauaCBrghEAzmna+tWD967iMEvW
InOi+mxnLarDt1qSBPEAwwKsskuMFsSA1xZ0f7tc1svszhcf8Rc7I2+pzzrXgNVYWycACKJtrfw2
yJULxceqmKbmizEzqbHoYMWzDNzM5wWxRKysAc9DwneOPm32UGnkfcx592L6xm+KYfdHZn+GFQ0Q
0ujSQw8b+kdt1t6wRwvC9+l7QYmflUodmUS9WIW8HNdsJ3ui/1tt8Crj9OQJnG4O15oavBvd/2xg
TJh5RaROZnUTIvh1cGi0XjS/t4dhugExnkLwcYQk3qICCs7vJ8VB9nV0JjDQrtKQbdcU66D7oAH1
LR4CXmrYq6fTz3XsP8LdGag21KNXKfoRPTMC98NUbY+0hPeqNWc1D6TLe8FHZ3GnGyh05IGey0pI
Ns2i6KQSVmp21nFc7zOlHHIbkcVh0bMacJxOstp0DOmhzVqcjKSqdhq46W7Uw8a/uxkpdU3ekIv5
36/3DCxqvYvSOn3gkks1nnRI8/lBuR6Gnax4dy8QGWeVexJnSXqvjiXBPBG2te3BDNx4n+7qKRbU
D2NB3K3bq+YypDiqX1R8RNesnTW1DtPeid2ApbmQZBu6kxuog6oaeYNxk44lpkzryjdffbxzpeZJ
js69i4AwJbPmSH3qSqbwIe19DmPGfsLpJ9UOdEBivBUzZWIXlERWCLFb/hvj+gvkBG2Q14L5xEJO
1cE+/ZHaBTGUjwTLNb+vfOaMJo/eCZCT2ov8Isho4L7QfSG3Itv+OphG2tWkqhlkHt8MFRUieP9y
FFj1SQWwnKUUeytw/B8bLeCHRngGXGiWIqtJ+U67l4wx6DDUNjK+Nn6JbWtva0awpv/MQG4TKyhZ
TbMYVaxsoyJJr0bnF45imK8+nuYGhD3FivnHcIclPQYEep472PzU/2vr3jQoE3M9D5QDlrUC7agw
exxlMrUa0RNQePx1f3lIHEfY8mYLaEaF+SmI7uaQfHElTMG5iiI/YlDSJG/ZE5fuVZ4zoZTg+onQ
4TI5BauFmSiKdCYc1BE46f9D2zyCYOmbABSdv1UsaS/g0nU54zEEdTmcF2+XBJmLEG1ydil9tcQa
WbxqONnaZJAIQsnJVUxcaZzlEVWeUsW2Zn8VbjBOmdl8N4SqMblcNzipZ4JiIVjvUEWn0mqr4ijt
fNv7nmOCG6Gf7tftWBPbWDCiyxhxtyaH0IlGsptsLI+yrYL1xdO6bBOMAEbMuheooR7WelxkCtvB
mLboJUMwg/Djs8+gPs90UNVCYdSBFURIuZwyoiYZYKnoq7adsOO6/+KbVSOfJ2H9RUl78+J/kEnA
0JhgZwd120ajN5otS4hK6+DKiZstm63REY6jPU2KAgyUjJ/qM6VRh2m6pefcbbwayXdVU/yMpzZH
oEHJu1QLJN/VH9LC+kLsF8h1eZvmAEJYXmczUcAB82CDxV/OyH7YivCzAFFhG3OMBAeOb5HMzstN
yfWo2X6XW0z16jVcQ9wOrwB8xSdbfgPHGyG84HdHm0sXbPRbwse3Xa7ZXxFqRqJYjdhHDnxEASDN
h19T32JE045i4GYkYUZLjZR4VwarH1pTGNJg0f/owyDfGGK03Uwl1ondbbGbP6r1KPbciTP+dvTk
erKZze8j4xrNYjDbpyZKh6qZ5xV+WtPL+0e+OUIxcHJJ2PS1HmMbjZUCYIKUMu4v07XD7azOkOu6
ZxMjtrKIDZFyIR7OvuC1J8kuUlxZ4Ze1tNk7SOQG239MTg50L8laEG4yQN85OsLd0iEHOn/rDljQ
LPC23RAIdQ/lmdWRK77lO7K6sZsEgAUrwnXM3XDYyqUx/lnXmiE/eAr6r1Lj7KR6wIA+QLrIL8OA
tSI0UTEkD+fwJQqi6f5EAXcjIF+eoQVm26hth/M/IRmk/J6pF7egsUrKZmMxm/qUDr0a+8cA7es/
FmXQ61dk3x0gnrU34fTZPRLq2cGR2is28/d0fxpGN62KLOQ3UJ7kxrn8rNcXF6BdZ6JQd/fF7XBY
ojuIF3ASNp4bw32IiAtBuhPgG6MYKrlZ4f3LZhxrUGoPFpbPOe2Hb3TJ2FRcpUXkfQKYZL7ZlC9V
IgNpWD+Du2xWCSgwcuoImm94uh2IMb9sSflZ1a4ab0Bf8+jxuMgPAzkzcpDYqx+Vpkah4LiH/G8O
Nl8Ben8940S3uy+3xtMcmvrsKv1VrChLnBqh8sFC0l42r99h9M6cvdCKv9s7rEkbdbeECyCOrUq8
sA7LbFe+yhlhawAA9HA6Aa17gfwiRss04RPCChigJNWzKF3tp73Y5YCZTzak/Js9W/ntk4GScKhE
J6s7JKp1gyFBi4kMX5Cbkrkv9ZteSS08jOCTYT8oIqBOLFJGEuZMpsGI8S0EW0kXJnIdwXfWWYg2
0uVTyJY1CCzhQh0y9UbteeIlig+xgljIQk3HqahpCiWXI3ad+FSbSm/hs8XavIglC1JldFT/Uhf4
pu+tXuk2uyEniDfbI6VhQ84n3AM+w5Ay016fvO78x21u1txtHCJOH8ul4LY5ekvqS+mqoD+dIstz
yWKH23xqcmrpdIfrO9qnKoKQXSVAcf70ozmGiu0zCzyNNtGnVOVbfGAc93MiU8GOyxx+euhtYdxc
7yVYIQFjgT/wNN9vf+mXVMwJ3GuQdasznBDOrNt20Qvzl8xNFpoB3K1hSmlKDPCHgBzqjMdgQZTk
R4Z5d58Qn33HJfPNei1+XleJXlMbQ43eI4xGbtSwsFWrTWw3P2Fst1q6/s0h/39fUsD+99KOUEvy
YCnx1Ha3CjE6eeFEhjjAcYn4tOe8i9fNUbYJuRhm71vCwnWz7auhM3HGzfFQz4WKnA5b2dYv2ptv
jKgTUhbqjjNZYeK6epC7I6YaMsKwRXUtxMf8kfKU7zPJ9o064091fSafpTqm9A/V8npR0VxeH4fv
uS88T7F8rRzc4LEWk9GSXR52llZ7e6IWSuZq18jokNFar/M3wEhIXbF2LbyTzG0Gg8a6HlWw3Jc0
PYVlr1XUPNaTO3izTI/kGx8pXwCqpLb45qA9N2nBCVqf0UcqSxYQUEV4+8vQNvsU3EoYbViHldlA
30t5aabngLXiCU6Zd4+PVM9/qEeqAWjQIGx2p3WZ98xBCGYFUhVSIhPpMv6tmSSbVZUXA5vTsqnv
zMxuxDbSBBgZ2HjoMNy9ZYZUiLljIkbqkeF/seZbmzGwqePB6Opid3Ut84Fe22FW9lzLJkuXcexK
l5wcw1PlJYJvaEhn2ze79mdUI6TFupzh8JON+TG0qYOvnNMdWG+tuIOQgrRcgnqjrHqvlr+NhCN5
c1s0XMQTNqridWXVNwuOCPBJppHgJKegsZXxJC4PaPEEYODfiLscDFspGu5wX91F0JTdqMHyIYzK
uCJiKCQJq/niuEplQR8rSPElIE9EPugG4wQVTEfwz+x2drButwqEbxHNAL5SVdh2GtWgD+Bdo2Yc
9uHJfKzRS5krAbQOrj1OR+PF7xf9L0fAHQb/HWKs3kVt0VnOXC31LJjpI8q8kjQ6gh2z+XPjpAAU
1+xJbUGO57EzEkRaChQ1XnVdkbrjQQFZfTC0CMiWQx1bjtXsFdvdAhujaOmSN2OyMkI5Kg9i6OsO
+HWSHOmzt1fU+X/k+Y3bw1q5AqCsvHPrYA7DbM+o9bdNTKpPxebNaPAUJi9po/B6sUbaqHH7oaBI
cjNepC48UQZg8xRHmfKdus3EoH7kKhBOWKBINcFFWs1d93/UiEBCIr9ezngxmdmKXotzbbbk2Q1t
GO7YhFWN2Bn/TUYC6NVl5Nddxc/GlKYeS+il+lFy4ARe4Dz86NUUGVpsrACc4B9Gys7P+9ppDykD
Ggyag7JOy0Z252tjrDnIw99zNFGBJiYLfI38qLoTfXqdCwj/F/5elMPPaflsUSz8gCbCM39amsQo
e8wDwPFsz+54I6awX/vm0aDU1TXwy5Rik/PSiC/+8oP10+ywuNw1g7C4qc9Y5xX8O4Bcm1eP3Ntn
2pSKI9A680PWGOgUlH3V96hhLWV1RsvBsQ0BbKHIDKmaUjnPQkHFSZBQ/F45PDSxVa1cBHXJuIuP
hDa8xH1fEaTgBWK42+YEI5RhXKLx1h+Ebaoy4U2MnH0c5fHC3erMSrYi8MdVIo1IET5pUeIKR7AS
IK9I8uYv61104yOIL7s8/IYG12dNUox2Cu6P+wd7add3+ralJz6i7SVDVrbrh4nJo1Q8WyypLRDy
npSu0XqeLkzcFcBrA3BPFFkRTDIr/l2/cXrUVkGnoE2u/LkEwIzd1WPHnPKCGVc1LUrvfr2NV/9s
ZATM7TERPA58P5F9JfYakNDIrWD42yNdt4do7fR7+2f7RiN2R9EYqSDNUICJb+NzNddWjvt72ycQ
kh8ebBA7hHKJhWOcqr/a+RHIHLuJmfkk3fC/PnNJTOb0HzbYYc3CsZi9ude8mfTkCTJFNvK5ib7w
1SteiHxQ22KamQhLu3Iwos7Eid2+c+0J1MY2c7X/I1gT08NWWQMsURhIcpdXbJpQHH90EtKgLu8n
V9KTturS/vkmyfRbt15q30jPS3Jxq9qTEX+rYrMfsQIHmOv6Tty0znogUYt1hGVV1YRMc2T9zo0m
aqUPBetZLQrxgE8FcqVrwgfypUM3zhnGHJ3VrFwWWVdgKr9DDX95cvR6tv0+RkIte4ABWo7MTN/G
wnfqH63Vp+UjNKktXhtuqQGKXli/+bzt1f/t+WkHvfkzjkbrcgDQ8MuBJBSkC6IsYsqXyJOeKjgd
G94cXjhAQfEE+E+4QQCbpqOd7vv4UXe9E72z69S5FGOcf/l3q3aCd0iFxKbcVfPpkHI+UCMHP97M
tSDRrc+CGq2HWrdJyHMPxGLoSsMXgAKePwgbddlaq5PJf28tdnTGFrTxOgF9Mb2+oON8m1L2AJEE
4Cjq4mbm+K8o1c0s8OnQn3+B7sYi+rCYm1sU7Yn8EJ1Snmu5Ly4PeG1Te7yXvwppAQl0DD3+T1Gz
QH5rSgK+zV2ykl3/gAKXl2jOd9AZuAKIcH5rTNzbri5ZOgM80fre7//szMC7C74vHTleVb1Vt9oW
DR35HYhNtzTfFmXbJrbNNgfCy2WMGdPNOR8H14GR+AJBbTYCJn5At9WNdh+ccEVz29SsFmVKIN8y
x9u6Z9r5nKtJ2IWgqYcqzhip26yzQvy0Zf0kvosgAZ/0laT616p3MqRNBP/4k8NgYyXLez4hdHaY
1psjkMUDjurlWc3Z/39eMOebeENV5DdS3gu5GI2+CeS2eLa7b1zXYZt7FByUSoBlxvDEIODRsm0V
o7ugWmC1L7jpT5BbngUgLg4iZDvnDdn+s9KFoM/oFz/Jelngvw1lzEaf+wJRl7GH7PgZFABm+WkB
GmjVAt1nSLqpp3BYeriMJXI3edV1FwIQJKL2kqo+aFy87gV2+xm1h/+K2faF1cI/OngDvCc9W97Q
r41SQRA3FRswcK9dWbSCGIf4awvOE4i5nu05o8dlfUBWypwn0WbcWs4iKWmEnkl+rRRd8pGpwXjI
id+LVG7n64Y7Qhj1PKnmjAVosW9yK8hCs0yvOTghVBxB/sJ9Jk2DX514zKv9+Yl4lFAkz8wmOrwf
kBXXAWQZdGQYM2CVe+vyTjZ11OdGBGLdJyI8M9OG4ZSsbQ+NmUio+/SkebjusAXeNEJf2XByu3sr
OkecJV44GBwtBSZnx35EltnYznaZuHmKjbtgT8VBN4ZF+mhXQ63D/F6+sYvzcYSkXX/k/M4Sxopi
YYyK3/CcbIqUxH5L23j7UPJDLLZr0uIf27N/lIPaYSKQeA4hnaFHN8RsRYRw5ic19Tl/txMHUXlQ
qVPNMvlqJ2yShtghKISj9Dr4GmgmeJj54wbOy1tw3Z63o+C9TewJZKK+1/zVC4TYMYa1BJDRD1sI
KYteP8SScDldD17dteS+iVVdut+Bn/i4DC75vUSfRf8fVjQP6h/AnRmgi3fx0zWp8douqYSWysy8
pBPqxwkCijaLTGzTEzgpMaPtUZmEUquGdyRBiRcQPrtq6IV7Y6WmQehq0FPqVzt6QhiKcY+ujFWI
A6z3D4zpPbaG55bUnGRJYDcGqJ+IyKrznETC+mEvQ9VN3YVO6Y465mqJ12W+XK0zoise40fwqMX+
+0UR2+f9a5c3JTmPrSqwFI+4Wdsmv5PEMj3lNOpMZsYZMnFchPY2MAsdXGbKrVOHqBPTgSxSISAo
oUYYm71Nj5ScKQW/GbAriy7Ahfv1Y0IajCZQa3P7JsiNXpg7WYP9Ha6lY8JwQbT9X5Gq5+uhjisn
+j/YVY58m6pGG/JcKLXoeGv5SzXNY1nPpST8fVK71JYUhxbTEo73fMhyB7zm4pqXoIkX8Lh7DCSk
3FXU+ZYM70Bxlk+L83EBnz8NLZMVnm8I09SYNbL6FbJ0RrRiglznD/5idAbX+tTNN5H7f5LReMhc
KCbwjihAL32gKFTOMLZyILiBYuCkn7ZoqUNfCog+dOMFpwoTnn9tkfsKCF0ON+Ij6n4VuBXr+XtP
HxF/prX3QnPT+6ipWCwcnDIN0obR3v2lD3RFsdxuA2xeNebeM+x0pnqBHcRwTyRDxYTJIc8BQRlk
Hrf1hNWNuX1PFeG3MaIxCNJ6FpzYQqFW+oodqNDN2t4zg3m1W+DJIJ0DT+NkkNsBYck4Pdqz8Gre
oI0NehWpqSuni9FPi3dzjGaiweWcx+3te3OK1vrSWvatmGL5yjWxupGG3j7s4bkI7yuRTQGQXdxn
FwELrCvfQO5j2P04GdtHVdD5zcoqEZTZfkDnU8XDM7MBuQYgb9A5Tmllx7tJ+wqg5Bfylf9ibShX
Q0+3TuZaJ1EZYiPaJzxpi+ePBPxLQ29oA+3W34upwtLjSUkYq0QpeAnSTMarJriFqV6E9Ev3McPK
N9EMvcU/J1NntjFb1TdX5mcZOj0GluwXUiRSt5ZByjDM8UpTEvsKMiDqma8NMwlJTPTNLv3bEsfs
Bjya1eRHBoGh3NOFpl+I0/Dq5eYK/Wp1dnjjylgSdm6Yt6t67HMKBbzwNt9MSnb3S5wG+RfGdaBR
7xTYvnmmYxEOA8bfO0ER6po4WB5vUUKkLyFV9hfuvNZWmWOT3B6Yi8aJbmMe3c2V0IdS3nSXr4K3
ShuN12qhQ/WVfDk+sut1/l+X4iZzuk+4QnUlhAPfaiVUkpb1gStZc/g73BUfJkN1OrRIwyIh5pai
JncgKdyafdMelfgWy0R972YgrwdE1fJo9/Fr3dJg4zGwp9rWelZILgIbIPWflk0XDoFQ+e7avRsW
K5nkxjYNm5ZFMrSXoMohskkc4l49CsHW1stlAzzZOHQBKMFQ1RoV+XBA8neXJX3uGIdTte24Llh/
tE35rS4dfE2mjaT+YYDVCP4YwtBs79zNVxRrKjshBk5se8e6UsORQOLaAlruSo7uelc1E6URvDcT
MjuXuGYZEbxJAgejBI2MJGgDetepUB6XHhPUZt93ZSPqKw+RSC/fE1zCNkFeSqmJ3eLbSIawajbU
+5J7P2lXs2uOtmpOAV67XJEZ8u4MUkic+IE8FxwWnIy1O/bH1JH/Cp0MWDcreMskLx3+LHvoeDzL
lt32nbrcRtjhsnOFqseEEtbepTCLlsWER4ik7Xob1EeOmjTIx6wRQKQ3FUrY0oZYQdDiXrHGA2LP
s577sK+/st4GlqIpZxTf6dMwbNfzTnXqT4ZVmuAiYuqs72cFhrlJNXux1/LyY4PHDNFKKolvWcMQ
rnIZeAR+djltWhiOqztmD9Nmp/99ylCqH6Ek3BZxrNBcK6KBVctiO+55aC8ET5IuHDg5bQHO8YnT
NB6RUACyMVaBf7botMSa1bQO4Rnm+SllqzIiOCFec1vb/ml7xYVzbmBrzWyJNUPi6nrWU23BFUnu
Chz0bOwymO8JCQTbX75jh8p7UJPsCrFVqSCeiN/lr+lN1jYOEPUuu0T6NmFnzEvHNcOzq2wpY92U
OrbaBLjgUQOQJ3eyDfRMNFYCyVpfuDdZCuRHoArODHHjtZ3zE7f2mPlgsPiGz1P6o9U4Z4KeE9jr
4BkApzAPZXwI62m1me+csj2RaK5s4p4Yrch6Mn5dHf/Im7L+R9DblsqIbo8eKxuPgCeh7YMT2wsp
IEaFpaJNXP6KbNGMkHytOeK2YspjMKevmdWRYZx22YlhdBxa4QkMW0L/jekVh5NJPLeCpU8WDLmy
4vjFC32ovjCw/4xDN+lEikRwKgn/SF7aIhMyonM75x0MNySpII02c3yA4gfq4RLDTLBKmLV/nyWA
6skHy3SW7K1OeYhEMfHC/l768aIgmfCLE/0I4sJ0TCC8sKPvLmeeDK5afP9/TNQjkEUYNztRCAjC
NVs/NHH4TzBbb6E3nozmomjqWbj8eqSFlwADcsExspKNYLyTJ1yVseScriSb5GV2SN1fRCiiVIgV
f+PYy5bAZReNU3ktKR/GVRA7kr+CpKS4XTUVasrcJQtfiGJ5MHOdQKKAtKEgWrNXMy8xuhUDQrUQ
iCRZP0Z7faEMks6mnmMTqOCNVdOTDB8+s62xKyMatO/pTCYjFeB95l7VP4rH2w2/VgvFTSkWm8gx
o6/3e0Avk2ITnlauIJdZBUIHYD2PLuKC2bCYF9JPuLKPgPmHoa4FUvGozlAZDpciXnVAKV4IukZO
mCaN6ThbIWHrs04v0nXI+vnCq3Oarbf9ymTJzWU44J5lMngMV60DjABEKnsJFvqR6WAsr6OWrlbC
RYbBShSsypclV13J6mHCZvquNlGQTlRyn57us8UVCooivVw/mUgLyCn5Js9I1bEe6iZTsGj5CSFZ
qSSs25S62gR3wn2jZoVWm/GKVA57krYHKsL9B82Sefov1SoARMcpC3Tl/GbcfRsPKMnFr0oXwYDy
thpAb4x+hadCgqt/59dqkU552M48Aq94H2wjXCQQovF01LvHbhu5IJ2Bj6+lJ9JX4H6ltNrCtCuU
dp2xAUa1RUrSou7Yhi3KpriOxbhCxlVll/7QeNTM4wqxl1118twlo9iTA+xYxzS64Tsgj5BGSIyV
+Cmw8oPaCYmIOxqKt/YdsQwbi54ebpSC9jeZnFdV25gkqMTVc5/L5s968jbwXnk/yakjpWPyqGR7
jogGZ6QBYIzzAUxRp7zS5scigIvzPYb7Tag/mi56FrlD/bakJ1GJ4BEpPUNxNtzxIu1yh4RrB2Of
qnzcAs9V2v2SSNDNOs6CoCji20ecbFr2/hoCjxa85A/Fsw80KMlIBtojfyujHzPZPtJKBGNpfLu6
TP+5V9Pu4xudKMYCEp4fepOgcxu5ROwGglZcqa90SNHirE5bnnMnUave9b5LMF8lCPtuU3QHZx2X
Chn26umIIIifu+rsBGeCetUkSu29UzyC7JL1DFiX/9OE3Y0GO5dD3G9YzcUFbzP3annTgd1Jqy7i
o5eR+99kf2xBxJZM+3DNtnxS+krioVaLLyemZVJepuWp3jFfwKzaTJhkBqSRt7J0TngFrvsMtBHZ
4A77n7GQwRMQW+xXkI//8GLn1FwQnx/1qcSX8JTjBDlmHYNmpZUs5+Jf7YVYzbd3rcOoexmfNMre
m584Jg6wOA0fcsv0T7Uq89kiE49Kxo3WZ/YJbczKZvsztPP67EGJbTO9u62521l8LcSn5HV5CA+z
2Wu2vm2S2JAVcKP36OL1ayYlmR9kzHZj8As7cZynZFjBZddotLgAb6FlAXaXkKUw8U0q6GEwJ4cA
IDApvfSpLi4NI9/dnrlnlN1wtOFil3d9yk6nD3AmVkLTTBS8LfUb6B0sE+dwthqHp5jLDBPDw/Op
2m6c3QqeEInEQNoN+iVbgsQE4EYybPdAXa8Mboama449SAG9H6cxp2eAuNYHrdm1qBJ7remnzf37
/Q41OCsrtnP9KhOCuaSgfhN4DCweLgrPYDu4MEd0GTWk1if7WNsXCjctnFpwCXgtbc48cW0OwzZc
Ri0wYzGVr5wFDQD5+mv4bmFh4z6D2M587wHQcSfSd4Ti9mOigdQ6+pZ7CVqlokujUWSsKaYyQ4Sk
/6uDNgWQdCvRrYTdXCGCVgnlBTIVJv2LLy8Kzext2YHzHFRKuU7V6u0FrK9koxoJJuOSu+I3WmtL
pSocgYjsoEgLYWU5kji4nBUVEofzXlZkY+dWL+a3XACcuX+iiT3h79v9rVE966b2tSy48LGLWrUN
HGeRk4gf/h0E45HxXqECaVSD3ZBvD8nfSlgMuh/DVSXOa/4PVehVGxgcQgUNPcXsGdN5A4HLxKdP
9DGJrW11gmgfbds3Z9gM839npL3BhEkHE72lWLY2NiUD8zvhOb72gl+og46hMSsY6TloqdDx+TWh
RjirLjy12At1R52/iQR9Ztxzs+UhYN0brHMNgOn+3FlebtpsgIfufgytJTsoKRIB6/CUv7auc7aE
QPbct0NRZiiuoBueIZWfXddUMCWaZNjFNS4UGdvXxXUECES+cO/20dbdTpZ8bMwPScmkEHvTsLoC
4sExbJeg1clqtHBmQ4ePNRuIg1xmKTqQ56kMpXNb4p9EkX03+8bvqtLaQlNVWPPTbPT6zzgtXDN0
dCcc0NCkB1frMw93J+UYZRuzvnmhrzbhCZEwM2NBPc9b7jfYPTZQH8Mm3TqOUbXGiMyiRlpxJ+NL
YgcbzmyEEwPunj+Sc/6ACzuwJM65KTA+Dh37QB3oVS1BW40L9WRLTfyLiUVtIFvaYGCeDncl6QHh
Oqg+XscSTE89Q+rSetUrbOzCZ8Be7S2YaNHxoUIszNi5hYyF52LcT2LDMwAKEY4Nk7zdn86m4AJ8
TQn7y15SX2LvNajeJmN3XFHJAGA22rTajN99ZLyE6XlQhYWqtzuP/WraRxB8FpEhSBgNDboZosvs
4O1tVTaY9zfib0H9dGTx2z1SG4cFVJI2Id0BH5IRkJeWrO+EfBaEfIGcBH7VmQJGMGdhMzyj6mji
N8zhQ0ys4VXMsEY9WFDZ9c+kV1vKcWuMxp/1akH4BtZmVsnzk3wCn8Zc77dq0C/T9ced9SOqdOp3
ogKQ8O4bKKo+sXekYCpqJD4O5IHekh5oUi0DCLsuWYniEBilk26rBeWzF4HiIGijD3v4F/WIt8Gt
Uonlq6xgEzYVHMNs0V0DsPc7Oe7U36+wrn5Z6ykTorER4M/6pwxmV6Xbpv6XJ4dVH+F+8MIZUoqJ
CIHOhAIrL1AD+fWAnGpxuZw/NWLvxWw5jhAIaRJKh+OBtecvzHuHehXEgK5qjzyE8tQJQViArUhF
7MXYG9QGUiKRJlXOxu52tgvbuLwgTcgnZfPjCn4sFR00ri4DCKK2TmbpJ20KIl8bw1d6do3o5UVE
wbVStfqJiZ9jb5JGYR5yhgaium3Z+fNQUZC7rmmugsfb3h7SiQ+wjeGo8izD8Q1fkCwZG03V3Rr5
Qqc9zBEJ10rF24A0YW6hiNpcAllgeTHuZvHguEN+9fI5S914cSZzdFjy9JEuf2xdIXCm739lwYLU
boEGq8Ok9JddrVdlR0BHZdJ57av+w3/QF0sCizVoapp+U+39Lc1T+klinBAHqiUHySFnohi2WUH/
abnUKj+UsNsCArgy5zC6fzZXJvFvMkRlhNy6NjbuaaZ7r86bfhS/+IzRGgH9JODLImDGwM8SbYmW
dFHNYsv+FuobDOu/vdeQcueG87PL4yu4JDQdeGz6R4FnB+rMOY9FqBaZFBFJWqQArBgDk/7UrguF
nFgFFaOhjaDeahn+LRUDTsDyJOPbHVvRvXhT0EMlznrOzg68ytrmQW5G3AKLvwAY0dViNoRqGdpY
NlTLMrrR2KGkidjaM2+qg0yVIee0g/bMpvx0KQ7n/vh6M0hrxDWPWlAMKUV0dxR1z/epg0lQ7kBJ
CImFgkFl/ZEVLNkzS6ya/cy43YWRMeGLRoH5z4s3aaeLQ5vmAUT/PLBlM6LeGNs1YKomn22Bon68
D80Le3vMCh8BdhhQ+DD/bZi7vAxHxLv/hkfoSbCGv9/RPnAMGPwIOYc/OI8awnFeJs0S3ERNsZph
Z4Dy7djekxVxTGKI+Xjqfsrb8ikPNta8Idjc5LQJjnN98Fm2PUmtbWwzDdzLBI/Wx0vo/vzgu55W
kVgDebLqUtAueLsz6IjpdOK9V5Rc450X+K6755aJkTu+2vAcnx1hRyt/DxYCbojVq1nJNeCz2FWr
aJvl2mNNegHnnC59mgrsg1jiabmAiQ3/4YOFVhmIx8Ow4VrL7Ju3LbXWOieMd7NxtC/BfHO0Z4ce
p5KXa8xzE0ilAWwOJmMWT801rmeYP11p30ZxKVtuLFCaBoPsPbFQpwCaqHFXPpoDOhp087kWTts2
x81g/j7hT7ICke/Zf+LmVwEPxoLiwxTkVbJUw1gNn8Jw+rGISBaVxg3av9q7JBdJLD0W0+L7Ibh5
NDoH3QMKRx34OAPzMEOQa0KXksits9t+teAN48JqbT58+H74UVU0cKpc4gTnoqzebcl3AGMb8KmM
rofDeH5DSw8i02QMON+4wFHLXZbvOwVvA5vImpvxQn/4aTPcC3tBk/Rwy1Zn5gXiBQRv6SSCLB5D
NdSMxnICB6TRPBMwuEzuK1lHa27Fn+u7N4AxIw4bvsuSHACENS8kjFniwwx/kgTmcxUGfUPqqD6z
q9vD4wXzK/XgynscJvW4UP8557XtFryeLU2Pti01rn0TXGp7fMzHleWkbA3FMBEk0Mdh1uqbkXvY
gkYkxB3fXUszzjqYCrFsWTbXnrwuexCUb38rgRcJ5cDAiUPxZpl1n5mIlj/WKhdYfyXV/7ggxxma
m94XzIZj7HDf19ILe/GW77KwKgeoH/0rHb4hhO+VZQaCTql/RVGZrqZunr5BgzlfKjjNL4AXlHhI
z2EHN1JamT7hButn39oZmmTi99eAm2lDBJd2Vi1GlM+wvNTjm6B4wDj3XGNZU3jgFDZCsrQGbq/8
MiizW1SOCV8XbOJ4C8V4BSYp0k29LN1EVHXIhvseO+anKrlBCzRM2scD5+/zwesmOlyBV8r0cQu7
0D5vmGmSxDTrob1tOWPyucDnuGRyFIDCmI/hOSLXbHKNz9jBvtswbkMgAf9AnkrMPPOz/7WZUT/s
NnQqYTVidll+6YZ3POMOG3b0VC/MlCCKM6GXo9QIvxwXdXKoWr5viM8F9wpbHC/OBGASDEX8yskf
+zDGa6uZ4DvzykYF6S/L/3YEfwfKQj1xmB79okLEwArLE9sBYeadrmTArx96OnZtjzXOuwZbkk+1
JYa5HoiIac++fWE9rBysRNAM5Xa+MGh2ZGH+ZUX+dRxcqAocpwiNYCwkZGbi1H/cdtiyBzp1UbHG
dAaq03inAXfjyM8i19uSDPtE7xp8ZlREaGsyELKK0FlcRtj0cz7l06vR4mqLHCenbCbMGCYduerB
yMkTCvlsJ980ACTlT+IgidDN+Oy7RhCjfZFSF3nk7t2wKk8C53Su7rCDaoVDrdGaeLcWvqxqUI/Q
Ne88qm1KhJejJc8qZ04JKO9hpBsrzqn4+3SMiiqixUThaZgLQ3X02iuPMRgfy1H2S7H6XhUznHV/
L50Jv15Shix9TX9OUv/u8C5rRp+weAyz5pgTVlvZTjhF6GGwYcCj8VEhBtCScRCuYTbfuPw/hAC5
kmIXHqg/IJi59ewLF6R7n10Ukoq91O40WS6JqHB5Q0/AWSeMOr1TN61itL3dbnqiFxs82EOYRIu5
ChvPBBwx7tp/3ygniSycJCWegRbtZ31vJbkVIdlkI/TTtlvtKvR+EOFkGohgBENuFvNO25D9DlLR
8npFEhz3xj0BUKYtMq3Xamg+HloaQB++8OYriL2yDuxrf9unLhr8/wTRYiScNPW45G1AfNwDEDh5
Lep6vwhzcOXPLPMOGNyllu5Oa2hG6FGGd+FIrzqQ2qkr/MF69fX3NDkW4VxedeSZEjYZX2BHmM1h
uckcYFaOZApqMSqCDsdu184mKCAzoXvdy7ZPng+v9TuTSRuhuExN66MUSwWmVwU7bmX/7DvdQq7y
l7ufl9VyJwmVkkUCRpPPJAwr865e1MGF1Wi2mzu+0Z4hD+O4hoNwq2iW3wdVZqY2c9UyaXaTNqG8
YQPAfo1DCZGPVPXbFsbnGjnLDyBpRxVMJ6+JjZjVP4kZjzyLTDHwKlY5cWriQqMQDstA7RhihNV2
HPiEtKzQF5RS4XVtV9H4O39Z8QLE1yauszdtfwbg1gV5FgQaCrNeUGrmb1RqQs65UY/EVDLOLmq9
pXDXimHDgxRoFne3qP6/tlR92QSPm8S7f017PP6HvsUXbDaXOpkzBc1+RrgS4oTnOeAm45Lps42W
mtbW9j+4qbQJnTNtA+2sGJ9Ql2YXoZLhijBqCVvi3z5WFTGsgQh28M0fAxIC/rRVeBEBRgqho5p7
tutbsqYGXi0ViNAN6IRGU6f1YYX5eEY7rcAJGwp315ZHol/DzvV52z39hiz1q7Ie5pEB4lQ2yV9b
/jODHxJORNTZhFCGdDOsMpOQCxBHlWlxJDi/W+XRkbzVdr6PCzmBoEvpc4kEc7hJfZbz7wuKVjIT
KaJw2MjG5dBYK5LBDEX27oIB6G2bajS/n3uIwldw/IsyVlqkxZfCfo+zCdnY1rYONN8kYrFitrNK
ZKqgxEBy0Ey6XgPhKLFhH/fr933808H2x9b65lVH+IPBe5d0a9Kml3vjBbrjRX7iLHxXEkgt9z/z
UybNd/fUsz86BvAnWeHbPJdaPLNPTOL2JqokzsR0PttrJaE5K2X7CElbyfmFgJE0rjuJ64Kn0nUa
uhPsLQ01diBGIUnuHIySFGsOUvbeOGD8FieSvvdX0nlBKmaUkoP04o8zeezZSVmeLJMMepIF+oQR
+IHQZca+xhFefD3Hji66X2gYRtFeQpLFJw7JgZWNX+ZgnvVPSLetKUq6KlrBQoqG1Eo+YWtmdDeg
k5hsIrYufqCzR63IN+c8Zm9jS0X3IpcBE3JaPV7bRtBks3ZcVmfE7dzPwlHtwh7mVfJFhKpIPNfv
/JaXEC9d1YWgiVbiT4EbsszdZSLm4oS8QJKdeT886yRIyvvs/6fwvLsRiHQBIU+mnpwUG9Ow6t91
R9cTIEvSMnrAMpbIP8Be5kK3DHzVK8jXyZYj5d0pMP+TkoGgQCVth/LXSXz88muy0t8Qc/Uejdbb
K5mtBT9FWpyTyqpPUskRZAHlHTU5LtbmvK9FkhCCPOCd7BCGf94G8VGOZfxYRhTZVEfMB/QkGBu8
73AzLGdVyo7BwzGMvWOc38bpR4CA2saPF3Y6uP0mk3uvHz7L0Z2ZsZe/f6+z3io+tqyeDABsv9f8
MurrDYPsI2WY2eWmdsy02mKkayiPF2yMb+zQ8tFXznc00WCn68jnzNTnF1OmOoImExR6Ogvkp7vw
BxErfpJbbjqFbUwBA+i9KuC/hZVFFACjtzoNDJeTHGfMJoc3B2ZDrzCHX5gJlJMMGlhVZAYePiVX
VJtXFzr+M8/y3Xy6WytmmqhstnvC6SM57aMgxHNcoHwHoQWWWnDJ7FGHjWv/NXPLNsIOlVcZD+FR
3vdYT79jsWJa69RCz2D2Vykm9OxOebH760cmhMyBCS5g3/HeEqG6yfVXWdNaHjMFMzj7aBsuSTDe
suU1D2jzpAGx/sAszErfgIucbHi8yAmwOutLt02JNUF0oWKaYW0zkYQWOY6YnMbT7tS+Mid/AHlD
PxDxDd4Lb2ycaEsp7r78QWYe9Rzo01olZL42sq5wNw8xpwpM3iPKaM/Druzx7Iz4/PKS1ChAPaS4
Jmj4/YVVbJ8ebmqGMO6q9x/shQUoSdgyWmPPlZhXIt/QGTYuIUQau30/lN3fk4PrM4txsEC0qFuz
4tr9m9vXx3809GyqRukpfOeyTvlamotJBcSJquWU3p56jo+SewlsjoL892OII205nx8KcuhqPRnP
z/xK8KvBUfKuTPfnyOZ1wjk251WWfayV6505CPkrF03uZ8ufrGmVoLVkq7R/38YIL2JAahDPgY/b
kyn3VisadOYMpM8OER7T51sGcBCE3X5DgmadSTrbbXqtMmMvsqL+QQpLKRdvnfjeIR0XWsyn9kFW
D4ugRdrJTrfL3KQSuyTOqgg5KCJ+T+mYG4u0JyMXZJweBdw0z77SFwHeH9kjqcBB3euW2aW89bZK
nMJWXm1l5E73lnnsCniizaOPJgonxt4Dub5eZQqRJby6ratMit+Vl5uld29S2EqlizxKUPjfhyIy
70JYCkKj5iQZuJj37AI3JDqFRw03sRRXnfXym93hYkm/EeK57qRt22FHxKHDu0VQtKbWpHQqOzey
EZG+C0zw33F6/X4UVqaP14B59+m0EQ87zwq1xMu+z0E/iDGtToOSiiBmOgj4Jjw4kdcMlmvdRJFC
k3SiU7JNcHf0r+vdtmcELgHMvCWCCHXGqgcD+WA4vNFloj5ZFZg0Ml2I3wq5ZspUGEMwy6WoT67t
iWH4310AL/Wvp3y0iP35YYeIZBQ1ZzpRhUTd0zsfSEd38DqExV3GvlK/8hrhrYUMINdqPmICvaJL
oe/czXQ+fDck7Av6N1/AKcN6nb6m3XlMtlxlqql9O69xRkyg+3UlElBnR4E7RDZf9xRcoHz1s8U9
bBQJl/c9Slm+TYk4bAfXL3+lN2zId4M2DWnwESebKro88SAhv1dR+9NyhVUoESZShpKhvK1rJ9Ov
0nrQBS4Qk1Yed5dCNpDpJplU2yIYiyVxX7oDB9yPiCXHcua3aSb+BaiwtADiv2OduyE325jizTOC
wn61ibgULJ33fRcYiP602xPdIUWQJetd70SrtGeHUgy5mK8l1QZSaw24ex6PBba6mxhZw+gVxwut
niR41pIUPpUQ0SCp6tzM7Udth3SIhIXek98oieqWUgoExzUtfPF4jVoFxUpjOnulD9QU9V8yF4MP
fjAQQijVNTmVczDSwviKIvfKr8+qHJBdAdh8pVXRm+PKeitRKAaYQ2YLNKSrHPZY0aXmWzPoGkZg
7U8rNorVWg/TeyjSIBa/j894wfdIE1NARrwMQude7QcFWR+ztaf9+KC5cU1Dq7tjFPKBZSHHhPch
KjfPrluJHmLeklyHuS3i11c3yDtpFOoZpn6HooTHRbE+znZdidcd5qJ8jiBF7w6AqdUkF9mGb11K
GjyyZMM+a8/C1vFQ7lKVJ3ipOgC4Qw/+cbEpbtmP5BVRxGX2tmlVN5mVu/4E/0Sm71Zc5Ev/oncm
4A4S3u3sz2G+LmqJt2XGgQpYAR9lu2P37n0BYsFqMxLPhWYAgqgfAAv8szyuri5Aqe3ryzBh+/rG
UPI2gZbjpcNFVZV6awbZxK7phk/bAkmwmPUxGlzt3fBX+3QmPEiMObE5vR4cN7DpQCZeCSXOGxst
2pru658A9dxZ8bEfVhndhnBA4ya7Owirogvt9/EgfB3hIDCS8C0OybKGyi7eglPH2UF/ggR5epWm
UEEeVfz2vtRpkMIlS9r9agvuzNidIDI1F58m4DCyKAMe0gx8nw3li9cnIGOhSum3YruLUtWIa5og
gKcsKw8o7JZehkAcNEePiBkB5JuwZCUpVgHXTgAyfqGrw0zoPiWJKil8RrYm0TaONiAQdDF82WYj
FyxadrmIOgE4eX1/+Pz2pZokDLsfI1Wcu00EiBrghdFnG29hy0P27l9Ubb1QDmBOjBgRZQjLxra/
ddg31kwfiNxbnsvc/j1YEY9SgvXip2QgBI9m7zpVXDff+Ih2W+/3hDSZ3f9lYdiNtltlgODWb05W
u1ZMnkKe6iNrxeMizO1CKF+0o6XaLHtkWsfXAcjlKKgNwDjjEe180QClaArI8H+FcRce9GiHUJG7
dPabtfvQCOE8hdYNmxqYB0yL8pCsAjUBZsNzgSWpSzCVwj8exhm5EocP7nR99bvEN+VK0W3tk40p
EZ7rCSU0ybOOwYK8kjunszb2HwYiazicgJHS3tvZyzaxyNwrLI+cBJMR3zRY3m9ykbVi7u/CmwXL
FrQsOO4D2EgLhauiLuxiUODmurBOUCPTvnVq7WdwHQniGo3OUn75rnMG8QzyfCEBGxrlSNmE71g6
4fougtxdLkCWhaWZWFoyTO+8edsW79MQ7b4B7CReuoEWX0PKcTMuAOT0jlQkJe4f9afnLgnrjxx9
AEOM2pXT8c5T3HsVEFAqDNFLWdhp0HhKK7JlL1o9pyYKkhg/90b5hQMuXnBpVWrMWsbL0GiKhHzp
TyxfGyHgptLQtT0CJ3oa9uUv70e7tullPlfIaeXBcMQzEVieiPksvTd9RMVFDF+y9+Q7jOrAAXP3
BZ/abxfUhL70ayu/qDKnLx7J3fEWkSm2keRe8sZSTsZuV+LfjUs1PlJyLS88CmoDJdsZsO2KnucF
BvE4uh2tYC4SoBAboGIARwPA9qmmNj5HKFpdkKKlZxL3etno+Msa1kPE4+mdOG7DtokbTW4WawSC
g6gERdeqaNzgwriuvlY8GWEXxqXJBANn9q50ePwzMzlTPGU4QPIePq+eDyn7faKpTspe5jlL26aE
2kjxe8bKYYiIFbNdQhqiA4sgfxAAkG07pBbLv4JS2/RwfNh5hzZsbsVkkkzAVHfVBVRQw8ZAvvKE
/iDA5ezMS+w/75a597Oms4VI7tp4fq7p/neEgOFOTH1+U8GjiJ3beUH0Oq5yPG/l2T+ZShrAjN9v
N5Q3S9elWpzCxCP0jN2F0p7UBa9n6HozGbosW4lu7aeT4p4KD5OrtJohh5in5smM17wlab9oDr7v
YR5WNxtR2osQdMb+ic+yBGHodB8sp1Ai8LCGSPH/dk/Jk+6QLAg/l8yMeb24S0QNvUVbt3BpIlFA
2x2BdrUQE72oZY9myj6UWgM44ff4zJ6y+oYFZWI3wnw7XOK2f+1tNOTjv2KNzizkUoNbLN5KvmnR
kCDwMOHT1NLjK2tshqU5qN1QlP6OY3O75Gbl49FDc+DobJcGfJfKhN8qYhwbS7NPznXcIfAZjGKa
kiMaKFVIefFaSF2BxWCYKfneDCphTZ0ErHyMlllCpiPbbYqXnn3cyVj1vPKBLSUdImyBVJBhM/3k
wJsj23m2bn9EpyB2vjowsjRGThB0fuF9wnboHTwqotZ6/Bw+Si2ZkzHF1zlRBkDlHP+BdC7khvoB
lnFbC6DrPhPEMKQVKNs4jUYYs4xMIY52cw05Gpd4WoRBTdAbB3l4mrwRQhb3rn7acwlPefc17caL
DG9zK36lL0uxs07wy8/dy8M7oCoYK+NTCEjaCzN3KYS32h7SGoQXsqEX0M9F53pc75VtVPN58CmM
Noahk4XtvZ4gBplDoeYEpiYeavr3FukWyGAt1kVs6p5sRqcCUeuJczmKNOL4Cz0R1S2bPaYXv0sS
J5y1a6Nwd1Bzr9kzWZqfufwKPd1YkOnqhHqv1pWJ45Wr4/5fCcZU+hbB+KcTCzmB5Sxjw0w4qaPw
BQ5Km1dS7xWPJq4RG2gGCaiJjdlzDeEj26wMhnSw+aGIk8f5BRhIuplsTG/e7JtDkrdB0gKLmvkA
DyLq06+/xndR+ZdfJUVQrnKA94pqI5WmU7BwT0SyDxuaQvASlWXr2P7NBnBndziHCNbgjU33K6XL
j4hktatUtMKUUD4mP1ApPrNSnjYLiS7JbNsOc6fyoqTxvtRhwYIqxevlrlPAbj471NBgg8GiJDtM
66Tn8CEWDVes4pAgRRSPoRhBTZhRh4In6E8U6rRe5DP/I+wMNryRnwuLbF4pB5aadorM8gWQZFEI
Nlk+7kOt1k/hcG6SosTPInrxfcJ4AlCcfU6qHI4Dopm5oKy88gEBMSiohm0Nq/6V3FGI7A0Ma6o4
m1PD+E6MikiZc0pyyV4t67qJWkNSqw1ho/WjUX2qx0/YjXH8RPFDjMCyKG39ds/3bjO8GxZ1zOXa
ehSHRVV6IxeVSfoXxoPrYqgQ3QgkM7xkpf7zQ89Q3muEDfPQqnGdQ1rSu5l4lNYwxuAKCvUIB0bx
oMnSOCPEYQziBxEr/5Ehoq4sDmeauVts+kiHu8coC386m8inY5LJTkFHuyg43+YccPENGOrRIoE1
AcP/3oy7PeBcyDifqlAPIZAClIyVnzygo/0qaSDovgmQ0QIhqsDYzAiHGl021dMGcSVmW+Ks7fzW
NROOUvlVmNWTRxZWkA2+yjbN58VBEwH84fUyyN8/s0qiwzdo/35UXuoCmX6gmyGvVSJGISnUInp2
H8l0nf9KH3y9Jy7FHqwq34G0RjJ+BMyoAYoKtC2svFi1N/DvE7fGKEhEJ4eHDCY9yKTDAQIuyjk4
uTnuIK8RODqz7MWPJenBVhmesMrufZNRnUweX6wn2tjRWBa/v301teioKMLyxlxGnYw8r9hdyV0G
RPaGkvRsDzFboCDlK2A91I2lHAMs+psRY8G5cII4l5psU2WFe3dS/aAXA7IAnfnx1tNYDpipjnLM
LqUhy9tJpNf0Z/2Fba9IHWQv93aoFNAGB+twmKq9i3XTiPFoMnxaFV9AGXz6pxC5lhjcHnznriyW
sZ7nzHMv8A8uQQrrilMS6Tq793tXHt9N52wFYbGK8crx8kzJmYuSSHnNWf6tO5MUHmZfHrhDCS12
2tOVUjlUI/Yy8gJpKyBajWcsIF7shWp4jgHtPe+diB0VbZNuWxXZFq8gDXLEog1uoGcpz1eDmuwK
5Xoo8WRHDQf55zAWBFiJyVnvS7fiK9WQKiB9oDPmWE8AH5drGZAArkeYdmqO4PNHzd4fInkSd1ab
yaZcy/+oKvIUaMJUb153WgTAHvDtgzQfbnnlc4m1MCBV5U9WjgjF2ZCSjbeaiVVOAu/yMQEOrVrc
LLMRQMYzDXE+Fopn9kj7wPN1NfqLqJFxsbtUeATI5FChmT4Yq9RVewWZNhdZtzThdRFDnwk9dw71
aSxa6W056cmpMQYYeyWTO4pVZeN6+zOED4hoS8A9AtCtSUnIJmDu/4mv59Ve6fqYmzYQEwuQEw0L
BBts4OG7hd14wAEFAI4QkxUCX0zNVjxPWRk2FvhVK2SMLUQoa3S2Y9SnT0ZnYBuZWziKAJQCM3IH
CPgd4qvPJ8vbfl1yOtxn4Tlsu6SmlH68j+qTlnqVgIhkWIfBmvPZ9snqNOJPi8sihtPDfs6CqiU4
/cOw8MhFkNgOELw3CT7wpufudGNVb/7xdvinwk0sccfOk27KFF7c+Cu3Tn/Oz6V3MmIvmhSidpnZ
mIYw/Xp4zMASIGpcvtVC4jxfrOsNt5vXhebVfQLvz25EVAbTFHrY5R7lc9jpoRRfM8JIqKsT2FJN
SJ4vJJtwe7m3g4BxbtfGPywTAOjmxgpnJKYBzcO+MQDyUn08obsHpsmHj7mep0j05GRmSIC9n20N
DEHSq1Jz/m8tjSagZNK6fhCGd3+FcQlJJsFcB+fFed9rwLf5yTyTDAffHtotfKKWacV8M9261zsa
p4eGgq0N5qptidJn5vcMcUtDpaaJ15vNUP48ntT3t3BZ9z+A1XmscMGCLJBmsx3Ns6wjG6LDNq8Q
ojPBRUc3zBwTJ3k9yZYj0+UtQ0SBhbgxOlWHYzIafaHmn5gR1LgPJtm4NIQhr/6KbrvFePcwJmBR
ZdETEwX8cBzSOIsu14uw4Ot3QhP/NU6KcFjWMD7EqNS1wJUTgkfDXcSd7Z/w+hmCB/sdL9ALbA6T
buViUbhd3RgoU/w3J5+QFko6JAyl3lKeOzMOlFAnKjKf6AKfNdLsH7Ib/PJpWluzg1qlLo53BUdA
EmTFGF8vh17Sa6sk7rlp8aek3tXLf+2zxsiQ3E+iZeCUbS8QdwZP1KLdg5ta9fLLBOGa1aWhoPxD
rUrXW5NEPag2nBgon2vwzS2iPs0IfzXcGe09V/UKd6MVQYMgNTxaDoQopuogYrMsMZsgPqZfAE5D
8AIsjLyGzbUVXirejd9+y4knTBPSq5O3p0ISq2IMvi21oGCW4/fTo38u1JGnUN7Hg96zms3LuuJN
P5ErrIVjYK1jc9GhoymEJqXUbihUSLIi7ejDohUSGN4RUvsOXLJnsUGjFmpk3nPdaO6LP1SqIgAf
R+Ef98VXJNj8sk2U24IVJNzIn4D1HffZd+lwmhlkafQpXbl1hwRwF13GFNFPNDfN3Ltz83ShwMQC
pyKTEt2tDmWU2WGuMlO6xPV7lHfGtQWItcs1BSWI5iMZAKcoi/S5QCaRFHEo2CAxxKBwriAZIzlU
IW+8ePB/iqbTt1CG9bJQ9zlLyPhcO8o4TiO8XC8d95jd5LkCdHLvsxW3e/bzyzxBIZqLQMO0vmAO
oExBb9cljkLzVjo9hFVFIefXs+1VF/WqquRAnK6t1C7GVx1sMSsDljSjTpEiZp1CfHs2sdTpuAZE
f7apyexEmI31x9k3ZH+j86vPRyVpwJ4MitYxgPFeqf3Tm6/3w7vX9N8Eiy7VVtpnhZNkd9tcisYs
/kVOE4ZnqBcaO39SrC68u6hLkdba79X8MOR/heWIj+C1+hp4WcbfsZwSHANt6MAPYMyQYjTDSwbW
MzhOmAY/1D+g33mGmry30u/LSHrMtpfonkqch09ji1r9r36Ioa6i0ozbfSXN/h0WxyJ1IgDkxVWG
4HHe0kSm5dEv6lZfCJmBUzBZ8amnvDOkthKOjjIQW2Fqs/Qlmfyf13+tpd/vnjev4Mp9cai1wag0
uyulAuPRUenVzUugqdkcgDQj4+DfGFho8XbOwogSCJt8Z3R0zMxnklDtqUzd8VnpaGOoz/P+r/0u
sQVkx6C8Nv4BHOHDPqwYNvcwfyPhP+tWoW/CxTkZBRwKLkgL8BMo/OmpDZisAmcUymLnHAg/5Ryw
GvxC8L3WnltdaNvaCGDmH/SzG6zsO7+U6q53W330EgRLc8prOVJy1yVIUEFaE2OTF/Fp6s+/748x
oLKHVDdiA99kdjyTR74fqEydCcFJhfzDfxqDNpudwUSoF3eMSDfOzOOS8UBnRcm27RdUR8kZB/gn
VsI5DSJsa/71oOh6kLS13WAA+6n0S4ju54ZczISkFYGttuYWogtiN25swbHyPS2qRjSBNRrTzJqy
hSlB6cU7VQeUthE4Xb+xNxNS2Fe7FvEmqRKaqbhKvE8B2rGQlosnQ9uEubwbgD4qB8VM6VZ9jeld
H/AD27tVVGSKzJcvj3R+N6nzNXxz8IuDMW3emHrxUVS/aWWpu3bTLoe5VvkeV0TqYNthzkaCU5M+
h4wSGYt09r90YPrVl4AksUbIBjHOG31UazJA1qB5xGOToozRmQKI868j5EbZgH7YqQsRkvHBAavm
gl7dxZQuuVVE4P47y4hYkZApTP16SQfkEEqRjpQ7UEQK1MtHZgZfUA8z4g1aPeaS2kjqCbzt3Z0I
Xl7r97oNtVuvnhfdWaQiGwRtmLPPI18xH8JWWpdVOHQQV5ztYcEKEHbrkksgOEzUl2hEmsyRVun4
/rMsivnB8eeLzucNErnBu+4yPpISkz6WohwjFLlkJAnUuVuFXdvwLaPBFNvQhOsWCUn/6R8+uJy0
idF2LqwWd0niNh0liWzHeHPVQnvmAUUolgEx6Gs3iJ+islyvc6yikB/sE87anFLigH1Wpiev7egj
L0TCirrs/0551jjBM+lT37ZP7sTIBwEH5u1gp3Wg0t6d5k1cduJSHDI/civvfW+Zq157mBD2NdSe
Dbe+GEuD6OYUxPuEAnQuVKYChxY0gwWi1q6iz2jZAy3XqnAonMPdjJRePhCcD2LJopJd5bu2bYyV
21Jj16/TCXVgc8Qac13QKXuJUO+H266Wv0tUV+m1/1tCP7LmGK1K9F8sHIyeqBC/L6bFKSOFA1S/
1EQUEBu/X1qxPJrSvl6F/oEQfYWSGfLCHT/+o6JteE0xaaPRn6pgwmJcJP6PLrcv2YJllsbeQpub
Fdn/VF48fLU2pksIzGmfhxcpslXlD2Feyn7LXVRjnpusPurh5qF20nF5tAtE7OMIadmfc+Z8PHDn
qOzgpPaOmN2VlEpR0ns29UK5MkyK1e5lLNsPpHW11QYVqBoxknyMJ88oPbO1xJt9071xjtkTavqD
00mF0Yhy45zR3znIFIx+meo4TrOsJE4rEMok6FX/VWdox4nD9GDhiseUDnAZt8Cq1Y1z0WCMX83V
MSP81a6TYfBxr7nSmArDscOAObOZvpckvmmrmhL3UOEorPsCbVMbSwIN+uE2LVoqRU7oiQlQUy5Y
QGabxBWQkk4FOQPD6mVGpF1LUgXTNc6aoqeBriWybiNh1uxjgTdHBntm7Ft46DLOg8HSmU9fvjn7
rKDvbYYPr24QjKJ1GtFQoQ1iXtJUZC50w95OOkZLWs+yQsF7AwocQdnvdMU1hdZ0xnEc4zdtEq0S
re9h0GNjmERWgWUsIeCe+eqE5S21jRsamgZg/owO8RZ9iu1X6XHU0qUonW8JjOcAFULr8aRgN5ar
fVGRYIxQPSF36Gn+3mhJXOVeNdPGGBTxCERa5WnMU9Nji55CYHVJLkzPAYFNkBYOSsXnsQEEltIt
v4k6RhJ63mioXCzf781DwUz9r13CIXBv1q4IvMKEEOgTF4liAVBllLRrsPr7RJjZaRI5RWekAYzj
cPgxeo3wbxRiQuRKhFexDNiwsjiKoUToFu8ORI0GZqiSDmrTHCxP7eAUmmkuoy5n8jBZkQ3OiCSI
s/HOroajiWQ/Hz1U2VrtJ7XyD8K6kbI4PGy0J2ANN92zBTke6EL7ZbK8iLSfxSr7j5nw8KFI/d0+
B5VNVwrZtYUVC7ObUmU7rqn8pjhUSyCKtv50Vgr88FBWmFp0kgHUEF258+F0N6vss5SlT8nMF4NO
h1mIgiLRfdcvvWhQAOzQzf7ITDAyl4VsXAUg+GhUiguYqrLUqd0ZZmh1q/ZacKgib+QUcfH7Gdmw
+KhbWTfxIgzzXMurcxyoGvfrn9Xj3mikhZDgpzVWfkPOqvxiE6t7HaRbpljuq/KgdGpMQacrhr+A
fLD5r6m7XkbTMxPKxrVm9aBI06fccNyMkAWxzBYSEa8Fttyi3G3OMT50PKMmgOmxWYCsao87gkI3
kPI8Ob38aFcdW77fDCMbSEV/Sdj46KNIsWJynGEYeI0WT74CwMIxP1waSxbyPD8sAOtj5g5zGJ+C
UI8FTHRqaPRuaLIk0/5NajuXeCRj67ddY5x4ssvLrk7JOkMgYKcnnfKQTovJWRjjdcID1MeYwgwH
ayVjkGBVbZ2G1P0es8e99P7Qxh5s6FbDIv7S+7SGpCe0hzOAs4ghQEm68G1NTQOOZ4HN2TY7DyaF
nF4EFoTLmoQQY6XYby5D+X9mSBkua/+pCaFJYGVYukaefAuJpzBeLMT5EFRIR/CAoXhyZzjcLKoU
lOH16yZYR4PzhLbG+37m/1ioUjxhBTogmL2LxQqFUQgTR1PIC/aLiPAfKB3UP2jo8oUNiOiGYxHt
bw9hGv1ONDDLRtYdk1JLp8rvhX++W0FwhFSOnViQUTysNUpAuUk/GuslKqm3FQLFG6U5gcmULpPk
RrFUGcGey/zKzw/yypxzJt/N6rHwPshsAZBM/QrUa7cAolEyngsXMJSlwxxR0WFqCskvy+zpKiQ+
u4ZqXztSrtRH64po0yA6FV8Euv0kPg5BFmUjg1qIedD77wvi8ujPQ9WP88aBx3zkY47xWBlsvvcQ
cxPj/Z+og7R0TLbKMhPXgAQi47eEjFoZet3MBfjCDQC7FU7BhK4tWAE6NdQKuxDGuSZwdP7AfQRc
4GdzeYTDDOnblMqhKbhFU1jK4IOpnku1zBS5xU0MK+2JMJqjJsxlpSUqBdBTkTOUvLiRdo8IoyRk
zQ8SpwqiKBgivTsV0lxJJTBCX/YysSsIgo5yE6SNkVL/VgRvc4phKeqOl+8bEDDDqrkOFUFzKgRm
9Y1yMZb3WadhVg+NYpHSXYbCsiPdq8Z1tE1dJ/huSkNT45hLEyZY0dKTV6cpzHKC+MuDhVGAh9Bw
Q5ftmyThhsr6o2dwap+9OYne9zLVhGwNYK5vE9mEcnORZLGIonjMYMcomAeCMsvVjit/JPAoMM5V
zjaebHQ5h6SBzVsxhsuSkOveB87DO7+8Yw6p4WGD2+u0E62Kro4WMAE2s+pU6Mkw69HZfhvSe9ok
JwGUotsMYuB4mX9BdV6FAmeHtP6qGkWFEBvSTfak9FMBEQwwHUvtOS+3fhN/cFoMkJN6GNT/fKV5
tJXHubin0a5putIRUDnMLd6L3XV6YqbZaIJs+61KLardbLrsjK+EJQ7W/ZXb7jYN62K7HsmMUED5
ru6AZwx9lIH1aZLT11+HqGsRD6aaFE9EgfyM3SnhMiETTg6PTeGZHHFbLQY410YYvJeLocLhBPeJ
QBhY7d9aWNY40opvE1fBa61LzBASZz7Z5ERHfuEL4zqk9gVCLwE75Q0rFG/Yd4QqtR3wbx1QeBNe
Sa3DXKYXQCNng6uWCAlNh0msZ1kTmJPI49jmf63XX81xo8Bla6IiiLQz/XvjGoVRTm3eJ1tsf/BO
9fZrAj/ojY8tz2hsdUpx0rx/Yr/YOh8dT+tver03tKYsIHIXv8KCl6yru6fP7XoHadsnVwAQh07v
G0eyIcNW1UF1GufWeaGkOD5DAF5FSQIvpqt60iC20pPX8+aIua9J0b4RIfZGfvw6ub6TN/mUGrzb
TDQjFQqatIhqzgBdY5ZjiQAGMj4heeurI25gEDktPNks3I4Esf6cRReKGuPCVUgt9mtlvPHD8QvP
mmi3sswU57/98UFf+LXmasLc9T9poGgcBrd4vLWtMS6TvYZ5pnXRKjk1l0FPgd5cvOdwNoIksHbA
PO0QBF9tQ5UwTvmisI9Oxdqtn5wxbbLK/TFczjb8KJcM/d/0FG4BZ4fqSaeu6cdTnf+JCvov4OrJ
qvR+B0SzXWh6uQc2M00V3wS0/mwl9uP0imLdMVQEad98t22z3Cw8X3PkwbbAiF14UcslmoYe8iHt
rBOkBi7LTIusNQbsJ7O1f8yPJ1/HrS2cdwlOA+plpn2CJ/Qh+hEZBEwVp4xoBGaPzPuOTHkf980I
iO18oRb2qay6Fn/3OvoMHwXi6/jsX8kqmo0uYGHRF1uuMyo5Fn2zxkCqBaycg77w8V1cRcbDpk2v
FNLa3PT3786NGGKXNg+uUbssVFVYM/hOgYrSzpcgnr7vQoamHlvyzZZTO4xjJp2vVgLr+DQiNy7l
11l2FSOkvrljHyfqOfMYj8krIOPtVz8A683Wvt5kOxmWir780wM+pJNy3RibDn22DpazRQIg1QrH
apGFCQ53aAHdB6xKV4skpqX+BdFxtJ7u+3F8HRxc0JvKJUwsIqNFwltj3gNcH4cy0FRnrcnhcvNc
T8n51ZlLM5ZGpG4zASAFnaSQfHsFLMZLkXgJefs+2SJjimjjJN7u7ENYZLEu4TFME6q87P+pnNsI
6e0XjWpMZvy2QcSx2C7nDT9E6dAaNCUzwsNt15XtSrn6SMMlu+pTvEE5VOcHDx0+jBAUwZ8jmtWY
4Qfehk1zLjLeS8mykLb2MBZ7zC+LQqYG0x0RT/PxOQWvEf+BY7G6KJlQwxRSH6PW6C51VDNhBg+3
MZHZuYUvivOuBPBNkkObbUOZba/PaVMnmPSXJM0gk1fJyDroKYVX0HADS56jUOlkpkGwqm3Z3n2G
W/40hwl1X8pWcrRw6YJlOSNjEtiniABFxw3NmCMKgRkOFmKze5SiOjTIlv34z006nrKF0FQ8QWs6
RwePvkbVh+V56VlkPdzcHP9/3mIlgva/jKGb0PJHFYAXuvOlL2II21rU4FvN+6tpCS3clm5sRB03
Xndt0nKTt/YuM/a+C93JZxQK4InsmSWjghVdyjqvQHs28/odaaUdvsaxlewpBxfBnZyPYY8oq525
tOrWLb4XfCH0EM+8iyWbmljFv1q5mg32BWs8iiujUQXb6pLYrOClnRB0z/UN2a7rWixSesAGObLX
Ii/eLEniAUOKr1ddwvq63NGaTyFkt4ZMlu3f0el+6sugWK307A9UeJO56oSjoya/eAwc/JO9rqsq
WTRCJmaih0/vGydi444pL91IUYFqqiqfnbG1fisdAbkKvqOnX/3GXkkUOgFy9JwDNaza7KgpMoQy
pVaXid/WdBG1o8kdJQKpft13mas0N1N+sXh6WHtFPPvFnHnFoG23BYFxhtAjY09UfFHzRNdoCdqn
2Y8qdCH786kBDjV8JS1N0VzBIS4J96eLZ6ruY5wE6rI3qiDFDqSlkTvpL1XYixtxaFt/DD5ZmZKu
BDwGHKgPxTZEWJnByNIMLKKqdLyeTPtBnzpLgX1vfY6Z3msrDVpVN9ls7HvEaSmHydBC6hxjF8zn
+VEf4G6FqYdmy2NpJ/+IBvbYBQw+XeFyp/C3+CEq3Ofgi+M2Oz9gvcKMX/K29aVsh8+Hu6myfUuK
nEzrjEKZrNK+x3RcDNRRxLjmM2D3L4kgkH6R3OmWn+VIm7owj2vytnw2LkeXwD0bvY8CKyTLPzCw
6fWM8/uIUWI+Zq3y8zuXbA5FDOPWK4Lbzxq6QXTxtGL9S11yI6+IJjDpxJPKvFqErIG9zRvMGj0S
NSFpG8eIZBVqB7NFMaiRCabaiIndP8nv5tv52rbTXdUUi0u6RdmwHX+UQs/NhVkdzfbRM+S1RR30
hkJ7IVSww93HpYBBNjTfThzCYwsCpjPR10DvU884bsE4mzHVJNdfgthR0OrFH72u5jw56zToSlMO
TWz39HZJ0BLPf1Bup8OiAx4Y1cr9m+3zxDoMm225dDkZGQ8qc5Rcm9wNJm+mvnemotwSNntk2SWi
qRHd5GsTow3hwx+hpY6rJ15JNFVRNrIBXuhoRaxYLsR/FC0r3UvacRVH/sgWsd4Gk0smKMl9engq
OAJFcrxzS7mUFCDxoxQzxIKBVjWjafn0sbJHshS6vKxdBJPbRJIBv+DiUOn7aQr6qietvRSSNPMJ
3UvxWgD6rDPBvyGzZIvdeB/67u/Pd3vnJagX4rUP3eJG+hgbiuzuSMdXtojcOL/GwCQesiP6uof6
k202KTH2w0JE1+wskfxawcK1zlz48T1b41b4f7Nu8IC1kUHycrkQ05ekgU1NCaFfQcJBewH6Hbpz
9FjM/T1f+FYpuGLAW6xlCfxsQzVzEz8an3Mrpfm7h74T/LL9w2MxVYVOnAD926t6rgmb5twJIvMI
/SgpqNoxBsH8ll1LhtGas1Te/rd+enuuGAP+ECzB7Juw9YsBN6CT3iiytnyZa3uKz1Xdm6WdlhfO
l24tw4dHBVl+AQUYmqDFrDsoLt1MAAmYkoHuElK1YRr2k4mMTufbAbN6Bf38qti6kD/7i3+irGJ1
o4k8u6PLF8SPtzymUpkrSBhSTfr6sct3870sdDUXrKkAPmqcq4bZ9338iTeqF6gIyHjTlSVzWpCX
tBG2leVcOysBHHr4TNa4oRa2cocwcQue5oT5MG+sIzsRCJyPX2FGJKySNNlaW4aOvH2CCYaPSjmK
rYUDHFSv5CaepKGG9MdgcMqBUOVe6SNcGTX6c35aojEJ4bC7GCQb86VOzZ/iwjQ9h+vLrhdUCgZM
Dpw0ikTZyfjmgfwKorIXYsOyKS2EFQhSBAWqhzvl9LYsXrDnY5dcWhYDELQ5ftNT6Oi5NodM1g/Z
7lcPgA9nQxMq9AzUk4BIKiym3RWXA2ar2tSYAXP5ZE7f/7GTas0vHcNNNaHifRqdyMtRzJjDUo8d
p0zHLMBt3hZETnBWkd7ndj7p7dzO74xTkq5C0e03UgrVsikcLGzWBQJ2fr+jp7au+GWqCkTKiEHo
bKBwUtgjvj5cseccDeREy6KQfsZ5VfC43TJVFetgW+tG955C8g3sI5wTgKqZLubmU+fhuzg05W4c
V+8zj/gO6DrvMCZkpzqfgwwGTrVcvabK2GCgTMk62RL/WzvrU4QLSRsXPm9cPzFZUl5Vqig6JgtT
3Vxp1XbqcFvXhmxX/KULXb/6UK2dFUHH9JNA7bXcG1m9u4DQtEzrDy+Prt8G+wzy/AQ2inhAD46f
2j/gzJixjhKE5vZX4KI7yCfXBcCiZufLI8oXLxGMoe96vOLDAK7c/kz0BjfLtZyG9TCOODy6dsNx
h9iLyqok3NTMtubiFrqDSaGTnwWDi24j85asHnLEmq3HdyiKppCa0DCWAzmkXoSp5m7JE+QfAvfR
QgbEVUUA47hP5dEuDQuY8+XnM5hAw2gVCwhpnLb1IMOimA5UZUT16kXI89qROVdnU0PGIkhZGhen
MkiF9NjEzojapSDbIDv9oE5yWPvPn/53xFT6rma1kd0Rne3ihSzNQ+DKSZmFSMDXZKpO7jM7AepS
FNL/B+NyJAE2gP+pCCxbjITV6yAzWdZF2v5wJkrMQGA1I2dWglu1cAw307k2S9GYz9v2jjIR00Lt
qTWSb2lHHG4KSENw1YN08MG9gV75KaQpOYObyy/xKArBrBpa4pQkGxJncBejUG1R+9W529MZJul6
kSR0bIkn2EoIrL3Qfw4q1bDTZDC6snh34AzbYxCyVB3oiKseDLVwzUuiiOt9uu7lBxZzY/R4Bi62
sbFQFHklWeyLpAOV1RDRXb6RHxBN2G+RuOK/BnOs4Mdl9e1lJSdmo4BvJb/BuktRIHB28fPGRmeJ
my7EXMPDBfcdk1Hx+3m5MxmbwFMgzz5RYAUI6Uy6MzwUJPdjDDLCC8fjdIt0bdOiqbYZJ01KwvAd
ZG8VkoOajYjSkbFZK4u1aaA+s+XZVRD0d2VhguYLu2PGUT5CW5tgh2P3k9jyOFdCSumfZlRXigmy
SXf07uOKECBqwku0zwo0OJfGES4sF36QNaFkhy/tKgy4USq9DE6OBFa4bsXWoSZ8627NLP9BplM0
6arM2Ad5qs1MjVdn/1L9WhZCfEJRHOBWnKSikIAWypG6bO5GNeA2W9055qqI7/4lRgdTucjELL5s
2SigPsBDtm+2/Q3l0pIKE9DoQ/Cawwb+9t3Mcoq216w5fl9pPvQrz6rCxZw4s5qY/o5AwnNhWXzf
DjVT6mNAW4KeSXOyVdj6fvGAznvc3gq1xa/R70EL7YqB2A633bvCgMKdEXuz0rRHV6uvDdvCTSr2
hlsJd73D87XtLclfOV1W757TZfgmUcJDMpOoXbc9VIkWnimr5ZVHJHj8by6UBd3qjWVazKhgiJr9
cHRqoXGMEUvLEXnrEVhownhKzRPr0G281xC9rWmis04U7zLI6qWqNWXqyvvinxuO/YxpayMDcbP9
2xZuUBIj+QS9RU0IxOTN5j+dNs3oHo+b1qYhV8PyX1Tqe6+HWic0g/oM8ABCEnCNMjn1Vf7ZchUy
qMDr8y+hMVSjZCPuYeA/ekxqLXufikq3PxtL0bWSAkuZOF4KYSVxJ2/BALnLbKobBsZXJyW3eu1X
jCXfOKFC2nF8Sx2CKxSH1mQPBvgkw1Sjln9hdPCJRpC7GdhKlpQOKVdy7cAPDo4C04EmdiG/wzUj
jjxqu4PsmJ+oKv9B8vxvg1CJiHkJ8ZB+L4HSrXvM4Qk6atTuwIHUtuGEiO2qtYpeLSv46QsDeXqC
bEQ5bblTW1X6PZuJlwtTasIjGOV86ZjlEQJoIWP3FfHWfXn148ht5brKGLYhMbcEaYOupgyH8uKu
SIcAupOu7uqPik14ET7sGN7JdvmrA1Isqx6LmXe4OLxIS3iDRPjdl/F/nwKi3yaxGioeOzoh3YC/
mtaP2JZ4wni+b8KSTHnSeDP/hT04B7VmtLFiSjoVSDXZsBlMzZewprxKw66Qop8SXUPrw5kRNnnj
8WLpQ5nC3FwHEafADx1/7AQf0AIzwoYQ3u4kyDrze15Iwy5t7q5KrDPPlRQcaBayq55Gzptz46T8
2foCawy2EIRgNJYfmXLInNwRbXs5XNcRBXQG0J99+gs2efr2s+ZsZval8kUzUQka49Ka9KA6HDGP
sJPK/fkJYFcIdZtnx6fBy9nH4CKjPzUvLP4f+QDRLDY+ipxQ3CMIk6DhpppiNW98Fbd+L9st48ER
636FqPqIpVXWWhKU4icUn/3P0cqYOtcnHOOY/TEcWbPo86TMuWm+Vi/VmOy1WieP3yPf9Jcyr5hh
YpqZ1cI6UXTJpnk1Js5Zw7SFoY1IDGpW2sq8IzrRIBw/RfOJeeTB6lvxIlqAJXlix/USFuaSYMSZ
s1zo4vJSwAopZr0Xf+suxwDaO46zYP7AWP9HiNp3ViR+hSdkcEAKETK0zR+tq39GNGR9duC1rLSI
dD2TV53UH4hFs053BAHFI5ARZ81/Nwt8PO1YNKjzyY2UVnBNxLO4FRln0sBPYP5XIJYyRLmf5/bo
l7u7n8plXohik9Coq33E8TawO/sSMV0k+Wf6HiCpK3ZFoJI5IoZmBQyxv5psJI5zTIAlnMyusVR0
GxKLwZzPVIWlemo649+M2Q2GK1DWgb1JocuRSml5U3lhHgN5mZqwmkt/dWJ0b32srKZFztPE3iVa
j7IojPd4rVz+urGnRev5uHIbcN7cogf39tGxO+ExuuV81gTLMsiJ2RzQYiCzi8O4WA2G9j7Ttn/u
bxqPHCRnGF0QPVH3W7i3Z6wMuxazbWozUZT58FS9dXVFUu3zxrl26O9nWvkqBShO6+PsVut5oigb
LPJf01ZnDOWiWyreQb6G+cAq4xNV+6VWqMZ2OKSeGb++UvnLtMq8IxVikbZaPpSupSBZeVVy42Qq
C3PwQOn7EtTE+1ETnCj23EVZqioDe6j2lYTO+sI3MuL1XB6ZbMEcvt1qRmYSLA6XMlvJxpKnhJ7m
7I4owEwB9po3QduvQo0IN0kbkxYTglTy/qDqgW5Eh2a6yoXJ595gxt0vvFoybTer/dUJOXlyi2ZJ
bmTIGa/mljkkCPgwZZB4rNMqTL9JcHQnBJ+IrVJffZK7OY96B64jJaLZar+RdwYeM/Hk7ZF2X3Hc
Ui04hkxeBv4eyTSAf1lpUsLYK9UgetgWpcDe3hdQT7hRoqFI617N8JM4Ptsyim3mnJC1v03+v62y
Gwf+yrT/60cAgnFswgBdiWbMGgIkzBzTm7ixXTBZdEBS0+4l6iRPNjcQ+0lX4rldwXqxgYJriS4T
I2+/StW3L7kMvdpBMBI2S70swiXySlDUW2YYfvI4LtxRCIoVsJw4CC9sTp0ioH8G1iMJxy/B7zvg
BhvlXgxLlziIXvE163A3jep+rbcPondERyDx+mUKxiMnLCqM0l1i7pK1u1VmUkBpMxTTK1LAfG8R
rjhrqHn5+oq0+bgAKl7cFqTQU2JvbB9oqi5pQi1wOmhA1lBqzH2BXzeHANHH/dI6XTMfNrWbP6ve
cCtroFNgloYbyLO2BOfnp9+w6NX8UJrFjNtZm83Y2Xc4Mk861GLkDRE/jHxgrOfkUzRE3SL8l0jZ
ihP/Jrp9WKDKQEi3sGOLfrO34o5aGDrwdCvvBVJHBFmKzBO09K/ZUMbnqNSkK7FpnveW5HoKcxUg
xGFNehGrl1fnccTmBMZ5U+xT87QixjzrqvgRysPv7m0I8l839o6JFCoz4x+iRIK5PRGoAMtNmWDN
274vAFI2g0+RzbR2xT9mtqIym9tr0/4U3jDPMdS2APDsNW5MmHKEZrbsfqaDFXiivwzPbkZTIXNN
LTWdcSJc4Ti5ZWQ0nrKZ3KiuROpvlAvqWqDbd3dhfRZ9UZnrLQLwgz9lsB2jlvNY2o+AH7mSacNT
Nx/IlDVcuE9WK0WTIieSNMYNfG5VY9jl/A52yIv7BrAylSJrRJO/b4GZO2mQ8iLw8a/+oIbywbcX
MQKnm87mllrqcbE2xaoN8sTDTPUdorm+e9I/5Sjb4Tpjf5NER0AtjJP8vPh8FR8uWGl9NUlQb9+B
2F5r+pyEgt52AnYvYxUdqInl8TkyEvAhnz6XGG7CnNs9ZcwLCxk+meLRwHhvYJk8fv1Hz3/xaeza
T0EYVhnAYolBpnEBXiA5hukNM7u6LqLpxOjfxacLS35VnfvjpjfjnKwzhSUrB6BtJYpYT7KVYKSd
sMRNlOsMw+9VMAhBtEgIHNR4oDjIQ56uw0ashzeuf1SxTVAtrVPMkTe6gwwVO0J0sTne91I6KIo7
7SKyVB731CIcjNjwBCOcSm0eNlsMR4vi40/kLWK9phIHVxjOtN4lH2K8rFP+qVLliqRmxbD2nQBw
Y1dLirP0tk/BaoJkMez2oIgcSozSFQyeu/83pmC3Fn67GNMxkiOjF4uIA7yxOU0vu1va+RH4vu4x
sxHaj9VTFxnsjHSLFPoT19tDg3aCJnkUbZmBSteyyv1kXMu9jgMibUBODwyPXVn3ZXW5UrpRziZ1
Gkh4sC4zjFC6EKiWJ9ERa5iXauh29vb1aRcChTMyXtJ2cR2wTMCZ3X6kGDjUUXuk4Dj5K+hWJwbq
kTx9IJg2/ygJpJZDFVnXLu0tDy9xB9qL8gvYm8RDfiDwZF9sNT0SmzGBZio1eeoUVN4lQMe2R0Fh
otoJ17nqSUAHGmWBZ5MEcjwiSSu22ZsS1AYj+/XZbNto1GUZ2nHWOi9u2gJW//ipzaW+xGyM5CLY
TkBQ0Bf6hy1qC5B0FwVndR17mRcvWH2tNyjMhpwfSNksQ1DrWdT0UmbDyocYH9zQn47w3QRyoznN
USP5N1vm1B0YRWSL/necEnwmzu1xa+Zn9oKvfvjRwv1goGSb7VtSuvWOFr8XSezYdtrpLK0O02sA
4y/AteAJGYg33hro+/8SNW9yTq8BSyhpR8QGx9D/NFn3OERXY9aZeMbJeBbvLs8I4gRbGDz1ZWsI
eBIDDrLFj24cVl5Qfk8TL4kAPtr9mrmbcPfpem64IZt6DU38VpXZFReD4aVikaKAHPWAR8SUu8P9
NoNM5M2CnF0oVGM+wBhsdiopCMjuGV/OUvHskjmQDuIocgrBUWTIYs2+ek9+/BIGrzjjz2TYpxJB
TgRJHC/Y0Tr2LM8DVRcQ0+49ebxcMQ3D7KOIuokFBuxNnnDSu+nvwjS6Hj9ktRboUvFZeXPIWLTF
+4czmGWOvznHHYMNXyFsX+nmWlDnbnRJXhVoOU9GVXMMp6rqfQwNjpWUDonFy6rD2aoYlKcn4WQ2
e+E6zPI1jJNiHX1ThMoof1r63USemylQWCq07rlK6CDvto12fd/6o6OjRJXNkHqzQjVxu8KlAnQD
dMMuqQ3WX1KchwdYCj6rlcKKGY9HVBjkW/ceoMg0G7TTHqgOi7Xxyx3MXQvbRDATzTzRmyGa9KH8
8aVaAc4rNQE6uUBSNF2RrXG2OzxzixOep7ZDXeiwSEj6C0IGnqIrw/ncBrFBTqlIZgcEUPk+aar5
6ctZ0DuVm8Rr7/xIbbIFJPj5v2zqwQgUX8D2n0G/BgoteNm0w/0qeXp20lglFDoyGg9Z4YQ9Wxt1
4UHVsllblwfps+ppAvWoZyV7s8JXzypXrtB/wDL5xZXxuRzmlz3XaxC7Zki2DAd++yYgXOqMW5dc
WxYLDGD2JnEwzxCT5qjKdi7PEbw17Rai9Ra+B2dDVr8nG3LPLA4Buno3nb1eHkWb/TiZ9Vkpf2KI
POOFeJ/MjWcieI5lID27PFvxG9MWCU6/w8QKDehmul3sgc3o1xTabqD3X0N42uFS3eYE5/6uMS80
qkxa0QRlXARNTj1XnmKRycmT2KIzcuHDngTQmi79kiEbsP4mQ4O+mt4XC/OiiFJwnN06Ljt9NWyd
bNnHhftjyVsTsDK8fE13PPA2GjhQ1ARa92FyoAwqAsOaRT0nMYpgUGT5SJ5uh039Q2rEv+Ng1L/h
U2vtCMBeCDpLd0HhhcvF35knZ8FxWduldRIGgD80KZ+DOZrkfHvwynNB+Jne0e6ED8wIomBHAdqv
pcRofDo5JUXM0MXbZan6pbfiCoG87ojKyBtgmI9PgDoJ33zjUt8dZHWM25b7tA7W973ZLqmVPbhz
fcbwedS2m0rSyC2QArpNGqZDvHL9Gxdm2Alc91GElz8bbTvSdMnA/PRiLMBWWqytB+oQvz/EPSy9
/dTrfJa/tQUzl10mqXr3gIUFeF/cfwVti13VH2h0p6BrTWWFTpcq+iLtuKtdZVr3dks7822GwjgI
/xOQ81NL4sK9iHGpuikyN6jV6NZYXdFRrRJXnYaBjse+8fL0Bd0b2XAHHA1VYzkgQbmqumKeaLUr
xKpd/navVTLVqlc+pFjoXnAgrqAmAFY9nxFkzw2J76VFvS5+xTeGjmO7WLnOGC9B9OeBy/ijDDFC
nVaLGVNAU23Oahy7O5iYuZOTSyUqYKFIdJyQ5zASItDcz6zX3WsMbqMH1DWLVzRyQli1qkvPh01b
g77SmnQCgAKfp/6TRjf4XoTGF7TwFikAFnjsycbf9su7JYeSPi2r90bl6DdiuMUyi3buQlFOlD5L
8uKxA1n5bOgiBDoKzVqCDraT+SAhmMWUBbaeX++r6uTu5nd6ONHewud+IC8N7ABEN6zFJtp0E69z
8ywnmrIcfq975T3XRAPG7p5dul30stlD3OApuzRN9BPfVPsLmX2aFCJIQ7bDARVtwB4UAyqmXcH9
yhKIotWAtJkMxHorqdGqz/15o0s/ihwewp1UjU4RLrXXWRS8akJa9iqUKn+XyFPOdqDEAdSkh+ve
wO+TpIhSAORfbk+34CtJVMbN42ooAe9Ja7wOg8CgITyVrI+OSZPeZsANMVZCkxNE0VKO5cpZ1bS2
i0ALOPr9S4QgcCa93htCXc5oHlbrK10eWFW3WxcCKZ0BTON3iY66Xf9GdV0JptOAF0+qRuo6tSpK
BQb/GSgi08vOuqu1F3C7FZ+2eX0m9V6a9c/d7dxOJMqN2ThWwCbCu/kew1ZUSBNI7JWACfqjdIKk
S96X5qQp5liKLV8uygA1XHb+injJTEUfDB5CnUoVdT0Dc4xOaBGsueZDj+HYdhEsUBhOMkDoZM4p
put2ZR3LI10SdmE3Cfjhw5yVcg0L56LFylOQkHToWviJbgH8+whLvxR3m63aNS58wokqjFcpNrvN
4PHjpKeK2CmxfiMIiMF97VHDniKImEhuBjKJWRhW+Cx8KrfLYQ0dRJbqcYFQCPRs51MQ3e4HrRNs
junjFvhQKNXHrKJu6x4+lsXIr3ZOoaXDIy4NBLFsKBupPGVR2tLPtv95WyE85n2FQAHwEqm/TC/E
IdbX/PPIStAgpafGcBwnOEMSH94wTDI6UQ0t06Prdj3FIBz57qwuJfmIuiMW+QLT4SLYdzv4FntO
Hc8OI7p9L/uhGqpaa3Mgtro1qZ+9b3G0TZReDw3j0pzCxhczkjKbsGIuSrwATDF5vfK6lb4eHRIT
ydDXKJG8E5c/8bOqRnQcGpcJis2patyXmIMaEAmYm/7FTz/OViI3DwwegnMHKFaYhl3qraezJjMh
OzSv3NqJnXK3pxavvKx2Dm/+sIcoGTqwmZPArXm/+CeRKEsVMZTmHaU91Zov5Kk+6FWvMa9bW/iP
VkF0tN2ouwN7KLaqlvb7Xt/l63lhBbbdP+00Fe6KgtF4h16kvFnH6v6gB5xc825Flr+HAXn/ducR
PFKJR1faBWLCGx+kXA8eLkFq4aH5ccPKyVKXEQG4lhrPPfsgKvXBDOO7uEiPCOtmbP2HpIuhg8vD
zvBfrxaIe8VvEzLoqmWn5JOzDQmThFc0nKMGMcUR2TUr1OVtder9FO8iHkzNtPNlQEPmEH3CECxV
VBU7/Bha5Iv6Q5SjLaQDnVC6WNIvMpT9zTTR4FBCep3V8dA4CCizrbkqNS22EuU/KPo0a12NFiEZ
wXr7wLi1JnVupCpuSGXqG3RkJ8GB/7ypEJqQPSnefYOFY++3KK8Y+zgzKkLgG/dgwj2S5elptTs0
pbQmTKcD4BpkB/rr+K1Xo/M5NAhIIYHUoemduJW2Xg3t7x5BuHtjG75pPAmJJiez79i0BX5EbG6o
UC0iaAa17R1/qRTsHmNXJPWfcoF/8x66B9EX+bncFDM7V1wDoGYSgRIP+FvhBebtIIuwSprHIgop
D3MLpWeasAgAvcrethCCJUqLNJ6oEU5VNCFPIQBbsIBKKoZHsUPnecCv6ViM2exC/ss52E7sMpl3
usjLzRTE7xGhuK9GcMofeX7kDJC2aTX3EXe/OpOEIZs3QSIgBMJMnGdV5OVKn+whiRZwi4wIdzka
cbpbZnkfM1AeWroonNHS7z0ygVqyXx6xeY9q2dJrTMq3agdEesF9zZRWkULoXigd5MFUlZlB3Mg3
EovTiKQG3GnR2pdvNuLgRDZxcnk0F/D6at6b43fl/Yp/FWGKM15i1lnD95iKRnsaF0VyrIstVKF1
eB8D2shoMYh2U8yndXsxJfOKoUq4Ma49mI3xuuLY0aoTex0FWBz8+m0CIO3lRQdNTN4R9asPfYJ5
HsrD/h2AaOpp5LoHNS6orCCPUbSFBzRR3V14YgmzNbywhaihUaZby8t+YB7ztlazMHMsO93hnJvR
KgWirnBifaAyrhHPAZ3Vpqk0qLpnE0WKHExOcV9hGOkAXFRfpAYOWOFgk3MYFYTiLdUUAATeb7Ph
Cm0c+4Cm5krQwzqBaeiAxazKUgD1maWoOYdu+0iW6yJ0YcQ1ltEMSYI+Mbh5iUBrFIvbLHw4W2Zg
AyCFJS4x6xHlcZvxICk9Iysb9McPwjtoCC3CmpJhabFBjFkrAklmGFlcrvg2uWiuQGYKcU1V1FjP
6VFvbQXmatbVVWfhZdIdaEwAjslR+6nQsby6frystH+zaZ0g9m9GAT/6JZN0Ax83o7V+e0ttZzta
184umUTnNaYviQjAX9Z8ewJLHLaar4nXDteNk8mijdCEvdHolBkW/j1r4p8Q+kAv12wMsr2PZJUC
NJTQ75rKcOlOBpFfZmO48RsM66JFkHohuN7qDzgxth6WkJqxs1zUS36bzS11XaCOtS1r25f8KUrE
inpulryADBPLU1UAMReNHWaqHtqryGwoOacmzOhHBT56/egHpVz2XJQ7cbtvG/1RkdmMn6CONjeq
/cwRKLa+05nPGXlpkaCa2YFEJgyJOtx2PgqPuDRGmvtqz5qYD3DRtVpTt4Djavki4ma4H0gaKHQf
pYOoezYws9CQ1xzvqpQ1Bhqtz++e0aNYc/S7fQWQBJ4j7jPBfok4OUqIk+yqM4J0yVX9Tt2waUhP
oUn+SS1/aD7SVKp8XQ/40YbCFpcPSid4nDaKf8vR9c5QFRp5rGD1rCsX/EJA2YatDzPNuuDMO35Z
hj9vlN9YVSZoWQqOBVPyexwV7616M0zxKRlA3vZcDJsrliLYMPj5LRsNk/DisjANScoQ/9Lr/D3x
vhKJ/nGIdqP9T8hmwVJxaKX0jKIMLH6Tl3k59CPaQdAmq8cT9T12fhkLEIa/JFq3uMU3F7wqW+DE
jMolYff/CLkRe8iFefuQvgvbfTN7KYCbGjAuc9GKLvyv9k/LpgkOlezOWCNKhRJLkQnWwGt1j9Ye
5ytPCwzE20jayWBs+6D1tOPESIc8sFM+P3dfleKeI608eQ/sQLbV+I5I7ukRX4A9YILNMSZpc0C6
+4z3Vl/g1s0X0qVWPtnpp6PshLv19re+WsMOqnCstjURGa3dj10CXCjbX8VGan2fTbEWmfbuu4sl
x7CGIu/Bcbw29XN4WRy4W76Mh1U5NsLYOB9g4g5tcpGaffzEUfiVm1zBX1cOzqjfRBC7BvUK9OJm
g/7xCVEj6aJ2aKlBnWRGQVFtAi9haCv01zmPgQ1BRM1nSMPqcojkpHc270iZhwfHnCQt31iRoq2d
0sq5U+pR2Gkrymg/oUHZ87k7qyvzY4Rret3WuX5qAJj42xVvG4cVuapMckCAKGaF2sTUv1z92qrR
oYxBkzaNUSNz2CI37kOypBq3RscovsZvJFRLSLjFaVwTdEWUhFwHiJ4DXAVaSiv7RESBoq0QVXLX
uEZFxEa3dQuxfqFCamgPl56HvorGQ2jpHcCJNkRZ/ZyFBEKXRO2ppz0Gtv22lbn6yOWdXQsckALZ
ShB6v9TI4EBOwHnSuT/f/p30/Sh/aOMJ9I36EvlKCVZPjUcbIcHmEV1bOgFkwKEwF39Zdhk8oljc
+cL9kKq2x7NyZORG46sRQm0vhmNUDL5S/1wur6tIoXjQ9H8JLY0/jJJb++us3c0dQphW1LPkxzif
jZyPloVIH+8DcJEZffF5nUegwgCFlXnGMDLoTWrZn0P9TM4POUqqgeJNRxxxtwrqzxkLtra99Rk+
StbNYe+V/0pg+Y1OKDhKFHVytEPw6yKZI0c9mSCs8TBrtFiZrlAu3W0wSal/taLJuEskcsj465xJ
FZ9Bklfc3yfp+DvuB9Qebr6biR/38ZXKjCL6WfPDwrOYm4SlkVKIUKTBv0AvkJLkq/YPEKuKm9lt
JPIShWQrSvZSOiFnKGvJFSP3i4AFJ1v/E6DfbevD4tSnhI5BC0a388mXjvn9vGse7dgqhhIrymxx
ViGvcf1BQuL1GwjCq7WiqTG0gArNax5e/RmgNOPLWl+mxiDmIggeg0AV+52O/E6jF75Ic2M5E52W
9o00NWkCbDZkv2Rie+KSuIXEBh82yx/JQFWuVJG/7LJoLOZc5zswMo+C9cvkGpQieaCgDS4HREyU
5F0pPsgfAXYxPjxc3Q/LllzqFgW39xGjIUjvn1AaRKoa63dv5AF1L4QH+54aJmu+gGGgI8J5Pzfv
loHcGAmHopPW4PB9Ff8cZaCaofAEfd11HfYSS9ZcLt2sWpLZXb85hOeR/5F9zrBK5faxbmk2DmF/
HkcOIvKNWYuPcA3kiqlyqeyR/pCNpggMBMMOA1HZHGD9r13G1X/oOLqvjK3P0lGvlzuUDLAVxm/m
0vlwktU1jscsLIv9ok/pMhF+Yg5d+c0HFAeWgw7xxKriWxSrvzT+lWqyFe1G4SJ8tXqa20Y2bVl1
0cJmTg6+dVXkSXWYqhMuvsnZZxKDJQcHetBilYmaUxi2OqcFChdi0Ay/lSdn+VlczGBIehe/xJut
JuVolyEHX7xRhaCuSaMwAgNECYmNtZX13Hj7B778+InRGTPaAeS58vYdJKNbcRchlZtOl5HA/tmc
Xi6ar5AD23vFbAykvnfLbDdmoZ2FgmncX6eprpA94AwxmwZzuFF/gbIq8CTN/pvc6MotYh+7YgPH
TjuijqszizHokNrSoD04waNmHzWHNZ+1+GWbRpJUXcab1nilCEq761lYpDm7iUTbflk8uLJDaoO4
ZnbFfEHXglC73Si7RrTmX4I/+D4uV9jKgrGB7R7gG8Wk2zSDD8z7ma3BAGOSEn2Ameel8Jpf4lh8
MZafxskMpNT4QBzFMThBQzAnz46SEFLohDX86Q3KGRX0u1aEj0olEWI6vosmk+rr3w5ebd7s41/y
NmeupqdzwtXtDUwKW56eYPegTjy5NeRGGzseCNRWvsO8KnsfhWOhyMCqHj6C/a8xQ/RdVUpihTWu
PA/wRCpBblfnWc9RiAdECNN6cGqmSQbXfmEXsYXKOgf1CrI9AEabe1zN3faw+dI/TxSmT0bX69dK
0FwuwNUTTSsRibuZF3T+GJxuRtgaGt/AcFf7RTdJj3rsgDFPBE4ithx0OOQk1cTIeVutuyZl5bA0
bfeszC3JHMK+tfWniD0XO6woUHH8wkCMeNpmPxY9O5zbQEbxYmci3xLwk7WajYXRl8lvMpKOm/77
GjTfsAPY/JkPTEDVPJr99oVBj0wBlLvDSiVyyaEoNxQG2OsKQY+CCPg5rJdJNEdmO8qZFhzb7CcJ
6VRj5GaJNYUSRwKyEL3ekFiQaCo/ZWZq/Fpc6ibmbKEs6uPhOnwL677F/jPT+vl/gMraQRBYEOQs
UnzPm6tu6v9HQ7cCc210Rf2UMjSD6i7yciqrAgbGX5b3wJhx/FZ2mKJH4Rs4ZQXGB/GfMZVw/oNE
8Wf9Kaojm3bnWSkQB3OXvU4ox/z/5ca0q7elqP+l502IcZWkAccKT6yIETmOjbsYbQuECdlk9EyF
78l2CB94X8KSDCkixTsUP6BxaBB6F85JY+8TAl2XdCb9DG/bd7NpK1lmSLfE9jE65RkSDycX0o6/
EVw3fuCJQuI1QlUaNWGps+nD76IhXrHi3cH2XDrLQHctuvIJraBtJQ5l934NhXlEqqXinmLraJ2I
ON1/vu51wFlKK2tPkdzlFsllWEZU6V56f7xSkjrEEYgXKDnHpFOjUVo7SZetNNcZnO7b17R/I1tG
bleVZSwfXUJwsOUpfHyhFvJyHpUqINoJ4mvwsoBCm3Wvvv0XKsRCVNgN/PguliYIQf05OvXwQ2SZ
eEC7TeAUFKeCSVr9I5/tKUFPwKbfHIwiO25KwvneAhu/HnNmwe/H7yzQOYPOAg4y6vNmCyVbnpHT
DJ7X/k8UFKKWUTW89VBlsu++41XySPoag4dyt7ghRWRlZUtWU+yrBh0zy00WiaNrkb6+XQScCscO
NGLPZrH3/PVWpRSSwFAZipFloOfLbbW7JzOn11xamF+vzFoyK9eBEYewDWh/L4JqQ7/cidkm0fel
F6EvRnafVRplE5i29lrYvyCrDhpaQdXfxeKffWC1ORQIl9YHcO5qMMryOfljTYNqBAfI4ACfbsFO
diCDRUfG3KlyKvm7S3C6iBM3RpOGWKcEIf1vKMfA1pjPxV9Key5nsLxKcluKMVN/SFRbWMXy02o3
PuAiWGN9ujtC4/w7LTShK6p2wQhWW//6Mn+52sRzBwVAhqyZAxONzQLdU3V359sKabkTEWdrRVHv
9NhYa0x5Qvo3Q1A6sMPyQCNtuaqJpKul9i7Wg4jhz1fe1iIt4Tk6Gp/mF6CaGCoNzokiK3mLHfyQ
L0dIA7WvFjyA7s+cMQbBIHbq4EsMTqQR8dp80QwH2xpFllOMfT+m1cMzeUQoswX1ATZR6kzikgSD
deJeMAgcI87qihGtVx9k9swgaoKjhsRaNhGxSojPI+INrCwbrxsb2y7y1ifPocILuKuIe/Qm+Q2T
wDZbXYFRD22Vy32Sa0Z2EHF4BtZv+tUMHfelHXs5ZMzYgIohMr3epgijWLcL7XhbnuGPSsgM5HZL
AkhtulYJaCTQMh9PJlYfvOGxRMM/Ika21dx/lxU1PvPyPqzbs5pgTzri/J8CoZbwkUxXGTGAtSvu
hWuPYFh4WiP+fnRusipbsYLa58KvYICpagPozCmgP++g8tPgmy6ruoMXylcchhNSDgiPamJ2nPCN
3tg+UbMu0wPyiru6zMaPFxYOiX+ijGFIdzHRpIQjavSTZQtagy0ijQ+0ZS7OmDjBUW/cokb+HIrn
rKgC2mwlwY0++CsUh1O5p3b8Sub3XRehVVlLXdCevZ739q4GX4k6gkbtXmeyra+pTOkcMGvkFeIi
ZzNIJA6KUTbPpDUPvjzbZ8+69DYpjUrqERatcnUFBchz8N1mctQTXt4sHwoJ+8d7R0wbGZXg715M
W0jt6eLt/IgIhBal+S9tG4Xj9Awt4piFSSq8I2YXhY2TCfOCpyz5JSWfbUa4M1ZSs2yv79PmMJyP
Q2ACiZGzQtxCXvd/N4oL41NPiCHJy0BBwfkbmpWAyemD/kZtkUo/r4rQaznCeGEX/WC10MBiIoff
KG0hk+FB/iM3mlVjbE825tCdiutUO/z70ffGxFX/EwmW6kUQeSPMnWvrrRltlwrdW6qwqFw+50N9
T/pzKiBmpAx87QDt0C+cMfDe1L6TA45fCWHc4n2H+4TEoKVHUv2RRCpUJ+PAtw/xkZEZHNiW+f7v
aYluXrIGRfX7Ue1IV2PIh1mnpzE7orZfESydOhP/lTJJp3ukVXJAwWj1mRaCI0HyXVJPpovghKZM
iYKoTWZzxCTn1IYSxEyeGI3Y0vD2e5SmrVLThHzz/xhXuq1ClmfM2nHezjapRoQ4AurkytPQ3tJT
DT87Euaa0kvzolibTBZt2badIAchOcaI3oDbWpfCVioZzLd5f5J2/wH5dVf8uyC8UCBTL7Fy5pf7
BrmKzcmdz+cUcyRCoU8uXCwRbSgzfdccClaeZF5bQj3NpJ42AObu7KtZJpsah7duZQJqfYXnD5jk
NdCviZ7nr6gTMcUsrXP0DA59bTLT1zNVetxCsriG//x0L3VjJ86S+tV+fjw1SIfuAKxejaNcya7y
IZxjzFNfs1o3SZPCzsLZ6S7KU2JEhUuBivOp36LSWEsJ50sDZvsThB3uP1Sn/l5VSb5VRY3Jmhsz
XYnt15RdX4lgNcSWTOY3T7c8g67kApZukFA0kD9SuejvtqP+tdxfJLzsizbVqm+D8DbexRQju6tW
WiCDAIKU09TB+59tsuTDeE3avAF/v1lpXEOu7LyGBlIFZAXrSvsQUtKnP6cqKEcd0y7wtRqAqDW1
rSGrblDIIwk32sIGkCGAM66dp1v9WTNI9OrgAutKinkMIWkDXqx8y4a/81pGbuuhdCtVTJroXdhH
O7+oERgR9iM0YiNnD6NrLy3qlTyp2bOcDyO/C+96vH3nppM43SLecWjsdI0Ch6gaFi9o3N69tAQq
pHQe313OADWafrOj/HsK/HHyMJg4fmvba65MXh8KNRrgtyeziKm9hK/G3kcsR9oq6ugmmpjjeGYK
FRdjQ/yULDjGbx4YQlNGnyLW7gGSZ0BwaPMMl/yj87RwscJj4M/bI1jQFFY4axGIN5XUxgM/4K05
QShDYtx736TdMR7lVdK0sSfMdT0I6H/H7WQ2yFfAu2bZZuzKcC681p67FvRF4pxtx5mlJHiT/okP
xRJWnLw5+7oWvNRVjmFvrxwb9hctE7clScp17jj9y+ITdAgXKyzVCdqg4gs5si3KkQFqQ33rzBKh
Vm2YFvuJ7O0zwKeasmgNNifDRCdbzonwuD3sbzi/e3QQmp/mtNgNOHm4KDJcGLacIvdgRGfUKIld
1vJgu/s9bJaYBvJKufRCSG38BBB4w+6dUak7vsvxqbScu9Kh5iTwrRw14i3gvtrtcAEZZnq6IFSA
bdtT1Mjy34F6xyMLAME82momK9p2ht9E+wQ0ETp1POS1Apmw5vViOhqpaqDkjfspXNKtoCXdR0d9
5di+PV1CIkQCxWrCrU6zwwdHRXbVNPzDq4xTwb2FKlEyy8oJ2Gzv02r0SQOKa+jtU9uKRS//1NmW
rlFTUO+2sCUpS+92PUnj8TXbEqg2McxuFSLjkcG8nH+KQf/yVs7dn7t8DGR9fP4X4NRc78j05PsN
yGD/JR5OQemWgIFmk98ZKeqlqTtFcC0Jhu8J2O8CAwwWiMIaAXqZK/kGksmWDKpicOuEKOpeQl9z
zzfh+aR38LFzKNoBg1qevN+9QQpNni/digj8FtsxKM+8OPgLJu95+X/WMlBCPgo0Mt2pA72nJeWE
PQfhYlktiLPawhWtQrxP4q+BeGZQzPMymTTIi7/PyFA8RzF8ba7y7uUUdBUb9DWSbp9eW930EW6T
xyjG013NL3ADo3K+TTz+C5EZshD8hJ+mio3L7ciULZFKI/2DLP8VZtsiVg86c7UQk9N7+sPa0HEo
yJr8RCA0mrHw0pPqHdmOVNzBuhwBaWz+MxZ4NoBkyO97DFqhFPujL4DDeHPaT6jwBqiojsEc0Mvc
cWExMwNYh4f2c7+GD4sEPHGiFrJedgUvuE4yt+6VHMcr2ZbqC/gZ+M7PQcdgcfJWYGk2XOY/GQlV
KWXtwbVLwHI5E0zpuTZtGHcLxgoKM24yQ3JRE4FRyG72m22jB5t82KIvktHbehVETMf7+FMkj+hO
tisCp5njhJtmVEZC6unxyLZ9R1MydtA6DuBaFGOyZR3DRZ00O4Fr9YcHJdxYZBsXnENZnP/QS44Y
JIpOquwg7JpPdOZ/BxRXBNQtM6IgFHyMbtExZh0u31XmiOZ+kza2nA6dvCTnQ5IchAA1D65LSoS0
Fxi93+FiYPzpxGO8FHsUhulxBjAyeYT8ojWvvzeA09e0mjrq8QWdc3KB5sGv/qiAwyivnc8TZx8x
SuBT6hLvYcP3DEmY24WQRGnSxWLzKg+OeyYO7Bib9VNaRXu9CSFsjQn/u2de3iC1qmZF9FJmQUs1
n0mY0bgF3qwB2dEuGK/Ieh8IXh/d7N0fwi8AyhNPN+TlnQ7BJJVcmNrJDEkiploWQGWOHXTDQvJ4
PSL2HBnAbak9voHn/DHGdQ4J3eaFA4dUtdCM8hKJ6e5WhUrd2T6/Mc+DYDc7zoBSRoYnMjOhPEqw
t/cBP2dWzeci9zUf9NHoXbjLqgB1ZvhL9+8fyRaEnWb2ze+cy7ER2ocjvdx+m/sunUE2I1fNf1TY
siufCTU+E54lrFpZ6oY8ZKfucKgI0ucitAGf44qmD5k7Gqc37weq6bPq3bzRR2zJvWqP5uQWrCeG
hWEnx010SUkas4od9BjoY77cNNVKaRenwajt3jPddD4zXrq2G3NXov1xOYdWHdSpvo1eZIiY+JbB
Y3iZMzn3rwdd39euwoBDd5gfmuT9BZc+O7pl4fSzeecSxQTh1bJU8tJjksuK6zPbtdgMsY8Xjpr3
Zag1ndE4X44dWxITSMpz2WcwTjw6emCrq/DjROUUPZ2Lb7psum76Iu12bXdAJm55Kzz8auo2Kiwt
Tdnw9pJV2B9x2TKfaFseZHK2aMkKqbPAJ4hEx53+a11VRqWdw0/5Qoms9RdM+fu7mwclgYO5+IB5
sEFogWSaf427prhH8OT5tqmqpGxto5yOZLajQS0ssfdDj/82l+bG3KPFOgKypztPXmOWdZgW0Jp7
BVbmc0dBKR+LIfvoPW+d1DVRFIJhqv1JrGhKtd7dauwPExWOMUmi+eHb+A2pf+FKO+LjpdcByfrd
q/IqZzlD8jU+bRLYweI0OkanPaKNcVcgZpx46Dd7NjRobAfdobxq66xe5xtZbgvkCXWF5JXSNryp
SUJIdfjfFuhGZurgGQ/JqJvs+yaIs7LxNDh93G8U4jzQRPw3NcIR1KtZ6iLzPAMWy20v6iiFwl7L
NNylXctzpKo+n9trVcGF51WtpzgWwK4ZE6amit1uqRuL9U6bs4QMQoC8R5wWCyRqw3h02A6cc9e4
gZl72KO+v3X8uRwfrrcSjj3OKqlbMdgZ6bT4RaLMx+SfyiUYLv9tAiw3BFH85dBciUnUeYt8JtPO
aCs3V0IwUPoFQAeRC5UsmTQpneszBQf3fdjJnB8NrCi+Bv8gREQDVJ8Xr7sL0bXuS1Mlf6Ug2t8u
/QD7sqlo4Vzv6C72a6dbASUGNf9n2ON5Y3CxbsKprkF/IwaCb6XZWn7haPIH/JQxQxO2rvcjznaY
qeuzoAnBSpkmhULbepaVIQMnWgpDXie237yQaVDbWuZu3VpLpWOxV1jUXvLrL+OZucbMa3eQIuKB
DzDWaGARjOjPssgyeS0XZgWJ+6dzV6FfBPRoG5yCYJVma5Dl+UeuG8OW6UevKFzGl2dJpLFrsoIR
EDCSvtSjbRMCaP42i+WLgz+yORZj+tXuW3NuUT/TyFtR+H1UmGtgqgauyDUjuNUpCSHBkgmwiPKg
qMzfItnIVNf5d5uIAMFQI/bGPd0PkV0Z1sNojs63XNgMzgj+4eno/edwFIBLVlBeWSh6YUKXUNe8
GcJCBtX4Rln1tcQXT0b4Fjj5NoeaUU062sp3kRoEIihlXiBxthIUwWnxFjgfHrGLil2b4zlDGVNJ
HOzMP9w7SBr7QhX5Xsay2sOaD3FcExm+YVvndgWewvPRat4Y5Rm4tqfKAR4dwGnyZGimJ6yGiOTS
R7y1PWNiBEeFYAJh9FtJWY7CSi5cVWs/6fW0iADnwUnQlQ9TZs4sN3R4xjl/+CMa/tke9woTGDw0
5PQ0++SgpJb+DzRA6iHoVf6/Zo0plB80Fa3O4bT/q5mGWDAat1pETBpdEAZxLEaxN+qv1kGMgHft
9OiJAsSpQ28l779kuIKut+lfq94hn6ECiyeO+Tirt8H4BhFjinQFmglqE3tyf7NaXOuJMU483LU+
31iJUckstsiXtWMk8Y9UQIGRiY4mH0R8P9b1BsVcCB3II/gi26pe6lvDkiKgeU2DGHByuzFFzqJ8
nEj6+PmK6jnyLY2EMDTSKaqjtKtCCgWXRUCUrXJ16/Tp3dZjHGo8LxjauNNoQetcCGyrPV0QhLB3
Dx8Q6Hr0x3mfQWjTGYFQufwjsA6he0VNdMQvm9YruYUdVe+8ORwZciojVWivtO59tytXu3Lk0JWY
VTrcJchW+61J8By4LMfOZJ1U7qV2rtcPxgJ6XtxGMHdmnOvtp1QFxK5GDHCf9nfsFpDbWpVBk4JA
Q54InlaqDR7TShkk7/axwqxJgK5HuRLFzvJvHn/iUdriFDF5oo8KYjNNCMxzps/x3vKsoauAL1nE
C0UQ/cfpdFRi2WM90v6YcSaBj2BZSkbioUKptKxYjH1b9wILLHzllD60SG1LdLjfHPF59xj732EE
Orec6CKkab5XJz6o+MAsk9iVEqFpJv1ZY+NlzM3IJW4y7AGYPpqwEEk1N7NEbArMQGMrjf6g+rh6
/NKzsmpKG7ZJFMINYFj9oEsXDcvrGg37iI+W/cjgLtEDc8vMwWKPutd0YmjGWvhXvJz9WVHQAs4X
Wr5uJdW6it3Jrbp0uTqBVvHcFjbi9XX0I+QbPYABep6AUzS9ZFp04cdqJTfEVSRUigi3SF5Dvlc9
XF4bi2FApytv9BMYVUqWBdXR65x0RsJo0KTcSt1St4FCw4bSD4IJ/lULdtGt7YdWDjsv+7H4l/vx
W11L9OyHlV/UBm+aNFk5axSxvK5b7suYP1OzFhLG1rgrHJss5kz5qJpmOa4Ngtk5KhVyCM8fLQ0r
DiBBkufl5KHzpjDWngqcTit/VXtUW0A2WSv3oUKy2gM7pi9GWARmP8tW//wRx04hqtxruqjT69WX
ZpoJnCNLp/KKrJxL2WMdR9CL0824/2ObYFMI6YpuHRjLxTadvhahbrlRzOYHWgxqFa82h61Mctwl
aGTOtf0tgSlZU3jmBfJs8YzwbSXx/FRJ6YXQeQYnpgnbTL1vmfttgCvMhlsSCh+6tpan7vqBQVo2
SmKL53MUF3Op3pzYBkSrHtM9fdEWgI3bwPKJnIQ/cX2KWkVvI363GzhqOZ/YcL5v6s0XBeqZ33vB
i7ybTLOsZCbOJfnAX9cv52CR5H128oozhCpeS1y2jFP3rH017+Ba3Gjc27V4VbVVj19Ijk/OPxsx
H6ouJi+eWg/ok9p+SYV8P0D734HJZX3ULtfZmcFhWOSdw7Q+8p/B2c7jfplGoIdTU6vGi6Jjj4fs
QyfQEOUuXn+ZQxaBbtt4sHEwg6UTHMFw3n7zHm4RhvgL1YwxBAmxauSupp4UTYTJt/Y9ibMEgIPr
tgl9/fIydXTkksVJmhgQUx1ZcY2UnJ5ZH3lgWqeLzeAL6UPbJdQ8unJFjRk0icMNVASF/9hW5QwD
oIw+mW+omjDk2aVd6iNg6xcGUH8KNMcFuW8Ui5ogl3FIrBQgQBeG3z3GpZE07d5TJLBkGxO/R+cp
z1wY0eXiRvtB0YsbOCg1YGVOU1dZumIMRDpILofZNyfkD2shUuuoxEJ+2Qd+MVXbuKer6d9ggYYu
wjQ7KkVYCAghFLGraNvHm/ewEtNm4oGx+NpIvxsUC3E3NnNoyeBXiHd8lspB1evkkIt8UDY1qNRJ
gttTndsvAcV5Y9n33VFLRZdB7fKGVm+7rYyZaamZAsnMGyrWaCrX+bDXX67Xo/IAd7AoZUPwVoi2
bZJJKCc7eO9DbKxU64Led8mVU2iPo1Gf5W7jQj6YLkS8mR5fvONMCKSLaJp0QYOV0cVh5pF4Yp5Z
jczGK2vysWeQvK75koKrW6yIF+E/1Ph6+qSmG0fgySG9L95U8FyMcku19FBoLznrpITt3tfm9NqS
OElAvksQd2uP8LwuO4L0ALCFqopVT33rvJqd9tict0jbTXRmF7qvuqTXUTsxFurn88iszsfok0+T
bFnBknwLNA9mubmk7d853qyZlh3qX3CCj1pyEQXw1LD5eC7IDvaOnI2kOczqrUwO6pFPijgEkT0R
OdsoD7xxvGa7I4QKFqidc8iQS60IiPFymEfnleH5Y4tYxNTQDPJSnlO7PM9WtjBk2MBbdaWogdTr
11KXVbU+31nauGmBfVzJ+2MtGFCWrgI5zhcAFeuBToWwbxHHKdJ4EEnib9gwhDnmv3GXKUAlFg40
U2TAPh89wbB89xsXRYv+mAkPl6+F0AmiRKyRUSNJ4a8F0CYoxPUdTd/it4AmN+Y/cunuOwbUYSaX
G4ZsYDGWpoBv9JR/ZrcYLg960bzXqVNrzeEoWWe7b3qdjbKInriuBY0tm5Sp/QR9hJSH/xSv3KZ7
OK9KKcs7u8/kebVN7jZ+1X6V8DuPRfQxItfBcTRCXL3Wt/CohzfP3ZG0EZknVA0Fu3Vu79EfsC7T
NIWwiEaWjyGI6pOV+v2fvm6eXt7fIFeycA9O/kVuiwM0yf1HfdcTgFNnaRVul3I7RhN0tDjnkKUG
EamjC8o352I/QMzu9x+17KYy2iYA5vNaXGohGZFrsNlAAC6vWMWvzxSjOn+WojiE8H2MF6KNp3D0
rrFlTeVWcJAO5YI3+fQff7lujcMACgGIDVspANWvLWbY2f1MehQxrhDOadKc6haCxk3DSwe32/Y8
QzAvMpOJ5gr88sBYfoN348eiQ1mGkoXwedLDHLwFJtYwN6Y5Lf+E1TfptylGci/bZfgKB7MFmLrA
L6/vZjRMVVzjhbBozCmrvqU4EObcAUltVbmnOg2nLdAWkE+JGfA8SyHJR2hYHcpOXW01JAm5AR4Y
RqH3s24AApRBhr2CMEiAAHFN0PCrP97PZwNMfvYi0z7sJ7qRqOlK3u3LGK1J7D7T7Q7/VNE1iQdy
8s52PUSGO7kgy3NjeAsT/0OywKH7rFUN3I17hyF/CHeMQ520QJUPRAPFPHPogxwzDJJNQytw3dt5
jrgMox79ACV5rnole0XrprFSuz3NbQrQBqbtZmbm/bya9zZB+9YqR3OFRBhSu/VKhUUAue2DI6Vp
ug5TD+ltMP0tq8AQmwwuokwh/a5yfkGf3+kqOSd+vVJ55p1OrL9YLVfZftxxGxlLGyZcJ3o8oMif
9KfN+LHEHFG+9iHDlSA8dM4xv3wr+Halr2MqBbo0eyxtMF7K9pW6QafBW8YjzlYrXlB7+ELketZV
WLQNvz235MG9F3iOBCxSoaHwmjdN777JhmH+3VcIStG4yXgwTh/arsXcYtsgg3K2CArW3eEztfVD
MJsAtQnGNZ6GpBUGNgWBLkTbByyiTGRrys4T5CvPmV8hSkhjx7ceM/quBcV6oeddVdX+GrhxRLcF
tju6/+XWWAcrqRldV2iZouualvNtLh19uOggm1o942anaY63meRHPDh3qk/wVtdPWXRibctqTecT
p6w5n9ppfjdEUFT3d6+RY8dOaog8iEp8Lcp3yp7uig5hmTpajUo5whi3WvvcjnjfXv4GILfE6T1v
GqBqFmasJzrThYzjcfTyzzFGmFTZeaiWm/K5BSvROFAar1HfciM9pcFzzExSyLhWqKS3r8q6IO+l
6lbQ2aCpfo4gKuJ5m2DTyDmASlIK7YTcpn/HBXNtgpbZVCEEmfsL+gy3DIr/npCu98KdrQXtJYn8
9e/Uo9y9s69ckpRRLPuKgfGWmXyy9Gd9wSkag7pn95paSJ9ZqFRCAqwKdvkkGscAxvLPlgE+zJsW
Z3P/qiz78Zzhlhd71JmeAWPRgowXpGFYZQ1kR+Uikx9boy5gLFNP+82xHqRVWpZ6kDngHg0jhDHd
RzNDdMVeMhpZMaJNliPCjN9qu1itOqEEEcjv6CVKo1AKt/Qb3Wv0OzUvRApQ30zQIKgZ0Zk3Wx13
GZ+gb3i6nb3lmflD0wXql6lxvseoS5wHpDtUjWlROAOArHV6AJJoMm1kLj7JY9cl+k0CBEEzKskn
IPYiAHvs6Ux80vAX/gwY8ozuxrKFJ0i2dozfXu9nMH4VcoZf2peup+CApgwINzmJPyHFJ58SlsVU
v6hFmUwNfz4BQ3CJHr00Tqg7KiRpaexEGG4/BY4RPgnBTAgo9+aahD9pJ3kcxQspult30rMLqPTn
uTqus7hZ46EIZng/JU2xEXTlKnecz7gmPaLkOZu47VuFjwCt5yAnu3bU0jMYjF0fGFA2Uut2eozc
KJxFveCUKHiD3EFS5r7XwYZ5aIsluZ+35xaebg+SSsfW0VqXvYMg6f86eSeXva7boeauroZfidAk
uKDqAPSmEXnNOPoKt5LuQw0eiBdeTiColgAxUSfZ6ymGlHfU+MI4lMujGZN3eI6eVz8f3WrEnUFD
zimQmtfhAVBbM6MfcUxs1uTpa4L87Nb7uPLmioJLzBXvEs92pxgvdmjzRosY0kQUYWoW3nwT9ypZ
SxSy1B6/NpFoBLKz21qYNkWZXvEp/6LWCkbn2rr1bJwLqCmjNYizhE6//j05h8P5D8iQP3yRT/qm
1htZ1Wbpje4pSHCMN6w2nYi+e9+rmmRjoVpXL0tLio4MfNTmy/R4Z6jeHTHhBy9evmie6rJfTKMl
71tv7IiK0R9XgG4GQmZYduBKuG9PmZv0WkjGcCNRAa9gcv3TrPmS52fbOzilk3Bjd7nVcZfhEAZ3
kRUoqzSSyU1/Xk+/8cusCj3UioZtxvQaPgw7/uguqL47VEx2RK9nGoVeUeVnJlwWJUImz+U6FJit
HLOpiFxW7rwSseOi5CJfiJU5Nxj9a7f+xb+UyW0/8247QhMzYBJWQ4Gb6u005NhfcHKh9swD9MaS
0hl+9WMAxgCcxmgtatcSOs37ayXHCbHFV5fe088Q4NJ+0P9XmaErFympJYUut4aRNSZv/lOhye4p
0bmaFXCx/8vCG9AlRd/WzmLt89JGwTUUusUMrbbN4+RsdprcdCV8Our0Hlsmrh2ZL7rJ1LHdxebP
ur1M0LyNOKiQhK+kgq/p/q+gp8G74gb0jqo5gS2pSHix1s7dnzHF4n5G/d27RWIoOGoNdlRsMbpx
69udRwLoueg1VIAub4pDuvpZGWzFi0M/0tcYJHOrtf84EzkCE0wDB+J34WWO4y4SDJjHldkErhEY
f7fshutpKGwX9MOOqSqsATMCX/LeGVsSEyRCNMiwlAoLWmxfMOA+lSEiwzhdEQOSSB3OLBnyb7Hc
FOL1JixWk5zLTPVmMDj9Mlr/aZjCArzy9GLu4H1+z5WEQ999faZItaI8SBdsFQSTHw9nvEm44e/p
cHS6wtWhNhhdFZ5ERPTXXJ/UrJRtvO4EHTGBhkqfN2hRE+Y9/rHH0SKWTZhoPVbPSI3t2Pp2D6B4
iU/tLJdnnm6o+C6xnK0C4MR8aiFUZJIk2DwzQjkWClaovuNEpVidcylzG03x3RfXxhq/ExTI27/y
jfS6vqteuqtSEs+B9x87HsiMWY68EBRXh6FNs9O9qHfpK27fcmuH7M+ALP3TQL2AXYJCsjmNX9OW
UqHyBVz2NQFa0EeIQQEfaDfWL5wn6VOkfDvG5PiY9t5ImTFvzstf/+C6qMPJ3Zhz587d4v4aHnFB
lWefO32nP0Il/20k9mMZ7K3pps7ULkLrAtRzmk+9CKM0AeUrYbbJrOMKAeOOlwGYMt7I7coggUaK
EpKPleND7+AWjTx/48CvjeQbr9CF+ufk1/UJhUD+GlvMnCU81wvI7jdJt0Zv1iHKpsr51eNH5nsx
K3awlvbFWDds9Jm1Rv0Y/WaCrWTLeWrfY9+AazrkAmdVYwW1wBr2ap1Us+8YCeT88YfSXuLL5ZSU
qvgeauN5CKG6MBMzIuuCqHG0GkWMl9bgxKLfGH18xHrf0l4HPOLvr9j1hTY5/ab4Fn8jsVrmw957
nfP9zoRZhD5I7rmzkjntMkWWGr9Sr2pqig2Dn2aFgQdoaTDnScNILn2H0d/pC3h+30TE5u0NYjXm
1nuxtrJuuIpedE+UkXfv30GwZpC+pYjwAOXYiG8+VldpljejMzTmn2RkhDNLUr6pO/Sq9JDcSSka
umRr4+1fwCOpn2awiOT2aVdhMozqZ4UUBPOO51c67lNUlz5jjZ0s+dBebMTj025Mw6jJfQvcLpe6
jmV0xBqUFT2NPHdRQb1cmlLHDp4Pujv+Ceelr+FeuyX/ew3tcwnmIzvmp1Srb453sgAb+vJ5o62/
/L5Z+3gQX/aL67nhhVyyT6Va1hZXehdEd3tKqXhkPPx5G6DNxMDVVrwTBcq2UlicZfjX4QpTmU3l
nCLZMhLv44RCMC8Xg91yuN3Q6NzBKZouCixvrkchq5QGN9C1oJIKs8uUmWKJdb2+cRaKDjm4BH01
A5XavZd/nruXP7ESQtpsnBpt+EhFviyDMTk5Osgy+Mt9+ziC355Abu49iVIXMwoqbxmggxI0nxyd
Z/S5g/zktQTOPyT4ofXZuqxtUyUwcV7UyxTC0QVL6q7XGJS9pXqVM0Bf98BdeSHQNGUx4jRlvKxn
rYgiFPKSluTuZFrNvHuF116pLrkG2W8atPSR8IZSVMfGiYwtd+QSllcX80B6FWMyyKWMgWgdrVwO
L0xxcyoSC/CgPM3iJeI4jkbx3Mwa1UHK0Ia4lEy9gmtgZpyLLfCx94H/UvdVCx9VQT51ctWXeww4
VrMa86HQDmnBjI/wl1AvKj+ba4+K4pOuQSDLCG8+N/MuYnyAY58iQQCAdTqxC5IFcLPLS/lH/gh9
qHc5vJ0fR28W7NXdoxvXpfVrkNJ5eLs1ChVxJGLm26AdfJlY4ej6pbuz3GFUeB7ozovATQdvxOsW
j4AuHj6w7G78PeNzzlXvFPONI5z62OtuMgNCTcxZ1Ipkkq3xiWSDKUHlvCTKcZR6cY7JJNXLgw7O
hwsGwNmjqkp6N2TINRJCSeLWy4LWccZn4VcruTeUICPUHsnDBc934qBwewdNeA1o4wFPtmlIaJrB
qZUQAPX8yDEB21Hn1SC+ejIhjL8sf212bJDvNxDHz8Kfa4jfG9QmrimbXjhHdCxLNo4l/m5a09zx
NOBFRDzvLOpr4+n06oUH4j2KndwWOKvaPcY0OprrH5gvhg6MHWGDrT5G4J36OyN5TzmZ+6TJzE5h
AdYaVRM4SMTeXILwoxDT1GxoEEvQkw1QN5iHeC4vc5L8gXDMNqyrHFilbWqgAUvWgA2I45FPUoWz
x10JwYYW5lQRqDpxQbOayWX/rG/c2sa8ysUdLWWZwtU2Z6Fv+e3U5CXMVPloVyJB/2i26Gy8FFDX
LF64agCAKR5FBAm0RYVWi0wgDJubeIC7NtYASeI8Hm/ZltJKfylp1ZpW01TLBX6SlitHI4cCAVIF
5FMFoNfyTEHQ+vm1QwUZDE4vEGkViYPApN8zbrVKBsl1eof+aA9EbdAcDSqzLrNTJ2Px+fSv5U/I
gsZbe/gQS6NQblMJ5Fs3DQAeGR/rHJKPiIQ7pYeofe+pHhfV0gHceFbm7KCHVwH9buBogM6AK42Q
neBVPFLvyY6VdiTmFUvIHBr5+gy+vttgybo2ssPIT4UmIqTGxe4T4At+S+SZG7LFxawBrVfkEUzo
LOaPG1/zdtLtf1Sq7WiXsWwfDpe4OdAEApH8C5u7tkF+PG1c1H28xDmcuvZVb6rzANNG9w9WQZJD
vZz1e3Q7ijm+DeOMvSI2orp2XUDZvr+6s2FwSOT0LggLvInCVl8xSEreaPkhyIdz952xcRA/yWXo
yxYJR8gzP/Iu0gkslWXnkvhNvNBaRYjZp71bya92gPuIgSAmcb5lMVHTsP87Lx0+b45Vsaf83VEK
eZNbPXT7QpLp8eFG6MsdSjdOSEvqS+wYiiiBXdXbhJwTJ21QuKGuM1W8gYkhBnzds6UCqwlKVIN4
z/VDQUsKSQsl3hrWyLpS98A9COaOMFMbkgP9AVAthcqwEsoEYDJIdwVIUeh7E5SfeEWOxu5eM4qQ
NSHe1ZyPYoVLY1NXH9KHc1GaTVon4C8Tbq6P0fP/1/W8Y5Q0pqzA82re802NgfK14aKOXnhHvNlK
9giJopkeJTM8J/Hc4C1OJtdzfPFm/0u0M2xiPohVnttd6sd92vPvzZgAZtEnIGKXRWcGdAazzK0p
uhw9uaROYEcMjfjtn9/uvcaphutK/Lbv1iTdoq4Q34p2sSdIIky78hO49nAHRYK41gqM5yBbCSxb
4UFtYpR27mpMx3d8XtFkQ2EWV8qQND+eEV7YWSLK1fY8FvSnNzGhzi6U/7zEoRTAFTyX/ypMf+a4
/wdf5P04+xDEVbJ7DEa3HMCJdQIsPc+02Xq9i+8dqYAoZp/kjCPzaVLiFzBJlMzAOVbAtTKVxLo7
Uuy2f9FMhwX4pBZYLYOR/s7XRxGVrWU4B4/tjdPVLpYfEzTN1s+P0Z+3d0wgLHktF7zOYs2Ky5gc
UMpqajvfTpNc1p1O0Svi+I1okAY68s/EQltVazR58ZoJmknYSFlZvtJUfNse4Z++JgmLp1rHmMXQ
E2C8qmLVIufbTVE8L2+GH5eRLO9hnQCoE5yuMcwiEp7pcskbUWTK+lkJX+W8Sqg9uqIYpBbb9ltY
+bndeN9lKe3X14UqI4AXupuNuZf+L6zZ3fxIKNRqE//KAkDM/R1uaihGf1xMaZoCpFaSwbUIWwLk
rHExAJlb+C9RmQRl6AVkX/xF9F8ddBRUyin9GlbKTIrsTY0CduCvVigWzZ1kYGNIqh+jFLYFQkpM
TQ3LrUJ+sTdr22CS/FFn5bCxHwL3f1QRJcv5HsPH6ZVxj73pbRvik9Z2bS9R4Kqk0RjLknIp8XwE
1744Bmg9mYtUbsiAYIQqfb0rCz/AN63cU+LUjLBK93Up1KeFwF1OXVGyB7y7KXIEoDq4tFoU6OiW
+Db9a2om/7ZkaGvvkf6MGmFUHUgXMvusDhH0gTFenKEbFMD7y8TEFNEF5kwc/JeLuaWb25Ngr6JJ
htRn56HkdzYGcc8MB9NYyO/Oh+ECfS3jaHGUIsnpt3sKHvUX4K5cc15E/2VksvpC1DIpfm70I4gL
612BywbUPSICZz6M+NSQXF/K4rZbdUEHgYT6TBmDQs5gS8A81EqwLy+xuj3hMW8hrfSkh5WVQ6pt
P4EwDL347TM7n5PlUavVtpRkoxyo9CuhfWbkvQH+N3wFJc3pYegPf/pKQSSJll0KXQS/jlyaRvYD
Em2YTETpie3kPn/kThgl1vIqipvVSqqaBW8ruaW7A0lvajTmEspfGYCezkx/8wdBBvEp8FjjRYM6
t8REDPjj+juhrdWfRRyr7VHiUu81NexSLuKmx6fSsGjnMLFL/Xm4cgGV2QjRymZTWJloQdzuBqyN
1uT/ye6RS0TrfNRhdxofniPun5mOi2O7ELORWbHmTp1tfRvbjQQbsA9Md3EKvDzzB33cL2UJjCaM
1WXLuNkiLlpblLTIDsFrx7zGLQ0kDY+d/y4D1YPvS5hx8AGB8TM0GTSg+6vFYnmVMCJSQAK/o606
Vqafk25ROPVHsiwr9p5MbtMj3oiGRUvnwdrI5oqiRg5Rn3HcXq/p8VGQrSMs21jbxllNcXBf4V7b
Xq+ehcAbA8J9KH/tnYvR2yfsMcOP0Ol6ZGQrPnxpYAyKX65LjCCLvBnX25WDLJ69G7QJjSB3N0T0
5JCkfdL1grArY+OAE/a0keavdCTU2LIMzhRYlaE59zjSDsxYZOLHXbhAkbpMtYs39+VMdueszf1Y
NxHLG7+36B0Wv1W+NU0sYwsgWkiim+WLVwLOh/8wODmjDbEvN0adT/075t9kzuejtqIpJR9N94G0
Sks+2hOf/LLzO1EhPrx1InkHkC1p7bCTvB3iZ7wQxRftCGmijsZzBJe2vnM41vj3N0KmZQ6VqFBH
S8PZVKvreSQTwmNismwlcaWq9DebGwoHDeI7AHU/09YHxexHQLvNUDBE7MOVTv4d6N5TaXMnp/li
zs1sD8UE0p6NIVo5PZr2YMn6NQyRS6Zbp3BjndqpxFxZf0pI8TpOACiGfLFGZm/3ymTcC4Qqw2aL
rbNEmxL26yOidVsZzQ0IUO/XC+YpacGro1suy9aOpEmtbMBBJJdkHtQ41biT0ioxpxKelRNHdR1O
hYzKN6Qvlna2DKnkJpVSyZP7ePt1nfSeSR1xvCBLZKBWWXBgNvLhV6fgCwhm5IzU/ee5NTAxdt9S
+7q0UwE0VL2IkKrqZ+YfbF0hVmDH1+bSuwkQxLnH8Ajq8Pyzao0E9RPeyzhXzXo0+27Lrm4a5lhR
AXGcKgAWOAhltOaszO0mjtZeFNd+naS36dDP5YzLuTOaeew4Hqy7frWBGqxN/1jbP0RxL9UprHln
lW22tTl/3KEg4gxb9kpnqCRfLzoraFbWXFedKHhsA8gZpdt7bMRxhGwmoq85cFlYK4G/3NJieKL3
0bNfe0S20q71INAEKp1VUh51U5d+TJ9qaXBlJV+GHg5OV1CYBXVfA9Ed5g0CfV0qaXabr7jlDD2n
p7fTFBtYkNfh8bPJCVrApn7D3bciXfEjVAAnmbANlN427E5f9HlK4cINWCk8d6MoNs55dlgMnywR
G5OMFl3ER+Wdga68e117m/NpyqXXZZVbaGhizN/Cg+WysN77XEMb6e7yDLxSQLPCETAClZ023f89
bRFX+ysKnVWn19+nzn2h62zdy39A3MgRGybaSDfIy4tCH+NWkC1YFfoQ+ZEIOr5jAXHcDdn0vpIw
sOqQIOwEvW598aov+MlnVpI2BssqTTGSdAP42STKTLE34JWVbvV78xh20GGeQg76LNrYnuwtvrWJ
WLyiNL6j3307sMfrSLBBdNBxIcz+9no36uVQkUMOm6PXcIVGfiXgMsaj3Fu17p5FB7y43F3Y0wRT
1FKz2udeyzLXXh1Cv/ViLANEQHO5IZkQ/rCjE3Q4zh19XrnFFezRLXpA+Oejo2MQzlE6STyVFf86
oCmwL5B1nE6Ylf5HZe0tVV6GmIlPiANpnIuWP8ggXslhfTS+wfneGTXwhpml75BhFMKGfrUyZwJh
3TEu3l9zwMeahzgJkX7oDjFkOC/7+IsqS2ORxyI5N8Y6RON8l91ctrt7a767QF/7He8YXnkL3XmU
Kqwi6AyEiZ3YTek7b/tuibI+SURcPMosV3vt/tgRvEVepGpbakLCB8hvPeB9fC+R3RFYHQ+j+Qzi
hFCvFULaTIqNy3+BXLedJ2mxWhDCAuhg9kPyXmlIFsjC8e9AKAj0xsrnrCejFFTfm1t1+EXRh75Q
o1ALRj+M4l/57GT5A8ibzZp5sl0d6MccAP3eeVGb9JORKXj/T7ut7ky6aa3g8qsYYxzADptpHDa9
4I9IpdzWQvbr7+ymNpuSf4qcZbokvDJs/SYHnGoVVqaeewMGEB6lfYF3DPIBNFDzGbbM71JT9NUt
VqUFw0yebY0qt7NDPOtekpLuM9WGVRvtCNAoMx8ZJIxvOvj9UIhwd8LWl6WvUp+LvhPcYvbRDnRT
QiJmMDTK5TOQkzuKHaE6c55PhAz1+oFDRNVGY0RYMFJot/2zIOu/Mr8Zv8K1JXrUORGGU+jNEnRA
6JG9aHBcVGzStmcWAWF8Qc5kDrQ04T6mLLQ1PqnFUaIan3pKLXWmYcaXVbrSX5/XxebvVEZcDLgG
KG7HP05hVX7x5NpsodEbWt6FG5N3ZBBNqfw82WoEGWkdFOMQiETuRiO5JJATz29w0Zg3enidwNCY
FxpSQGB7rs8UeiCZMOe+uqL202+reAj8F+SgkvUCljUxFg3+FnZe80L80B/orVY8Xn1e550XoxcQ
j+kON33fn57MmIK2gC+cPq8a54Ff02OezaW/FtAQkjHYGRuJmkI9/sC3GEyPpJxwXm1kr2+5coGO
NFOidnRCOLCa4M8bALT/JkZ+jILghduanqXr6lE76J6fQH/fjMzu1NzHH+8tEGMQTVTtyFFOiiui
mCRztnz0jYR7cLanaPlqQ/kKjKGRV7it8puxB78H364eVKi+Ucs5O/DYtTo2mHmJ6SO6eMm0l3+P
iaNW6FM6grZzPaHqlyw1FkmU7Bo17dZFuLQXaH7TXN7R5AoibKzwr5EvEOAKVTWy06vQdXUJYolz
YLU7zSUqguGRMj/9ApsrnW80SjZMcMB/w3eX/RPDzkslg+4I8zGoNejfm2Txaq8/JpTShzuA2pgg
MwYdyn6DNjB5YcfWGi7g1wTieC2hpPZS2pege6PKTnpIUsfZ8dwsr7+zA2LqomIjTD1gR8ctrIM2
mew4zn5PO2uXGS7atcgy3T0Xap4NCGLiNwKEEv4OjfMJVdJFzdcahQ7wPlKyky9OcOs0Gg1V0d9I
GExJQY65Ts8/pCEBMyfm7+TdvEAEjYZeiqyk9QU/uhr055HOsFn8vEU5jr4otHBGJOsymdy+LWZF
tFZGZrrizsiSgJbt177cNbxPcNVv2VNlnAXwTB60B/DlXsKfZfUPISAgkSQCZe/nZzzStnRGXvxn
qnHEaJ1ymb+hsSmc1inxQF2apBEeF1TDOlYF/ccX4xOO5wMYDoHcAXdt7DkK0bpvS2Xt31EuLC4H
GOuP9JCZoosKijBqO3nCjG83JRgHERJr7b4toKz+dgJahJlkAsQNrcksHH934QKV8n+2kB641q5g
yYTQJQi0MO5MvJi3cn+/tAHidht24q0HUp3DaSrtTPni3BbBJk4/ocCnH+bolluuumSMyh79+DMd
ot6YFn/cp9EePfjJ/XsPbFwZYxswoVW2vhIGQFn1xRfj9yUuSYJZR8+uowfba/KNyv3Q5qNkvyOY
tWtcNp7ZdYT98vlFrIT1N7syVrQfiCULHmJ0Co3CFWyiR/wTgXbSGhzfQkuYHMvuMcoaHNXFAeiH
WPSEF7LbqvPah2UPz2nZdoUtCwnSgeIMFhUbQnKnacIhQdceVOSbsfi5/6IFksYSil6p8RF6Mjp+
IIGnPQKOebbgWihxkJ7tmsPxExXDm3EJK1hsIvW8ZoUOCXNhFmjnWuLXrGMKPseidNKWZqFV4FGL
oCfUlJHWQX+iESDHlbnJD+go2maVXCI4b53HaxQWccQeIoBsvRuu+A0O1ucRjzsZwQPuQE7X2k1C
ihw40dkUaeQ120J0sqBHqoZrAezmHkl7drRa2NcKsOEqoyBAkPNR2ccuPaB6mrRkI2SMM6obHFzs
t2CH3JbVKMzVtgsfuEzjU2C7IimLtge/Rp6maKEEamMuDOE3K8YWyDUB9MGZh1sSWfIDi18RkjbD
wqYkAcoD5nrIo/Vc+g8esALHWCGh8RYzu6GcvG2CatjmIhstXfmQoWvC9ctSz3d7WC4eEWnz/fAc
LEFePLLmrxTzjTzrcq+xYz5JPNplxmve4usjW6iPQGyB0ECjHgQEtAo0NsWrdLqwItuql8d27+Wo
pUiN8iQZVL6w4P6J3uYUX55Q4MztHgenBxp1C2TETvohvGKc+3nBJQwcXbcujqQJmj4QyfeanhgB
lZkRQpxBoJThrTBuV4XjzLIVPscLeLeXngwN/aUcPSo+6nS2EupRRJEgEd446Wkpbj7WQ7AEvSgZ
PQNhGdOwWqU6HeFAWM7JHkvDo+GKH+ecNg12mnSrjwDdZXrnN6lOhbgHDVVnuNYC5eweX3MO0JPQ
T9ChPdwdMrL+SaVUqMIZYE61+JP7B5vGteF5X5xQ6ivinpitzOVLskIbSVCVqdt10siyuHlixZQf
JrNo1+7mfZWGYldhHWYpOx5Fw2SCM43Hrc52evnZtzW45qh84MuOODa74SJpZULwwls4QL/UNZqP
w30xx3xWsUc0xSHpA8JssgBDp24nU6KWmV4xT6b6riSg3cHTUd8ibUBvNJBeXcdSj1+rTI2aFFKH
8zU1fAOnYfOX3v82wyDYEm7wVgpxmuZvsWIAA4oSsDlvKq1VmKqT3Y4ysjNaIokN31LhXD65b/Wr
jr12fyzpE43Z08RHqh8r+HD8X+DjV7wNhsmLNvYJY92ytLQh6+7VHr/MfAn1726E9S5sfbZtaGpV
65e5dxembq5bTPvFV0wBdTBOOMKQ3qOpMyGAmEqcOX3DVojJPMOxF0MV8C2OOrCsmh9H8iwUCJrr
8rXKTU3wKBwAY0aQ1Mnw8wIOsBU9XSUZ6oddJXdvsmilQByvEYpdtO93VOJGFnEcA126jEAaIMEJ
/C9A9Tm6Att7djMxqUSNRH353CZUPTH0Z4VEySLuqzBIQwWptOcgS8vaJ+0+0VWrcrbRG/+CnWRI
VE5x9vTLKD8/grOKDcWCtlZZNeIl9IIxe9FWr4jzhjzujdFS1SSJYNC8T8G63FZ35heBcqzgfF3d
Fz0JKJSuNvkyzP/7NXssTBj8zRh33uxhx6XYtTbqKaoBcsuhUIscc8LPkh+sQbLMtNlAv/X5mzyU
u/xUqy88qYZElFyTA2zVC3WYWpxmyJ8Au7QL+u2kxUhzEr0oBmAOKYstzfp0NWMam1FA62mJTnbe
I9wbIFoS5LmBpHxF+JuEQG7C6qY3u6rdkoximmVO1ycMTicoZqfULARySfkZVMosAZjttjnr8Xw8
lhY77godiJLnYFTGgpzaauMYs6aOI+ZEaacUN9jvC7/wqDfYQjMc1UadATrQU7JiHJfcE5rEDezY
HAxPxxllbyVivE6AsxyNX9XcdxLQqRRIlhkJVi/IxQ6dNtYUpPCu3Rxsnff9YTaGwF/nB1j6PGOq
WK4Y+83UU/imcSlxEgECWqja/q2jLmcl1D19y/ACEWB96XQYomA+5QAxg6lDu+hpeu8uaxYqbAa1
AtcOhxghLH0F+PGhgVeA4IGCdeRs/AMcvC0S7QLRHe06q2IhQDFEeBBEwJQEXAKBGOLplQqEHfga
kZGb+pTZvn+GiBudURnptD5x0/qKLA+CCSj8ELAIgc+VkXtTbEU8ELlRPEfxqGImcLq4WA+aB1O3
PSQ1+maT+ceIkL+FAUghWuimta8by2qpgsYNTCpCp2G8or1L9t8485wcSm5I71JEvYEvYyputX1L
WRBRUsO2Ru9iMPHRAss7EZugMSKqlEMBLP7DDQjxnx9IzN0i/cCmZUTxgc5oBwMgAjOprXmAmqZ0
N3dxHlP3F52VBhdqVaPOcGrKnAzLjqGy9p4LMuT4lhpV0zXVCbieNrIRE/IQ4yhwWBgjZ8mSCtVm
u+t5Ka2UPgXEwq8Nw0kOqungT6jKifEnq8lH3rALsEW/bufH5a0Qu7LMoPOtDOiWqOBLHNBV80Ih
bUEzClNhniMhlM6Wn1inWaA2Kr5vMCDRTBN/SuEOEczwKqnmrIDacKUgEwr0ayyKooVHpMfZTD2N
HFNpDlsNzSWA2mP/t0+DU85aVrlq6KXji/sM0iWYJsgWIaIk28pmdTShUe74P7VnI3WgKXtK4voj
yHs/3R0TvII8qb9e10R+/T/xDCkgyfX8MvztTxx6CYciyz+UB/nH9Xm5oCA5IVtBdLK3yOQPn0W7
Bi3DpKtZLKVx8jxThWrBDA6rDdqaIjt9g2AyIUVfQ9CiTAbrvAqtmyPqofQ8AJVnTjA8wB3FkgRX
zzq+DygHj8LIBYIWrtFJpk5nq0fbwbuiTnFWzCSTzgPL/ajLObxl/2Pr6gEVNiaUtr+IE13xXqk+
2PbZj1brHDZtKd6aXIrXUM9e6J4I4X2HOV9nWrsFPwUYHOCTp5HEaH6nm9BTAgL81PeSrRL84xX9
17kA1wG/uyPTjy3kU5SUgAy5/SnF3/PLjB3k3Bph1EnoaMf8YU2Ng9O3ONp/kFSamVFtie064Eze
6957Zs25feWgUe8JSzNLbymNksVyDoxrLstkcI5wVqueRTIWUUCRRm7r3G7jBtn4CVudjRSL9VcL
pO0VXk2zpnMoZSNDYe/GrwRzsmXFFtLuzdC9rEOx2lm4qZIIiPjdTExuolVOg3+KNojkIPaSVo/A
r1/3Ae41NtWNYpIaisIJQ3wVuyBycZL+dR+jtjMwR0hF2xR1DP1JGIlzyVQkTEojut4MzgGqKYna
iE4N0NXBVO6qPcBB+cV4yuJmXqp62KXrZgZTg8TbRwpm8mTLhMS86bCEWg2ggVV+p4ET0HFYrLNH
7/2ikX53pYXnOOTA/1Nfshml/do18CLTLuXx+26+cb4s6FhcF7hWDH1scQApSmgcCBgpZuobuaWk
X7r+jnTAuDrKq+UpA0MqV4yeSmCC4blYGIO47Ad2Z4vs18NdF11fm6ubLCOCPTodcXc+muM1y1xU
2NvWnOpA1Ac/cNNimzALRQobPzIQjkR3uNxr1vE/ldorhsK9rPUdgWfq602C2XtfFDRPRwCq/KUL
B0CsPl8awe0l39LjkvlBkvbkCXE+0ctd8TbJ5JrMJ5NVTlBwPBXb6uElDYiOK87qfpCK8tS/tcLi
TEnj1F2OQl5ruP+GTuA7JaMVTR4wsUrHw/zZx2FAih1CwjiOw0xHqLy0bnEQ9gf3olw5H/p8buY1
BHOv7HT4sc+/HheI0AbVQpV8lDLX9BpdgKC4Bk9aH8JmRCkN8oyxMLKu8BmOsZ4e0Jiov1AJB/ZS
8bzGht5Xy4qhaLt0KBoqGs/q//JtXcO9RA2grCRrzd2JzrkjmUShPbGlgaBYuQ0GDy4rIYxlQi2h
jFsGBqzBgJJqqbiQzrN9VQ9mJ9m+F925Nu7rZ1sXCO67BBDKNTQmLxcic/0u0F0RGC1jwiwLrJr8
tXaXDyTD8XL8mLYU2R1dpAIHH1wBZaWE5aLUptv/czqJ6/T2bAmpBDYSuecT8wacvoM1Wb8qLKpb
dyeqN0R38vmHyWYtQd0gCoUK+OsKWDwQsnnjdrwlk6smdE3K20rYvh/xL0q0d0t7VzhY0hn3qaSm
CrwXmim53oJ4QzN6eQDUCK44K1oBXqWdfiqfbyeyrHvxCnur5iwzZMRIe+kFwYbdOBjDhlIE7xR4
halOOgG95JH9wr7bThcDx2oXL9Z2p9QXO8j4M2SYRG2Yd4zC6FjsKFYpW5KGxUyd/YaFsScrhMsy
7hME9pRMgnkEbF1fm6k1DR0HKO3JG0+R69v1mGjZ40NHczCaO0qzUCy3QGhtSblKSMB5VWcRZmIU
YxLIKU7e2r39/J430anZsmeuCIy8gbcFD63qVQ8Uz6V2MugCQHBInbMAzZbxssKba78aglRAYWKf
Ul8ajPA3O1CkTT54eaM/yzmZfoeGaoZFLt4IFnqUsAPgzEHpQJga068MTYzehoyf8MhQNc3oOWnp
lmQXqIF7Pe9hbe/v8X3ZpRyW/7wDSp4ODYmuSHtFRSIyyMZnAsyqPh+JMRsHtPWptLKQ0ghbtk/Z
k+GvFHG9/C2zPpkTpA+qhjW50ReRxp4eBAOCK78IUqBWGExTmmx3QpXmpjOVfWajUVbiqFsP+ruZ
RBClWoh1LUWbFhJIaGECgSky1w3vCJzebGqeYd8sIPN9OkSCgfu6Kk/ifzU6P8hwW4edgw460thp
I2DOJ4Xlc/+kI6joGzg2wr0miJhkbFBpoKpFVvrtjItATfJ2uSiHsOG6Yn3J690RD8gWQCB3/CET
+7a/anQacoLyBMyDbzt9VjSJyU1DXH4orWxg3m6TLkXHiBOOimGvvK5QvBo1J+a7XJYQTl8I21zO
DODiQkSnV6kply/KsfoV9Pvtsr+1uZhf6yamPgVpZpmhX71aDY2RiSDlfkMtD62HDJA/uAI+rS9x
zbXlrO0PIBPPdxYUe4bWYpYdMZWEdqa0Tx7B0/amB0miAXax/jhbDwT9/KHG2GUrYrciUsfLvUr+
rg+0cwkGLPxDcWuy4gJmZcXMwHu+FUFuAeKHRBNdiq4k/u2mJAbHWK0rlCuJOBXOIGs9u5mGrm/O
5VTFvVKhaHejYJFARCbP84xON902PApZfxMK/TazqGJB5QzY4WpJzWvIRDY1l1z/Q6rrrw27foH3
rjs9rPOXoIl+unQNMk90SJQD6HpjZsos0Ji7edvmRVkpbSKIBG18Mc0ih6lObV8taiCNw5vWRgla
qX1SMs2n4g3cX3O8f91Sk47/2WSTXJXW18tF4lTZ9quwJ4KBnhoBrWbRaqWHTggWOvHjbIhPPdQ+
B+PoQTY1EITB5Vc7FqIk2TNZ5EdY/BGx4ACk91IR732DgHf03fm2YeWcMOqh0vCkZuCMcl2JBZdn
Fqbi4lxJw0QoFHDS66No7Ncts1C6X4fnwDGuOKZfMElxe84rJekXxZycTicH9ZnSjHeFt6rbsQCZ
YlMjqxAObgvjQeN2uOnmhR02ySmdHZWprWrUqj3T6gXX4ft4bFZA+kEkSLPzwsv19+pTlHtNANOk
irPOEVIa62khZKUbxw2VAhHyQ4suXT//N5Zr1SXyRWQVVb5ewOvkAjoin3phEKk9aPdkSKSK4wU4
xI4U+O6dRrh40iV4H837H0fgecWycK+TrCr4+RkujOwfNKhcOoC9iTupOdgnISlYMTq/7BP9cCQw
kt6jjDCwiJDZ2xQwq22bjJ7mYOgTXwOBPJWDzDeHNMK/ue8VJJR+pCLEayZ+ZuFp5z6B7J8xapU7
uv/Wiy27U6u3oaFAZfo6x0EP/Cco1UhjpgtUR2A5Ka5AMSmAcAtukiIoM/JhpUV8Wbt611OxCrp6
uEP4GrM4/ZC+tip0MHYkLlZNB6j6loIqQRchUtRrCUxsVPpsJRgqqO+tPxUZZ4AzUtfvQL9MZWj4
YiqiQFjyp5XI8dUW5otv9KCXrmbtTACJzUW2rx22C533tvlEzgoa4La0LuRytKLY2cw3kW6kOMw0
6YIczPGbHVyAIIikVlTpYnlwdpj/HmyaexI6hFo6Rc1svhPlCzHJrCtlotZz6sq2XrihAqvxm6xG
FfUAqKM+8Q5t+gQfI2Nm2eXICD0MLI12gOF6qDNsJ02yVvq4jFlbej+iHiU19baFamQ03jlsersQ
ua/qGolYpjnN5z2gLKUCR5No18NtYchogu+PjbXSW0pvyAsOcEUw6u+Cz/oYOX22AO2Cg8QmIlR0
LyprlmF/XDk6tI+eANBGrz6NQgz3FB4/J2y/tFeoRhgw72CYHYWmQSjCGmiiToIhUJ1FvSDhYCp7
AeLKjeFchTPXx9GOw64LEJmf7BMs5SltAlNRYWTYdYmw7RdZFNEHtK5zoct70wXITTg9SbrxPNzG
ouCr/J5g1c8c6ESF+RS+/Gm0gUCVXIYSrkb16OmMzt9bLaZ84DeugnFToL1+CST3U1b2B3/wKtEv
B2GYJ3vA7q5O4Okh7Jt/qj+x395cIs/EwWl0pzPT/pqgDI1LuXSAZ0eoWZHGkHUDL47wai8EqmAw
zVafnCVSKr7VHSy9WFKuA903GZw/Urb6yj9jhlbdso7/HLYVUf+Rj6ZtUJ/jhHBLbzcFLAAq299N
keSLX8iaAPL2fmvsrJYfhBfoiKrh77FYyXRykA4XYR86CYYzqR5rjMJ2ucsKSHipKLSCCJrlN7yk
SCcTcp3ye/Hu9knuGlucom8orrkg/PYYct4ratWrzuqDT6oxPGGyFDH4yxgqtS2yGMrJ89uqhST2
qy3feo4JmSOPx19nnpGj7JTS9vGtSlibTh+PayIkTUYMcRN46mKrfdOEn0i9hFxzRHYc8cl1Tyu7
XUfKWPQdx5apQ2vmHAEMaRoYecOniBTnSPXGt7+aBSqTEAnz8WVmZf2PFWqNfPuWucJdc4XroW2w
t8G0w0X5wwBCQmVBTqbEvJyRf/EjQu2mM5h5I5uKkUSAUEqMWxTj8STmSAmYTXmrhyUbPN+cJFbg
N498pD14Y14iAzjg6TrAbzSukFMD2dEN2Ka18kL4JEs87CFYM/nq03bn3W7fcAc5XLEDIzIyNxY3
L6DG1iXlxIE1C3fHMcq3qh2onVPp7mJ/yDmDx5HPOyFU8+hQXdeZQka7bT9g+SPTnaE+MB4ZB8DT
TXZUg/e+qjFTqeIZXcIgXdEd1LUOXoD/uitaKHTnQRASWo7rRXdUFdUhZrkA3FGg8w/63s8JwKu+
qit8LnU3owh7ks1uktz0XupDYlQSGQ3Xn+AiZFxPox5KyuxSfEcCEDmPzdgSf3uyLlR2Xq4WVDCb
mDELNFsTjZvrry0XuksmeyZuTKC9cOsFSMI03BfBTOdIJBTRWuF5VpLfMKLdnjzKIJVQPp1lOAaO
HHP/IkIzsOtHnI3/Y3bHGd5yMEvOAHXVwRPPBkxG/dt7Z5IogmlnA7gWQSVxt7PP/bon8IVArnBF
k38dC/k9wILjJuva+GDdepvZrRk0kDBUvABovDL5Ym2MG+MmfiSYd5jFyjZT/xo9XbM4/PP7xI4r
SwCgw45bq8Wqds9iT+N8lApbch7QV9bPzRJYc16qRo1s2wKv3Su90rR1ZGMp2UEbb2WNKjWMxass
iClaczB3t+dGMI22UKZb3kH1f+0gKZBLRR9yYpBLJC2G8ox7MpWL98mqmpFhoNL6vCg+V2kGxGir
Q0Z3VayMLoGhMd+uTTfk3dFhAoBuIOQAo4CJv5af1iHDlk8jrFEC4rXtaD5diKrE90oyLzHg8kp3
pXlkhkNENYnM1ooaO0fdRQnb8l6muV64OF0MI0LCuE8YPAewgaYN+MUXHS6loGu+7pyluB0B1tP/
4vgR7sVmNcH5A6xQ57p+XY0QgUcwgMtMozVeLDAPYW4EzhgUd4jQrQKl328J8/VwQTjceugmQk2z
pR9+P3+f9BslzeUEKCU4fHja1uThEWcqM3tsP7PlkkWITQdysLrFn/PvpH7hkpFg/UQGCjPkhOam
HKjTMr5OWHIKmAgdJWW7vogONHUeYT90WV9OcDPtl2dIawXe64Uq+6S1S1h8l2yKeSMyRwcyqItb
j38d8gGmNm+T8HOp3Mj+JzEEJAbOrF2568G011ApKc4HCLtxegzOeUee+yLMHhwnxLYFkpr+keuN
Z0DFVltt2oO3on2Ph7jdXfZOngPuWDHaCiHhkvEquuOFzw7TWw4+JtF8RAdursTOEsSRNMLpWDMW
PchjShqwlfluuVP49B6aIN7VtEEnsyGewjIdzWB/wlHS5uFU9D1Opzwk5GGWiaScIYUkTsQG0Wri
rZvENxgh3BRKCU4FOPjJf9Ruz1lyziVyMNV+dm1xCt5CGxXG85S+pu4JgJ6DMMR5fP2Wx2Q/NsrM
cMmvmJAz6h8CzFKDZA5jPt324gTk4VNENEaFzEKAKWvm2tQmkUC5eWOvkG7uLzCUEP735d+fZQQQ
BxnxFLU3Z3HPyNL/cmsxrzJPKJZrjmz3/mGhhH3ELCrzVI88WeHp878C829FOtdR64+g4S7s3NTg
bCZ4qHFDQRRz8TZjPFwBjTLc000qO2/aQ93qtGAv/jI9zC4zafStOS2ld8nXdpXAtS3R+8dMKf/V
dgaD8V3McALqWqbVPNk8/jsCwpg0AfO9mJPWShYXGztWxDKSlTSRSnTC2qkYHgnkT+OK0WseyCEx
2YehXMv+lz4iIj2XHm8f90b8usPEpzHMxdG9AruWczOQGScs2+GiMGsY1CMctZ1OEfY35KblokK/
WcocJrFPQ3lSqvk5V4wDDGo4bWJW437QzdZawd1PyN7+pdlUwonf5XFUmRCoRjGlxLbLXZM+2yJ+
m+Tf8Vn0oZUrxMe/AD8qnaAn/UYIMqIY0h0vbg1dFc25POXqFGMs1lbLDN67br5YOp3DU0KlO/qU
Ou/3EVUiCu2JN2T1H0x6idvk+1kObLIp+I9phTJSkjSbUvEXX3rlfFaDPU8XXWOhoPRBkbxhwr7F
xbcn+myUEwhVix/6QqhgYkg4NCZkpdm+JSRP5QkeXAD0o84XY9gNjO9pKQzPAWpCMr1SZYe3QzT4
5kkXUvT1qkgdEuIC4PDqE9+LcUt+AnieUqTLF7TzBWmnHQCA7ZVc7PQ+pRvxxKuveECSD2YXoxNd
Wpt7Rxih8hE7BjaJzTjUoHtV4obJLtcPMRqOieTbmZyXfsr3cfLuHw4af8ar68nIEmn/+dYfHY6n
OlqSNIthwZ0X/rQfdV3ZjKMd5DgBNew/k6KFtcJA/tb/fJ/s/mKWHK5ZsqkozjGupWUIoD7vbZCr
k6yqBSqZD1mA8eb12E3W47CRInsIc3x1BH+SVSR7z7W71TF7WjPk1dPk/XCgWJZe4E/Py73lso1O
wxvaYrMMYiZYplEzw1DRxlFeBPn3jsKYrn02MZ6QM3RBPErPsrMNDOjHrbzNkbjgzl3D82Gkl9Cg
jYmyDCTLnp4yeeyNBbeavRhL4WT+0qBBmILDMoDwFRf0Yy8+dldx6VIlM5azUL2txo7JHIAy4COi
reEXyyeGIPhP2Gyapg+Q5gUlNJYME/fTRcFq6XqmrRCQsEA4SPtyIrW+ziScm/YLcnzQ/e/6AoXc
MiEYj4tvlpKpObknvXGb2KYRixkb/DCeEk+zTKjWUNaUFM1wOwsP6AaJfG6LVXhk2Sqm/WgWCGl3
YMr8z0IN+Nkk/PQWKSU0hhzGR0OhVmxUCNwgtYbILz5s8pCX2BNn1qsB4MVo9YC7IBLTzwpONaA7
GQLsi83Ul+gZ3lS5qqcUTtGkRCBHdvrleqysi52e9aoyAyicFWf+2kD6JohXzKgiXTqAPdj1JVTL
ciSG+GiWsEstNBuQSbbZrh8Q4jy+6VdLhu7wVnkNfm7TTMmCzYUovjeVaOA5Ps6Iv8xGzauZ1SSO
vWvMI3srOKsuXBOBsFAo9c0w/4DBLYCPuuUia6Kq2vasCIky2DvOcsxJt0U28uzyqZr9lZX3OGlg
jtm99/uP3ey6WeH10kQZ7LwLsbl/DQdw1zlMBwwPTYEoXsUxf62ZNFd2QqEW988o+NiNXtNQ8p5G
7Qzy2QHAGFNyZGJBltXFca/5UCjyoZQlL7EH5UY8ccm3sR4jF6Pjf2sRDfV6dqs+O9cuJhAXMeaS
G+A9CDCvButphQM7Q8LFn+nQ/1IH+2ZXcEgZMWktosEcIjJc5OTLx3P2Y5ns5EIdEpd36gmrGfXy
GW1CcCeMfofiwKoBeuLDy6SyXI6YW1w4kHxeyMmNMNUmY8vBIiRYRj8YpwGZXUt5SBjvODZ5C7be
jnXuTwIXqk7hAmvGsW6NtaJq7KgxME8MNW4kDtragkUjvKJxoizM+Tt4/h0pWOSQ+lCOqJ8WIj7P
F41N9o1xhV2Pj2ROJj1XoRpPoCIQKDTWBlhMIxO4J1yLUaCaNbe3kS06lcW1B5/xxRmzHB74+N8O
uZJZyaLVEeBhgDOKzDsI5DdcFnoTDVubN/2366dyloZDgAfVGLmFSdN4+CtkPwe0xJytYV5Q9dOe
2ula9lQ3XXrU2J6AtHhpR/ddIyC9W2onFtrthH/lMnQVH5QPmd32SbOBPrX0ZeECCGjtZ/KPANQG
2zuCMzUrvHVGV/34vy+qf3j3i3qr6FvZieP8FE4qerP/Oa6Ztfe2Mpfel3e6jmjtJcyLTaij+VYG
MoPKow8pl152Sfwg0vNHxV4QrnnwnDk4pja2b+fLvngWhF0Syv4RBOk/vY//xvQnyMpFYZjhzuO6
KEFimksl36sO7bXJMbBdG51Weux9bYRhfM9ZahmvUNeZPZ0hLuuUu04TSjudW9rjk0Tre9FGHFmE
QjqW6X0Vc2ErAyEvCA0pp394+x5MZu7U0Gj35u9E+6RxCW8wJS3dpPYQBAUcu8bu9p649bw8ftth
UY70vvoJ8Ro0sSsVL6vVN36r1Rve51SQO23biQ8FGGomh/Fa4s1hjsRXyusaIvvN7klkWuJrBlG3
SdDDxlLBkanITFRNwWCLpZVGZ/JuhgaOvd09YGNMa9fu0TmmvyGLZ47/qySetKlt/5gikIkuc6/i
gQVkJTuFN8WYulkGVlVBlmkhxf+kPpbqrMAR7TrqVrD/2EZib0ChYwpFGv3MUtcEKYiyLUmVBL/6
EvTwGMUKxw4Cm1IJfKsD8W8gKpb73ak5P/m8N5pvH/y3bSquirl893Ro95CPChbHmUWkgN5sNJ+a
neQSPKZlmMIEpGOt9iZ4yjRwYYKK4FjpeTaQ/pOSK37jCLLovRDvm4SEBCQZLzqpfmHGyS79u0+m
ZWzFMa+lS9mq9g2ASzQAmtEyPBFcWyir8vAs1IlrZFDJgqcOi17QlHvnhyVWG5rrUxyw8LJqGZrs
/OhBN8cyBrdmPwPheuajVeBLwzToOwxB74fmvw3j7aBrb6fKMC0ilgDSYbctAYNpAzb76rZBwfiL
EzUjTS6c188jJ9PY+yn7ljfkgxqxMWWETBsf1EkwOgeqppyWsY058etAO9OSDWhbHwRF9A5OpgJD
qmRqa82U1LSmVN5qWnWI/SwT8rGv+IdGUVmQr5TusYgDGDynvJNhRGexmwmJWS5hd7hxcbBhRXky
YDeT6s5Q5Gew5obHzRDfiZQUjsyPRolsjnPOoY4hte2YldB/NVHtkxrDAy3tSHMA+V1gzThp8R9p
M4m9gGSOo0hX9wvNGCmmVpvIpMMd3zteVt9tTTUfgItMknD7Rsk/XUtPrskqTkdfiFGhHjGypq27
hpkTnplTmKVQRRgT0pbPDaxE0HXAVWRi0193R54tF51YXpR9tf3oqJXSlrGSmF7m+o0+0Vt7WGll
ZAsgpY9jpm+xLekQ9CfN18RmtwNiVZb8mFH6O6ERgJe4iJ7egGo95nnp16FHob44DkItCVbKpnp5
hPvhQBko2+wIa8dN48b2jc3Gu7Wk5viNH6p6PAn+s7hWh/NKqPPFxbnJKW0Au2KeZjQEP/rcueqN
JEMVJVqCSdgA1yDHqwv+BmkyIanmANeoevsY7meV2uN492mTukWoSASLOySH7jIhI2C+QnlU43K0
dktkDMP6V/ZotFVo7T9xDcmKQbI5P1UtCTltYy0Li8DO0CtNgatdNijDTGNQYgNZF5EoZVsNCpGo
5BmKBmecW15/K6hkcKjrtceiOIISjW8tOgDwCd0YmCsYYxIiB1MpPue+AUb24dmMNt+2pj06Iq5Z
B1KfTgaOcI+LlB3wIyp9n/oRAa7gup/XytpsCaPWpdPsmThZBOWQCZ+rQakntIrjhGqg+jX3cF1E
9XZRarb3HqCNj60MJGOmA0viPf+hmjF910X0s5BDeTj5u7fzAtWPbbGvCZB4IGnw0ryKQvM3h28W
Wn/wcHzQYPrWzqkvhH76PwZGno7lrPbKi1DkA4NTeD6rVUmZpGUDsw+mjh3CmP7rRIKUQMApFPkS
R6keWxRVAFFyaZXvLeecOXcc6iytVRWCMWK2ki6UCudX2Uc1zplhL0K9kj+/wXuIbse4Uu/5kyDK
FCY5JfSY8SjHpSOjbCfvmPKggInTRL1l0vWiZ4/f7OYA1jIYA+WmfZiEAuUr9ggWpES4u3I90q14
y2Lxh58SZASh9JyYPYhQAbvPZmx4F8K+ZXSOpOKvZtHKHUsQHZGU3J99I20qrdsgdFBnCyHJRGcF
GH8ok820Yee3GELXcr3srTpUmPjq2sG11UNAmYwcE2R0HA5Anlh+ZNfouEkdCLbu3UAIXB91o6sz
Gh3/pADzxZKrJbYsVLenr52/kJsly4ii4BTSqzPzbHSy7oOYLgmQVf3ttPgOe3vMr7rbvhCezDHV
ZUePuSi2zQXUzI2mbCH1+3oVVX4h/AwWgJXENkBBD94TstV9FHFbdTgRgkyrF9fSdbHtSom+xR2r
KgDB2nsrrkWU69dBj5WItPiMwxyL/4PhC6lrrPoxMXJaqsxkeC1Ci1z42rRyX+cq2k6Pr4ZE4/oi
M2J3BfbRkeedK7aQMxlNkRbxNb5wTYJigz4x9l6ixmvLFxXtOoE5uPIL1trxZckRsABgIa9CBKuR
g3J0YZekDU8sHOzcbRXFugjBMppxDRSvmtM6F92AgNM7SWgkVFKUSn4rGGo2kScKgNX6kz21b+V1
h4yEd78WQnTIm6p4qkFjXbk7FbSjUGbZjB8KtPm5LmOhKAn6fM6uFiYbCBLaYnmXzFXJigyi75mJ
ZSq/LlP00bSWPCnYL+SYNfjtmLDA1gwtKj94+dte81VxnJmzzF4jsGvQwSMqghh0HUiTt7a92Gh5
Ry/gUL7bA+LsO6hIdePbcBT0bNlKIQeaRGRAX8gDMzLtPS/JZfVdv/UMQdIb9M74pKw6d2OmJXmE
a2laUy9U5TJCMCzsq4y7rR0k+pRuMxpr2yqdW7oou/icZmgX8TnJOt+PQBPDvQEMXi2O3SUdiXjF
MKfoUqyep1OBjh1rDlkjhuG8qF5ZAagso26D9FyzsQ4Te3PK8cxV/qrF1vn18Kv+6gs7yy1chpMN
Ntq6o7Eskq2ANfqHIbFb4KHIDj78lwel3eTDTkjqpgd6TchNTVWtoYVGctNWQk/ZvOk14aUI3hxC
KD1Ayyme9Zau8PIfSWs50qp86cjieTxa3Di+Cw28JRFprQf6kp38dNAuKhN7cBpOP3XPcXxQ6P39
B3lPvFv1MMXcrJ0CaXVw2MGwV6/rihTvvdIkqrxDe8Et5UCf998EJAEVRKBm+p5qYhcP1OIsWFcT
CjygQqLE6a7y1uMDO91+sIrJ5beMiXA0tcAYpyv1fCi/PvN1sd0POi8owf88g8vHrAgnLZVzeEZA
Y4jFYg8YPv9o04Db6we5ZKdos1to25266NheNEH6iG9hwQhacbjCeCgyex3AuckyoK8WocGRobc/
yvPYc9eZefS24Ne/Ldtg1QCuibBfDiPg08N+dgtaBPvsaJv4GOfZXcpZ/bVxwaJiBgdrqFtwdlQZ
JOSFQ0MZYHuaG3RP74MiVhbRYdgTgJXs9bxNIguDO59fvIBH/yG9Ji4o0ew4Sd/UtQLDtmII+hno
ntNbFgX8T8b800NvoA/kQQajqwO5I6TqYanro7q9agrX2jvdqzTdsejwNVRTDlGfQ0NQkXP7NeDl
rJZ3679LKNrYzECISaqUso0LPSy4GmSwxlOR5eW0eS4M+iXInV/9mQDJmVvHSMPRiPnal0IlUkYj
SPMP4s4d0GYvUPPLdZw4kfSLuoMur6Lv/iRdAf0YXW8W4j/jzWRm28IChkXSisp+h5aVg82Y9riZ
zEALzxz+yucgHu17KObfQOfKf88R2QwPyWfoNVz55XfXUPZ69O+3fhElVyXxxIeQBVrQgT1hsmGG
llBZbJpIKBXKfeb4hjPu7bgozwLSqYpF14tg+Alg5Hxc7pkPBXMT4LOKn2VxiZukGyYn+m+6yLtl
poeOTHrLMDi5nnkSYhwdZvz0zexoNdE9GmQ4/mjY1oB9Oso4tmk2OqKTCOs2iq2T87TK/pOxSKfO
vYw02JbB9t+LsRGJDHKZqbGjNNc8OEdEwIfSmVxuXZPWs78UD3NgbCNHQIQRlDBukwhgDvhdLHwm
1Q8UgNNZ0G3lqugMYmQgvTpcf1QiFlrmCPIqbg3uucSGBiAMFG3FxVvL6jmqiBRl5GY7kLwjMXIG
AyrwJl26wFJPmC1ltK0V1KysevhRB6uM6YcAS2lE8EtXoX+8fJss0w2La0ckaazTulDLPKf+2Jei
AAkEToe9Iu3P81xQDt28fHZ1Haw0y7g3nInPyEgrM0o2sokEnmRI6jvgkfkwNewmxPXgbiH2LaO6
8GeuOe6KXeK1R9roAFXHI4wRQVJeuBMBtUHdDRqGUlPxxIjcdeWC1KcsM0wXyyTIvR9gmqfRKjOZ
8+GKA7C5fwgAACLRscgg4uwscVLz+cFPUp2IfTMywmw0mAj79g0acy3XjbdIC7CF1GI+bmh0rlfz
Kj2sQ8ZMxMjJZUZzuFOBTUsU8m5Elkb4tthT70Xzxz+rDgxHJsRnhIJJl1zWJsXJ9HcokadxBWzR
rCm8sU83UvK2AwMItaEVUmqUQJ9TWCkeu7LvKTcXA9+gO+wWdjiwuMtM3jg1dSA27KlSUzjZZ6Xo
ahUkhV/eevPbxcDmsfkV7u/IxjXtPHddYDQqY7iQ/WE9zKry7zFJa52oQLuYB42i2SYKqtcjQcq8
OG9FSbPWc4s/2Tzv7CDS7wIj8sWeCFiZxVzQ/ktPz/GRHRvHsPBYTU/+MU09yDpsFdssri1BwIMe
U22vw9n2I5uzSz7PIUkQYQ2Ce98hl2q9HQgU1jPCubIBOl0MAW9d5P4kit1Jz1Umkzk+N0uTx2lE
Q5T5O+YYA94uXWdzAMM1vI8EoHKyoqBAj7/nXrZiXQyvQwJ0I9VwqZjMfC8gkwiY+wxz2fkXQtDV
pSVHyCNq00VFbc+kFvp5ppf3EtG1wepD1ex8ZnLF6phjZ1ZY3gxdvNS7YtbK+K2W1KiAyNdoFrVW
4rwfxnZNOEq7FWgTzvdJdpSvzFEnFlHfA0n1RfYfMhnVafuildxClGOIwdCaEFyHVkSdaeRsF2Mj
JZBcDbdKWfQespMb/Tr4nUmIHwGauHLnsR3XUxO0A8cyz2tZRICLvdkUBPJTwfmjX7XMpbr88gV5
JXoEI0zd9DqF5ZUkfZ+5nqjAoFTbfEN6WuiLBv4XaQ56o1cRvdWltnVnCG6hz9Uu/nGfu7mgUSnH
Ic73SQUAr1W/YagjeHRwMLzxQZ6nd2SfrhPFUbpxhdDlxVQnGHZhrOu6gqoiyyPbblWlxbl3tenb
6YGk47FSfGCDx2HusJA1wdm8HZRvu/iSAMKVWfp5gny+N92HctfoKk+nAdtGXFLtIWJffcFX6TcN
P13UQtNyGRJftSctEmIVoNR/IE0eBcmjhDz7nEypiow5L+FFsQjnwtpEZTyCPrGPJDeZo7eTpi4q
G+uzp54y5zKJeuvhhWfe06EsT+F7xl0lUiTOueP7QeqtIhYCS8QOntpV0k41TVah3yLFdUi4rm5j
nxMvbDqSQHgULS+9yWGS5CPouOPG+MJ7LIfEQh6f5JXpWl7TmFCozpDAlDKWizHhIVv9F77VPq9T
RwMldNNs2zoYykjyxqJrNoGtFtlhkVvxj53zJrZz159S3PYBXwBwcjJbVaGZG/UU7nfj2XIH+2m2
wJTPaltxDu7WitODjlRn5/bab4KKSTYZ9i6+Eo0/QOqEP4hiNW/NqePNm7l/v6buJGR4bBjH8Co1
lMvYc/wCvPhJKG54wp0Z00dylFOMq0ndwb0RdJdUQ9H82cjkZdK2p9/wrRiyzEtDL1x93pZN2nsS
djHPGJf5jLWLNbXVSnZNtU3xMY2IXY8adSWN1Rcfb+kx08lOlFNKEZxAqds+61wKeL3zppMEhJrc
KZZknwJNa5UY+Kc1p5NIeVPjG51BMMbeby4U/nV5RVbCO/aGjWzZ2PuYT3LxUO8GsLNf/Q415Nk7
T2QNGjjn5UMQEuEv7aiou2sGmKWuk/iui06vU9bpZN3GdKdSr4uC9l34iwwpTdKGmcxOsqE/liMZ
Me4sCbgm1CxBNHMqzpKWRcKxgmDKpevoKIwrPIw4gLLsChDlpqCnwT0zjScnVufJFxC7/cyapNQJ
NIoO4/z/+p8jkYrrZqqfG3kJ0LmK58NEX9JTOkxhJ6x8N3qkZognwpBg/jiYN+oLpRIrlz9h4ZDD
mminxVrSXEARurY+ein2dHhTOKyC0sLAu5zBzK+oeXwTolDkdFKUd27uCAoCzxIKhocptzcuG5Kf
V6WER7+VtmK5v85L2wLqI2U3rC47NKJJrp1+kG7Rl9yHDtwGu7X8iwlleP1FcDIbwRO47wzNZTDe
XDnoPwkUY56cKBkk4UkPcIOrTA8+tHNX/BcdGmGf7yjFTDp+PuME+yxJgKZaKAhcK56eEbxUd9QU
9nRk798EAFk7gOhEnTdQ+kyOYzpZsj2YuzcWgI788+SB/+hlZom+ql1vq8BmTBXtJYzn/GHa7Sie
7RvuyhmNT8mEh10zuc/cliY8wrLVL4BYwTDOkf2+mdwNdXfmOrCLN+1F5bfX6qXy2pQvb7vSJDN3
j09haHXUHmVOQhGzk/6m6B/ydWIsKQ2dJ/x1IKja21uQT5EgClPRNAWIpVLSgbpvhv00vJ/Fx4Wm
dl3wt6HdH3kKaIZfsY0WGdLtmkU1/8PACKlQRMPPgAwyczn40Xm8v38h3HSVR/8XGSFD+1xUf0nH
NpncL7+NNAjlIH3QANjmTLR6WtO9lUXVVgt1nD7kvxU5rYUl8h8EbxuzWMjbLXx/vOMWfkaSWB2H
MDSCAPHuNJ08fHUpPDxofA+YJ2EsA/iPBxpQ625wWiNGHw7eY55Nnv/XSPYJz+HWTGeDpT1+Qmsf
V6K4ItXk1bbd1Q8lj6W/+QzztzUUyULgXkStV4lqwVk0lf/RVCyjtFCgHASnqKrykS3K/8fUFqql
F30VBTK6E3KxQp/Qk1B7LIt2DumLnFOLNfn/oUFtTKVo7R1a0yelU9mMI0NuxR0Evnr8TlZpk+C4
XpOa4CGQwefoJ3mgZOK0nXhd5wRlI4ieo/K4wds7dQYHYSga6mZ7B/SOfuzRxkkyhxzDt+gU2zHA
KIFB4ZgXWwRHYGTP9NNc5cXLlDdWLzoaiYnoykH8UIkkZ1NDpb8DHtOdID6RFOzs2hUfahKGunsc
wQNzAqxIB60CgpI6cpfFXf2ybcTbAE3dp3sWQA3J7+MRNyvd8OY0u2tFqXeETRORySgihZcm1igb
aphlYAgnyXTi1dFlMZU5VIzJDEn+ZGeXiKvQQRZ+SHqYKGYh7owfzdodMSq9GGvAQCsk99SbQZEf
4o3qqauStuEgSnmPbNzIYDlSQ3U5kqO+gynsMNE7c19B2g8Z90p8D/QF+W2eZ2DOjQfSTd4Q5oHT
j8pFI+KfXGNBVj4AFqHItM3Ury0RNQOc3BQ8Gux8hIdBPHBCEGx8B8mksZxiRLlXDNohsK9FtDcV
ZtrVQf2LIa4B3NWgaRc5XpwKrZXq4sZqCMfhDgTp28F5StucPqk1CweP4E2rjz0H8d48/+DYYkLC
UxMGQN7tSRnMxp0Uxf+4ELY+4Q+bD16z4Jq86jiz5ZorNR07AWsPYf8WNiSn//LQvSkzWQ31qA+L
jK0a0lUr8hni+h+Q69Ebr2q6tpPlII8j/LPhOxN9UKENwby1Gwb2PJ1ll81nqXwgkbz6rtJ32ktU
hOakX7OHeO6LIVPTj35qOyTO6H3x2RUSmMOxJC+PfNvSP41mVFPr3QuoVz4Gq29H1cr9oldfkD3/
IOCe8NRN532EfZtEWBYC6PbBxAoCFjsjHjHJSbtdB7J7zNgQabk9oJzUMQuODGuXtIUTrjRpVOrl
e65lU53SZeCGIzpHaPZQwQRncHDRVSrmv/aTgGfTI/9Ce1zRVp82FXHAPl+MZvsPbe+e3igowff0
TEQFnIihr0VRWJm1W2Ec5dvdiOQOUBbTKLyFwIJvJZ6Y38HDcmQHlRZu/gryKIiHoGL0Co9j4NZP
MsYubz76LIMBgI9jlxSDBuKobyxnMFw/dtTS565gFWZfyIu2MyPy7vnqVps2kjmFFc0+ARMPaERh
GQT6xOHlANKnfWoh1qgzCdyxjuD8YQQOEpY2l896jIT3n6PmiNlCl6A4h+0QFaZ9ZupOOK0Ry6xC
W2M8ENsGyAuWb322nDrPNPDHXHoJR/JGTJfFpU4MqPQqX/eEI1DeP+6ddxC95iJlBjHZm5Vs1bC8
5xiKe3/9oNdvyayZEpZp7m9B+It2WYiZIcaXrWMjTsdXjJL1rlxt7aFFPqlSZTvf87WzGWzXmn1w
QoxnKv+ZhxBc5phKnRUelbm507O32XqnzcFysmnPUoXI422l4Wl0S6xlNo11VEi5wNny7S7qzb4p
fFEsdzwMSmBmS/w2JsFm60CZ/5pSKUBiH/d9AI+1Y0w3Alu1528pYKED8CrUqr36AKNci5dnsaDv
siGgUWrFYs8AUjYfPtdDtNcjisCuGi8FTPSA6G/D919dVCD2pU65EzFJ77z2vYuoTr6ofQvHUziq
Ry/iABZkKSy2Er8axP4wPOFsDZ3T9fsoH4eHKRD+4LtZOrCbCKWkz30pXoAaL6HCbLHJVPG30cP8
TygvtkA3fGZAgHi35z9bd0WGJeOgQ49kGMrXf6Oa3n6difkKhCSmaQsw9y9fsMXVjLxp4l3BrNOK
RqpVRLM43C+PZWx8IR2ipONiAU7dR31BzAhdZkE+D9GtUW+njCZJh/1hO3ZWKDuyiqunQtw1+hD8
EpKKlg0xwAKkSrRLzE6kkS8MV+qjO8hVgoX7dBKU/hdkIv6vQc4T24kecvpekI4KoC0pdWkPKjsA
ohuxL1fGACg0n8r4oxrmd5NNZ8//BTCcL5cYphFBnccbhAGVadx9wbBjepUgKVEk8a1dCydOmd1Y
zh9txrkJP4+mDXbvgmUu6qpVOfos68kdHvjpSOnNvNc6ekYTYdmsSQXX/A3kh67ZtTQC5r4215gp
2LRvVGrfxralGGBsshYE2l5f085ubL45bK+x76UgRrRB3LO3kgYijgSCMOsKSVSkqMl1dI+ef7qy
5dFQQeYvJnQ6WDi+682nnEL1Nb9e0eyz35EIN+mB/QTogmckCpkn9lqnpWAxso8D88Wpe7x0n6pQ
0OvIIino22RuIlIoVYLS+zXUvnoFgzVZSpLmj2k22r5x+NTATIiWLLj/2LjY7NTaEWP2y5ZP0rVS
B/j2RPsKBUgBtLKjYhW/cTZCQoORDX/dOiPOkoHtzjBNX4zWoEz1cf3d5YPAcmsoaPgBP6g76rCn
mzv66c0dcfhG+VVBYcN+uqXtULAVW7wUUmngdN5ejYJes048raHdOxg4NXvZaUt8F/eF5QuwvIBl
X2LuAahTJI2gbx3C0a+CUGVTHfL34qIVeD68GG6poE9bQ3Ss2PuB125KUUGg8smsmtRZiZn95xJ4
EnP9YUw76qWd+ifMjAm9zjxGaIeHFB8/gm0DX9ncx7eggT3PAGgRaytrspv+pAfGY1gk/vYOAo/i
bGiHUwlKDzDW6HOOkK+EVBjP4101Y1mGMpelAJSN2ao1u11DKaJdW6zYQu070ENZPdQerWm+4M73
x0o5hiLrx22ax5outw5LoveSI9hQhsKeBlYx2GmXwkrNl6nPAa1st7u+9Pu0VyrZph8g/54Q37Vb
RKgrwrCiamFLm3yFIuDAo9cqiOOVEEm/OeDOMtxE5eq8E+GD0EAfBSdpw9YFL4MTCiUHpBj9tJdw
aH9N36VlYe+jbmLZ3Iab/4mrK2xFsXAr5hHTY9k1Dtm26kCWLnCpX7SyWYX6WkEWzwonVAAFQQvr
fPkrkpmmwyDi3ek8fJ0/mSQ0v/iKlJY1raE6ljecvm+xv4PWN+osNWBgfh3zqqjAZWbwoF1awC77
VFwZ1+9DUpaEMSPM/nQREEtPxnIi8V4piHpTikqcCuNHpbZ94buGFovo7EmvGWEuP4Vu3hZ6skOu
cj2Wq/ouzGKjkRaplDmgljR2Zn1u56rm5H8s0syVOem2dm0GwKKZLZg0GtAOtR24ksNBT4QuyaHP
X/DBd9qZbAji3xrBZYTLQoKaMFJGNGvXJlLBKkgamWsIRiuXM5ShBj8C1kpiAdjCrvaCG1bWkCpX
BtrIvZN6eBd7SqLLbp+Hih4q7ymyDBzTx+jQSVlCOnXr64lVUL3I49GCFOGQ/pSSmIBRd310zxJj
EZ/C1pnFqEeJAKbB4iSfxsrSlRBU+YMyyb7pCQkuHqfqQZKLCfcEnUfrA1umFb8ZrgvARvBzBzvZ
JFJi82ApNpT12hm10y+7SdF3yW5+zzHxfYpBshf7rFmROOR2vswbJIlV1Kt0Bu++/9Vrk5yRuFn6
MJWh6UM8hRDCkn/GK3YHSoO0RFem2aGuxjSEWIJgOgD4weA9ilAyh8EDx7eSxVl4kPqXkaTiDDB9
B/73aIbicntVgGgD0EFSJvnlCUaW0JcQr6UApZk3wCoAbEQsA92goIvn2oz88hT/Zbue3UBfO/kH
uNbruxTehzC0GaaORyisH8wbwJPYcYwxC7vi4nGxqrxvnlxhkUF/6WRIYXf9DsTYTDnmCPhjDIbs
OnEPPKsqwJAi+0QQejH7gpaquahOXc2PpIFtbeSwIdpoxf/r2O1t+JAzpbDgCz0NItjSw5HBCXBy
BpK5t2rxPT+fKVK/Z805DycaBQ6bhf5zuaamuCANzgvE5H8HNpuNp8ByesPeoFlW8YTAtT0Ct5Ni
cWKNwiR8Zma9/KCEErDCi3p1k05vyESXgeSdt+OwJ0jTaa34ttbexVrYhSpA7OCP4qZqu22xnxjV
UQDc9THCtFJJrBKhVrAt02sQlEVdkW3HP3fm5GdldVfVf3UYzHp/ePE/k8GmIZ/b3Cz1vXAGfcww
HhS5HdXMujaB1ZyusVkM6XuI25tS9yKjftEV//HQdun9QBWLOAKaKAHa3DXY0io327s5A4hAiN6d
txprpVlCqqGgX6TH1MctCzOHPWSIcA+Ve34K3CCLLAetMn0MLoXEFT6/gZdpDh813SUHjZWclT/j
3q6FE3LDYBDUIY2GS+LfufqErFV8woYF9gWGMz2e8C9Unx4dCD8OBYOLke5F823y46Fn049AWuNe
j5OXnCT7EV5BSz2ofM9Z3iQOyFitHVC8/tQJzTRUuYuwKJU+SIogTq/oek+j/Q+031j8Bbakq4Sf
Fqo+uvCj17wWzxQdkGgMW3AcMG/2TOeWmNh4q5PA477dkdxBrra6IhKaBNgr2spM93HPlqJmuGW9
24H5zg1vMdWoBV5Oq9XDHq0lQR9Msw+3PotZTKdc0tIrpz17dP1nn9VVltStX63jnn2l74EEiZKn
7SNbpllfMZapuiiXCuZ9ufm0L4U66xVItk9mR3RWuVltFe8fNk6fCtPQ8S2yccnsa6GrDCFZnsHH
IRxO9ULBI8C5XQreQqomNOdU0F0M+ilNbTD0vqkeMQPhBp80Zxegkdycp3lCpIeXNB0LBP7ZSYmx
aZe7EopfEiIUN6OEeAAvmVUgLMRgJZk8bLd2vf3A/iIjxAvJUZ9gLvAyzbqT98gw5grrQnfmhRWi
1ucvSRka1G92MmdP/+FlZXTHaa4KaVNRQIjl2CVIZCOnKuP7ZfxRYBZfVjDnTz7u2SeO1DJVpTpm
ssEeMbUwcsK+t2QOjfYqKgjWpjbrELpCzBG6/AtzsJgaDiK7scz5tUeKk1fsyy9fY8ChMJKuX4l3
QeMNEaOz4mObp1P/avfheUWSFZ4BNOtLnr85K0h+VxM1mJjulDO82xBSD0LzR2ImEnxo86pCt0Sk
vgmLCskJkU4YJh5Mp0KPZBC+uSBfRHwm0zGm5KuwrCbCpwEhNv+TD8WPfR9TfrcHpuW7seltGMTF
rdJlBnJc0e2FpyWrWj4TnHYx37xPUuV16LoiC050ADupgmDy5W13roXjQ6QN+67D76/mzC0L68DO
EcsPK2QsDDjuHzO0aWuHKsm2mDAVxExInQHaT3foj1Xcu0RCVjiGFspl585SX7/8WvnnFRHyWg2R
idxe5QdO1wjKV6Ng0Mb5frKMjoedZSkDyImMYsx3cYz1FTsrWgrrI7tTb82M44y4m3O3VfzUiGFK
ZwzI1D9pzo1/XnYLaRZyb/K3yL/ksvg0evt7eU9+RwOla8RfisVEo8k8myKp/HWlVDWFAbekJgCW
dQA8UU/9/SvczORJD5sUQi1t9yCxzw5DsJWm+la7YZsvAkklN2B38lYz4o8FenQNL88MOh5nF7Xf
oAhqy36PxGDc/DlXAMqQC/+kdjcYfEE9CuzC0vTwXBARPNvbunHynZgvk16S7mXTzDByyCVLZyRH
UAtc8rW8loLc+74ie+PUm1zM2U4I9+M99gtAhMggvHVk430LOKe7mCDndRaLbtd8BWN08cRPwOjJ
ylCUALsUfa6kOcNLhj+WVj//cTZGA/RC0atu36HSJ3a8R/2AlbF9hUdvBLM3i4c68kl5ZpfT+tGP
fBwfcaubbua3qX66xddYCbFdvZuqIG+IF0hSROURz0jmvjZm9vQIKbbycJ8oTD+kMXVfm6ERXYs2
MDw7Jqs42gxsf+HrgkTCCYXaBA3lvRKPcpFjvPDYPogku/qxhEOKStPHi+h2meLVwNFuec0WoHjR
n3vdWpbzvWpDFAmj7Zd3nzF8T/xk6/VijRQimE7beeRPxyd6zEuC3YPy86IMtw5vNRre9H62/NU8
8DDwT/V6Bj7CK8HfCklJJrt4+nT+mbc5CJ29/1RkW0Od9c66acg9tovmOyLSuDi441PKHiIKWquP
NqUBF8/mNX2yGC2aZ3CA/3ja/URoSDoBA7t0tb7diWi+UTX1kxBCQWbqiySsTPaD3MoF6smDNkJE
hqT1wknU6Y87faVBYrsSdWAU1ZSR5vVBtEy+kmB0nX5o3VajC1iWTUZoXzmwJDxkyTYmoZ0GFniI
o89m05P5SnCdJGJOcj6eE8EoxBvQmHzmYmgj01Ax3+XAsJeRprJv7cAQYbS+XLOBdgl+xVjfmQWA
VZnBhXIYLAZWi5vV2YV4srMxGrAhmhiU9PFZt4xjW1TRItkN+N0lE5TMHgeaF+dfKF1INDGzANTM
Xc+7eRTauZgU3fpvv0ZhY7a3iJJUpBwjDUkwAFkDuURG+U9mN+ezdp9gaUwzf/SwH3KUZTaOqk4i
/oPMgfc6w6QJ+cpjtUPY3jv4LOTfXRZF3pNwn19BSqiMAVWufPF5qk/mfMXTLGkoRDT0kVbzD4ZA
3RGmSoPXu/0NqCzk0CQeL3suNPC8rOMDGM7Fa735pmSasuZADNJge7lMKM5WmTkI4oI9QmJ+Vah1
Su8keu0nE3lbSN06uV6M1RcxIulnTgiP1K+tndw09QdrXYGr8WDJ2LUGXFdFS4djxxt4qYtnD4xQ
e/rjj1oYavZBV2/7J8lBRE8asYUmNoUrdKYqN/aRF2w6epY5RbG4xRhyH/pUFwQHU2reEAP84noj
Y4+jiHXCw1ZsltkYULu0P9Y3+pAjOXeSQP7A3LDUFcAVEENOZIJxmP5NekwpZzzBIAMQAX23D4xu
rS7w9Oepp1HPEqhc5s6LzsyZT34Q/PcBElw0nTuVKQRJjP6lMCIAQ6IOZ6PLz5WSBsdcCS+uBt8H
UBrNKgcPYBI/THvkI+E8489UZLDme4BM1dvZxLCx3syWWkH77WuzHrZEynPA+TV9eN4ZkAB8tTfG
0Tjvp/TTnabAwwRJZWJSXJGRrmceZW+ogC/IjWztk6w1tTpHl2Y/eoTUhM2vfRY34sCGG4TjO/zo
+zVGM/KAjtRPB+yiO+/keUy7yR0rzEuKdXyIUtcCUiTqfLDnQp/hcXI/9/S2tHFaacT+lZmuT7d3
wWX5RJzgx5vcqNjXcLw0UJnCQR7Gv6dJrycHCLkqqUoRAOhI+Y0KXG/ZpFBSwKHJTp6oq3kPr5KK
wVxNNiwbsgjWlSiXLeHIa6j6F+bQHYRGUNPdXo0CIIIAcHZk5+9aIL/hQem/WdGtlap1klvbGK5s
wNOPOiSRQaS3hGlA5aX42W4W7/VNDcDofCGfJKKpOtbCH9yUhdk6hsIqMpZLP3SF2CVCx3YAYAaF
KQMlhRNQSmPRmcIymWToJWL3wyWY4sAkK8dXjmQjjLOxiOonsRZS7c6bOlAlobCkPApM4c3paGmH
r1aDfUDag9cmuu576GHpMmyGIHPFknl1e9aH+iOV3Z6NfSWP+BXVkzzbKh9nw8dm6YV8SY2+5NEQ
DgftLKUWlETBafxPjYo0oO4If20jWZKfN+VcUCYDVzLAcbPylFdvWnw+po9HONtScJdAruZY0xjx
VasYaxrH12sPPFgIbw0nZJoE7bzhgZa+z6ReX22LnctY11rHuRtD+gJytTPy/pERESCBZfyKoTsn
UPL/ppeOH+fHWU7jmG7nPV1bT/R7SjV5FxCiFUa3EsJkYl99dieb86KmytyCVIip1gONJ6e4WKh7
FBBkSAPmcNpWP2I4EDjMqabZEkPPYvjwG9cJSxfLTLqwnvbREhEgIZl/8xyJ+4RN2Ye2XGUaKRQG
FLq4jvc6KN0td8NyjRcj3GbbmhJuDOLO2wCaEKOVW4xrHRiolTBgh43YfF6RIQtdfH/ruxUpgk1s
mwWjLFm4Mnkdh2KjfC0FgmcRxTKByj9ze4D4YIQG4p0jOkEPSS9eWfXeJO54GxdgWSJrOHQRkT1C
JbPzBQw+BzgRo27Zj7NyTb1vMT9pDdy/KBVIk1gRXtaqaO+1If2OdugkrMylo46/L0qu7VZCHk0E
H+KmA3B3Z7wNKNLlFjFS0RdnD4Zdv+wvKmxdLuK4hsZ95HSd31B9OrsGWlzvUJELmQkUjwhId31G
6gBm4ZY3NV8XqLZhmwf6aQgyw6UaDR8R6m7sSl+pLHm9cjBB4mc6OCMQv6kFDDBEa7Nx0uIXGE68
tI+o0kwMHa9TPz0Ys/Tm/HK8ZtMsmyDfVzeZ3iqT4pzVVygIV1R5XWgI2w+dRrtSsw5akkzwql/a
uj81DAMm0aLqrCJVyOXi8orQTBlu8a97r4JNOz/roO5XyjluqTuy0xj5L38z1DMwz5i3tkp4alfj
5aP2VMFc0/K93GiCsGB8vG7Ya26F4rw/YUWLlPiyxn07vwiR5qeieLOpk2QNl8iYJTjZeYdDuQfC
q1GQqjF5hC5ol3pWKZjwqEt0yBJS/6jAbN3zvB9zYpGV+8UG1OttHUkAU0lUeuS9s/FGYh+s6Di7
4J7WfOMvljqepka/LLrtICfNnzLI3QTNkgWODHfe2Y+WgbXUS/i0pHOY0lrszfXl90O+DrwNDBN0
PII/1+OAqLZneflWlvHgOr49NaHG/UDsuEEt1nmL4bMChJkyiSzHZGNEYBZyM2AhvpNJkJ7PgDj3
oeXNEmEV8N3BvHOLywJkByiLfTPdw0WbYpDkR48bbp1hr4TzWTWuu/ayDnJyEU749aBq78RugePl
Ua2MF71aPO4nt7KGWl7/KLqAUBXXgk++pj+Uqsf43aKJLLIo6ndo01Db0WpeYODHGzNleAj84x50
KlbDXK3g0QVMeWsZj6kY0ov2F/Ju/rUkYOIfMxxcyyHNq8MqARDfYpwYZT5Pu3GuhDSrOjyQTkPW
JyK3iJkr8umh5tTnp900rRYSKmXAtUgZCMrebpg6v4GWsPQq7uvrnL5FAtB/Iip43ZRr/+EHCRjW
NdtjEYGeEQ+myBZa9HPBX6+Hu+g8B6VnxNiHCet96y8n5iH6EeKMMLt01meC1c11iBxyOEvs0WNE
phtuvzM90HGnORhaETqsiOIEcAMBWKvCZOXeAOEMxE3UkZTnObzTxhydqhsHkQw22jG8YQh6gLGQ
109w7ri3VaRqOINuxVHiCXmDrve1REKLHx1vfS2RxOGElpoKnhFwCrUqmV1l4NIwJD0EdnBaFooW
Q4xi46OFTikl0ZfTo7jXOP0S34visstMG9uhP/zwJleW3V5vPoWJ7YOpcZXYCGXBUcVnb9B1phpS
3RthcxXyaPKJ3ui4GCEGNDnKc5dXuHOnDzoaBMFDv5ex/P4fzTD1mK05nPzmmmkPPKeB5lHcGjv4
fhhQIAmiVget85XQG4i8BAWu+2iqEHt7klSwlGK1+TAX7uLpoR5zqcbAlVoaWFiY7uttdgn6eXwV
Nae82fVMA6XSEbQOmTcQZLDWw6SVnoCobMl0Y3eqysdLgXIJORQDiPD95uIFIoXI6ZyYaCp6foxl
hW7w7/dbFXs508/j3VLWSa+RjivmsL8Nb+/jEQLbzGhjfUV/HbsW8IXwwqcrspMT9kDzaWbp2imF
Y4VqGEWMvdndg/Mg6ajV5BdtCIwtZPQdMUxe4JgDmqpWH9WL3QtYE/7pFr6+4ip9tvJQIuAZJGNE
d4Wrrljw30D2inYOt16ol3sNBnrvwW9O6pqHlOcHvLN/moqSi+xiVH3jMmikCKIBTNZA/Dd5a+nT
5uhz4825eqbFA2zPYYXnGMyPYY/xnnOk4rY2IOnVbkGWKcdyVsj7C4DSyngO4cvpSAa5C2qtmPAf
S4TK/TnVDqdf1pFA74cIXsdz/ddQiUMVRBze0Sr4GyML1ndDHpQP+J6ZyOY4xWoUViaO+mGCjjND
WmDBVniC9lOuimdbz9bFgjR0LZBsX1BSN6tSPngESg28WhXei9I174yp3MUy8e72zEv4Z5+AC5X3
0DLjOzsL2YalQrQ+od8WB8yx6262wg8fgZo3QKnq8w8C7S3GzJ2Q2QGFAATbD4ajfou4wYkI5w/m
A4eK9BEGT9N5/H0waN3xIf0xFSP37IbbaGflk6YpU4m+RXCS3PG0jpUcn6kV06+5r3Lec0kSRECH
xPBFtgfZCx/uKoxeuB0kooQy03UgYYZsiZZ7u3Qr3EZ8Ns59OPm2r0QSWtYJpLWzia3VbFblpx1h
CqNw5pszPPco4UqKl0WRXYhuiYccXasTHYZGJCVA3Egmv1AU1oBS0c7jeJVvVIVwpHmnamCR+UY7
EjGTT/pNyUj90rW0XgWPPVbhl2rBBAoYiEXxc8ld/eGirzf540hg7mQ23ZYPAcVB1F2V+5azXX9x
6Llqca0D1H17v/GNX9QF6sQjCdS73d9zFfDc0oAROMCgGXESfXem2gf5rHexqnGHizHQ4en8B/sD
/Gf8/Us6DjGRknm5XnhTpQXdanLdS8HDjRu5DQzwlwltLjVhYchtcQ5ApkM1gKoIZHBEjl//Vae2
xZv9xX4/aMwKg/aC6EdWk5Z0kQEqAzFfbgRg+KTpH7XSCYBNeDrDGVw+WUXosAr8aPPc534mKdRp
0we1OskSgGW2y6MCz5kW00PafDpP6i39QNCAQ5/napj34fx1YxVmAUHzTxaV27gsV+pxSK7Zh4kI
PWX0W+8GmRLUV8J9vAswFEAQ2Ipemjs0OUy71mTrVd0SyQbfBxgA3k61L0fIfeEQrcb6xgVmTCs6
nPZZc54T9mcu8JbpehbgBC0ypCG6vUmtInmSB+IkiavjkAMOfEzAGIrDfE52c6Gu44PLoaxCfxUp
PavJjO1AZml9EQ3YpykUyHkMyLlG7+y5W70RTKBIVq2uTSegv5BgyZG/D/tCTwY6kxWukf7cErwV
ZTCBl5p9hdVu7KFFSBERNdp7eHC4COZAEs88XCjS07jXw5pGXp9Vp86IFVREtRapbJ15RrzKUEWi
1WQmIYNKPcbkppGmqSQ0x0GZIL3yA4HD5lPDcThDPStIvcFsaEv0swYPa9I9h6v7SBHfD1fN3T3r
btxZkHxLlN0DY+lHtBEtthteMLj1oZZ+mHVwcnoflSuvjvHrqZbAGGhJ1f/JudDLDwIHHooALeci
YOGeehhfGuBM17fPC5jDpK4RMdAenetwEs29vcx6jpixLiwiIHDoFFkfTE9SADQaAaQYd7o0qrW5
a/QkZ16AxkA3f4oW6Y6u1Ua33+092em2p4az1dQo3A7fnaA7szaKOaMJEnKT1U+VOdkyYrqOqKrY
srdBeqHBuuvuVsDqOpbSVolv+pt7FASY1D+exTtKlsahSTt2CBttx1/EKZ9AuOO7h7CoZGchfq48
eoYVNFlJu1QEuNgdAegEYZrcndM43ii+oVQ+0mQ8akJq92i2xslLcobJ6YxPmZuiaDM7a25QdgqW
CGaqhA0wXK7r1yly9pb9lUKfFzthJPzbpvbdag7PsAzlSUH8uZepVK2N503s+UaDjj+NHGHIUC42
tFjZki65/Yb1Qpv/bCNc5HacpGUjM0yuEYerv+e30pMafXX8Au1Rae1x3fCT6q2UDekgjDQIbISi
VRpbvrmc+7Fj1ZMjmMxXPq5jEZUsWJ3zUUaR81dfj9f2PTITC8ZhTcLUSISDU9Tmn8Qrt1Lx9v+Z
TWdvbKTaa1nWyd7QRYUdlUw9KR1Ze9Ckw8CBHZvD/r8I7Sc7m54094B1c7IYMFj78PMiKppuEQzO
3u4ddu20VGCzxoctXci9xlfMglE4LYSBe7xObCR267jWpPlbAXcWnZuZo1CC22tlmo3vVNPYuBL3
CLjdL36fQ5/omPGpZvy2n14il5PWYinaPp/KlpORSHBZDcLfaWjRsZ7uHL788KWPL8Wz3IjwMXJG
1RAW5gyfmsz8ArjeJo3BiOgF7hlKqm97K1KbUYtx4b/+/emj8e0bfHsNv36f39wvA7DHkqLLfgXc
H0ZSS+JMQPF9Bi/qU8GybN23NtHUdJfFxepNhpvyLMA+4jJPowAiD6f2w5kdCDepy3OJNzu5epvp
vMdFLFeuResQMoXrC+niuNG3qfFbAZhJtWLHDIJB76ecfnP66O2Dy6GhDXS+94qKgFvRCoYHZviQ
9Rwd46c74W8eECGy+3JIM4QlCEZ79Tw1UPtgc3lDNMBa5y/25ym7H0vTvvyLvJ9i9+XR+AbmE80u
9/xtZzGsymcNj5kvHeGt+uVrVKcqrMri+qqEtnG8VcIwo6/8lzOFlpWhbzzByDvT5HL1NzK1RRH0
yIZgyYqn229tYs0siM3B59plKUDEZomCf30/N/lEajM4CynrN2b0QeO698GMCpG6Q6o3JWgcO+Fk
iIFH+j81kmklVM2DesN8+KmBpb3PCgcL9S6AnlcjmR0Fr1rqc7UgBMds8koGGOQiDsjRs3dq4RGA
73cV4FUrBpA+bFlViFDk9AasH3Gs1gAhqE8rVDmwEBRfkJma/zAFQ9cW4mkVeStHF6va9/gqCxR2
jguA6qc8hxLEBjE2ePlwHtuxiXQHRRSl3+hk1Wt+RiPbBypkYAu6lgpGQ1PhYScMWroxN3o2gnr3
k1F2tqvI99YU8z9z78mEit7pgo9F6JRWz30xAKN9QQEua33QpJOyiRIYKC7fZmiBkS3MesxdFmEb
zQ+nsVF9h4WIhd0q1jAqMfn8wMeIhiAmd3K4r8FHm5atfHG8wVRzamOHt0Ab5jn8jaJY2X+fLtfH
5+yKCuMJK/WwXdpZk5jnGoNpMkVboLgzzyNOdGRzkCHaTA5cx46h2pSdj/CE21IABHaBI9mFoSd2
Y13nI8shOd50Wkr801xRTthrtTeETPCkvQ+FxDv9fBIHDF/qcnfMXi++YKae3lIyK7Z5+FkQgzo0
7VFyFJei0QSMlrbvckzW3lukuB4JWhvAycpA2qeZc+V0yHCRv7gsp+aoPETJpwgloN9QNrGsihsS
uHxr3dio6NRfqLJgWFU0q1CQ+LHK22j6eEdmsknZDbvoddGrtfpBbIW0nB/H1uYhGBJ7Xq6KoU0G
KHXL7Y49lsngCbfjx+hMVsNipOCevAInR8ZOY2vYh/vKvfR+e3YAF9zhAhQAnj2i2jR67hKvmRkL
Rx5gwehMrWo1yXvhwRI+VQZovMIKj+JBD1uZaKEJX3ggGoGEm/lq2TInhEMwSrsfdyaJEAj6Rlks
+lh/S7rJPKCZBnjuwD6MrNkIM/nRATGjl1QpbH3s2UIF81B4/3Sv7Sg9nWhh2ppksqmrDi1rZk4J
UH3jXy3YU0U4Un2V6BzfFTflo1jE4fp+n6M7sVH3BYg2GjrN6su3IL462O/diEsH5qJa7fMW+Mpd
jrf5kSIJ95JZNp6ZLWlSKu/qfzfsF1EUCL6eUwKyze7bIc06eHj/HikB8PHxJ5irRnbbmIIoh1LD
gZJKy5z92ly7qCyNHSbIhbUZUelvLN8Meirf5A+vsTzG6Ryro26mxXusMuDZ8EbLvVYPdc9QPLXC
cYPG3VkvWls65RZW1lswClmF47CmkKyFxQvB59vZFNSRTw59VNdaXVGBb/6IITS9Y+GoVZognz+A
RMtHty+4lkOcA/gXtYi9VWfAUZjGi5jDDpGxnHjjGzAYS4zHKoWJY+e9lwnK79SgfLsqcLOkKKgV
JpLOcQMPRT5sb9hFUI6+Db6uxvesK+LEYB5rGeYjo2CCYadYYD+IshKk5sskyMP338C9pXYTtEyo
722cP0oOVWjJoQvUQxYA0YHvHF18MCgfh4BMU1Ui88mNwHwLGVhayb+xSqDkom24UblCiYIbGrNm
8nQvAt4ZvqkY39mM1dO7h3uWKZ1Kcy60YeTD6aEmJgRRn4rm9x1Z9SMZs7aCMuHHMJszsd6W/4FR
+GbY7Iw64sIA6vjDN7+Wp0jIoMp1vTNgDLVR54hFH3+2xXhfQaLODr0ZagD3q24eGyfadrFur4Fz
4mHHE/ddNgMDoFfVwa1QfoU3t6DTfY9yFkgCW4GxD+sK4Noflug1jH8sG47NS9CuvqdYaAgZqmIA
iCRyss05x7I42IS7IkMxczihi95y1Y9VnCOvM+0WZBIhYYsj3vr1WwOi62SCnXzgR4WF1+a6sKCj
m2OfxZ1WYRfSCmk6V0QrrdNwEc8bcFRfBk5KOs/sA5CEMVYV/PGf0KZrL2dLjmWwjRcQebdDaoZg
Wac8fZuxdGFVeapG2z/zZQvV4s2sjteESLC7xorzwBaqVqOY22iUjUsZvZHMtFONxIX2xC/pOuIb
9P3Lfik03eKjThTVSTRhOiPdRmo/NqfnCcBJkGPbJy0BzmSkp/5v15fLtjTL++ZcAplaUGa3LB52
EYkvDjXVczu0LEIsXrfyGbgrqsAQATu566LYWhkszwnFvVW0HUz+iowZm+mY7ydOxvMYORlf8q4W
FeUnCTS5ZB7b2YgCJFSxX+mElcekQLc78pQEydyFPyiE7mZrTChtBqtNPmqWX+TM1TcyMKdRHNm6
msCKMj56D6mRIpIppEMotMmnIkjfKsBr/XEoMBkA+iBrRPz2In7/8cHkAOcUJiTJEKf7DZA3VA/r
XyHvuAEirTrNCofLCThcy69ynFVgXAal3Tk0xB1cAna18g6OBB6VG7NqzhweQdHHa5dY4spcGOFX
1+GErPoPZ0moKMavC63jPTAvgUHGOTOfqatFl6u0aJwhq2U0CCw8e6oIG/KEeOXFlUq8Q8Zq/xJj
PV039r4P6lBmUmxdRVKEHW4h6sPbtaTfs3aJNReFobq8/Fs3tJlixOH5BxFIPkhvZ9+7zO9WWFVX
ZvTA3Uccgk170LbM/WrDEWDr9UQ4nVG/Se1TcEWT4KavyStQfSfEp91QsnMcXgBNvMS6A5+WiUkR
OwICHUDH2k45MykeFdKjVgUsaCDDx0+mpFm8ABG8vkZodzBrx65kQsxerkSJrlOcgGevUY6d9TH0
5BDWd7y+rrBZveOt+5VfnPX4OPUU/XDe0Vd2TajR9ahQEhGbLMCWLiqzKMFd39m+b2U5xGmYBrgf
DTGAvzG5V/Ug10bMq1R2rlwpEW3JPdUiF1CYGLjkV7q89KyovbTJMaMTTR679Y+T/MuMNYg/LNrn
R+3IsdUiuGeTuGIQbertR8wK0s+WCVNkBnXUEBCdCMaU461WGyGSDU8JfC0qLHKsV11EH9Ny6+eO
YelxO/cEUqyJD3eXwg3fqJw3Fn4J9VFYK+8tMFgek/+9f9Pr1aSAlciJX3c5mjGRWMZuo5x2TXze
6Q+cilzwowJXXtZ79E8ZgUMRRMqvAD78Nev8zFJoDY2mZCZ5jJVBYzUGSG3kblPu76LDVqgDFFXw
Ey7IQUASQpKbt6hsJpTV7e22Z2phoYhZDWd29RcIRRDLlJufjv2RnBYX0eqh2xWEY9WsgKp0R0Ro
qULvyMSit/DYzRVL9nc55Iy60QRKhC4ifRGad/yFnNMxzcmnHDot6+aVZQD1QSTqEkaCawz1rEJH
MlTusjpR4TtLPu8AGbd9SB2t8mVwoQumesYaaTwPohzASex2mGPIUEyFHYA4QTS2lJFgmpIUihX+
btOe946UDFQcEWa11W6PiIl3+zoHuMM2XBUuHOC+gxSz84l/pkyruhWFG9hWWgFAYkZ/BnKS/kPF
SNTLYFbuznGC0D8dRMoqiDkXWAEVU4tDGUJx8AzhUq5Vfb6qxeH3pNDV2nJtxiKyyvcXaUxdhn4r
r4Kpunbi5yV3k24ya4jWbPdJxYald4u+3AuiFqUzskVUPL4zwqMascV+GCFl7FxmLYfIQYGGcQk7
px6642wp+3ulXxSaKh+KhmxER0hl4WNuWFC5yY6I+R/swA3cF0EP0yNT7i1a01RJHDUjiy/zMG4P
6ri8bVqN/jIzWVBuV+4EG3bUPUpoGGk7b47g9KVMcetqsAPONT+XT1UC/4VjsmSVlXnT/IK6rRwt
D+NWxC9v0Pztrol89+B3A5iMUzN33UI4vDdOwdLZmsdQ9r5k4dMT4BwdDNs6FPhpnE+Ft7ob6R+s
h94x1H4fXqSHZhPQtj6E+F4E0/q11uiQmez1aAIZic2Uhr9RImxdhj91T6V9sGLZqWoLGRg45LRq
mREXw3rBTWJzx+H/FiJYMhF9uKIME9uPST8SjWbztvex0MvXSQK6e3LMw6x09a0dTy6Wr2Zvoysi
sn+ADRA1uiKKLjIPWF6rhLKeIG98rrTLxQZB2tXMeEZpFh1b3Wse5KFovXco/AyxCTOHjoXaEsXN
baD+A5P72KHssdkgYtHAWJjhAOE9+8wljTFW8K+wT2tJFw6FnXHDa29URzcKjtCJ4CaXY3c4xiI5
1wqfEp6Jyq+C7gQTHjOxTcDuhli7O/YWe2hdYLlLG67IYVltNFhz/M/PG6NTs7NkaExghCqhGg5X
QcQrvGPZSpAeAE6yjihVCWjw11XLPhB0tc8OMhyTjWHn4wDl49+PBOZUzUmp1uSkGmGzRchFsV9K
OtFLtJ7YIO6a6AuWQVDlXt8+UB5DY3d/J7+o9M+dWfouy0LOFK9UAXkk/TppgW6to+rvLFCquHio
OgbvcI3GB5T5/0Cf3zfx0c8rb9iqFxaJn19+rkGEb55UktJjMOvmvTDq7DrrAQqro0oRolBjMXdI
3hew6oRJtIp1BCBwvStFBekY7Vm92NR+UhLknYVCOZoH3ayvqftbeF/SnYniaAUaD/C4fkj4LKdm
mNX/1OtZKbhoxRYPEZ3I1CqldhX9S6esB+58bLFAGBr/HWalIy3BHhT8+qcY5JoQ8DaNrpInWjfv
2pm/NWshexWEmmU2lOGXgIRzUIrUJ4GD5RebWOYQy/OoIwNKbwqC90V2Lb480s5Rg8+QIdJPlr4E
ykaudTXhTU02nd9uhN1N1lydCJgSr9AJi2yt+8sLyZ66adO0zbi2bRJxw9Geqb5Ka2B1Fchgxu8l
kHuP6w+Y3AEeruom5xOJSwEwt9fk3ZETQu3YqvPA3ApXhOzlholbo7PJ+XkfNyt8C+GWv3bHFWAh
aBTurQ4w6VbpCanSgsaL41qd4XlF77+Qvt3pPpnW/3M4u+XcUu84PLf3j4sb/0i3wMbMH32V6cvK
4BSySNCne1eR43XBvTSSzdiFHIZH2H1ydXs+lXvNCVKoJOcnEz1lhVGuOU1j2JFTB/ynbEgRJ7lt
GOt3EoyAPmvlIiSBFEHRfN643AcNTB8QjA4Qr5Qb6rU+oaQNTcqHH0cDcWuwuFtUu0rSmKQw/nyb
FB4b/BFOOFkFb9lxFRD/Gb+mWR32phvZDjN2O5KW5DOXr+SKl3Rvj/9NLgXXEcw91qUoOtoMsGN1
DIw3AYxVMrnWGwcXorguzXJ8O9I+NGg8OdUVjFgMWkLsky/OQQkGYtlXiwbsQpXLzHPLkNqW50cW
hBqt6VYIpO/Tj9UdWbP2NrK6RnJMKhWCJIkED5u2RrHRMRMxt5Hn0/CTxn5w5hcbN/xlYRIetCIR
Z86wCLx2/URrPygb3vq+1QEGnjZWkw1/WPRUx7WPl+TrpIqAzIbltjrDgic5wdXe3jEQpLoPtxZd
Fdj1Fc3yPx0Yq3niYrfzLMDNaBnXxTIXbYJgwXa8DArz7HcPysVCl/yq4UmSXjWUl/xMYP5LwDRR
5X1NJvCHfXXiX9rOtpH2ejk3ZYVFRgkZSAph62AgK0m/SC6c0qNE/jXaby8LkBpqdyVZVGuCVvhz
P3eb1PaXv1xScNL8BfcjfKqJURxSg4j7nX296Ggu49Fdo3dC1NkmTEw+tDjpx/5YcFK7GnuBFd8y
YEkVpX5bnPD0Vfj+NgEjMPZi+4+ThThRAaVYEPpx0L2xhul6UBEO6uCsJutJMh0rARFL9doScsWV
IGxdIHn/nVizQPVm2hm1TLC0RotjZ7iZ2HHUvipTCT0ScWXhYllO9NXdd8/m1m7GoStZnIwYAEJZ
naZLJoo60SjxFJ27tECycsuRNrKCy7Uu4giYbScMZup7n7qpCIjpGIJ48lhW7w5Oe1xxS4FH4rmr
a6mZjEUMAhdvy/A/4B333knE6Z5VgG6PgAlWrQCMAtjgGIK+CMljH8Vbv+Vv6Xjmp/jcqNIsihAd
KdYVbrbxLov9tLUO/GsBGNvL5qY0N04vWXQovl3iXYmmbIXN9JQF1P70faSEdapXevW9PnMfI7wq
pBMUTknCabYXqvkec46QKgjfC4gmWXXzG9MwwtwId2Gh2vUGgojy5VPXa0dwqkJlmFKGiGknURgb
o2XcsAFNUSReasvnvb+SWI4+9Uy5nCxmiWjm1F04yVOZjTs4Pt50pSl43I9b4N1m3t2IIkv+mjBJ
xIB4oAtSrcoMJEdpC7XTOQLbCRP6e+op+vbA6ktWcJYUd6dPyc9i8tQEFM4FxvnP/7c3aYwyvdSB
cZ3QTcWbgS+nWpu+9z7wXjtPz3H1gM/XVIAeRMnNG4XHM10VM2evXY/gyswj4FXT64ZbCtpCBJhT
bvl9sZ3MJDL5YF4DuxGDxGKLiXKZRNinWjnr9+Unws78XJFOshw59bNOmQZXX5C6HQhewFPYZGPY
ERKcmB5n6hRoUdogvvdhXkgyRswU9RZiZBZfnz3t1QZkuDFLWG1yRJzBnH3Q4w0hbPP7bIcVp68Q
PSB9pW2DBjsnswbNRhrNUlh2K66BI/kUV2EPGQNi4nEShOttFGBTiJb0Bct4kfsawU2xv1lXQqGw
ALTmbg63x3X92LobsUjLshGqcecj94qXe11OoLHQLLaQ0icbP/hPIkURXUB6mCy3jqZRSkyHdQiU
/2SRWNXCVK/vOZ0rO0APS8Pk9PmX6XukIVJ9mwsL6r3Wc9Dx4ThTRt0bkiRIzHXX7k2JokRzgU/O
aqq8EqxQK1JxO0KUi2wmEeOI/B4CHsysXMvsUpBjH1wkvk5vJamz4X4LTZASL+yJIBUdBHgfe2YE
7cJ43SaD5hoPOsGD8ONr4yiIU7iyumYumDj01jsCxQ0HXUI3Lwckn+RerAfhhjqhY1cpLwSEzGND
UDR8CLwEDjaWZ/s391RXeFLyC3jPBOduWXLJ7sXJI1EFsa54mfixMh0RKOIA3Ews8v6qv7e23/R/
k13VH42BIkNMWnCAtgY0vRBHacmDYaBhcY2GzZ/BMUYsqMeIjpzPa9qyf93dXnvXuMcKTLuZ+bCS
CxfB2KarW+CGt9FWtSIQrwTaa4dGe8RdR+dzx195XYVJNFozmNUAiedgZELW9Eb89fF20xb0N84K
T6Rp018OTwrSoDPZ6fUst4RK+/j5pfgemJYpQAC9MAbB/jYg2JUxTb0Hx4kVwrJxMTbrbsKqE/mK
nr8Y0QChw/5K2/u4EyxtDC1wnX4lYJ+axrzll//r1vPEAxRNGdOZHl7dGE+0AHRCOx6nPhufJCof
q3uIFcp8F1CBGItmKvjeS0gm+BRQJwV7uULybAz/QXsZ/DVHWJWIONBWxCA45V2ZP97Ba89zGVfh
zbSHE6bid9rpVjS0L0jrJb7daZAOQUS5TL4xN/Id0fE80r0/AiXjyCbEwKTDIuFgw7Bg5cfILVj6
iMmHc4kvvEX3/tLBzuOEoJamjVnoj6Q0Pzgp1+/dk6VARsv28LZhayCc/6EwcMagc1k6vOOo/HGi
IoRyZSy1VPG7OdetfHBIsjgJKiggP7oPpRVgHUQ2ew60JCvYLDZyQszWhaqEehf1mTkRHWPj5gMz
+N0SCYPzPBpPEujTJlKPOZDKa5aANBtLhfSy1fWOFduATvg6ezJUYaBQWNkN86CCbeqS/OUr/lMc
X+5vpnvvTmNtobiFrNAUFNW37PrB07yKq0OZcCTO8TfbS1pt0gtKjft09EUQlXk2y/qCC5Bp8+Df
0CWmKbluGdz/Bc1PK8ZEjRE9YHipf/fVxRVcA3kII3oSED/oPEajj3jSCtA+921BqpNLBpBmY/C+
vlCmdzPPyC4bfv8DQLg+cvOaGSccWUVN/qGUaKnynkBKkw+2BK+I1/7mFZ03ZbgzKegsl41ApAx/
XEnhF04Rfj3FosBbaB5FWSfjHUhUThlRsryUtrdXfpkgdnM4tSylO73Dm03cbWMmXrj/iVNDzoBR
5U941aT4CpL2s76HIc/J8lVvBnLeqZA2NiaYetfPlxCrQOybCyYtdDLz0lB5mmTIXehXHsNdjILc
VgutHCJEUXTbQt+K1tfk+QCVrl9WNeUcbOsvIPASVzLr9Mi1NqEAvlpfu1qW9GKLfnJBHvj1Cw65
hmK9gEzlx4mtmvKFPW4Xzr9Gl+8MxNakjcqJXJ0J8GOMIfz3chvvPDNW+9tDydxJP+aqXM2mhgrA
tWh4b5refzwJ6rFXp7oIB58Opduqx3aT+Vp+PxYYuaoFdWE7u9tv5EGV4A6QOF8H7gmEUtotQtE/
twR/0VK8UOP95slhDcihB8LeXYK/CDUHShuYzxXihm4roNlH7y/azQJhfCY1qnEoCn8rSVrkMK6G
76hdAvcueW2NhTkcLFVPrGI1mML7kzY0WVT19qFIQY0EZtkwVUM0lfWt71zNmsBTWryW4NURDpMh
9zwsoYhGWgNMdjAdEYs8Iv9YT1EnkKwzjWgF0fXytj5igax+jgQK8O0r4jhflkkcvzdaQU8CnrCg
jnwUuPp7zLprgAI3JBTsxd9JUjquh9xjxu73ZBSPEMUfVQB7JPZOo0FLAUE+x6rA3OlKbTV4nT6e
PXO/xYUC21PgpQ6NlJiFXI5jRZMmS9URUDJnhICF1VjYbYFz+b7mk/GmzL29WBE21Yh611e0qyZQ
1uvXboS7fEoIY70mV5HlVfYMIlKULnjoLyzk94bGd05KZcM06DShTcKWNkQD90TsPK3JgoLdLJow
V7GSwNK6GoRUi4FLZlJCOB7oJZRLoZWOX9GzrZdmYPJ8CGOUGUkqwgaGmipWMnkR2CTd5AHrASwA
9F9aWPBaD9yPx4s/1W9aRsvKtHS4UeC89ubxnSlL0vf4V5Oi4rInnvGy9SdGk7rupWRAxQ4X0VB0
P97Wqj3lI1ts9yFTeYfDLo0k5pAJoFjRxkNL9TC7x7KFlbn8qSIghwFvGzsYyDQ1Gt6obIxEc6Bf
KM8yQhN8Z0LT1fs6L7gPwaJb4ZLUMavitpjP6qvRVweeB8ptvHQTu6myG3xX7XEzxGewsRtNwAon
C/cmZ9jfZMENbKTfBOnkS23k+flCanXcgWcVdnNEBVO2WPSwP3WTRnMUkF8t/3mt9CAggFN2ZEig
0iyjnzhkx6sYabkqFDbdNtQNfuReVL7jP4eTYkAy+65Jb81bqK4vqizuiPnEQwcFg+cgtzkzzsvQ
gLK3WAh+ZFMeDXP3wUE/cd3r18rewtx6f+HwLjLo+i3lZxO6ycMf0QX/I8xU0Zxo9IwnLcBXBw1K
NENFaVtwMysvcGL4SrgPkq1xx5IKEC8lRH3H4440AHjoNJGjhsk4BBG1VMmPRyHkxZOkgUZtRacs
3KABqrmCp108MGQSzr8E5n5sP90v4QSfOBIkfxHaI1koNmY5my5aTvhhUg2ZLwf+2E3LGChxPlF7
xOPV+jGvEe1I9KupjL+nACaqz616ZQvmORgttA0r5vrNJvww58cWAn8LknmW5r8vMjRg2mX9KESR
QkKMCx1EceawHZiuaRkccrLXfeEGO/3yueJYN1654oCPompGa45XO96KiLPE62LI/HvuKm7AC+Q2
77RgwhzbYrhR4HqzfFsVw1eMorkG4yz+rmXoIq1keA/O1VJXjUeY4KTJf8yOEebqeD/GGA2IB6zJ
pJ1nGWl9HIduqfpJAMKD2EYDmDgZpe87d9S/STXWGT8fl/YkIXR1SQ5Ab68Q/pBNSHNmLhLdFO8i
ZRuZusu957hI+yCEPxWyGYbwo1dnQqOvUQX3c5kcNlbIt1O/isZeH9RhFwU/3cznfmOWv7kO3Mc+
39P/c5+G/LiSya17uIUgUo9NMyEJQRjVWBxyXHWCPMOdbTqtBqbci7F6dgI1ScP8RWjDI9hlxo9S
uHN2PDOwR5wcMxiY8xCYBz7sHvNR5FlYcnEIbOOOEaPgomjPgYcVWeCTwXvchQbyaZ2TMQOF1lRj
knd5oJw9B5dlSedml6r9QnOXfQ2mCzeDI+7j/5Vbk6b8QG7eNG5EeMf2pPDZPH21hSZMzUL3bI+O
aVnhHaX7yNfN3vJnj69hDuWcd4UHNHf+kf0oqAeDq7OD7YvYMpGKn05wUW5OQ17tCztjHy7gJrOk
I3jjxhiUFr2Jwh080gWS2qbp+proKr8N7LscCLMhd3HgYg3sgPmotZYxtgm8GVvSu1akQaRPDj3y
rvGtja6fTEc4xIvVwybHp3idv29PD1+KiHAgNAmjJMX7ZvXJbypDOQxZ0jiUoZdFAfJbXm7JR3J0
mxdNeN+MVvJKDWRy8ioTOi0Pi/nBAmoZeCJk58HQ3WaAyiHWKRHD91gGx/6jnSQkvchoGTPmsS0o
cZ98ot8YNgJyoalZ6q8KTD25oM7U3ORykTWZ6pyarWpuINWW+t/7iClm0Hcl8PAcOoyVfc/NVcR4
Nvt9JTycjZSZl0Tmx61DPzvqQbu3Bd11SPuGaIXz23bcLfrz44hQP/MSWwSK2w7YpzotJ9SeWEp4
V2DAYBsqZEpHwU4z0opup4n5xxegXCpXmzJE+5C/GaoJsAaNSNQ1OcW8DQnipjCXz4EhV2VmdbHV
VhwPlXLCzgorfWTkRtzcgYmDA8GEtjbY3vy06j33XFr2lO1ZJhj3fSx72SWmnbwQjius0qYy17MQ
daSr2vG0XE/FYpMy3nX/99KuId0kUzw77+JPqUVxNLsNXUi2z3G052+3R6tSuLPq0dFCnQGO9WOd
+jOD/pJyiKHqQjCiwhW6iHZ1gcMyjEOEbmKWvIEGWkI19g/nd2PEp94zdgHEgMS26+Y2YG/ZOkOA
0IKxiw78khw2jWmvAIvKqakp3QIBC6SPJU3UDpKaBdRZoHrszEiGAdN8HoCXRcwddYumBrMYrGgh
EwN+5i0uzo/AVo0I5at1+VgQXijtLKj7Q8AUuLiQMcCAmZd4+rFdhBzss0wJfB4PgqNpB7JTV7YV
exQXJNxvlHgfRbp7hyaMG1v4BQCbBtJmV/UIWwHYklsXblFpTFo67kl6wmAkoEilFQSMBq5tRp4W
z3O7vC2HHVNC1XppF0deVc2udz+rm0aZOESUUUYoz1EidrCt406v8jDcZEvMxV/kCh0fvjNI4/Et
QnJBinWc6ymJ5JIu3nxy6xGUwgtw4YABJkSFk5phGqJAcYuhoUqiA3NC0T8j6v6kWApFq76CBIDg
WNKBRp8CBEaNw7EqPNBpAP85tlcjDp3bFyM+Ql1iF9rDdXINIGCRm6RpWpf0hpWosuJscBDPVKbK
xrW0MVOsLRclwdtYGmVaWa+h0F41wof0UtOB9CUN2PbPQ/DpjirFmsAAA+eCO+8bGXSoqswwDzyE
QVcUT1KlYPvPCYf5QDqW3OlbL+9Bb2xF6O5vG0w+vI177zk1sgSPgUhHS4ajxLB0vQzYl9Uk9ga5
NygonjZHx2BPhv2Ao5Ou6QzOwji+V8L4EmT5g3FRLIBFx3rRLnx02igrX1tOcRRb4zUraC+YL9BZ
oT09B2Wn2AwnBqyRDY+W2Bizh/KZ8MVfoEeSuEFmVT+uPLVT5DjnVqU3TFiLFzCOcQc0ntxZ3pgY
ekoTSaRZQxKLULdoVnOc11Cs6rr8zv7lKQCmkjt4CgKB5+8aFtAFoBUo7CpAZwo8Nz8dkW8lh+wg
R9u/tV7xoEVv7TxREqK9eF4xEeIBesjOJQHDvj+ZqqpfCstuekM+xunw7CnrWrg5YrrHQh7YL10J
6CDL9J5T2lQC52HboExKGZaeD0oehgdlzaRo7fWB84M7YAZ9OwIy3PK+gqzEtOg4mq6TD5kjXV6A
riJSwHhDF18dA034kLiq8YPxUiD8la6adNyGrG1hGFoGrPZzPLXUockxtaWVgxN/2H9ZsDPo+TI/
k5fL8WFg25+Wk0QL+3dOySZwLPzqTCkb83asKfxDDklOvOGUSOW6Zk44taQ/OIe8wMKu8bqXyDru
T0A2fLziNSpe1qPhMknallKWoPBIE0EjNLjUYaaYOeOs9GkQTtuMlWiIjDFght4Xhl+BYHB4NSZq
mqN7R4cWDozG7DyhrxU2MMp+SBfjiC+Znvjjw/p/UiYh4kRabfZHdv6woqgkd9BaTifjA7LS0KWu
qyvU3EfWyarAhpiKZzbwrVnf7L/OmWKx4mQxSK0QaPO8DeY8Z/MBSmgVKcdN29S/B8wlQ9WMsEw4
6WIIvClo7oOYmy4ijNGi90v+CMUlq7rsMqTFDvYcPfbBhQ98a/7q6V2XIE7WM2Hcm+VnxOu2+lmg
HCLdOP2d57nL2FqGU8Iqs4m/Fq+IKctHT49YRpjRxNJMA7Xf7SI469lFG0OqVJIf23FRWt/iI8OH
ykQvg6/2iZ4Saz+uwe3WNeDv1JpnA43wbpp2s9nB89qVOLiKxGYpbjF/TVca+MsQ0QWW8RzFVCql
h5C9V64Zq4fBAqy2EgCxonVO5zFVWhYSM4cnBuEia0bBa2CUoYZR1udzbWruU4ZtHyhOFiFuuRM6
sdZ2h/bgtgRvyR6pLyul3S73cTmbarqipoI/iZssKLdQlOgCQEt95YAW0csLdNusJqDHfDJqCK56
rjaTm4s78Y5veoC3irOMbMDRd+jMKTptNPRvoChBDzdZgBep46S+wCGp9Sg+7yBeAWJYs475M0RH
O0OI04sVZSTQXCvv6XXLcfTQf8lRbkaLakWJsCvjA0nnpHKJpD7fPWFmQjCQ5Y92cWN99TJoEldI
LzANKPRz8YHznjgjMUjMLgNMXz+VLVwTColM7h9hE/jWhR0gY/lF6I2lN+j5QirrwIcPkxyTZmxS
gSCvF9KcI/a7BUNA6lO0L/Uuxokx9bXwzcyjOZAwJrWsUMGtUlWCfRKgKnmjjEOmS2laFbxtPxiC
DPW07WFRF8G5t9MZG8iSpUMvgaAHjl8fqKeWRUIhCrFYfbicbsyGqsTQeg0CtaXz/FxOpYPug3vm
82QipAxEBF6K6cvQm8UfOKj9McbfyygqTTSBakGHutBhIE4nz2gIeauBIEDk7aQ3THsRmbJuDOrY
qq3fWJQXdON6Nsol/mm/HPleMfiyO/94tHJfHWhTxE7sj+Itt7yh3tQd9fzS13aoGbzhzmnYNSwl
/KQ1VZK+N/dlWD4NiwfFH1iKrWVtCg+4pwHV5jh0L7DY4A5PfBCd6KNsjalfvOITyfHzSJ8ZEoyu
+tYIWOz1Mjx0KTzu5kNFhAkVD7z+su83wZKMWEKB+uuiGpw9YxC1GpGDEHbo+JMDpvPyY6hFzo0M
rbh6tyhMhY3/HsLAMfvtVYsxe8KHY/qk99PvUwCLxiVKYW364OyobdcdohossczjNV1O0vqZ5i5f
LAysdzujARPJJs6Ico6RV4Jk3bO6IA3zS+48uK4SW/yYKIVFyEiAYh6o0HNqtdA+iMXZVn0urZh8
YSM5Hw6JzFy3LNs6HK9KE829XzJiXKLDCyb0GNrDzPJJ5Tygd/uV2s8303UCu5kxfOCv0kV0mjz3
g8j3wYRTZ2J0s+D0/Pq6QiqBnXRzahMMzpnXR+rEvlc0YDIJaAp9cUtfPa+9+LgpB+PW/M4jTSWc
oYzl+p9TgdjYVVjMBZQx7yP2fcpXn8lHhSbuYUJ31vKmSh5rBEuNvBhonOh34n6x53xznQ5rZwAZ
RaiOe8AkLbWWChrUOaZYYjcYJ0TncRtRTJU4wq+M/dya2HVCTSVP6whFLPwVlu1ZxUnHnG+oI6eu
/mvIPKBxoFsEnWtqBObA/en8+tGGvkhUj4wBizZDGu5WcI783N5yaT6WMmnMZVxu8XZjkhWZyc2n
6Y0vL21sYByqUAM3bF5/2YEAoqJU5rr3SKSPy9UZC7++xUrQbCIk4NhFI1Xh8JJa011gCIzvDngL
tO+GVIe+1Lc2Inw+2VslKZGlic8QU1NlnDwtcGIyWbl2bvQiwBmoWfLkdjQMPaymeePweajTkXy0
35ovrizNtR//YnuE4L9p7xMzufoeRWtm15QdiYIcTQzl8rLHi0RF7Og6AtQJeu3cLPwXzgdgabz6
sPnUSF8oZNIOzOGVa6Zq5Ls2Cg8W/dnYc3ICbXAw+MYkCAA0u7sWYhpWXMU3dUMQTursmBbeQZRZ
BrpwIGPD/Ao7cHsoT8N2cIldEbpgWZHkpiNbKi4Pl2sXT1crDP/1oCDPRPFQ5Gt1hTfVTyDrwKMb
S8/DymmlRTIF+JVHt+LmLGxKjJjAvHQOJ+RjiGl0rYAE0jDEtKWJgtRIHA70w0wyAAOoLCjb/5mH
EoIHGyzF3dTVszWgT2tqDG6YWqf7BsT2qcEpHvKxnyyAanVqoGYHlfrO40fHOK70ic3mL29PSeNd
GLB04iomVMjahBEyMJdg0Dv2DpDmfEfTKOQ1VU4a+PIaJnWRNsseLU3j0jI21xv6QV8xuzFuBKVt
xBWbRdBqD8JLoYkbxgd1IGMyYI0FwWXmmtmzFHvjNchktHz3vFLr0mDXxRSb89mF91U3fwwBW8Mb
FR0Ig8Hx9CTfQl2Rxm8zBFVg+QWzQl+LaaXYoAFhpipGNUMceQYqFTok1LJ7N7HAr+hrIkBCpOwr
DyDrJmRjpDCOvif7BHzcEMsQ9QgQz0c0s4GUArmPT31tlV4JarWvkgd+XjqgMZ+mTnM7rbm0WPgr
TNU72srSDmSD5N2pEK+Q7CBXOXcxI744kB09FMg7Jggi3aMJtAfqUa4rPw7b6PmWf0VTWJPZTOuj
/+1NCTPB8imz9SHKGlsgHye+HqBMublkf6Si67lzqw5gkrnsrI4BRFWcNs2ocr1ZJIIWu9Uw0L/f
GU9lsT6SyxqY/BQ9lNPOADJDGRDRJSJ2jJQoxc1Xte+T3wqEcfyk6LCuu8o+hN6E/D/qpOr5Zrjx
/r56bS5mO8Qg93VKVALWD0how8MkJYW4NgTcNTLNO1/LzdY4JgLkqetRTE95gFMi/ZLeiM38pOkT
LkDH7TqGJASEdyASTFqow0zcsxWvLcak5A8iCPEkagrLUxHRK5UBHXOOZIWTV/mBwm3p/zeCpjab
5iQJESaIjlaHgrESLF3/x2AJSrbgNj4SP1rhBxMii69t9LuR++qET47C3mLqls0frOJcp2uv9JQG
Qdg87EF1vtrQMw3e9Miiohmbmy3yXK4mZD1VQv7jlOp3X1qduCJmUfbB1wH42VpQkpWU+FrF/V/u
NJSsV/ig3Mm16N+ZQzap19LwT1kSoNvX664B82vlTtAP7oUAqL6I9ElddF2B1SGIb8N9c5vIps1L
ei43U6+QD/6nBao/v2Zh1imOiOVwwRgCWfScFa++Hos0RUmvxQQGDbZO41T7NVLkgGuJ//kSUFL1
KFToDJaGp2uYgPPlbX51AwcD8seOSwKbWBdI62vtuhPJRGtF7FH9CJ6Lltb87GjArAIBPAJ+Dt6k
lhD3KB62NOUzL65nTVQt6h0pF7Fp0vn0RqMTT5mfg/KxsDSSvN3HWoYNYZUh5DkRQoPv5iO5t2Kg
n6Q0F7GJbBjiJJ1yjb4/nNfMKwHHwhHZh+KzLQ1P9PqZf2V5RVJBJ4xCld1nSvXyMDvKaoSzzc1j
0QgSl6HYE6s+EAFHJyIMQquirya7g+8QERLnnCTEoX1Ru19Sj602yyar20ejWmcCB61knLvVh3Uk
PGIuK5aJZwg4uauaLZsoAPTo5Yg2tmMmaz+QnWQAnDkbVGIkmddOwRfNM21Gsop6ko6m736bj6iT
P0O34x8K/7B+1bBOhFl5m5UsvSUfN8tNhbLaUsG2sbegP3u8BJQwm4e/25oU/+cjlTtGIGZ4F/wB
l54b5NWXZ0UQbJpCOH0Hh6h6dja6n4ALnzimO0+KAz0puoyXPRkg8pUfBNQIVE/vN98+3UOFzpJE
adxXmMiDwtlgoctROV2moZJ7nEKs9F4jj+ZN3y61FBAA19E83pqnErFDGeshr7zXeMg89r+KV5kr
IAR555SAwHIxha9njwKs9L+MshkH5hAhnqf3ylb4aida8LHlduBosIpPyM25LtAw1xhhZu+Dw3T1
EKdgGonLJGKUTU65iWbMSxA3JMPXBXFZ83bMDvm/t6rR9Q5ht/Z+lya09T8sLXb/oDmN7MgnX2qk
39Ywqzxp4fUivjEln511GsjNqhJp0FwMRsDPsjqwwt4uifng0ASQ2tBrza6ktPHTuJmP86F3sRmt
QSDWs0M+ID7yKI81okVXLuGdSWpPsf0ednFwGrB3qdxOoYxto/AYqXYiSj+26fCA0ZGoF+MWtCsU
rcWVai/BWHruptToYGEkf2mb45C0AucxHhToF8fPsyBU2Jhepipu2ef2kacPF7WK6eR2oqB+FNfU
PkZFDc6bSpr8K+SiGZoz8RUMLhpJCa2vIoOjs3fkO/4vBah6HPqiNjmeMlTNsUB5SY6KpGgb5K3f
v0Gt+8lf2oUGkjEZpE4H9gelugtLIIv+KvsfVTlZSi9r7GSx+GiBLyvIiWlpjCc9uSyibTMMTwr9
UpDKvPCrHFI/7prNhVicmI5DD54PgEXIUfPCEgwYGXRN8+IPwBrihdQq41m+V68mPnB5Nw/Tu+lJ
fNYbIyD98Qwmswu5Riu6Y3DUqqDsslkkflCrI4OXi5UIrOxtCUtTyxPJSC9FoCWa0ZFGXcQDIEDQ
KxFBYXRIo3qKKm1JD1hdWU7HCrLM1OEf+NxSj6uAEf2f3lw0i3Xb3AKuMMm9nEZic8gJKDaxUUKs
QO3sfW6lJxLkjb94XukZ8HNzI7lxUjJ3T5RLezk5kzXzJojmVkuJJup+YneWmcDkK1V6H5dNpxp8
mRI6S1QSV73sBJRysKE0lyBzVe033NPk3v5Jk70k0wECUEASopSbm6Fr9E8m1qW3V8fk7eHE5eRe
/43cO2piyRBijpX72BDPSrRpUa8TKvZgyhg24gQNFJHjyWiTIM1iON3TXlfnOzb2hzs5sVrBWReu
PMIcFjMRCOvz8r15SkTDFTNflJXjSMXGinRf8OpDSoYW4En18w3IDLKS2pTk6Vzjows5ZtNF/s8G
vDnDGtxeiqSmZT7OnJRacaRII1lOwhIqPd17BAH3TEUN8Zfsr5tTmK1oppZyoBxc2C+J36R3xPdU
QlbwtBAWUMBQdpst5QBFYOpGgwKSWw2qZTKXCS8DGPBYzKfnh+0gLUx6ZKGdAvbPu9Ep9jf62o8O
k7vfNbOXC9VneBTdfju1+zkDTic3x5UO/dpk+/nBwhTIE2rXc0s3jcu6BDmdiTnaObOycLgBt9Zr
vAtS9JHwB47fYccyGnsxUgU6RugSs4dXKlFLSRbxZr6odJHRiknJ5HAFYTZl/FenlgLh9VJgFPvS
tKQYAFl8ofomYpj7m9tCMDR0gDOFWx3Gfhk0T73gddgBF/YBsToorvvzY/b+clk3ZxjYmhCd7jSP
Fllrw/Uqr8ZzlP59Sz4lpXXXv54TBxCQj1Hgshs+PhUDlduu2nm+rT+HJ4zaQZYE83tZP/POgPNq
ICx66sV/y5lKIFSF+vojI9nznvN7BJVLlJIP6WMMshY7n7b4C1IoZfWpvcLlbxzoXDMRndG+YMPj
wsQxPILbXKQNTr2Vn8gSvc8OJBWbcLKqgp9eyydfe4S8hZWdKsSvB2dmA9GfYPeDxP71y0YW9EN3
ZkNqlpTJnRyBjBJY+czFNRvvOSxm67DT+6SiNEI8eZ8jveTc+slTL8FJIfpbkh142hvuY7J7O2UO
QVb/cO4TbEFrirh7G8io60UKcTD92teQImxzKletYdmeCT5YYheW3XxegtX3fsqTJBuV+jKgv/gS
ms7QC73BVynjc1cMegcW2qP2ACiPPyj0wqnuEKr/FXTbg8Giw3Jh/3qQVBvHjkrQhqX+pp+UPsbJ
lTbwgewhQRjK/O5ITeR/WPTnG/XzgxydPEO/BQ/GdkdHcsmjjMAn+uyyWWi8dEwUECaGAmxyEyt5
Z8w4DRsxi889y12eLGThmmxvnoAG0Xq9l9wT1Lz8hAhWGX4iWSqCSqheapZkU7DO3I91KI9zY1Kg
340RnE+kCs9YlLVZeEHzGH/Q+LSKcXS0EAkP9YJz78M4abDlJIji6jokqAGFJ48IXsVlBtR6CDrK
9GdSIyqAbmPCFcQZ9CRpXxFt5ON8iyzLbqhNFq18Uvo8Td7DdHU7pAs7rbLjWpB/EcapQc6VLF2K
WG+d+10FbypeF+DxkqLJbUg3K+PwfL3/nBrmQ45v9gDPhXbt6MAcdhCkNmtP2CILzvtU3fswmqw4
C7DqrkwEmxQMtxxMGYkuPBlNAo6y8+ILsCWp5o3DZweJqy1msauugrLF3i2rsUZFCWZ19QHEL6jk
4DV9NRluqUD9wYiqbCCH0dJfNFWKve7hRt72gjytdRXdJ3S/Qh7qJQJXn10qV+N977ctXcOyOBfK
4Nkw7WAT+nUZwVeyWYt+bCZx1Av4oVQaKp0rpq/8uQC8nfzcaXTvvyL0JWfk4d63BFjvdQyoC/cJ
Rw4fAOuLcvBW86IAfy4cyvi+8l6PiZUXCAJYheP+QAlrn7VY1OYDmdtKkNLSu2ODsYJsvITkxY/0
l9f+NIYKnWLhZdyN39wjDo0HrkVkh4QL0n5IvtyThHCfK/UxNQbBt1NDB8FqTqRNOO2aI+LuHxY3
wE9nJcdPsw9NT5PHNE4DYVS2HOunAooO+oKaLfTsY597cOKeo7aAWUx2R9qDMYfklbiF0slL2W7y
v7T1Iy/Ysbs09c446rUTbAbdjkmMQRePY+Qtx9Cgr7IHwpvQBcDlmc1XxS/NHdYWzGd8SDbStopZ
57FdVmGDup+FCIZMO27+lOAizE1TdjSzhE/JVDUAznjrQaaLpKADqraAkrQGf8RWDm6istqqJMR1
1aSPfR6K23bKw5n9QGi13xnM2oBvI33InxfuXqb6sgzvylKSRIKnVf5vZJAAXw4DVG/2UQY30GYa
60droZUSKPNimOvHgcCqaQBdIZuYQ8LJjdmdg+CjGt+DMoAhYBJ+EYYobpnTOC+X70zlVQg8JwzS
+OWg3b6DYw0wUOVauk3NkGhpdF/KOuCZ8tE/HXW33/1H3SUa7Sj0NwtiiPw3I8iSCl937Xebq5nj
otmhx/LOTtUU4o8JKxMFbxvOFKn2u76tYT3pZUV1a3nTL4TBEqUhxa/+eGBoePBnU1uKEZhXjkUf
eDT22HM4oNY1mOxENH411nPy7WDZ2uYjU1GFyPU1P7AkizVBUiiwbWMNEO6W/QxECeN1BomjsY2T
Z5VvT9gwt445vNcBha2JcCdB1mN3HFSK5Qc5JEv8ep+FJ9XLlQ4SmbmUy4zQee3jWP+hh9JfvjdT
e2xiEdc+HVAAWzh9uoDtvxDD8h3vm1kiinbmGwm/RIrordMAcKnueGdCswMFGLs3/+1YneQIn7U0
d1A+rqupseQfLy8StQsp6rfxlqLZ0jo+JfQ13iqg+wGLNX3yk9xGrTqj734EQdVX84mpt0LTDUH5
am+LHNuAhnoYxAPpI864oaKmFITL99viJuC7/HlW0jwG7If6pOgYZxGT5iffa3pHmop+JCjxH4DO
7Kf1TqX34EQXg58mmfTZyZqiCzwFAyjm+01RoQfRUxoTOdUdvquNu/PLxguMKle3hSWSvM2HNVwa
KOAyP8lQuQ95iL66lDEo0TCUDhM/AZExGdeFBU88sD72IGexiWO/3GaIc2I2c1cxz1Pq9QXoC2Eb
PvphfNgRL6vygNszPjBOyw1f2reX06AHltgPbm9wiyI4lKSiGSXQ0dZRkuCSwqrReyWnbXtvyjMj
GhxTHPSppq4nS5Q/4q/cREoWsKtzPdIlr3hjOewLo6bJSQH96fF7kn4B3sIZoGqwIpnWs7eqIMcV
dO9g/RS2NI2sNA9Fn4creRwN/ov0vjZd+lb73HaKsJrz6lPwUhv/QdS4/EmLbrpHtCijqvlLQ0js
gX77G3rHBlW0jnbg7+BN7alCNnNA1ZmwWPGU6eynF2xP4wbFYGGYnMDgicds57p3eZGbUmkn2i1B
UbqcWtNQBOkS6grjRwGugInTnBuhIGyggDwr3FV6qt5mdKaa7IpWoex9O+WTTMhAYOB9t4x0xEHu
p8cenVuNOw98IIoVfIE3SzjBDnE4YSs6dwQyAOBan8o1Mk2etJWp2gQZzfB65x8zprlpKK1RJVNp
uPh/7babwQiA7zTcfFkxmw9Ngj+8LnMEWX1kLpbzg4RuUZGnhmstdR+oFETvypqYWedX+NZt328U
ARFjLD1enbVHWRAxhAe1NJYcgjECnQWle1mY8jT6qRUJggKPZmZlX1kK5WRdqP2rE9hfIWnzILy5
y7LJ3S+dKYbAsvIzjo0aRt3FUJMM0P5WzrD5qfdXpXDjy7mCZLHulEp0gy5gjiAs7R+k7zTHGFY+
HK617O1ut/AxFvf0gMRu3a9J89ye0Fj/Gb618YtUFFgghen9GrBWL285dKuVFZggrHaTMWm1sVd5
sNxmZuJOAZgVz7QAtJhLl98EqaL9sMg5asgAPGAw0gR18d83cGMjbogD8j1oFdMPfLtjmPasajwU
IwCN4TOVuYBI6zLjdkEITRfdEoc3XWxvE/DnDVf9bpvScX69Q7KtwOYkyzBGFfBEX3KMYrsM8ay5
A7JaqWtO5kA9zgSM96aVv1L6sR1TL5MdCVxxXVoV8M67VNgydmi9nt2P+hrc2w5WQe0UZsCJBNH8
q9dMu1MrH320ukRx0GLQr4bXM4cssq8q6dfH8pSXpaJbw31PRlwxU+zewys9BeBunxcFI0DiQMHL
EvIOxuGPz+6Mk/g/4Vj2zSGh6aCNjzR6e2UJeqEHtbHd7fIqulowFE6TkLEGpmhFC9RkpYtBVxee
CCe9smgi30mB6/+K65bk00TOLUUBF/QjuCMK5Swllq27rhdopiWq8vDKBWYqeHWSjurs78k+oCT0
rEwbTjwMpkhmha33wEzBWk0MXbq3qrT4lc2p6fATm3P0fJUh+SBu2rPfEAfK2p606a09jmz/Z1n/
7TkPPLKJShexs459AwWFT1pGxQAR8Aj+P/+dZyKBUC8FY6a/v4uhxWk5XpNq3NGEZBvDxuOj0fmY
R3PqLf/Pl5DlrgGPKvIdajCUno4peyWC4sl4GYcpaz5GtKudD09c3VmOrhs7zzvGiDeuaqnCfh7d
P7LQ2HY8+60ywSUyooKcakiS5pZh/Q5c0uOn0lU5P0KLTH9wuN0h3EeWXXPJjpHBoiGrPD7Tpifl
jW2JvUqO53cCI7w5UeKkmLkKdT2DYa7Tg6uQlLy8wi1Vj2zeNlug/BNALLEcQrNxdstOAn98ECc4
Fc9D8NUqJte9btvk/QmElbLd6Fqr2wFnvpKhzOHKpxeHGnNbiyMsTc+AEVLnEvs9qHoxGszukiTD
0A/BsJtJWY6aOq+2M3IvNyELyyZtW0VVEk7Lsn9LmPkoASagQZUdKJiUwXQ5knZ9lHQLt4y5bOlm
S09zwNyq84Annmx75B1STrXYqBBMjCrbmO2ygvI04kDdwve0aGJuw9CGoKtH8DbviGFikczNElVV
aATlAQkAiRdHlP9p/xtv3AEAfu/1dZHvic4gEDMOoOgTCf+G+7B4I/Jmkbt0mIwizlNpw/RWH/ue
6YE7PsVud6nU1iyAXfqmM6WWjmJfFlUXmOw3QJpsZ/qD000/uB3FppWuCxbHwhqFgUbwEGnO8oRG
cv0PVe2TD4uMgTd1lusxy9M44CHKZrdAlxxrlS0XaSFIeGYUloFdXKBD5cFLwplqdYHI4IAh1eKL
8nX66ITDJxMpQU3r4IvjkL1neMiXFq8Ohj0g4BDhISS73tco1+fjOCgbec6r7EPFrGne4yTui4dr
yGNFbn+IUcW/XjdFa4X1iD0sjEsTXMcQwiJLKU5bowFK4zd3kvznoPpgm1J0ngT4d86UIWRWRRAX
2ipTz7SUMWxI7OksmXRAzzAnwlFL8TLExmJmAtrEKvRngI3RaI6z4Y3UYBTeevJPg6/riVzbt3H4
BtTX2h2yTQg3Nwbg3hPv9duIHiIi8k4iUl2MLQYCzsZcq/6sTltS+Ow+HfxVSYAz0x/HVMb/oZKN
XqzZxHpGW3xd4MgVbPmJJ+d99EytLHE65a5BIMykCj5LQVEZFVtxfN8NYOP1p6qUWbwQa7pGMx8g
Gh6EpzOJQm6YYZi5MsLuKtLl/taxNdzO37/JHBb+jkUuqycnUmYDBEo///nhPdnzSJyeYtNQf77u
JcXkiosF4WBRwiLch1cjKP8vJjX1vOTORjSrdmXtbMU5Vi6gWiULYZAvjpPIFEWTdrEfHRa1drzJ
CT296YD2L0iTaY9EeWIOTRkbhPeSaHGLMffBfMaWwaxUJpYu+632kjOFRMn7YqGFr2zqVMQ6xpQN
/PlAoeu3c2IDmVAQPqJeynJqn2hfieQIIhBOV+GQsdXxZfDnQGkEf0b4lkYyBaVgae18Wg8Ro/h6
rBqbjrhXSoQFOjrTTztIv8zxKOw1x1iLY+oDG3uBG6uRUPwgsqvTwvmqegBK6DkjiC9DpUtN1PlF
hfGeHPludb/Zx9lkiUQfJl4TicKFqwXHsfaIx6b2ZR5+yOmX0mvo9+bXTZJVHGWdniiKrIg0qcLi
vGQC+oBeVYsGsbqXoBVSBl64bfV7hzIOjpHroddVZsKkDeAmmyb78GcK4ILL8DG+sDiYnzY1OLRE
L8OzWt53IYZsoqJmputUfMznyH7nXGt77QJ4rWSBBKkQlKUa/+GVMgl/PPKlhw8nV1KJTDQMwgaA
nXgEPoZGpDEUpQeDL+kW0tMCM7NznkdgMv/5ot4uI1PwfF3R1vTgzrkJYHQ+KdRfpIMq1cd7wbZm
VgdfW0kq+7ihoqoNh0PpmXWWFKxXt4RcHhlwU0oiCfWnSrHwwCUByAQ8stJ21PRvwVX56cboTXFt
U5mB/Xpz0y7vBeKM4bnPtuzH9QuT39LHjBqUfNTY/vrTYD3oU9lycvhWXmNZ60XrQJhtPzyV/Uhd
cyXiF1ZeMwhevjpT12o+OTKyddKcRhOVMq9qQbCe32rVX3BHJ4czxthrmdVL5r8bCo1ODka6TX5q
GONZx4D+V3we5CvAfqgEC7jOX3wbzOvgNaVhzaO58eh50Kb41kppjb6HhZkmq3qDd1aB0GudxeKZ
8JHfZpajJongzHlK6WG7uPk6Iey4eTTrC8DpvHgAzMyr8cZt172xzc6NbSDgrjV5CDV6TKlUAeOu
hpaTgb0+5qSdwAt/20kADaca4ElZiXseQXWeGZrEf9+jrTh4LqEJuEwWL5lC/6SrzUqrno0PHkWN
lkd+TtZK/RWSbGM5UKt7RLmMsQKYhrd4HZpgRFYtO2V940ENfS9NAYHcKMl+UDTpANii1rbhGlvD
+SqeIJB//Lxspcu4PJXiMj+EmYt28Jo/Rd+r5fdZjWS/lctGYiWW8QvMtPL8+kNHLe3sW9IxwM1i
3K9Cakydx07gZxU1mYy3j1l4CsbvAMOvotvN50Am9vMgZtbWsc0R5yO6EfA490QPC07J0xdxGQ47
jij1Dj8u3q5OQAnyQ7iLiyM3W/QJbuYJygvLiKdL2kGQ8DyKZko6zA6sY0GIM8hWPVwso8ZMlFwL
C2UrsslIebsQNyWr/QbXCWGuYxJxdWK9bo+gMtRVHgsyyQnI5qPC/8nWqWGBiT9ebyBsIDiKPDVm
dSZN7/Q3T8n0tiDFwhZhkx7HemYwFB+gv+sePK1ZOsfq4fV6zuvJ9mMJE+gidmePGchGYJTypNPv
tncagWs2OItGv6/8KEVT6bi3UP8qhw4cmZCB2JlEqYleKEu7ByC4Cf8BBpb+UWy69tCMZp65yOra
eecvUHUDJUbKghrA3M2GbC52P03PHHuA463kc16j42h6sCWqd4/Ta/r6ld01CzIt7DqT4eVUpOux
tbK/e6gkIw9z18iuTgDlReEo7OZOapjjczCfmbSU+5VBNbCVB8P5tbgf7lH7Zuqa84ffcJ3RxobR
vY43HuMgilFjv1L3WxsvP8h2xeSOHrIW2KFpTjDvM+PkCLoqKgyyeL3qLue/bXHHsEpft2JTulpa
kKyKSCX61hi7K5qavXJDDohaVWmE3+wQrkkmcKl6iq1HyJ3aRx6IdaSNioyG9DgyHMQhsMI4dcdt
c/MDlgU47pkXERRbmwPsDvVR9ZwNbIcpER56uA06TCQhVnYEHxO2t4iYA1svkhDWySwlqzm8vvwt
HDxIwc3E6iC+aUSYuagmaTKQSPlnB1TSODy9UUkVtRTJ6wf2AOfGHeCRnTlSsLVfkQtifhvsbKuw
CjHrxO31ILxubZolX406aGgvhNAIXsE5FuHqdjCqmUUwSIbpPX4s/3XZFH4roYCa780aL4N95IJG
fTRv9aXkXYUPGm58pOSmVLfOTVX+tYUuMDMunCKO14nydaolKCD8B1Z+yjuKKaJIQxtaxZ9zmytv
egyCG8VswM4srcN3JZcoxxiNuE37QLIcxUhEv3T4pXIhQ/SqMsf9LLA52mxPvTCCd02bNTLrnuwp
xhrXwhr9aNEDD8Zhuy5TfdC8qypafxedfVyjP8+JRGxk1PNzImEM6UQiRFQtoP8dUkrOi+DWDzIH
MXyt+jG2IQCm0dYIgEOebuBlKQXomFqPl5l5hXr0VDr+B3DK/IpILO46V5Vzm4WCqrq0BDfoKp9/
wRWNfqQpmVhuhprJliw4kVcH4iv2ZzjXQA/OQ76upmNVU58hzw7BhRGw6nfGgak1spT1+JQ+4+82
bTtC7wLfIEob/MnFR3G+DxnCfS0dk6INY/Q9745UTzp7yjSpw+P1CTVL8uXxISLmVm5O40mmDX7y
kLilzZVz5RCy7jlWHI4hJKPVVU1dkkg+EkVvcBsJoGt47SP0f9DPP1leD4O48m2ULj+FONH1X0Sb
Pr34uZL4LlZby6ACyEk/VsiBbcVYd+AVwxxtihu0G6FKD2KZFhkXHW9I5fvEr/1rItBdaGHR+HTM
sBfodHSOBi+Fzq6GZoeXlRdgjCJTmS9/3egHl683Yk1jUtjRPn9dbC7cBB6wGlA0wfcVW/4bpk8T
CUx/IIe+hH5fiI2leDCwagBFToF19UutS3BTpG/NsMTfZqj5rba+CUFaAIVmovi0vzZmEOY7RQis
u4xrfsT09qElCHp9roQWKK+M9L199Ayme0g9qoLSne2PJrycKNRiRrD819z5GRfdt3TybRWen+IE
N2eRBQV8pBjLtNNzLksHNw4x3P1hNC9s4l/gveAvLNg8YBPxRD4bk1lYvAk3cJcPBoUF2QLw6Qhr
Zm/XNlOFmCLfttZBoaHvMiI4bCAZp4/I/TPxGFFEU5ll5+obYGoKfmbTPsHnvyTE171yxLIVUeNY
VFrhd2fi4AEJvNSnv+//UCmEsFGGTmqM5TbqdXOZl7oDOh413mX7bENnV88MUPDmLJPSRDMAZJlT
MxmKSZIjagxVfWc6FXVb3SvhOmXZTxFuTY05q8c36xKHrsqjBfEJ1I4ep+sz9bEI8QN7LSHNBLV0
VxSPuJCGsdA8/YwkOJiB0Xmn/0Cvw7m35c/wTstI7Yb3meyCQM0ghVu3dugsATv5bD++8Jd+v0m+
HYwMsVIuqSDoTeuBU3JouG+XWhMacZ3ym7dZYg6rJKSkYjiHk6oABwzN8ZFvEOqLW24yfIQNXPeF
rh3LlMhFGuma9byior2p5zA3x2NdEwycwqNH7IiRje9V6j+hYskEcYlxZNlyZToPFwCbbltQar04
9GufYrsFsTx5j4MlOztFp5W75Cfucd2JLik+HNo+RFTDX2wR6u1fQVtixEO4k/RRX+ED8pJ1Ouod
LMWxiGvBZ2PNCG52qLPiwf3e5Rp/GdpBuNhAZLTQnU9LhN29DntKGL0cB0L9a5IOsthqjt8v++kg
ukkRV7vkzFQDGLJAhurp/uL5H5pvJEUtzD3lvnj5sqb3bnNONBWB3UFGYEhNhj/VyEWuOtn7xXXy
wHJg6+X/jxPOQKZMfhvODJbYkMDgBVxeO2LY7wWLeHuSCp7QcHSyUf2x3r7cs+nMKRfKNCHlSh7s
LJLy4rYnsdZFrnzJuV3XzhP9txmDdBpTEYCXy4ASGEOEQjBrxY8vnNI8naRJpLOQH3ft7wmejSSZ
s9G3RdNbB+b7nTitLNcIKx6ouJ4NlFybShcYRrdRRxDAnKklpeMjrJFOiqk3B0ByJghr+zYxbmFs
AmpYf6yXsHakViMYzrDWG8QR2hZ0eanbuwuSOtwQ38RAMwDkcMIlkTshrGFq/gBN9/XGUV5HZlVA
+IEV548q+tFLZBfuKSS/xmVxfJKpXK3J788Ca291FEBZNdFIty3VUBKI+ZOmODubF2B0yfe6Evo6
fTv9+gQ5BVv2srk7lPHd5ijcJshD3Ox9uPyqz1X4Sa3geIg6iTRuB0vQShSKQ9O4aI8PR3Ndbxgz
Mx0gym1rwsNUDpu6SQ0ungcxoJzmEOyQgBAc8t39jLmY7+PE8+WFWwVgTCIH6TGVwzUf4fNw9b0i
uCfV5mfoW1RiGINfGwh5d5qRNBBwx3h7odmhAtYdTex9STnjZQLSoFG1YKSom3vsEE/7y9FkeQlu
e7OkMgBa6xSqTt5T8Ll0xWbJGnNlmBQw0ENLWt7K4S+DQYlCRkqQADVy0Erz0EyJptKTpoTuVNw5
ZaHgC1dr0Yw0mqSCmIodK4018rqApn7F3kvtmhDbv3ZqaLyOH0G9pYr4dnq1IJzpJg4Cvu10u+l/
dscnpMHD61Uzc7rimorPSkKZTa5imYnV6e+pnk7j1/5OAbAytsZY9cPLWuHLpM7Wv9Z0zJ0Ieq2l
y0yrEL/GKuBzcauy9Xilva6iMBLOSoOlO4IQSN4VbZQ5vMbAUO6RLSUJ8ZbAfaJM4lrrpnWozqU8
ppC1X2VGGUZrIskxsserYC3i1mZJ9nAIKGUMWELqFKeNyI5WazvYM+w0fVNmhrmlSkDZC2Osb1RQ
t7wEEszQXOuE/uHnkEh3m0PVIoEwSaxTdSwTybdEnFSS3UPCkrqwxCtkBUANusgHTgbIzqYPtj20
4OcGUa5mt7qC3KrhGrX6h0QVlGYoDMJoOFFzlmF1/nEi/iy682h7OabKZQt69np5aT5bXULeoRF4
IE63p7rLaU8Yv0OSUnuZF4BGrpJXBG4Z+yhKU3tV4BAeTXaNYMJS9GX2z44JVsDr/sg3ys3K9Ypd
0OtQ9I+iH+jQ3dmRBAmxybbSa2rM+YDVyK7lupNumoXnar7HGwcyc281M9Ya0RZc7fZDo7Y0CLyo
bouKO9edhA/0LeIhgASoaZvMWTGzxzSbgclJgOmgiU0M0nnAoItZEX9EooU6X5A2OrENXDNHAsgF
ljJFNiQGspmlKwNbILbPOJPE957wH5po/7T4O6tGK2kWggRKvXsmDPUdJrm7cU/CUBxDvQqz+ipA
bIB/OMMj982ne3ADfvLqJD8k4F+TxPylm4qolu8BcSsht5C4v2YmpM2Q2huA+AafiF6u/DEjxnGB
mC7qyGyDLgWiPfeJ2JXrnauctZSpbuA7TdwUlqGoBAHIEpbWchKU2vRDH9msJSOi/7YrVKbrIO+r
+Y1AnLOWPpm2QY3J/CJ1gqGWComkk5g9CCZDL+4o53jT71YdqGYHAkBDsqJ8s0MCYk8Eom5re5XJ
uf4hTketdUJE0TedLbNuhY3gBfuJhwnhYeh/nIu5TJvAO1gUIFBtMSRdlzefMGohTqkgdE+a7Wmp
dfaqBIC5B5J+b8Erp1DNJ5lUcHcYAIfDNRSS3jghCWhSKo4LkJT8RXOaNAzPWKou888nlt8sIcME
gUcQCugnvOkt8+NMJJxk8og4NRVRB//hqgaRzml3Pj+UXvdokBrsqaWsMFIuhVsRm7Ai7X6vFP/l
SDu7LEjfkeBhjdl7GSG62delc+MPkegFqGSWxSk5KZSMm/oW88cbbOtlLJUeurbW9uIp05yguhfl
AplenThnPrK7j5YjWX3IvFNdxNuBbBYM1mEyMzcqD4FDvhLZHaNvpvC/vSy8+Fws32frwEov4uIx
O1Mi/NSdJF6RjGs0PFw3utBbdJk6nqYIF2UH9AhluwdnK5/40VQ0gnwR/GIDKFK4suG4CGV3Ojzc
t6Bv1PiP1KpWxYAKXzdy3b2n2BRsR5r15A4VBjaY50Cbww+QtLuM2aZ2OcTYbfe1T9MvdBy2fOkH
Sjp9lczYVDCJYmW0QEQ4woQ9kgDMFl9HOI8/uBMWVbiPulvl9SHs5xU6Jyy4t+GdBWxJQMXTECjX
OSmylMkzoMcHS0+cSn5v3S1NhfrGm1R2C4CtJ1EssZUqD0HIwobovBkOEN29qal7p1hKu64PjWxN
sFBu7omH7+RzR6VN/T1TICvlvzPNwlth805b9Qq+DaE6QqgCU1igvSrO70f/Sj/MsH33DnXF2ECX
AqSAfXd78bU7oAWKcwUoPl1Wf70wTduya54r8eWcO7wEAt0mlOOqBngrazRSp589S39FZ+ATlVrB
Y2AERTBEjkEJdlZalW4MVA09NpvR1TSLgdBxLthnKsTZI0NcOK7O4YTo8ETl4lISTnFA35J1kVa2
d4iL/Uxq5QuucDOIHtEj+a1aWxCm7BykAtWQ5ouKdQcE7L//XLPT4Bixg3lrwv9RBFq+L1FLKYhm
qIrrP5e+tG7aunicDAPNYov4z+k98IIu5t3jC6VWX49utnQF/m4gJkY4ansf2ZVC9ZVr2rZqWtrL
r7yF9QwvLKUbivcL90JJnknUAWY+mi6XWsrUxA2ez/ECt33xtgHRdpAv8Qq0gEYMciYYrVlUvz/d
TLads05W8Uv9mcpyZcCGCoBpG7OpuDppkdqXNBPhPO4Pqlc5GhJmihMQ/ycYuPKfkxI79FQYqjuN
PI0xN6kQG1XLrbLC6OxgDn6XNpMzZXVhH3ovtGG4RobsahxlRQQ7CX4dmXQOeBWMHb97YRFghZYB
CrKSzzbr0j/xH7bT+SyjJvNxsaqsOWt/AiJcO729IgAa9YklVDd+xmr2czt07lo3jme2T3q7pSRk
nL82jsfBupLYyBLgYNLFpIB9t38yizXBZzS0ov6W3gWF+EhECn+E9tLej4mSsxsGmxC4I4CgNmgb
TpKNN/Zbv7w5JQJsBJD9IxPWj6xRRts3zNJaKJ4OqY4kqWenTIFnvEA4hRRYT7dwglMotXkZNPUY
vzAs1Fc6X/Uu9eSIaiDa/WIqBVrki4+DRsnwf+ZEQdoehWZuTRF12bhPYA5Od33XzuBLcd0VCSOQ
puZm5C8YbfAf/lJdOTEd9iHysp8qX9WSGW+0WzI8i9d6LcpJX5I3gSRbSPVLOIMYfCCiM4rAwrgc
1TwnsSbw361OXbccpTO7DAbyWNTbpnjE+OsccSYgctHEXLxm3jdszH+QcCAkp7+Jmkeqx1PGPCyH
aiyClWNLHYqUhIcnZooXWYF/ATV1vgpxvudwutRHXhIXrnfaaHSau36Q7UsmYQlQEI3TJ5OgR4OF
Fe+VkFEEyPgJN5dvcMP+f81aUjI7kERxKEMpewodWrovWKzc+rbpnJ1Q1zpYRupA1ZyU8VMQy3Do
kDK/ACK4R1736CPR1+vs/IUp7fUuMrq3tbDwGnSJLPcOeb7ofrIGcVjx4M/J3aqka4NenqD1DbxA
WRjtmOqTf7c8VTXZJid93gCzWFIggBabjmXqZj5eZ8YZg65co0I9bQX5nKpbDBvMSpKz1a7vBXlR
pmg1SmbcIxloczuFjcyvk4sNm/qHr4GP+8VioKcG9iHg1rpnwqDn6RXjJGhHCzlD7uFO0CLf+m1h
uPWge2k0NqJeSAqzJUkIG2RVElarSgsQad1EBzlSplj07b7lAYjqMcezuSFUKyerprNfEC4WIP+E
JiAWvInHKqGmKDtX6xnYDE39XkzBmPlgke4FyJ29NIPOPb2a3fLE9j0S1pX5RwwmkYpdOkrDlD8M
JKp+890lcuu4p8luoJLp7/hRUhqGbv9VdlXwUUoodM8Q7pC9wiGvUvvmrcGP9M8dA5WP3yTfadnf
ySqgOKLMMWFhcA2j+/BU0hmqV/oUAQwRVl6JhO2wn/BWuXGpaTed4yXYTTow9f4NKFt1uv+EYM+c
APGNP7GzHbJ8NuvNfsz5APQsOxkrVdW1N3YmLR7Bo+uTGRLEnoYv9ginqjV1y2Tk1dVjZ1ROsmvN
IXC0DuHTn920m5bd767KTiLdthjKrW7xaJ4E/LLu9GpYcqQyGbaiSN/42dVfyyVPn6W9Dpep0ktm
Ls6T3dM0jEE2klmiElKDqG2vnrdqylvoVqDaDOWRnwpV1wtTsimHxmTol5DxgCBv4JL/fD9+t449
uvBvRE55xf+lpFzXWGLpIfCsU+ItbIM42jc3Pf4uvJco41SoPzvAs8AVWLHPsg3QAwCe7hTUHrEd
9eCo4j+DBgW2f4KjCRYsfj3FXqbTqr75UCTUqJqsNON3fL7SpAh4LWJ48hfvNJNozX/VqyM053qq
4mHhHrNsKTzFkaxRm1d27D7GGAbrH/e5W+zRw35KanJwreWMv6yE7hKuJykJFeaFjjhmLBVJqPe5
QVnr8NX572pcd5a3GCgfVqD8UYGfPnaXCg56Re7icXok0obNiIaeJVno+6S5CpNfKRDR6bLJQJQt
0UtbeY8DBghPxHWglLI0zWGFtTqaR5rVd5Ii4moJ0HZDafxI80YDFXBMk91B/GgU/gf9J71KrnmE
MA9as2zVch/Zdbbd2Jr8k77K5hBg8+kbq1Ir0b4soIeBrQ+k+Ts1QX4kKL77czykyv6el8Tf2pZq
3a0cX415rXN8q5S/2K7t+USH/8r7428UNqQOvH7jafRCcE0H87iCyUh0nP768JWz4+JBpf+DPv4e
NcmPZkRuJWLvo7MZbnJJSxPK7f7SCXbcqGhQlWwrgnnnf0D9uUmNKpUE68n1EkY594YmLeZr69J8
OcA+yXavsXfAfdc4AReJquLUp/QkXwxBmAc58IPdBcXg7SbN26s6cinMDau1g/tJNz3snuShdoSG
PKqMltifBIJT3vCgqrUEapJk0cBl4jaKYPoVnVbmJmNJATePjBZSDG/TJ2NOHFTEOqnacxOYveaa
Mb9wEMAoWKaEmdQSzGxDgBSW8lBVXt25MCwZuNhpbEovvpmlOGlEBVfUqjabrDThRyldtK4Q6n28
l2r1U5B8XuWwdnwXkOmSGG5739gxOpDUyQdzvlp9g6ghERl6o+157vQ5oEAQ7iutGtpInADORd1k
trditdll0Q2nBFoIk4eVjgeW1j/YG/RZuW3wzZj6RLHWmGJHIgPCk39u7HQjrpJJhUZIY8adDTHK
qUUvN/GXqQais3w0P40cZlt1myla3tP5wqq7qUK0aE0OC8V0VGG7g06+J3MrMXHqhjOfXSVskNYc
gx1FRje+tiEagIBlXXLhsJn9YEsU8zsKxiQRC/i2osd+ONYUkNRbTOnsDNI8/rBuGqzsCpxdmVsg
kDzLJgSziW+Vemd6cfAb94/sINUkxVmRekLxbQ42hD0xn7QlAC0FHoJOqGcSY1hxkdKLwQB9d08d
W5B4h9HdbqnegFRbB/X+7Y6UGDEJlyIHERXaDizU9cxc2gggNuu0WeE52fhKtDXtMfOGCOvthOiI
dFEja4k4nCagEYFeZCFssfiBUpjo52eOT5XrLRE0r16RoWLbAe6jVurQYbA96shZoHWEPZmRfidb
fOSUY3j1R+bXWSNbQoqCr7DKb6yrVLXReLoar9j6RqNcaOMnZ4FhwtD0jqtOKuRMmU/86aG1EKCq
0xTSiBoALJxgjXFX6pSGOMn/vhM0f/O26Y3avsfaZ+sEkI5J0Bs6xIktqibiSE3WhqM75gZZdhKS
IEfMq+X8/2sGkiAODav2Bxwqa0VU/bGX7Ji0NCE3XkXqO4ZpeevtNQcbCtPRmSGTYPxFhmSOjxeB
DdlVhpvwglHimXOdpHtnzpHg0T0DAH/LAFYlC/Lz841rhyFdNqujdDhCQWKqZR6QjEQPCDefkbwi
xhzxO1JP7BsmWX1qmhB+khpPGONP0skkx4i5WEpOv0w5IgLA/+/nm7rq7rLxLYhHs4P0iXXozWvx
pq7kVxfbk5weEz8bHtDhsM0J0Uw71XZHcH+7/+Me5JkU7MHsAC5BQcVfPa5O+C5mu97jtf6I9tOz
3YANe8Jy7S1AAlgXKVgX+I52xlFwnQTVXu/1eBgF/8NXY906sIKof2cZMVoTslrO9qPYcySc1Yms
zKpt422nayX/u+E+U3ur+o+6Nk9Mq/bVQbyO9xEe0XX+yrQIMp5A5plqJSz8zScRsGskBv5rNcYb
dggfZPGKY49yd+DNQ1BP2HiiOnll5QF6P6MnWX80VcC7mtQLs2A/h8j1irb/5FkdWbIJQEpyuiwB
WNCNEyYhZe3nMS8fSdDHz47d9xe1QgQoIyPxoybeCqgaRzmU8gTxaqhZrPTLbPCnrTsq5uDVqvN9
OVd7pXzBef8S9fhVGTGzkAPk8QT6ytd0D5qbukWQDBK2+ZTR5K02QRTP02zRA6DdJ6mNxuKOlMVi
mwwOTH2D2WeYOeDu6SzI4EJrN3lIYndL7GKlvOuVg7zXVgxrmil3MP4ONXnnf5c/WSa0a4HlAp32
/Mo2w8d3vya8RlVgYuo/pv3UQbaLJROw52etzrHtmhs+4YGUnJ1wjscA1SgPX6dUpet7mxhNgxWx
2PMR4l08KnY274edHYzCCslXnDD03/IBpL+KyVvzQZtp/PxeUzXpCoLcqfu8j6KmGKEBv9iJatlK
zx7Z/exxAaYf8IclPcwkzXp/XxqiPTuPxCZuDqAtCydFb8gUw3zv5hmXrLUQBO07a/vMOd+05Kpt
OyhrEQBc0rTNmq3WmnlY7TeLK+n91KMKYKf9TiJmHEGxTHRuZzmfdZRzL+AgSjp+79LWDHVbw9El
/fn7RuwDNw/WdeL2UDleiWYv6bMVIOowzPIUSggB6f4oXO8SVQTqlS0rpKNCAJJ/Zn7hE6I29uLP
F6AfIqqMv2K9GZN/O3kKjEGnxMpXZJJAEH/fPW/aqaVNBTYdvMANpEFR8OjunTdeMlrmn2RtxD2B
N6ncb+Z8ItqyFe3l44iS1EcZGIxOsYkLxks7afTxyK1MK5m8ipMWmImRiQ4b+5MJOF9cRz1FbtKy
Xrbs1+VS5AKV4/+eJmeyKIi9ypYzbRcKAeFw/MkImfu5EvtXv9nMA6Bid2YANGeYRzUrWSt1093Z
XZzRFkhxT5SQd8NnfvUgJjQHQXI2QZ1k1lTwbmCgAJnXXHwSMAiJVWD0oPQS4onWQMBcCjlyVhvx
Spm9L4gXZ7J4IlqWWSirnZZqjbBKp4hP2KeZiKuKkE3YSGCqSigGRBwN7aQVBPxsEG/umFPOILXF
CHanXMg8GgLitIC1yhBkYxs4Pn2W3H25HCLJY++oiORwQT5ObdoiTf8J0E021hBb69MeQrXzzzm3
QqzkedwwWOXllJGIu3ffM1O6XcbRkYHAxMf/Od2BFZL+iH5B8ZcGEfyszGr59iB0OR4/L6bS0Yov
HSkhIjw6G4Yqq9Rkz1hyHL6Q2eBm5Zpv08jtVTKq+5woEpscQIs+d2XrrHY+XS+iPRRI9uype2sm
OSPQMwu00jdjgzJ7Pz1+l1TZTBw3W8J5Ocgz3cI+JjsZTxuLp6svVid/BTzP64KqkdFCqqYKPAkZ
LY/KjrByWTKEAv6w/sxQQsWUXZnNIMoFwB02C3sCpqHxdNED+Z6zZPRYvSp//KZJmGRtVLAxVqKt
Wc/mfGC8XHu03F8Pz8ECxHtRCG5JbxLuJDWSz0PCPzDvjil9DhOrDQ2rqHRIZJb8IjG1IjR+QpEJ
JsNoGvnhPx+5FUz4JLVS3dZEOHPnWXELcukW5kvoptHfC03sV+hZVwFXRPZHQLzHnTWixQp+2kPb
gHMyBxx9cyzuk9OatfKuAEtLEd0fEqv0s7/WEw9Mt+Vlpo5exiDJ5aa6mp58jPYZK1333mEIZWlQ
Dre1EYn4ocReFmbSynjR7ksB+tDKZ04uM9fW/TNvtOmYqvmISUI40P31Udja50MMWQee6oHnGUTX
9ReaqmFKy+bOuvuv9Mx52zFsd2MEFGheCQVydVFMglDTRMy4vb168jKeSsQbEUhrwM4H3Dwkjw7+
gTQCp52uOTuyxSuFTLFSKeLlxfPclphT9TixisgIMJCVc1YCgaOqrnu1IGy+w6iUU1ovCBFdq7hx
DmdEIx72TeIOhgtwpR/AUa9ua5vJGoJ/7Ht3OCmFSy8tKxBmUzjV6+i3tggdcgBf5wbZCu5zBpl1
dXHS8o7TS2EAUYauOUm+0+ndNxw1Qle0a5QlA4sD/Nix8ck8pNDa8byCwcOospq/x+hfTmOhBz3H
PGhCg895mGwGHyn2eUPElYgMZDs64HcfF3wcbE0780kVdTqevRKzrk+pJx6+gtC4InUiAhe0hXXY
DGIkO2tT+AT0iLg7mq7U/JOJE7y35AfzHkWgv3m7yz0NZIkUXT/+HRsr4Q+2JXT4r73isHY19OkT
QJIjGLs2TXQeyvE+m6oBu5t84VbrISIEZQgoB1pUuwsw45onsulcKUZ5CEBnKZGqdc0QW5zrsmAm
R0Je4IZA4Xm02j+Gl4GKYG9X27ikC9lEA8e/qRp53FeD5oSuWdc3cAtFUkExh0S+aTcSvLMhTTeL
nltmfofAjYdz50K6UJiadxhA6yXoNKMS8xUF0AN+xLo8HqToYbVrIccThOMqAceRDo+RiMZd5X16
5Xt2/f5bcYMjZNTch97tNMOV2deQ1l/iFrFP4sobj6fFRejs+euYbU2oxRsrUskl26zZFgn06Oge
wGiGM8KDkzoz7O1zupmxM5kTkbeZsQPoUg3F+p8HrW58SSEE+Kfpx9b0H2grybJbUgjJZRqmczXr
Pc9zAIFHbvdXokaN2SmirmAo3nd+LmjZczcUeX8Q53bzSqxMByMNPzmw6xkkOIXBMyVkt1IwJhnm
gCftIKXhkm/gBqqnPHopBE5iE/rVm6O9878mNerrRLVUoXAvGH6LdaJWTQ97oJr4D6VhCOiSO5RK
Nk609VrvO1rtInkNNWncQ2MKXoDnjjbWv4cuuxh51hj/FT/AYLjvsMs2S7CPC2KWsaRJhdmjcwV9
wAUnnhU/lKEv+DdfJ/gJm3S5K/OjcF0pRYTdU60z663FMYlGvtY/qZtrp5A0Wwa3KYf1D/hO1sRm
15JMumCQYhsYqSxLGYB5mOYp+jl0MXLeIHHKErMW+jggSByp/XWfD+LeLWF/REpTkvlnS/dVw+P/
GwuEnGiZbR7yadYzLaVIzxMkBy6hGAlwaDbCfuuBsNyuvzPaN/0uXb7cdwxBlfcZDymRhpFMT9fs
+M0EXNRFp7COVd/dr2MSS4aWCtNHyhsy5MQYJqHqBvWUrqMSzFQe0XvLwAGTchjrBDyBdQWPC+DS
mjZk7rKw+fLWQuIiCYwR4YiQJ/fvo8JtTt1KTScwjO/leQId5R/5tEXTipZ2yf5sLP5IJes4JfYV
g88McffAiFgfMr7A0HUM84hazthLRynUpT5mNSDfOMzUeMv2czDik5XcjqN4m0RLH2MPVmE+SVGT
5hy4VMJuG3FHUsKUJCGHD1XSKaZ8Kk9uuUSA5V0Eo9nwlffRKE6mgms16H9+2BoSlDmhOPWMlei2
MPRh0RGufxstId8edACj89QJA5WKlmO9QuRQid97dBPnw3b5fWT4yy3GJJ1H7vg3aUUENLtYqVs2
FsrfX3oNLXmjtWccXD2qbE0FAjs+nwNk+jAf1hOzZYb9qsW/R9tA8iASxkSY38j0JnxfYFrDSp+w
mdEypGPTKCFhJiRykn0onB5EIjKJ+2jhBxBnOApdTqGkz+wnoUNycZCK2GchCrvwf9grQtCwoU+q
09IGK5xz3DQehETRDzwT7j5k+LVfPN9aIa7npadUj71HFWf7Li3H8LWMQScUn5Ob2gEX25Q9w6F5
Zdrbdcffy3HA5OoNGknFZbEIYjbt28ZuUWg1VlF9SJ8jSQtbNUOvwggVZmylR0AxJt6WTMV1zRyR
82+4n6WqMSDh/ZZ/yqFjZzlzFSnK05S6kdotF9zbfBv02ZYW/tI1mS9CFutUeItX0GXZWDpsTdrL
VxM9thdHHm6GN7NYcDPoKB7BhhfDQWPGbD0WMMof7a9nGTAMDYbeH0xRTmFagXAcd4FJgTl1YPnz
oRbR78F//FUwApcGl3soZiEgG50rONVdZy8I2k6cUGJ7Hvs1se4NfVHnBBZayB5yCR9usCX+60xK
SbWcpgPwXsHKOB09/HdGluypDKYiRquMS6d+d0U8uKNDuEEdNs6qtNFfHqIzxVrcCPw91dAraE2F
8ylsEDBbz/iykoOuXP03SGW3wV+mnxqgC8OtA4g/OvSR03FCZvAI2Mn0qUb8H7nhx2BwrgkUMYKX
HmqGb+mAHPba6l2denKSkl6p2r0fzG40H8LkqpM4zu3VZHxCzojYowPqaKTYQbyRUMPVnO8asJmf
fc50H7tKDEChsoindboeS+Yw1VeiZBqD68xG+FGJrFKpmt3TWmVFQrPMNLLOfqGS1sxY6mepdj3v
Oe8RvZFbs31J9BGo+l1z3BBnnVRNyhGKJYxNFgEdTBTOX9/hHkNHc6zQRCFql0GV0Od/8LYhsb8w
ra5VyQXVZy/uvjXGtu5S4ByfJ4SdfxSW/KCkeWR4iKvy7fBhxGzrq+cKw491nIwM15uQF9bisloJ
DyGDrszn8AclZ2gakR/B6RaJvkN4vtAUplHAGEaaTKlmXUk4pijPvyLdXNBfLKSTce8UHvmrDm/n
ZYf9Isp4y1uL/rUe+lz52YVd3tziv4JtHTz/qYA+1lUTFyvAf4P94AAjUiGwGY2uWhc9IaZN5SaC
/Q7xWfeo7+zgW1ZFsl1zetYNlRlbs41+Sb9YULmRzusz63pmLSjMseoHZ8ZHlp0mYzCcDSaIxMbN
DmlAKjs5iOJ0AN/hTMw8QDwks3rv4ahD/L0mNpwfARjveyRRoQ7hvyH/gTQ209xkDBNd92I81u1b
4KC4AJIgZBBTfzP+hpz1rasz84lxrsBVfKbxj7NiCnn++hLUFPnotSuYPNBgU5kznq889lVLx+P2
1exB6UirNt62I+rD5OXaF5vXnusKppn2V+sRGTM0b2FEDn0bmfuCAec5f2FhbJh1ImoN90oxw3ms
3SoMaplUQm22yRPmFb4/UR5Q9BvKh534QagTecCaPgev7W3Mtb5N0jbMX6pV373RtfOvsvmmbyO2
EPa8Mbxg5HfPzlOkezVd2hWF7q5rYgUVOnq0hFLfd9btSE+sBYvRmhrgdz7J393fxPkt/0AgljcR
+YFhiQIshoH7k3vuiREcTtbfccW6RCKCtExtGMTUSdTIOJdKGJ2cxPvhAv2CTVybPts5dyLG3lvA
rxN2Kdfq0wZqCvB2FSY/8dVcBWvWEaAwfaCrnWHUAsiqaDlUIgdLXE+BtZm98aqcqXBnHFVih43M
ctJaaikgkqiIqLkU8QlKBXFudkHIJA2u864KeRW7DAtHRMQQ6LW2bRrVZKMT9mdayfyBHVZ3d2+L
jT6XuJRWR23/6jjTsmH05KMubMJaowVCN1WL+iSjp5r0LFSdDh0+rkUDjdy/uA3vXPJYhrjY9Zmt
rJMlqI3w9HGQbWwm9xowvTLvpuvL6xOW28NDLpw4sfOA1cJDYqqzQEM9PgykZ2tBGH3hNwzxgsAg
SrLDfl0j5DOkP8aen4McCJg1yVMdoZEDC9E7OtZAtJFF0VsPnZhWPpqY6dAL9CABkYZw70C2FVhq
D5lwkdLisbxAtZDD4t9zj9SRKIOkphimYCtx4MuXl4a/RtqR+HxjinCks1PLRW8YqKYqCMcPbXDM
bIfH3FY6jiwqI8trFbFnxj6ExzoFheugxqneulbAKW0tJVOB2amZKQwrYa8o9tzGKBFVbaEUGvF9
wDW/ix+7CEH6wPmDm8YsS5QOmiYqdflDnVEihDMbHDTSV4k10/cqZ2cjJtjcurhzDBCj8pR+73x4
VwHV+vMA4gqTo/vSz+FOAH9FPfAO7BBl/2O7ab2zZX6R6I0n8V02id8vfAJQkK2W9u1Ou5rWsvm1
t1m9H3H7Ons3n6ojg23IWh39rqPgHz6WctJ6C8jW+NFx5MDqC8Ozqm8j0h2PaQrKGdxvgN7Se0h3
PWEPw54xn7vjXFTW1tR5AE9Q3h8wnvm3y7J/gtSGABkC28QzT0NNAV2w/2BVuxIUuAE8rmP4rUoI
JPcijqwB1i7vMttn4jqnPzQ+y8HvPZvx4RZ1sDvbzoZbG2enXPFLTIGnZvB59I3xPkFjxASKYq0K
e/ZtWeTpcua48oJZc/lQeVrjd28jRfieDUCaq/Baocl96TeyeNbVdOAQ27fv6JMg3KNeq5VCwLdL
gu81M6KU01/qJLXcBOEEIImnJkbYz+9dp4K+60A8gCENIZdTk1HW6j6fxM5olL3I+uaYGK4GU/ud
q4oDJCNUhEgfYBtykdEBdlAsHZsU4Rc1tpgqqaxQ0Qp8JMF/5Ub7EU+c3kWXgxNHKe1NFBal89ln
DiLNT+YwWWRmX+vANDtQ1gJUDVyQC79ZI3GYCIJPGWNuhDCFlQPGZzX1/Sz0AhdLLixSLFHsvoIx
7y88/Xk9PfFZoIFJhF40Gu+qQOS9i9FoOG8VPXOZQyKemFp3yyezV8b54BsumQwrA1Wy7Bcl6SEA
SKFjJp8fZ3XsC6p+1P7WLy0WQSmbFwp8g6z28KanTfKSB6wbcnP3bwB9+SL0iK80oPieCZvq65mn
W3WEYd/Iv7wMQNGWZy84iX7ZvLAJbxwdFS1VlPgfPOCgM3P5YdhFIc1dLPR4Z1MfFhmMIWRHnBoi
VqAcf/edYnV5f7Vt40IPSIqDJQkwqJtcJVA7725GYFn92yXMyPNnuAR+WzF1WigK8hKn7KU/X8GD
d1Z3q8KrxxljdtFtmqxL/QHAckcEFEWCTqC91MWig7KqWcruaVQMV1m5C1dt95LYKznT0tdd/gvk
hkr48FNlFHYN2U37jKBASI16nTiCw+UQi8EkkmwCsy0WcCJo2XwhYk30Nh2opPsHXXjn18yFRZBO
UysiGel0dkZBMGDkI1/99Ri7W9C/GoW23mt1LsfrQ2mY3EcF05B2cVYNZw2JfaSTyNROS/uRaZh1
GPrBRY6tpe/yaC0JuStWergBIQ8Tj3jkDDWi6xC55pDPanGkE/Zh0f0NrxKYGnEfK5TBE3waAoWS
jkjH+CzvueR2iChNCxQ/anobz9RqPPPg2VKKSQwFupTC47vB0dAnqy7krlgXQ9UPzZiJMrtKigVp
Pmhxq0RvZeUg2qVoAzTov/0Dv3gkQvgfeEOPwyKe7b5nJSXZVUhXaUx4MuHHLgY+3S0QK6YHJ5pt
KHa3EqdTRFNI6ECqjlGpmtwQhyMEeKfgLxrqr6b1fw2Kg2XMGztCFohQlsliVDbAMp6XpYvR/baC
BpB17ODmzn/DPq8QSOqdta25LEU4nHGXi4M8Kj4iNSLrsCYuFBGZwwvH8mwSs4X4zcfzH7qb9+99
DyeAfNYcwBaCNIGwqG2vw9Hp4Nby25a7s2n/L8Z4XcXpYOODIa0ALoHkxZBGr+mj+HO+f4FPyqxU
FOiSDalmvAKulDjCj2RrXvxYlv0HvO53eRduRiGDqGNtFSkEzNsoIUhl/s1w/1viDU82JySsV6du
FY2GJ3ojpyzM5khXuHJjI3AbBBuBvb6b4kMMmSOdYxJOxlTTgljC5OLJlBQUzbbSUDIV1qv1kDpp
lyLfqQVXk5Z5uXqPWB6AwvkM5K1UoTHXJHFi3zQcOs+HDVkReG9/dzJITX5re9w2TEJtc3NmfUfu
Ek2F73wgDzAi3Et1ubcuYceloVwmltnhv3PuLcxYlsFzF/NyaezPkGEQBuzn/pGe7NiJGVBKd7oT
cThpvK/f2CjSFja0fCE1Z8TF+EEL1ttqUfw8Uy8qPAyotP8zfkQXxAoZkpQ+szgIo+mAyXYVFTJy
Fe/ld4U72p9JhmrW1s0X5guZ1wGTJ/LWjC5JPM86Tx4wxwvFLF+UXgRUZ2H7GjX+jaWUKCSQzYh3
svpO+xK8lIyRMr9DFH9ntg264cTsPMpUq1xjeTw3KmUARw+Xr9TayR+kITQ2jY8s9axzdQ6nYyee
Ih6eaYV/h64IrLl8ZllBuLCjJ14vqMHW5cwyOmTxcgCR2TSP2U0DhCQrlRlL3jn/ehQg38+4YwnY
LBBIWZjhMMVE1vPRgwWzEgttVt7VKYb7YfKKS7VBSnSC7EY1DBAWGhb2/OIa9RKY2WIZBF+c1B3J
Yaws32fdfh1ZX2HLUIBbS/hsZFAG1jguPfEJRsX/MEh/ZcQDA54MXQJdUkcFFiZMBlUIrM2DGgqf
qbPepqCumhm6deOv4V3a/b8XoVwstRmg+/o5WRoMvNLws7SH3FcLEbpyxoqAPV7o6BwRB3GJAOfZ
BF2hVp8veY7prA6dysA8O4MnHpWAeSqWJ7PG5u99G7VuzQWaRbpVpnJP2qEsKfbPGJAqzulKGdP9
7+EyJ4QNC9EvBtLjoqaQRXAvztHm4eGeJ8QQEdLSLmwD8dbaEt8PyhCTstS6p9CDjKPYruDuBY1Z
6LSPXGz7xDJfZxK6S35rI+PWQqknSDP8glGbHGePk6rKtrQpHleZekimtCoYULNh4PWp+jSyCEs8
w01+0g52O5UnwTMKopIJW9NChlLqBnDtFSiq7rcklaqOwOZUi1mZIGAgefADcOYagw71TgHNWltt
EPE0xtI3woAMubsVlBHYBVrowR9LkhSITyMG0ZzRu38GSlIQf21AXXoss6kXnAQSlouPgw0sXIQN
A9SpHAf1KSRcJxI0/9QZp4K0+lhq/A3uS2M1f7KxDUgBoqbrhoOYXZ8snSo2lai4JvXZxlq6QP5I
vSOERcpLTuuEns4M7P9mzG/Lc5rhfNHQ6+ER+325oPOHzHwlhv5mpkfI/Ka6dC5ANbqIyXfIlJAZ
X4+a6N+5I3syptAO+IK9qWI4eP6XSscL3hYJAdF7g6Qfq7RfSsQibq0WmH70pObuPHVnS67nZGyA
QtR06tyna/CqXey8lX1JwdB8H4lBUBZghfC5n4F+KuXsMEI+4iaT7/+brCNlxxbcZVvN0mG78mHE
aCzhjHp01jC6VNAeGfA+FlfIEckxONO0rmWZ3dQGhyagJOTr23bHjgFyehpW397KZ2fWEOGG36yJ
Yb5tU+Pru9/BP+K19+vtlHf6z9uaRnhlhOgxXg21L6g3QfgMRRFw0+3lyVCcrAlcxVeCY7sE666q
XVsY/rjpNgGPemqpZbwQvi82qaVpEoITYMzR7EjpIOp77nEIA2DcJqXz1YrkdU3UV9RVY42weY2F
eeho++Y5+V0fBAPlzj0VOcXg1zfm/VaxBIY/LtiYy24aR5W4Fpw229uFqfFanBLJlMm5yk2sECn3
EtFeZocAu9c2d0momYL1MlvbM6dS5/o9imD0mGO9FEq4wMX8f+8BHw7qVgtFjTzd0jpyIAI3kKiK
RhF09DsMYHsSnRdomCDxPeCVmJsARvOMiXTJ14okYhTEUaUkk6LBw1cSB0zmXtob7lNJJ4DPzeCf
qQrKxQrX6z5b5YZY2gGPd48YEMXYP+lH8RcwObLXH/fI9h4Sztm8zwDDY7hGd/NozdTGauO470vH
JbsNOcvnGnM5lba0qQ/H8Kr+zidvigA/bbKdAorowyr87a0qqFrZJbKDAPCHXzrb+fHlxPNP0ds8
AtYuxj0pltqRdlJrwnTKsUTIAvxpjhKYP3WpqN4TPFwTY1stN/5G23zswlAlDnI+qPVUXcn8Xp59
A1vnldcA47F4CiNkeD/nEnGd+uffENAFvztCKg1Ox+nzNhNtL6MmwdvNOfjJk7pA46vlfgFrXTpR
loa+ZCqhq/VzN/QBNsCUCr2FvY4EXgVzhLTQKueheV3/eQJo7g7cZNtKJoVDg5azGyefrdHM/V2a
3VI9PHP5cUu2usTCC7Et58On3EKMdgy4m7seEQytqdPmfZ2cI0F8t8sczbkrCTzUhp/LAIZjPCJo
lOcnsr0ksaQXbSQIrCsc2ekmdmRp7k4cylEZJuCvQJr/92WKiq+KYQymPjHZuITx1vNphdL/wQu9
pBvGmPKKCXgx9NMvRCRq93qoqRHQe9famuUAH/54bJJxgsv/az9PIirDLa6yVuwrkgsYvvGDsn6w
NDEv3LZkWLv5abk6C0mcT288sBLfwna07TKHFFy3pTB+VOb+dATK4HS2T+ydSugluKYfbg8HcO3P
jFhmo5m1ut2eESZV7alPsqJ9EVXqfo3W+jhhSQK18Dmb5GbYUNFS0yvkhfmM2O2EzjiYRav852sm
IYn9AUFRu365neMEnpWF1O5zDQFTqi6G4V3fC0opUlYTb0Zt8kzkhLEtk1SpslSPnBO2OMfJJDPl
QV13QVRL3lg6RbhVHyCtUucGiaPY+WhmytIbP4nxaN9LQtTRNgpj+IuVcmIG5fypg6BrR4GuEt7V
jVXOpdu3vehq93NkgmBiNv6Occ35Fr9YjVh5bdJYQUc8327qa4gx3omAC6xKLCYFFJp9ejc9N58k
YlNY76Q8nYhd37mGua9nzejJKSjaMgFwYa6+KaonSY/yYHY0XPiqf/7JNSTP8MJ2f6WjjkItJryS
7gDDE4ae866o+K+90HEJAix+XnzMYUTei5+vRmniDmiwGD9fkJbXAINP6aN48CJ383d3QbfAaLak
HH+wt5eLr/DelPsoCXy9GkEyqvosDraaIJHKZBCdQ/N/hdW9ahqjRAxlEDUxS6QUlItDOq85R6HY
/5jEVERIpZNS5Q6GeEKVbh5vOdqt55IxR/FGEh9lSAr7phwBZX4N+rxQ2BQYzocXP8JOcLV6dEdz
63T5wOu4MEZY3NiFEVLTKUk/NyZZYKg1ZrEYnpFmTBnRegBWDaPOj9G8ugmXkVe8Uv5bG1KTGMCj
YpljS2DLIrhYRLufNyB4jWYIoIpQqu1O+x1j1R03p00lIE3MNjaMlwI1FQxPZmGc7dUAp7Cd43Ne
rnkVpaGymOlnO4gAs8sOeJHC14by68de/vTB8by0XQgXf3bSVIeS2tbOxC8mfEu3CIERjXMfEaSz
jQBGg+2TQafm6Y+4qIQocRY62bhXE3uOzfj82EsvP3nJxjPyeIVXeY/tuovedRREYjHoW6uiU613
7z/gezHkYmbU2Syz6eEyU6OVSDGfgKyONlEPOSgf20JBJLyOke5GhKtcv0f57EfJXG4rhhtuYYW6
RjCO19IsLga+zIRZ54mrIl7pdpj8aStft5kTqGbjYHPwW1FTaAJaCZVb4FF/xAybGJ5+b2jTwL3A
0UuvVUYck1V3H56HBlKxh7FhtYeqv6UojurYo08Vy15YuRWLdhn7mN4h/nTxUsXlxJSupWuciw7c
syNKgroy8MIYZwtoGd7vi4hqgNNFr/+AE67wtvoq3ApfyQvIuWKYxztJ08t6Uo1w6VkJmqXGqNpi
ot87o/1adQa4cbrGT4erqjY/st6ucQ1wtuTAKFJlgP2ji+o91VATJKwslZye6gARudhMvzq/s+iQ
7dp8/DjTByteiSDNhjk/gHtu0y9xBOmns6x1aHhU0m7B9sM1VH+FeVA8aICR3rLJJc8cU9jjfyDC
Bv6udREjtJAb++mKCf9eRJmI2iobTP0cRdxpSy+n0FZFVgbwvjlwqk3NLjFB1Bcb98RErZYx9tDr
Zu+o0mIjd5XUPTVsj7Bs/CMT1ai6xs0pBtJwAz7bS13i7KW++eaJ6IFbdonneuqaf4dL6LxcyL4q
1RDO6h6/n5+xk2BsQ0MI2TCQzHw9lZxPywPo/SNmwzv1T1fT1JfaqJrvsxv4bcp/WpOmWRWKduOQ
HKq6HIx15u8AyNO7RZrGEazf+hS1kHOIMsamYGrIF8LO7ZKAuEyY4siJ5NcpjehcZNiTZ4ozc3KD
6SlNVejPFjIj9/lfrk8Foi1M3pUeN8nuRqqxZgURvcPMOPLhsapHIzA7fEB7lMHNm8kxcOhlvPe2
3P8aSF+V8zDs+/hbeo37YMXi589i0KpMFUzp0eB14Hsfzepd2ip9M9JnxiifIfej6njK8RzJMkqP
e7eqRM6TI5pf17AUljLiJ/+12drd+mDFfQhFn3zXN8NRmGkon+D38FHS6tmQbYseZJGMwKe/88Eo
KSKY2voRcbEzwm/LYaFIe5K1MMR16tlr/MTXv3ZV7E/lZrVJRTSeeDzmR83eStp/hsv0TWCNCnOn
j25g/lk0oVnlf6mbyWbmGXKNtDf9AXjKu9CaTXd9zBVipq0jHdpBARdyyLQoH4+u3u2UMGNnKe4O
QWAsi25SrvM138BhUGHuoCMb2jwrdTjjhFxHCvuGAqhdFvCwkcuaB7QkfLyxrK2noWV8xoqB3EJY
whZRwqi7ZGkAW/9UJUG+z3dqWD+roDFZPmFwOhmk09gQaGNVtLUMNaU7XQIGXsaWiqt2knU61Yvf
uYBcCiYrC0i7CRpkO05ZGIVAlV2L6HXLHrjOkCWBfloWnO3I98MBe1geq7kVFo1ic5xMl9MzkA3c
E6H05l7ALF8rGrKnHc3V1WY/+duws+yzgAxGlR7X3+5+je32ycMWKwvRj8s9sg+/SfWw8bcbNQlb
bD5aW7CsJAxUDM7Ixkmro/sCn7N8npIO4tIIs/2CH3Q1zRYn1SRNhALsULYMBxa23rBrYGNsg6yM
/+E1jJNz3RM1qaLjBpCekY0csGKkXkRa6JL9ZFtFuTnOHhB5jP11FfV4UYkTS4WvaoygttEDbMrq
9Gpew6eFD957V+oC/g2v9bo5J6s3ckqlrShlG2l0gyTfbjfF1LXESASJ8l/WF8Lfv78rL9Lqr0bu
WmHDg0NjC1R2buPBZfnFmTeTmFKU/fXBYj7cA6U5AJM79NRTTt0NK426e4JV/DS166ucAblR6TT/
OJUK1wzjMmu5ENyM0BRtxM1clvrzd8AU3haclOXG4vXP9RxMczTSAJm13C53caKRmE6o/UKpnp9w
q6XqxQOlr6jAycyVvxvEPeYHVYFnTJeC4Vs50AJsfKXLvpoqvIiC+SW+QJrtCzM4umoMgxK8eiqp
nvGZoAa6Mu4uxRaosHgfaRnBgipxEL4tUvkcDjmm++Yv1T4FFFX7/bBdVDQ44jq/51qjM+FZ11KO
0YCp7w3wtLW54cpcNiWkEnjbmOyqCzh1slNACIDQXKa+krfmRp4PwU2Q8UzFcx8Hqr8bVVCY0bP/
3klP7MQMFeeJJvhhC9SOfadyzt77RHvVKYcu/EtLlH+fhXbI/ubmd3qwy/tlVmcAwP0XNuoXcEaV
I32ztFyURW7wzEF7ZAW6kGK4Pq4qpGnR5OfU+M8+ED0LvJs/+tsMmcSPU6iu8BzGugUA2gXSMXwI
9utSr6SOWEcFdI7BUTZc5WxFQSu0Rhyg7CMj3JwnGDOi1ItfFuwxGKtAM1e5n/H8zOuI+OTHrdu9
cUpkXbuFr+Ab81occpH6XYbsxUdcRbUgYp3YmDVKBn1LfVDOzSWXda1ZHyU2SssvsQOErhrN8eEZ
rMUXOxPhUTLrty6U4yFFikyKxU8tGp8R/HzS36/cWLlQwbQ+0ePzfRW7oQGYHqv8LVllvgVT92DZ
n3CDdDFcbpvadSeSMHB8ljlBSvmFV++HhAWHwvwpjSNfnbaOJrThKuEmWP3o00xjFddot1pyXs3Y
AEmhps0D8YhX9/ad42s+Nrsmmh3W7xLwLzDhl81hIEzcTQlMphGTUpIdu3WRMEvVdwzcAlBwSlnz
pfQfQKLA8ySvQz7RYp+inPqIPimacMlnny4uxRssDmMQgHkz+EWm8/DD6PgOkLh7dwmjnJd1hg+J
HImo2mMkiTHV0GfF1O61r6+VIrFaN7vcM7261kqP4W2T4PaApbg28QU4ivuM4nH6djAeSD7PPFx2
1wB/2skxsMRODWC0L8b1uJQLs63YYRa2Rvb8DbromqPAyEGwuvnqnC310Kt6Qwk9h5g/sYd3U1q+
UUiIlqfXwhI4HjZPAL03z+3+4cDvE1zGObmOZ8LIwCFTdUKiupriFaK45qOGPMivHvKolb1qOCq9
VeQrg4iPpn46trfW6/Hd8rvyWEEv2vvI4uT9QVHv/AM3y0GnYuk6DpKVQKtigSh3ueGVZ5DOnm4B
SMV2yu7U7A4ZMb5kvQspBUxRT8cZVHjXYGg7TiIOiC/Pe9fVK1nY7mWaqSUQ1PRiJNwI7BCIOB8m
kXytgEWFhV8p505a3xRC6kOAygu3cv7BxED2vZkJUq1n/DTqYWF80MIETsKJj+8xVvRTNPINcb/I
28nAcN15SdoEwpVFlbVbVwLJ7JV3DJt7tiyCWDxGdPqRl1htcktX4HysfuYj732RGiLnGwRGrG9n
oEXg46n/1T5Cku52SUw4WiYnT6TjZ0LC0WWxWDBKRKhLuoK9zGnrSm0hZ5w+YSlRRV+UvdTKqZkt
/gzm4C2EB2k1jD1qiRg25hmCVfCbI0ztGSNN7YlRgBnvUPKeBg+l65f9ug9y7SX3DslhoRJGo4qr
gmypkk5CroEGVOm70Uy+Vg6HrTOhFHN9SGWyPiX4UgsBmyFqNhH/8n6eo6yPVbU/bevQBJ9wCNFD
U7akudM6n0jBuEy/zz3f2Hu3WbV9NTjgPQ5kIXyJG1c5FHbOFliPzH2Tqy0zzW2/OHKhHcjILHNe
Aj0gS7issj/eqZc467tXyGVm0VGJgsNsh51NbTE1o3f/EQtenwq0NT7WgeCBmhtshF55QcTeohPX
OdVu5bJXl3LCR7c43FY4IbQTKyCevJ2BOnBFOfHQgDgICY+FLjMoyH1xWIfxpp2nH/4bGYb4l93j
zgxGlyGwwB0kMvBn49wAOgLeq0XFhGQJ43E2TSqTgRKp8dw/BML3cyLBCQvzSFCbzxdPq/gHOJ+s
7o5/IzgkLHYN13CURGKK/qM38v8JgAqO51zAsEyUeSsiBO4PZMY+08a1Z+P0Mz6NFyt/YQud5mu/
Jo9HdgA2lY0USjeXoFxOtW8mffY1LH8h8DLYtbKIj7L6Yw973YsA6PG+YYWLLe4PsJUP6HioZ9M8
MKk8HrZey/9LVwmMMr8yP6X6c92b+G1SOio1TcYaVvTmn2MhYtfbjoGvo66HmJMgEuByQPKMDgui
0KkjOAQ6B1JUR86uVsgOdp4vSNQqj9PLOLkpGkKBRJexvHySgweqokD8e8teZqPwdZv6NPR+tl34
86lAGF6Vp4b24a4sTWZ1ncpfYv1PD2+KBbAy79CxEI1cfjm3pvpq+w3XniCS+Oh4aMw9ODvC2pxC
9jwQa5nt4iJjNBqstIcR13WIC+rYWHi0D8yInM12ZMX0EW80yonFSvwfSs6hJdG1N0PS7VaoI/pO
QyJKZ46kNuvHfBfGn2Q0jNZEjNksRDdVafWjIuYoinlQ2E1OZwQTrtrruQt//GecXENq2zNVnOh2
7d90NPGXonnRNsZvrU7KlVJrdUyxNlaFN1maKXFfX3oJQS1K9EIUPDg9a0zCHVgESK7MR9ows756
FTMndPgGAUzb8CvGfwQkcO7TxHGv3Pol9yAaPZsrMDZGRzSPZZ1VEbhs/mI4yyGr1HqFV1H8t9t/
Yt51F++nLIekjJWzLcAcg1dE06z0Ts13u6J/D3lGfvyPWuga2e2ZIyVjOVTPLgYgYCFYJoTqvu+F
KFiRhBNQjayb92S2jJQR6qKX7khtHzV+Q8G8xMnx0IDigAsynteFksZYBLPU6UHJegAHHd6cfXsj
FkRAmpE8HrDRA+rhegRZ7QfImOuRaeAtZ8BNl07MXbN3G4FpzmI7bgQffKGAisbBFx2J9ujtMdev
E6NruBWTtUNhSkGxenJmwrzvXvXIG8i4Cgz0oWth5AcwckDnARRHi2EniiwjJAL+EmxnRgnTpTGT
QQfnyfsWan6t29qdTxo4svMIKP2kNg4jrfQF6stF3VK0Ak9kKBKfNNdn5VIiKw4eNNt2iy+yXof8
nAkLRqmh/3G0HChJqeNeMjjrsOaCrrVI/2gfAYqo+WYd6sfnJ7a558shFNRNtVsTH1lagCNdsZ7J
2sSMYP+itQ155HrEJbiWq6DLPpDuD1r3iyAApgUMan5479kczwHDROBzfPN7wVCVBsQJF8KVyKfp
0KXZLhWK5PtYnUdQIHagsqdjbRehtO2t8n+WcFxSBmRJNJVihcPcZX2W/V3Z+LagT/gKnpUfcvJd
gU0h4ySLcDxSbwIC8ewUiQjmcCMDoPWs3umjVqGwEiQmIPyAFo7AuvhziA+3KvmFMKBsi5ZyerVW
GTCK7NLMkMP9JmdiAk+sqU/gtmy4pvdvaO3y2xoUEombz7oEsQ5bh/2eh2cjlQxvxgs9fvjlcrCH
+j2L5Yr+3OPlMsqTOLomnrpEYKBdXXTPRgGnhZZUuGE5hqvRrfO0tj2Iq95YTKfVpJS6ZcwhhzBn
StgDqa/ZQyUZ7mHFrSJz2Q7sCM7rEa+TESWOgWhh9DTXm1CNnUUwNX66r4yYgpFrtKuOtCcQOdQv
pD0m72BSopXzwJkxJD/2RUfoho7E/mFkfDu7gvs0aQPSXNji5m+jWKQ433+IJQ+9Fnojn9yPpwij
bHiP+Pg8bZ66HCtZEO+5SqqYNz7FuWki0BhO4WnuEKwxhIVe1b04jgvBpC6QP0csuIapNe4oAko+
w6i9+jxmSifkYY9sEJuXdmvcIL4xJMFcXUJeHq9w/HV+froBGBCbxKkFTAJMpiepAGPpy4iGAsKd
kmMiYKqSt8n8fGWfyU/67nURhnWUqAbSFUbzYzsxnQeQAhmB0eOLl30fppr3YsTY/t+bbS4/jZkU
dOtB+CHw0+HlNIXv1vMTiuOBdHKhnoaM77zmMOR5CiYjWEMtHYdU8cPqSUtxxDDPXU4GdYMwoG2V
060tAcER+EcEMXP7uJgjKpNVCJFTsO5rtZoe+7RGQl/PwWqZGKfDeUVM26ZGD+1Q/qZMqBN9IqKF
t6E0h36kAU28WXB/BuRr/gaTXIG/6AiILgqGKqFD3aGe/OHMn1XXNc4rdHk7Rf2hdfZF/B2Ib1mC
obZ7H5y0omdiMSZvdOsrq6PyYoe1fPiyXasW8DXmW3AbwHUzLS+mDiKx1FmscOw0oeoP9TSiMd7n
Q5fXn0pPu9n8iqIt/DIjmrTCqZBg/FNO4WizcGtW3VEsv6i+i3a5EFQe8gPImoGPLoFYScWLB1os
hZopdHIsxoNl2IyZOxKcteY6vFDsEsS11cgzXW2UjKHQdNcb7AGPv/2u9oBkT3X1ixKuJ9QTkz2A
la0+h/tBuEAtO7kXXi/yHW7bHRLGIOCB6BqAUutpw/JP5b/N2uSpm71gXnHHI58oZjoNU2C5M3fL
F/JMHoIq6Lo1rcEVVOS2WH4P+2CkoyLgZfi1sX2p28U126SB6UDHGKtoH28yOFXDrAoukstIxVQz
BWQ36N87Bwy+Ix6QOdSf6JtsSzOpz7G9oDxZbbkQPNnQY5o6pLOX2rCXqdIAcdFGuDcPTqhHLPkW
octAppaGexoDICdoDfFDIQpIesEjDhUUddn4PNqkp1uL557vPOXzP94dONuj7Lidrligj+3Awmlu
y4VrH5WA0QvQKqas9PWvdUCk+plzdf4NiOZrMzItZTChwS4q+mhOdDIUFaCvxeNE+nsFJ5jcg/55
BXithnPAuj4T7kcUyQeCkmtZOxnS2dPxgb62hC1P+iN0k4EiZO8BeVIx7ENYodVtK4KUWTWTW8Cy
qanRIZg3hxXounP07/Y5vDJqOXPUUlTszckUTlZXuQ8oikXVx+zGZp0HSUi+SQdSElmMUTCWybzH
/K2DUwauipPV5BETK7qSlvP6BtysP5k0OD9G95CJAUVMx6TFvJgcfIIP4hbS8nREt79TvDaF/t7R
GAFL5t6VKzNpTiL0G4eO6UsqvQfCfYOYpC1m0rHqv3bYb1KVpxtqllFluosPhMudTapJqdOOmAae
khJ+NHkQYkiJiqkdONPJPqIcruVn7Pa0Up8BurVvng3MF+vPnJQNzt2ud5gwplugnnb110a8P633
YNFjx5FxdrvU9oHCxY9Oc2zCWonFSMiQYrrys9YBeU/m/AfvELAWQ8ja8qhkTfGHOHOwgQeQFs0T
rOjxllFA4F+YLKurkQFxC2EQsT7co36J7o0Qkym+fgNp0FvF1KyhmWYdpNrRCDER0MSWzYJs0l1H
op3V5deXMcmJ2O/qo4fw4VqNqdEGdzfVmz9bkvbt4K10UOAGKhvoAYnns/xJ/1xIwSF/B/l2gIG9
nqWc17WZBqh0vICdYSSH4peDriF3NaYzkYPZa+IiPsGyJ22i1EZe9BkSyzsYzkHYaWvk3tAtz8a1
Wfj12UAQ+u7uymE7spu/u8wXBMVeuEFxsEQOYlWUJ4HXnyA2Vww153Jw1xnmTseIsFp/fAVrNQRE
gEibko28Jk46GvNw+grNdGVL40COTpdv9S7eF3wC7oj6A8ta2pZJQB5ddlNCc1xJELcSJ7cRMnaE
F5rVGSm0tSsy22Y8rWy4rp6HoMuZANu8W8gXIzi21YffnmRAF8qI8G0JLB5IZd1RqyhVGb7EgIXh
jZZclMl7QokhxQAbON6saYsNUd2Y0k7P1xb7dgY2yYJ3lrIz1t4HsdNjcrsAv4Dn2TcTk+e7HmTw
r8EtU8nn3yDPv+bS4Nrj6w3/60tt5W7ASaUvv8SP+EhBBiFUP/3Jzgv+PqBcd/asL7VwNP/oRRwG
cK1U3TNWfgLszoZmzntbAD298z5/CMvYzWfmV6YYAgmzI9pwDbGL1QNZpcIK9yrTWK88k4fXWdN3
vfZ2dbkRFqXYDVTThs+WEOuSxa/P880CNzjUW1ZdUbpcxkzdN+UNo6kzoO/kNuZfzft/1f9ay1U6
ijfVQO7xcNRJEnzFh2cKQFL043rbyxPK9r1XoPytfXm8d6eQxO1qRK7y68ASve5oBA03IBIUX4Yc
f19vObFbbu/3RsnPOKJA75DjGpMdMM2gFutvkvRwaNlpPxJfRTffjfGMEmSErGrfyrH1pC6bw35s
8V5IObYylvP/PrzRLCaPA3WfVelV/pqOkgAW5fBVeO8FFEwr4qfYGRXUH4UmGkzXTdMp2hiZvpTP
FJsXlj+XCAxGIY49cZkJFWaRVearzEkO3VVT1rHqtqc7QU73nmpmdTYXtD6fg70O0SlsbBo7Uezo
pBs9okFr9ijAaP++XnMy+1I3qYj8VlWeXRsLSeT41ZuwlzD7qIsR4nyzkMOwXnsXogSfv9307okD
xIqPZ2jowqB2fTCx98iCvyu0k9gVKXm5Dd7CXGSYaERnzm6ovzLqWfWiFHPjbJy1i6JX63+abeom
Yfz90l4YayIw2k753J4EcR7SSireSzBAufeqDqOoxmDcrFEz1T2PDd6k8qhNmhY6/hB9Z50Ig91c
g81go79oQdIndp8CNMCmVUYoKlwSQt7VSe5J5XICfwxhwqlVFUxiB0dTXFcVR0nXh2Z0qFd0/MU1
TONY0zRDjjjIUtxyvVhzDQ+QiHyFn6k3hSDY+O4JMUEsUwo1BqKkIazCEj5CzVJSN8D+Wr3htRBP
c9msHB/uIZhiE3M6pKn9Ts1T9BmOUyW2LrCuG2JyK/yY9AyGn9hkrDyfYcui9tBS/fkQ/Q0xMbPO
Fpn5/uFqJrn6FPDaogJQVQ4tfWFY2lm008TFCKuA9EpA2iK3C6AQkTxlJTt0yq6uv6t4/5u3NO0Y
8nbXQd2u1VScXwWPhLEJ8wHseg/RTa2gO2DLnB+jq7SUI2ZBZgbyBRnhilvV+fthQN39KEokDcCz
3dRYYKGWNoNwXqogpr/U11o1lsnAabADPG3RhpgQOXTa+Ay7mxuOIkjpscVXqS6wwquk8po2g0eq
yesZaPGtzyvuxRcvgBNYQzsaU86fDj77QG1G6eJg0oXw/jXk4pmegHJ1nH3V7z5URCan6eUUOC5W
/so0mRqsS//Y5/owaJ+ahEh3fOKef9+Q0NRXZ48f7SYUtHJ8TYSqLdOWAg26y03I/fG3LFI3C/dI
roUeamcYXuFHkcUli6Szdjohcw4g8dDTDEOvGDKaZXqPzJaQ0K/r50PZyN0oRuvVrFDKjMs0dqDh
DD9rkVeJCvFWmKZSbvQBz9OHzfbo73Ya2btEYfvRtPRLv2LQbVu/3SXe0WHkaKCF/2fMYXAOv/wP
AvSuX55vQS6kCLSv+zELKLBhL8FMqMiGxnIn+Uxm7FMEKuhDjglvcH/2jt/AX1b8qY0QNiaI0jMz
sLcm1fbw87yF7vZE1U+tLJtzA1VYnPvueoROJbS39gZsoq9a0Vuo1QcShbE7nx9R2YNOEySAkflZ
bGyyQdE5/vG7S7C54Of/KQSiDafq53n8/ZpFsvQ2dJumYwJsCVw6NB776Atx1VN7jZiUyvPkTn2a
1aNDO6ddfkRSh/siSQJnuotUpIszF9bv8RIyXRwe9fZ3Q6s76c2HRHl4f8Jb5GG5AZpKGya6EP3g
JDpJLb84I38c62dcy1bK41p34MTY+QN/62e9oGd0ZxD467NgYhRE+0YenzzTBFNrYIXCgWl9hJck
80brA469uHA/ZvfNBM76yESMWlJF5udwDGNgM2aWL2ARJE+3tH5DnqIddUHtFigV3+7KEKst6IWc
OvrtT67MKicpk1SaFotWjgHCpxBH9mj9a8QECZPqYtEDXtXd7XAfnEaMW3Ah1sNslfa52u3vk0xo
C9H11N70UN6ye6pJ5m9Nb/C1/pLbzPgJ/bfpWmlfUTuZaBOPYvE1y+J4TavJMqLiZBUcmeLoxgi6
rimcHyqowZm1EKFuRDuRCLKD7klIZNS+wjo3bc48hNVdsefaE2Ssk9PzoVfvKKOKGZ9X72XmvVlX
ilpDY3H9z+nFYV7FmwAoVoVGI9CbYUm+2eNI7y9zGUkjjbuaTM+wAHpBaXIOXQQ6d7PyIeb8KENh
anr1m4WtDzH61nd/tipfnbpq8wZfpm6isTvQ0QgeFXo4f2nkgQ+nTDAQL8YgHNRDLHLvNYv7a5kE
npPZVZ2z3ujpGECFZflzF27kytiScC3aQqAwqT0/COtrTrVVZIwAvfBJUtUfSlQl3/KMIem4DTCu
z2Y+TV2E6JlAXrDk32MiwiU825IgbK+VE+J+G3CGHb4Zsn7rPrM7bIO+WmnUnK19cEEuQ4YFZLRB
KjLzbsILIVOEoj1Qui7B1l5YyX1hy/MB0crqWU069HgJ3JFHs5OutrAqJ9QdUGXTHD0pZV3e2uZC
fqepuVAGVLwvGukT/mBc9TSTLvquNbBKcL7U/vFbDcF/uhCRNJP95lKDzTgyA7p+UHj9ihWBwp9E
sNP2JqyGZEAnWKUB5aLngjbZhedQ9WXAnLp4D+crN4cb7w7gUEpvuB2psESdoUQ0/l4ilsNAHjk+
JluPU6Ft/xFQJ2YYNut8lTaotDTjYTGFHrGvoOKAYzJWzOGi2YJJQqzvd4ENMzQv1hfxBZAlEBVo
eBnEHglIp7AvsUp3zKKSvNcttOH0cjNKhrAgnN/qsMTCctq+B0ianiUyQx+DWt3uAzZ+lwb8CScR
T0pSpj9oBYqtlQoGbXjxKRvMtbxQ4Gki+JYUZDW+bTwDcTU3lytxS7y/WNyvk9DT0ADiv5gDH+hR
uDa0YY7F35HYGU2RubCuChVqkcLgxg4b+TSc/ty7tynnEzxabhrzMWR8oxbgHy0j1kgPj/34Ms0h
x3iCNbM88G+qu6ZFoTwqmQ4o9Jm44W5ZACQML0pH1daNQ04I8mfSeLlSkO7QfBcGTkZmnLtYsSiG
SlFAlhHFbr7CejeraS7RRS6m3Fc3UpuzxNgSA/1oLziPAs8Qs+sohDCefGq7mRJ4EVgKZQ+jXjDu
uIFKtRiA1MsHM0NbTkQK4GgX/7ZN9wr5j9qUMeQ6lpXsl3v3F6K58vlONeVKvJDnXPIpeG5ptulP
Q6L2ewYJiNOnGuP2/DgbEsHH4cqb8mkwu5AC+q+MpXmA4ou/dJqhZ4XXNIobrW/XDu826cRtOL7A
u58cx8QztdZmRhu6ItOzZ0/mS+ZZJtPlonPsHyGk8rUDDzCnIn7ilExu8ziV1UmJhwr0xDGpC6Ut
6AWt983micvWFIYJlIgm+sdQ4Yvmb8gQLYc/9+q/OBaR4WpN+/EJzwQl3KLyoPH/TIpTP6jKN+JO
9Lfv154vRLN3+5h+ga0032PwBWYGM9q3kwyR6+Il5ulzwGLB3vcI2cLn0Y5jL55PKKKS5ovexbwU
z1DU/As0n4Rwwc6MTzzJBmxZwyH/HofqGPI5HL4h/8dom6jWnwL7uWVDGYBjFL6KOKCzaOd7Bzvg
4yQJW2D8fomNU07GEFQzdsqcwxgCFjzrFMdyFwfppynuTmM2/xDRyF/l+csb++YcGr370aofrRIW
vWc9CwI90aCD9PTKFnv7O3RvPMLu3SKordCCo/1lAnLyiEmMdQsyOCmf0GHAkvAf4NqSJlZiCGVY
6x60bU7Dh568ZGX/VRfw/0KnApD8UXsgV8yp1jksOC7dP/U2l9phuJefdF5+/JCf76J39FnEDchr
YqkPvlFA5KCUpVITqLPk9C4ClN22Z0SzArpTGmnXcZEzxK2Ij6z/HvwSsY5d/kpGVFEtz9f1eChd
/HaI5VflYiO2tLMbiDVlExtp4Hq4MEbdIQvM6y35QyyZn3j37NLf4W4CX16/DKJNHsyMFpaJlLSO
AFWbuAXTS6oIisk2OO/zzRX5hrUQb3HanXplkJRlg8gkAvPpV/Eqov5c3X9M4v7v06kI5i1iTi2S
Y8ZjSHIeDcgQqIYR+iAc4hhA9WO3jB+Hz/iKQfwUm4G0KgtDPd2W9/NvntHlI/9WilvYvzEIKN5o
aAL7cFL6kuptIidgjbYrtTYBJ8Ptwvt+8RndLV8FKPCv9P3egt6sQrPQtiZ6ks5hFnpW1fICYQxe
MVxGM1AN6HzR13REOjghIMR9EiddbLS0taf1+t5yJl4kHnIgp0u00FNYJbJOEeupSzHCC/8ot53H
NxFFjz67GwGE/ROM1cIcMjoy2u6iPJ/TuemhkEeffj9LNYDH+52PPVN51LRuTmRXLfXB5PzdWR1K
WBm0EBk72mJY8c1xbK5EH4FDWz8dKT6CUAa5JKeOej2DKctzooFfcgLvDPOetQt/v5MdeOsyN7QO
CnIf77pay3ifU57ZrYQEUL1l8Nxea76v13ubjaz4CJSR1TDPMk1uy72S4GoZZKrVghtw4vyqgvm/
r3wN/ZjSwi80NTO1xywxbMBGO2EAH6T+jnoCfoI1gQDs7U33gJCy45+bs8sWDAU13vaVW9gpoGLn
tLyFZrJPksfAIt3nPXZ089JJmq7WeLUxS4vAbOTpQZxaXIFoYEVSv6ewR9m9+41CB5pg3X1SWMe/
TmeSz0/1LoZrPBsbPMhpPRQ6RdKinS68EuGfPkY7nW69IpF0eeKTatZFFnOYYrChrv4rqSXILouu
+KGk0N1oeC47gEqbkZbmKZsCiukb/bVuniD+CotCxmlQVQY91QbR2Nr+RVCeZ2qbIhr162R+yZ06
57XLIIM3hZxWJa2K9TYHB75HTcKMK5cq7OWzWw44Wx6sCPjhcjzGfWlU4R53zrj3fYnA2xyeVPD3
X7z0kn2escTBop+QNe+Cj1TNuSxD41Hq652vHrSziRjoixwd5dRqWFhoUp5ELZnxHFFQFUuzNVDF
WQC1kSbn95txqQDMc5i0KA8rItqgY3VtmmuMHaG230z6MXrHpHz8lKXBRmzeuGzLV7lB30vznVAR
0VpiM8eYMSrOKmDno2Ch0hjlw7FGkJtchExtWUzDf1nZ0vI2dT4m0YWYJmwqEFoxaWyDWgN29MS6
NQrzn/+5dfsNHPn+n5GKh5GyI9AqQ1H7fYjEzMaUD4oUpNV6UZ8gzI+WREDjXmFK3sWeAtHHPpzr
LW22CKvZMXlIvAWFlX0vp9+Gr5szylSJMsQPUwbEocLh1t0m8SS7s2rB6vI9vAjkgtFPbwm7hkKf
GKyB7sxXdUmWOVGR+hQlOpsuWf3Z9qIiKtWZNt6YBfub9WzmypHSmsVjWOw63gcct9nWbYRDJwif
aLaeKbHYFUK2nXML2lpuRlAQ6ar5dZUyw1jBGeC8KuPzYqz6DqyeEMqLO6+Q5RIJUm+9QmAHEeGG
UpZyUwiA+k3vB3snuctlemVyEOxgUyXBGFG1IfvUjzW5Cl7eoGEUB/sge723cwrujBz0Mv1wRlX3
wq0Wau+8u6p3tO/nRYvm2mFBeDI7RlAhbPdDN+yR6UcaLp4za83iSGflt6BWeU9luktB2pTUoDN+
GIPDbYZKIfrHETHwp92idiKoKBhevEOiUwNMAU0cu7jIDx1vm/OKwsdDobIztHiniZuVCKu4+YiX
hvllFh8Nn999/o2eT5Af0o02HvvT9vCR4OBMTkXLuHyisV4GPTV6NKg++w+v7I9dK1/rbkcml0c3
u2v0aMYpKahaB+zAkV2IZcCvFabab1I+eLHQy1HMNVOKqtbKt/GzjdHP2O8i31Do8y2kb/WycTsC
LkgMfvKxRRCgF4VRhIralpRJ/ZbJ72THLEaw8ufJCLEN1zH56mymoeVxQ0o7PcpO31Be7rMqxU/C
+C8p8LAhf3exhfvB9PPeah+MoprGxyJ8Uj44vYfhxgjX05u7WEUZz3GN6x2tSgSnOVrcD7Brd2oJ
ENfRChTsuJnfQ4Sr1WnYmFddZ8r7PD20lgNw6hgegbzS9uCn+ZZPZ/LeqCKIxcKL6DNTggOIR00E
yueKwSYHnl8+VuESOm1ElChIypXGfceDhPy5WNElJTpdNlLYoEWrsB27RO8z3ykRhXjyB5Ps2z8d
FfcBu2T7S6VS2N+yyUVzH67V1iVXsXbE3V/f/W6q7L5Q6Guu4M/SMbBM3MrXhZTuaXzEsR8o0aqy
1LRW+ON8OsQweB6NLrGzg9IeO+rQelBJeOtpCfzfYFiLnuYi4tre7Qk3nkfo2e+SyFb0RarovMP6
1vqFq8FHTR4HluuF2/25Jvm4B5wKo9tCrnr/EkAq4XVXTLm2CDaF5E8/7BRpqLzI61uqUKBJKRm+
P7g0GZwezEu6dJ+Wrq4ClYbeo8IM8Puh4K6HYdpYkciJOQk79tTVjZfYTtJVia8QyI3iCm8Q6Rig
TJDfR6Fv+Ill6Ui5eoAx2fJagOCeCsMhGBajDn/JjBdw4bUV5knJihz0Vejl5KM2mwoTn/kLRp58
l/2bBmCiLD0feMxr9phSQJLXv1ZK+43nXi+5wm9YkS/hjWD0qffVmRlILOMKHUzSYorl0V2XHdUp
ZQQZIDQFSFGHUESAlsZJLAFRwOH2dYoD7JgJoVpD0yQwnheSGIXC2YrLcRwVZw0nXV2qbQjxdf4c
Xx2opmu7HOzgDOQf7uedcMOsbnioNWMO+IJp83C7yNAwXfdinclNAUUd7nyf+sd37Z0WNwFbfKKs
UH1ibbKmcHrGqNZvj+SVK7KjYZhPcdu/OryV0ySxaM6cCYXVBEgMMiaScwPIzRBXKp3JlUsRTE58
ij1XOyLlcoB97BcXD9xsZa1nAFRTScFQWIaxJ1qLwrvJfhWmHZl8bjA0xXnTrnDwBgEKxeZikMvd
j8lPS/sGQ2wK8+g2Tgd9w99vVD7+ZRmvu1X2V/GSSuja8wpQsO5oCjmZR8ruiBHYKPZuoUIyWcnS
8zbOagEGDcoTKXDLhulvzy76I1COeuhVhPbha0eAfMnoPfYd8Dzs2oY04aqZe5veKNEUekAGR74S
/Ykc3bv8Dl/tnT0uBj9TIcsrlIY0rwXXzZPPKBMqckrcpJbDTALBuWn7K+ErDgihe/B7Zb9vu1oo
tKfHl0S4E31VBjwm9+O/krnec7vFhTWsoFZUoxYgOJdzI3QTQi9XnRvAHn3egblkNacewnca2Qut
TH70eQQnvRrVGmNGMrVP58MGI6nYLYxlkcqb9kLM6US4h57qn2j75NK/1TL6uHtkUbaTyi2JfCpA
qTaTDKQOBb1q3G6aaAqlkNHLzX7GUyDDzJ0WeL45w2Sn1SOTEmUK904Yo2HTQIx2Y4VjT0pQPF34
iXsyzC+8Y4trGUA1Zytm2t4zv4YSfBb4U8bJV63jwmjJOckNP+XNOW+91W96DU60GJZ/sQBKcly/
EeOwPvxqpSqlT5KRN2tfu2AKguw52raNaIRIR8xzI8g9S8qflNrDumsQ+GS0253a7FxsCVBuA9b5
W+Wl0raloon20qoG3sWrsNqJ0/sI3Qeayx89TX+Ym4wV6G2UiaS5PIhjwHeck4BifBFiTBNM8mxc
pNkA5YwYNLPQ7TcMLJwe99/CzO9/gilRo5+OO3mAGVcWRlTbmSy2+oILHO5lQFc7lqgLB3sop1DE
1sHqITsSbdI+G123KklGn5RKRtpoh8dXmEW/4yZwvNNuLQyjr7hV2c6DjjW7g3Y9ziDzzYuh8E7c
6Q6EftYyaKHquHDx0EdKEZpxCzFGaLq22oliJcQodpCgR6ipmcSHkzkRUya+Juv9PA28RdWGSSre
d1itihAbOcn4KprxMWOBoO1kNq49jffS3e6fKj5FjZ8/yp4yNAMiH/VCtZ0b1JIa8OTtOSbJ/uYd
apQ7CBuTgDJBaouC2A/642QueerLfoZBir3jeKjx0Sj9RB7fo6zbsl5gpJbw/KsQZ4jNPgk4te3R
0AJrhWTBbQ0ZzqN8zLiL8RaOuhG3UBlJ/31zIZv9HY6RGAyFeXH1nmzZ0IMgUGQ3L1Co1OeJoe1j
KQSuQfna6wXpXuBxMvBq8a3SBpmUi8gYcfpWGWxoGY6gT9uusyMdX3FI2E8WlBilIRHqa0BpDQr4
070BOSnvCq5xgVEqDv5PefaP74NzImwuJR3dwa44HztqC/5dXJqa98wuCk3ZV6sokAa4K9yH53XD
zq5/PkLI5N1Gn6gEjtc7P/OzIh1czMEdRw4ITUKE82Q53uCeVqxiVk28O+G4MJsDkj3T28gqC4XG
zXAgt9Uq5lBtER3hMouedRD+4tZWvZKJPlrn6y28JgfxyJO4FgUgyV7KU103Y0fi68VM0AuXP6dK
zWLX/7iBW7T7UVeKGIZb3WrojND3Ep81Jk/90QJ3diQDylwIzSRia5RmkRIoBpuqVXU9rZZpI0ME
QWgoHK4MVQJpoH7MS11K768y2ji7QWcdbFBpsvnXJ1WYwmwAwiPmprl2r3d/vdeNKxr53LA776gT
Ls1WLb11HDVoUtfD0xxaPZisqKwqstQGrWTcdJiHsQ8sDYkembLSSbriYIzIX4aWjxGUrQ4k4ERz
0n1+eg+xWUswJ08IN6oaHvJli1FbZ0kh29e2wlchC6BOWsmofwi1l+zMpaJh8sSkV6aJuX2fWj/z
Axo1BBWEtSjQDshjpL3kRjMU8H0W8GHoPPqJ6slnLrobcntEpCEke+/3u1J5UHFfyrmnpRFyECkK
1DUuTj8e2UshlnCsPg5AKC7O63DmlgBof/Bt121DuNzv61ZMurjwlwV2U5cdO1f3szWOQXfSXGCw
d/YL3UrSfELFEbK03su5LeLObFcUK2+u1Mn/tr7Zqi0214fq9tNj4stkB+JgK4DhF//QW4Rxfa56
mLtABpWoOIILG03f410Keba/zYkFZR5/flIIxvZuTeFTHjMTJnMcUhsoL5lIOb0HJXkfb7U7yYZM
X9YmnFqvz2JsOiLloMdH3xxBZRdN63dUdhqCZQqp3bPukQUzkhb9QMlPO8kaqIFVXgCFpxXeWADY
pt2EfzR4yZ6a5YdaUv5I933x3EkhR4qZTBo3dFo65zuSw0DQso6JvLQ2hImcXO2GjSuSQedsLWyx
lePwZ7zGNEWGf0NRWVQYko0IKtaPCItxJzHPG4AhuLOrDRFKYnpWySoZEocWXV8rdF+LEfnxC7Fl
/rSw1hQH6k6DCL0cq6PJiFlo3lJm11PCaqvVW2nC36z7KCXpaod3apW7P7KX1kQnWpB45a865BCN
05fd3svZJiTUOKxlDwugId0I18Ryt3tBxZ6B8dktcYqkbVDWsSiw7UusMqA+VoZ9LsS2FZ5NM6kt
8eIHueHKa3t3UWFoGtfKKvIJ2eymsYsipSMGs8iY9xNI6efol3MDJWPa7eqhQGlunceASuwIIMUm
2UWLi6liCZ1aXpZzxYwRgcuYCKXbh1dkaJIVmxmkdk2uvD4FxFuI9rcjH9hM20yrWwr1mKrzuTUI
m9I1dspLdekRv4Wxr7qAPyr9rQ02LGVj+VafxY9WdFlBDaGODyQrddRsjPPt9+3ESaCxRmMNMyyz
0E36/XfgpG+q19W3Y+wZ1UHvtl1rj//YU+zrYj6kSwGeqset5LU+c9LL1xVZpGmuXUQ/pJ45c7zO
xx8yozn9FKDTOuQOCsaufwihZvNgY2UUc6Xf0Ih5xGyBT0/Q/TQr8wjCzNsOhU1PbLt9gZ1MgYl6
mICIyzgh8lG4KWbfBq/TazUp4V6UieUyDsrI+ogbZm5nfydJoGOxSskSgLCiL8ELRohUiPw5Q7vI
D4UR8QM3b0MAqYrSCBHUbBSAQxV8Lw5lkQx1bs7/5BP3us/hUtzUJNMt1+XPb066dZyTtX+mdOzd
JUdw+OkATj16TvNOOl28Erb3SkbQ3xyclcydfKbgcDA+XqSs0g5rN9Nw7Es0/IPqVBEn4w99A0Ox
PvoPAeT5ECb210W/WBum6QRREmlStpPLQLg7dNHcnsBsRwguZrErgFgY2ZYmY8GLsfSucG0Ui1n5
ORcTuk16AZLaXFlFvRgYgCaBk5eZ5iyBGxOvk/0++/OXQ5tXJi1Qm58HAn05IWGpF5tVDBPqnrsf
kTNgaDEDMXoPs82QDWPXHRCneRltnXlW1i8w1DFMhHec4o2aC48fDpjaKZbrPuwn2zRXbMGrM1ox
70yUISWd3raQV8QBYIppQpONzlQt+lqM0b3Z/WU2GWWiRADNP69k77GjuSOhD/RybhrSuTXdN/ui
/NyDPaLBiaxk6ldGVs8/b539TClQGscC9atNMIQF+wC7KlzBv4KpMVPs+Jj6/wuY4zKrypKeWfQg
iAA2O3DiryFquMmAJHO+RLWZeerwbidRWCcEA/3RuCaH2Sk1OJU29YurzH6bgblW9ThM6q28/9Xz
NEDWSldp0TuIgHFZW6Qb3CJQcAwgiMT1/kGTxB3xrDE3GAPOoipJNuN1cd78Vsv5JTB46Q4LV4cG
IxltO1C1PH7chbUhelDiKovhg9x2I5tbJcrVP90ixh9h3ewbLXhMgLuk7mRN1WtdERIM/IA/48Hi
TqiPOv693/MzGqKjrRr7I76+9+0powbZ0k+MUGPRVpNrZdq2EqqlcSVBTAirWXLtoXVDWSru7ydy
6cqhstxA2Kx+gUN6qvHbtrvQwuP9cciSwD+tH5Nor2Z1jZwUTLMORB149DfIV4zZNrI6p4yJZKuR
eSmryzpD75a3j+jdsfcL0bIJokDt+zWQtzZQVS7rZQBeIMTGc+SnU1FB+U4armN1tJdwbcGz8uiQ
UoJqNYSc7iRQAas6C3NWZSKnzUVS85vUCgBOwfrxastlAIOD5UPvOUdgbIlP9Rqte8A6b8/5Vd5x
eR4EggY9OhAeV3596po94PASkrJcuackzqi3Nq404zQt9vDqbfc7z35IQZ74xjkUt+hsiWIjQf7c
F9JWHUi7sL5lHDc/Ke4HknCerQm12qUCLJVkgVVTP39eqHGv2pm9jKhkRb5U3DDNcV8QNn+B8eCr
8KIbXaSha3jssM9k16ethHkLcYvKD3M6yRC6Dre5Fx2SptNls1p6i6CyS5PBsoHnZ08AaIYUFTrQ
qF29vDwg9JhQgjCHl0oDN9dVMrH2o6EVxy4z+cZ2D+xvy7xv250gjbl3RLUd23VIhdIlkihU6Ojv
ZN5g/Yms9+N24RZHeDhu16GyWTUu9gFazKBsGu5AvbPomoPVSthI6tt3ksHBpHwUTrMI5Am98/Q0
L8hk3VwZA1I+ucEnyTTVfLrTFzNv0b3pOfS2wYJQDn+rWKG6dPCSRMluXrE0hSZOvBMVJSFrn+CJ
QAbcmfWO1KOcyuEUVYYXK1ykAD2fQmyBueXm9IjxZbwxp9iuDoXcvWx2hQ6+aPRbSrNFc7f/JiGQ
7Vj/MYUG2SccOICQH3QUOCnU1uwVry82Vj5pH+OiMohMX9iVPjd5QBSYjji6sjbXVtX5saBcaNxx
ZCcpdUDyjBH4asBjNKhhqVX5YuRCS8KphecVfAeuXSw4vbe5+yCxkvLPNxwsVvJF5/ERKmhluSv/
RTD4wi1xqqiTXQ9/Tipr7lElsW1//5lhzc48q3jYPUyL24ogsieiSDEs34K9mPuBuE+AUlqaqs+Y
8YTPuj4hnvx+vxAv4kc1uKZorsq4Rmlg50jmPNn1PYU4CEmyEK/xHOkHHzki8ChqCbb1i9mPbCmQ
6pSKy6Li6dc+skswrYJJZTGJecEgONM13+gSK9U4Qh7CSXvaBTBVxQlDHyKmnrE7ioEQ3f0aMEJQ
W3xWzev+ud/P2KORK2xFNyvmspQRSqVsRph0grbbsjLHJKXm8OittboGP8eq81mCpqIaCs6FlwFU
vdelaMrsSHf4rj8oHwqnYLkIIXcxqsT8H2DCr6VbrCfZclY36W9pEna4WocW14hyfp8og5NOupRm
kIDUPdvKaxq4vAAZ/o26BLGcRsNNwF2AWbjL8oGfRtMsWQZfLVrLf5nIJ2twjPsO87ZU+zawwO4k
7Qn5inGYMcbSB9doRhN5/0FW0gpJZt5SOJw+nnY+gJoHU/ytI13BCeA7jKfhvdbQvQB+H5qpbq8O
W4IgKoriTcwwjg7EMd+UTnBmPTwXaGP96FAQuquxWVxtVYneXX/yeBY3TdIsIRztT4I3Gh93P1FW
jtu8j2WdEzFoOXQaTat9VgB97I0mulcNz4igUmYmWfTLsd0SK27+CPNHOsDfC77ZLbfaTr7YGXq9
Boeo9YM1a947lFZrI/ohWwB1FHWKi383rLO5p9n+Rlu6r7xrwgjMjrC89+tkHXRZCRKvMM7smHRV
OrjI76P0Jq7u0CpNIA6PnEq68mDJTXrzJxLeyAvqfkG9SuY5yr7//5DKvo46eWGmLNxB9iYiQFp0
+QmhYcUt4lVrx5X6fyKPFhipzRk1U4TV7SlyTtbGgf7ogaWTawQLCRpxuKxzRGtF1AXmlBYT+nbe
mpSwizZshbcnL1+VvBAyj9RWDCLXvIIiEGEqpEmPF3DE+pVkdjhr7NTZnF4PvVZbiYXebeERTR39
eLdPB+X8iULJUOk2aj6h5q/kXZ23Pd+0uhOUGEz4g4RC9Z0yzW0yh4F35EjuB0mikaFbhk0AO0rq
vbIm+CnGOUNwMk20Mz2f85yTVgelgvXdYEgFOVNh69hcaFNg47EBmkdAAwF0eMroJ7S72qks92Od
ajAQaLZMztSbOC73hglDCYmaZYZVkMtNfJLnBLfgquajzMOERTCjFS3CJc3qbyviSYqkZZ9p52ru
t5urS9Y8aFs/0ALRaJIbZYZHEuZMWrt/L1y8pnP3oLs9EHeUu/pSQn+SjmhE/fnKr55lPm7dsKaM
0bH1yX5hj072c/iz3DfoQ2cIcbVLZoyQ5foAHWAgOj7bpInaMhmkTmUEiIxAMIcrlygYGTdkAAtP
qKQ0QMhFE31cHqBsHf07KHJ8P9h+sGsCQM4ZKQSv0BUqSQtxuX3vj+8L5svojS+mnMc6FSphCEbe
cIBpvtxFOjA1s+V8wGty6Agn+ZIeZQGkiaVofcDePFxIh88gG6XOY44+I5PztMyN4S3EtGAqDDTM
mkLWDj6IFcuzXDrhMH4SKacTUxRhLh+v/qB0121O9EH2nPNJqcJtQ3QTGodG5FCAi+I9WVSQFayu
Eo1yWAv/wxEJYKGCOgnaTiDrSJjQiWGWFcNdBCVCJLYabqmaRTiYf5Cxnf8CsCNIQiopq4GqjfE3
Cl80PpzkZslL4aVQvox+iDE8KFqwWgs8DgDW+AMIJyIJMYG00rGQn1GTo9WWeuCWnXIMLQfSiOEv
osoP5HQdB6aPmwTJMdayQH6jAt5YUTlk9Df4VcC2L4OnLCZyuR1JeBUaJhDnZtYApS80Z8hdnKu9
T8xHVfoVSadUqsbNjhJmmF43NVOy0w3uBoo6HV+OR6ihqhiuN0zsFYQYNoWFtblm4/rx50RSpMEo
WZaUyV0J/ixg/xCKVRxhtGH7ImzX2TTBdpnonNtezoK1o0hvuS2wZhbtNGBvxezizV9946tw97GQ
9avzV8xIqdBJF5o8W8GAf7BBO9mDWAzk2clSnL/ju7FNG+BrmlgDtFc82NG0XBj8pof+s5r7aKIU
NWx/R7U/Qjsdsyp/T2BgHv9WSohQiyB2t9K5fFPJjgwfDOOhO8F/1rfO3qQ0oqLHcZx2YP6vReIM
zD2pCBjUNH+nFh5SfOEC3BKrbq3Q92Cgl815UgW/8aNlxk2fURJtjl2zAm/XXjXOYNrUgUVsM1Qn
syYeO7ewTDzPL0mM77nJixZAHaQlbse3HGU57QTUh2p8ntNGAL6aItaXAkspNbq8xLW19Nkb+6Rg
qSM1aOu0qsE7v+ds/TT+VB0KunsmcmTOy9HYqUMqzg9Pyz3HDSso15xib/j5iLHmlukvkohi7k3/
0g+D1K69PrhubbrfqFhPrDFRL6V8JNzKfXk46tiLB4/DIHT45cDmnZpc4ponwFhT0GTMNRqOwynL
gZQHzrBo7dwP/tvFPtGgn7zUioKaH6ehx1v/imG15vH7jUi8M7bA6BsAsQkja/CVtoqlIm2SCyEU
Mh89N0mI+XC5O1oJJ4QZ+Om2Y/In9OzlTICOCkQmn1bZ0vMP+kJ6/mqW1Rk/UzRjbmJUvSArrSqK
vgnYIjftexFtleMzxXI1fzJV4LCuYX8a2NJH5PtjMwcuJAq8j/c/4345eg6/amN2xkR+OedpotLF
xgIYfpoD6gzqc7Zze3FegeVC3FYf9exhcbohM0kfvAJiMqDMSwiZs0Xh/F60swkRq37Q4JT4Fda0
GHdU3+VYr0x/ItRmYSBdaxqx1HyW5mizvhNTVe9uJEXUUbXX+Sv0xV1ZRtI0BQsxXusSlphuyKRW
6PZpKcdBlsjgGLlMROJunVs17Wimdu0iNRthlB4tIyOm4NhJSddUAOI8JD7ZKzP4eJ0Vy2/E2kUU
g2wsspexK3z+J+RIo/5jkvfdgUiOGg+kndtR4Lhi8PS3g4HM8lyLED7BWWWeKHB7234dP2BdP5HL
qXRqkiXyKOiXaFpi2dPVsC2GXjB2oBUH9gXD9BpRDpxXdb5v2HXcJ/erxRNWZrN5CXwwyjmSb/N+
4UGTj13tWAgy6a5m+VEndV3bbWKjX7lsVKNH2G2tSBHWK+S+lNkJpiarPeMMYfhzcMlfnQ9/HMJN
tiajQaxt+2Eyef36+c9qDqhj42vRPGle/Mej0LdOnaSzXjb+b8hXalU7Gh3J3p1MlTP2/6arhC3V
Lvq3dE4qAGnI/iVmInC6/Dn6mBeWawTgRDFevo520DokwERqorZpqYtoMnA8miEROrlprp1btQiW
i/ciBf1gSrtPoncMzKwFxVk3RGpkk5betx22Rfyyh4+TDqK6K6znnnggXBhZGsGlxq0MOYbF6mvW
eO80PI5u9f8IyB8SXL6p+LkvSApCSSRsp6Zahy1k7PPNAYX4ryQ1BPEj0mInNB6pNYETpurFo6rC
M3vdaFyhMxjahS344Cs1Abq2kygYAPOL6hM7DYCw9rvGNCgU37jPgDBMBP095/hsavAOrUDxARK3
/2lBvUIaHD7WkE18QkAFT1bENQXSi1fDVufMc6rxWtgsLqdnFeZp4xU3uMhudI5uAZnfHTwbiD26
Y91/Dyr0NAWEplMeRGyRZNtcIAESWUivrgehyhSrwdcUvKioG8uLJcKi0Db3W1UIubWNtgfonVaF
OMYetvYY/czI9TwE/z+n+xxDyMggla2Xb0gQ4x/0wrAjW+nK76VLNCxYt25HNqUR6/Id8YHNfXY8
0iYbdtLkFsxaVKEcJERwOjS67DRKfMSUYWz7Oj4vBi9sjXvhQq6YtZKtClJA4pcXg5UGQ24BVVNU
w/keT2PbB0r/30/g8S1tqSj9fcoav2yq+Dbi4nuuBdkqu71t9i62HXXpeIcpRELtMlNHG52K/Pm0
i9ByY+1lamnLlR2eDbKMyZ7aTYRNJKjFCs/jrcgWTGvDjlrQTgO0L9O+CklF1loNUReqLFgx/19q
vPbzUJViaS2bM72tBxhVa1k0HFesxjE+4Mc/MgNNfVvrYrK+ckFx2DXTjDN6oSmF1cpkVLqxmaID
LwFWaM38Tmyz8ZXo93pLI67/2ve9cFs5+b/DTMwDfy/Kt8nlbNRlAlvZKI4wpjiPvVtIMcy6TvYK
Zpr56xhWA4KbZ5gw3ZcCzxkTKVfuyEUnwGMwZUnz/S82/52SoaOxFnHf8CvK32e3lEEg7RXlGNSP
kVXxc3ln4kXs1/iSOrYyYBDgql2eJmgjnKAFGJSz3xywuZpXXDbSf3tF9bNf1IWLb3OxagjwH0o4
G3UstKFrB4gJRsrdHn04lXdGWd659fd86exe8MCQXbvXur+08j8KHfXTZr8DXVnZA6jWNgOFWZUk
ddZkrEbYRm2t8lUGe+acITE/t4K8Ph+B2hWPbwItH+14Da98N5B7Y7G9UhpPScPkcSxUhUmllEK+
k/0QNVU85YvdMTBeuXZ/RyR1NQcqA+idwQsFx4hTRcwNn2H/07OrNNzbHRXt2oZT3TB8JVOPJ7+6
0s3h2g9Xv6IXXjPEvBL0hL3qxbD3uHX/C0d35+rhT6Ykj6bjVENFtz8ZVCqkOrofHkrEbDti5r64
YyZTC1N+u5GC7OnvObT7Zlubukf5d8COvgr4EJltKtgudiJVr/Upk1kBoDM3g68kH70A9FcrVHxs
vlJC9yeRRvI28Ch3QO+H/BwcvDEL00Ld8T3jXbNOK5HHM934LsGtI+7+yQ0DrNxOtlyJ+of0bP+V
ZjIRFTWJhZUfYun2ul1wMzsRARp3+2v/DSjE0CtF8yUN0he+FDL8BlrfH3mL0vUDjvJdL6ZYIsVr
Gr4NVCoFH1Rct8CkjTN2/2OE/lv17TmOtrNHS8l/ETW/aw1xOJRTqacsMq500cp+Vr9GslT6OzL0
6FX7cJrxoS2pVBSq1GkH+E1lZW1Nz8ua8Kn008BsWdejJrdb1KWgTo7stoqDjvas1XRckR10/HW3
X7x2kOo5t3xzt/aDU9qDoWRM3HCCXDPjwamAG1SotrqVkb4xelDKBnatbUM623NVU9bu57d6/Fn2
dGqc4i29nx8WfB4Ml+pu1M8wrpY3jKhceTBkR7Tryr9gAelotvCpL9UkwpPBoaTCWpliv806wK/P
GbJoj5uCZL733SLlKIRtvcgteySK54q67u3UVfRcPXdVp4dXv/25+6TAx3K/XrhDusnnmwd5vZ2u
Cx+sSOSKuIl9P4VOW8wwdFExBv1jtxM0ZEL3utD0DEJQ+giezd5s6clBpXBDV4VaEP3uwosLR7Pn
L4vK812HkxE6P6A4XcpsyIY34+422C0X6uDxAuKK8jqxFZRpmJFvO0WoJwN1TVWATo0hcasxyXkG
KEtJ9NB4mon4NSCphFsu28oh+sAHhbiQ8nxPFgrDiEIzmKAY40PLiI3FPolTkN8/kamS31ulmt08
fO1M0jPdNocbTZO1wTEP8JCc1ftBxTexncxXeov/vsoMnkK09+si8iQBaGSmspvH4hrLoMTVasnN
yNnhbzW6FebpBdgSllq9yfFGX+bvUuoBvhT+4FsVO6sc8f3Lzgw3A0r05JKVTnfDuJ/fTx2VncQC
SsJlzRAOE99Isttr6JeRYELXKV0nDukfW7fhAnqR3uBDgecTsvGWSOfpYhoy1AkjVb8YLMZaK87m
F57SEGyCr428viWCIosRBbRKLYTXODt74kYZoS6njcVVKx1kiJeKem+OzIzEmBNKf0bxkyYaBwVw
CllunoKNAQpdhv3Aya5Kq/sZGwe48FfGmub8t+iydWDvgAWF6BJA2aEYT72C6tSolTUl9FCmLlXm
V+H54PmpdWIlVtajOjyWSZSrmSL07HFpt0xpPhL40H+glbFibZl+oGGsGg9MUNzfpLuE4jn6bjJG
a+BmocpNx0SRcchDZR3GVAFixskidRnL1CNY14nnH3c007X8E+CpTOo5arSWVDGtz/28diNX9nJP
yfNK8aq7xiEqv/JcjzY6IodJyLl0sCuaFjoLmumLHwH0HZNh4piCodxO436k+1FR0La2MzEkiuPA
4/lKl8aD67RcEXwdcJLrdOEzFTN3x3kD33KqS48W37JXEUsJr/KZlL44pEjyDRrSgh53WS2nk9Mn
HgL/CvXJD/+0CZhn6sgRm6Au0wRZ5HsdhHmWdFbb0pmhiZuWLghfRG+QTBOQNj5up9yrxEILsp8w
pfjcWUsbdD2WsGyC9GZlo+U3NC00GByv0U3/fUlamwh3TyTPv4SYXFOw/8YxpWDUPfy4GBCov05i
fb6gdo/wDMO+qImYVLpHMEjhDTNPzet4gbEEDAVzqQzz3A1EYnCmOzb3DVBAnlQKUd9hzdccazWo
oFOs8LisBoLOL/zmOUIi+Yp+EiqDdcXHRxT2yLeRGVJFu3y+onSj8oQQjj8BLHeJnMbhPQTeb6b2
fasonVuZfRVNeSgrl7wWzNB0EtNl69fwNRIHQOG+wM9K96eAUqhtz16SQ352eUx9NUnHXIhkJJwc
nmUqOx2i6yOsRDi0O9K4aAP/ExfJX6b3Pz1PiJyUVcbx7/TBCfDHfGx13C3uqnfy9VUkixqlBvAb
0ILm082cSDdiF0Z7nN5oS5cEoXpZQF28XIEsYQJzEKcY8UvXrD/OQ/wuGjX8uqANFFZjtygKLnHp
EdMcnxjTbqmrYZr5vdMm1ioSKz9/Fr4U+SRdO4mELekyMwzGKBoZmpGc+kI87gHeSaXIb80bBjzA
lPRllFIh9KTJhWPM7uKZ51Wbn3DdiWqnlvcNN23wgnQOWKWyFkWmXAMS+TrnZVEvLsKsdTLxpxIx
q2l++kiYvM/FDpxX0a1/zQM6Tf9eEjbxg7PKqAfzqqV8j0XmqS0z3GEM8ACcUUd46OvJFoXHaZ3V
wIWqrMa1g+MVvh+Sa17oD3/AyCtjik5NY1t1ZcMu1itE33XXTtVJK+jLrE4gL2yKGKTWHS68szow
FHLAKxRJpLC8n/QVN1pcLxk15UBeaP3U69LAGeFnC8j+LcIz0VmjOLCkFBgx8Uvg3STpryjSCSQZ
khrhJLH4i4fAhWRdRkgDkDNA8i5ChJ4hKrwLPdaAsHg8DY1PPCCfzus8DWQKCXNjXec1lYFFXPHj
cxWo8iNRaBXkpxQL9d9CqZ8KUiMv+b+qeogjk7fl4siCb2EJl6KdPqw/fpAnRVBn2dEqCZ57ozYW
lD2OIkk3GoIV3NYcDbqux5U7WfCchgC1S8+IOe1tuT5KxDF90Wk3vkPjMAUbuWKh2qCYKpUWXTM+
oFfWoPFfwbLRU0pudKsoOLUToJsZWu5OaIowXaYcQ89yfZVAXjyAltBGduXo/Z5BVYofKpaMgBon
nqc1ouSUvBONt71XPaiHhhuo76FGvRk9ViuEJGrGVPTpMw/DWUYkO+xX74bNWl/zCvay9YFCaiLQ
VujsHMCDGGlIqGeCWKtSI9QyM4ljfl9ZBLEhP0CEtDuF9RJ7m+zfJOtG58OT2rP+9s/HbqBacNpX
JYmPb20l/XEhhWSYl21IjNeiopUlCDJ497/FzFpj+j0nIhQ4dtYoMdYPkSMB+S4cWXeTp9YSm9SL
gtxUpaqiWfwLOHANj0AFIg2S2UhhlCuvElnqwHbb00GaYBBmr07uQE985LcCbLauj27/Uf44WdwT
oqiFrXRY49Dim0I0T9D2MphcA5O8gwVEQFm3gbVJcDWaPTjpednirQ26B7Fb3fzk4j+v7NuzxpTT
zFnsqOsdWmD4mQ9Zz4AT3VWRcGv1cwmVpshp9QFDpv87DyvLuHe98LZcleB2V7EQy8rLwmU5901E
FUFdRdYPQm7WsN5OJtr24LirNbYcXF6HN5RBsjVZ62wKeGgU6bnUIC9Jzn6nYAMxuXtSyZMGU4MX
lc1RlgdA16YYe91uRpsjE7oW9SfzWALVOCQssO0nuBJPvBvOK5iPKqiF9P83D17H7RBRKbn3liA2
rS3IShYwiE1tU/vCElvJOqb0F3ybdTbTLyfIfPk61+2mE4fOX8kGx1PgzkfeNrEOBunugQrgvOQe
rCPYxVIdZGM4efh1bBr7Hn0p6nW1L+C2bsqSJQ1KE8/4Gut8n1uO9aSbNWDWSciyPc3PMj7F2HBu
2sFzh+D+c0nwE2882XeUTLgGdb5/8hfUCwlpFCmGurYZFZ8IoXjzDBmA+ocQCsteMS1ORJtHqbjN
VL4C+Be1gJD/rNfV7tOH1psVH28Ds6mDIxaByZOFmujhDRV2Gf7kl48sMpHj5CU0Zjy5RMDLq55i
hrQWxj3vxSiHAiLf/FJeNVh9QEgTrbqpvY3SpCAM0YlNWGHlW2u562ApYbUjvkMVhAzLCCmQKEyA
WFBWqppUumNh5vsVs893riitCe44n+ZSzpxm6Rx60yRKlmjWgao9SxE1v7bfWZNxNP1dlZ/muZzw
UgFNp4MH/jj+7xLgXlQdoqXQ2oIqWSW6jsqgmHytnfOgjX7UrYmwQJ4dVsgwkLUCx/1WvCBVOziu
kt90fkPy6IVFaiimR+BcYt9+kM+fnaRV1AmXfYOq7bPSWcknH+uC6DV+eQWeqMeyl2Vfut/UsZiu
3P8RlLDDnJbEqIp+3LZht+/1g/po8dQS19UV+mKUQP454/GD9CIebuNnsSkYjkLqWq5J1tZJkUR+
+2wwyqUEzoUamRzgqFQhEPk0NzF5YH1NZ6POWkuPcdqkDUDAjWjXTN90oKzNkeTGpulWKdcEExDT
TdLWXPOnkkXX2FbmdoBtzFIQFlPZRq5WylpptJ81gYRDq1HUwRkLYWuBFNYdqL/mE1FHroDc63km
HSxIO0ScT8bvzN6ghjN6bLw0Dwe751GXkQZdsJp/3nggpOxrBHslUvmeLaD128ztfC6HXNcXUssp
B6lw0jaLsoZmvZnfcv9/hGR7xLeGzz3G0JsXVZoGJDoku16f9giiJM092eGvFpYIZ3T1snaj5His
ifuMpHUrM9M2CFur2v10MgGGBkDKHqfXnu2CjpG8ky0C6Rf1gxByysMD9f3b46lt2WFGcqk0uHf+
5yqW8vJ68dx6JIcR5n0MPaUd60uvEPeXF51XbBqOHvpUZToqcVG5v7xORnfhcM/d4fBgJr44JuGK
ZVmEHIFx4P1ZCBZZPLRt7uegFByerphPxrGzHpjeY21iGuE/lIu/a6VGM71fMvFdR3ryOa3t0SRt
EeMpTVCIr+k6SgW8VNn+xSgdDEQmUzaTEZajXKqCnI0xitUtqjfxbtIOmZyh/HntUsf4F/7o23Gb
uyRjPIr+awA6IWiZJ7/q9gX9cVx3kaprmRko1arXCpFFWz0ZBgAuRD7KsbI8Af0JOJmlAJoOMB94
hH+bNig2YZUMksJVtJdd9DcP1CxSTXcjl+/ergJ0CPlkK7ov/VUeAh4uH/OCY4OVeh7hWTnSKf2K
x6yVIAm9Db1D5GMYYJ8Pl6zZJXkx9J5UeSFEthRHnksvHpcYpDpJZq/dB01bu/hR6+Z1WBve+02D
eIWlgpuD6MjbpiJOPMRF1kSa6LoW9+35gFUHrwjwbwDsQurMFhugTQVrDbs0y1DeDxvtkvrmbW1Z
O2Bu5a/N9GJYpsWqWua4Lu0+VDzrMTyDgRfxFLIGDj7vhQcp6vZGvyJLgwNziobjUO2P81O2sH5I
1Ga2h5nJZ23QUII2oUEJWJzZtn2viTsLXnmMkRF/a1xtgcIVAH76b7hsIXhZZuB4vRRb9/O77Njx
Bthii6XXyHJZbUp1/T8PjHCX+la6oCyiQqI/LdwqKH5gejxCyew0GhvcnqzCCS05RPqpEfDoebQ4
galBTFpk2+Xjlx3hHP5xi4UCENrPSHyE38YkhxCBG4S3oEhQJ+9OyUUkwFXTsaov2IuVW+t9hZTh
SaHSUZuF7Mv+NhptFbidspq21skzqoUGfmEVwX65Uhl3VywPfUitd9n89hLPrEjnf/v1vym8WA+X
FBrlg6axNzkFqal/T4aG3hPW/nnGr9K5VosPwn7dOpHP6HexBRJXStsInnE3g8KEnJnLOAHQUKXQ
GvJVzfEn2GO7WIiVUZHjbjzO/z1zf9JneqGegF6AQXQeNz8vbg6wpf97Fypit40p4sR3ZziMIseq
DeNg8twO0tAJ8KBqMW0EeNBxEusaKefXVt9tZZW07Okeuz9vUYjXKtKQ/s8dN0zHhglm8bGVJTOA
Zg8a7JEI3epTrmazSGXpZlh6ZrOt5Vpe4TzYGLhQapT93qpeAxTBNCEj3V7fmF4TXzQk+j4Q3EEh
ooL4uAD5uHYvo5brfIZXUfCDyXyMETXhb24HbY22l4YywbiChI58pbqeZK0g47EaLmfKPHbjAJs7
aB9v25JJq/HDtB3A52CA3OjqSBq4HZZNeckKgbSlv/EkmMoVMF6vBW62O+QQfVd1lzDgXoRNMV7D
tqAx5Ps252EWnJOJBhmTrDtENFeXKmqXUii7ZvKP3uPdLKGrnxVJzvSANEif2L2C3ZR5BUlZKQL/
h2JbQZxGTD+zdfv5K2r6c1V+mxxSQN0wdD4Z9SXAz5xvox1pIq70nFi1oN4BhC1ZCcNBoXgW4kh0
jgr01eom2q9TmaTgPHiCtyAxkgqWOuxvoCzwNOLKz0b0QE3ez82p+EeRlcEUmgzrlmAix65FjstB
uEycfXKWiMCCHhL2WYn781dBlgqvGM5Kty02AEnsV8nYB7jNViueJSmHheDd0psQQee5aZF40YNk
FUtsQYQtSrd1dDkR3VcSCYP3Ti2mMBwTAzm1WjGkqSdXAnJ9kCjlY+uZS6J4wU+K3epzxPGqpcGG
IPSMXr79iY/a/LZ5Ufmbj1xYMfNnW8X/4hnvEIF+GZHQcic8xsOAGKaZb53O2+ueuOn/8BmXhdmi
5RdFT854/6IbxzQ+9vgxDHVTXFo3Dq7AC5I2CU1yo8u/9vbWSzXIpxz2f7IhaTvhew6eh5fEjdP/
HgagptBISwtTWS4OcWTM+LFYiSrLHXSBYY7HGwWPVqm9PnWu3pucUbyR+tSW6iG/MldnwUJYPOms
GxDUUoS/qbVzOrMUUjPPIKgY/eqjhkjtpxvl7344Jhf/TRBo0HPF+CQgSHOBnmKiRb+jFPHuhAXL
F3kxt6migs7GdCctd2SfLh1SGp217JGuV3JNdRTzAbTpqLljwhhc0N95DjLKPZFmxZzZmskxDd1J
0oLcRwOeZ15G0ZTCk84weCnBqLq7GXXDrdp96Y8NyRAtcAS11RDM3l8JxWRxVi3e+MzyWmwH/yS0
St3AhrAhN5qluRn9U2auEf6T6m0eWw1LyutnX8bMkkJg3OwKqaqwCXUaXx3Ol5CTaudTjfIlX883
NNYo9PzaSVprQYeI7yePPbpBfjSfBw3xMojNPeOj5E2rtXGBMFw7SLwqjxeV2gf7l0C5DUJlA2/U
tAjecsOWUPCU2FTUUywzO4bB8Ph+yDKQN0X0iHkDaRfZWIn9v2VSFZRdQfdpwwiW5iWIVr/vovtG
WLJIAadWsTYTp69lOxSIYRjyojgZM+LzFU1+7v/UtVDWU6vNxgQG4cbivIQHmiQN6hAPTnjZG82s
RISSvmGiqJ4F1YAYnm6HDGHP5ByrvdS5mvbsEsnVsX2Wj1+P2iMUHV65N/oVaDOOsiM3Z8IPrJZb
CBj2T05ePhI1JNDV1fkJ/Pu1Y56iw6w1FCX7im5DpV1uKS8ef/ULfqvjIwbery/9PS436OvBGGUZ
YfCYtYOJT9WWgPq4DSyOPnqkgvqNv/ANLfMZxIw9niu0m3F9xg/uBemHDa8BKEsZ2OqHYv4f76QV
lc6s2rjzh78RQkJr/9VdOqVMpgfhBXId4ZK742zfSqJn4RMAUgRMvWrwXzkAJ0VLSFUno/cqkjBT
xK6gZL2S8+IBNSPlJ9xC5vX5yWvDO+ACDEXag+gnVr/mx7LH9SWnPxXCsYpzVRX0HNu3C0ZEh8kk
Gqx7mrVGgFoV+t6sGWvrnyf+mbp7ttuJhtiRoK3KHtWQybRAhAGRoAQNSLKbISxFYn5EOf/IA7WF
72UQ3/vSS6Iog+xG56vBz7BuKMAEyTAXxo37RrTNU/sUWh6VCmv5kYNHRKU1cdi6r5diZyojVn33
HEMAeTrh6uX/0uF8UY/MmS+3AV3/eyLj2Sbrw2FxDRIRSxKhNojyGkJVDL56Do5fdPDN+vaK+ETN
zKJL6HO9wkRhOa4/RkUYzV6kC0+35C5IoB0xnGUthCBQyl/BBfnOmPQI/J5mFxhI+5hyEn8vlCV6
lK/I6LjQFd3ZK0zNLloZ8XIPy0us546IbqMXMz80CSJCoB++UF6Amhc8no/B/ptsahR2xGrA5Iuy
vCV05/PmjJAynTJP4hwXf45GwbM++X3Is8tK33eMke7mFcoh4HWtLeSee/74YAsYfmnFUqt9OVkn
C0DDBFhOLtTa7daHVJ+IHZtii//IS+d/qe6gxbQc3kslxXUGGzMTViz/j1HIG0I5dpn+iyg96zXE
iweSSaVfycWyNVgz9a81xJIf6exg9fKqE8M+HVOQ84qM+h8AAHgP3Cxm6TnaJEVcgtttkVIlarbZ
RbSfzbDl+65oNSoeDGLGQyE67fFeDu5zRXI0ZG5jqMG8mq4ijpiwIJ49N8YhGiRV8mDZbP0C3Rl5
a7CjpuIg8tIMd4v9h2TKNFd0Z8XFEljZq7/DSs3TgyGWcJEH9bJJPQy/npiLk/ovB7JXWAkL0Pe9
d0VpRCBCEsRYMxXFa82an9gejyARD1HuniqF4jxeAOatUPBKQFXJfBzqEirTA53sqMRfgcyQKKhc
+u4WomDa4A/a7m4wCzWrVibLF3G6/9jP2bln8VAayZSZzJith4b2G2tuRecK0UMFjcgH9s1xdotz
detOjCKAgh9bWysk0yPoAXMsyvQ4pOA6ygG3yKDmzozTqaXCprTc95y4Iadp0+sKQkRZcTf58uoe
4Nq0kAUEtT5I8RRZZglXkIKtiMRhZvrRTpW8j3bsmzQ9yDpY8tX84QwK7YKXgGwuozzipZdkyhgV
Z5P8ukFU/VBUUZ+toJEYozHrQlafdeOXkEcCWSrkZyRPgNQl5hH2rPjNC/NSCq7a+wjHrL+fek0L
D1AL7D9YYlyS5zavQFIB31pGS5s0rYVzzfYxbRloY3Xz2CZTpyEsq7SZbbNXT2lEobsOfrwiC9mq
JFb4ea/Hn0SW0SMX2r3TUR9pQiPWDtjzyrMaHq7xc5FyZFlr2JHyLwiYc4l+IMDV7vJFGMpDZ6+G
CkITT2NeRGHR/36AE4T4uDWzc/SVy755amlk0QKv/7bRXKbmGt5gnlg9ioPxZgI5T85+DUgxZ6Yr
q/YZk6QKtKc8s0NCumm9ppVI4RtanYVtzviRHVFBTj9dG/cHl2bW42mfzh+i8uKX9GQpu5FjUE5I
LRIqMxenAHi52/X/W80yRdfZaGb/+2+sivF3l313OtSvgBqGHShK5IcvWX4N/dTeY6derjdgc3dw
BYb4A80ccVjbwUtlFGHPVlr7a5Cqz8v0QDfLTL+8RK2IPgxneg8U89AN5kLr6RpQaXFo3UAGJY8X
OzkYNEhdbZ3h1k/aE4Q6OqFEAUbejiHyMBNqPAP5QWaxB0F5nsxGrrCARhUH7GfDG51NueHFBStG
jOa7ML4CfG7j4dF8EKUo9wg3vxhx72cvuKjTIv+j20E+Rjqd69lEDW9TDbNF/ptslGYgFb4zi6r2
lrs4+nyxP/hmhpy3568eSuxXICR2IC0SoP6hb0xTyOLDW6qG9bzMUhG93lZKxB4L8wka8a1amxkn
iaMSTGUZDo25+cXPAVb9J0V6jm3fjH/wJsENuYxlejUOxQlfOWimkfiWJGdPLlFq6C3BMARDAQtJ
AOTroQwYm5IHUs33VFLI+Q8ZKI9c/iBAyT3ks97WCJwYHLuJOVjR1h1b+MMYfWta+5f4GJh36Vb9
gPfYT9yZRo5+h0lQ1BzOmmPtFg/1+rHbQj6TKLKoFonvz4Ngcu3Ly8rMVQNVY0Oxak9EB70AjI0G
dG5X/u0gc/2qvUjzrnHsz0b0LFYW6gn+wY7QS5qYC1RhGhp1BnHKS1xgMXLUfejS20RfyRaL/RQN
xP67PSX2wcnQGW+lBDBjXttHtjDFakv46uUXbdvasMGcAgWgLcRb/tmFCFKDFj8VIoreu8OCg3xL
7498kP56mdjzA6zbVUGue+t+d5l4hvlJcoatcIGdTclbEpzyvG1Z0kug6qUP0kmEpZisdH0pBEwV
Y5VxWK38wO7MAb16bXmwPJfo9EYbCeo1HoD/KIOme+VywosWnFWC8tpz0vp5+uYvz/ntTV8eVbd1
r7GO/4WTzj0ahnPYD159JA9NCx9nHFNfKxwb5nvckZDYfVuEMpzOZhCv911mOkvnWcfY0unOses4
47kPwFZoOvFjOtK4AfBJIvpfM90ptd0wZqIjyDFeaXdLAXr+GmbRzYN1TQJGxHpM72gFXxyD6sRt
SsZ0Gdpy1+Tave45ojFfEMVb8cRqNdZpr08qcSBx2q3f2aHnQQNRFsqKNHKG3UlHHhgPdIskvYb8
XEdudOOB/WQMekl/FehyTdX1NOO80ONCjLfCv0MAntIyHsHip5oJSViifwc03ro/AHOkiDDREwPA
mG8xtscQGEmD60RFhLEtdHNs8UNiPXcwPJ6iHlwjhk7aLzzX+lMmTwEsehInTKYUkp9u71ihWgDR
0vnSDT19RL+MVO0QhTlTmDbIEQf/dBiCd4lzkPbO5I7ufA8rBpUE8Wb9lHhvzYntPaxwOkJ7swf+
MNImCqQw6wO10vMMKv4y9k88h8Xuel3Dzu9jShDUOH+uYsUwZDTR2N6B3bWYOnwfPHwH/XcnfiT9
pxMvpY8EO0TfILjvBj+9EZCol0l4+ko5oP9cHLmNQcYThD3JdmD/MtS50n+X03XEqWt5UlC0Xtup
j2K6P7fayVupR9rXKpseFKNeoc09zMPbengTKj6hLHpcvSYt4mvWT1ZGsBoeCkPMOMlRhN8Ualqt
73uKtIgwxyUfqO/UNVzISuljmOjpb03REfaLrnP7dEVjgxMIN6oW2UGVxDgnPKPXdRLFWmG5kfDR
pf+KgWkPo68mOXwh5R/zqialdC8YdP+VTUGPkapjcTcTt7VGcLiy8kguEtnP7OfbsFK1hAoxFbXi
7cgC+He9Ig2Ayygepds9aJqF5kDDIw3uBCqqa81S6WE6DTrjELBZ3vbj5N7Qt7fBDZqpjFvPZXVJ
jmbrvLoyvx3OOu93ztbcBQ6ix7mK9+N18QF09eUdyNCqGb7Yzjoo5ABQNzMcTKUXki27kMscRMbN
YFDuUJU3fHxcb5q+UcD1ymTmOQGuzsQaOLn/+O4oLzYdU8N3Yo7OhFX0a0O7JicZyRRi59rkEh/W
v9IY1yGIxfAHS9N9z7fT+sOEEPMmnQqm9dblIPiqJMJPRJnTN2AvqBSdhSiM6R4fnBg+mn4GPaA7
u+aBkgOyBjMxzS2tQP6HeJBoRrDHarFaLO/8rv0f1IfkgqZOr7fLuGSbJB61yZEBdKhb4+P8Havc
6YOVnKHmNh9Z8s9lVeuScpxyixldi4M14mai9DQD0YRXLLdrLlttJ/UIXcHi7QQ/zHexfvoqMhEV
dLQU3M16JQTJOPgbYMQ3J1XAG5lYND2QFUee2LBy/9qc9z8Mk/vy96zxzKhwWkoeEij5+c43Lzup
XUoDwbQLGzCnJBsCn1zg2a30Y4l5EmlTd5TnqWcfAyrPTN8pNkIIpOxqcXw5NK9lGQaaKQuuYY/w
V85JZGe0jHmIvlFjBqV63/viZygmq0Fns36klMZ8ubKDug1AvT4jQhLFEK+sc5KkWjsMp0HjJHR4
mgp4B23qVbg32ktEEZQbOQBrBmJMRM4mRD4aF/LO6+3Sz1OcOHgogkF6y9CFlTDHXkXEGpt76Hyl
kudYOlCebOg/xk7WXvM+J4scJrW3vo/eRA7031+YdK3cZTSbUfxeqd7z8jhvR1GrFhlW0ndJKEFL
Hzykvwod6C+EWgs1T4Fy0Aci877Q10LbckYPoCnmdZjaP7AsJP7pndMD9itojK3PmvkqJEjM952A
q13kpQ7AnHkBdCc2S3Z27YwATJWKITVT9hX7vJ6531RG5MIYSVrnG2LAF5pED1xTpvRopZ6qW2YH
uA1aVWdiy7A2fYsW0+iUoL9eEIDiwxvtk4lNVdCNeIDZAiA/kKcxp6I0r14V1qNYA4Y1yOrp2bv0
kxVHeH5tlJf+NQKbFGvIMSNEg6hzVMI9F6k0W+Qci3OkZ8siD+q+4LzjpCJKh9w7Cx1Q1pg1uQVJ
gMAsCuI5L2X83+CPj28YCeE5qqGm6+JNKRRoyuLk2cC1phXo++Zpys9tqJFB1j58eMNHL/0by+Wr
nFCzy7lwqt6VdLqrDOJXPcNLdsFieQN1B/iNxJh5MQM++a9u0QMG2SXTP0LQDkh43Vvkwn43IYWV
iNtavyahOtsMAP+wtiWjnUPAtQzkiqfarcF8oN2fGuQ10B09/p18TMV405dTtuiZh7DgMVgB01no
7m/x80WR77vGk2JCgCq5fzQqJVbN2EhKeVtcjxkb/O8uGvU9zr8Zq7yeIbzM7FDAoEKhFB2OJrAs
dzLSyN2oqK2vEQuK/WHJuZiAs3NncuVknygysel3hHKyTSuHP3ZbqJhS+z4aZUvDbaZkIgzSyUi8
Pm3myRKXBnmGsee+msJ+se/SUTpIjNw8l9Myh/f7UOz7J9jBs0ERjDXXCgloJMmp9vbAJMeCs9t3
+h29La4MxUOJkkkUdEQb5+hc5VcWUe3E1fBIzh1LdLKIK/2734EnWXCpwjSAFT65YtaygwITmBkn
jToo6+kaaWb7xq9HtXLlhI9Eok3cXRum2HwjT93OUZ7DWmjuhVe4Dj1dxnjvWkIpcT/ft4Qorgrr
XrAegMKEws6xVlGwDUVEm7SkFYsg/+HeFlFshJ525oR/GciGlds04/sMsZAeW0bOv/V+7lHRwoxe
7kfJaEyaU+38WsdZG0wQR+muMFuKmQ2j76SQxH++iWTSVooEJCf6zxhfXi2v2pRx0P2ItOJhYlha
zmRgD+jq5y+ojEf/Jk7vy6b2Cg/5/hqs6met5TeRhNiIUe4moT8eXV/LJ1jhNPpga4IBPj6pMZCe
h7wfjnQEXZVdCTKZMf7XRU6+9f7rP6/W9MzM48zWd5jrR4tFKFalFlDIDaOBy+1OBm4q0nc7QEGE
/BsevdJ1g/B5Zlzcdj8sYW+Y9lbo2Udla2u2LqwB7NiS9CEOukOCvfMdan/0QZkUnfmNNxkxTt5R
bPQ4EaIrel08vBan2HXv4GLkCrBsFmTy5EawTMcRsn2m+vrtghCQvMhKXm6oh1hVWrEjPoUVJUW9
ccLb4qmR0/XqHVS0o+XQumL+QiCJkoHCCFxKIN6ZoReGntubbq1uxRgb8D17/bA1m9CGBemu1YVD
bqIbiXcnV0BOLH8UcExz3n4wNYmsu2bfpO1KfGwZcazE6YTzdJitf48NiaExHFxjhhg8IJY15I0H
C937FJn3vt5eNYK8GqD9/tOnOOnE8Rhhl5mJz6DWuDlrVFhicf9U9SRL1mU0wJokXMu9MIJnRfqf
VaYhiqPReADj1OO0FAODlNlSHCXTfp+RgnXIu8VEHP2LKkamoJW3LdcPuF3tJLnomQWBGbJwOk7g
6Vvnzjfl4bSGmHo5Cfq7ojVsa4u32VSQqSCR7M5ptkt9XNz2r3Ki7sTMOz09z9w9Whah5Kemj/Jz
QYaFTFtm/E9bt3S54OPh7Cl270rsAgCmoVSjWWqWz6SKPCHe5+r5xdWyNoW/wHgZy6foCa62zjjr
MbwHWJnvzGczNeRveYb0e0aq6bU8uRYgIsDiN2x909bdLZ1G3vg35jORiBXPXzMbgGyvxfXXYD+N
RVEbeEOJZDyi84oEkiY9WhiGsM+kLuUYTQrXlz8v1sd6VPUpOnm5r1RW0de07VGiwZuOV1fVarqZ
2GBnUunIwFzb4y0vE6vrxNhgxstQlpaGVhoJ3dWrFcLs6i5SaxhQuf75OraZcw6rPP3kY5ahdrXU
aZGhYRIGm6rs056rnHQCTkbZO6PHJ5r1NIvxFxM9boYeHVWs6SwQNeBJDjRP9LqjqGqH9JTH1tO6
czHaDIZb8K01OJrpqmlXrwRZDi31XtCqJrVFlSr0mK8W1fJcCF9XsLJA+RrF82C/AxT4aB2YX69m
UyYzUxyZN90bQqba6ETJqfuGKVUenV6+IjyATE9IhlqSXmxzx9tNrvRkH0SCnQ0oYUFYCh0czurT
y1KIMXK+/S+YfBbEOq6MZ/HUSnPS2DoxEslGJyLCG0+G7gQkUE0zOuBGgB20aJ5UU3MVF8aRGhUB
onQcOtDCrPBjDhB3M0LuxcMTFF8yc8eHuqDB+0paPyJOOHvGJ4IqDr4U667jVZYQhrP7bajFPWFo
xcmp/faJhO4L8WNsM75tpV2Ry7za7b0su4CRMrByfUcWfcykkljSaJhmiqv6pyNrqDOb9ZLoL2MC
j4gF15Z9pKD0JO9zmxIXEhL/udOJ5qtysu1jG8e8mxdIv9+whN64qtIJb5BXM5kQpj+GSLWtrVZS
EUdAW5ZRSJaLHS8/DhWj1NhPSQpU59LJA1AeIU+flv9xT0+YldcVmAsyxxsRsaeAbZfCuykttX/A
7s0x39OWTX7ESj/N143isCiZkHdabcc3XybHOLPXV5s0e+NxEOL2ac+E6kwOkwLk8weZhHl8J5uk
98nvoNnC/ioEvD/Iiool0C4yUP+Bkd/TibdDa1zVx0IkpwiSjWqbYcKqs49HYt8FQVlObAcmxE0K
Ks1XtRnZ9ZquUlkL83BXUoXRmg272OvBhHAPphUhY2lWjYwzNJP3gqYGvxYLpbLJHEJ8rjXSfmx1
vAq2WWNWhZuDgRdC4CpZKVesvOnjYy6kvil7p2NdMzznZ7uDZS/8iBq7+pDg0rUFHy4DWrhwDfRJ
xEyKYUi3LrGteoM3ObDgAOyhay7X37brD9m/2TdF0WbYQLKEQSYuAZwoZPod/irSOP3Kjtq4uQgg
n6VJrpKICEkNZq6yfFZEIxpDj6ip4x5/8L47XTxEotIzyeDvbfERzYGYeug5QAzWkfmzN2O+NSw1
GMAmDy+z88w5WMhttETq96NHNMo6CI/m7qx9q/UJZdy6EiqgyQDpM5ZzgCSWqLHeSdKWEZ9H/Zll
J46ibzRckEVF8EA3h9X6xIzqYJRAOuym1dDh7QCAtST2tmjQdz6HjO3LSsJM64OH2+VK3LdhWwb+
m2hRjgeqkF6xMwx/O6hg0n7J9f4HjzgtCerBgwJ38/0d7xTvhrhjD4UjCxi6JsolaEHnhfbRbYn+
/l2UnjL9BHk6Fb+GQ3IsJmQQcdAT8WHqfr2i08UG9TbVqc7g9/c18XFvzMACMPyltd6LfZgeRYW0
riEU60FP2Lr1ogXtD96w0YMgssUYi4tWBIDnYfahyxddSwIjFC1SchPcVf7rcwHRGZBYWk5D5opU
hzi7f9E0PoRIb/PnKrJNScsz/ZFpSaSFQMstOAt8e/Bb5+NaqGrYqg5xVaIK97XZfcll4OXvRqx+
q49ufVPEm6gmlJmW4nFrtBwOk6F36v86TUrcLJ68LgKJ9qR8r2FUGKIFJRIpDsxIahv6wGd4lyjJ
kWBriIR8Y8vexp2eEfrvbP8bVl0f/2fRvZo7y2T+awotF1BH522ROBjkWFD3qbYs+dCYoYijQNm1
dgpI17CbIUwLsXXgC0TCT2LNqEthkLabfun4+6fPDFIGnah58bwDCyH5YcdIVpJ61nxTroM1ob29
6jMnb7MWwViWvJUzHt4COO8h3DRyZdClEKyabxFJ3ho2mR813udfA5XE2w9G6UssK7io7CQQWWIk
xdjtrLCj+ZN1/IkIWugy3lIuryGQCmCFZIOWv9VYcDPlJtvBYKS3PDa5E0UNwg9+VY2GCy38hv+j
18vzOnZ52RZ9YL36D7SRUJFoFpKSZdmXnkeF0qTP+mtfKkydc/KK02nXgUIAhT8VuNnzmEXL8a95
V1T33t37hf02k+sf3W50ikClxsrETMrB+jaD197a9E2aMlqTVd9Flc0/swSmrXm634hF7u+d2r5w
KxLSKGVuYw1gBV52xGnj2/Ab5m2VVDpMi0MigIl8z+yIN4TvQT2RArval0PBAJG5tQt/SiBfyh2g
nQO43stu5hVRg7sW5kwDT3dukA8dUjw+lnvYGzzH8ERhRdDFDM3aCi025zk7K9YmzVl21HCFGnsi
ONRaXMSG8fFcWVExW1J+BpX8++2qwrwmiexsETYNrUKMAdvnBaHPvo1xZOuvGJJh0iAojqEcI1wj
4CtugBt+RH+nyJPTeRop9j51fWrD/T19FUH8Iakdsj5wX5rWqD/eA6RTo34IUzYXAl3pTUb2zKBn
n8EUzSaKY/PcbNq/vwa8fHzfhEabW01C+yjpsYM88ay+gR6PdiwZuQInHef3N5Lg5APzZSq2BmyR
VyeIawg+BrR3q3ZIuCwYINmGprV4v1SK45G6BtVUx+TdPBa4SpkhBXvzn9v4knKXaNXIuazlqcYg
GHrqhXdiw54UCW7yeWkjBNZEXeJJeBeV6frBq1JD1S9NXAoSpKftXnhTtNgmX3dUsu5uHFJBB1xi
EX4hUE1XTeZ+z0cjqdFJVubMBrs8tLD4HDkAlGOKlCMMSnsCcs8yOmL/LtiTxAEaZN+V5lgLzcvV
JJAu8fXrsb31uSggF2idxMdRfjaWCrFwUtOI1t4pFJ949iFErjMXWy5ihIQgQl3Puv7IUgQ+8k0s
ihP3bMsrO3/YZubOJaOO2C7pHgmRP5P/Zm8AkozFIY3LDhJip7keebcYQvFvaHVSUbb3XgX8DgOl
1boLYB0tKQTa6mWsQD7q9LplFEOPWMBHTEkbGo3Bvi7HWytUXsj57dThX+HJwhqt40XWZZx1WM/D
U93n1inxyV4r/iYSNah6V4OOeHHk2qTfpybfQMMPxKz/B7HrtJA7F+3xkdqgpf6HR5O4/18FOMnH
PiWi4yFeRKEavHG9Hq+2wtELH0X04u3Sugm4JCcXLadxDd2DsSutHBM8wy7ZA3D5WGGmg3oA3S7Q
fV6uXhqtCTWYIwXOq2OJ0PclJlVzJPbncPG7CChkq9GJtur3uDC+bS9br7IifOCRC44/8Q8TD3o8
9uKyegTbNjH2CQFO8urTWlbRdXL6kMJGRmb2HvwKNZMzZA7twg8GOf60CFyyMmCA+HnxBoE4ZiUy
USTQAYak/NCKUwuoo8ltzYR9ZZNJNJNeJUrvCkhBG2k4fAwQB1ITANXpioKuMQQDkl76Iw2IHuhO
DKoXDidyQ1olMDib5Lb/PlmBc7nc2H3FjhFfsJA4Qn5aeKxRyBPdtFhXuLm1km2m+dM63cB4rBUw
fpzh+CJYHzOoxuLt0Ext0EZT3BxDYZDZw3I3JxYsB54Dk+XfsNwJOn9/GRk+ViYp7bMQ4YrImk6n
+ckGwd8JIRsfEzY6mYE9VuweBNReCUewr9TEilCu67WeL/iNQ6SLdaJ9azxsJoav3mlUE7b/UCp9
OmsKB8/vUFfGJ62Zja/IeVFg5+MFnKyNBSvOyrGv66DCLL4Gmu1c1/h95omgWcYruxa1+PlJze1j
wPig0IgXrMeEbbKsSfnBEusgVVzKaEOE21EZh0zJEhrQOfKB7RBD5kuFYgFm2fS+aavSbOel6r6B
ydeLhh2nr6KvnOuA09iqgFGND8QgG6ssFzm8jL0LqrzGgak10XarwGB2byhpPwVqsm+bH8t8GphX
3aWBlH18b3apSgnSljSr7zwb4Q+GxOWAPgk8xYQyytm297p3rrjCCTGYdJ4YFs7IieT0mEFJHTVD
8Yps7Dnxd+T8Ow0WRLf3aHPZjLIEhn8wgEJhujY8zC56YsfKq/RpvmRSTk7luqjN5v6FphEJtovB
10WZIjJ/nLFamPgSF2CmoLIXHWHI0fHSr8u5sZM2siY55gi1LTFwzRfePWrGILbJl2+7ZGaENqK1
AeUuPzOxnnpyR8OyKbDwDRtpNuR9viDItAeSwCXUrUVgJkq5432TIZ6xmCAIW9I4Ev0lYImKXBh2
x0V0eD5skp3yIP4zdeXAsWiDuOSkyjq8NcUTGS5uif1mpKX8S3H6jWzS8gdEmeDouzjDkj0JMIu5
Mhl6sx2RMJD+XGHJT13ukZGWc+LJnkmo2xT+h98DkisMIBeuV0HBLwj0UX9FNc2L5B7eIssvGsGD
b56Z5D0HSuLvKz/Q+c9DxkoczvWQlHLqtYAODUmMwsClGLzo+CZgRc4/4nBNQUN0D9uH9WhL/TXa
OGWWNsLMNWIpXUuzQdCBb/t/cti4jsCleJmFSLWD/+x08meITwZ9Bvs/kqsuuoVgTbpoYfrpwyfa
lSB9BtyKTRKbLfN5y1p0oDTYTiD6t9hhXKEwuRZmP89gn8BWwSOwfCrqO8n8qJsKMAzHZRDm7A1Z
aXdtAehJ6PtfkKJpSlWXdMezag6TM5CM5Amw8ji5IO3HMufTFb6htKTxXF6eLB1q9CoeqA6BXFGR
XoroG/iQYq7pnbt52Y/u+LshSs9Q9W9yBpj7x82NjqHKrOuwxDustEuqMSdLPeglgTDUnSv+k4MO
+2bTIxo2fNN2HYsB0xTsaZLzBoo8DZC/bzJPOY1RylJnUvSJdouZoUlxDtFpetEeVJxWHcsAXkvj
QTNJid0HvppiQgmK1Zp4WLNiUzTji1C/ykDtGJ8/TqF1uY300dnAyDO9RCPG/viWagonnozV4UsU
I03reQz2f1bmiyrFc51b4j0qK4EuJcrdsyxzMeXth9FDwjIEiL2uUvpjnKu1IUpHOC5m1m72bHpV
9zTbc/e46UUa7gvAqlCEJLQ/rkgBEquxUczlUwk7K0sG5J5JgOniX9l1XQU6vLB17Sr3Wuf3z6+f
yAChydXP28+/sHzDh4IFXBTFsKyZjzp5JMGGZaQ8UrgqSm8VFf79fwQCO6jtpSTzPyoMlpLf04s6
Sx6B80801oR3fDL5dRJWFpOuJEtRgqPxg1uuXyzcjS6k99875ZncILpY1q5fs7bGmnd/TPC+nuZi
DSRY2ehrbLq5LxTB4w5jQLzb2olseqlS89p4GBhQs2CXlOAba5kslQEgxsW3Ryr8NhRs3ANxLDBw
8FIYQ5n8A5Mfj/NvQegV16EB3la2BVUbWDFYvXqd46pRvN23fCBZnXumyNDKnrJNmudvBoq7EOrp
VgAy7pqXI8MwEIgBg4Eh4e2KoEZT4JU1IQsroieZ0bMyEgudRLdwchYMg9107VeFopB44TPOu2ML
wT8XYNrL7mez4h+huEIRABS/oYh/0iBmadhh6vTQW1BB4q3R45h2N8wScdjbbJpbsLz2X/702u1K
WImulDibqmzPW/c2IPyguAPQxHGzVNKm8TrtJSfT1oxrql+RbSvnum3EVPcmgNOO5nPzInOMF++/
nVY0xkd1dX03jc0n1jZ4mOjm3uYDI2IY7qCJzXMaCIgnhX/vl4yFPQGYKt13aooGZRzAJfaKa3BX
rATsWnw6+Lw2AAHKBeFSuDVHLuzfEN6QGkLefltNfmnvaA56hxvieMJPM7yCPJ0N34CdONBNdA6D
ZHBYkQL7k8k9mf8IqjQUl8ceX3K+61UjiFh8k9fRyBQSfQlBjmr5o/VRerpzaLrf0X+qKdrLw8V7
qZuCbFU+mv+9EQfrcxazOQ9fGQzEqN86NXicNyAA+lGVO9UjPeO+D7GU/q7gYv6bebGaZGFGNnFk
L6SMR82jTefPkwrApXvWXVq8QIri5pIBPt+h92ZtB2LsueAotQwvF89bwt+v9hCSSFHWcxE3q/P8
R52xghv/65IK1KsRxxehQyAl0J7u4TMErmgVnJtmTugPh2Hg81GUZ3KlDvgmx2SvxEgnqEe85j0W
sYFIyex4UnBqmqmAS5zGPhn820MoOW+vd5WZCoonafOIhe9dal9KIUM46Xa1Y8Vf5dTvdnpKn782
BC3eP2pN5l+iwr6Pgt2k9hk0Ai5fRYdGxZJgUOyqtLGzKOI9hzllM9auI9274hepcXnl9wGNwU+1
0804mo+BAbo+0JlM+zeXFm3BaPDLSH1KnxWGnsDqlKMpEVr52/laVykSRCUBVCs+lMfKL8bXfjEI
AUT4cbC3KuwdBHsjrayxldZ0aGZt2SjBN7qpaO96NQejMwyl/MsWPVF6gfr1D5PZ/lLqGe4Xt2EI
F1iknUwQRx/adDP5YhvRcLsfgd7qGELvefkDRJ+Vi2VSusvnifVd0m5XylXmji9jfeot1WwZ5AXK
g7ggx76DKu/Fb8lUDl+Cl4ZSJlRqtp0MyUXT1khZjQkxLmyiHK6Fg6Dn2IbYBelJ+n+mZ0H+8PWk
9zMpclkXDbiBJo60Vi6+4awGktkMAUZcijub7OqBDluXfLAQ/fOeIpWZARSB4tvjCUiea0JuCAhm
U6TpvN6zMKZZTGuHbgn/U1IPpOYSC7lbPMlAXOoboW2kdeI0qK7u1pMAmDcN+iJBHwjCe/dIT/0q
E4LaYkuiYb1xp4oQIJCMO2qCHZeWFQ3eq1KfXto3LOW84WbJE3SXxzVeTOAGxT0DcLvVGpsEBu3u
I9npFQIBbG2zth1sieTQL96JFZqNptuy8nad2a0DyFCnElwuo7glMFv11EREn0ZHdsz18UCtMCmT
4z1MIQH6Vc2vRkL/sxgD3i3foUu4hkfK68rlUTbdfk5LR5ipqsBzdKCtVVxfSgjDE0ft8+KlP45H
RAgQ32Dd3qY2SASFwWyJQtFv/TRIXX+2VLofI4WL6hpvff2OA6jajItwm1mIipU+bgNyF0TFRerK
isgznSblxYgIh2L5xDQpck0vRemrZfLY088CxJqYr6NOEDcjvViOMJuzNUWoMC7H52iF+1klcKwf
MLXOASakzjG4w8s8mJAj7583I85tgX5QIcYQh3si+H/++ITJLW1K0DgMHmkXQsU+5YJHMFE2+cXN
Q5GqLlcAB+NudDUoVaZgyQo33MiT8rgflG7nonXdzzgcVB+HrQ+itkHaUAN5/G7AKRY8/IZwfIJM
jZnrsCu5yHvJmB26mVzvsPC3kRnaXoQq48ekeF8NPqd/lYhcQIYlyXLdkS/L1ZWv3ushMahAyWbF
09H8jDbV8k0f5ZAvli5+aG2C+qj6UJhAdfWyEloGUMQ5bHKsso+6UIqfbgxFJMviNRhaLdYYCfIb
iKYR4IvLTB1GrDBIj1+wZ5kZbrN/vDeBe/43pl0mrhMQoD8nrQh8PGAyuev2yieYA2QzD5ffAv0e
L3hmTNWvgIOWg5m2ZWL77vfjtXt3CkWX9rrrIH/C9MKi8g+5EQTfkben1mmT2NWqZqd96ToHLqsV
bIhgJ47qpuxP5X8FXs5hvC7q3uiwq/rqF4Nv7YD8CJWz2aS+ayo2yYDH/jxCg6VuAwTOCiroGN1D
ubudCuzbHjEwHHJf5VGOtBvB0PAuspt/GVAnvVlpW3GQisLdePbFBC5HKVEkcSPrgdc9omKj4xBO
PjYojT3xJeIoXe7R0yGwUjuZ/DVVE5EU+kSd9JufeDZz36IqDD7//FasOQwQGo6RxUHWOPM+pfOw
LZFeB+QBn/QjIioZ8tnIZjg8JYvs5v9DQihwweSeanChiKDs/1fVWw3juWLCvaEwbFnB+p8utumd
X+T8cG9+7WikeVWax8J2U95GYtovdR2vKQcHNWlZjwPlxw0Zfo8o7fyhJ19OnkjAwPNbT2TBsU3R
3Gph3cnlIX2gDRhiZavRnjadKNAhbpMqjZCwcoKEBtN6An57Dfxb8e9PZC0lzymx88Xh0frkR68q
SnqOEEIHOwvIZrIsqH04LUtyKz8QugtVGRlIPkAa/53hqTQ0E2FhHATVqtueYel+dhJDx7u0mxoh
2mu7I0TItpimmMCaIPewZivUQ0GIe2On1/rG/ooELQ3Kpss0yXnw59NiWW8CZyEaUkkI9nZAfMFX
n+OEbqF+/9oXLb/cm8DssZJHlbypcKvrs8PZ5nGvNW2FN+qxKluwSsSiI9iMU+Ec/87m/7IHRsEe
f8bN8dZBxP0KQbH1cW8dh7eoSYejxfQ6j2YoX9tsagTv+cGtEWO2WCYud4YpFVrNoyQ5jZfN897S
ePPBmxZQSlhH7rTl/V9nXuOF8OMfqvsrXqKP2vIV8HVaqucRjfP3JwaM9RUD/l8HaQqtr3JcCrnQ
W+8QnLLARMF1qy18JQjW8tG3BFoIJBub3NFnAv0l/fyIiHz9OAGEi7Xg38JvoVBExycnhHwL3A8y
BgsqqYQtiiWXJpJlWv/97rlQhSmzMPKG/7I9Zsny1UXVyI20Rqu1bkO7SKodJYCx5a4A+qe3ZoYz
6PhXdsRKeI93nY2rqqtTCa2Y8D+2yB9/yoC6EgdiyewRvPkZGG/O+PWe7aFJ2GuJCMXJ7YMNgKUj
0V4bPvddy5lvzp5w/9lOccmHCh0JINQ1yNzWW4i2Q6e5Du7FMmN0djYGI2lmCQbqnYA2hDZeod1N
LSj696lm/bKbvRhIJtbLHbftR+o2btA2IYRt6VK0vQMLm92Y0QxBULYAScgQZmHU5yVBbp/IJ0RH
p33MRLsyH4LXRFaKYkbxj05GJNA0vqoQWa/ai2qPTu2+V/3Z0qH7PP1Z7yg5lpGJzAM1+ypUVf5e
KQipueUQbnhtDtZz547XjwKFecLw+JO4IFYVIw3G6Sx/4uv9HE1uMX0Gk7gmi6jZ7sQsIk/Hciv2
KebXV/o83wdnUmiwDcamJ5wMPu6Mg4tcPzMlFwT6+xKwCAal9l4af06WWB4sOywL6cP9hmREPk2v
Th6qS53YJO4BMxDj8eHNhCx3l8KDgPmMGGrPn9r0XG6PmRFnlUEI08bwPXoe27jmknymuEhHMXQD
8m3RwNjrt2IR0Reu7uEi8b6ZveB89UnKWNmu83gNE5Tgbqe83jOna4R7ufs2oViZNNg/YM3DgWzC
r/y8v4xG7acAMYJcy9VKRav9IjBHaRtGpS/9crDXLd+EEoiI2AC7YGmTBscjwNe9ysxgVaP5qXl1
xJpn66qCFFU01gTzeQSEse9/soBd62G5WZkM1SVTQMk4wUmpMJE2FfieAbe/u7mxJ/y8Fp5sA2VD
MxDSj3qvq2mch8OMpWzcsXT7UWi+HI34KJzA4kHHIXLbgPqemAP0Gpa0yNtopfPUp/9O8cATV8cc
BYLtA/GVtPZG3pPCDkMRIbdTxKftNYWLiMHGySuxsFazMHCyYxE3rUTLYADTA/mX7SJTxQvwZuFp
GSCvkWb24JkOuFu3wULEfofsx2nO5E43jZ5PcX/bLCqmhIwj0m3b1MBxq6yVBssoTA9RYy7cSPem
hmfRlYS9TBetjK5udaHZ/aoJN1S3R557S4QY8YAcS0bpUR03QxgwXXl9b4YfaAIOXH+8CD9kM11r
iMG+oCh3osQ4FaKrNclBLpL788PoWK5FUQGf1boexXb9OcHfidB83Lh//VXur0/HDUm5UcslH+qj
6xhZM6gAPtKzjOF87/GbyD1JkM4F7tP0FTsocOfxmbe1Q53/BXNSV0DB4R2JazOoGs4D8onGI9Dg
RY1QVgsV7nhueCjA9ioqSx/WzR4xtejbebknH/UMTAKO8/rIdwUs3O0k5ZTKIdsvuEY7uozh0IMv
iG9ZO7SqdvShGZj4yj/zMbRA8lc3FYu8TYX2j7/mPaUvq4DmoOPxE2eJstOsp9BLrxY/rM4m0xfu
lKv6OACiddr8QcPeLpkWRPPOY8AX+Rpj7vNZlgUXwgRUfMda/jfkn7c/6z14UXP6frOt+3VSIrwp
F/RzfnmvtRUYc4DhvY83KiMvC2j9wr3+j42RZyjvxALMkWOr6FQki8GiHxCgaDD+0lqVaDJmeETs
e0/224ytsBQX7r+gMTUHzim9aaw1vbp68ibUeYFdCocOAJOSaaJq/ZDQZNV2aEoCa1BiIaTZPuDZ
USADbu5E83pfQh4oupLtIiKqoMSk8DHqEdDIPBelUaTYnSHFc6ZmqaDknMdvpNEIShFiDAgIjjz0
oYVAO3QrhbOFsFFoQRaB0/nW3dDbMZbLxlV3/gwRnaXbXZ7nrKRTHZSJ558dKAqPs3IiGBvbfuQq
GvWdrCEfZFei3gVdsDbQF3K3RG42C4+Rv1NfzSWdnZnIUwmyR0Beavo53tegAvhkG6RwUqETUhLV
nT/H1eyJhnWCnOp1hZbrZ3EkIZSBsDOq+u5rN90g8PROcmW/UZgiuSMrsuSDMNoIcTHF6pEGkAA5
AuRIuVb+y4lBCV6YiF4hf0GcrGtpC04tl1xVbRD7R/EevwRzivxZcx/5C0m5FHKezdgBm+G4ipBn
Emh1TjfKWaEWrBIC5CsC8WWpeBBTU6B0RZeXfo/SHFNr3j2WdIRktgWslNvSXKl8rZsH+lV/5Ec+
+DjpUfNm3G1Ut6rVpqCeyX2CR0/t8YDoTj66mF0IjSkJqiljdpgA9+bL44l96HALfageAEtIyy6T
v5I7Rbo4MuYIHSxUOp+AVpR1pRrWx6uoZb+n9sz75E7zlLEg3R75vd+IMa2VHfSWYpJCJtDdy7n4
c+TzoQYGVfGgWswIKskXoHuhaV5f/z1kIzuU1N2ojJxCp0JFFZzSTVJdSGsjQCjM+259sy9vGh4m
NHJRMiS/LJD8QQSBp+8hQ8jErrHU+FjDyL+7jKyz8pWSq4tDDDn8sgwarJ2ZeWtv4GX9nTQkf97R
0WnopO6iGJylP1PKN2SKa5Ygj7p2Xp25oRoIdj8bhui2WRT57DmEg+mIewGVUggNimxR/jVWPje6
3NMOacuxQdQaDAl/X+AsbU9m0EQ/c7mYdqWROrv9olEYR9yLBahfQT1F9LxTRxkvYsdBnL5V4c4n
pYxltTn/4CLisI6Ed/gKHGf062i7zDyno5nHKMP5Uxd5Zqc5LBUR3gHiRXc/D7r+fvE0dmKltkqO
6DWwcApvuTfCKrlmZ92+ha2uFICtJVxEpOfxdl9Hlj1EroimkringZMA3vM1bvynnlAucpRmvL7O
Dc/kjVZPi85VFX0OKEcfpj+1K7JlWn//X/QEi3n+UpfFmCxPa4EBpDtUr30UAiTWudmtYA4Jkg6b
tY1XSjVyC+ZsIvlfP33zyfi7P9BA/O8+Y3MjQ7KIxVIm/9fA8JOETzgD7amCJ2bsn0y5ABbzIKO9
Y0V9Fe6PNqu06knsRma3DZD79yO3mSJfuAOKVZ/utz5JBi8jfuAWnhF3GwlBB18qDcR76uHAxyAS
cq0NtSsPuTybuu8cT4/fP79xls96O3kN9yBuBYQSYIE7PPbq4DCOeWW28JWPMBu7xOAbG6zOYmaQ
fPmLlxUfcSYkJjZ64BmtSbnYXrilnlh+8zq6uUL5t7+BLt48WRqjArl0kwF0ax1n4m5HfgBeLkEg
DNJSXuEOq3LiM0wgWozA44H3M71A2Ui6zLMvamwrlGKBjQ1bIdRBIRR4HxZJD8Cz9JYmK41jVDXZ
TQdzKw9T5I4OpcjePaPTedGPVCdBHIutIVIa4i1rQy6R58XXCEVv8CQ9vtLOjdg4KHcX+Wu/F9MS
u2dy/TMN7d87IFFPpbRo6aPwYQOXu8fEZ+Ri3fWRSvST60El09a8zdt6ad1KPtuk7qXGaXdDiGLg
b7E56bGhiEQwOXbgUlokPr6PCIu1p2CWX9M55aylgHtvjKFpx6QYWz8NJ5LlrvFmwgAEwjT1WwW/
oFWksuWaCauG5gCJBjllOCo/C1fphrCXZMQMCaU/Ljh6qDaw7Z6Nts8bgfAqX9ISrXu9TVvQIISU
l+WKTRynMF/twQVaqz/ujoXjuy+pVlDv6ZYrhHj1IFiGqnvudyLKzfh+OpAI5SIc7PSz9o0zzl4X
mCxdmu+08/aZ+YC8u1n5CLWXZTA2vvlHdDLmi7fLfFtllh8d3ycRPmJGuUq/47RuX9etzcULHkSM
94jertywe0KYJDj7dLmpKaV6F5FvcRp7BZS7YySp5V/q7hM/Q46ZLwMuxEyJGBQ5q9CNRJVbCGKU
fL9jBBzmF6GQE6zfTv/wBE7fkTqN+Mw57ED9Wt/RvGMv0cDbtFEBda7lDZ1Qcxqj6maUAObWMMJ+
MBabaIg6TRiAIp1oeHookb7je5EBVSwjNBWt2zpTm0oqu3u2o+rGO/wns/J7dta89hcfnmoVeON8
5r1CopaQyS4GkDRTcAhJ45hVgy/hGpMerVL/h8xOhqmqDfXyRwUslngrQHun1CHgXEkBVvPe5vWV
moxwS7i/Nlnn3C2B8bZOiLlQiHMRstbQD9J8R2VXLMyG1C+u4Lz3Zmk3uzt25G2QTFrqw5vADVnk
LBPGTz6zGT5gQAe7OQ2GWudFXrvj2bLzFmzp/1la4Ijon0mNk0LQoEMNeBqxmmPuMSukA6aFCgI9
0Gu7/PLu/1psZ+49vDne9H9GCPDQnrStZKKr8H4tpCCY24qqAuTRSIzUL5kDlZH6ot6fmU25cHUm
boFv9UDcsgSFGtODK7oi3IWHi5tTRG4e/ny6CIW2ZDkEhL8rGWhVYJWaeOgUD3oT8i3m4dZ2fMmr
tuCABCb+1ntMI9MNgJWUWCYeiz7zEioHIfWa2QgoYCwNTS4CP0BW/VaFj5xSjzAFctMZtaAm/8Cf
cw9tbatAecFCVdMWBjKX2Cbs9+6MdPQ95Hhr2nleJWLv3L+9KmG/c5bTkN/LdHgd3Yd8Syoc+qyh
szt5vxsimwIfl0uZIe7JYzYNwPmoquI/uap13mS2J0jdrgadpjAtlhnAHxROXRYlBvUWPPWaoMYk
QdEDXKpg/1Uwxlyhns9Y8O3IK2vueA3RcnzAl7OlVwLtsGlX+QCk2WOrWKE7GiIMPeJ9Or60Fh+n
IuBNmF/XVbA9iuJhQD9iRQKhoAsCBeU+b+zwFx6bfxzB4SrSr+NFYqNLPcwq9hyWIrZbEe5dpNja
/Filt+EgkA7fAKvZK92Al4iiUGC+mj9q0xrMLXoECdXPUFMW6Q+gwr7xyEQYED7b0ujpRt+6mMdl
7fkaG3SzXJTv1F9IFvvCmZCmUHbxAlce8c8PzKdaCbHFtseyRmlfDxT7948MSVxIAlfkwffHNpRH
vfLf8AcEbZ1hSpMx18LnrX2XMsGAY95SIJbGulhfDAgyiJFGrK05Xz6bkFgt764B8U2gZ4usrDXw
YR7J0nSdBEhKazV2J15vvSdyjuykKwpTTVGK/9cvyemu4pLtoWqZWirG1xm6P5Qo8WReMPkWHWpG
6rMjj2L+wMFfOcq7sKjN1EFjoBSv64jPi/4yu4WkRK7+rVyeuu+AaoQgUeRHOJj0sDHaAT/xDu2S
ItVXrn5zPYyLnLratK3oAoo6VmcChGR80M0AnOnZhJ031HT6YSEieRLpIKatutTGihsTA4bqrGHS
GT2VeThvj1+xi+aJ8nBe0hRBfRwnH9CVKpmnDlQ0PD2Vh7EvgcxGVSfuJycxy7BNnVYmP6SZamPJ
MTTguzxq2dodHhYUgQ72kA2ebn6I5t6B3tQCWCFGPloXekVgO7A2If9030vL7l2PPU5MMop2BtEM
Ny1vzSo84l1CC8vkVBgN/f3AlOuXZ0KVg4KMfoiJIv81U04QCwnQxmwlLRAk8HksQVICiwl5GnU6
FgyHX8495W0yAPDrD5EjxIu0Pei4NV4z49vV2TxcIQhXVve6vfqTTnl13mBfShjDgMdYtsnFipK5
g0UQvNBIpdZwY6MYZEMcPQ/WwugUSr07rYpG73B90yiz5Ad2TGO6f1CQfwd1j1cEsRuM8vE48E8I
ItP3k2ngzSvHSt7ot4sR3KdSJmvfdDSUxcJ9kczGfw/Dujrzwg1bI7ooTWBcG1ny8Q+aZCXbdufP
IN7TmmdeyJZjtxMZILMXds6eoKF2PWVARVzihaK95C9YVIuy0I85khcF5OKXg0pFus6c+8JMrHVS
KI6QHwnKz4yFDz31IW7/JtiUb/aU7u6I5HBmeaU4Ru1d3TJUGhlbSXd6mcMtECxxyr4FdseeMrMY
0Vn+ueiHlfQ0FJY5V/m28mef/o/Y2KtMmohNye84fwn2/zf4w0W/6kNRWp/NRJ5jqXQ2OlYfwVIA
FS+1CI9aoOaQG5D8/REhrVqTgAwFvv7/cbF/wvT/qtKUErRpuVWNW4jI6yAopTIY6fs/LqKCvNyA
TcoF4QTc/CypWz3bAx+3Iv1ug7TugMkag/Ujam3gzQKg385NuV4+DNBNZNv7l3loVwcN1Yc3EHFE
Ej2DLw4IK9FXX9jgM1UABxDw4r7Wkl3UtekK0qKg2RKYD5PcqAD948Ds86m5NzWFYo6HDrq1Ms6B
PBVaYALy+8M6HlsxK9xgwVP89QcWIDZFjwzvLwdJKV9nKbfKt14Apzp+8YlkNNs3nzIABuXhiKiI
b1DSung/KDyExZvKys2Nk/4tUQ1E5QaXfbhwGuxztlu+Mi1XOwSjBqUUpxu3lnkvPVZ97FaAnVPP
WOn15mF6/7Dxl7rDJKXuv3qC3LnLVBciMlJ/3mY59ZSArcwYtrap26R7jEPoZHc/Ln/6Ulxg6Mvs
NJWdivWpY7aNNxuCaNz16ZsLa+BLtY4FurhDNj7HdPUuL3TnpPMD/fS4YrihIzwCVBJeChScbWy5
t/N2hJz1xDJNd/ZfpT+Ow3Om7OB1C4sIgTG0vjPyjjtP8d9PGrxmwAripX15iRNHfVgEdEmgoZi3
awibDzjGk/7CEcBNnhTG+W64HDo0tEz9tov/U7TbGtoCd/WiUBEjmXvkR9LtcS9ui9ZqxPcnheRc
gp2wgeCHfiP8f6IBvy/tQXA3f4sIRSZiZMPjmpDm1ZkwZq/FXiC3vhyxJg6lcLr1MR82ugpLqvXC
Hm4/5hEh6IlXS3bzn5dsG/a1qt7e+2KxOD3hJqrP7oGo1mevXsw+G8vv9M7Y6BnL5TnrQPbexT1m
aJvff2Rkwp8/ZwMMiJw6Ee97HQzV3jESc0IwKW3X1N6xU61uVI8XN0M/qG+sQqJRHnT86La7XK4p
5SzD8Q+V9jDF3FJrPB8lcE3HX1iQ0aSN1D8ljQKaJXisYwQKzPwaX8USuqUtnGlOf80f4i9IoVUU
M55+h1R9e+Cny4uabdGmqaVbKfONLAuW39SKxjN0FMB0LdH1U3Blee5dhpvfnYPa3Rig1QyNZKnL
Rc3T539pr6f2OQ9TCG1ZionYMTkXfC/iDlM9Xpe40Sc5ujtMi3hEtuhu5uvEU63UIkb3JzlQ6f92
83P2aMPo9Rjw0kK+csxGl5lmFJbgADhUWuzlbvlUi4G91p/FNHn65yCiYgVotKqyxCKOOngy04Lr
OaI2tf8nx9LM56sm30QOR/QInigW7Hog5TGYcjedBgJlBHLfY7ifuEIXL1kOl/Y79uKNuMR4L5EY
zI2RMUf/9VOHd6nWHyqcLs0qiroFB1HWxTRJ+BK39j8bQ+lVWefRqADbyZp3HYHttp/DKSKlvMlw
HtJUbN/IKc6KAiPr2ohnAmggwW2u0aTfOOp44qbnG4efQvvVjyMjEp2Gz9a7CQ+6WtI9xKqlLz7q
5MGp9dlZ+eiAinsPj4Cd/z043jGdJQXgzFd+Y6Tw1NG9EoRPhPCV5tAyXGdb3/PUb+hsB4vNA1Ai
Q5nUibwln1/dO/8gGqDHaHEYcdy4/DRNrNmaBqWLBZdibZ/AaTmXDUlph8Gvo7SEgIJR4DoNuwPl
H5zXl+33RYPclcDXx+Ss54XVpr9m+oI6Zq75zmsCiFSimLMf9cloKQdG2DxkNIfaiLl8rDeU+qmo
yBLW2VOpZN9oXAbxIY4Y46XDYM3PefC00rYQBCZ9yHlper0aPor9dsjCDwncK3iRjSoiW7YpRgqj
bZRq94AkKIx/3KB7srnz54QV/G9UvfMcgDReYPrg6C8l/meDsNovkIT+uIw8moCA/zq+E4iUbK63
DY1+ffh4urSCzaBqNObvo58BTEbcdp5Kpvt1LYWIWWy3FsnrSOcy27/RLMLPxq96GkqzZ7RPmYAs
mW7QxNsNRHFcDSiF7nCJJbRNCw3rP/03V4wqt+bBToPwkTLdlEn1E7HIzXSRG4tw4rRTKSP2MRFx
Yyece1I3Ldm6x3q6uVQpq2cSlZpdLZ/hkZgOZKYb3xTNWyttre1F1HhXiYE+I2iVWrCPIytShtl0
4x+eO0ca+jWTD7l5cB2b5WJg10HjPjzY5Qrjb+IAZZoWEB7xZMV6Mr3aN781wyKGvWnAtTrgghtR
nM5BJGuPrvDLwViFA34JXcwb4p3oO/S0hLfKKENKcccxPl0mYNWjQ4ULOdBvLcd/3QPc8ERSAGNH
vokDpvIGuMZirw8Eua5ze21A9CUwbLV+bUDrwgMDJBt/ES90gUQ+tKxc/55Tm9qSLTBcLrCGajYk
APkm7FIS/boqhOE8uBiYMybi01k9ioQWWZoKGcV91WzY/HssawodG6mQr2/GRcrvWypeemBKmJsr
iezVTN9fHCczxI1RMvY1Ofcr1Vi5rMWrNTbxlDi02YlbEqnID0WtgiUCzuUbM0cTnQ3I5am5VTPq
J4mPc6zigpSVjsl1aQOdW83LcYdxzRwu3WQBrR94DBWZhfio4ryv8vSCPC743AOHVUAwvc7O6b/R
D7OyEhD95Y5LM6oiEQNsnZnhVrccMk/AjUzXJIzLKAJqwYlA6kSqeKWiT0a+zb81/MaBsuNt0mgm
ZlBBkoT1K+ECNNeLngl+WisLd3uJbjx9hvTkjXAoMvWZBKRxTawsOuaRkhHoG1ICH/x2XUkAKk7D
/KVlv7Ql+l/9V3XqE5X3CUTda/lY3VVW2UE3oKzdcgZr3TTp1d3CwaC5m+07zYKNeO81c/8WnJXe
0Cqov3ZEpMv1xj82zNIHkXftT9J6Bajuk/oEjPZx3Dh+IQRe71zWvpECcGhAPOrZ0aG6iSIPD98T
kTWM5hrQjhbbUNVz4HY6J5LcFjUh8IrXn5bZ+lyILFJ7y/SjY1umkfI5Palhq3NUv1BpOjlTcqCH
MagmEVvs+4meH591ph83yaqd4qoxxo1luRhZV1GDWdzWPrPNEUbBU6EfYhB7gDdGH1BwYk5wsXOE
S28Aak0djWo+Ljqc2kSIbl75eNfLLb9gmjocohseO6Xti31TAkkytXxTjFo9I0hpFbpNa2euNL/9
LP+/umO7eI27cQfSlxpTFznVamUS8iVT6RfMVf8qRhKVHC88x0GsZ7fZwPvxWpe81kh+td5VLLBr
bik41ZVE39OY0Eg0PQmhTBYX511dW4K7nlPlG840W7FcOx1s/9UWPUI5Dn/udJ5tq99RPAkeHSfl
IbKQpoBXR1lVczDKsEo3+wx0/KIbk6QJWBD8sHzhM9Vs5FVxR6LO1zUQFTlMDXksiIzQXkQE4VkP
vKxT4a82C6TEQdhBplKiUDrjyk+vUgDF25nYfABrl9EdKm+fxtwkR9qE+jEVpVj6RsWlHA1f8evV
V1fC2RuoHGgwPB3YUrMoeV6nQ3R5Kxp4m3Xbxr9uFqUvTIzJdT+fI/MLF591Aprjph9WKuVZXRfp
9nlFvmFZieAFSP8aN4ydvIDpnYFCw7CVZQ8TRx/uXiJnESE3Wk8eu5FRnQeYswEqMkrRD6d1kWUx
8Bwx/fY0vyniQVv+105ZaJ3D77wevcEFfymByD/Ud0hE0t+M3ZA6bLUiLhTZZxObf+iXMu0e/kJx
lZEyoODitKwZaqcZefMM/CF5zV+/CGwAgUg7Cv7VYw3b/WSExLO69e4PPNTz6ZCvbXrHfDyUqTNh
xHP0x5fvmMZUHsynZVPRhFkp6i+YQeleSfL41/rebJ4fN4SL0wk9nJE8Jqd0DesWZEXMV50iZ0tW
UosecigRi07VFIjq/EJCpVGmn4GbqLloLYjM7xC9wu0+K0RX8kMR5cI2ZnX9y362x+H7dbfW92HH
TnunZzz/1kvQW2CdMJZ9wawnoOI5h11PV+Efe6ulJ8lkvB/3Rwr1lXuqw/oPr7z90LMDDWgJz5Zw
zoWWhYKqSZ3WjIEnwPDkjK8e0XZhnL6jYo9O82Ek1tq+KL4XvbgDYjNrdRSoBu5tz2efXVJxwOPq
gVFOoctZJn9GAmxdYUahYbsvag0io/rVFh6jLkA1cmgrqS1R33mbhSv6Oxyarl1aaCIHLcxiVrnv
8ETZe+zUqZqW/lSh/k4YoZF1uW2Ib8pme/05/ZWnUKcqhnWJD+LbW7HkqqI2elEUzzWwP3U/833H
5UrpxmIma/AV5bL62q0tS3VD5U3zUtDbDrN7qCDCKQDA3rF5Dqj1mLWwPE1h0GWazqsg17GpIJQT
N6422iK/8TqKP8fPloB47whMAHb8ZRhPPWGFxQ060oxiwaOhXAlWAcaknO42yGIeE42W21DzfMgs
lAT9TIS3FHMbLHQAThqW/BhYN/6ppXgKWFf1CjT6nsLgDuIIgSWcQvAg3V97klx8e0PpTmde19lK
Um+QtJgy10rQFVnvUUVGyiHiNn91CMgIN3UTZr9CVIWhoQLbv2ZuhCDoVqJIO8cKHIpCKwbL7nR4
snOoNfceNp7tBycMLycGo1xPuxbquYRUygsTBlgdIbZqNUMmwxAbgQ9kc/G1EXKONg5ANDujoD2h
9f/06Uz9KJa5j4ZM1zVc90FHmFXMTWCYwA/S0n0P6Yqxca+sm8KfodknadIKtRI9I6A4Sy/sNMtQ
/8A8KopLzmkni9h+DX2cdcIpkRVqdTykXtUp2ABcunHlldIK4oT1UQAQzkslVUYnmlTrDqrdSRLa
wbWozf8PRdMEBqKV9AX3W8aIt1EvIW+WCCefCIPxlb4eE1m8chNXQhPAeNES9nryVmZ63bx9UbNO
HBjeeDnZN3faqZubqDw2VZ+UVs3BR7Trr/us56Y6gHeLJYB6gPqUm9BKJXi/SjDUOj4HNXsMf7ui
WUX03llmaf8YaR0rdJkfotYCbubjMCIK8stKqINQgF4fWalSumv32nfd+E5e66G1u+JOQwDhCDc1
+JDhV4uuDjzOXvFHIs2ssZGvJMUNqSq/OdUpVQ1u5E4PV4vhu32I+Y9qswu1DSC4ueUzGlGbh7n+
3APv9KG/1onu89y3M3YNyEQ8Ihdx2TeeFN9jJ2YbZvfnO9wqkDWlI9YLr/+OTlDqtV8SVRfvVu9s
IrNyUqgjLdnyKacDk4xVpHZ9FKZk6G+0VTVT55kkf2icrnVUGaZWFiEh8sB6eyz9DDA9cWnuBZBn
3pZf5e7a1vI7f+gsKOF/LKkPSZ/v799oM0anWb/1XI18Cdo47IeAsZRrf/tt/vhz/bSBmO9TcODl
CxGED46lxl43N0PqrlKA4RBbnxkbEvGPBVAmaliHeU9tVowu1JPeeveRKNhDhpWJd0BgNJpXU+jQ
tjfLxpLJjRLhtB1PxlM1EayuFErMY/lbtIitwgVVRRfehJRCLkry6NQ1gIfbBF5W+1F2fTwMeiMU
G90YtxMr7o+TNC5E1YbckPoXhKjBgUyb7dfu9daV1beU08YrLcCnXDIMej7jtwaSRaqmWWnWLLr+
+Qz76jQRkTCzTZRlTUIv/EHy9AZ2AO6blhSlU81zHSL+mhGhThIrT4D07Sn/vbuCJYOKhmbHn2lc
SkjpWsMAGHanl/Aut5wlJ1EszPW8dGdr2S/mGDevQbRyI4O5FA4E5DnO5/0c/zfmzGFxhO6eO2KU
4MvR9fXTLwKvczCAeF3DwzTZ+GEqR04Fb6y8E42GBC5v9klLP5r/ngbl+6kXXO/bQ0oonQ3yRWYC
bbANDBLcq8ISjW8nA/v9aG5GCPj5gfj4/qk7FNhCiq1Z6eYuV81uEz5K/AnsdV4imItDqJf5dUkl
P4nEMkteGPAkQ+sOf8o0zypr1W2eI+5bDkw9Pa+a5+P1UBylvejxkVs9o3iOtsC5GzWtfHSkg/0E
bmUkESuYRakVaTJN5TEMtRNYZ2Q87Rc6bty+VYE7QB8bHqVJoecjoNQbJj1R3bt2piy6V0AQCAqb
yVFdRK1aW2pe3QkC4KD9V5/mosuCypDFo8VpsfyLV9JXJJofqvJMZqfOBNlZNnyxJHWlexN1xidA
rldFDUyAeZx4xcZm1DfGwe0GkP9yKvciRdGrCj2AqlPgYcemqw6wb8gVauzGbw/5AR3GnQHXcZ4N
cWDh9/Pz6gzQpIop5KbMyrUhur5rTcLRlvfui297K5t62Wcka3uj3XqsWVltFtOb91+INHLrKClc
bM+roZ19Ux53nZ0VQ/lV5mYFELTQRJFcIRiRi3s4F/xnSKfJF4QNw2qUBD1uUTleR5M708I3QIAh
iNESn88C2qJd9SCEpo3Gw3c05u2SYhJttyRbLK7gttxucgUgRhmhg6smSTN3IMbuBhaaq1bKO+Hk
gMJ4C+JHO46punYyVWTZmcVflix7UaATk67ADMclAtRXIGZGT8BHr3gAA1yGYZQqoSySxu0SZJnZ
sXCqojYNvgwzvPphSjy0Vg0rRHeuvMCAPYGaHuz7/tez9YjW97+pg4tYVAtYHK2EO9AX/KF4pqjr
3icYX6bHTjkwsVr91dax85uX3xqMn48eS0kjNuWCBlG29WT6jYs6MSn+ZR1n51U6kRWIC5iSxwey
bvMkQuhpZUba63tTaZVLf+GB89GPFh+txBkQCk8pRD2LL2dk+TgXvwR9xk3hf9Ejt4LYgJMny7y0
pNh2IxsLgdFVetpqFZ3Mkn2UUp4384/hEGr0lou0dvC3vfduBnW7/5rTBMkJG6Pk9Lrxynd562es
2T5LzY2cgMDZUZKYJ9HN0L1eDBuNYhihYGQX6nMbQU/4nzrbgho0cqlOis7Sm7xN9K6Kl9i0ySE/
cwLgUHGygKH+ZEq3b5xCvC/MbuPjpN/KXrlX1JQw8WoUp5NadbDlu2v0LKkNmrkhbNkmGTwrj5rs
lRalq2c/6FXySe2wMhqqUyxVGLE0ommNudpIAuXxSooW1Kbx8eWWoVbuTbulGqPdtjz7IxxEvdQ5
hZXUpRN9wIxNuU3NQF/O7Bp4CFo15RwQwCO+4HY0oQtWzYfHQ78Tc+N4XlIbvl0vR8kiceUzBzTX
SxvlaNRn9syOdmochPR06pdo3nOr4N3+YsEI+oDFC7/ME+/DMzxK2iJ1s2reHSuGj5190nizgwed
10DuqgC/5B8UsobcYTJWU9o4FX8g4kkB5LthecROvDdIKw00Sd9Us3qZPdDYyCfUU78olfFKVdE5
Y1XmNbbtRV34qapGhf2RBqpvn31F6UZgfYGhrSknlS0U8iw+hBBJ3ycpQ3InsmI5nt0JsAFI4kXi
rr6Bx+aWeXEn0HkSrPEucSK6ccIn3AkwIQEE/NOsv5g7M7+cPU72+BIGBpnx+wQEJtl2oLPQvc8o
ohj1+R1dTFbXOgl1rm12+tBFcqwsYXHBJly+jJSH3ttespFBwW5kHh1jsOJoDVfiJCu2BEXXsxnM
toLSTM7hKDEzIER5Vc2pps+pxk1nJbqNHkA5ne8iRFoTios3YPM9q3GMMRK+BLsJ2iz+zBj6j5hB
txYKrL/v7GGpD/vaWnndQ3HK62gOyPNJmjUiaqE5xZR+U7FwDYUOZ6awDTtnicluRuY/2Tg/zrJF
R0thKOGXGHu9EAd7JtnSDoQtbxbd3Ay4KuSx8uy4L+x7vdGrPgQuUygcBLJXzvXSWS5FFwJdDyrR
WurdgmuZrZpOHBcJ5Ic3+OjRcYYSZsaO6C3mwiveCc8WYByQx/PsUnzjx1LzhSctFG/T9PyZWr8X
Y1MNaZpUlcu1ZAHc58RSx+l5KH5FvfIQJop2Jo0kG0qM39aUisc7wQNYulKElIgfr5VOliujsk76
fwWF9XVlUrVusyrmCwEat9zzKOcQUUMPBYcSuqntXd42TPQ+F7F2A2SkgImDuoPbZx3oMmEofm+E
Z4jgZ8nLzVI7DSxl5FsUwQD/E7XP1XhPW/iLeFGh5+lgP4jXdXQF9U5Enc8ewxuPCemBRdW+6w7Y
lhcy3d6bRje4wtCK3pr5szTaaC4t+VFBb9CnqqfAUXOURIxYbReIqJN8qPtxJLKsm0PjgNjxZvSv
0OPV2jsiyMHJXYnawtPcvo0g+2m8lGBL+YMvk+HtF72qRvzFwXAgzLuT+4pGd8p3251oFNio2rpt
WMH63qyz5tmvVbZC0UyqjvelpACdcbVfo++3LuXOfn82lkT1ZF5H4oIfC1GpgBE6xq7Ii91kv2s3
+bS51H4fU2pnhPSGUXcO7g6RGEeYXva9p7DQ4cK3G8PuMFaj0qp1NPGueuRkfArvuEFiwxXMwbnE
OtKtSC2eVVJIBN54pm67hCmBK8ZlvRh/5mrZUInl7NwpZLFNgIVB4zxtbzTn4j794ZEUHTROkS3T
tXKemGSHfS97TgFOl87PtFrSQyQ1En2nXjyKWUjhev7OTjbbNqgxtHjsKGXLeISLmygjVCWiDUdu
HpMHa4F8ogSYHGv2eYN2eGxtp8sSDGo0QKkfV6DbAGFVrMijHK//pbWo0zfaqqJT9evSu3B6vpaT
gEMFiPy9UlFEkZHgTXF/15JJgt+7NLkwUkn4lts0/1It/7MzojlXMoYkEspMhNnQ1qCtqQYO62r9
mSEADJTKGYhOPwkChYFIoYHOVw6P1ZwZ/ZTZ703bBeajmjG9P3rXx07UqLkJFpHAb2NW2Roc6FTW
LnReLRo3LVb3r1s7BaMl7RPIEkuFBPprq8rnUCCucMopZabH5OOplf4dcIagOucsSFX4hedr+FN8
2d9fjtLDPrfe73lsC+dkWskYsYcgVv0tbt4DZ0wrlfbApEP3hdhh10MtXr9c8ta4kt9yOl0Yfx/d
x/pgW/pqK5eA9pifx80T4xlIRlVrS4RmKK2KTMpATHTa19jR0BS+uTyvvylm2lr5AqnRY8rt4dQ7
ICNTrlXxKDdHb73nRWPpfBqMsyTyJuIkuIdj412wE11HbaS4OwqDEpRS25yzjmXY6/dNkxTXz0lR
xxE/xCmFUtq1XC5SMXYr40PtqW3d4kj4UeQfaXbCd6Pzjn/X60tVzJ3ILepeKs6Dm0MWbld3vWmF
/J/JWR3Ledy0Bt6LfKh/KnA9bobVIOzhWjeVR4zF5bL/9UH7QCtbYXhA9/HdBguF6sGxLrQhDVD5
U5mabt3ZjWQREQX8wL3FKMTdxAaEeOBnlg0yTJIVclZ3UT+Uy4PNPAo2/AC3j29cSvup0UQF2bdF
CiIV9diqurkPWheEk0fSoSBfj3keIbAu5askGXFzM72djBXpWp9Y/GSTbe7rzQvB5rVW53pAIpbq
h4HrdfgyezOfdAD7x47OnBAguUkkUcN9zUSyd25ctrAZDcVhRbFuLwUfo7QKZCoxK4eN3pZSdlZp
WKdz2gH5/lfGy8yZ1SEyWJTKHErtU/b/uFq50UHMtq4RVBW0rhiUSMInIeg+nWWKKHh5A8BntFEi
i5qelMfgr8VJdAuiAGOhSWhtCbWyEtcF5/T1IMB5f/M8DHM1nN5CfQQSenVg5i0zscNKPnCC3fNt
U6rbpY4fGau+yQyxunk9b1CHp6vduHrJWScdmUFRUVPQIpM8t3yuXe5FBsu4ASwBAMktTPwABV7W
hg/PHasnfGleajexgyBBtFpdOelUgCDQ9pfAGdxgx+1KFfgy2/qDyRvhEQ0v+lS6i0+v48J+BzsI
qNWdbgr4/7/L2N6lq+tPJdk0MQO9++U0ufFrGm+fwqjeGVd1IVfib20d+sLBbyySuXCRgHkgzXXN
WiMKD+blDOKxlFmT0X1FYT2Pvq37xh/RUjziu5hJ63x4tIzHOX25f2PPc6SiEbDlWIsnenMJGbxT
QJPQ0K2gwa+4psdvWj+VriG/dSgvU/W/wUFabamY/+FTp4XQbQETyl1rZiUAVbJT9ql2SqYqvIAl
HHJpcbkXbeBKQlyUzozXbnsWlv+hnNy5mJRJnTYiP7YsK1Pb1DgbvvN9AyjCYxbSaw5O6MHPAwmQ
RVSlDXd8cizNmEO5/K9qZiLfGrbafaYLvH0kDMx9rOV9/6K9L+xgHUT2Ezo80xmhBUTy49EDNCCL
GCPHyVp31DqNuARW18pIk9OkkoAmO1KPg42l7NsOFxlDrHWT5i2QNr8U27Ca5Yir7u66+DK/ECNb
PFVMJX1CDWUG7+dIIgMwkq2mQ6ZGQWPJ133qFCnuue4E2dTNe1YG8aC/Oxh6V+8DuLn5Jb1T89L5
ivtEqKyzznF+Nx+3eRbMCNW9+edjgvUsbcPxxy1QbqzCc49RmboOc9S2+9v1mDJORJBWi5zhlG8c
KBy8P492p4xrdf9Nr0i+SuZ2j+PVu6uLyDteLH8dfer+3KIAH7o0zvy3jP/RgTPpSILh9icC+ayn
vYfhtUXOyt+tqX/NXvdg4U/nbnv+ijMZo6RZ2Z6+sVbpaNzY5bxYtdmBrceYDjwH7G1VliPnjOgr
HHgzFtRzFEzktKj+/twUb/DFNQjjSsyNEFR/tioNbtLLBGlvwq0qsMUd6EggzfGVY8siCva60HH1
BFBXd5ZuPyDVOp+z3dIjd1hxzOoL+mxF1g5+1YO31N33bdLrMIM1vZArEcsKuQLy1lRddLU9Y+SP
V7h1m4XEHrI1U1z8vJr5g+sxaILRG6eVB7uKt6CIPbtgdcgvTRQSR452B9FOOsNO09JYKMp4kHa/
jyfqJ2TxD9IxzHqaOfzYViwTfBVPgz3zLBUQ9/j51I2Z4/QVZ81FHvDH0fecGPI52FxxgHsDj8lv
svuF+ojbjlBon+Bp6b+L6nrY2ET/A2MhuxS9c/1+cS3JujoUpWXQCtV3gWaqrTEBNPQMMKeuwt06
IhUT8lS8LM8/GvQpiaZgmy+gWg0eN3b7UpB93ANB3GYqjwjeBGzTNOnPRNSPi85QbFUBQH8Mb2gp
VHqmNlFeztfVz1vYXIG8FeWLNMhcoB45iUVZEWIMeyntOJzYjdTpsd/P5fW2DpNeFX/QQxv6WQ/i
RXMwAo6j3SQgcT9uTCKHbajOET6wHkPnoWemDrjA42yPyAKZxzs9mxjART89agaXhQ6IGIGKVfXa
yDddqYt4jd1d1Ts/fTExUn/xzOSSuwJB12aSjyGCbN+y2I+q2idXbWVeovGX83Zql3/P2lj2yH42
HBxa+stKbLtoQ20KK4QChFBrTmzcquRA4kEzhkENWQyHRtr32aiK4HtzIqeqWfTdjghswhbv0IlO
Drf65iy0WeTlTps4RNgsTW6yBKnWyfJvWBSNVXDyudQxiIXOHun58M/WbkpGT482ypZ4Ha2TLS/N
60G3W8ZDqfJzdEpZ4F15GwvGYEyzNqOrQI2axiIg4W6MOrrnS9jC8bGQFGRGoBbnEOs8ULsXMIjX
3k33P/ZMGljDT4ImMESeBpl7N5zt+oTTZ8OU0zUhGARlZ6lhGP/xtCHmtElx+nH7wdVOcDu7L1mH
qnsnf+iImVLjBklkFjR/zK/c7l4naOOiliZJ3KyhDnkmuwVjNqx0LbGLJ1PrH7L9NuWuWWCD+zjB
8lGyn7IC8oEGnHzjrmMq6uU7+/iopuL86Wfp3nLEfS30T7ODl3lNWEIE0qLt335RFR4a1TB2w9br
uLBCJhnQjEoogWPxNftPpN6dSxm4R1YqHLvt2tn0Mo457UajY0WjDuvE3+79v/DkSkeqU+QzYHpm
TDvOwOYUm1wOuO6vcw1QCL/iCJCBGxZI2nnBHlTpmxfyrW/YvHpQEItyyTynKJ5KDEFT2OHKJ+aN
tpPOHFbkwgAxoDvHzKH5uzRXA7IcNZCeaHpFsosxKyuvdawy0uCUr7V41P5fi1pK+FbBNCnACAGU
JJQ4WDl6bHwq/fVEksiv/m6sHnXbY4pkRvG2E2TR6X14cRtsMfxEIy4w+5BpRs4ARhVwx/owQRvx
rvUUs6L1b3XEhDigyngOMlqm6jakPz8aOWZ275xXo/3jBvmqnamTaYosZNFKpULOYPGXOqpstcZa
OuRS+eyhnPqDEcgsB0lKjyjDdmjgbk5vvJAJ07uTv6m0fD/LvPGVgb3rHeeu9TASXqhiZKK27NC9
5OQbzetnSnSWl6EXCsfvx6aFoqdO+fxjgfUnwWLqgjgwXGBanLwiPWf9bHwVFHfJ6Ba5WV10RG2/
H2DEhzV+PJNbTDs+29mEkmQ8TQuIJZVCW+ZaQiNfIOnFikF8Gie41+6SdZVGrQI1DLU7y0rHS5lB
NwxvaS/RWOIt60NDwniQU5l+eXylq2/72CdXkMOM8+oAS46X94j+YhnThhJ1KlhxLOl54ZJRuSDL
7qYalyhO5cP0NXrLz0ZYBXEi05jrcYlGiXwiipmjDlHPV1/UjWsGlxLLdcYLgnuzAVP7NCBf2yJx
ktGw06B+Mmzo7Dag///4dQw1QcsbIXJQr3eK3QtzEUg5+QmiROdyACvFRMibVSFawrGU7qaP6z1U
winZoJO/yDnOqioE3CvnuYxfe2yrb/Q27APYiiccLG3cjKxAR0GI1uSCUQQNV0rKQHU1E24P1Wlw
Ovf24H9eNdJ2Cca2VAtDKHK9GJkexIBJb7hfMtLZApl2DKsJaEyXe8GypexBmmopC4Z4Exc9fBQw
qxyYORQNf2+CIx7vfO6mhhCZ6k5yQwAqrlc18MOIrxlxe1GJhhbcq+52fuVDCXdpWwOUHXtU0Nhq
CLUIXHQ45IB+5B5mvK5DMYa3KGSeVAZwKvuEU+02lce55qohchtyVuMapOdXJYuf195MmCPTqkci
k1YnhNuUaqMhim1Swtk1Mv7pUosmJZzciBMhPVl0IAqPeGLsR87imEmx+VRAJW035kW5EQxt6kQX
L38TaGqQHy/eMOFzQjvsmvihm//hq/OHED6dt0EE6s31dN2Jn2kCzVntdcMH2jUOOMiGxJNFSArV
uOrHWBD11rdafM5eAUcL+KMm/ahGHdW+FGbo/9Ddus+fjcBnCR+epy3pOsr5nHpjmXp8j9k9Kmqq
Ju1o98RDBdUZ2fIycM4wKKgvpmjNQ9WFMNEYoa8+CfYs/124j1xMEO0tBc70GXWsEJ0IYquqnj3x
tJ5GzbavdxfFxG4z8YqOJzSq744pIWUYPJK6y00jeZyYaNwJ7wQto8F7JpYztIX5ecsMSJWkvekB
C9uJ4gkDudaWupQHPMx0RvvSwichvacLUfgJ3ltvdYRS/uHCA1J6nX79RRCSLZfxkirviKJrA1Dy
q2Ay04/lobVhOJiZx/qbQ2rCxpeZRXzQX+rtx3ZI6JJnNARmyDAiukz/Cb+Okz5ECJftDV+zoB7O
93ETqw4RbxNvilR9FeVd4yn283dNlf68QgeQm/ZuWXptH2uXXUfCPAN8OhDMZRdtVZ4b4R0/Mx3G
pOm5jWh8rQWmBBYIM20jvUjuK/9AlVIsigPfx2Da/H7d0Ecmaw0HRWINgdlhCQXbquXK3chjYJyk
ZMKrYzKE+3S6r8D/NeryAb0I/qjST06xjTLaj2REJAOXIeXCjlwpsl7GI2mpKUohbiDUaJqMJP+U
UBO6bVD47diD0CEc2laF4DWEl5KhdsGXi7UG9HcuBEpqVbDRCVDAsb+3nCC/SOC5EXCE92AeQ73p
F5PsnofXuv20Q6WkFUuyRphFbp5PcSUcXLUXkVeOZcZnXNtWSGun+fhtw4QlMG5WnGivzl7lc4Iv
YCnI9sfDBiZjq/BuLoRwaOE6z6RxrSLK7DAnAvFI0nVzSWNoMG440DT77P3nsMjcuKYkbFQIIQO5
h9dy5Ej+otF6Ny2NiekLReC3y4Fiq3MZkHoGX3JN32Hrm8FA+dWzhkiC0BuxD2H/4jDGSRLqeSrd
PacMTqLdYPv0HOLX4y+ZM8osd+WbBokA45Gd9zrXg9/0q+MRP5mm0dYL+6yNXL0t3rDH7Cmrsjuo
SHugU7avzyDtFhLL+Fk90mH1IeJegY+K63CrwlFpbwq+XHDOJ1gIEFhR3oZXz8wOdNRMC5TJP4M1
X5J6LFsehNbP49+mKBriEkJu/1J6ftdpYUvfXHTsGKc3qdQq/QDIuiGhv+5HTsDde+hpfzPQNjkS
UZBFGvad15/GRFinzuO8Q5IAU7lf8nR2oFuf09Td4EdnzxPzAvgqBsgHl6LxvkaB8IAgADxAWjZK
xa7rjGfFFlHEgGKv9aPbNYHG2+DRZdVhyHDyCQffP2FoaEf45SsXY2gw4j8VurczndbdkxtWx+GW
UHx11EuiSF3etSeHGPRXSljX1yqWzemns58uaoH4j0uPQdJCufid4CIiaZKWvEa7XdtcX2hRgr75
KBX+jag/QD7yxv/sL6fk2EqFtQfpI9wwbB8PPSG0CkFm446gALpiXcU6Ya3VC2usw+We13g9AH9G
n9Wxua5pBHW8VsWYFK0Maf7vCHmxuiRL/X/R1LeHFn42wnKJ9E3Ob2ejicSwW1LONLV/yk5pVQQS
1QHslhKsJwixnuFojG9vsWHTOI+Ci3oDGn6qT3ouVtPjQQabGZKraoi8QXfIdcgBNNUR8VDhxWPp
sXcPz1PYrIClzal+h17FKP8aCKt9fCimX4rueprtlxvuez8QPbcT686bAwAlXVMyQ1oNhFtwrrGT
SO/105CFzZUyEdlCuzYvR6NIbxORdsjoEtjkU7/g0u6uY2VFlAXVWp0a9KGM7SmgcNP7LyTzY/We
LgLsqQwZ5MLFSelEWdos/BJSqIlb9+wPsU6+OF6D/m8LKDRHGfcQ42kIeeQT6GNPIOH76/kJE7pY
Zjj2lfLSDCIIW3uj6ZnhJbPM741xXKFQIZqCZ/AW+scd4EC6BeMzMNRMoHvGRCKo2DlSG2aadqkA
wR+Sb7zXia+K7MpU2GmZGKzPVOdTAgUnIYBPRqGACbLb0zrJUKL8MYS3IB7TbHKepB7U5aWToqYs
YH4MIbLgHgLzI3uGQM4Ood3i2o8B88U2IuuP0/oN5zXVRGop4xHl1cWSXA0Od+UuHxM2k1gPDIQG
gLf/HYfC0h4SWHtPRQTrrNJZarFm4cywtMwQyQLjffiskmRMPiqq7a8pLFv2jUeF916Y2Pi88BXg
6SjxM+dtPh+Q4yEXYwJ7dAjcsfcORqQmDwpgrjDH3oEk87xCnmfGNKnMgB534ie4cKRTHRU+kKgc
actTaV/DruXcqJKv/NAw+RDYbriUk+h2zZMad5rXyCPDl/5yJfdhsQjTmolcCJp483+4UV7o0xTZ
YdqYde8TO+P6aQMkYFkZk1vZ/gntYkWOkX1SWhH63Jr8IZuNmEwKI2CoWDJ7WKwvjI+JdxyljkKc
vvKITew2e2iUeAnA6+iPKSD8fZI7xRhoT14q8FsLKvL4zxz9p4LhxaFUnStY5cegRh3HpcYMNSb7
0vzs0O3N3/maNTgJsU16g3iuGEFoo7igt3eyuKlCmQZ+Cnfy5FqqBvSHmPWbfdD6lAcu+QhU5aXe
tQRQfvqzYrJrI49Lr6u5w7s/Fyus+FqI/4PSbqyY+pDdqJm3/FXpqb31iQ/WDumM05Ap2LOQIIiN
rshekpO3FQjz0EBel08Px6pQlqi3F7N2BY+eq3WxVImvajnZT7UwIOX3pShulcTeRI6xcNTb5VfT
dKtMBPVX//qvv0CZ/AzVzlNxZbz5OgXKRmXw3w5kNFuEi0a/qOnsY1nyicFC0XddRRapAYgfmwgz
Iwk9NCvmwbSylsXV71TxYUlpkT/y6G/uNG+z5Bckq+ZbcJL0vlNMdxps4u2yT54cm8zRHmI+mRz6
NB92RMXI/kfHZ0mL49aK8SwHkrsYNleZ5+yniY5zwakOcdPD4TG1wwIgh5sn6CDWdmY02/JhJ1D7
kCcb8OLZqo9U78iKUdGzcrdUGEMk3UvhSPj1VsGLy1g7MroQ2i4iqD3+mvaML2avHOCFLE1q5pK2
6kxQfahTStZ+HOy7NwMBV9BLj3T9dSBCQtjv3SjDgNFGyXVI4krM9cuFigQaN53Odj4Bxa3Q2Sv4
aAAdcJMjxQw/FqrJ39EwLedBTSXu/3H1mDOc0UQWER9I/T3AvAbLEywJA1w6o9uBsDlLuWwAh8PX
Z9QggIKR+4j8kYzjtRegqmTijay3aD+/zRQNv/ZLMCBitfe/IEbF+0Iwtbgi7db3mr8+h633Li6K
8MEaJR4+aw1MXjH5IdIWxSSnZNHsYASv6g4HI1QerztyH5T5xUPtVRajC/4q9ft6/Nz0oSYLMPGx
/H1swaqSx72UlJ654xhrTsfw38wB5WkiqDW9Hk8LoOYFjNUEvnhYcavM3zK5r/RRL0tRdE3XQF6x
TXiJov3sAE0A8PMUpxDfmfXTe8wP/uLwcCTUiNh6Sz7QBxlcZGCGlqq/lPVXdA569fHrOJrv5oU8
+rwj9XLzu/AQSnthSjZdj3et94vgJPEFBeMTT1mP//uRoZ1axixmGExEQtckGinC4Cspd/nvESBh
MeaYx4IJMj552VKmb4vZUKMg/HnUHpx4L9owNHPWGPBIMBCE5oNoXaQF/48yJPt4PmQ4V5YCpHt7
wLnFuqHk60XfcZQ7KXcjgM7fSCOzV5OOMastEX4vXutMiAvLQBj87o6CAYFPlCeFtWs5mzBBS6gx
XUCNtxlcTXpGAwMfw6vY2yz8TgZ9WBEyWi+2+nwwMHHfKyF/4ivj/7lWh9pf8EEJzUlLmg1DuxQW
k9Dltf17Qnj3rZsXQgQ1QWPue1whrctGY0WVy7inkSzYXohOg78gNWJRj8/rTFGJhkTsHLK05d2X
UhLrnRHd6PC+f9DEf0mVlPuTwrqEQUZFkSyWt7JyfGBeiGWFVgZxqwTCcTDuNC0guWZhreLpolgZ
D1pgapBnHKZdxYm9QsXbjU3MY1/trUPIw96nR378TnYZKlCogiB3NEUpQxfN3VRlmgw3Fc4MkxLE
DMlawPI26zWcFFn7ft6f/lHpLzz1f3SVIEY9pnW1fnTAIaI1wPuZviYGTXAAEFIVxTAmOEaEKdvJ
kcIO86JR663DSgIGPWP0LWQUBOLwnxQiEUfrKY9Th9ewDTW01xPAYTwNlWZElcNeOX8mPod3CISs
CwU8z8hKirrSjkj0HLdWHjR3k7sDdwLEEbKIJ8zaC0LTMFZDWWDmfManVR+vutxAD3YamGNJ6L2G
Zv5xP21S1ioNAkvrEIqfDjSNVLO9XdSLxu8IY/yeVPYUU4E7Iib4xQ6aXUHNllxnjt2yzoxef+q0
cVqnowu67l6yCfitQXjjSAJmeaQIWyU5Nta8YgzhHK89CATkT4Kse/RnSoKwZqP+VR2pwAnDG3L+
5qq2tHgXQ1b46eYRGweO2LFM6++QFev+RG43QqlzxBbtUVSQXRYzRCGA7BD4YO8f/hoC2Orn1ja2
Bq3UuFSmgNFAyv9r26s0gEbhY1h8i9Jdh0O0UL+3N/xytj5iYNdLW8eLS/QdPmEF7mO6Q05LNgep
pROvyl8GsaldCKUmCXOlzoBvp979krgfIbMdyBHbPKbr4V/+dm9qH063OeZwmIFEIi8RP7C/ehTn
k3eO6l0Am8/JbwLlpjuRlzE4aK8AKhuvbT7ids4JFMsUkqi/XiHkZ7s+aq8CTojLD4qDAHrGjKOl
JV0n1jogkByflSCMA2hBBj9DT/jxNBnthjirJQ2ZR5smLKkVmD2lcJrzhGMfNZaO2rmwKTuDH7sU
GXrnCRD4n711xfA2D/6xfORJuaH0/4pxXHg01bQgVpy2Oxr9LQsstBoXkWXcfVEA4Ysd+UK/nI+q
0rY58WKRz+nFVuqD/IXhRbQOgr86mlQIAVNfAXBMCKL/bv+4zF1LnddBYFtn1S6YxBAAkocBav9F
c8bq2QRtbi1+yL8TycouhFeo4nFSxnh7V5L6ShSmDMAAbLmrVyTNEljzqkvD7ijkPQ8U32aFBCxu
x1fAyq5aZ7/C/J1lqOLuqH1K+tE1Az32cMv0CICBeZ5t3qYe9k0Kg9Il+06gtbWPJlhkHju6OuC6
5R2HfDYj/JVcUAogpgEVt4fL+IeGIiBjDT7F9Vj0rtBTcQU4Jmoa0dxLbjSNXFJmJc4OvUODV3lU
h6RXyBO0BhHVd5AuDaMwq+kS7S26yGsNK5E6NNY7VDffTSdMa1EBaf1cf4Ru4GkrnDJsvqZwwzLB
5uL9qwdu4Ivy9WAhfa4iUGfuWVU8/zbIoWmPznOyoYNPGb/vOuAVlmGyh/gyokrYMwltoPKSZ+z0
lZFElmtKykn7FYGyTxaxkdvnfQUmq9bLvxW4pCAz89KJAaGpPYLFAuMKGRcYesKvRvtyOtZlm2YV
zIHu1VNE+Bh8DVvmv4KuO50qztPaIG1VecPGlo06CQBmYaDmiudQF5gFmI+ZjH3Ncerq9DwxV7+J
y5PCYQN2a01DEM0FnFZmSfobB+Tt08Axi1o9l/S0syWYz47hHXspWbtYpm7T0ooQ9WvTR+2KajXa
8sqeYrn+ARf7Mnw4drZu7VZRxmQbMu8FXICo+7wdCrTgw0LWqRqA1YUSkgVGIki/PrhNzbpay/yO
E0ULA2+WtQO21N9+gmPb8E7RypQLLq6QQzm7txbP0bTtPxd1oLTFHms5YK693TeYE81AEExQDkoP
ZAdyH1QAhBMMNukSR5prD+SEVZU4r+j3FPKlMioE6aSNIzrHCZAcAqm2G/0w9OChKSkI6Yr9KWi0
BcTq/ojTvEnqhGgxuSH2yTGvAPceBi5bXXZQBUqFVrP6yD+Rl85u5azAz6jNuAFd0TGYcDGjg+VD
dTROF75vwEsi1LQqVFvn2rUn9Vv6w7+unggjcAeSG9FLDoO980BtHp2AP59rnCJ/dM7d+kykKq7O
SzB9M8BaYA5WHCnQNqhzbwryD94YHm6vh6lzmRLjZkXHbnw/QZC5DchUoARFkgM1wORSI/LIwfO4
LWUY9SW3Hm4rtWiCIZAr3war5+zpCFMy1tqkizn8qkrBQtvIRV7G35vfOya7p6AADe0dWpkwSYw5
0cvJuSgX6Qdgen4OzzYeIs7oN5EtsPXvcoSk22sR9IGA/0BOnJrJ85nxs5ksUETD8QLYwf/Tf7A9
Sy+Rq6zsv9OEgTPYajANErgre6Q2SSUPcnA8ZgqixL8uyDDIJOLwh7yTwPrkTgMi6ZzPJFyNMOy2
5raaZOyEJ6wEimxuhu8KER7U20Ykkt13oL8JZKFU8PY0kebFWUwWVoz0rMeZEP9p9oWnrTo/Q1x3
g9Nu0Y5Pzxyvz2X51ZhQ4gi6x6TGkiPYq6OrPEDCUqD3kPU8pcYOHaR7iVf/8P0PhT4DQ1m6lwa6
LiQUzf0nOJ/nvSCI22jim79ajLnphlQcs8kErFo3+5Mbn3NzbU5PAclWDUQM3wys718Ad0zvJHap
C8W/XYW+jgeVJhXmFxF6EBJVqBPqW2TYftzW6NnGfwhvGie1UkXGO1W3goZ4BcOyIzWLnnpbX0ds
yd/4GMOb1mTmk3b4crYy9EYRvP5rgReZ19RuwvhR7r/axGDvodVrZfaqsGiVbgI15AJVAsqptwA9
Y/6Llzvurcz2Ti46pYeIoern/bFmv99L5sI+Bd148JkX596UTutjjdl8pD4ZUazRhfKz/HfyrG0n
9QbSdvO3gH+/9GCrozYMovFbPHx33OJXcToTL2OVzbDSnaIxs2swnpPCindBNMmuW5C+Tc3N4xmp
AZYSJC1oc1H/7JRhij8c/Jl3gYkgAwl/sqdqmkEEHOIiMM0pDg/vZc0H7ofzvtMCxfuB7WP9nWdv
ul6YbLR//7NdE3vtvgQlJ+hPPUneqavYvx+lJvLHFkGHiFdbv5az07BFQyQ9m3VcCo2LPfKVvkQw
gWtkA7xPSnZ0x8kNhezh3Jo67Ur/E0N3i01bDZmlrffheIxQMjWhjeYoLIBEPdMEqsc15mTQvqEq
/3qDHQEVEO5DPBEkznxsBX3LEHt0ACp7NfOZH3Xuwun4KfO6ct6ospErmEFQioR6rQ/ROwLW6U3c
2zei0390xBL/eXj7vaZjvwZx4Wlo53yD2L25YpNliFiNDTuirqjFwd1h2cF3bvvvaGJ5sDplgFBZ
iXbAgYGFdX0c1+ZovldFnJCPaPQn2Y9/BZBHWxyQLiRfW7ynKL/BRvi8AnA175rQRu69S+IZ5jOc
Sv9rPmo5tE7ZEDO+sqhPfQtfZ0yBOsee7la7XGnlOkARyF+GgKKF0v8fhMWmIzbMq54VLcQcq7IV
Jd5JfR8Dsb0Qd5Vv4lCksmNgWZlaI0+7NYta61Ekup82+9WeUMsb7Ed+xMyEycbyXcaEIel07KtZ
bmhdD+330cM6M9GnOWG1U9/xg0nG8jb5pLMt3z62GaNvgZst5T3Nn32tMjvBAzW36oBjj+hm1DKH
0WZ+I4bPkBZy/4DEUBOmJpUUMiv+esJqIf0ezLm2aerv+xytVB5yMzaOvEodD5vTvz9zAeTd7+3j
vTsvBmqGXZM3o6V5XJ4FQTcS4LkqAVbgA5E4kcVRESkh2GISJyC4uubZOUHHXN0lk6t+2wey2Mit
pZ/oGw/BsAmq4xVi2f0US4M3+qN6zU3gGXfaayBDdgQvyfi/r2dMQGDxm/MerAjSqTonDTVjFdvU
ARAjj75GOpVWOOzKUu1YEgQsn2JLGhDgoqUri2pwJ8fOCpBa//JOyl8jclDZFbnB25rnShpkfv4M
ADCNfgy3p3IbXzPQzRWcKSwDVZB+/Qj20LNNmw+J81NkGM8N2fOa18AA31hOPXR/FrIUpMrlIKt0
XkGBpkapzjOD30HFhYSv1C+bQoTALpRLz1boktFgG991XU2KnRrgv2+fmbxTHGbcIGlOTa/St1/5
B4k1XSRkipcJxJ0Wqc6nJGsHhRrpBOwkudDH+J/soski2QRiTECExWki/HKNpNfbRFMjynpvXYHO
rMd1d+xcIwa6eHXoDq9k6AmUMfEZdhtAr0GcnACCHzXMcxIQgVzuGKNXxwQ6Rj7pFzJXTvpKISbz
VVwyPrWsEq6btY50D+9PgWlzDxJt+lrwYGXDTNPad0R3B4EHIcmmcVRWBYBNZLX0E+9GT+6MDZQg
aGaQdwYd63AHHA8rAxQQpcmdQ+i8TVAYdk8U/RJo09288pDNj/FKlqYVGSSHh6hTaytrehGkdSut
xHkNJLexHLCAylJYf3pKo0s5eqRdymM9wtNv6UdxyvRYUzvj7QEenaNCfVYoQbhjthxxBN3VKer3
Rz4ls/y/6mEdwrfg5aobCIRGIVfPj9W+24+G7TEx6ON7yp3KwBWPRgrZFwruzudbHDJVPyYlxRd1
aNv97Kl5i7gqwG65wh3MiKpCDtqZexB3m1BDr+TRa9kFENOeJx73MO5nzlFQSFw99IwmENGIRV6B
VwxHURZsxZeRkDO17LQqcjBzdTUbrd52CUqwpVVd660U5c57ncJeHgChA6YnqypoXCtyQBa0uDZm
7+IPJjbmvTUEb5GVXb12mQKrK1sMsDr7PblpAbUrrwS7zFb+vEKQ8XHxBmbixUBlhzC31teTqO0V
dOE7RMr5csC83jELCR/6fGuLLtpdr6zvD+td5eV9jqcpNN1oOyHibsndAjBfz3J0VsBBPmmLt/Ob
6dZ0MrAxsIfYB46wZKJdgnT6IbiUDfz7ML8QdKaWyz2gc9RaXnKAlUem3aCIqL1uAKUjKs5Lj5eu
6VgUn7peZl0z7nBkECfeE4G1/j0biPDJpMLCY7HunscOccHjOWNH6+sLO+qYf5+kSjZddOhCyT6q
EjljlHFpu6uZDod3USoiP6LTA79BCv09LKVbqmudyZ+uFduvyx3C6NTyaK2XRi29e9nmiXqwHpJw
d0KkE42r7vl/vYCr1Lw5xYQYbLBiyMxJWo/Q4LLXeUF851HHDFoyjroxC9p5y8pfCu8QGRrRJ+mr
8jUr7aEEaUc7kZGcCBoAx1dj9Sx3qnCA1+3Buf3Ms9FAoVA9JNooN6Kyp9Sv/Y4lTRyoFou1/Ro8
9H03/p5azwRN5k1A1osPva/fceTiQe09g+KMHt85T7P1f9VEBtQigHZQCs4HPZsGj9Du4VqEm/cs
MNybGO312A6HbsLlK6cZciNrCUrvRB8AWGy+5wazD7XoplQbzbvpQG5WoepeqEBOAiFksX+bpviC
/sRpCjoiETpPskpgxiiXD+Isdep8JYax8XKK66DTQhniJMIzhIFNtxE7GqbpG2PF/faZnkT3eCAw
4vxdNP38Dg8QQOtB3AXYvORyEYZ7KIbZPDnubyNM2J7HAhKd1O4zvgGR4ocID2Kwi/D9e0Q1ht73
RAaYtz2ekzuJVQTW0tVkD5zdfytNCXfRPN8BDGSUF82TyeThZxOjUt4buh0qtA3imET3nVW8ki0s
gQ4yzOodMH6hjZm/ypDDIPEaCpQ5PR+A62gEIuKa+b2PMtcG61xGFq24SDxzKZLHR38XF4hFirUt
UkT5UJmZN0cU7RuC+0oifmB/tEvGN9wfTIj+Eb892s2uorxTij78Iq3WcWFs1i6B/xtW8ao99zzw
2C+4h/zJW/Ca/WrUeX2usfgoZweXDTbeXNXpOiBBhpzpRO7mO2cAFg3b0ECF8f8ZRL6/TKFcjAzi
ZasfJjJYnWz1Fem5QOT9IUCRSDmWiaUOOdtach+4lMcq5/DDFBWo4Ys17uOrxjhU41z1bSXoY8OZ
bfwslQuVfLQK7gtyyz0mMUlZZIY/EaCe4hsI9pW9Q3Y2h1pOcMWg/LS5z8dl0V32Agfl7SG2kmI/
sPY5FQQB0/fPl0M/FgSzwxwf3L4ADga0YHDrhRRrQeEFVH3RiBYC2pUvjFicir/C9YM5FTVrSrUp
KlL1C4pg6j4IhpJIQn8cW2f3ePDScgbZZDk7jNivhZhVIGoandqwFuqCTPcRqhby6vxKzFaTI2up
sUmKxTLmeW8Ilf6yPO33CqSMmFTZUkoceUnJnQNO7Dd7kuTOgMXhxKog57uUvuTLrAxJ64PUDTOZ
DXdE9k9oheeOyz6ytm+wLDX8NLqIciuvwLkcjZ3vxrq8TD0XYIn85MVfBXDkTH1wb+Jf3Bnka5q4
Uq2/UIGNoK4gHlcTUna6hslLu6TI1r8Ekdh9YakJdTklWpZSoIsQ+N/v5vLzMObeTfWzxfkcN+rG
TmithD6iPi6Fa6QHetvqAsR/J4mSfYqzRe1rlOdp5bqHnu4TD2Fvb0nI4vJb9TsAO3wGReTxchh3
H4a2wNU2CamysSnUY2fF/DRcdhTdangUzYetrebYCjm704Kd81Yi56KQV9c1iPcBQJ7M8zXG5SqX
taJsvGsaFiswvLmJG0r2R4t1kpe6sFo8GH1nAzid0qp8AfLy5N8HXDHB4B0aZqGPRYEz7kWkEwNL
r1NOwl6tPz0AU4omB9bVrUDfYQCrH8VCG5UkVIYqWUFDjQqf0iIQNt4TsOkQ2DgCyrYlGTQrTegC
e/dbJBF5Wn1VgkcONRIgMblIImGLhxZYXLAfqKt5V2FnwAOcXh5szsZ9pavtMAQ+YPvrFwU6MTTA
G9fNqa3LMnnBBEDWVKSTelHo63dvSh5lWdFmchUZLjvWdppFU4xB8XvAh2BHbDXNKLp9k86hgDyj
4LYK5N+2DOQecbXTPnLIbpn24OwNbJEAv7D9dcX/LdsfM1Y7N9eoUQjelOuuZI6epvhHhFDfZO9J
A1nZ7X5IqtM9rpAiNJgP/RbUCc8izyUmLlTnKJSeq9Qyi/LuhVihXTPVPk7IpnmU7wYqH+1Eotsy
W1KPvtVedHsgDozVB1iguYDHRwYyMiCyBR7GoNWmTfsRu4k2GM9E/382qik1tX6g/WEWgAYRRzEf
vFwmZxwdu6MKpZaSUWGxUv3PhAobeP10FhKsDXYNbAeQF5KBfZf8rGlNFOuDmqoK0Ar44lXm+hjl
wQZxitHyqT8wa8iVrZaoI+B95H5htiQxzSKuJTYtin3ueCqquAV9T2iAHWL29rjnfh9kdEE1gUwE
wSyx37oPtgrWDXLsXQaLq4vc1K/6pRHJ/VdbYml0YkBQOVmPPDchk6lwTcRuQYzAbxjzfdLwecRT
gI4SQCYcovQZSmYSpXm//Bg5wVIrYXyt7ABKoXZySty5j/VENP1Y/hKxfmwXFNGCkxf3SByKAn28
iKl8e/WLuNegRb/QfRTVTLOwldWPw6+m/qHxsqLT3yhvXHWHkxptsaxrT0s=
`protect end_protected
