`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gzlNRI/o+WlSJWhwFBMigTc6roI3H9Eq4cxh0Yjq3EyaKGoFt3w9Amrs/JLP96APFsK0vHtkdg2a
ZZo6fXbIrg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RmVnVNyw57yQwRkHQO3Fv+xqQysCFJLLM2qg1cCCSsie/6K9hkSLpjN97tI4xc2YFKu1zVWGyTLI
l+gOK6YOClZsGYmEerd5eieQbSWCoiKUGH+je06Bj1Me4a+mIoC30hApj93+JH/EMkC7MCuVpkrk
M61bZJ0LXrfuS5S7kY0=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jn5OPQk6FXg1L5vSDcf0OXQvFxivX/fUM7Tc6MPuTLCKR+Yyic6HVq+tKstF1wUXrTL0KkmkoIvk
Pgm+CejcGCA4zrVmUAiLOOs1w8RK/P6CLPOz2CxvEbvrlOVUGBFQZiBcw3fNzDwkbsHoCEvXPQG9
+ck25pZnPUJxK99XClY=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CiCIjIJG/4MRRfS6YHH3K1UMLPnTuW7JifxrTY12IV32SfChd9b5tVWMlBC6oyk5oFhqIOQHlSpt
Nz4JX2lND7m76Goigd6HH6eqULEtujtNEquDXpvS62+ifOdScMsipAkafMZeTFc9wn6MzylDlvKj
P1tp1I5Ro7aDTjvJdzzY+2MJFXoEI6lku7BQSFMTrDDjB/TwVFwe/1dJieU8N8PLCm9ZoQPVZtjV
M00qa7FNcDBMzm49MWsRtfcJ1RbJtqBAH5Pn/rGRa1nPRWgFrb/WvYiz70xor/B6NgxXRqaigVos
9c2rW7XoR665xde//Gx3EPkS9zucYA0xAfRm7A==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qBj9TFB6Xf2K76TYj63S634lJ+cPy8mUjTy5fMf5crHJsXbSzjl3jp5lFPoCqH+d/iZLZpJQ1jTh
J9N3FacW2gGLqSSvMlDn1p//6mTdA251+fq+mOEX1Yj5SD2C7/UztooxbZLo/OPDZPe1jSyDAMr9
7vmpcJGfYOEz1LJzup0a5glDfbX08a9O/9lnkLz9fyTAt3D7ckNs7ua23xEI/IBc0PNCatBff5MZ
4NFLHSIBoZkHeUYfdaHiku1pyP/Yd+8BqDq5YEAruLRRUOSLuVMPlZMzTtVHx0DRvlsGH/RbwjyR
Yznvu3d2abtgTj3uSre8PPZ5ZpkK2KfRLeVVmg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mfpnxAuBiuCZebC1d7qO8oF9i20HDcksl8wFI9KM7wiKRZA94cTdy9SgtHd5ygxFudYqYyd1dpSS
YyqsGveSVICZywImGlNSBqECoi12n83nw7r0RB4EyKIH2d/hTbduXNstw5RxKVKYha0NKE8/njxO
rVwwAnXcy1/SXdaMu2eMto2AcTFzwrj/JFitjlOlfO2FL8wEGYCtLE0atCYZmVDOMJUqmDbaeyFC
hWz5ZIKGIQza8kAsFCN056qUfACxKNgKxBtPaLryuBMX7zgv0Udd5MR92Mw1jOpcJTYM+BbFB47C
NIoItJDQt+Sz6uE5tsLlBwWlXWKVOTT4LU13BA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 610096)
`protect data_block
o5/0z/ZgalmuVL3RcvIZmcmA3VTGBFpwAwi5cR5iNPZK+H+Ngsv5jCPWxwOk9lmswReWEPCIDKpc
A7g9j4L8VwRujR10ggkGk7pF7v4kNENnxiSJYt+SsC23dDCUKcZLEsoapCRscEU6rNiZ8WJSFyI9
yAJudD9C61W0+IPIVF2B8qK09BG2Tm7PEJkPIdmfQwJm0nCISZwr3tDqbQ7gWj5IX9rHvIUqIxWE
GqBhbfk2eQQFHQpdvY/90TvXelHqBFd1pmQ8a2TdxubMIMYciQqIT6M/OnwUgveu1CuboJaG3ivj
IwUSj53anjvepjtdsQfQ+ZB1FDWeZ6qtTX7vcTCM1XRoxVoUbyHWU4/1oZ8wdlJYY88xvCiuFff9
XiPCdBj9tADbRDnN6STP2hYoSjzHXObk1Z6rBoJVENZic2bC8GYkL7ZL6QTNBr6gorKp5H4VMAcX
nfUzv4H+qIjWOzZcrmoDDNhDM3guOQGyABXMoc6L75eCGiL7oiJzHRV4ZZEPo28k6AXADpiKHe27
LKmfTEtQkS0GMvhdN+a5sooOwBj7kvWcxRZyaQajUYq+b5aDQ9NkrKj0GnsEx/s6cebof4/BH7yL
jPUGgIM3PXpKphChzEGkkdrhtAZWxg1H5ZqB2Rc95p6QpwaqNLowxYgTN6AIA9+ZwrDyvSPCkkAW
PuaL58LbAVBmSE8zhrLXlkbKGGNLXFjvk5eVc5S4vHBRAc95lIdz9I7pS7CVjSxTf6tLK6zklGZ9
xnMUq0YtqFI4QiFurooUhFFf69BD3LWh+4mh9b8kbegt7CbMpRIKGPgSmzkrWYFnmzPBzCHHbRSU
LkOtiVyx3lp110KGjM43QSldForZ073Ve5qFRVqggqSlOJratgOcNYdtllfKNE+bKqwQzc2ADXRw
tXed9lDMB/tDcP2828aZDT84gjP/EZ75yIBA/W5ew9qeU+GfZehjmMR4cF7Ak0yHnuoH33r0BToO
OX+lQaaDA8qIo9nDu3FnI5Jpbq03hNf8dADuzVEkKKp2RwM6pL0kUbx8+LgH9iJyJkszfO7hMCCe
DQ2ENYQcNWyb5o4dAbOk4mHE9ejv2YVLX39zwXas0DG3plaV7PjWwcFFfSm773eGDrzVk3SeOm67
HrE/fNbyrxZXgbI3BeoixK1cNiDoYpMUrme1OUZYrHRTGxEH2fj/+JXaUwEGrRRpmL/LLHtlRTYH
Vbi5aP6KVrz22oNJ/kpusz+4b7Wh68zmsEB0ynM13YQ2lzu6bFwkRKShXNP6bnaY9vDQIeBCavoN
C3/pxwjL7v1+bSW7pAH4MdUkLx56kFIvL48+ocExFZHsp4NN0nRvy+PFn2vb3poAHWpBEQvyo4zW
4BLxSuo18lxbQyDMHUbKQI9pB/GJGBUsWzHk8z/8N0xkR31lPj8Bv/crEINDGQSxGal33SUgmiRn
4J5S9qr8d/tRD/bWOaMPaKPG/TSJ3YoDZgv0D6zgdw+sKfnose6pPUeP9y+SsgMnleMgHI+6LaVc
DIhGfuNO3vJ0hmxZcoJtwhorNs9O7edd0X0XxVUd2TlXLt/+RLNIbDxqTZ+x+zLKxp/oc7Ig2mA5
27zVlEV60pWvUJgIgLsYD744WQHurMOrkl2vbSBetY91nhb04jOG8fMHF17n2RmVHuYpE/2igsit
eSiXw5P9KnKoejyA2iXbQtb0IpB+r/JYm25tORyEuWFTPVMBzq/fch1xiuBc8PASsIn7vnOKsi/S
wuOypmIgb1I8Tl86wpdK2rGTYXNT1n+E96Sb1dH/TtxzCdsqt5fkwcv1nIJlJC3uPae9iOkr3lUE
w29JTK9g8v117B1jWDW9uRwyIcCxPUw+2LdPwJlvRjcBf/01a7ieBzbyHQGphzMPsLoXN17Ntdax
zmnkqCKgpsvK4r1AhXTWtfev94PZoVY+1cExiR/riFly0Mwo1bOJlnJshsn9x6GlOKPkOOeGnAhT
c2iIVEDr0Of5UPIuNwDzr+ZPKIec+xWZ4HnXc+kuo6sJXn1uDZOOyvTftQzQieGOeWpIglYXURLS
ZHIn+UT9yYqH3IkgOyo9BV1aWV0DktVpywy8mzBH+WULVXArECNtC+FyRdAthoVmKhra/Sk4llgS
XH7A118vj/eJ8mnQ+Hyi/DheA1TKQp1WCBVV4To5IMn7EGbv76EAIT9jCC5gPfDMutTURbUQtfZs
5D+8Xqiyjz+hSjoxy/wietJJ5c5j9rF6u+lK/PiIaRNSAY5uVfjgZN7h9XWFzk+f+2i9rz5wPGJb
cG1IIRTwi5N9m/XavkMQQqsybcytTeiEulPfAlGVC6Zjtyb55d20xZNVl0NX8k1IUmmxxg9bi8aC
+nr5WsZ9sCcbRyh6Qm4viFl2M5vcFR7wNikXApqcMgMWB0saUm2kWC6Rn7qOzCNFHDodiseVN00v
ZokK0zKnpp7IoWT8eastNPQl+cBkIqDGs3DFgraETa7ch9dtI2ROIQz6vSdnNHt7uFcxXt37BCZ4
ZXxtd4SdUdzI9zqb3XooSHJDxWU93xZm/iwb3Zj42gqRwl6bAxqMEhE54tsGdBJmZ83cycH63r7w
bQ5fgBg2L9AvY0nCeEYa/u7wZ+LqS7rOUH6xLroPBbJ/ghjwhiOS7ZOJ9n2Y5tne0Wa3MCA/t27s
LsCUvBz41rLQb5fYfOIqt4kMSrKg4TstIqnUQ+ROmeZk+BoSigidn7mMM0G4YtPXP/JSp/S5s4II
CxbRJLOv7oe5Cvj7fQK2TOmSOSDpXIrR/jJcfmD39bAQYFo1EqKKKuotQjUD2QKkR2NdiGo0LKqt
WcZhuRME+Zh4i1rWuxcl8wX6tPvRzeb03VBT7R7K9YSYWOuVldk2twgpL2k7VvGchPndF+g4jMTj
ZDbZbgGYANWIJ6atWqhh978jLmkT3v+40qdQuRKlkhcHrD4so/+finw1CqC5x3KFG1EAA442gcLF
VBR7YzwtJBGvQDJg7qkpSWVMld+16nHEz9tOmMAKwWqNcxhXLBZQAeNsvftLTp5IRZekJMfJSTY6
dRV7oflBLlDkwuIpMSw5G4HnO4s8AlvuhQvHAulNhD2knLf+8Hl1vvuRSX2xJVF1XEdVdNc1Ig4M
e7hwrwYEL+VsV3xi1DcDGO39ZpRrXmCPjHyFMZpw+iKrXV3Ypm0ryu+QbVUM4eKiU600TP7ei0zQ
l7bJgQuW7YkCOzdUVD5dkNI8CuUYljwfluyVoN+W9pzxCCaqEjABvEpBEQ2BNxAVF8X+8Q1E27Rg
H1pSHSu/U67/38ZZvB5sA+8yPGZcuKfFTCbbyS8yFFNEaL/6EE9d3uZ7Ud9W7TUbe0NcEqpzK0ZS
0BnM2h5wuJhpv0ybcexa1OLqxmZJHAZGrkrsoRajP8VLLCT4YhfUAqBG0uJw9S8sTkOCYn54vUp0
Lk1Np+pBVvp3vADLvQphor+JB21dnFR4DAwg4obCNdJoY/LKnqAeFn8yonlAWWGSzmi9zFotsW6x
uMiNRngjglBFjYhyceZiZ919eWgb6hL64O7SuV0hKvI01YIHWGKRasWYFoiZ+NzS0UQ8DntlXBtU
jGwg4bR1K+Abbk0r2otn+tH/jV5KR5EWYNfEeAUIEhMy5OxVxe2F+so6BZRUepWNstGesmOTK5z+
iH0kiNsHbPk4eH67Gt2XUEuYVXTLAKFPve2NA19JHR5gq+Ope3crcDzOT+OkmH3TXt+0JkcE0dIt
de4SDAl/ndDDgCubYdMBSVZd7/Rd5M7UFo/pl7rlyBLZxbtHmgcfT3YkDcgO6AHEk/l5Jt5rMKCg
0eoaTvmiQuh68BcypYGRJSRZWzalIIv4TVIYFXSmlKjhyhzpin+RHvzO6AE4Ws33YGyURsXpGDyP
3qAFDTqpH4mRh8TVj4lTYXDi7sQJL2SrWpsG/d5f9gZmqIodYtXmdv6rPPSecCny68LXJ6P4lK+v
bvqJZfrEe5ubBQr98magxDycbEc2nSuvdFU/5zGdv/6Ui5fzp4gzNW/IGqjSgasqd9/tFwTLoKmM
RSIRs4tKIOyJzIC+1wpNW4SifBej9Dj/A6McjkApx2N3u7+Vyv/ifRciuk7tF6HpvmURUnZHAxoz
IlZLuNrrj5TJadphARPZ2h8ueIqV519hJQxPXEpFd6wZxQunnjbybtjz0MrTwANJMMXvYPN3lpOd
db1AASexeWY2GCGeeu9Cxt5VjfNULaklbjLZHJ2K7yBHv0S+vOIHMxsz9vtyyQnEer7lAJ16aL0o
+Nj9Y+K65SGnGq/hzFIUq2KkxwAglpOXOmwSbtVU33FrinC96SaAJIgvLrUzD9ngNJZGyzCBvyrT
c7ZhT66WBgT0T0kc/WTeVoH0egm3me7iKHzJEO2869jLkrSZzTDxBxcCHN2ZRD3TxnyYaeeYf5rC
Xse2SrCYow8fvbLZmJNxbrVADd+muNE+26GUKAKZVE9G3PdJ0ds6EzZXVHLzmlv7l1vVUXd405Qj
mFKuiVMVRmuxtbQ4aCI5R3tB/a9F6FdWLs1dfQDrqJowJY0qjBKOkweworIGpH5OHCFmsss9p0bK
5vcbkfZeupSqKTtcxZgh/t1D1BxegsBC1ijy38VGroAwDElxtvRcU3RfcpfaHOQ66mp9Lda6qwSB
s+5/UD/63+tfgQ8iAvt1qdNaFHer0ZtIY2EggtaY7xrCubK/Jfp7WPg0IKVy/p2BNt0TG+jqUO0V
n0E6b4UT+zxKWgBlp+o4I/Z2iyApfkLNSJLM5ARcWsAHYEy8vJpkMFHdspggbq2PHUfemDGphYEh
hkVaLdgXFf2b+LoHF+d5iNoZfedUO9WRzVupFocvkXufmhLKR+oVMU2WzEF4QG2wmQ+zkZXmmWIc
EPVFVsC6OwQanxVtr8xcQvQFCPeDXObKN9JB/PZFhROxkEV95M32h/XKXE4iSsPUFkqSvi+AMIc0
VpFPbZiTAPLgnH4QAv65R4G1DPbJ3ssol+4Vnd2DeHUn6/eHeLio1BIcFpIbEQgkuAtvwZQsuyqT
SebiDkVw3gfzdqvORmGOc4uocoz5BEFH8SkvLRwGnpH3skBB2lYJrILwYIhr5SajzXPiWZjecERb
QYanydMXi1fl2MWz1JyAcqX28D+VQqiQ+yJiko8LvNEwY+BUNPjyp3PqVpf1N4pv2rcQOfGvTyzS
10R7Ogr6jy30LLudZMDIRZ8ueO2te5AEzNOreUv10gdZlbtODdI1NTAmtMNYHXkxbRjX/zhqKmoQ
VOmT3qVvD2phhFOds9cHuH+tL4FPYq4kWjhHdthhk+wb9TjpTMr30ywGXNHhCPkDMQs/YVpNTPSQ
pAK+MUzD/T11zPYHX1ICFIYQxRY9VAQ0ZW60rFDVEm5QK0XW3u9RzBB24nLEF03AhsQ2v3flo0zV
F1rHyWPpcPnROJYsvPtrRjlAZhFEVj/uTCR/sDWHx7KEI40TGHgcaF9symLmiChKGRCNr/7C1DPu
Udic87pymA7f26UBtyKV838L6OKN72YaBxdO0gz+QXN2lAvViLIW1NI/xH/ffwkgPSty0AiXiGIh
tW8Hsn1oJhHKfmaT1tIHTu93IrrTiTtGJQMVXR3hoLykUsu22iyUacEYFjQj4q5FUfq6vEEnSikq
wm8LT5TqJQJZFRa0rKvN4fmX0X1WE8/XjU1QEbccHvGl8Y2aeuznEVLEbdoNHZfZZ5g21KhXUct6
0gsiXeGoayl2BaF+7jCG4JGwMObtZE40pbTfJqhTh0rpY8mBxCrgaZnf46q3CKYgJOsw/bLnn9KU
43A+eOF6c4SFNyvE97DwtIDhH6P+37BrYLaxnEEIa2Lshin6I4oMsRBNVxKmYPzwszlvAOM6JusG
oolGmfXaKMOcnXr1Fhuyg2LL7xJmvJfAkA8msXa6XgmPLhE5kp8+8OvfoWJQ48ax5b6Hi1S2OeA7
cna8wuF/ECcEP/eV6fw6RkYpL+8RDz/pS/cC5EipVwCNmNRmS3fD/E+ESzsbOrmWlwJ1BAwDbE60
P/+G1Zf/IOF62t6vKEAaC/V5m2IBdeur3snrLMFcWQh6clpKVHXTZLWQglgnJIF3rXQh/oKpdFSr
Iz0j1dHCza19Airg4DTLXgmj4nTTateFrA44bXZFstITvA+P4/gsbRLLurgv4vG6FUmlKIwCb0nu
qrAwAfbYixveQi+BnvGVkela2oVLKtRCutF6GXzRci3dQZYPE1ipXkAs5JfFKCAeMtznrbvR6Udm
u8f9UB2umzqt2pRJ4kQtm/BlPcitOyx8G6IjF5M314CCx6mowvVKh1ThT3GY+vOTNDz+dXUZdKtJ
yrJ42pF5mZkM0Sci08M6wDIlwoV0IRXrGy1FABF6Z6SvYWEjztaLDIwybnv1zHgjzF+Q0Xiz0WuC
Btqn7ZVETZcYD9Or0nq8QpwIby0TgLlmKCvVj+Qh+lxotaM8/yNcN3mPRyQgI8UxwavVoe9dQnia
pb0Os/dHOt65tg9DqiWC2arZmvPfJvatFvBFfDL7OVVAKen3Cy+H0y1mbIOl3EtvojOCg+fCiBlv
rgfl+WIWoNxFpIJgge0mN9hy98KHP1c3RqYrYQYtFZHR5VObihYOR/Z+o0MRZddsW0iFV+xiSaIG
tMyxMThENnNpHzFzjOJ+SZitK0odlqVHQM0Lziact0XsxJwpDzTZAmlbFpBuntquh1+3aKW8V7Ac
4zP3XuCUSxwculjOMApVQMfp4r3aJhUiCYMUItGqVGt8gMPZUbrQbHC3xiZEUlnlGRA8Yqoiootq
GScuwyWUHqFpQDqIXitAlxo3l2HoD8VQxiDhVFtU6L08cX2ij7wj2Et5bmdQg+Vbra6GtHl5y8hI
JJiFgPStBruxN7jzbcy410KOaJdrZ79HwtUuyCRBb432FghRyWi7WtpyCvXIaM2Ly7zO8DHJgQGj
+9TxEg3M3WwX1/lvxCUDJjhG3CSp5U306wroqazivG+IGy6HR4hYvOVD/CS68SDdb/dSFIZbB70S
4IQ0nPrl5pEbGVpt74VYodV4kmt5q9hSgTpuJb+7YeWfLKLqgeJrFXiOvXyneCGS93BSawy3RPkW
aqpL6R+pEX2q4i4AIOZvtOWa1D5vU3VpFarACpIpvgUuCt4pHd3Z6SswV6BUk+OTbWXaWkYss2P1
W0yi9OU8DEYXomUlBvHOf5hUMbY249yzc4GVfHc01rr+GnTJLlN/awcgQ2CRWmVlk4iGZYJ+Cwb4
By6A8FKjiYTaa3IK/jZOWZNGx1Fl63ckjA8d/WCar24po4XSaY0jWVqpahEkRGY8TILc6sCVpjzF
FHp9g6XmPU/Zmxzb0Rjyn5X46Eb1F/GUysOh42CPj/cHP2PSRDk7/tksbigeeh695CRy0PLG6CBS
9fjqRTctpPDKUjvswW+lOlsWmBObfYkVARSk8ioStGL+1gmIFgWbl/96C9tbMViyfphq3Gaaf36Z
Ey0cMtvLiJ8ey2qvEYs4OXhuThE6PXcfWrzJuvqIR2QelPAi1x8h5ZhRrpARQev0QAXGISnHi0Y/
79W0Pz5w2bWGSlOnNfOYxU86pSAErC4yhJheq7lT82jxD+lGvper+G+yZReZj1b0VCw5Nj31oDuU
PmerlkyzEjEn46Pg2ayNKHtSq+++HnWQkTbuZj2NDI+lpByhkKKv2PCP/ArKPIerppFIkBkdLXy8
HXCQ4+ZMJ916bCuWo5DaEb/dNpy5Gm6nugYJb41m7zFU3mX3A4ypjjfxVe/U78Yg5E3pxecxLGiR
UvSpEGs3wpj49NnE+iJUZBf/fu5V5jK7UAHSYrlPBo+xnQbu+vmRVspxYa2DCQgCu/yOO5IW0wFn
2BJXHfj8ONRvNxMMK1PWYPKpXTrDwdzsKjWJJqx/fEFUgGbDCNrVrjQ8BqBtiEVGnH9ola3Sj73J
dpOaGEMrZQaBFWGyTaCUiSWyFIVIWbVoD/bgtEfCegVFE2OwZaOwAz2yFkHMJrLtQIZREWHgoelF
nNL2x4F02PbEWNYYQk7mk0kNKO+KhccWrVZTZ8GtQnDvaSQ4wuuRIoBCDmgycwpBylV5O3kIu7cT
0ytwQHeF533l3RDCh3mP1FBZNekROsrwFqPjoy5jESfGeS9Y/JrdpvWVRUOzBxSW9deJid8SDkNa
uXEpGLBtEZweddBGZmyfzzZQazLYa3XEU3tBX2cqTR+S7S05xN2v5Hq0+UyDQtNgSlPKkVq0KOfx
MhP9/Z/yEmxBUCGonN4q0IfzIgEeuwdk7RBB/6K82500TubSyeysA37NBlazaMwZA1D5/L81FbG4
9e6gYtms7UT8rbgSSKcut0Y7fCPjrb65UBqO07zX01R7+SbiL3xn3COoyBbZ1HwiKm8Jpt2s3Xqg
3t9lwM2XHdUD3XCT8btfbbFXbA1yKoLAwtr8iqsMRxfSeWE3Pb1qzz0VPh6lA5HRV0yGTtmZGMBk
nD0KOjBtKyF7U2BGxeb7WpvEFbJ2IwQlA1BQFwNE1WSmbLN5FegGbglhaaYzpESc8ER4gjo/r5WO
PZIGhk1VDpjXGUxB4eMWLcNLWNSnKfEOslGHhWASXWOl0KE9oU8jz4PQABsDCNGtetuHnCaWkyNj
K6gz2CK5z/4onf9DidQX8PqCnro0yUw79o2cmF6/HO8AB//uHdSR0NQ4DXUn6xPvOZ/OAN7NSP9b
3YqWnD4QL8sjvweHm8BZr/dUav3NCAm7fGpCK0f38Y9c5hkJwncN3SeL4iexvriU+JkLb6ZD+7BG
YIpXWI67jaXJoN7PObO6LDuaye2RK0hIrni0P4iv+j720hq3JV5dtuZe97QfZ6zXfXUzFVv4kFWf
1/GAswRaF+6CC5sJb0f4QFmY7OjyApvlHLisG7Ca401cuujeDDxxzqI1UnCVdBWYyqscorLPEDaO
M3d2XLqFdqQHiywUAozDEI5UTD29yKDs4fPAM2dJa0TS7baW/Pcs/1lKC+ULMoUk0guLdad1C+Yd
9fJmtrO7sopN3Kv9L/spzIPFIPGFtGZ0P71twm6bUWz3mbkPj/FpVM4lN5gtk12gK5vOYexHdGeu
dQrFVj1AQEJpnzYS1gUiHJodWJ5iH4WxMP2zZ8eP6Qgtq8pPX8LtTVxXjzuM4xAlLfjuBZ86gw+W
o6nOX6PP3KjHGZ3eq2hR255X7uTIT7mAXHOjvA7t+E8j1u0dlePXAna8l0MfKmeXwQIh/nO76SmJ
bk0K5FGGOJCRTwJxTv5zjQ0/J18+bV6f8ou1MT3+pqIFbj+Fud/gWpNzTS/KPbqmyVMQzXQ9kxKu
ZN/HmrxJEMiGvETDQm7350J1ynbDe3CynKZOFt4z305BD9j4XRDIpTw9ejOwsbEKSkdcESS1kZyl
FUmBZNwXpSvAKTAfY3Q1Pmf0qLBRT1FGOEjStK/FFFsd9nkKL9N0vPiwxwP9EcmMANo5yMCgeOns
nNxBEa0lIqErUN9jA98YW3rQQ4bKyKfnhU+/ws6EXdxABOGPPdE5nSgF9q2VTbUHueJaAWn98qHp
lF81TI157hlEX7thf2FD7hZE2d574DorOXvowo1oh0crmdgUeQaMBOFv/35tdmEFEyrE7pFsIbTJ
e+kCo0b7HJJDOShtL7sIblgG2XL36zt3Pv5lUymIag6daZ4yFlKxPYhZOm6SV4XK8O5fXeeKgT89
kqWFOa9VCNSA76Fmu4G7fG80EfLaytjmMPf+mVLheYgE8sXtv6QpMB0kKomPbu/fMRX/noqnDHLA
Ynd7gW7Bkj7aiIGLjYapJniZZA5SPuMbWTWLW4LGUxNnc5Hks3vqfrzjywWWhoFoUibetuFnlNdI
0fZDAaayKS/6ZgDOwBD6ODZhzZhnLDXwlJ+i6QmdC1qZ7TYtriOe6EzpY6g0oZT6ltYssBLzt/bi
826PC0EvQA7DIDCluHYzNgxE2XxWPSsrkmSM1RYDhfL3RZyWtW5XhIdRYnWvaWsicwU1OPWvWSqq
vykL9EvQrigTet1ercsTQ8iqyNrSTpsaKulZyQiTWIBmsbEMKEyRA7o2HxrzfKs4zwMWdNYA6YLK
WKcQLHz1X/ZQlHKV2MQjqnTrknCgArATQXyBQFWJZBDYOjjWqAlMJbWIxhYzn7kQr1Fa6Ci+wZmS
4FLuOMb9zFGetuGtGFpmapXutETq6byWYtpCZD7lKJ5V8Kc+iYtwdkCeZSzeuwMiEoSaw905FGFY
Cb524pwmOr66xaJbx913+p+wP8oOD1C6V+JJ547bYt7ZDIQb+olVHZQXE431DNUqXNuN3kHkAQNP
KC8RI0IOatIEek9+eX9lMl/PMhg4Q+yGsx/U15/ATLudvxhJor3ABVPiDOovQ/4wcS513LcCxYFH
EPK9sI8Ea1Ww0fyn6HZd8lotf1ItXcSCIBvrocLfKl5PuA5rLdstRsR238ixm1ajo8SSflGGn7T1
27fVHHVqG+c8UOxakhq9cEavRRt1I7s+5mLo78VadjmKyL9uAmrrUQInNWR2Q9ofaHQIzO4VoYUp
JZ1holwXpynwMvX9LJ8EagLgWHDkUxddskst0idh3NVZO01lg/eLPUTn9TW/FzQSszqBvmmnZNva
u6TpE5ofpsR5gYu8qImiK7cV3OmY/yWX1WRnLjFwTjq2DE2XJDIPHLLMFmgdTUjqXsAjk86bIIcZ
geba8oppOEUJxQfWceLT+SIYFVZZyFxAmrLeDIURQdAItYGea2SJOLyQtjz5BabBIWwteh5gfEQ1
HTX3f0l805E1EkwRNGTnnqhLGxV6yrRabS9Zn/53nQx9jSHqPVYwjMVAVgbufOCAVpOJVYpLVz5T
WrTp4ioHCzcSMjOg9LM5ecVNwdEh278aSyEM5yuoGEMJ5nLwYHdjE6Bo1DS1wE5tNHnqVmznyf7J
x7mnZOrAhrQYpv124hQ+z2RN8LroxHRvy0N1NhBT5dUkVEjLfjmGfGkUX7McLdBNZcVkiQMTVGol
jhGjzvw0a9O/W0LWgTcMzJqMML8YiK5IJM/QomIfhReXB1GkYxU8zwxUpQ1nBxXC55qrwa2/Vovv
RbEtl1jWYevIKa5rO/XvXJZSSQnWgN1ADjXY+1gfvRWhPiTX3Wjc53FueTlVywvkm+X/uQsMlOnF
R/rrKzlMZVvFVAsMf83DGM6YtpqRrKtyIo3ETdmg54dtKhJ4rrZsSQE2uh2LuW7TiqHjzWFkmPWw
lna36tOZFodsOxELlZcOfF6BCujHMrtvR8l4GOa0yaOFtXH+5nXuEe9LD9gfNU2+WvQ6V/jlBWXD
Qf3VVTw55G61eCJ4Ru6AHXhbAEDDrJvBel7UHJrqc0PWub3w91JPj7Gbuk7CWhrcdp8HEXQLEv+M
hLlbO3gFZO2TG9S6gKkP5oRlyicxD2mYzF36PXX2MLdppZb7JFj+Hk1R3razI/4qd3bBfxFLUpin
qCOetjhmWm5nKqd79OUxOpO4ZKpxHdFOI1XSCAdyIlAD9OM/RZj0RUKl+nrzQshdp6yY8UAWHzw+
faU8+BxT5xH2uu81HGf3kKgFZW+/bZwHVgmbFJn59y0JxFd0Eri24nRfq+g0TKzewnaGpJ9hTHWw
HZbd6LUhj+gqun9C721ozKYzxqg7I0Amt/w3dwVh+FjJ95Rw+uxFVoe49TFe01Mk9XL5QdB97I/B
OqZzuBRA9WMq0rnHIYo3a7Olx/YLpSqPzbLqmqN64lIVQVW/+y85t7jpmriojjBHHTKXwHpk5rgX
6cbH2yZW2UZJ22pIhBmpdz0GLiPXqoU5WldYl+F+O5koK1hvBUetWMvkwl9p/TCApKX5s2DR3B7J
bxv0dhbI9qz7WdEcMns1vT4DtCWuvmrj1HUdfCOba0lrunUBvpyRC7qHE1h5TismV4gwSqT4ZfM3
aGiQuPQZ6FI0nzF8kRwp/s546nJyiAj+OpEhxSuYn046KJdVCaEPiSS3kIlU9eL7ilvzzZZJTth2
VvYAZDlnSL74lbjVnunFMMjr6cqq48wNr5OPGBWdqqG2c/cwdMOse9dmQhaXR03oqb2XBiaztXCe
1MhRAuoYsXorV5amS4Y1eitOUIQ8MS5E+K0eda+nRssg89Fz5fl857Pl7AKG/DDrhaJd9Er8Ynzm
DqPa4t573OYvySAHsoX5HEDLqOA82FUnlBxWhcKgs7AlMkxMivYt/Qv+dfzza2fpb/U1CQHV5dWD
f9w3dTD48H7FRbu3cdL0UyyJDrriNCPlckudyKSFB5YXCGuMu4/Zt8sUgvJL3oQy7YvCh4pejPZD
dMN2yT5sXmX6SbuHfXVRV0M0e7kJTVR083+DIufMX+77svOsygEnueqM1n5JDXPQchQcFXO8PX+M
5eqdCyLK6ozfqzGrYvrwZwm0zABTdA+t6DVvhmVrQ5KBqD+mwuECJeT5hsH9zXJt0Oj94zjYDW+l
krPh01hwt4z1RgLunsufBucSvI2jItn2jvslWi1OUjqPpXgcbs1J8rM0L7gYF+4C2na1BZNU/Nhf
rGgpyBHMy7DTuU4ILrJjA41t7isqA5szwITNIbiOTKvSxWIE55+m30sT4U6cYMN1p19DTd4G6P7n
DPBV0idNvKiubidrGJPrTRPM9J0MC0QJzvhuZJeEsqpJUoK5aHhOiLWi73045zsfqRfhO87FLJ2h
4fCeZS/hfN7ikXqIK/lIVeRb1xi4MJ6hfqQALTVlAsJ9QCuOiKU5BqZm9Miz2ynJp5J7tDAXo297
oRL2SF6kGnNOeTjD4HU6Nr5tmUL4ErGzqzOqVUYH/wlEcd2VmMD77gH7k+x+XiZ0PJ+P+ty0RYJF
lXVEmrPmepu87UzEgvdLsnNtZwGHpZe/4nD5A+rqCA1zY4eTEFBNC7Wo+5xn63StTIuQ7o+tnFO+
LEIGXrDLIMfqjTmmIOmY0JqWicFbahS48pQzLz7Xp+DFlh/+pEtsuwXyOqo1t+NWMzb/bZfjyZHn
d4+jxqO9XN3E+kC4rGkCj2lG19CrhAdKoisH9Y+DcRujp34bdRehnU2nT3rhSgwHsIhRZ4igGub2
JV0XOpAO2Jp3hMleNnBQKsJoTki6Ph4eLhCTCIGXqp67qdl0L2oF9HJlUvgjsx2JP/fj3XeLSCZ9
VTuk+Pu2mClx/Qbqm3PPlKo4DR/XTEcw+/7xsigXAfdTag4lGOGTYoQIl2sT9gTYaETzqLUzgUtY
JNjG7iVbhj2WSbT2l+AqAQB3abjirncb0tkN0rw6zKiPlGeMR+njrwj4TmPF7zlmnnh3xrqAfDVm
78/DbkjWVY3jFTXtUQ43wyNSr+YFHbpHjVcw8GfMIKMdhMpWSyHGoTu8ls5R7y/uZHbHZQLce6ZR
JRvwkQs/8MghrUEdM/D99a1xtNId2EYH40PR+Mpw2sGdiCDo3iFJABoO7NuEIWSmPCyC2NWRtqDZ
wG4Flk0f3Zf55xPSDqCfabRoWxVmrDki6iqW3WYmUeisrgH9TEHBgAFtx2YTONfZAB3jvEE9Zrdi
l+upL6nP8UuYANyuMATvnXzmEkreZjVWVCgy1/Bq0QXLxHRprTbeXQL/VW5XZnPe/i3ToB04kJmb
M9rOv/aQQ2TWx74QRq5tE/xJkdGKmjdKcT9CEyr75/MMP2ZxkIr7ZSKfpInSzF+cj/Ra9E8zR8Iy
J4MeQwaChYN1ijWhf5ClvQEPzVPLT+rdcWldgsVhu0iNi2z/kmnWEONLJkgw1utQinBSX70jhzaI
70VT7DrOBtDo429u/7eQMUxcQ9VfcG2ZiIZFQDJIeJvfc0js4DfDiKqVi14yOM7DIRlIGWbtwa2I
laP12iPCPNqcpmoIKzE0hgoYAuADKsq4s729Her89qrJDdfElrGnJ+AB38SAE8pSfG6/Iyowl41x
4Us+AowXmEPM4FUZvhz3itK4OHqxIBjmkbgjbhZY02lEmRaxz1dGMFX2td0y77BFVyEjZn4BBjNW
tkyR0uDecHDjBc1XFb25/O7KSiya2p1lWpkdSxMRK8vuezWNKSJYfpYYaYs0vcCfDjhqDyQx0ggQ
PvJoDCTn08Qg+dMUSJdjs3oClsYDDGJBQJV57tWakaLWSROzdf0KnXSC+p/exW1Z5ZW4dh9oRrX3
P4f/EKMogJvU+1cqykxg+NaCj802Lmk1P/ybLFJZTveHP91JCJCPnLLdIOs8McXAp3MOqzY/SD7H
caxSu6qhxkDVI2DkU5XPzd8cf3zTLy08l3fu91mAvzEmmYSmyPMF5AtFXjjaADuDAWRVCJbq5052
+aL9AIcYXuFhorSfdP7W2VAhWI4lqu7B5AMmvaAHMjSaTEnzIhGJ/8M6e9EylnwOdUj7NdubLRSt
gua4UdnUwOtfOgd/lbjmG40e4bYYf29p8+9/8mwMYbzSRxu3L/9SJw3Hf8ko9XT/1VdmdSBVRrkz
5IYp0UigEdpo+eP+/MByWiPHLim/GJwgkrqZHWAQ3ogWKlkdOhAbBVoIdQPlZxKWfbNhx98L2MB7
AgCpJiiWAd5Nv8oLZOAqdOzTTx5yak1ep+3uy5FPyOt9IQWH+BpoG/dSawVrPusJjfZR816IZ9j5
ExP3J8IbwM8hXRUpUQORi5TfrgG5kUeROZsDm5LbI7wUJ1R/X8AIWC3YaYVXMCrajGZj5sIzFW6G
ha2Wqkeieh45yoYhFBCEwU6zR9+46v5hRwjJ3y5v3pMSTURoJ8ZTLIg1HXbQggRL44af2cdjLtsg
38DQDWQTQgLaCx+HOhNTRJMw0V0ZgAaDYw2aup47Fcs98bZUh93wL7AUC2im1X4w8xnlszmRMHAX
WFExpLFNxxigAQg7kxLEndmoMqi2A3hpSrGocM6Uet0qH1AdT+Utjmu9WIGkjCf7kU9ixZ152RUn
ihU1gMOayJQBfPj9d6SZZ11+VlZkGwaf86sEu02f1VDyS2EKuEx8bYea5FFPBW1m5g7PviQd3PdV
u3IO7eYsACSA8F1ZLqvkeHGBYr0JC6Tg8eTgJdMm5wEo7Z0yF1VqXhLdu5bIxK7PSvX0+J2Wt5Hc
l06wSLshlj2fz3TJk3sQ6kotDA7qXj/Up7vWel7kNZ38dwiZSb7GC7cq3f1Ktl3HtYOvMR+AUyen
YHJkoWdbfs9n9U9w+vLdnMjQ7ivaWbZjGGbrAd10JrvOMh96iM4G5I5svK7LsllqZaBIm+8hB4WV
5hi1GLAVW5HaK0k8+Qua8HLos2aa6JyJuJkXXrDetaHH/xlng/2Z+9q2xIgi8DYDUWs/EB4FeF+S
NVnYWgr4sIXexIm8kMcgfGslADBa1LNn32bl8+CskHnIRex5Jgg8AIrn0LYkNTGyV2nSSH5imUos
sU3bh2Uxdx8MXlwLWXc6Qxw6fq5KyF9Xb3E+lyyuNvolMHXRGI/eimT1JDX9m/zICFXEGGPnXjXE
Im38hW43HNI6XUJMupenVWtWtrDeSqrNz3cS5C4pGMl/Zii4SnHBVMfbR77Sfv/zULZaMgCxE761
2/Mtctpi323mk5fvs+QMueMgBwcFuBQsUWdbXQIKRYpkH39OGeGvgj5idlg5qPPrBEa/QFNj//Hg
jpC+O6BIJsSsxJk1bBNK9rYlvjbze99+DictwA6Diho8RlO0zRhaSctQ3n7UrJTYZrGaI06CDah5
7jDA2yikLfXPdMTzYKULZPPQZNL/gDPU7YYuXuSV2Ppla7pOUKolpxTmEyiop36F9miH2n6RSc60
wFddzjBldvQC8yV9PTP1QmVjjeOw9yOuR6cwfGjJBRGFZK+9OVZ31bkUCUnjLZppNep8H2aMgFvW
6FvxC/v+/gbJjoxcVMES5yAg7gLoisfd2gICHZ4WU75DEJfmFfiZuFTictiTjtrJPCsToWxeQSEy
d0QgPp0lP9cq8aPQSbu3j75fVIiueS1DzFfL3U4VbEd4hUS0L1bPXZirimiwFwGCNAhTQUQkjjbe
qx6VuVeVxxBPHdzk2Y35imYfuqATHjIA80Aad8dAaulN4fQBXOeY6Ppp7Yz6bbUlU5WRh6SQ+qgD
jFkGFZa7eaP6avTGZR5nhqvArIdaEh1+26ujDuu/aYqGmWLQxlo1NRhmblTKbecRSwUwSDTJNWZk
uwnOiF+qiPN4w446IbjeDuPnpMrBDXzCgNFkxho9Y+Wczd9VSSzR0dTtgJSUwixfN5Y4qAkGyiWq
E1gBIAh32mDRSqoOYoGBGsYs8yW+TSJAO5WkMnuXIG8u50GWz8xegvvNjm3Z/Ryv94MptGK7eu7t
Pno00bPqIxTGRIQaQw59d7lUlXujn5CkTUXI30TSBftXPspz6nhlY7YgCgiEu2s5b2VM8y3rCngA
KIphXXvOC2AqTV4mjRfQG7dcKnG9+zX0RcIGy4cvEc6M4d9aGeblypZ7BVwn+e3XJWUrlmPxQdBA
4IqJm1uMwsS2oA4+8wwRXfYp+ueNc9894CBekHgJgpbttFxIrvCvGS9yOgqh+tAcXc5wRuc2olBb
9yCQV337I7J9cEPVGnlqZwawHOJ8lLQHPP4U4LNQb+OoEwkr50jkiJRxtpev0VgxTgv+GJXDYvjg
98lGG1PPpdzG6Dfp5rI5A7jvIritu0WzrcdnU6yVA9LzDueHJ8DgXsoJBhnb2BEmhcOtfOesQcDV
NbkRlF3MLE/a+bJxmmI9bWphYz3cPvjg0pvUYY9OTvxdlesxhqWCAyCyfuxUhiRbbZzDlkLZYDBt
QS5b5WWTPqimfzq3dzRsVjntY2/fVL6ky0EJbFWdzu7CqW9rCyzUW5FiIS3OAUa8dVHAxgXcJTM+
ikZ2BlpVnZr2eOc2zgONl9CjML8aWnv5rABY7jm1boJUWGapxkKCOm3nWf3T1PmyA9FKiI0lkgdM
3sB1TdLEyVLfogOK9gR7NGoOb/bSG0DB/XSeWJG3Lw8SmXqnRurlzWDWDnopii7i2YX5n4IZpzMm
VngHD29ATJxIWLMALr6Hgaya4eOkH0YqZR8tT4CKMiJRTX7FoF9mFVHfCQNls4bWaa4xEabY1HNY
8SAY7LpCH0gjztTIJZ1GVwJl770/Vu258nHm1RvQtpJLGUSgXd57aG34GSOG/GrbuqkKXcamvF3e
wJTsSh+nFNc/Ih0ZsVuejNT/6pJSaWnZ6F+8DAcKb7IKtksLoWxHksLIuGtzVFCbJu0khi5mxfcH
cURZ4CLydQ4V6WgF6cVgINA/ezqTKBLcX3rMWoZfS5afC+8iGvMu46TlT/oOoDLr6AD0orE6IBOv
vvuTRwNlX1R/iCHi86UwZVjiv7es/FWfnS6lZk+6442WPOGHZ/p0dDraw/UKeY+KKyixCHlu2FPU
vJc09g7btTgwPiVNmivvftQT/mRiafSnaAvglA7aE3sJkbDt22O6nhnHyDsH6DkivhH3cpRubav2
0Zg6JZOtlrNDq4Y0TR5yi42HHiOjpyhSuM9rO/nW4ptuH7BihSWYK3TfuZzydDsLfmDg5bYyV/lp
pbK1oIviVXIR6PXDZrF93UqHpFiKsc6M+LipE/WnanmHKOq7Fv+vjMLec+FVVhy6N2L7VFtKRqxt
P9mcOrhRJRdEQte3TQdux8iAhvTUwMVfJJez7lD9jq1TvqC9bH9cyIsm8vB7pIyXiONO9ufB8ksM
BmuzfogxAqhAgxHgPiu6+BtgZXC0nWRh+Mex8QwcywGojJJ0SXLUu3EsUksZ00Q4CTzIqflldsv8
Bz2d6zYajN+KSrmJcYByLy2bveIQVtIPuDAf0fnxmVm0LvA4YbtVlvqMcbf+fQMEyLR/ujLLBk/9
D27GwpfJJ9d+pO1seVjB3WQNVkuSr+Rdkf3hrxYcSqFn8Xzpzxegkrz3uyLJqfkWEI//EcnfVP5Y
yfdf/Ck+YOenTYHGV9F4JB9pZVwLPU2S23MaqpqOQIa9R/wfxexQ6VJImk4bv4vdKd+p0ZAqxp3o
5I2GF7daj5V7DWYMwaqp1/9yDxt59Ivpdd1y/Lsw+6ZVhhBBDghjd5OoACsb5MNVaZbWu/XyieNv
9TUxqhjsDSfFLQL53nOwKemIGb1KcMdEvQciGR1iX89XAB3BJ5Q36Y3VolAVsCdtBqlAvT6vhZRW
cqMNis+fUwfCZosO/2h1Tpc6hnwEGCpqru+oyv93eH53XAV94ugrjmH47qJCFGD/N9DKpHGtr+I3
1Q9xpfb/lONo4J3Qe5FVaXSlNFC7EOiRq/IK53dTeX4G4LJdGIgdNqnhbfZwtLVeSqOE24GC0bVw
Dp08ptCqBP+Mif4tqMjuZV+xshy24gsyBMcWUwnVUY5eg8hTiVXhdj7TtWHuYBCBbv2nJhsZv7G8
EwJ34i2rCTCT9qcFGv2HfMf5JqaXoympxkurtDxo0G6J6r2TPoKjOu+M3qB0+E/VJzo3Mybu1cVH
XBgfrpb6ZSg213j4gCC2Y2lFj+l7Z784XCAaaS0HE01gpwojFCm0BWPm0MmXmkEsjuVZyzpF4Qxp
diwqmMucolUb0VCqtHveOt2U5iLp+8DjAs2O+HbNZUKkZEt0FJvOEN7h1UIaoIkHbvgJoyPeoyFJ
AxzQ8hAdfh1v5n9jpEuUyetviweX2c1jljyT6Kdi4AV/woxBcav+qofsl7nuEc7ma5G1PjQFUPNI
spcdCd+5+a1/DvjBlXVoEaYw51d1EGu2A/fvv6tAkCaJllZwNZEwIrn2jsw750zynqvbeXZVm31A
2iLeHUZMYCeSM7M/LUs4c9lbKeqccgkDLOOqmOxopGG5fr6CSx+4ZTSaMXB619EAV0XM1GyFTpXB
MuIkseKdm94KCmQRUJb/UxhzZNn2JzQD7JHuVzhJCQ9MH6Ssu7CFhAlOCHm8PMQ6R54qL3fh1LU1
z7zqPgpiBZb2GRMQdihtYpH3ChYoUcWqd61GdVHq+5bOYfXPmf/tIfDxvc/hzTwajYIvNfASw4U7
uNIiqYGPFGH4+vxUb7D4MGGq1gsLRuhumFsOHEPGhn2hskbDEbAwHpj1sSp7EPI2PF+kGFC04zAE
0vPsYyaCJ35uofB+iNDo1UJLuuDXf687pdVz3IlfVE0YOLsi9QJzYAgQ3j79PkPG0hK1aOyVZCwZ
C8T5ECNiX/GjgtQ6o10AYED0avKDaml/5H/Lc6eeRKw1ndZMQV+Ut4wPyLhZ+NEB4s8CaDGbY4DY
Zy54ahxKLUulc3i+Ev/aibacH0AsPpXug8+/g637duZlmTNjz9tT+hyXCw57V1D4TaJzNQ+H0Znz
BekI02R6cGg/rTqLKuV9UFjZ0+hNbiG5NlAd9ZQIQzJHzTZTW0agHDzg6Nc/jfmYyTTIjWGjMaep
1xRxDgeUWfn3lVkg1q6snuOqmGYkOHKT8e9/psQDdd/HpgtSXSQ6QlrXIqOqOu8OKu8CIfDYMFz/
GejypyAvozgja4e7rtYsCk8eMldjGlQwP55lcmsmP8G7E68GS/sFDzp37Ts9jRHEs7wUjEAkZy7B
Y6hEhn5dm/9cBhCXkAYMV4q41ks9qQ1jSed8Q/+Q3VSn8Z0XCWcLABwDIStJ604kYY4umJuqH7B6
a47yA6/ZciDrHPFf8whfo1jXq7vz8sm8TbDK3GXs5jcAzWMC4sgKyLu3CwWlPg0aFEaoDIR1yVlI
oq/AykP8f0mmuvFKGEPBC3iTJIwy52cpJTwtvlMt01Wim+Prv4w6+AtnaAYJDPK4Q/9aT8I+u6P9
jQq4P8bJvt0SdD09TcOKi73oyO9jMdY489nGDa3C81jDaHhlRJLbLeKUvMnFzAWSYo8cR3feXEMJ
6u588m1ERhaJVK0MWou6KA1vq4sv57JEEtMem3GbqfOAtrOCapFD6/G3LJ/rMIeoNuOEnxpf4lsR
WMUEJ1aschng8Jhb3xGyhxGcBjZZTgF2c7dOIKqgigDGc551rGT1n96ATrF1wmzM0ANCXqFi+jlF
5PuFKDNmNY21cChLpO1EdFZRR7k4tOwst+J70QFQZ39iyQH9px854Bt3pPZZXwKZpFuuMbAVL0zm
dChCIzJeybh7K7TB/dTIzyCHpPPKJkTF1rH1PhXNud8I0vu2vG7ppZCY4AMEQUnomLiaVFN8GL7F
eeg+/M9JIy8Dll6cLKQU9YkR7/HT4WhKdOYp0Q+DoRjkqgRRabm+x/MZSzri0Kinej7vegjZXTDW
SmUHuQM+xaTScGwZzzSa6dC8tk9UwR9jZl8tOZtAQcQ0zXJGVCWhI2nmu0In1oBG/W4mb6FjrmpQ
x3VazU6qpuwZOOTC17aM+Bu/Sdyz5CcMEdYxA2wtqKvo/hjxXLoKLa3fpWlYkJDnjvsQwr+c/bQ+
VBTeNy+eqSJ+MDQsSa6f4gaan6ZQqGZ4Lb6/QTjIpkEHSVRi9/lRjGJTIdbjXKHQ32+T0Pvqho5+
le+NV61hkZVUh2Pp+6GSsOtQso44Ws7duiLqfn2TGGVIBMVKTW7yMRNpAGe2E9bNn9g8MPkf34rT
f5MfmrL6b6Rqm4XiF6dE4rFP8Zn/A8JEZUmaxNBZiEow+oOHDwQD76hSUPjo1Q82L22SXPD/PwXg
AsvTxi9YFAehpo9ZOM5XNSBr+AB0yt+em7LdRCX9DcBwVVzc/+ede1koTKlg64U7wzEcT7fgUmW9
HoCBx1qlnkpfBz1791GFn9XHSOg8ZotseuLuhv41QZUmjV/Ga68HCtdiXKyimvhXQZW10Aw2nEQe
7yIaLZy0O4A+3lQFGvPCuDS1jifTcPXVAshDq5aVLjfwAnXLvztFxKFLp8Y7UJ/wvbYYUnLLkQN5
rvIWa+0MFHZKoU1jFDVLqTZh8nFQX+S/jZw/075SFdhL1Dk+O5NrwUUiCCU08QhB8nNaj0t1nzZx
keL56dJ9zUGcBae2cA7UY5PsiT51WuBGFW1p/L4128Mrjq5bGLXJJWm0kFeSQVLoyKFmx0CF8iYh
HaC75RUGIaRVNfIGxnne1jOaSPT76lMfbQAO2FeyZIZdhyEIF1ieG6R9h/fhQUgpzZPleqzPRIdF
4drhRMKPPUWskizH5g5k99asEUsaacV+E1fxl1eRFdQoz9wD4bjROM41VGtWAf8yMIdhV5MjubN0
b+9ydZU5GYi+a+vndPYa4KEAGykGOT5hIFQs74ii2jsrjzGmsrx5l7kdh+GOqODgiik6G66zrnAV
QfEGHOikKQ3lFHsY2ckAvIQTLBcZZJQG40+Awf2F3KBUto0mo144gevV1sgpfr6kQ8Aq2ccSu4RP
rF65lo5ZG7WKXiJezCjJikr6wVHahUDaI4frFb1z7CBwIEDlkgwAv9XG2KwAnDw0JaZEg6khtfW2
a/PH+LtZSuEe8FpP6Mvf7JeheB4spGFx3ijJRmhddf/LADysqBFntXUMNkkC0Wo0Gxf9WcyJZOCy
yK+iQ0hJkhL8jejgBXZKqv827Av+rsWH7DpFD7K/wOFDCurtRo0D0VHB8OedF091h3boFlSO9d90
PAPSZ9gA+tc7N6uRc9cA7RFSpz45HuxakZMfY56+2xIB8BAOoC04rgI2A6jA+tqZGgKC2YCMryYM
k6bYnNfU5IVvpELi/y00WReJKR+Ep0WEk0R7h4GqPwrCB7CGcjsiIlS4dOVAaNpSZyH1gZFidTM1
wKfUP9FT26A0GzT2Z7cHgut1aNUIcR7puR/ou/spE6j/iDeyebx/s/FY8yvGDAbyV6k4sNJnqPMW
Hm42f5jTvQ5nStQ/+BHicEvQGeCVA7AUO3BhdFgepFB4PHpoDJlUoaEyLjX42MLA40YQg3DN4fUF
mJ8+waMq/YId7kiqdemTCcpmeNNGqMGemAMsLK10iSi2Xw4iqWB6e9AHGmqJuVWItrbZ1Ov46S7T
iNedWCgw1bZZ9Em4OOOV97g544llqBjECh+TxI8irSmoeSDZs5o8rz/KF/AXomtXEaa3v5jKw5nq
GNmQ+pccHKcBAIRs6i/8S1f6k7oIizHJx6sJGvDPbyPP24bjsxlu8tb+dMEyW9u1S8cj8lHM7KXD
AxS4GiFi6qt0+pKK666DWEYYCCpzD2BBsgrZHz6UHcqU2Lf+ly9/d9CMDXmaYpY+sX3tBwi21I3P
WwKuHcrQYPw9kSCRHiINlBic1wLDMdx9ddxS4BFzHxGDc8FUAD9QOfIDTmmoUM3PHRYae8wlBSMy
vWDUFjvq9/RSnp6Rn905vlSLPMNeDMihbrSpQihnL3S4ozu3IT+NULa2JUJnuzqQWkfA/QDaHd0N
91zDDhvUOUjvzpe63DQA8QP/vsl6CE8Xj9ZRyBAFL0RJ4dOsTnVm5DRaFM1iSzPyYQjVcwYKh3L3
EkP1WDulyVLRH46ESy21unzb8yMfq8fo87jl6sqlM4v55V3qiAxIjZ57SHkCmT98pEPvn/Fv+EPq
iaWbY9HSwZvfcmUUL1WyhiCD/chc86P53zBeaS84XgYkfBr2+SuvNsB1HAG/s04/+65j/tMlnxTj
UCDbWa++91Hbs2g52TQZc7i0kiF4a6Xe+Nkg+OID6IkVGjEG3blzvC7wCcCECOJfwQ3vJn9LS9SM
w0mPEsTpAhubqUuvhC3bVNxXDhY0uv3pCE3qDNdiwtE/pZdvv9ciY+w86vp6+cz6JYXqY/m5VRYz
cgLONRZd2evAUukOs7a61wCcY/LPkOgebIp8k3ba+FZn6lY5LdA3+IPHUiaxFf0Cx1JaiJIvlVjB
4cLi60EIqSvQk47pAU2UX3lTCX5zbrXn36jeY8WQ3BX1Y+kcsFSCnX94J2g1/PJmD4DitZLldFjm
khqsoCmQlPoz6jW5BdzpMNtv++0iEhulQHVDt+EWFNN2cu1CyPiueDVu4M9X3SOmbmEZFL7vvAIJ
bVfruyVKYJ6jXUntNwgHhVxv2MU1q6DWNj4XlRSUL0I94fVxbKU9n47S20pyDyYOsfM503/aHrXz
RKoMjdb683JL0t9zaFE5IIvlDb7UQbWk1+oX8Uv7HlkCoc5JQakVZoX57y+ZrBHjiRkYJQMAxbdQ
gc1MSSQQIxsi453v+5zG3dwv5BZNZAnsj7PeN61+nkNTwYxX4r6ybMrrYaL8PLHGM3lquPniTVtx
LTHJzvl/maAh4j9yV88BgsVvtc/zgp+rdE3oPmmwpY12G3kr474tHHxhMNi6+xRZD09smGOn6/HI
SCL2DU0WAHZfjwd8pL+/at1BKvBgbSVOOHdfVCT4nYbw6TPkiYx/3Tr0q3xDJBIo3R5TeX0uTw+y
D+jyP6mU+pPUTkfDKCQiKHsQce0GAQ7d/B5KWm/A+IwhB/KbeXtfxsfZLf7Y4oQPAWEyYRUEmNi3
S7fkFUBAcPJ0BriopqOfVgIjbsHCNTDJ9BXl9TbDgPY9NPl0bAZzi0P1I9NvkRT28cct68O3tvfp
Sf+aVxtCdsHBM9EwxZpRkhoxjd5tNPOIpR0cSxV1FZjIfhTNYMzu5NQnLAmgZYx7zK6HraCG7yzH
ENqZ3lPBCSP8Q14aGAj7NlaIvb5WHJY6THFYH9uAyzGLBgrTYMAUxlnUUsTs5PO2CURDneqEAwpB
RGMiWxUbbm1RwpavcJeEwztLnXYJhr+yvJSuB7NY8kU3Qh5c4wteLukUsmBmJODbEpvd/jS3swoX
G5jJMvUBKcL3ul9urrYNvXBoscX0cYSv9+hd+Xq5rHhUrH2IKF49NAD+PviQfwfwUDQR/cEn24Ob
vyEM5pcuXJBsTsRGHH5rk02JjxnCJccvBo0FZA65ahghdkDwruCsN31voQnPREnzNpXdUbOXDkjT
irybnSFB1VWi8fCqAbjMj/nIlorY9bR/YDv6C6dNLF7H4YzjxHab0Z101UlPhiGXpMq8YTFnOUtn
PHBrLtCIMUziIHar0w37utewnqkL2A2QRmIvB+sU52xDFEwtnPiGEFVY74VMc0+fg5Ckmz72zCKt
NPfRB9WPq+FwOqVSApgvj0dG3EH4K+G1bg++4alYN69ISKpidkvk8NbtimrHs9FeKtU2aPeU0MAY
y73GQCTOxjYtSA2gnUNkpjpF1MwEPhK5i16xD8a5XVHSvouQqcSeRYWWGQH/EuATPC3p1Oa/sWWF
OjOntDiHGJdZXI/9IQ5qzoUKD27dNZFbv2/VnkzbunKQLneh91/WZeF5OuFfpIOTpfARwW9dKrIl
rrL9MtWS7jboCZEmibVpwkSmfFX1Ly5GqhwqhNgaahr4GAI0KwpulgDHWOnPrgYfbQMvlwG52RGE
emnwOA53O5oVNxLC+reiq3Yncs7jMwlgb4RWefh7sTVLutdAfTxlBTgbnXpGn3lYlL9074WoAS/s
XSUZMMddbBMFth3OFvoyA9WyjnsOJ+qZjODGklvImNfb9n2Dh8d9RShJFREupJVlKRP7kUFvQjXr
djmtNJN8e5Ff7VCnR2qiEd7LXRoNFx1KFi03TPcCGuyDiwtmPM4PMFlOgB5ypohttMsakc6vCW4e
SXC2E2X5PjrdPZFGoa7Ukl21GuCiuItujMQf7FWLSrHK9euu2/HgoKctPelRG/LH0G853WUDDiXO
IC6PSUo9RLNAYoWVbBmPKkfeRJGAgCRPLKu7h7uihI9IB5RqoyxMLWkTJXWv17coNC3OSt8C1Tpm
3jo3Oiy+TjvoCpxe45giDY3wP1W7jWZwS+x+XBfdfDMhCAR5PwZzyEVF7vdbvs/kWA+p8LhvgxFl
IrQ3bRLWshy8KcaLHfIwfdwWrjcvqaBWqZwajisZsu1osjk+BGK9OJWdEVawWmrSy6t8ptpkvznC
gRagp9M1+FTOoy7jxjQkZNlf4NwTgXP/98J0GdCmyjRjj+8vsdPWbqLOQKUNzJ+VBVJjjfl77rrL
i0FHc7QgzOiwoLTBnwqSWrd7S1OmPe/abKqswIWj1zJNo9TT2ECGVsl/Ejuo/PpnvEXqH6RusRZy
7Xu/YgVXFVzODTT3HO4qWgWUENePLfg0h0w3fvZpcZHKUnoYJZ3j7lvDoWqdhb+K+cAb/XGXKFw0
6FhwNIQCfdS6Oqm1WRfLzyD0y370HQBWJNA8nRY5HvRUPNNJ598foxD7Qa0ZcvZlYT/vCgEex8Yy
s22sA2YSKVCczn7FIeAdNAdG12A9NTR4undeRAh0bw4sRy20tzRMlNN/Ywpxla8Tml7vHJui0+Sb
onvWfgKjsSjHfYOIjCHdnRc4nFl1VFvuL+rnbER4fwaXNn1+biPJ/k4Lz5EebJhUwofTYdauR1YS
5PzfFwZo1VT35hxyzBpBb50enbeErq/a6h3WjcPXWvGLBIAwORWSKzwLcdRA1Bn4J+U8zYhbZXcR
YwItOcXfChZW92OkAa0oUmRJ96kpJR0wd8i4q3CxlZt80LnV/NaY7OP6Vplmi+K4zWHffCXypzJL
CJbx20ytOjcaItZibWVssaoBptyNQVgVGhSGDlSUySplrk7ioc20fSkC/IXuQAYOqHfSV7ZTgKCS
twW7gjsuTu3CXWGYom/u+Fvls7mXuYPkDCIrkU4r/Sscdkc7PLaOMFgp+YZVg2inmKxSqL0Kcnqv
Ns38jrW69KipPhB2/hP9crOCMiA7UGv+mVABrggWXE0fXrTidfQzGcfSrN6rwpKb8iKdcmQ8bjzg
W8xXxLNb28FGPq6pFfYcGIQbEJjHl9yOwhiaiwnzwsS4keQf7N3VTTJya7bWYsIVMlBUBsdlNjGw
gOw9U9IwqYNbFMzQ17DaJLrhuouDRtEVLWZlJ67t4WpB2JhlJPCDICXwDlNmVZ/qnAHJ8bPUbR++
5xIo2R1tFnfyPUHf0UTFy0ZCbXQ58p7Di6TYyrbRDyJ8MRNMMZh3HP6L4SxTUJceN5rQrkhEsTbA
7d4YkPUJL5kt2q86hxKDpPwaL4u/K4C1urqZy6qU5KP8hOkG0i53p/qoUQ9iJMIwR/CLo84Cy/5g
776+ntm2ONOidH9CrzFSEKm3ddG+MllPMfOHVd0s6eyRBSFTHi5/Y6wislPspXoFnFr0We0bzpvi
oe+4NhBioWo0ypc1sazupajF0bw1Rrl3lb8q7RAdNeMpuyXABqqasbkAo6lvIdySsGq65fI3UpL+
eSL2JZkkFbd0qBq8YOOfFiHYUXUyhYFBE1z6qsS16+tDSWbcyEpRuqAm+cQbnrpeFfvZws2Ej4jW
RcL4KXFwYsP/XeethM38oCivLoG/nOXgdtDR4bkqMMOYDUHmjoPZV3kUljUJ529zM5NuV/YjzYcw
gAZ91x+/xm7KzmOfKSRZyLYsPnOjpKKqcl1FwCmVLYuFDA4UiGrm+FUEizqpro32312hEkCTRsrf
DMxnVVrYsVrncSM1n2ry6KEc/xcZz7RI08s3JvEHOQik3AVpfSsmb/G3fCF3aV3g7rU/UXm6c3i1
z46M0VQjaE9mgt+VLGZzaYdiuaeHI4wuWt8LBIQxx3zr8K/Ai27SkfEORBRcsIA5rJwKTvmMXnev
kAzX3T/hmDPF5MOyMk3d0iSu0RxDtxydJUI8OoRp6psmdwDq/61CmBbBf4wva9T5n+KjTpBR5PO0
dBqTFS0pcFbsuliOp+FFoGIUmJHkXgV/mJFfYmwiK78zpEqH1IRnaIAsw9Eu/WJhGgnmrZUAO3P7
op8wjtviKBn3YoW0JBCSWI0BsxAztk7/9a2nDaUWY6GE37G2BaLx5S+7yE3mXIT7ddXFoouJm1l4
7iRhDnK/h1lDWoChHbBNoe17603E04eb3gLnZY8/urDYaDaM2Rr34vPMxrJj48KxmzNzagu0e+rU
BG2d7O0OhtCsXx4B82eIwLTkGeEUodgwbe7SKgr75bLBeLF7//e8EgkC0p1Hb1Ig+2nr5+cl0l5R
yBwNQcd+/KawzvoCU4bZM/WnTcixEa6mFxiIc9u8wb4viU6aCcd08M7SQT9LjFfIHtCkECbwh7RL
7LDhX3D20p8Vc02v2ANeEc+4nlnyDmbcNyvA88O2bYzkAMmw/bznJFtHYoHVQh+1A6XjF92Yj0CL
wfI7ejqvJe/OEwyr7zfuGWEP+rkTHieyN4iKnsftyiEu0UHgNehSxL0t13P+N/FtqgcscgXa/SIl
QJEviGGVWE2fkpz121ZhG/wglJJliBpIb02QQGByQ3gpohthFV9718Jim73pXIUvn1GlqtAKp0cs
MBvFQdtZsVIVlGAv0LO8y2PuVEJvDKH3l0xIsH+mmMsNe+DwwceWJs+5TMT7n2h8GE9SUvvi0Kri
8pEcnUMfLGG7CkIXnAHxKFk4n3VwplPTmt1flees9yAGyHDSd8Rxeca8bl0ggX0xfX7kHtWIOs9w
XREmqJ5GWcNxZxs52TV1OPTmJ7QHmaCAe1Wd5BSQ+hZNbeBepFzFkhLTNqqxGt2xz2t8XV0Orofn
wGUN/7PKAbozj6aTCSJ8gqM0+woDWxTTn5gaxVEmxkYNg/uqA/+sIpBtJL8rQOzB4qWOjauTrjX5
D75ZJhvgHF7louqQ5uciMNw0FKWpgBeNA0BTlBsQIVq1EWRYVDlXBNcGeKFusRjqeptdFGDY4tFc
pZEJPP1krKx/d9SDJ9ijtERiC0ospNnejxpJL8c+0I+jTQ/vb0WK9/zV5xtPvPLNakm3oxv1tTBD
bLr3wrag4K9bX4yubaEeL9T2g1SWCpseNQ1kZ5SPPbfa9UHQp7r2684OPrmww0iiNsmFCO7sH5GT
ydxk6mJeH7C5hptffGCLnkeA6lHAYe0LntLUGpmcJdYw/zfOZlWcWr6w6xVENTxZXkZd0ARmCJqA
SXxodRvFmh4kAi7QSSl5znqC91L2UPpMCmR2lNGdu0CvtqblRSeE3qA+al5u1IFTgQbVCXG6KjXG
NrYYq7jTNp4eHyUL0Gj5P6FwRN2l3QmDz7qi6mpQ25t6xph/QfaXCaDL7+GeWgUwve0TpHgzHj5/
QSpsivQiNcdbOOV4D5LALLUx/rRB+UWpQIBQ9um9mmOX7Y5VPNbxBICf2//7+NvDiH1vadvFfa7h
qa63hPqyqM28P5oa23XRshbDcWUV2um4eUWfUKINrL0lWrmZHEezPmruPU8OEe9ly/3ehx31P4mT
/GPLFe4rT0jUjKgHLZBHVJyYTgRgYPY8ntGjhW1qtzjTgTKcvSuMEaQXXEIzWmaAWGhIi+FDWW4P
IM4BNIKOjy3R/aKk9Tyy4o9wWt1slvluD99R2csYsTzBIV9s7LMjy/nNSEAS+kj9DJJnANAR4c2e
PLu32jrp3IICF4UrdfsagfiWkqUf+Bcu115ep46oXy5acIU4+r1HbclBrhbq4x25rYbD8Fd7N8Vm
f08LL1zajMHDraCMAZUZMqddnY5r+DR73hkEiKduDbMGqF1szB2DQaXdVSygMdBUvWCoTwVhDlpU
MRKqvYZiQYVrVqkmDWvquBV9zdf+8iiiqGorXZloJpCrjpBpcNOkq2Qwak11G97g29GjvB+GA91q
usx7fhvzFGMWZpLd0tTIhUtImZ6C/17lTwqAvUWCOTg2eXaCVrU00RH4hoPhppCQGSy+9Qdd/+z7
GGgD9Zk6FvZySUIdJlKWOq/uOT14DK2ZnLdZK2/W+g/u8I9hXPBMelH7avknU/HEoNDfyvatgLK3
jVgkAgg5//hrgRdujFjlhjnn7ejkaa+3ymHQtT8h4Vk+aT1pVR92Z8raV3kbRbEFkOjloN9aiGl9
UkXn1m3CSyFtoileZakhO+M9g80KHUk7YKS68pN7Wup/WRNCwHUsg0e7vVG2hQleg8QlYaXMdqxL
lknzRU+4Blyy2ajTPYDlqdNvsTmX/e8WLGA05WOhpIwkmqHrnzUddoDX1RhxkY2HRtsV7WQvn8JU
wdxbBB0DhCGLADj5D847ZniJXG+yc/Uy8VFNWFjJNq0y4gGfGg108OkxSlyj6e50QkfWT6qPWr3b
8Sh8Yofa0ryNl//MazHSWSU6MlbNxiYxZQkUCSF/W45Y0VBVqf+X5j4ZgjF4dwaAazj6Seq0kI8w
4A46SDRyl6A9tzHXd8WQ29NHc3/6e1WfswfiORLvAin3dLDdOhK5MbUwMa/6IJXv3C13MZcyy6ZQ
DIkbkTK0OpNEs1vgYwpw+U4tc9fD53RYWRMj6xXPGcR/SwwIksTxDYNZCxyBkaCs6dLS51ByiOd9
2fppWPUUCGVcPL79vxOZWeDkwPrJ6A07JA46ErFd1wIie6J3GqWRqlVImarxWAe+D5Ny9gHFcHe4
7mW5fjkYRy7qMkCN94IsYRuwumAWPZXlU6D5p3zVuuJiudfQLwjh61PrwXO7JBxtw5vLSC4MsC3b
NkrULkzu9S5sRamKXWi2Tiu9MMDAwJEg/Qjm5zpXiz3KgjCcD2jB2CMHIoDSr96Nqc/81P114bKE
mKLyFrvp/mFawTBXNAmQiqWiN7z3W0f0SDL0z3hm/sAGIfCZPnsOJaVKjzF+6NHnLNb8+QZa7/XW
4dlIOeIV+E5PiWpvwPpGqUGqKMbTKAxkzB+A4xtVV5lv76vIqy0ev52v9eMGLc/Q2xu7VKEf20MR
dAG5m0eZ8gPhWBJ97B7ii1+XuF3ixMhqhWK84zclVNCTWHuRuAQ95gYl8UQvqu0bL/dd6YCK9Uzj
B8SuMSo9KST/XDZjk8K4e1N2SYKXbDRlsR1Qcv/E7GLCClXxx0yagSnRpydi7iuShXEtAAvnJYg6
/K/5Nzmq2GEoHSK12e215VJbXIUwbpPfCuNDIMYgTxZ85cdJOCb6Yz9cuf9Myj9MrWjqnozvMD42
XEhr78AIQN06t7e68b1WNbcAdsEpn9XGZTTEw9/NHzwrNE6f5MlViZliCBs9q1ohTQdAJm44FcJH
wNnRWOOLabuZZPKtR/Xe/Ka+0liwQfBOQDj/L5XO8rus7/KBG/Rlj+xdraZiIiGPg9AA9M9NWiER
hZKFmMzuFXk6VsdcS/cDdatBvnsPOA5VRZ1f2oTZWfUOPhxE6OnkRXl2eGRuIi8HnvTg9Q9ZCGH2
UIDi80ndbkD7zomJkntu9oU3wi5GHeQql8eHrDArIUymWSeKSLa0hLOsFc7s8oTJhm85vy26BYwl
8PVTgO2dATiGoB7sl6zeuMTlmiVplp1zGngbxh+QbCXXKNg4J1BUUOJkZPRqQIj2iftMBn+GY8ZO
pnZNlA30bW8WbcyQQRKjpUvxjottBIXvYcGweezTUqA8chW+RTSc/7h9i4IiohIfkWJmpMXiqObr
j6g/9pVYxbvtMpbkp+dPXWCB3iWQBymKraM5FT9EsKg6+//7vqZD4vWtzHIzMrphwQ7yFCpYuZbv
iBfeQsRoSMbbdzz8cS9eZ995Hh5h2guT5fFtJfF06iQOExPPY+h/t6mYQUZJ6TxjFdRwKcLkDtyX
gmys+Ufv7OJmJrVPB1d2uLuxoVO+DQYtgNs0KTFJIO/diE9oMut6HChDWlq789ZS8rS8lHzU+OXg
0m3E1JfJkQlbqXBLsrMn68XuCsvp3AFyaro8ARUi/82Apr2l2cot2yL5vGwqggizYFrYR6q6IogS
Hdn8tK1qzbEw37uU/yUVvzH+2zBXbJKGPhF1FkfKQqXpj0IDrTpBb0hS5tQhSF7seTWt5NIiRhqK
ZtXxPq4kSiXJaYOFiSg3H22EK70sDP4xUGc4TC8W2/bUiYeW0qb94z7LMjHJMRp+BjE+k4adwm8T
UdxOliRBx49t1lLmFIyciwIEhf8EeZiUx/kd05g20Tw3ta3AswAvfbxCxpc/9Drb8S+39su99yq4
azNYmWcqRwc+KTTenfI51leLikGWffGg4lafw78I4Pq6nvN+JpOGy8RFgFM6kEK/6PlXsk/uE+Tx
yH3Z10Zh7Fj3PQD7GUeH8MDknxMlMjqgGKiiRFqkeyCY+9znHwlI/D/b+awMsa6mIlUdQSW1sU4o
PYeWnloddFyuIdeaP94AKPxQ93REEkU+ShUGQl7YLgciZC2Eklwgk277SJbfZKqAFgrH9FP67l35
H1nlsEctEP+7IZj6bT3DYGKm5Gh1DTS7euG55QgvkjImqzrZ/Hx2AcL2Dm3capluYsmVHh8g7A5s
iGUDrZWz0V2OiAhmPonUllk7wBiNLG1iQHGTVy6qiPs1XlFtZ9JHvUieN0lSuI8SLGZoBI5eKNEt
H+/1gr2Ryo/66lkmwJWdKWYSIj4dc+aA5WU2qAIA9ztm2DAmodwjsq7z8KoGW/t1ut0R0tcrdfq1
BNiAXi5Xmq087z3hexPHyBNbo7BTnaWGK2kaKFCrgGgXuoCa3yMwISm0g459mzxfeNcDWW4CnPFl
cOq7mschhgM3owrsBmT8y8iZ/ma6252v62QerXAJW8g7SsoCJq7psC0SINsMOGj8wXSrQSSdxBmF
41/D48hw+VViTA9qDLfe0cwWn0snPGtj7QOu/NVvOua7iP3V6XrUl/8Ix1T9KslnL3WIl8g3d+VQ
sATbzgM2J/QCul1shgQIADPdanoOMIUfNd6nk7lO20KoEIzqcBM4ySYQvDcV4hVNuEAa7pElBzjz
+RqI66/B9isrkiOr/EYS6Lt5KrgYq1Mt6eg1vwcD+vPgsppibIoUpHQBP4p9moEFSI4Y+JbsiPta
zKbqhn8e0v1Sk0ylIFpunZYcxenHvC3ZsLx2MlqRDdHxODKdQqu37qGISN/i+4Q1g2v2PJLrbQ5d
AXg/GGZWsokTBFnQwRuQaLZAK/nXtXDAFbOPMMrf8p/5r0pe6UJ3jlu06gXCEYkn4auS0I8aja9i
qnyua9DskQRv8+2BnaFnN2l5kDzmO6XXY4WWQF+oXeWY5xCwpkmypFWAa94P8aNUVQ6Jt1pg3+4s
Yo/hXLiQ0Rv/t0LR7cLCEXEBKY2QploFUuhSULgz5Dno7P2OcYIXL3G5e9eyXMtnkjsW6OnWSRfy
jy2Y6/ipAZQcP9wbCmyLD40Cm7y6/7Pud6jC7ldKZ8slV/Lt9uDW9/JnNpZxx8rpxIlRfuhWJRG2
SlF+IuAAiCCc88v4ZskkMmXVtAtEjQhmZ5MIyPsJrcE6Hzx1e5u+blb7eHi/v55phxvHkF0n11zA
kc/j7GxQm9OwW1MckT0oq/XbI3wiWzwhiTttkCpKH/DaKt8qZlZnWuC5E6l4nQNQOApxo6ABXAav
NaHIoopVc98GKhHovTTnCdKOjY3yWVLuDhI2IMpEx6YkUHdQVqBblZfqlIPd6ZCppgpcbgv9Q+tK
2BcXS02L6SZHnn/NoJM5ZdI4T+7NQQzsROTFwO6NV3AXpOO44G/Y6/2cHSSakCAI0I9+8vaH3bi0
Y2moVeuol9aelxMnHQ1MDFf+2I8MC6Q3q1G5rr5ptLoQlxqaRy9vZRn+29uqm46O1arKeN3HNyXU
dgAebytRcm2m9jnxIhyReC/IDJ+ZlB1rq8ZDWKrXrSLXEY+M+SewkJfVCXAD+tWAIb6OP+XZwKE4
gFMQiuutb04IdJJSTdnYsvQqna4NzT6LnSXmluE0AHNU+Db0oMQXNJMnalDy8LZUHjCzb+V+10+H
d/C0kGHbCrWrLxo9ROlWbyWo9qbIRhX3U0+7q+5l/QyahW33h21j2HGarGHS/g5wwQY7kCJ/nc5U
mrtpq8KE9R7cxeSPaJBfEskrclwsSZDzuRgCJh6uFtKv94xvmob0Mg7YjY1xpZ8NBnh60sKbcswx
kXy91ZiaPPDdMdUjJ3Uh3IfvIYYnkVay4Y93NbFw3Yfg/TFcqa85Ki/xZ97BTG0KhbrpytiXBEwe
f51sU1/uPFuVPMDGTv2Pbr20UCUxcSkFotx8Fj8ku5Jh/GGTJKkf9YhEOFTqGiTDvMD4ZX4zLLYH
tnTkA3nTOSo+fhfFiHlfQbpzTK5dlolv65Yo/46bihYbUsSfy8g/0V21WZE62ADjrt0n2xxKjm4X
xB9trlQTG5W3IVWEAMB8KhlU3PERmirabTucAVpVX5byqKul5xuinTmOI3/PSCNaDhUvLZ6rqBU8
4JpCE2eT0xSAT1XLvdY/EbNJbEHcCnfHIUbJSUe9riix6Dho8lKV2ZseRj2tjbp4NzAwtDPKvbza
MVvTOIVcAmhKzD02yjmq3ZHFMgVkQnexzik2tt3tYsYh8Zb+muDr81ERlNOqMK4WPqvxH1mbmryV
ullsYaeJsTonNc8n9k0ZosVsRXkP2O+KKK/+tNCZlGymIfdl3uIo4LX1MJzqJVRbHAThBJE3Z3dh
wu1+SJLEuhvDH3ayaPagHH/Lf9inKtL2B+sGLJpYZ7W5jo6xvQX0gbXmYJVtSv0aHvBLGm5rdgtW
/HVSYm3EAK0VKd6RhmUcAgBrHd3U/EdLawUmtsc8c/lSDPZXLiTwcZncido//vDEM2ulacnZEGMB
OxoMIgG75wWUQEH9fLrxWWdUiFOEL5e5LuXEyd9GYb/HwBFs6NaqUUMBG/41GKVvi8cLmTJmBTw8
PDbVfo7wy6B+o81PbZgMEx3w7ZsGuXgB3Evohm7s0ikRGuIOz3wXCkJtk6L2g6ostXN6OIOuftFj
7m5M2q0WMFbi1Lxn0BP7J44IPY5I2N4gwP/UQOBe623ZXC7Yl13S4FaLYiTMWfbRpVUhjfTtZ31l
OCvmWNswH+G9JuUKpljPQ2/mAX+/HFhm2dOke+9HecpbXWL0cX6QgWxXnSpMxEnJlW+YZHFWHqBj
JXIcH8t9EHXRCIfah6Xm+CWS4vQr8B++i2WnQaw7wQpw2RJmpm5cXR/WSvtgfBbFdRBHxAtc6KPP
Bv1iFjXnXtw0DA7LigbxZ45Gg/b8uEj4BDePJwLAV00YuYKPdatJs6RK3crZbUIFtVz6bKFfcCtF
HI3vh/NAqkEDbnroN93PTKZE68ltm0DWTs8yx3ZinO4ZdIDtO0mRwFv5l6T1Z3T1t4OYB2it++61
xzxDQYBEwg62buNBV1XWRDyBk3ssLzLiNGQADG+0fHpLMBradRTGIQ0mcOSdYryXOS76GIvlV6E9
aDXO0hGWlTFLwmrXgvTmhOmvbWKOxmjZTKh5kJ4VFZMCa0tUxrESbwWsG7gHT6mxQc9ZvYGpZrr5
npROyRo9G1OgAcFvJn++J4WpszYm4RR1JpmVbVWLq0JDIKfAMXw56jn6NZJibdwxunrfoFI2KEn5
3EM8M4EY49zPoJ3i2whLFmSUpx9KkGNLpVulZAZ4A8fsM5Fjmv4oaOZqmY9dq7XJd7w/QqEGNoKW
7RcqL67snO/K84yWSHWIbGpjSOVozAJ2D+wcanjKYzM5b9umePGUjyUj/iU//LyO9cxfmufq8oc0
ko/k2lUd/KIACiY/nkS0ltHLDARpVT922AmrliUduHaoHUyUDRY/4nYGkJcy+AQv4VvTXACRP3rd
Q0N27utXNdWkDXKfekkNsR+2ks95Bj9bUNNDSg3J9jGfrKNwHmpvvOtZDDI3u5A46T8otzA0qay+
jgDtIaSvpy4KJ/wWMxIcUakoNmZYEnbXDT6oUFSKW7R/hhVv3HRDEr8AZgLzc14g6GfEQEaE1xPW
+afnKGjAjF8rlYkxxYmTqXZ0RPy0kGmspvKMpEuJkL1dzl/SxvpHu+Y1SPucetAL23zXdQ14NZKS
Ik5nESGtx6xG92C2L8OqccQa0okqZcAnmeVron0EE6GQ09BxSKoUeb6uRF6JfsDRCpsHPxeS15D8
EdT1n8TevQ0CMosZdHtSCUp3owySlEdVQjVK8N9hrmfrV2LvSXOikceWUI2RXZI4pQZU6wPqWRFZ
Wn3fe+bpzRQdQsIjvUVdLYE0f+A3qzVSEXeONLFZ4//vr/E7PnTPmaWbqGCCiXbfHsHW87Sc0bdw
i+7Qgyspb+pw4qJgAcw3G8Ann7MKeFKRILSYH/b8/ECPmZ89KHM4cRsl8KQ4OZX0l0iwnbf4ixca
4ma9C1kDtUp3jblyMf+FhHV5NAY7gtl3jLRGOsQhwaGekqqjS+yIjg5QbnZbTW5bEb9zRrHqzy+z
Hth4ENo+x5nK4vZaibvtNBzKU0eb1rKxFV6K39sPM48a5RL0iTsWItgCRxdpHZQLTIIBv4tTetZf
v1KjAM53/Rt0YY+XJ1LLYeLEW5JOH8mUaj7VbK4pLO/Yqwo9crB/71+tgEYKloi9AYBbtuvPS7qd
9ozGB7Q8nalm7ffMW6GCIG8Dvmtziak6EA9JldhpbOCksnkycDVaPgvRxPIE9N6eFPM5exc0AtF0
DpyHiS3sOCEGB6jM1d1FPh5FBA39N62V1L92mvm6SdU7pigCZGhiTTk7njdKX9MCCnjsVOb/pcbz
tcTTLIvsjQ37V92CZG8Uu+9OhZ3/6rw8r9sxbh5SM08ia53Hn4CODXVJjGaWbJsO3htF/TN24Qe2
Zkao4imuIlpHM91Fu+v6YtyC/TwA2MFhrUlKMHvywa+T6yEhOeWjmiLUVWYC36apTCFmayLsF7R7
DGQzmNwHJLLDn/ScNIr7phBtQdolbMMUn31T9gcKnS4ZyMTW/B3PNOaSxleGxqmFlJmowirJS2f0
c5tTygGrutKv2ca+j44m7JRsb/2MqybWk+nMI6OIZnrnJxnM25LQyzDBC+1w2IbRCo8M1FLDQp3t
gcs1wzP5Z2U4ZmZMIRdPu8MHMh1kEoT3yqYdz86gR52BK/RCCF7jipHAo4epmLJGU5sBD51tkjnr
CVcxISkfaCKcQG5Tq2TaZ6phSbotXket7RwkvtG98e0ST1Eh090YpOq6/YFZudXk/Mi8Cw5DfQJQ
pvWhfluLcT/EHIoqBUT/Bflp7FC+jAeKqhe6LO0XReuoQS2fTN4Bvo5+K5PBHPB8GR5LAd+DEEN2
V/bicLxJ1MfESHNF6HLXJ//47RVCY9jUUEAmOGxUJVUXBOlmp6U1lnq5OgKmHefaC4/9WPJlWZ2v
jzaSOqu7msGFmglQapEhjIyNJxbRFBDY3P8L79XB8AtKsKvdsQwTsdJ5yadq3uWib6WeT5e3ZzDG
DYNg9NuqqnaRaQ2OyzbuQeQiSh2H05KdO2DavJcXoWAg+Ejid+r16IW0Gj6Cw5pxXJ1nz3eENESE
kNscVFqVKcjbORCFDMi8PZE4rOpuHTpNV649YLR2MpaTi4Anb08N41AzYfv/000nic318VAsavB1
ON70i009QYOVHc/qQW6YYiPRbodpx6bgpUXUbzpNPifDHkTeDXPtkkCEQmDOplI+dh+U5DGg8oBu
0f0ADFGZ1bAqWBPB0hXbrk9NW7IUJ+85PaE2cAGYr57BlR+CB+XPx1bTbEaie4tt8VJ+hBc4iSHa
jOIfuVYoSiaTf12Bgskl2w7ydIPh5qQl4C2GpSA1jzAKkvGnWHTin9O4J9oQygQg+JsBr1uY4yP9
UdquLziwSvWtgI4mt5PtsHCJ4mQRZZAmyqZBe5TjLfjMHN2z6XNTQZTIJujWpG+JvzqP73oeWOBB
bww+WJJ7NZBH2H8ezDjQBGqusZZIYh7bCrB68D7TYyAmOSLYCQxE/8FWh1mzn6s11UXQzQSewPL5
memr9AxuU7rw+465ZBsQi1Tw4n5iQRIyU4gU6kn8j6apMVtTpAyxMLQI+f2w0wsA7sbCgB8wjTN+
2f2C+NZpiiU0sYX+l2yaN73eedcoQFHcfakRGRnY4VYBa/8tNItwlQKj6zyTDLRzkKTPcgllmFyt
V/lQtrVlb9rWm4ui3uqvdwc5GZ21aqyGtwEaToLbtaWEAgDbfM7LFu71YisV/rjhmwtO6gc39QIB
t0zYNH4KejfrAkpb4Crbzlr6V3d9mCTIKtnY1zSH7L3E3179NhLYBlEdHxjDNNxSJLXARNREEk3a
TmBEQTRQ0mPuIDNB4nIYq4qjR+/6S67lyVhhT38YMLG1cez27nTcn8Qp9KhhYF1OoTkbdHWyyvSF
G7HMrg4go+i8S3IHp+5fHDcw3RhtmfCGuBF3htEF2PkRlmD3qp2YMQSLdJ3aviY69GS8K8NGVhl+
IK2vFo+G2niflVMb1QKiUFdfzrx0DGsZkKrsGAbY2jzpEkEn2XG8JtwFfi4BveeWhMMp5uMFk4CY
fsk/y1TldnC7QGRWxiLV2eOtxAibRidUEDPLLRhCaeuLQH0tli9M/2KGiQ4/HqLxFg85KtNjwLnF
N7b7Bg4/oziEavYFtWzR2MeOWY8IUPkbDHbVRO2eipg0j1gm41X0VMLxTrXglig0QGUchy7QjK8x
tPyNeFnwGQ0OdVevR4eNz4xeeoumpF1OBWTG3Iu3hKqEc+hsmpQ1PJLI4dqRcYgkUrXN/sbH+2sH
sMKZSX0lfELM72ZdvDvgnhcU8XJ1ZFjEIYFs8pYYUatW5gPNUP1Fhke0d2owZJJZk0Vs5+9JIOLK
PxhKQrH9NLqvrQ/dRndjhKzEyOnacpgL3R7qvmpEEtVsKhG8rp/oTgzgiA5CRJGefbuyxx4RqeAL
wwLHezo4k0Ohu/DfOh532oBidS6hIuHe7aQK3Q6odyNtNJd/2QnIiUCpCcLrSklL2STstdW4yIa2
uJj9wiUiAIP+6oNYiT+w1cOJr7niMMN+5/7on75AR2s01YRkRhBV3IBTI1gsMw2XrqeojZnxz3XD
6LOG6KxGo8l6NZGK6QR4qbJxABzOpYJjbYNvATnjp2XPfQdO/UiVOP8sWBqVaLeP2grrpVdE77t5
T7Pue1rlnEnI8bW+yQcasNM3HFKzMjU466vBdOP8Lzjm1s1naVf25UirEaiTv5UKbL+W8joiYHB/
QGGSotQVKKtU6NeAFOpFPD92jv+PONEHoU3fxM3sC1bQvPNoaX1sZPLdQdZXARYv71YxzW6/Jk03
WhA4O9op/wAw2XQa84Po00CSTaxsLk6d6P1w3iegntaOit/eLi85C4V7LmX9yf+74kwM3B96xZTP
G/z9L2szF09RBp3YDyLwK4hF2qSjXgL6NVLu7GrTFv1ugOMLKBEaceM31UwTt2D+FZ3KitQdshLC
WCepVcnS1LYw4qw5IB95V1P+3udc0WNU5RfIib9S2/i3Z8G5rC+uYOJ9DjphWk1zH1W7N3cN6WgV
oCL2/SjWXTNVQHlkSWTn6DNMpDPGK1L+qL0Rb1BUHgshT/6+dDGft10JJPLL5tHKjBlIXGTahXbN
cfbiCr5zx5zAAM6T4AEPDcnuebW5Z82ADDT2KxBN+qabn0kfpwT8pEDoxDRiAP9WWy4AtIoSgA/2
sTg1FvT62D/gWdmXNdeWXY/173y+7EpogEQCfBdaXPXeMzFnqtG/UNmIqOCAMiVIuhCcf5Suk38w
AD/9PnZn5KYrPR4naB1OGmZaT1WOpya4JAkhRzXinEIj1Gtken7N4vDxJ6w3705o6u6anWRF4cZw
SpFGaFSgugqtJ/QuBLvty2f2CtZb4TZohWzEauwdYtUU0tvF0Yg73A0HzR7wY/lWRFZ0n08pNCo6
5gYlPSpbqeAv+VAU2NNOsnqmqE45D5X3gN8yVElpQJd2I0l6SxFQW3nS+xf238s80oqo+Go9EOXm
mAqZGCl1Le2iLcl2RPwe7A+apMDUiYksTzj6u8cq1MquP63AcU4egLQ9PXIQsHEiUH8e1xQyJONg
Augdbr14ULezn7XCSAYAcxtnAJlLhDnIjnEwXTHal4pPG6z55jPtBxH5qLtAEJOu0Qdg3WqLCW+s
DquxHa4ODN8iNo7/SIw9JNvYTPyemHnRe0TibIiqLYm5GMu2tu9x02FDLiStj+dgaZpwDLWShuLv
X73blc+vSqrb08mCsfZVhxy/u6A9mt58iJ6WkG/4P5ulJFfiJCD1tgHdUMuH8smkAodP1jYjcdtQ
n56wHioTFSPDGixsiYZWQD1wQYBS8gzNihXY5pZyiYnlD3+M3+SJAguQV7fjy6zhzjAFBUYTcFaD
E/kRLlh250HzhnlxB3sMOcBkBZ0e9XLfMy50DshRaBJDsUOXrlS5NfTYT1VSC9jV+tho3lG1ylek
SeKt2lZqWEaYHqcmGsm+rABbpFYMqfScHpQtPoKkFvP1SmQTZNYOhxZb/loA4qnHr4jgPw33c4US
qrAEsTsClV39/t7AFO802T55pt+914q2EWs5T/efhgI8mM3orIRjAolWaSKM5qRRL++wSHYj2xnc
UZnIF+nu4+JLxjj6XMEHCR5PuhUjFp/B7/rOlBVKeUqAZ6pM3kAy58ebMaf/0VbZS7KEDvaCVPKE
GAC39JtVoEO2m9n3u1mHHqSRZG2OzvYytu+o4ezVF65xa+Oi8F4PuZuC4kGcm6k19NrRA/bszuuQ
PG5yop+C4aCXKHtrtwRj2g3ZE3MxFwRBcoH7wc6YBWtWhXIfCbfwfWSmDSc/gFIUBsfr67Z8idOw
FoU+wRb/GOWfzWVQTumWQhvDLyf6BumLMnt3TiWezLvqh1uzv1h474KASnK1n3OwRMh4kHeHGz2s
kQiM8HT3Hy31A7NQ6U3MUo90ZB4n3abJpRVGfugkMEda0ZczE6sjepbLODirVJkgyJ+9hVE8HbBI
PSrL7f9oHkdmM0zq6QQg7HCj96fpe+R4WcbZou2pXq82JkkEzCaGp9oCvS3kxpbfyEiR2xoFlqZW
wfGcpDwc3a/zLQAtD1G/bje/lUp7zAylVDeXW4LQCduWQXs5YlSepnURapPbYIhHIj0cCtBvDSqQ
01jBuEvnYM6YoTpd9klAfCf+TeDs6bq5LRByvJh14be/odMEH8ClRC14OAOpUYaFW1rP2L2kMU3G
wmifrTfyels4r1McpM3OBUa/Jtq7WJeEDZxOAwrGQe1BcpedcDPT2trFmfwcLzJRz3QKTfO1+ncw
/YPPPaxGKtey1v/MiMoJB8fo0QPsSQ02kT4XR5pwE0NX0LqrSQMi5aDRKTPBR6/9JB6DdbnYl6qe
WIoWmNN7AT9z5T/SmdSqLwZ9cWQMyCQFJB9QMnUY5Eoiu5W9gDiwvurJQI9OGHa0tGEueet9JvPJ
bRIw6jyKfX2ixDrsxtNvEztwxlcBU/zqtvMM6RIxI6gL1J1KwIRFvUSH+L1rKKQ3I3bb1HT91UbM
bEkHCGyU7DoxpgSKtnFbvObHWmYBUHIdiiJqXt6Z0ToD1OB1xbdH+6psV1C+JicDSqver/WHP/lF
y/gZv1I8bgMT9bI4tb7l6SfqkHWDNUS90JLzFqfJ3gwwgjz8TJ3Tof28AqGpJbP/XkRvLYDN5/Q5
EQ93Hjjp1yihkE7SWe7wJEKmfsGOIexcgf4fsNz3lnqemRLRaohJY4aIG2PDbWPryfAlaWNjzOpA
4x/eBWqJ96H978WUdagzuX+A+gdWz/y12D3jTKOr7wlfHya8kftqrYNUfu5eboTFCHBIyQzSeHg2
A2LQd91obwEKYl7m217ZYaE9TWQJLEy0I3TsrlmocIEjYswT1gnG/oaYQKExAZ+UE3MR+S0u/bsU
1qPf4WtJMbfwxlHXnWie7Mx8C1IHfaXsVPyXnMdGlZoe6WpJNPPIh59tY7RolgXHHa0MWsS3JxeO
QJi7JH+9XTzdqSnspmMiVwQyYr80OVShJoYUTboGMigV9oU1bKBQF3TGh6WvdW95K3XCHCl71Nds
J49SYsJKw6Y2gFBTPX88IGSLcXwAgys/wK+HAiofIazQKBu/oqLgxQ0wXPr3aEKRfRMoA7HniQ5N
XZyU6OAxA4lAV5CKSlxoS9996ud38vlSSZVWbMC4hnQH5WHAWDq+FStw9Bu3X6u99klmnGfEHWJm
tfEOcd29scJw5bF7az8+I2lEttD6WtvD14xd1BFJzIjuKwCPSVt+EhRBH4DHRinukQ+SZCoRBWq/
txK/e84di6q0FJcKjD/ATFuMjvTn+o7kW3LTZh/hffKOge09AcF68Sto1VfONqWkc7PulwtymYV/
S48/rBgDkVfxEfkqrEwu3T0seivfgK4sWGfHQ2GulNX+9RHoLdUK6XNKpQZtp5C5XhiuzC/E95ok
FvFcUJxYWvYaMaMrHYrQ+hMBmY6P+PMSJos+gmuXYDHdCwYHK0pCBqqV69rAsu66ULXiS5LJ3MME
q0E1+lOevig3GcXuDVfxgRxwA7wUJ56MUnfnW0KVGUQnjzrlddReFjL0zavjJ1vwLKN5T7AUhRHO
JQFO9NsijvDil4PIyEeuo6OuEbnvLWMiP5+R/VhvxiC4ykeeZnBYYGszbv/hRSKu7MCZhJIF61UQ
v9KnFr6/cAcpd82NUwPu5x3KmVPIq8jpQypYiGyfWi2QzMTx0ganPOkifkcQhZ/HANq7CYyVeF+g
I2xSZptjl8Xv4+9WCXg0DX8Uso9mWbxzr6huSMhISPjO7EFUmCSRHXgUSQAxgSeOb0ZV9HLoGtj8
ZRnMDuvzALyeAI9+kv+TVe4uy5hxFhI6uzS+jDURuoWmSOwnwqL9x/2lYs3Czrwaf31/8X78Kfiw
kb/yXVebg4h865dh8Jhq2DQgedo6mPjsK8CoJQHf/x88AYxBgg0pxYxp+J5+JM2/qjY0qmlGeuT6
k9yJ2b+L2YoncOUvBH+PGJ43wA6vF2/cN+GIOxFH6KQYSvF9/W1iOdeAElbgdGU3p/3LazRk9dD6
AjMB/lgQvH8GGOj2bq9uHS4ZrQ/6fkgnghtshsUlSYMtzHLNv19/JgZ4XSvn/VGqokvHOYQh+tZP
ZgPoG4t3Rgz3i5SKmo5wCnZmm20WdSrhBXWYvsKhYMx4Zkw9p+cf3cKn995BTys0KIC8c8r78U43
2MDfWB77CHJL7zc5ZzWWxQr2kh0twxB2U57h05Qo2N96eDPfd/5JnrFwqkzenUP6ZAv8CMf06f9S
8eNgB2zID0an0erXgPBhUrrR8w3/MD5bgjHYmjCtrMrgalxXOEwIbg7RYhasQUdLn1ZCoxRH8TUj
Sd8SDvdoB2Hd1mzTPt6/hcZvlcSuaQ6mcEjGTXB5YLmb+kz7rGRyzCu3YtAIzDPh1ZRl3gEWVmqx
7KK2hRJiQvJ8/sop4Rkt7pYV+qD27GkoiUAQGXs3NtMPlkPwvCt9WUZBL1G9kQG3EcSMMcYcc8if
lEArhMCNjacvSry5fJo0/siyylCxr6+9WPl0aUf4zZlfwpYE2nNkAaSBZSdvkL+qw6q8UZ4MCbL1
/ZjU+EgyN63eEgu9AoDJEroH+1+WgxI1xDhskwr7+BoO0OHAGVPJ6DBSLk7xBNtwwfGJk/8nwJKa
2j3yrqsXe1KVK7VeciS/x91VbFrubZKXwzANnaNofZ3SDsSTKJt5vNDOJTPomIhA5cZHd1iMfxLD
bRj4z5jyZy7pVzf4QZTt5x0Bt61c3kLRzSI5I/JqL4UzAbPm7whUyMxF9j7ZzbCZSetHkUd8pB/A
fheFHMQTVtJXboATsBnYysWupw4qsOQCIE8M/ZJ8F+paozPv1+NC0UMFdpMwNwmtbBGDyfe+LsFW
zYD5q1G5901e2UVSzQ6M7FheIH2KFS/QLI4eSHgCJVbkvquJb04OBgy/zBfaYQ6R6+BktmTJpMxi
ohuTclFg3re2I7GSqbKu/7LIGxJW14odENaRqIBL9qnHlX3ebwsiNtMEV8LeaGH+3xtD3WIDu9HN
50Ea//H6ZtU6SJVH+QnBD/IZiS4JWbyHFB4nGK/77m7OzdD5EOIcS5mJjv5Ja2GwQ0eRKIXFzeMZ
kcF5+5xbtMvxzvO2e7ONPPrH/r0qQNgGb/OkKaEQeQfOmuCo/560QtCNv++2Tds8CdpgumAUMXUM
4ciip6gqeF6c7HtLeWgUhe8ZvuJXkvLGCAYUbWEMXhn6TY/VjP4mIP5bwWsK7XRVLz8Zxl/+269N
PvcjBFBlD6opviTyCIc5ycKELn1PAiZBvw+SkX2VRkIl48RRyACze3DSTpWMe5ZxtY2HU2mm5onV
xDwwZ7rm8Y369sof5EjGflKJwXJ+38pxZnevA5YNm8boZAdpOY+7eJxXOpg1ehAvB6lL4qsEtgsJ
jnIz6T5bg1WZuipEAYxsjBtVQm8Ie4Yz8IWhAEbQ0LonKIYZMnA19W2p9SQMwSvD0dc+9/tuHoKR
mVeh8bn4Xr3rG6KYh9rAxJ0q2zS1m2J5DCmkUdAk0K8oguG13B+SyRUfbQH005O/XgNXacppfH6Z
LbLmX2A6r6hmn4V5AVJbRPG7f7UaVqvJxmMPrsmS4UYBRCusoSSr+fRP8/WgmBl4+qGu5HqA6/ID
xWuTJVpEm8+SCfatEkkSwtg+liWMzyMgWW7aMt9k9D2QcoeizW7meNoP8sDOtzHjUWCeDnbVmKV9
7dKuLRnzF0GgoemqknWD+RIXeoeqlgyeen/jm1s/+PWzsuRvk8tVOT+Ge/9i0qmZVoms8GOfuq97
f+m3DERS0xQ/jrc0tqSUrVKTkX6Sw1j9+M2hE+0yOPkcvi2WJzhloH/B3vrr5VE1FqaY5NnJ4JVb
/voqQ+uMFSklNAcbPGixbFJT6JE8oPVRZKPUDwoOPnnC3e6Ul8+HioRd+zPSHtw3vcftdbcxJif2
iUQlIykjcegMxuw1AB5AaH0aBRxQbRjYjf+L9tT9s9ER3/JcF8nh6XHkaIMsKokIQskp6yFAAyqE
I0YbLOShIP6lmTbpIx6jkIqkYpSGqSsU03apBtxFn5HigUqgjDSFWsnbkoyr+abcN4QcjylEcfMg
qIK8m6b8mWsjrgRxYB5sHBxSqbdzf4oh0Jl58Ok4xgqlqISi4Newv1O10VhJzWfC1wgZINBmX4/F
MpOkd8XLMUVRLXmoYNZpO4oJMQrx0ezVWh60BtVsmlXGks1QEO9aS/7A6jEB8zj3jjwlT2wGQTQi
BPKezTUJNrSTZXZbSA7pdzVraxcBu0AX6UaVgGmkMxBRS2/7wbbbIVHA1QEBIq5ByxMVw8Z67w96
b0fUHGaB7w+NDiwK4fmmFydfljU5LZlbhLqotxNhC+Nfpnm6ZgXwoJz8+7DHZF1DTkDGtqUBJ5LJ
n06kdCFdfXX8nXeFTbP9yqt8fBPmBwwvop3OuSnxF/0nTOkBlREQh84oqqSjvgV9kzbImYZmmlj7
xSmHOzJ0XFzfUtWjPnbVkG2jJj8F5kK2nOvjYkCoRAa4jxvasObibq7NbtDmODvU/acOtHNnTPWV
4fpCg5OCjf1w67gkQPzJBZXfD9x4hjEmX5kiKBhnLSduGvwTQYy+mg1pyDi5HbT5dG7vYZ/PIHRt
cvkw3IxUL+F5LsB5/thPP1/WecYOYWmhFP5rSc3dAhdkmzYryfPjse1c44cpdr20o9YRE+gqD+5W
Gnym4A6PRZGUaerxV3LDDgyx5xrXyvL7XforBtiTZ1WmyvQPquSRq56/Lu6P6zp8kmrGqMX7TBux
+LrMgoRmf55rDCgbqbFPhw83b053xfB2aJSxpL1FPfDTtj9qjcRiSzYdrzBBIl8VW/S4s5JbYj5r
Cv/tn0VrTvbF5NB1z5RRoiNh1zKL0xRK4ie+IjEu8ETTyPo9WGu9lYwBMJBNsrzTm6addctIoRx0
ZjmL9wTkvKo5mQQ1V6orERxChgAd8zqQQ7HURT/xMpgQ+ZTWleZ2ODt1W0EfgEG+8WQPmiR1CITY
7sKc9I7xc2z/ZzwXiEqgp+xobPzXxuLYR56KH07xzkfGnv/1RQ4xaEflcSNPQeEjlGTimV3zqJaP
NLfvqusqoGTH/U6NCf8de+OF/DmLTjOY/ubKgIok1gxniu5z1YakTxTgFdlGuXRN4RUkGP+S0eKc
sd9YNDDRzcPxzWjHmg1kYpxz/3Bu4Zm/Q6NNbrm/17PP8HW+ET1sHVJj0S5jG/uR26TyJBNJG0R3
xRnKIVDft2twxwG0fl5G1BF1ruT5ojNF2WPtqs7yLNrS/KIH7FcoWYQd4fl3PVjDb/b3f0hvvTmL
sgJrAtG5xg8xMhGBlZl0YwRq8OIjE5MKwbzoQ4/Xb4svDt//Vmt+2GBxdbNRsHMGXqdNd33rIeKS
08yCtH5g1DNO/xFodcGAVmrHMrlGu15f9es0gpBHb/DKRkR4r5VM52WEzERSF0fvBUOtn1XFS/Jz
iBptJedekBx61KEEkp88oFQtFlbLDx4jDrPXfVB3Gttp3e0k09SQgrGxc0eGJfCb2qTIOroen8b7
C3DQPM6t0n/Kv+y+x7WAaiMmFWTKhjakDEQixCRF1tDFr1UrQ9cW/jiUAYMX2hPlH2FpRQqsqfX6
/pV9ZbzuVdjXgHUajA4e4CEykaBknJUvMxVHOPHtZwQx0KcYEz1v2I2Ip+ZpI8kwjTEEz6WOA7is
LgOLM1g2pa7I8ozJ9BxGpi1iZtGafGgrar3vXb6MBiIeM2PcR+2SqLipaNo35qQTaTMBSUDf4rO1
8Q3ksHoXTn3a+LCivMRB1tYKKjJLLVW2e154gRiHtFK+yb7+il+HzQSaLyJvTfLxSvtjYYTaQ6Ta
mbB1sCquECHzS0czjYweAL5QWqRu6rWt+loxRiM9NljvBFPefmvX5fKJD5IUHGCEuYtY2kAIiKZ/
bIl6WUcijK24NYoXrHEtAyZf3Cep4HTz7IVHwwPwkDSbxmvTo7K0GC6Bc2mZBgcb19OfG9crofB2
HOO9EU9ZGE7MENrtLutSePgG1W4NonzkWuq6tfYdo7ZGzYWlWabuoFKtKtxqolActdmDo5+3jxmk
0k782VXcD7JxcSj+SydUxsWBEMXY80tgffRzlDItwM4EbAJok2zzumOILZZi2JuJNv6t3nry1SsI
YYcNOb9wPee/PU2wh2A6mOch7+ZYr89pBFklE4NeSuLhSnluT1agMxiffsgQBGRKyny8OeHlzyvW
6mXMnHbenl0W8nC7gBnACIXXPPm6WUtv3+qGZufv9ppPRyUwXsXiRiAdjEto9EQs6gzEb/cRZsrh
FNZOjXiORLAy8lA+i8xBK0FufN6tUrmtmVR2arJ0EGKqEM7ydfXOWweOF/0q0j6ZHpTPwNPm16MW
qL46bYKVkZBgxXso9sNN3rHoGvyy7ylgPb6NMPApPQ3GlQsRtWcOtBjaRaNhpboxNLwiqb7BVMat
iENwEd1SfmZUCjinM2UZRVEabZM213atUTiaVbZbkg1A4vXFMHIjFGbHvW4ksEJke7NteGCJzl4q
u0WVe4Fke/qhmntkUgdtaObz5XNhHF8dz1y3FH0RQRjkgd7vHAvz9yJbNPKzyE/3eTcm0bqhp0YS
xBkgCRb9FtvGhDJnDD3tBZnGOJUu0IHUcyHdqBDgvv4VAIF+vMJ4S1xTLgXdiIAp/k4OJjSvhLEc
RRnIVK5DVhBBRYXdNwWTZqp0rQs0Vbl6Ke2ESkQ+vnkVaJfbWU6qs/T4DIdmXAQNYVJNBRil9xdT
2OlW3iMjJoRglmkNaBqNtYQ43hP1hMGdBwoBlvtVkELe447H1IO+4R+62h1VqFpOg5qtOV7aJ8IN
V8SdnaIzPF847mbYuprWDDFoB4NJhPlmq/VGW1INsx4JapC/M6eLCBPtAAXySgb+gkJ6SlCBpz9N
4vE1GLzKj4Fgvw8OOuBFkibo5kd9oq3y7EvuyOhh/tkgR7Xw001bU3uJfYwES16yd6rprdVcS9Fb
/mL7aCMKYU7i2CBe5GVn6Uzbodt0pzyuPoBpraxaaJnJtsql4nOxhsY7/aCXbOCu1EqGY8l3k57Z
DxHdTiKjQwnoMHR/jdWu7+xbdBjZukL9ry/2VqJdpqVbkfsvbANzn6ovIbTCoRuQqMDyWoQgRwbz
qouY7t7AkNnF3Rjpldu4wRGjPEkmtCWjjVFCHscEnwNchx29bONOFtpH/J6R1BrLSHFoqmjZKlpV
7xDu83JirWuQzkW6q+QdIBsEqjb6/G/xGzJTRRp/PakHM8B0wrtNJQ1jJW8d/XeSvdVBAoY/JokQ
+nbCYEdKT+bXwEMCDNm4nA75jzw9B2DRfKLb/Oxl4lyUDtkZrTcyxJbVaVg9lcfEpUR106kYZIs2
QmfvRfhBXhTJn/zkiBsjujyCcVCQR4HHb5aQO6ajhit5VtuvP5WheaNuzTpGu5kK1QqXI9rXJCbb
B9608Z2ReSATr1kBSo0xg20BoSWHsQ+lLL0roFN2biisH7grIJfSfkuS6GCFpH7lLr2lqo5g9dIF
TKww4iovX/LAPMWwcIng9Xo5xOhSdXLh9KnenVG/k2F9OcLdD7YzhzBOPrEn4Kh87mwN62yOWLB7
7g0/MmTg/7XI1m41DxXGsSvV6DHOJFfWC6HXdxdY1ZUUMKajXpFj4FZokgou4FUdY+FlgOr8FcX4
6vFYYziXxERYqX8zuovwL/LJ5WRNBOZEOxTiinv7w+uN+Y60zyiqom8Bvr+hjOzJABLF9LIkqJuL
bVY4EIAdZUY5BLdIz2b4/lKL0IMoePcx8EEvD1ZiUYGhZb9w8Ipq5wM+93falxcrcTRi9O4Ko+C2
1K9rGEh5aoHqmHVe0CdBrbVHqSHLJXDyDQrfRHh5h2Hu7lVBUiMpNFVaHKh3UDS4wwYyiQpkBm5W
51HlthRyzQcdkEISvZ/xTNy+2mIUfKC86kHhhSpaxmktdT5RbLVwuPqgGQwb5zat+wQXNnydDaSX
QVF/CfjYUPWFadwwP4H9S23Hj47vLugha1hKjk0OeBivI8bfHFVClYz9MNeO8UN2s1dy3GCcb8Zq
WJjRtBKwBOay4ke9haQloz/rf0Cofv0KrdluYAK4gaivUW5QpMjBQC/jCZNK/xuiXpQmd11jcs7z
VSmWWz23KeF94KfIhE6Nftd/jrPTgxCNk71cdROYisxFULdErb9/zsmYEN+9rqwuzilUEFlWAT+R
VsxYz70S350erllHg2owzCw66koE2dIW8xis/mYErD+NlfLqMjAG/BcIMLSW0kGg5UqCsWMXVjoL
0c/6RWsuenbdriBzIh98/mYLrYlK+ZXOF3KzQwKeEc1+CSx05PqX9f7gjJyP9M9dQFhyVQ3Q0Fyr
FfS7HEMtfigshqo2hsEdr217eapqZXYaDkce3+/SVsh9o+fSda1/OvWfxgiBPgQpKAVKzk+Xgf7j
snRwDW9wa0uh1mP289QTbJpMwuMVzBa3n0ekXr06dOXaH3NEBFN6g1FOZo2kzOdi+mlFk2nWchmo
uapgZIXxn1Lkc0pHEvZBKFiMML6iwoQDjOW5yjRNJrMq4HFOYyDbk4WLI+r5Pob+zcqFpXRibZ0i
Lsg5SyT5E0VylsXCHeRXJetIj0ljLk7fRFMDdJgagk39RP5VgndLtubhv930He0r+uzbKNk4rUPL
mN7vvs2UecmWicohnJUxgiXr75blheoPuo+PJUIR5v302obDfq8XH7WUIJvdCdkyQFUaEoFPAb45
j5NOMEPGzvthQXjfoSIEPEJNdaueb28cwrukIsvTKO8EQaEVXcD3LnkQ46QSmSe2UmNeGY3LFVv4
NgnCmvOwZ/5gezkS/sAza38gYsvOrBAJbLdWF74hLtfY0HC/PPz2DV3ii6v3fZqr/wkLc8ecD933
z1coKXNZDyVjbur0k+GUIP2l6bo/VEgWtiCmDJvC8YcckOFCfWpKVkkNl4JH/ENEUGA5EfNrHLtM
4I1pj8BEDQ9uo+erG80/WjsgrILEUEYO2qqvpeS9nSI2xTG2DngapCfGli4T/j1CHtm2Y2D3NHCY
NqX0AU0MP2PnN15OjTdLFuoAArrzIWMh0lcx9S51oPE26U9cesaVqt3oXGf+V6MX1Wt13kd/57mW
L1F+DAjju8E4FfY0+PJbd3CA3unLaLP8BoDBqNjQD4ZwERCP1f8i9Be87ujUgcoXAjswqTkzekza
JeaSSwPN4OUx9hOy3L+A54miX8KiMtVG90iJxW98f2TSakVxXcW/bZOvcwHT6/Z4yOucAFWifJnz
5wG598EHgcQcFNkoT1w90Jq4lrqcI6eiBlXv2261H77yTyJNGf5KrtR5ynV7/Wd1JiZAbDzO2ZjU
ih/a9qAGzWtqqgrwG8D3X+GYgeiSoPQJyVGdf0vA2Hv5HEVBL/nQ1T9M5gzqHZGjN55mJgpmIJw7
XriYc5NAEuW1DfesU6NUu06yNX+bk0SiJ1Nyy+DZ9zLMfgoxzw0smmIv5bMcbeoTmGR2R7HiVJo4
Rob9Jsac7GlP0+JfbWqL/7ZAXyVVxJWBCe1n7kv3Uf8ZNF3atTJkvImMkDmeSuLgUeGSV3Mgd+Zl
l5mvIc+Q+qOxh2Uig2wsvK7N4ITmzugp+5Zx1hMYUqmmqJsy+kFQddis/K926W4GKTDU5sVmX2sZ
l/wIPJQJEpro6jC71mqFug8+MktA6mjAubVTMS8fcdtqO90N0+3Qg6lOdXq82h/c7F5OPs1cEAs2
Nzi1m+RUSsms7vecnGpObwwsHevjw2Q6FCBINSKgwfVBet0rR7KESChdY8Rwpzwu/x4Uz16WGmuf
R5U7bf3tpPu8h7DZoAAoeZDgKS3jlwzxLfTrPiuN7zl8Jhnn2ijS0sDRIPNbteiqfabAX5vhOg6+
cV7ci66arxUbT9kBnbD9sL8mhSOO6bQzn0aYqnvwXcaqQr58Hf1QpHumF/cleIy/icU7iYXiBhUH
fCNV4KTTAfnLBaZmvEt4nBaPXqLn/D/lAVl98xDnBXV5ekABE8mbqrytqxJvU9Wi2tUazXEbXjt7
nFI1+t+ufZ4J3Zwo7pxnv6meeI3tCsf1Jkhvy2w/1gRL+z+Wa4H17HJ/rDqQiIP0cDOp5c83vaiT
ux/SuCL8RvIj726YC6vBeLfnL7Ka1EDKYBt9JgDOpcnDFru/mf28cKCoCv0NQLUci+7zgXJ+PZSs
ScRbiG9iTwgcTaTwbmz+k4ERAgnU5uV5cQ8Ul/9Y9yU3tZJ0QksZrtpmCPX0Ua0SMM3Fm3+xuuf2
Ni+UHMh3WBUByPwON2l1o0HLJzWZB6N2OnTLyFaYputpUy6vT5I5TUZ9n5JvV+SzJNmM9vnIHede
2OXkMvwKrXsfvk1z7ZhocYTuqUcyk2S3KcarBmMkixPOebAJEWPboswxxZbJ8wR4gIFYnD+qoGg4
lIWrZAi5EfgYCkqyX49HC0wu9fg5IT8oZDrkHHrgKQmYG7K01oEs16BvQyiUmdppwAOZuUKP1c8o
w8hT0Ynohp4q3hcaiVLIFM6cSSeihcrgeBd0f+LqsRd62X7CS0FilCVQEzV4XaSEaiHnSvG0tfps
cg8kELKev3L0CrWwmlkRbY+uX8evaeFuztWWhsbUVPHU8oVkHLf33m7T2PFU7g98/JoZh3gdLt97
K8cVue6BS78YgPRpy8pssNATvYIPPceoqO+5+eV4BUV27/PB4mMvby+4L36/MeK3RQTXMI0By8yq
N+AwAzTYCq2Ly7qFDTxIrgYeP86G38QDTPk5lGX4mYECcmUl6xIl71M2hAHj+bHizwa1OhpSjHW6
Lvrdk4h5ZZYBr1yCl3P3ULXqS3/9wjEYue2YwZUJ0s5GHjfyuwG7PueuVFKiAhr0G4sRCkii0c9r
1tEjs8x4aiC34PW07Pmz0uVUUU+avVOZYkYUGdoddeqEDsO9aZ1SvMhHXSsp2Ah3adJvNS6si+0i
I85g5zhwJLbdbb/GyfyF7AN1CdlJGosiod7B5D44G3qK+smQPA3SCB6iP43okpG90ORIPlycSF/3
ZdmIdedNFuaA3qeJdJXvO34UpAIu2vMByzqI5Ma0pvUfJSmUeBAwgeCbO8x8UCF4+cdJo3czXURT
t7ZWoW65QwpVi4zCI1wbsH7fxaL/u87A+BmgTYS86h0CXp0ihFt9t/NHl/5pWzkiIshCWdQBfSvN
ibf+3dL97h3cnbvU0zwrx0QnlZ7JLvjomr8c+sD9kGAA8lzqGAMiU7CKHFHiQLb46I74ntfkzIDa
G05Bv5tGQuoTtuoB+R68ZbViSjF5Hyua6Lnz2nYHmIfpFu6mFSJAjOCayGhI74c1UDcxZFkoSLTc
TOexML9fn7i/h0nPUTgKflXDNoJRl6FVlYwUM4Lmhwevd3hOB5L42Y4ANdAmbhuMJnjXgPw5aBDn
kCG8buOd/vwjfdEWxBzNYHEhczMajbeSa8Biq0wos031xkSACmP+2GFwGQRk2Qiv0SIw09dpPkF0
OJEi29D+cKTrZ/qrLktPLjZ40FTBAQNWsww8CGgE1+rqH2saC4ITUQ1eVucTTKplDM7KaBHmVdX6
Bf/bspVj/74rYreDJIdhfYhVfxRWqrqL0uaK5W9x/MNevGqVwjCFzzbAmsZwYr0s/+JGKYtQiftB
4YZRIupEygY3NgfEcI3xY7CMKZh+NyLe9h0srv3gN/EvpYnYMpXGY5eB40IOfOCyR3zG9e3jdGur
IcoIZP5AyKTgdizBpSIHXVN8iXKy/cVcRMs38LjyaEi8TVSRVZFnwIu4j0n8osE7ZzQMN3lMtuza
52yRFdha5PlzJI8HXvvx6G41GhURhu61SvS7GvH6yR0y7t0vMZKtpOIk+Bhdm5y/3vbn01hVS0Ie
H/VYM6FEKUruJo1PRngwvxDzMsTd3pQe9HqvnyZ/5CXD3HUZLEm6ujjHo+VhRItLT9ydkKksVA8t
SpI4NydfP9ySLkfKFWDGjn39a2Vg0wB+x9Si5J454c+IyTbMrNm7B02MBo4s2K0mLTlC3HQ+BNl4
EKKG3HSfEoQpYzNd8UWVu1+vgRi7JjEtiezKlskGb/dGVxz5sLk4hkAvDBBhhNJUfka8qeZHEJvP
nggkCx4wcVqwHdJzDSPFQLaW8SzfPMmGwCBuU4sswKKMVbws4HNuJr2DT8IumB5FCgwRmBrrfrNn
a126IJ25pA7CKwXawoDXEWKWU1etcAoBVu8eTKI2YNXghQg0rSCHpGC6wLratud0h5Gzq6+TpKPY
Hcg+J/sL8KOeabOqQhdT7zonh3Sb5yUG37BBpG3N5BmuJW3RVPePS7NjleaTeGnlJfuSpyv9ZXGd
DwrC4g9FTQYGSPa//bwR2nja2IHTpleUyrJZp6/ObgolzJ+t4ShlndQWbdzkZHOu8GzcoPPxo0kC
h4L3k+DzSjjvniX0knCk5JKDH/g01VyWse/6vThMK/hPPrRb0GzUT1ut8KxUYb31fCT08DtXvbGE
DOGTCjUto+lshdw+1bCpysHQ+6yMIj42y5sz5AvkCVKu0xa7fQ2frU5wzcDXir8Ai0JXUqtn5Gdu
6TdUaPgMHaQ6S/S/AbXorwOcgdYGEGpsJVVHql4Agv39WOAS4ulc/tFm1pJQZE58MmvfTOfL5V7t
u+4Z9GC43U32eJELLToXa6ouNLO31nCTMFRjtbtuGFut7ACbjEfZXIb/zxWAQ/1Z1X+O0kcy6I4F
QrJ0UIvVtQM/Yp81sLjdJLfHYrr0XOm/Z0GkWs9aZ0uHz9ZUf1poWIA+WBcr/q+AfCAQZlDDU5tP
eSlxigBLVfT6gbqu0gZ1QSgQVr4ngvN19XrKy2wuE4gFmeO2g+A9q9E2Scv9GDUnWxS9SW36VCJo
YklQNiH+99xi2Zz3+EvuOuvNJFa55CjYMPx9pdlYnKl17k/R8r8wYATpWpi+9ghQFaDHuwl2zcE0
YoEhTTpCt0IgzBnoLA6YJbzsvoAli6Dpmj6svFrYScJ+jY5HewbLBnaWcVq6PBsTH3O6TlvO4AnS
8/cFXPK88udAijYr59n6DekDHrazRghksWRZIm1AQBa/hmGRtJ99vxJ/pzdgsDc45v+JD7nR6O7z
I1fH4U+8tjcJW59kIgLewQBpjBcLXQvDD1IfYHCiszKXqgM6EfN6/1x7fcmp8OnbFb/P9uGblSrP
u5YnTlBYttI7BEzdgu+eQ5OjeNL1JX1mH+6xMMzxNLW7Oa+BgQJerpdQkvGE0DXbjnWDc3sSdVau
fyYP0wR/rKNWhIywzCakELmfCjrsn8oUGp81lOrBd8fJjHuOCIhlz9kJ9UWp4vwk7dzF7p8B153C
0/c7QSvZJ0kzuILvEWqlnTBDpTfcq7Skk9svNwwHvo4v2UOU2tb3M+QcSBQuOjwg9PkHGu1BXOkH
oH61Qpt6Cbb5CDSsz3ooYTsqnDe5hnpWw57jaeZ51nyJLTq0Droud9dbpS25h75oFtiJVU5gzMVC
jO7SZpXFZvBD/iVvEJc5B7OxmOJqShWa3mHMcd57xuBYD3g5MvdIMSC5CKIyrTbZCh49ThWPwXv8
gqhvX7j3cLD2+yamdVI64PDVAtY1FEAhxBPp72HkNNGq3Hq5a/i7/uu8gl9swO/Tw6YZKHgVbg6B
SGpv48KJL6xwLiM5ts/sTCfDRK65ZyYL3/ephm86qx0AQrvsgA6ljRvDRXfHFl1kfKqYk9R2nFnp
fN9cQWAr+afracjTEXz8ExJeTGnFmREU+VB26mj4gHpbKPw7Aseo/FHjkJe9iXp9/9y2m8TCI194
9N4E4HYyRlx5Vqyvhm4beyXfSrvTl02al5eqouprRaFrbnPyWTYyB2CCfuiYZsEjmB3VgXKsoGar
9zzap6LM2BsGZBg4fEAe7iwwPLvbHHT6CaBFqnDYIkdI/IJcT0LFssichuV6PNzmeZNMa1wC+SwT
KWRtBuMx21zaTGqCBgK/sRSK1/7Cn2EeElxsE/dSIOctL5mNQ5dCABnrmTWwNL86wzGQrUJm76V8
CGphgZRxP6CNv47gU6Zkr+SDLvJr8Hje7MYvdE7tINLLqGAKA6RoVKB2vrNlHah4AaTRNU+oobmx
/5BQT/R6xRs8AwuBn+9m97MLOH9R57YWvc4mvgIvqbjYPvNA7neAUHQu2P1zDxUoCNsrFLWt4FX6
w1o+f5Nf0WBhCGNcFQfGbj6JSDM2NXwjRKyApXOax3cTKw06fv3y2fq3zKiTPA+kqDXs0ztJ9szs
4K3iA9C/xxiW4mm4WUp+tWloFktG2XCEydEr28OovJO5btzqan3O88pJ/YbjPj6U8TnlIWyXrRSb
oRiJDWEfEIHSQqM406AMbwMoMiD3DPMglyB1CDH+ZmYSPOVGBaeiC+lnHyWINY9LI/RQ2SAfmYKR
l6Ugh2U3Mn+cxflzUECEcwPA21Gp/CA88kaC80YcKcxyucEDu4zKfNRwzg1q4W/+ANVRjXq08nmO
8VyMyMlww0Kz0CwFYjNevHMoACWI1nYfOM/OHbrkVdGb85yfPZ8o78QqXuEDYAy7z1QJY737gBeI
BZKA12l7lgaenYCVcLHnDnICTbEqJbLWfJpNts9D4h6siLHklyg7N9rPrTFvUr7vvzDa4Km/E2zh
Xkqt2WgHV0+4yyBcdVekjrJTauA2k0+WCV10er5J2ospgRe/JRGK/MHRYLQDGgX2fWnhLWL6FIu5
iDRpI6XiYUXWhTA3lyy/B/+SKtFId/kgW0JLQpqRoTLD0oIFMxkUuIIDcolxOe4lbRp7U/18CPNb
/hsuvU2eIdZ9unqeaWRLzrF77HYI4HFBSX8W53F6HLgCGXhImVTfdYHHfuOpIHwn7mt7ZsqBUlMN
GlE69hC4/DfvQ6oPbBzL6GyT/ncyqa2vbDkrhJ+AWAGgMC0Kdq14afW16R0omdSq+FzMbCf2wzoH
xS18gJ+8NXe/DBCJj7DlkkmmjiaXj2yJZISPX8GpoWWZ2B15Kslsd9u+Qlu/cInCBcp4W7fscbyj
n4EdVOgFi6u3qIDuz6PiR8p9Ha2Ee5DM9gx41s4Wb14IWjP4rumsCVoFCk1IDLdxwTj5rWQi2qdp
QuJht95J4fWm0jxCXi2rgr2BtNfJfOb/8QZKtx6Kdb4mngd/IvHtJ6MsKqO0I/KZYVGUut8nWiXN
styip7fMlagXjlP2oR099373+B35qDvW7187pqVMa6zDM6+BnyzBLgg3f9d6AFV71l+jV3cnu4wG
i5/td8hGNc7LlncRNqVbhvuubTMXTNbSUOihgIINWOtI5VKf7D7GvxFaqOE1BcVzovQsyeWVMpvZ
j+0CsHRDlmpJuBPXN1oJUJVU4VkaMLEakIJSqBAXYEJp3Rc35tm6t89zWBF+LhKwX/vm4QcHDY/I
Qni2owENGeU2HGLnCCN35E4d89xe/J/E95/5fhH+2aAJG98J3Efnq5aEQkAP0NT/IgamqnCPVHwO
AvtpOEW068R3fvJNCtlZzsGfz6ciCxzcHYa5WTKoJlVt6dJ/sDoL3RLcnpO7WJyeEaHzH5tQ5xUt
19PvqdOsZC0jEKCeanZItMXnr4jPG54tHq5aB6CbqPTcHjoLlOFeYNIdPuzraU/vHO5dCePe1TYY
etYjzkFyREmpQOuLgTJkFPpMIocSghAyS/yTnIwQ0wbTFxeJMYtvkn9ep/iwb+4CREwHlLQyPlI7
3q+018IiFJ2D7IMGIKFpmndkU8jVBjZYhDEX2H4efUFVF5S+LKgNt3p15e02djjxTEIDCXCCVUny
VpTH6RaS+VEDiXwzQgyeZ63SZFSviC6pc+u1WLczsv7G6umrWMRHqJuUm1b7zgBn9ip5nPeL14yt
LU8kbOMfVosXKkJsL66qBsLE4MBodlmTzPQIpwoYiIbLDEEltZt/FmUVdHnFN2S5jc1BxgLb4+or
YUJXgnmxNIY1FyCIa/NfqBISO8iW3vL2lDi0VlPMDmUkc8jwPDzSEwD5LXfgVvJKcTi+74Pu4O1i
GrP1s+MI2wjyDJF3eabqZliNdIJW5LMVAziHTu2eQ725D8j4fbC+SSFPYgMbbu9rtm+MR+euyOhj
BZ3n/cYGEk21kgXYLUtDHJGV/COxo4v+sLic7Cirj9fpaUq3Hz89mjRoD7rDxxIMg2JiYMuctHiX
N/s8Z8s6HLoVM/Pe0DxjRpov9/azL1NE+KfFqb9JirN1vdOMm+g5FdQ2J8ke/bN5o6aB45EV+7Tr
v6SKbUZChiYYrWxam/4eo32CkN0+Ont1vmLQ1ZZzNUrEeHEHwHRITJ5MCLvs/LAOA5qvG367wusC
g8JwG/t2Qj9VGlZcG0ZRqs4GDMCAtz5nJ3J58nwO6ty2T+HzTTq4rgT5a9+DvAYZB+E1E06mcUZZ
vWCNz1DjEzvUvyz4SyF5jJIzksfEnUVQPfpUaENonmvHCQ9YI5CmamKgf78w2rJ4uQQLJFyvCSg0
SSmjXNLIFC96lWpPxBSUhLCzpEIkEM5OEQuKCBoAXTU3Wmn94vjp+70TnK1yiecPfSisTqoT/fDR
t+kBHzmRIikFul0U6CL0OI/M4hApI4r3WS/axktPOKpAy3dMj5g0ySQ18px24zFsIsE9gcM5CD4L
6c9pyYGC8DVi/lpfHnc9z9yJJK969pa/CpORiTsd0b2eZ2ZsgSyQ5bg+8+gwgiEBjpC8TgnhPEbW
GjZTYWFzD6yQIFZeP49O58D/Ir6r7Su/OX18Vs6PiD+zPIohJaxQtxz6e3fM/u2TG8orbmrbTom+
Civzu1zD57s5rPAVQiEpCIs9LcjTlEH1m22h4FoNa3S6GsRV3qKMYGs3EEc2WXkMUmRCsvv9acgU
uKItVPsUabWclaFIKZyuMiAYRZp37Bin8ZmF6jxwH3C4cVKLKKDxb/fymJHwDxqr+Pno3uwxywrY
F6Qfokk4KmXlIB+UcV97PWH04Jz/cGDyfNzeRXwAKLXNHNmfYV1UPVZtCD8CG0o0SMdmSR2N/98/
cHdbtJmEHDhHjTo1xMxMWF3tr33rfqJXKT8UMQcCG864B+u40qD1yuziju0LTSH9AiapWfxhXoGh
iJ1hwGXJoe8/JJcJJIhwziLt53zjn32ZGOkJ3kNzwkxVEeZKFIW8sWx4E0eK02YiXjoWD1f6aETT
bWLLItaXdL+IAcDA1kaJCrxghsjzq2OARN9+KhUPHGEAcHPDvmhhU9aQzBY7iRnmbtOzfkxVJq8e
80VQDiXpzAdCUbu8FS/m/zuV8zdp9DgQJbCdNzoByeowvcsP3daFyiiA73qIBzkDBXm2OANANiMg
KfcrwWBNfAX7/dbqP9z9JBDJhOqDDosmg5NrELcy7EO8sa+6KVhvfdIjlboC8x3bYaWszb9L9UDS
YmNI0WuJzy3WnvI9TGOpsOZKvS5fq+8tvTFYTZTVA++eKi7P2DEye6FNXXfJdLE2g6SCt2YdVckC
cOE2FS1+w8jCCwADU7j1MhkSTHkXFxqPhKHK8bgTSGY62B4kj/xxPxyokNStw0jzYPbV/SEpxmnP
Obht2gL31qZAnRt/Gu+jPfq5RskQy1IOF8ptugQ91lZRujgYt0Eq7CrCe/dQPbdJlFmfG7EUBVBE
c9wE3kmJPpyL5bLdIiPNVr02RxtOmtnUtavTVSgVrdBnsy+VelOEHqoD1DJeWtJlilB4JZkCMR4O
kYE+xeCnOLCeNZGouKK8xhb70LEqOCaeeLrnT8NOMDKspH7173eJ/iwpwkk54tTW6NXZkNBj+Qyr
6pceBok8rS4eYxiMhCdiGKvPdfW8Z7i6620m4I/o/mzznH/q6FOub9RaZwFxvWiDSog7KHZsY8TO
OYeDeHjk736G2qtr5K++VJVtNHlDWdvaO+m2c1A1GPjEHxWQ6ZJDFx//KwVTzOX5UXH2XA2edZtk
qjZK0XYiG6olkW1MobLTmHToQwfxpKBoJpghQFIcXYGo4S/BVThcRNFXjl96Mczr88FANccTnPdq
xQrLQtvQnaC2CxVVzRrJ/lm4D0VpZWve1n6e59m5qOfKrZNW9m6I7x1/xUJtiD3VZjesns4Ow75k
RjqJfDf6PvzfrcXb2ks8mLa0SveHxVv92WbMJHA0NbVZCTYoZyjTHE9j0gD5YaqoO67VM5xZhdMN
slvZn+16mTUwGcY3AIU6nvD4wDmt8pIRdzf5ZticCTc0HH6/uaJ5pFwDwhG0EW3TgOwRZmqJYBuF
LrnIZvn54YWgHTjvU2VK4MXzKNLJIxaxqnlizgAvWsHM8zvqtEV+i7lhjc4H0++LRjPNmWeE8maI
F8OPTU7pGt42Pf1/KD/Q8n7BYqztqd+gph/I3ZubyGtzw/A0HeS+V5E9PjskNKL/5Ip9Q4e+cfP/
sk32a3GQY8ULCdjQLYOpcSENjqhhZ7yoCtjlYb1B60e+PDaLtJWtkQImrIJcA34DoOFrjCns/FGq
cygx36BGkFPIOhoyf9cjw9iQ4YQbZ0oa7BVhuUy5Z9V/MPWNlYV+s0RZ6nfHwmZqV6gDtygYcXB6
ms3vELkcrPX7DVtTd3EoYIqU+XiY+2JBhBfGyytmauSJGLyQUObBdFykIokMduF1glWyFvTKdJqI
MdFpiffbCyiC7A/yWo8fWlqrOfykChck/ca5ilYfvZWLFBTmqISYaYcM20msDWG6b4hCYhMyo0yy
ix7KaewLItRMxgysDKieDWFyQC3RYE+1qr8y0+yd/3X3N6eiFho1mhy/DL9+m+K8q95iHSXuFP81
JpmX2pT8NxtozMa9tkDVgZFiE3b/8ApX+BgKtLQmHqCculcSwuOJJG0nrxrLs6HlLHuuUElEWG0t
WxQGnYm0Zhijdo9ll2t+/qA7tyFj3uJSdtfNtH9A/L1Md184+PMRMdg2Vk6w+QUtKOvipkOsytw0
lZmrn7aprY3AVR96tDbfuFkTf8xdPIrPb4S0hYwlDp7wNGTYsPBJxxFQ0ewuWRYjM7pzbaAtCanv
MUjdI2yaXUY7cetZ246Lb6ZvqRf/fTe4HLoTdu52WS2xpHDYBPU0G2RaW/roG129MF28KuqloAY4
oOmhDb2BC/NXgcfT7LwhH9jtMo4gOE6zkApkWXdsNoc9sqoijmBLyfq47LX3Ev75hl3dMNofwvfQ
NPrIj7ObIRqYa+0cAjmg+RA09xtM8mL8y0hqNTIcv2+K1x5qY2WTCEtqyjnFvn0K14HyXuALUbXg
jZzuPLcY9l4WM4QJZepNx+bEJD4V71yp+sqUFW6ANBKBA/BITeaYiC0i+SBAstmXBJ7+IEGuJh/B
gH5/+IJM6GrTmzSrKPf97uc7GUWqGn+PKJjZxx1Evji+ycVSGV6FRezfQte3uXfIV3JzukNsFwzO
nQnELpDOkv0l7JVEAuRAh7d4zP54t/Rp/alEHXuGr9nd/V+sOncRgRTSrx/BltqLeYSOiOM51ycS
jxDpa8Bye7/WEzS0XJV+wweSrTDVDr5RqpqwZZuGjARfNSavJTPkGJEY6tyiTgM7lfH3uQPt0GLw
dgpQhzg13X4n+iqOw2i+trJ7PeVmXTJLdXcaWvXNZcEmKrdeytdMpvBLVQpj/Odmx7w3f69pSfCQ
3POxkD93pQekNqnSYDfs8tPbkuYqLM+hSmsTI8jH8aPXAyBzBeoudJDAmhgGjHQUH5BCNJILQT2l
HxDDcgoajknAI6G6o6UbO1iJBY4QsuttIYmrgUHmpJvKAwYmX4bUpE5YkZHFe7fq9sZG9+uVknoY
X/IGMpSmpbV+j3ez1vj5XI1uI+4ltLBqpllIXIvcTh9oYhQ2AiBWpf2XoKeeWz4lzbJLMNMcqnWQ
CZDb9mKE3DVGDVMNIgXN/UCK9a8P2KLytbcGDZPO2HkSLLPkpesQZmgvxPEIpJ4t+H5y4+7arxLA
+T/aX1smX4kV7aVSJGNAuUvKV9rSeTVLY4IUDx9OtU+KyiCcx2S6ZI1pfMXEE0wzU/qZriPJHD5W
7HU/SHVRiF9ur7vYtLaNRjr1n9KrMpBldxDGj2OaxsfYCmMXjG5UQEOu7yrxtIsbYMso98epITo4
YCcLOV76uVORa3fgLjzsXXzvpCfWzjpZH8lGCmsklu5ybP3oAO410C7E05JixQsJ9j6z42wM5dpR
yqSiBcPfhfMtBoFe/A8ImzAO5q/DdDKuSOoNYfeR+TTnzNzFovkaqd8/nQG9O0JvJnjJcuf7V1HQ
nvemxzHMpuVMMPgLa2OAonOmGYcxT88hZFsrbpCCM/olneMbVOqog4V+jormJKp+PkxSyr3sDY8C
Q0raL05BhwIzeaBQ6ZB3ToUoDdrSRKwgNm14kl/uiZS7SBOd6ahaie9z+GMXqlVwpzrlukHcvB/S
Ows3tHHAHLcCj5w2X/MLBZcSOKy8C6sqio736UGFc80nIfkmh+VNzP/0/TNPYhJWRFvwFABW4c5f
Q+OQNVUhBap1Krw76DKHbY/PTddyaIMs7j5pu7nlXzcuxFo4z9rUmj0/JqEHYGH9To5ArDdi+xrE
VEIeg7k55Ub3ExUsGZj5KZ4TGXcZMISHitiT8L9YubPK4B1UJRsZvJssSr/Bm6nH5v03msAJza7j
xkidMGx8GCaP0qA5kOgJ2TfLhcy5jEclxpczxvlMVoTtB78GLyBNU9W4Ozgo/qYjtOxgVzimJ82u
V9VNxs0MvuRwg+6m2UR3Tpgv4StKgZS9bolUV+7l/kEg6pUeC5QTPG6lSbOIcjV1mAFkYcfcSLpC
Sc9l7QboMCvqTtsKnclvOhuKOXsF8mWGjOSCTpojMwwXVN8a1kuEw/hIOmRvq58owwBEaVicK2ej
PDAKKiAelzc4Nv23ezBcG0H0u29R1pd0NClRM+37h6AcgBv/8zrtTJXu4wVSM3WMbtsUK+c2OGVg
FPE/fdj8p3hT2qTMeoNfhyQCBmKtj2+YgFceUIjs6UzmE8VHI5tMWdnxteJc9Qe0fMmvjpunXbiu
n/1eveO2Wg4AcKB4dlAdu8IrAuCpq96PqHvG4QU19PjtRqDMnLE/X0iA9sr/XS8djVwfphXVg2hn
ZO46WHyfuYNPLCGOrBYyp2/XVJCjyYSdtdUjgafrT1MGixnklJqxi0rftfp6MVj5AZWvCYemfRrJ
UQcahF8KoRxEFRO+UJ1bm9cLHatHhFUS7r2rxtBF561916eCt08Qm5lXat9KhhMu9FzI5QgtEzJ8
3TDy0BzV/BPhwzhAxoMxwj1NwYcHKXLX1uD46sgORbKOHkxiRYvXIsny/NpMfsOFnlTezzIoBbuO
ow0LSgO31jD3SJQThBT+sdrMHtMuYlnsxVPMR5+17GHzl9Ly6YRSmsyoH0yJM77s36qF0MZiOCJJ
+6zR2LVxWJcUND5AAAqLh/fghmL9IbLsF+MOo62kcJFRpcwM3pioc2cZRNWGWAfuZ7Kuy58mYlmR
bowfOhrcvCJQxoof3z5+k9hrrhkjL/9Uc505zqyHMST90izwYI6hoSU/h0q8DSxGSFJt3K71eMb8
2qdYv9KWtR85VNRgsr9WevonvixJsmVCeVLqYmoJjrJ4vqrYLscbs5PKqt8tgHOv88+s+kV/4MBh
HuYTa0MAaenBpOxwpbiOTAoxBAwzxL/pd6jww6I2Umr8qUbtIbzdV93ITcIRy4QfPPIDDo09no4b
FnJ5RVghWebLkuN3KvG21DWaJiTNb/1VRzhTsFqLSRbdkgAA59dO8jKfNeT6o0k6Bumaizar+zbD
uOV365HYAVaodgN2xhdSXVWQaaxh5LvlwSyPGjiZYdjGqIvkJxV2g6ecSOpW1DMfTjpKIXVBjqZu
j60mAYG8gGLvhPa28hnyrBlvncSTW9C5f7ovU8i+SUsL75PXvyEwUM4D0KI2pGV0Snko65GF7Z+o
CqR+B70zB7V/DST9ghmmSkh7AlrD0y7VtUniP45zmEVVA2UL0SnaBoSXU5OtTdRJ04siDy0qjooF
bhZEEL1W9DRYwFLAqLXLdt9uVdFTkObxfUlAZ5dnadoylcBYn1jSnp2Lj03wfgSmLSKmhiSTFebU
vSQHwgQswntUfl1ov2NO51Tzfu0RBleNs46b/TbA+5RSazDJ712s7ykAtzqRSJl2AviY+FCt/gNn
LDuiJP5GVMy6X2bskeUFfsJ/QHoHIh6s+rYcYyyf6GN6QOVC/rxGIzBy26L6F2AhhluE3WN28zqx
WedsVGlyobu78l7RPh6b96dGLPwi2vmwYDnwu89oqE42srjVjYyhhVUiht5hXXQMY9XlOK2wYQkD
FgY7qb/7S98RtBAqsJ3P1wEk0oIX1DXww6+g/nCYonYAB2Euxl+0w/479QrcYA2KjPtjP5Z4lOq3
BdkSZJXc8d7+CACo13mOM4+XRkpZMOpxqrJ7jeE7N5x33jUyzCgjRrWc1y3+n1/dFHwIZZ8U6JcD
N4SrmZvauSe4tgM3NBk42seBCkZmP/L5qZBZ04xexzceDKeVBNY0G1voeMoRWTGC7iRztkxLNcEI
J5uLEHYdU9BVN9ja2Jtkh+d1bJIP2InJyee8Y7+Qb0RZmGuOB5OClKQUEhEgB+LIjKDWGaVfv6t5
dzyi1TWeh/evpM1wfCwJtME5FVPDa6689MIm7aXbzFHc9hTs6XqFe9UcFPt3aBiYmjMEHsDiEQMG
NhQjWs+M3v9SHz/Jf3uRQI2dRHkVqAkqqFqLfOE977y/ZCIZ8polocWO8a9IkaONPS0r85j+9IuL
d7AztYyVuk8JUcetbnk4JoLEUYjqCsC3zcWjoPCoHNSSHdPLobrkEz8n/gvZEr4KPb/tmZKYEpRb
OMERE/O9s0UliRqEUg+O9jjgoDmyd/seAOKFCArFdSR/B68RJjIBFn/NS9sOKabT2SCx7ZY/hVGV
FBmxDcR/nIWwaKevCHn88KJnDkS4BbGx0FwmtF7j3gZzRWVOOvgQ3ho8L6+p5gmn/Rd/M+pMl4i8
TX+V2ioS08okbDkhz46ggvQUR/LjOqyTGyAZELJXTXNHTEpJnhNkKrSaDEiIyfdfd68mZN1/LG/B
Eg7QrszAW1UGyklNtReu+Qta5ADiqSOF4n9eNdfvNkzL5n6Jh43XUL0TijBC3drAU/aS945IG5DG
XfmH4e7MGocOOeXonQtIpPRYLBJISNDc8kR72+RIxIw2G5gKHPRfMlkKhS2O71P07R7/6VX4tvax
ttiAcxlw5C2t9gYKa5YV1Z9N4zHh8nAhBWZlXvcibFzwCEY1uGF6bJEKz8gHMExwDQwKyOURLruA
gJ5Rss1P4yTXbdzohcZDWAiiANMG9IKRQRE+WXvZJhMPqVvh0dqoUAkLQqX29P32EUs1orPeIExV
dGJOqvpcV1m3p0LiCxBlmZDdy7GfK5xdsu+ga6cUE7ubSuYc7216SEPkTiolZrBCRjXyEtPpE9LU
6k1SEgNCz3+TwbzA92vPmRaati3YmRys/B7pEYw8BwBnMu4cdRKxqfHysJpSwFlm9073F03iE+5w
ofZRkIIsaMpT/2S1vewQcuVS7u9Nv1fcoNbXbM7b1LvhQUIbOeTghvbo3bx1V92rqC1Z4tuvs4EG
giIG9Vcxle3tDGCebzmYUaBpf1zmB0yjrUGmLqvvmp6Ojs+y1HkdmuAhM/O4KybXx+QFNFeMC3zr
FdJe1JEi2XXVrn8zXWu1iPGsQlKWHBLPMWglgZlsStBBvk3bJ7yGqRWfz4r8h3rkqhbVXsZaTdCW
CPlmbbOKcXSJkM3nsltFoV5+HzT1Y4aaUDH6048V8iHAddDDDYQUxiexPW0CgorwmXpGe0fia5Sp
qFtcE8tWB7oBBZwG2YZzDnn7SJ+Pis4yu6DXSjgzkbWC5d8v4HyY0356pc+HEdgw85+q4Nxu15Ri
duBQflDNOnRnkayB5aQlJBdNEYNwBODk1939ItZU9WIkblCMuDll0/UGb5PG1LMrgkrlKWXMp3TK
lxPMR9Wb3FSxZojZ3J3tuPR/GuvYd94EYLlY3QbspGiSFBkUhM9t3C1rm4dlf5zUNL4IofUoBgh0
e3fLkWuVobninT+0p/6uveYh76HHViiCIXT0F8TrM7hA8h9dscMTQtKBE8UhGW6p939aOUnEA8cq
l2rDagwVIW4V7QPjmBm1LEz2Puz02RMkNd3sxf3BU3khlRiR9cr5vHy2l0L2du/Z6Xk7DINxaBir
05Qz2iovTGF14IM3XqpDAh9DF6VanBzxdUhQGcpexiKY4bzxZaZlimQpwn+SOP5jCmQ8EM0DM5pe
aIgfuAe0URf72BvvTxJydtneE58zmPuwTmdkYeP+Fs6X7uvoWxDilhceGrja6RoF61L8Ps3Even8
pjFrlzglydO0LbaeWMilXY+KiJ/iiyxbCjxGT3wp73VluC8nvkLQnvaopnOCUfdfgIX2e6Dy3c5n
hHrCcvFPQ/Kl5sJwgnbi389VNjzl2NWwv779XzjQtM0Hr7Ayi1YpAptYyYbZPJUm5BQ8FRE+Ycm6
srnhiHzmZ5Bts1CxSfHeSSbS3aAxzdtxpUNnHYoeYygb1DwkkgtqU9jdU2PV15lH4jISU+B0z91D
77MTcsywoaemN6M0UorPFVR2kFf9cQ4AYqzs5+aiJSJgqyZZQhA6s1PJ+VApgR9xspK2Jn8yEB4v
I8bteyCqctKr3zchupA2wJqYWT1B1bbI3QVY/uHbmVwHbuikKuWNsYqKusp1hQUXkNbhVQqAsAsb
3idMKY2UoNPI4/lmPk13uZuISDWSunwimr0hc4EVNmC40/f5izcJun+fV24kVqCuDpNK2lvMwbsC
e3ZyTWC/RKdy+OVAi8RZ4l+QZRe1LmZfvQvcroRqkbDjFIuGumsSrvcM065QbgU/KISVMaHbZLTy
LIuKAJhG6WEifN2PMN0hYH2n/sf3ns+Zf6JMBvdejKjy3YzYS/2DUr0yTsOrBqF1zIRnOrFiSEdu
rEouIAD40WzuQfIKsVdyK/EsJSZBF8ERSlDBpJQmlkC/FCsqCxw/T9azT7sAbB8q99zmQ+6AAxBR
07pqWIf+e7D8cW7JqMFscVcZ/IYC9Fux7CkDpStGFTT3yKjuzqlC1PaaNfyLWXYHQGA9VUIMJh+Y
eNZ15GgKwlsXlXIgS6iTae4h9ZGx+RhigV5OrZ1IoYi7qqCLKhCmxvo5iTyOUkVtgTFTegWqKI+4
JPuH4DFl9s/5QAVI8aM6yxKg6jQtcWyZwYDNGRAaK9lFxkfGcCMs59kUC79pmpPV0CjErO1pUb2m
2JrYfIsoX53yuUePSeYrnxqt757zwF4I2t92xTIfS966etQKqQ3YxgZ8YnmKGc5g73iTZyuc8FmA
6g6hjkmWZmCXQOTu7tZQ8HN2oj+ADMS9lpV7mS0jRQRWyoZi7JSXXH46VuDoim6yZE+B74wVDGLM
yVWEXoTiCT8DVgdSVDhDcU7zOiwZAF/4BH1mlzUAjpGIAx1LESyWtixg0Hp/GaHHHjCt6rcGJbKW
T3Y5skPG6REFE8CUGwoSAAAW4Ll3pvQqNqyv0qNSwDYIXbXfJjWSAQJqO3topado/a6PUiaS5tzU
x55kQRzNyDBh3vQ6EirbjHpXSRSMjVekdh9FLW2Xcq1RHokflV9h7hm5DeEkcUaKtGNMA+qsxzW4
oK4Jqh3CEZJ/g0PZdJyCCPVMDvgP1w1EStdhdWVj32Ta9nc6iu4u8O2px10a64w9PDcHsZb+hY8J
2h9t8ixTdvVeIUtMSv3qhEc0NtrHGUd+Sk8KdbrlAQswEqycSgX1TY0p9fjgJzZ2+e4ZDTVoHaJQ
kYwt8ixHi77LHb4pBhi6KWXwdhRQRtSbqlfFhUuwzS5GjI92o7Vrbys2bVQwfS6+7pfWK2ltzyk0
v7aD+eqs7P0nzuAsmQjl9bw0hmXGF32mMfXDXmua+MczpUOaLF+9PkvSjg9TWu/HFnfpuzJadWzK
+U87XfiNpil396UK2cAH26qGDyHJh/4axmp5/q6n1kK5rcths2zPODajNqo2ewYUjgP/2uov+61t
OJBhQkIvaLA2a8tEI6gepVwh6rNtxNY6Az8NCFw77IuBmRoUmWVGwY4asOfyj3qd5ABwm0wZeti8
yACM3lhIP+2IBYMA1KqYssw4Xhxm4OsFzeoXeBEqiGYTGELJD9b8XQOkbcNComOIDRA8iQiyNHX9
Il06gtnQ+UPeq88NIqIsFKSXKm8+LAoMhrCwvMV1GQcLEWkSRbDkvxWH1zh6t4tbS+6W4BibAh4P
bdYM3vnPulBhBeD7E/Oq8ITqPu4PDfnflG4LVmil7FIO1eVtK/zvqls/xwyB7cYyBGWj5TRItfL0
d7xhIocs7TcmfpuCHd4/3qpQ7FuPAKMdbCtOdNI7AjQNvCUvINYP6Z260Fim7gtwml7iXjy+AbuD
fBWfzNIlkjuc514X7UO0e+G8+nq7i+kE8wx+hznJZORD5IOJi7ECjd6tmqcAjcISm6Weo52oEAim
eK2NN74an2Z+8yFGblNbyYvTXh0fgw9SeWZEei7AbeD/Yddw7R1IKgOWCNoCnu39eGaterUmX2GQ
VBMJ293eMYE4dBIQtNZQjOeezJqYAmIiOSlLbn4dV1+Zb5mb9EE0EgNaaYsm1eKv3qVgRehtoYMf
OQ5FUsZN0w4UWJZ8c5rv/T8sIYAXowAuaymzcAXranQ6l+6CsMsg2aTDwXfDdcAfsBavL59Cd290
9DvUBcF89YmGc9j/LnvINnN8hjO30r2UzJE3+OpHuUCgBg1AmcnzgPjfEvQUUG76DrozVXCN63HD
xpeV2oxOPMuHv9H9GRgGS4lOeF1Ch5F2Z07EsNnSzQ5AYydNlZUP/u/uckshNeM/AuJZEiMG8MlL
hxvTnezkg/ERAxffx8UAsJgwsvaEIRafSGA9tp1eMIrKEuqFVR1OpOQT8svC6hN2rfALHXJxwMSF
BMN+AR12JfOqySsfvxjQaT/UlabPdCAKOU7OYefy4zjL9CSLnCm6OxekiyG0Xv+SI1H8oZdoyDsW
AgJB77VudES7CqaFlcJ1Wk/kwvdfCS84/phDI9lDeD0nrm1GNxhcLjKpm/1P4ducKW7Qv/VF3dBw
7WPKvHE67MDHe18LJUyb5QAj/ZSzS7OSpIfnMjBt7Jbtaei/E2Y5wmyxdeiBTQHQlIb8ZlTtwwEf
aqpqJZSfstV1FoV/tQZGr24i39Tz+Fn+VdPK8kW32nQIeVqMfKe1TDODUrzIrjyPKsaK7rrW9Tu2
peLCzi75WSAHHZPoweL/iYcHXUoeI0HHlm9AX/p863hEbCWpWSbpbnp1IUlt4CP6kOVI5popwqhq
qoT4wTMRPPcqxxkLbPv91FN78Lm5aLtU2KDIiLcIP369BuMZFtL1CN3eiBM0JMg3EAE35/C8xaFN
uQWn7IiARoYQVp9dFRLm61w2dTqXFH2uD2Ep13kE7i0IkPURTxdPB84hQgJR2JzlCFgRIbBHzhXL
9uzK3QsDDiXyzdINq2Kxb3ZQZjPHcwoXXm59P0kIXHlnHWdyM/+pXRltrD9EgvspJHVGwnOS33pq
PQTWHifoqCaCg6EHK/G/DXQcG5plz9Dnyp5gj9oHa6pr6JuCu28LTdwba6gvqedQbgNxCCOiuyBl
YbGU/BGBnXWDR3wOkdPb0ZyCwI3MDvrC6vupxQaSI2FV/7Pxlko9OpYsCAsOcth7J5Gmd0hftEmJ
F1TyhfpRNOvKAT+PA6DTyGJi4/JCQt5+sspUUBbKLgOhyQGZCy2NH0bKrBfUqTyBViaihN8J+JIb
vZHVoLYu1LtBtQXqNO0U7FBf686BE9ejf1nFlO9N0dcVVyukkZICLc1PglzbwgsiBTQTtDbMp68/
cDLQb+xob71OzPmRCdUIZUt3cvT2WNCFZagoNKEi1IXy34NGfL51ox77+UpuIAOH84JC+f17OM7b
wa+5yQfXDNWSjxnWDYmXj+vSZ00NQTYSWH0raVsuqYOrjKKmIcttHlrBFQTknXWXthYWoLrB+KST
D0+pfVly6epV1dOtijwkLnxEytjxxq6JxjE5iW8fhWr8RpUZuhAfLmMycHGnJcCPes0KHBB0RyvN
778Un2S2OkL0mp0Z7o5IBLdHNPZ7wwwSRWQpUGTElzU7qrYF7rb+5oEC2yt1RPdKClG7YikQo8RK
U5L0xm5hjRgJrUpCNIwlFKNiIXetOlAT2YgOlx0iDnCCboWJw+koQVQPhmBFHKQfC9LtoXDftUc5
ALe/HyppehfwiiqMm9U3bvCP1Fq12SA9tJgYYPFgoNW/r1lfZhDlmoabPvLoPNJEFFo+qJeYxTCO
Bd2fz1/GkLnT7Q8zCu9UK3Cwt2vuxAOP/j8O4k+QDYginFP+UIKh9NkC5O3kpCNKRrqrskFPt/gG
/uMpMcyRpxCacKE1frBnHZQgdj1OJgHGA2HEIlOhneYkkJcXocG85+ryfAkM47lTcgpz7qJ31oEX
nWBya9wyYN4jyrmGEgKMwfwgE3C9A6Pa9YngSUSHqLoYz9hJ6G+ZPAX9MGb4TxTfyxZ49i6sOiIP
pw2RvFqw0BKg+5QHPKFgp0+0v4uyBiGKVuSuVEN7jG/yoEuzl2WOryNRsXC/V5eHZ+E7DHbgNA7g
1ZmxXTwILmG4CmDSiwfsvDX2g561EfTPVikc3FXEu5cjG3mp3x8DvwIQTg5v1ha6CRKwd0qL0jUz
bmX2ftMmEJo6ACOnO24vCYTHqivwdM5qq90tqmi6mQD2hlUxjW8v8i7pV1oW9pNWwErzwf2B0hAi
Kz0M8D80RSaK9jtGsgcTTmcyRPrBeY06Wa+E6nSFt/x7Ccn3diWJre5jgXSNqnwv3/MHg3kS2NT6
eilTTwooPpmVL3ypSkzMi7hddsuOhLZZrVGyw2/sU2mZbIlnHR8zLOPNG5dks8h5GeVhHtiJX4An
9SABPn6O64FGEt8RGTt0gPYs9wmYuYuBh7+tgKzVabzSbXisAgiI6Q2vaVMIrUBL9vu6DdsIaVU4
12I5e6JjQ99h5Qdw3bZri5Qp56NL49Pj1vxyejbVMKuOLqIAXGQhojWHfRH8MI24fSE4Glg2woJv
yDKo62Hd4By7zUpff8my6vJRWLrPRsnZdn2HMzOFLTo/gDF1uJeo4U2m0/oPFis22P2zvCndp2GK
FOqaSwjKQS7NHYEGaCn1oFiVEm5uGVb0r3Nq9RuCYrybagwryWbN215egAKpU5+t6Xo2XsQ4Dae+
8aWhDCBrlmfE9TI3wSudv2iiYCQWEvxsa6zW+bdpTeNLnPZD9WI+xv++2v66OhYbaTdA7jyRyU2u
hYU/SU1ujUBNlcy38o6bXbF3BHjYL5nBKvJALhVT0r+lP6A2ng5WAC3XcT3HQ4vHVp1bam31Z/Uv
eKIrFm+0oZX3TuXYuy28E6uGXDymtI0kPgOnTUPrtV02UNQ6ANCMZaTtZEAWqbRll/763WCKd0cU
ghfHF+rLtdEQbMYS0bNkVZPWTh8cZZBCfEy1RyVH/gYFR/wwO58pyyWvMlZEYZzZBU/i5iQAdE9s
qUYtwWRKttdTsJU0KZVaULM27Sh8GlPQTRjlpgSAVyCNEgD9dHwbqpXpfhW7uCgFvBi0VnGW3MUH
4lPV9IUduZxxAt2Do0EiWfH2SSzmsmnZ4T9dy31YGokgICql0LFF8C401yw2VZwxP5TOL73BHAWq
UDR6UOGx9LmZQzr/1UlAwyopTVKzl1YGigxjzFPJf+pnYwVUF7/cdgruPMC4iE0MqTMZyUkYXoDT
PBIygsBOtyd794ePvFuza1UyTvvJBqVp6RsSIg6bPUnti0IjMsMQrnF2sGdeIsX7SsMVvJtcd7Mc
Qcu5yT5dZGgoPmHGMIA2vXjlZUqzXVVr9x/LkjrdcAQmXQLHc2KCim+bOeLR9yTXesjZvvS8uMDQ
Qn+5u3QrKnFE/xUo/j19avB8PbH87d6QpC4SNuEpXEMC+DTJYpZF85Xgb58iLMwaXVNyxIx7mpKu
OfzeFUtphEgbcuv12R6ZG6tQ/HyuXYe5xO8aiPIT9LHdLmZU/E70UgV1Tu1T8NKpDegiEhUhV8++
cggGgUXXaKCDCvOpOxfX9fMagNs3oIT3GdOngFmXRXuRwWNZRBGafxZQ1fwLhBGdxbRStUbiPYpW
mcmC833U31T5oa3/Lptb1++IZUV8RHGC1mLwsYC+S4B7/gHuOr2MJdGV1MNDO8fW8EPnIHyNcCXJ
rzl0REWEudqs+iFQut+Iopz4zh+9hpljt9N2KyusFHFn3CDL04bB344/PFD5j2/7QAIpOArhTPN3
ULcXP2g19Xu1TfZDnGwaPc0A9YMdVmANkJz7DGCa88WR12GycKh+6/sCCtYLvEyp3V2IXUOuFCVY
KKseHZYaJ1D+UDV8rJa6FQhvNjf3Ai3mRVbNNyiq3E6Lrlmte6beVHulJdlX28aq0eMSuFu3hxOc
osoXIGb4aKHlgh69qjo+nYhToLaw7fTD/qoHJYBF+OJnIglRXLH82sxxGCet+Kb7/zML9bjKr0qG
NyaMSjZD1cHBT11uczqwfija4NXCb0Zc8nt/PjXVAIfz72w9g8RDLgNNPQmkLL7tBV5GjHqWuZ9f
K+uoRPhdmpKMyeEhuPThfAixvYOlZquwFEpenCn+Y3ZLq8NfpJCOGo+z6Bsmu9WXh5ZC1biwfloa
B4LUYr9a0LGCL2xMeGWJj7CDe2V4AXck4PXa5LvNj6Xz2FM51KWSOxgKnt3Fce75ajQvux+xal2j
AP1ALVl8hKOdnLXyJN5vCzWeaGj6JpG/liFNzHd+9S6oTqQvVAX4G40JXkuuMqG3vix9FM1bUr6i
LVZLcMN05vNycHDXcDhKNSEIWxIRhObtkK8Av5755LIKeLJIfiyTPMtY319huOC6II9sV+iK6JJw
qtZMhPXisdhmsUd1m+6iBx/K5vlh8PebPZnx7quFrFCG9juOB7LPokeB8hmBEX2MwkSPznPvXdYV
U+mhVaNciaEEUpwIwGEF2spAPCSF3m2nd+4iDsr4iAQ75iSvUjNZMJrYAQRaPNqwqfFOaHlo/Rmd
x3RofwG7Ie0WiFktnHfbpLaRLTLCF7VBPsbWpkuJDmJ5xmXbG56aPvmuPsTFyIwl2vqqGce66DPC
sLIHe04IgvLFcMWvCSrhqARN87XlkNis4aVRqnCUbcp1AVd5SgvWIVBgVGFn0udynP+DhsAvRfMC
hvq0b1i3F1aVJjreaXlcbNihTCqtgo4KcOZVo/W1/QYRrxloL5egRHLSrByg9yC8zvqs9EzMGjoo
iXGz0tituCCpgRSlmu1BcrX3wrr8LbKCiaRN0UzVyfkxwm1el19TmT7KMrTQLOCMbOdfJMkXyO/Z
5WAO2Co5MHzjbiYUhYmFBgHU97KIl/pYZkj1aN8+qyc7fpPi5kxRPA5sNreqq4qDNVQsKhaf1WF/
w7DREq3++85ZUTaHWg0WTG3fsrLeZKekWTHq8Cg/jOgTDo08bwpDvqy7moiHdBWxol/HpFYcb1/P
UjoG8TE3Yb9QG+Jvvr8Af8NA2Q2XSajqjg4CwaORS/dLikZ1Bnr+el/4o1bS1RF4Hw6FRoGlfP3V
vxuvg39LabH02/aY3f6WPI/8/JvVye0W2bQfJiRz/H0TEoLb1byhYSL9Lg182ar098lkwcSJtX8Z
MEqiO54AxoVSchkYBBZZfFjtO59zL+FND7uAzHTTQEEaDES6XAgd0aSUlEGcva9bUfaAOQjbkLoy
rAr5wPW/FF0jCYHKE7PWHw4MBRjftYxrDXh02t6O2LR33PlOgzTgz0Pt93WLz8ipfoHH8IKk1RGZ
pATjM4dtgYDhSb4gaxeCSQoBeigt7Jm67loqtLHZrqF07JTx+8yX3xBQ0Nii6ZXcouLiE3ikk6ee
qfJnVAs5VXKclcqdzvjK4GVNWmVKHodTRr7MPbsEar2KmcllFTrTNi3rtwT7EDtvk29bYFcls+YA
/IX6XiXnoR+RA8ZZeoMgCxGke6dpM8XfQwSVZKwAlWws/+5wX/GvgwVkPU8NKxJypluwhCV/EqeU
p+kATAvwiXXEBzxchM6Q0qn/u6WW1ocTJly7OIg+P4zhyBSPzTZkYqxjO8uGsGqQqZoesOtlqgNy
/3vIxpto4ysnMglWUaAi4sU+OeX7LL6YkzM55poSE2GqY3B0I3wQy58QfP+yfF/NTrGjw2KHJ+gH
ZP2zAa2uj0Zm/1aSQuAwqB5WEtzjamenY893zMo36JE8LGKqkS/FjJZf59Zw+jnjwM2YG7ST4lXt
pQfCoRnfA2IBMUK+XRsQckVbmyn1s0+92uRs3l3Njz0id9dVEM1ky0b5RlhvhZpMa7y+0yobNTIt
qWoQqhPB8u9oht05giBG8GAb4kLqYkKjkcak+zb6rbXBG0D7PYmq0m3kWVgDBaBcezIDOOvDUvvj
O2jwv2FSFkaeEcYXXD4KhnewqBjZ5BpsTSwvJVN2mBiVA2E3vj75MvKm8nwtCmU1cmwDxqAgheUE
NCtQE2+WZ76BdhQcjpEMlKRK+b0VY/cLIlhCL5qKHM2IPIrpQ+reu8V3By0IHR6wwWs9mSFz2kvz
fIjwzsRuQdXkeEn0QLOjF/GR2hG9LlpWRE+K0L9sq7NAGTKt1U0CH5TDlHoBkcervuqPhD/6puTE
s63NkqyY4gIdqatDn5oiBbt5fI3A7mmIRa5YQKZR+Hj5xfbIbUgZXze+MCZ/VSIn1GKzLETMiULl
0pBcOKxBCshRWv1S2vSsMN9Tij0F/70ccqq6Tk7YkhVbgvgcXmoBGXwmZsW65MCUo4hqCDOy/AaT
arK+Z6xMpqijGcmm0lSpSQvKfLlaQ1Utq5lB1wSKxATXPDQ9ZMH7MB4Xh0jeENCUjlnhwrixddlG
ze6rSP1N9ylzyTVInX2waCbs4rQks85c+VZOuWQggKIeVkqlGYznYW6bOeT12XA5BSvXniAkZKwc
bfahAKgu/GoZavYb7PVKIU8wb0jjinRfTg+6RX7uwiZLlchfUu6ylD9XkbdestgJFhotbvp053qt
w9b6fXxXIvWulXHfJvEhLX5Al6r42yQC8q7Aegv7apow2JJusb5rvMzXI10Znn2ks/iZtyaOmrKv
fxjsqOoFSdpCv5LM8fdpNQ66tQ4q2eJC3GBxUOpahLXBmlQhYoUB7FYXdhdKeM+F6twIL0eoy4Q8
oKEf2jTriHtxRGKTUxCK4sGBe5D43JONPQXU6T1LcvGkKu1+JxtAjKLaW4G1eM02lyHL0NMd7QM2
KgAWTX8otoQptkTqwX70r5XxgksSaZqh4SZs7DXItnNx5R0oRfsYl+3g2s2/nD1yaf7oDGOEn8p1
gi4BQkKmaMkyyDW8S1SU5C3j0QnpZzytH9PTgLRzZ4cTAgq7eUk2TJ1qazxwIsLSiikO8u5Y78yD
kX/oVK65eT/4WGAhXP47u1LKBToOYBpKqblAV4yd3UjNoOed3ykNzgeGoU4NYDW1pEftEHym4rdo
R0/LZS8qJ6pN3WCuVJl+3Xepe5lXZnsI8dO/plxa2/HtiyD5R2exI1QcWY02I2O5SAiNOJLNHcPQ
lA3RJNVEHyRMjViUJTK72ZpeQ/xbQRlV5wCKCF9TVZQ+ZOHIC2uTCnRc7qJgJNGlBAYM3xgL1LE+
71h79HaiR/BRFWCR30M79BPlFvKYOz6yz9Dhk1w9g3HW1sc6o2aom+IRtJxtvsJsvbC9T+pUkH95
Vd2j9it9wW4lSNMBvKFUaI/T50hqGhZtlFwsF2f4WQKk/2d0f2Q3rNRzz0AKq6aBmdbcxyIjRPlV
DaC87QKqlZQnnkWJux/tf59r+QaQfwbIkrDkvcc6Jhv+ZfII6EC6Pd630IjQCr2m68+mKd5yOKK1
aVxWStHvtk65V+/alY6p3jerJBedKs708QQvtfiPdgsLjvDshMvb5vmUWOcg4tOuxv1FVtRbulkg
S9IkNh51Cs96NjIg4aU1du2jOZRutVhi6dme4KbQ3XjFkLJRz73n+1kfCGCq6rAYATRvON4Er+cH
PQOe4KDKor/VNERFfqmAwhduDOVaX0zOAs0uKyVQ599qBpMRrfWE8tUxtExAsKgpP2n59+I1UbhB
SVWUbVVy974weE4rhjOFFv4zGrfyaq6eoMA0hiW5niFl5nlns7tm1oh3ySzTa303OkYlrFYFnGTb
rs6lXnuqtOmRmSeUXQuWNm3oMY2joU5ePzK3NWZdeIC+TXAJoCGQKT8jTaTYoNDvViuiziqgmpiV
zTn6kEDwWGQsmQb65S8YDAEkqpEgaJvkaVB2QTsuBd7ugu91Gto3hfDT0EnF1c7cVxbXXH5Ci1B5
BHti3xkhOUM104ywJPOkk/ybBnRXMk2P5S+/JsDaOG2DlZ1/z4GeT40mfR61lsSonpSESBKArOgx
A1SBc7NkYAF6e8lEzgdYc6h6YvnsNl1ahUGsQeVZ5vPtdxz3Vbe74VbR8wG94wBCY2YtEnzOwOoB
DaJQR7/G1oxTVf9ldKv9ClHWHbkq5PXhLg9F2/NUUszBB5XFFq/03R8AE8N25jYlSBOIGq8vcSdh
Ybqkyq1YG5eDYVGzBGupKf6BOnCDPrTNhLZ8wmnBHGeZozVtRYMtNK5QGzbrDoA1z6A6q33T5MLZ
OK00IVXwqdZ2c9aW+37oN+hYd0uZpnZU0T8yS0y2r5bl+TsvTSru/GODIgiB6Q/AZs/+ETv1OxkN
CM7U+V6ptDiGMr016TjcvfsojOpJ00UB2GwT8kcS32cf+mGzLyalk5Zuz5Tj+XWo8FveslWt7xuo
ANVryIIrRIEudqVM2uaPVXIbJv5S41uyNj0w4WspzFTdZxx/COUIEnrSqgmxsDnvBU9t2qi9qsHf
KzDpjxai9L0yl7oyGbPec0LynJxB2THOG5oFBTj5PcLl7+Spb0ky44cDwN8jFWREfyVIY4+LF5El
UtRSF73p3tZhBWjxAWFxBXMQCnp9c9accp4smeEyHnzO1ZT6TE3TjCRNvr0CYrhXuXVMuxiyuC8B
PRrl0qp/+L6H1+xiR/fxYhSHmelZSeluBX8hqQQ+T1Lp5S8E0jJMadvnoKAt/QZDGN7RKq0vWBul
AOczX7Zmf61fMVTeAu77KXacozLcn0mujayMd5kd5diS10YFqsl1U+PTGGh+8N8h2It7t85KD9VJ
aNFLnRRGab8MPNpVqPji50azei9Bb3zakHLrsmcaxiXi1V6mpJDSMa6DsUKLRe49u754OTtWBZCi
wYPLUH6NSK+LIqekKGo5CQCiiVjzELD9INTswUM0deesjxBIbnCRJ5qy1FFIhQ7wQ94D1fo1q8YC
HsBN2ZKRQcjbWKyEOT8pI2BSO8+/Gw/9BKoCGi6dQgCVFE+At4lzF5HFIjeyJi4voddDk3m+Qygf
/geUFxBpyISBORLsqTwnD6O41nF1WAlNg1ib3tmEDsoSo1MxwftbrRYF+sLsNdD9Jf9aDLbjTn39
PWGENljTChdCX5c0k0azfvNevMSFN/ynrYXgntZXo3oeHTrMYOzY/hEitA6Fq2i9v9kYyVieCdEU
kHb2ZX6SxcACn19e2FDwhuRbortyhvVC2n4zdRtCKoUH6h9lFVuY43m8qVojAC7QFL43oad5Y97U
bsGbsexMjA+CzVJxkTc/5BAgq8yrELXAo6jBgzIyzqCVQWa4USXb13hN0FI8iC0me/fCXRspoFRL
lnEE+HF1P0gCUTMjH5k+NZ/586SB35i+z5qb3v6R/HYN15BYH16gW+Wrv450Rgk1vW9E/vTgOjH1
xwR9OP205DHvvUWbUxVKIHRpjBnDaxSP7lheVXR+bKmwIfLYKGLLfdoACtU+Wq+Td4UXyZD2nO0W
Yh8V0w3BZeVDagEbI4daugOxRJt/eHpaJ1lN7n1xsEgiLA0H4V5HVZl924WDXL0zNHdZ1ucgX3Sf
lyrpEMKt+zJgSMtixkduI1lVI1UCkyrBC2vYdx+7aWD2Qw8yeo0H7CllIGXq5OQf7zEhb5UI4Dbn
jXMl2gdgwuNZs35QiRP1EMJvxN9z1e2yXXnEUHRpImyLzO5iXqfoJfTlWb29Qt6CJujMplon2gm7
BEvE9NIhzKmaWOvwo8q7Z4y1vU+QPD2J26lHk1RHgia+m4PoGvc0B+lGPRA6vNpcinQBrFM3TfQ4
erLqcKsgNp9u50/Gi+deA//H5N9yfoNYu3Lkkxw3xTFdWZmy0YRymgxiPF4NEMOEtILXyQ0kKIDN
NamVeHwbf9C9mF790A4f0XaPeMTJeO02yxBHm331eMyFQ+AyYyk6O19hG81N8T2eu9erX8rn6HNO
nhQNrcGb2pYwZ/1pHEzkolni9le2PWkCon1lpS+vstO1ToIRYf7ZObpD2SmjJhfsyutFfpLP85ZA
ZbtYGR3jUtU4ja6gCIU5US1F4kAXgohaB8Y61x/PMtPd0AIv/cjT7+i1TK3wyQ0KZd8R/osl1g/O
TDp3qmY1x6a59ylfZexw1Oo9FkYlpFPwcah8dLTWMJsPEUQmJHQJrFBs7oXZpg8JuvnxI2S7sGLY
CQKpoj1TmBlztZW9KwOmuQ6j8TSQwSxcEsUc61HgQ+8kt9bHXfJkDSQyrzZJqZ3iC6ezL0njK15N
sPi44qiXt1+9IXj0j2pj6fo33uldb2YnUb3S7Mic/UJzqvkeDfIACtvf3joNOzEYAkGNlcXTJ6+f
9h9gJC3Lg9o/tdD1Px+3jR0V5LJjDEMtQadk+kpr2rUc9+AqfHqyVwsWxYvn9D0sf1xbghGi/oy9
rtjMiDmxoRpSUoPJIE8Id+7pGkutGnbJz4GRnj4/ABDFEcBD9iriUCTVIRIfW3u2NaVTYolFbZXt
kv0/GYiB8BuIgK9T78Pnq4vThM8luU4Ub4hFnJmzcZ9jRMx04+rpXwjV/RiBxNhCIetmtSRF5KtK
KKnwxNVTkIJk9i5i+m9Vja+DHEe7heO3sOL0P6kEsKoY3ksZQD+509fPyHVb+wEVJuQPXZzYGTkr
2oARIvgy3/Ayk+3obG+hcAFpiE6cM0cI4vFm3eucgsCxtQZM78VTz6mn0+s9fHROOTAbvo2bL4FZ
bjIu//Czwi+eng+5ma8D4OO3pZvM0I2ov54qh2jeNHXyFPCIryp9L7uLFKvc7qy5Xcdnj4TEO7mM
B8gzU4GFKCpxLqbBi/RXeKbIeRjjHnexZMl2agdcDs+NYUFhipNEew/oXqED05aSQ19ww6UIoxfb
pd3TS+SyWtFW9W5ylcs4sHwitTjINjj3NcgNzFYZLg16aioqgfidHWboBKcv8psXldypN27Twk/4
ZVWHgMUmTzY+LUfkCu/ADizPxtvqNqwoOBwZpyW/+VmQlTdTbF7UF5qydaivf4qpgySFdFP0D5rF
4jj9ev8Ct4UDXBqXljY2TJX3b1QDDl/AMGomrBswNiQ0JttQsWGqYKsokepB4wgiyrXqr/dAt8OU
01LS7iaKWbQeZNCsy1/22CCwmH/9Cnt92oPAG8WBxHnEI26ybWh3c5LgdIiPxdL8a8q4uX+H22bh
HbhTPOEq4kvdDuwJHUmMAc0IlT6gSJDJ3YjEmxYXk3HBTgRiaRQVgghkxW0up8QFa/WEarXjchDi
oqVNhpUIZOtUG1ItCXMdj9TjYLxNH0NCSPsTcRv5jj1hITzETTESdMS3NIQeLV1zyHxRYFfd+gCq
PgiNuIdKpOa6yveWpHPN034NbF42ePXhSe0b72QLTAFtnYwo6r7h2lAlHz3MS9ZpWKYlMpB/LKv4
RhLDsOqhuKf8YRU3Db7RAoWVQoNPxtum4jA3oLG/L4VHyuoASrnCbKB3suP/n9zqZZU/zRFlC/hv
Tjsg3qWX+YmXPv92MNu49Qv7AalAqkKjNjRh+sVjlQqqh5HTEgd/alC3ye0CNF6smBstjB6lv7/J
C/xEvXTVf0M/kPsG/ecpYBpY6Pn/sdoq77l/MfU9OVQmZj0T5bsurCud128T/5zlTGuEO02AKajF
r+7zCGkjGhbgJc3hIetynTHn9DZHKCKNCsX6xlHlrPJQ4lRDV1xmExxkg94ZDV805cTOaix9xNQX
j5eqELswSihUpwOF5kn+cEs9XgIRKPS7OQgfboxj1zmPNXdJDLhN1WNiY9S1YBgk9437EgAxr8aU
goIWTRKyuIdFtB3VrCyGdb0yPUtnDIwdk7qIHM/MjaDmOAy8i7LElsPuw/uiR8OjBDh5Ku3YFrJD
ySct9QfunGIDX/QNQckMh7mqeJZCVLFO5wVWmV44ERAEie/SeRTbk7Vrz3uYspJvmqvyTH5TmK0F
aQ0ObisZUSGD1oM1iKOhRwEtFyMl/G6myu6uaDfOn2jEtKkH7UyfPHKPxEM9Wnt549S0AyCIEVqB
Esd93ZDyfnn+llzT0NC8dZNa+bv9/GIdAGfhuQJCSXCvI1RCaWaa0L8iJhe31b/kJeKXuxTFDBBq
T2JzrS5GeFf6FB7k46GpKJL6FXV+tjpQ306JjlbP8jVeuVWinuzSqYLpmYXbk/FfMVNZKLC6U/9N
hTMonNmAbwqnFp9xk5oTFLqBG8K3PnNrWA6Ds+bGnc9virdmjZGQCzxbcWZ1Y7yfc/Q2abXMGd/9
f1TjT26ppFtIZjtktyl1Qdf4HGgL546mbXEVWfZKKZqSQUmfpBOZjy3XfohbicjAYn3P7mm3JVhO
4LZIrByLj9rkBZ281Fy9J9WCO8GEg6kBKiuya3VLdG3c70axJmzbS4xpQpwkART9MSRsOTv4Lckz
ITeK+WdQ6EJkOf95KNn4xhBN0g0Voz68hMa+q0RfkzZVsQ/3EO9pvBOKLPKMbMYzqce0aV5MZIiZ
cT96SABKa2ySL7xWttkvUNxB7RqtmWhOBNyLHPA2FjyDi38K5LmLEOXXI5Fe/W4SryZ0TAbq9z7v
qeK94UCbH2+8jQJQb6ljFUxORyTYNNQZQR+xoDdTSORgjVJrgjGEc46D0FhRiwceRJa0T0bMu0to
dFZ4DMtEeAIvysDccvvruwX/9tqRUnZkUV1rIhkaF/Phz9jGYSx5lfBwpQVIaHddBUwJyPY6O64P
aTVjO/6WfjgoeQI0vrsZ28sVh8uWfkojfzGj0n/N6QVK9XiaXu3YydsE1WX8se60WLBPo4P7Jra6
54JAze+Nkhym8r7eDbNv6tK2XMSiiylu+K1boaEKk4kNStZDHI/0w5v91E4kBO48OMWDNoZxRgtn
AU4wrH1bCG7Y68+aQjrBIjnfruuO42zvAMe5aNAkYgcfhZdrikwzxohJjWIHjeUUDXisyhNftaH6
7BH7ptCcqMbaf7aXK4mYICWwpNBpkOVhJ5yu0MNL4Vk/qqDHIxeDMY1h6bvyjmLPS40w1tnccnrt
VNx8yZ8w6eRHYD3dgwjGEYYTgsjDpRmSpYfVLMCdrjRif7uIRjaXzRzMY30OnOwUCkCDdctSAVOy
lftPpJd0kEgylXe2c0rW813kwyWC1+WeK84FxL+wW6iXDYltMS1OGFR98cstyPAKW4yV8RUEBv62
Q64xdifBdr7CRM7vMhPIpiqpruXOSe2ycKPzVXQzliovSem9IoBcIb+yoHKcDIXekiq6KHRv4q2M
Bb40szCXeZOSNKEvJVJA7UO5iEl6tJ8bwDFzDn8WJa1HaFe1tHGT4wA2PTCR5BPFFwMHKWfdfMtG
aPJLs8ErRxHpmqIN3gGSBOpIEJx63V14PcBm3MZznPoLRNltY2uwbEi/W6papSmpoNq9aXhxspbr
AwjzyPhSoA/jfx+F8qsPgfzejHg1mRZfJzpQJgd5FjRVOw3cIHQJPWE/cJd7qqoXT3lJg+gcEDPg
WTSAMGDake/+DsFKIoBfl9cPeqOLoDGcPz0QKAaTJxUiWdfC6xm5vKyKLfoNTtNFGkMUQiPRIscP
QR/+AzUjooCx2fnQQdUzMpkGV17V/kpwKAwsYxvws8hRE9t3hF3GiFB91pNl2QuOd+M/rX+3q4Zp
6v7pZvm+Lv7tzfo+vyjBaY6LlUSaIa5vevEipXgjwAfM+JlsUIz64aR0iurMoUeF3KmXkU+cPMvF
NyZ242DdzSgWBxgHtqP4I6N/zm+HI8Wz/WKSrHO9EnJyzppbZf3m5/O97HIouMKnaWhPbHjhr9Lf
FHzsI0hpmLP3ejgCSH176feQo9w1a1LErHOR1T/Pia4X9VOFHC3s9m8wPVkPmKLeCN0lf/ReAJPr
qskc68GNJp1SmGpnRsvLA+Sp5nxy/OpQiIVK0X5HTvFTupvf2k8ui2WuouITYD9a8gcqibngGtxU
29DkFE/isByoyIfXNmYOtmbnlTrDvx/geUgNL9Dt2JojbTCkOTgR0BTngZmyxCHQICr/VP8I6jjB
n3p7u9GR6peA1o0QulJ4KL0dThpM7sS1xCcSyl5XYZUsub3ftz/qkJ/eo9WioKPV919zZaLawUZz
nAVTi9KkHMWaxfT+1qVMDHjBjI9sVKC4GoLE8hXsiz9Q5HESSw5i/gtYzE98vtV4zYWazAXxuJE/
J9GBbFp0+PvMy0JSwDKePsb6M2avf0BQi66Ec+pWmXqXo9lK31ipl4sTihdVRfOsMLmQMqIV249w
vnJdOjvhMEUsVaqsqnHVwLaf0gHJd3xQcZVdp19KcukEqy02ok3KyJd+uXr/oE7lIZ/ekC4H98HB
u8akuLB358wi7bh800CZpKNtePbZMD5BZyxJxqrwSjyHQBubWq0fF2onT3OQk3AGXi4+hflD4SX4
kl5D3JkZI8xyV7V/GHI/y2dvh6M9N91eGf4aPTIcdq4kSfr0zXy1PzUdpwZn2YyY9JI6ZslWSKQy
28RwCEywOn37QMSnuv5TDSnds6xEOZc89jKVrwJcNnzKqxi40NQHAe6uFVEA9CQlqlnNEO6hhvBu
HEpAKjWsa7QZd4lvQor8uXVxmHQo0FDiVJorB9UfeVw/C5Ec2DHRY/a2GRMukYIxZjSsVsqUxMLc
IjLMJFLsAkitRm/ygM/MeLmAxoBwcMAigAghS4wRbNf+djm6RzAzkfj8EEY7n0RH1HmcukO4eZb/
oUrQHQSi7excbaNN5LrZX0j+PvkddZFBbGPhebUQg/xC3yJyZ+Rxy1VHCoYG+R2aUjujjL62qztl
0C6KgBUWcZPdr8Jptou/fU3RzJARMDaMauKjVa9oalsgiAcgc3NO4SX0OzAPu2X8mdiQ7wC4J+vb
6BYUcOMsafYaLH0eZ3LBp5yGY5P4XIB5EXZP0GM1Suoe4zI0+q93YqsRutceZ8ZRuXKz8pfIyQST
QMrjg0608GsApphAO9b50sFC+GMcypivbeAAS5R8brjQLmUtTY4t4kIqjrg2qiN6rNOtXRnV41EW
P2MZ8cvkboYHZQqa2vNP6yfZNCUvFVO4SYK9bHtajvoV5l0UdNL3OwLaPe1NnmliVS2LrDKjTWrM
HnKVOEKlYlg6Fio9i9nVPVeFYLX2ZmWuZ6Knlk4Xc0J9ms4Ww824Pn9S4lq3MynoglJquXGmI01N
OqxwyjXIwR6ZR4aEyhtAbgxycjam3oto01QI2XrZcOnLUlL4uDdvlVw4ToiE102c8dDv7g2LjWQW
+5JxaWc3Pkal0Uv8QXGFFUpmawVId53JITp1FDXaWnlH2EucBg/+gzSB8oXQjFCjUiplUqeks3XL
5hbL1PoC6to9G5N4InJ618UJVGiSq9t03xqWand1f6qAsssQAi8o1GcDfzbpKAXYqm0AbxgVA1r1
raTp5QBPMRojorJNsjpsSzzq6/LQlZlpk4etp7mlhk+glhT/7j3QP3dji2SWvkFt7klNM/mANc9o
HWGUfxUSHS6USzdj+XBhIaShY7pVymBDBG0EKd0seiD/t+fwUIlt2aQ0IoRrb6TrgasEfKJH3C8x
Z8Co24rD0gRrLlIiBWz/zpL/XsqW4hwz1HCAJll4EdmQeCB4FJxMyl2UlxSpCaOKtcwGB1+6gMZU
f43IMqpY37Ywpg/AjZzz7J/d0zv0C7FnpGW/Xb84U5LLD7Py2OxTw57OUc9L3YUMrj1iaonWIRXh
fIVS3/gUGpY56GjrAmotByacB2Os5JSGLh69vBRO/UuTiKIp97Zyib+0SwEgyWAAXzB044LElbu3
9ydXdkfIc1Qu2sGu4N7axV05b9rHTXc/83kmX9x1kr1HtsuyW22NzLBJKE6/DCJ+8nX0qSPOfvm8
r/ibzucD08M3W5aP9KuBfFWzSeBoG2CTilOH0j01OXFH0uE3KeLWxk0VMxUpAoSZE3nnkNOgNOcl
kC51EDAnfJ/EwDGaG7uzLZFOTuI9kzPq27j+QbYvnxvVT56Jr2CpGKieLDVTHaRmTLU7LAOHL8H0
huB7zxcyaJha+FeHfxNUSE5VjSB2PspW/LHr5F17L0yaF8ARwWLLCffAJAu4XqQF2B3RcCo4sf5F
h9Fiq1Qd4u/6/3LOXEJ2j9So3Akz1w8Er/rHe4BM4TcrhuGBpU7SPGYZPMsvw6eHybNSb8CYLcoi
Bux5dwc3UK381KHwDhRNW/WWTxp4QF2SVahXzqCUc5nQnPmGE1hXKSKVfzH4Cx6fNn3enXZ+Ln8a
mXM3LHH3kC7wQUoq3+j9q0Pzkq8kPpwqmLCfPpyLwoau3Yd8CivTI1Es2Eitr4II1kZwGPwhJNIr
HR8s9FUYOrPfJB1uM7CDuZz1bSamDPouEMD5+pIXm5NBXsD9kJb8bEwvM9pSvfJWL7rkTIhHnMS7
vsxYGOGC5K5mM1ntOEFzHg2ryomPl0ym1qBdoyeHCHLS2noWwCu1LMujZWA/DBGKWorHMpz9aMQW
YeazRTZD0YHqrhhrzCrEbASqsMQDqQPhU4JkX/Fl4cdwCWNcDijZyNZKi7CrPh83ca4H/QDDQZlI
x+FnZBpX/aoE6hfvq3aYtu7S2vHnr+qqbImzKEC5RSQq793NcJaNgYhWgrAq92p86jihFylqn8xl
46CJTZ+/NQtDBi/ivNd9e3D0YkGDVSkJ3vkfKg6BTQvVTGwLxjMXi64YaUxufLb0ZolQAzNnjRHP
Qg3OJtMjyd4XGcj7PjEdvnl92x/KBG2NwKWrGhONitK9BmDOk/66hT4TURFYk2KnwiqgdiLye/9N
GX25yegSSGGEDFa8we5KkCrYKqHixA+EH8hhTtIh9CU4t4b1dBngZvBsuSAirClKC8DZsFKxXu2X
BtaFLsCwk2wKlJugCF4t7OHkGukpltWAX5ikz3UtsqsAdC8KAUGqONx/EzbFkctYOfiKHW3ELTry
QOiYsDYYh3gGfCiXr6+hcR9PBsgeuP2vihbkUWmy0cEs1xcJIm3ZLjdjiu0/5iYXtQP1UUk7IOvW
0tglUGADj+YJvfqeMWcVCuTjLPA8xjqOeswtg84RVyj20Ia/ebMzX3gW0zJIp78GuSswQCOe4vyO
6Un3XLIZlANcWky4VWyFhEeTSVptgddd4WWiBXlUSZ9vKKxc96EIkrpoeREZHOLgdQJLtIRJnH2s
yqJQGJlP3RqN+adrAdlFJ+H7FYgwU6gkx+AIHjGs2w2KSbjTzNl1iIbPMw0MHf1Eu5qjwXK8GB9b
oSSqnkzfRIZ0BOSy/+qc8AhWsIQV8RYJ8MWJXs01lduq68qrLaf+sivPaq6TSxTF6RoyToRD20kk
oFvRaR5LzLyQ4RRxZfiEZFwdkPBSJI4aIcxibQLUnhV2XOFWSouxHE18BxIaawuPl9UwQcXnp+cu
s6UJmxsfPZbTaNUISZ2t4lULygg/qk4OJZsY/piXjbWrpnRgFYRwbAW+d6Dj2wND1vzHTnhxL6F7
Z2BZIDfUesdxAZNo5OBw92H45ImnjKbI/S9qBsm39lfKiTqTyZM53FZNskjJeN1bwCBh6VXeGfV5
097quZiQcLXHk9y1L5I1NUaWPq4l0Xpr6xXSoa+brYngsUDvTrLKNRHeOFCN4GjGxWOqi6GrLKLR
MBxQRCQ4bkYUKP92BSUTaf05WiUEmPepP4pbZD5VnIQODYk2J/DpScrjdxMPEh0ggOrIbIlgYlLO
o+Fq+0ee4pIKClX1h4azTb+MsSVU+Y2yhG9auXDXbwhue1lORRE+rNKbSszQVRc4g6x9L09JcXsr
/M3dO5PJnXYBe3P0bmyvSdjDZa+LpatS5up45O3dAOdzn0ZD+I/FTLp+HjIP8bh6RvuDSHrEBHGV
maXacQLb0QQpndwv2/akP5+WA+Zf+2lRXnj0h618lscUNY3E4Oq7laBxWxJjcrakYJ4FFhZ4ri1X
lHkR+MO0shs341OajEHYvf8zZwnx2vRRoxN2txbOnN8VR3OOWPGLQUjc41oqt4s5qxPV7b4X8Dyt
KvCeqRXiOED747kAKA3xDK+NozNf8osSZDQ86pvHnl48hbCVmj/b3SUATj2YT00pLZtWXg4DxOCL
33J6WcHkvayf8CFaKtW/JP49DbiQEU8oJRBDBoP4U1hly2DDNRkCmBNJOmdBh2YO7wEIZ876OGX1
GawbdMOxb90TKGDN1pVeDLO9Bx0IiZXDW3g4HDoo3Qfjjtuoe7emvX8qXp4SU+vn3A/BL3fGYXwj
VbF9AH0GYuISnwJDOHi3nVNJtqFUeTtssrZBzjiQcjRrpRybuJfNNgWPZic77VjQSAvQOSMYe9vC
/CUQZkxsHA7fA7GXIdgTrzNd5tfotdX5O+ldJM9BUnD8zre+2ffVDGGtnoC7J+L2jqF0P9iFD/M/
PgFVHRB2tpe6pa3m7KeVvgytO9NPQTt/AKvccWQDj5zRW81xIK/DkXVQD0DyDExvHQW6FN1G67NM
JhZ3BiwmoOgvx3btnZ4pcFhr0k5VTLUQ06kjRRkkqU7d3tgwoYrWgwVik8OFf/zVbpx7alpQgw39
Xxhox15q9zvm7K2FPRgbr9qMPZUG6RUoWirBTG7yf77046eDGuOrnqIw0Iy7KU/9xbTM71YQRttO
ZYM94oayxGBceQ8bPIAFCXlNXeuonGmLfnCGXU5QdLKbJB4AnyFRVma+CKRTIXRXW8YoFquz7fBB
QASK8cmwzRZbM+foVM/nMV3rPaPUPseJlCVE3c7RL+aRCCr2iiHh2qc0LggOlzXe99MdiAtaGpAE
O9nrMif7HRT4I1wifz77xIUHbHWtRRnAjAJ+9ZfD9oXMw7EGKLDWYTVlkVe7b5CS44/gYYbmoEBH
3UsNOtL1qh0LEF4n7gN2wL7vVvDbBen+heHMnrQ9J5ZemguH1sWJrj547as6ajM/LPQXmpcL299b
5X+0uxEsyJ9u9V+FUboaXXyB6q2YKd7XmUIykH5GRlEhvBQgTxgt5wI7QXSqDkPq4Eulsbn/LQaO
XN5rmvHxw2URN1CIB2KUqYit3kHu4VobHddWxAjPGAtXUMtGRhFRta6VPO1FUFJvbOnctf8URXVq
gL1mM+9JVpfcFmdCNMQmnM7Rc7CKO3Ck2y7EzS3SeQrtlEs0oxysCD8NFDUgHGsMXZO27i5/lD7L
Cd2h98TdMy6/JE+KHTPmBWT18JMj6KEZ0U6Brmo7pkwn2mmyqXGzAiPgZ4Y3P+R1+Piz283V6Yg9
HiF2wv9ND6SO6mMHszApE6aPrpCQ/wxayeGL0Q3YbCrL01pQXxNm3UyOQLf00YRC4dY3lMXXq7sn
oUbdTdrZCxDMQn/l0g5ALm1nCk7gqi9Jk/3jQyxPIg/kbkSV0rJc8H45kI7YZwTqLbtp/7cCiq5K
TyhmnMjRS9rOCzS0cjyhdprVhTR7FFIybul0np7Jvlx59L1LJxiMNUx2Ou1GyqRw3zSSGdDAB2V1
HhNq8ENV+DzfxRM+Huo1u/PAQ1raWlSPkrkJvuB8R89H0Xa7fzSS1fraDkPhZ0sXPPcDp+xm1zpd
6s1IJYzZbiv2WrretZogpUzltjUsXeyCuFJuDPcB2L/4QyKXckVuol6ANNpJwUm6bna2UaEcwOX4
68uGhKcGgqVLdQjPD6tQKvbjjgJNFcvB+4Pn2TSf8mhtHkNdDVjrFE+Qdq1eO+7e2ACDUfi3JeSN
Ofqm+4WJoyDUQQcth8Heo8R60eAGzLMxFgHeROJPRkGlX0fe2tgK6OszlEYfwDLnwhgUw/yFN/MR
ZLoB+GrZ3cHuRY2X3ZyvBqhXxhYvTgHiI0qWrkJy9jQwesDWKiZIdCRPTVBy/05lSkQfPFL9zQEj
0PNWJgHLH4hh7zcl4Ud5/9T5BrFMHB3/qiSMyO+DkY8cbrixgt61Qmg2hn4Y7cydA1lRbmFF41xt
AQ1LZ+P5dRz2SeRU1+CSzTFBU1HIU/rX/8nGeBhPfOtzhpSlzEn9hfGfBssKnePVRypo+29JCfwp
ad8pv/araf2aZ9/cnnEaMkNaD7Gxjx0L4nhajUqkb9PFAdIowKmT7sD9bEEjx1Ayx7zum49C4Nbx
FLgbore+dHEQskwM1m20y7n0hjxbJoZFUn54YkNkJBAy4hRQaL++GnTvgvTCpzUdgr8MfH/h8wUh
YBSVY0BPKRL3+TnhqTIcXmZj9Zj7lkI2BJFj9cMIw/zeT6v+49EkOJviuUBPtiOFK6pPCBtlfcq0
M54kHjzjbF3IC7rlnJzigGcAicDUqwoZxJx+StIfomHJ96bxhghREUoJeYaShMciho3gy7UgVlid
3+njgOMwUrETOZnv2zuLRhXGYprLj3Wr9IFvpc2eb2+iW8/fJs2usNKMFeaXjbU5P8m478qIp9uz
5PDIrAABD7JW62T651DKp+24PyyRfs/2dKtqJOmWKGYrW/t4zrC6J20P9krA8WFUsDYURVJNtp1n
a+6uYL+nBWzu1spOdbqoUA/GNMUFVXvVXP6a9wrqpsFMT/isq8UiAK/0zxDRKYrijDC6l/yBZXA4
JfImIAck98TU+5ge4uuoH40cKTf/ADxFVw4Oi0e3Okw8tLxzwk07AlabDjWx+SQSeVUNQdj3vhxn
5nPvN3oqZWF7LFhHlwmcX69UH0ePIzxQCYTrRntapwPto7NBSDHO4TrPCvQEl18Nkbnyky+0DfQ/
bFMklvUi4tMzkZLnacZDoe0CB8PWS8jQhZIeMLljLQaTlDOdTonH+3Um7/jWa8rkIaUjn3I+OZrq
o3Ke9DiqaSIyn1h7ZItgt/GAncNjN/SMVihwY98ytGyCyOxwh7/ImxpZ3GHdzN47SoiYlI5xB8GL
Ol5rdLWhTGkMaujmxZIc0Q9zgvNNWxTcgSSpOj5oRimGTNuOh9ctw+XBT7h+gMmvA/4PesUa6Jbv
sUjb7wUVbu4XIuO7hgpFHEqJUh6e+pM7dWF0V+MuRtCCsF+qARpuk+qFE1q0Vkwaz6ryxmGrrFUH
J+X15BHtjFYM3lwINXl2/yATfoDgVwMyodl8OxmrcNl4NVUMy6ueNGyFECgk6occAY7cqH5EwiDx
EuYzZayhOHuMJVtDZJMrJuE/9UKcVEk48xisibqb15bbsNyzCxnnM3g6tywb/TVbs4F+SJpNqVh1
WdBYz13JwA42ZdlUnTRzwQoxkEgW9bStgYoITFTp4aXJMsp6ism/CUNursqT7G94SszFyAhJ0Ndi
QSMEBOSr3IPMJ9GyFcDd09XgiE1djPNEfeLSSTZxY50KAcrc0VhIPlEIVS+V+Dr6w7AnqQONs7iq
kxHtJ/zaOUuHjNYvrWnmJwsY1NeRa2R1GVP4n7jGRhMzQcq5coYtmEt2kW+hvggLF100MNzUjy5Q
JDKIQkliiP7RmVO7msJFtDd76erxUk485Tac42y8pe3Ll8FBzBAvRDFUs8JXnZbb2Ld28/NGp2e9
fQTe51rKL2OxYaPm8sXT3b3EEz0HQuuHIyrVypKYQOdaQpR/Mi1UCfXA8IfDAWAOWKAyAfP+pDgO
il5ddXGDE6qKn0WfdqgLlTPl3lkaOG7UUZ07N1xmf1XuLbm/nCuJfLnBJ0WnS+8RN4UU/sTrXS5r
Z09k70ir3nX9tBpb8bwJdk3mO9m40u3fMOTcDZeAQGUef4XdxHghTqew0bU15Pik3vfGyXUKN8h4
4DlNoN/DcT8GpThpO/sJrtuMF9fsesOlw5vxrQzRnz3z1hxS4zxD8TJYo8G5/7U/Bp8bWvgcAPAF
smjBMr9gs+JApgSujaTgoZ1cqpXve2RSEtyuszRdzGOPLk3EUplbM/y9QIitPysZMXtDsD4iVt43
RTg0b0Ktig+94zMQcOSBf1eSybGdwc/UB3T9XwIIPQUHa4djt4EUnOP4SIgAkP5mS7gtTKWld74a
TvGBYTa436aSt/lRTaEb73FJij5aVW4v/zaR6hjEGBbOcCfbRXx3C4jDfIv9klVgYLsGOuOciE09
rw0BB6YBrphwbkhGr4k55QMEvKW7A0pOesrLFkoa5JsilBLKG7PrV/q+19zRqZ02MX9tBs4YJyn2
Uj8KHnjN2OyqaxbG7K6ELvmkpOZ4zLczPDGc6g1wUNuO/QJLOijnIrkuNYUWCjrT+bBsJGERrgGM
k+OwG+/V3K1qklG8KhqRu8gaCr9VyfsimX6JSGb5Yrka66bpFJ8hOEeyg4BbffzSl+c8ObwpdbRQ
LAu3qP0txRzdbYTEDbwY6wTWfIxtRD2bJz8s5LGAd5e+N7WmvukwZ6IAsknoasqqmcWsMsxcDz5+
FoIYmXEcajzFfLnruldDzokhPFeBDbTd/M5+lX8igdZ9loVwSne5Sljka5rtt8ZZIU7aK4WyBGva
BOdZjdFysErZD7HEFTMNUl0OQOWXyt3JRDXsPoZbsmeAeiHoDwrD0Udk6+J23mrFnxPGgiNjNnPF
HMSQ7dmuKSLcEaYI60zjVyrV7BifFUatQlKTRCS57CDB3x/knXI+KJ7V5yusY1kY/ZvVQqjhiDde
FbVGA0kzFfouU79lLL/y/5CRzsdsa77R/Jy3WMpDMjDnRkEvbNh0X2subMiQzE+mOzxV3zvd6u2u
45oBRWJ2elNM7eKUABrAWfa2pR+hHbyUBcOHgMLChW1MZnUjh/6KJ8sRBFxhlCDFPelxg/GOktP4
rgctBn9AAEo/e/yC9OHt9dy4T0NsNEaHmKXN4Il7yOdnMemIDTZCMxIZTKCcy5n0UydcUMZxr9D9
++49yInINZwl1/Xjd4HoEqL3OICfQ851Uf3gClgzq2ts7ylDgaoUORdChhNg3cMfb7iElsvd7y2d
U1X3EKlm26TQc0lnbIrPYBrxnbSg/TdchT9G2Ws79BpVDIre2xulOZo15ninu3sgX1xcdgG9AsBJ
S9PP3EQdt2jLE3lonRVpTq4y4G8DbTNcuGiWn7RLyHqMJTnLw07KPn6wKLgS22PwLiRwaqiJw4vN
6rO44Uo1wR+2U/Nku1fY7yfUEz9HZFneawzHU+2gpL7Rt9NFbHcy1Ss14OeMcQDBihM5CMyx2TCf
YaREBH65OT7ciwmb/9NXL+UtKaSJgajlesiFiaaBwfo1+MiVIPVXzVfQr0kZRVPiR9OOvrb/eKvU
52S/iY5ubwK4Ru9bZqtfQxaDvKvPR7zIL6z/t7qZUyW7PiJiLoa+qgbW7pKKPjtlFvii5EQLSd51
MbSBpSEvZXe6ru8tFYZ6KI3BVKmPC5peOrvhCRJvHcw1mtiocu1phbBugykTuO1UvZXAbIDFx0dI
4oH/JBloknH2XbG0QwXct8MY4RYPea0bgTbvf//G1ewjqJGJxftJnorLvwOnhLSW3HU7vtzyUS8K
oUi3XG/PvVT1DZyLQerEKxKNut41LBDfkTVvolyLXNRAnuUeZc+Fu/fwNssTvuV/ufltnLJ9WcnW
fbjYcD8abfvu67gYv9pcz2sHAquOLdY70URUh+kNqUOWsOljMMVcZu/T+487kahe72BTZG+5BVuP
Rb8vebdI1AKCUIP+1QAbRD462QWTUjCOfWzOGE1y5VEXcgJ/tJfAe6HRqoqAt8pgQo6y0FgYtezx
uKvfhPmalQ4cxSt6ZQCZUyZq0F9fU2uQ0Njc7l5yqDXGFIup0g/CiCM5W0hZPj3Ov7W2lmqKQQSx
C/Iy5YF5cDfYaSad2yTMIUweULwfNX08+iyA//Wli1eRxrqbVb8dkH95uTL5wlgvIAMLglLcdVlY
bSjtGpYvap8BkRU3/pUpKAHBMcnIKU+o2w6DO/XvG7fUIZC0gKtGZDPbK/Why8O3aWTEGsmCmLBq
kIsm5+7kNoBIwMaaAs1804flneA9xlz9vF4+lBgDTG9AihyHJuaCveNxwyJUjQ3z7w5blpWbTbcF
LQQgmipUEpoJp/PCphKTQzI4iLmeHdOrTHijvqVAuRm1Guu3xUSriOWj65ynJB90ZouyauXbtK3E
oRO7aveO+BShaOq6AhrPnipp8/WNEWoJhxRrUqNYI6sBIwgDBbEHEFKBejKSFY+fVbPShxHatieJ
9L0l4Os448oIVIujA5JDLkFSStN/qT4rCmcW0kz6jLehvCdHmVEKpok6zY9RUtQPssTjqBb8Fb9M
p3wb1nf3LH70D0R0rx7Jx9YiA7O4pCBIbgkB9NJpwOPbll5DjV4AOmn/3HnFCc3TcS7bdA6bK0Yn
V2t5zQYksDBfW8Bg/Pp3HVV3ft7J6fdiVps6fF+rsy8pE5Kqkfj1v8m6EQbTFDgz/779suhjyPya
wiLDiZ5mzyonPhrxau2lGtGTUuC3bz4M46jblOAHD7WJq6BDR2mJvvKz5DfTvpF8sloQsM5DUXxB
9/guHnTVPieHDkNL7K3JjcLqpfJEr2DV3GFXGXOQwlzLji3gfu6WFSmIjWioq+jOHAw/RdHf0s7s
nHS4opSzfl/OuPcBV019eNp0oQZUVUnYwAfWbIkLcxQrctAF0ThYSeLm2rhIMxQo3WNOsRZBnfha
tuiap+f2jkC+RBhr0k9hrvbgWYMUY8NYnsm0srczVR2HsQn59CQ0dLfGKl5/Wt4N3RQLoGb/juOr
YrgIhiw7Fv4ly0PZ+ccEDlDL+7dhBLEpwnqzL0UlLy0aH+rzuTVldVFlVVpPfbiGaz1WqslnPe2/
eU7EJHBPbpBeDLEObe7uOFDfO96CMaRvcCRB6AQcnxPykfs2o5PU0EvSWNCj7xUZB2eRIBKI5BXJ
3dHnx/y1ATAxNFhmwKrUfCjaTfJLuohB3SFt+aMh5NazZe7sSyGT6KgV1tRpvr2XaqkMNtyv8A+1
+WNTWUCOjI7xaLrAuyyXNHFZrLHGyAFRJPNw0dOnnuPIMrWpODbaTPT0t982zF4Wwe7B8/ioC6PE
xGqGga4lqd9KBpSehCXln1dDw0JWTjZiX8uxWWVS+JAnYJBe3yr7QvrDturxcVPN2nU3kiPkldME
GOzps2V0PjqZ15x8XO30SrTdb/VkPTBTqpaRzVzAG4TlluW9ZCMD14W7FsmYoQN5gJt0PCZu26qO
WLBs8F8E2mBDsqI1ZV8epXJdFy/gSBNmVaMT56P7iqfAvu4jtQ5g1KRfRQeD/y9BkNodT9vOZvBr
UZje58bDMiS1Vo6G5es+z059gDQBsRJbxc6JEtnJxvMLcyn61l72BkuuoMNmNCm/ficyuPp66T1y
Sfd8582cPA2cL3nBHQ4D9InKQj0Xxz5RAZMY7ijNgbRik7rqe9P7/gTlVo0D6m09F+34TEAFB7ka
gBSK13NrarEzKovhTjyjZ52EXpmm4DK1Sz8Pr0SxbYu/t9W0rfL0CkFRZ/gyBmBtEIOnipMQ1vy4
iPBpQOL/lYOckoHxi7uBPTOj3coCxReKAvk58Hp+KdTjfotG6bVjKB0Inw9d2V83BRZRFw4RpwQL
I9k+xNrfnyE5u+HnwviisdFPglfcZb9F3rdenQF/4t/q1CKWZb0sfNT3JCdY+FKw7Xoxw89V1YL2
+hC1B1+Ngnts2Ik6s9MCwV2S/FGjQa4vOxFcB6RwDMGom35N6/Fer/V6W8TB6zI64OXfQS4oWOtV
8WUOy/PytrcakCcaunjkP7xQosQYb699ofpaJMWW3ZcFDKeBn/F/vmnGK2rK6rE2u0ZlrnepyeKr
V0GSkBp1to6APdanZfzukCW8NhB4eVuanwpZBu/aU8i/OL6wPz2YlhKYCw29wF3LiJ8mJckdOd4e
xlztsIc9aaTugGPI1dE1vi9JCCdk2TBcoGGABVD7Ceg5tJDGFHa23EmNV2tf+QHdkflRyRYTkAtl
7/jg7eawBx8u3fp7Ua6jRp72tLml1T+feD8wE1ERMT1Xhnj0DPFHQPL4B3rjbdB7V5a8zHl+fuxJ
5ewyeJJHprXb+O/aSkBOwWsBPfcejo/XDhKfFJTBjYyKq7q4rf7usXUJo1RbfiLB5Fb7ZzPDZy5p
YnGXS5NzEt/mFJh/ffElP3ot1j76H4HsqukUaauIURttUMFFKwgA4mkzq0w2reuGa5ysVy8t+hYi
xRLX0aNHSVCma2/DVOy/qThp3ElfEdG1yOO+kgDrp5T4LoKO6Mx5BgXnICLTpIjt/uSRYu7KnxGZ
i6QKwu845CV1Sk37Iah7JyoZlopopKjVJcclAxlogkWaB9f2WBYeeAlGNsmo64da5EWat2l368LC
Ql6YT9hC4aSGMo2SCgJA+7CB1qU1SMyjK5wW2gh+zOPY8QvQAbU5IYQIFVCarwtGqnnF1csLwh8S
+UWthi6yZlRCy38A8DhLohBCUtHlgUATgpsQDrc328MYMCWQ/VkIKck/D6NB43Sb2uqhZOdMvd/k
7vIxAVcBt0VVdHIvuJo2L0w1ezDUPE9F3Nz230ZcKe225o61mbLXVNHZ1XNTrrLzavAoDoKH7nn0
eYMFSKv6u5eYlAqPiSFoMTYAFkOeSeO2kjYa4YZSAZ/Tvxby2PsU7PTB8TT9ljWB4eq8E+Xcrwqo
UlPMWSRaIyc+3q7DQpKhnqZqU3PPh5m6y3VGG5jC0hwASBLjBpH9Yl5zx7nioKCtJwKiWBJ6v4Vq
ftgnYhZAjztQBnsMyG5/OFsF4cYMvyNecgW/cJPv48fgKbgCZ/whtJ9DppfKGFCiW5fajUTcguL3
jNYZPh83051PKQmhqBtYWVrTWSkY+zDxSaJhtCjFQL+fpG7khmXleYa2+3VCx7b1UNrnliNgjfle
GVA5N32dBhsddHPwR/cu+WEHkOeZlFxwhdeAtYjIqWnaDiH/3j2t1KR+EoQzmvpqn38uj1O4aZoI
0DjWB/ZiARZOPBu5vomQcmSRIwCFPeVPC7C7AlLeLLq8KfYysT8wQIM1oLIZADpiRRbid+i/3iAL
Rm9myxmYjcoGG0BFxriV40OMvNeD119QprPM3yEeP0gODZ/9IQkmyrYpm1aBvULb451wnm0qEvnD
qjwvVHFVxoN9nGIK6a7xy80sRfH+4XBSac3nDXDmmsukOtGXogTksn5kbcnewgQGRApbeWOrs5mX
WTJFmwJRUWsqbnA6BwukbfCvPXQYIO9GpJhEUOdiEmg9CCtnNJ+py9awhD3hwR+Ll+7xMMh7wf6j
dcwmukexGZffy/yG3msK+t3bpP4GUVrslcx7J6U2HtRfpBki2va0TQOdPrnO/WLGu87RzB9GzEcU
FhXQRPrZc2KKX4TUyug5IXOm8bhLBG92A7K04h/PlTsn1xTw8I2vkTUos1FpfyI9knZmJlVQi9/o
lGQ4B7sqXOUTegFBeJV3g9j2+hxO/DGxoAcdNEJBTkXxOFHAxhwm3bDjSAJYz5GhFx8X1fRhBoUW
0G3PbBGuUZg/GRwrL0C4JVuiECjP2WMgBa+PB25TadOmX6kJ+POjBrsqvngp/Z1OKcot5QKV5MQX
vT4r5f4TOAqunFNUUZVfe1fg1/+NexCj0x5xEMJqtQizoef1TfHj9oR0E9QV+04u4lSLGv8LrNkj
W+9LwoMvz3D0Xk8AIwmtw+HFJjDQlmgpPFAiP8xwjNc9Ad6eI329Xzsm7/f083/8OmHgMlcFUXUU
rrhwlKIUOqlNytoEEeEngd7P5ptz6+HyL7A/wHJbnjyB3vZRtcHuvZ+A/bKUhEcBWmS2Ld0QTwI9
cjCM9QxWLktMzF07OdSG5ByiQVeK3IffT07YN57SOwq8FIomvMIDrOtVdR2Nx8qTjvG8BLk793wO
Rr7GwmkEGtQcV0grv5eSiTAwhmmc0FIiocziNj9S4Z7ZamCZ0w1H1EyhdWvaAHHcNdRYNu6Cx4S6
qQ04uhiWj3dKZXjgWydqoIusNJUrr+z98TzgyDlrGJSQDhYzetIXUeTHZi1Bcl/maQmML+AznJc/
3ggJA/M+PdmKKx/msZYRQxLsyKzBHbInqWqA9lqsV313ujRNaIqfoaD+zOr2IZBiPQ8LaSbwzruu
1eUJ0U3vv/NjyNqgkBZFIOamDsff/cCbEF7jm+lr2odRg1Jb527McVFbe/pTnCQKQC6IxPcg2TOK
7hJqMIb1aqAFJqVkzoQJCa8LSv36S+yiL1bClWlL0xvpPlAlSTglzEyeOJsNMmSu/jwV/0x0bKeM
wQDLKMqWjXAKEb2mhO6aDIvXs9VCva5PtabDwI7xlGzRTKJ8TWLlinQLFA06ABudNcI87ppuGuZw
Zi+su4S30VvJEQ3QQkIBJId+rBTIP8k/W0rpHVIcr/9eIVMqK7FJEWKwYy5UraPs0ZAnId9vGWMt
+SnUjPPI7YZVfcnTOSoAgjNb713l9zX0cngmDaJVcgStrUWiBjBnrOl3s3L2gDw1EiFnNnGfcPax
kgFx+cMvudf0sUOwDz1ngWvIesiq+oOubDqbqEuJ/wzH2rr/3M4qud5QLoSl72r16AunCljmbht/
aBw77dTPHKBjs1LWrAmzx+YK0b58688gbn/gtfserlyX0fN2dfegkvy0lZ62lbyVdTxB3Ik0hYsP
EAeYnzl7YRF27g+eQOUaPGm/CTsjdQkHHkJrUSFOt9EXvQGLruyYAnMHQn0GhF95xdFVaEe3fjru
ewfQNxue1Xv3P9xKtqZuNuiVJVc6yMfDkhLm9WVd3ESbGfweUsrVMssj/4FuY2BP8RAPdmq7SoGW
cx9DMLS2UkYKxCK6zdHIsFBuk0H6JfpwZCNdImgETeZQuRmrHd8Jt/mDhM8ulqn+QBDDTsbGTrhE
gASl3Q+fqrP1HetmcCy4v5X9Pvzuehy5C1nVZNADIxIABFaNTkqycZzoJcK308jcyCfxWL3UZNAY
dDyxdqil4n8K/KlQOtbEG48Zlls4H4NeksOi+kdz5IuvLxrCjBFR5g6VkCRXIjO/0N0CymHQjn0U
KjhQusHHUQhRnbpNgiQ6Ey0UQSSvvZVMPex77cZPIfWx7/Dc9V1EzlSoYRHGw5cgKXAaLqEza4E7
JzT736XjrEsXFNDc9q9e8NnlDKQ0NGCupiQHY99oCOLYbq6U6pJFVDxeLrA+RCMnXbqTboyJLi9b
mM9pq3qWwuz2baR0cZuP0+InoP+OD3DeIzqB8kgTJR77k/qua6eV1ZUP6tM9EII9fq/mfvX4NW4s
oqOZ8wnS2o1oBYyEQgDR4Yb06glYTv+f/o4cTzzCKAFlnIlcWpO6q0kgfzimxHqn2fug0EOHYa2O
L9nbTRInTwuahv9O20VCoXIkfLWllJctMvVaVnJIFRAYnWftqvC/+R1CG6OTO8jKQut/nlgSuob2
+PtRKwb6J6uPWQjSSSdAtQDJfvbLG01LvT+uZft8bYwuIScKPnZw9Dxi1kOQjc1ltTEH1TzBUcw1
mEGFqJkXgFr6j1BKCWy+eD5NTyhT421mXmylhliEb2J94C3rT3V1NeEtgkpwF/TFBInigVOZ/ZlH
Se8a5mX+Iv/E95NTIFQsPBExIQfl0S2rE9fulFYOqfBZa98IgfACVJRQ2eg41iZHDmy5ZjCWNAl5
lHuxCchV1wOOfczsjW24e57DpFZtH4h2DChNKewzY5QPgho6oXo3wyPEzP9z91gwQPr/xoQqqSDT
hFV3xVmHVuc3sWb3JDFE36cYk1EOeGA8Ph94f5xPLbZJfvj7ZaC8XLltG5PhAIfByM6JeHAjnF+c
W73pg0PpOA900B6kmgTfc0Usm4HE6Z6VtoYLmGkj45Ap/T/+LhmZ8Qp3atywllP9rchj1OagMd/l
aoOg0KC3bo/e7W1VrQeR2XhWyomJ5YerIqIQ4Led3dj4e70skm2FFb/L1sl+sFTnT97FdYRLKVtg
X0q8ph+fsCsK7vMnGcuMW/lJCIg0O/OitK32rwDBeC20Z3Z9EsgU2V2oH2AlEepkAyddr9SJRfI8
3X17nTz3xwJLtGu+LPr8fUAzrmZqrhLAcUsSKmoLVCwIbWNdQcL71nJP7/S0pxrtymA5e8dQlnGT
zdTNJcElcxixzWaaIlN+G6YNhons3u2bnO8/PaQ0SI7stADOaVaMKW+ES4S8U0Jmc4gVyG2/kNB5
HYoR1c8Kij883ih7A5FEjrl1VgSJzyLs56q4j/UIniTzh7sx9J5c5kRQztguleg6rDtxToxVthW8
h4oKLP2YgJV3gBLz50DkeEroCu6uW+MjQOCuvzOXaIWmziqKMC28rLgYgBDtoha32w1KXgLUp8Qh
v3M2sT6JB/nyiMW/7rf6/MvqEnoOi9270p2gyshlocgiz2NjPN/UPx+Cy6PxHSdW8PYiHoCdW7AD
Q1LKPZffm95GPVyvQGMh/ebOFQSDXsWVf2LeMplARLaVf0rBgGCZdPCI9tjB8Q8+cu+hQ1RM5G7y
cqAEFbPi7FbOt4+bOGtSE6oF/J4XI6z6pKNn5DV1kVPzfOUJpceaf2mFCekGV9TbJ5AXoUmCLe6W
5ywPsP10HqDejEmAuSrNChvKCt7O/xAzg3hOV3fJNUoOUOu31Wd/lYgx3kZb3embrXVjLuqKtof0
CFiE2L/9hWtY3cDCK55vhlcCe7EU13T4wDifo/DP4iAiwx74Z53oC/I6uPhyVXk68k+8iFTgdrxs
M3mwrx6xmUw4XCzkHk2UmHsy78i8l+EAf4imht7Js+B09lAGzVStSPwAAmEk+Sk4IpMm92jRdpyN
P61qZC5Vfy6LGJkx1amKIZttKYA4/3tJSgaQRg1HBk569wHO0L07LuuBqOxxytNMDK9bCbohMmJC
vOPiqJlp+BYYGr1gOHWJXTLXNTcxqCEopY2BOzoriNiVVkrYVFICeU/7DiSmszhgOj69Q8U0HERx
SETfdSyq5V+QzAoIO2bM9Ug6ydqRP7A3wvVAPcpoEAbh+JxBChAj9KLxUrCzcIEu5p6euEHuflrW
SzDUAo2NbGutA2hdu57vBV/a2ZcLNaXfi9Mf2iPEh3rs0smQW7Z/nGjodEWbY6RRU908dBVW00Ae
mRN6sW9q6Tfc3oe1HdmZNFkemweHXZg2N4flyan+MfcybGi4vwYbjtWY9s0OCJXqk8JBEvlHXxun
9pgqKLCPZ+qi0Pz2zgkhz0NP2vqrs19J181wwtpbkUgVxyba2uZBUsN62CZnOiIf9SW4UP7y1FPb
Xw1Mwg5Wb9SfVRzvJloqH1B0MIknu98Vw2ZvdLZ0aNOOY/QFnnIxWPN8R7crH5Inr75x4EVbeC33
BMd+vN1Wnh3GScgwZOjE61bu1xNlwUAXNKJ4Tq6FQ9OkgmKu4ViIatD0tokGWBEzkno4Q5q66kzM
aOdBUh6LIRUHM2p+IScaXCwXzN7GG7WHvjT1i/vIN48bz+f1rPErgOzekmXT4vUV9GhCv4PsqWRL
qbu4+7tclwUJdu6LmYxKKXGLZm1qHtCRZLk+jpGJekWXuxqOvsHSonHKEDUoxsT57YxB331L5/3f
2HDikDUtiCfOYOmM0vQLF5gnFH73gP8MvR67OfbEnUARIk4bzSK+eFs356pQTb6pkZhv1uk1t50T
eMwGBP9zv/gQVVOVhGCYYAKYMr5gfkWJ8o90b1V+lWvdpmt6GS/OZDXWZKR8Z/EkBkjI08jtZalO
4yYrUwuf91ZTmDbE1GZhz9XW80LpBjpLWPADb90xQs588ki3tBBf2eW1gr0qZk1493tebGDoGXSQ
vCSrm4uuyrxZaUFN7dKGHwklfq+d3SZYGk4+L+nA8QqCLz79sAAPv6xXyUbuRI6lAYKV6b2BERdY
ScIt8101tm68T1o+GoGlHGTPv/HOUH4MnB5NDRfKIuMXox2JrXFBbMvv0d0wwACpY6oMyolnv7gD
ijlbZw7C4stzJ4woeYfzq6QRi+UoLsrRvyPYvxs21C86C/yEwAM0vZEJ3I+KBOq8ps+JKEn9OLQp
HeG+bvZTyb41m0AtrUpob3Fcet51eNgZRNxaaxdqlnttnHS/Fco6VV67bdhwLgMh2aGTcKSek3+6
HlizJOhCo0EpTRF40Jm1WGIpXnwJABr9Wt3esSuwEOJdpW1QEd4vg8m6ok1PP3j4UOA434bhaTSi
biNxTCbDbirnMzbveJ44udY4Zq/nnP3VurxKOIo/p8YzFO1oV7zQVEK2n77ZK2nw90F3G1DubA1Y
0T3LfgZgv/+XIh05wzu9wX3CsTViXZ5um9kyQBpF+vE2yuP6op/58aXGtC9Nu0cSPzVPcZvv8INX
ENNSColwVYAJZFehy8ZzCvYRVi9YdkHoMs0/OcOp3HulNzWi5DGLqgh+0ozEFYsJwEooCgwQLZfa
S7dZUlByjRmR/Rv3mNPGN1BWrZcWkmHh0et4wGTxCA/VXbHkXHGnwJ8DLMLDCOOEZ4FjzmkKYS61
pTH4l7YtxSMNeV5PTXdIBpKeXFKbD+JDiQJc4sbDm+PBlO5qbq0oWWILUZnbN6RlU/QkMEHAbLNx
EeW08GNbpf1ujYtg7HCgXucCn9R410gKu+7r+vNRDslEC4giRkPmYKkH1na1kZx7xkshaE1rVpYl
ulgiOx3zq21K+VsDhDoSm702V+9QxsEHyMlfzFwzAIQeIODK4CdYl44xPVLv4JSrUSgtLo+nvjEv
R7l3svZ2VWfm1Brw1SqAzG3szKO0RyTqtAWYFpq0hznHT1/Em15qMo7HFnPDZRQIeqs9FrJIIU7Y
o/NzuWMU/R3DJuzWy48Cf41BOiElqk/miLKsg4WkMYT8SKSS84/+5BfjHaDhDMR3u72AoqtI5aZT
gUcZ0HOs1BTlrt38Byg3GU2vOElWHsjPTJRUXYyrARhDzZxOKZdtixn8AJV3dQGI3hpsdjnDBny5
bimfm6RuB8zlLfyWnvHbRwMbD36BVNlaCu2yNznjtVwAjGMcFwW6jx6MG4tepm6NN7c79Y7ycSNk
e7T2yH7ZDwoakcjr3nFtqogdB3pKpf0nbl7Gk8HLhETV04NICJDRpfnJkmutTgim1Mtx0VUFbgbz
T1WPnh89nF25JbIa/5wWSqfekWb8PSUvD5oXCabZm0+RJl9roTHgmUne7Uvh+P7mZHj1/sAC5yES
kwhV4npyDwQIV2GFNKC2Ee1gca8PliAOGlQRcQpQM9ACctdX7da1uZemgHStCC2PmDR49yqtaSPQ
43kai7m9rC3foXPVAGL+zdGMMvnCyr4g/VrlrArYxPoyoJBsADl48IGU3OLxL91LTbFcgDT4kpJQ
KuyovnhxmAyXbE3wqQfjeU/jSyBTqliLfZ47AfQsmFXQVnkPvwG/JaOzjnRweBacq7ue/Ze69sC5
QttP6fSM1IhKHUxePeDHuP8bTonplVYlAYEOeR2AoorjbdlRoG044VegcQFxzRAe26txxZwfc+mD
VDmvxfgzXMsNHp29BxuKBkUnns2R3qLjofaPTWZaKAJFbAjPS6Ksx/B6pxltX74oFsJQutvGb9Jb
rpsbU9OVxODTrvlKwrzzO+zBLsdh0vtmigU0yaJjNUZWshyAovLRI1LA4M35VO9jFFmR2fh5YaGx
XTZ00179WBRtDt9IW2zmPj4EyLLLp/b9HLE3+YD5gRBST/WjRihbu6vMVcWzfp5U/JLGVR9nIwo7
1T1jRDe+QYraveTPfhcCilFoZK3YldbP0uB1r+awB5aDDrUR15/LzvG6kfaYUlnxO6PvMp6OT41W
ettZIzLLMmPCUzxKlGtFb7J4bERkKFG9zqLGW9odCxjIgTgF3+N8N3qx7J2JjYbLZjIuEwXq5+Fr
oIXEkCf0KeV7HDtQyGUxgARAsFDqNpx7qgN+g+FKklXijSmOJ1l8FpCxYcoFCuGrJUX5R5avObGE
DRe8PXB/P4u13+HNdpE6MFoXkgizzd1E5yfn4/UGeMm90k09xmLuh00l8unI8dBM7KBwtZW1042M
UkKMzs9T11pMZXd1inAAp8la68tBl8Bn1W+AJWErw5SMxzpj6LRuNmAhSdFtK0dug0GTBZ1OExAf
MQ9T9n0X5xsDelOCV7XP/TgWvUkK4M9vIFUCkKkXNo1t+/gqIl7wqFEUTqGb9E+eyabHkFvceXR+
2BiF7ldwovPfR7D30ZZL1+rBcYL+qKAZC34BZOJJUfopfb8Giy2S/Jbv5hdkS002f051cIvFYsc2
wGMxReBR52yGEUrKdJBb13G31lk1ctPU/K4iMZYEsnZprH6AFM3vLSKQnXn1I7jf5H/ESSVvb6vA
2d/Ozh3AUjEM1KcPhs0kTEttA9Ubn8/uJJgCPqqYyAZRehwg+mTEdGqIjotWp0AHNlZrME9huZQ3
7nX8g6NEagelFlfnpx1h94adsZhpq80l8AWwWqjLgjkwmTU2/2zNvVKoyxGyGbqHL1rNazUwBuMs
Pv3atJjhurraOQOYYTeIwavPOzUDB66AyFd80CHUx4UOjHupWILabzT80F+Xjh2t1qfNxHC5ZYl0
FgW6sDD+VFvWXKhsC01uoIcmZKLP5R1cT/KXdu7Ym0jOAcp4pxA9T0vuEvBRRhA11LFLidwR6M5C
ooX8TINqvqI0huyNMyHx0DipDw3+Gnl5mtRww7AWGY93M/mEJK+XgsncRfTCez2o+2xFltAu0Fd7
/Bir4yY1rznd7wBjJPAfrjuPfH4u1GfEhvAzhw8PtZjeTqt9NGXUfJdCEzzs057LYdJc2rBgXeIe
RbiuZVhRv/5ff1x8Xf8+Zp4zJsoFPPM6CRogH0S++VA89kSpXSdsLLJAK6+mYGReA/Z81xGw8uJm
HA2LE0zP88GiZ1Ynvw8cv18zwELb6csuA0OF7NzOfWz9CNfUooKw8F4cJ1NSzN8PB5xjFl4KkGsy
PReF4Tyes78oFEbz3Rm9ExbeMMOb7ZFdbZKkOl80et8zwUtIJSpZux4Am/ezioehYb1HlyHBAbD8
hthpB8E1CtaOv21ErHxoJ9alitMTSjC/w4ROh3NGy8IVvTgVKfCoJYxdriM6g120D8e+Da5lu6Dj
aU4hX0O2UF5S8PAbpBopPDrWvHw1t3XdKZD6bnyZ+nWJZCqqAg+cii466ETr0gRw1hFfz76TyDSn
La1q2Z3K5P4DZJpX9+RHTzXQ07stu2njjU8Vf7RGKevNApiRyK8zkwtZ5QjavCfhzMpKcGtjftBQ
rqA4jh0qzhD1nr+pk/WvUFPiVIurs4rVUF6vxCghdp07M2A5PjEibmova8VgSkUx4ZtT5C/jmX6r
y4jW2I5zLM9E1aGcZdfVmUMnXUhOsuGf8Xu+tHBVSqSOrDbdPGDBCzKsnq32foHvlstT+hjmJD1b
q6FgnLra92U6NG3PvRdqA5Q7pIotDnfgle/c1dUxzoWcXmKW+uh81KM88lGgRsFOdxg7vvIGcHEC
bLSa655pwLrkkmSZnY7IOAFPWlxVAj5xXJNIDBItcpoAtlp1lXGTShR6Bir5iQDtffhzlEr2edhC
rj+LhDbTRkC1gHV88LTsnPuO2Etopk/DO23IlTqqNyREXG2429CzLl5VRNDhXqckTBfTqGsmGqY4
Lcm41DIrrMDVmpFnrjFDKMfQ2CiIsitOjNBBQe4AuA7uqpnzhZi9p7LJlJaDIXIw3FPY8BU8N0oV
YRlPfe+gwOwQpRneGFSRIgLKK9m4Opz6ages6igK5TF5KaXV1mRRdBKXzQjvsHOr2PqCY1s2x2Tn
T4D9t0y0I+4b5daTtsZXdp5vPMY3DmnGj0Z1PvoVvyzJnsHiRWOTAkdMm2PM/Q4DZTfrZL5uAi0P
0zwQ1ihOokQGPX2fxnf0h1FB4O7nkqE+w5cJSSZWxmsk2GG1x2zImQ2BpUXOane0Ky6pdYwmDu3L
IIwRKSgHucs+e9ljYQ6KpqUJH/8u4cLAqg2sCXAqr0dGvAuPmdlvmKD1uQuOcyIbZZr721yoEDMw
z9snjQcdYbedTw5vJXC4VW+oBQeyBLOnHGxuvoDlaIprVqu4xL8d3zGjxFkUONJ3Z9iFDv7Sj93i
D8s0e7lxSXNMjClbikxbC2ddXsXaaXOL3fY8kaiBq4lA6ZRDYU/AIoPSbUcEYv5RL4/JleRG7t/k
+ZI3Q6Pjk5TqveyWi6pfNsAVBaUE6idsHHA560IGLNHjovl4XiKHzr+Utiq+Wix2C//is/QQyWOM
gEro4W3Oy/atiN1BVULDE+xuGS2ZtuduWYSaoQpnHL4/FtCzf0iqTA1j5SmM78B5+i2ZA3Co1Tx7
YAzUndKxWNaQyrxaqFpO9heDEQ2cdIYuJeSnt+rHuQ/C3VKddOiHYLeFItXYr0FSmwAbpNIRqBhq
d/7fxRqfQUIegC/X04eL+xxB0YwEQuJ+uCVd3yKLSCRGaiBX+8kkhpTQrEtc6AHXg3GtyZZle0Wx
KbGorhRHrhVB8kHnu07/Tnmw5hvabfbjgODS97hIXW1i3Dz1ejaL3VRUBo8L4eakrbGhZDMtTALG
rYCSdp19cJw6hVnk8LLdUKghCbcZjeaxkDDU0eSIOtjm/tsHvDsZXLgemcAWK1/3X17Q4owIny4g
Bu0t3D5Bb8hhsUa3BgOhXSxBKDwpoR5IvIn66TISDuBEuiDwb8VwlLmqz2gHPRklSbSg3Csl6KTG
BMj//E95GZX1yMYKmNxDct5N6KXNWyK/v8ipT6SP5mcUoNTVDh+r5PS0kBAPAYnyELMIC2qJSUAn
7dSEbZIYWSOYvT5nJ3Y/frVsgOvgjAEQa7G4yXBLkUUN1anwuChUlV5xiywGE4rIRt7w1hvlxu1i
qNabtC4/aOrEWDEudW6w3WyDEm1fsOQSbOW2fPhhKaxErGTe+jklvKRS16XWj5gcW2bsHTCPkkFy
I7Q6hhEHQke6O26YP7E5/S8eXydWPBziaEUzeJVtYuknB7O9Il+bSNCSaulbPjzeElwGNY0ipTWX
gozxmtvxjPEAoE797r8VELiZnSUnphTuqohlRK8gzyMpiwhRuPWBtTBORUJ5qa9eN96KJNatEyPE
JCn+Rz51C68qN9soa/NCk/P+BEHgVjtgReVuZo7kq4Vm04sAq+19IFlXM7pvZDuFygdgI7Vgvf0o
E2D4TwlMShFBHVbkXeZDZyquA4cYQnWx4PpRrUcDkMBqYo+yvdKhRgNI48/vxk9E2PB1SbOAgaVe
THEpDVP8S7i4gefzR493muwWINfLLLA/RvI/X4qz1SL5HE2wsScM3XurCQYwz3rbimOAvlDGQH0m
c45vVgZ344URQ5QQOjEbVrYtgfmPTjKYKBQSGcN0bDosK5bC2h3RgQ317W+8GAZB48GVtlcJBJ1t
AzfbvFgYQXRCoVnBgDm7d3WO7aCvTwm2qr/0iocs0bVVHF8/biDLXF6/OcZWtSD5pKEw2yzmPqbA
nVTGetpSItRXEsHz9PHQ3raqpJPrR2omrzvsSFp+4/g6OpQgjUTHW8yWPjetTl8JPTWhY77pCDAQ
kgTXB94SZX6/LbxZcJwjN1ErwoYUWw6F+qK6t9gmg3pHZ36sqj4u3ArqcAOW/hhM9B4mp6iyMmbP
QNOiCCKsWeQprKLJCoogDZW+zysmf4SwuyWfCZPf1sBMuqBxsxhE09r2K2rRxWHgUfhnJCY+YpGc
HENUerqMayhY1prlsu2lwHhfb7iaMQ0UlgxBmSbxL4D+jdKFUeEPkxH3n9PaBSeKmFzcJOKj8dtq
ZGw0wApQmICDZqqjhzqfjE3PMjDTBpTRXkLDy+pGNyGYQOaP0C2Uh+eSdma3iF35J3K4TGP4EdZr
C811D0OU/ASZlQX/7fDG9tmGQb/1VNAN4yy24hLKS/s4rR8nzrwRgf4D3q7Vw25RzNoa5jIxarcw
1wjEnBJop0hb0BRlp4PpDHNd2vGLV1VSlk/7n5xT7rxsMZVhFwQuagY4lQGtp5cru7E2xwk+UXy2
fvAGvHasrCrrVy3j/FfewrfKXoAaFIasGvWZd8SOpju0tbvWdYbICdFrAjTyGo2Sh0V4IUEyiQMe
6+xDno5+Xc8zgUWjZv40b1k7/xywF5oz3Vz4Aek1LhIEF9cJ6rQDlKnWy1nW+LIgD5Dq9Dxd/fZZ
oZyrmsWS6EUU8wgqsTKCr3qCmbGSVJo6rDVyaO2hHb4uIhiFXfyLAk4vNJTF296tDhHN5snrcE3I
bFDqmfYQjHwODqgMtCDwS9NlOfkQ6cOEFvoHgIFJleqtzBeQufgOHECTVf05dCpqO7ZDVM5nes3r
n/w3F7ZQVjqk4P7K+UYtNZRSQGtgXXxWDnTVqzl2rfoeYPeKDka4kzFaI4tEM2fdp7Zz+4wXGtVI
HR2rEI4vNlrKZw/6qMnp7D3BYUr/b5KyzFIeQVTFLVVfI7UPzwxNUe8VG5pLX/4UB5hZeh+TUhtu
mBu3nKRA7Z+/opKx4RbCMnDJV1CT+ZVOrNLfVLNVx2GLfmfpAGcoggWuTOp1til+9EqFpZPn41I2
27FTPP8lAxe7DpJVHXtUm669bCA1USp61gd59sNllyE0bkoSzBZlk60h6r/7nA8lWq4mVJs3ITEl
LuQL87/eLCv3wn7q2KcmS3f5beTFvc6VFoMSHpySF6WCVSNOZgWX3Xp2S1isFKAEyA0cgAP1M8u1
CXgJfXL1bKSe4qySkNcmXG0qCTAKTMI5Myav+NUHYAB0bBCbIf90yXiVgnq/C5CL4E4UFjZWTdYf
9xw2JG5++BHXMqGOYYwgaLK6GWtYAPTQqJYHUvBayGC24uIHP/5IC5vkOsMMluGQARVFIyt6kNK8
2JBGaqFEbAIXHprkTOMa2IQN7a4HiJCcQNdo2wGDW55Sb5dsCIjmxic5yz2rtoYioniO+ozINv2v
7ILhd5Aalonm6hicWB7yI/IIjiIWN62YLgmet8CnfnVK27n5D179uK/UkzRvnw3CdDjdgVD+Tbj3
2V8swqvuzb2++Mize5LzGiuo978IjBsSIOv+tll8Q6e8jMMf0+o23kb7nPBgHk/F0LAxFTJJeseo
cIym21n6yUb3JsnX5n2YeMbpFLNz24JOpsnDrQGXq/tEFJRI7OA9xCJF3OQ1XspCRIbkM+OoxrSl
LxxSiyxp5WXeWEoP09szRqzjV/BrJpmvffPXZi7u/GFOSlbLcRYz3dv76OM6Jd24upNYapaBUwcU
MAIVyLJyEQqndJq2w0x4SKoY49nJRrfZmkG0KVII2drRlUVjtPlbuW30ANvO80Fi6tkfv75vwzj9
IcLDDoHQm0NkrkBcX6sD75M7GQ3jRRr7WsTGn82avLAMXbBcJmlHhVefG+bT9CxjbYBQtTr1nIWd
cjkbIEgGnd39uSheSXJfGVKq/H8oJJTtU7bNpx4gDI4+2mXaNUuFKy5hhXbnDA1WSNQ5Af1T6eyb
MPSAdSmfqvzF2WZ7kRn8hhDncCBsxWckp6gImsAGRwTfDpvrpQ/WGgoqw4fKiwyjHHdJbOoLw+HF
sD+oN4vwKEC/9iTjML72j2Pv51PIQU+FOKldcbxWVAQdTCA6efEDHcH8x54oNRe7ECvpt9Fztcqe
sDryvZV7S5rb7UXGT/GrfYAWsAx1/5qfzBHsfxlXC40f2k56TqC0bl4ZFcOyygyYzCSC95HiAiN3
uMBqcUDRg9a+L/DE9Kzo8qgTKSl2VVuKVUkiLxB/3OqcnR+ImL0Pe9MvkzL54eTe4YpSTQSVX0Yb
7qmkDAqfJhpkCDq0/alSpTOto/6dB2xpb6lnz2RZaiBaRCH4pLwPKmsz4XJ3rVnK1hBKKXUCedEA
3lANOBUBYZ+U8/9bD8H3JZXij14dZVKXriwr3uiyyZFqodqv1YiWz9cWxE7P4TRGZLmFlGRhjIE/
dX5xlFfO5WoLgwomyeZCjk3gy4H0E1cVY3maLBNzwvX5zSeKpp1oWk+dfPzMAbTFEQuUYDKefsn6
LF5IN2Ij1fkrS6Ish15PM8JskSkG5MZzFy9b3rHua/78waGAz0zG0BT5p5puv3/IIh3iBBs+Y8AP
bMH6eOb+gDR3rkS2X8Va+hM2sTyAH9MkjuUC3gU5W4aykuJwmYTjKW2DAzvmRS24DdsfM+g/HRo9
ppS88qk2p4y0JEaEiibcN5BcpprO/WxpxucyMKTuq5trBs7JND2m8H46sTopuzOWckVJFOZdRQ6X
ZEq/+2ziDxZ+D9KcU1/tTz5X68eRTjtgmgQw7ehR5/SxU62gSO+66PuDgEFk1a+Nh6dBNhs+br4q
vY5y1WiwGwL9+TQYasJqrfC9FPq4Un8gAAqPoRDOoWAwqg5iq2p8ca8umso6WghWZ7ZhhgyMdR0W
rnSIEuB5SU5Q6233qu5nWf2cJ/QkvQg/lJcXsYXzGVJ6ke4WXTfPqYgqKXPzWPmyLvi52rMVwcdo
hQz3ePCOTT1suyTv0sZKNb1ErSF1Zp6sXqvAN3fj+AWY1QwQpb7dXTVkZR77Kwtc31plNf0zQM1t
oIZr4Dua1wjMJB0ZRgkVthFNhqJgiwE5EUZ/HsouavaqED/drk9JyaPq4a6g9dELcjeJjc6gSg4b
wf9YfgFmxeaUatbfdRrSRg3gQpDX3Dtao/uJNiyz50iaxfKixXU+w9GorvaeSd28Z3HtfB/5wVzv
GEZj73EiAPSb2whXeUUSxwItC95w6Xs0orlZgJni5xY9JYK4NRhUMcUNQUBcQJhpEwWXrp+qGl7V
hLl0RJ9emduXyVrzvhLPhMddyj20ffgb9K0c/71DqI6A5xMUcYwZsewuxPiZ5IFMTuvf7GQTAptE
mD+AvgZaX8wx5BkLmvaOj/EFLV+pez6q1qsGk1cRgjDdHNJu6E8x6IX1UqvRqebxb6BV3847xm0O
RiikZwYoL9G5xUNwo26beGG9DRISMdNv3yGwqofqN7MgZFFEQvQVU/AsOSOPcmiXWFUbeksy+vZX
6rn1jxNATyIFt3bRnnhJpWFk79qLVCpeYmoCRnHVokQCHWrCsV6KvADkzeYy+E1F3PKxl3fi5E8E
2k8Zhf4W4qRI+NjTooRxPOrihRJwnxZ/Wqd36eNSCSn7alRgKiSX3RdnDhFeCs2b2IaDood9gSSl
z0coKeJnqHcUhcWZ0V5/Qnw2KFOk4pxIpV4arJvRBwXN9FhdJmxGXZaX1Ls5+WeO3fPtQSiPPcQf
C/5viTcl5+RspodBaniumJWCCs8ER3MCL/eX8nCIncWAeSAwHyD9xRPDyIGUbbFTPWhay3UXi/tJ
ZpofZuNCgdCKRhtV0yeyl0bMrpEDD8d+g7vqmdqYtl4g+RTPWBXrwQlIJgyWYuUKpfKubBqctSN5
YpTucQcwD3XEwgi+canCkPkyY3J3QQxwQB0XeJSQcor8FHvUwUc0EJol/c5T5zXpiL+S9JeAHffN
FoTZWHQFjnZsKcO2m17mhP1IYLd4j+jkvfyviNKoUao0yljbqOPF9qO7IAbSCmv1qHxCjSrOiwDl
GRQV1s95TK2g1xkYcK14dOc+Wvt3LDNl2yQqiH5aaw+2oaeI8R80VIvJFPjKF0X2fWXy1i/kSwuq
X83Zxl2QYPLDq37KNodlEQz2eEWEztQvJr11d6ALCwuXJftZeSQrdjH7yZJY3zw9BSLIVZmPlMVe
UmSDOQB97kwQaDmwmmhEAOl2Vy+5qnJJNRjJwxxSN0e6Gk5tPzPFFKwcbogL8DbUsozMjIGDzuhB
iiC+1k71IAFbHHmT6EI7WhUjWeaJ0K6vgE90nqYXLVK6UdaGMedJxeGdCi9+zlFZVHTj2hyhjOwO
sp8Cz0H2qe+5X6TLns4w/nXXtHTBReb1s0/RWkpFzsXHhm9k7YOm7ev1IJYTQMgedClrnT+v7qiN
h+vX5igXxph4hrkeqcqFYS2BODDRqZtWZ/t0jIsrO5Z50NyUZvt0jh4GWTgAs0/dBJSE/UlzERDo
7iMR5p+MPGByK0M0ittIjvFFlHBKhny1W9xn7is+kgjQcTt+6+kg7MOu/iOBTHgVY8eCUE8b6m6T
pP9PVpQ+Cu7dcBeYB5pU5/rrDHoZjehms2kCFTk5r9V9g1i+HgYPDGMlZPNtyKuvSzt8Rtgv0III
rqT34Dcc5kMFkQAg4QPNJJqKU6ON9mLReWz6TeqN05zWywetzM9yNzEVctEFJLuAMrt09gjhmNy0
MJ4JzhTPApLMDVlfYe8Vlj20OH0E9sMqMT5RsdINLitlTzbWOExk2uNeAAWERO1yAQIbVFeojMEW
a4RWv4UrHcKVjg5wnd+JNAIIvE6lT94Irh3dsfGratNJecbKYzgYJ7xH+CpIflUEdU7ya2PYGCWh
PaTUzgcM/4Da7ICehnhsR0z9FFBPL0iYN78+agofXPiwZms/769XsJr2YiwyPYp0t2g/rwkjWkrt
OG0D/AQ9I+9f6jKj4Y4UJPYKdlpH3UzKt8sZ4Z9xDsI9rkwRjrKaezd0xAm1JGe1y/Zr/IytGG4a
RUklU+wm9eoX8h0YHyjOb9N2Chn4vkdqlTXZ8FfuXiw2bGHxkGBoZ4xxNrrZhhe+GIyFQv0NyXqe
i914IurW6fTbIv8pC+XZnL3Ths6TgY6oZ3Zccq0Yf5Vp+gu3C/VWZBEYpXwu3b5v43GcQOFWv5jA
Bq0KF5TWnE+L5juwHJAV6cUEKybBHj8EEjqk7jHgO1K17xiwxJjnezVzhQj5u5iIQXVf61nIv79f
YorzGuyXvaCMQfS5wjXQMTbN8Wf8BlQnP+r7EVJ4xTTi7DItNotXNawVKJ4WyXhSw9X9L+0zjwtB
ekTBWrKSyWtPMIm7/Zm9CgGM2+z0lxe10jrPo4a2otKy4oO3baskpKnanelU1qGMH4eXxR0pang8
2EBMcRc+Pkvz5kacTwsNetrCBtOnlEvYkDC/fLmyywkXesftm7O4VFFeB0s42Oe6XF/jmLBMIqDm
UTQ88SCfYTIO4mNs1gcOBYu+W6rbQF1/d6L/H9p8ekAGT293bmuGgFsMNaLgHDFCNXQN7hLrtdxN
t/BfGzicf96WYTI6dcY8vRiM8txyW8ZaJiOeTTRjUp3USv/jFSj5y/TKgk1sHMrSOm6cV4/v6Pob
G+0DWFnLQecR+s2NGTOcXi7DnOOfmwIOvrfBYYLTGDMqGLW+BPqKvHMF5L6nMe9TJ+vDtVD7mL0k
xdLwOaIGbHw62I9iZlGjVCg7a4RO7ufq/yO/8BNBjqzXAgMGrApGBs8lYFT4JKozu7mfleM0psiD
KuBeQ2hlLnGPncwBmlV1pfE+y62+SmexWJJ2aVh5P/cZTYhjJ0nu5bpkClo/cv2rIKQ1o59CH8wE
enjCL3rAKj/R53Sm4lQEUamsbqE7n876JtF/nj3cIsmOG0EKpE+RQJupT8+49ydCXdRd2BymwR0H
KKBpcRC7amcK2sMvRQSGF7GZA20eZxfcrXiAMrxvqt0Biv/Q4GqTQ61W6Wo0uv6i6hz0kZy6skkS
69PFVVX2m0GmTELGtzR0ba7W1oiQwBmZ++Z5QrqbvkFTcCtI8MMCLWvoOobKlh+DoJS585F1V+DS
UUvlaM6gAo4y+ro/c85u6OkJdT7RiodtcMfdlLYb0XvltI7PGPP7Ui0GeyXgFF8nEkVTowmAc+2s
svekarjyJFJZEy7R2LU5ybbvvgIqEMWAfERXmABKEqeGI+85jGW4h1cWVO55qZEvIF0O7Q/kaBS3
wdj9zf4WbVI43r1lOP98arcAFkh6MpKUJ5XACVJjf2z2DPQR9Q3QKnULVC5EIWT8IY7QH24XY1Oa
YI911abnEGQKxSbCElseDNef1S3320hdAaJaZ6GdZ0WTSGZQPh37PW/9mmZOkTC+Zqn+X1iAz8je
F3G343R4IurbmQVWnpJsXNYw7AvY3wsmzCISb8FspRgjyE1+j1DnYwfFm9XL4o4TJkZCHGtBCxRI
EwZT8SUVCXwRMhqY2O9hnIL9DZfIYw93LWs2UNFi1fTsqjnrVi71Xg8rp5Bp+tyc00exKA6OC240
lDqwbyr+8SCQFb7F44PGK28VM/fvSaGlmBxf6IVcc1qRgBYI8K05G4iqQWgWU5RURe3dkzAoa/MM
nWDVYmccuBLIkXr1UEjF2QNNn2OgFy19jGW95KqP1Z2zpROaGNIkVLhT7ZlJJ0/mImQiJ3zA5lW3
LVbzsqpF/kGERYj6fsAqQmcIuukOIC4kaX3z5BMmFbh4R460QjctgmHcD44AsnbC07C1MKnTMp7w
FpG6F2al5s90BC0bfEAuv8/Xz6kMTlopEjK8xh8u55cfyw8IBvogz2XjMdiE3he1ZO/TehpHR+BH
geIrr0YaIlCB8YSfe+WAh67HDDqoCPndD+dqjrDU6VNNvwrQhLMiCtOJ36LVV8SvdAD/+rJsdRdp
qcmrwNZ3XjntQ096h+AR1OaxAanSVnWWQtCJO5YIlAFqmUmk+s1DpeIzZqNIH1KZ6it4f3tLVWbd
q5nyTtePkepMlG14Q1frJ6DQkGwWyjGogLXiXpyHUbO4FhHJ78Zeu015Cj1sj/hklF9ecuFmr2GO
TVoQ/TqaKGG6LxxcaNleqRh9FSMRTev4m1wApd+SS4au6JDFJBa5VjlZOSQ6HqpLD5ZZVQfdxOxA
D59vc/krMgO1jaIGJzMpyCqR79jWYY2BduCzlz5L50Q1iAVUcBASxIavNKeTK+hX3OMOTAiovI+w
F8dZXIMCK2ks99aSScI1VuGqIhI3gO1+1taQ4Z9IdZUuIys0qjE7piHqlHY5lFACkzNjvm+I6kYN
g8HpxvenKZSt0zZMwwYjNhXl/E9DNvFVztZLx8cGfwhMko6p7/isTxW9R5e79QCrDgSjdtoIv/Df
QrxbJ4EkeClevR5Wb91b0aWvEh4GynPJbuu7fj7u4Ix0zdisO3R7LesB9vyWqV9wZnKHbqEiYMbR
fujXjkk6kAleZWrS6QBf3plxrS0/LF3SL9yBM+JWDfxzRjNXlxNk4IuXUC1+qr4P1dIXjprYuquP
lKSd1F79YcDRlKhNKzMabNYM5dvnVTOzSmfIaZmK5o1fDJbsq2Hx29loNIoH7tYxwigSKKvmD79G
Idu7tXDFaJV5c9gulcy5GeiKJW8cXEmbc2F4x9N7J6Jy1nWzFT8MSMKx6HElYvIFXcQmwmsz+fuN
t8CS1259HLGtKeL5scUqIuGT3V2TcI9PHdISOcn/b9mPD8KhKVwGnoqDIhJWc8u/k66SDFYcYarr
IJxAmBuXohSw1FnZi6DINf6O2KyhhMNBBmx3IoEzpg5Rck8kvIq7ZYNPgysfVpLRoUEf/VludBSy
frjPNh/goEU3dirgE2cHO4MOJYZyfQivnUPMlQVFdBBqjGU0a98TtwtKWdieknw/9SewsUD6i9Jr
lZlr5AWymWltSfuhvCQmOhhSNxa06xFcyzCjgUJWonJk+7nNPrmoL/YM2EM1efeumqSEdD3Ilplo
kpDWplyvuvhrq6gQbjxfYLKSIO2MK+IYXNJh4imIpAjetKMekDgVtWGCVD7hqbCS7R/hohIChmrC
5Idh5+2YlDW7xga/0t1fQzdyWlqTn38Kr73EoN6De7ZqGxFvqhbObZ43bUosD3mWrw+2IZVuSzz4
qyExuSaAxZI3PnRYxPuOls10MBGuFeZ7sT8hBJwxxOeFWktalb3r1HpfxYUSeFV0OKV3G+ZFkKLx
S+O4P1Xs6BqfZsyzgqAQV5T7aerpI10sNK13ndv8OK3Twj7wanSr9Z03FYxQ+QjzJpHXLFCb9P/Q
+aSUPippPobmZa0VytcTym6cCJLCAkQB/VPzVWYBB4RESnVM3Q07xRua+ZawD9ogiIpeKAJHrYDG
vz7hT2wNOX/3KoAeoS7ISGiimzI8B2EiXHqHiG/JuH9nB4U6XqAoLPKDMCMp5CtPHO+Q5KF08h0o
vHTuMQ59hcpnp9kLcLj74YSMo8Q3EVcQehagj1qQDczz97l1b6GNs6gNdV98KB1f9l73BDH2X0UA
1VAdpfdFx7nTRz9n/qzqBCp9bP/Krom8HEUkaEMKAbovLdBYjIsrdN5Hxn/NH9mdphnjKiIDSHHL
V6yK4OQfOM+ISpuaujGxK2YAxB53kNgNT6Q3Fm1sVFD7M0SHalWB5oFk3IaI3/mlOkau5eK4iC0v
Oefq03NJCN3eGd/RQqdU5KOwLXhkSMgMvpF/VhtqmXgpxrFM7gAZLgHUCFRLQvNjd6ffcX8nYNXw
oYbUFJQEg3MMkNqxlzqwqjPmnE9276GmFcJOhSLT8DpdPARIhYbR1ozWu2GfS3AIhWciKEVUhgp1
Xhi77p6LSgCBftP0XGLlTY2QrWufqcEgMixIA8gyhCWIWokzTvOKpZOv6VVcu8D8JlkuWfsnsW0C
wxGxMn2IMsTPSre4ZuU4Ph/fUjuDYZFAi+Mvpss6V/9ZpSED944BdnZQv0WZlYFp4ypsDGZGkCgL
3Nyv8LeXtC8b3U/GeLMZ0ji2ImQeSFBFmFy8cMXQovx7c4zow2mfEKTZyDJNb0Gie57u/edPPINb
pN8+DFvjx5QM7ZAf8RDpqFzfooZSJOGSDxDl3//H7P/sjw6ziCDSBjTIgFGWTLdRC+XrFiHS/1m7
ev+x/Vjzcigi3Vm1Nl30KXotvBP7lExcvMVRd42rWnDX8SA5x85pJarAtYE9vLTXRU31noAEsHt/
BezNRu4dhTqy86LtXOSwKSMzPI+HiQ73NZfwlcb40dURXjHU5DKJ4xjzKkuRxHxdMuwLwfLCse6k
D54IN/uyZSCNGT9c2ezy6JlkaoI39m7Fb6fTDyd+EDleEQqio0fq0bgW285nbsbve9lmND9A9uBo
3H+aPiuHN75kCdILM4Nei5swNdC+xRjoDcorsfoslZdK4Vw+S69GDHSnWL4UeK+BiSoUd6uLs+jv
A1CV35MWdLQEQwets794L1dsK2xq8kMTtud1bUvucRdc6nmQzrvWZIfx3z+wrD6PTpGljkVEs1zX
Hi+y1h7ItsT6hwdPVJAGlFW0/KfDP0re0fjBrkZozrVd9c084pBKBEEUJlLZdV8JFjWKbU1kwFZr
rdcYnBdtnh4ei153gk7V6Utk8EZoUC8cqRzDTRa5Vq6DbNpCn0Pdu3kavZv9F5Yn6vKp7pnk0o55
AuJ2pkTUkBGQKm775pJxDCWNJLhMwR3U2R2uOxaZZpz7nmlm4jo+zOrste/pvWIwdQtYNMnU33ki
JVwXqxXI6qDdOL1Lb6TARf3FurP+DhvQdfI2CDqwPGGPG93BFRQddeY+9cjabjrbyi36j9T9Vwbk
QA7CbsCMasv/oXM/0eiPDgJY7Bq1gvr071GyStCYmgX2RuzXEB+gwAWQFM+MJImbL7TJneJg7YtC
pHO8L4lSRXVmHUYqPfy4pgfg2Enm/SwuddbTpWRh+5FG3VIy8R28sMt3GtSkvKVXbEoospmPgQZT
m9eHADWToAHlaFn9P4EpagZ/fr0PbVoeG96Xktd30Xr6Rznh9IsdRfN4bs9ROfzguetlW6i1x/Vg
Y+Z2KHEnQ+RmrvI9RzI/w+QJwTCNS0Fv/pRjkXt5ZYhdIDBLbdRJkI8FhO3e334tVJvEB9AAkr91
iJa2qouL4A+kuFlqF/lw3pSAbozxheXFUMPGDjNKmgXJh94o+UpTR5ghNsUbaOvfoWbhkmHYdfVg
KhZc0JVW0JRwRVuvVsBZ9XYmOa/r5WhApeQzXDuWz0pW5JFH+cb6RqHRf0EFb8a874cBRYHi/leF
1B0kapc5pHjqoiVlvyTB7RVoGa7LRqxPq0b9Y0MS77Dmnf5RbW8bTr3nzcWjZXZA929ggAXkTccd
Eirfzets7uqNlD5Ob97r7VCCtQATpo7Ph9ZepA8iOIfttUuDZBClHKWrACEo+adIHR8cdlzjvUN3
okUfA3PV3QAyv4bePKPphk/xiOy9f4QWUSFLAeZ/IJaBt76LDAvt7Q6VGsP6D60utA62Is2Y+zgK
+Mzm3QYGlVoEaZWbU6sG/+2M0UYGpnpfFn8QyA5ppM9KW6gM6I6/ZblYfBPObJ8gDMQUpqGu04FX
StYqQPFZA0dEnTmi36ZPbwlPR4eEOmLnJ1kis0v0cpw9/VAuQRtBsGSFjrHkUydpn12eKHpvdLQ4
9hDXBQnPIm75Eo3AeCMl7tmEysbXB02dFxDDAKIcFcvaRMBHkbNHUjq25vJmE/4bi/uq03WfVS3o
l6nukIeNU0KGh7FAHkCcFv3ixnI+7yCRGxbtwjYKqcm0YVrm/6kCIPTK6cd4kCO0dxSCA7nWEAP8
3YzQKFj3up/YfTflkMGWPnFlt8C9HQfZFTFeCKs3CcI/N2HlFFXN1yJuxumRCCii0pYpaVsacjdr
TffiqtbrL8IBErgd2d/iodcRi7/VbQ2jw7Gl54TXNqjMObqWZa7eENI/KT3kESUtx3GPufKK/Dl1
bmln9zKbtcajVH6a4OHuIIx90HMTplOBWYlCj+01nkHFCAvWgIqgDeyIcVQIQC63lhYi49BdZeEk
/X1G7OZ71skS8ZAyWu49FGHdnNnk0qkVcO1R663WRCROdvROZTxq+8Te0AszJ/ISEfeOOL1DTpjN
yRmPYBGHMDzAeriMinFFAagzQw7nC5eRJwiRLv20kEEpygYCl5syghrW/3z41HGeg+AIOFPP6rtL
yIh7lOGaHNbQKR2xYvFadTguqXsiXqCICgcbIKY0k8CpAxgG80gT8orjf8IXu6XVygWyhI5EChGQ
1lm4sTN1U4arT/0sowMQj7Klsbja661uhtPKffzSY6LJOEgWBT5MMl8XGM629X5iWt5+zolnIJYW
QBRf0LRz+80iLitl8UymgVbwPBLRcX0ovLeJlQwoyjTU7DJcIyyWXb0oUIen7mitDTdxzoXSvKdS
Bg54E1XbxQ9w0g2jCoNmHFH3eunO6HVGZ3i8uf06VVaebqKs60MMPVk/9Lz9Fx4eZkCAqDmfQa3e
0i+co/60zRjqRVNngfJIIJ9iUrLdiejne+y0B/QdPypJWy60Ofu0D7haa3fkByGEcuOoOkk2WUcs
DgZimJ0r4xSKb97Ema1+DFiR6ElrFWTz6Ug4v0Aj1Oej+WrgXyfm3Pw8PVEmceE2Mmv7qG8ELatD
Ywr6wzkCNbWHr9dQiIo5wk+V+JzRLke2pwOKirFry1rrvk5lMic/IKhztOmCgydEgwd+IYqnQDTV
CoukByi0AtHuAVaPLH9oERlZBrbZ8UqasitvFMD8Fo2NhTpsK+4yFr/ot9wtY65+lEbXLawRNoSk
5i6sOnjQVZQ/FSywGo7nStC8+qIx6WOJXr1/YSec6lJyTOwI3TsNRDFUY8b7m1FUz9QFK1h4vDDn
AcF7fVoP1Uak6BJuTGiDfsJltfg1VYFbTO6TjjH53T1PVz+9XN4mP3Ar3Kkj5nBCninvGY87JwZJ
Hf+KG+Rszzh+bQi7buU/SbFHD3lHRhJe+q3XQC+1tKbav0JLI3yDSaDLJf2/YvfF4O+3bIu06zuk
AQGu/JM19XT9q2Wp+8pQURQIHBEFalEQK46j4GlzkwsRRCyzVS4QqlIeFNbzbv5e1Ha8c3gkMZMa
58iTCW35zHQs8OokZ3Jke2XIIHx4MAbkwytHhkVbFAiXiCdLiPTJPnFHzzj8NZ0YmLNObm5KMIHT
B7BdFpqtSFr5iCMVMSZ51DiBKeH31rr+Iv5IWmNcPLUgJyavZ1p9BzWHdt39RBYyoSuxh/JsjCN6
dsxchiUHsOglH1Z9dQE5yD+DDLacVnXK54iht5W7vNCkpsfr+G8IGb2DOC5LhWmSKI7PjLROh9Jp
nXFq/9ZJXKfiNM/I/u1jUkSvvvNPf8D62RjpknCKLvKqFLR85R6Bz0UQSNHzi5IlrQenobXQim7+
/yPFRIDGfW8x6z8KKuWg3p/uzWPSD70v0y44GZBT9ZQHLa6h7AsPEiZY7LagHQzRj4xbbbLXPy4H
5ARCohqXgDfHoSAl+K1Gwh2vYUJa3lpwnqdAAvchWpKrw2MPxa31PhwVi+xHS+67wG9CrAqtU9Aq
08ZUlRvagjq7+qkQelLnZqomhP1IJjgBk07pqM+uxI6YUpXt2w6EisZVHhhZ5h6IN0lLF0U7k8Mv
Tt6+PNHC5K4fK0jy/FFoLlc5pgpUFuTl+tzTFslNWzdlhTKAB0A4MvovmtZxIsjNBB+xKQy26I7V
BlNmpkCgJUvrvtnVV2y1gh7KYzdRw0OwIzgOAR5giYxDDCoIccLOZgr5+xrAG9LDg4LU9f5HENe+
ozNgzxZpTRER/wgW5cpmGxobXA25+xpuQYalOCvAb1agj9BBVBU74ApoqLgofWaBELRwGZD7Fk+W
xeKYm+/WIsXUdVJUktLzq7m9/Y8APD7N5c/Rak0a00njYuwLK2kfMRlFn8v/BvU4i3Z68r/0RoW4
RT9xg4XfEIgqYCtEGuKyZdLBbwMt/d7aNAdhlqvcC4TplC5rrnefAq8Mmv9iIX8dmABo7CL+2E3r
ibCi9WTEFK3TwDHcWvQAXp6p1aLraIG4oBEn+0DR9yRnihEO/50DV701iwYhIFffsuxn395SvXu/
76/fGNIRBaYpBWsbBEhFy8mcayZzAYTgAfhZ0YjzaE93gfLvrXvkYTfXlg21ALyoyBPjOeabLvFm
Gu91UhDlhocr0aVxvNTFLZafaBEZ9CgoyXMpUXUVhp43/I3hFIMsgT9x7hWcDOaCocKgL/l3wXdf
VaoDnbyw9Q+9CeD8iVp9ULgEonBtP62RvwBpP/jpokTE5o6CqWG0Wjvxm9s02yBk7dML/8Jgfosq
Tv5eoCUahm+MuyM9eAyG7fDG3FmMChF9TP1EYmsM4PEAMOxba3xAEeEbkdN9QzQuAm0C2tewOzJE
tTdik0pCKWMxui5TbEaaENzxYGXbWPgWXQKpjGvGOjGXaOnYxWSDn1K3HQb1dp4R+WwAGklrN4J7
ptgYHH0f6AxJx/nW+/7OTuJVQTZxr+GwWxP/CbJHe3RC4P8Wi0LwMhFwEv9Rjb3jO+adRMXzqw1q
3LxjsKUFStr6DszMP6rt0DPPDo+/qHXt24wRDm0MJ6nWErxHmkiuI8k0gKZHicLhrNOutWtGJZpo
SIWMTNVa8rzuT0RAptyT8hbxui1k3kmkjy7UwWH/mZqy7rFYVWgDOiJN7zYpYy5FLvdyO3Fwx6xQ
FmZoaLqXgcRLU/MGvem3sUS+6Gg6GixPSaWod2t0U3SfiT0AUl2iONPbNpPd+q1bWrIcGfdWcDFW
TuATwLWzKoBlrfSp1FQFaqYNJ4Qis0aJ/Usvr+iBhtvrdWcktsUS3xl8hO54KJVbJ8n39lT2ZDvP
PezeogYNehUnrdXOzNABcTI7coyBJDyFGIgxnd7PVsyKRlQGQcPe7jjg6dvQBZTS00PWVNxhHOaq
p6rD1kMrQJG+LPbeuorUZnV0wKuf2++E4iFthaL1Fd/A1ImwS77J0+1H3pPdiGJRAM6BHem0/H/V
hnupVQAiArlHMA2mSEgjKYwNPR5i8i+/eoEBiJ1y1vN/lz/+CkTBtgDYdwrO3hVolqFWV73h671P
m/wgZ9c7bECitniLeqHhr4q48gDVWxdMs9W59X+uRNS72ZAEzOunltRF4rJA8dkAMvb6fVcCHOka
7aYv89cTlsB0mvfw8zelnXRTChuDmVAW0I0fvVMrRlN6F4sMon8x8ARIMUxO4VBK3+wrWsz2HCmc
0Sfe2jSlOR/XdpanLG5GIoGYdLb+3yBjyETp1cs9C01SJJkYAc5tGldtumJdQ0WnFwj/iplbMNlb
obcRtiSFAZi65ssPu63GETfUz9bIFwe00yVnvDHsL0zVvLnVsgoA1n/R0q978IZnN/FSa4z/NGrC
7F+lzFAIijuL2hGKzC4fzXX/QRgf3sj5ukd6k0ozh/Z7zU/T3j0SWDxk4D85go+QkzgcfnPGKn3v
qNvKGiCRE9ANCptEB6amOBiAGuCEhmF1GOw00ODMX8wAlAJoJykc7Rs7z6QGXx+dZWPqVNjpERsY
WUO01lSy69H9Uxo/Ug0XSytkslY9ytgOhQg5MimR6vr8L4hHtTzmc4ehOllV3Go0KdI4xtNrmdpv
XPHMnWVhU3DRYIkVMsDmdtH7Jxq58mRfTdzE9+PdSKLnme4lpw36knbqQHWBL30c97Ls9Wn1qL78
8HvgVb16XIgXCDYhvhrW+4SMC12+EpruPGm7u9HRovOFCpqmIhgOX1SUsemVTgydd5kIkVnsANHb
dI0LVBnDwEEF/ThAM0A8eIPzAbV6WZnl7F8Xn2yvOpla7g2reekw7CmhH3mLtH5fpuH8sC3xyvfD
OM5S60GeDAXjkEuJ0lMzYwk0K7lu/y1jyl2tQ+XOfnsRdivrKbtBPx1LdVJOBMS2tKv703m7kxFt
7SmxUgqXTnnIy5740kHeu7AUaU1rz/OCxArhL6hri+OFkFRoe8MFFwxwTzVki37YNzWcmxiKzSzL
yrRr6Tf4NNa40GH8cs8dYBohJuBS9xg5Ge7rWIMvUfVj4Tz7k5PfLnOjL9eDQc7DhOHk7NSLRUIV
DH2TiYe/vGdusbGtHukaHQhBX8eBhXbnTZTkYXFb092FN5/wlSPjntlI6qTW3GOpZTCFPs8lYR2W
KRIPdAAY89Zp8ekwPvi4g1zImMhhfhyaUhuky49KEF3RmKzy8YWhQzB4t1hEJDvoQUGP9ogSUtzf
nZnRWtNJtg+tmTaMF+dIKDleRWLXGFkYyEYohJAYdRJ60ZzObJMUNPeacwz1bpJERe/xYx4ijPvO
HbH8BBB++BCgy3zrhgguhIcmrHj0/SIIWdpbMaD0DMUdGVN+cThJyWGV+qAB9K3eSJvPzO/LW85C
z+8ed5qQWvmG/gmXkSVJlapmALIt+XWzsXqV3ctVtxLDWLYmzwk9hmiJJrSIaRchB0/OQjYrumWN
6NxkgigJzYyZsV7yYh5nK7rGzVNmMfePkH7iabOaTZfji8gCHoxzYYdhx5f7cvllwZ6SrR7yPpD+
in56+QAaC48o5ntPim03EuizTmiDTmInKk6AAl73lEAJbISx7vs6Myo/TiZ/W91/mXsSQDdLUxK0
J+Ef+YyWKjRRXet6wwBbdvMFMwKA51RC786+hnUKceoGyuoA9OgIqqYaObONatRuJLSuDe6jAGTt
8/wblET+S93SB0B4QvfCBs3Jm4aRe23+13TJxrpQD6gT5sqQrH2AYlnEFFql4vxWQTBinbpcB6b6
sek1HQ2l3waHfukLG1SooJRPizraqWqkkzQqRxN/s8wgEk+QtZ8Ljxn/muvJLYKuZpM1bJPeAhNU
j9ZFJZ71atTY1cPmcH1xM4a5otN2JYRK0xV8ZdtPC8vHwdxhy/nOoLdLEfOOPAOpt4VnBL6sbQGp
SjlVxFMRMLhuTSntK16xqsCvemsCIGAHgJm7m4cyAsUhAeT/12io7wF8u9iEgE4HLSDUftlZiqtr
1E0ZO8R98HFF8BNHtG2wt5nj1DZU5F53FgDocaguyIftI7A/Iz8OOh771U/Q8WbMmStJuqt3iO/X
4R7BYnfUgNy3GhJs5NxY0iaLVm/I46D2xl/rtdxZ6+M4oKUo4oq7G/eDtkP3ZlwWJUdXgS5nzne4
qiT0WRuOskSieUxDBAzHa5GlLpxESDTpfqqZkDJz7XX9MdMdTtUbPsEOmaXSk7etLW/SizmUdXk7
t0zXt4/vnnaTAtOwpXeQmb93F5fVKC40kdZJHDzEm59oCwnDWGqFyFMLQYt7VkYE2gODV62dKzDz
n1u9XueTkdLAtmMMi5tSW0r5PD2uuHVOm+D4qZFGJJDO8PHkAj3YHS5tWv/Fo9R0b0OINS9TH5YK
G3WnjqE67RhsASqfdxLEHmJacPlepnrh5a+AZZfuxHEB/irPJwDBwehgs9KLq4xSOxLgG+nNEvCA
MREry6QXOwh61/9e+zJlwigSEVSvpYHn45TMgdB9CCPHIYHF+dul8Cts0uZmLH63zSNK9ujHJgnZ
861Ovx1CsN6kwehubPdgNnqv7hWZfc/iZ15Plg6WsiZAajSGGiqaYhvYLsgE/3ZZa0Fhzd5z7ajy
Q0GN/TDhK0K81PLzyNM3eGczyTkELkoE8gL/tOZyYPejr03uxmICZeWhnOH2VZF3ucbTcpkTwQMV
Bwf/iXcVYirAY3VMQK3V9VdjnTMfVWAiVEyQUYMJfaa/c3CpeboOnG78LcrPFfzr0FRUa9ctqtrX
HPckT2d7UEe/1hWGRFOipjQWRkITOxb51AjnK7QICJZ1Hn8JubaiTRBxuiiaPt/Jn4yvl6LeG2oL
3d2R9fnYvJ2Lcd/6IAItdAGcvTnZkAj1NN2Cd/mfD7xE6U4KG9hDkudlmBI7Kbc0IvLMpDhrIYrP
16sqqAJJI/XvKqoQgRedayWVSzcfqJLXRcMnJGLW9vIawsWQyAN5oKSnKwjgdvB6+29g+sl38zOu
2d9Mfyrp7HMUnoSCnKkDQ2GfZdBVbqfOH0/3GbqNFQ4+rdo9PStvklgjedYG6Tq3rLA8XFk9vhSP
oG+MAuW8Zsx0Z0h/yRChVAyDPof8vX4pKeiV1cgpzDX9QsQ2Y+MgC/zGC9RvzdrpXtpH+xAgaTeM
c0HktE9G1HXzJnqG260NlkNg2pKGP4JdB9tO7LzQukvXZ9FG4kUj1bi8wYpaIC+84U7L6KbWApPO
6N/u4fYKRMbfQ3PZAIyaGw48NVXawhs6cKWxijtmrNROZKi4tTOYhxwjjVoaQJwV+8KNdWQGcJXC
CWZ5ozV83NummDSfLnBVsBembW4dDrEBIvRptDOYw517WDnEcQ0/ekagUN0ApDTyCJL6FlHBIV+B
0jxXYvKn3mp2PaWmFZpnkFO3H/lU7qIa073kSP7udcyUmToMf9Vf3CcOZuU6zW5dsejGRAH1kmci
J/JQi4FsbwrG8XUZcbU1KwuW20V6ODIT1F9Invor4XjkP0syU+qULqdR3Q9EURuqHxOSrvJfueY3
Af2zfRsmH+3dbnLTMfud/8zok6G1szqnp7NnPTgn//uLhg0yTSqon1Cougb+CvPL6SAzkRbKdKpI
sWlieYkUe2EiWCGij3dQ+OkHSUgKr2ujm0pK3EbwOhmuKoHAgs/K7mxtY1z9Ye2Epe5KJPhYTz+N
pysLh+BmR2xC1tnLG/YDib993Y2aTdoltKmn3Dup8IRJKBxmM4RyXpoq3jFM6GFA4d/nHACTvwaF
WU34P86t7Bar/nwU/ZXODEtqbxf+TWcbxWihHjlZS2GtX/r7er7ob0vkXfhsv6LZqyMTA0OtMIwt
cnNeQ1E23k2IVsjfJqXm0GCaiah/UeyEPD9tCMsJUV96vSrZrKdqe/GXuUsp5n9HPW8fKRD30C70
k024GsI1fVekqlqg0e892ViLy+mbkga/BKpo8Rs3lQmESNu9F0kRchCVG5+W+FXjwYiG5MZWHcaX
gBxleZw91x1OHLCQWQNRLrCl53Npj0JZykxrhhprO0pa3ss10CJR8RfQHdprqGw2lPeafKzpfuZG
J/17q/vgD4XcI3PrYRdoe9GoLgF5mRxnueoh+ZsJv/4WBAL8svMGcc2Q8UFz0ga2Ze07cjEXXnsl
q2ZekKq8tycQJe5hIRpxI/B2df7EtZQfLHV8Roi0uJ48wFOevtNX5bSYLp6SaBWzZOAB6JjeZn+F
sf1DKAGQFDxscJt7MFBWu2rWDREEKjkMMqocuyV9PMdCHWTJY/wFjZiPUT5/QPpjr4DCmtmfSfxn
sSI2MVUG6snIewaAzgMg+2CcGokB+cRklRpiCiEm5gWwrN4Xh/BvSs8zqrmvYumjLg1OLQTeWULR
CchY1iZJHVCU8+QJgg/LRv3nC7h3JZfG+ToKopFCxSXATc9lR+G57WBnZCd5SwkZddiy04HkQDnV
AUGYfP/MUMHvB4PaVyUhgqBw77q/x0tejRKO198wFiXPoPBYE+BrihHcnYZJuT3We2yhNqqWmYtf
fWN8CJuoUGI7TKuZsvyWEgOEj+FsaCKiiclpv4K9bHfaQKiMFJSImcpQC0oIw2/B/ZFoGQI7QJ6O
8ugwJm+SKhVmuML+Z0nZZeMYxlFyg92SpKNd1ADl1cDh50LrZVWVSW/PeUEtYQL5flP3fPPlPkze
KXf93zODPPBKDu9lJ6nDi4AlqVZLoT7RzaqjXMfMKScmsZvzxnpyIgMU815nOMgsZfYsHB3IY9SF
O59go3cGh2msYdFNMHbcjpNkKGEaNMIbGNPS3LYwQ97/NTd9q+fI6UECo6bJIYAc4Ioci0oR0Eym
xq7x9SDA2UU7dYk46U8veK5fAHcP36mgmTIxk2QYZdo2XPyfl3DXw+tcaCcBfg/TqEmKYLWPVmUf
+JxibvxuRLlrogI7KnVaMh6iZnpGiPh1fo6TJk8pU5uir2i9dfm3prx5haZkSedMpAn/A2cpdN83
M2TiNirBazJSUqMDi+chttZ66FlBK8U0lakUDPckwkrcjhz7qMR4YAqM38riyd6EWySmG/TbON7a
79144vhAz0asyluxY4uQC5FDmIYw+j4ib4CL1k8HezZPTUALxiMjDgRkElRrRwEAMYJibtAd3+AE
zIMKP/+3DVo1Cw1n1KgsZRQsFFq27OBE0atqVpcEKPXhGPuZ4rsLqsHX7itPbEpC3DFHii6L1hs9
aGn2k0J6YJhT4uVU6vYHoFOILdvc3OW9ovSTeNiDJ/qwNUyvl0a5m1o7SpqCOOO/h8VpK9RVTuV5
mRl6CB+SuMHBBN4Q+v9ik7X1IaIP3f9taEOVBaUkoBhqzJ0dE1p08mP2cZPETL9X/+N/l0BHifTo
GnsQVxV3b4rSdMyMvY9aBjXMHHv3x3KGjoAkkJlTuUHd72BfvZcc6LXS7K/EXSI54bmuOB/kAUSR
rI1cpFDQhKuSt3SwX4Ar6tQU/ZNpNd5zwRwsod4aXpKIhSuXYot6wRhUjqD1rSIsPEiymZFwwYqc
QQeGpxXeeJZ7BbXipvgjWcezBZkrQEEqdDly9N+ZRhr8oqMIJ3O9U3wOWW9+rU5fc/AhVwWuzg5X
K0DNeuBAzHFgaq+T5bJ4vqVYWGPQygRLEEJaqKe96bTPZRxOYsmlRRNMKyWKYtBMT5jVoZ5Nt7eg
V69qRySmvMrVcceIsTsV1+tdteLn4vm0Jani2Sh6PQMA0bvKGiYhIL7zTLjsZErc+GesXQxF+hUC
I1P5uJnoRHQymmb29SbzOBTBuJpaLLmrUTed1CAWi8hAjxF6aDksgYZWqt79aPyucwlwm3+a/oQa
uTvBzt+XOQURWIMre4wC8KCnfSKwO/Dlo7MikwXcPh8CLpMbxB08QUoIRSPeHw2d1lzbVQW0hHX8
cVQ6XibIFhdPkm0A5k6DUaeWYVw8nZ8iE5s/TD4EFEnKQf8/SDo/QIbQVmbeT5XuqA7AigIF9S/+
zyoXAsnk2IBiVfLfTjgvtCUHXaPhGSE5pGY0GzNZAl+TJcGKEyU1ktVR6F4NQvtwOL1fyqdBJdHY
KXkRYI6g6hTNpiNXCGJ96loU6mZqf0FecZM3J0sbiWbUHDLVSFKQCk0SOgXOXqsKYw3ESHmeLbPx
5qQRTqFezDxFDNCCZsAkRr446+drA9MwszPq9TKGtTF2IS/AJu9wlIuyvlA0r0K9LRrLbh6QFvtO
p7oTYyPgM2iK0KvnR4E8LYkxl8WQACWHDNAspBaKeHzjaDfGQjfGqkDSvk/72I5G55ThrpQ08YEN
ILA2bhBCxCSjmKUxDU8pdnMd68f1bcLvxrLXhb8fLffOFmBwIGe+R885vR19TtW6Sp26inm8J3cz
/s+1E35fBR8HYrXEkPF8Iev3czN/AzxWnHR8XQoUXZ/kgowZ9hUXxVWgmpJ0Fzm+vgIfQ7E1MFOO
S5KwgE9UMetxKFEQHXpjbPeV82Pze9UKg9Dz5eq+w3lXx7s08s3jeGWpDdbnt14FtcC+E/9z6RSX
ZvV+OfJycjoZTKa+W91clJP50ofof8dXbobg18hwYa+MnVnYCo6z8dEcoyD/5h1uR0kOmO/0GFdM
mzDUTBTSKtoBJ83UEkBgC/g+Bgyaoi6alTCWH1t9uv4uNwQ5jLbbW1qG7qpWY4p6HpR4TrR0O+le
EWesY06cIklJdkgPs44w6bQMIFXFleDYmLaIfxxY7vGdi5i8w9bexrTq+BQfYBx+w9Fxiw+KbKuQ
sSZ5DtzdDQwTDFbtuZ4OyWaZaiBIUunABCv2KoMFkchpTlcLTr5eE3YOqufnW3UHTl5DhtMA0Ssc
cRfEMv91Ijuzb9k55RCuIwPTnBvvFxVp0pbGkzhKhET93banxoZWNdhPKvs6x6IyKtNvEIRCrSiN
hlwOCouRYl30PeDVK8YqK6mnjZ9RCmv0IUXnfinufcDcaSZzWF+JSEqyRfU/fiP0zG+xqayNyrMT
isbpM/tRmH0qgkusXMA32ep4WpqNyzxnct/1ZqLdKEAy4HJD8wfUuvZZqBr3YrjyOgd6kFIOxKSO
gusDTwsFYVH9rvQ2op2MSqZxoGO0EpfeY9vp2vGt14hT4jw7A/ItXA+AAG36qsaikSLCs3yJw1cV
LPneCjQwGCYXMwZfpF7t+xJPrGUZO6NHRvqKZBjOvCTOQ+HYVdJvyo72rGvzdviJpSLe83X0ZhBy
BMmxpcvoXkATnSU5gK+KYmtRsT91W91RkrnaQK20ZaUt4N1CWGLmd2U3aEXgiBUNqGGv2fcpSI4L
3M0VVFiR7pn+UAqYFvazqxdKT/nEJ7uG5RDWNg5rO2ch+NmphaBYhJRxm0Ai4f1C3N1uhPV32yYv
UEAus9Y4wCb1e47B+f1EyPA5bq1DQ9RTMXa3gcsm0A1vFsGKUTyJZlUbbSbiQJx3Vxz7rCsto+DE
UXq0x18YiuBjtsI7CS0V+xE1cV8sS+sADQTjprfyLNUPJaRjTXjAhgXcPO2xEY/euHsT4jITzGOF
QZVF3lDFIWwidlwTvZDcog4LoaBI/xdEDaeLpZOqKnH2G7gCgLMWj9A3QPAE+InO3GFv0B2xIn+t
Ei76/yzohjClVmAwv/jo76p/t3NiHfGd8qwUnV9CZuQ2lFy+TMFfYrxMG5MudSALpE5X9O06kraR
nTRWSKRBlMuhp9quMirc9IHOFvLPW9CNHKJIglG5SfZGfnwkQyqejF349Q13Y5uXjQtmp+YzY15/
8D8ETSqI7WOjrsLr1dLOW8Bv+nfwFEfk1494lu+AFNwiUE72MBzzvs6pQCjojhfzTOk/OYdkbkJM
AZBDGRHz0JPA4EgdR1Fv0/VMY5860fKNmH/+mdbe5NO9o8Nl4CWOtCAwTz4ot35hg/CHjIRBfwSe
FpOEY8eQjgmzW7DAmL16eZ0vfHtZL03XB8L5HLqYd8mq0/SwhWvf7lmUSgovi0bMfjmB91kiaosw
t3z8kMnobM+qnBSWb1Qu4deRGAdZ9JiKVjoyOIiSFvursMmwcvjvFw6gVnh3HORiV0nnKEo987UV
CFFk8Oz8SIBVYY3jKoLH3obUwbIpoAMe3k19BOW1BVHMMGfm/R5UMgw54zxwZ39/9bV+/S7DC0bE
IMZo6wkEH46JNfA6YWjKeMPnad7ltTcR9+je0XR7u5ocfJZmiR6oHZAfvqy0E31ltkKeMfd8hIPp
P/LixHmPhrNUOMcaf3jZpCTDpyYPUB9Vd03WalcUkWAMvVLm57IsJw8vUxytkVwJxicDSd8kNLYs
ggC9DU3vnZ0dzp4fupEbotUDnI7/FcRmoEK4GUviHxdPzdisW48b4S1iyrLcAVna1WRPetso5WVK
MMmUL2feoUpxspb0JZqxFq7sXnmvgolSF6O3FbIBwQABBmQ8XY/H+2rhyKlReuflbPZ5Wtr6sxXd
Uq1yvKk2VibT3v+5ZNGNGcTrjKZ1E9ORezIlN0ftYDQhW0KF5x2yBi0S+0TGoaO85DkPNqLtvasL
3LWCLmoyTiaLEWwdUqDJQXhZI5m8SzI4hcD6mF0nKJzW9ASoAaPkzwxMQe986ZjAm9uqF5D/285J
5IEskEkjsa43jY/zqCCLCvnfnjEgNSJzbRj6i/pkLjK5DwtGDvgmtXfcl0UwDEHGWdWNjO70M9wV
SZz9LyAGYrBMQn+GDCzazCj65Kn9nYOHjk341ihI478KNM6fNHBaOvB09v9aBvOxLYDBLb6kKtsJ
EH40KEvbJl4Kkscy1UbTKxaQWFDJikarBMuQDbmabfKZslIYkCOVJjIqIrriY7K8GAPwwFpRISn1
J0i/xs12+bgIWdEi+27bo1qTtyiiEfrH+3qLodKBcb2j2QF3PM+d8A+LPD/eqYwfyJZacPYF16qb
MX2okDZEQC9Hsg/pZZJQ6ZausSuZuA5WDoKMMcIwOG1gHaRLg4Ply3U4/2zeVLQ6nPIV98dxaV/G
zYkfGKwfixTScWXTAgUmEG2aVdnqBaBEUHQvbtgFdQUcuzuc8CYkgmdz+I6tH1cZRSFgPSLHZduI
NOJvtia+rVpeK8CzJdhNUMxJRv7yzGtL4eBo0fpk1tPkMpngDum79DUhdeWpdxciFcnnyCUGiEKE
tHnfniAFI09lqgxzGV6Bq81TNbcJqDHCTOjB4fip0n28HvKHVuAMVCWl3pduyjJ2jOfNHNl3J2Yg
J+TpINBvzWhovV8VQ/QbAFjqT5NntPtiK2gTPGhvXIdhryqxljXln+SeNqyEG66n/sKQuBOVUCx3
hPixvff8WLlSrfRpspswqHjR+Kd9ClsTe78FrmbplQ7mNJ68LDfa/3p0LGrhoSwJcOSxJDGYmyfi
JgfDZXa71BAx8y2RL9AgwthISC6UUgWhcgUKAEKqgYlTOwn+etKXzCjreirtLjeSGz9QgLfb+hr8
7eM9CZiMTwGePrnbG+V/v6k8JY9aIxYfjZ1q1LtKdHF6prdlLQ3pRCMC8uGHnDmBCjj8tflt+Gk5
I5ENpA5N+KWZ3Wftj5PbBhhZ9shwyGnhHnPb3WtH//Ihu5eCWfQ4n2heMlsTFiIggr0AxtWw9heB
Jh+lbH3CY/SP9E5PPZx8c5UZdjZJ5JSuaDltsu4r/nGCivbLJBTRR5bbD9+I1KVTJZRzNmKoxs9B
DR0BJ/G+kfMSxHoj0r46xol4E5XbtbUDy38sqm+OMqari102CJ4Uxu62IgiZ2AxOOV9/N8Af/xSd
JmYCCwDGW/qEIZ3zZh5/a4K09nM2rSkLd/As9MxrAqPjfSTXTaIErdxAI4bDsDwOyx++NMONqaZH
X90L1BnbupCY7cLHcsiFEJtgV8qBVwivxiM7Nd3doo3OZkNKktGlnZCqmZGUX7dHIW+tdR7kJncd
PI6b4pi52O4ynSMs0tYMXeu1pLFHymtKI24M6PzJdcJ/MMRg177xSrib/AcVhLPZhJeojZv4eaMx
KmI86SuGqrRN4XKzfzZh7anyjoOkmDlw+8qWddiLLmVWqRyBSxAUarOsGL+p80wJNJKf/xISt12O
YNCOa4jqd0qM/oIFinNl8SQpqBK8LU8PoQnIk4b6IIcLka1jLGL+59M0fvNwygqypm1ZoIEsuJjW
Ot1IE7LRggrv9zAzIqym+YvmSkpQVl1zSmZ41gYZ/qzAWGlK1AbC/vJxVwKKDsbIkFc3JIwAzXvK
b30od55KMMmVZmhGtkrIW96IhkzQl3Ql41QuJ/JXI9xM2mWsLqc0l67TScurxr5eZBGd7iuNOhTH
3hyhbi35aSni8313icEnrAr9tPDhirewOnqXExXP4RqLb8KWYFiKrA3uLxSxrjQBWKCqhNJPBKev
Ulze5NtKsBoAjdg3vtAypSFfaYNxFKAXouWvqF56QwTpdNc4qcuufvrafrW483nCTcpn3hRgcQo2
2/OfSonyj+6JxkXkVPBtstqZeurHFUk1sbS30ohCZpZCwz8tBMFOKeq1vO3E8X3xnxWC5HFslmiC
wA2UyHYH38wTjTTxAE+QRahXqDZPLgfhz1Yr6xTr7rD+upwekUFxIS9/Kmbp0YEgXHMdK3TqdWtb
DaRfm/MudPvI+xO993T23eTHfFwm5ab6AxRhnMuPWgLe9ZyjkHEIHpNAIPgpSD2VYSk/DY+izrgN
3rl6quHL4Tuuzivin3xQV4a6vmsRqUkI9pOnv4bg4ZTIrk0Dx2xto5PxHsauNS751TXavcIgf/F9
stBU90j844JQrvrqxKoqMVZAzlRoGLZ7MzyM9sy6YCLzIfB9ybepcZU2G4m7xZwHRR5uIpEFESmr
2a/NGYR1bw42cpfBjb/Diu3pmnjKh+ZSOCBppkVUWcPl1QVixN6KUld1Jd5ZgXUWbsD0GjmEJAL4
J3oZM1AvOBS+R3bURGiRrMrx6WysvpFdsd0DX6QBz1HNBsVqdxpKvxDl5wd6Wg79An7mU6JpkQPY
796ItaWLxpaL8acvxeO6RENGOpnj7C9ib29BNANpAFmsM6sByBFOcx5d2zWU96uyk6eyaEb+7NMt
/xvOoyMbKZL7kiQeUF6H+ebvYFYz+45egSn6w2a0sS8Cbe4Lf1zBOmKx7qgJIWgIaq16SK2SmK9Y
Ui2UMhhM3teJ0YTym+uei3FbGOFVxwDZieHgukAFyJXQ0cvcNalZjg3zhwuTrGMOV97eHDxjknnA
hf2k0w6x2ojlx11QQL7GzWErro+UTkpJkxrTLetVpIwAElxrB0drsCHwvpKJOsG+ki2DFcsooItb
0ZMGz/9PDcop/WdeawLmQ4ShUT5a18oKygOf/szMSqJxQSEBzS2eAmS1DC+E4zQlld9ZhusV+48x
hPzJkXOcS11mcPd39j0IZKSXCquuGQw8JoG3dq6NUY6cEI3qeuCZ7qGSjYmzeAJsZmQF1qT+yWep
XVSju/EgikK6r9akjXpp312XTfY3DYYUUcgjI0g+kfqxCWAod4fBZzu7Q/W3Glxyp+//wfw3juU9
pBUYqY9qzJGs5Ouu4KdESk9+f9jSesoykTqOErmWrq+kdfInKghENbACFz0LGFuU1Jipbd/Ltc8W
6W1c6+YfeWYop8tZje8iC3SKpc/gKQnQzbN6DhNhruPpYwYhCt1gbDwl41gEcQ+FUklrf+tqPcq+
jvs07QoDjyTCd2aMbedfsA+BL4OL/umxbOmSJsjY35b7xv+2rLPx+LhfwN1aafYTXBjTb5TW+Vux
/tk1cy5teDTMeH+GuyjOvTlV5P2S1vIUxICiA99WoIk1qOB3lQBse4yIYHCxcQkUMKXs5/VdJS+8
CxeWBNKvGkETkOfSGs5W73GvSbheqgCw7eKE+FM4bNHUyfLcJYEQHOgooY5wx07kxY2tPOByfYtT
9kyd4jPOmFAr4pEugFdJ2MD7jqjhnPZKGVG2Xw6/bMJaLQAAAV5ite7H+PgKfVBQwE6ZykQcGI+E
QYrbHWRlvg5bGuyDXTvxXktpDmdyjrtZMb8D6gt/ygnyAD5g/tv6RA4T7yKlub/PU6wXTgMMa1eB
td2poQ/PYfELxyWvBtegSWWDT4vq02Ig7agXiCKHi9EZ+pt6WxkXKdof0jEVlowkWgFBq2JlcgMG
ERQ/5VZBRfr1odxWjFKRqqOziE4As/kc7oUJm2VL7Yz8Baxc75Em5O8lC7QDQhaBVdDGzzzTPt0H
K+rUfFRv+bbq21c8zNsMiwA0rsTYlXZY/kmcovCl5oN9C9ZfmhUvRDGCzxZKrfA+NDd/YMkAqlEi
QErdS3+EzQzmKN/Rq0W17gdALhECSdGuf0Jgu9gF4ga0N6s9Ar9e1gWujspz78Q5x9YqSv2TX3IF
ZiwWuwRy/ZY9iC7FCf3mQTSz6i+sJ+SWN+/TunJeE1wqTi1V+AX1JUdlXxcvowk70H8z/gtI8T6V
0TWJDd6/0uFmS+ZhDIQiGLJCcbo3xQuUaiApsRNGMRptvmpuifTA8DGAO+qhGvqIT/II9kYDrOwF
RAWiVGc3jrlnf3UsreZM+JhEQtfiQAd9dhl1s27HDsYp3rxFHSl/Spk+iNcqMQkgHRC4OoF4knB7
4sf19zQLyVfWQ8glGl50GRnlwqOgLNfQZn8DN1flh0oPlEKYoUIJZRDAtuSofbI/ABPQqCiWB2Vo
38tdvqCpirItfgv6byoAtFAx6EvMYD/vE6HAPObZYu+NH9GPdXxHyuM+WlKHTMdXZ6Vms2Wgvh3S
GU4NmQvy2/pcdVEs7bVAbQHk/Te0u2BFO0Hs5fHeDX1WXr7479BdJ86bxwj5pVS99SVyovr30oTA
G3wgKsLA6Agytr8wzYMdCy/kcjLad0KvL4f9QaNaNUsFAF5erTZQV53oShSKx4akyQZgprW9A1Da
246EgCUZRuBRnn7FMzUFdnSu/5Fo3PD/ju2i/wl8OsA69ba2FZqr/nQ0v3l9Ecn8fEutDZWCUa3l
mFuI9OodqhRK8/tiIVWVbBzoHjKL3yDx2OJSpgXrDNpWhTOBHA4e69zDk1EKALTqnYZURoZEkEqw
AId1EHrLpbGQpnu7MHAU8yv4Rtk8PofS61OOi6PKXMCS5CmHAxlwLPiDfhjvnlcAK58YkqYKLRzk
XlOQ5XtOu6U9BOMg7w3XS8hkpnwGM3OVbvtOAeYKYMTOIywAhEeGY2S+tv4TurT12hLoH024coHb
c8D90nOAhaDAZGm3hRyYsawN5wPUB5ZtiHlt8CRfg+K843RBauphG/UX7p8gBPrRvISZP6ZMhiqq
69voRCFzUxdL2158eyh4HJZ4XI1ZDKcSqMmb27CYB8/QU/KShZ45HJq5W921Rm3PLX3vN/0HAQWE
Yooomakcb8hsJPxdiq7G6YkPS6v8aiKvK9YacKQQs6HVn80eEvOM8eJfF3JnQpe+7B1ShlQP+9o/
z2zB1ZGM+Xjhu3tdXi6YnhxO07uLKzp2RXFaK8OxpIpw1B7g+XWm1ShBVYXSl1rOBBcdU39Qwhts
TuxEOoOpxyOpnIib6clO5f+TwKtXTHa1LY0NIoR3iLAjjtkljAzA2XzMB6fAPkA7lQBlIDGSRv3J
Ti+n1XWjM/0sQS9pHGHft1rLW1j1T0OEuF6kIx2EvhK85fthm76kpsqENQufygF8kHw4aYKWrlKz
E2eCSGCAlkHWUKNb7cIU5cSqwdAx/8TZUX9VjrOt49jun8qfQsAwhwrnDR8huQ6ciVBiikPnThcn
SFdKdNgwZAI5rHXOCEtlQx1JOoLAeXFdGCCzAD0IHrw5mNVKObsvWf82MiMQ8q8cI6Y+UEBNm617
3j4eNxby91DiIKjYVkI7BSIUrQmi6UyVFXyNXXgLpjsMvsW3MVWFVkrmRzujBaMdaORhBEmYbuDG
rvR8z4REGPh////w/Xco1IZRpgvvLb+yIoYkYQgyCkR/53kyna7e8MUvWjeHQDV/Xm9l/dTLxScm
++KiiSRiyRE7nd/P/SHxpZ4qpTT0N1SjecSTGeYjR7zI3rqUB46f8ePub5x480GvKH4NpMw59x4O
VR9AEnZNvCnToxjOlVNPzh3txl6jSxONFyRsuP+VJSwuvNqCdSnJUVwrgJQBJJc1PqLYLuijL5Z1
cQf29REBbqa8wqcTEOF8ZFQejAo5Hro7/3tiPvTUHoeiKRKeUm4QLrghuEXesNPLPOiGfw7BaQbL
x35Lir5X1jGUPMfngxPvKEAB8YCh7QnPob97pg1wieD2iu7JBiT0EiDpEWBoW+GvPMPrVVFkRlwH
MidF4JFMzjy0eRH2+kykNoA4oE0VnXFWAc/8qmH4Q657fjgex7bfmcC2Ub5nVcB/G+afm2kSESOP
XVQSg03rWZuToAEDe+7Fc+iVHxHhJnVZraRYB7Ybo5KK+jfYree1kpKBugRa1/HBZ9JGfu9RrJxh
EoDOHX9vLU3GlIPaXquoxaS1q74dyzEmnJHdAsl4kgpHqXrdzF0DFKe99Sv+78y0smBJ7vbHQOO1
BlZn4KMtOzQ6dNqIwMwNDMSGVRq/NgnWX5offx/k8RQ3jeGbMylXaLhPE8BFnRGma+B0zkS296f6
qAdO8p/sAfJ2hAL2qtD5U44A9P9l8uqpBq6iplYJLU9/OP88go2Se0wOPAnJMA9qjjWcwcrRME29
cuHWDhjWWkDPYljM0DbLeWnAr/oLxcPWxmfHpwkVPTXRYX+jMdqJSKqN+qFsfmAv2wYLvUhcF28l
s/0nKV08MihPWUFiYHtjI4A+Hq5cl0QcDxBrXWe8Ag8a1vpqFy4/BHEeFOKtQAWuuamg15OD4oxC
ktGgKu19k39p6oWAdiS/kSceREk6rB0V4gCEwb6rNRoboABqSHVqqgHTjJqMbQ5IF/1imJjlCty1
EC1k4ZmKp3XAxW1MOxZKTvKtCDcZ2jsvWTHXboMAdQgCFLVwL3MgrHuibPjPFF7XVTfr703f1M3A
4lV0/KI2S9faxj2/R7qhq4fUxIqu0HQUT6TIuuC5brxxAFSWmRYbWre9R1U7/8KfXt3C8Z8SZDUi
dwwBL031Zhqb4m3AX8h36Ncr7LMwP3JTRiyni7sTh8bJiDqAAymNwneTcaHqkVzb4CwDrRalzZHu
8QtBOQXogqv+tNYhum9tWRHqgDrh4z610aWpMdAb+p8+8FB1q8NVNlwI/c6rojG/zKPezT2ibROp
cZB/ZYmObZY/Dkc3UbMqE9Dn6xVAkhBZ9bzBbKBILFbj7gtQIDW8MJL4oja6Nolq2R7GnRa+fzfl
TPIxPvm3oCf/p6AvZTMG+WQcF7k36DN0QOxgdI6mBXqNMIQglWi22HOKbJe7/3jggCPhcY7ML0Zc
/3DZidImvRi/Sr1WmwKRRoKdE1EzmGjx1R05iAx+bgUAQCADisaIBl7jHqgSnMolt6JuUnvhblgF
YlGb6qZeDHvA9Gj96V0wN+SOhFH43U7a9UoyKHnAqZvj9k4PAC2d+7buuAlSVA5pedTHc+JYVPzV
9aXW/DmVIUgZ0D0QzVVEgn/4a1TiAJCC7apsmXD2tn9GsYC+lt9CzLP8/FrTg72SgISCT2Kwqyqk
yeD8GRt7zaQZCgcKcXUyn5WwwmLCCkB4FbPvuBz2oQA6gfnzKcEYwYDmllqUZaYhiOKw6q9ABD5+
2EuFSxZ0v/9m5Lw+B/2cboPnjxyqw1mDGlSRXTE26n0qWOr3w3uyVyy/aBoOqL4/OXVv+G/BlBPr
W/QBOLF3zeZ8qiKCISTa+rpdgH5UEVZT8uS4H5FiPh3aeaEat+ZIgBu/RJW9XbRm9ZICVA0O56x9
mixI0rLKRizM2fN8evYRSJ2dzNOz/TH4Ebc7lSALe2bFnfIgyCQkgDZ6XJfUrsCozsaoeqBkBZNe
5/3QNCjehrZkskvK8R3Jy+4zQmmAIED5WmGL5MC8SGVSv4/DbhU675uPf1EBciV8UxsRayfij5m3
FcfnSSvWXzYxqzp30TbzLBPx/XT+tDqtzQ+vU/62Q1RXqDrshwI7qSTDusT+CF0wjSSOZ/tXdtEi
Zm1E2XWCvV58XC91tJdaMlHkDXOtU/egmCuNnTbdmcArGwQPePGZf5aI5Fxj/YdG56mKrOxvorBS
Pguig5ZjoxJUIMCTAHqhfZ+JR7QALYZj4auChwXNmNxwGa8PTbmyZ6jxo/718q3HN6IwESMtVTos
/XbTG60LhyJvz/140A98YP5CogdGHSElHwQ7zR+tUHkv7zpZ1iNn2iVJRC5qwp8L0/9TVe76Mgqi
I/bo5866QlQyWtHfGjQ+U/suYUP5m1FuEcFXVqhnVmN8eG04njtGFUod//LIT/MALB279uLPfkpL
Mn5eULzE2pAsSiFk4GghLuOdK5cmVbytuEby5eMh1sCVsoVWA7+AcVc77cq77Rrs7JQRGMzUZNbx
qX0OPyvhFyihkFLAwkUm8KZE1g5+EFAramIn00cidSccF7bVkJQ739mV0iOVDikMBRCUCHY2qPLj
8bIkGi2jZHSBMqfM1puJhr99Q5Qoxf2r7I3tKW7KA0K1oa0ZzitBoMMbEzpnjm1eQdN2kgL/Ob3Y
fv7otUH28mlxzZoEVnKzN6fMGTwQb28lJWp/u2ng7IW7NlAL1n5yqt7ymYCFbtdaBy0XJh4pno85
G/xszC1Gje4NDFxbzxHOQUv3PDaqQG+tMDxaHzbWM4zoaor3So4v77x3nZLLBH3EO+LAiQTg4ZvC
Cep9UqmIxGELiAzbLh6Vr8p6qN4a8YvLCj56rFxwsdca1y3zN+7t7Ax13kT7V04w9FEAXha3tpYs
c/8x5LkyyWMPUizzpqLBzqilon86Q+JWXu44+O0kcB3BSEswP/tjWrTCvqSNhQulDw/5fSWyVWud
g3AM3NkSZzCEjKDsRz49XNGPqyDDrpDSYufMP+EBzWzkGUF4bKgG3b6RKQA9V7g6QHrQSmkvWluS
J11TM5sF1AaDsXbvk5JxtenLKI4Pp4f/ZqcYJ5JumcqsFHjq0JbvAytdo4J8wZ2i8blVN2U4jJ7o
KdjhXjd4fWwo4zvgR+TS2Kqh8WNBJsgDm1IvpOApUhwqqucqEKCzLguFacvNaY1CB6XcHmSUClLd
0TwC27vuFSFoJnHqrh7xnZFmPsO7ZzTIl8YaP+00zHgQkhG/lGT96LD5G50xijqu5SjRhKHaoeap
xQ0xJ7NyvtswMTSc5cZVumUJgKtXc8osJUU02ge5ypC9L5o20JDxzLLB5OjhTRkCtUgs/ES2cnst
afgHqyXdwbUilSrxWtntNPQHqH+PD0se84eNiIDgOMTUylY0yc0QWF7zH4X3tMIGXhmNam38bvl7
UQ2JjQ43dWoYoyO+pOcJzy0gt11oCSLKbaHj3wyx9PeF2khvj98t5q5gppvA++VX50rxkX3NMK1u
z0h8IxpePMOuqOPDPu+omB+Q3l1JDaDrc2Zv+Iv7XtgmGhraOuig/o2eG4yh8g5tNeboDSfVZdnO
fQwwurIHOVvZZXU9yTQx7OMa1AHCd+yllL0evvCQucXW27bS9UNMjG8JXJ4M0qiYk9ho+sHRbc7f
107Cvjb79+lCLzY9vdgz1uE8IB126p1bEUBHR3m+48JxttDyXteRVGxDSdTOIzP/YoChTX8EtUpR
tgmXo80riFSXJpEpJz7/6qBX5Vvk6OGIKrtweiqQXGWXoeP2GYKm0f78W/GxI/69jqgWM2X/eFVM
gyv4U/P8CGdRDTQbgxh06IklYvRU8ul4c6ByvAkipsGasQAahEAFG/np4tEgpuK24VMkI9lf6mfR
crS2JZj9EQ8ViH5ASiEoruD1t7CDeMAhZv5UwrC6WZPmNYHV+QgSvE7WP0+pOZWBaZjE3esKBQXL
pFP6vJoPUPoADHqKV4l8QECU6AhTrfDuHp/SYIJNU4+8FjrYKB7yiLyRFnIdFiG2Dm3scROm0nL0
hfMtl5m4lizLUEybwh513mD8x0JWaotVP/PGxSKxnIy4hwXVenRd6CE8b/5FdYbdupBtjIiKylZo
Hb5mblNk/GtdZb3hmUJAlB4aSM5EUfAxAiSr24Zyn0SBm82U8qztzcdHjmcexJOh2A+KCeIDJZ11
XW1KvUOfPKofjuR41zItgvmkiCmJ8H26tlzaTeZ0Pwl1LDRlG4gWHrjGQVV9XMIXsbdJdq5lkEaw
uUy6S6gR6oD24n/ZRiAYQt+FVnloILZseYNqJs7KrozRSxgiPHY9SKjUemk3UrUkKiPg3VQmoPYY
26FQNVbHcFKDn9GB3HBmFLwTiX/JYL2U+h4mfyesBEN6IH2GnebgtoqUbmy3To1tU9/ai9Q0s0bc
8hf7RvKQjVxrQjYtRrr68Zh/vZiSCLMG295YF5zksdj9V+K3OsUbc3WgWUSNFBuvV9+7aZmg157t
Wd9MRf8LNLrMq0pT5A76Wqx47qasNh4ipxGCHwgWDX0mSiBl76gyhX/CUbmY3p3xxG1ON1t0hGPg
4Qf3JhZbg+7dR259HkKvPa0CcB1u715KxPwnoVDmc2OedJiHMZ1nHUSVdTiXgGj0B0vVHmf/aT4P
zk36h8VrJuQMrEuWc3S0O+/BFjP+5ET6aBqI3GgRlzkrXFlAGr/Cl+fk945HnSfJAkS3SbgFm0ty
jzdgnRRx7LeUayZus84xT/l5ZywIK1O+jlso0bhZAQ28AeDIHpdCFLpqpNvEjLqSVzZickZEImAw
4EzxfRUGaid9GtTMHkJ9n3bx14TeXjUlCgfSd3+SMMsAvAkwhsJa1dT/nroS9e/3iCCIGUipp9Zt
FDDRgTxsTEpCVpL8IQ1REiCvU51tCo5rhLWVmky9j355a8VCqkO3OqFppQIsPnP3JH9p84Q3C7mX
RI4sipfYXmkSZiujFF5lmCuNk8yjlm1ciedWPDgi2KnmC2kOW+rfuAtRE1PlBsnkGVdImeUJQ3Xd
ra0alSypqkGqSb+rViyqIH9Mz2e/I/2v145F0isFR7yX2IL0UTBh5bBVcd8wAOC/sRzi80MDUI1m
doWKGl7shinQVu2kWG4D32piPH5oNrjp4yXAGc8g1VoPXbq7XbY6afROTHxSIblF3gi36ttkQN71
5/JAAJrQuJZKI7tjQpENypDSCAAkC++2ztQ6dLo6l+TPRHixcGsCNX5L4zQTkJieobTMTSBPTv0f
XKzQIJKS6IH2CmOsD98TodwvVvjFeiUoCyvHpI39gKbmrGyKq7nPP+4FpOWYxH1kHjWP2q4zzJwm
nLy7nw64YxklFiap4+/sblxkmfmq4tpqdADc/ei/+9ox8LhK47oLGzgaPsOdnah1GOQ6A1q7oGwy
ssYoMN7mI7El9mETBJRTWNHe6J6MJZMXnOZCcelOorLOko5rDTJ+4XfKFJDKNOPHXIHbaOC61pBH
MLPo1xH3sZHdHY45gRV+LWrEC7fgqn56hyLq+OrXoIk8zmx4p4ODm6EL1NqEz4wTMBsxWTdc6Xhb
NyW7vw6hJz1vv27vrmcOi+Oj4T+YVHCOL1TOwTzNMiJimSdChOGKzVWqy9tN74KNGNtP2qR3l9b3
PbFzaRB+r6vsc+8n/TIkvwvGnFK8dRmAF8hj/9YA4FxsWEBrj+FMjxpRdrR0kiSAWYtoQO7B6Cdg
V2SZqdawhkTxbrX7a1mIIvY3VDbhf2m9GFyD7tjX6+YLoc7P6SOPfuC4x8f0WayOGA3/7YyGFtWV
55q8BWwi2hw/ma4cFttwaQMXU8mBJbG3Ne8VXcK46yJEwn7GU1oHxO9WfY3jJs3QpLUtArT7ttWS
sNI7OYnpBqmjpOM3+VMJYyk1i6D9aQjVg3x9P6Rw0TBoxr9Luhjg+JBEIg37Gxy3832lb1sjbmqi
lBcLEiqboZvMYZ7sKCvCFvrmMKaCxb2FtPwt7+2S/kkNtK3SUT/VLpiBvYmBI/xEM4tHCXSjLXhd
qiecvXTzM9fDfAu4pL0SuqH5BgsvCLVjle4Lyb0NhPIDT0PDmbgEeVKUDccbO+pwZ+JtUiBLg7Ga
/PqTNVG4bYlMS2UEyZURhWPyetEZC6UyRXfdoTXy2el+OT1d0WOijkHinMY9f1ZYfAhBb3vtKrMK
lyFpGpa/OlvL4DVSH1btF1POm82ncwUfk7CsQvbAQmMs+TIJJMZPwU/zLigw07sqrWLIzFD1ajd2
H0tYcDiqkwCDjavp+i8jSC160EA3mdxbvSyBdok68IVyuCrFItyRp0mVYd4zFXirkw+VglrCUz+1
5h7X6IoYR/NYBVJ3XwPNbR5tkY0vuce8tcGxRdRzOjauL6anQhYW9mFHyYH7O0H18DXv/+ShIU5C
QyrImttrPVdfx3T02Iv2cneKH2d6iKeq0HYMf+DVHnCOWV9LgyFzY45pOtIzZhEQFT/giOq3RqEB
6aF7m2KaztPOl7Dwy20PsISx5syAOVeAF19p9hD86Lcz9BVQ5GPzbUCyNa9nJlw+XlWLNFXic4BN
p6XN7YkUd8QsJQNP+1TfH5aeIpJ1t1bc2Evd6kKHC6Dv4GoAnmRPyNcOrBZAyxDR9dHQzbcJg5OV
8dBTA+9WAsU/7lqvzj/UNh1ibwElfx22vr7M71BG91YsZozjK6ibrfbii6bpamJzREnqTSAgN3vR
omqyPvm2TbNaXejjLazSn0p4Ku49Ao65VNQvakaQL8pmyrlnTrFba0JURAFJfJLWDUc9WQMi2Zys
XCz2R0TbOXgTtuYeJqpGPVqo+WkazXvvQNFj4m8qfh4MLqycd2ditSnRlYU4gmPpcDl/G3ty+EpP
kzD9NaQS0V7034SyNzTDtfGU9yJ1DL0podQZBhrruR6McJF4cSZcK83E0MyTAbF6owSX5qIsPRmb
pgh3pPE1fLdnQN0wX07DBanEfbGk/7WgjXTZtV4c/PvVuVg3zCaNEJIBuzgjj6vkfhxpzG31CdvA
bH3nlFuOqahrHROHlb3TMrmQIC9YoW/u9FlJQEuqafzyA27EvamA+VVye9mJD6ITwE8bLOhJJxYM
uKzDMMM6KIToV3v0GVqBs1o1ji5nn7PJkrO8dZI2zqohYzMHDPK7l92xpJBje1lUFGCHvLnWYr57
I6eS1iUH9qnxNKHc9IqV1jKRcMQMH7u7RZhOhEZIvex18lJIGMILxZXliDyzVgAPcbWXh923ZvBj
DcvJyOgzl3Bq2X+7seD5OyBnfEp6cg6jZ/aRUpaPn+59geKlo+8Ln2eP6Oxygl8p9c4tl4aYBefi
YkpfD0X4x5ISyp//LvF4+DV2162G0ywwomeoRmHR/bEFN7s5zB9quRYLEh0eDa7ZyBbIbK6uAq67
jIWCU2ySj+TypFCvSVIazzA8XrbLLiNeDq14oaPrCh7/ZAa/UiOCmuPfBgWKEeNYRrTrmeDlX7bf
qY7KNIaAiiy+VhkGMlW2fb4bjVjMFU4wHl0IM4P0GwJEl8tel6lnXx2IK4gxjvVoxlpiRRlw+mii
aGU7MhOGhFbDIG2KKIw7GG20a/YZBrx/hKvxKS7eQ04c7YkrZ0mDde2RKkGDH3kLMtxc+fWO54Mt
XLEQVODHPRMw4xXHLXctFU+DmMrDVCd6FtZWTpVLNl3ygu44SUxlSqybgh7qoiFoEWopsqdtlxtu
MSu6pc/OGFvmpCQFmG9XVTHzzmc5VhJmA+c41aMOE9F50TFPZ2ARlZt6dqLftl7afzcp+IZSzE5J
F2dt/UIOfMDJSG0WOlzdGJSvYNaXQI799y4wiqGKBgzlpb6RBYprRcRwjHIKge7JVFWBZejFvLkp
DD5hyDT1KBkH7wDFBGypQSAx6S+m0J1gAGSPh6LWW0bfWVcFHCvbpI9Q+JY+Sc7+MS5tAXOQBxWv
aHeUbaCnQ7b6V1XKyRge8RhtygIuBZcvJc3x3gSHWgKY19NAoGBlSd0UJRV4rckcN4c7FDwOIYVB
0B1Be73jcdh8htck86dwUM5XiAmh5mklQP9CZFPCXakvFpw/nIwzDg3mIhIHW42xJo9dqDHuzuop
DIpTb7jnT3mBhM1DhZvSkFzlcEp2PoWfwuQKIb3TQuTY5ZCmtXwzWZ1QH1nnU/hjLJRbns0/B18j
WKPLjhwqtghBpFKiaO8hOJlRFQLuuX8YnM6h4V0ZbEBcBwE/hXbfT5t1FWsL7yWWMI03tT9XichK
iSlNxv7nuLK0q9dMmaKZIvpgM6YxRMVAccdgSRzPrx0YiPzzTuCmePahQsdHiqpGUIqlyDs2g0I3
ftP0WKJF/JdtmvaIBfevrBeldIVRAQmZV9fAvHBd0pzz2CEmYpyuNWk4PfWkPSsxum8kXteIsbeK
oUfcIRV5JpYUgd4tLBoxTvDgp/ibqgV9x0KfaaI1LuUP/0lN4onuNe9EZ6M4gS1awZTaRWetIbE4
8261hLiOOOsumStA7qASsxCL6vMspcJ+mhIETjA6D2sfV/STfl/rbihrLS9iROsfjK2wXHGzSTEz
risOKSS+2sj3xy6cWK5gHaXxSMxxGYaZsoooYwgcfOqSyKMDutl/tf0FnS1Oh7KTaLQ1EveHOKw4
iCyV4mgmmdY3/0I1qTEwFpMeJZkfwj7/3mckXshE7/aDmXlMZnm6yed6YrmC2XVOHOHwxZU6mK3d
Sny36jLx9hlI0MWXn5NCtzs/XZhqHYfuUUoJNS0S6Rz0XgVYM1zyyoapi+hFzI31OwHeOZQNhzZ2
qOxXHq9QyAUGOeH5KpGhzAXuFPeAl73QqsjfTy5BXzxRWEq0U7EZty/7/7dAOG55pYzjmMMsR0VQ
g+pj1ijFJFgEwp9aQjOl8A/8+CkrUVmDuNoZtUwSg4j6ka2nAcVbLf3+D4dJt/hkl8yCblB4PBrX
Sd++gCy+JMKTvM0/ZRfEoJZbMlh/6kjNAoDi15RKxy7Tu1VtDPAlPSHf98aT/RIrVV0mcpIPapSC
MVI5vzByNKK4F9MOpQN+aFf3eHJHHMeQiWX5TdzzZWxA+Wpd6cBHDosXfaGTrxv7B1rTH3OhaBaW
A9z525qAUZpP/mag/OnW5J28GxsbT7BgmrxGEbaXLLuIm5c6D4cUqeREmwDxa52CFuE7hmwhlAMy
EkMU/oqiKGQsBfId9A851e0QqqLOx1Sp883VZfnUwGOMLpopVcReeGetghbmnJYRf16Tgu1GyUst
uVD+yJY5fyU0HFpQ9oijiGso1pmKAXwX7BNthRWUkRZrylfa0j8fBxH3z88u6zDuETPVZB5JitXY
+aVXdQN3eB8X9ZORXMj17l/XmIrofb5hNze9a68e3zApMkMg5Q7FDjDpqTqDS61e3KuGKT920FLU
UKI3D83lgf5oLSrpW/DheYkK1qEYRDVXRYU84/G4x5on1T3GmHiWBlUwvFxViCO6iPyfBuqt1pkL
9GYJ5S/R3BLPgi3SUPZLPoHcbIdunGXj59P+CaiR75dUiQ3N/3RqFfRltDa4odHsfSyElyJverD1
X7oVyhPGBTeSTlhMtYcNxMjwlK2pMx9fICemO/DDeJzKEkgjvXP2tVNEmO4tZ5Sj+DXJU/Vg4tuQ
13deZQe0fIZhwj/lcjLU6DftfLvfdl+ZovNn86dJlBe8GWJtXaN+vDf7ka+vekcdVrSlOrcI0a/l
x0WLpiZyq5v/039ExgUFS8i6SQVjj4whCIm4Ee/4lV458IgvGNnbVmEuuvyKg5TUIbyG1Pc49vQo
AWyTdMFtoC7HPkdspP8uv8TGJzprpZhsabMi9B4jyuyKedGP5MfarfmjwJxgZds/jbAXDb0J0bdq
H9rq89Er4kzoi1oIGHOPtmUoTYUkPVk+Z/U5neovPPzRtgINrLTuD9dOoRLfdDcMbASeFnD4gjxl
XmKG8KnSIaN4qZxdKqtxKe/hTe5HRmWK4jFN6JyYS2Up6Nt5MT4WuDSEnbimx7Qykn93cw8G/Mbo
ejL9oDWIc6fyPudNnotQW7L0p19YHwNLkfCC7IHVXsuH1FdwzVkxC7VOhaA53QcMFmbLFJmLW9V1
ue76EqFujVkPIagBprPn1eMxB4mXop5qET5vbYG65CAELaiIs5FPxGAQNutAW0+iVqDIJtlD5HBy
YN0IHpQ3+h1DctG4RpU4u5LWuStFBBt76oknZn3Tfq8tBzdtsFxpCbzYREHflO9VIyH1ftdXaKCm
f/N7Pjp/KbR9AnmWkl4Fo/fwTYK8u22RIjhOSODp1tpim4yOmeqKWFRqR1IV17DFlstLWecN7mSM
ZvstK1EtQc+5pNBZn9gWAGmcsKacI3eGCibjbKt1+t7qge3icZGUlUCDq/9w9l7t6pHKsMg8LqJf
ZL4XUYHfxcEmkL6n/lq+OBo2I0yOA+wNDIzULnOKcDaGqTJpRklf0NIq1AJKVrPlA5QkpTsLzq0b
XyKX6IOMXsc5kzMHjZEUrVvCTR+WX4wCrxy4pY/hz1we7GAnIp4CN1TRj8dmRXGHQmH1cMDrrE/v
Db5o6WXK4oL1DaBSuByy5nDE591OV/NgcYAy1HlUrt0gVWKJCTs0F2CYwshKvLvuVnFjxWcGm4HH
RpGPjHvIv+/1k+usMvFCJkVAUPoqn7CTFoPIgSf/dq1xdnuo3h5vQ1Ew16wmp/3C/fNlqm1Uh4nq
AmwufQ7RdYv4eYfSZb4bAnQbF9Nux7FSX8W2XJaUkS809779JuzIdkaSseT0kxZ23p4uQZAJH4BA
KS3PSHhCDzYD3fZ/fSNuO7ESyGw5MWM6Yk0WMLGQU46Vl4XS6wfyOBnyonHfJRhrdt2nfEr3Kswq
Xt4sOeeVcCwJ6zzpFizrceQroIaIIk1wN+vb6GmmOqsRgBmSqvf+l6jPi2jjzUAsoskFkTo2JHOj
omSMeIF91ywrCwacW//J4GjvbV5g8Lyb598Zx00ePN+nfWmU/dNivRgJvfWRU2Bd6/FbxX+ed5U1
BAN2KIJxS4h28er6Qhcz8S+ZCRT1uoIVahb4CwqZPBhdSS1uYig6JVjqAQM+ERwWTdLZPXZepIrQ
CeVm00qaYvH/1Me2gny+1uIvXcGAFEIlc5/rdAkWY+qFsyTzCrQwBlT3FImFOb+2F4zsLBHifPaT
xjeSsRw/zMd+cT3fF2FCyg6PUiFyBTuqfdZSoOeE5s2fLjgHxVl0me/HLeu13m9qeqMKsI2cgfI7
hSH7d0xo2ft1cCoh/4JQ5FZoklXsYQnAy/EWPKMGQma6uNOD2yxSFejDDYxJvd67a7IWJGPwuge6
iRPhYOxG2/l48Ml6hRU56qTiHnQTGGYVidxeLWO+yV45zNbD+GqaK0nTQzReGXRcBXi33ukTy0xJ
QljcL9k/3dASPJ6e7BMUmfktbettOeVribmCZneq+3aABfFTs8C3FoTujXS4vFRMl62e6Xn/XDPY
XZIeCsQg33wM6AitR252uHUVSfURn3WmKjm/Fg6e2nrOAFxC+8+3q1JJ/SCtidoXg1NK9MAOmo9b
pgh64eQWPceAZHyPAUCuEJirMnYLTDpjkuRjCp2/JxDoQtuOsX31/QPJsKm1WPWOCmUCcFVzf2pa
A6cEtjvfsrQwPNTgUxXfWg98YmYrXrJSZfz9Mgrowt/21DtNCo9N1z0S88/TeaWYPcj3VZl2kDSm
zqZ7w5odd5RNh2MtyIS9rAAzisYddRd+7JPVinOhf3rVHf6W0u/yo8UY/QLKC+tR9SSbPJVKqlpJ
AD21GLZ4YntUZ1Yyjca2+zRvjrrIUFCp1JwgBgqXmlu4tamEv0qtT7QpxDVMuUM5IlXQ14hk9en2
LPyZVZvlLMd7dqVKIBh9haLe5Y5P3l/SvDC3KaoBnQUfn770JBYTmigFHQDlVFdFrDv5fyUPiq5q
a/csXi7cTm1MqHEHcjIV7QMqNvaYe3Mh9w5Cr2VFden7lvemfDt/eBsyYZfeRn5P8dWMDHGTa7fw
7V1vLIJT6ET5Tzsn2R0g3D74iba3cIrzm3/XuWsEui/6xehPBlOmqrt7ZtLyM3E5duetYy/8DNHg
O0Mk+nz0mmnoAdpZLz7gPeAzDmBSyb21pMOTye5BZ1LrioioJkdkMcXUdNKxnT6qs+DMP/H3V7XZ
Qfj/h5mZsW4QSL+P766RJgwGx3B+6tkwnFzX5qjcIyRUIIhhPWxsYPBnCsfavaMRZvCZfIBbS7kn
u/0W/bSiEbkDBGK9BcQ7aVgFAETHS1fFmmz07fFAFdlUcSCg+xvOLxn5OIj8zH3+I6M2xiIzUSJC
vbCSy6VgotbZrCwRD0ewUYrrgfiPBcDNY/RGMBQf3kSlnX4hkEOZA05kIXKua3HgkxLeZrhzghZz
mwzwRW5MxrW0VnXhe9Lrj/rfxPHVQR6G1dtbP2KARrNBNflRrSMIyuYDBmXsBz5kLFd2ck+NT7nO
JpZd3BXWNVp7LtI0Vl4X3iiEPS6DdFwqeV5RsskaI71lC2bbO4W/Hi9ePXr7N/YOmyJICCX7L5Rb
a2c2Q/23/5I2NrgR9L7RwrYdhQg62cC+hzL85zm9W6kXAqs3kRiO2uQLUOqlOb5gHURIrEWJ2YAo
vwn4VyOZ+ugEs1xNZqs2Huo3FOuGL9vVwU9fePCkC0L/4UDw/EAs3Bg8dt2AUn70zabibj+HX8g2
eV80HLyhnXxwnAzl1bfh/L2rbwZEJzLnl/1dUPIgQocAE5Bq5Quyq8pu6rSJLrMruTlEjdjqDjXr
JBmu8wUWBeahP7qQIth+oDsHl7adoocLVFdIua5q9u/ZUWFowYQHP/VoQiLMWJxNtDg8nl1jDSzG
1OUJhQe3hjBD8xCMOTabZcMPBpDVmhaF5j7pCdU2rDGY837S5iRTz2Yw7r6VjL41qv5DNJ8hzMyU
9l3b9sn2bDU0uORK07w3jClGPUaerIJ3h2ylv3yLRjCykjtW/kVbIzCw/rKxC8IiYW924Gr/zMMb
4jg2HKfonaQuvN9ByL0Y1XKzGxTf4A+e5q4gfAbHIrgizOwVhEKDYVnGb+zg80NvMFn/G+tCfICr
33+1AzLj1bJhlRc6dyXwRkv8slo9Oi9Yf3ah28j731hRHyoCAFC9tUSJtNJLCsW3Dzl8OTrzS7ux
cBxNDTHpYwmghXaGfe7synasUHaJ98MLBC+L3CaBM2XFgilysLnfsgTBq1zpUbNeUCDGF9CmykIq
YAnbEEjTAXk69e0IzkzYVqdbjwd2wIM+1L9PACWwExbHhuK0n368A11v6Nb9Kx+bQsVsRl/CEw1E
Y9hQ99WPrIESrUV9wXNfosC+E9kD571pgZ4sZjergxbuaK3kgiikkKkEJ6rZ6K17fUsqLz6nhroO
Kc5j93xdN8XkFROx+EGeD32H/qo3xsDbi4LP1jmRUDR2Sr6b1jVHe9X1zqVFKLZ8LKPmavLusgEz
2RVGfgNflS6WX0JDiOuiUGlY8Hvn2ZaeW6BJukWTWPYz8h0bA3kPqoWsar53ESWxdcEZlziHvtlf
Cf+TpNwpwY6LJOUZKFf+8NYVnGJaDVY3K6QIzkNiqaEYYw+ucZ4UFJoKkgcAGWiJIO+GoBI/FTLT
RryxxdmaL9nwKNRDJOwZ2xyF7u6W7B+cV7Fvf68YtADi/iEQrxWEMdV7y5szsws8OWcWBRQLdycd
tIr0qNyvAleqUcdIvCJsvCPz/hWnq6EXOpvZwKFjiO5z990135zpUQnFChtKoCNxHnFk9ViwBC8c
twek0yVztkzYTrtQtV9Iw3xvi+NJaj4gJEidyRzpjPxJK+2i1NY/lTjqvt5PDJLmNkQFwZ61/KrU
0n3WX6hikyYvB5CK3Q5kOEpF44xp6GETahloyGMlZMnvabK84w0UYlfpqgSuAdANFC8PAcqLK1QQ
NbRr+X6rpFomq3n4GjowngWvJcnyQMqmBmzujUZV2n6ivgd+VqpVcU1rZTk8i6wXCVDf0Z9IIxha
5iHMEiHTlbZeNi+qHqlMVldCkkam5lYMPDv7G8PWZ2P+r0j0yViUYJ0baJc0hmPv75Pro9ja/BeN
1cZ6+W6vwB4ZaIgyNmJKRaUIqW94WmC+ZdodUfyNYVBBZK5Y7/GSdCPjG5kSCvPFUA0fBKj04CGW
uvH1knN7FT07eW3B+ALTa51EL+SmsyJT+pFM1nd095HLAyn2dsNoou5RifPYssJMU6QKMCeytu99
U2jb3LltwiEsy4/yQuvreTZA2TPd5J0AOe2HEARS6pLhj4MIkQKPIyiapKefsI0ON02xEQM/sYpE
MtJtkcBZA1OD8eoaB5wLDrrzL/PQhXA7Jlzi8ee2H+De6Fss6ubCC49GhvbxdG1cdeI+19Tg0eui
K3ORm5zrHqDSGOwPi3JS4WoM6rsut831Ld08LkPgVxDraS25Vahe51uvGj6MkamZZnVU08s9Srn8
/dWu+tIeYoOm0vAbPLxyT6uGanRhqkoPA79rROHk+OiiV9BJDDo0zHA4qW85NLewoksjM4r6i1kO
kR0uZ4mwkkCr8TmfNw8mkAkg7JjHUzT8mbS+QwwgdOGhirBYTG7kExu+O3+hiQ1InLidTKQ/hzim
rlEbZEqRPQh/K0IVeZ8xdeIfRmyFNrFJ0Gx3WJ/itNgBpkSkxgkceM8v+3jNz5aNyDVUoRD+nBXu
4NWRmkEkhAbF7twQlE2thAQaM5gnC3ZZ24SIdYZIhHswCDoZeexcgcOBf3L8Bqe08CZ9tNYjJubR
ULho1eCWNwdOTUyOUvvQciPian3da3N3wONsFupjYoJfAIjYTaPF3K4PvO1S31tFDkdq1VeJWsQ1
pw/TQbfH58a/Ln0OIy0smvfWvUho8GCd9/C5uB+ieK1J+Z8vhvXQaU6b6Mi+PyowU1x/aPOySPPC
cA3r0N5iSZiXjAdsVS7UgUDWPBygwznk7tvH1bG9cOmLoinRKXoXvF7Ncyqx2BZi7FGCaWf7svvd
nAwthJnwphjegOzDiVxC5HaG6Fp10pAcT+H/0vJ0s0bjE/pGTzNWmKOD0SGFD5nIkO408j+ugO/j
hVYm1irgpkMe6qpVN6c154NKjL5XBhVSojV0u6Q8hgU4M5WmwDVxBsjXbbXz1RRmOvdTw6jNeQxo
IZny1NxxBcx578jkUKgxm2eDCWaIX8nToGMBRA5+UgfTCmKjwctSKypva1qYIzp42gJtoUp5MXk3
cz0LRKGQZRS/1/nz1OdqKGyrT8EoD68oz/BuyDAgjYOqADglGl64HVWvwTR1ckNWnwm2y1T4SONE
+2A5hKD7xMT86gaPsz+rkyqqbxEK4AFkbHU+KOcD8NTF4rLdEJFISPg5Y1/XPeVyp1/3TQ7zYnlP
vyFGIjKtq+oiQVqhqkkjFF+xI0hXTiKDoUB6mtom+ds4A3PZ+kSTVd84mSnT7AY9kT6CWguNzM1q
J0jHEVfZQJK2hAbvzJ212YJiaCYa6ZIu5M/yD2bkOLSzMMR7DcjhusOf3npOT2nxSh8Vj9qgaw5s
QuhAwPfT+yu+6ZmxLXPsuiLH7XmB8wuWMA26ZXhdDGgfZGdjS3On6qlRLnh+DhifmOC6U1awRRGN
OArON8XrlMIImVfIHK15WvIi/u48s+zNJbr7sxPfPcQb8SD3uRvy4Hsfv6rfQHjttWvczMMTewap
PfggmHyBnIwIDThnYWnF5edZtzXybVNyUmZqo3JZuyKmRDZrq4+tOUGoy8cnbcnHsgD69lQwpxqu
dWbB3Ftlb9T9Uw7Sfh13J8xFDpfHpdjsbkw2n1+3jYXz+n7K3l4VOenF7k6f/AcU7m7kup86uvNO
Av64Y5jQEc7zRXi1dripwnoeInHFuOkNkaffW1DsCou2jLMg1+6z1X5JYIrMelN2T/9cDnIelg7k
2bVdpZc0dRyrKiaikLnZKcNIkLYYevQZ8Q9hHF+zThVSsiuD2bRdk5frGENobyIjCltSykXsJ2fq
FsPeCq4Gi7J21r0+y3QcJT8UXtqnGHL6i8xzVjJwctbT/G2nyp0pb5nkx1ikPdKncMa9UiVcDy2+
OB4WHlUD/7MEWUXMFpmSmbwfNAhQFs7ptdoyjkEeaxVZfyfSmy/kk5rtiHTwkvNQrsMbKBoO+oz7
vED/c62ltabzJr3Z0anNjuB+/SNHrgT246m157bI92Fq+H8pYGEmMPUQ9gsTWFsgzFN2dUOr3ZIn
vGsKcwbMbZkudQm3fezDXjxpv7WOyQ9X+wlVNeV2GCnV7YM1jt4Pb+SQCZLnHylLOI1OzC25E30K
djpea+tqvoga1LphZJxq4tprFt3rpVYXOzKUZuiuaJ0RBAHZQwgzd8cjllFMuGVRXvft1US2V8Ic
LW1Ttzw/WJMHqIMezSddvPwYVIB57z3spE/DPK2iwnQYsqIhQ52HryCne4I7HPwdnAU99Qv0o2u6
2QzOACzTJ1Q8yoGf7yUB+vjORGeB0cdAxDBEJKH3DKEO9Y19W2WfPB9tVIdNhWx1BfE5pOF9qyCp
vsfQmzEdPD3T+7WG7I4acr3SWAQujFQIaZ1k+hyC4gsy/8AxYDjqZO/PRQXHpJGMNQRMdF0fbTzw
CS03ZDpX88xqaRQd9L0zqFpEBbvhV1OAVvWzPTZqD+x1/67a/PU3oZ5oEyTH1AaNX8xoVSLEaJE0
ZQF3SPE1w5YDIdg9HTnsvSC/AgVqx7h1hpNqn1q2bzVdWaJABdkyv6S8J6zlKWziG69jRRlpGzMb
LNK+G04w9s8KM5BEn9FktzLBNCVcbAs5qMW+YXXnLssJgOxql5EAXdjwzPjqKmseAOgFlGIjKS3C
8AfNbC3qR7f+JBv5Cen1THPtBcdCapi6Be7bdCF+dIWylzlrKIhRPl+rr1vex4LCapM41M2iCuAF
SR8NRBOZJ625gPVnscsigwQALENmcCyCdx+PzYYTD/DAfDvnBwWAriDmNVB6AYKmxA3BoR73cYRH
ZUx9/eI/fWtTvX5LLIUyJI4pwQMb4fJjdFspxCGmzQKeCBKwrOqjhKWg4tjRsJ2hGrazpMKvTKcI
4tDiWxNK8qFbYbrPMCXvilsXt5gLjQgK4RT3tw0IDLA3ef0YdYXFnVvl10gS1XIkByXooCXLPFWO
mgKEGRi+qXWME49Wfa4v0XFCddl/p8YAnU+lYEPTO9fCvpazG4Z3lTqXGXBqsTd4QsPy+5cyuAK/
DjDUy8y9nugoS7iRa++MfBX7/acWkVT4XJHtdzUbqCHCPEY1/OUKjkKgNHpLAPyk6+lyTVtQyPel
zH5GvvNFPTLVY4zTodNSJRvkoaFSpQIWhKR8n/llzEEGWYtSAC6SNghhsnuYctREJqMpnwfZ1avN
0S8ao6T2z8J/0bgQcsqHipr9s5EMGhU5I1b/IOYJUHgB42eASlkKefqUmurmWXbJJ+HdCU3Ub9p1
iUgeWpwhtqPCCy2mlvaEvzxkyQNezh0HOl1DDRPEeifUWno7WTKSbx1sTgr3XMVkAKB0z140WU43
wSiNHrkaKe9u0z3B2ty9FfLTLLukJkvRZwfJRZETHXPUHueUXYFlgcxu4VI4TDl3j2FrFy0XwYBz
VgDLUYkeifmGi8KekQpPzKUewJVsAccIlPWRJYZMvZHaJykgXt0hSFB40vpWodpm/r9/V1h/TlPM
ESyOwxk+WQ8npAWZmLIH8fKiXLCaSPo2mc7UuCA8bSioHGfuy/GcC1p6EXBCj6jePgWPE+y+C80S
i2KJ3RHWWuy5m2CUtY8bGoSwqgT8KfWXCzsqOOaQAZoOiai5k9qvFYc/aOcQ2sDyo6ax8X1duQQY
W6CDEO8jYIBu1DOSiO3PuOs8AmfVF1Qtc626C9Z39VS1cMpsbgRk/mMYmtU8ZD0iHlhi8nkHHHI3
FY+ZhrVuOP6k1Dfw7N0gOKKugnu4eTMMpvL0YawUgPSJmMAwF5hzCUlBsv4wJmQf1HtLUXLdaj7F
N+u8zh6bIzpD6ZVM/qZA1YJcNHUYjM7xkSa3VA6qeBh6Gnp8rzsv3qqeGczPEdLBuEQiT35dTlGc
IQ+0aun+sfk9Y7dm54NymJi8esdKhfgaGlg0LFcgy1J/1eOUdSzBwrq7LWi8N2mePa8+sx5t2WrS
gONpgR38Dzh8685vvPPzD/Ff9RMQ47qbjRebEI63NouDyka3AAxLVVwKo0g/e63pexY5xMowmRG0
DzO5itVXxviUz4xSsYwnAXY/J1WuLpe0lqCEC0L156/Vmy1o6QhsruoD2jRT2TIg+sJacVW3r/EC
MvDMYQRlpIJvTNjQg2Ees8ZGX+TJsmf7Hnt1W2tR959Ul1IyRzLMMRvSuJHtyJ4w0CHdALvkRMCw
JmNN6yXdgzYjz1ZsVQM279k/DtNFO+X/wcUp2kHkZUQFxFb2DT1Nt/JUK8RfFe5dWPG8o0m2U8Kq
p7dYxqgSNvv3U0ANn3Af4iKV5kzoCyk9PTjMKD/37T4yvJfcFPCodBvB7lop/Z+O6rREeuRP4jy5
2tKB3KOiIEVyoCBg9avIFlZ9XELFbn3VBmo3SDwWKZCfbCSMD9I8EtctpQ+pFZN5/qg5ClLqv+eT
0qWrEOw6kgi8xQWXsERv5Jdid/DMKCESSL04Chh5HZxN6NqFq8LZTjfqQ8jfrlL0CTxRIA5o2t/x
deGRzGV55png7zkvpBp4uxvsh2DOxXgLjbsqxoexfuDdFYvJb4FJ3qhPCSIdWsXV/uwsq3xuYcxj
QaXGlzNuSxw3TG6OvgA56CHM7esqXiZji009TA9d5SyppSwIy9CGCHQUCd8uUREel3adG71z7Ojf
AVmkYtTbRvunDjwxnBDyF+5fzKGOR5oa2ZzQxgS+zBzyVk7Xoe5o8jlyuhPZpvYRWPzBn71S39OZ
+J/jN0bAhilfD9zdCOu+8k2ZNIrty8aZzYQFEzvj6bm+OBOVF1vdHFJJlsFWVOINLlkzjS0DW4Mh
96Xg1fxpzNUEVkvkFuhS/LvHZEBmoJVejNC9YV22WfPoeOf7hqLR1f0SPgcLbH1NdFu5nXRkY9dN
XSHRSCJBgU5LiDpFeQwYsQU0+YQ+lwTqOM/NfAveQFOQtmw/YE//D7X+L5rsB8g4HUMgOIkn1cyC
bPK9+S0z0bDI6JYT1uMxHw+zS3EyuplaAxA4SkzNOvNr6DPC09zdS3QUaQ4V3SwdNFTA30Xa89i1
ISDEwxD1ILQ6yByv53u4DzLrXPyk+bzDJxY9kY4hFbnUYzLYjNEUPQnIS2DNj/QYH9YIgWAEHXRG
iDP6jVmxb8oY7HKVuK5/mcALBqj5HtSC/VcvYIWTAmh+tL+bTp0PRDsaxo6svGA+miIgqPCkhtMN
66TUE3e/1KrQtzFoIVuARht6x0COHQ5KhVR9OWYOXbO+7ulXzvkvpuxA4DZxNz1tdv5s4mMksNzW
5DNVND41+Z8dXct5WFpizNVyBs3kpJ7NhTtLgs/BXDe7CuvLXG7B+2BPslqUydtMBuvPBg2b+5nU
vgzozNxVbXQIGB6Ocd4GIRpJoFck9SCyI3estgZZDEdJ/mnI/sdPiItxnAlIXHX9FyEVzZQkPYwq
tDiE+uPXfYbtbu35J6y1FHf7PAA3aL2VPGqGnGDryZ0Dd3lq/MP1NEw559VU82kYmp7Yr4gyBBbM
UXAybYnhPJghYyntzFt9ocyK//1fzfWqWeRyBHK3l+B1wBw4L2Og97J2885w09ejdRSoh0ZNhNIG
ij/z3cO6er2cxgnoQDhC24yVJnnMxQ7i8NmWwVpcVrdbXzMBpdR5AYhzmtOM4RKLo4KGj0qWDmKz
Y5XaGU7a0K58hi8V5YBdo1asFo190gYaP5VwMATRRfk4rm/uOIiUNtxpia6IszFSNq+8z1Nlkybp
OzuBdHdWty7w+dcazrwxqhkquoleRZ2XSUpI+OzhdDZDzI9u9cx4r+BhmBJUs7HzZlJ4pOQ4+w2i
ASTspjaWhO10Akksez4EDeXgO8c6sCqu/xg6/bJ6jG8Yt8joDUCWG1UVQDTq74EcV2GFzbImFsez
QmZUuG/jPaDgy6CtCnkWVtRn0OvHpj9OJTXYAq4Fzxxi6dIwICBkoBMKXXj2VYNUpEC/WtS02f7K
eBciifMoLq5WZ2zN3Rp7Xee64XbzfSTtGQ370vsvbvtLzC4PogUHnScJ5L/NqMPgEtFBJm16DcYY
7WploM8I/7Yzd1bbPKCBGmtIcPDYXFJiH3G5nBnzwdgL1tHsdQBddMcF3C54vBvmuN1PfTzKujre
5br8Xuu/F5bSlzhGslC/xiNrcQU00YQdlk3/vqD408z/ofuR0ylCJVn9/MgRphfV90jnkQwtsULh
5fYOPdA5RMRxlEZcMPw3JIosAvrBh/RMkjhLMjxHmJ/wJ78O1+w0CTONw/1U/QGsLNQ6Nc3EXocE
i2p2HKDEtaV4zuQKTaWTti8JW+GS1vnuh35MNXr/CfJ5oKiYPg25QBnphgOsjOMOUnn6i9XYIV6e
FhaMJEC1uXs7aFA1MO1vxr5iR0lz3o9w2LCCWTynvGwzLdJyXIFbt7OozN2goFZ+Sy7+zopRpKPw
13pftEDZ37ebXHC7aJIq+9iUeep7sHVrHHhgExsYaO3L4sh45t0gOfthxJDt8fTWketwXB1S82CV
kJCRzxAVkHEFTdISwv+x6hz7F98H6C8EXOXKOX5qvklOVl2CiajREPSjArRg8iK4QTsBFAL30RT6
Id2uBC0zkhE0S2Se13mOQ9rXfIsNTM7Tx4s0WmIYP6gnrEaHdcMvoRQ/kr7BJJPzQIvzu/AQvpwa
FD3+hjTx1PW0Z+pVDAOSxQVq29t9KtXQM9fJorFwjWtSHjp8sCjsqhqJ34fItQuhxqmpHCdkZF4N
9tmG0f4jUN6AEjDkK0fCcZjQxwC1+g8QZKux/pt3uCw5HcYRYneKgr8d3s/dWDbsqnIuzEszCrEW
h6mH8u9P4aCBd2bD+5CVLVnFryPVoUiBObbxCkYJImMBEl+zkLRbXICNU+kcOklYSJCH7HJPMGHF
Vb5NWq2YkMdt+xH/QhEiEq9BZR9z/kcHGjKyYTdKGrwWZ/5kUIL2612fDARgWA5rCodSidmleh/A
A3Sl0g3blUWL48/Cx+W8m6pTRF0dNbekIThBG8wUktbap/0enlFvyzBkQmKCkZon6dfTurlPnpce
L6ap3+JBNKK0LHghh6odT/H7R0r1qwNC5RK8yqfx/xoJwHB1aP4iT5IkDyGZ+ai44RRzmOCVlCxp
4oieOSffd7NcDDR1CEqbjYa2855fQG+RP9DpUwK0dXblp4Wh4vm49n89BKIX8R7zmAGPyLasoFh8
QGSn9Jmad9Sjwzz/EeFHcXqrMEESE5r21zyd/FbTIHoyqNUmtnm9Vu9bQAbus1+cgvFlCc/TRRNz
B28R2FogubU/5IuXv99Oli4V7FZ+P5me8XsvryVGPIkMU0WH1TlkJdLsiQS/P13xvMvwF/YM1o29
zTinHT85tGDXKIGdp/nzLF/8oJeElB6oKZjmTHA3cSuATavx1OWdyKsCQ6vR+nN1Gn3VceebONEb
XFnyrrqPQ7Tm9LwluGe1Qi/G8swfd9WUHnixYbtiILY2eDodO2jXTlBIGI8c18H43BdRX4uNRmjE
05Vd+OboroltI9ErjtypTd09MRR+04b1u0Iw9XMsEuIFEo7JVVVEf1ovOe4cCOWa3ISHeFX9tW/0
SJ0uyV1wKuAp44DM75HR5t8YC1I4xcfQQhm0cGlDviIOu/QqD2WgMVB/lCi528ErXvOQhdo8Tthc
CyUq7Zxqd1TZozjZ+sjZ58vNbDoXZ6UhxdF2/sr8+AyS2uJ1loNSlosXkNBbIyzFum5TSdRSzcJ3
Xwocw1hzhitmyiCGMh8fQXtU/K3Eh4yjW/K+/+RRosCXyaAhySI4VGi4l51P4eMdJSDpC/jpvP8U
JDRI48ngsMHHRbBCv4DldPEh/JcBm3LRSMzehT3LrmVhUtHCfVhhzBmXfwPD7IRXDXZy3jPENFuV
rST1hyu4L8Hbn6AeXI+QY/30q3dGNKI0y3HtMd7+PWbypBYjo+pvCUM4YqFJGHA6dZdmOAmPz8Dr
D8xpd7IfWl3LcxCxBbkBGW1LeMBsdFpZKAEY52FetF8pc/KqDWw3a9UeeUsGWuwkSCysNwX/doSu
vFY1259p/d66Lx4VrJpSGV8+g1gImrS/mK+jkWLa4B2YZKrqh8KbJDdWl/bC3f9R2kykUOV6fRSQ
K+JNGTyurqm2J1wNYazAclX6s/TXuH4GpA53ZAWpxuV/fGgN93XqhJJpSvkSbyGg93DYEjtFK7GX
MV0h7szXU/3pBQXlWi6M03VYbLo3SJ+9GyeiY2u39LzMACEZcep2u5Md7tVj434WJLFko4icmtsw
aRtdy6kGdEqknwj63vVIdQamRimFTTVzSg1lxwfqswS2DPkfoTWskmlWr5k/xSA4K2DkvEqwC01y
jONYMgpday+AGMZTvu1yA2E2BduxFI3rHbweXv6qofB89u1awyy+cNvArRnY8qwlvvKvLKi36pwA
MB/dThgB6vCARurEl4KLpuxQ6xyUjnjVo8js/GhWeEf78V6Z+lWA4KUpCKCYzPViaCxZhDbtKsT0
s/AnYpG+CYdb6EGriMwTFChtfn9o/MHTC+7W/JUZWwcq01FXDpsjLQj2MbyjJ8REOTXvApWQ5ytJ
IgBY3KX+kkDe78/ir6AcHL5Hpic/kYJTxLIcdBidpoVIYjekecW+qYsfUAfdmOwLdYe6K8x5jr36
a7KyehHyYOsCSmaotjnMkGQAVJousRwZ6L+CpsLehqKEb8axrlVwDQeuY00vLXit5Q3c7U3UZpGK
ohwp7Fn8fhiz5NmWkPOI72LhXwK7h79IiiNTS50IjV0AVoy2oKwm2i9vWW0rhQvwrOBGVfpvZui3
2OcpGyLstCDJNWBZVEzVYpYH5ha7L1iumzWK482gR7fHzcM7FO6yd76NqmbpwWhhaQQXTit9nFfI
/zWeYMxXu8LHwrNFmm2jzvi8ud404DmWQ7RtoneB8dUJKoFFCihcitHZHDuz2mQVCo2KRfidZm7B
PBzu9WchQNlDQz6mOTZQ2GW9QXSuH/bnaSp2UNDlqGIS0+0hrrTg4fAqncEktxuCGLKCzBrK/xPC
CGnwzo7kN8Y7pzOWptJQfjlJX6YShSokvPCoUIsZE1DZDOgazk40NQQJb7Hs5qVTPQeQ/P+sJYew
0tet6dTa7/D9KhDDbsWrCHysfwwtF3Ovmk+Pf91f78GFhwo/qSXxI8MIngJxZxu01ZzaEBrITIl3
Hes4Ij0kJmtgCYlwK2RsAA0BVQyns7jkzE/CBnQe6m8UCegpKtUXgmhziK3/BjQbnrOmS1DER7pC
btM5Jk+slkCzTMOf25TDAQx3mlicPeOpx6MBgbjYvdes41qe3mlvyAt9xRQjqhQnmhLOgjy58wI4
ZRyNJKCg6wIx2ajn+kQz0N04WgBN8dIirK4U/mgIzJUWdiFE82cgB+el1rforc83iPaSjCqkgcM8
BqFLGfNd8YzxZMNX3qKeZ3GS1j+yFlf6esFo0K5j9b2AqobSRpFZczFnXchUtlTSppA418vesJ26
nU7IAG0Eoai7yUAJAf/7+oiunVdLlpgPD5C8+MUAs0yd0ky+oDJlGceOZUCXAObT37Kern2ckl3Q
cLQsYRt5KsXOjYAjI7pGVWLJZ3bVSlzXOwbbu87/wwBGsSrg4soqvQWvP9lts3mwaXnUpD9VlJTh
4zSVJDGwx7ZrTBsTUZmPBZoiYlKAaTGtCljzOEi0YVPKtQOdfRrZQ4tBnSGcRUZvmbN/cXk0Ztxm
yQlZCWrbH5azOy4gCXEYnYwCMxLP2XfDcrwVP4X47sLPhJ9ZUKCVpw3dmLH0+nzL2T1Hccc8Opl0
MyJcZ+BPfHwZPlLg/cWcUhSaRfofV/OE+0dZ8lWpt1N8ue5ASew8vxZyODCA/wmtyAekM9ebgWNJ
uyCBEsXQuiyBPRLk4rde07wc12EWH/tBVh8N4bxXg7sQ2Lnffgf3fVffNm2edbsIVbb8WVQxgMkN
IFl4n6nGioKW+mAcUTs95wfY5IIhTnc3sXBgJDWvLAn+QBnMBPYBcffNPm1arS/dbQiw8GefqfJn
wzOlzkf6ykAAtnhm48C2gJRc//GZqKWzU5k1F4T2UGTY/7Uc42WANqkZLMydZrXLtjtm/JFzWc+Z
xkqIQwPCmgpvX+ny/roF+EN+VlJEFA0zixpB8XB6DXv4D4iAE/ssksl35zOv+fmXtqPG3kloWWuz
N3cu4VafzymImnXqhD/7dFb9aLjztwfK9xVIhFiotPash4ZBU1c+HrR/8zIwgKAXnu3nBipOqnF3
LpCm2DGxmvGgZkuevFlBczno90BGyztaMOchJH1cMeujHdLp7aFzlEjONRmFmwMRkcCsVjjfrEFL
cy1lyMw8BMNtoKO3vX5oDecYRRaM0+Kz7rBgI6APYHN45UXIXtkg28uwoUJJ1iQ4OI1gScJkBI6/
aLyLOFjdTZ9l9p2zUev2ZCNCDAnmInv9D/jYloIa4K0lujcDFlZuWrL1mrAIMGEuIF7XoSpumu08
7XEIL5+IT/xhVZx1LLNfEUK/O6n7ZYnC7P/y2dL4SiVaBE+SMMKKWiiC01G0i49vjG3SGXNHMlJ8
/B16J2oJohmToJzw6PKY/dSSrvFkFyPJBqp0nLh14a9IbSXvkrZV+8Ejtv2g1xIE2eSjwsc67UM4
F3SlBdn518aXR/WM8OXMZ50J5HnKefxDNiTiBx72xMMS9lAT5gkccgvJXGLOWMVzfJa/Ot1t/OE2
sklcp4aWl94IQVyF0kg53OYk5eKmPhLvNGHDadUC/a5Dkdk44IYgSOdq3d2vy9E53BNGExI3PZ20
Gtj+AtA6WPH47pAQYG2oE4yQV3VuAX1/KsCTpqQzZbm+/1j5/iNsX+jr3JDF1bfKrBXFCspyvheM
b8XSZ115V7+2SbDzQPDw+VSuyq0U6YlXVXFdcNqSHrSZo6xYJpeg7bYLrfU5rcJjrZRjCDoogqEa
QszRSl2/4KJLQtPifZOuh5Mv6JEiOcKsM5gNFFKNJrdjCm7ge1A3OP4Z49sHEVCUZ6A6o+FbX9K9
SNkNrheRYyAGFSRFzwIIXAnM0U0UneZb331dxDu6Rq0G8HJhbM0Ww/bclox5p/UlHHS3wsEiV2U6
j4//HQoknI8tyE9zY4rdVm32XzkYXFVNjNH7Qv75ZgJDI9EyewCsNj96dK56QebpSf2F3k0ZYiCo
RPmpnoA6S+7Ylzqe2Bb0Q/QGSoVks6+djHWrYcWpiq4AsDhXj7uRgntkiRtHru+zcarJJiz6B6PU
mxBhaDUV15r4QtQX0XfyxFJ8EjFr2zVB9t0PSjoxyl0KJmxDJ/68Dn+34hLHiHMqFTuHcY9YyaP2
ZKG9/Y0GG9MHEC8IQTBvk8l/fRw6fbXUOaHX/wpkfxGKg95mP9p0qxoGK9tiZsIwEI+pcxnWwV0B
6FfC4Kgj4bh4xkD47k4OkErQJrNi6wRu3Tjhtqewlaqja2tkezV1ed6o5rHGvXbWBr/rhMfBD5nt
h65yTE2vBghR289Av9TVwpSsRUPRKv4MrB0LbnqJ9w1dXN4ekXXWlrWwhLcHTyQYLxxAuA7Qgq/K
TTqwJ3k37Pqx4Isvv+mxksajj07yHw3susxjrJM4zNWLSwXrp6oJF+ymltcgZUjRTUDPonkQcpWp
Mu6U/s477B3T0eB/A1IPfqN1+qWcEEKRXcsi8oADfcPerZmUXb93kPm0tFX870y/a7cH4G0zIUIq
/Chy3LLIT/3uevg2FHKkMhQw9J3JAJvO835r8hHsyyvOaMUBUCsIYdpey1Ee/wzU69wKNzoJgJ9t
38cf0xLdrxkWsdy/pdk2uute6O2Yg7o9O5ThFmpdDQd4oKwJ1Ix3XcPSXCExPhwAxMtVi2TSUVbc
OL6uox3CC2BxqhDVIN8/b3jxrfNfoFEILbcEdrfk87uR14MpAiZMYU2gEebL+yy43INqsOCwiz/W
oq6XHwCm/7gZ2YHlzKsEd7Vw0x2V6ZSLJ6Q3HYZsnCXA8ZDTEg/+rtccdwPTr3GgEdmvzEy54sj9
64rw3WbKlCEtVmgQl660xf6IidpIv2qqXFuZ3yRhDT1Wt6+bDriFeC+FSoknYtI+MCrgAF4cFVtS
XXmLmqfoNghpuDLK+8p24iXDOusQJqsDF14QSc6C7DPyYtiEcfwTpZNHFo8AmAOGSXmSlaZeNSPj
xkN8RPnI1Jof9c3BmisMc2MzLoGq4gl/mxq/ZmRrG81DhSUp8LC492GL7F4U0bZkGvMU7+FfL3VC
B1GcpbXwGkZrNVugp3n2bjeK04HZrAHGuSh8vsxtuPlF7CKQ9tLU5yTZGTnfQsGTwfleTUdNk5WW
3ZqNUCJ401ycOQN2Ccl1M1Vr4o8KM4fNi+wqY4lIFVOsYe2unp9iFMH4J6Hzu4M7y7OvImyxMo2g
l+0IqNQ/uwkgZk5ZU48uTc6CakpLGkae+Qorfvh8/P3838RVVBykIGTBrPMnByt0Lqv2jPZqE0Jf
rEycxgg0Gq52De3QHzW3crpMUXLKPFMHEUQgX9EyyHskasxglR5MzSbyr9N9MgF0ByJ7i9O/AsQP
jkzd2jKXgrDalYlBYUGtKQc33orRKF6KjIQTGJNSr0bu2HwExgdWqpogROab4uS7zOl48s95huIy
LycHfB2/1gaArO6OAKL/WKqRRjTittojZ2EQPaxcvtq/4DDKMSrm46PhfMxzj4Ppbc4DcKSUmK5Q
5oYB+3k41YKdwAB5ozNz7RebHb11luNuZXDf0MW+ucvHsA8iMZQ7IAaf55Kofb3kS841/uqyaxDm
736lr+9A6lURHQseO/SV+7SG9OodE38KwuSTDWyPVXl5DHOdutD4eELFUqBxNS873eViH1FB5gLr
HDAkl/a/YwD8pTVSbSK2hsVnjmUiYrd5mWNeIRYjP6J+6ksRiejcjux7OSgtY8k0DvGQuPt7jsAS
X0YQ7/Vvb789yYXn7FUY2gv52jeiIDVFla1A216jK3ehyTCVEkaGDn3s3q/OpBbaYqyhxVOzb2nj
BiQuEmmBsUU5T57pjtlgkFoFgmu9Jao8fsqnIDxxHXFtvynX9YsRWGlDtuErChpBId6pkHr+cQt0
f2AF+u2xuPjkIvckENEZjorMcUAfRuBs2X3uQ6bi/sbvTipMVGweocuOr1ziUOtRoWvu5GBg7XUZ
Csf6WCTIB+zWo6aVODEL2m54BTyhzjX1e6DWjwucQ1GB1DAquzNXNvuZgm/k5aO5+2I2JP8Z1wdP
AyFzaY41upHFuCG2eWR8IO9T2fWED2ikkE1xP+fipvIJOkhFi/UAy3Ai0dXrv6NQ1ntJMStQ218H
HnCzmUXm5l3SEYvRPyy4R8ATChIXex70LUAL+kYdxA4k9qfyJ26+PQrHiyoPkAWVKlJQY3uJOMSg
2DnAD4Mr63p4tRw23RZ6eoE19Br//pIGLBmhybk77JiXxzJ+DV1hYFjsUQDu4zCkLxmSDwRYyevo
P1iWWDA2efqgtkes2M2Xe0asgVfyd+jbV+TonWzgN/LNmPN6tNBJVeH/Ja9dNPjxL5KJuzyZ66Jv
CCEiEWWIoK+9Us8xzhRwqz9FmfP4YEA+tsj6x40pCcUeE4yCsF40s8lP+k+LEyh2pfBBYmuRrQ9c
ccb9lr966k6YbqznGiSo6PAicO8GBVsrv3QkYH8xhgotRIdF8fgzJnN9bmEhoOw+UNsmUSutcK1h
A8Sd2EBaeU8FsxExN+duL/hWFfTbGZo7omynWWZCBZUr4T4s13lcllYPmWOd0QNhKdaeZ1URrUTO
/R0vxcjKidW7xePHKX3J5o7v93GMzrU2L+oiTSXedTMJN1RMeNy7hqXOV4Z51LHOdYbj0mh+v8E7
7CITSC9WFAAQLjdZiMNpJqbcUVur8wf9ouzSwg4DYgGyjLgqWIh5hGuSAORAq64lUFGMIhKIU90d
deV73zdriKaBy76NP3dM5k+M8zQPP5EsEoFq0Pgii8SJIPmEruDW3LJB6tcZ09+DSx5pI0mbZsTo
2Lp+k7q7ZL292udVQFMTJsSJHO1RwehFkU/C0ZHNntDAedob1ZUk+tw+WW2qVBUoCmUX940iJwnF
NXuq3xuapNv9DStHKZajoKKvDi0K1qIf4Eid758rkrlf6D9u6qHwQwYTiAWkfmuIRAwqJRx6cM74
F9A/Tzl0wEM2qoYNTsB0n9y6sgmuSTcB+kHREUWuJZlOfy8PokAQSTIbONaib2+a6QKYfIGPimTp
BOr2Npa/kfn8DX4MQ+XJ8FIK7AfvSdb094Npu61DEeX1xzSI/TgsSg7zt4D9/ADhUPlUUWXroTrq
CoSuCTW8qfP/rdswmuYXTrimPWEXDoUvSg2z9DqYzR6eeHq3p0Nv6loxkCWE3wdgPIGpPDyWHa1S
vZe3Sp8MjsAeBxoJTjeVuogMndRXhPVGRtEiHXlOPU3w4gfX4ZC/Uaf1wvSOCV5a73yKiRqIDkvJ
J4KMmXR2kPdxqbQDJIsE4z8OZVD4iMrUHDpwnISG809vsV4VtSDdblaylW0UMM64ldjik3+XVsQg
kpSwSJfRAaHaAnn7xe2L5/Gn6e5bT2dlRTDYrzor6KOdGkqcCQorpRsZdas8Yc+VReGn92lbjEdP
ZmUVHnU/cJrggqoQrVmknTvUvfZsXSXFePRVAQL9Ihd0aNXItNg57EAwxP312so9M2l6ugUpx/Pt
+mSm7wVQX0kk3QYUdSMrk6gCBL4VBmy+hmkd2S0JuXJQ2W2OwE1Z4OM6a2kn4n6+GP0UL/OlDum2
79R8Nij0oyWU7re5URxxwRYNOZiEnhUhHJGzRFQ+7hsPxszBpkOo00+utdimZAnUkQoTyKIA7Dka
H87cFwJn/2y5kiEmPhkbLY2f1rRluIGc+MkMx66KJqDPV+VZNUkjrpdWG2dFrO1qY8AU+xIXwRSJ
vHCDL5UsaUSjNDA3qNuvc8teOgIK/cXhH5tbpJgm6SUDWSSW3kHezzx8YNOiLruP0FN5JXPyf78V
QekEoTyEfefo6X9EISQinnIIIN9IhaHTeMgh2S/XSkflKiU1aNZA3cVBgPw07Kc3AwkAix0MWSMM
NALzEkNlUkDcNLL6FgcM5OKCEHBr5cCUgfApXZg8AP0fTRk3XzmV2Mhy91cmAAqUpkhuc9EoeJq2
M4x8DY2sgQexGarXYnkWvBCDf7HmaMtNQW5vGs76LY8XjC/6sdGXdbEhtyBqrft1NeFXjolfBSFB
18K2SPV6M+h+wNkVRmPkg53bE/1g0dV1KrLBZ41guNvK7LtzwHbqYqSGQcfH+veb7SXzFzD4pmRp
wYXIxZaqz7UUeCG9bfCYlkNcTJA2s3+K66Z6c1qUlXwmJRvBzVpJyHCpoOaqVLVF2o+BBzFasFxh
nR11FGhs4hVkfl9bYSI3GHfWcdeAWnd6RSyFrMCyml6Z4qQykFFQc+pGNpbOKqP/nPc9x/4QxkYJ
8C4+2w7HZufMRdlSzsdhpCXIx/ljIfgIAgJgRHbz8DAu0duDN6+jYXCxBQXoLqffZUDe+WUyxyVI
4pbQPvmuxQuDh+b0MimOODvOQjfHpLtVqw2HsCuLa95qwkir/DhI0rnXaj7fPUjiB/vpGu6gVnQS
8qq1btK6GNWr85lPONByrsUZT1BU6Jf4OFzRY5kYL3emO97H9LfyFESM+clrOgnvjo8wEK3aS5Dm
MwCwLCY9Z7BeXiLZASArJ5M4mHWDCEwzy8Yb/lpOGc2iUN5i015TyC3B+9vlXb4BKOPQxKF9MA4r
TvJKN8t9e1tZ3wukXRJzQUX/acH7sojNLSSId0oaSIZbOEkF6K2l/9rwZALZFlE8r0sBe6u4Q1vH
lpKuGGMd3fqgkUWeUI+3HAbjFVH63v55chZT1cZWbMJpWA0OZ2ZICOrxj7CQnLILnp+nTGUf6l7x
5MIGZ16IaoMjGC44TekV1LR3yucrj0Oxdqo9IdSmsSH6UfyEzqdrqPfC1Z455U2Xt/C9Nw4uFgoM
qug+trVFcKIBdouolg5TLG6OrhNUStk36auaat+ooiKU7jacKD43toZX43r0PKKPI6TilJC2wK3u
6Ri3ZkMI8iWHyZRVmpuoC1g1AVvZJ+p6boFUTV23HdcL+P8Mq2jVjfoq0GsUrf0D0OR7+N4Ui34y
MNsYaUZ/dLYFBKnzxK86qiWyQLAiDixBDWle0N2T6Gf5NGJ1fmJRgVFrAAi/DOY6rrrOZ9HTOMkg
W8C5w443z6jEEMj9wiXfE7CXUpBCTofwX+IhlA/yqOka4qI7dc9xseA0q3zvCIZZy+XVfIHy7XBh
laNWZ0aSqQOpskDKjCIv4JcrDX8D3CBagcaZLvxxqF2Wv7sRi9wY57WnKZweyIMZk1QDk5Z8kPOE
++vcV3k1QY3S8YoZvvqayoFUgMlN1YI7nBheCwUOVfJ7CgyMCUd0EvmoZVP1jrfEGmjlGadgLxqh
Ebjk6gsb9Ugds+U/TypKP3eEjXgtVK8ny7+xZd12laZqkjT6QEtMi0nIUZytjCO70kH1bOkjIyEH
r1UbYgtksXhwOdPDAR5GNfrJ/8Mmr9Gjm4GguIAK4Do/KXZzm1B3WJzfB04GfabhTHNR7y8jmbqt
uYmxJFMA5ySr/bTjW6MOscbylhNfc1KdioCzJ4TZr1l9DuMZHXZGQM6jJa1k7gPo00q7R9PtoVO6
3dKYohAMCzLgaOXGlmp9kcc1VUT3A7Dz7C9+ctrNbB6roGxc/tO0WAccZssXA5UYwVhFP62jg32h
zbCq7tPQVgW1BHm9yAH/lB/W3pbQjRkViFwpS4ygouRu9met1DpWECrZPaCOo+m8tZnz2GxmiRTS
V5imIuiguwjAde1mGAe1vZtjJ9aSEn7g83DTLvxN8+wAxwiEnnHMhvwlVP9+aQrDNa+1m5Gmhmd9
oCDVCQRsKH9QcqxuG196E5ybQ3o3RQRQCSxYfrt5R8i7eE+aapfQ41sl9lm7444AWTvxwAS9hOX8
wpEWgthtjV8gaIlP6SFs9qNj+fbI+YM2QpSraFTSrEMWvxeaC39tB2NMfbwBum/C5W2c+gvZCWp0
WKCe0qE6EC/Gy7nCNklXudv/La4Jyi5hTRd37s0YirZhv/mJHqNTtbFLS4ms+IMgAmIoBeHV+2lN
CugEOddA87aOQOnVVLHtojzSK1bIZwUfJFNEEOasB5F+xrICWnvVWHWrbIJF0AAEC4JdtjleHeYV
obK4XfBDJkL4YSXq9jPa+p67NoaFmZ+14KS9PB11Nnoj8zPMp5+R+EyeNzWNDdpTIyplWXMEKvkI
WB3FiyZ45KVTCVI6/bQrcfWn/QwQM2pyRRFDtvPHhHrUXFmAreSr3QItknIy5R6e4QCuuyIDOEvg
Q/VKZ7RfdXtSAP9sU/2oAT9pLvrsRxTVTjnCbmxmzTBV0CPXJ7K7HNoqgxsBbyOIrBaRQc03LLwj
pfs7TsoE04IA3sUlUxG2AV8pvqigLtoBoJ0rGmY3aLEkyOoTVcWkDH0FW1jbSBLjhp4VWn/uiyl0
5EtEfGUYp0DeS4GzQUMgH6GJQkp0Pgo/3rHBPoyobLiSZo5iMYnOnjSVI8P/jJyRJ2Ms/4DWvomj
6h6rnBatinyiK06k5FbzyTqTRbSmyrmXxXrD/OXRxU6BR+iXe8f+sgnrtZmH1q0MmdIX/JRmbkez
TUxge/R0tFSuj4GlD3jmrbBHlad9YEF8vFEm02Axq83cgmWm0fv/faTPOMhh8tQOaIB5dkLIup9g
MLu+WcITIO+hzesbFnsDY54CJCUahJ9DbS89EnkVDSa2v0GZCgxCKbpJIM964nZdas+DxE2K3P4L
GC28gH8JP+ViFzu9AEXWJY9nGBH84xLe5rSoNL3c4IuU1JOPi6zc7Gbrs/lkJ24lVZiKqxOReLDS
L9dW0ZGA9A+3HqQX3xBR1kD2b2lfvBBXs33Liq6QTSoMCzW4ZU/i0NzuMclO8XMb8JHVSyJmo5ez
e1WsJEtPUNfAWcUB2qVjs9rz2BN8Y8SsHUXvCa6VPOVpSLVxLYPZ/DyaTiR44HTHfC/9jjpB4aP/
SA8WJcXQS5hVuPgfotb4pvzKuSjc3pASVpiQqO6Q2kqdoU+D8LAfGy7GkGMyO5IRCNc4fyoJrvLu
+oCO6AUsPUBDl29xZJ9aqCpCi9+J/naYxB8YyA8Q6UH+E8QHswd21q6fzSRKlU0peeqHWDdS1+52
s4ZshkgZW4ZOQkw09PnqZ0Zh/ySS2MlWFxTH3kXC7LaOzosSIj/97g8q177yadLPq2NmyzR0GLk4
1OU5FJ/l4VLMCMWjsOzbUwUsAzmEo1VeIMeQXRYB10gJ362aFNrqwQH5kp2wHPaRp+jEFx0/smzD
HcYN25ZjZrD58Nuo6YSfZXlOBAmHMz63VDnKCfYosU8PVgSSFY0UiS0R+iOqs+8UqQ/rt0LFhSio
j5rpIoRGibm9bpmHE+mhCrmiirGDpWVI0iwD+fOg+fr7wGZKOUhfzeZVYxA0x+THHs4lTuGvRHuw
szrJ7fP7qUEcLQCePcnVebE9OkRE++EDeerDMvSfoD4rru5QYQuGZb2F5VQLLPjg9y+o3S0cholH
jclPf1oFrAtWGrRlL1cq2JwTnxLklt5jbJbNhJgeKJ7qHFKX5Q0OqLRQ1JSmN1ROXeXD5PNLtz/u
JiGd41wKnrRGexLMw0cH6o7jsbzCtfXM4gH+iKC9slvKpL9FjHOw4E1drtQcQ5UpitPUBk50FEB1
QKiFi0KElfbqlZRlW8zwTXPS1Okp/fGcN5gVf0cjovGUR9h09JpsEjTfb0JBKHHv/cNI+gPRve/A
LsomvIcYE1nq5RJSKpU7i5S8CikUGACuLCzhJOpHVsQRzTQtek2Se5aVAUhsNmTyIk3bd+hlfso1
n91s/7mtBxX9bgfNZ2n3V24UF5YqX6vh6shNIbqYFEeOyyaNzGiEguzPqdmRo+ixMobHk7INb3ve
yyqRXi84O1hpXbGN4qgtSekxC6rELRKGKkILP1R2dq39gNwYpZa0CGu+aqKN98zqb+lWfmGyMNix
gE0GcODecMvpavzMoHrG3m4ro3H3lOV0S4bUcTWSWeSyoY3l6Q2KDLa9U7umqeV2pSuPSP1LwLeo
KMYTLxDZDgynu17+HmlEg8qQEVgqusJh6y/L/4rBe4ylvPq0EJiq7VcJdqWG5vFA+3uhkEhVkU8A
i0ZJv1LUjTLXUFT0EaExQuesrHYfMpBMmaDeXnhwkhv1yfTHOcua1eP02yHnUco4lohsQFHsxiL0
s8ihsHNiqguf+wcu+8UHg6WriKmgUn0QTM+MgJCr7QOTETt9qmb60iCLN/XNAWlycitSYJZDYI0k
gbQ7IrWCXtrb5rpBHUhAOigtZYTWKgY3u2HwNVhkXAdPHVsvFZg7LWVs8Ta0d3rWLHEJ9qEnpBSp
6gHQJvbYpxX6iuWutyfXM3gh1A+qWmwNeLK6fomXguEd1tJfhkWA5k+wHO2rrgxvYm7BV4vU0H+h
/ammvWZv12+AeQd7Ll/KcOX6FnzhcyNa5q8bj/7oNvuSbY64Z86jQWhyWmK9X418LUzcJLuoUap8
faXxr/cU6kwdVR8TRjheWZpWb51s6d2sHzKY/LSY4pRHvzyekkBstd4FuqeYL+7/Ljd5niwg1igt
GWeJxN4P69PNqrl8L2P2RhFYg765KHwCxtFuPC+9bmn/61a/fje3Mw2aPC6J6llOOjj6LLHcDLGK
AMQzFwPmFIc15/e07MMfvOzwvFvalVxpc/GMpGEKziBi2KxcJQv+TM3zrEcm7oWCaaWnBNvz7Xsv
xCuBMG133fcmmruKCJktONz1EMAE0ArlFaIKyWe3iiA7/wGp6tUte7G9FMPK3Gnj3M8bie65LPHy
V4wwqrNGF1KvVYrkbBqPbweUZ0LXCXG0UwMBRfvOJ+855XO5oRXJEF+krZv6nBrPmvKuaXRYCFFZ
9QNSnEzRvkDO944SJQZHfhJyozxshiM6ZObKGWTRQEUNsyOtUlMlNycfkT5DmMz2BPBKLEpve0eP
1uVvkfDq0Eorsrg/4U+CHzQe/LGLasNitMZHoHEE/qtkVHwb9ep+qI4PUz3WauJZxQHnjtSHopgh
asv0R+WNnIXdDpWOZLCHWTOp0mlO6oF07j0kqXZbKPVCuBgzj5V9+GrS3b9CPJrswNDhQcKiKhZ0
rv1uMa+q6HS4MSRV9IZofd5O52sIgDSJpeWJ8pHsUzMNwQWu467VjA9WsBfRaRYrCbdUdj+T7pEo
uxEwfBr7zMdBv+ALWSZx7b64IqQcZczSBw/1zc8QdPFrKHr0pZ+7IRmQaMgEkEtP4vTVJdxjjMyM
LneOg14cwK0uA1ZuGgdbRmI4xx91pAlBZyT97BkIMH99bVV7B7ProMpTPYFR31rD622mJ12SPu3d
9jru24b+O3KWnmUH8BrUPIuIrWChER0CpWFkjvgY1x1q3BXTNl7AtuSe9iJaXDOyBr+ret8fO4XM
mve+jGaD59uGD5GNHqRfrUXDOHwQA9KWi6dGLbly7oVHk9US5TTGacAb9VGLjhoJuo+OHni1jFEv
QfVYeq3qyXFTCccUmHBKKyz9irBSIh+LYJ1ovmPx1Tb6NSqEhzALfLA94laJs0PT4uKCEnYn4xzU
K36NpXYJf/l7U7VasfJXbae5BHy7VyrhMg7DACkv31+vrwpOtIGIsd6ndRd8fVnNV0v8/mJRbzEi
O1up2kOsIUtzxgq0BxErO8XvKiONnaFmCRaFIfg6J5nxf/dMhLUaOAQaaYe033EsJCBVUWcdv8Kv
RKXBDfxO5GFbAdBHPr68z+lhmc4MjUsfLld5quqh7Zk12dGHNbq7aBYIm6mdz5ewQBCoJxNglwl8
Vqhg+7TwxLylUt7nBnFObIu1Yu659rIxtV0Mh3xd3H477zLRmZFSlWk2DCy61vM7oK6rOAk0bas5
1gUa8wqZ0LGtqWjFv+Q2GRvec5wNzzWNx4Xg6HxNp8u9Bui30Pfo4VZCUErHwbTXtRpkRUI+pK2k
GR4u4cS7b+GpRm5wpAbWU1vMIyxlsLwAifBarGj6Al3by10C4nr4gT8oFIpP9qoEejVlmwqYjfOr
35VFI0U7DCvWnBV5zh0fi0PY5RUWgpmQNgvYU+EdeEonWhby13dbo3J4v1CRluiW8ngovrURooOh
QFwVVOPe1AgI86OTZJNTOInipmSULDjvUHdDo8JYPhGKuOOOU/19Tomxtptu62PMZ1oQF8Hg8Owh
M5yx09TF5X2JUixyR6nMrwJRrCTzghKHx1Bc2FWX6250ZJtTJbNyWYQ26zyXTAmeKwAoHu6FAgXt
6MDjjwBBiixwjgOlRELhDUh3pyK8oXiTVpoQx0Avb20qwaMxB5riQ3OtyAtOCMESqkut1LFlCZlj
d5EcEJlq/GA7EE0V9OQx6TwJeBEXfMYfUxikp0gyLEFd4RwvK1Ho1s+Ope+8yqTfkHthuni1NNFB
9/CLYUZ+ntMhRV3qhU+oMVz4OqD3/A3kKrby/g7s14Om7PUoo3oMMUw2atfKfoOeyIPnIHCYn9Eu
WICcLugDlr4ZTgNFjBwpxwCxNJYJU8OF+6SL9wLEXlDJnSbEfmbeaIsBRP5agZobXEEE8kHsRIst
kGOrRRHzyESUuCdhweitdNsp5+8GCJbBu6kU7Zf+iKHZWKwvcowXUMVHvImOK6myIv2DHXZ7aZKR
+UzKMthKpOYMOYFOmMl5zoShxEpApHxGlFCsWg6pLrZ+ryZStoI/2tSr+nUi1AnkvvfbLftYWPVc
3F8HpfhGx8Dm06nO9LKgPvZ/1h9SgioDjHgmBQpWfDANlQOYwv2zPx347mxe6DMFsXGBn7kWkG/d
suztPQXJeEPY7rtBLalUOCl7wVQ38Kyee0j3SdeHl0m9IMr+ojJiPCukDFhfYYj0/Lt5XTbtuDgV
gIcqgC/u10+yZh/WLtCGWPabasrrNmLHY1uFkJPi+85J6n2rd6VflOgLyTBTldFMCgJ55zHX1uqg
SgDN2QMvMvW+2cwlap5Lgc8QkUBojWGOcmGUuLQqIv8M6tjmhDztbKnznkDzwdfV3AD6cHr2z6Uw
t7AT0fG5CjhsnZxLMGLtZb+QHoXcM2Jx0bH5/p0hESpL3GpcP/qJwL3odyApRTxUdUeqXSqUdl6E
TzCLhEtf2+f145mtZ1SikuN2BMNWj3dwMTJwke0d+iQQCpODR8eBOc3+aB1KKl3dNFWBzBAwtAfM
RltPuIl14eugzFDBSx6tyPLK6b1BGqrCJhUAow3aYaK00pwDqR/b05uIwv3tk/hCDgYB6LI+Y8wo
DbeMYXLrC/9UZuz98eA8EKdAIYmsvRk5A2VGhT7EebwsvFNxRrNzBWTv9XhFWTJuFkFSyqbRl0mv
ih2hoA04O3604QHzXOBfPMOIFwL2NiOv0/v/bPujTrZdu2ytJ6oovv14AO3IlbIlaYnZTLziAlY8
vwoZtzErK/uzL35x4r60skNc0VaSqEGfa2XgudZ2A3xe5agPkhEufExYLA3cU4JPkh3XA69RUkEG
+DFHGZoeyWkCi0Mg41urxCF0avN2xHxM9woWgq0rJoluxfSvs0snqzhBvqXwmOqURwO+wQL0774w
8GPJDD4ueOkHnHIWcSJ/Ild4q9rf5/igUAc3RCLbJT/UhwQf2BgUkY/YQJpuEshn461T3SibjOQR
IDpaHpYVB5ujuP5u7Ck3wRN8Qks9yEX+peykaxNzq/9X1P/AH/vgqBBvlm5Wr+Y3pib76JdbBS9/
K/xu6Yb3lmo2NHBvnhpgThGvx5GYOyk/GdcBPMkLoRmwdwAigl9M5NkTab817KBwQ6p674V1s3Wg
2Q1bjnkMTZA8gXn8e6b0HG3AX4WmoBadUdhPracH6f9e2YaVCnNJLJ8sh4qurGpBswXf1+hxVUVa
jEW7snXCTVf99NJA4VYQdKmzAKl1dYLvnQX98aT+3pwv+FJ8SljUoYj4zBtf6dmPOzAX4cTJYHL2
E56iuQEq6+2nKBZKQYYpnB4i8Ojv6Au/OFHB29BNa/Hog+vg5dfPV0rkqGCDF6+GY4EGQXu8DaEa
gzh31R5lVelZTd0njRAudZpKuhzEDX0YMY6UY3AG6+GXHiBzVM+weD025jjx/yFtJ0iC/aHYopDu
mdb6h6rE0XWPl5eovNc2SlqjtgVCWrtZKze7A7fgavHDP4mjknc7lXY32lR8pyPGnziFWT06gHyc
A5hgNe7CShls/vO73S3MlQgM+gm2vTfP+8bV0CoFMLsE1AV/RlMpCnfkV/Ki+odZUC2Fk0y1bxSC
F51qD1RKpLioRGiloYk+V2ghQA+2X/dHPpc582Gqcu1wg2GG5ph605RP73R4zgTIsxzrUoE7TfAq
Ao9ppn/k3gI4pEZ4BjG3TQ5OKdcpbms/5p3oAS0QPVZXb1LSwwZNrXgGcoeqHKaPnwfOJThTiWKa
28NdRYJqpGgzFaJpHwu0wF4Ukq1g1+YuZK2ytLbhkWdPh8JXMolUxXUvklWe1uJdcCp2iZ//wFgP
woZOB4WsBxpC6F8MMh7v/3di/22z/zPsxePfvQRL3v0W09QP3TApvu7wuhpS8Ga57CwUYePi41Qx
/CrJpX4tWfjbnXN0QXsqu9KhUkMNPMf/cBQcBUy4jFEtzqZLJrRsGYbmnxf6nXy8vzJWPeFp0Q0s
7iRbhW0XmpmBua/mJE1dw24oZJwK3SQ30pp4osCvGhDo9P3XxCU7ZXKKJSSR3cUqc1NJPmw6FmiZ
Ya9mRmSTeoHveRUk0TMBcGtEMVQZ4lFiTnAeAYlDU2GyVdwFehJbQLYJPhhFE7PmL6eT5gNYiH9i
GwNcKRN8awv5GbCA9CNpGJadc8+fknFduquW8U3aI9zBLDKrs9uzMtneB52htarvhCk9r6fddCIX
kzVwv8NvCi9eEiTOaK07EtadvZHiC7lVTjuDBIUFHRP8XjUb02Y24jKYO90RAEXUQRCqDfNUDXvb
rIdJxBGKLViCuGAN6zw3KPtRUeo32LTnYEt1edkAxoqPabR7K/7VfkSjlizbzWFazogptqGVJKHM
mX5Kyw252lAEdHUVpcGFvpphpFSgW5BrUjbn50LoV9K6vdIhSZRyHZPTitqPtiEXxRbRzP7TJbvS
01oxNjDC5VlFTQqfpahZV5sspH+FI5ahK7WUn3NaL4RkSF6gMQ8KwAjEj1NDyG9gjSvTW9Q641ra
bXC+XV8oAyOYz8KC6vcyzLwprY1qVUVnmdqNOij2oZj+eA7CfFpJw8oIJHO8dIY4n/IXrC2gZAu0
8QkGfX7k1nfDSuHSattjCk//UOZr9J1zGAG+FoFvFE62S54exVoXd2uH/tXZCwWLAP4V0XmuQ/vs
VWuWDIceJ4o+qa5pqQ+iNy2vPOQ9w7/IUqspE2fE32wsovtrdVO7rVvglI2nEot4Qk5VUGq5EWDu
zgk6D4nYxaSPkfYazqpDKsccWcEfV+7J1woX6ci8iTpWR0nRCo6ilFV7NrvKfh1L1OpPVy+MW5om
5k6XKvURLFepabKLi2hWcNnTmspElN5LOcvFAwxTPQd/rTRp9pHzNFVzSotV0UvgqNR9KQHt4Owi
1+YBXoH9ENgm6FvyzZl6uTUEp8jwzUEag6/2c7bHLfvZ8Ik0TD6xTGTxNkI9fSw/zH6zU+4M25C8
ZPP74I4zp4t4Ds+aTCBfWEZv0IoDCWEVrsFFUuCRGMR1LKfFQCQ1x9lICR8X8fAUwrqRgZnQweJV
KR6uM3gkZ7k2qt1Wv4E2bzhu8XXmZR++QHCyZo8A4qxuSwCmCbfGqG3KJVmut3DM5f3wvyovspyL
581H8T+BX1edCMxEYkCiCIatInitrbQw98oIbQ0rJzgtAOn1IdSKoLE3hjIPBttg1BoDSjRoZJki
rNhDcRJEeRw8hNlCnBTCWJBaWMH+pdYSf8R0NXtAkg1cOzN1XYBdz6m7dzUboRcrVqg3r0lOt+nj
jOkXqgkpU2ieCyc3TefT1KrMADPG/fdawEzhgtBa3XktJm2rKlGHwQa7qLDbQfTJpFtyQSRCWXC4
H5E+D5qJQUerqo+0m5vKo+JBAsfgZ44FLBscTpN2n6TwLInJbx1ctWgHrYA3QelhUzgQQRXpaBag
nBh1AJKqkb+UCB+2s+658mG81zQTBmfbi66HfIQVDK8BjZycjlSIEXuaiq7m+SVVFNAK2HQUdb5r
MiQ4u9V1iP7AikVv4sd5S5WGolxQohV1MyOvSS496BCA6y48Sr/DpF4SXD3ypil5thqaXEviIEco
CLrVML6mEauUXTXbZkUXaJHO5FNXuXTPTpHGyOa0/hICcpQ69GJlKMDsHOuZYugt2rHcHr5A4gMY
r06XCvMGiK3XXnsregp0o2YoYlu6yylUBKt2HQumBx30nCb71jMQjDSYNJTwg95uJcICoDHktkt8
huaafYQVPKDYAWvSpIviHZgGJqzsgFG7N+/5yHvD8Y+lmqMN55KHI7mE3ElSleoZN9RmycONk4Jw
KcqsW5b8FOzaQn0cdFQ+Hi78ypUCZ4gBLpaSzpbULWaA/lNyxnWDNFj5Yj4Fh/AQ2kC5+iMQ3VMP
VaA87mDaWLQY4g0r+eEhAJuGcgaS0nFZilOP1BFt/PvbyIocRaQ1PBHoYAK37wkjU3dOMM7/wiKE
X2lpHM8b8wTXOV4mrGM3SZJv+cc4ww3A6hdheGz2S/awaWk191ZaSyDVeWHV5GxtKHkIirlfn2cD
3/d/SazpsjQ5RkoGq5As7j0Amaic17ritUTapuqk13eWPx6EfQoTL3qd/MhKOLoPXly3dJL/HNS0
AQ0TeRNR6P6xU0qZh3ZSZommTCYcpnpBiONfOs3/dze/aEVXlqsdrZn2tL/pq32RydVd07V+pptQ
I7/NjCGZEySgYQfNA7rxTQu0etn8/dMKMiv8Z88hawQP/7ALdRV1eaGz5L+lADTOPtRfVIhEw69r
/OtAxmo2787BWkCtNiDI5C++lWM/E6+aHIVeF7OPzvufKDO5iZUQORnrA+uv24DWjIK+f2+VZePG
Br+nTWH7utWpmrUfeIFJyO5R9qM55Ikc8PsNsMAhMH5pQYNCz9wmCQTfqpFKLQgNNNEj+yWgDdIo
JTKMML7Qw7LyDB82gnr7TpFa1A5bQ8rsbSX0kYZTiMbWZVMmb3Ty9IeUhyUVswAnQek2rQIG27sB
G9awXHVXc3VGW+UAxvMf2TrnWGzPCwa7s7A582z1PLsvcQOIp3itVmacvS5DKV8nhtq6KwQUNuDg
KDgGvgVn2NHKdG2ZpGkTmXCDDeqjCJ++2SIrpGPd+5hsw6v8/eZz9a0P3BSbXlbNqR8SM5uMEHqk
rBd87tjzm9jdxVQ1GTQZyPHVKRtCZGIwnY6W33PP0r/syWsJSYyR45SXet17vvoo+JhP3vNJ7YV6
SQZmgWD47MPfGkRHk+jSckqiGi4H2GQvd6CRVUZoSLkcFxZIdxLs4gAGlNkvBE+m/sFTFwIi8wia
WOvPoUMMnm3UfPizxUj77yKPDngJJ7hA3HDmVfUyi1HFbZBbeKNfnU7UcLo0l7iv+ZmENNz7c0jd
q29K8S2jcpnGIZDcT9HdnsDmjL8Y8qqPX8aM9LrGKukqBMY8On28wcJUaXzDwlk0PIZck0JkmE06
ejZfWGP80gz1hcko+699Yforl28PHzGnG5vJ+dpd7l1F8Tz9BNj/MbWhx7/jb3cMWtvSBkBBUysz
L4YMjsZMQV4ETaZmQJmbEzyW2YvmoO/iWNm1UiFhqoMHmG0PrTM9TGNo5ApyVWkSXE9kfGkm/0eE
tpPPtm/huuGv5gBsbeAIi41pcPbiMONPI/BZh2g3dTtYXkSMQtr1KEQFI32FQRdVh9qgwwH3B8j8
e1ev1AShmkHELFrZx/S/iWes02Y23xQxD2bmLPV3Lps6VZ/0VXQLOsaiKX1JxUTjeFOr5mL9m+fI
+dbd+XEdhIE9tC9R3ZqefbgUkRgKJHEsAFwtUpJZoWo8csM4fA/XYFAItLdzZQe6l80FJ5zcZ237
L/X33cDUhtlWxnrXq0cBxYs8ouoNJx2Kd/fPJjbcssnUctM6Gf4SeUyjNyoEYvjj4j10uWYuVbw8
5iS5K2ZSfKEKLYhF9MDZawAUOeszhaXPybq64nsswSWXHCUjIuQXenDP3/E81FVsCZJfbetW8uQ6
t0Npq4FGvTCedFKc3J5j5Be5uFPerFkgbvIDCjoDCE67KYolHtLZrP63+GUvmZkvFp5WU4203xWe
K2j1tf5n9M2GNE2C7MpgoDl/79o+zNfdHO2RN+hr2DhQUTvFmMAmRK6vI10rqdUeQ9FImJEHtXjo
FwHlLIV8l61T8cJUxgv8iEPSRexhgFA63dRbX3HtB0/VmeO7VHGxV+C4ftKHRnuUGRiazsAtcc+m
3PdwZazXhxhUGEIylrJVrNdNLjxZN9m77gabvMn/BHV4timTKkcsh46xJoDNJSzSKaubgnalOl3f
7JcfBdKKLBDUWFCdR62kM4K0c905LpjhMCfNZySpQMl8NPoXmOZIqUjTmUNZ/hUJ2ukV/9f2qB2p
tHVXMSisNiMDer9y139nxsUu6Ewm/6cXvxc5s6yMIcVPDThKDnOKWwBulZyOTij5xDwm3ZbkgWzj
DorUcQjTQP1kJzyIEQcafOrnRU908ORwWCTLQ1G9wNTlFzd5Ibr/EJo2QLtUJOU9liCHLPCaw/L9
B0p47negwRXL32lCO3e1+UtvE5n1ccs10loEGLz2YX6hYcw5XiFiSWS+Go7kFv2aK/SwpPo26f/b
AtBASE0GNPm7vA9+pf5vZfX373npNEBUPySEDHo3IvA1S7eszYUgqvRpjzOVMiXXAXd8Bf/BlL7o
RLLdSEQZM5RCgtcrNpHCF/sqlbhNGQNxlMrihcAAWVS8j0UNbNVwzOgbJr0F3nUozTQuyTz8foEf
5kq64645nEg3ohRMXZ3835A898ki4sBqKkY3wyIwFYuPoeYIQZ+BmIZt83wJ/h4SvE6m6XiSls04
oaOfXSHlcfJE4WOAXF+oVXzp+EeQQoM4koZ0tH2cgXX9K721lzcJOpzXHoR4t0FuZYYGbkQ6tA+e
CZ7MZKtTMwY7UFpe9MoEhcMqxIWBBcbIiIX2VRxeLcIrJ3vCHJk7lDqZ+APiYwCRETqlZsn0HM4J
I1TA3NBZdR6sZ1K2bQkqWUbntaMG4PBkir66q2J5xeyxv08IobStHl8OTuhPZru770faw8VNyYQD
Va0o1N0lMRoZoGl4fUTo7idThulyDA4/5vtnsuBo5Pj7FOHgIjwgYhehl3bwtP4WoUC/M7asvtio
4CWPRD4TK1QRkDaqI4tGljyw4bviOIxf5r2FzoK9bDsfzE6wz85G4prXCUvBiQ+bIYKbvIzABoY2
2PsgBv+kbc3QYnGASb3yB4kcp9zz4fJ/bPPjC5dDEB1TzhcmCz7P7njgd+vT9335NR0KEJgqScj9
6acYUhUzUYXI6ieXMqtKeuF3DDy4EounR9rgzggWlgF864xkjm89sB3mNl2d8NV4qyVlCa9nLGrJ
+sxo8Dy0WKXqlNmtBGBIaAwPzEVlHbodWzAZBkhPpJXBOqxffrpJD51+CbkP7GOJnH+1nMWz/Ead
n4FF4g5FCyj5Iuz8nNDXu+y9FkJaMqKAPJUkoaLcQn7L6giFSGCUcAOwN0QYPItfmWngVbpHhN9Y
rA5TcPZVkguA3JE+rP/l43UfYYzqGwO+1t7df4nb8vNaMorVUaYaw9cq6TG6uMvLJHnG8yF6++vl
yMHShkV3qDEIG3qc4x8DN0gx9TcmzFDi/Hssyy4ZkX4lHaAZxxP0u7Ly2Su+RpUIMvXnx2Di0DRQ
OgdTgAi2qmsbITCJO8bzt08cUfDCKE3CR8WKuERb+F3e7QZfFu/OyB09O0kkFlu+QOxjtLJwQAqq
bkel23q3lBzDYsfoEUShByldW1SPY7gMJHjdd74GGXc2VngvgXZAp6EL1JJXwZQT7OChJAkzBsBv
upNjIl5MYxO7IzDbn7G06ZQJSzA7HKN0GhgzPzS8fKxJU8sG3+iVTtYKs0q2u7Niy4dnj8zlOZ7w
Q8u2H5o/nISzrtsRjuLExNWZdkgpAf0hJt3Lfx9lAC2UsrDh8anQzFyc8agBd+b5IrHVuLiNCdff
0s/xkqV+a8AnnQJ+B/Am9vA40tTc5qWaUFO12ikw6EZIVIQm1ZFr3Gmz768KlQos7nHxlnD9H9Hr
rURM3mO7vJ1nIS3eKrPa8aXmutl9aAAI6tuKC9veAIE4p0kZbFmCElGdeEM2eETtmXjnUilZrjD7
uNx2U+bXuOEe38n+zSOiW1e9ZWkZbEZSWWS0JctifMQdOiKx7lxe2yj2zMTwPKsEC7Q27lyj2okd
6gZJfd4+aVWP4a2dukw0A/pui/kWLmMpFrhrWOzx0LCvpvwlF+pKW9SfbTF8V99ZFYMNvtuww6BV
pEdzdeEK+zLQAoAq0sSTwV7B+GvFrDrp0JcF+RymZvsomRAB2i8EPEKqtKxUonX8o1ft7X/+kVCh
q1t4auRm8Um9CuMouSs/L80N+B+E7fQgCpFg8Su2l7iMXDbdcGS5+5ArDaZ3+7je6azOjJZ4N9NU
9ILBTcWO1bVWj8osjb1fizQTD7wu6k0c8YCAto2pERlZFifBlFl+4wblrlmM9xlPhMNPyZhVqywU
wmF8gLTxd4acKCK3Jm7neQmjwJXyK5hWc1HjLXkyU1l6X37Cdb4fS6iTCopALrQAjvbbh0Guifk7
PtfMa//3li+eEx5glQId2SDu6f5KshKd59G7Iih+yZOow4imDiSUo3RaeG2ZyiDPcARWoxdQcX8I
KGRiu64/fD+ZrUqK0bDYP/6Jyxe/1g5kgSXrnt+Kab5D/nF9Z73xGVLZFQtB1kYwjhS0AHzgBADS
loIydAYAVll6HB49Rij/tJIWQqhLQk06MO3E5x3Jtg0VDAhxncLITc1CcHNJUEmawQZ9hucY0S61
ve88ykLk25sdihX+KkdO6qibTDv3PjnhttW3FfkNXgrB2UkP9Ewh8MxGvnaPHxIua4Fs9nc8yhA7
Uh6dNxO6TUlicMKhYk/Yxuzzf43HgKPy+/ritx+d5AGjpF2l/ypZhpoEaAPSDzoPg4UpbiKlRbfy
lWeiPB520XmfhTLfo5FMGyqpwn5ZDtTSoZ6KCgshJh4qaiFDS6MUZXoEChYA54DPJP0xwNhOjsyW
irKfL/L46x4hbe9lKw75j5R82tV+xWmhCHu2cpqW3KiRpVRvc2oESd6tXh2QnVeMNbwfPe2qRzn9
1tSv5IHfWcQgqbY5mhwsVrHUHqj+zFZSZD3TXahFW7pfFyf+OMMXI+yyl1C98NfFupracAlHL7ps
JCoypcN37fyilaGZxoJ/AO2eHdgM3F6+Y/tMFWqU6n+liirvwZgnmMMVQJdUj5vqrEiKJ/pPsNx+
Mfle38bBJ0Mv7vilIItgP7vFb4kU7YvZs+GPXnHMwKNe0qECGG467VTiKEfvtYVICkjqaLNocv03
/p83cQE25Xy2BUfcz4a5p+v718Ixe2OiuLtiMlopON1oUQEeeuQn+JNW3eXeZmlY+Tfpljnmcq7/
1FGMorC/xqq/5JOtTEnPdERaSVTqwVKcGU5g7tFPYpZRdgL0C7cHJ88EWkMTJA8qqiUo6X3CsbJ+
pFkl5Eap5Nbq835NAAxoCEDnmHWnwJISzn3EDxGj1RjTpYsv7l+2tr19GvBpER1q/qvVPxUCjtfK
On0fpFX94dKpqNY320jf2vbDZL9ZD8nx7wfuLWFWnpPJRp3HWNxNCt88hiCRvZJ0bpbffFdACUct
NwokMAypfmxFMtbrAc3WcPHmuMW3G6+/g74JavTsKBA7pbs75Lvul/laSr9cF/UQnFTy+PzjJelJ
5qr4OBomOpOC4M8cMC+mJbzQH4/ZIUuC8yIGMgahZ5M1fRa6KapW5cMksOEceWssSCPuLRyBE97n
N1GkfnSd5rbwebw/Db6rXQ0wbLkre8WBhsG22BMMkknOKQ16F02c/SooT0+rq0Sv+0S+k2Z5vp22
JKixPjCmKNYfXjwITgRipdz7kMlWnFaiQiPh79BkeO+vKlOYzMFV94NWceE7VRJ1qSD9+bEhz5d1
elOEbRsLxy1WDQ3/lddjYZG39ve9aB8U3CsaME9V6G4Bomu1VkaKO1gWIX/uHnqjBEkg4zqzjsFD
g2ZY81sLGh+xVpfYu/Ixmp4augqZFy9VXiSrewb7ermFodC7pK8a1hAoup7EuH4wweBk3edsZDCf
bDZGnCJ8N4r5LDoqQW02k9N5vtSPLAYqtmfnNlz20+aU5jCNdMUiVtGvWKG1wppjeiAmMSj+iyf+
N/Ad2HP8N+xHZayvmY8Y+7mdmokdc8FWMhOLFeBC9if4xZKM1VhnwDhGgz1LbLS91J9TcrS0t0L9
QKNSGJyhHVNn9Xs6IPC8eu886+cy7/lBHVa7BmG2sBnYxvRVn6fMNKWEEDPUx3EiI/Psfst1kK7Y
M7Cs0Z5WTJIv3IZ+kgzVGJLSnUwz83k7hCwHrdKkcDb1HVf9q8L37YjVDS70hndd97buSYmVg4d5
aawVMLmVMr6g8Nl+Y/M1z44TJ6rCkSshzQE/HgAgwO8uJ3SL4kwTuY9M/KvjnrSZ1h2KJ3cnpUSC
Z2uEJPckYNLeuEwBnjrLcVUPh6xwDKWGxPmavBNDxex7+kyqHdR4NJrYTLSCeSWPKprzvk06GVMW
PVZIKVPcU/GVXvBkc/CW90+CYPCDujbUw5d4lVMARCHw6T/xRg5gddSNqecGWC/oOsLq53/7BAAh
iE6GW/L+3m2Lq09oaGCDeV0c+ToRqpyMPy0u/BPMUhy0xcY+9VdpXm0I6QHkz47PUBu8fw5EmEU2
G2NVm/JjmZyYTYYW5dAlIu2+yj6gCjIZRWPye4Yak+288BZw2iHRs9vBhffY7G6WgBG9TC6rt2CY
SpAOXDCIziGgQBLI7uJKqrExB2QVSZrq0aqBBzA2C+YskHj4Z3XMTA2zn5sAXuuf1oOEFV516xtD
QQRU8EByLbBY4BTq/vi2kHPnXIf5w2nEsglkCuDeyII1eZ7v9KOFiR6/ZNmsgpU6O86TF8FCvAgT
yRfSH07NibPoc1hLD7QPc5wemmPMyN129Z9neDNf9NiEDoWCbROb6yUQ8CKIYYg7nQZ9IBBqn0SF
SnGc0xFmZT2VwlxqGn7Mk9LeD2QmuTbyOZz++XS9THGZ2cdJrsW8fQr0Cafu473Oh2racODg2r2K
VNhq0krLtO8EuPCG1ptJycbH1weMv7v5/qEE+pH7zp91MzZxQUvVmtJSv8GWKrtMxOSdIw9KUHoU
BCTrFDDOQWKKhZC5iLbh74LXKN5enLz6rfjVoSg1BlSFezuFwSaxDIsV8wW2xgN2ML7JptXVSBcA
X/QtzxROT4/or9Yi3E70K3caAwcQwISRo6mX54zLdBGkWVDI4dSXnW4RAMQ3n8ZH0g4hh8tkc3/D
2McUv5DiclwApCy5LtfoGuZX6IBu6Ir8CAN+ke1CIH5iHLWjhCanWO6CaR19dOT4sF+z5wOQS5my
PjKnT+AQHS52uNqGuSWb4bprGOGzhg8KsmK9SGyvh60PFe3Emshlp25dZCkWO2sM9oDPCRBsb4uY
AnK47j5qGPAwTVs/C6uimTpmjvvp7PkX2kFvjuIZkvK7gDLOtXHTGBl1LjUqYNZe/3lUUQzUmO7g
sLfu5ScNlrPBZj5SN+TR6kG3Fc8HpV8QkTosiL7DuncrmwoICD4hybGdNNpt/6WhE1D/GnADVVQ7
TS7RyjEuEKCOCJ5TnsLVs53CmdisWaEAzO4mWOyyAP4dre/ag8kMJBdgUUbHE6mv2dAc7OE/V5z8
oD4Am7OHyjTO2MaaqizgZano3Z7CZd3XXXf8hewa2DySMe4pYAB8B/y4BRlDJIjh+kwo6Ay+utTT
cERUrr94LPH7Wo06orOV8G0SztMoTy0GLZy6Ud9ULmXyZ5gXw1HiKP3lTjYJAvz4O81jrdrHWggJ
8JYeOOsTzJH1cqcCIxfY0iUpWzgjFDD78ECJSCaH30XRc4A9hyEUhYU4IR8RFqbtWMq3PhGMNYRn
K6xQR4Btz6DG1/wGhmEVBGCwV0ZkwyIqXFnioPjjwyl77dFgt5feg980T4itti5VyWgJDp/PWmFL
7syDS+4qqPxhKAsqFLcv36DH4etErnP/Q8wHvP4KstpaXwuoEZRdT7rtlWoxBZk5lw7sRlec3Tt4
uPvb0Ldowh6s8YS9MGywJl51sCdSgKTgI8sNB3FBpS0yA98LYcEV+dxeEzxnzqvFIZTAdTFtmPuJ
5gC1IHYmeQBJqWpnN8uKa5CFIHyN6TqkhFxUzXi0s/XAYaN2ovSKue0xwVBKwiQ7ugEmLQc8w8mM
h5lQl6qnh6nzyC0URdVnywlRwKt5lu2/BDag62vX7+kk2q7Jr4xjijESqJ/JQtbMaX5LYYSp12qQ
VFTJBc+2t+sKDGWTtazA2+E2Gp8mCao8eHfUDsj26ZInbQzfQp3xvvdiXZgzig2C+a5X9uAAo/oc
KbWxyCjr9YE991MPzWju9V6QQFX9LatF491u14MQWq9xiSEJSjms9F6bofz4E0qqpJm2YY6m/C4I
9scGidLx6R54hiN/KApL9eSLivLudmZgSi9smBrI3XBekQl160PVgK9t73f4BJw7GxPyeAr6ItGd
/q+DT6UwzxX3r9HVoytgnCFPB/W4oMnblDnLi/PNGQCmbb2W5LJtrV9KEQp4RgqpTsyrQjM1UXk1
wTW/x9F5zTp2nCOwUq+xF+DqY3iT0Fqp7QJlaaTaNe5JK/oIF0yawhQZJ/LrZZjkg5hXwLf29BuX
TgNyfDmjM58lnrHQtzoucwlkD3RBYF9KQSFlc6R/els9CrypzKhXFjtmoape4DdAb0u1Bhc23/5W
tOKB9g9WsPbED18H1wL8WEuCovHZp8Oa89Zsd55YcBVzmdF0ViRXuBUzWJQpdarF0dQHyebOY0hV
sGrBEFWtawGyRoYKqI/UqD3KEbw0V9bynl+LUAyNnnSGZkiqijDqXihQIBrMZQKANpgtIe8yRRO+
JAZCGgIliXreRmkWv4aQAIZtAszR21obz+Uy46vXd7nHd2gRpC50OEVthWz1263w5nzMDB9bQ07t
4ttymcAa+dfpOLbd/Cs1Sew9ad27VNG+9Jz0rT5jeKZGATXI0r+iRZ3ht+rhdARXa39jhTxBRXG5
q5+K+GK73/ruwThE5lpNy19V3ooqzsQsk7gzZl5glQA5a2hv3DCjlXsxzU2quQ/RnyDj7d7sSqYs
nVEah1e/tOUoQ7p3GfgdUE1hQnVu3qiZvTJBM3OvLsSMIo82FZx4uuzjyyudYNO0LbhUxRiKWNca
LoC+CxjUk6Mqi6iq78TFX1PjP8Gj/mY4OSSDGuJM40S14EaCzhWJ8GPLLzDHMZpihUr7PwMJKyjy
FBLMwX7SyQ3okcoADlyUbX+RTqoxTh3LlZGkj2SoUAERgJvKWfGOBqHjRkueTgw7EA676etYk/7O
Wy4+CmbDWz21vzkXiDRjEGraVlM/5ZKDBxF2ffjG9qc2lULUZgzeaa01bq13gVlnrAtd+R28jOah
S4pDzNlmNuTD9x3mSjdzgm2uuT45anBfXNnXUrpPFMDzaRPeYioLlxdyLwzxv7SQsNs0ww9UUCR/
cB2MNDRcB+q5kydyvrkvRpU0CAKCvM9vGdPdvGWNKRimbe6ZMfP4XrsON9Im0gWUsKB6g/UFZ492
GsfM0TV34Zn6RVcL2Qr9RxoqhOhRiH9Nh9+rdSc2XFN4ktdOwGSqCzf9nY+jF5ZyQfhv/QY5kOw2
psObaeKAtB+JPbJVXkFgH2FHY99tJHCZHmUoO+NETSKfCTSkxHYW1a+ZGnPrABe19cWSDoelcuMW
DSl2aJJwT+PdgFw/bHTuiRPDoEIfPaU80KlMaefoPEk8RkzcF+5v4fnm5XmZRy0RQSNqnwfZgeZz
ITETVth4d8RbSxJfwSpOaMVDs+QtQePaKm5jWDe2RN7RS3AmqlBV5mrtK+ne0QAuYSoxtC5WypxL
mfUE3+gKCucX1LZ2X3XDwGYdvZT1z4Ig2F5nsfZ+nvYSFuieQzJBaatZta60k7Yb1R7/iZrZAXE9
eBaFVOe7pPDeT0yCgpQ00S1BMiVp4bDvR9ZQHhOdrM6jWP5vERHdmqgizYFxiZ+0gHb2KF7DW1Jl
ULnpkjfTlio/nKk7RlO9aZarwB14vOlpYQGdCspbr106zzoE5cuFeReI3opja+qkzjQfepmGSb/7
mMvHXO4BWtOroHYfe+LXRd70e5vdwCxdL+Th8CPr4t0VSa5BhOcoYqFjN0yEjCneORyWFInubx9b
eDsCA6/l+deasFNhSxhNFZqGS2KB/VrzCnjRmjgq0RJFtIKF2zJ8mQSy4oR9xJUCU3BBY7HLafcb
sKmDJz78069G0oVqyHtblQ4BGjgEcYlIoVcAkqLiryEQogWiU6y2auXE338rBWTUpxWwdV64t3DX
iMEwsF4VmUBMQ6rdh7iypViiQtjH7HOtbOOP8JZHwZvzNxuYu/U7RPglVaor5QenpImdfci+7+1r
NCNruEdPZGZTkzgIT53nEvoc53T8rdv7a8kDfuUlu8wtkMrGDDW8dbAIoGxm/bRp251FJdBYlJWD
Z2N4wf3rKIA0b223rnyx+PQopvaNX8ly1z+AjgIQw2ILQVZYZr++cZ3fJg09PmGf4yCd4CL3Cr9E
FOz+lNUQKORf5CgBR3PkSJZiRznF8TpoW4etY957ozJpSXoy/qkmVARMgVxbVvm/cnhb5JdC4zpF
VGFb8gOxAw2WLv3K5YCttBCnDgrcFALbMUFcoXXXFJIF0jb+OnmSUN47ht7ADxktMgvJhCugZw5A
eJ//e7ITRtpy8CLSrmOilqNFRHg/eCL0WaAuEhtjwN7Ta7XA1kfNFAmN0SMdHgb2o8WQHbr0oNi/
YkK4wG0DqAhL6pLdFubNVtbjEd80KlQqQRLJLs+10ZWgtF9iOjK8cXB0acuHlwxVq+3lLEWxAXeo
EUkCjo9sa4qOwOls+sT0cQHK3qqPYfqxKt8qQt7eMkFWixsbMKqHsCMELcf3fi4GALC6xUjNUGSN
osglyPXKwrRNP8pmB51Qig04in2pbtOXMNj3RW4F179mvM123APKSVFrGHeAcbs0lYdCcVCLXedb
lvm/6Lx0kQSCd7+Vq3YMTkLGnWEkqnkWOl6rSpgvwAya1h0tT2z+hYSnR/jUZv6sysKe70XROnEN
7GM9Bd4aMmCk/bnYhnQB6iARMSwPMXkxpog12qaCrDdesL+8R3cK94JEWyMLCdt+hiJO8R4KuVv/
eCXauVwC+h8zfkM5ok8TtOGoukO4ozaAqlfWOy/vxA4eW5mnJCpCEQ4mJBxl+/uNgal47pQkUgMn
VBnX2a/RjD2c4jYrbAa35PrHqh5kLo8LSs20eP6p7wdUXS4ndpCnMO8iC5dInF5i+aDfr33HzUbF
ehZmfKSBBkB9JnUouYbLrOokRhSLmMElviwEqJQc67ssZnd5wHwzru9jWitOnKTybZ821COAajkz
HUvzDFVVLKj25MVEyoYJ1OXHcddgDzAbWeFNl+ZG++SWw5QzXRl7q55d8xJAEgifZ2SsaQ38rOv4
eS+uCxHZuIU1oiJF2rJ+LnhJMaevgYCsy3NFvVHcsdTShnImb8rfC8YPo9hr4M4nMV/jzmJ36n4h
YpZSjb5VXsflEo+7fJvCxbpDnwaH4O/4LHSDQdlZPORVwSBA6Qe72n4ajjDk+0rRiV8aGmSDfvQB
ybGCaScHishaCOBjaTGa+/BgYyTvCLgj4ihv3dsYIhLRlQ3FlBVpSDD5hLdLg/199lCA1oMGCXdo
2HW82pDU/14scAnkuhhwAxKnHhKkg3S5OEBtWIat9Bh4L9g3nGbtmrT5VqFyQX5ihdmLzVLxni56
HskWf9xQ3uC5YjhqEShiclDsHI+GbzZcOVr6QWE06D4IHpGdcmSoFP8d5dg/gsk7eGsL95KNRLjK
8ykpUtNOdPhMjdFtMX6U6yl5GycLn+S3Q3dajzrA1AO1tkAsujmM0Ma3jjfqxcADwO9AZUVc1mzn
g1MVMvZ5xVaV73NNZHPrL2SBGtb7INnxABcbVb8Z5x+bhBkhvlD2Nwx8edJ9T5GvPHtta6dq5+R7
fQWzTUpVmytpr5PmgrfVqf1y6r3DydREaXRY7OPn++mnZACbMc3+XSIdtddXWjH5Z2WYoGjVcwHl
3ZTJ89c/jXLahLA02hfoVyEqsUj39ELd9/QqMcmnQ5QVEWhISZb0exPvIywVZUVReyiBiCBxDNM/
uujFntKUEprOsWMVsH/ia3txsgyqtFWI7p2pIFdfzgAsBHc3GaAd9NljH767y9CIsBlTJdygH2xg
mRhMfR/unZFxlWp3hbY4Vn4ZnlKKtpQQLKgSeSiRVjKgob6MDJUzMfp9ax69G2S1m9u7ldjeZoXF
wG3HJ3D76i8zL+Fw3idOM0kdVBXgvXV5+il4rlZEkJ9xt1eplhSgVnFGVRuAb5l7gd3gyefopIwk
wjexxaOgIjslzTIFUsruaD3xrztGuPRnhb3BiC0hV2zevV09jy5kgCi2uyCP62S+2evA0QQLDbCo
VblPRfFcJiRXvE39rbDSfMUsrLe/DbQvhiczD3EfckRHMrLRHjLP9CuMDgBjlEpGZI0Btt5WWhqu
Zp+Ur368nW5yAHEn0tqVtOMlhcAArIgUTp3zNY6x0vPzjqfOPO1kbxW5MouF+jmbQMG73mjqnRDs
cJRjIsnXqZ84MOh8wYspzRMNG4gyNPXhLs3u0mEXVXRu4y4CwkAAWj2H/dIcgRicwdYBbvWQG92b
+icZZnoYWiaAehz8dCqoW8DzB26Sa9gN3ZejeU5sL2QBdpW/qZHrYLXbeCKUJWIijtrfMNpeg4iz
tPPwTHIzbX85Hau5qsxmKoUV5023Vh8D5m2ZHbq0hIzmd4xJknkFYIo2cqZYu5/V6NY/jdmO7CMf
BJmfqcsqD43J0eIxiK67/iS5fvr7UAdZtUq5Sl+Ba8tTjSqoVqwAs0236zshHZUAOGOSQi8xdt3u
V34Ug7GKOPwfjWLGRdNKg74DCM5nKPraQtrrN2b3IUcen9G76Fe++I/7kn1Ay+4jMPFo22sBN+qd
G2OWqEKYGYX5xA15xHDNFz4vFLOxADO4h193bEozrAp0e2i2S3IQXNcF0ddI0APgGWvHi63corHX
xqiCpDAXbLGvJ7maAE5h8d3BiseqqPx8HBUfhHcSjwHfdANRrd+8u2cc22hT9G7bxc86t0SXlSnv
6TWGwn0nfKl306VI9fhbL1u65JESthjnGRD93iRNl4ecgPZ484e43qmA6k/9JyY6JOJv89pNL41C
SjffDpjCVDjy8YNxA1dfaoPRbrcObWdvHerJWzUT78FSK/++TSXm2MkFKYPoj9QHVvh9HDzmLx22
8Rzdne/woQZ6Ro3BWQdCF15cKqF1mIDhzVvuLo9YEQXgGjFFsqYLUjq9JMoOs+V2ugpB/imCNf+F
Q6zFpWp3vqB5xV8L50PFjn/nC383meuYXEs8E74sVQ40/H6wQORh4cLWlhnxF9sIqGrKXob0/28y
IdI2qUOLWpqZidi6m2978riL0rJ77PYGJyJrkIBUMNA83Xg+JwuN2WY8tyZQaiNQS8p06GVk7FwW
2bcpsPWZayEU1pVEgcuk/uIQujd3O0Vl832kwH4KSORamZSWZvU5CX3f/o9ruj7M/wMEkytSpTm5
fNV12vC/6Pe7MAazv55bBbgFQexwBgJH+pEmCKqufHnhxCHEOvn+9U6AogU3AEfevlFuQkH1yz3e
1NxDWgWgOC1/n1T8+cxvUoPuQS3+1/Q2mlrkMBVu0s4X51AcHh9Rnt1aaic5tjJouhrdlZBLcHN0
FqDKGil7JrbFc9ZItD9/uywlecp4GE2QErfWqaxTbUeWdlmgWffrgPGGqgmp7ZGaSPvQNZ+ctgmu
u8aubVO07CjlWuHK9odbwvDoHLCThu/fltsvjk1ry/qTllG7qajZdtFkpx1RzmhkrweXVyDSNNs7
qrOSxoqPKTXldXj78GFNZWXj90UmzGLxPD5qI0MucIZEFeeEXHzKLcUcxUz0N5utkMdYKaO8xpU6
XsU0HMtPj+HjwabB7i/w6WEXajoRkqXzgyLCQLZRTNQdPQIcK5dJlSDGyF1fy8ZKUP8flRh0x8zp
24glEJDy1a2RTzQz0IaWvkICz/W8N6qKfL5/A4pfEVwLeud1NjHE6teHETRS7wJnduiYET5wEQ8o
gCZPDpSjVoFcTUlEAN0v+ChXk+2tNenVVdpgV8vU4qEchZRqgWpPcq8G/6Dtwg3So/irkIYWAWpL
sfYNx6BEW80+l368jr8NzqZ8QO0ac8RjazaZxWDJ3ZEehqxVzi5ZSl/9TWauNJY14MQqeRSsjtrq
IKKt9ryuUbui89xagRUjDFHeVl6CZpaUwQDHGr77AeNQABhsjcGF1WVYDuPxOL7atDRvom3Q4G5W
kGrqAUEV4JTzvg6FZfGWR0JWjBiTex1So0DW3hQoDTlaAgjOmwGgWMieWQdMlqq3Ha2VdYYwUtEL
0bmW1ZWqJ4UqVvg06TzI+btxjWiJUXs+u19Syfp+p7iHDawA84hja9ey7Rp4R8nTOu3XTqFDa3UB
tRq968JC9dObfVwFpcR+zXjGmkX5YQV56XWB82zSp3Yygbkf2b3LVXmPkDtaMAEYW+drILl/yp7Z
XCy/FXvJmubmctVlovQMy9ry0Op81gsz5doU0xp4BIX97D+qi9+90relrp5FgY63zTeBNmi/SPBF
dvmX79CeWswWT366BUcHZN51A8WGx6IvVWPHMJKaN9kD4YM2sPLyWuBV6g0B9Dew7vSx8Ez4Pegj
2lAexm00fcQWc9wJCVraYfRri5ayqUn2+Oz1Zbcg+wTYNqK4XJL1qKk/fu5QAgeff/euuLsc02yV
rqLqEzOvyUK3GWd/W+5MzmC6I1r30mHTzk7tv3x2gauZMuxjlVss+7Wt0TkYf7E4MZxUT8QsEL9m
yu+ODquKVfhXiQy0eLehZL86mU6os+/bGHvE3t0L3ZCeoyPsACN1tRirRnCSm1xCykCgXQ9llbkA
V8J5/uBorJYKK2dp8NsOK0WAp2GgO+DiqiM5rPf0EjLbNLDowKfpSSS55/07nfgmwWhQh4bf0HHN
rIW8faRvSPNzgYpXq1eoZav4pI8cZUnJhyyQwUItCLkdunPV78LDxEP0Fh7zyjvnBSgjfwAamJQS
Vzm5DAJezhn+bh1uAvOWaySRUNj2nmsUw/dQMRthrkA7GMaIK08BhOWTRzaE5wtPnHGk/XNGSKwV
CSdcLMiWhx8mD0uk3aphr+df+PDAUbGYwmvoV8Ahi1sbNHpj78+baAUA7O3jZFeBf2dj09XOP43Y
UZTFxz3nSXPBvhP4x7LoK7ccum9cu04bo5NFzCP0wB19AVatdKIsO0BqJeBDPQJSdw0U4TkXUz6I
K9/ndxePqdkYRfwAgqE5jZeC+nujemQjGAi7504AVUruXMlcgfR0ml6wO481cnU7ioC+Re5FRUsg
bcH56WlYoKfQVYaOEJlPD6a5ZX0Y7Fk7QKqW24yd8tGztkPueLpK4akR39tUA7KabEbMEgvHO6vW
m4UQadOVCci7SJ6Kxi18ZnSCr49oE/sj3qxK0o1QuY9RN1XU80vk0zoSkpELEevx5cqEwe06k3Ur
Yd+VgieWJhve79WgGULJj3VkFCJk0qcZrInqseDyeeELhTMgbtdD0F1bfgM9ht9P0Jf3+LSFg/nh
+JbL8/2lSP0BhdrPGTDycBOy0iLWHn4K5UY5s34CU+uWK82HVybOmKPOIEFwtlEhUmlV29NFgeEl
JzhszFDJYX0/FqOAQP5JRzUK+zi/dIf/zgHM4tN5lf68F2qCnf9lP59jQhUhNy1vCd5zIG+dknqQ
9fwlRIpb8Ly47HlC7SsLGlLnPHqcq62dnQka2Z9zgluHUA7MuoirXtcGpHV6v8dMwD7kCML8lAve
jDfTIYrZPIOnktZdchqmAbg5JXDSTsaBAukBuwqEWY5VMiOssUof4sycl8/axcUq9JE/fRkV5wDs
I/9qqTesh0TW8WcXmyn26vH1DVx8SYIeO5jvTUGmF+cCgPRV1T9ImVTQR2HdTvrZsFDMsXI1gOGT
AzURzNRC8J490DOEPx+A97+d8K9qvXtwYBtRS2IAsGZPxBWRI5j1xLEb//eCouICjX/U3dW6oUrr
vZ7GR+FtlRhDySC/ZMiYDDtoocDsCC/v7ymvIae0v7ERcJl8b6VDoRrjBq7OLwT42DQBGgkFhHOo
riVK0EZ81WjgjKuy8oamOj7AWx7uhxui1sKc5vKavdHzDn0Wu45mNPdG7wBvSSoFqOHe+bimAXFb
/VVcPcqMDmDqFwRCRlTVeFOO5sn1b5lwZOomNlHGL/BYWIf7OR0Z8a66GjP26uP1ofgrldLyVkb3
FZLGLTagdSqWgi35+QmxO6lDxpd+4evrEXCXW5+GuWzEv8k/3tXt50HYDWUe4rGgHw+RavQ4s+iQ
qPCCRrdSxnjAH92SWKxQjYbmkSMDlyXwJ80v8pvMCC3DnQEkn0Og8wJcocJbknVCwGV9g/6Mrj2Q
/hnzRVuk9inYmlm3SN1pBvqMx2qXJtjFgc7Woxq2uD24ymHTdFu++UwpuYKUZmtATdSt/mRqhK+x
aRTyis4ZXXOMqpkza1IoeQcZ8CG/s0+Vq6M3fH8J0nPo0qYzKpDhvXNsKqMRHpZZwno5yGerth0I
YEnnp+oAx/A6dwwxvAKIPSKtfFbb22OfNNqcYZP1arXq21BAxD7/cIN7Kg3g+REo9ViG8Yh9vO2D
+a8KAmYmTgxGPxFaCHqpnJn98wyocQhAE9mzExZ8qzWkhzVvNRlTdLk+OhA4yHp5dsslxz+yPsyl
kTh0WauIJYX/SbHpIjJywbzR4B+srRFGR5/txlxHjPm6X4lO/zjl49VmsMkuZenuhvF3krJUYcdL
TDPCs/XfmJpEXOfkGOw10ohS7qQZhUq7qjn5gQ14zf++nYDUtJAnCGWGVBja7wAROVnD4KQaZIHk
61Xv/vO/2s6sxCBuxZgbBFX0Y38rTOHYw8vbd1fJ4cxRRWni/Y6s8VzKFrDz8T6ldSEf6w/+/d5/
oYKILpNxt10wbBWKJWbdQ8fFoFQYvYQ+9En99m0uMjXZX6ZyrWipqu84xK9WaQp8mLrvnHU+SAor
Mpfk7uo0TGyk7SIoIooY7nIuRMe3yufgq+Y16BhT5otuyaQgVUOSCPENFwQBtBvhlWxlHdhdqlJG
PAMzFYU1U5L7cZdDu5QB7sookiVMmT6k5YpiJ+tcR58SFZKa97/a5F+AgPm1Q0Ei3UhZzZ+/Op8t
HgmB6dYvs5Ru9jpwhVqGD2XShKri5CgbXa+jqNBbq0+nJ8uk2zkZ0fuGBWn+/vY5k1vr7kJQeXZ3
48LaBsx48bQRCSPc5JEpuQzfGtR1chksJMT8s7eRArxhc60swx5re56fzOWOKS8Q8fLKNlefnh/T
8NBjgRz2JmwcYn61TKG8tenG8uOPh70wa9iXFA4GHLc+tTEsUyfQaOIraORTfyT884d40sDs6oOV
aDTvLSg2+v0unHsa7QkIQJpnmBrQBM/okVl4yHplON7O16USjo2qHa/pUMYqjiynmTni+mCDBjgD
dGZ1IVYGBiHu8Me9CEb0PgDmzTbGbI6weYxuH2UIo1ulh3cuIqZOiiw7DIMTX2Cd2NnKpgVh2ZNY
G3LuAnL8VypFUxzDaw7isRdEYpzs7BhRJspz7LN7u/6o3XtTRLE/XegvTC8bdzW2AAY34GS+ckbp
y/GmItWItVm7DzrgxPniDfPRnrDGdtJ4d5qY7OcGP3ddYbb7GSBIRR0vpoA+OeIf4Pe2YfrbAMEP
sj2Ua5OwyGYqGI/AHnlGkwKwJfGwWS1SRRqTOugCzc8yI3xKLWbgQybrrqgGr3dluI/KW1sHgOz0
Aw86kmW31dhi9RhaCxPFlf9/snosrRBmkgoRfNTWZCMV9n+1rvEQA5Np8Kqefj3luB2LdPR/UOGQ
n82lBulpsf3ULE/sqDYpNqzIfEPds2f4gf9AuonSgCKaegteEI412A4o0sHFFzbzRBqZtwHy0Jpf
bx2ynHhtJSx3eJl0VuqdH0w0JWmAuYJjNBKeUixK7dJbYSqvdyQtsIpyJdiCJP+BWG0Hg3gDW4Uc
OQOSeeEb7KAmlluyZ/VeQCJJ6CSaFNuMtFlMoW0kY6TCtUX6HDYcn8HYlIrl3O9qzHEYj1SAFCdd
B8lGzmepFAXTx37nMZaZcba8cQjEUwPIE/I3Z0ZIVSaJ1vYUr46L6uR3pvphYpL6n5sYVW74Ohnn
kylI3e7yswbKNaW4606URFzpmtIPjDlGexDrSLF2XrZfFwi/1IgIrGZb5l1LRo3QZArNi+TOCQSj
2ycP0l02xGZWqHyBTYBNLtyvjnto5HMC5pwvzKbh1fpSFJmIWzICfWeQJZ2D06iqY+6zkVCymSjI
3MjUz/IaDo0XPKFn3CM9ayTTZCqI0nnw8X03U+/OPc3oUMo0ppMN4TK89zpbxb+V2FUlmXhVbaRT
977NfttAJaJFYlVX7Y+hd6/mnbZr7H9y168Aa6e6X/OgayQVu8wTz0Nxw45oBbcNzqh6OWRH+aV6
QQ5WEbopF8PNVrPUqSdQX6D1qVTuS/7Z3DsTfDMiUpjY9L/5QszyQ+0586h6nCe0fqFipt38U6Qn
9tTSoCJVp6boGsKrQGFXQ1PNRIRhs350833FXWYbe4nQsFr6bOCPiy5BCrHrOFm8wMCUVrhg06u2
GEmAXFudgYISoz/BbbimWVqd/4wdAZsSgW6YCyj2lY/tuyjf0Jwtk+kFoBYoMWbZWdcFfmxnPikp
JOzcS1BEEylXNZSG8JH3MNtHZvvQrGQKDmn+F5PkqPq1LYHJs2rHsIcVPCaLbsxH+TSnq3HtfPK2
VNBCbVQ73LijDUB5+E5qgwtoiy1WYF/L0anoqPcw30OqkZypw6I3hU98BaUib2ucVUJCd9HQaef7
TA8jGS3MFGbKKPq4FK0SAnOIrroYWPgJjOhmDF8/cXOTg4/Arr3xN+qYKRun3Ch2PLPcpqdkT4gC
iFpiC8WB+iQvaJga//c50w8diIbJaeBf3wkXN5zrvBs7gsyxKLcKtLQpA9GjLdyGTdqzvjWgz7lo
QhkQ4CyexpzhsZcM773hy1b7v0Td3oY+8E04/J4YT6AJq06j4EOdPzKGJEnt+utBKiQvVvpYIsiA
66KNInbcKQeU/6EPa3zugfuv7qApwNh6VJkQBduy56TlHCiQE+Z6o9dIabXkXZSuR8oVIoG0VMH7
yAZQC9O0Vfh9+oNPcqgmDIlP5xw1tSRCNr+wrZoNPELvrX0SdA/Tbt6ql314DEk38tauqGQD2iaA
AyqVrPJXP1U8KGvc0pKOlSXflOUm+D1H7UOptR/AHx1lGwF9pfErtpg/Ko9HzImj/Y/bo7bWRRtx
vliLQN5ZZ/jrqWXrbLbEvbQGLVGdnC8qtsAlN3x8xtnAAh1m2znV6RO2KgLvMopgH42LBerbgars
U+Te60oqkzbL/N1p5WEmKm1ESzi5WUMoHxRgsAiYrMiBqIolJWB49difyr0DsqLqa8KF8AZ5OAxJ
IXoqtWfcfixwvEyP3cArXu+kqauNWR/v80fC0hxzpctQtD62yuO+c9UR7S8I/NBHYCoKxNoeD1tB
DIXi+r0BGXgzGYf48Fxuwjb637RwAf9vFAjeCRzuxyg32BSm4qOwgrvyRP//02mbbtstJnk5vljO
9VrrEldRubvypV22odTolNBbtxJujIWB9T1H4qSy1FP8fkxcgDjn4siNkYsbZ7OfXHlnXT7GfG2u
k+Y8D/44iPXwEV4exlhh59jbCa/zpMrj1pXYjwy8rvpI3dIH3cSeXIu603vds7FMG87mPFB116Lh
3in0nLzqoIbFjCHmFHUpW8MUuVDjOZhjoDVWcsOjXG2iG5vivpRlgtYLYdHJHBRuosE72SHaDX6V
mXH9MXpfwSIkfiJJ+tJNf7ZC69lzHxWQwL4CYoTtveVqKYzwmTaVfvMtniswbw1/H+brGhcP1UkP
CUKp4zQDTJrX6SiZ5ytYpTNjZfi5HxeRkzR+v5xfEp88bd/CQbi/QxCYq5Mee7kFSZqyZREJr3Pu
ZmLgciSEuu9R7WAAhAjMzk8pRyEHtJYvuU3gMK92zkWXsXg5oUSMLajrqespUUDfUov68t/4nk2y
ypkoVclFeDN3ws2ITcWLFhCgjVz4cp0KRYHD2PRb1hmsjH8dIR2H3WbDMBuDPfmlU+RaJDtb8WzH
4l8wuFDhx8d9xgWb046xQI1oVfqen08+wf5YC32E8+4qkA1PpD3dukGSaKe9zjGu3bztzEBJkKT7
HyuneuOEdO3PbW6+Yw0j0IH0ILdTjP/n48gtnaQymEKQS798kEf/kvB1GO4jgPTZi4qDVgfPBtWE
jgKu18tpvPfmCVpxpCg7MNR99c2OB5meM7cjycfqdDtnl7pcmqPhRSprX++9Bayhyq+vVbrhipWa
0jY2HqKThNBcLYeInO4c/2mN+VuF8GC4Qn4ZoDiJUW3GQBuLGqbrkTH5sjPKU4APR1Hd/LZFyl9v
CqqhDwmzh1iRFhHQx+0FXJx1zkTd/GWQCtsiokpKBYTOtpnZxeoh1j8K62YONsrIAa/O0Rr6T8F4
+6BtZN50ZNStm7Kf95E274zxhZ1OI4d5zqjpdUJnBZldi6FxrEISREnX/2yWS1SLOBkz0sW4bsIJ
y5eX4ghvXsquw0bhmmdH+om2ELbOMUrkTXxf1Mj93xJyLma6E79LCpov5niM3eaRsdSAnDuC377q
LLAMpflZ77+iQFvjNyST5qYKt87n74ymUu7/Xhdh7lVDspbHq7Qw+Hraunv0zZ/+dvsnqi0TknOl
wifZTSMk5cnE3qQuTld8shw0G9HzX7sgVb6yOtqw2rMEjInLDuLJge12MeDYcq3wgKbWyvMtFA4B
DiBGtYYDVmM8AmA7XsLARWrsCkCXw/XtPste1/ibvj4WAWKlP+bDCu0NyZ2YWzQcRDLoiFljUata
gT3WqEzaYGL3Dv7GF2mb7pRGVRAAk2YN459YUthrXcXpP8cp7Lpco8EmvW7Zwjq2BHZnzkP9DA+K
Z5sruJUy2XAheJ1pXTChHpdVnYs5LU9OYBKhozA+OGRSfqW2t3YQyFZO0Q439lyKxUUkY3wLScVK
j8LtWMxfVM3+la3pew3aeMjBdF+xKokCL3bm6t4JQ9kNJHE6lyFaWg8De1r8kwX1Q+kCnXMQGGi/
5ehUrTapfNLlYbU56QhY8LKSxK/nt4B1KQdeur7/orZkifOVpF1h5wGYqkQIA24Dia+vI6twETtp
0sRsdRFbqHWfEbSB+ARTEdBh2hvTTVxggeGZsRHhD+QkpO/dOwiHz5nT5T45XCCvZmA5imU+S91P
BTOoTtajjHu4OzIHI6zZDCgCmEFoZt1opROLBj7LgN3iD0TDUQoMp5lwNUbjeYTDk3NmI+9DLCAD
O+E5gVePDT2mtY9EivNoNXa999ylZIttjwpWwWkDingwPR3apeSIgqMCzGJhZDdirw578bB/knaH
g4w2MCkahXAWee/rVXz+U9sAeo1gCSU4ZJIS5J0jT9mtAwV47eTCWQOPAtvHQfdBd513BolTioqm
g51uFWq5+KiYe90dptvJfi8yvNKjUL0ec/tRer2GoqpGDO8M4Wt+kgjLUUhVbXVklUgJuNks7b5Y
C1KYJ2RepKzV+ua0Gskjl0G9kdek8PVNOBYowojcyM9Mk5+zA9hDhZqDraVzsly416DOk0TkoOKk
V3+UzkvcRjEn107fs3Y+hPJpSWCop4yV10n/Qfc+pKG4BxUR6KkFu4N5RdNigW8jY9uZwOko9e5N
AEOIttiulVdsKg/iZCFBvl+WKlWrnIF0jxanoYLi/2PzaeDpBetZaYwT3fxeOxe0s6lyE5OZIs1Z
wTn0ih8SL+5GTY4nhFaymaJFpGWG6XbBWmvOMGZQj0tnebsrM+abLmEZS4ahkGrkunycWbHdPrm2
3zTHr2Fl3oaqsnxFKlgKFassxAt/0HK8tKFxVTA5bhZiGJkiEPQLJWMFz70TuPLl3K1Roz0qb40H
zWPowPMpxcjbe9WpMVUYwVSZtjqsLrPa/PX6VzLbBCgeFUdpR4GYPpxekFqcJTtHx3OEl1Eekf4d
U/9v95+EveaBBdGFWGRiGwegCLafzSUno8zEHhOQle9NA8zAg6uenFRfdgRoOLMHJCAqedFYpOK7
SZk+JrAxSICZC8swunCceqS0TZ3b7B7dFNQt9BRhMAsPl+RPxBKWcSvaielf9KnfD9FVxLRGbQCM
SOfNWAUu3VlE1yA4bZOMO3vxY5qBYq3OUFN0DtxBpm+E4zNlflvAoqVnvDktgEFXpXFulzwEHrPc
wdTHATfW8fI2Cjxl/lAkp9mtcOzG4lPvZITaeg4hGWrroWf5HrtXPirGjFFfkRVwB/7Hmb7914WG
gPHlNi5O130TMgY1L5Hq79IvN51Ct7sBo9ZxteaFRa2lABYsAfG3CuJgEDlvfkpZhHZe5cytnInD
I711sOAVO2QYmdqEKD4grumfOg+OFR2sTsuyJsGj3kSs7KypnWSfMxUTi/7vobzJy/gqbO2eRuo8
AKNJdgPB7wJqUJYPAaQhNrmrnoZo31Ua782TjTzoJeEnGaHWNR9QDs8IuovxjHg6DNxtfGI5Zz+C
ZgzLZNKrLSBnk2W7fM9LgNLp7hOT30wPgRDHKWcgP1gM7ufTiWAPNd8mgSc4YlGplgKn9ZB7lpYn
RRjfUgblm011ra1+3ZJ++hDy/1MsV9OYzWBX5LlwELT7qTnXVv2gvo4hksH3rB65RKADiHyFgZ02
pwRGFaiJSogfW66Ju8yeergfbmd6uPa4Db4wpG6tSHq3Gp/tjH2kQMmdFVkPQDDEXVTBkg2VJYAk
41sBeM2bxL1fAa5JhDg1SCyOVzQKrilBzt8yr2V9HVD0CuIw4NyQN17mnuztzOO0WyH+kIWgD4bm
EJyVs/9Btpa+up8XwH8NuvpYe9z/XNyo/uuLMI5vfLtBFsy+0ACR4Nn+kmQTorZFpth8X/RhnDD7
oCwQyaq3ZdfwegcKNT51AVrEtQSPcaXMOiehWmjIxgxAA6uvic4NKbUpBVVE4eeLV5OLcJQrRlzx
Ph73Imi1MZRLtTn4fyZF+V9/a5ACQ7xK/xZQhOSC8XkG+Xhiuzd85dvnyBffl1Wl3O++yw1Stkct
CPYHV8hryaSMgw6QPGwt+zhNBb1qfEV7KfFNFGQbejGyOwKtKhHwiIJYOLKiMidhba2jeN36nQ70
eYcH5F2YjwovTpTmiUvEwFcqbJPhuIwnyCWC9c7pTmMoVtTOhblOoOI+6eWob31s9g94JTTfomlp
wix71szJVWCrd6xvFop3ErqqX48LrFpTHNlTMfLdJIGTHGt2zBeg53yIVTDp4MAvuLyP1GAsk93r
O57Z8cX9GNR/DuBklarZxPpSQcst/z9VWw8tXG8E70vlET/tML2Pz4pk9XalK2KYbreDSdDb0m5h
PGTgkf5z93Pd1nwu3ec1T+tFTexbhJnRkYPWpXYkzHgxKVof2ZMdIDyI9lwrbxTxsKyJsi3ao438
+a3477S74+84ustqNtovBmldmXQGHMIplIojXYbsqYSn4wo6uC/OxI5a7eTM1gPKdxwN9UigQjTo
c11083XyPFi76sA4po1WAOrswcjC8BYKHAdvMoLqQGZMuH0ULqL+8J6e5TzaPDaMN10CYcnExHtX
0Y6Ddojt/4VAjyJtA2P5CJS9IrKqER8q+teN9z63b6ROtwZgzx44MWe7LBbahG5UnS113SvshIpb
MouUA2sAVn8FwLm08dmVdN8KDvFeVYyb2YgQ4lpLEdatPldlbUKpTYWSP8pNtsBioUOzwsJwRQCm
YHZ+hvNBT7xYI7RATg9N32Ca0ckVeZ50wV+525WcohfUFFqUw4b6ZwnV1cxH5B/mwhbwCVuac7sP
PGvyomW3A48/zaj6QyMU09a2mGRaKyuL67C+1UDJ+NCTGmgOWkKN5tzbELWbN5I7jgD+QCMzJ6i8
yy2HHNBvXAbaDX8W745mjkL9IoYDVGVLCF7xWFuWAIXGhVkhdM7cPvvRdndgkkJQwwtZgnGMu+gF
iEffSTGxmCjWbw9D19iJvNFPQZCj8GokDIox11dLzSb8w1K2hnAloFZL3PGV2ZcBNLWCYwUJkKL6
jH3/C4fZqBqjoqD8tGLN8USe6/+h/1WdLOj4KuE7pgmcbnnMUPWA1QYXzdrMIP/B7E9e9qGXDXv/
2/MAl8KeXWczDHB0jHT2Zs4T/ATfVuYlvU1styW4w3l8gvKomSuee96Z1/RFa0zFk/imajKfpJT2
KnNEtGwUCzn1OEUfZHH6PqMJMgRtpEvs949zt6LfPrgBRPhGuiuaX+O8AG+RJ4hdEu+Tl1fJ3xyl
LL8j5KPSG99tm6SxoJ+gFjvsVDfS73y8DJ9HczduQefYSS58LudufaMSd2dPdO1Ojxn0w3eCbLAz
MfP6ZucLj3kKBwcR8elcJMBxzecKlrBrBuhrDHLQDuOU6GurQV2jiD1nLfMp6uZ9+NKCBG/HEl3O
pdL5YBUWDj2ODOQaPrgp07gSjuo54eVpkxsKPLRMUWKPJz3n+i4dI+GUsJtChG36NPQ5dUdiEbmp
IPcG3R68Vjw37FzWXdCZNCprxyMuKspPtNr3iom9RV9FFzgb4yZFZZ2VwyrCAz2K6jLdrJtc9GJB
STU7acjYeUa+EkaVHnyNMmHgBVgRw0aJt/dEpy2cyKOz18zkCeQ2QBfbRd+IwizjEDv70v50J/4S
vmapWLII9aK8dEaIJC0Nu58zCeDij1QtQtpSyEj9NOOcBpOOZzqMRh8augfTqogVNYY8scyOXDhp
yobtIeTzWPVX2zvZvFf6zQQcY1LoIxfHKbCNCKGN5tVYmtTkykMiIrHk2KDuV1Pk3BeXdc74xwUy
akUiSfFGfkOYgCuJzT1cbgyGe5lTyzJtHKIpZeGnpL3482Kv+0WGVPY7GSD2ZXVR8Kj2z+crRyeK
kiVF2m/SjYAYx8VHP24LEvlhwVA0sZACqfF3xndGwyU2fOOLsqA1S43WjNU2gGTLZSdsdtXJnZiU
uR8eOux8WHJ38TpV7DPCHbZ/GNs51SMHbWU6C95rg+wm2ZR4v+j2S5e31WLB2S2cSnu5rlYWNkna
2WljIKG+2SfujeR3schqr3oyxfp7oSrIMelnwHDMLcyAml+G6KR0dL9Kk1xQGF6QG0NS/tC7CtnZ
s4eLqzYcuOv61AcKKG+j4GPCtOn68Ugw80i6FGFfwDRYEUZUgPl2usmHRdTR5vtsABa9XmgvdowJ
QTcKSXP8Nktgl2AUjvsqVaMyAXc1vN6W64u6HuX9lTuOOYiJJcn9fGga6HpQqqIxjLwyie93myXG
SDL6WSqC2O8BttKbU+d/4ds9ZFZMDP3QSvc6aobFKGl6WvdfiT3s3KparUfht+TW2qsFjg/GYYmn
GzveAhsI79IrDMEakTpbR0lHo8a9wUpkRo987xgQ2rFfWZwD/aEnapO5UPRkYdO+a/gKSiL8Q/a4
IGCM/JpKZlj5g2Op/pr27nveYvbh+4Q/3CXBes/uzWzWjf5bsslfg0CXKbB2o8xZWER7eTKv/gol
6J12TTLkb1kYtfjpAnEDDluNphXsnxQvDrAEOPkAIdhuKtLAAerAgXbJvukowz5N8QC+clPYe3Wh
WQc1aU3/vOMVAboRTotpZL+TCvJmLgff7NRYQsy6bdj7QM8zP5+AW1SkjOCm+YrvrotbtA75/+i2
qM1qCZXa5/NScz0Ju5lyHPPg1vCH/ToWldgMSTQU4w/+KX5NU6g706nO5RBpgtPLhrS8DEIzAlhh
7eJyytokOrWlwST2j2aoz4ATd6mjW2yAZYWk28Im78i90AzzF061FlOB2A6p6mCtZPEWtqHWDWzg
FH9Gma7F+1MIm88kLjSh1vngrjAcsCxNx/3JHIUEg7xgYRb06/XNrhEgDSukHiBsbETt1Edy8L3n
NDJUD0pdpoHsGzxPvmSeEP4ccYAJOB7ArSN1TOFH1cY2nha5olGrSj459ml/I9jDUlF+GQp1yET+
CHYr92JXUn4Pqc9dgyTZtM5GeeTv6CnyiOCX1hM91XZzdrXrX2cyKn6PIB10lPWbdKvn+PVYz3DX
VmI5YDKbjJJvQqR3AQO6pk12f3ZuTZGB1Iumez7+KjW1es4jPTqs1lr8JH/Hz6Av+AETIkpHmKdA
Td4hOMrrODnSnb1ECmztKZkZGuJMG7Mj7RQgLwJgSbomaLNI5tl1BLcwtlK1fi09YVaOqDA53jAr
MU4G+BcEUKxApfjl1Zxy//AWK/iFG15DfoA2cT41dm/xGFOt5bjv8K1SmBRhasqwZ0fFHhO6sAlb
FuAvaf/b0N5Wq/S+JRbreNQ9NQI2L7GWgwS9fP7mwbdtgBW32e6z6LkQClPgCwhjK6oBOK/mzFXL
Cp6949WdrYhdkAaYNBA6bjHoi1yMz70No6ikOeRGZKRcRgi2F2V/PvKioRzkSMtRipFI6i6F9NZR
js3j6n4epN4GKhWt4sXITTPrYNiTO2+xUp4hbJd+rG+gW/1kHFYMY7fq4RTlKWJcUX8BVgp0jkVd
5NknX2vt7CSM5DR+UKxQW8WIxnpyMtnHTQHCC/YHNvQyqOs7OyF/xPlY1BNaYv3hDYl+cr7cRqpk
LdsdFybhi+U8072vMSrscZGgqSABBRMNvJhAfsyO3UQKNJObtTkBHeFYX40x3OABMzwWvZ/42kUW
qBboMkYpxTjyYGVEAB3cbJwvRcvDyjnFWOpSzafbCtqtvsppU6qmNiEFj8okYfB48Ba5M5a+LJA5
+SBBjB8QvkH6KUT9F4UU4wjJh0y3sRQunQyhaAeOjNvBkcgSDfyhqUNE/naGYLYG/XOajLeZzUNj
1anFoKsLdrh2fehDnoKEizRxYeK4V18oYnxdctw+9vBMQ6FXvZoNZPPvOoS8h1hgjbQzdtZ5MN01
PgFaDNxIQT74Fp+esqrexL2vktZvhV272A/fIv3EKupDJQbhT1VTc72uhX3sS3zxNlFK1IT3YT5S
X6xBW3iCnGQ3RsAMPc2ApLItMNrqpRInlKsLM+cml/ywLq0KIUtn7c88vthQGN7Lrt12NOtL6mmm
4GDsdTqBZB/9nUETe6yRDjr1ZApG9lJhn/z93+jEYSqcO9SL/8ByMuWanBgntTnwMnO/MMiT6wx6
vtRUUd1uVVRf+z1yP3VT0ueBDXVMOmyPnNKnOFIEe/q631PxQd5oKnwbps1JiGZH0B0RfA1WRbDc
GwjN3X+XTCm8mzrBv/ex+AfKKOmLBCqLToHul/ZFXw2OJgGbxfk1P/Zrc90tTvzks6vglD7Fszub
F2zTMmzaCJA+944DdyKdq+XejszG78GpKRBd4SNwXELGPBkCkIdF6waNGQ3R+Si3dXSiIdnlXdIJ
yXY/Gpm9bqB9r9R4TSjvxFE6E6Z7XV/COlA6OmOHI+orrmAqz4ZBylkADXFc6JH6lUQMazCd+i9O
LOs7W+OWpt+zK/WYoBc1rkI8lCvKuM7kl//Fxwrw6nPh+EnqSBpcj6hhZWCvgzGF4KY3pbzMw+Kh
jjDY2YYSrGMH78di5cDJH6VfRpAj22wvhsJml2HnQ24P7hEVzighIkp0W44IssjhgKxBdAukgZrr
QziDQYAsBvch3PrqrE9gH2On3xvAGu75p+jHfDfozT2hg2smTI7gBndTV6I8IOgvRM7Upr+Zjf2I
Ivnt496DVm6PoSWYCQg7jm8/YpMFr6q7UlUnOPhl5TSMpKsc5+gPO+D0Qzv8T9pJDY0FTEVHOsda
G6CM9R265idnG+7VAzB0xN2fjiOYhyjuEribgWNQFwlp0qjGJgYX4Q7do+bXTkYMswZxQkbZbpxW
VNUCxJz24jwkGEyLoPj914DGFj4CnXQq1GpF3CjWeur9pcTikfStN7H50eBNYTs43s3eI6PLTqUw
lQnPRO8Tq2r/W08dRpaKdoVOHNGCLeW8W8FPDDNRCp0uJeM3Nk1yfPEZ8DqDR3wI6+kODJ68Mcaa
qChC5iyqqIDcA7tDNccKdRUMhiZ4OMxUWTVLODZaDBKsh76+ShZOk0fLLDwAdUsMTX4s+el5RKPb
lOlP9yEg3mR2bpOSBirqrPSHCaZ+42CSbvkRSVp0XRqTP0f+M2ZZrLvpcDLXPJZee4j8yXnxtUrS
MMLHIz8r1qEv0mb4sMCHOHM88/KTVyhg3Y8gqzPTsUE2ggGTNk69xuYb07pcrQP+oKcim0KWRBA0
0E6zdiNaaUt796i2tJ09kV9mPzPJV9EWhiXsnWgSS5SCjjrtdbPt+SjaSbxK0wxcqSrsklscuHX4
ZGQMP71IZFjt6MbMAdvztDuVUQcy0dwXDRzN4EwmxTlp+aIySDd9mhxgcxlJDpKWE3Dc9BIazjZl
4l+kQH6scLViVWO/kKLMkixik0tALrBokiSmhjIIcPxzWsEOGs20MnusNU19D7J1UsqKanrRSnB2
7nACg3IZoWFtceIiJFESG5KAleclJuQAF8IMNWfwnqqbEUke0H7cHFVBYT014Dm6NYF31p4ZmPeo
f9hXkCL2pOtNUUT6iV7eSmyKcU9gr0RYRLv/5l2NyCa61XlQlhAiZ72J0DC8zsCiiQkacRa2CF55
KDgPdbclBvq8POkPwkW1+e5RTFG3c2dvZ8gmn/j3welWKtQbpFMQiQZxI/Vg1LkMhiobdBfOwaLA
fXBuS3NOz+xes284XJ8Uf0F8pfAzq6VpTFa7ENfdwybtCeep6RrZ88r/0eG4cPT0fcthvAiRho0X
lQwuSClE2W8hk2CXpj2ru4NTAmgJsCdQhIjwoSjIlIaKRxa/yOKzpgjS8F0tdtNGf+vLwj1oHeY4
thS85jlBZDz+A044xhV51fWHoMVUaWhNLZR26aqOJmb6Edco5II1xyrAe0V1aWxFHwSKv/9N4A86
Fq/E+YflrLcZw1rc+Xx6TTRT2Hf2DSt0lGvVaGrpGjzEltYjW8imbJpjpsbRmwJQhXc2deCdoNMP
F7Qbkb3mdhBwH1JvCcI0dT4f0KGjt9KLC6eAj3wd2wduCg/EGrGbOPXN1oSjLiNw9y0vyjxNoVB/
S5B2slNBGY9TfCwiBFZOPwANOpJEl6YRvWcEMM5P8c4DdNgyDM/BY34UAauy0AuD0dRh44mx72QZ
5GrYHExE+a/nQ683JZBUIONXRLgtbg6ssBys5b57K10t5TQg2eG435bf1+4x1gp4g++8Nd03i0Lf
zf6tphZ0ieT6MqNrHi+77/aK1ZeL56rzbg373Rn3tovFrBYduSmqPhltxKKEj7fN6jU5/aUBe4lZ
UzHOpd2Ei0JYaykt1Zo6Atj9Q8APAskLSG6FyIDxn9ja4euPRMb1I7CxT5OEopO01L3vRaIbb/8J
D8c2GHWcdF+ZomcgIe2k9NWyPpreGj0iRyY3ae3SiyGq0Sab9Y9/pyB4QJV4iwZjAgDmDlJB12Oy
vua8Trc7lyXk3+qnmOEgNQ31RFODsQNwwa4HEbtjAi3C5KYQDDXIB+T6X0e+RdX8g2gu97nAt3hZ
YoqqJZoxWQLYGZkyeVfjHBMUBJ+xbFG0v+FT04M1Tq8/3+M9in86/fyf4SUprRHzvxaRhSbDOmv8
U8oLeR4jeKbavNTI9cTaCYunj6UacS+RNwLR7IcdxDxD3sJitruxqhyU3LDwHK3yCfYz9jaLXoBF
hgfJo6tdU+ddCj3pjb4pUj6kdBeSf1oE+k7qldA6KDrF172vdpAzetXtnkMO5G2jlSY/kubH99lq
gqIHTApC9NeRAJLUIxcFXw+IPAbP8/QAxmWya8vgF3xMI58pKHNVz/Oiu72qWkWMdDUEwY3GjvZ+
0mRJpCh/TcJWuGgVSki8Ctyb92vuvmIL4vHbuFNCBgw1mqCGF8xwCjsDN7fTG/5RSTY0MUaHsk2g
/t/5G6qnCoJF8mnHARMEwxRC9aCDm3WCae0qgrLEH7rn7EUBEA38eQ0WrTNhtfihz9s8I2zGQmm9
R2qM8yZDZrdmfwJu8Ep17SmBOQ+foQTSNGYtot6/VV8utOsD+hw4fiyeH6pjpsKyZa+b3kaDX4uV
t49GqrJeM9BJyB0bkH4SHSJk/hAIW/PQyRVXuYpeZ5KhHJYRKV8Lp8tJgUzWXIbV8P+65CKClUql
/o7qc2G6x/LtMqcjrHtjhRmPkdhUVaFSQJFuFizkkSwR0T7ainhSMgFuzTG3uWJCiQDERjMhTIFB
Kdosmh/IEHiROcqQIvopXwfBBmA/FxA8A2d5tRkhCsEEnZBl+g5q+uKHvlErgglmqBnpFPddNYQ+
wz0lnchYaS7QG8dIq2H1Aspwp2jynAtT46MaahhDRfwdQO1y6TlWZse32cZ9bd7u6/yylTQNhIPk
x3Bz6zT85HuqMTstJzK2e8ayMKFYiOPuAPAH36E9g4hnQvzD+rGDqbVKMfn/iweM/JLw9HJpR8Iu
zRnlfG/48MLegkcJAcJagkRdOBBnHH03ptyu/UrsUP5zfpWd0nqgtq4nOmnx/+dXe8SkBbqIasKR
ZPIt47c9g+zF9L06VP65Y4fUqZB0wjfkiLh5psoT1Q0JpdSaAAfDNmNibYQeuvvT+46PMsp47rh4
PeXKjzHO4syIvZtdjzV+HBrbyAKOVS4xTNgGN9GjXHPITT7JQwE5JbBsl2h7U42h0cKMBkGWbO6X
EVCxsCg2EsZ8qGe0azVtBf3/iKosfKhpgR7nHAHLhaAxAknPmhj/TEub2FyXeyKoR3RPxSUdlXNl
kVIE1qLomgcO054Ka/tC5QlK5NSE6M/n9/MLN9p6bHdQw0XMm7aA8kJx5O7+eOTMSLnPi6eFd6Ek
hpii3nE7ve6X8NiF+S+Kw8SKXr/aXMDxJ/V5o3NWKkZQFHwztmH9n78V7maRW8K9CgzzqeTbT0hi
lu7RIr15c7gZ/dHMenV9P1t8Rhvyv2nGWFXbgMVhFa7UcN+EoPB8kHE3H98E07Ht6gnSnkpjtDO4
N5n/GAZErgLTufkUYIIweYGJiFvjqF7ozC0841QtrJ013hL7XKGlpRCv7f1HpGYCuFrgjo1Tqv4I
r0vbYFvT0byCZaQLlUP/iBQKSOQSqqLEZz7DfxgfXhmebMKiz42X4I19nJF/TJm86zuCdLm03iw0
psKQ3zxp3AgHRENDkbX0ExNdRg7R3qXeDL343m1kbn28ArDO1JvTeKi4rUEa+s3GqzAHgHs5J9td
scTdjvU9BaMNG0P1yCOrpiXGQLVnbSsOSEFyt50z/jKajMCigpXEmJgjV1g1ELltUsHSf/6jsJN8
0tdQR5+a3lc6nud6z6CLI1vYPo+/7hxJ/cnjwvQs89PQmx7/IsLr57jnmhR74rqHQbvyVKKsQ+ku
x6CgC4u78u/VSMbuCiKG2bpyPHc+O12gIpAePvkGib3ByoMiQmCDLTRGptf7X7oko/rL064/Afwu
gzxEmNNBhrYzmer+DRO4/St5PVFm6BvRjzh7S4EaRG9hYz1LvYLTYsYKwyO3eqL4hQ9B/GlUQgsE
4kN4WFerkbNQdFLldsJ86kOaQdRGZjydREzJ9Qttuv6ipCCx6cUbCt5QCQan+I6J89gfnfVG2aUf
WES+8zPFNY3fPJmpoCXt1za6TyIs24f1TuUSSw2qePD4HugdNTIwUQq5y8zB2qPKDSvH+P1Ha6LE
+MFs1BO09f409TkZiy3Yph5NLou5Q6MjGFLNDXvUAb+5dUu3b+qxBFSeIb0H3GRjnobRbKII5PlZ
PXr9AdB50CRqzN6Xye5k5pqh7SVbOKEaQK46fnxak0Zv3yRvoqtxxprHcpXhJ/N7SX8IWwVy2IJ6
Q9tBRlcszHBYbA163yO/8/N1hzs+0ICJXNKa92gkmShbRd7JSXgKt6pzV5b3U5D14zS22npvFgH4
2875dL0eUwHHUl/+3QE2lOWyZRonQm44jCK9FBFf4hRgeQt3WygfDvSzYnDmxE02SJqvQzopnqAX
5BMpNR+hF6cfkLMC/rV2tN8gd/SfW1G80pEmeWn6aUUBK8R4FrmfCBxO0u6xMuP7ryR3rTBSBFyT
UB/4OSL1yk8k6jw8qeWxw19llF1lAVYy7utNsAggcTcjqqZE7mwd9Ub6mpFK9T9KUvYOZMasau2P
cNrysRv7+JQtyMh7cEmr9IW/3yA+4kR37Jwaa5kvhxERkn56Xjsvl4pWm2odmUH8u2kkpHL3EV2T
UpNNXLLoXKtagXYa5sUFwwsa8vRAzWElFQ9hQGuur0pwgYm7dVmgi3DUIk2OQSYMAN91DEAIbPfJ
+K/XhvXW61LqmxfG7yn05QtMU+VLuwbP/GiMfv82waPzH9NG7vSXcWNST0CNx2fKb0NKws5nHSkZ
W/hZO12IllDkRG41Bcib31l1v4JUrI+qT/Cunc5Gl7QMJA9vDxFEv/fIxHBkiA4qIpWBPQBh6fgF
b85mH3AjpkfN9KeGYrsOe1euTN7L4QFGJthHn2LsGWq7PkXwU2Xz+Rda52LWngtjYRkZCz8pDEhi
Y0MrReCFPJ1udNuWljbjnwJ3pJbFn+Fo400Vxdhe/CoPXQ0KbABN1JAwusYtoQMMJTuVh+6W/ubg
py7XUgj5c+yITXwEo1xaaG8/KxEIKSmrPe+NZt9SCVChUYxqPULpQYdbCtzqXEm6I/tkpNrQS4N4
uRJG13EAD9n9w7Hm5G929x0Z6jWlG60bgYJ7f/Dxiuw/IeW/nUsrAn3BwUVyYzl51qaWP59MEg9X
sy2HJbY1cMqaFTbTmuKd1Jv8uBnHAZYqRQukplKXrqlQaVOfXTJQ3Lj35xUZlMm9Sw0qyIY0wOSc
2X18UK9rFbyV2rDfw72j7Yc+EE8hcT5byCxtYdPjpCdoDdr987kWlvNXW+Httqogt8mrVfkMiGmG
sMgvQ14cV0d4NkuVrj5PLj4eX1aaEt9klR4AaNOMty71RzBGWE+VQ6MlQ8ni9VfJqJKSEcJ66MYL
syCu+OiO/WHqOwF58HtiTEEL2U31gR+FGYCMapwiNqwG3yOtgk1Znc2EomCa3Z1lUM9vOPCZ2ayO
ZGjiEMxf44IHvDhMQ6Pwhm89g0y2k9jq+c372QpMBq0euJ7GruE7Qow+ck22xhfuOlBOuyo6kkFR
pq7Dz0yWA1HDI24+gakncRPCfdy+scWowVCcEfLeujQkFPknfFZIQSRIG9Uk2Bbe7osxo8z56Wbb
YV7U7Z6PzNUmj1jPMwHGWWfl/9iAvphTrytnC0bqij14bHqUUmqjvAkw8Go0OW00tEuTUN1yQqat
N2zyLqJY+pNdEVbw980pmzoRz4XcqOHTjtBVwMYWYKq+dNVv+FSWvbYJT41HhWDSEn0/b6iunHBH
lLNK0hr27nK9OqaZjrLNAy50Hfj1H/dLHqfW/tT2Aq1WzjDm5uCywWqS4DnVwrd1bBdJFdkqZCS5
GRFiCAS1Kn+mtfkq9OUwXseufT4PbK+cEMawiIOMFYwe9WxHNHXgsaYg7twor7pNB7gbeVVlfE8m
wPZRlpRDuByTn7b5+4u+gi/pA9S1WNfovQO5y61JsNOUwZ8yKpkvC3PLA+MAx/b82oXjjjo3ckyS
UQ2E6KkM4WiN97eOiEiFwHcNp2sy48wC5gF8NMRWjwnpn1ft/PgpVTWb3Hep6bbvWedgOT8r8U0x
p+YUHPKncNPBEJ9TwKLts8AwCdbysrY7cY9jZtS6rLR6wnpkArI02zzviM6FRIyB1QuZyAOQWIPd
qPjW9I95Hmsr4h+KVnrMEEmkiWGr8tV4iDkhy8ElJySfNKeaJYPgoHFVF4C7ZFBu3mr73sY1w0ZB
YVwT4B2/hrir4UVL1m70ocJKTerlWdrRL7Q9nDD9vkuQKf5B1Th2UqaHijnKNWUXwxkgwRyjaK31
09MEvVeVyWx33rahBvudJqDWEaZvNhy57qx8nZvaIc7U503oBae7ezQVkhO1CDNehNZ2oBcNc3iX
qlYz+YReWLvmgWR401eLbuonefPSO3oL9l7GDPkijvMm58NZvT7YhVNkkCkIUhRhe8/QKP9yLXce
6F0VYGPd9OdKnEgGqPAc8Orwc3HXoisBlEYkrTN6nxiLSdFCI+UGixejVZ7CBCBI8gHQHjn6l0JY
T8i26vk0HOzPkLdDEIFkWYU2rLH3xF9Wt1iEDctMgQRzV6HasOtLDpNvps4Yfp8rw4C3Ckb/OD+o
1y9soexJYLucedKqvaN9W2rLHf+hsbjkPrmweSrC7UNKa/kO/tmu9SJ369X80Ldikz0Y7sFgtK0B
oV/eRwU55h+lxNweYBd21isvXgQFUrU/JqJ79QkMD2lGuZ2oIx0Dy3rFMXao/1kwLoJP05mibEQL
k6Kt7WtaAggM+fcXFX0W9XKGR5cQWhqWulJSG0zx4aqiLX9PMc4wNFBIevSi9VZTCd8pHoSXRDOJ
EiF9l4xkL7ikefaAlBMZqm32gf8lI7DFHLI9OH2KmUM1SQfezfUTgUjYQXZUBSnjO2gcnLqLftSt
yEUEHIKI8x6VAiBHFHZWP8+JAy6HCMbH1zHBdtIjyqEx0MhjWSXzrKhM4+ckDlglfPrHDuAGeQw2
tT9Z41hE/SnY++eqf0Fu8m2LPhrzROD+DFuz7NWfavbcNKDA0F6kBjPW1kUmZzcAwuS6ErJTR/rL
DhklqQJLZ6bZ7rbHxcpuLTWEDx4+u8fuw6dROFjk0bg43mp0zSlg88AZb1R5VgeIJocEN3AvZPCv
Mn5iTy6Oq74gskMMROvYieK8OYl4cuq7xMMo0D9XUcirJdvhdJGYMJUXUulEY8V+U80fCYnfE81h
yrmrR5l88+fHdeEgqkcJi3a6MhRsMokNHDENAK97ZSNlF/Iye3L3L94cVuA4g4BFgacd7JVZmTp1
dwwPDWsQODDnGpMyiU+nu4PCSV0fCa5+89UV4t3g6gBzbqvQl2qdSoxlf9Z4L5z5OaaxFFSLvwO6
XDjohhnRQtdlXxZ2fLBGviieC7sBzLLiFRJ6UyGRumYBErjsh17HP8cl82G302jYubb9V3CFvpfV
o9LZwlS/nHsJ9w1JROVSDxnFGStwWq0sFdqrgA6ZE1vR/ckVyGZzANACdf4HIcIG272MWeDzqNJE
Q58457tAL2JEGJkX2Jxs+HJUZQSxiJo5C8dFENGOkZ1ymoxY9TO7hDhrlVD2A1lmhp6JVPlxFRua
FiHXZa4V0QmWxXjedBf5yj/E6ON5SjbbMAUpnYWnQQIAr7Zn1nHYHcyQdgRWQu3WamiuQMe+dUEH
JpDYMFNPZEYzYIf77beEl4yK2S/tJou9wFN2NmjgsH0BJ8r4LUSHnwWnOu+1TwLN0JhyxUSzpzgL
S3GHu9a0o1zDoj6quuOsp9bKW28OCz2H972eBPiTOENKsPNVwolo3ZQ7lktitSSMuYVHMUJshkbG
OGctlJUvTwqY4ZhrgKbSAP+cOIwMJXSYXpjQIpl3bqhJFE1ed4JnccKIjtbr54fFGS+Efv8d6VUG
tURelZKWsEyRFa4YSgWSAQVQE592CsVK0B6owfaHgI1R1m8+psRLDbgbiJgswrYF2YGUWzaZUiil
NxfsDWyrssKs8WvHZvwZe5d5b8g+aZgH+GPvPIwyC5nlmY2vL5YYo+MsWPRbaqBQPXxQdMu+ZfWX
ZofSVVmWXwHC//GQBjouIGbn+VzmppBwjhBfv1Y0rz6chF6i77Iams4U6CwIHmpzGsm0mv9SZkZQ
FRVNeBiTa8d90OdgSdqYZVef6wErbeQzve5b7uipilVuuLhmjZ2fGDHtvT7n7Dk4KdWwSL7rK5Cb
SNv5RyofhkCnuDTwiILirNPFXwpJs5jC7PyFUylTZb6N9UbFui23jrpmbgwIqcJQIDmMF4QP+iMZ
SE5oOOl8qsvvBmPEemM+gcJkJJfxzD0oe1WbQAGBDMJv5x+IP07mdhKvA0uwUAtiyzoB3+I+lTKu
z9YKf7LVo0UGqR5s4V+OpsYa/meE9SrKGZ5RHat0n/bYr85O1jpYKESku2WgnIqc7q8WCzbz5vpp
LUnAGVBGw1LH6bpvg5NrU7TPGtjetdEO7roVGQg21fpDUo1xk/4+DZvZCRPH5aUOE2GUJHn6x+jv
uNdzds/QF5YEBb2mVDs4KPMn2baStOe4G2L8o5s3W5sOOeauzw6kfdQeRFK6BY6YxzChu5xze6S2
sKOqEGliu2uBefUF1Hg9Hjzlg0SXv7u+jLQNIFtdISRR9v8Bijl/KobDYSQT6DJqCJQ1X2FiVZx0
ogG73fWIa4UDB5ZYTlp8u97og8lo9Ymbw1MJt2kJttz4d+Stim2RGql27B1YAMcqLxGDI14UHnbe
/K/udoVgWnDP7a+J29vWqAd1fWbWL8sYuzrmIEY5KKazy+kBNlc1OSkp+G2nNVK6a39xVWvwZ3+O
Og80EoeXIarDY3vfTJVV+Zap/9dyfv6wEFPpCPIZv8nPspwUuvd4Wr8DG2jieqb/0GelE4a76DYP
em2NnF6LNJYjSNlhS++XFO5r+iaE1EK92yvZOnH4BoLxXsaTkC5Tc3/JY7LeRPJuYCmr82wiNzHA
oRckxCabTdHlW85Mh3eqpYqU1mRa0O+Vm7VKykDOVpbqlWiirSrhbzrav0q/sdhFHGw3qiBUxiMm
s8j1j5YOvy5JUsI21/Ayz99lhthmgD7e5KvMC8G24QfmZN9aWMLaZ/MO33fVpvQ+fNDdsYEUvpYc
yz93C8Puh+EGDGB1+08dCobkextER0dMtRUrjHaGRx1KuL2epDTbK12SXihhYcLtBsHCLB/FQsSg
lWVB013pOxS1j73bIF7+l27CGVeozQMWUbWKVHqbcDgrdsCEermShHZ6E0jlfmiyCRKoW1GODDmt
kiO1SKErVoFoSLHinjih+wrq1Txo8Ke0R7iX23G+LJr3cbfwAwbHpMfvnJ0s/rhj3SWbNTFVGakJ
BHSXPRx0jhqBxRiFptz/NzwNLNSmQMBRSep0e0Zpr559ZonJ7CkrL7tZepNKXZUwAzucqSOFAqIm
GPisxKfQmd4wWv0dDmo4kJ0N2L7IwJrRslyCLcEhtEiVNEW5MfDbPXJD6pkQ9Npv6v5cHLazVY7M
vURKhGlU4qrH1SiXK9FUJ1o9tcqwDiBUuh5vtm9kZg76O1fkcmGJ3uy6KnL2j0FTx7lF8az/n9PY
1c68R9ZhL5nsfsE6EYisN5SjaHu8hDllY212dkCclvzzH9oq8Swe1iUKCbxsmHs37HY+wnVcv1W6
Wwu2OTYnxUZIKMi1GeIpNs9+N/8lSu/6+CNB+xNLv2SmrZRIL1skbmTk+wbBlIh4LVAqGh1/Mu7W
LqujtxjrFEsYFVa1oU/Y33h6NHbE/tsXepKNSjeuEmy/bJhq5WnKgZ7cTjwiLS9UKb6sM6RmCQrM
GG9tnwlnYoq2g6Kb2GWA180ITMHQv7t3JmKOC6au+hF+JOciLUOUlmapZIILXx2Oas2fhTGKYySB
ZnlnAS66NStGxIh8J7UjbmR7A4/CyfuoL3SwzHrnxjKC1bLgfGHG3jUkaMXmLJb8oMNor9l1u5mg
nkm4RtX4AfHOIVqrZlbiXVvRFYqMMfyhsb/fI0u2XF4HjQpAQtO51eM8eaMjWSwz/0+qsUvJ65EB
s82HvuVS2gg2gWV5+iC3J/yqQQ8wwnhhwuNwFuWRvnolNaWWGIBDG4FeJJ3JbgHuZHqDx1vKqdLi
M/bz+KuWd8UI0Br47x2PsK77twGDs8TZM2IEaIJVNbfoenYU75fzAyspzVbeA5zvqxXpH48vAJdI
NDg+n8i1+oluGo0LhGxq9cU1jmkf8iVynCe1ZFqR5V9RaWyDvKROXp+w1BCp5Zg7a8r79Qxh348e
a0533oq1vYiGgIY8y9nm0/jFa6g+Zp7KyybUbDON5KRf70RWcr0hiCKPX1JkF0gUvJG+hKMz9rLv
WW6XvxCTSDwk3ULo6+wQqUR1QjNcG/VCimmNJuLnTEsJHyzxRtZAjKaT6dTcguuvTkxPDrEKewWH
XtjxDdGNfPVWB9C1v7gq7zB2BG5jYV6pjz7XjRLKqy3zLrgi1nl7XK/Jbm2iaXaWazpzXENIqyC9
FrPip/jojky/q1qMRbvQ8Ds0yfC824TXg76+gXDfNzJ65DJWrpVkdgq8zZpqKkfbPE/HlHEqJAnJ
m1ftOF9T/ccOfkUcuLwxUf8sU9t1vbuWXBDic54Lvr/KKoVxno1n15Cy8pkM/WJNVCMkGkMi7Qsz
T4XRNWAYz5dM+dl9ZsrsvSnomr1+pFUHZWyGp40BVw3XZ083B3fVG3SBsNvPepV51Yj2AzHhQUEx
dDQvCZ271v9hESyau6gpDddAlgyrJHC3vERnMcEvG20SaWJH36iYVUxq/EyFp+PoaZ91GWFmPuBh
bAPaCuUynn5gS/714My896JoEq7MFL33f81cszQkJ7qfhWdzL5p2YI4nT3i4ffoVVckkPI0sXe2o
G7sNwsJNzl5J0ZlMaQn+nPf4DTXlfGYXIKc9bTOQ6grCpXeDLc2pIF1G78lmH9fMOnGRFngKC9kw
5QmbDaI1qm16DK71iLdYcrbKHJzFa1YXfgVQffs6CabgWT4G/0fr11uhAmalqSRWB3rv3UkqsNKV
mzQIlrVeL6kfgbejZF8wZb7ICLuq2gy1AaBLjCeyqLuRg8x1wr1kscLYEusuS0NtfYvXXc/9dlKD
lrRcJn+FV755Llg/oIT7HblPsi577SNnlgBfFpV2uscm/Can2zmODifgneFs2rzqeb6UEUxMDE5X
bmPxRpEMzjV7aMUOMBx9qFxQVGhsoV5IKNB08yQjJa8MD/+1hxOJoO0r3JSkWFLY/Y4KvCCLJQN7
dq/R1pKbLta5rOMsZMYB6rSOB3KKgtpoP9AS6nofRvrVeQfEE4fOMzdTSVcAqd1jGn7S47FVWZwh
JPt9Skre8yAklMdM3kfuo9bb37nXkt/BPuTDYwp/68bJAxhzklvdzQbvp/sv43xuwUSXQVOFS7jH
nJwQoQguBMRE/BDZuDTiThZCsKfJkdRAG7HylyTiQFf3Ul/7/goYrX3b+bGGNjY/BlutEURaAjpU
W6k2MzJOq9x1vnYj/9dJSAfWDzmfwDCBLTpV/GcE/D+BdmDAZJPCpCh4eLAK87wNB4PfHKi0TEHN
uhy0WEOKz4kZJz2gs5t69jEXKy9PFvEwFL3yTtOrX5vh9YMg4vrsM/gnrI1Ua2KiXBc4bBuH0FEI
vG4ExQ/QSorPy/K2SCUQ/FHXYIeDRbFxpxOTrUkOGabZ0cOPpn9AYNf6YbedNDJMDzlEd14QnYai
h5V2Fytz5I+RfbTziCH9k/a8RpJcdKV8Gt4s16YIofhJJlHPpcgGk2p71IAeGLYMO6cz/yl6SIjr
XUhqiUh0pc9GarkxRsX7kSVRPTP4ZNp6bG53HOxs7dIQaScO3REewggU6TVE+LE6MQlc+PD02ZDb
/P9zrvySXOztkbwIyhBP/ygI96s7wyA/OZlDbkWnhpXA4sXaeZyej3yOuDByXvQs9O/ORt9a5sV8
dKbl1yKB20rpaFx4ZH1NMW9vQmKVbXIl79mtG1hBPQunqsWeFdPDNN2vpJOPPgruYKPZMD3Hrlo9
lwWPT7qMIRt1SdqSFOIf38tbHa4cTK1uy6thraEzWj/8tPGLYm+ZB1waMVlLv9kfHTY7WhaKcL/s
wLw/SOzjxFghzLbw1NGpTfbfdrZ39P7cxmSZlcXD79rLgXD7M+SKnlW8Gop0LAwCgyFuTKJc+aLI
HtYxq92PLir/Bg433sSk5bWnMtE91Zp7+tFtC8eaF68/Jt3j1sc/LkvJ9sAWmbbqkt8qNcz57GwM
qzGfINfv1270k3be+AbNwh+sQltcnwObsftCPA9/xHa0b2xorRf8bVuvpmVzzCPiJ17TCTuvn6hr
t5LFhtJzsNOjhKzGKMrMsdpl0wsZEqsCAGsRjCjuHrxLDDfyeHc9PT3oW3QXFUtSWubYCEIFeF0h
3S0FHT1Rp8woh10tHVSGUvKh4uMuXDK9C7HryT74MszjiPt4C1a6X9gfQzqQ3c7PGRLj2AFBox5N
fyaec2zzqC3djop47T2EkyxKT7OvNd0fXN8YNDlWsPjNCoOKyR/6SikOzWApmVOUlYxsleN9Znuv
9fdPUHyh8GkiTYuBueZF7b7Cv5BMNar1ssM9HWEdLvZUIrvHZzi5C4rttnCK6BzjW/m7+tpoVYhT
lGs1FOzHmlvswurGh35gBiw5R+iRrnUDFOQMzOzXaO+zBTr5sTWd/fXtVnv7WyFCdHcENYJQKMjB
Jp3J0PV/mg6DlXYBl7HZBSS1aSVxFljMrGSFSkz/uBvBoWe78OlzkwJU3ZZ8tuEDLsUQ6RC5xpkq
Pfc43RF4RL30IpJDUbq7Vzaw4MmyifWJllXnKGJnbJzRdrrJ9wGPJiHUsMBm6ZU5HySXbwcIs26Z
0iv1QZmn9R+EexkbGnbN0jcdnGLQ74C4qgBNwdEXRx0mXum/GWVB2wF8Gj/n6V0lmkmG1mK/IYXC
EJpUaMREaP8FDRXgWS0cMiJYLPaM31cxsZydaO/tygBEVPpbs6sWK/WoWUg91JOrAsYgqtrFSzsK
4noF3UQ6b8JR+xA/KI1M4Ye9CGkH1WiUR5JyWyoIO0cBLyfR04+VSmZHRROEs6/UMS58XTgnh5qs
Y9yqXtCYEoetWbOwUtHzpmnufUBVhafEL+UYTWV+IzOTvYcK1ct6gNSoAUNjX+Z2NNsGCdSHfzaN
wn94yDt4RBdxTeN73fZpZvC0E/skM4/k5S+GuwOWvH4I2bcBvsXHKbkl7D8EQsoiLmFXk5MfwjAk
BC+Gdcyi4h7UYD6NJ7H2jlxMgBO81dus7ra157jqqgiRSiSmLBy5jK1Xo/gdbZmVakeLH7rBN6d3
8ULR70kPapNiYn7hca0aE1xjjGfRk15aHuB8gPRG0F36D+WTuORwtS0ukfEmeoH5z27ehChqZZCH
TNn4BbMi0OYDxL0SsdDAVmJ9ET/Mz88Vha0sim1YzIXCo6WZ1xdDXQtVzAl6J0YrRXXzZwPDSnpf
APjw/brTFu/sLbR737/oHYtrmdn3EqeRha7kcRHv7fVIX6n4Jct7kqhGY3yckeRWYgg5UAhtsGAF
d9as551Pnqk51hhDllrvWuFceGxRYrZwahcMDAoiATU8yd6XgUVEra4CRMyQL9cOEkt9wtN/yipF
7Zy7qMKbWTVtGp66w++RBgwPLG2bA7W+8tKWyn0c6kbbdCyEGNNoExeA28oklU/2XVaW+0InlIqq
3lI3MvXfEszJ1SIx1gExRYXGG1PEUOZC3YcgRtvdifay+H/VjGPtqiYpq+fuZaiHsmpkkGBcZCsl
ryVdEprqHVvelMan38JYdIXZA6Zott+V+5fOusoucbuOqg3PZJVnbv1zUhcyNuskE5YhOuzG1IOa
NtbFl0idQPn5qZmbmnFmpATa46FhKXC8S/zEvmQbgvami2Ur+qreQd1vv1D9vMAteevR/pEtCGy3
tE7nEMAmiDTVJKEW4iiwjX8EmtZ3x7NaadhVjNja9c7EItuwvxSLlcoGfrjFhS/Cw/JjAJRxRS/7
LEMs9iHBr8GFDAOIqgX55WAu7OyVeoOUA86Muprp5dVy/yChHu5bGr/1vqHiInZWwBWqs9A146SP
qzf5Jsjdfr6NuR1lTbpjVturKsMzdpGdmsaQ2HDMU3MSPugqCqbyefWCpurdDqw0BHeke2G1GQ7d
mD7lw2/FPMovTJksjHPkBos7snBJmsFCBw5p58cDJ3RZl/RbT6ahKC1pONe5/GvphqHrsmDCNXdD
GvIIQ1VF1dp3vMdc9BQ73fOXfPoCgW9c6zzop39LRa35KhOs/TdA9U3LdSKd31svAUQJtor7ytxK
fbASJRT8d71u6+bbmgguzsQyg29Lwjy3jEJdUAqbjcdR9PPSqQa0Y2o4SxzpWL5IgTAbB5T/0y80
Rtr80hfyhqP7wbrnNp58mdVKD7owXeGAcewH3D0iIgIWRloyyVOnUE31/bfBH0mU+bWexyXPI1/n
8O4wYBWEw2GYJ/42HcQSp0gnb18MOlbRVtitrN4C/w6q1KxP/Krex7x7SG2UeIZk4CBx0oiZnD1R
yHknnJf0W7Ns04BN1XLSVKh0E/jmfPQxemWh5maV4sgtJs05lVR2cC0XFp7u9c9OqVHg8RhDywqq
UXse5ccMzdpI5iw18AhCnfY7jUDzNurJO6J0UI9a/hTAIosZmaUwdDjOa+z6pQpU4CuiBQbBo3ng
NmNpzGR6kDNdXX3+nuiGGAmhC4yiAOtv6yuXcnMn+yrlTSwXqXxvw8Ar3kUghnyAtKCgFaaptDL4
IObjehvJVbmgjyoEmEOO+kzQ0F4VGD0YOkT16H4uOsbRzfRfvSGBP4AFINhY7Ww4vkXu1rVAnM9x
dPk7RTk+C9N6rlPIGsCsqvkSfTTDMKnAvdbtbs+/0lmw4Xn2nuWppQ65zf6jBzDE6NJcW/6v+gZZ
IZXlFjntzpVEr6e4K1E+2ykFkJpjhrzI4K/wJ8YP12GCfo9SXhfsiNkPAOW1gL5wIWdAM9kmBokw
K83+jOji2QVYMmGx6F3g13nNG1joLDYzXUohC9sJHCOgnP1veuz13OmEVBHcKi/dSnjNGVQcaTRE
7omvm82+UefrAEpdt+tLC6j+S1BDoYQ9vwpwLGiFkrdCimt4tu+KllUTeHkCHziC6M+0J4Tjk3rQ
Dz/3xLg0TY6A15RO+zpzl7D8Vmv8A/Ri8b0zJWWjmlCBankau1lULsPIJWj74AqUNDy3RUdrIAZ+
5hQr2EKVkZgiJOxbohrwpaZBFRm2eavRAEdFrhKNxGjlsc0fsXtRtlDpqtYkW4agFJVIlCBOnlwY
GixoBDt/YNOIGoZM+B8e6g/BO3khoG0MJcHnlOPwVrCyGQ7EeU340wOYWCosr5BtuJh65q7exhcY
/yBwUWV7KUi7HumCAyqO8Sc/MsA+yTTYq8Lv0oH5YddPeAmGXh913GQjCAF0MuiZe31TwBouAD2l
YmELU2TQAmwqwWBU+bp7mzdoFvzfNxR4QPR5LFkKUoZDrViJrzHv/jj9wNw7Ks5S9ydpZtdkyytQ
LJwZ9rY9KoKyjkgWPnoT/EoYoKRc8yfMpMWmGd03FFEWyv2+0QqFHDVRbo9KSFBMQ6L/moD1VUj8
Df2+8lK9qZP/Sb4oOL7jwIHdFwKdbTHgDqty5yDlX90zrN1WuZN1vHV6nV9Fq8drQOTJiG7iGtMy
WBlxNMQ43UPwu0HeeEUxjj3mHBvePRKEMRN5R3jr/6l/4VJ1U9CK9GH+bo1Dt/0EJD6DS0EzzQ4w
yZfP8zDQUV533u4Y69YH/ldYMoAulKiiRywMnVtmNZfjSW6Rz+NRGLcvOhrjmiDv6Ni7NXiv3K9h
JhosBhYcy78/1YwHX3tnqBya1qn4PduzL6sAN1TgIZwmkABZljpDo0GEv88Qv3gDX6PawjR4IAkR
Mv9GEYlVwypzLjBR0DdLfd70fCJV+b6t8s0aYX49/AlqwnH62RR3CfZ7CtL3KTFB1Gi+SLerFUAq
K3XNt9HLMmwactsiblFgYrVI1N1efy4/iAyC9ZrpwIYMU9C4d4xi7fyshTUaWf9N5OIimGTxpidT
GzId6FBs8ZsKP7UqP27/vl348XCHxlu0TszZLyThe+e3PGUM9BiBKfAH4KNGe/H8KaKbWmcs+Iiw
zPQyOlgiLSmfttJ1Wawf/suGPI4Lslp4WLAVwcy3Jk2j3miFe6FBnrxaEWWk6hg5ljqOYl4IQONM
L0QuoPxkf1hmA3OJltU2CC+l+mu4jyqRNiRnqN1DiyWrzy8cBuBr0xOxEuOtIoOobjjKVUmx0qn+
/9lOg817FsPVY0GN30lolE5uCNFfwNGAlWooBtiowvdTkdwuS+qHxprPjm3Tfw5e7sFIJLRKyaJu
j1Y7iwGyEvVZXASvnqeILWc57jWGCnFgVcmpAJ+X2xpdeF2DDnizk5U/W49dzL1G1H+r3sEivHgZ
vY2GIKVIbBNPwCWA+oQ4t7nGPT7EZGGXMuZho8fn8mOgCzKV2+VRN5workYyfI84qsHIWq04a467
hknc0MGFoSaElWEDO66G1bO4KGyriVV/MFzGDbaHj6LD58AgUpbUEDN9Qn++9WjSMIlZI1N0nQ1N
uK59ZSYcMxU7HruxLYY714kCRPMJNV0V2SxWegrQ0UL+767Hb8d3dzO+vZuRhUcpPpTFbK+Ws4EQ
uXzjlDtnbT8D5SeM4C2c3mVuJaCY3yOS7mOGRTT/VwT86/BhJ1uyKn65KTruU3IcuDDuK0+RCiUx
b+tFIpaBvHlndAEpIjASgR+Flic/RjXwzRCNsJp5kNunV6b8nIfv6zCpC4OrDUWZ0fLfQgRjBqJN
dP0eZrFUWyv9iZBFmGjrUwUT6UOXrYjkQ6HR1Mc9jZqEEH18Ce5kcAOXFdz9hcsdyK2j4BDEq8O0
tXbv80EAqLETk6Y+z2LbhIMMU/ZFjShgUp4DSCcs+5wG63qXtP1dHFGDqDFo6SeX6IOCNnzdGPmU
bJvpA/bl0dpD/6sx2AIAJAh7+7Q+kPeUYdONUg4P9YakdML5FT0UbOTwAAyHE+p6Jv32aPwZRao5
KmCeFxdUQXoD7jggdr4vwJAv0Pbqt23jWdCStOxH3m0N4r5XP7tKzGAQ3GYS0ABSKU1Rz9jG8B5b
XfAStLPU0v8U1t64TNSc5zZu11FHpEg/3flK8ERTa4H08TIfLifqb12WZwqej93VpVud5ADbcbKY
6TwUfaxgEa/Ps64c6zE0pfUArDgWq85WxoiBZvblYwk/lNEINrb2vES80jPRFY1P8i2Op0L/L3Cb
rXsIxT+OD0Y05YynU9mUY0TlQeGHs/dmVPCJ0XaHETl2SogDVs5vdnOE6xMAfxLARGYDekOLkhcg
4u8ASW+5Sw/RfTCaOoQAYUK1EDAZg4qNQsY1t+Ncn9nWPgDViT+YFubVVozB92KncemvL/W0U2tr
86E6c4DP4q2zKqX5RgIm3QINiMV3KOBxQa243fxkn2MjN5WEZkZyIf+qNtm4zMc2Zb9lffwiTL7N
KBJcy4E9ku9wW2f8pqA+MYM2JBJaub0bdFEEM69E113Tau9TeTmDAlVTBZp/2GCQLhNCY8T1CM57
GSIVE8Eosi739jytBL1jFZeGfd52DcIIIewzkoA2H9300jV0JgP7KcNxkYo6niwLvDNCOauRVpgW
ky30yBa8OSJ4RmdRenx4pwz7LPEt6AxoKsFZyS+y0TJQJoHAqmPR7/nO7hD+tcXnx5T/U7KR/h/W
1oaTPvi6PVe0gmjj7DSU23vCL+49ewGO3FmLzS89GOD8q+XeR0Abm9R6rgZW/RM6WeU/D8txEJFK
rU9ULr0V6D7iVP/zBW6j7LeEzOnuKjcetGmyF88ijXCxoZsWLcoqUqk649pdIgPLPibqctI4p9cP
MfHV1edndTVTrVNN9fnaEg63wVQv1Fnhn8MpLhvV+fc4wjymqyF/b3WO0yhlBEuXJZ8AxzTYVevN
b8I7Pl7xDenwlbzLSdwS7HWnSTsjzyR/nwCs8PXgy1f4cymcFxa21WqRxvArET0V//ejBfVN9j7i
s2glZWO3tzWWCL1KpJhIXmqVmCU6fZHQne8+l3sVBjoJKwsd6kRSjWhiEqTTT7hoHbJ0KscTNAdc
xmIk+mt30hYafsK+ZSnIQroGfjLbOqRXfDu6OCNgFc1oWvKvUmNUvRWRGeoOP/PPGrjV84/+YfOs
Fin1xwYYSs1zNJ+hFHBkoPKOubn3RLHo/xV2rwgnRMxxl6yxnmVT426Lnal9rSjJxzoyaLyjXRh2
mlKyHZ53yNF8wdANbXi1fawJXIQLJkUKZo2kqxtX2B+Jc69BuGzbyaZVrlScQq8mkV6xpBTVD2D6
B6Cyojo1wlD8a9kb3KSV8ii5D+qApc9d8pWneMYpHALdm/Yrxtgt8azEGnsvwo6SQO6j4dmUGmZ5
3S5duSRUmh9vhjGOw2coBg3PO/x5hq1M22NcXMDDoglQbeuwAHm2350K+7fAAcUz6YsBsVpYR92O
t9ckLFqAN17yPUuHIDqPUNNj9i640WZ4lJOsOvGCfDJMVBoFrPUaAyZ5bpxNawfM8YHXP26PUmsb
40WDGD3KGv2LkAdzmOGuszVnvR9wC2SBbIFwxTYSj0baaxOuVmagQrq4awr1/VQ8P4WLxXNEIVla
a5Lf7pfTVnGzYajSRiKYzgQ1u6MAfzopq8QQ3I2MgA22a8m2ZPWfqjDCvCr/W2ELVsYuiKRpy88z
fOzcabzkV4AvFPYcM8uodh27K0ZzA6I/MOpY5TnISy6DaXwbkYls97WzGJlgYCdx4Z2iJ9fAY7OW
I612kTM3NfxaYpTzQw/mOujTIzMqFvL/SutINk4GpnRdjgOVoffuli1k5NTf0hCa4Z7IS9RPzUN3
kP5SYj/6UuZywBsN/5tH1YOPlGJepCIRkz/o9/553qIF/48WwYOA23q+FmwcnzkOAqPX+r2KUGuA
IuIKinui8BUuMrnyKujYrMJWcjF6J/y+QK6OKa+0TI78jxtIPKX7rQ4mYLtphALSkICEI4UZc/85
xuSPQdw0yqhch7KlLGRVqOHmbW/LMhaQZiqbd0+kDHTLpKUe3CsRb9OrhQST09Ouu4/WGsJN0aUF
qisuALxlmxCujwsU8CvFSSRgDngxchCJUj9uW5++eaSmMuWYFAqUYszeW9b4BEtdoP2yy6tbYboE
ZRZDRW9Al1qQ8ZVyAuQVmdBuv+uWup8VXAV8G/5BcvhE9xa1FZKIJ7hkrTxe6Ldk5YcmSPgHCBDe
tUn2GR8Gwy6N9eZ2u1D/LAy9Wt0uF9AD4JgflhtMEwlw016i8KXBM6QNflWpTpPI61DV3v38wvWn
w7JAEYJII4w3+9Da/dB5RXkMPzmmoV8GwFmR8j9aM/L5oRfoefxNq6JwdDz6ye7JNURxeeyoXJMW
jtyWl8bK6JjGRGofL53mi03xojfKThTtbKfhBjyDmVu6ae9whvBgJw6um20gZ502nkYQkSpmAgCY
pBe8quutJkAfC3m/WbrGk3PlNG1ZRpbYcqvlvO7Qght4Fgf2NHEjuiAmTCKN0Lp3uZhr0ke4di/Q
Y7tp3ZNQzLWA7aqR+F5LndnijLqAafmEbhVkWm+Ekw5W9+JJwhBw3NqXJfcDpGpCT/mM4N1qN4V+
y3Riv1yhb88yc6T2HE3OoDi9Wj+eE0j1u25Q95cSRh+g42O23Wjq2keGIvpCdoAj2FLxBFNe7DeO
+Xk+l3LQYRnPBYRVOKa4KweEO+eTKpRGqrkUObh7kj+7zl5bxBWfbUyo/mVjZaRZiL2P47CaP0cD
b8KI/NLa909NTkvLs6bRGw2Svycge05Bv8K6IIDpCZo5NIckRflqVjRjWPNh9mSVMN0rZMi7sqyL
2IUmO8EPv2sEzPpT/ObA6sq5O+jDngKTOZCOtKQUSg03xs6D047+PRUGXpEbYYhyvMwoOeIVStEA
5JW6qw8AqrcTUxsNc5sOvnS3C6vwt84LTvfnOEItqU0spWWxfkXAzUo0XGI2M8+CbW19rlFZZfUE
YGqR5hIili4DHvGAGb7ubB7Z2I/jctDxvk2c/in3YLLrV6yKkoIR1YNU24TVEbgTd3Px1laseOU7
amsep9MYazhHtC1EbYRtqotA5O7E3YvuRpL6vv7D1KC3ZWhyB5fyYNF/0FkvY2PSzIIgb5c8hDn1
Rb+l1gYYeePBXrOBpKN+VdcgUr8g3k7jScV63SGK6L/Pg5ECdV9qoseh72JyADwR6ADBY5wMcZ/s
U8dy8skg65xlQ4Y5D/ML5mOrBDBCHInpR3SMneUPlz6oCrpwpG2syyvyXeJXNV2xiE6wZL4xVbZM
KupJIjB0R4CODF3j7kUHkjfmxyJZvSmfWD8TqRLPEvaQHPA+zDdfHjIOCCcgSvkPJAAJclMAkZGS
qGcX7OcU3tqE+/xgjw2z7jXX29rBOT4cfAakAjg4SKcvGFfd9tUbnhCy46ZH2u+TJqvXFEz9hw+c
KmBQzgfjcSPNig+JcpGeeFoXKPWDeNBXQdwcLLcWm9d++b/ATaUZhzcWoKvq7QgfpyziNEvtDvV8
ntM5tfuyz57wHUJl3WxJlrgDnFpPXEq+24MTWTRbthudKIhwVHhcX6yxU70u2Xr6V0kRgQWbLouo
AOFNFqXGyDhLNH9MAMYhk47yXDMvOkxJStMm37K3xI21tgDHqVAyfxapabntHOeryS4bcufXr4J4
SdVq8FveTV/uADrDjOmVtTCgjCK9T/8ppxCilXjvnbBgESIC0VZYmq96uH+rdcroGlc7t3+wan3K
Fd1QBleOLNdd+GkUBXRMK26xsxbbGx0e5dbg7tjkOF0X0wxoCB1qhsPxonY3nxpspXsUo76aLDAU
HItXu1+hNr1QsZwSLyPwrLEIHkb2bYn/lRIalskj9mWwZkR1iG1hVXmnX6gvuZik2qUzbNbW5Pv2
qKFssjAZmzWYGM/d179puACOaYtOqPNJtUo62x3fv/tNv4Tsd8s7HoxpEAcagUwxKRZBaZB59x3A
FzGTXN2AzVs/N36bN0VCQhAT8VwG+uh3nXoItLyc4e+i5wcsKoFO4qgr2qIeV8+b2gGfPxoXrGK2
bS7cx+mb6VX8nqeNzVNOcg3o4xAA0Qaz+WpvuxqNcVU6HrMLcS6peYBBf8Mi65sOcC5VsNPJ1wA9
2ZZtjv5bi82HFLZVj5qiXeFTxm/81zvOVogXAOc2DId637x0hvRT0FxPi5smlFnVyd6ZeTUzSHKK
YV0BN1VtwDIwmgG9+WTZIBBaElSFFI37ZAfE2ye6g95ieC4D3jMrS4B7LXjhsoIsq1nXa+uOW9Ce
Pi6X26B1p0phxx7zFoH8b5rXj8hTkyW3OYJCQQ9FQo2MkeP8hj2ON6GEZKzVnNew9aFZGsojb9Yy
Bx//kS5VRpycDudJaTxguyMPrElrDQjONmCgyrPenM4ijIRExQvv9NZZbNm13LoxsXnoijhgGjAK
WtyMyeMMGkoMWPbCbysVLY2G4M98uIJUs3PWnPX5brRSStdUCByU4O5zXbwDV9R7wVEQFt+W4aYk
jqpKn45/hpZuapdekDi4WSgs6LFAtmjF7o4rxlWXHCOmfb7kmdbdayj/P4MaT3KI8ZUyZNJdcfCL
52BX5UeLiK9ORtYk3ob2MZpXUe3pE4dmi9obE0K5eDbiMtqkQmiZtgEgIOLsrze+HKRC9KRN/zlX
PSvN9wqMCwnYE7G8qKFnspG3uh4f/Lu8/XVXBVnxeWB0SbFPNMExTERVeTppOD5ZUFvoQ3AYfTb/
56LYwExbRawwO8dNeGnrk9PjxxbtrQWaKWr0cxhX/U8DoCVycqnEJP6Ur/VZ7IUf/RhlVt/wgeGq
aQpTVRfjoK7OVMU6st2ec4X5GfWbrcnLfhVIDWs/sHKqlImiv0J1oHqtKrlxT5NAyC5jKRQRsc93
hmx5EzKM+I0H6CKVC0rGdHxnggFYnlBszlLW3kgZUXjRRBV5Rsk6DFF3sVnvWmKGLqRQBLo2haO8
se5ZJqePPRVlJIqXQQGlZ3SVOrwohHudF7fW47UyDcrbaQu7yFpmzaY2AmbGZxiuX2eYrTMUcyzh
JkAINiAZpf2+0VdqMBWERgiqWWi/esD0aWW6JYMVOZZwuwz/s8/NedPtzuM13Q0z18dPZGqD37Px
ZvHmn+fhWRGy+VYTQxoARKIvYUHq7wfqV1xZtNCI7pt7rGnnPlTvz2H6Ekf2LSD2cbcz23Q+jc/Z
Tie7+dFR+yMJM30zBuZ/I/Z3dgMa7VyB3Q3DDzYGf7cM6mCPrC4oC18m4yz56hnzi0vbUQsJJnue
pUpIwCjmtwsMH+urraY29r/WMKVCbNw5BDxdBIxPcUf52NXrwK7jXd97snvR6thUBxukwetRON0U
3zwRZ5u3c9H/2Z07ewj/Q8lBNLqbFpW5JC/f26kgrqMtpkgVlpqNWLxgQzWxYR2RN/Z3L60pq22G
mmVr0rMG3+6n6SohCWTGU4q1m85O+RNum8mUjMs+iOxFCXhwqBDbvl3Tpzd1kb5muj7yb2pMTVAl
QGTRToE7deFxUn1LJdEr92SMvXQjnKlr0oKa8oQCfqSrpangxHy+Cqbe57/a5ZNHrJlzrMxFWEXx
u8s2J42wZiW6T6Vdu0h+1rEied2UkBQwJw35ZXicTpnHECgoIUw2DrcYKGwsXv4birjW3hyeTfYB
GrgjvTuu+mof3VgMswXxggshAq1mUfaMN0eiWSSLbeXwBtTEoSvHpR/kZnY9ea2XduATOOt0PpBo
DM6k6CjtRnABjj8ItQstPXEC93UrWjMk56+iTs5eb8kkAQr9fOYgwPMlVkh0tYo9sRTdjYjcO/is
yMflDiuH23z2YzV50wZpvcqCpjbdpGwGedqDonyOwSwiwLt71+ZBYfUYYXOYHxs5RDSCsPHdT80Z
r2P+cGGr0kDOL72n116lCS+k5EVtJ5iblYVn+AKGHTS/hj/2nd7M0OJbtCz8SsBsir/1q2kS1zVc
rw+WzGAKGEYjNRNSo1m2AFRv1hyiDqSM4nNDBr8z08vhyJq/Dw4l79ulFswRppvaQSlwx3g9jc5E
GDaTevUcCybeL7sBjIV50Gn97qNnX/VXDOoKMA2R21JLs+Nk6YX3O792+d3YF4bpgM/VB4F/sA5l
fwxILLNLq4f87e7BJr1MxeSG8Gml3bw6gVV+EVj7e6F/nxPfWawpMTpuXKNCSkzdbheLHQpSU3o1
XRlefc8rRl+taoUyXgupVt3UxOZYBgRq8qEGP659fjwXGz/ryf+lsQcMqkZ1WHRJTD4alo000HC6
wIbHKpmOYnfCbq05L+BA8UeabxZuUgLqc1hf6MNVpddiX6pxr8n5zwLDi/WNsV1zcPTruFfwkBCw
ukOzu831K3DALbtkvt9FqEB06Te6ZzhmQsJRN06remlT8hvcUCLxOyVM7m3UL8JQF0GFXG4m+N+b
1+eV4jYfjXtutwrtPWqiXcQ7tisO51QOGQesPcqTxIitWwYAdz7tby1LFobukfu8HrmwIyGT0hD6
DOtK8WeMY06YysFPZ4EWbEHEeA6htMRokdR8zzObTQGeok6Gug6vRt0+Z2UeXI31gtN0MjY+xdJz
cFJjiPDJ2BnEqWFfaCWrMQIUtDU0ggFXlELFR4/VByx79Rw/ywb38lmweWAkIJLnxNsRgyvXYqBQ
8WdFi1/SsOqouTFkZPhJ4PmPSb7fP4TwR+8r27wbuQRfgM1Nf4LCwASng+6kMHBcyLgmIwX3NoC3
X8tBum0kidbAIWn24DPfY+UmfT3Q+m8IW89cLnC1IyTRNSx0PdZkY/wSUSPZMqCO15mUjTm+TBGF
tdrUSWKFJg1qiIWtDbO4Luo9QVgZ7We1fgCOERu2/1562An2C87MDTMPb8r9croKSgE0S33lW1qf
2luMdLnfOHCl7JfsFqsQDB98RRT5l53C3AC/yxqcH5/mxdfHAGYsVyVJjCMrzODDMPSiI6AhITcR
FiTyl4FO5fofEW2f0eun3fpVq8UTVvzmM4dp76bNx7SkF+my2FjoO+kRRZ7wmt6rbswAij+YCvrl
Y5a2nJGKntfFzkSmtTra47cH3fGsOFzD+WgMk2vsrEbUyeGezxRJPbEqETcQhQpeJOL2acooUOG+
6cbUDpYAmbeiiNLuX1v/W/OztTa0aO7oksuVwZzKkJCfNUlG+uwY61DCHSwZipmyizc2t+z2RyMy
d7vMzFqAndiFF2+NNX+Jg4XeYEHZJVv+2HtrvM55fuSPYVOu9oW65h/Kup4kFbb20L7nRtgaIyJx
o1yfWEEat46kX7yaPL5oVP/WYeyeQMpXcapGK+tko4Hqm5cwirg85kNoujdblCfPDQAPPD4fF2Aa
2gQgKhSnn2tLSiw2maYUaKJzCzLwGMKfGs2v8lJFpqzByBqYe4+Ho4cPwd7owXpaC+tPqs6ce+D5
4P29p5IYtJMy+a9zXzjN3n6GjsClyLEMWtK/98BfWoKOFwbgHJx0pWlwKl4bwq9pFDRyRrZEkAob
gHV4/ck/N6KEN1FPI43CFHUUXN5UJSQ+8tbfu6YH6FGKHF2Fp7w9Ru8NFAJLYnRQSSkgrAgPh3/y
z/IdYDTfHOXU+AwbmWDK22TKVS9eH7MP38xImRyW898DSDsQed1UbUqiHu0CTeE/7KniEbPFDJPP
0g4ew77ZNMs4cBn4MdpfcNS7t/5FJZ7xwHAwV8FJ+hS+rLtQIjz5+7IqFu+S9AbSLRlRMd1jQTOd
b0zoKchVmWh8Bigf4TlQprQBXc9fTcFxwlvvFWejJds74Sa+PY9SwwHsRmgFfL0xs3XtnPh2gaWg
CGqSaGlwWCV8jqZpRshE6DAELCfiK9ytNXGWzERgpmB4Dozgzar3zduvoVB9FmGID/lGABCxB8Li
zIfaKG6aXKAF5idMAR9hZagw8Ognb7D0A0HHBF/Atlp54zCnWrdeSjs6wp/tid4RiQyMr21xpwox
/oerlWkCNcQnS2BE+5qBxrRdtCC8bz+2uM6tqRuUiL9mZPsLMVSbryjVxyVbrZtfP2dPKBLO0HtY
/4ZVNhCl3DVgh9PfFZt6myYTyI8Ka68AzSgplrRI7/3J3c0H6sGFzNYZf/Vqlu2jysSSQZ5hRoMp
fRzYuG3s0rXEVdph2OGFjRXW6V1be+5V4zLvf6htuY8pXihlYakg+Kq7U4B2Hvk1rJc2WamFNXMA
delc/7cS5AgMt64hUjIce9Tu3gBPPXS0Z5qfMCOq4kfOqVbEhVrv7/oI138nnvCRBZHr6FpxRvOh
J9Ivtm1C0/wEItyXpMvpH68fuhag5QsMYomBZFa4MVOS1Q8SMYnb1yk4OBxCokq3422YtekCex/4
gzvWNnl0x9a9mWwzRykTq+dxIk8Xo0lspmp+Vrb1ThX/BQ7OrlkKRSni0K85uxZXaMy5ReTS03d6
4plohd5n3/i3x2dp8J3yHbOTPGVWtumVv3hqvVSYroO4NUX650AsZgHx8WZL/uQWkF3veYvhrNGf
WQgbaHzXl0ZvuWGxZfQ1hvog2M14/Ielnj7N6zHhVIwRTSzlkykHqzn10f/QjE+89yj8RgD3YmdM
Neol0u0r1qgOjAZuxNUhXB3Ek1V48cfmV6+VZJv+PXYPHL0gEq8fPggq2ktQCe6BcQ5VazzQTIkv
aDD1X2aalWzCnm8fbruoBn3SYYH18wQChjSpTqBgQ9zrOFplOq/V7pLtSrliiCngBRo7cYifsomG
MLlF4vAztftbaJ0syK1itDziLCTBoEIMG9jlWitRZW2XZPBen/gVt2x6LewbLsoS7EvaXBxCaMF/
4VOfVZngDKV4QAnItg6dkXbKwopYX7ICYXd8AAA0NG1jqO/rJpez1WCTgTX9xF+uuqeZkjnwEM1m
ckEnBKHZq91Ch+2exA2EM5ceQI1mlVm1sLVgbx+m662aqLJIOwK7IZFoN9HJtN3U7SY/qAXDG1I8
Sus2I6uMwlNYW02t0inwV7K51UX2l/Po8I5+qteKJ0vhMNL3K0IyF/YP0ScCeBarbqndEE3WZx6K
3AMTnSVcEJbjyZwLdqFTHlG+NT9YngRcmVJfDo9uL1XZm5ogQA/MDak0dOUhFwDPOEJCMnoglLc4
h4qTCA2vhrGleJRTo4y+9x/m8ymfdnE6wiPm1CukilquYhexFeANO1zbp+uGoJ67TBsUNH2YzHpY
hSrLaSpyfCp7yM4NGK6YvQNqEIcFhZ37joCeojSOR6F36S78Y5YggBY/g60tciFEKJ+zFuhXntBd
B+ApzPh36dwSuAijSTgErDVHCftwrJpYOpVG2XO4sDcXOAC4raqWw0T8NashIiUjpRn3QntOj/wA
Iem0ijUUcHCwLE2EMidjDGjp5kUkC61I4+1quuYSrc/STKkeW7uwSvAwfaW0e0IYZpQ2v/Niy9ZD
J5NHTOdK/0xtUYLwo8nNyU8QNYYxZ3Po/evb68ERZkvsh51rXGuI3H220rE2xE5qt14u9VozyHo7
PGPy2E4M/uhPS7Pkrb1bmC3wM5oA2p07vh0oG0q10xeUUXN/kFDlWz7+vKv6xNajt6z0tiPB0SqR
K7hxD4zkFzHvci4OZlqLCSEeGW5aHcRk76Lg+294NXMALKY0IKR7Qx+zdFozICts2WOvoK6ecGRM
yTGDBVoR5TBuQXEFywGLUeoGOrYBt+QyZQQ5au/lJ1pWm8gEfnO8EJI4R86BCFHLujjnYaaPvEdu
t7az7Uaaxwl5SemAqSn8MBt2mUTLd5RnDLoer0cpB8mBdQwSBWmzYV6WuAPEeDOlgbgbjKUmnQID
3Hr637pzWmr77fIR/dWQCY4ECcYvyYJ7C1tH7XN1ZxueN9MVfxYcZRvrqh3Q5AxWR+nzZFLAui9C
55qBVA2ReB7qpQyfjk6Sbljdyi9nSBfNgb8dONVuDX3AraM/e+Gz5cS16B+calESMRIv4dGfZXuj
PFhRp7AtHzaOpPKFis0Ocib6WPidc3ELYVBVTVoqz16tDmvrv2wkCP1EgZa29TDjoAWDUUtDLWMv
qH97bU1y4236OjTKDcv8hCPKquMBwul/uN+WX/SnJA6/Bg63poC7qfJZDRekz0H/SN1LshiCN3No
unXm9uz5vnt8uk333E3pKhhmAoJ5K2GnKvvQlxf8cqZ5ARGoNNI4U9h/kG+eXdrKaIpEhoDn2lBQ
W808OMwfzNnpMgpDkSO6IImJz83Kp5biKCUSw34Nlytbc0sLPDe6NviunJ79gwCHagbLStnKtn2j
8TT8kMaBo0ZQr+TsNDZplqXCVmuZgRS4uH+Y8qxm6NW08I6/Uod2NQ6uZXlVTyPqcBjGXCftLb+t
CQUkZ1GfH9Pwgh9m7zFQGEqSIehHzujfnVUa71nKN/VxHtvGA/TjNAHdLvWvTZz2NMIsdBbeuREq
VGptbVzWnIkKACAl0g3WUNosp2Dxy1oCrGbBSd18J4a6ZaG2dRISSoq4OU7WJNsPMEt2QpdGWUFp
paEHBDQUmBMUp12izGEMF49gIQzORqeXwV1Mz4990/oyEpDv3+1t8AEp7aRKrTsfAGH+X0+a8oEk
JGBuKh6qKZ8axX0ivVMmg7sARgdQL1WerBSsjqCrfbocLT5QJ/oFmkZYvexhWizD2ZEc4466KCm8
gP/K0DU2/RXC4mdRG3Y7zMpI8y9gn1M/Dmb1azmnhbFuoq4wjenK2v2XeLEaFHCcjCXLptiVi3PQ
d2AtC6EuaMrEOUtJQGMrd6V8suUFKsqz7XMqvL9GucUUhYYEKolezuAJdvj1dkn37xrAKoD2nNXV
GgFw0ZG/I+Wj9s9xb2Ghpa/pA594EkK/p7YzrqlfhIsfds2AfSMq2Vc+dWSyHsgF3An42gfpSsOy
+4KTMmz5T5++7gqIaxLFhopu4LT82CdkoyBdvanLH+ryElJmFD2m7E8/YQSTB+Grv9PaWz4l2nHN
IBJvJvDakb4ejyNin3dERymQRwR4GBxYl0TBG1AAVRxSQc37KCk9DYXPqYKS7ZeKEBStVqGsR+s1
KEmpc+P4hflm5YjGXZVOgMmojJbY87DHFoJECvJ23sKaB1epnqBrcYb4VQKGAvyBxcHpF/eYO7CV
ykoNUvRPAkbG9uVMywVhvwvshtvX40D/xpHIwuHeJI4GEqSMEkbnOFHp8P/ZJAwVlfO5t3aZreNU
+ZyEgJ7LfDbu2ucNJO0wIp5Y5t+bmUkSHfWLa0UHPoO7GlM7bShpkLXNRmiE/3HJ2sfXRHHpOgzl
WdrdtTEk9DGalOY7mFnF9B+hUS+d+efJISE+JMi5bRKeLo8ve7yyAC19J+oz5maR2RLTgDraaw4z
iHpJ+tu5fTOsclBmLcG3zdwjRpqvTH1ZRU96zla9whZcP1R3MnojbeqaQPHgAkr3a/X40johuOj8
0SvF29V8U1mTQzlUfoqZldPie7Rwx/Rwpuw/WR25sQ0FipPOMMt7CfvztrsY3nOe6KNe+xMMm2pd
r/forSVO6GI5HNJMJEGvn9ytO+1EgFk4E/8VFKhR//zssVsEjSD0UXICX71PneDugYQ9QiMXbAKp
OM8HcRFiOxQR/fGcZPg+01Txj1SuWtPP1XUuzMwg7mW+OYdlfKo8OX3PehAePT7Xat807wO1Cm+1
Eb/tqX2tgUdKKNM5/9JPDK8KxGTgwl9rnjsur0l+Cz+JNko+uqZ+Z3UYwwGUG+x0utaUWObaRd+v
QUctKR+D7PbLoDWlxQrpqLxjPxHD1TMctVM7bSZ6RDPlBMaTUMS3IzWRIZG8507RnuqsGUx8cyZV
4guRv0cWj7RHaAwgfzgaUFoYZzjGybGVQik/bRbzWQoQNAGEWl1qisTu16oGzEUWkT/Q7dz+ivHU
YYVfX0yDxo4dvAnKDqPX79bmxnGjb8wCKKh2oDo6B+47e8WF3RzbBEDtid0UVn5Vg3JgcrVuBDM3
H/PuVgj3w6rhiwud4xCF4DVDOqx4TMVG7vO8Jz5rFO9qyNaAuaxNaCPMiIwUlytiVcJVYD/X/frm
j6zseX4OUD3tt90TFfkNYruuHX8MTVYlc6kHdeqX6cYk2/RnNW+W2B34lqliIP7bQYuUkalU8m3x
oVQ1dguk1BZJAgTuN62aryrYkgkzy5gB+IAnSgj8yaBJAM50QT8AzyASbCXX/nabt+n6033RmexR
xI8xMQOUE6UCPdMYySufP65N5pMqAGotHkNkdtdPkt9cwOSvAfZ772laTahwofkrYarLb2za0wtA
oGl7vSIqI26U+NWItSFScyqF7wgPXrCPw64KG+y+YeseoGy35kRD1TtUtjgIByLMUqnJH6PoE2ti
5ifdIWhk4wcZi04uLCYZst/WDLYu3XpdO5++7Vd00RJMcxSMrTf3EbJemqbYKF6K6QjPa9k1J/6C
wIwNapuwY4ZUsR+Nm+G63W1X4/t+UHaXdOe/IS7WZSFkHH/cdpI6jKUWg57blFbT5I4pz/K8AfCT
20f8NHldCFBg1os5GBES97fCaOSc5c8I7rH/efe8HyPkBWiRoREqekloA2RLGxOVCWcJYBwy/bro
iEbtfc7qoEUdw26o6QZ+TyqKJDW21L9+Wlc5aBVTgw/ZhbonguLObwN64Pc6iOfQ+9kyhmTI6kmF
TUdi8YDegzNR6xadsriEJnDW7kJ/vDHs5iltAm0TMjWrxcOqVL7HYDd2qxnec6YV5yWGzEh8Wngq
TOwGoJ/Y1yL2owJMqkgwvxLaNrY5i6PaCee25fPxLEQbPcFoJeLHZPO+6zZcuUh8k0eNWIkWaUJf
HT7sbpE+RQAz7bexgVdgOofleRJ+7N/Xezj8F/LHlK3Mb3eaidFz9DAzic/barW29B/m3rO75fmh
bnr95W/Trwe7DMXD0y2FcCa0N4bj09uouICEQxgCwkCU3w7bv/hHwa+0HqzIiGRQpMjEzPRFNJFH
wWvbnUmnrARaWJ4Wd2q5hcs1T9vNrEvsbvI09K7RqsKX/ZZxogK7b9AieFy3Kx8tOuKqYr3rTlvk
+vhTfM1xMIXxtxa6ZM7HPtF4rlMHlGevYYWr64yh/RVe9EagWfF2bJJkOWSEW2c5LKfaNjhFsSk4
p88E6YWDW+dvKR84NE7nVW2aHa7Q9mwHqw7VgoJ7yMqYmQt9QMhiPv1qWTMohd8cAKWWfKDvjQ9+
TB5ulGASoa3ImtI1poe2FquEHOVaimQo84DnuvcQGq1GuJbrmAfYzoSN6gelLeW2pav6iIhi1xyC
7RISB8zGZOLBGQKqlZnuC5QF68B5ViRONQhffsB+CoBSiT0Vk4t6GTWY2+y+2lQHyQ74UvaUupJv
DSkyyE6LOILFP7RX8rUaUQmn4qJWjl4mXQ0OOegsFSw+qfr3WoYvunN5XsetOW7qMHkIjltjUOP4
HFfyR7CBxrrHSu9O5dYBnp3UxhjYzWY2q1tf8XvuAi/hTRAuOLoCAdE45DFTdSQADr4WZUtZyx/9
qVz3JcM4YquQIsak0adSL+A4rVbL9mDDpLXn5lVZow+N4nGW8fgdrVWymr8UbzmV9wTndpABAmKa
PudJR73C5ZiaEh9t2gfHnuL0cUvtgRq8zcdZnSJZNwlZmZplcFmnJAVSiV5RUJbPhwQFvEZ3lrxC
wbOkgK2HdvsaLmm7AuNyIRfsRNdMd+4kNxPkXFmR88QShlU7ZTdqDG3p/Xany4wp7RKAqtIRNJeC
Ioh7PDhNyzNVSMVZ50MgAGqLhnpvezBFcYrIjARbEWJuj4Gz1Uf0MjSKsl8poAt03x0QLY0kdv7X
9cDpTvpSHI8SN8pJL9cZnZS864jEA9SbYcWcdxj9WD1fIn3rlt3wXXp6LbrYA3okaHE/BIFOZHjm
icO+20+QX1sG5wV1+WFYHNEaYkoYdk3WBd67XmYyG9byKaftAMC3H87YhB1H/xoMDOdJX3vhoD4m
EJLTZ089F+apkQ30RBjYs1IltZ4/pqAe9CkDX9+yipbgQMqaTIfvGj+mP67FYdHaukul6E0fJ73z
D9f+N8LwslwhLE6l0jpWcShpU0xHXSKGksnMO+IQXajABAuNcwspNa3QxZznwVpDy8Y7+2K1u87g
3cavYyhuu+tMVUVoZrqd+jG6qxG+rftENvNYU8S6FHMty7OaD5qHLDtznwOwWppmILZC52tD8QGb
pD9KT2WdAwC+RRaa39+F4i4Ev5pQwf/iCmtkjLgQw1QDC8+K+z6Yuw4uD/3fmrNKqHEJ+154bqtd
bRFRqznsaikEnGT9AQAp3vCveeEn03XrSLdhzE2C2TfWG2WToXV+JAkd6XSrHFbmrem/p91+R24g
eqxHwvtQH8LeZyCJAX1HBHYmT9hj5O4Joy5RqU+/W26pG+rrPwJ0pBilcZCCcjYopb9q/dt6eNVx
OlRqic9qTWzlDc6S2Iolmi4y+OMOdjoobYJpGWEYO5Ef8TgBRJVI4XpPTP03HK2THgkS3qQ1IyaR
GXtKYRHAjQGFhadxWfH8MQU6EjF8CQ6kV94bltiD/JY/+kcJZE5OchGIuJLI9DJ6Qh+ZtJ7TzsS2
kKzCKEJojZ82eUO5jRgQWpqg3KAMzvTC37JVwp1VkKj7fSCbRLgKdpEl1ekH/zjwzYAbwg4c9izL
LX8fjzzabPJHWYKxGR69AQNAcKEOpjdvZa4B+1qhEz/UYa2jJS3ZYT8iz/Vi6qr6HIwgI1z+yPG0
PARWrBfFXetasa87xUj4kZTcKTXLncR6VyWxos9ZzgjAXiwFFBc/tD+MgsHTnUtEykle0TXaV9ee
VTtCt1+nUUogCM+9cRh5cdBMs9ktlOtM1PUiHAu4gnHl/K7C8kE6SwpMNQ9s6brjy4/MezOuRNmk
NicIhUCJs697/sGkyB0KblpF/02Pr7c36HNeugb1CbvXA8CQTPLdN5nQGEcVDPozaZXwN6eX4rGW
ucpHs5M0TUfPsDGg4f3fNQhn7/T7XzBRfFHRCNT4KGfEpN0UtjGdr0GiP23nnJXKjb6wenfdlnGD
i00984iHXRXJL/q6oY/KSV6MmD2P2gbitp/sf1Fr3TZ/Xnf4j6fpqyo+ses0SJN7ySPSsOu81hQS
sP66ufIXMcwFItYrfEnC/6WmchpxKI5BndmNreKEGGcYNX1uaVTvIqeCk4R/5JotgapF9Xhi9rre
oZmB7VD8AZjfpQhbqjf5604g6LAH8kJZ6zzGDwE1m8AGexJyjS7VruVdm2FPD3kqRBOFFi58bRWS
w/bwSDgdtv62w2xWkPKeyZWmyV1QHd3rjesOoWbrhK86MA75s6JNNKEpvk/ryE8OqYB3t0X94Lsy
6tdakAQM9hViALypSQf0W8Q/AI3ac6Mmi0K/n9BZnNCHUYtM041SBsRKKiE6D7D3qRViinaTBKp0
qgCsqcc4IuZDxFPgRfMZvhKIOyfItRvpTjnPdZVtodWSePb86bRLAq1zP+KyfMH9jW1lOeu2YwAV
zJmC2umWuVl6DOR6Xy1BwRJfBU4Q2PpE+XBfH/AnGPxn/HSD4Al62fvGyP6MiZrIi6I1wwhGMd0v
HuoShYAbFCNMAFhiRIlOYUH0vphc8RPG4O/xmbEmmmnW6wiSHW1B712S/bn/Y3TXnQsLQuV7epPv
R6iexcq10xHoe4Pvf1oghO3DwD36zg+nhfY1W1/c1CBp/Vi0H7ov2kVwf8oBTX0C5C/HrkOUGqnC
pvfeTnN8kg+UirapQdrsm2jb3lQgM99D+TrEqA+aPM71KnlidtEUr27iCOUF3eiaPzEYaHx3vHf2
TYt7zGkqMkqjRg5StJBrnchiQCUOk3PiWdK7/DXSym8jMzM4rmE3gqsNRzA6AY6iVEpq1RrHdBLo
HTBRPwSczvF34SMVayIw1610Dpjx7SMw5xd7+w4Z2aYHs8pKfrFMjyzxaF8jDK5LsouuazQCfiqE
l/46pZIulSyjA6vZQyn2Zdf/1rhcjpTAKgVVGoeBXv0h5yWLyaTkD2f9OkWb6POeYJPONmvnvvj0
Jm7GjpoyqvR8vvyYgwRm9zmXnsH7JM1h1CxqRXinr/4/ZixXH2IJHFrbiBakMbpdlLH0EtnI8YQR
SM71FPXDBJP5+NjRrb5mlWsMX1C47YnKDUjjvQbceJGBx1g9NLoqDIltwXZx82EM9O6fxaGJ+SZa
QJXWFxjz04sJL0vv3S+XPFu594NCqEBhwOMgdx2B7gBdjjp+dzM4TX2hqFB3Y5p1zGPmrqKy/0k8
05xkul3pGeOds8uZHD5UIbiNJx4GgmW/ocuaNptsjJKIUCOVW6utN3OgmcnEJ/RQtmLbBXI5Jgke
FVjTZpfBim/ACD+ohRilto0MJVNezFobQ7+pueJZz21T4/joQmuT2JdSlBlFyyW9HdahkfM0MSqu
vVrFzooF0W1Ipkc/cmxSOuGlvYR2D9ilOFybzowrU7GDuaf3Nb/UbAEMcGlB0Nvj8Np8Fyg6189r
YyeCp4JPV3aB60oFu22Fhfl+WLMqTRgOKW/T8VRXwF05jncLd5UiZMdnZwxrSEV6ZHUQlAk/4lXD
ZIA9Gfl9euVQBWGAURc8KeXp9RTMKm8TtiUkyq6nZEb+g1QG04Twx6wNT2u5ddWVznhyxzx3A1KG
KZcjd8ord61V7BqNXs6oDYK5yltUhDyKBqXrQ0LAYO4kyjAbH5sligHO0sWvcGkX2aKk4hGsJEMp
VTDIlb33/XDiSUPvPwXWJpuSpqGs35ar9ukWuFYP180BohrQX8eb8yeYu+fmcUBVZj/ZqVkyQ6YG
8VoNQTIwA471Q4FtKpEWmtZrtQ9TBTVNqQa7pmcsK4NPDVT6LF7Z1Ld9pB8ghsuOrkQsiX9qyJGN
hWZlneUp3bhITvoADLV+BzpnU9Oltpx+LHEuC6E3aV0ehbXfpIDa/WLYrkEi+EmIJ5Aa45eKAywK
2p5XhHaEZ8c7iA7lPItxq5eqAdVCOo6K18OI209t+pLCNDWI2PbKlKsI0wQn9jGqaJbp2WLh/MMw
xcxan5ofP71OK9W9N6e5K76t8S9oRzTAajBlXZKGqB7veGQ4tBKzA6gbr57QoqPIi+WfxRbtcHFr
yvlym6H42QJXgNtSrPCsrOk3qD7MEMNq5gRpb6DgNMbI5W/EincJuYSYF+JE90DsFoplPobGHuR4
EYBHptS8pu0FsbpoBCQ3Tyxt71Wm4EMfA2lg21+nJdV2HRAf4K76wP6A7AR1mAOsMRFf8l224RRE
XsihOrii76+8QNICU/4kDF8oFW1FIFJFjJ/zt30krwwLDXY5eGPlVpwKbKXT/gzKSGS3I40g8Key
x5Rc1PMBIFqTl06KV8fQ3WsMKdq/YI+uVxss5l/GZLM1WFVD3ws0V2UvthJdsEYaYE+VbAPR6fdH
PyEoT3FGRHnYKd8vjb0j1+DmDBJUqdtvVegeWwDMoS/MHRMJ9agRwxPhqM+lbE1V//XidsJoUIKs
iUshSNUpbit5futo8gAobm6QXRZnLTAOMFETae57sgAT/usD7oPM+3AIMRXNsb1h5QlFhxNxYVrD
3RGI0HmSVSHYy4a0O3jOmPxS9qjE3Xt4+mJHcEFy+Q8j0Ski0tCyJyrpFQUN9oxnNFPP+X8UMzxK
/lZl7MVDRSRq+8Fwtfbwm8PhPkusSHy/qPhuW9vlq/Z7pMBQZgIRFxQ/B+hKL5paSnCeZr0ibF+B
8hXG8Sq+iHtxQP0R25EZ+5cBkVzGxKlcvFgR5Hv0jRXUAQdsug8GQdpYl+h3h+gxveL56hYsmpZP
AKveO48G8VCkZLSpZN4AegG6v8Z8qMU5tcZIuFQhHr8ZyqR3bYOXVLzXTDSxL3PP0cM7wrhN24Ya
ObRbbyLyq3ThH7aZqFWXiO2yCUSV1pbrcFxtlsfik1Ct53BEbLAT+4Xx4PbFgn4TfxEUN4H3Xo3Q
XlOWwvb45951vfMX4Hdt1ZbjEcOpnkt/QmgZGTVV4XPVwGNcfXvBOy9w1/VWlI5sCOABva5TaoCS
RjwunM/HwGycq4fDXHx34UCXxdUsWANdJlmCs1JLR86hmJz/qiSW5rZBrv0ZqW/yfvvoKRkGXhZM
0my7MtiKOx9Ysnh0hVAljEFKLSNgNxrTt4Vl7mdpomcwm8WL4gmd3ELpMxPE+FoLTnhR4JkSz75Z
urLA5TAcHV8/Jy9B4hN5i1R4YxGmccsWCgf8fizxKB05PHluWJyJrcVWVPb1CPDzocZVaYdtCgVm
6xrko3WiehQPR+vlXpqhybLiFaV434+GUun1w3Jz2YQ5kqTLueF+LfeE6ox/1AK9Wjt0unwbiGLQ
5nTiptRgB66/OXWT72K/HTjVSIUqzA5EEGX4LiZBd2qokrJprgS6JjWBCkeeupvFQt6u3MVC4ZV5
/a7h1u0qJQ5xZbWaNbdJOCO7edworPYjXhqOevXbwaBHjATHYQ2tUyldDf1vQfbk6EpgMsT9mUDw
4av+iw2FZXbroCMOw31ORU5fYgL/HfXiLkqXOO4VHr2lJk8FlwENMrR6wHgFBtoLSYSk5Gdz0lk1
J/b13fYXz2SbcqgAIXmtqg6o7HUHD9dbi4ryZXYWFlw57f6LWOSXQS9LV9emgs/jci+PCb3QoQcr
YtuhPLvueVpFoXU2cDJTcXYO5J4k+TOhtnCEmYGLwYuZJxqrHIwb8YT1t4zhvE/jvToZxGMCc3n6
BwRS8LDaSSNdLAYQlm02IEaVSHlLz0qRQsj9ZyB+yIUq419wfkTKGaptnIYVRSJlc8Q6lp9ypAQJ
Ro6Nx8hMaX/KiwNusuGaD+qgS53alO25e8GMjPizbVFDsw77yMQwPjnsixgDJmW1CyFxQiOc2rRd
uNAbjt6m5nW3tQddKV8iI03mUvaoMqufdiK94u4TIu1Rf5JG9AEDnkciIVNR11LrSqd3/2jNUfuB
8UeCqCw0zdpdh1CxmFncW7OBAmwmMdcVy3obthhYFZytvYgzLEntDvDHE7PxI9oG6olaUkYQtIAg
kpCL+b4UltgMlRowdJdFW4JZHFYm1In3gfzJG1o0bGlU3bIHTm/WbYdR3BxQUjUCaVJe61US/M2H
sibVsvIv/akLh6sJA9K+Ie+F1bg/dHX6PpjdQJOzlgFRlrmg1AVoXhWHrIyuItxugfoKP1pQ5Lzj
gvAP0Wfh0K3FZoyqdEV7DQomEjAVq9l8vduw61hbLN3EKrvflqFAaDwYozghmXFM5Z5VBMSswmCU
6mTek/GV1Bv9217/rbBhls4gfPBeqkexENrJI8uOH3Z8iQnavMPHaE/1RoFe7kxuwbxLSYqnjZqk
NTmzOcbsc87wfMXtfTY/IdUL3t15hOSZYKNsT8LLip/MYi6pqXgYAKpBSDzAv+gBX73QI+UcpjL+
ObOsEkvTKx9PMTws1T2gAU6s2o8BTVFrWDbz86ox2gAd8iNzvs7MiB/L0pTWnNKMYAfSGO9HFfHK
Of8fZG0Dp/qmNI1PqwX/PTDprS/5X42xXKKYHJF9srpz9QLJO/0JcN+c20F/qpoY+iBXXN4c6aFL
aN8W99huVKdlC7/iK0Aacvn5yyybbVly3oi+iYp9+DhQuuWKVrS9pXDPuG/PAWH6C6FuJR5b3Yvm
Fb3vl8ZYHH3AfYusQiKXpKJAMbggrhSjG1my4l1nk3pYD2KTRr7hdfrzfLBrubd8ZTUOZtsuRpUR
ZnI+mIy9fgC1i18ISOFAP012kivs4Rp0MSpxf7YiETGxL+g+xjiYJggjsGyLHPJrh073g2/kQasm
ZaGGIrK7aEB1J6xjA3IvLk3DKj/IPqfU5j9beNI5o/T3I0uh3gVnWl6dN4eygBo2RNF+IQw+NJHo
h/uNRo0bSbbc+31cdPwKodmUaLUcHNknFpSh4/xnvN9cZgm30k0BBXvIhGNTxTauFcMKB2YIdNy4
Vsrkowzna143aGyUb+hAqhF1FoBhyvvkrYsTDPzLsIMCI8Kqwc4T65O8cit44gU9luRPDD2Eqt3A
qsF0sVqR1xNVlTlRstzFQtxqH+vFt/weiSJxgxffztUinVJhot+k1UlA1yPDtKVGViqqj0ZMf77d
oYHahMNi1y9f9KxqB0mDQg1yYd7KQMYgrAx9DsP7aDEKh47MwY3EmlAylHLP8CzvnRh8l7K+wKZY
DmdIqbS3vQzw7a5v+DWjAEO0+RkXfvIIOvYW3fOhgD4awbasE6uZVNS4f3fOLKqIrwEFfqscz0ya
An7+HwTjxygrvLWK0iEBDOD2mCOynLwvKy/Fi38wEe+aIod6wY9Ni5AYGiXHnb4dhPlZyPMNG5Id
qjQanlk5h+XQemAOBXPCRsXTafFRpowc5p6JpuzHy6V0oTZXcMtII1ma1oNE5Cyt+L+WHxOQIkDh
5oqTFCDFfR8YB2uJRYd3/yYuhoz750QkWbmRORCtC1cs/+oxeShUz9I8du4fOv7WjfyVLIC2SYJ9
hCGs3CWngCMZrFWXB5bvr9QkULsrQx1dgGjXc2JJjTxrYRVxBlvloS/ylAuuPsrSXKOhAbIciyD2
njAzkxBsIhyQTXdNK1BExbXJUVDf2wXYAt8UP+n8IAYnm8r4TYApEgbCsyzpzWGN6uRdR4rYDhDp
MQPCK9HXECapc3HKb/4nxalDoPr41RL0tPJ5BcG0TH07ihTKaUpe73ikqFW09HnCCZxy6JTdBzKS
sKHj5JOSK82DbtNcmRzD00vqH3DZ64bMY8ptsxS7fEsxgYTozGG5nXqtgucy4sp36MlY/fWaNGuR
OOS4T8U0QRPaB7wd+l4eoi1oh3dW0vk2vmy09yLxcAkxJgjCE/SHSwwN38cb0dJnQQZH8ccQ2ZGs
+kVzAdvmUnS3KpZkpuTGhg5JyMXH688bDzyXFfZId2naRCIpPPKOCqyKKNcKuzvuDWGAttXgFXZw
xiRUUZ/nJtmgmqju6FjOJF7FErtdeJdr3aaiwAASaMJx+3Dg4Kk3KDnNE+Eu/UNMyAbkT9SFoKAO
yT+cxerO6smKwiBGtOwR9Zny4+6Sr3wXZ6896ZqOuLpaJJz1GbcpXIq63ChKYUzkI1K2mOtjxGna
PsIgKNfsWCjblm9AMW1sFCUZB/IEzoZm/zyqnbgZEukZM2G74tdkMIoiUVYVqYfPbk7dfEGFZUEz
SACuE9V60Y1cgzo9WAx/AKZDb8dnUhIn8eqCrlrg5U+DPw+aDq3ZjJ4cho4ehXi3NuF95ojSHGxB
PYiVtwWzHGBAkfiMWT35Qe/mUNRZYMQxxS5y8zbv8G4AL24as2slJhZxp2ix+qyZkuJuRhBlCEvJ
RzChf9ohIZilbHiK6zAsPgpEstDmDEdOCAd3adO6KzfS+xIdJr4GhttOAY512wPP4nR5k/t1MD7m
Yn0uQfLlAICogS3mFd505vKGb1Xw/tNiCnZ/cfXyRsPE0AjCaIFmN+prZOU+uXtKylGGdyzcJu6s
vPc+LLV3f2uB5hLmmLbq8X/YpwT44ys//k42+X7Ny3E2ybmwBk2A91y9euHLqgKFjdxswwBaziEB
7jgHcySDlv21xUNgqoCBOsciGhnMK1hpx8AUIb4yWeXTvfOmCT4vhaGwh+HpOZXpjQb6LCnvTnAK
v95+XHPXzSjtv/R7c+RD1kbnGtbUsLX56u9NaJ9AieUCzntMYCCMsT/Y7zi0IoHcCmdb8nTVSa9X
JL2nlOo5xB3FQZ6EXj0hdeDFLwyAdpm8AWSkTgJPp2mZ8ylgNo/oeDNePn8doxaGhi/mA7Rxf2kh
MvommF4bPXc8vEzJiW229kj4qhpQ6RuJ5DvloFytV/oG6GFk1/6uYVO0O+B1KwcVFdNSpoXqa2aL
/mKgWgZO5JZQZbXypy6oLL/s40Il/lTCc2f+3LsR6GG27VENoXSmV82AQwQ7at1p1+n8e6moayKA
d9NrT6hqsZiuz67xCrs+Feel2bHWFWzxg36MUGsN3JNzU+iJ/o9TOxlz60qxPnE/lRY9vXCuOQT2
nUKDfekCZztyq9MQmvJujFg6+Otxk/m7+nIRuBGKANCaxdqbn+rw5406g36BgHx9XpzsZpRv1owz
tyIN1yD3Nr3A0GdgeuGsDVIUqN8b55GU4WrRPVZADMonKY6sRTwiopEoW1HN/gcb2dkulH3CyS61
SqdzoLIPMQHgs48PLCP3fNArVxc01eMb4zNdDq4Le+LWhAcRByLWIOIZ3VIm5eSBAH/JsUpd2Era
AU0XG8pacCag8WIlP9mr9QWoHaDCp2qOeR2vFH07o6/vWJSP5sqQCWdjOdRDd199CRP6xGxEMgIJ
EPd6ic3i/ROH1CD/4NsgVt7CPnGI9VL9lUfg4dg3qj8D1VdbS6wAYZFY+rXISxFDhpd6vdIzWfP8
u7VThOCnjyimzLfAK9q0DgjULNFoCxNYQGpDM8/bVEmi3BT6Z9r1O/tCt3r+f9/ap8u0jB1Bjsri
fw3UWx00E4khWqHTX87CqnZgebr8kegm5l6FyKLcQvVbKi/jXmP5PfhxAuTOaS0j1VxTun8s55/Z
Md68RoVOjJMZtrkrXVHGcqY9OuItnH8iNIfzOtyIwrORBK/z9s0UhtBq1KzY7btanFSaaXvDuD+q
Ucoos9j6Lt1N29+ZVtvdaQYRNWBK1SekJFf/lSoIoq/ZVE5iX3OkFuxwf3+cU9Z284CgiNwZFkjC
Xsr85GQdXB577a94dMc3Ss5IuUuo+hR7ZCjaSU9AyNG4DOZaadTYeZj1/9LfK65+uBcllH11a+fh
DIU4QY3egykq3ppjCh1Nw2RX62QGH//clS3m47/PmgbSB/G2R2yE/2S5XNcBrUsU/s3tFL+GMut1
czQj6VfG7PSbZZZSGGi6xIJgZEPaaRmIqfOgM8tFx+/VOWYISr08bxL6pXYMx1o8qu+K3BY/NBDo
n+5DD22q9AsIWbV6Qdd5RCPDg2nwRVouiLagENFpJxDgiKWQi+pW3n4G7J7G6a3FSkNB0eGjc0WB
Nv9LFZdg8xKeOzNZSImD8F6kLNw9F9HentT50jTAdrRtsOy4OpA7mZkvKge2DkuLC8SZinIO7ry1
/u26lx8Vaj0cyKu2TDN/TD3T9YEWv0WzUYmUgOjvxC5KxhFEVm42jCNYFCZKe46RKwAOVtC/e+al
iuczW+5LlLRfMCa8d7AuJ0AdnLLr0mkj9IC/7+qn2u0YIWXcx/Y4KWXmwrCC4rdTyNUaEGhgtSQ7
NAwjfJlkjsO1Dw5KUtQOmeBHx7KiEcK+R+ep6vKyT/6PeKpLlIgTMxwveWOHqa6IYlKW300Wk0P+
KWLIBBFj1354ujJd9snrJ0VNOga39QkCBZoqwXI8Uz5nmx7QXXoEiWkOvc2KPTD3T33yzD4F5DUf
g3Jx1D8Z5W5LmO/buEtjVnQmqHwwZeZAxT6ACU/rXSJ2dGGur46kXftHp9r9RNdYjGVuqR65xzys
UCtkfQd+O3CF6AG2vzZSK9aNxoLDLGL32ydhWrSDt+58xejgrqEqZh+t22h1OCBhK7S8klPO17/C
0as0JuSxR1nzwtO3Z8MhEUCrDntTAO+GW4rFfvjqnqMlGfztHXEbo63ORHV8dADMSFSXlTzLS0KD
ktKD761JsPfzrBncFvcec5ct8t6YQoSE24pZAruEWWnVbAyHd+hrDhV+tECpcirSThtFMXPXTSMV
TAAt1QaFeu3RNEs+9aqi1UHjzYg13TU2c/gsyL7l9wPnKSrvISAyMfys/7DA/2m0kqgDoOQvSX9O
tyQh28y8LUCLO/gx2vILz67H2JWR0h7kadgcyCQU/BN+ssQnMcbsQxEUXZecIvxfnYQi2vC9gjxq
bQiayUU5cQxLkEBUe6raS8cZAf4wtoPSTOtkz0yR+AIqxwiRgaFDCuRo+DhdtpYxQbK/ZnTdYfyB
/Ky3JetbbcMf6iKKxGDDMK7jpm7LtE6Yg/7O4lPGROEq9ep0EwipnMwZ72mXPJs5epNX5dECscbD
spRiXZDY9qecdLbH/AwNv2kGkH/m2NpPY/r6XX0PN19zVV8g//EngogHWuRpPlOAuzz5fijFeChB
bduTr3isDlEv7yPXY3eAQSvjfF1xgt5p+y1jinpfT3q1VPLsYOSts/UUoRi5aYcLW7VGgKD5Udpe
1tl6H6OkTIXQsa2uy4/Pt0hmKVZITECnoq/c2H7vSZ+aSV2NIJg1u5I7uvFVJut3FaLOX2tI2rUP
7U+zao/TD2oGa3IoZ3xX4syGqMBnYTTeJ6rw2lELn8aw+prQx7AbUVtD9zBM8r/5ejd2q2fdekGC
GWQfoEubr6opTBV6YUHMz0tLc9PmNxTx/FhBo7YWZzjxuvvs8Y/GiFNqMLMDd2LwqzmecyaVbOJN
Ni6r8DRxQ/ZClO0yd6O3ouuWIG7q6vOFKi6ir6k9eR1hAAlYQhaHH59bXrsHm8nKWLwzBIl8yOKk
0nzyAXpc1ietI36igT6Qw4HkDNdMkjVIt6yA6ycL+h2bU181jqbckx8jOE25FHr1Fy9SZEpDSZnH
yUzUlAmL6XDgvrrDtJlk7QFwaWYGh1Q0EzkCOErdZiMzuy/qi3b+Rj9+Q5Iu316MWo4NIR91xP/1
DCqb97rhIpXah8z2Vunj1pZEuq+vNcZ5I8EkwqlXZwErqb3ZT7hdjZlZOclN2ioRF+ZV0fohyW2/
RXUSRRksjrsSsa7S8krCqRijY6iTdF6dL/doGORxpvz6goUfGsi6YHMET/9Gc0r4z4RJEgJgYED3
YMB36m/KPMdcgCinxGsbIvi9fT1gQghJVT5SD0ncnevPI3wUsfEfJE4Iptlj4T6iDhhQk/luG+PF
zY8D+iGBD5GRYXd34vaniCi77KgE+jzRq+F4v8tGzszOK/KzE0A9iKQGXczErzqqjAsS6Qb8U7Hj
LjmNDxfuV6BI1S/8s4vtJi7GcRObofUpjs1Sl5+EVzJyePCr+54AKDYrh77X7R5RNO/X7AzUiVHe
9dzp4TfyrLEANw7Rqxo77IrmGdvsVCoP98A6RhXIVqHec1BKp1AsH1ItcskZ1DX5LbkwJ8nxTO0E
xawjNSDatgp+heIoFmTsE3hu9JTBDIW+En8/kqAwGT+gycg5lgqn/Exq0P9yx44AIwluy6BPKbrH
L8qSD3YFITN+QRDKnEfzRIMAM59OKlZZUhe0rPhy0G33NyOWcqOj/K+Mzs/aCNqmePKGZdX613Uz
nl3gZAr/l4gIXh2R4mNamqhGa6xDVJwEk3Rf5971zaAutRz0mBABMz1nCSTesG5n1qmQwN9EcO3c
ztDAZOPKdSuNzuFdBl7/DFjhE1LVX3OpXQ+5gI4nkVruELUduQ80XklFaGAp6H066uMPJU3T+j7b
uTHwN9gUyGlY49y4lpDjGCdqtpeY4Vdoozmx7wiimsIffMnSpbh6BMzpQ+xmHUyDD9R3wYKC5ZIw
FDffjpKQi7SsCvymUNCDEncoDcfFMFaFd/FREad1q9XlZBCYLbkISL5EYLhD0wJ6vBMuOwSeSQ65
ssDymRP67lwRttKLmbXXXsOH0k7u3PVfIFdKVt7VSQ6+TLZAtwrtNHwSmlX2Z3AMV+8vnadfKN8g
SNciHWy9N+2Em9aVx7CXJII3Rg4ZLR0xbxw+lEv1fO4+aE5fgaSRl6Fz6iT9q5rgtnk6RotmOxCr
7NFn6gf9w1bTL4hrrmi1jziqqo27jtKtd3NXcE5mlrzrjXJwC3yHk667IxDY3IlM3iGIQoP4rUA/
Ramb1jonOPOq8bV/aGf8hgvF4JLfOULNoBrSmQM3AMJbCcFMeDPyzS8bWdrxIBz7sk91y+DJFj//
Rdl73O2QsyyL1yqCxxRhSQ6vo2M34wKFVhsUHS9At7Gt1+AnVEuQV2+mdydGwR6ao5e6XG6pUsWj
3+2b3ufW63qT/n74oXMZN2Rm3RlTmOupUXuf0rGONO2qDxKA79PcItObbIOKf+yFc0pFB9QBBxi3
IpilLH5Ntobjz/nO3MyUAed3Ez4rf5f5c6MJNLvLsTSL8b7kQSfX6igx9Uijt/XHUaBatD7OGy/w
fAFZAeipt9wxd6aMFmVPEnjdFStSR8u23vhxiwm7USkIo6G5/VC1WNxt0K2pR6XMMTh2xUgsSPAa
OD3BzsPdceFap+6UiBcF6o3C0wsId29rlxTXct01s27iJskKbuIVSpcDSDImpyOWwjQmN1Jcvg9H
eOoTkY3PS/KR2vAEJxiWW8SZDo6clhZ5BJOp/ci3lcFLkgVDnR69U/xxEQkID4UgA/x26Ufgrhcz
BEt4juhxhWzRFd/IaAgV0FM59G/WrkhNexl6K1GQ63qpO5ohG7dHemXHGxzJwmZbCCSqEH4gVBlZ
5pEwq6FUFcX5TVsm1q85GtMCFpOWFYuJgmHWCAhxlwzDr9YnH3GQTUwDen7/nzZ56oOK6sAzdj62
7wq+9euu9xG25qnNlNiW3bNuFbX4Tky/D48PTwPspsAu4+tTleZj/tnp0VHreu7cPnvTKqazh9l3
8p7an0cXWupr4DUj5fAfh8fa02EFJoMhrO9wo1rg1EVzONfi2s7I6mkILvOnDGpTQ6d/6L77stBu
aMHJAZMVpYwFNkH27fBHRq0iNL2nzf0/8vCOLUHl4N1eRhBdf1A/tblYbI97UCDdjtge/vVEsg9o
gJShjl4ENk7Ofw7Gc9HVXlRKAuEARjnEKP4p68BOYUFs3P4j9qP/Vce8WTL+eRxKcBqcVgb3a7Az
w/382agagEgrEKXGEBm/ClMzPxqY3ZRfBl1OBlcftgG0oiVhHd9NcjfCRgkNuW16GjGgJ3tLpNlf
iZhtmeEvwCdwbbDaKDsQp5k9e/fAeSQVHd+eCNR3T0hDe3+hBck+3YaPAYJQ/CK2RJ2A8FMhFrCx
Jvd2DZii50CyJqugOEKHLq73+wXB23wcEr/4LyQbMCQtDtU0pbRepdEcDb6HUTS5thxCyIeEG3RK
js35fQMRMno4xjJQ8e1/ppvxHQfsU1oCTqdLU9KG8ECfPfoxaKEfatTbwpHcWc+BCrbOuzP2qHLI
FCgYc3DSki/KA8Qw90+TFkfT2KtZh2gEs4DTVEmz9aKO0pfCiVYy3joHEp49jupyBzqQzpvlOiQC
enYtDkvxwKl2RXriSBGsULoGQK+Xpa1su+e6fP9EuZTfVQp+XSu4bAuGXBps2HdvAGiKaDnwSSIj
+6/Mng5bcJNsGW7Su7x5TJrdfyE6/j2Rj5ASA6ebZlyO/9mO6KgZD3W0AnSWUz+q7VhMJSN4c7WR
72Jw3dYtBIW4GAo7GCcxa2kTIZgoyVBe7FdSUA4gHN/557H1b1pdXL+WqDD1mGwqfuE1xWmu58np
tZl1SmSqFOZGRvvkmeZqc9VTM+EdcDecDQBJ42jaNGy3Rqf9Plw5CkBkCEYac6tHC0HrI0KPNgrm
TnAp92rCd4K0VjSjWiLXvbWkAToK9MqkcbV55Ec1bE/ouIfEk5PvE0XvcFzA6kDHvQJrYRZRKzYr
dA2xPcJVIDKL38hF5HNa2QZJdZ02aIjTusI1tq+n8WzMdqQbPOcAnT5uCZk3oN+SMhooLAkk3Gj/
Aho2NlqKBb4wrKm1NRTHcuCRPDxmUpaoHP5U6pIn2QoIi2une9AotmA6mqZFYEuxtLOaq4Q6ONjg
zVN7UsrMnLqQYWOv5A4+8LLku9Mm5VcuG7UiDcqqG4M0syml302IVW7Q7P1GUU5cLvAL7Cay3K8G
qotR6zDm/dE5TaBzqY4vOd4X78a2+I6pcYVbamdgw7sNH+vzgVs6xlTunYVCU1BwdzAKHwS8k1bu
7DqDglIRN1maMXH7DEoUnR3o3TTJiYwhZUOIfMJdo5lnAZeI0RUIUBXpjTcqcQ/l7jBa552Jc5PF
5hd0gjyJUeoJsbF9ZYac9hC4spNl4dHb9jITJqOS0moxk6GkexhH7HweAvz9d/vM0Xgzz1/GAkS0
Qka9xLsdKh74HjS+SqRUsIMtUJ0OeAkpb4Cs4hi7fFn95DzlAez8HuSrBxViS3xljeCq2vq/2t4G
887jd5xOQfRhaY8m8JvPojcRzcSdmb0xj+8L/uYyVeja/+N6cgUmYO7jqqnTn/VKGOYks+/hx2a+
pT9p/4AXF1PZ3HlSLV8I+Utj4cZMV+/rYmdyhP1rh1Ax0ONtNKx17JMw6FatvV//53gvDcCM5mbH
iLzx5bNtD6eRuCrDjXeskRl/UTZKn/WagOiCAeGWHX4c2YQJ/m20F8A/qnnQVyUGijMArJCeSytI
sjMzO5Q+Fk5A1NHJKoOpSYuy+nJhJ25iQEGUNKAz1ZLNgnp35/+MCmrrNl28yHabWNVa4IcPxh2P
9RfCo2ryd4XK2U74CNxbFRUUEdSjOu7nNlluN970MCLmrHwMQbVj2OmhkBwrn8m7OYZZiaVgjcFt
o7goA4Pf7bmnU7x06GjBCNdixrDJ0s1X2zguM0vvRB/LiINbnjfvDeM1FLmVtTYJqPgtlliRJLVX
gnuqrJJ4dxxhLnCnq8zGNuthachqoCcnmkhB+cHtu2c35dG07UyBL/nv1LMNX5uY9UG4gvEvKGzt
IKoxD+0R5iFxNdusEmj0QMN1ScDICzE8iJ1Cs5wTk95levC5hXpv3is7sxx6lIic5ondL8IxZF1A
DFB/neIW6ze+XU+IGLl30m7kdq0Sa8ShX5+BiKJ1tynDFkLLcHOjNLhDrpZNPY+PyPaSkimbZf/K
2rjhqo30c7i8p+KkZSYmmJnrej/uOmOZwVHUZo9Xjd/AHDoKRVYiRFreEatRWw5C/s2RiypJeVb7
vt9pnHfSVfhUYf+A90pkUF4fOjf/oW4ZJ+L2hCkXm4CiahTrO5p18BF7OeUIvWv+i3KuNfHvDDA6
EhiYSuePJN6dalTdZFJNByBwSxXMfGOGv7vpj0K48Y/XUZiQKIEWO1UpbolgRL5hjgETfm9qf0Ym
usWUutn0QLnC5hFjSWLHJdEnlbh4t1xjQl7E03iuclRJ61PMJNXF6fSi6Ov2y1xbwRGiKshKfnZv
31/YsObVRK2WQZe/GHa0cIro7vKM9cHep5Eb5vKUdKl+gglNAI01/rIbU1mT3hEVLIuS3bOhUStX
KdydjxsAcxEUy6F+tld0FMWKNJ2b+NoeMKo0xgWSuUaGmz6r4mdM5/zCkI5emy07k0t3719K4mkh
0QnmiepfI5HoCRKla3bD7oDctRGYh+LEKsZMjJapnUbHo/jqLb3W8FebyJYackAFiWMi3Q7xRwcR
z7syY8vmu0arAgn2oQI0wLesewx/1JXDlo2B3YHOS3fOO8cKEbx4G8ag92xjr+EQ2smJNE3Gv+9U
vBVGKBnidGXR8VwpqG2xCBDXXB7SSBeyoFvLFcopRDULn4/oT4oz0u2JCT3lijARHERGQHJM0Jbu
n2fpVR6QrKWLCWEENd4aF+8XFF/zyMjTzTNCYqDBQUCDMjdqLgg/AVUB52l5HCkMt20yYQBsk4AW
ifMSs8mVPpOgP61Xgqg3Z5TlCWvTOykTNE3hQPXaxT0d4LEfnrGTPiUvW/5Q+viBGt/NWVNNsKJW
tYPjIm2XnyN6ijSeujtFDtXeyQWmK5Yw3OAr3pHE8TpSUwWYqo0MR+jObZaJn88FfsP2Kyhc25dN
zbba2rfKUO0kUs9XzXwQOdE40f9OTQqHRdlfFVNQCnLGQfFhZFonheL4TiGYI+v8aXLnobh+Ib5c
sYLBsKyH/qOyfeBSDfubyW0BoOUiuHpIe9sZV9YlagQdmbhNCkJNTZ7ef0os2a9rbO03EJRxQZiF
0YHPJYUMKIZxtNvUmlqLY0YQgZ+6PsLgCGDXghisy/Pju1HQBSAD7bzd2yn3MM+JY1oRU1n+cCEo
SjNl+oFKdJbYoRYgbAvPTYK5ysdKA7IoTPrJSWFbr6K5KbpV47XXBILQ9/1IA3dQyvABOEdKmYlK
g5IQQ+DIdsuzb7LCs+AaE9eC1aI21bQB6lEeTYgguyt6lT/es1Xr7JDMvtOrbce8GGXv3djcl8V5
byKpvTfdD5kJ3+KdHmSMyEIBOJ29ox4ULUu4tc2Kb6SpIJBRJu+2D8aa3xR9XdvGCmO45lHLETc+
pDjsIpNlt7ZCCpNPgLJbkR8c6DubFhFrPWyZM3cV3grslODIROgsD+M/+g42PMuQ5/YlyCMJFvXh
bWOQUay/5Fdx1WbzrVZMtaqK42YR5gNEhcyG7dc2/5hFCfHMWd+2ZqhOSL6BxPvr8ERCLGvgY245
uNH874Qe/EeEgBhWq3biOP+irapAMsytk31OgFCtlceikX29q3nS+lvyflkLpMUOpuSbiaDh/bNv
sApX2mWTApad8E/pkSpaUoMbwC6xF1Brvdbbz0LGmrtp45gUIESIBqgjkdVNPo3DhWXubHxOflnk
gp8eL48BzNUxUnO05SCUiPxJqsXYh6O4giQ/5dUIMjE0o378qoGI/dMBpGMyI/2vKGi4IoG8i9Lp
LcdPUGPpZmWg/9RgP4HUX8haEyQIechDOQJpTYMA0zHvPlncKo0xSc52tSERPYK8Ao8fnjVpMdJQ
8rm8+RTuwk1edVNLsxfCZCaKADeKumGoJodnQmYpVbRoG7R+uebFBvZNAr+vcmux6i53j/mRRqF2
xp2us35wbf7P4fhsXcRIdYImr6nSwhaDdClDPDiNkMZ2s1zEYXNtmiNF9aXyvuqWDPhwOEZkb9Pf
krlOnkPCVlaGqWzz5VMb7//Y3KWN5z0YgVW2wpOnl+diK3nvwa76RmgAkOFPGoRt7jOEWJffbNNC
YTtxnyKOY0OnhLZJcIRZObKHUj+7V941h1nC1OoMndrgb/TONqZv890dECgrkxdD1Gq5LnhkcYt1
8DMXc8UIpM6QFRhZKVzYFQfCZa7XMxrtzxD0qZ75MI2mQyaA9svYJv+nSZGeuouAQmCIDBnqGqjR
nEQsLYoO24y0LnaKICkrqq21oUQSONn5jbyqI7xlayLytKWPYylb0kTN43sWPuckAkaoSDTVO3WS
hpgXaJkNSxt/UcQYIl9nuSLfVB4qdTN4RnDuhtLPglHuLIKrIS7lCQj3EHCMi7XMrPlfE+5e2Hqe
0jV3hWSQMhpOTFOWB6sZJumEfpmr7TAmkbj6dyXljQrKN/R1k5/RyIX0pc12syeJ4pZQd5JlcHVk
+j9W8knS4nlZiBrG82JkZX8KGRPS95G615IXDGs4/OGCfMjNkDx0FAe4CcdfuuP8R/cBk7Sb9wdY
TVmuFzT7g5WNpR+XNhBBtvHTx3nRPHey7iVtylRniiaWtY7WkBNNsOsk5nACXmA4JQpBvW4Onf8T
ioQT+rCnK3ObDsOn1pcR5TKlbwxP4i0MTKMMAALl/l5uaB/dbaKWHZzS/Yee5BzwgA+1nxy1Ipjv
a4eA9GBAgiYS4FXczq2sgTIlyfydf9lB1rf4gZI7ynhEsVK831W3H11/AywJM9xjk04VbqTQONps
4n4pYCIrNtONDNrgIuhcpEh6nymMpvqSZXUR/cNyuZWes4dHgp6MfETZS9C0nYmOv+rgmBydLas6
08JCCFO0kxMxQoPMW5RqoGmCvl236LYc5GHo6CUSlQVEHde5yUVwPR70DH+DGh2mhi8Ife7cJfEv
FOQH8f1toGgBZ3hb9ZHPhlqsySL7mchFHbOZbYHznqZbtko/CkTtfcamv7TQNYZn1QvfmJmTIYxw
4OKLK2dTWTLVFXqwnXunbv8i/BC9qY7yM5LHPuRBqxNEXQqSLVy0ecg5BbRBIcek+cleFSdPxYFz
bbDtA+hi4vEOBc086UBYkHqfNOmkDqQAlbs1oUugdBnnj24KLuBtvSo4XhUua4UVoUoEAGjKpgyl
UIAcoKLewmVKfdLOzhGbi5YP30M5xYNn29rIE3AAwj05F82CD0+VfjcHNtrEHOFtyoqhRhxGIcJ0
N+jIwu5YPHFb0LrP+vaWgO35rNq793Bpml/+g+wPdHW3LAZrd7EW8sz2pvaNc/k8E5BDtwgvP0uK
7y1ILJuKfpHaKbEOoY0SapMAxJ9ZslsI1fGAA0TXacDacztOX8Oy82mUe5EgAXqP1ytw58Za83+K
lbhDC+J6+wFOUpo4n9SHOCrHNuMrbiOQ9x++rFfkywFER0dlB8TjYyaNg1vxzBwwa34QoXdO5/kZ
zVRFxJMTKFbuZuTQLtRvJ2IyrH4p4Z3geZupkRsoClSOGlJh45kDcQVDKPFqm/8S/mSS0jq1Aw6e
aEAYVV9SL/HdofpmUOnoGNS8Mtp1Ez1V4qbt5UeN/d03ZdPAsbTk7mYYvaInGuP2YC829TELuxj+
dDS5xkztrs8QnsCSU9fCd02pk2oX4nSuIA7Ifkv9wbnU0lcDYv7SAPd9GRQu/iAdhkQdnBI3CGAq
iut2hheUxXoW0zSI2WTuCA3+nU0aLOwJUSZ3bnhSiNjXDT7j1U3hNwRFT8AqVECfUPr00h6lKE1I
9QeXwyKipuNWiYB2ydHiiw4ftYKxQQk1yA7Hi1Ll/XltYpJQYCj5TeB6ybTDMZHaVEQwa1WPmyeY
yRqyeStIiWsjSFK9iSkGxm6yNgahBpk4cY5Z6X2U10Fcc11Cewl2UoM6eyP7rInhPrbPQzasCq4E
yEa6cc177TielkwYOsxvRpbeveDyADYRJCZ+yNmUfsplEzrsuYRyPso9XpqBBOYvlN+cqrqkhaI3
XbAovQWEFmU89+DUQas3Qk/NlADr4P2nE4t386HFlMOnflbsl2j8uUxPliwySegnGwDKjcUmyMtM
4ZIlptNdUsWedoBB3h7BqIGfj2/7MQDz/KhAixdct1TropSDe7hw0Jz7wbhniBYOV7KiC17pW03q
SXAXXtI4rJSXdeeGHptA0qvD41wN0SlxTNp733aFNQTceMTFdvnuufN7uur89eyqhOE7WKqC5j7D
xwE0rw/oCZjCAMgxcAlQqa3HniHhbwLiXfTKvlIdaHXQZ1WLaoyAonwYVO/Wi/uAHeCFuo+/PrzW
i7rlX3tKK3dfi/lxUezCjRJZZfLfxLs5O1aIZk/iswl6oPuxwCF5pw9AkHPF8gxz13U3px1oameB
OU6C4VAHCVSGPFrHv/K+P+6p1te5VxuXSLy8PUghzR/sb7yMPPMFo1U8PHR69pe5UW/ObcIELn5X
l5TDdaZCCXs8v9whI1z8AGMp/OFHylBELzJoBPsjQHnngdbqTL+uANqwpLFlqIVwmPGu8a6gWIXT
IIAr/xwglWwzAGdzL1OrBCjiG5ny+TyUO43aRnLJwznQZqbMVqMGPNUjVO+fuyADYB71EryCu/DH
sMSYNakUgs96rzQuvm1S9xOT26ImE9VV4M2jixzRORvVFwHMostgKviuDuk0SccK4zLNIkSCHXbb
4vZUITR1THlm2sM13X3u65YWJuUT6deulJbSDIQjuAK/yPLah804n1iu7m24C74qoT3c3DXBSoc9
HTnoyFyUzWDdUu/uqHzxdsOAB0VO/N60r/SNvXBzQ9Z6ZbkFW7VWbcPfWqSLaZVKRRFuUs6Mjk5F
8ZnSIcqCs5bvzSnmM1dxunOh1CfWWJRpM8pxAUHK02Zvf7Dp78vq7KKzeK6D2psgdOIyiA42Nj+2
ZdeexANXr92yMNIULXk5lZ7k33p6cW2hx2RDFLJgArFcteCMwk738razA8Wu86shlsHQFoZ/87oF
ghMQaqXq6qE3XFlM6GB2ujxzHN61ZwKx1Go/LLXo3Q+N+w7Zu5TbxMis+MQRRmsFnpzvQqI4guOU
cshR3xoFro+wnCJjb1tz6YC1OEFl+GfMoqmOfGGC/8lxbXwdRooS21v0lQUuu1FOwMwqsfPFSDko
JblJwoDvLUA5KKRhFQ7Q1kI4aCD6XMNbPCxCuovHXjtgZ8opERm6wsuHd7GeDJLxG/pG1nS0pCc6
fEvkclMivsCpohTIr/btF5QNRb0sHiolnB9W/QSsjAhVKQt5USFTXBMtXhmfvo7JzyjRoQY3CSUj
Shs47o8OqaaQv9EUa9EO1nfyJ7nm9mwhUmxzu2VLQS1vUuN2ayJn8gXNZjKb1Ztm1PNxdHWny36R
cFjAGA8qIoAp4l1NfHamVwV7Wb4DwPRDYpR5v1atLfwaqDWo2wOtHGF0iWIwbuqx1XuMyi829b7w
anpCTN6PKCdERu63DKQTiVRPAwJ3evcpjyCa5lPZiB/Z74gsmLH9EO/C59TiBZJ2t5h4wxyxILpG
js/yqkI6FB5uWUyKeGg5uT8IhN3iixVmQedrphlupYxcTQBcQ0VxLFPiVOAjgT6orVF6nr4NFsAI
zG5SH6CKxOZ+cSj10oU1MgQkPKep0H+VS2FRGVsePdYCvl3CLuj6Hu5twMKF0MBjK/hAabxhm/Jp
lqH4dsq/fkPyLdzSDB0me0LdsrWnECStfA570rUtMyPAeqJYCpJD7C95yvOcs1hbz8GF0J8fb/0z
YWNl5UVnyesCfzksxKLb5ewvRMfjeAl4nMIWEmOFCZFzEIHQh2Br6CeLY2Yaf2v0qetyIE0PjWbi
J/LOgzui1zl5ie3sp08IDahyaKHCdJOJo2RnCCEo1W4qWEdSF3Usxrpc8V5CQGTJ9ppDzeGORJew
NkK0mEBagoK3C9267onpeEX3b4oE73oUzl66nccpwFxRP0u0nqQPw6x1pGbcQbCLYEhpTYUanG7e
07iuBVRCXrJHPbpsi7/NLlyZ+yIUld6Agjrzi6GN4htA0j2ql9Yxntuo9hBdrwzweuHE0U9DALXB
dQvBa5nOfP+SnhdM0Xo6xVePJUeQQj+seRQAiVrkUHxNoFUyip7s61cu71Kx0X5vPV9Lx9cbkw/j
15lB3ZQYvI6VsfNI07BeqAa5ut0iCELNCBSwpM+cXAy2RmOTyL7H2o/XqpClzDcwYSJD25AQVw8S
YX/Ybx3GJFFv0NukCg2dIO3VFnc50Fa7jDakzDZc03sga2qcy3P2hu/UsPanjpQqzRAcO9Y3+vju
f/UyiOb2QW/sthoWCfZs/6x3YVpHMZU0aa9oJL3D6idHUeqq/Rt5J87ejH8wzPkf+fTT4TJmWonA
rbSmuwazFqw1wyBbLLknlH8wgpIS2bIToxtQifchv2mW26aOZiga5RTMHn+jASQJ64IH0J67YPS0
3EEjwqzw5/4WvS58X2hJJcZm37Tsja56CPZKdYXmZUClnYh/69adNM+NZYSKJGRmor5RlQqP7dzF
awKtsjTv3Y5bCaElpcLKfrPVrEIyFkIeryyhrsHF5RVdh1ac7th6chK/GJHagegEmmWvqsWkhbrF
uSG7LwqKb2RodAgMD7P15jaJh3hXLAdg3kEBDTG7Jj9/6KrYFLBxf1kxDQxZBMuizuunLfaDs4gM
bvH0PBxH/4LRocCyc7WxZ+Y36rgCATR4XxxOPV3btww4s9tVa9keaMCaGzx0wsZ+FbwWHLtkhugJ
vul+aIz1JRBmk2TGB97lRsJPtdJA9JGQqkSd0MA9rdhqpT7spWy/Th7F2KEFeNGRsQN0ATt0MH0u
CA91gp6PlJge5kq5dgvbpoXRH9DdSfGgH+BYsIfBiKfCYUeZCRdIFZJedr+xuICHgQG99ntgnnqy
PFdQbXDV5Mx9QV9Ze8gEYk+lvULcR9Uuy41bRQnHPFx7/zPnxPb4iYeaMilJoEhT9SyCibEULBNb
M8qpHbc9SYOuxE7OmNPYJsVfy7WdzmGkvKVoE7YgSxlCBXpIlWAwfRvV3Snow/Gki+NlitLN230R
KjgzQmTmcDBAEjhO2S2jauNij4plYSkyqw1CrdgMktvji1hrxLE5kD+slDMZVwuYoI3MByV39N+d
YslG1ALIlW6H8VJqwBK65mVFN0AUNRa68KhoZF6K6b9zlkVncTsOmszDDTk3hIUHXe/RMHX8W4s3
7fz9aKM7oJYfRCvjPUKT89aJT/ngkt+LRCmKBDIEOEdvvElsHccD7fg5fy+i5/oHadIfloPzzg/R
pJKw4vf290rSgDfg6TYvFmi0HmYezTAeAdKS8AzTtkZxR4M9uBv6k4hIK5LAbYqR6QXVIlnGGfE/
u7lc3bgi8ASJGZeaI7TF1VRMaK4fgn+PgfUuB2pUMR52/2eUHSN5BI7dlyNc9rp/aNwPdDMJWSZd
FDnj1bYu5ANO+FArS7ZiyZ4aeiA2fKAH+vinQw/pAWBxVfXYEy6hw1BYezPdEXCwSlxmq4shPzz1
ajvUNEOu7TsPMOkRGn1HnWCfDooR0JlRqsu82TrnKcXmLJRxgw0wS1iXVT7L6l+NPJjGkJnKkGX/
K4tvXO+u39JY7hzNiyQ1ISCJ6xkq/peQRx15XDUijxsucK7gFYjHNElXHbMsoiysOjXpye616S9Y
IPkdzV2bXsEit1mVH0qG+K+9YhZkZmhoi2iDd6CKXv6BbF3o7LirZFMlnN1V21S/u7zy8ZWA8Yvo
9Q9oE31pUzlZc4oe47489QODyGW/56nhRo5n8Eluumk8PF7ITLwKs96mpg7U/aANiySONUkFbcQO
iiAa/iJpw8z1pWoCPeIcXGaUPdG2g97qu6/5qQBHL20qPXJK2eAmNMMUSuR6owLVaOzVIgMRWgGN
NqxWV5rmGCiwU7KsYj7MYxjKpOYZZ1iTjCTpj4y2A4hbUSsGhJlqZeghxEyQ4Uxa4jlq7DcWX5eX
BaAJGGd7MtaamdLiy3GakfaKWawXlWbWZlLoYU/0Yr9c8cegodoQg4SMHr12b2UB6ZOPzhz8Df+C
CC2OIqyxWF0uSOL6APZa2mHZit7ag9BMM9rUTLu6ptaaTXB7uWGxL7ztyr/iEindcnGwJqD8Iqn2
2TWPEbep9rMguQ1FUSulFBeK/Pmdd4T1Gk1IPrKASDOyZuLsOFZXx8r6QQ7Dl5UisfigsQewljnI
ActnMycZdr1/bs1rJCa/mTluG7YeVePAslQz/mXOASUvaf6nHZexbw1zgp1Cu65bn5uqtH3EvAV6
23kyGzo2+LgOrKN5TBxHky/OtmJJ1Uyzt77GLWGPyL4NQpCJ3qNs/lqH9XksoBqfoXuY+mFhRLF4
szPIsTCtHFMvkcdN4SFn7neZ2G1hu6lNB6Jse3neqobTpByc81awsUMjvQVW44mXY9B4CG3eU1A8
JS9mnKDil5hDkiQ0axIgvb9Zll9A4fzIWiamYPey7dHEMS81ETuuDAn0PRV9FtOe1VAph5nFLKrd
akRdlCRtWT8YzW6KT1XAdHbmwmqMeszdX5LvY1YhHhB3HqtuPcbnUZ/Q9LzRqOWfFYDMNEVpu3yd
sOR1LLCqIrEFMgd1XtJlKjDCA4H/L5FBJ0ggGJjiHcHiSpmvfC8rOMfe48p2cyPiar9I8A+ERDnN
j0eKYAuHkNzfO135V3aBbhaBXntTlVAYSBniCs6X5APyWTSNOIbG/m4aC5n6Xtc8M3hy7O4ha8DY
yrJkMow3lHPn+sGcHTpgVXMsFn1KOrgx+sGuwR00DrQ/RFgaTpa6LP/vHhM46E/56+UOUqpBezJl
e9jUpKgr4cqo/kv1AscrAy/7h5NTNPrqRwSiO4/SsK3KCo9V4DECXNsn8G8HtQEihuKv6zGacF5Q
a0CfpKcpJJf9IfuijSejZI8HLNw3kGOENM2v+DivKPwakQ/7567xsbiQ+VlNsw+lo8pjV6Ara+b7
h+6Iv56oIBaUqUY35sSM24KT/pRgOexJo6pnG7F6FkpvaBRKpdOWlH73X2EGfw7f3117D7axfqtN
SBz/urY6Sdp9hH+EeyLsSFqGqZUUf5SUqKP5pFAHe2kHEcZPl4bI02q+XbuvxQeCX2scoOmc+rsW
OlzxAuoRbbIH1z4VBi92Q+/QbQI3+hoe6TzHUI4ROs1lo/ufWvWpZLMNlzjWpp7IAvLuwohwHicT
qNDpUFTFSSKXHlDe5YRvQf2tR2SR41fNO5OJjtxstK2ijgeJ+NSjtz1pKhbA/F/e9IMswLJPp+fw
W7SsF6FuP5M6lXwnphnsQwQxbOUOEFow+Fj8139xaguR/wgTx1f0XN/RyidhP2J/ybEiPrN3lcrW
8F7ltoaJAqsQ621velu5hw5KCAsUEpk8eOX+h22bwYLtGAtSEaq0W+KokZWqRiCqT5zbwW+WxBr3
3M5O5XbxQfXYZG+90hZupc9AC0hIeRp/ayF7CSvtoiLLPeMVLkzsduLzPwHJOtsAkELWESPKNKeS
j3Za9R/+5OghNT3cMsAKXUUQlwEzEBReULysd1rCfVBNu+mf6KvaE6PbhM93wSVGWB6w1TTiDbzk
+lvxgWBGieyHiujEdtb9fRc5cX84MZjywQLD78weyBAKBr63v4Lyc7+V6nJzb7q6G+6TmJgkYHSP
783g1L8ugbh9mxeqZJb1pmSRRLzvbM9ib/lRVO59EAEk+5vSAnHguMqQft7KXdkjQD/UOtHyh741
BO3x2mn/E7oLXHvID48Zw1Ub57aRTqYC4sk0ycUyV9GQlho/Z8LTIrY90szPsMJAgbVvtjuspMw1
UKvOtSrFNKGdTs2p5NNfVnZ2xABJz0VkKBqrBeIV5sSdq35Iwsju/IkH5n1gUquJaaCmNjXFqVOx
9osbqRTqXcNvHKgyuC/BYW5msTLaoD4cuMAxWy/CVWi30j/dNmCL+883Pba3Z32GIClC0R84ho01
0VsHcJrSPeXiQ+W2pRjW2INPQWFBKpNIQG0JeQLdMFTrSLviMW4a+I0LZAnSrz/z9HfFTt/OYgZY
6hcp6IfUGiw6abJM3LVq2jVHGuyFz8lUjgTRK7lCDSKpRXpr0TcQcXN/H2m1JNkqB7oQHC54Hrhg
SNPaP325EqimeJjozuq/L3HXeRVxme7yTonesoPV9e9RU/+1xpKXJBX5mErUo8SaoAVSLEgifRcC
X7yJozu5NfwBN1pN9g1trVJtHSzKTvFMnAfvJufpdh/FV2dDXsYhHoGfYNGRpsV0KWYuGDo5cWpt
ZEOi3O4tB6mvNUD+FobeZtiab7fe/SLLXdNrJmTkC1DxK+FPwI6z5i5YOX/15I1IeWE3Jg82Fc6I
DhmfFPZh8fTq1e2RYTTT7SS4HwXHKA3OevAWByVW+WXVZnIVaevftTi/2sUmICpH3PraBGkYHJ1G
nAr1FtAShVR6j1w8j9D3rNKAq+fKQb4FxWH/CQsYJBBTJISDkiDiAVZ+F8KxIinG5xAXOdgfq/yb
XZiwgXTEvJmjHsorqAN4eAB6YIQ8+KECTf7hQ4pB5cJvWwpHSU4QfXzXSAF/wplfTe+gM50BR5ji
hTSZM8U09viEVfegKqmuLoeYHYA53+Gr+lSYGI1Cn/NMUEn7FKLOB3JPcCw0wdEB6j8k/YRroyCu
kspRiHoaCVYqRnE7FM2Ug4luN+pBJxOEGei1BcIWiJsxatDK72eH6zuETtA7b90pOiFJV1Qd1dFz
FXHIdYuQh5vx+nAigsBc46S0Me16/B9zEoDDc7tmZjRqmqaMjPVhZv1h4ZKmdoRMwvH+ENwQ7gNJ
IjvJmTVDs3Dyw9sQj0FMSYTrTvlMw9ZhtHWkfGgrPp1G9RAxjuJXeFb3YS/s5soktBZar3/aYT92
LC1DjVB+rtAptPlGnC9FoXsnYzrYG09w9c5QlCZwt/2aLXA0Vv38Re6xhFjN61ijaGzGtX1TTtYn
Nd0KZKWG4u38ACdJ/X7aKaW9pdFa3NtQa9f+MDw7DlAuzbDZ6Rw1BIrrhdh4/of6gIm1Y6AURd+6
XZ5stblyh8to6OiG4YW0mzxY5uK/wOPEFHLupCzID8VBvRrCg1S6ExrNyEgyIcoxNLiPQMzWrcbA
z01bQCVE4IGlEqo1QTKctngJYKt4ZCaZRTTKk66fACQGYkyal4rFe6sKsqnZhN4tsKuavmeSmxbc
uvEFB5XT/tn7AIyQA/0EMWG+Df9+qSWYdtEMR6uk8k5Eb3BMEmjsmdz8qxrWRJzMDiXEtTR414FI
qEa7oTNcLUMw1+Dejfp/yUknCkFpvjDsiz3bCJoPy7291OlbI5QCgJYLAbRNXXNpvp3bDXkH8c5x
fyylEGvW90N6Ng1Zfv4hGX+2S4A/ig6CklmN6hXRkfMRncY6J+FNv9Lx3M3zE++hG5Xljcdkg2Dv
h+4BAge03zElnqOlxz4YFdxUjFlAFlDyRPo9x4UXLjShMrkUiwrPb14wPgwb86iPwaYd3t9g7gTJ
CtOeG0kJW83pJtj0mCaQaAzBBssF/jjWYz7+T6CtuwbWh9bOyYXZyB2Svl6mRue+tgEIarIwflyL
M1Tf4Neygh+pdC5ScoukPJNgfxw46fE3q2OyzG/mWubFv/IAx7OoM4RRAKkt0KKN8H0u5stgAWVR
HzScrN64FOQAYFFN7LLAo6zoWNPlpwshYHnpwVCrvWb4VT3xkHiPdSzfGlPCzg/AU/1/mhRhxdtg
XoU4rYO/nDHt/+3OOklcshK1Febd960KW9GdJTMX2fLvbxZCnWVhu3ehpfxWhi1grOn9KIU82VMQ
91MuwNkGkSbwD7rCA5BzQcXuVzhPZySSVm+vdTAkoPxFeGk3aCxTmEAOPfy3iLNAxqNegA4PSnKt
lMB/Sfuwi8rioBJNyOCm6itHJrahUaCo9cH2l+uE/qkjhp0T8fX/CgS1V0M2s+d4kN2qEFvUc9Ss
EtVl6HUN4FlloJjJZWvNpr3c2CzSj0Zqaf/XL3GbcFXUfY9b+UWmpDVO7MHvObnXS1oMdRglQ7f/
lY5rHlzVRZE+KLmOB3mBIAGmidcI47tOdWvk6VxYkKI6y5o/jLSP/dmDmggodEF5YLNb4HAhrbrm
bch4rVVzCjTUzVNrLGdFTH+8ta689du3qj62DLtlqRTr8vEyzNsc0VAybJAP2jADX82A1v3N7urK
DaDAKwBzjTPZ1W0YbHNluBZCpKKiHTL2lqaq99x2dWG7TcKIKaZiWddEtIMX3NsAS3x9uufrq2L+
S1FFFL6e96/mX4PQrdJW/6gmRiwv1JFiTGE7pUAOwpzX0lTBTo3d9hHT+mQBa0Dn4uVeJawfCext
MvRVP/3AYyNPHvJVEArEYKa1pPmw+fA0AGViSmbSE0PYXeyi3gUbn4YxBBzJAVfxd5hjEdVDhyBM
OCrUGEuhl0UdFwB2UMZ19rsGY4x4lJfa0pY2AiBnzML4cHVLS3U8fOVvUZrwt3MrCHLNqYRm13L7
WkvXI+TBjEcQHMn6E3dBZXbPMXwQsOZAY0aq3/6zB53eEpmKzGETPntxzsKIGph/15Rbe9wKuoGj
4bb5Ao1Nvw19P3hwx2ixfbZpoJTEFvZ7xy37qBzk6UCsbfhxB1b1lN2hQMZP9iL7TzZUtPD1oN8E
KLo2OaaYILEGIqLiwKGJ6GRDEpODgkFQUK5B5S0NwKbGwDn35YkctcTIFK7cbCKDLdi1Fe/I09wV
qKsGKiVTwwKu/dYSYTBa84dfFWHM6b20rxc3NRakdKIsrc4o8Muz98kwNsp+v7tTr/+v2W4W69GM
GTiRfdiBiWosp0fVtAzb8rzhwPBo7O4RENLNt2dndMP39EYhhZigF/Ca9LyfsZooKBCcimq46ViI
JOUEDMfPpc3I8YUNPFyAQNAm3qFglAh7zGwJRwOStyuTDzl2Tiej8FMVX/Ijc9fJpQCdz2eTzQMK
GIE2/yOjwnJ72LxZteT+S7pjJvexzaw08EJBwdoFkYSxFolvgT+KIZUcKpg70wikh38v4jzXEXIN
dGNwCVOr2LlFTJ1UogPirtLprJxoyF1RhZ6nzypCY3kcgVqVQhkWnRq+0+iu/5sZjyRVAC3igy68
WuIVVw3sibN8zBkIonOeoeaX6RPjv/4DedesmikoOMeWyjZTeWiR478YvXUZG9G65tzI37Y7dGbq
sqXIatyxToIxdhDiQUOAZmZ+mu8qAc/OVq4Ik8k7EEVLWWqud01JPtyPkPsQQG/p5s5DIz4OlbBF
NhbjnU0Z7XKtbv5W5rHFC4a5xVvxAeDFqTL5RkM8MXN7/LbkISwRjw/hcL8d3J1KdXcdbns0kqKy
fIyjKOfewc+xFIXfGXce+6/WvsnFu97XDOE7dcKraVeHl80Oqbw3XR8SBEvsAMNCnmH+1+F4RgMT
aXaG7Lvnkf1QczW5hz04UE58cxlPHkd3LZB3ixD2aXTueuT2Y4tDL8+JKZY+1GQ2u1X+oMRPrjxw
Zg3ozP03GUIrTVBME8EXw4mc1L7C3iIrq7micvLnNCQ2OgxVb524w0B74xWrcc2VM5FJUSO9dQn8
FsXfsASz03ppMxemO8maOcgpMY981JYvhC56ET9yRLnBAmA0OqZyA0/dNJOd6ax2Y72sdQINL7as
CvqdVkYiaSFb3io+0ZouEtbBODSHb4S1MXwKvf5QbGEcIeQfc3yPzS7CPabGa4ee+g3k/3XrbgXe
UUxAh/NYZvcAC1UEUGxfgAkbjhBqsb5iRNBlY2lLibsntnbHF8PjpVQ5ys0Abhb3bV9my1Z+9Omt
DuwB1lunQTKTl7Dy8fHBiKOCVlapDkBTPCnfPo4JJsLqyT9OH3R++lxE8sjrwzPGyHo3m03XDm9n
5RI6iznpAzF5d1I5jjf18VNOLUR6oRDLHxEybyC2ExY1F4OkkaJwrpdMVRXvhE/sPIIInh3z3ckP
I+CJf6Ulmzgf3/I0eJlP74ORvHKxldlielwdYhh9+dIdcMs/LALsl01rWIxXrY2oAbcBN7YeqNJV
5ZnRnwqP0CRtbwY2IeNelXi8OoJZmhUZrXl3EFq98my34TVJJMQ++wdBsQkiBV3wKS7n69Dmnbkq
lou9gvEWrwabCjU/qFahEbSC28PUdHruBPa8eSDDboLJoLo69pH3gexAlwRlVznpXGKssWN7PYmW
9HVZMB5SrSZjW8dlfGEzIW35a8ldb7cD6JQW8hEi9Kcoqjqg0rrMcWg+XQskMqo9ZSwFMwYNyT9l
/+T9DRRdOfgtHtqQipVk7tuK2iaG96KkkT0Ty+daRKqhHGTPaynb8npuoOppylXjyekyBf4HH3d9
Yd1TC24gsdnDDYqtTm4wbo+0wPw2Npu4BAx4Xt1Ap6LhaNp82tLz4yczFZUo9+UP6aBvbzqu3Qp/
OrcZiaPbd+QMW+k4qFfElJ1uR9wIge5ZIItJp6AfBnPY/t37aBrdpduQOvMrht7L9QLQFQ36FziP
BjyKbtBag1RyPqxzrd2xPBcGBO3thnu1rP9zAYbQPzCGtCZljhHgOVjY72qhvVPviJaeGkB0EOS5
Wb5MVcaS6cenoLOWQm+8/SdlVE1Fw9wZeFmRu3raFJGqh9iQOuGcm60kHKqWa5dSBXZ96w0LwjTF
ecsouLnCDo+vYDgPzOfWdj6cZAIGCm4khRCIa3V1isWl7lHisQnAiIRZAakDMZnkW0ZlK8B0W94N
kKiibFV5dLTf6B7evRMOd7oRT/LtHUgJyY2n7f5xId3dLI7SCjyf+jVuL3DZPlIYdaHtsO08qAKH
otLkOEJpURkIbNaWLlN2fx8RMq2gx0OzASCD8+YJjkM+iHTsVjOs7rOSqI4XRdtZAfto0KgF3TNx
veqNi1YxJ3riUJv3WtebqZeNyXhVv/VoyVq6E7fBzeIzfpI/JFAfYnGLnert0l4VRQOYFuBIxQmv
jpDOhTbNj5N3l/5TMvE7OXehdMe4rVFXEEIL7BJbe/3nEYAzdIbtRd3O5MqxnXR9mv1TliJ6QkDX
4f4jwSLvqw7fntdBW+ayxX8YTTg0JoKH7zwiTfUBKfh72TeQ3XGd+92+t8BLjF4uX3/nOHTZj/kJ
YM49UvxDJD6z/1jX66l6CPo6EQT73bBmehmCh5lGjfgXbgIUfa5ct2JN6wzxaceFl0MNLRP3peaD
ZKmsie4qrH8EITYdEh85Y9EXhfRkHDrWd3vr9881TfhH6MjAFadCI4JsJGdfmLS40cI49fhJpsMz
+dD0eymGNoy2I8FySRnzXYs/0T/sPgt4ZLrzH/kcHc9lz6drjnlMNxmu3VmtbsxD9DOIXCkYgm0P
ygzwqfdLgDDiSo2xF/wdVmXCmLP1Myitcza5A8+jnNqvthqDe8glSFdeoPvcZCI07LxQYR7MCTAg
6N3c0vU992hmFlHaTQYIWHTYarozB1VigvxMfx9sAKV0WS4Mkk1SmEOfYdul9Ru61qtkGbxNXwKu
Jb51xKka/fXxyzjAjQs2/eujtwUNDPWDQN8ekF9mnyv5UYotbRwLr58SRLUv9VaNx4tZ3Zree5JD
UQQwR2MDVp1jIzi0wiQrTlJFTGShrAoOEKwhzROZcyAo9XhToOXI6jPAzans/o2Nc24zQtPa475W
51RWtUJlNJs1KjSy6/ZKBXezAbxdCjC1aM4rT+24WhY0wHVRQuzNsjfk3BMSpn6YVFrTmprQf4j4
yrgDS64fYnrnZzOeMnSPYIorFOT8lxyJOIoKkhVwSLOjguYPJWMRVMHHWzICOGcciRre0P2rROIT
NBIbpGVtwyS6UXDpnZqvnK+Rtzx+iX516utB5PgVEcRSwV2Buuz3wkuOdRHADQvjPq8IS7amkCjf
RHslGARWlhrGtwmUAyESmU0UuBnlDuE7zUEd0zCwHiaO0SN+hlNhsH12zYQtM9zTr+t2XUhQXeY4
9ZlIW79TH6rFZjsmXohOXZDzLHCwhv551HieTuNKO2Pv5MQ/D6QNnILdgMV7dji3TN6zLZN7pxR3
vHHVhVzjNNP1lbqyTHQr3M54umvUAg5SQtCPACZ0Mqf4USgtjkcv5GNuQoW3yW2Jzv2Bcyyti3hk
UaChje4WGnhmLlvDPS+8rRbHnY9IXOfNGC+G78qhp+JNv3yX9ooyqq5PszfdKPlmmEOfe6WOrosK
+sWJLpKVzmoUy8+TTfjJCLWVkEqxarL0wJUnksuaTpPrzocppRK66IjF5DW2p7hPb/Hufqq17XVC
3MzB/zLqMXpZl2qH7jsr1raqMlWzdseezctgOghrmGSsnR6MsML5n6S94A1oW+Ym1aP3c8+NPs7a
7bVGV5mNR04FTMXfvIlurNPXuq0YbdW5ii0CqUsSUVMbAGXXrsK3J3Rir8sokmM36s81kavKGCrd
lrur1p9u8YypfDXJL3y/Vz7NDsd7IHQN5pTuV05GdgpEB7Gc+TZuzcl932fimtWKE5+b+vra+lJj
up7wCeISm8lkqQkcLJt8wqq0hvFszyRt3K57trEC3dE9tNmuguG2HMLwB43pULql1h8uwZnbOo6m
IrZGz0GsQS/vcFdJNhUau6rpEvcKEiyAQaos/xRcj9LvyBEaY95Jf9N3aXVV88WyHbPfqIhiLEu0
tKQniJeVaSTp+VVM5SATfGC4DWtxPvS72AUWx59oCzU3/1Is9cM7A5m2eu6PkwjAO1mkFHQAci+l
ZWCOwhPow1VgAd+326lh9/SsxvmCYZzTS5Y4f6iimFgD9E+761JWGC3ikQdQVZVUMYvYBpapyVlC
3ALXEug6+R14+AAkFc9UyV+v/Xqoq0N6nGVfWBASDs/+hkLVImcZSERUH+njYvIg6MMs96RIwCoO
NSulcHAmJU/W0qtJWLSXpRsPUP0ecpVJ3g6saS6PhbzewwuOBiRX32wvxz3b3pzd00YD5k9gV2Ji
Ku2HN3/iV26DYcfe2sRBL7i3t8E/AfJxMsltTpvoC2zzJuCrv3aC4NV+8pMYNs3ClyHuloI2OBbO
qnxlu0uCgwYlE2bKw+hQ0ffLx5Epe/JlnyEfSGwb8EdYl+aNfrh3sab20qapyUiuKrJcW4cCg9i+
wi3+p5vpdlGWZu5yzd7aU2geaU86HPPHFqs60+Zq7A+cdV5vcBWUQ2gTIc/EHPGVkx5p5lc/9z59
dpFb11uSwi8V1UpejVyIHISCVi5Qnc/GWEft+MAVKAq1EllkiqS9MTamRWMrenmU41H0oVDrtbPo
EdJafVwqdrH6G0rhOl0Bb3ur8RU8VOHEkwQDUFcz7rl5KDDLvLx045bOFi9//XQmpFSlJWlGKHD8
uCmdr8oWbk3rgkvK+0BiEWPEOD99fKplD2IBAbR/70497mbEdyXBlyZXsDr4cjtAbH0HcKL2fwdc
o+VMw2mZ6qC2B8BGdedg34iMjBssT2S0a47sIGGxfm/EBaiMrPrsk6WWFJQeeg2a8oGpjrZgKUSm
XwKGeCklxDxy30gdTz5N9a6r2Sk8CIVV/8IP30MMt0uzAciCYLYgD6D0G77V/hg7SmR2dm1oRXWB
WOuiJXihqijrPQyt6VBr2xf8h8CqxLKPRgGxMnLtpGAOHXvulMvOJZ5XBkT3UQHblt1qcwOuSXie
9LdpRxZUIanBYjo7i/yl3N8RSEYHNobQ3e/uTDz4IeMeUHvdJx91gNpBEaHXytwr6l6li1sOpUS9
RQdSUHZi72LEu4kzhHcaODWVNl7Eyh0N0/1wd+IIRrPMkjsMHS36hZP4756AhjXGwHqr+LgOgrN7
VXYkS6s/0V2WBBvnfC8+w254Y+bGj3DhcFftNewa25+emkAUIfLEUQAIoElmggBMX8NRiUFLRFQK
Rm1TXK1/QGB1Dr7Ujk2nAqP9htAIOsV5vQfBeXJmhnzqsVmBVu3FRjyCRlymJp6OJnC/FlhVp6hM
BGe7PNBVmf2fEsDes8DIcHmN6R2I0nG3K7+5UzyIbm2XPPQBGNlnzg43GzAtD2jXLmajjlzvmHu2
YAsGXekBUxTaY6t8ECna3l81uNih0kqsgYyolY0Oe6EzZd5+CiK/BEZTU6pJ+ejmKj48Dc8GljOo
qqDTQD4Re1s7HL9Rxeq1cLpcwNg8mJy8VzoD1Rp/wnoSn3FOanlaR6ipHw4yF/AeiKOfeHlS8C5v
ETkh+ce3e0Qn1iHkDI4Bn7/ynKHuRuyo7N29fnQBUksBSIhQBed8jJfvbiwdSqcxK0Yn4nzBljna
PKxrewtTn5NH0zVl6x5Ib2sKDN9ZJhZMdNl/QC2ohGjBueIUS2o41WkIgRTEmN7eD96vwEp4PE8d
ROSy698/6vZm9DtDRvyqVpR8bgIHIpuZZ5TCizi2FKFprUinbF9gJYcwt+/Rvh9/NCVyk+ORCCFc
l/4I+haTDLxXOVle+U5C4bOHptHbUg36akvAccI1+2wW4P+O8ZColfB9/DaPbsY9ws6nne81I7+v
R+2P1isrQaghFDebHkabUC5MmiJ9NzduWyrFRnj0cAbRqj9mvy2lqctZc8bV4aoHa+gERJ4J3wG0
qLfy9DdXT65F0QmLVFP/9n3BBmt/IYVnsi3O4Q0IoEquFcFateXWE3U7fQ+lBuU3P216QW6AAQbx
CNG/EEda+ZoD4LnuB10YDBV8tZh2Bn7pPeB+bGXMChbjw9wVNxk+Zrv4Xo32RuKcXL+MwBukDIaX
PplSvwl15kDbvNR4zc92SNUPkXRm4XyqC6g0zZT7zUjCTcaqo8GJsNkwyEaEwS4osL/St7K8BiHu
DN2yh5Q6yQ4Sx6KXDnK72IuriyO9d8QJCPDeandqMdxMVoWg82RqJLbE9EghmJ9qf+N3MLtLsq/P
QJR4gfYBiLHjUL40e16a9mskWItwncLFto0iXtx/K2ItKGZktK/8sbRGZNiEbG5+W+7he6cyn1uQ
mAoSur51jz2AJMBzSxPjGgpw9c19kHSA6oNNGpZyrjt9qVL3L5soUYjhMVJPWxelnQI2PQUVDDK3
bCYoJaS16RQ1FjuhT1uvO1As0exjKF+HDyCmOlUBUM5D7wM+Jt8Ce3SavNqzDbKc8Qey0zvatx6+
uMYDIopjaEFB/T52/PYsTYwu0HnQUvZ3qVfikIhxNQ71t7bJjQ3/hPnblL9QkKK+NEKqjJWnkA1i
iZvdEkn9xwW7b+ygH1kGurvpwFj9JOsIk+HrZnFbllmwPPyaV11+ZuYIy9hQClMBvtxO1hBBUH/+
Th38JWeafDI0I5xK0rJr7MDP1Ey6KkcCTzKWowyofasUzwknpAwNuReF8zTSFQPsgRo6mweBDFf9
iD/5LBPGxul3RgVIwfQBeOceoY6gSjaqvgggaA6zjw0AUAK6UsjF0EQYbU/L2HS6q5123IliKO33
CVKksybmoj9yHawssKa65xrMH2IG3mS7s1TjNohJSDVBZDEbb0DmYmsIoTjeHPWB3brzxN+RP0Fy
TcnCsY9aoUE4fkDnKhLRNz9ach8tI7+P7m3uvte9YOUYh5hb7V9B4qvScAJbXzzI8r+eKNoDIkqV
yECE7KgIercMgmjDSFA4RSp8Wa0HlYu25/ZMdn73LR7zfArwm1QIVV7VOg9HtBCHgey56FLlr0DG
7b6Om/iwjdL50/tOcFrbmd4YJ4FfvF8eKCNnNhShnckAAocFBfCkN4lnwaOeZ49Inar4nQVgSx1v
bIKwTvNKoAJOxssVSYp40yGo3IntkanxH7YjC1zW+ZmjQFhpqomSxKWOYSGbRI2tjc5bYnJkARbp
Y3GkHzTMJyqMgEC4bF4qcdqCvHYmDzMCnp2iGd+mhMGxrIRZY0YQx/ctIY45mM55KllntXEOjYFQ
bIpQji0MXdMZ2m2xXqJd+C+i3/vjwBWs1L02zz/u80T2Rtzvr4p0id35kXfOvkH3M2QGk0LsI0HE
Ux7eJmWYCDBtmpC8Jg4xWP4CLfeatUurMSH8K0ExDAIFCskyWUt4K+x2fVChhr98xrMdDHaa4cdx
L+9M6kG0e+8QXs8CEtnZ46270dXPyx2PLkjrX4p0e/v7chPuoSU8wK2OiVIGFTNiwtT7YQhfMEsI
hltX8GxJsZTzLc3qc16mEGJKzIXXDssyk+UzjoMGxsxNVy4jqToW8eBWoluJNuCu/HZtVOhNjfNg
qOuqhVt4riP3ZvEdE6RxdiQMuUhNVxiCA/AZRV2dM8MbQzmY2muio4I51tAtrJzw3yu7zEtuy5aw
kkC0ebdkXbWImQlU7KFxjv+VkfQ1+KBFxNGHOYw7Ktq0GrLg5ULPtKGEL90SVifJkIs8B/JlraQk
e2BHzqAthfc9twuwmEXq0eDziMxHKHGPOcRWxAgeTqXF0L0VAC7D6ZG96zEANtj6zgHp/4VrY9Eg
kfktddwAsbrdTIMH6JeFmQUYRrUddOw/JeQTDEB6pHolTcIVaAdjr+zNCIMk9mXrtGafKuGF47RV
dWhZ+bvjjBcrn0Lnk0VMYei7hsPFJtbiEr+6gwGNofRtvk1tJqJ1pzG/bQJlptpOBY7otI0VoOvW
cXkPCzXkic8j+uEdHbjmrIYv+QLJH9kQpzL/FJBdzJFRAvfqxBQE6eA3Mpko8LWW+unoBoztfwTV
PS6DAtLZFh5hILgcfIegVVGlJmVpuQCpg+RvAZ1+E6kEGu9TiP2nz3FH+WIQPw9kNnrDdcfCwrHM
bw5YnJf10PqeWNEDdh7pAtRgRyn9gH79x3EQdlJxJLmrcsQaNtrK6JgpYUNz0ycZJt6xztWLxCVf
9ePEHTqxqwcLqBMPX1DSkZfAYuy2rmY/BtfLHLD+ZPULMcjnzGTL6mQLzqCwgatczoPczljlj5mD
JXsBMFl4AK+JZOfPoeThz21Qvlemq83aFhHI17rWN2/s2xzB61pkWoDPGUDyhNlKnnfQ2qcGZPlc
vqoIQ7YGeql5H590DsBFCGI1c0NbNXt8VCzJ1uUN6OoSh9igQuRAO/mNSxp/CUAIfy9t/JAel28j
OteS7P/CBYXs5ZYgd2T8iW4fzEbNV4x90/YQZMyOuCY/4P9yVuXNWTChR9iNESX5Tuo9tjlmwOCW
xoqazRbLTGoz9b0AdIdVwsMnn7IIAmWacffXYvLBSvrjg/hLaTjEh+rHD1WiLWnl35CcFt3I0ymq
Utop50/xajrA67N9u3xwtRojf9THps+W5oeWc0B2USDPAAlnsCy3sxBmWkXuJATMO3yHLND1/2Fq
RM8LxN+0zuBolXAJEVuQIts3Hg0gESP10CSAKxV3g9aiyhwr3EhtgBR/ePuJp3x4yfBQohAb1sde
mDGTL0WZ6tFurBKpxWmA159fQZdIv2uUNJhfTvqBl8+vIQ82Yvc4M6IPs9iDyoMi3ZLXLcKHVJk1
EGVDJrQBV/3f1ytAao0xynY4SxD7r9sYsLCHAQJqXxt1Mg/Wu80ANB9IqoAfB19BxCQ9bmegMKEg
QHAbqBgqzXWh2vIZOL8HqGc2mZTorawnGF6BDVUgftvJK0+/EXZgugn9NqGRC++fcPFU2CQH/R0m
Iu8KpVxzv3ZpGsfo6JfU0I+e34/B9I4syeeDtfxnamVvG/kEymWlwD/UlSMF+jcqG2HmJaEf3+GI
Y3p08DorduoG9Pq0OAk5KtApP41INseDabekWK37OsdXeRYMW1aRuPneoNCsykO2EuDuq/6pF1XN
7QyKHIUvYUW28794B/a+C3bZ/G4u3aomNR4j6BWTBIB0+Ay/9qJKpUOd3FP9ZNQRMGfVOGGV09uv
sAzrlfXpirUwfNNmzlqCaTwLAkf5eEfGUtLwIkVZWjkwKFuspRoV9UEGsfnGhouAOMaidgrl7ADC
OfKb63kh+s+TvQiEQ/5k5F/b7lFLQA9yzK+umFEywabuxoxZtNPnTsf5soQwVws3Ca1IQhTnklBf
qm0/ljvL+KxO+bifpuKQazlWo/+i3lUpZc6+RDR6wTBac2lCv0woa14p6AsMiVMdAHUkW5JYoDrS
90Ng6A/f1gMudWOHH2AHjEmaZ0SX2bHK1StF1zYqFsRh+T0W0ZHiym2eH5i0BNjKGUSqzugWGtHe
l8wsfrVUUJO0lMtfMWnkWxvr2xJ2sV+Uixo3i6lAk9+jv6BqILQcabr+qxj6/KWu4qzf7121AQDy
fu7Kf/5aKCGDoNkbOHbbinKol8kRt5LgrHO6Ms+DXfly9yVU0hmzHWAaVpQJrEQfU3O9Vewe6qUn
n5Fq7D5iAwfM16uyYD+mdtxARjTACKw6//qJG3OPDBVcE23i3P/QZurEW1xckSAaboVDY9T4+ZNA
4S2DANiOYicZKuxtnix46GhtxIaMuTn+nZy+ZMsbXbjOMcVnMFfHMD1oc3RI5NHO7NXOi0xK4oG9
U3KJuZ+sI0SX+i+F6GJqB8BYxJdxjoK3sIo/saumTDKfhfKSLez7oIHSlelf/q1+IILmDSMbqhZj
pONSRZWls+8CNJtcnTBuBwPrUcy+JLo9vNFsDMmuFQFaIWwdLQCxpJInkyKYj94vKfOLsXkO3Gev
aB5E7ujWx8AjIKbVI+HZq8a06MrfIwBdvpqn0d+QnCvyQ+O8UJ8s36/FYYTAgK/NYg2tlWexfVGO
XYJC/CR8khL3RYXFpOhOVxS55sDhgbIYcour2mxCFM7qexyrR/nRVoD3z2AzxcwBcxWzmYywH5/W
FlSWJzI3xn2CeQcJ5WAjG8LLQLmh39/Z1oVMi5uI2Y6r+N3wgp7SF2vw14CtZBTpuql/YeX+/4jp
W8EtJFzUhxDeiBX1wkJcF34wDFLB/E+vhItz1Fxb/AvGdTh10L4VB4+OdjtUe9a2KQYfKUZFRSUH
R0HqEtaQizWc9Qr+gQuSnjSDIBy2Olf8ZbsF9kW31fuE3/wk/p8hQF51CUyDS5lnIpwZ0JDyfUDP
+OJ86uxg0rUej1vrs5phqG0rVEtWJ3EgakoeTspR8AmS8D154+UrkB+R/0Ss6cWbu5vy63cnPe6Q
q6Jdmi2B+wZJgS6UosMtZl6aSpZEvOQTdixnLCdph3k/9yrPO7FRpvtDjYAoYgCa09B8Ebr0yU4+
L140QOyQxciZb/GJtbzgFLWqdXhhuzOFD5hSEZSxDJ4ocxvcdVF7MSRdA8QtRUqq54kwInAgpmDn
Wf2MBGgEOEZRrqn0tvXZajW9Q9V4Fv/nzgag4xvb9bj9OQ7FfjO3II32S/mb5amiB5v/2Og9lFiF
GPf5m5t1nte1cAz56Qt39XpOHgtZ4SoJlh9l7dcQHZAt9OA89kD0I6EII+dPGFJzDKPx7Iw+VhGj
DZvYms0R/3UQT7K7rv7G9K1D+LkGNRn2mBVuKRDmrr6kG3l0kIjeBaopRnBXmBt4Y+q16WuOi04g
ttgJTpMIbfEcdRnAusUrJB0p7OewWT7nBVCe0tfrEEKiHQCAHXrRsTWJBIUMWR4TQfEAxOJLzGM3
4nIvsm+TEtgTgKkovfwYDgzwr2bBUW2qVZJCnsjDzjHQWv5Fu/kBePYVU1+7+/4H2zeE6VVNJzzS
oYJmhjRFywGiOz/VEgqXic0sShEysvUtDaGy2A78x/WL7q/gVqD61Tl0w7kA5xO0kjzwRm3t4LNi
sh7sh/AnLoRASsqjP47thgcMSKOyTAuNVHwIwPK1XHdIXPm6fnJ8MCfnuq2uRCugaHGhtM+hUx35
Cn+riTl/+3iSpnV0NZ0EeZbsVI/hCMBJwyI4C5LJTup/tvP+zZb/DwEdDIOuPbUXRYCHbUgH0CH7
c0SRfHmTsiqHVL/YJRIA77bSrQwrbjxsljZAJfPJL5bqfZfp/LehnWOSxC0tuQCCOjAf/Y+3BDhB
045TqwDvbYz+pZ7BCCdEiDHEduftwgAitMMSoATfpcFpTwlsxeoMxwPkWgYMSTCrJNDLDSEN8pQS
navkI5uU6f1rWUUhchJX3T7gDZlJ/PLqZF55gVVxbWBhS2s73WO3+Ya3pzLPOvgc2jzp3cHYxz8j
5CuD4jI+zMCb5+irRwVgLrT8qu5MUKVH66Rn9m2dv4e5FQD0IqQ+7aNnyeHCCodneVroXifTqvGF
U/pwH3UIWBi9kPcmB2w3u57mXTbGf/pkm6/Rn3WG/4wv+g07U2VZgWzytR5bKpztt/qTbS/k/ZA/
VHuW2fAfFY4RkhgilxpavjGB6ZqmkrXrzmycQDjfqVtkGU8WGyHvGFh1LLaFLivrGVf2fskMaDgu
LHJxvZFPwnXBM48y7yOhqb1t757NCp40+zuaba5JvdlYlZH0hxafc4zRIW59rxltNeUJSeBhO4sQ
PNxckCatEUIJ+QTmT+cTZCWhSrWe2SmpKHkeMECOUpdjoa7msOMBPed4FxJxnYjEbEhR14FWcR+o
xW0+Q56m5dMXtf5eyMNJQYToU2RLxFO22BSlu67d6Cjz5AS/ONDTFj8rIj3iIpU1xzaXIX79jn6P
hfWNU4F8hPyFYlWb1ov0HVj9nC7y5FcrPvMw9VDBJ3tlymOVpfq6KwFg5Vn1NzU8BhVnngVPkVxO
icFPPlFAVPDDON/7Oh4oGJ9eHc3v7fI8tEXIm8Fbb0Puo7CcJG+P3Wr2/UD6TaQc+VDCfAGogcur
zizw/Q8UK+AmGW4AMmiP0XTXwxl8Yfo46M5QIlocVY+GolEku7PmynkL3Bn9BrZ8Awc9qgaHXfVr
nNSC1+AomDV6Vb/PANJEWf/mqCUpsLzQSj8srsjSB9zvVKRxS6HzrC330D3IsJGkum6gGB2NszYo
CmuFhH2FV2eo6QoB+VDHHJ9jNoPKs9vT6JGbVRuSmfTdjRxN2b+79yzN83+GjGJRVw57eGuhwsgh
DtA+G4Fp/t38EmTzcKqKu86rVdjLp+ykmZ+iqLsvmX64NiqcsNlwhcdnPZJhutdPDO1vsJlP6gEW
fIM22VevY+W9djqqyjOah/STguulu4XAxJVem/hZeUTCHkiVpPDOaE8notRB9T9qFQJ/wHw9veYq
3CPWxA8Ok7BgR48tTh3ArLkRZDXrIxp2ZwoWhTC14uh33BGKbuwtEaePCiaCMmKO4lU00m4g199i
LHFU7YchtiWMejVH9dzAWLMalZcF+yvIqww3xmnGefk7zesvS172wRrksNAgTWPl64oF2s3weK7B
ONwPKVqHx7hx+CzZFUkF2iuv2aTxC4a7Sx5gx+g8sh78RKhOdp4hmrJLzwPge3XNpMcAPUxLzHFw
yrR5YRqQUBRBK+4+Sjnfi5ol4YX768NJuuzy+gDiADnh2UoXBQWqoF+treLwKFahmLCzYFqgeo9B
XDC7O9MkNVSWY2W72JXQRXWN1dFl9Ck1v7usaVkZw6C4Jspk1qVnvHwRm0fLdcilS8WQmbNnz+bD
8tfEvfvL40U8lhcV4OhXInlnGe/SaJ1tcKd5sRw2cLDBGIo0E/0cQJh+QUYsPugl2HpRkijqf6/2
eikL8x/nyx1lpf/GTCM4XCtabONwGPST4qsbN6TOZWoImR9JtHWF2KVwFQMkiPQAk/QdnDJ0Cags
6xQ3IF6WudPnq5QYANtP0YrLqL9PQPsNFecIDmqp3uf4fSd029y86nA2hTUVPUa8+l6F+YYvC1r2
RTRB8BGyddy4i7TioVOv/mBe/BPQYNNigiMJkIeofbdheIX5kBr/aAw3doZnEX2I5hQJYqfh2+RZ
/x2wz43i/V6OGVXWvmmNv/bEszlug8KBk60TKa7BQnBj3E+wZZ/Sbx+yB+9s0AC7IomxIuq/3edr
Aq9cdsVxAdR3WPJaWw6ZdETgbAGcU7dk4LYqtgj1kj+LOmqWjkXa9PDFLZ8uv2wWuiwoujQYhJV3
XtjSn8GEmFTPPrUEjEPvj26riCE4BuhoCFFXmM4wAwv+t04/DaFz13e2dxNo7fOgwIb/gyzjN3rn
WVZtSPeBCBzVLvGs9Lxq0YQl/m6Nl/r5YEbLutAS0TpI7Ri6NbhQkRjIXmVvuh/ON2oohIqs10+t
myZD8BctNWbvijEZmhIsg4td05StH5RuoX6lpu+yideGSRM2JaKcvm7QyF/sdzg+QGL17Hl7aqqo
LhZJPOWMWsNHzYnSnhZLsMsAaPXVO5cqWmRqmnPLxkkcMHZHK7VRW0/ZZ+Mcf8LsmUqTf11ls4SX
H6szqD0HhriNSP/Qoxmw7jOuPp4sHSJmgium2JSgTgS8pECp3fAVtvCFZVjbkKwnlF1fB6Y5iF4H
OnkCGD+9bodli7mrrK02zXglLzZMUyUmyQ+SUq8pqza4ZV+1xrFssWEWL42ynk1ikgF9Qx6WtQYy
bMcTN/7EWyDi2Gq5+gL2iZ/HCpKz7NPjHEhDUapyMQAR4T0fldKZGrRv1P7hK/2z+INrqGDY65R+
d5R0qunGO5v2n3pYFN2OHVlcavlhuGGRQAUDvAZuZlkwC30zdU8xqpsa6Lv1aunaOO4eMhSA5vy3
KhniySOCSO09Me36jbi6LWC1FEpcFQOA+eVWzbXCVjJwMJmIyHN4i9USfW3gkFbLbDlREVYW8SwF
evP8h0TTt833dYiXS2Xf630F6j9vkdDMer3y9pjvQakXr2huocjTHJ3YfEQM9hIA5PgaaYpTS4nK
5GUGS9+VG6Kn1BGq7fAM5iDPBo1KtZyjZcglbChU88WmcWd9lP0EPXzaJfb1eL7T2iT3gtFxQ7dh
siDoRIqcWgXejYL7rcFDx6si/8QOobgKG51xpUW3NiuIq9GQi0v8bk0yP855cuSls/FEOefjqRWf
i4DeivTsrhtOp4Y3lqV0xfKI/1AGVud1YMPAHAxzxFLXfgtuwVZzh13THdNAJ4uQrfRentSDl7tH
TZG1c+2UjsEV/F3ezNYB4b9fpzHIKMYG/H7pU6blBRFEVhb+/3bqYohonEty7zVB3IYVbqQLHWpf
Dop5J8NulUAeeA1YUS8qjfR32mmE9BIXF5JXU53uj1oDhYgKfyDYltjKvpmB5K0qkWvN8hkgngRk
I49Fv+dyd3xSh29cP4o/bDfdbv4HIheZbfYGYyDBB3nxYD7yMqZvRPW0TQ8ekydLSSrMxP0D8Azr
FY9h7+4UxAQt3v046q3YZcAs34Et10KyCXNzeNdryy/DF3ugHPfHcW3fCGVCPYOnhS/T41L7Kn5f
1U/l4UHfJSc9SBDgXK2bwq2IhR1zoUO6GAZoWpIwWyFAlloSJHv95VE+Js+4Ds13+lXQjWSo4E2g
8UALWaTgFxL/4Ln/TQ48mPos59cJ29UQlgjGQBlZL8+tqUfCpeJ/2gmsn6egw5QutOIiIv7+apYJ
VHL/OvSsQ49yOoIDwnsuOWyBJIoamkfx1l2TmAkKaxiHTrEWPxbL14hTO2J4u8agqg0ySH+ujGXV
KfHJDyjMml/est/U/T7e3rwJ5OUS6EYl4Jh436/Eaa6QRsSOow+LbZzNTTgwKO2BOlHGl66OYIGh
+NC582BZhmh4p8ica5/RCQxD/J6nCyrkCJ57g0lzcmz6hQ62puXmYgHGnFB6UkZWzRQEyS0bsnQ9
Ov++Ap36OyLW9e46tJShF2zMfPe31IOEzhNeRLjZ9qaDHGgHDX0d4Zcnvh3tgY4VbtkjIq8tHKAZ
Hf7xYZrMI7YiF/oJ+M6tU8zFIFWgqBGhBRDOL9xyejnrxz6tIs6ne3KZHSSVY/R/8vFNdZ7G4VAM
f/dXl/q7qWOV7VkdJWOdRIZcqBAKLmPDZLop56AxcXP2mVNJaWUx1o/EGEC65y+qGx5fvbf7TBI0
TZ/37Z4qCC2qD4n0RJpKgIRtF2XY5wBlVcrARF9G1AE/abCS+QyxrmarJBC7lAUApObOqa0AJ7yg
ZotkW+yhUabJPkRv93ERtBE5Ci72m1K6IxB9WLDQhGI0hAP/YkbzBBYoKgvXU0czGM9ybm1J8olA
pqOnp2HDyOlWfMETwFSINOVZLtUtsv5/zThjydbbvGAYcakFTIU5GjJmqpTUltLciN6MZwQLeFaa
ploCYtI+25YDRhq5d0I2AF7y0axI2M1PazDHLYSnMRBZ+kmY2jWQD/iscYf1DnaADbXuLhsHt6dE
EBt3qCYHkZUTT4OWGnYD/g7qJQ3D6cHAz1XUMlt1Ic3GWGa5HCPfbMlVXAqNg8MEulk09bNVXvYd
mcvgJ3SzBAWGQozvUDGIpx055srmY5KySAtnh8vzJsd9JIE66TS6gb8FhB8V7unK2L7s4F3Keukc
vc8LpSkF9HhSZm3dlB8FW3Jjzt8/+FBoNQaUXmA6f13G5t+jfN2EYvDWsS8Z9kQV4kqJ+h+abro8
ROsspagvvBnJVgD8bfkQry+T1JUrVmsT3t+TkDF7eqIp8q9gZ1VxEJ2+lyVfnlTmAStRrOrqvNh2
2UV98M0JNZggHKjfJAv9mU2NQmMOzjMvQBWcBwSSuOZKrx3XBDBDjsTwlDsnIxvOEDm3wF+YXafZ
lX4aqD2UEagCur6QDmdtLR7oPzRHnpJkx4c3ugNr1WPdy6PpIdiV7yr1GQDhS+AcOYnPnUDv2p2J
7JvNCs5zQGFX0nzSEif9VjXCowLLX8DAeLC1+CpfsjB4ZwkJKvDGkDdRmyUNiT0N09YTlHuJyKzO
iudseSSmta5ssyKucS2pFcuH0iBDJL0SCvedYJwq0IpIiV9ZePERSHHByL7XV8vlUlocQ8D7uv0Y
/uOOftwEZTvyOMuG7Oi74ZC8+4epv6Us72VqfnZRP5DfbeRkTPtpmzr+NxM/pYB1MSrF6qWw8jNI
aBlIPDWdS+F5Iru37upnql5f0il2bmZKOG6mq3WHwfrATUvuhAxmM3z5dd4ccbaNN7FNcYfl8pZZ
SaTxHWzRkAJiBfi4YmYJnEhZ3W31CMY/oPTHB1bJkmtdqcGh9og/5W7RsNqsm/rt753xf/ryzy/w
KyJ73C3K1rm625/5qPwbtNhcDIiQ77flZWKc5sQUsDiGxUN8KXlWacUkIBXwRVtUY6ZnSr+K8WxJ
10T1EBbX9WnSYgRHAbjCXvI/Awt1t1QQTcpqAHJuyg0PAj6LAoj4VhGzD8OViVxxp93/hfkrYVwv
KHJPI+cUHbgsUx0C8IPopDQBt014Zz+lgm5t84yhEAF1eG6whNTtV9+2T72AQ1mIoSp5Tmo0rTDF
NeWPISktl5jHdnb/10F/MMUBGDlITBkX48qh7UXQI3JM8QrJtzu3f+yrGeroaUPOBqtKG6kojYOW
G97mSObbI5jTFerkqDOWoUG4gkXHMVOltFIB743Zt6aUjvxDcTgRhrwcVMJQqaqWpKxXAAlpeICq
uz38oJ2mQkqHA3UyIvyz1bP3cr6mf4Jdc6Us/4vX/7QjPzft7tTOVbkcxhN8BO4lrQTlPJA7X+dE
p5DNjn6Me43TxKkKQDX/u5bGWjWIifvhTnOmQFPmfJwQsaygdmEDC5LrXeXLWK1pWNEROy/4I0HA
SXbt0lGDXMiwRbT6q4tOMhr3W17myQThtMNHUVp0VfZdGzfyCSkCrovCaiK62X0huP85eGXIF2qq
av85TH+97B7zKFcZ6bwlfbLyOXndcUoJElMhdsoUaWQTCrZaeieDm8ZOq4eyYyjLRkSkfzV0DCvQ
m99bWQuSa/E3HuH90NtLuqooYL7Mtrd0XOURq9WDxVznmTsrNS5mLGiKM6g7q96xHbFpDcVKW+/x
O57wb9y78tcb/aFfXzuF/vhOzYnTNK91hvwtNIAnQvP82VfiJlYvHGyXCT2kZgXDUcuHODW4weI+
UfCBV6Ff+1yF9NFykxIhVwDEhBXbowtVdF+c5fU+2jfFTxbvZTDEj/0E5Nf8LJWLkDoMWMnlcVby
ox7hl0VOLZWgILURwQjIrF02XGKSmjkb4rAb4R3/5KwegUSXoIjCDA/RZNPPxbQjOcwy1nOyZP9v
KnYwD0R7RnQ9e2UnUDWfzsobSWnjjEJZ2nqFwG3E18fgzKCXtRUxO0cG/hWk3n2MSKaOvyY34yKm
D1XqfTMXFGXPmoOXMLPFMugvd0aWrRRWSVGqj16iWllq/v4xITMyi9Fl9BeMOSpFiN92WFUYz93g
CdCAOyWSRwN7p9aWJ50yDZFaQy4fWLIc18c7UY5oBka6UiOTTcv64XCPyrHwLEI1VV6IofuUSW3p
ug9b5qIrVHg1ZEk37YQHpJUchlFwNn89BLHH+3E0Pj+c5GxcRhZsWV72LWgGIwVUgmGZajL2U1K0
wloX3bOffCeTRcAWDY1ikTfJBzE2ow/6TFJZN6mXhryAbl1wqPznqDx4JAOvo9PTpbtMgzS0Lx/I
I6wyzU23kf6EMPGHcVu+KIOKTfZCP4i1iFBjRbuM9hGQiAGmSn24jh9J0JsG1s3HZUq9vemTFTmy
GQbvkYW9Fyc4oqh2Lai2eB8hCNCbeto2s39ynaZQSSaC3xBFQOxZxVb01XGkeiaoi43XnDIOUBKU
JGHG8f+o1LH/SzaTwicIhPeTNeuWVRU8BQZOF+tq/8bfl6o+hUNkYnUOmmrLmKDG04SKICAxrKYS
o0hxsYdAY8XxmeERSeXTKEyMv3cadz9Dwyuo0rR9/HyTx0I2VcPlXNvhkE65LUWgh9is9plEYphk
byclo2c4LsJ5VYBO7ttoZsOjLFfGnhzs3QlxEeW17XxNG5j40LliEjBmVNi58BDJe+dFNDdUyA2A
wog6WmsbI9IHzgF2Nz1prv2LduKBksEfsDW7osG9Mtgc5rYSTL7Fk4tz8/9LE0WKA1riqMjS1Lo9
LiaV67zZWgxEMwS4MsfWVmudxjQJY7A32uqURnEMSNb3QqD7d4cfmpkUZ0UEQil8rhaKgdOBXUEd
icHMrT8mESRZRwacb/ZDYy5n+HDtPQx/ypWfs7i8ODxCXnZZttLW/8vNmJuQe/w2VqZ1y0Xgdnde
LmBPjfNqfabNvbr1zMx7IQ5I8iYaEesJm/5NgW4qSCIgTJe4Ag8CLytDo1vohzYxH/TwYX8vunVD
ouY4B/dXxQhoxNX9TrS1QOwRClzNgHPSfrevWpBCLKZ2niGqW5wnYSRBTVHSYPGBUaGcjxRCiULC
miqWBNPkpEEi1Q9uxUWqAk7Ovm71k9OTXAwzuk9C+LRFpf2/OMaQDb2YZKkY1eyrPnQTBO8XF2lh
WlwcOfQ2Fij+8zUMEIX6W36EFqvdmD2oE3op/A+qFkcBK+mUcqQQgKbf0q0yFYdzWZMPKxlI/JeF
se5HiR16ga8q3Uk00ys2feBNqNi9YnCnMZj45Dz9MQJV+2qlBxbTHa6wOr3iWJKp07FLEPbXd9zd
tdBYhpyXrEf40RjAIgmZbmbKGJjy5+ftn4fNZQC6LIy9MgdVWpyh6JBu3kxwEKadH4NZSsnUkE5t
Tsq9S8vKlT0YXQmQOPvmQmNjDWB/pNDy3aSXc9AgZaxOR1M6wqyWPk24fi3UUb8oTp/kmXMHTiJZ
tWK6QpUYFwUMPOBIRQD52xOAWE1IY6rqXLApPalCLdErylEyEnFH3u37+YX7ZvFQYq+lZLjLi1F9
fJStMWumQa5EFyMLoA67gP32A38NlZvETIQ5jKpITe87E5rgTIqzXzNieUbUniDozJnbV0kov5ZJ
Vu4738PmLkuGpoyGNTTeug38BTB7dl1ioTrbt5cOQ8YZs8PQe1MlnBJ5lcjCHlVnI64cOlpfFbLd
0HYOA76dTn9wf6xIjJt8geBu+39i2P13i3gil2Q8n67KzJSUdQRfLs3vhCl19IB2wiFNpxozB8Zo
lM3r9pCsijGu6OID9l4r2WohMsIUYaseSRQwpmlg+QMb6apRGoIZ0Kg8uIPgpibuGcPShp+qZtxx
AocFKg+dspMp2VbshDiSc5Q+GDWAquXQG/hFzOvxW7M6iYA6y0226hiR1E6ZmDYGHIUrGWl9aRf/
FMiOq07qiXr4nOIf6QoIQW3Ub8oSgj5xNWQLvBDXxMd/z3ZEkFlVy4YSQi2lc8qeIkpxRYAz+Rd+
tm0UZSxAcqmMf/hy5udxm5sV8Y51ajKzWO7AMtJoS5cdXpfa1AcaP9vdqDa0Dar1DhX6qaMS545o
vmu/j8dS/ykU8LEMvcUcTdthacwsu4zVVvkFJn33BYqHnYGB5M4TMjkcz243A/VN3uytFtgowHEZ
257TkZUc17F0uCh0y5iriWof3iX7QvKxPKT9q10BC3bAgYxQ86cs0YCwLrFMRT1DG0xj1ummpyVp
THtmwd07bnV08aO4oVMu+nUmxlB7/waJPwQDRm8gWNEYqsf7WNO9+G++Nh9PJYNmoKCbd1tTRUBQ
KGh5oBsJpqO0pJPmaKrRfJalGGwJtYSY2EgyGTlnB41Q5zbyOs7PT6ZFqC+96Kf1yP/gOSjva+NT
R/F271QIoGejazqDdaFANYfkP/mkdBvWALHVdr42NX7aJwVAgaIbhsjD7gXrKyoFq0vqVxA4ItU6
E0pLRQbRNBHv7Q8vtKXQmkz5l2HzwM3Kr2qrBx+96ycoj25r1RzkUOTTmLzZwUC0rNMPND6XrSTA
i1TJoJeJomdleggIv5xm6Jzgei7snD4wlh83e2n4d+LuY2ZUm1Sf1XFsVZCqQa5R2sXDpAHEVA81
An1rfnGZ7z3p2tP0tWXm/cGv8d9cSebAJgYu/cGSFc8xnV/Vp7RdaEB6EyF8lSDzbTbixwaPjOsN
0S7zSkCKAI3AmXk1j9mAg+IVfGif7IFYmtaa9ZbEBzFStnXw9ycV8TM9SrqyCg2Mz2w2MOy3qFpA
dlcBgNU7pqQRCDmxorfi83qOktbmNwSpwFww8KB5Z7c2Dq+ya6WUsNpSTKIkluPl1cH4I8fNHq8C
7rqx9nViWQqqWY3k9t9LuhPifegp7wlF+It3s1L5KosmJKoqYNjB6nIq0hNj6jl0zjaukwibwf0U
PKIlqF/UCcONGEnRDK51RcdThAOSZGZuCfqc/i+1n0YAr0LuJwxvg6Xeh2HBXr5xddzD4JNGlyVk
5DMp1xRKZ6go4Z+NkYQr8dNvv1WJhm8UVjoCx0K+LVsyOxJeFP5w+lymAQyNpiwIQPXgnIhKwb57
57OATZ/hLYBNoHBH86hsUyHcoEPaKP/GVtLFzj+0gfhlBcKmpE6ro3pyQOBPBrv6/RrgykaDz5Jd
lkJoqUDQUywpAf28bzptP8AkRL8ShuD9xGg+OZwyjzSnTFPGP8iE7hqst4KoiSB/sxNvNcTxUiLL
3jYiG7JEI6A6uWjHztwkaBSF8srhoeCnQdVdummWpccedUyugYL+pZjMFLmm3Eyo2AQ9JEfNVYP1
43QOTwwk61RzPYBton0e/He7xn9yOJVouw6zWCbimyfHpQjePMA/O6104hsDZT9s8p0dgJUXGt/c
F6XznEXYjySlKQdTclz/r1w85nE4OAEgqQuMa4Mf/uhW3Gh/YUGaWAHRkE3bBChL+uEzLUW5kxJK
zcq3hRkhtsKW6fA2JC9A70AuulEOfOeKIOn/QMYxMvEJF7Gum22t2B8saMP+QPT6Q9wDEWhKC9dB
X74w1NP8GW/CbNgiwy/OlyG0S4DO3+peRUoJSjGj36R0Z+RtceFjdSaGeQw10fvNYwYDwAFCmzJA
WsLkzRI2MxalhEtcvQUUaM/eYFVKo3+5n6dALbg6XmzKfjtVIjqHeE5ic+esEnLaVLPK/a0jRCK5
M0er1Ac0XE0tiq1i9kC0ENiqT6w0Jma7xAMH9QBH5KXIywo2xCsDSvglnCS9+QXRJfGyHvXN45SH
/+981Yb82HTSt5s7c28nshHCcp0/hZqSy4flx6yUCFh7MKZMxnnM5juZemYouVEIWjmUG3xJMm1u
a/7nRohbRvfJ9iDzj7XatJrD2o517iBXv9hY8QO88knj1top5ALplylmYFP1IM1j0sae+uqvzZ33
sDRP6ofSNdXpVRXy+M+q1wMOY6Fnbf21v9uRxEcSp1K0mIsCMQGCOkmCFj96mCxm0lXVxwqKqvKh
3JJH4Kf6HPxS083yr2e83G7ql8L4i5SXJp7Xt7dh3sJNNWbqeR9oOakwEXkpotzrPg6j97dXglFj
W/QjpzK7Gg0kWELhSSqpVQpexf7CmOKDYL0cyOtzYOVlHre5o4BKOhIXcvTube2AlxsFq8yjqmGN
jq5iIycHUwlJgEeTJRkjuH9XiNmJDmYR9Rt987H1kOUsK2nhv1TrvBvJKidD/rICxjnjIQctyifm
BxIE8Q1g49rhm2rb47DqXrWFVAuRUlMbQwCfPagsoYUwS3fsAjrQtN+6V2Q+PnjeXP00AdxzgTNx
r3slOEh8kUZ+9cTk8B2yJNKiQuNxwkcNMrkahWgh/Mci3N4TnDwt8dn15oTY4Yo3TU1byWGO4Mz/
IvTthltrBjcjZf5Q4ijQfDLoxHtKzjcCyqfa3+r6g0mZ+0jFoU3aT8dDIfVziIxLpm9Bdwn7R6Z2
NsFAEwHggyep36sRFT7YQRxWARIAKvKoWDgDnOuTuwzfe+chDGN38lEcZ0nX/pyloJMwavD+jH2p
2ivmLceAfzZQOS6d9C4pYJZtVxuPlYJdBJQ/OTlbPtnlLpeUzIrNEv0LRsj1ZneSAABn0GHAVcsP
ajpA3CO1nv4yNOyRV98Y1BgvGkIKIBtbDrhsGcGQk5p7wymMMJ71c2KMKANPN2rtxDGxOSFvpfz+
t+6rgqd8K8YlEt3jj/qXCCjsuIkf/inbmDl/72fX6/OSaSy6HPtpXWhx6Y2MX5NUyVYYHzB43F0j
a8nZ8kq/2UsXejscSJhtaomN9lEA1gPOdYsRX0YWzLDp7wCFthf7cXkq55yldB4G2gnakUJKrmF/
EEnQX5pySik98NU5LAGgbZQKH4mRukzn3WCHh7S2dsIUTuQGejsYA63V1qBcmHlWEAmVUMJscC5v
TvwBbxAXtwjKq5uHX8uiKI+UqXBqPerRV1AdWZTvtemHuZUm15hTcYHfRqqCkC604FTujsd2ADKf
Yahvn6UYjTN89xpMlFp68U+h5ofXEG23enyREp37CMCWFOQmbTNsrQg6NdjG0e73sQ+H9UoJqp4y
8pdHFc0siHPW84lxH6yvsVhdaXraaterXwd9nzZNoANRkmDsXt2eFI79nw2ZKLaDtx+9oY0idjNF
TbP8ToD7J8NBOqBvvCghsycMx+zdFb4O8utZmXcP5YNelMCReSRbcLgNQPa4oI0tNHT0sC2e2dRu
0CKp4VuCHg3vZFYuPBipr4kDfxTF5z9W1CSKnRdQ0J1wduxC1TP/rHp0/9g451m1J1fgaWjs1nn8
dcFts+z8j7SoipVPRM2jax+WHTOGITYGFvu0Z6uy10NnbDy8tJ+qfOxT16vEFUdeqGQ52UekAbkg
z+dPW0YOg3sINrHrtEp1d4A4nI+X5M4F+kpv08hNbGfogEkNIg23rFzuz8XBuoa5v2oLd0diV9RO
XLl5nHrcl/+U59zkY4k4rY+cav5cfsEchzcWBxYzIbqeuLZXv7j0NO4WOZLTYUZlXYkRe8DWQYz3
BctCLcjRihJZ8ixz7JgHQGvcx8w32UbB//i8MrbYkaA9ir2OhDS9gqSpOEv0b+McQTcFq6cttO6U
e5cqZeg0VhK6PKwwemFZJf5kulpaMYMp6qYnrarKvCwTBP9MWesT5U9/8O3XehU+zlo4s4CHffyM
87IcQNR61QCWBRwoE7v3emIYvjHKXWPaPHB4efRYgDYRDim09oBaF9fPcNn7rfgpEfHnVd7+xEhX
n7TeCgjB1ErfFXJVoQSA38aYpd0MkbD3mLvCUrjyXfYiGvkZsQNu0Sya4weFF7rUrP1OMZuWwRx8
hLFgSdQ2FmDUa7ur7MDLdHXa8cDITOQ2u5whP0uh4jElHQ57XsyrQUftR1lEblGp44I1J/3W19SB
ysaNBFghVkOhhmgc2yUYySLktzMDCX2MVSJrQbv4lD1WUmg0DszKpmfQA1UoRXV7jMks3x6bWydb
t++2E56gNcKA/doqBZdBXxJhZ+PdTFqFt9IJCjoF15tmMhh4NQO+84SF6gNCXDalUxFPOZwZKsH+
yKJbDyt4bunqgBTEaQN8/DtIWBUObqKtvTZvgzNyN5yLJPPLl9mrm83OWpXxcXI4UdoGrS+lzjuv
cv+s/6SMUE/xxCgKa0RxzhF7sxm0NEojwo9UIkgf2s/n1ai3wcWHMjaxkQpxt+6Udnrj8uUG/RcJ
+OK/uHY52Nl3sJ6uwCwSi4ohhrpRkHj3N8sd/oVyFXpTaBf/ibHbvnCzE8XNYC3DYP7TUT2cIS0u
wk+SsS9/2ElNFeNUxp58rUa14xPHIz9f0ckV4VHFbAKK7hr0aXXkxLkyi6c8SaSg44xOiBYPyGJe
28RHlQcobR+LrmEEyQtWNm+Li7cOnbWsVMevVcWpgXjhzgxtQQ7em3WseFkpgxRiSkGazCgX71kN
yQ/kTo7K1V72GQ3IyAej/FGfKD8+MIyWwIcSqaksFkiRplwQrSgwTO617jOZwN80XvpCKqloY7O4
skJHQUimos6HCauxY3p3jlzoeirmCs46AMqugz3i0ervB4t/toYpd5PaNRhnmuFHi+e6zzoIx7Xl
lUpvKc6hCIF1P05d/YI2PU3H5DUiiMBa0DJkHTI2GqtFRgR/L1KjRCHyOpQPY353vvbF8yLWaona
ntfaldZ6PjTN/JpHdm66ajOl1w1B1jgHC8Aj2ROwpYrphRRZldzV+z3cuKZZ/7cSjr0EN1Lxk0G7
l1nNu2yZmYRGMpLggsllzSLfjoOoFiheVT15SFL0NrSnJfDjAD0icuEAoeTfNOd+WIUH5tLD20Vw
qKuujzbkvEpLYb8B+wdYR5G1psPobZTHOnI+jX+2PFKRBvW12YubPm6gC7+sOVaFiNP5UrdWqedB
/GQqgw4SG/YV+oAzZTnBUyB0CUUm0c6QFGh0I+U7JJsla2m8IOSJXs7agWczPCo4ssnON5gNSxWj
xJWiqJKUSKoLAHO3Fimp/0mnR+hLOlZvssQ38Qz1eab77BKd73cTqvYtYIbZagLBa8gNeDDbiAEC
DgkbHt3BDpzgy+V9A8RHhZRhl3T5ykk5mQ7qUjzRLobvn1FMxNUlTdDMDdalL8sBWQ3nWYJZRjsi
HNgfNk/typtiJK9gkILr0jKuBhGhJxLUHZ117lo5ciUrBubpIRKykPbrqLAqObVT5bNmDOEUGcNJ
R0wIgjJMvVWaSgrGHSmwqyIsYhbylGOxjjMxvL3CL1Xyh9uRIEq6DecZD/0Iq01IuPcNK13V2K8t
k3qQc0L1omH7XDHr2LlEdarHmhkULlc3o3xa22Pg4iQwHdRw9aPWJg6hd4DpXNG/MNqcDAzk56kx
KIavB0BYXKVnZvikrA8isrkURnlTS1sgJF6FftwGH5cLMkMtObyji9BU/lB691c2QAK1x1uCcFEB
rX6fKfV6r7VdwpTVgj7V0WUWyv1hzGatx3Bo3khoC6srGyyQI4nDlxIuWFTAU+eB5oO+cXbT75nO
416Z90LrqfNcmD6J6Fu4WuAt33yqe0leYb5gesIg0iIYQQbWqIkDVhNLJYeOGEzXpwnRLrr9Semp
Mi6ffsgTF8zEdP5Vw3nyuZm4zWX9F6DQ+AAPa4FmsJTFVIr0PZ3dE4Yfd/T96dZAkzc2T6I3IK4l
Mk5LuUQsrnF+EdMiEYGx75+WnGy8oriT8nsGofBQba5bdyYhVkWDfZFLGERdcevHfklgaPVTgdcI
4zuVhavtsXXtUGqD3GYIhUz8M0MAK964Ziz4afSu8IrJQlEP21b2KZ92yEn3ml0aRX23c6tQcBCi
SaQ51Q88A/nsxEpxxSBpyG91WKeKdzwkcGLefdk8tTIzkwlu+AcSLdrd1UBHngbkiJKmi0wOomjO
vl5kO+KCkcsWrcHuc5oQuxwz6oGyY5/QPKrHaBOCd8weD0avFiPuquYx9VDCFBFlMwYsjJ1mdj+8
9Fg6ZUwZLjaWdiGlzVovF8SF7JeLc8D/K3VH7tb+OHEFfN9kTshPGVQ4mgZHCDYRUsTLsBHye0Tb
A63r/fUZHaWUjDbpkwzl056gqOMuLzs/F/cwHSzbZkHioMlIiQIm09qcCsw9papGGioo8bzejBtV
Msd1T2mRKMGAVUhsJJnqOfOVZXJaoaeK6uOYMoIqarMTJuevrWSZqBhB6wmsRcWLCV/k0bTjJIQZ
gIAffCAnW+6TZ1rlXPNdU19kyofE4z1Z46iNS6MmhvGlIu93FiZLs11sR1axQCwJcjyfxH4qU7gB
scxBpJDEf3IW7ukhn0r6kOTMgBmlexJTtbtDxoa+tfYYbSVlTUmJiVDmXyVFPNAmXR27sIu46XnM
ykvvwjirDErhfotB+drsNXjydQ1ZkVK+P4XTN+5bANRTz3Y0Xppk/LR07/j42uvGZFePuKB0NzoR
Qvx251LkwqT/kM31jxDMal0UTn2l8RSYKzTC40XJHtZFu6LfFLRvK9BfHObHvHD7XoA9Feaxyidv
rrBoVPbVqTQCMU7MXv7YxMed7K65H5a34SK5fVIgn+vixGhsip/Hv6Vkr6xif1QS8K7J9Flf4cs2
hGxB8BMjQfl76p+2olHeFbm2gCNSrAxdDscnv8eU/W8OCXmu0fIRhuRsTN5Y71gJaQ985vnVDNBy
AZxqoBUKNhQx4Rx20I87tuTjY2M5Alr70gWhx5QNswfBEFZNyo9ieFDR+AqpI/s2htaU39QU5CCB
q32rjp+dmuqzlcI/0RpSfVnRzV0x9IrxCAasVnIlxp9Pp1tu61BgyK0jDA6HIh4H28s+SninFAiP
bwum9sfvkWIIZl4JUt8JlLsGF8i2PRXaiX5mxuVB1CTiInjfDEcda4J5TRktP1pBXajKG9FQwMEo
coikM/MtmOzzi7n1re73hs0N4nS92wmQereHN9qvzGiBFbZqTMt+zgUmPt9V1kh5rnFWuDZRSB8q
utXByqOMYGfqATKoKkfSNjZCc0i0TFMDL/r5/BsetkTMo0ow7RcqiSQhK7l9LzHPufWkBPkMITjE
WElHkkQMm2mCr2tluMG/KeinneuMvkBz0x++0TMrIi7B/vShe0IyuJIwUze4JjG2uxrMQAewS/9E
M4Mh7pIASohPp58bDwOIkw3R53OcuX1iRSmvN619ln3fk6tie4IBPkbu/ub8X5CVQiokR6xfssPU
/yMoGzxYdb1mlDM5vcSOFECw4QUN1IODxIPdlnn4h+aD3fk6170UXm7n/zwf0MXtF2zwK9BPv2S+
omKQZhj43Ih9wSQeXepLr2ok0ahUIt3Ii3SVD+2a2WdF1Ds/+MeWB52qmfGSgbmemGrVInwWrAbi
ExtVIR3RGlSofxy1CgJq40A7nFMsSwESOrx7vhhE73iKc1fzhNnTNkfKKVLNjQ1I+dVXmzLJNKOX
v7Pi+VAFeIuTJM9V/H24qN0vgLeA5Utz1rbYRsNg792+WcYCHJbq3cP5vVxEFcCJ0GGJD4bKfBC+
Xk9Uc9vR7o7k35jV1Ul5DQxRZ3CF+PZkuCq6wTVSmjmgKHh/j9GFXKaUKIuvEh8F0CPVhDeF+w5X
IsLx+hlu9oN4WPLxvQ4KAHpXEYAX9SEvZqE34APY8guzFOSunxOygbLBWXwK2kCiqoTmdDrahRoc
76zu8aoXcGVDdP1mxM/tz0p47gM25+4ncoJfqkT6cR0V4DN9NreS9uoBPYLwESZQSP/uGNsb5au4
RZDY4S+kcRzdj3urQpuHSM+iZ023P/WRjJ/MMpQV2wDSONGWpW1UYmnHtRaAffJpN5YDAEWaFji4
pLnt2hJUSdPiyeqz1vWHuJehxKYQQp17ZzZHTPEMhkbrfm2PUWYrE4qtS/m2K3f7/eEO4nZ6FhzG
1mVXJAK/mEkopMyzA8CeAon3E1RVnr2SW6M5hnvzuPxxgcjnxWbaxD9qz+jmHBKXkIaBtFOFBgN6
vuI4D/nZfQffcXdX1hZvtgS7YXoUg7zh7NkiEODa2EcREfrXpcV5rGeIHo/fglyn8Z6it4OjNqoh
/v6/AE0hukwsCnegc8LIZLTaGsGAn2HynlHDhF66OT2X2hxDR3EO2xgk7nchYw9E6FvP8y+MJG7k
0PRd42yMOePSBwlScksgaS3tMFze0LpFlURqlzMVmdA6Qbw4MZzWCLRC+sJcYQn5c+K1RoHeRK+L
evhI3n4LGrz9gZILhKffmy/s39uLLaAuyK5eUqX8kdIJ13IOI4OLivE8rSjqRyuLUCQ/6o73c2st
hSBr/uYkqBCG9NOXZSL4FBVNbxH2UwkXmig9cUI2WL8v+aN67LHgUlskQpTfMu1TblgvaCGgbQ6d
+btHh2BQsZFRsUCak1DLY5QxHudzlh8PXe3BOiMHVICMBS6ldgd+sTyT5zIvOPepVLmOU8JphkOc
n6927WXhZvXusiJdJfX2VrAgnVt7Zw1H+BeOWeyLN/hYqEpvDWy8QmYW4ejmmpuyfbVOpJLlOwjg
vUSOnUgLTMVhggIaepihFBycTzzDcSxIBs6usj9Jb4SMRrlMzTRH9XEc5xSbsqXNJdMZ83jix9Jq
76uFr7DwZLIIY1IaBbcdzhnQdB7Y9dRppywuf93mV8jeFSQEq1Hxi1kxwhLS/AN8g8GHIst2/G1O
P/IY+I+B4JTaYHePA8yvM6irP20vAehNmiAF04Aa6Mo7Ta+iX+W6DUOspF/npp1zLrro8rL2Z1Lu
sMaieQcWaZlAEYPwCsWNijL2hYGCjUMaRPFebBb8xdqo9zX4vlElpjK2z/tiLzmFmWnUKQkkupbd
IiT/R5s6+FpznBavvrPdBlyLxLjBeAINrrmO+AJ3untZ+5XLdEHFOsXsVNcLuX5Hm0Yojm/jhnz3
wjr8Yp0FFpVmCY+4RMR/dpM8cA+UIq6hhR08JX0QzBCBmmh1ha9JqGTnDbf52iAijgmJYxl8yyvb
7MOrAhgSFjj+SQ9ucofsdOtrK9TUz+GvmH+bgHCv6pnKVQfzVPxYBKcSexTJM1TdOrBm0vhyUr2/
3MVoqcp/K7GEvkuqZtbtpjkNX3sjXJyGJFPgYV28sQguo5zqB2OniT4iv+WZb3FDBTLLwmpn1Ega
mzMXKmNNTbGWESZlj08ilz2wAG9pNdtS4I5nMAKz0nc9/tWucgGWqywr52Cfzm3oAjHtyDp5EO2/
SGqMjA17Z0PjBUaczqtC+uknUkM8FPcYAM7+7h8fhstqafnJSDB1+GVW3Aapj5ODYExjAA9tHTX5
L49Y7JDCJunHneZeYO0gEVx5DPdyTQ4pKeh2q51kdjqaTwOQ+QlhpwaLK2v9BqnkQG8acj7YJf7R
qxFljj5d+lhu29zRiddgY2jbOh15vMUuM2EE+Ay5CbAWU1Ag3CSH3HTG7jhx4ODHBVzKO1nyh99M
PpnMa7Hu1n4saCnKNXnZy+20NKKhdJb0fQzNW+K45x2/ooi5mb/YB9FnOUK05CfNBCVHawT64Uu/
+QVH+e7WZmzZfXedQVwRTBUCO5K5i6FDsddum523ZsfcoBD/K9qTsCsr0VLqIMNZzlrmGq1kAUi/
knDNaGwp/j4aYmDnG+yXZj2xIEl+rBbB7ft9SgFTNrJFo5hErIlCAPbqWNSVJ8FHOa2eqPtRDyHw
hsiLvBbIXgYYvto0yuqQIk23GUVJFu6Bqkel7jAHnniQcbkhPNXf6V97srxMrisig+sqY75pDG/Y
hX/d/f79z/uwHzmDcz1SS5DjtTM9hfjGsyQK2ULPZCIwhrxYsuYOTut0Y0UixP3RInb520RtXq8+
KK9N4PMDqKR0eyqvJjKddJ4Tv/2dIfo+nnarmYPJrzs5Fr3LBNTVKeZOjrgnOQAqeJgp0SHYGtwU
9y3mYlI0uXlKcR9xbu6QlDgfxg42+Fac0bZ2yXhITNR0194N+7azjA6sZT4kd3teZmL1+jRL8Htk
DTKpboNjbJQvQMK2iC8NS1rX5B+EfyokqyX4SpVstp9LlpauMxdkIOsiNMttuMuftSmD13AQsujW
0G27ZBJtWMtPWdPJVb/+iWA6bV13jVJZjD4cGLVC1mM4vJ9Mea9/x+jHVCH0Mt3O3lmRW3c1f9Jn
YYpfDSnwfPeQYPLYD679KdGsomb9c/iZvrO2Cthy1GAFnqkqwcPaGzHRXRO5TLx9GGzDST9GfSx8
ub4fZ9e7vRSs7DXTIkUK/e21showhYPsey5d93z0neo8XWgQs9Mv9HnLvnmyx3h6/QpdTzVPOZVu
Uu4eHE8e8NT+5H0QlvLhN/kcddVFG4z1dGH+sOL0O1Dmixdj39HGW8JqsnL+u54oICWQ4mXfZOxU
5z48dqK3rH7Yl9AXmuQwtZv6Ql7AkgOTSn5s5Mew/u8PiPKTJWtkBz0WbiUKqtFqkvA23N/Fpu/e
JdTvo2ERIUU4n16CxYjZahUaC2vzQkjLrnTctuzTXsWbw/+RG8erpm7U6r3Rk9jVjVnz9v6FtSVM
y1g49SxT6nAb3++bOzqWRuKxtQQbzsUxd9kweBU3yQIRyb0XVlvIRPy/I1hYBlJjTKGjj5ARTqst
v0ga/3YfCkdja04y9gxEaFkFO3vCT9EDgfBn6f5V12vRRiMEgb9mOcDLcNIvA5urqKlPa4+G4sos
ojlqluo5E6jOowe1ZZ8emDj+yvrG0lS7xGSVwJU+23hlij93IzFxHUwSyzn8X3Mc/fsvOyxb2AZN
tcX3VwAVSE+6KrAZ59vKMT9MJbM1tvQcfRogfuWV8si5xPMcVflfgfRuehFiMp5nw4UEKVbbFZbI
IryjdmyqiIarR0k4BE9Yd1Cfwvign9LO6ck5BIlnGFyp/kqmU3aNhbiu6JUJWNOlNJFjtM5ef4A4
oHxopcLSpmx6rCoKC/M4TEjFc9m+PN62TllPkHi7kQ7Ang1oegWg7uqcrvyo5O/f2lxHgILS4laU
ymkEg/qUmJ3Ps4jbXDR+NlQXAjjI0Xvtq38g7ujMo/TzZyHS/mvALkGEyFcDKizJfALmCKxzrqQ5
GWGqFj+jXhpG2rAISuLVBzzIGOQKkVPyCuFugPhSrLl/xj2b4bn2v+sl1RENZiyfGlNPcCiel6E8
D/vc4JIT9wVLLtQ9mkl2tGJiTrdNTfUX2sVVBiYvjOnWVRIw+/JqibAW7mWBBmkG8kc4Bg/1caqe
4L5vws/ttrFDX4qP8I9mrMNSM7vS5H39PHogIlZ6GOVA9/RW/L/0WOXvErjAym/KORg/vRK8Klr8
BckPH9JJ5vFMofT1SUh/2r62frA/h2GEb0Oqb/jrZ+Uyhfm+/zlhOf5NtxgCs4xFXdLlNuXkZ4Gf
sosQpCWXqWCEONrCWhrZ1SPd2Ocu9bgqMiin6j0o6CkIMM2Lf2pJQqKYHr+HqWwm7P0Q/b13nXJP
XtTjawLUeMgMY/hx4+/MKsBcuCwedSe7F5e5kuKEwPKhNtq9Cg7lMbMLT68VYP5Im7WmuACRxNTn
oVYbT7V0c/iORmw7mYryWgwpXRmV0PVbJo5iIqfTe9l7VMkUgkL1FI7iQq/fKYoicMFUkaIgvpKL
zGz/3KiJcyk1Emz5qq1T25I1JpQrf90Yg6szE404aUZpITfj680AH/7ew5HxVPsG57mSI0ceX2fC
V/l/adil5uhtbWekD8F2E87b/hthhl60dw1jEWgxvaI0lnQvGQS8BoUOfuPpmKulS5bL0gufx2/5
4LVkYuIoVNLy3dZt2s20gD9zEGjvPl5doOqjRe2JEBjRRrLDjDVSPmfLO1H6CS1dhQgxvdO9Lh9n
0FlcfLV/P3DQe81lVtpZAYaGQ0+g3IStnuJWPFUcTJJQN88iJ+MSdTSyYxgY4aCnk38KKDbTyTuL
q6yXl9fTs/T5shUbQSHzKgdxcNpjIvhdSGM7hj2QQz/qoXXyJZ3ZLReiArx6Nz9YpLiXPNKMMeQU
otdo1XFtYHhq5MnEaylTWOjA+ltudYKvZjdqJmUYsod7o2oP9XkD2BzogDMnEf9QMdCK9aa7Vqc6
InVUo9pnC7uwoxruVlGkF95igYkJPP8zw3oQ1er0rjLb4rzaF/u5NLXZotNjAU63WPwUWsQ5j7qi
rlyfiEIoGcBgEp880Yo/yHT3ziIAxjEE3ClJz2t3bsqqD0tQTb8MEz+kLzE4ZUk2SqqEsWp5JPC/
TokI5u+VoxkfqR1NwKa8cB/n98bBqzxRFUD472RaPkkIPJUuhQN/oa9Al1rJYw9syaC9NrARv9c4
vXgmzKoRgebXQAUsG2Wz4PZJP3ECPcYmyEr/AhGP4gxb9au5peyfuR3eX1jhng95sZyK+qzZOkws
T6/PZgkEcs+GnTKQq+wTR8bSQGQnS0tKggXVjkaHqWMa3moQrcB3mV6vORoi4Y7VBuskasEl4+69
FZHwrm92EZPnpCyG7nPcEXSUNkUBroiiX8EbCpT3aD8RaoLDsME2GWikBJGHBCuos2//Y9V3JEwC
Eg3Bq3lO5AS29ymusyWXyWkGsbitfxt/yffkJ50MvIbWXKb4OqV/nR+K74YphXyKPcAEFv/0jSCC
iBGQQqfAycQujzW60lQhwBt2OqqkCVL6OMIPLXv2jLMDqzx+ojYIaxtzoOIhF1Z1DRau5hILD53+
cSTzkieQmmqlwLqojS/8mHSStk52coBZPXc72vIoD1V/vN8zgYkSPlz4g/1TGR7K25pLDKz8DfXc
d19ZMOPcezqKyPc/m0PsK+62JJpe+2oqMaCN7dj/WHcR/Wje2UkIrU1Bfjr8jy5mTKnEN5s2TP3j
B6d5o5cxNlqXBG+OesvkHFSwjbY4FN7GPONZ/gklySTY1/sMDs7emNle749MqJP2jL4wLFmMhMnS
Jt6qVD6L15L79TJjT/zuQ+PRo2+WGH6d3/UqiWFnHjYpiIgcIkwOtBdM4Ohp7md6783m+ZHbMsIk
jvugnlgmprN5vhbgcXSxwR+BeWt9rhgPxE2olM2QF9+y6D4RL+LhiEjvzUU2lD3DvlK3Yew4dldi
yhaDgW98dLt/Hh3jEPPMyLac1a/pE9KlTPBWVx+nnY0USUwYiIS/ytCW6Jl1cgewLi8uKvxoncPn
DuwnqydFcLhaiSxkwHTI/Q32ettRu3Z0HMI+FbzIEJVzcEVxEa+sQR7+hikGzj+bUJbZ7/BlW7uu
PWMy6D8TAbcMM8JOWAdber2YOTPtP6VFyxpM9w+v9ohAnFaP1/U/kTAP2fuoumlHVjbeqQsWSZc5
IA6iH3I/v89z+jtfTYlIDCgQZFk4NlYHL9vsbI25zV24+A/z1z/tHncwUICg0xFM63+KoohZ+TNB
xXqItOQ5UUgi4Y5gQk7xWn/rU22/agNo/wM0sXy5ZjcvCWYNS7j9ty4jLQZ8isekCfxh27ZoiGw1
8hn0vHOn2nDLW2/6T0imiV1BjOzLXh6NfBauGKh3EIr2hWVLL7oMqSWs56L+Ky2Qy8lnJOiu+wFx
Dq60kwqmqMIOT7OYZIMZrEftEHPw4a190i7UbVh5JbrPn+0TfkK8/RaxENX7Z4BBYppmpTU7UJO1
FIuJ/pzwGogot/MBgPTpdNsWPqxe9e/tHl3fhJJrEhz/+6aPQHOxgBllQ0cBvmNbTjvDhnX+KsYk
Ey2asbuJO7egTh545N1clQ54vnb/t3cRhkxwVuyrpapCew5dTAG16WopVeTfp23Rn4wu1OWrLV14
Nuoye/j4ZRoUTuDKbMqqBuXVb7fEA5YzEYlzOaMr92oB5mmA60T6iAcXBv6DMqgApr2FyVLZ2HkL
jv2WrjhrWBRQOuGi93y3byc9WO8N0dgzWRDND84+hnU8NPp73LlGSq8Fv8ugEstZQ1WrNRNLpTiv
5AmmTiS88eAvQ6nSOZUfKtYBdMvdMhu5mVyxIMPTtwP05nQ3jaas99x0D6L8xEGLc6Fddd9dD5Lh
mP7nygDClQ3Zd5EWddVqUAZmxxkO2JsZB0juLsMnt4dE3YCCmn2rdek2U4VefQUFUZQklnG1lEGG
5uN4nAzFyPnVDpFDPC+CjwGOzx3botdicgO0+duRpY8NNxrYRflcCFB92Lll7yBXg4I82hrYZAQ4
iCOyM9pYp2is0oWBlp6Njh3EyET2GzIGo5Y+D3eJ4j1GwVyroLwtaJnmz9Hh1VX7sTCac9f3KJiV
PKk0wWwS5NY5oKJztxUwHSjmttqPW0BJIOJqux6Xav/21CrviG3SP8JL94Ezen7rpmVaIGWDujUz
GN5SfNpJIQ9rZsm9b3lfRtV2Bb6nRj7bWM5fsjeDroppLydBS/IsnPlhzf+32DMpCet8yj9gQWOV
IlUiNoe9YMP2B5J9F75llzwKY4c48EMG+oSR6GoiGAIUpBhz8k1RJ45FTrVhip1pGUiRS+IG3ZAO
MEKGT5Afp1VE1Y7nQttTjJO+ELX/V7s0auYXx0ZVEbMHJRdzVAcrHQe4rlCjfjUntzhYrpuHBzfx
LtErS2Qm2704B0rhqhdLrudz1TCkftCFALgphuJP9sLgda5h4emgygMzK7geXZaiiQzsGbEKdusj
VQRjFPW50dmi8OnUsQ5LbXUNyosG7O5mkOuWlvRBZLSyvhBTga6RMQGLuuYIJ8QHhIGBZU3LQN4q
ZQTiXnx8gM2r92+qL/v000NBJr8fbHKfXz7AtFURtCHncysI9j5v7Jtla3VMp4OM5vJIRwYmyEVX
LAlbxayhEXFD0XBRGzIF/o/SFQ1HIPUU+mh14cgceZVJpNu1r3Mqp6QXvV9Y9iLBZdB5Ev6m/NEx
Bpd6y27u/O4I8KInBrUdsAsy2Jmz+oyiPyFJbCYxjvVMWlnS53vXnE/o6LgKxmVZe17LWvBCedRv
4tqYnO4Jab4J9CW2aNmnuRbMjarrLl6Zk3PxxMYg5MH1CcHmkL3Drqr7LVZ1Duo9vpj8odMWKsYN
ILBair9eDQKhW6ifm3X9ZuFNXtOI0lLwML4TpkXAyx6Dlavy2pBje2rF5xr/rO8JC9CbnCdYgyq2
u114Yo+5yRQuXf8g11zaRmKb4FPWDAX2RDJnq0Lr/a2KAurseAqw4ZysPcrGB60GpAXQ2swvgLMG
CUozzLxFAlzmkm16qSUZEDQwBVLpqPZjidSNjJDzhM+7roOS8LuaS+KuPiwPNsjyYcIc5753G8Oe
WJO5O4HvILmwXKEKZ/ZRSgt3y9UU9kgQKT46JyNhBph2+9G4LgCWWbpYe4KhN4/pjxzixc/JToPT
Herpweyxth++44tWswDbiHoDDGSwqjPudSwcPXvtHlBnbDtYfWnn/tFsNClpL0vfpdxmgs1yPq2N
1Z4EoWKUSCBEX0fqKom0V341Tpd8vsON/WZicRTugd8rppLNKnbjNwpa6KH0Zr54lwjfXaifKOA3
M0rIaezJthQFi4LLtGmT8qCar73qPR9Paho+aXip1GLJJJKm4ZYn/aodvsmHqtk7JRJJanMTKioS
izdRZO687GmGngpro5qDS7YOe+3Q/VwqM0bvoYTey7T2O+b7vfgSDCrkUiATE33sPyDgdnmHyZeL
UKqxoytakMCIu455EvhkPMEh7jq+z+Nj1cySLZ6q8A7upQjoI3xBpEDdPiXzrWKpTQtZY9m9a2E4
sQ/5+OkFbCOxK/hjrm6CIsDLUZabZ61KEqKsM7dNMbVI0ZlJ+V+0aruBI2yfuVYnIcsgEO1UlcAw
pgTXn2vCtHKNk11ynZZ5DpwqHUJMsI7RqT7wg8Afj1LbJ2A6wKsfuF1tuZaQ65j9z+BCmmVdcgE1
gp3qQQul5MfFiSIgVlcbQUyIr1q6qAkrxsP7/qpD05aimYi8Cu6wLR/rfHSZd5H/wl3degebZ9/E
K/QHJNh4SjFN1XRoAGd+uUzp3Zp+1HIIdRONT4v+EDULGXZv+LLxyjNyvfA3Hk1RzLGbcBdnIGP2
CfERLs1xpvF1NWFDAaDqTRgRASMeq3ifUGsRYwcXjEmyj6a8XSF4/LMr5H5koU4ySh/y7wMi5wLp
jSfV1Ew1xaPqiLlhcuS8FGr5vXEaM2gBYleU6DtDQxzUylJlo6P1nE8P3ALHMdukGscKnRFlc33k
t6oOIphtfg+MPjZTK/A2k+7J6JkqdZhoYVCgN3cibXGUWL1XK31dPe1k9WQkZn4YowMkFP7DnVXj
fdxPl7mW5WkuG12VbtIRxmQwqEfLCQGmgZSTymNsOon782bVidkj8qmkC2YWg/qrPne4K6P16axm
89USPxdKZ/YKFvcsQxo0+WZ+/wEsgcQxLSfJa/ckBkUMVDj9RiLhTz5tSXmAWYAgG8mxafu10k9k
rxMtZx51o1Rk1Jz0jAQiMECsQ8Y3rAUNceYBh6fHKtr9zKmQK9Cr2N8r3THvTWvFW++ex2UJUq6V
QkI/T/Do+Xxis1SjLalBdbuDmINCYHUDK6crtah2lU0u52jmLrTo8+aKxEFmURaa7vYdyuS8PIRB
3juInIv0GUerpCdClcIcHEOuiEJ4pVDAbLr9l33G7oel4D9qyKdNYPjEUO4gUhucRXtnDA0Z+VLa
qiQ4hrTcRKmdVKPxjKC22dG9cgiRt7jupaoECHajdonz6L8TfugjG3EqsVwhUQxMLEltPlOo2ys1
KLeMvqVxsp38NANcBaNl7Thy3J/vR/2QBR+bCeyyGLxtywRDI+uIFSDMoztq3beQ6RhXzgBU8R7e
zxWSceVSDghHTtF8Podd+61dCS6yJ9ZP9MaMPMrzdawHlJCK9JxYVblRGlTp0cerLhAAvXDS4Vho
bLdsVf9EKW0kxDFhS/LeXd+LqA+dlWebbej7zBvO+PsH0EOCpT67RRrv40eQeaH1k8T4ezF54TJ2
+/syY+oFXrLBA1Uf8KVQ5P7889Qn5dY1C29AobwLM5/xomTEmJcybpb7OCUaGVrfMmah0g+vjt56
AeNJt9AS8WRIMZ8sONPaqgCQzEPIph5uZQwZ0f8x8zkRBQa/PIZZGN2s3ZQpXtgkkn1SiE6kwYFD
vQe9jgrk3xYQr1cqYqYC8sw05/5bytlzYj/wneO+5BC+cMRjJxHzq8db56UlRNREFyVh509uOzTl
t3C0iYIK3sp/wuFdkhyfwg1bi0f4+2zA5povOimg0S9038v92lB0X9pWKMw8fNNXgyArYB5gIjtF
ldCrNmgnh/Zt7ymb1EPdlHZR5YLo17mjToaxpQkMtL9QBGEf8zl2iAjyVbPYBh+RLm4eF+G+HXrJ
+XDdQTm5BSXeNK5FCqEpssTWTHvqRJVywcHK1WxTzjNUCMSma5jcNSEG+pVklChLmfBGyF7CezBg
UxZfiwVbm+oULMEL+lqSL9qUOsSGQO7avXkCTsC2Y104t29etHnaRevy26piFFCeTeSG7orNICvZ
DDp2Drwh990a5ZX86J8lbZGrLQRojk8n0vOvYN0T9CVKrF7XiOGC2okKMqfGxo/t1qokJkD+Jobw
dtg1eRSIWv+XhJOWLNmQKWIPt+zxmCdFSsP3v8WG15AYtzvAfZAX0LngP4GqIq4tQ1ABqlhrKfNK
YfnDUB4gS6YEYiRfmxaK5KnVDgF+yatuYymMH1eqIFgY4msqiV0qt3xFbFPiJxw92uPU4gl2CkoO
bk/o0RjhZ0zlHMCIMtb9PJeV7bQ+mnPJ2EsNkpbxl7Xb5cM/+ACt/9ig6HVaSP5JqgUwm9l8S2Wn
ff9kQznkNZDADtxONB9vrgj/Gblzn7uexBK1UPowA2xXQyJIs0euMdm8NspYMJQCPNiebgkBhQEZ
ofDUwofAyuYx8F4ERCmXQWeks4xbnNTNMuQAEDu5+bw+Y2q4/qfh+gagYaYc+nnGhDHYQMBZZSzy
wE9qqCuMivShq74jkore9qev/8fWkUL/bKCMvpJXol1CqfHmoWB9LBRVzAa00b3eEukUH0jOPZwX
eZ+7I1VAmW57/H3P3Bd2THWByRcrkDX5pBfk46BE4Og7V6aNg0jTPTBlyZLJNRSYYk+PTAISoDas
xTiJ9y1j65e1VQYCeR2iJS8n+n7hYe457KuIblM3mVm8EWGygn5I7em5AMqOySj5gu/8N0qfeEpD
Kx3JK/X2lLe+scarnG3D4+Y49gYJwq1jEEtZ4o1qMpHqIB3ifzLA4dOKavrdCOotc1fbDCiDAifO
GD30vmgjs18BE1n4zAceZvIu5bKZpy38bgxCuYL9zUgtvfdryrjBRB7QgRUBwgSKTAAj0pc+qgSa
bLy/YiBIIeF9aunIEebVZT9zqQnIa3ho43E2fqPJspkWnBbwNKg8iefrXMxWsyOEkMxRK2kNYwLK
dXseMqJ5q5Cw5rZmHb27HiazDxA4TvkvEnvqKaIZ7MjVpSXkKzoBy9+JFnQhq3qEnLhsJMrk+2/V
Tx+Dh6U+2ovU46vpy1LCNJlAo62KGhOX55dpS1t8eZpP/UImXW8DyldjqzeD56KHZ1edShYT6NW2
P2VJRdtO8psM412MCwOr19ZgzZrq9KRlPTWheWc6YlHKUZnBfNVGeW/ccH+PbTajqHHGMdBAzw5V
5e2yA6Dkgm/33kBeAQOYLrynW66P98cFMY2XooPtMEkmViO9kvaGajNB8OKLBXmohCAMsI+oRcTI
yhkGjuJtiliPJgiSSEOkBQbcjzj1MxSfEFiqwzo30sHZ6Ya3dJRQhScCcRKyzkecRS2/N2BBbkVw
RsI92hbBuDy6K5f5jDRJNhhRuPTfd6xrxU3t48z7m+i6qIjLYI/6nohgDzIi4kgXo5qUbDJQNJcd
mg3mAFatgainvBpw/6h3R4c/fBV1+tJM/CcxWZq9fjcSbe9vsv9BqfOsHSxQiMrJ/DToekR3c8u6
H1txTaQzF7v9Sn/VnoTorsa40+nQff6pRt0OVOlzKf3h0EFBM5OBz4IYjiI2DHZW9MZI6d0kcLFF
RMI4GWJ2nB51cLSxw4XNnNYNNYGscUqvVx6vPXTlhq33QIi7pIBsh6syVwlqnkzIMzUO+zzlb3Ca
nC4HZx2JWDsS4xpyvnFmha152gMiaqhRnHnrkn7bnL+SZRw6HbURPOwnxjbT6j4P8znBeoNXzvnK
Y61jTLZ00xJXHeRK/qWmt0d45ESYZOHRFhR7ChpWfgJMxDLotaj+eW9J2FawdWhcCXt0MKkD8rqj
+QlR9i759G8fixtpSAcre7UsJAqI+XRCD2eURYCXy9w3I3aJsSvtKnOgnBOLklTBhuDwDvcRqpfv
hj0+x/pC15ISxdQpZpV/oj3MxkfaXcthSyFEEnAmIg2duNdG1L6dsKuwa5eECHFl9g/lepVuqaWi
yNwTMdfOQIdYHl2pWNQ4Xl5so5yu3900gIU54Q6WxrpUTDMuNDW2KdQfA8e9DZGs4STMz3D459VZ
zUp75M1gmMYYFSr09sLJQLWn9hjetg5mpWonG6ku2QIe8Gkcltbviuy38mts09qx2QkQVMtN66pE
WMsfYAg/bBvHK3/9MqZSfxE06F86C9Hj0wsO75mzD9EOOkJDv5LYELekntzAhytnbTjJUlBfJXlo
5ILZ51h58fhXau8z29xHykcM1KBoFyfcmDkSAmoJT/PKCTgMxVpTofX7NcpsTwKB0T4fGSc00JDy
DGpqkIe7bt7wgAMZwzCSr+0qWZz+v46ZIN84N7czc5afxtf4F9IFeffJ//wSHStEXc0PIWt+Z0yX
xvFZ4GW3dh2xGlELYE/dfFov5eIeifkjKoA/87EY3fx0OAnpmTi7g8RNZhMES++pcCt6D9ceQDg6
p0UMhWfO2lkwEIvI511sPrOsYaHuzfSJiy+gXJ0dDmRqL4nSquMoy6a8UJ9OOsj265w8SglQIaP6
BmSgIg1xdYsPiNhXDAjYIUweFmo04IdAwlSD/t5Eqxwfc4ZlQbDK0955lQTRg1GzB0bp+ogdxtAb
Z/CWz8AijSc8xzpcHT9l8Yr7sj9G0W6qfySAVTliGFwfUabUJa+ZB2bJHrU2kdBndHEFZBPc8brT
hft8SfaR2+z4CZAd20pdbucseAPvZLA12mM+ImOoLYcM/lN/wYEY4SQUQ0Gu9YoP3e8z+GSBa1h0
MTUE9fUleZ3Myzk3pXyX3tTmiAiC46dMfrwYm9BbnvpivXAv4A4AzaGBFaZM9R47wRKGB1mgLiyh
vdJ21qkBr0lRkrO7KlDll4mmXwTNnVYKGUgODq0J5uaQ0Sw6yG7QnSlK7xyeTThm6OepNquAg9lG
K/pbiJTAQ31VIlvIkuK1dcJ6tQel5WS5drZE2Ak1aM0ac+69MXIqTVnhUXvuimTv7hqKgJl9Zbc4
yQdlJJvjgCAZ+5B5ltaKxKHm1T69QQNmtzCWjdIa8wKzoelkU+ERQ35/EusOaDXamfLA5ukMPBNQ
lFqcgoz7eI2cWRLYoSultaVm8/WzlxHEM/xhdtvvPs5CtBv8GXxeXaizA8DVDI+anjzfWMZ7q9KF
pVSM9mrwdyZukgPi5FCQyhsHca3B5NK9Uybbct6JIUMeqZoEXGDVoH1wDmncwL06RZyxhb/Idw5x
4OPpH4HI+2oLBto+UijalmojLQvEgjw9m97mZYo9Loadi8Kspry6cTJ1UZmU3+4E2v5sc3y6HGMe
/uVzvdbhJyowrHyP9SXtIzYGQ9hUtaLJzl4SS8HJ0GzTNYwTNLSwemhCe6CJjWffbAdddrP8C+i+
S6AKM+YiFexJDMCzhJ9PlXsh7jTUqzJM5396Rb867/2AS0g3Qu1owlDyLLOZij96zVKM461JbOc0
n5uLrM3U1hJNN9G/p8szuBmb2YEi1mb9o1olUK53F/5CcewjujTIKkiuRV6tIJhwmvAdiQBTY6oE
tDwJzrWOtKl2eNkz3Muz7EHLl42LEgDjnvm57fgLUZkOLYqy3nwPCA8vs8lUvqBnz5pI8o5R9oBA
HlZ1pDdW9GzImMuyNAZLkQgJ15j3fcHWUJ1vRWhcOn6IJy3KykwZAWGmYhPk++aSg0dj247rHnMG
xXyUPF1oGpeYsZqFFw8m0XQMI1n9Mk4ECfYBD6U1MGDunoUbnqLqND5gCTYc76eWNenmO2ta/oIE
8mb0nXUZmucDQ9N+8GpybcI7xawUqhic1WgPobHSmyEDaRsNWUbD6JeJ9AmtacTapWPAlHmL+9i7
DYmZ5kw3H4I4KFf3WpM7TzO3TmNjCf6hE6CSM9Cjl/bUISuwbtjLMmI5nsJ0uqFVBBNoMHuIt6KI
hp9aLO0Qkqi1gpTPRdxkx6eM094IqcIctaKLVaRPh0OJxb4d2BgLv2SJoAtK1dCbbFaIacBP2J5E
dKllI6D9q3i9IE/1ZPTMq9dO/tCMUyHWx4vC4TV5mVGkAjayoNVIScK2ge8Ef6gnM3grxr4Bn99v
W/m5d0FzSUY19RQCC6khM4+g/XRQQn19bBV+oocuAf+K6IMdROxkX/Kur7aU8BeXkiXbtnTvHJ4h
fVtTZ8VNyic8OIRrrGGUzyMAJePLy66dliuoIn8vsJ8fyyes9x/xDdzCkA2xsRSmnVrqFn1qC+UZ
J/cqnid/xitrsAYUj0mOMfwh64L+9KLoYOuSuSIea2A8rZn42GzGkYQlwCG1WYBjM3g5OnJvgjNm
FDvosTgvBJCbAquZGfuKTQEU9DTLSrDXdSBYzKHgMFjFBXBpx4Kou0j5q3Bj9+vV+PrnQCwH8ZjE
wy9LEffiHQD61qRZxAkiULH+96dp2pZfEwcWmQG1AthKDj2Inbu7LyawSSRPOySAxF8vLRo8C8s8
pNlH7qiW/QF+O7zzIp7leFp0p/GmrnjyhgGAwqmyOm9haqXmn1E8MgZSbauqhFs6fHvCmzBMl+cc
91pdZa4Tar0o/KwzNKuWnDkGU5TLJK1sqQDX2f56nLlcbu+2/4nNo5d8Ne/BQEbrj19Dz26s27Ff
7dMPxSuN9kU3daUfEu1qrtJH7zRHm1KZW624cZYo4uNvSUQjBsZhE20PaSpv3JXtwUctvYijswNK
DJwBSywBvFflfBuNpNgZdi3DiFOpsU4x32XNJW1UoivX+ty5c0vTxY2bGarXR5VUmWLIrMG1RxD9
zOdu9hM8IIxVPgrnymt8vbBL8cmhnVUWqar2Kd+B6WJlSvtNHNe4pV/wIt/q22zKL7sBT+hrbObl
WjYKFvdp81fG4IzjiOGvgUTDZkPZfSAARomDlUsw3HYI7xETDeafgLyuaQ+hgsGQkDSF57wA8bm3
mk9TOjQtk4yBWbacBtn5/93FFvPMn55zt1jVaU6/g3RaEY14RNMt8E4lNPlNZBjOVF0ej86FqAzL
H8c7e4tLMXAH0FuP6KUXh8pOX29g5QFiyK9EEIZMt0Ya0rwiLj5suf1qHkMyPGkw0WxwZ2fmR2y6
3paqd6Zn2A3TKV43dXdSw0jYsq3K6naAWJcDAV3qKx1oc8nnt0Gh6tDwREXK4TBnYF7xJdlVo4f9
mSm0/6mHrGI+tPyGXMfh7O9unLWX3BEE7JTzb7SzSdiygbUosqTCS29DPUW2k8UeNK5jge3bj77N
yGyemr4ngO54GzqxmJCuypsE6CsVNCnwnOhaut2NOXEbN5Pun+QRyl6+jdAWI7/fhXzpmN5Lq127
AL02Eg5Cv0N0IyQrub8Vfa7ZCQ6mE/QpsKt97rsq4V2LRvEN6U301veYeCBL/zk5IG8IQCc3k6Lk
FSnCBpl/lGWhR+q2k5EPvQn40rL90Bdm/70+glNwKkxl5feaHL0URG/o3giKKb5fKENK2kn7QisR
a0qxuBeIT/FoXTFCVXLn/KyjRGoaxc5b3rCAS9OwL8P6Vyp33VvCiZc+r7MAJipYxETQ8BvzVEDI
8gAouTsYLDVpB6kEzN2UYDC6TyO6OrXHzVXzNWaLVE5kWBCX/nkx+8Qv2/PVQcNkNnBPe8o6wx4Q
21p25hJA5LODrG+D67kDqLTUSwAVgIGFpV32InKGYZ9ZG1+UsoIx0kKXRUiBbV53agqd0Mwk49MZ
u+oODj+41R0n4osptkZGLLe+D2q6KhFFSd0H3HdzkGBePMb4Sr5FKZac09e/qkh+Emk9i5wS+W7x
CmomLK0Y5ynQm9qFdB+goip0y7TH8NMZ69O7I/UYNL76QmiueInoZDuD8OpMDHvoERr2vbxp8xBT
fV1ZBjcOPYbQo99VkzJvaREHYyN7gVNgeJNzQwGdXwOGf5OepkPCxkbH3gvcI6mbKDoy8B+Rphh3
J2c8BV6COapW2YPTakO51HivSfn866au4IDBb7BUZwBjVh6+PTWlOqpOitSZgOElCcK+Hdmv7VPs
YhKCc+JBaUDCTuylweyBgkFqgf6GkZfJc7XIJ0SNgO8b7nv5b+FGEOUMuMIpWZMU4D9Um+Ko5GJn
miHnaT4ZvZAOAXqdooVUFqPv7hyiHox7vdOME8H4cmHq21Y0weB3wcx49HkwywnqaIK0sgo0et5A
/NEhH3lY2lM5W2EYdrWz1V+IHiyhxL60nbMAJrONJ/8i8tGDfD7H1QoYLy09lCfAT/ScH/qc3tIH
4Eozq+04Bz57dUft6tWmU0Mft6m0o+W+cZlvfo8xAKeKS+tvrnvPFVIFGUnlolH5Fp8BaqddDvNf
FXDVTpB+seC3a79acZpcAXZT0dosO7xEz4XsK43ck/7yNz4sWMFj4DANR11cFDP+FXYg8YnIMlUj
un5CCtjOC1AdM5OaXjQohOtxMll9eIujiBCZLlZDNQLIdfst9Wi44URJ49CL7gkVltqGJcd+eAta
EUXbiOFaKeLbbeoo4THS7IH5lTLjI4y3SxVzErvpK47psh02Nr2LLM6yoNPuwlmCMkGiGFW/D9Ke
bWRwq/iY5G/+bcDafOhrucmeJbrbqduXpEag2rMViFOXO4No53EirZN4UFVVF0/rbhM+Y+XYX6Ge
6LMtoLgVstgjq1FZ559jzLITt6t/6cSZSxATbvVTLCs5XNxm0vt3GM+0Sm1wJqKfsZ5xP/QoMpyz
cEsWwH2jR33JVgR5J4jXgV/NX6M3frtSsZ+S0ZroY2RzGxa8MstG8NRYQCBxh3OdmtmdwR9tkJxZ
wpLkud8fSGMAJwt+5+hRZV9w3h5cBEiO8psFFojfsgGtoQE56CvD46m721nzlBEdSF2JNmVU6AZr
dMR7BO7/5ccBbNwaMvsnMsYUBo9pDJ/3dTSDBX8NbGv4RM40+xx9nmHg+Dj3QyPt5AVW1zMT/gCA
9eRL4UmxH2LOcG/+Lz5/HxdHEOf7EN+yrua4mWlKBOjx5tD4poTfzTBwYanS1U1+/e/VjOXbiXe5
ssq585pfmbxYxBDr2tEi/StuOu+abwaS3RTGkexw+XzPdwXJXBqcEh0hLljc8/XkbdoelldMiSTp
hK25/tO+EdwJd5MVaBwO8rbxcmaLJJX+SalWzpX0BZOv9RnSj8L42WfBn64mgzBJYF1hylBUAaCi
S4+dli7hG/zDzg3McyIhkZ64Nn+prz2z6WGN8iG4CeyTJ0VmqNsUYkO1QUako9pK//GxhZhRmtIo
l2O+FRDl0QPdydum8MMtF4hC70Fu5yOPux6JRay/TBZuyf0WqZWRSzwmLwf1SkLtePo0S84rrl8x
V9407s4pAUgXMvLj/CWVJQfG5wETCPHkFNDSzbEjipTVCEby/ofG6TkNkLAB7mfXgsPr3kAHCrNC
xl8p6lVr5VduJlUEWlvDmRYiNf4Uq3LKuOZwH4b909L33ZTWq5loONJlxTyyHE7vxtyktX97sOdy
YzmXH8mGjccJNxtNhgiVrfBcqPlv/3Kqq/qqRRfgS+RXMcnzfWDpb0wdzQh631mZju2udkMWnl/k
rrjIoVMdFdxnedPzUxv7zbiIDO94UvY2jVyI8tBNm+xiBXN/oyxf2NoG/ktegCuRpLOZ9dAgZonH
Z+XibFBBve/1/s1puBT5WrckbVmyrerD22fFh/mKuFVnaKi/oBU3AZgrjlvuec4mZBfIHtremZSD
aB+D7dH1V7gEGrx5OXknv9AQLbHN279VDjsjYshhUw3jGwbFzWN+L/t6LvRqeQSX4I5isrgxQj6D
QRrYJp1N6TqGrxgd77Eaj8AAOWNOtE7kpZrRp/4wk0Y+kZ24aaeS8DHFaWA8J02d1ofHeVhAxu3n
y1rTF3QAm7E2h2pTuIr/niLCQVTyCE9c5BywG2v56oDOb/g7034FC1C9yQ7hC6xDDx0oGgzIHwQB
Rl8PddXVj6qK+0YBdvM1A/K8sdGGMDyhSEsVGDfIvU4ab6+9FGTdw4yyB7XrFL8tqaRdIo6pZ6wt
XdcSx5fEwP3/fn1MoZLZ+eMukISibG/iUCojcp6IWf1EI7tH6I7ct6aZhZg6fOjvq3Z/21dx+tlM
O10TIyYT7GCmFbsjTNcI3sts3wTvWfLFjfIOg7Srey/F0lmA/2Cc1dFS2gpbAF1SAn2eZ5izs7vS
hsCUV3mYEN5R0ubZuFskb0YEexzDQhDFjOUNN0xZPogo/UIPSRa82DX3yamjmb5/ZEJ26MZANWqM
0OxjH726UC1PsdsFqwJ+FZo4epzc6AM1pfACq7qPA4fRRXeHB2uCdmG387v4jf3qcKlThZBbiPA1
a5JhkcuMxNZkoV35g6vaj1reh4qpc6nOSOKBWtFs4gZ3+SrWW8fRKVww6fuT894oISyJMZdU3gzq
xER5fg4Vycz3de2kyqs6io49JLHMi5QUU/tT7gwjvFMJSwvY0fAG1r5oWi5W9DZG6zU6gQXMdAvu
ZeGjvuj6701ML3EbvZoPH1ZWHWY9gJy+MuNUWJepdkt/zkziSpWi4SUXQLNlLvQ48qM5V1Q8tckP
QiiIsBw3irYLFzrUk4mfi2cao6gYiZSP2dR0udSPLEDqyrYU7iWtgwIrSD3hyKgvJru81idOkPq3
pmGp/O3IRfJMyOsbcxjPabFvM4zym3ds4jCrMsFyUncL0OfiIfrjTG1BvpR1x6vU/5gAGofMSkxy
xBKg0A5WsLQGqrtjYMNDbV+aAgyZjstpqZ4WqvXDD96s5pZkoOzQepnO2Yi81QoyFPDNyagdvs5K
DlTuR853K9OTqEjOJi8pDhTreXwRSAULmX9n2wNGXNSoY08OquERBegoCFlV/155e8nYCT0pHLXy
2SakS8GQfG5eovH4iaskWp4SxltksvjpvwpLTYa6vvkLmWx+G3yGwbtUEbPNvmaYFED/i2Boq1c1
Fm1hEP8kNHhDAKLFQ3JPpq1m2tA1emlMIpWJT5fE97AeF4qEARJBYF4aFowzqSwKJF7GRo57AnH2
7WySX6wa944EHsXEneOuqWIhtqNhYPs28Y3v1coBKTr+xSu60UvoGbLpUqaPG4DgkUr7xmyll67H
v+WiP6ddyeoTsC/bN3BATsahlbuNo2jkvacQBEwE4y8gVxvmVtnJ4gEKz5Gn4eUE3ukoZ+VgpMG1
UEW0cv9daKJv+BnMjHjTk3veDUoTVN30iXKRvuDkwX9eINF8IEBLdjrvsTG5AFP60ANgF3yJSSeX
46pYBsr+pKrGrAVhqX1eWjlbHj7m9+2jvOJgpDBos7x3pWUUbqv6Wl3U+EsxiZDL+T378TLlni9q
ZKHjK3EOjIhRuqOnEwXZb3hwRQe+wnLP7uGoujI2TPVFR0DTD4Jzd3TcTmG2P+BXoN35apNMKFux
dbhBe7u8kx2bRuwvKTOZAZA0z1WMKeZj75HMH9az2P80T2Fu77UE0Q5YA/hWoM0gF5WGhj5qREcR
kyh8nDmJi2BFvTUkNMG4JiSuhCS9539UvvrPI3K8wlh+ngMhM5A5kRfQ35bwuJOgd7pPkf1twlJs
savctUxdKNd5U9BIXpHHqJU0W5h1UzBhzEuulmnuMaWf/R7HHHA5Nl1ycdJuEvmG3GpsVYpT2k+d
kI1OBoCoKxVf2oiM3TSksZpawYYK0HbKMl0T9HnffMYRlcgFMB4iqw6T1vKyiinm2Scm5t2VgHzK
K4Yhe3fmKvXB6vpSX5ofyNFQHKDBEBEpfOniwI+czz1boSU1qthSLz22FQgOdR+N6oLKsexIXvZY
3qmuaDb6s7o2OnlSvt3unE2O94d6bbE8EVn+GJlEU1A9PXnkEBu6k1sJPwO+FMZ3hveTAZaLSbzY
wa9K8q5lVLX70RFca5DqR0k3v+vIVzlLbJ/XS+7Y1ER6UIj871Mav2WW2nXwcoXuYbko/uY62qF5
b5mjOoVGR33k7TzHd7exJUpyEIAA7S09CKG8H6RB3zEoR7TlD9UrG3RxtyXzfq7v33btzmQIG0Nx
dh6Vz5QfAsVE5F78T8oLgDqSZtkBz7ddlO9GcfIB8SfztgL/agKDZlmurtZ4ugWCwxlIjrWzKesX
g/mdcjEPFOWyKbDNbgwErJ0IYLLZFFtqwnbFLc9st9DihS9AiT44IRPebypY7yxv0kL2pHVVF8O5
iLJecEHf3Fn/sUiXLwafHWv3dKlZyojhPFWMML2laXRkGU2vzAVZPVd2OxidcJIdxeGebk4tfdJT
pejKshYgLlNQcAUi02LgVFMsBzY6D3M81JRgcTjcaAKo1uuqA4jzX9FIXt6a2Bxt1HRcOwzDh+R6
nEdwlr5+ONmfOK8DI+0Nd/uS+URbw1YzDKFrlCqWZAIbNqbc0gE59yqDq3agfyA8CQqTYylMzMFz
9mnnG7Zlk0XFF6Lf8Ec5rTkUiPpY5vDv3ozIMTy8hMWkSwB6V3bm0b242YrJiIfw7y6qFbWNo6ea
hGVQnSPM8/ZnjKvclykwFxhKNY8OZgbb7rhOGznac2K8Me8ZdDdmHUKhDTc8M7QDBSgn5f0DePLU
HUUb6a4hBYEk8w6t8zJ3hcPcBHyYsxHnub9Rk2gX6CvxbLlVRgbjaB1dqhXCQuRNQFlWL1O8EmkW
rkF8pSTpgu6y1LtsIqk8NzpdH+6lgGO1GI3S+aVeElkc5uU3SBAV15Z0RBpnBf3M9d2U/Q3faDCU
Ba11RFmgG+c2v3fD1Rcmkm2aQ6NWpDk2efYt7pmySbSTEKdlN/IvSCX/UUCtnRf4V2NMdEyXFCIe
ww11LveNUItGl+vXAYY6u61W3wmkz/VptssbT/1ReJllN8T1cylrWsPDHsUI4F+KUtfHKMbPytXA
CzQlXXVMxVziqe/JdOUEvjVBAfcll8hFMqvczACqs39qRk3kIgdRtVwDYKsrZDIpytIg05SbL0uG
pabam8mB0Dw4GjlXCK99gWPJ1O5I+5FrXZx/G246yP384PAfHBZ1pMEK+kAAijZHl56QTMgqaXwJ
6bMC2eo9uGKbf0PLO9jx5HwehG/6GOiF3r1wsrClmTKC+Wo5vTC2M3NqgB47gw7I3wMEOL8RkXeI
ElzwJ3BPFJtiElCk+qnk5kp/C/EZ0ddOtZZpUuoUZTu7+VH+7NuE1+J4VCi9PynVsnI1553iwE/r
Pjt49PbBPrPK3OUFqo+QxHuE2uUfeGtwzyZo7YAuD9m59ipzTywQRLp7DMzcxFiuKwvRqnRMR12E
0sEjuUDSKJg1evCa55Sh741hBQZYQ4+xru5JUYIa3GOgOOWB1i7BaWpX/k8OLZ01Am5wHHjcneXd
+aOBwXXbtkalUGLYIyFUTZeIKURJhE37wFPFhx6gJ+xI3KsIFGbJOfEF/4rsxX6Ab8W9TbMlw7aA
lp/yNWwZOPDvZ47+lYGbsNmOZOtDp2/9NCqLNzHnBQKvYziAG6/eY6rJJdE11ldGXa78bK2P0Sex
tXlJqzP680nmT4DIRqf6SiBqYKGLNvN0D4DNoiPlas3gchvzY9k3vG1bTg9JBeYEE/6DQAsWcoc5
x79sl3AhA0Iam2TeLpHBBxxt7l/PoOP54+3jmOU2fIqvSOihjsBqo1xE9CW+OYMj68hWUPxqWomc
W6YTCiTITBfFw9M04OPNgr/5DGCfEQJY6Lfn6mNiUSR4KEAWpTp+DXnJAJElGNuN4P7w4oiklgK+
Ity5LjpwdfkgT9a1IQ+6g6MjZQm+63esrRta2Th5rSCKkGDngA0/Il9aVp9aYT+5nevoCAx/WEp2
Z4LKjg7Zy7Jin3OTJzWWde3EKLZLvH57XyyXCn6vJQLa23ZNg/h9VP2Vk99VlpyPLBJvnvCHabSg
wIII1r6DsJQ9CpLQOBUsUIH+WchUv+GT42KupTOoMVSYtj1naW51w702fDdHqRuSlrtPMsuiGQEA
7kHWuwlq4H3sxMsAVEPj+/huU/HNb071lwoa9x1Rkxw78SVSqUhwtHkhrboAg6Qi2c//QIS3xDJL
uFuTwMb1Jwtfw2d5nTUbKRdPvCPt66zAr9jKiqBu6EUhBdLE0EBc8gCHIuQmsQ78VoT4/QVkKO2m
bsk5tZ6NLcFiocxZixuv/HHxartujo3RgkK1Rsb1l1GoTQVcllMBh8oYtVxx9bcntoaD4YY7A5J7
qBAKavjpOc6YU0c0qF6xYLkX60iwR/1dqlGiROBhdCD8a2dT5jJ94/5qIDBJLsn9rT1PrGeK5o0k
My8Tr9m+IZ9FiqBxnuQ1nlGdjEOgtPJUfcHeAz7rMrRkk5cO6IKe5VUq4510rM4k1smswFLd+wQt
K+O934SNgWX7z9/xySpjMwfkYzvvmz7m0+Re2c0JGuYtAvRzrTMf16lryfyUfWS+C5A7vKegPIUu
FtXNT/Xj+KtW/vGoo94/BBRbnUXunjrNBazvBLvb+WyqXM5+NiihwEXM3y8iN/J7LL2D6+PvDbPj
BilB/BI707I8cgOkASu9Zzs+baXXausiVjPNFTkOxw4JA12cKsOeSG4mNfHPymD1IegGwLyZxEEo
DK77OcjVDrMDUJeSDIwWOnrG7pdBStdzX0OWeyUdppGzOMA5IVirkpODPK4ATYAzwyZ+kNz8WzKK
0H+mHt3//oUzhsRnRr2GhXS5vy/bOwwGtSjD8+eecNShZFdTNtBTgMS2cfRz/LZPQnT5U0rDYf74
6PV7zAWMfV/takImv4vhwPc9R0jOqyR3gIOdBZKLRlrBph47beV9TpvbLC8Vh9QzGi6xLVTg/kgP
J4luQBUdKdbYCIBFpn0OKTVvk22ifEioowcFRnaEOwyWFJlFz4ra4QUNRC7B1mtqpe8+7Zq7sRc+
vZa2sbVo6A0/pMkiuNy8hpKQNboNg4YwgXzamYBnXboNmU86dIZ4jh0jcO3F7pI4c5EtUdCoS7e8
F6jALh1YBSQ0r5WFqZAlZAkYuShZJL+xkm621M8smwz+2rFovgA+SmmPZq8HXNlkEyhGKFnaeNZ2
+1xRWoz3FiJrkiMmuj8tXt9QPlq9UhxN8DcObkAtI/20yQKK3ewerbiVeRHAw2SAX6z+p8Gas5iF
JR+Ew8cLX02c0bvcFRU2EO3Cam9kehRIXjem51KOOyE4QAG8oNz5kSUiIv+WTcELzSXbUtPTMnFA
ANSWuEYZVa8l42dMv1AyXJK4gT5QSifRI7/jWBh+npmfKGliJQjNcw1woiD3X3wOWitys5k2kGdM
Yir8fI2R2qASB8QBGNEvFtrwQS91B2a0oLI0Q94BFOTY9K3UxioEXsAyKQoc5WpU6+afyxMhpeB7
kbfrMZQgDLjNOt1pJ6Qd7kOI4NlqvFwTBWemtQwJCoiIsiGOiMpnN3Asy8Au0UskA4/3VTMFGqDT
7mm+trQaS6aQfLhdae/vt2/jhnHK/hOh6hJ4BqKLWSHP6sSxxTCrey/iss4e3Klk6YWmUBYMGpMQ
fhVeBQAgu8OMiEg29sr71NYUsBNwEP4iOHC0dEAf8mqaE4Ehn4ue+i1WDMGweBkDdNyV7QpPi1LZ
2dCutHbCpd0DzE0IDWARPZxhig2CzDx8JkV+7zbgqm1hU8C72vxrbyuz7MVVqX3IM0AJIaByDZh2
Vpx1YK1dDVFZS9DqrAuakpHbPRUodpUVzCcedJRm4Y4NQGAxQJXD0zQAY01/SK7LQbAa87qkHlwU
5iCDCG7TdeIkdDL4X9l9XxicdOCUjKrCp3F7byOHjc98bo+/AYuTn98YG+idalEFMatMlElQXGXU
QuAggE2T2LPkYWFBfbu6tAYweCeGxlPvv7AjG53FhgMq5a20SIRkrnGlv2HXGNvNpsxeIV1qRU5K
3ZHreth5EpwEsNNXxr9fEqCKz1+uJC4NVj4o/EcBwo3l7mp6KZ+LeL1Aa1h+3+oGI1fIOwkaPYgB
sklLsDT7u4R0HU9mLD7EYP04HuNOvTY83o9WNcZXoNCmLZlPbSl8CsXVgmUqbVN++ppNaMUhZMHt
uOkfbd8GDiG2x/lr4sI69puxmXEGSF3l5S2mTQpCfdZz3QCEJ1kM4Oc0t+yRkFqkZV1Z+aD+HoMC
wHPlkE5Hc5WzaL9LW3uiOZy6rj/dL+6JOBWeH3WRKolZstpxhP+372TOvzfXUHztgL3NtxZrMqut
gbWR9JH9BCUTjdnZam+NxeiVC8UTagfU34EwXFoHExpjzkYUa7R7hHZ08/IyQdiPT4Ugi0BMlliy
Eta3CuX2D34j3MbaZdSZzeWYfs+sE2Dvg5AAR8FVTLc/mwfSZzYKENaPEHf6C1rmXtQrpV6BqCgB
f2l2TMg6XawPSaJrA6OK7OWOXDI7pnCPWKQQBpmHlMdVBzDKm7ksxwSdMAdXM7RD4jbRbzG4Wf4x
Y63D71csUifnWZiwXxfdbj0/wXfm8g6g6uYfIDc4a9Xx7aAyYDbR0w9VxsFheXq69AFJTA0U8NJx
BJqRDhsgrNmg4r55fOy5zStnD7h0hg60i3zArX9LYlFqm1AvufsKmqir7fdCQHuRehCSJIEUNmDP
IeKrZLbqTsyobRJKld3HqZD7dOXEi3cUp6/J0RazM7ZsbFweuDIu+9rUtYhbRQMCFJSkpLHGUP9D
7lBnMx9AMk8NCcWQh6RcOoPP6Q/ySpLa4uL0gHboeCVyz2OnTx4qDZleqOrJNJUTbZ1RHfxy60xE
kEBRMZOJoLPSGX4bjDOe7VVGiEPtkPifeg4ah4IxQrCPrYKJgknoUutf+tb10E3sQWZWD0LQvQmi
tvr2dSlzf9smwc6ffdUi+4HOqiMphw7mKkL4p4SNDCkbilcXYtjl85sG6TDf6Mgv5ap9cEJiXd6+
WxhFhNIRp7uNu7SznUTWb3qechFBu3A020AgVHL3DGN85Dd/Siqmfw/as5dFEhIRYUrw7W+/saib
MvNwOL2MG5Q+lLXJlhKh5khDu/yTDauI2Ty8h89+GfKl7U3eeoa7yJa8EvF/h5Zm/Kl4VYXPfhPP
OrPxQtnXMRjGslgJO9calV0AlvRvQa2UejFLpKkW8ND0TdiUaK9Ceop2pBG8dtmllSXHjgUnIuGS
tZbIFisnRQfV1kOF6mfsq5veEhmKYl/70QSMkIBfPfmUGKDlb9Om8xpTuxobRFcPWFi1nZzk2BXi
M7Z2/xXVno4+pb4sPFs43ZAlMv9IFDJZOEKpSEuMjf68z4vwvhOHdya1EqGxESujnBl1gyf7crtv
gtGukGBYmmJdGyPzMbqeJvJyANjKhtjR5LCjvBht5pp82TYgQBnUXFENtPidjBKPgnpsL8SvPQ4B
kRle1ZfdBOeGMZoqOVPVXo4uyrcacUK26wprTfa3KHauabytx2GhO2Z8OgzOdk1QCBrr9O6wfaTC
VU5rXODFwnM7IfwGg8uEuMXF5CC3HXNs1bWu4Xull0uIkfF7w5KwlAz4Dnqw8Y7jnTahwUgzzQN3
kJ8AosXYEygHHL33h8KuXj34BRbilTvdnvGc7DOEG7tdvJOCA4C+eR0QN1SAgsl74xWWfd6uEPSE
UwX1V5SuC6YZVcFc0sxn6ibA2Md9NOWtT/wLbz0EkV8Ta9OfW7hp0xun+7tltvl8da//8E6C7uto
9iB5hlzDqrVBxRlIJtkSu4Rm6UEUEyHamfxL9grqdrA6aEL4IHcj2JSGCymybB1y7nGtiN09pDh8
dRgLaRvYSKL0xXhozRj56/50EiGFAwhWXqqXiteSOEc2PC5k878VKo/ex4DjxiPguGsOHo9SJK6z
IaO7e7HtAY4e32oUXAkXm1WsKZ2dQy884Bbpl8fMAYyVYZtf+2siPDvg0W8MGJ1clboP1HCXbAEE
lQOj6+rBPa/RYFSmnCsNQplf6x0PA5NVx6aDkBQPm/VfJr+qkEwlui8ZORpHZUuF2E0ksVZbzxoW
RmRzDGMMvx91dJKFt9kchuw7BxD3jG6ueK7mqzcXoMLbFWtZEecAt9/VlLsfNz/yF0EuyrVdoAl8
L1qqFUhCZwxe8W6jhL9zh9imPZ0vw0aEcjVFlMwRJNOSsLVxnNa95xxrIIg6pv59X/uVeHOYeP+E
S2NQyRxF+WJKscFNMufZaTHWqodediNjoAaMvRRFpDkIJhwOhzV00CKyrtiCPBt/QKC5xGBtrzZB
UyTCPYcdZLQERUPCbaFnUMGUTCMArvjpdyrPM+OID1tVKsbvg80BUepOgDc/e7HZXuRdB/5yKsBY
vURdz9e307UYuWyZhKq6l/vcrwhFdIcE41PUAZzmOy3XAmvCWnJOHm1g55/bkOuEs/IV7n6oTr21
OIBDTDl8UjypTtZIl0ljEt3wHCJ/2Qt5I3zifYlDAnpMWDShmBGkJFSHtKp7HaJrFaPKiqfcHuMI
+M41H/fYivDRatQPP+neCaVFzISZ7LCTK/bobTgiCSOyAS7ZkmBpe+mSMV5wm7YqNkVzexqYoxi2
N21l6x+Q+205T9jtSaHICxlhfsE+ceSY0vjFlEUDYkBYU/bLRjXhDGnOAGeyQi01Iv5Qh55pIdWT
EHkut05Z5Owu4D0Z3fawlR7G1fIFOCnLMLIGZ88w8+r8LAWg5yQNzs+VZp4mFkBrHip7qz8vq9Ad
YN/XqlpUz3C99zMFvk7LEwXrAHUjH+53FxAUX7BsGsgM1uJQE+EvqHDAtLYpOMp8+OBiqiJgOXvx
3PTl7qN67knnHiApypltYHgW+RAPH/FumT95HY5N3XNWorfpPtZiEkwKriLcthpZiM8eb7jfcsp6
8AeFbwlHjwAZfB82WMnwH8YyJIXN6kzf3CtsCSkUmqKOH78YGxLUIhSq3CHhRrSoZWb2658VrNCA
2L8MiBJJ2h4j+bQSe2gSYxXZBEUrCn7YBICgRPEm0Zi4XRzQSbLQkxoHTf0mXt57wd60hHYW6ixL
tdAilE9Hh4wSyixeOxG/9rNYi7qrb2pFG9CyL7QcrX/4ZDVFLTRpEhf4fct0R3zpD02a1nJOI0L/
Dgq7mc6F80GASO8ssiiZemlCQRM2TqTPfqcFxzfUJqV9S8kP8ta4hneAfWPLrqHLFY9KMXMvynRY
E4vijW3HnwgUeuj5bYZCmXvxPsOZQKBhjBoGrKBHX2CRKun8+oWczLJiuuW6mPfVk3kl1evznuPn
QL7TzOqfYeEYl3Hm6+7W6Y5EiKjR09EaRB6r9sVRha2I5i3vJsAVaWHinFmsq1BrkiXs+F5l6Qey
1z6LNDdRvAVmJQM/hApUGgWtaefndzLU8qwd928RPgTTWR9yRrwSast6oJJZFBjhu/yS6XuGYrAa
ehZkzBcLuAdzCh1684L6ED/aZz1ExC22zuRMsLMKBZTy0Wx5pXH1y8n6nUJkq4zPmfb+z0hDUg6X
8GLuGNfcwsL2AQw3scacurfuzi85KoJqE4riMBJxGVZk4nl56ty8LtFyYB523V0lvaliYuY+0s33
WB9SfgnaO/eRJPe4oHGhzMnvJMuTv5cak1YAtXwilBqI7ULLG/Xo4pxlB7qRXrcTwkD9+WP2lQXL
83+oxDI47J6SZIfGv3TLiL5UF3uIab8B/G1quPoEmoE5x99MJneENbzm+N8GPnfY9k1vklEXrSBo
SmMitn2aPpOU7s0sf+aw4ZKB2j9DmskPKarocuoKzCmj9KbDZJMft7+/fsxC/3FMqtGj4rfrn+wL
hpPckXSEaU3PpAfSMt7r9qoi5ia02nMEknFHo+0tU5N+PgmEjFtXuabPgJ0bJjfOwB9wMUjyD361
IdJTWQgqma9GeMJhmilELVx5eS8lWTPKlWHKb5TuY4MHUSBc3JHdQQDzJa2pI87E+F3V0aljdjMg
v2P5/M13uF0gwsflFT/pgx2Yw/A2beCyljY/4kBdTYZ39597TOIKKMMHt6oLJs4r4kWq0sKtPiuL
qT9Up1Gx98QtDkUy079b5kZ9zA2VcPG8WILUHyK6RAjsfAzl+XLA4UjAV88K2/bDOx/9wbz1iIWQ
FdF96B2+76rSid9HTA3aaTkKhSIZbz/wft91nshzj/5csvUAEtxWOZ2hy6q2CM7pIyGHVjO+FyCX
xunfD+q5kr60QaruyYJhGJdMu9gcezmykTid8SXLLPLxzT6uJs1daYZsngJ1yd11hR5/6l+qUZh3
HUHKWcvjwV0y8oD+3+FENsPapSpUbztAtH4fh56ZMzCeOZfuG7QaZrutesUHEATwv+YXhdcIXkZA
893mY/g+wesGBvQiBcEkyJTdWyJzbCPO9ed83arwjabkysS2cA7rsj1jWOS5cUONBl1tHuWYTz4r
ZjpuF0Poe2drbQmyZBISSbnNnUOtm95iolJw+kiHfAobLWfT2RUITH2qiX9RVwe3kjVUDnSdjD3c
Qgt3df1ugYJ8/mkg2gDK4JCLwQan75WPiF4gWAxHAEYX3xns384UnmvI69cEQcYN8Gpv+bLlVlzh
LasziRcI8SlAghRArRd0q73xa7uvMbWbyqZh/EY/LFAGiD7VOQdd2NoBtBXB0PzTKkxaMXAkY2TY
v/w+A2cS5RfQJ83cCmlPjP0w4nGkGx4hbSAtDRpjbm0VFXS+FxE4M+gWX78a5ky4GIs1BwsneI8y
Fk9VfdEbu3JFaDNs0wV2FTS1YMOc314MqfQajX5j1kIvcHZVjwkVQEOhFr8SKRrhcEq8Q7/K9SCF
3UvJ7+MgrQuCTNR6ZLPj/BHr7agD07AeO9tm4XwVPFwQ/OHYbBrbVRQaVH31JhIMSKhads65IriL
iciHj1Zgul9ognZ4rCXBcCHzkpc3314mrpDOcxOYGfy+1AU9a1e4GyV3YYhV+wYWpi3E7F51KQtR
/qvEDEsEAfQPplQ2gLXYBDUKcym+rEg4cwEn3OmZ6Rz4cVBGONUdFpdhHvr7IhtV0ra7SGm9itA3
PqLwrs5N8bRCba6GrufTjxYCU3DjC38D+XaDelxGqs6MbzeTreDylW1ONybhnNCEZsmiXM61OvlX
j7j9f9Mia3eB1CLc41zBS/4kkbBm0cC1hpwGHZk1sUSfe719rLizBduIPtz3h0DOYwu61O8ZE6Si
TcvGEsTtvl5+2EZhca0kGJ/fksmgo8ZjNYpmeM8XAMvi5cmRskwY8bSMVLu58cUfgQ3uniylbe04
eo9NaNHeU2/0GrIJvmEDIIlemxqNM5BgNP9kfnLDBKpRONjRuhMSqODnvmK6I5ypsHb8YMnR//qD
WPilw51YytxTQ0qmHFb4vSRg4fmrgimE13nbNKTv4JgPMZmKaXS7PideMfLAQOBiZLuao9xLXRKK
+CIKSFkESb5bu0PEb/9ibYmtikiAf4TbkgWpti9mkC16/5KcAJuNCRlM5hL9DO22csUUAa2B+Vqx
kHvooZ/8MS0HK5Y4JenhXcruCF4oEAPI3f0abqKzTwlWdkzcobiqkkb3qPkakvE0GvPcdlB/Thmf
sK5dDPVJ5uI9MboIArVAPaizTH//v7PsppNwHgxxpS36LOHHw75hxXof4hy+pgDRR2r0PVF6dp7I
yqS72W4feGKY6SEEGyDsr8BX+OOHfSfxpd0ZYvs3dQbrIPr6C/AMLrsHKGLJi6XfaXmO1jbfxcKP
7ZOK7qsb+lX8UKEjI9E2M616WizXeR9RQW4Vj0FvRPhsuogHXhBK1IIUfgxQghtfkNpw7f6E/Wp4
VjZvp0XPtWEKF3SdsoAg6G/Sv4V5Y4cPXOF/jL9AzA+neGonZUexcXTLDs2m7UfsP+Y3k3O2Wz3S
dmsyIpZV13TSv2PjUcTvcC+1rmWgdQ1kj/70LKt54PjVTtpSY4AChrXBj8p/Sou4JefIceZu6nbk
JnIRBpJGS/EKMbdRM3potTpYyG6yEI/qi98n33zMTWefaYW7kEJAIgIAQvGv9oUfdqnbmlQ6j2NO
NnvQ/NMJMdQd9rYPtqkCo9G/Qu7dTHEOzqoVaSPpAAMxz6PXwZBN4ldzkfU3gyaCdanVOWirUS44
+Yx5r03XcFVllk+5+/Y3m5IThwM61baC+w82avvGrG3BWha2k9HJ7nXmiREHajCusbPlXFjbNKZV
8V83SgDN/AtGKVw8rkQV5jQkH/H1m026ZMwnM4VVK0eJPEpcic3n58fpav99u/BTCu7LBqVTRSbS
lo3Vxc2sG8dQFLMKOlos9vqYx78slRoxMK0eZ/5+f2tQr3Ehc9nzsyaNvQCHm4Kp8/hhXnCFSpzc
TntMXWdsgZlAXPxjLxEPivoOJLmk1iijn3g7nIcB679KoZVSoamN7JMAEyWo6hHt+8GaTiKrgMGR
2/Waek21iJtiylvDJFoNnGtXPFiE5BCwW6xv/HVAyOCVgGfTRcH7bRpeb4nsI+UbCzL8CTtwA4yi
eiKamtW7mxRg3ozyZVTd1bgPAcyUwZ7x/+upFdD2dLQJfCi7MIziPGpxkoE8JmM1uJYKGTrn+9pH
s0zthtR+/ce2pXaIwrjCHxh5T1ev3GuYsXaQ3nr5xzpe+Vqu6dSgCSMSjKtix/yo1+6fM2WgaOOp
XTIgsfunX2M5GKMkqqpSvabg5PkIDJXaLM6OOU2pP+3mzz2hL6plMh2wUJC4ZthvM3OuJiVV2ZO2
TmHcdBFjVZ1NPt79n/FS0j4pFM5Jx8CXlwpKE1Vw2FXBhwTTXfrkHmPSpiuV8YXa6tNCaZw1UhoV
/Pu13SoXxrtYDeW0e7aSheTydi+F/xBYiL/7ygAp8h8k6AczUAa/mppqPl+5orz5aJL+yffDHYDR
AheRMnt/WX9N/9JUrv4WXq9tcjSP+Vpm12MeDbqDxK5qN8m+jB61mNh4zkj5q7MHu8IDXqj628Ke
vUiEQ0/zuuvJWga1j8s2sfGflfq5GaKDxK/8VzWQDMRcCdPVjG+S16v6ippbWnrhRieUAdgb79+F
PMtnTSqMp7v/rhU78QEGpCCdiEfPMmC3ZBkhsUK2qpa+ZpYUhM9S2aBd/MMsvMX8ZkswT//yd6Eu
EXUTD43sJ+mgFHn0OFE55O2KxVmFxz5CG+PmALd/nZoHsf5KSXPAKHPx+mRTSY255S9qvORoseJX
JIDSsiAyvs7PUWSM/S8TZrmLKq8eaOK3MKGw8sgcCn4Uv6OA0ulwqjiWWkOgRABBZWBzrz3uYKYY
noqy7YzE65y1VmgO1vWme0/M1whu3nRQXpfvFP/Fup/nsSnp9zpsepgLvNqWDYuzBswjUUEpqjZZ
tGkuwMJp4Taux3zPwf9Ogg+WSP6/8NqTlkI4CGc3cs/Fo6HDhCqXt72tXEIRSIfNLpqZO7QN8KQA
Sxa35jwIKRTwVFyOD1FAfsGugcqYh6109+aRa2+StrT12NamFkzFIrsMIeHf1bFavq7bAETJiKyh
y4wif31URnjpqa7yl30vTA0Z0J3QWw6JfTD2fEROgKTLBjbQnnp76PYP1USX8JOhKArV0qCqa8Dl
j5nN63y/UtU28J/PZdWGgcgBcXnHzeeHJoy5egL9p2//0XJdKT9t4Us16K+tMc01St4fgimrAEtD
JmzCSLd3hreH9leR6LdXeaqEgCm0Fc0hRtoNO1qy2qv9gJyifpiapvXqqgm2LEA/Snwa4CFg13EU
KV1zluCZimi9evvAO0pSfPtJiu4TDhG2yR/998EWukoTGtlBSZifPBgmPeyX3MrsF0CsM8cbDJW1
2gjLYUI2LfDIl4F2yvur6CtkXI92+HLCJ9HQSx3p8MGuMx2BE2zpAGgHyiajc4zlDmRBVtrt1/+m
ayPk1n+OpS710vC4S3tXMip4DTUESgGhmOV8XoOVBI2GvC3gd7Z3O/Z6Xm0VXfKkccnLjOUVbENa
A4S6imalhMVdu9OnYbiCEvFcyJpxJn7u5IB0sT/GE9hkdkRbUYZ7YI606QefauXjioT7J4x9pyld
ucXfNXelKPmCZGqn9oBuT+pKB3z7f45nLsx85xlmCrWw4gHmWMpn0RRiWdX3HnQWaYmwmTEgstCe
//z8Btl6WwTYEjMJ4QULHPT9n/W8Gsprrh6Kb6XcHFnbVMVccT2YVrES3F6NZ/L1eJax2hZEJKbk
58ei1jLjJppscxMzEwrBCPzdUiWhtuTlsv/NB3kPPffEUw2xJZu/BEeW2AzuTqHTpFHqpMqsxNPy
7kzNhEVRsWXdKblwG1A+EephUWizX4FOce09jzjdGtAPmIthKwMsXpgnWHO5jIO+5PejR1F9+p6I
EKzgItphZBjRzYzEAm7LrS0cbzRziId1bq7t/UtKpybvdMwbShqoV86zPLgqr93vC/sJLk1kZTXD
ebUCwKfPGr1e2N3PnjH85o+6Vqwo1hL1QuINbDvPxyX8OYilAPN3eT/DERxXHYIUS/0Epl4nmu6s
v/+qVuK6TR9LkSgUwWZAFWwdSo0wrIFX+zZU9t7Tqijl8Ov3wgPolBxqCgNiFbTz/PsscUe3WVLU
nwIH9vUm53Yp4qgCLarwq2ASPxCsyCe2yIhPge+5isUbofxFU2h33MKZdC2CpEzW2V6NxCgorzGn
/O13VU6MuqyAIRPakxZop8J/UljgWy9WEsnLTD+Xe3hTtIsc1lcSDU29RfUGNKBE/mZvhXZ5ssef
q+bm2oE1Nn56jdf3D9WHBR/KkLHZcqIoZn57w5d6Dm9a4wVRefqwIiiG53e6efC1aqZOiseGKf2Y
0mfKZBHsnonD+bavgWme523ndYiOP72fYx4X/l4MdEzGBzSxg/iUUkWmeLTnbtVBHanxyYptsZ2+
0g8i/YOD+K1TdlgwuQloroXPoiirKLGF45DKCuk2y2Nj8Q+H8E9SNUVislyoMbE60U/y4G9vAlyT
E6fLbIgar7syErydZfasKUJwKTFANc/vl2CgCFjw6Sbr4xp9RAykA9nwKlIrwVAFRolPksp1FS7G
p3FITxNHIIs81Q8ZDphE37xwVwvXJuw9mj/sVwddo9gdkactSx6BXDolTWrVlTNh9Qj5bz8FUBYB
wK5TYgohzR0KKWdk+2wgDKKiSpAo/ar4VpXrRjMhC06TuUNDa2GgToz14Z2eho6v1+JV/KzHIwYw
KTfBx3fEozXXgQP7OY4u0yeuKjP+v9hBsp/TRi9BFO+OLf/gb/9kT0DGOdAQMHsR4dqMAedpQjiK
Y27JDuGLAS8rp84PbNN+rz2PH++IlfX0OiOzM1gVOJnUR2jSTcapBxhmh7PxX4xZMqJVxR3Ga5m5
uq/tiZPXuePYW9k4I+UNCUn1v6bF+71pYUydzfeoA1EqbcRMbvUMDYraeZfmrT8u9Jovl/fk5N/1
fezkc72xiD88GXfKDfFOYbUsrWO+MWDrIkHVwRP+1SN86YIa0yt1Sor1j70MvCIXrmemkVX+crug
ZCBlZylbJcods+AeDoiIed961cVT7aqm5YErzoWWkpAoPo/TzHu5t4RPLL9WnTjwO+B3CRRanX/B
Adu1AHqPw9BmM0ZJYG64hDtMRub+2TcDcP2yW5xX0Ju7veNZO7FHf63jgQWpr5ZWMJ1UlI0uUV2j
3bc0xAtcqZRFj0YWi1EgXG+/e6EIY6LY0kfudEXNG9E1EyakuQ7254NObZizsRIERT14Nv2JgG5P
2rO4eDHjoXM/V7mfE/mKYxVv1QvwxIyadOqSsxLZCAphU4WiM5AiWUHp45sU2lTtH+erGTfqBEyC
EILYQFj2EybiVyPuZ8+xWUrphQ4VbehEYIZ7k9lpalblZm2UGdD7IQf/YU8in2eNMRWLPe2T3YmT
PNlsn/vshXMpRkOpA+eqRcAn7Jzn+x0Ha2mEt4GGwnHLbryj5fiAyab6i4QZuTsjadQrRjACS2yX
494E73EvCLzvKoA5xAImcJMWdvro7n77IDqK8PsIlhZKcyh91QSExO4p6jRPL8faoK28Y9rK85iI
TgVsTNDjea+eEafTInYXT5WaaneKG7e2h/IkQtAZelXMcy6VQz9Bvt0bUEthPIUegTjHV4oZ6PR+
IrjK+a8hCr3TbqPZ3YN4wb0LOp5u9R3hjcJWlIz8FuqpeCxpea71E6TUSWfYKnGmOe2bUfJl/f3B
Rr+xXAeNO4DAxiPUSxIEu6jF7GeCfz+v5a02a7JV4SoOCfEEyGs3HRlr9R+D+j5ivEWzbKMDEsin
TnArMJQTiePyEXXPDNksPrpws0BfvctX17q/+T55yW49D6OIZjFxUTT6qL5LaM486dzQg/ZurVrL
z92Uatl3K7Y65WiC50ILEecXn2gHf4xZO9h4Coj5dnLMgX6cFM6GReQrAg4pXQDaxSThWASdImRd
IDeplTNH0M6yvn9zMt9arh33+DEMd2JOpMLVxOhSMuZ67czvBIzFx6L6rVM45iSv1URxQ2sYbxGz
jyYnZOdNkLqTA9utyKK3fEKsLJu5RCUAXKoFRypEsRRWpR7JjwhnrQUfGLMeQ21er+MAyzG+L/uP
JW3HxtdqgONAg1oCZpewV35le973GANAgwev928w0wbYeuJ6uJEQfXpIETyfnfSr34MlR8yRJYdy
GxRxgwbRIcZ+4lNTiXZXJbwjvXAW22FXCELDA77agOkRrZ6RZniL9RX3xdM/tSW8Netf2gsf8H5O
m7+XOz9BzodtoqPD9MKGkHJJPkEr9IcMBQlwBTXHhBm8bDsmuIRExGZMCiVwP9PH+s6aNf5gW0ZH
NME1ZmIpT9OxripjChish5OedOKm/PPcrMqT87qY9fZ66aM/UyPuntMESZXBDbhdurfmcBXw/D2d
H06deudI9eaVb8XAV++jOtNy8qCMMG8qGp4ffLkydyw9YH9Xoi6Vc2SqCzGbZxkhmzfh5CKPyFzf
djRVLH2/jhV3ShRXMAj5gvgP1yorNCpl9fJw+JsXUf6kpRB+UAHkyIdEic5P9LbY4PHDF72OuFPa
FAmhs5LVldi0fnxF0XBuJinszi8aefOaByG6jEWqBckt4IbhCkBXohvOQze9jbJhvq0MlbSVFCdd
8gD/aVhtAbpHpWeWVJDwzywiYlFrHh+TgfqwZH6nyheDQIpyw6BArzMc2iXjqtZW8SXL7Yja0D9i
zsy0clZuFAwmeMxxyPJFH/cF/sHyVGI+0//ZupIYUoFHNQagHCZ24lgtGpUj0yagKqH4RI280bYl
7iB9owmh7WXsZWc1w3ARwcGBtUSnck4+IHYTPUmAj7rme0bn2Q30uM21M1bzioNgR7jvrD35QQZ6
5f4MPxDQ8dIRSpHJtvVgCjPiODzBa97V8BhypJZJ564Y1lE2dfA1nU9XBXg9CHtjWyDt/JPWiAky
cNt9uA2KFVChc0e1jd+MHmkyKmJDXz6ny4sYn58Shoadr9bz8uQr0lppD09B79kaq18cc0bwIve2
HlKrK0Zi7Uwe4fJzKLV6DyWeA3nyTt+7YLLVau5QPwlq95kEDQ/i1XWx+mkY73ZeZX3MVTVM0pI9
ujpzhBHpk8MUJgXj7+A3U1WFWg3N4YlKkkY4lnR7JZWzmSEhr1jNJYKK3VxgnCFsXbN128uu3gr9
c5AIaEeCka+zVkRk3pRs/PnaGDZw9gmNzW5ZEKdLGZ76uCIb6nSbhtwg09NbAF37aAw+ZmltBxYU
TXpDlf8sR6YaKxJuAmCwf2O8d7PAZ9N4DNRlwRjnXyNDR7iS8Gyc3Bg27U6CAgHrVe+OQ7cs0Y1A
oZRDa9vqRf2AV9/BQvoc+pebgU5Zs9F78qV0H/nbR/2G7eQuQ81AD+njqh7wQ4amKBktueQixxcr
WP2mPinRP5ZpvAmOXRF51GwnBpwfrfC1SWKRjfyN0vY/VZtd7HhD5kBAkakxAqr7GVEsAuou5chb
A7QeMBbriJPAi6XUYHc4/HcAs0Nds2Sh0U8Qw6noBKoBcqYA593pQ+zIiQ3eY9HcQ6ulz3kYhdPc
QBO7fcst3N/VIaCjI2IUR9jwDeecEGbF9R9SQcfGPSxTCof3Sc79UbnTl558MQnT7UrhJq8uQyWL
qjQQ+NmyL96kOu9SY7MgeaNz71cUKU9Tmqsq9nD8ehSqYY6QsXi5NNWWH+lt75o+ZfDfaTHo3U8M
+bJw+4Ss7eLtMUSSXaO790twnvRjYo4o4mkhhRpFZsUgZDDUDEdtv0LTMZRqtxBbjJ0d/ELz9Nn8
KiXdFP9BT10WdelVmCp5rTbYPLZzGTOLEutvJDQH3MeJXqPpmkBrf8+OUjiaP0bLcjDCkEKq41Nq
sbZkZgbqqUcaoIe8gDau9NTy+Lo+niz2mJCndqhKI5e4mRtynFsmOOR6eWH52zbJxOLqI4xe2jT9
1YNNqB4eQkrNK49mRmn64G/mR7l8U8ZsYu15eJ/L+IMBRhEGhYAEsNVvJjI+l5jegPpPtbiUcB+N
3J1YThjxTVFqCyirdpmfefL3P2Gengxn+KGNcv902YQ6CJusPdaaTPLVG6a+C8RmX7xxjHJpLa1N
TWe+Yzf/ziNeAPVzKQ2rqFoF2qriSnuPYv4BTAWXBPPjhLevnV1R0Dm8uxmK+Q/6UZJxFg9PngbP
DhCc/8gmEFUspsmJQmkp8jXa0xOf0Vlk7CtkjW/DwtRZ4eaFAdP0uImdoUJzGiKKsBEZ/2aPli5S
td/C//8ZeyU0pOYMjYJjBI0eiQALWPJ9fYdARZhfHFdJafMjLTJKB11SBFclDxctC5OaUSXymHfb
TT0UoLFIigcBB8eZCo7kYJ9paLsK9uAQul6yh3Wnk3Y6O9i+Q4017WrcJMKlBm6zoMgOSmqMaoCT
BGThXX2ey57rSOxxAWQ4l3EUumOc5c96WEH/aeHV1dNF1NAvHRWtF3uVmx6L/UFX4GRiNwn5UaUP
8SWUydhLV/6jA5XJJzS8hsb458X4/Q0tLn9NxwIW/jJQL1HolgTuvXqZhoq5/dN5+sYF4NakLQmo
dcviZEGgvGsKjjaa/6jk+x7BAZ5PgRHbhcHnUvvVl6TRTHI9qqyCk4mP4ZVTTTkOZ3leqyUzso3y
Eu55o3HABMOiB/b+iurmd2GDE0Ytlv43B8nPDQNhoOYFbKjJtTWWHD8WWoXJSkgdhcfC7FZyBqyp
MUXaKuPPxCdFLVL4tLnI8wq4gsvXEpmTBkOPgXg2KlVmbCPbf8DR/YET1VPdXSEUVeBhbMV+8nT1
iUOUJr9CAY8ChnPW5XkDtMtmLSN8emOi2UWW1d9GzYwO2z4zhdVxWo4XWk30CqbaJlgr/CrPQN8L
cQG7PPhrlyX44IygSr9OTy85efJMDq1RGzZCuZJ0BS9WnF+wzFrqtO6avFSyOvExUEdzQxebX7ul
lZ4n8zw8YejaBl50eME5oVHnaskJ0cOrUxkR0lbfajBjfFWmtTj4C1LvO4YMw2Mo9PGyCJMD1sjs
MOZo86rVTzuJUU8dTYZOI69KUTg9iXRl16BjFc/4cy3LUnI0/6BD/St/FrOMZJC/mMCrI8cV1s9T
6dT0GRul4wZstSQ6IluJkwCwsLaNdB2HiXfT++QoFgBWcm7oYifb27VHvU3qjL7xKR4LwgQxtgOn
nQ5iqjtc5LctsMI9hpcG/2TR7h1gEywEnsvYh/AfWxY22YWdDKzU0uxlUfHQSbuy2eeuELjBbVRS
7MXqAf3YGLWxo/xyN+ih9pDzDBVvb+zKJ9snT+R0G69FLMRYvjq590jrK4Cx7cSs6mcKRjKsm6x2
gWmM4FP4qlhHOZ/aDvJkTvPR98BXgJDwB3YfO0voAO1Y2q6sKcGGwPNPZS5xOoKjCkQhJv6Bqqyz
oln5Xc085r85FGBCe/H5UEb0yDkzKl7KcxU2tdPoDmDV8FaUKySWdX5+YSGA8BdjpSk5nAE6Vc3G
/PpTRbZCEFTZSxGiwW/qTwH4ZQTqO3ST7smzx81RdvnwzwPe+APypTFhRZ0ctpDBLe8KkI90MDll
rNolGLPMZWvOeL1I1Wa4XiQtDghrtJOK57joIqiPwZb9OfPyOercic6MtWlsrJ1Jc0wjyj/bm9MQ
w35+5KWD9lXQClMNXazJlihDD/WD2msDCrRh7SElLaDAtZyjwGMvfT8D4Ez/QGHA3TpyXyZc37UA
ghInpkcVbzBn1ZkNl7QvX940nPVMGMk0n5P6O57MZDrfDq8nscJN96xIp24M1fjWMUdmJGyJPqAF
ufYTZ8kC4WwoND6l3Bix3C9LtsLpa8mGqa4AQ1wUAqDi8cRzAoQ+ToTGVgqq8jn7bZ+3ZBkOKeSg
AMOwnKmxizOSc/4ImT1hvmD1xygCuhLt78L9x1l1B10GT1locKX2jHUfkcGHtmrr0khtzJC+D+mm
aHHBSV90obu/RhCm5BjJ6giKpPHYmREbRSdaai0pWdRjnW3JU1yBaacQSOGOmzvr2KImBIrLyOIn
62CJAfX9G55tBVZX09Xw4Eikswvx44DvBQ1XVYZB8A206rxJxXUYvAwIxNqAN583Htu7zuZQYaEu
qunP9CQ4bncrJ/hTW+di5qSBjlUj3NIm3zlVto9+R2zp7ywmtYswe+xsAnUi6yJaezUn07Ue5EDm
rduZeZKHQ/oSETJHVymfkrRsGHt04a67qGWc4xq5+TJJ1Zk4Vq7P9U02TX1Gq+DxC6ftLGnX6gaY
p0999mMJtEFOfMSPaUh9aSPn/OBhTZbgoV8+Zy4fdzeN9s7xv+OYIeEJtS1Y32h04g8qlwiD8ucl
ePiz7XSkLDMNp7hG300jOEv43kID1u5jJ/v+MGJU91ASAKE+0o1c8WmNNBT0/PVNm2OzLqS+xGx5
IKN+3SbTmTPsMDRVbsDMs9FbJZBtpRb1xsregY/FsqlzJ/Stoofic3iWe7D6ObjW/xvqR03ZuqNV
QPCSUwFgH2PejST00+zsWOQgELK8Wx8dRA0V+YjMj6qd52X62QzLB/oObXz4I8TSujNRI864m0c2
ctYoKxk91lNtlfcbEy2VuRD71pfr5nY21EVdvvMdHp2C9RJtuVTNlPTgAPoIN+D9aErhVkLRV768
p+/EN4EqpVni07+mAgADIAVcjvXmhvvePWHVvYCtyjHGylTUqU7DdHGc1kA0nY/G4HnEtz1PGD/c
9mSyVR8zd+fc22nn5TScTVymWOy1bzS7bOZtnN9vyopu9X5c8uHWPvcNBRG4/BHysjmU+5jOL6uJ
5GqGTEGQlJd8lm3oE6iWSy747Ili3giNJI+fKJJJusZk962pJ83xwOxwleWQOPzgDwIoiRMCD9eD
Sxt5+qGOcIYlXVYwQp8dG1Rbss8mLpN4i03Xx0CU0Y019djB/gdyfNktK/c2GlLSEx/260BbYgil
YWkhevXJf75NT5e7uHQmt9A75Rk+rk6tAPjmy3ZxXSHwMCNpPGrKPdWD/54WfaMbJwErkkLyp36L
ErsqzZmTVSzpcPM4BLFhE0g2KvRUoBxLFrnaPBzxU7pZdInmCze7VFWLy3kEPeIKi9XBDeY1VGpG
hXq2X5Drsz7fdA2mIMgpTUZF7YZziY1YeIENRcsDI88B7q/g/NUXCIM+M2d+5S+3q7lLOtJTGIDv
SWvkGqiOOfeDv/F+bVWqOHmwM6fb2abr0KBWO57kYxQhNQ1XF8u1GKMVmdkCJonPAxjt5pG6EmtJ
eCYkUrlTzW6AzgRw+x6ZUVy1GHQSFYsVnA4bXXGSCuE2kO34R0j/HPKxsCQLxD0uwcKhHhhDWv5V
j4UiuqGc5qxyBGCQsc0x2GiPq+gFiIZ99Wm42+hX+0lf7wpn74osd+/rcTcVkuRxzOxP+4DPgr+W
42C/zV+Xf0mciECvBXCXNeNWqONTYCn22un+F7GXpSwpcCVR3N7J1fOXp4F/NzYpTxv1E//1wxs3
6bjXngUQ3VYrt2dug72YG6ts45Q6uPWDC8pTr/DHDEiGchztXnvKfLInAjvCgfpd49nXndjk+Y4F
y6hH7g7Flnr+A0ULMryP+QvGvGf/hhNib3WLD+GFR3VddDAyAi7MpRjnexTMeQHygsYGxocvpty8
frJ//VU9isV0KSubMedXZbDOh7xDNuTqXPQtJ3HIobg5SlxtGUdhaU+VHAqslG9GwEzlOqLb4IUx
ubi/EoEPBIak2uCOw//xOVaJb+nG/mQqaPV7wRku4vihVE3z8cqcKw4pVoh0kXt3BmE2kkOQvgQ5
dkhvSD+YZThQmTOgcUkwppDhxum+NQafWVRwC433ASQxHiPEWIezneiRc/fUVOvmhfnTDyiVJ+P2
N/5iDrdLZlJcDYM200MlbW8i962rEN78WznTa1f27mvDAMdCva7Uw9rHJXIba73Cx1kyhoCngGpE
k08oGot6izhMwuaLrpoYpBcupEDbJjz0AlStxlyYjLBf1I5ihHFZqNzPctzq90rDpYyIzL/64ntF
5CjTnVKl9bWx3S2dmTusCzdgdq4IrRGC/bsDJtfyU5ENERI9Q20bnGXSA0/iAjqI61MjblG413QD
7s6kOxsxSpk9omq32B5BAbpC9CsVigbjGXPAuEX30wzl9wxayYTmi4nPMo/gIdscSAv2jCm25vdg
1l04CeW7xelVW7JRXFi7avNEVxJ+MyasT3EFDE0M8XguMmfavjtbYAwvT9oQFdGw/wHR5dIAQ8ot
yEcrf2IVXRHti1J+2iMqKAwVVareGTRJAO47v61eb5PsfamMJHaNziMQn2i2isnWjMZNrZbl08YQ
QBiAa/wKNUmacHtPYWsBwXQIfnEVkR4c7E0YZNF+U3ZcxQX/jTRBe0/JkvubHsJZhCTw39Z3Yw+P
o/VA/soaGXedBVJlSCpwNxNej7FuMpcWRNTHKxFLU4KUw9OQJEphZtoVYFJiTtXkTBb23dXv/bex
EaH82l5OBOABsbe+zOxBRhVoaLO2WlIoCKr9j9vFjfm16nUBR4LtS7VzwBkTJt36YSdcss7Xsnvj
9lpTDhDcczwuYL4wXRKJxKHabP5crDXbDVZdr5bjXNqdo6P9T1xtrYNLSZGlMrf10W5+KVcrlyVf
XWo+xRPKDQBocuA3KMq72clHVPAdjfldjIBrj+oyL3IQhxKrTisQ+CWBZKzdxwFJvxgDYKzA0HBx
nZ+XnH9r8f+pfXOQypSseTDoGUQrFDH/GooSD7JYXr936kYr//WJAHUwhqpIbJjfgF7y/B20tFaE
l6lp9LDjyBXMNY5no4rzA7xaASmbGIAPJNgKY41EtScqXDuz9dugw07ZlooOFwHogAnV/BtZ17BO
Tm9egLV0I83U5k6Fc9lcxxjMsRq4UjbpcGtsf+WDyeRK954/nY8E4bsRS3StG2AQpdpexYRFqNzu
Bwgzz91bs5zelpJdUnaEAEdyyrDKVCDQ73ReRNUpzAscmmb3FkV1v5y5gfAMvHaW6AXo/5B5eRg+
WVAGudSNGcHam7QTnQEVM4elVIccrbNZG2KnVqHfSWdkcqmYbGVRRcBS1isi5NxqMTsBk40YlbkG
oPftv7KFMVbjf+Ytzft6mbDNTSkQ7B4B+/XLTY1YWnZ992rDj+4YA8GVZfzB5p9r+uQ0/4I6Faci
uUmdu5iceYSlOGu0t3ByP7DB2WjxTgnksS+oCOWkXAj30YPQ+v+8Yl3o4840rqnELMhszMJmzG+g
sc5CRoZblpffX1BtWivPUUjBLjLZsVQo1M1GL+EqDj9rvrFOkhBo6rB4jTy+fZUXYvwLeYsAaHoi
Qn5Ud2FsRllOP12PqdPUusEspNeuZCI4P22YRchuWepqjjf83DHoxhhNugmGnEhBZtPtPaoEVp5R
uz7gQOEYif3a5qnBk5vO8dh0IrCKQEQsutdQGadFi9jY6ylDX0g7Q9Pf4IC3t4A+9dzOBfdVI3mz
Kv8k5vYapg/F22F9MH/x+SRCiNHGbNd0lgxkLAtfgygwzjYl0J9rkv7DWrsyNVByvlHBkVhdnW1E
i7TZPmCoIY5WBwexP9MaMmiUk1lPnYajzpDzav3QRgrFvo6kk35lOZosIJVs0GP7O4xNpkOkk/bh
KkKm7rGIm+Jb3zA9RFklkTM1AJsCPdlPm09fqWMsfbQngCKL/6Ze7YXRBxVM6mf08OUellDCZSyb
0CfuaBvNBw5NrGp9lVliDt2aqaew7xnWgtksx7GdGzBwlr9qu8LeEy7fraMwgLEtkMaWrA77XnQQ
ADLbLB3/m/rzHC44PR3r/Pvl76mNJI4TspBQk1NkaGxqIQFE9mYH0rtOUsQdALy/tVSYW8GCP/6B
53RFLR9Jp/aKexLjIjK3Z9y6FG6RKZaOojZwLrIwRYD3Dta+UZcJS1Dd4pTnHJ/qWKHUaod73lS7
9YRDWilkYQtePHQ4+HwFWsdz6/SxwvT37/ih6EtYjFWuFv4qbL2xHsru/AkRFovb2mP69k0Yczf4
e+MYpKLvw9XgOl+d7KtdwRoBDUNr+pjlGkd+yszDtCXej+AFW58d31SaxDPd0nK5bnEreW4bfLjw
2LgqImw8pVVgK2fkU/pZBzXGEChWpYd8sD+fzdoRXlzVkdgCt0GjIXkk4aVR8sf5+VW62MMR1p+n
xiDbPz5oXKbJbQ0rn1iDR18y0T6EbE8XVC7kvpeyBQy6jE1Pv2wLsiFtVWaNuqYT2mOSz/nSlDcK
o0sQ2yVD7XId6D1yMAzu2YVmruoFITPJcTBuvlhoTBiYPQdSAqZmmpJB6QVokpKcJmRK32R+zN2W
5IKzMo1kUiruC57oOfk7ScivsYf9LKYQgfJe8L3YCN3FJow9wJBNLT3bKBMjdiJlY6E4oqk10rvq
RYE0IPbLQgFRFmmKn/dpDlJo7EGaYWJVduBWVDMIimZMc4O1wzGzjhFHrv7pYpS7OXv37gUvrwZG
z0TjZ6rLSrk21dEFYwEsN6kTgfX7wip3obGQ4spX1xHziu+bHxjaU3iVudNzWTyBCzkEMhF6DsOx
XTL1/r4Qgd37BqdNmJef8ILmVw1m1NjFlxlU6AmHdIQvOcPkFsb64tNigZANovWucma1LJhMfjXF
lRb2vKBLeor88fVsucYtYnVWAAr6kgqUXAClnh2xv2Jm2beDh/aUuo1Zj9EKtOSYhwA0N8riJMtG
oVX2URt2UkqnmbJ48erT8x6mNB4SQeN0+AItPx8PH0zgL4zjAG6NK+uuBTwDkIp2Hvb+TfMyW4+H
satZ41uu+pJ0WU5XOtJyuURpDHtnXRkYtIZ+aH2O7mGld5cmnpv3qmWA+J/DQhrhpKJmaAC7TWQO
wcyAJjb55enZB+5i36j0XXAHZ4md1dLeaqvndlJX76uYs5qsySmujNhB12p4QcpucjVwqM1ev8o/
x9T5FwV1JgzraWMDycpHm+ZBR6y2szPye7exVxO4vp6XUR3PkXf+Y0I4qbqG9yGZZO0ZUmMtIZCT
5FY5HOhaJ4pN+8gfscyIi+h2DhemrySeEm7CKchfaMdFgjqFCN1h0E5m4hBHOvBr4nYyH/7rQbiZ
tlUDCrcvZzcHUoKcRZgnWtXoNscimnEMgDsARteOUiuStZTYxZrnv29DyiGYacJ3cG1pTZJ2pmtv
JH5Yc/Y1MVx6ZgDcF21yTQh6HNkqW2+xO5lyy8ZUMuSGwHhM0yKR5yWdCVIEaKUoRBI4Z4HGJ1ij
LBAEVxupz0caaIvsqAwbVlYik08GV5dbDhZkcHUIz8fGEoLflU9tgJ2Es569Ufem9HHmnaDlCZVd
Jbcw+0JKFSt5Qo9IDR+zj/9q8KQrSbUHnT+XxwdpBE7FOW3ZTPVkKEUI4I6wCmQ8nxC4eMl/aXMa
vFYCwr0pe8i2GaNL2FnW76NK30Ozumj6k+/U3IIE/AZDV1KpSHwqbHz7mnepwwFRLvzoHSQ6q+8F
VlzP4TKaAxfWED1yG2FHjAz/o8N3kcBy+/jAWLrg2te8H31/5GdaZlP17Xu0zSlvO/W1yddVkolS
3katk6bkI8S6HMey4ZVYJFURgRTN07ot7g0eozteFQq4kgVA9FIPdg2Zz+eG1H9tY45Zsv1rrl+L
t+sm2ar/jbbk9mS4DTe17Kya2XV2MRYrgM74hcjX3/Utm1hRqqeuicF/xFdTEKvNugEnNMv3lsnj
LJ6xm1ybwN4b6rucXKNqdjjf2IbD4UlVDoHxEHo5khMXCxYlOoZ4tVGmPSxLfKjdlIWl0gGNvFuv
fbjqeF2iGn06X0eUZ4CU6MjUaYHVR/TM6STAUa7tl8Ja3SX5J17yWiYLCCaNpVN25AspALWw9cYo
I4aViOGXTGNbd/IpcM2uuNCWd+dpd9EvCrKiy6iCm+VtXouS9IyzmVEJVJ04+sPyR0/M4y4XN2Vs
f3t4iS90rNPRM7vtwYC7svnEJtnxWls2yELQVhaBnWGNe0tE0enfmNNu9p47SrrTeysoFCo2gc6n
/FamJeP5k1mK3TkZpk/wO0Vtr6ykfS14XoPAv+ddjVx46HNc4cF5tYV7F/TvGz+yfuWNYj6JNIen
3kJ+4dT5uUoDfUJAWIK/4wp6P0XQHTE1nEh0LZqvzxrTpfMeYYx6Dqcnasx5jEdzeVRBRCXkc7p3
+42VqTjoGM9N3WKpZs0Vk2AY8uITIbC1A2SRspXxnAAHIWvKHEXevoVxnszMI2ejebVRVZ2/VW+1
rqf9QLZK5X3QSr1+eX5w9ykw02QkM7ZK9nRj+2JPPVRrBv3uoF72NRtIFDWFkHK+U6or+dKIrcXN
ok9cYGCmmRtyxevN91siIV6lI0GZ4je0uN4mpdddF7Lxq4P8Ke8k0U2DlNQNOIWdGNCEHknhZ6cH
h+qmov3nRQ5tdi7XaCy9l88bbH6PTxujvvGLyRu0u4fdquonPZgTOf16eMuz0+5tSinLKPL69gXG
3NMS36OPQzb3ead8ZtP+tw0M8IaAxo7P6atHfPYQl70iEvsmjyymajWvXheciATIjNeovFME13kP
GF73755Dlx6B+C+LRIJDolgopScaRY1VJY85oYxCYHXRy08YxBMKxKqo3h6sC4ENqELC5PQ+BAW/
SLeoEUoGp/jvcGITqmEhJVM2NTTef3BxWEwqgGFJf+myoDtWSxx4h7TADuEhckJRV8vmJm7QToUF
PoNajaIKerw33Zz5wDzgE/jHnUa7EmBm7/QLigszeWMjiaK9nOQ9Ae9MsqNqnRsyG4KRW8p8S4z/
e2+WG0wwCZdqRFkPcgPdXzAfD1mRy9HgJYXch/U9PjHCdlr8KmoNsy3dqR95hP32jBCMx5EJNeeY
d5KRfVMdwnhMqNzpdtXtP1hz2frwTLt7tezdYlPRN0J4PcluKwehTFdat3P2DFOYFNUu6Msc5FZj
ahG/67kZkFz4ewLcYtzQOQOaTl8Y0CtpFvO0nHk/7IbrEhDuVkAmrt5UsaJ3rqVV4dlqsz8Nnkx7
UhLqr8NoEHhFq2ctnoT7MIOzypvGcSwN8Gg8uv63hJzjyeHprLqUT6KHov3j365A/2sGl+D/Hw0z
bwgpNDRiOfJXh9HfwN5qCbUiI02TX1XXZn8f7RKDmkmCN92vntno0NLBGieQmqA/zKebzFqdxgpM
ok4XtluQ5Th1GhbdbEivgYEOraDjVR/2ZO/x+JeBXAUXz/nLHTAdtiRZTeCd4N3yrO1W4HM4Hv8x
AyQ3vV5TZ3jk8xYUj/zsyqxp60IUuPQQEHZ+tbjEtgWUlwdjtOxnL453ZbJxYVmX9qNf9VZDNxlu
1gv5+7hmMSWilkUBNNuCukkIzWrBX4DKXmnN78o4wW6Q+Nh2KV6inhCriyPehwE0Dkv51fRNW+na
7/kBMujLzF2vGRBAIgMKfKZxsyzxFqO8NYf9nBPCn0RxlyzGcdg4HehQwQyuwaKeQgdzTXTqerE+
6cEWbggCsK68SbpJWzuXYSD7B60A5WDcwqu8vQlV+1NZkGIpfSGqSljDGVA9l+dLVPqTqA+tFdq/
uus2lgvfqBdBg7xGsyFfCAh9bWyiL5p+zVjeypENbc62Fuer04vFgL6qk33quRjyNVNuJmoD1W4n
X6XhZiCnmYGMvtYmf/dpkuzMF+1ZVeeSQNkIcxzW2DZMJVwpkhA3TQWA6uzKN8NEpwXl79VLufHK
/mKuhWC7mcn2Td4rJgH5hRr3Rh7qaPIv78/ZcKoOHwmOuYEtlXWo6WoIdfF/ZX76vE1EjzTC3o9p
EpK8ChQ/l2PbaleHDLMaXudq5bIfNOO4dQ0B9lz7Nl+1rMCOwJYF05d3s47nga7rTjEAUj93umXD
MPQ3xo8irdoVTR5AYPJlfWHMnpCtF8xFGlZGy2TIfsaA/d6icQuA7BLWBFUQIOku3qK+wE3IEMEs
+qUNnVxAgb3uK7QgTSU2twKy8RQZgjzfTB6zLrOdj/+AaUYU4Xm9UmEGLb/xwMGX1Cbm1asvFA0x
fr+6sKkHkJVp+5uNWPYVBHIv+gMmTgPquRLZZLgQ3jNICinumhXVSk0lEv7bv1qKXcTRmFSrwYUX
LENEB4B0cfrvTUl1IoTGKFfQZKzHIqTv+ph852ve+9g1xTmKUW1I4J3xC/7f7+82uGz4UgRwrWA9
IxIJ2VlSIhkIUjDqU4wrF08t9zyUjdRAeecuYvC87KMRJquHLl//VvwP5VKbXB9O8bOQaLFuOOdm
lJ9dxn6/oVkbJDEdx705YiRvtrGnRxQmg0ClM+SQifmcuEiYvZl/5Z/VuVwLIF/cA+O3Nz/vA7xj
OFWJ8OH0DrIWJQrYTJxE10jXsdCe1QAqZ7f0gLegY5+aaH2DdtZVkd/l8WPbeQsTjoJjRXAD8O+E
fT9pyB4BIJdPe7ygUgdhfO97acAhY1imZrkxYaz8pU+mqvatRwk1d7QwJZ+vG6jHdwyPnaulM6d1
ayjuu3DdaouI8jFXPeziQfIQWmVee+erSSNX9Zy4e9RQ0wuQuCNJ9EqcAUqDgUySQDz8HBRxZEUu
1lomqvgJxLxIxw/Ib1C88Bqin2p7cEv3M5WHzCshCoDtshaHGesVo8qGGcuYcR9kv+uJxfyhuE/s
6spBvkDi17fLSgt4WaLlVIa6kbjkxQxjqz3PeXUBt3JpAxMDsv+npPqPzeN6RHmnaKFTyl3RzDIK
2AB1WoFt7A3d5It2o3M8F4TXisQAyd3rJeFXP5wT3ZMjuSK1KCs9fR4RIA73gyhj181fACK+EdXI
IBYf1+ItxdpiJCfxp3ihumksJmUQMurffBRBh8zGHnRt+gnGPtDqgSdLNAWErqhVlFDSarOG/ezc
VJR+9cHD8+B5+k+IrSS6A/yzpNrY5A9n3qvKuwAfBrnVt91LTm9sGjanh2osNExSPJ3TuDME1D0A
34ytCpNvtF+k/AuhY5cTQxIRpz0Fs1zwo1RzutN+8mz6HdL/YIKRLxCvcH3cdIwFv1Q8w26gQKpd
hzytnjfmNvpUJyN4qZoAV4xakXvG56nlH4/iJVZIC3oNcBBHmVZcDD3PzRi7DCRRl4eQQz+SP8HJ
MkiNvYpr95nG2RKXo2JNti+U9s41fgGptD0doRxAWJsjFqYqoCw/kY4Pp57TRVF3+RhPPb6D4hU6
FhDqS5AUuN03TS3RLxGCHBepnPDAUk2nl2VtKWDUY/SNXVz7majunu96ptodRfqiK6w0g0GQ1Xzk
wZ11GcG/3D/Llc1M/KZBokb22A1VQoX+baJpcah7AtnNd/Wuu5ENV3l/J2oVVZtAVrKQlAEc5mRm
hg4hTiVurk/leBH2lBo+cX6Wnj21kDiLzxwpLImZfd6PK5brBL36ZcFOwWJJR29aX1ZBEl7OxDS6
Ak6S3a7sx2On+WDf5nqk4umjDQk2QPcLoXlOMsnmo1hhwhmV1VrWGZcDNSU3OIQVd7xZ6rZJRohq
PLYkg9jPHWKDzD8g/6AlDmUucl9kr3gMpdTo2yqItiM2TvHqCjoQyUjoF/VkrIQgWK/isda5QDZj
bDzmdXPiCAY7ozTxBKNXOyzREh3WByZ4NQLtfeMFelJEAwvPH6tt1Hxq8E4Sli6oFPt+Y4GgOY3y
U331jPWa7MkBg0LMVDc3xkqjMw2TeSXaKI2TYVjyxscwb5ZVXFCkFzaNMAip7WHnr87eDrE3RZkC
si/faAHAb7AtQTtoeH0M2owcGN/gAnG5gHF+ZmH7BoKQJUNsGnufj2bszkCP6QTySO1xve39xHVL
FASL8CtKb6iwKJCc2Zj39XO6MDf2U97C/ggC5LQielqo9XIsupr/D72uBwoBev+qkYNMDM0ggfxy
Ya3y0EFdNythdbrTlJ40UwRLFFs9r3a4qzUd2nMuWo+TbpSMdsT4PsqUz1xiHdptEuqVYBvZemjf
rQMfWrHhfUEQFBC+Sy/NzfEB5VI1EMzy9kfCpqZ3Ra2XosCbPD3xDFKxO49aAok48pAmjI1sd2tx
4+0W9m28akLwhH5X7d8AvnZR4IWqI3IWcu207kJ3dyT6u73t1x5X3D6ZGgYo6/s3GlQu84d7sQ2k
mc6xCi/JEjx6fTaGDhlyLIY7nJTXhivrJEn7G0F9Hrk/EDV4lAJyN6bZYAlOyJx09fjytJXhRwjw
ChdQBDOe1/jrP1dv8pDRhZojXRQX3CNWt5ztVJ5ebCBIP9bjawn4DMHGAicGhwhqBgpx16okeUDj
CffcKtamZXDocMVFlYObFvfROvRYVdDw4BqTbGxqbhN6U0FNM9mc8bby1+qR5PJOjVxa054pYkip
tOJyh8Q28xShcnLwY/H5rD1r9qiEDcL70U+C/Mz5ARyB+1Wbpqu87ejsXIs3+IzNR5uC1MmTh2fO
sk6Jj7CYorVnfcRwQvkU1J6wVnlW1IIrmsS7UyfEnP3e9DSVRBjX9fgg6bb9WtKAs51FjNLpNppc
Bfwje6XdnB5oJAwELlE7SlUbU6/a9L/hhwQojFnBhlk3QwErV3C1sjkGfnkG3M1YxT4rSTmxIO80
PVXIgdUFl+0UEslyABahRSQNoArcP8jP4mtoSlbCfGrO5qPH4Yck9/Y0n5Ju0W6bFG4kV+cgseVg
i++u8mMvP195db59aoVQ7Ndk90CUHfLD4dfJ490lvDbG2pMjCfQtyTniqvWovUkSdVsJcNE2Kxo+
PVkQS4IyemMG19XwEPVDTgXMJQpQ8Xm6zv7pCYKVveO86XL4dpZ4HgEYJRgmiLumjoJxc//KXx1l
DSwjzaI56IdqTrnM2DOHTLLkj7z6K8guvEtEQnK6ShBUBj+QWSZ3regwZ3lNrRqUNDA5WJRGCLKA
UF6CC5GzJayp9DOG89BijAp/ZvY76GZvxpCNbR20DJRqb0h23K6RQvMU3D39z+P74TIZwqNbdqrc
eR1tYyeGnoA/51iEPLsxBIqHsF4vr/FFKD5ocCOtg33cC72/d2Y4IyfgqBiy6GDiIdza3ySa9Px9
DcC9j6SX0wt08fGMbX90zSAUClxo0MVIJUQGH/Z+Irgw1Jh1vVtzs/I8yccm1k1+OteNmQnOlb2k
hQzoaGAvX+8easQ6hIyS1siq8FItrGICzsznMrlHh2iy2xRmYfq0vSUxCdqGFIPsfyT7uOYdISCm
MUeHwlrOtHFGUqaCMR/XqHZW6lypJ+8cnFQnVa4/Yp8T43A4RiHoc6PUJCGm9E/KqlDVnCDxa5Kv
+ACgfFg/PPUn2oqNPND/xLG13uaVaNAhtb5JdDHuioWYJmlQ6+rjZF23gAtusd6q+7ZFfIcf+AFk
bxihRRXpizqyLgbUN4dBQh8H2AgBPYnMBRrkZHFuplFaAhc+YgJ3NZMq05VZde3KSn2E4AuRBo5t
IYlpkvAYo+qH/iSHVcMIK96gBrrAX7NGGGV/f9C5XPw5GwtxIlT3jdToBR3s/Ef20YXF2elPOwSm
GTr74VYjuLnfF/OK54sRJ/EfrASW7UGxYii2ZfUSoDvTTDcoKVChxFRAFG2Iy1bpz2X8CpJ7hDno
QGZpbNyq+KMKO2wZ9omTQpMXAdwAuFWaZd7knl2PPXF5AvMzO648fWZ1rr7NEDoIT46PuN8q/h+S
KJ77YtB3QmPntSXMsOK9ZyUKXUdRy55xE8x35DauFeXCRSuGZPAE/JVqsTsenGaDGt5GjElsEbkm
/sFcfCXmcrJc/pmCU9qycOisFWf5g5gRjwZy7z+TRxOrEUDZFJkHVrlEAVBbjlcYlWDckepHP+2G
C0CFSqWht28yAtTC3az/u/HYUKCNTfKSkoWFwaJ/ETxy1Kv1xuzg2/s8iEdDc6nrmYCLlGd11Fmg
dosJIB4gX5H47/ucv6K+qVGgG6lBV5WwNbxZxBIoamczF3mdy+dt3JSDfamyw8VZLvhc4kfUf5wS
Bb1MdLGx2NCHJH2H0JijHcFJLEzcgIf8jI1+wbb2iouk/E83SvSvyDoCV5hIlpOgK3VtUHhzaMEV
n9FTUw04lxp9f0TgihJIPmychZyYPVmjJeqSRIR/5BSaUiLnvly1Ndk6jvhi9M+oEiB9SFGcmJyC
+2wYltYqKwbDj8hrRb9Q3UoJgQHaUdYDnygDeYQZkDfi1m5DKsnVIp18rM/NH2af851EPzT4qYou
xKRba72gEGmUOXaXHRhmUFhYa4Zodfuqge6jRXZgA/qwpdtG35kKpRwczi9EQuQ/96d9p+wRlmxK
j8bDfdaTzgcp4zHkUuDIrKqGmfLYIGIqEuC+QgwgWJ8Pli/rM9Uqxfrubrv0c1VtuusbYSGEnfVY
qkT0t14komWP4ut4+5lsghF0pqpTWO00vH61kgn+Y1Vcf2Z47ImIv7vInqJK20GJEmgNzCluCy0L
jg/WCtqj+8Gmex7llYMla3WyzedXmXn6ZusTrN/x2lMJmmvLcQOp+FJRFRh8y+1IARXuQvKI0e6b
j3k+bAvlbhwFWjKMGgaV7AuusVNNQ2Vv18/Gfkjf8JU+0ix7utntNPhizWss6ERhEysaxQu4Xbok
dlR2hJgYZG5tqPGGg5YWm0QbV6DfjN2r3HddyGziPCelgaFYKyk8yvxG2BxICgJyMUoWDogFes98
cTY6e0p5Tz2E5xAnuwMqzowZiKOkpiDgI9qz+laXHPIL2bvi50wjKIj8hxxEK5IWx+5vUmkNMEui
vPQvw3i1lDAz5RiQZHLqm2AMaed47nQJ8Lhe963E4sXB8nyaSqhDNAzYuTqmR55ip4JFSVV7W4hM
6gv+VHglCmK6UE3j2m4ey05t/nekeHyZVG/+Pq4qZlqRMRS3pRUy0P5M/gcf5pDxaku5GHN6OjjO
wrpFcoHIJhczcOnviiR3aYP0wnuchrCGWYmdf/AC9rVX65hGOoJ+dSeP7E0drSHz/6oNX/hYouq4
Th2yaEJv/B2FLPYPagSjZdElZ3nqxg1mAsNllaDxMIcwqraO/thlyIqHCyNvofPQHMqqfuHAOXMl
R3avBqNIrAgSu/9w80FLFPdobjMrCUjuGKeHTfedIur1fWk6tF7XWZ6upBjmool5PRQj2p/qBHfe
LSb55QB+uL7G+jFg2IkgwoKsknbRIMUx4yeiWHzNRVGHY8hdGwYTFfrfnmAHOYrukF6nrIc2insC
ktpPA7tUFDwfjL8cLFzMDumXWBpQ4VBlBqG7+T9oq7Ea2+MZ+krBwY70WH1MJT+9BeXlOncr5o1W
E6halrWUIfkl1a6y0y/cQowaHnYFYo+WON3LK1FRHZBM9xwnSm520Uxa6Avo/Y59f7nkWt5anEOK
+76fNc5iuVabFEgDOF+3rTQR9oT3HPSgKKc7lB3ipF3m6LQHtnDBDS7skgMDzUYVmuEb+oAo6DyA
ARDBdu50SP0IKi5yjRMcPpbfUO/e+EiGE290ClmCtsHTugNFhSBeD5pWNiyAbpYXIvSzpS7C/+yu
uh9tHS7H/mUTa+O6A/zCrXKOZQ9iMA8N5aKB4cDusohmVlr5zgDmKz0OJ0sokwztX35EBaMKNInZ
BdgAv1IvLqOY81R1bObQ4aXJnGuWgaWKHBAPhTMHdHEKprOkqlwe8iZXTdlk47dnnLhkddcO/GMt
AXKW/yHOwInlOYGhPW1bDmXVNDTbmEn0XFFws2az86DDq5862jNNAxpRt2DzuLjwoUJ5VNAVlYmA
q14HLx+NK6lhP6vkKJCXaS30I6NMigL+m4r18QZ+qdTfVLq4DsqX3pohAQuASNkPLxO2NGR9enZV
fcP2dxr/RTpuFWhxjHR0uZAuiszIbv24NaNN5n6Ci0OwNQD+w4cdLFp/9xt/kp/PDogmiTfNjixU
/NlEO8Xao8fRMVzNzA9gCyH+YJa8UUYAoH3O+WGASDf5+gSgbG5N3K7jwr+xaL+zOb8q89pGzssT
TftAu+uja6eB/f4Uq1Bb4c/ibigZpA7bIFwSQexeLUvwBDor8Ik9FKMUoAfTVTwtqX1acO3b77eb
6yZ41l1r7roqDNT0eYLBQpn9lnKDGrQPiwoeVnchYD/lvOLkZmctGTPQas6x2wsUv6OJxtduxa8s
rmUAgNuxSyIUDs2sWLwX0jitmHdJVOwxKFViGyl27TXm5Syt9dwrIeERtQFBHY0H5Y3oCkUA66o9
bIsBW5xY9DT5U+zlNO0sZUjVXSC2UqYHKYn3FwWmOrHCziuE+XZZ+r1gecpXMOGZiNITKCG/faAz
GXLp5HeQMdWhqlPjTG9FaltyL2AyjS4qf0MVQL/7nmGMWfMDT8URP76E6lQmULPaAAdz3QEfh3i8
xXvgbMXvEkjh6MuAj/Ws9iF5R/wy/iF86OX15a1uWZA2AiES1uklszTrLQG0Wap6YiUpylSQJcPm
WpfqCQJBrxejLNSqckySt9+QfFWKm8EgmjybrnOD02TlXcKdi9i3yx5FuGG4baKLahWlyr/Lgw9C
PRhOV/AnT1gYpNq1+7IyNnCBWU+Clz0m8ABu3VElgp+lVp6aSjKX6IJhcP4mctrmj5P0cPEWFYf+
0+nkXBos2qRHIaJG17Xy7rqvMcdN28i8PjbzcoKpj+etexoTB91UXUkYT/V1DNJGdWEqB6198AMv
3gBULKp4ir3r6K/bqiZZ6WK5tmAGV1dnYwPi7dCm9Y00MYJ/UkytWE/Ghr4LuTpTRAbLrPnFN3dz
JfBndPApndJMgGov6O2r8E+Tpu0GZ5pSgPAMUtzaaWlx+YQHAdHJ1kd9bbHG4aNH/gn9Yp/IWXLg
BMjbI1JavoOgE4uK1IvE2bmBLKoiUaltn19sFLaxnvs5p3LFgvemeT6cL+jBEGD9lB3zNg2lXZ7f
NQGduiycnqrBYQrw04fGSPMSQGmBOVtj7OgE+Wx5MLUvGy+Skhe5OyeEPIPSDkxFiL1e7E2xVUQ2
KburXNEDNqdvm7aUkiyD561JYhDKsCY7sMI7fZyaXZDmLK1HUW2Pvb1UObYhLQtE1ZRCUqzryNo/
pP8ykk87ckXbGHowm6hgNvtirXep5i45dLEsaeFZHk/xmyrPG+fLBo01Oi/moZAbkCszCco89g5G
22KTRB9LnPfsvIw37Jq0eEzO/dTesi/Cp4wV6Y+88oFIeUzb1woLlG+JTP7uSgW0mm2FbkVZjcQ6
cz89Myk4fdZqgQmX6sHYGanRaYpnVMj/HG2dEnTepcwQJhUCwTh6W478hNp5AEJo1r3sxXcXgoW5
u+Wre2IdNoN+yNpN48FtLw2YwkzKKj64je50iZdPs6xX1/s+25Bf/QudIFhTDPqdHyu2JwjUNfKW
hgHrwVqWWlW5KtLjiuI9CG7UrPETVmTs6WammujO4NMtOfEAZcRJGQ9ylGtpUAlU3su9/YEF4od8
n/D1WO4g3h6kvkewcajDwX9oUwgGhGtm7YCSWdjv6f3/h49Ixv6+xE3Yl7Y/PKI9zkO8C7jxuaxP
h9bgLD8Qk28JL2+oBKydk9myHD8KMU+sZw7YX0iasKPYB1nzpCRMTEYMijACxzluuLzgwvdUo2ZB
Kmkil5k61ncDBHQM52e+8V/fQak4DWHL9NWQJJQVr+zTuz0TYmYbJp52/xW8nOTgk3m1yvGnH1SK
Lhcx+qHqje0b4aU4xfQrFJLqPQqGZCrBoGPHpXQ6xezUh1I8A7YA1hpxG8H+KY7Nzc1xelRCgK2h
q3tEHgXMbCpxF86X0vPRrd8Z/Snyn66OAxng2DCcAVCEB9OKsgeDlGJETBhMvAlFVxgBw2YYxPfW
s6/+dEfPY1c+n37VwA6eLb7GfeUqfEl3cJsQlaq1aEMgrKWWrYMIG/x4tDYdqWu6CBII8a8Gy6H3
c9fyfFqKZNCmQdaCX0Sr5lopfS8rCa053KfbTim8R8ntQy2g+8kFb9YyrC7Q40dw7VgAyRdZV7Ez
KqNU+8ZiBinV5rOvwy1czSNfeZ4BRNhv9XasgunPqXGcIx9KK0IyYZyh/lKNvZDykheGINYZIR4m
a3SLFuwS5UhYpokHPOMou4TSnYeQFebN+yctSugmRiyvRUq1YVMEg7vXqNZT4mrGXxbkx3DCCJcn
wQb+q3RSN+YQhZDaUrb3Qf6Y03tpKcpZsTYEKz+h2sh18vK6yFvD5b6N2P/NoM0POGg6zob2cUjf
R7B+FHgtS/EQ0heQVdg065plinT6JOErCpucj9Gwdb/T2yq4togat7vl8QogrrsrfhFZA2KWtQGs
rm9s82NYVkdyRwQ3YrRWl1T/70A4qOUG02U8P3yqx2Qtw2guLWo5ISmMVwO2/uRgimiystajc5mS
ENmYbsT+99otgJKShKdSwaJorZ/Br29pP+g8KRDNfztggCWUboYZBeiUE4MIxvbVi0XTkoAyV3Yu
NOSgrVvyR2McWU/hrG+LKtA7z3Qgx8hJpp8Tw/4PbllAWo8T7hGNMlx4Ely2OKx/8I6PqF4HrLDk
PP7urDpyVhJbiwu3OeybbQ9+1qNHQ1e/reNiOqXqLmoFl3PX7SoBnq+4uSC4q+sFnbkialudOam/
YdsE4rfRF0EXzGdAgs/tGQxvc1n/hH+SS6Dtkd3rJH2EaWhL6AUXntkRapG4VoElmEec6IdB/bDU
LygoXH4k+4onIGPIOdh/7Kmkb2caMBgm12ciuvRLUGVbODTsNDj7YpazAVIvcgs+njl5gDWdI/FD
iSCl/ljrZJQJTQT47WP+4GjIM1QJooRRxeXlxRlnQl3ZNI2+jj5Ai6e0+gsIV8wQML3Wc8D0jFFE
Z0QDXyg8H0CL1dWEuwFdfZV+Sj1LiDZUci0a6q1eT+TBRzwT9/gcrMmnZ4nJdTzXYd7CIB4b9CZ1
ng18L3aFkYU2nEebefmvgLsRy2MlOoKUmM/IHuwAg/Svbvsc/QNXFD8PRRGek662L+4sjXTB2F5E
uPYzQngDHnZK+CG3LeXrxxXijau2vKtlpQnaSaAmYZ+cW2seLQyk6Xz4Amdt6D+WLu3P6jkKBzzX
CJ7K4Ih3+z+5uud0ykCH8YLTaC6lOoLTOOZHhxLf5IGAJsTGCtVWuUEVB5l99qtztUthg/+VrAI+
EsoKV7OBULDnrEoxEGSCLRXsn8bNhw3WDWkI+SBVXu0p0lF1798RvslGRobdpV26Kak3p6wbwYfq
3GnJbybl2gnSU7ua0/a57+s+6TcnVANix5iQ8vupBZOfPLz+AySzaVogIw+Nw1rb04NwOZM7WmOG
r85ZRMtlB8WEZ1TU8A/Bq4+fF+mG2sDVkmC5RCxsxEbjOJ9asvsLLFiKclDiSVqsUuTTJNa+2S3K
66RvaMQYdb+cZD6vxxUYONbFFm4NRMKTA2srZFKT/yWD17sqyRAqqQFNQvLzE/epn5ELYoobl+1N
77kb7+okG5fjk7E1LYfHGowfdBcRrvGKgoioqQi5VrRth3Nki+jTrQRBIrJ0uY2cqw667em2rmMz
RHO/r3AijXxo4xT7xMXtmzZexy7IH1gjUjThlAJ+X4Y7WRzv6GBX1xT0gjGgrRy2Tn2bs8CT5nnW
DLtf1k2/vAxoBViNJEtHBbBK6C0zfiwZcqfGKbMQvIp5l4O6BNxDNWtQjD2DgWb/6Or88HKJJ02s
9BQV1h+XKERirP92r9wNyIz6WgZbXckXWV/p7QrGklHde8XqlTDXSwZihkxBthmBHvNu/zaYjWyp
HRYquGdWZnDwlx8FKbmeMG3v7FekyQNR2syKefu82QmichjEDX/EmfZZ1bw77Ctge1fEUHS2BADO
xKVg1IaA6AZvi+V7MZw5ezTT9T4ADxInX4PYz7LJ6EbakGWSVNHb1c1RPGL1YiTDTyStHzYLbBNV
QgKh1Ki2UemDUi9TH81nn2B7jpnu9VqCJG1Kkekc6YLhA5tYfkTwCtRuB7gt9RTB5SxtIWnP+2Yz
YBUAUAXo6EzuNinvdn7UXBfhktPqx6OKana/VZIUHT4QDfKAnIb8qAoxrKZ3zR783D6p3xkyfJ2h
X3i+o5kT1uglP7grk4XhohNetYPMZp2I4rijP+m9PcpAFMlUck8FzAeEpW8qNmbakMVw7Cd+nVq9
HUliAjQleNvpUFJNkm2/lNJjme9ryrQjzUXM28Ydrhsy+LgLy5+yAG+kSJ5jPwEMAyIbNPBMyeqU
lpwQHWcAQjPrvjmSnxmys0YlndlbboPxZ709Yn20b/JPFXX9iQZsgCSf/ubtWhMP+iBqAXdc62iV
m6M5owmXuARXYyWeWzcZLEP7ID9ZHl5C9SH90ObwemgDN69WvKezfxHSMU4tiUYUzundHpAyxFQx
KfwWdcDEBfH0swlowzok6mqTlrH0mfn5Xi/DRAblGAARWwC3dEKaYa8+bGnhdoQDJ6m3taMKHZGH
+Ic/sXeBAvrsLKq74Ib8dPMZ+OuTcWFlrPWnFvE3z5/uwMOex+XzWSN8LpoEWJdhJqK+ZaOgQWgu
/G6RUWIyeth0O2jFWVpd6tG9gWkka8l/+C7VDbS/bQlD8b/3+Cxb0snfngwFhXWiySPv5duiFoo/
QYIzA8F36tBagmHpbg8niNdfdIu9IOIPwJPOT79ImshPi/M28DoGcNT7wrxONzGS9s6U9iqx2wUG
K/qRU4Jh7YKAwtpNzzTyPd2dTlFgVVvyh6py488J9+FywSl34Li0AaSq15HTJi+q0spIkkUc3Gad
lfriBuPOJVBCyZyHnfk/lRN8GXMJ5GSmZLf58Jdvq7RxW39IOihbV7DHbh2yoCNWqcKrgyJVuG79
7naUmdF+D277098GNXJYGHwoWrK7VzlRpeG0xIRucPVDktuRKz6P0q2x//ms94FfKTsh81CdAOCX
Xb+/c+t7z9jfubuohq9Dd1+bg2AuFYYlSK/+aHeZQgE7CR8f7RlNl64Sq7ueSWskxX4uCGtCGaMi
K0Jen0Vuoq4lwHxo6C2Wj1QD6gXgswH46kueExr25H4/Om5IEmQWq2stOyCTW0FgQhwa4v/fepjg
lQ2qwVsMXVZ2zMoQQfgZ/Ymh/dgXAOgxJCwL8AgjD4udAWM6zhowK/pr1ts4RQBshPhAGueCwFb4
hDcPmLDMzoDvQUr62TU07buYebxU8SJ5pKh9H4tHG6Fn5cQLryrn8hhEnC/Vl6bAS8Hw5SKyBUdF
cX/g5tCESpnIBvcO4TU8zAe/5+kfb1igRJIfkJTkavG6s2BONCHJCBLBRy7WM+8coKbudXZqsTIV
Xxg7BBPsxJPL5jBSkzdYP6Ay0iZbK1dUW6g28xrvphXS5SGGLhzbykKS84OinuWNaagoN1rMeP2h
c8nZkrIQoZ1MmTqUSEogeZj8TmKW9Z8q9fm4qf0HsVbGtHIiSZ3qY2ziWLdJBJAw1a7pVQYc4FC1
L7ZUm/EwQ1jfZ4Nd9Ez7TvBOGGpP/vX8x9ZE0cYVDZVgapx9eh13OnPtFpJt8UCrjgK2VHKSgY+l
DNfoJuZvToa5pS6Two9HHmhOKwKqZrTlpxyo72UMLP5y+YsjGigvPLmW+S2zTe1533KTw4S2xTaz
fegOdbterlghzgn926X6itmYxlf+t+VARWlb1glb6rTXsMEufmlMPQe/aYXNbH+5lW32wKXcvpao
GWnMJeqWiGLdrz2I5w17W2sXQbAYcW2Ow419KiFyfQ5fV7OPcuuL9Z3ET4kxplX/9skKtDqJHCjQ
D7BH5qKOCxEikmZ2YURbdXORuU69ZbxwCMtKxOXLM75YA/wbSDdpHs2sz4i4Ui7ZtdmtoxhrwR5W
9eBJUkEQBY+TNEroIjI/MIuTDUGerF/mSAdUhRUo6pKWarpW9I0RxKlDJbnLsfLzPqGHwmBprfTv
q2ImIZuxaymhlFrcuR1x9x27ARTgFveTX7N35uPWNU/OF7kpNipfhJGInvlUwPiD6APDRmdyXmU0
3489tBJWdfMptLCQCGNwl1STvhu1AOEW+7oEos+LrCnwrQvZ9OiqGuS11VG0HpznxDxrIx4un5yz
/9mTx6bCR7kU5+3+65K9LDxnrPpUIc0LUG8qvbzEp7Kb+tEVGCCUi0wdOs4Dhmi0onfEGljZwAzh
yUqGvERMQZEMVJqpN6Pb22gq3L9yPGxIcbee1rwJTnTZQ+aJNZF/IcHqBZDW2obT6AQdfgP0xgid
NDA5eQBc9VEYAj3t4aNmh/hYZ9/wM8OatZA+7vHeq5QxYZ09LJq2QgjC5sa1LeNBwOAuotaGx70B
sqvOPNR014X3denSbSmI6zCdM98dbhlKYv5A03zMUD5FPVtqjWscPJojYIJJkxDGcPMN3I2hUXhi
chhZkn0mYQp98DWuBKfdg7sdXJFEOE5gybRqqW8u3yno2LEWYh0TUBixelhWEGOGtqmQp7yK9aTV
P86g4qyAC6yBYnPLS4wK+qOOJnDnz86X9C+wwzqqKTHsUW1jgBGL2bzA29snYMmoIUQDafCdl29I
qMTLGpdEbrNhykj1/L8bb9nA5IM3/LF/EypV+J7jnCjjtF+jjvOdzZqWRNRQBSvpDUvCLY6E/cfQ
aly2zXeO8K0Qe8oifvJMK+KW84jC4HGeMm/W1bCrJv41xd27m6LU9D7iMcT5VcPBnJAJs8Ib9fY3
eXHzdmn68gFgANoFcABF3vwD8JqZTsBxYshuWatfg/G9ByJ8VwHOmhiS2wGQE3o3iLtlENQxRSR7
ob7y3ugLDZSURWjyGkpmiNPY5glALCDRYxWqUM/oZTps6lwk12IQ4yxsB4gRzeXdByQKWDqvwBxU
5XTwflycj0/Dq5oQKsy5goAn85jUWn3vr7vYjRAh9QYB4xMFW7DTNN7/wlu2L+htYNmlxtUloLQ1
EuepupjfvISI9DMKuys0EBvtgyrnZybsqOFCrx5WQZxMoUVxqThW37skFM3m19n4yFTQ0V6S6efs
FO2qNnOWoR5vGpEpA75mxYLlefcf7H7BriaMfc4WrDJOLrqU7JPR6sT6hiJCl3cnKa8B/daCFOjn
PMFORS7AtwuvdD5L4uI4OEFlqz/XzYNd0VOTW5Et9o+argR+iZMSV5ct/jDEYoTXuiiSRo54+8ul
O3CBS1BJUDG1vwm0NcSojBS/quRLO0WqS18fhgIM5xf4M6e0i12Mz+i9R07oWnrI0wlB+QIftA1O
mYAnkqkPKsz1p/eJSj5sUuv74rEpKkokGH2B1g6a9JY4a9aF5q9GLqus8RqwKxUNexDR7LR00BfX
IpYn2n9NWF2fIQM3WhgAdC34wjjdTWS7AYyFZ9Q7kx+xsiFc6/enA1Z/jbiMS46Y0mkdJQqRAbse
LgeEE85JQTILsQYbnuNvOW65wnbdRw/bnK1xWzIpRJTOUY03+kl3ziBgEsQvMwo+5X5hp6f6UVzF
IdFfImGkP7JgTFPGa/Ge8qRp0/ef1F33d9EVrLtYxqAOFJulpb4D81w9sd/mmpRW/aIx+tvSdEl+
bjN9ZRwWeySUcnQsOjEcRFeDt6yevlgUxyoFPg41VDYopR27efZCWYV9aktT5ddk9VqEeI9toony
JTUHYpOiBWat9lcNxSTLzGjUSfWpjJgg12mdzJZG/KoivoXt9f2kzRQl2Onx2O8vtC1VKKAUBhIA
eB/EhBfXQfJQ7FE47UAlN2Cx1ZytaUzOFaxB5KGl8gn5/RaQtOqFWZtM28EAMnnrxq54wg6YCul1
4I5JzyYFWXgcBwyBL+HjNdarNidvwMVevkkmPgHDiHjL2hmMjdH4EZKO1hrdlEqojUl2Mu/pn/zJ
OqoMjx1orv7ncvdKeNvy2w3xITRJnlBNG3Mf9+Gy97Kq3QsdO1SqOM3aOvv5PH19MX42M4Vz6bbl
+/9gY7Wl7wzNDSZNZmrmmcoNywC+Kdq1dq2YxaZEgp8gqW2+C06Ebf38vk/fZWENShYwoYcQEWsg
8UzwKKAu6/F+k0iKV3bi9SYXYp7r2J/sPaX/ge4mTH8yWTvOPZQqlvd0ibTdd8s8KU+s2pf9ZvAl
Y+L6p5zdtDDeofWSdkQuKo88Vmfz7VjsbaP9ToRpZhDWHLQgCls0VZqLC/tMg+tiaBp80m4Y0NNN
xLKtv1g6+If40vcFYYrDwJoMl8jtdP6qrjGmGqfQ+QUeKfbbhCx9VXYw3E39KhKq7Ci5b1DJOa+u
bCjk8C3eKMCl9QPuiuR5fwOvaS/L6Qb8tHdE7eGVj68JWMBLbOqsuIeK75m640qQI0FJTpb2jCmS
yiN+mE1T6yKij7TiT2Qt3F/lPmUfvRuGF1Tm2VIE6qNtFQg3EvMslkKGOnaIroMpzudKXPBM6DTF
RqpawvR2dHJUBuCJsyaca7D8CG9KQm3C9j2OQdALr1zeeKduUhc0jhn0d4pspUVkRV7JVfCuWrJa
4k047qKeMjW/8+HSi2hf+5SwGNrkgMk4YgGkSIQWtOgOXYrtjtND10t8w9CmxSwvB5NqbcXD7tl9
dzWeILIuQESIWXU0veCkEiXX++vohQISFa2gpaJ42WqMxRaD4HnqmjANObwosrY3TyTpUtMSAnAd
GHjHjO3aj6hRIuR5FTFGzitzPlkab0Ebaz2PPw0OoOUjU73dqaF0IqYrRsZf89jQMW4nBgWwiexK
pUE1Fbe3YRQEkyLeoYbbVzmeGUO/OkqLUl5/lPj17xjT1woda5AiwcBwRADIPD/3IP+cZgbJ4NBJ
L0Ynqbjt37boShFRsOWIjuRR0DZ9ii7H1FVo7OWu8eCnbcAt2F5SWUXM4yVlj9XwsC4zxz8oHB2I
XW0eJcBfnXDaGWkMP5dz+vIpIWyWnweCeT426/IThKqI1dOhd1AUjn0BXid2fXApk/mfXaAvxP4t
1Zaovo9qnhQoRJlWeRomSkr6uzN0hCxyJ41AWfXHCoy6nGCzujMbRliss9hY156VtrbIrwiLGeA5
94vdcEB0xWIVTDhcJGZKcOPnhzUY3eWGcJLJuwri6TQ5kIBLhSdkEHQM9U1gsse4kWrgbAZ+pWQI
uttMueG2PsdpVL0YfP+0B8XdKc0lU1RueiJ6c70Ob0c5kCkLHuyjhPMRnTYfIfK0+6gj5Ie1+FY6
bYJkCY95qNs13EZu7pStrUrXTGtAA4P4g+rpbbSMmT2d02cWhjfglPJRFxxBF6z69AV12DcvlB6w
BZ6rkCaO+n/UHXHWVftj3dCUY7Mr0Qor97JEF3c5yxSJobHNnKyn6FNII9RfeFbhBJC2PaV57dvF
+NHtFAh5KcOI0Mvyyv724pc+pBtuvwIu9KkL+pLa1vEMEAjlrU7BnRALPgGAFZDowgAo1QovnXJl
JJmH658NDfjbll/AozLKzVpgoGy+UKf3MmdynWUumEL+lnHE+bMcsGAU7JW3MfriXB2msRO9qFT9
AYfYtdZNRpvisQ0JebCdZ6ulC2FLdFGG/vzoN7kzgFNtSc7xq3/ezqtLkYmo5wmu4/VYi1IXCPL2
QAiPDH6xwsKW+Q+JbjI1MFCAVHZzT8jT2AvEbmsTjQ4B4xaqHefKRaQiLClA1b65sE90fv1YO+wx
X3ksQh8NOCvJrdQ30z3guhWRmwGQTIMirZ3DZsv8hHQAo/pFNkIrn+2rLw0N5v0WrvMd241UOB63
TZCJGHc4SvLSh+2tEIUYLYFWS8UvLLMXgUU66rEtsRAZwSP6k6zUR4uxquiBxEeU+OITEqogUPCb
1+KYuUdRlpcMlKsudek24Zgewe0WIZJ2iB6fjRjcDPg4wqTxMK9yav/eHOm5AtS1+XDHFoB/BddS
QI8bw1Cq5RWxSKxK+G070uf1ufSCnfzYYNzl8xrNXDuHFRp+HYtXkH72+BrYlio5WglXaL5Xkd70
tPhjyN6Wxx8X8elrIYDe19CFXiY+Qu03/A3eOHxcFH0n4fNpcOGFzHHcbtk/CJLoeWazcq09s0e4
fH61V1YevZ4Hba1AmCZiSPzYn2jxS3zKGxv6xE+/pRZ6S1UtX6uhjuwkKCCho3ttXSIfkQj8t8e9
eAOVgKl1ECUj6dEY63n1k2ceLJneqKBpA1H6iAVdrngqV36InAHmzvdrkYymC0YWXSt537KwZr/u
7dZGNFvCdbw6PTn67qLr2s/BlDakOAoYq11D2Hm8Rt/dZUZzEMO8HQsXmJxwoAw0IQ7Oi/i3jhWc
bgHroH9wgPl38cNgz0jO/6d5JckGIdQF8p4aW837krt1DlQsWDkwfjE75HehflkomY0uFtk9UKGC
skH3Y2wk1beICukIViMFadRNhkT4y6SEqx3zlvDsMRm6uJ91pandNQn7FUzzPHt/MdU6xJWCl2Dg
P7O1+zmDcWzhRnnJt9horM7cMrXTVomIsUjFGhtQnJgXKWzXUp93/NgFFQmrbMzZsvqfb6SiDdTe
EqRZZOCBYqUcP0gKpPK3D0P5UX30t3L+55z9lvLiD4w0bLEaiz6vXjXIkpOOPTtAb+kFyW79O4Pe
wSBMHD8DMDUQ7DMEujfZWQYPUOHsD3j0aSwxbb4SUqpBgvCc2qWXSqTwx0fEp380JkvEkq7u1GmS
FRIguv2jXxqIfRPiCHAiL1+SbBwi+sU7OGDgaWdGs0itt4MoapGQtrO/h1Z4APFCL41yWX23CQNT
OC0LSQBxg4xqLrjCDw4Mmc+Xi/IBmK0xP7j0F7Wt8zuJQnO9VhGFIBxSa345eaQ+Ww0hbhlRPaTm
feeZKxaGD2fqngObRDw/vwgR6arPdl3z0QQ6PveW+2suk/nh06XJycyfwJo8QlDK8yzuhx/zS/qa
67yKKht3KEWjhbpIQBpxyiJ07vDLZaSXCrvraUw/k2zbLuKXlxPvR0shWVMEwiXolX0eRliBCxzV
+YBGpTBUYVxfU7u0bSvc9MGoCEpmo5r80hVmrzkeCo7FyONbK8w+46hdsNmA/UtJzm1DBo8W7dsK
qiczovLIRRiY3C8dYWopf3bu6zjSbQOJqnN1oUBY91cEyOX/tPH8ENbh8xBln94q0Ad8me/vbcOB
sT1L6TcRcX8N35qVE05hqnjw4W7iDgYjQKdNIdM4tqrQ8kfS/DH8Q7IMvAhS36Wk8dzLtDsJU421
q0gNWFNAj9sYJiMy6mwgG8V/ougb+xhHj7YGC5XiSMoTlo/v2QWwODIKm1nETr10mB0uT0KxQ6rt
3qRkaZPqAKvAh9Gj3TTFqsJx2PqQKYjouPPplduUKAGA7YW462wK6TUdkKhZupTQClGw2kp4t0BA
YISmbQMZ2o/h+epdqh9Osglasp0IWio57hSVPP3g7Td80wuNfcJJarRYJa4M3M1TZJB9YVaVvzVI
XV6O1LJRvkui7XMV6VyDGTrhJM24ZJ0Axe0gUP6MaxUiAqlpUpFGCfsGNpthrxXrmCA1N7hat5K4
toHAd2f9TsRHLvrLRgXa7QnCe5RVJihMSMk7hRFESdkvSGB4fj6SwcYwKXcvi+gai0rXeEasbAfc
B1QY0L8l1LDigBpioxLtIJy+M2tAZPEwtB75rvywuEITaZ3A7MmXmRoLuFjZYYaTLFiP1hlxN99D
SyAhk/Ueo0z2r905yqM/WXKDnOmmEvv83PnqOVvz2/7CZJ1NqezrpmAeQY/li2OmXfzcOlYFvsvo
GaJ8J2b2PqQoHdUbHnOiACPXAvjDZciqSl1YOgv99ndy9iyC9StYcFgm/4wkz8yvri2AznsTv0OG
3b/MCSb5t9MHPjxTNdwXlXuxQ8Kf5oBXf69YNOIDijZ1VmT5fOzReb6hNxaE9E8xn70hJwcA35Rv
i0J75f+kI43bGrJ6H83n1hBhH0zEIB8qRm42Ir2H/woI/cJnJoqywduwwNJS2KIfgWH3KoIOyYx1
89MCJdHIjT0D8LL0ewQeB+CbooogrIbB21PE8kzOhkd85lsFFjSlYfMm99A+XgnqusnhxVy68+oE
3oeUJzIV4oCF3HAZDJuPS+Qg1luX2g8JHEtIh9oxNgBs8Laza1ZC0jEuQhjNJHDl6tpZFbzbKI7q
xl8Xjwq8Q+nSaCMi3yLnxESB0B6+KUGh1J0YRZSM4tfVqx9etqGoveP0SUWzSbDyhgJW7xuZLjtT
uqV/EfQBs+FacQhetwJL047B3AQfOWKZXg+BmiEn8JiXcKk80fMdQyPJivcXEnQUzz+cM2kljfoL
vK4ePlP2knw/pswtHz1DK6JvsilpilT3/cQUy+Ee5LfL45kHT3X6OLiwqTEJF7gHKJg33mF9kk2F
nhOJXSDAsoXRr5N92U563vyJhTQ52jrNmhH3aPVmvfIJl7eiQasBcsj0+LrKzqleJH403hdcAqIE
X8znHy1+JWYEvCWP7o2fuLMs39fLWrYrmp3H6nhOwmMcWFda8bdRLjQ66SiglYsSCdZMB7sIoqgS
70MxnZJTn67E2PQU9zqZYRJfVnN5OPLHeOAH/m39w6RBQktGmtnh5ez6on80opGAM1bD6eN8sYAC
HHtbGuP2g4pIS8D3vf7TaXRe313Cq/hd9IcDE5bwVY3nL8NXoI4ehz4kRYRvBVCjtxu1r8dotKga
cdEUWtucg0E7mzBmesmDXXZNTcSY/ehafpgFpKty8Mpegw4D0LL5/ApJFm4l3L48bb6wrBgbTynB
ErH22CHnx1/3Vwt+p9VZZKWQLfNkqgDERx0sj6p9xq6f5vfjRycvafP+snUjZuNbk/x0ymZ0N3a/
8b3Qy8BvtCI6sFf+cVoR17nZxK/DPDGOnJ8oQ5eTI6ckqzhwt57WGyGhX6+tgT/anmsaflcUbVZ7
9Q+gKzzFxe187KZ4+/UhkzQqAFwgawts7hAUOfkXDKLMZki11AJCBRz7tqLHPq8kNpXz1AwOkQMp
F7g3Ut0pqNSR2zCMOB7YI3BZgtO9BIHBQg1SpgyoIcra51uX+rc33LiLQlpLa8Koiz5FXx8Q8cKj
NIjZJVSiRW/256JW8EKrMv/RixkVtlTZuR2daPYTL1qGfVUo8PZxLa1zX15S15HZyos050froWCG
SgZz9UIOXDnhyzAeKanfdYBHM7eifeOpWUTT3w4OYfNleSP/A5Y0+wTUk4M0dHfrdn5SmFO4Y6wI
ZS0YBU3MvkFBH6BF2Pv3d9H8+taK55D1Gh3DA5UrGirZCv6aYx/lIjQAoIWDwF1r3PU7m4fihiHY
PmDSwC8LMxgVK1c1wjrRszvfqLqrtkc5WUQuGwmlzufhPJnb/mzFry7aP3Fx0mbpfgoiDFxgoiHZ
Pq/40sZeQhBguE0qghxAn6+XA6GDpzubBae8WBf4QKWiSpaopMZt/PCqSLCTjn9tWcWHpLDLUx4i
Buc/wLG5riZ9mDaYKqL/TmxDXXxgT+KJCFwq54vr0+xDE8/K9qZwkqOtzl2hTZvKW4fLWPtA3Ddf
gmsMco3sTu5OoTZtxRRhQ7VGVq0uo2zR19PPAlPq3v9brFX+DMNxvXveol5SaNAG2dtSkDejjMCX
y6HdwMh2UZCVmMwjVN5ubluD+EwtRq2T0MpgmbAD3/5n9x072HFjSp8esnKouQSN1JiI54YPv8bG
IEg2+zFLGfGrD+6O3aa+WYx1918HWlqMLpZDk8QjsVVYsMyKkngtdQ/jfsj1bloBkWkF5aHyYaXG
RMqctTAytieMRbIHDPCV/+X/GZYJTZEx05BR8pAeYf8U1JwSfKDuowiXi5QMPLxComjStnfLIWag
ylSibC8bk87LJX+y3YPNjMOu4afuDQTcARlM2TXMJgJDMm0jO5er/ZP+I798F2xz9JQmSHkQyLjB
JuaXvj1Wz4fkYVP3tXcD8jXU4yocx02tpLb64YDNKg6+qKQi56zKuEGKeUgZa5KxAqf36ed5Eawn
CVnHUQ53t7OYAwJkYXIzIi3EFraxmwR+mDyh5atlE5p+Re8c2IzQ54RZo7G58njXLexVsGQTvYZ+
TYfLf/yfDqoCOM1a4vE4kQTgvhYqlnKMEj+9FCKUXhe5e7rtxNUqZc4JkV9VJChIeg1FTFPon74m
IAlzNnzgKFfZfFYRxm4zXScTC83Y7rMDntJXnf9+U8p5OxTxfB2AjP5rL8Y4jCfdP6X2+BPjAeFh
SPJu4/Iwij9XRx4kfhBH6l2oeS2ZlJ6YoBylFjhU50rcfCDIvj95zN7WLCiOh//hc2sXqjIrllKA
0m1/lReT+ISaty1TQibKJkVRQoD9JgnRMombRMGR0Y9UWF0PIM1+YYz721d8ZVaTS+FlIUqUCOKC
hi6XLTCGxviL/XLvPKBjOihBeGAQnudF/5tApLcWj+YwlxBWJBKbYUokXWHojROYTgWoGRcvHqkL
HgduLRcfKyOjurlfmEHXM/cBuskuASX8xbigYAaAyC/Rf5BId6iNBbJCUckvqrs8buTEJL3N08Eg
eWCtdfQOfn/2xoqm3B3fQtAO0woqW2be35bBBPkTXzH8/q7OEJQ6lPiNt3R+UyK8zFBpyNcXxKC7
1/Gxrg2DRpMhFHF3UaZw0Yzi3kgnDa+1ySrcfhN9Ai7dtxYvkeJ398bG332UkfWKn3NWzYq0Yvuk
xl0Hmgg1zCgpKpfT1NmK3koD/WAMaAwSjH1lTHOrb2i05NtQvaOMzlB1NNBHCItWW5phd4NqRdI5
z6ng6CjODamVJ68EHbRyiAn/U+MdW83n8xOcAgG+R00nrJa7qnfibTOeVU1ww+YFH2OS8GHmUCHh
wA8Ly8HKPGX4Eq5ghRnOjy/2f4t9dQqQAe6ayLVXs+BqzurxG5n5bT6TR8ivu45Lvd3MGCFDk7s/
g8iuFHT7eaeFFkgAOblIgiBa48GJfRVqcvz0sdvSwtnxMwG5pRQxM4ix8ZYm9V0QPemkcV+Tc/R2
Oi7It+7hHtofjEb9+L1598tRXxhc0FfPWeq9VR3EtU1RAXKIe6vnfdwXaMnugB0+IP4fsJYFQZwK
RxZqv59UG8sQL6Hmx4yGjsUZ2YTAIyv44fWq+Mj0hbXjKQUxKCXZ6s481z1UYu5vXS9fnaTZmjof
rGC66nGAKJ9P2/tYbGu4S1l74a/TzqI8Dvlt/h99KN3zZ49eKt/g4hfSMoA2Pawkp+lO3AV3nqzT
DujY40rt71WIxmDC9QLG1LFuf0JQ1KRXcQnAnprmtkKNBIpGW/N5b4B4xD8kArMjvWk1KiqfkAt/
6FLNvyF/Wfma3UuQXyMcC0u59cN5ZB1YfA0OXjYUfYr+3Ihi7RiY9rCkAuQNbKJhFAtcZM9QHSBv
H1zMWPbnPcx6CQ8Cv7YOujphFeYrK0BpU2XJntgVe/junPyBbDcpzEqw7YcI3ED3QawmXkqAon1O
to0josB/MiN70pj7UctN3IRiOPtEAesLSlkFhPm9aa01F2jVx7ZlMVvrQ2cLn+be+Gc4fViY1yhQ
OtvR6irISH8J+//PI2nqpYmTyHr6baijkMX/jCs66py7HUfz1x8YECxDO/TxXSQlJHSK7HofIXYr
Z4iZLsP04rCuX1FotwHIfJLnAHpndEeZK1MOn/b3OF5Xko5FoSZeMHUZG7pHW0myuAORT8uNWZ+U
ezVa7tiY96wP6JWaw0ko9/cFQvL9sN8oCRoSyqBk6/ryQ8BLtE5TqqV5YIFmdFZM8LUL9bN9Zyl7
B/GKPTb03uo2qm0JCyPK13wRzB/SkykpvyYXVLXVhIK5ucEY7r0CL1E2QEIrYVjR/YuPJ6MTKVKp
wudMxSGZ+YU43ixC5WiSXAw5OkDJq/oDpPjQ5oO407PnmBHM6s7zsh6YR2Zea1VdgdJw+eJBVJR7
dG74xthVIJgBLLjfsQjExAmtuntWp5y59DFyzXgD7jzcgvV5j+P8d3dooizA86YYtRGhky1h8fkM
HsDc2fF0NnXQC9svO10So2kkkca8H5oVv1neTWY15jsDtm4p7WDK62gZPoelU6APr5lSHyGLbdIB
Hv0n5I7ymMATgqh3QepvwWBhrGwZOCyDviMv/wYalhArsocBY5MbE60oDPTF4RX+XJos/XHtO7wq
mY2V8a/8LHq6RkGdVrukjSbn0zI3+eJ5M8b7Q4pOYX8FQWmhPL9lJTUa9pu2HXGiad996ywl9fyH
8xlmdJWfU7Xjh5Yyx3f2ahfNDTM1vxf4CBeI/M+5BRzGIW/9qf0JzcxW9guVM8F5n1DqTwtsiZO1
+pAme4EdCy1TyzboxZMIH9ftWC/9S8ED9z94mW75Ih8jRZP4d+daeG0+B8paDiOPg2Zxx73IA5Wb
rcoRgX9/pDz8udaNveCK2S+rw5aYu+ac5iIQiwy5pr371q0f+u7bVLb8RMFvueVP0hzxVKgzNDfP
eDZqtCvDQIL/7mn1QOjk3vlJC8lAQ9NdBbdVgV0xsIuEi58+Zffqvrp+gyz9rXQ19yZX6+iqXgFF
1ukTdijN+vWuagz/cGdqcssk5bWmS4HPFlwIRRZc3Z6P0rnIt03GkjSGta0clV8SkSvosENJVr4t
fULsZtHiJmvik6wDxANs82FN+nw9HkXXUaQHN6LmeMhpHy09xxfAMC0wS5TzI93zY4eyD9yL+/Bs
zAxX9ClUrOvVQtoovY9+1v+FKv8LR9HLgjuDqfFSGG4VamlWpK7ZVZ7RMNYW+9znTH+4/uiHNPbZ
GMcL4Vzpr4I0n8loCTK4VUi1AEErLT55UQRR0fqJb1Hyl9yQ2iRykAR0yCe/ZtIjsoI/vtXQoICS
OLRRvOFqo+xSBKPqoJIm5YN2+RCYhS0T66m0Wgq0kcKMPLmTCxWoPLaq7Kz8xRPux51nn9PzDSQx
DmUgkLIT/jJ+38p5YHg0Nx16Br4LXrCVX0COs4Qj36ETdv5us/xetrzSMELwwUwLALtSv1A63XkA
pL5fKdsNJwXUv0n6Gt4/56YtaVfhJcvt8q4+5ghT1GR8fE4KLDQRcwT6HWIpkwqP2yAJ8XvC7YJh
Szg5xRWgBQUUpKUHXn2lMoAMQTOor5vme40IZ1XeHHwhCgRJQVgRfk2pLTT+QeKqRG8dnbUdyLZI
SSE9sEZ3tB5S4722PWzrykqZlD6EzzWAMVKQkXee1LcjSqkE8lEQAfmXOBlWBbhTez7Q8qWisy7U
DMUYytDJuRjnLEuqLnGgYNQZwAPuK0lRP3ftTEC6FK7GSj78oX3ggIMfkQkfviGvI2PZgEGwnZaJ
On3Xj1gnvqR+RiSSC35ygVaze9ETaaWjSBD1gTqyqMj1Fb8c5+SY9InKwpsSLZDj8EOxD3s9e72T
+ju85xXsiSpE/JHokTWbhk9fch+jE6/4q5/NPMY0DJrr/fzIk7PWOpFvOsnk29q3pbEOfiCHoziW
CmPLQtPwk9bOWKO3PTgqxxDK1NgWkPWZWvAfQPzp89IGdcXV1iPm6VHIayHjKp9FlTxDj4JnVR4b
EWP2KejW8vvxP4tvA+rOiSarODXBVuJqGSrGPvOwMgu8y3vAuF4TXSf/7x0JBKGB3F44Ki/YyE/h
kMCeUbcWR+YE2F+05/tP1wbb9E3YwsYsTtaYyS+3xavpqx5XQwFqMt79YVmyMOcUfR5Kr6w5Fkuc
UCDWc6i23xn8nZN3i0lhmc9GXPQymWkOVpGLzr+Ub5zCy9UsrIg/pSdUb3j8qmjFEXU+LvMGTYSf
wOBZ19V8yuuD23xdoy2YPEwHBexe3d5x73zYm21w7lH5QJeg5RI+YpyFo5fynqTCIev00CB1YyFk
4eL1ffkbJBoxQLGfvT045d94/Osc+TsWCBwkwMu+mSz6ZkwKbsQxfq8Xk+hv+0u+Csg5NLzS+b2d
zq0twczgPBJIFMNvYesN6Ztr0B95NqbYWOULWZDZKLBiahBKyryq2oYT4tZmuvLpVxzqD+rG3WAo
9E2KNXKH8rnHUX6TOPK/ixTKUk0gY/dHx06es+ljneRJoEzyBtsXu7XKMPOczlF/+ltU6x4AWRzu
wbZ7RoRRPSIneqMMVQbUP4TyhhPCgU7gHUc4uf0ec1Ky3G0IqQvxmsRCH0J3haSKdowzNuzpWzSW
IXrf4+fNrn2JiPK5y8680kR03pml4Zi54a5BCRyUVqOPnHKI+JpDDDhLozezApdEyil7ZSNOQPIM
ej+OWiJc8L5mEwIw9mFr3WLOkeXvysO3seuPRb2RwKbr6XLeCHW1xfXyOERxDNzx0ybWo99gkVzi
HgB6UsW2rJ32is10sGRXHf1S6HzwtUfEM4oBjPYJyO+EVGpVRIwC+Dkwrg4UU4hY2fmfLGCkbHrk
qNcE4/NxrClpYfja2n3FTcvM6TrfAHFq+YEilNs6TqOEm6IVedrrUxWM6S+pKEWXHWTUUAftth5l
25kx5b4dMbxeLxCdWORXN5qdUJRFDkqBI9yz/vLRWjitReZR+jcZuKMp2F5FGO8df2etgkPqJtLD
rmAJlEI/UMrPpFQPutr5QAIj/OMxv1kpwLx2g97Q/r3iRL4el3i+oY9/MurulQ0QKAfKFKpn9Fop
xztRPiqv0aT96yN+6zTKaSd5cQ1O3byWWMBmGqszUriJy/6dgDPaH13MvLJRJj6uvHyMYzs4zbNu
5/q6vK5G4NfWr015ZW9vz6FpoD3WwCDfQ3esmkdYZbLjh39aha7hMcQAeDF7VSZ4No2xtD5TTTu+
N8g954m2rCPefo07rZoQ4A3iZcb7HKlzd37pd5l8fKkgXCC22s9ypdDhj/pC7o/Ev/RV9U/1xF2f
GdzgfSZc05j5r1+efLWrX/iQBvy8ivqYPT5XTOFioTkmP/2SfS8p3knc2ZDiegWtWZyUdoeqYW2N
DlrdbRkO8490DfgTdEUyyPDdilbzH+6fN+1AY2+pAC/mV6u/8lTCyaqC246pR90S2aYxpNTd098D
BeYXj823CaNB01G8ATo7YOWzjVYwSUGTaaj5z3Vh1C5jmc569yyxtaS+ccEq+mxJ5ElO6mYBn9Bq
hmGT3vLXikOajl1aftYrZ3ukY1xu0MMWsva4c4DXNREW6EqyJS4eoeFxWelbKiyzVUId6AWzOa52
bUHWv84Ivupzq1BJHmptLiTEGisf0t3J7RYHncPcaQaxD1R35x4kSd6fEWhyApvUkNM6I4IqcO8H
gBA4nHp8fsJ/gw61t/B/IVGY1VNYM96Cl+E1VAkXc0RxGo5oA5fjWNIOscZe4LOar6SxP+aiNZMT
LxSeVt+HuNn1vsphJMEsDO/BKncHhUzXjZU99oJCUwWySoOrO9Y4+9Hpth2AV7zbNgaO/um6Lk/8
3d2e2WP1jxXmF5XVsKOwV/2Uq/QjvwYBKcqrsvO3J+Mrh1G5TdGpj4Ng5LaNv/2BsgQhyrY37HbG
GS6feksyHuB5ixS3pewYB+q2zbygN4ZL2TVMLNxKGzfjv4zz+iQISbiV6mw9VdSO8Kq67FN1hCcY
q2jbgik3VYBqMkCfR3ovD8HyAKXGKbtS7e9xELjL4eiNSQuP1DNKCMJ1Td0ekZTAFW1P/vf96IEF
wDg8kVQtmzeX5CtPYOou/32VdAdpsZ09hFvS8hchFSKmlZRgbijkh6NGFaPAnddBDAWOZlqUscqW
vJjsAnyCoE+88RIAXi1KsUadaaAFLs1YXMTJ0qTIiOw/U8yp34HNOGLSMUHJkA6lZuOc0MK3EzOr
fpSbW2hxv6uCX9S3L4tiZ+kPm8MnR4MpNBhaOv8QLKzEiHAonUCqJXiewNEdekt1fuzeCR3ygB6v
Iz0OuzN9HzlkkROfpX+HdUQFScLHAQ1VjOlR2Pt/vS8fiGHPMkEtory/iMVfhqVpMfYU0v5/3SoB
NzHjNNnGuP0nvOa3VOhznI0edEn6dNvtD+/Kxx5HBco1r7cfyagbfaSCe/EqsdV5ppje9Ep4Idev
OG5481gMvbWCi/XDoF0NJpLK53KFW0EFFZQYVaV3hQCMHkm/BvE7vYfCDo+QsgneZLQ1rzXD9dUi
KT1R4AERELIDaF3M+wLK+3KSiXtrM/nrLEkZfS1+SaHuxgprqPQqNOvt3Mbx5JwJ3ThHDRoGdAd9
IiUDwcsrBSlU+UYP9IGTYY9KzbJJFV8jGI014iI2F0PX7cZSHpF6nGn3uekdPED0j2Sl1SF3qKd3
61ZjGhY+6JFtSEwbVCeM2zyAxVTx8P38AeLprZrw7Ew7Q/XrN5aHcpR/EHHvodISjpd/JKB/0GRf
YNoVGSpcb53p4I5rZnK9apAsBQy1+7ybNDcp3+7hXpezOpc+FGdttUPOy+4rKWnM+MhA919WuIRB
bD74079biEZ6FH4EbwKgTcdghVBI1gaFfQVG04y7/Ksj0D04KLwnEYyvFNiNxEMATKmCJmebBqHM
Q5pblVQ1nhp072khyBjdsXqALz/ENSyH93ucfN+KuiyzBGSnh6jHQsBUVQME5ov4EBFFIopJ5qAn
PZ1Pz75hXuLBdEdm4KU92I+iZ0dFnl13xWBp6yFITRPu1s2szKFWjy5Q4iJvljtHvbjnwep+flWY
8h07G1QJMFXe3oEV2D/d5t/CpGE4qnrtHA1GMEk+B4G3c+FZvRfbZ2ILBNwgZjMBFMPRxsL+HOkV
KrQL+8X5HOt+wdAqwbvgR33gW5qZz1o1ZyEpJcjU2ckBpD4YWVddhEASdpaGw52AI4t92I/Cx17D
u1BIPTr0mtWoPpCBEfgPnHEzJtHDu9x9jPTXmhfNuZLH2m6SnVtdazuHdJJu2NDyqSUnibTx6bMx
9MhYX0F3oDDhmm4oIfzS52SAbTMXKI5J/5k2z5nqX5fi8+4DEZo0hY9eDurBVnpjPzzymnSEkYBj
lRWc7kKN+a9PyWoXgyyZi7LK+DsPqwkwx2wcQRJX4YtFBqx/ZKjwanTNyRjg/u8db55ThMe9mmIF
ZZMkjjSVsqqwodgLXfNor2kLsekfS9uG1EIzoCVtyltvx4oM2HYmZYaWwZ1rKLvnyV9p+AtxAAwz
JV+ut+snvOAzrVoUlQs8M7AE20hthV/AqFKpI+nbtVpgkCBsf7D00TEN94TOCeNNuz7Eh3SANC6u
STlgNqm6dcS0IJymkNle4kJ46ZHeysvRVGwGbmZe28CGnMn3levdVD8KS16grGXvbcfU9OGs6U6b
jMjMKj9dHfuf/QUs5/nNRcwl6pzKRN14/4xQj8/+GFArmkTdchHfqfihkOfUYnsSJtdAQhfl2zeV
7vsd0cwcw6vb8BdcxqXjx5nFs953DBSb5Y1mA1O3wY6fdJvzucX6sqg3SFYRCS/PYk5HBmZ9USW2
xjVTXxEcFWGImhPDNjWY+fNMnNF+h9Tj0ry/xe1kRB2DXUl3cWYS5mpxkqNSDE2/6ruVtc4FGp91
oDJkhb+43tt7j2Jw7cn/o4gHmtvXdo/Rp9P41z2AfdxNdg43zyO19M8KdvpK1bQh3JgTZYMnF/xi
+lO7uhzOa4TSTq008/fwdQwOQgZ+lIJ3+mlwXKye8nM4rdOJyc+4BiJT83v7NPWIIY4xV7tfT7Bn
wY+ynmHtojtsZ4t/sTL3EkD+Pg+AmhJdnk7POepvvm/Ry3MaoEYzkkKJxijWYXsqt77K8PmxgiqO
e/9g91MY5iiRKTzCf7Pty1e29bOUkttShFZSNT2FPR74ezDf8Xw3IEGGYsuO1dchb+7/jWMYCdvt
iviOgkeXRnV8qoxgqwlrTQeUi6zvrFCjiNVicI16/scjM0jUUnroDawkvTgaINdeVAil94C07j9J
Sxp2NCdW2Ghi+NdfLUMjYWrEK7NLq9d8EpbY9cnXax0avdTJplGCtMV+UjNq2mAvJ8oyBxchwsjG
U6j/qLSVgR/grZ5vjH+yXvkOy2w0zfBXbxc0Km3HUKOR2SoXGfG4FS1ZaBGRuCMFdlEMnYbYA13H
77msgjjJ5ci+7gbJ/WADCkuXv2eqW8d+NB+GC6hysuh0O3CzGwoTIDsxiiXY6m+N4HP/Miinb1Kf
p+jUzzaQQP0dRWWxnbrO3DjEPSRn7vOUUV7g4dFqxv5jwFbKt9fp1osf7Ov9TeJHzKkfHraZg0Ly
0wcQ9FMvymml67ZuuWEAz8RjLsPs8dDGwrvha8YyW51QToYTYIxTGJyT7xgUdysitTv11ykde3R+
RgiDX6KEchP0/LovmUUat7JLbOQyjqCi40NI8OH/OJ7W5XFXtrCyxpTSCCQuMENzCrYYHMrfY8Dq
FC2E1eGqzP4XUEAmYpGwFmolv8OywLU2m6qStPpacbgzmZR2nsPht9FDNsDi5XG5IwBdxymi44Dp
i2Tne7lHahQ8a2nvWiGRK2ejswOAYvMSh1DvgIVbFJTUeNbAsv3p+eigVK8T5ZdrWTpRiBv9a08d
DBf4l7/M8LkFjW8xs+wo2ivf7Us9wMkskHDFJ4ss047f/EayPUjo32U05RAJKVfn8olh+nTNwTHY
YO35u+ROmWvnn6N+qDKztaHy/ia6Qf2ik4m9E3bqu+/HQQzsUffjdvrkUp0kKw+kncCHb+ZT0kI4
4ICvTMPe3ZFn06+GxOaG6b6bdMf2DTK+cJstvH8D5/XHRoygNMItySPaIAYDEwEPPPcvFL/QqRg4
A662ak7488H016U7/kpQahQ4JBIuo4CJYS+FJcM55GFlHH50aXDcDuVVIPhn69emxkFTkLKXjz/E
R3PvhQlvM6YTwh3e+swiNOBHtloWl5+EKQSX5EqiH8UEIvC+XEaAUWq3vPCLLZHvDkqEryS/ilRQ
0/h/DLIfnIISgkddiGXJ6XGwrpvZS4UX2i4r1WZZ85kA9am0ldwnut9g802hfEl2pYCqZCdAQQ4N
JQixMrNAL8U3AMYnf1tnlmW8C/jPWr0cpZY/Ho+6f0YYmnIhTtISMw38Lp8FrN0/tx9STb7/+4NJ
S8Kp874NO/r6lIqUfy+RkARs0JjN1LfW7rQn0FAZeIRNnwgSZuZPEY3B8agxJwc+ZXixm7hLZt9n
8yX0K+QV2mzl8XHh71uOqRVxw5Pcdmg8lecdzwp+ldE8F6MYZsiG45tfmoXl170vqt7uOW+xPCSs
/E3V7txEoDhE5ZcNmB2afzXymK35DhtzFFuoWjhUhtrtMkKFkpiEsBf1qAgO3wWP1f5dQ03qr4dU
yacX4qavUpaj7nurlaE0x+9i5kDTflKJe2oz6ifZ7lSNvYzXjQRSaZigZKb7xFQedyIVliy06/dr
DE6AGhqdHjjDLb2Tos8PzzSN7YonhJI2kg+vWI6tNifpkbaVLOgna2fdEbnV9rqDwU+d0RKPN0xV
1IuBc/vD5IoLUZxWGPr/6CRKYnNd8NwbnxZSY3TC1S4WNGBaHpq8ClVnCOCnGIyYNQ4KjBSmpNCK
b+DRgdbORMenoH85xHdGlM1rm3fVE/wmRQDXhykBjjDXGLVHnWJQYc/fW1oDp+DSUltSV/i/VSIK
duwPq+qoVFoYMd8+6Bsn3usXEYoMynbMHt0KL1WykBKyU/ctNKLoFvs+4tw9cjB+IrdJllP0YlGT
Et/UYWaY6XDlpcUxalDQl4haHBshhHrXBo/65Gjg3nUN1DD2KH5oC3Iap5Z/Vm8Bz9sbsIgXU3vV
N/5Xf5CgVkSZhJayfUPDjN1NCYw9CZon3XSQI+uPpKqbDqanYosVIOHYguZQAZ7Nj7LY4gpA09UO
+wEq9fVkevgZnBr2GgLd27mpH3MsyQqxol/TMRzVA4nKfVWQaTvfB3rEvjswc18fqJwFqGKJG1A8
EmKV4qsouQBurErQqVGi0TtzuNtnk78WpedF8jp9OkiwbJB9jBW4HsP9Oe8FV2Hpx/h3/+BvyhVA
HpzzntfQlzC+KxHwUxJni2wHWcMNVQoS+iKhJjnsVq3dMwpXWnP8W9+AN9Enbv3jixMTwJa43oc7
EwdQidZsuU917QY1AmhX6Nb4rd8ms3n8TwKTMoOH4Xaz2u21gJDjRLP0Y52Cx/d7nunje98CJ9wS
FpkNiZ3MNq7LkjLmSMPlBJLKmIziI+niKi/HnkLtggHqlkHwFHQmoPNkW5lWuzi47PYxnH8KJGOy
f/lmw+sTC4TtpJOoayqx6V3MIkjpF4t/rw6/NdJcZX9tsqSqVuavzWfXJld4K4PZ7tqFeYx8pVmh
0fyCRLO37pWs6342uLdnCnzefyu9nuohn8FSI9u02gGOOMAuCJOQvH2g49oPP/UdEthtUXjVXxJb
SrIy2GU7fgZMbwFuFLrhE8d7aWU3QlD4x2QBjO6vvCIj9VrZbVHH/w7Ws8o30a1uh659KhusF7qm
TjOX3gkv9h7IOhExPTacp06G8+TUN/pcjWgKLv8chKiJhsk1gnhKxs59ZxYqE04OzwgCvPeJHMsQ
MfSO2DYo6Dc2LWCL/WEBRxoMJIYDhm+p/+bI+ND11fp6tH/Vbi1De5YMOyEL+C97hH6wY6mpmoyg
uiOs/sJctQBMECh+a7a0lY0KGUIW6Ye0K6u+CLZB1gChj8Qh2KdpR3dQH8iIu8OxkXyN4OkvmhFc
YtwNbVckrTTxxWCembtIM473Pwz5bKeJFRF5ZVtSXfF4aD1BB0LJSrhJC0yLfpD4RySsw/ibqRgE
1amAj4kgun59KzOWlT61Y2EPSHdFKaoatZdLVQA1itEaetK05dFgG58/uG47Hfu89D45ZCVm8sOC
f0/lOvyYgUbTJaCTnUH0lUooYpmoQQc/LqwRyGYKjxxsJTOJbWZdCZ6wu7YOiCUJPpxdzRnMMkQR
AGN3l3YMYNJbxopfj63elxbqNHmp8WIEPS07NMwFoGFaIscyoshu5Y7dLk1+n+ajjJbma50F3/b2
22ftpL4wric+vS7hxDACfZorjoO+yPt88aEWob++wYCKeQWyrNcO3sJPmNvLuH0SBQBdvDhL9pNt
VX5wpSzSiLy7IlRj8nfQ5AES0Bmp5lLkjNhRx1Zay8o6uLuN9svziPIKtIfkSobYLe1mo4i6gjPD
BVPqYLBvoJubcyE/aas05dve8GfiL28fU/0r1zR+R9bfaNLNRLkghz7fEFUMn6z5r9//JmV3KcIs
8U6X2GX2LX1QlvrK6tiza3Lmg2lSdGn7fy/SpEUDo/gqnAlkKmSPpNl7ph7f8IeNx5bifDRsCOZ2
19ZZ7HURfYxDPlkMD5uTSLSklY8itk7Pmbkkl3JWDsDJFmnzQ/CghgpLl468iS77enil3LsC/vxB
Hl8rhu45+kKWLdAbEfCsWNqGv7RKmFWrl8f1oHtdmpZRO6b6tV6fVIeS8etVobXjfYxO3211vPml
ZD4Mp/qvPi31nd/4Zk0zhgS5aVK/vtdgsOgytcWLNeEzEFHh16rixAx/mmI60/OYQ0KvYBgWuF2l
z7sqO2S36Uu5qr+CMhtq9INCae6PeORWux6A/wWaTt00eZsz3qzzU2U1c/5fFm8XfMKkWzxCqczn
mIv45xbKZxQxOp8nZdX4p8lmERAtW1JPEku6Gunemd/E9mfawGMJRNYXYc+4ZH/8wrWsI0vl3QDj
4QK5aNY/sSkc8lkjmMT9+5DNuA2cyQeu9+kPz/Ti7PMC7Jh31ZY81Yw0sA5jwqyThWb3Vplmwg/8
UBrHxmoLqDKBfeXWOcxD02MWvHGrO1prvfe/coFGODk8a+CUt544K2b0ukULKsIujWcuwptfICPh
0yojG2FOX2RdDV48LFQJsxHHPpDwtxbbSdd8RD6yiP1cPvHKE78vesXbul7lsXJVMaHqC8sjrJyR
hBaplhQRtE/ggTQ4M9+DAFK4XMlliGTsLuxTcI02MfvIaW4sPC5siDdXofO4aQbE3C3lHWqE7WvJ
xm09fiCPQKLoFOutgalGVVUAmAH+6Tb56FnPEX3//K74wtUKffT45lM2HWXPbzzefpftzXcIsMSG
yx3J5DrfTRkHmOaO6LQqLNs3WHKmi9JrLeUckPaq2u9L++/zE61nN9BuExMcsGawEWxuRtzpX7Th
LzIdnNJY9YIRtUV+0jyiPUdbe1NcaCAXMQQ4dYLZIq5rrepjUuvrf6oOHn3UDO4988pGgtwWJT5D
dV6ULZv64vJGe1ZVwqFm4skGtFbB8ZRdSpRHUvIEiLBM+H9LrdUNkiS7Gs+RUAk9UtqhRD8ssats
OyoC3TCCQ0ieYlefBhXB/NssZd2zcdNO56FvLord6ZN/7mak4iaXbccCz5jSiSUmXJXMssG1F+9L
U5iOi5xdbE44r3BZHkhueLTQC89bieKrHwvaf+zlo9e1eaK7MId6E7pDj+r17mNO0ztfxZ+q+mSI
zrLK4Ml0YaCzoNXdCFyeNYWZHtANWAHkmTgbj+Kcc5hg5/5HpDECNuxan5Jj3P2RiLf7l6biAydU
tcvMuhjYMUrdeeAk9h3Z5NymKsIlyPS5Epc0rt2oBL1yvxSQFV8FJTpxHeZmGJ/UnzY9R+rB/0IX
GbEbcfxDt67bLFGEtvA/xPaeNxezJreJVSo/PHreqlWT16aQ9UEBnrmOQRQ7D3llBLk6O6RQB8IH
am2RG4bN+4OuK0HgLVCcxYYnnn/p6Dj1/7l3DJqsqVSxAPom6Jy+CJApCjlmadSTXeKlL95FD6oq
18TK9DWqn20LJkE+LHUIcD2fxWRkzW+lZgGdaelTZyhBdxwO30xuyIUStSxFEJl68QjNZgzwSwYx
q8eSEFfWWULyd4HHiGWbRSCWhpKZWhgnwldsW+llIq17xGJaY8MzcX5QRrNGEImPGVQ3+2xuDe55
HSRWErSYoDtVo5Cfkl1w/sBiPvCHZJctxlRSPSvLtN3hV+OriO31GCITL8zOYIcG/ud3O0igqCqh
uhERbblreQ3R5AzW4cMPNcyflu/jzINmxXihJW2X6Edj39RXLdziTGoBuRXJk6Yaq0Fs/utkkJ1F
Zu9wmLidRbTd4muvw+CzMbfDxYQkYSnEYG58eOjsmMLDowALg0jMwOntrevDEhekw+7obT2qrajK
eIZTruCw8CjoY5WDovi+dpqE/N1RaO6cnjfjQJ5Bot1Hyt5hMPZtIvIUugLxHqTJzZYia/O3wjvk
Beay48n/cYLReHaMLCZ0yI8xcwT5AWSccxgwrro91QvdNs3fPqKANdL1/7mprpga02/lc9crgfmj
lymN0F25MMWqBiDN0VMZ/aj9nanejxIAyHW8HXuOw0G8EjqRvHY3EJKM5nhF5R90QRsBian6009r
bAfekoFEdAgiwgm1oFzqYO/q1H+gMQ8GumWFz//GlocJayBg5vPSrc+fgrI54+GJL4mzviRkhrR2
r0Ccm7Ow+AFzzMDSClog1n9Fulira2IkNxzhMyGiZIyxZ3kVimPc7zuOfIeAouB90YUKSOiVfc/n
hM50vjCYrTCJyJPwNd3tzWKAG1Fx8dPn++FEqs5DYR4dyMKJSzmVixb2QVL6BJUKvp69D4cu1wmY
W48+j6xZTB0qOdF45xWm4QxO5QtLicwWu+chaMq2AX4/QWh2Oyg7fhElefx0E23ZFzc3a+kD8Wai
8zue0iECqNDObkXLzfDu1rygidHzIu40CbSjTgndKw1kFOJqq0mEX16x81YVJW34z/H3YUhYZyQw
gfY2B/tFq09UwtM2mLZAXAByWCD+ATuBJ2kCs8mG+HleSrd2P7ealZtwVPpTyjhT2sAA0Nlim2GY
1xEus9/coUgsqIuq/yCBgDoSoDU7PQj3i0N1iy9ky7qkuaO+xd5uNj9TwhEJrceasea5aVXetdoK
JwCR+jkOsnCSMQGpgGLs/YsvAYmoRCP70z9OOzFg5UdKdw2JKxMMha4AhtOHB7DxwcooLLuIujHP
7t65czeCOUTJ8iPNYa7oZNN5MmRlZQXajv1CD8c3q+r1uHBq30H9iamS5nxTVVGZhKWV4AOY6XSE
ejPFV0OE6aZ253C4cxAhR1Q4QT3CyhFyg5WkB/zqe792BDzkGJwrCzz7gyKIacZMqhg3MrzW+LCp
UcFl2TMR2sH/mAu04cmlLYhcoFcIeKV9ZMBVkRhihiVsTTQaU9l5vjld/h/HJBMVVLGrBcC4cHU7
WMglFM8oczcWermFyDHxFUIYjghdq6TcvhKNsuOhfrDQ8LzRoVd5MBTwXwmm4dNFZfyvs0hONQth
MFqlJ9/rAT1QrwJ6Z7i41nd7vDaz3Wlcew5IU0QGu4c2Z+qia0G/SJTZ9QhU5EaHSgPYo4UdENSQ
7SnjkyW2qNO93mWXOGttt9eAoQWhk2UK/7Z8l9VjEgOiwBoS3BQMhMHCyCTTdXykD/OIHv9eNHpK
Ed8IFR86FWjviVCfqNSG0vOtdMI5tkDlJeub9ne7co4Z6T6W1KOYZcwWj0PdoOHeg/JCPebOgzOP
zNi9Op401XdiVGcyVtepRW7Yz+oUgD+UWTtNT937SGkrMnff2EaVScme5eaEf4a70zAD6I5s40DP
HS9rbcnbbaXVWsPJkY2JsBy6+1khNMNIU2njFISUBzN/L6wSGIySArxudb1f4oWM0y3NhGFai2Os
n7itlQ4dI/yVVdgdLZJHkE4CQ8yDOR90zZL6Lq/AsfSRwOKbpFMIN0exidyAMSYVQSP0R2BMm8wT
sg0V0XVtEEmj7/6Qvv/IcAT/02Lg+IBuPZ6yqSaqFUc9Gbj8Y+ZSuFECBw6/c9NGZBwon9/5/Dvh
NOlMexLM616r09/KukIUayCxobD8m28/5HWil8TCPvJMdmBt0vgwQRkBFdigJvcsOxLfwA2kGMsP
tMJUwDbdtxbusn/aJoYz6oVZ5MFoj53dXFL3Jr0ofUxWrdOo64SkzWdkwjFsmafV8tpUAzlYxR2L
Se+MBPgK2pnevrEWkPJ5e0e6Ae0z5XQKkXx3WclhjsCWxGhan7WyNGh5ZLc8NVcjYTzAEnnhaQJu
t7e4Jfeq9InFif9Vm7A9J8I0VTVZQ6226w/pIURHKFgHIvF40heQdWGQzQxhVcl6P77KhWPFPaCB
pKVLaX38J8JSI7sgacTRWeQwfG6eXexJXtCH7p1/p0tYrc4JfMPNeNpSh24PDzAo6ZcBDGwbc4eL
wGOdskhopYU8ydl3UDBVYQAp8WS8f5A2tWRDlRurlntHrAxzddWqk0+qbFQxmzC+jVtdS/OGFW2K
YhupurK3Cm4oWoPmOybl4lfPsIgr0xGMTekaX4kaiMVpEAqbNB/22x1hR5WYszigrNl6FpRBEFvV
2lOhVS8dzAf07vPT3xYDtONUuobpLWSyJ5ah995pT06+1myGAlGVrN/XT7ziFBqXcJsUWVHZXOv9
yt0Hw2YCfUkIZQNte78oBxLP4/5JGeMt6mGRmztgcRTiV55ujBF+gtgcGKn9PV4D6qBUlRz86tpp
CHN5WAcP1uo/w4tQ/lIb+KDtzUxWmmZ5SATVS/zsvSaQ27FpgvpgnJTiywDkRb//cowYC3np+klv
AEdAxEWvqNKMPaT9aAsfSnafCsjnhyTiqKRaEaB5kjQuiTRt/BBVf4+XjkoZ38GjIrbdCqio/CLt
g3mC1EFkhBHQtpJDrlAK2YiOKqklRvi9d8iodWB7B0E1m7K8pxcMQhuUPBYgo4Iq2VhFVbqlrRgE
p66ihjiTq7S9cRUhfRlw3EpBrzCnyItZUSI0I0ESSMjZbavuCmAuwKkwQVnMH2iDZxYkczBxzrag
PyZxFnqUgW41bfylaXepjYYGWKJDdD7Ji5wUPFSyD7/3yKfpEnrZ/XlPAaxpwStURoOXYTQILB87
+UJQvyS23vsMh3rXHswQArbY5ekdCdw6HJi7dXEQDRegtH8ts5BI0Gvo/WntppZwoHBzNWCGqvRq
2Q8FO8OB28M2j4PA9A+iKvpuTk325qg8NIXo7U9RUysdm1W7wljLDmPxk7mDhXC1h5nQw6UYzBmx
E8a1stYHzJ7kKlZ34HH/nzOwG06Nc5FvDsd7b9yiq+UyDK+gw3OfNKcQQC54pmNeFu/qChQ2SVy1
Be3ETe8rdmZTvGDv7JJHJ2HsYtDnQUbQtGfSsfnsSSaToMZoUzkv3u9WF5Hz802QrV1yfJoxWukB
Gr0+mkmAUhSIl+LxDMOuDyvyk2cgaWaE/IZScMpnIJEqtMC2pwccStmYRcl0has/XjWoGMoIvV0m
wy6w0gh73OjpzXrqrY6xr6Pqxl46TnpGJxQ1oHEeTpfQxEHZ471kqIG+knwXJrYdzTskxWaxlMIs
2rpJH5LFSjtl5C8zx1oHxpjoqu7kuWR/Il4YXlWZPm3pt/Z3r09fSzpYXgACdpinhNmJpA/a4ikJ
XH7QXUznKkTvW71DFkWC8uQxc9ppmZLNmnL7PL8HlXhUZWeF7gWa5EbEKV4FFPFp7hxo4jVFBrDp
GT+FevJ7Xe4GdGgIa67uoSALj/oo2C2RXp7H1KZw8ZfBeHuCXJltO6LsHCHOzWJE2NzYF43k/kKc
Rc1eiKzL0+wVGMEwX2qHbei82cs8uhhypxf2su3u1eDRiQ7nagRI/5+fNayjAFLZYMFYArHeiDcX
Qbi0D4TW3LRyUvmve0EPHAh3ZfwH2UK8bBHkopRQFYh5mwPI3cwd7R3uaBWS7hKYzgLCPAUZHSJy
MyUF2uZHktAccFA9bJ0ju96B4cgTmBAfqXV11G3NhwOaC6kfqvVuC8DlpmT/wYUXpnFNfXeouMd9
lnAncCcOERFc9d5Rf5c9OztUHubloS9ljps8c+0ZG2Rw7p0/I2Uc+bMBnVbJWhXg8U+w5clSqI28
DZph3cG/Sk30i34XttRoAAdmjqknThmOopfR7sKHlgnyuBgObXijFBz6lbdJMLYIBTlMIdeiOQP1
SrOPQ4N2MPgZ1rDPV+tpfaec96zFLN8SADDmTVF0X1exrBYpsAOG/TOzHPpxRSKo6FU+u15GQPG8
3HUMaEltwkYryeJ5IRHGC8KsspeNr1dUWST5PFWTWYqk3HiFKd4f6zi82WPrGyDzWMO3n/LA4zEN
sQBEmwZGBk4PLD7jC7RuoHAk+9Hcfl6YLlyoYxD26b9fFjKc9RuhkJ+CKAj6HueAAER03BMMo/ov
rJsFrShLI5Q+gdadymN6QHcBx1wfRCGHpROuKO+5ikDz7IrWEi2AYcUkj/3793ZblCDs0KiRe5nr
tZxM5Zk+bPAh4kknsZnzMyfIyA6MYj2a0Bt6DAbcZCKZNdp5HlXwq/bjd/MFyr3/FAfyo/d/eixj
kEw7Q0Xrh6/3lU+vjXhO6siyjuU7qUKa3Qf/gNH/D2aeLkTpxyEn3Sil+EsdAiWsuApMldcl0Y+A
qYzIgmrON2wK0o3UwHHuvO9QFDnOLL1VijGJL51BiOoNSQChc1yhCPYnORiNdinC7+nqNiI+CwDk
iKfUi1r78RDNzzEX0v73LRGANb7T0BpGog2MEmJ5HwkcfZvquGJplq4RNdP4EqzvQ7i6skkt6TRq
WruIrhd9Q5qMuAt7ANxb9NL1zozgB3JBPYKcILPy7boT8s1KozhAwWvszyOroVWHD7RnnFvVtmyB
LfRRa4YAR5+OxGFwwV/QlMLRHwOM/vZ5jkqDuikvvzykIvBXSwBX9koc+Sq0gQOvCVxWUPiUCpt7
MbA2c7M2NggBsmSRe3JEDwRIh3O38+ZY4L+soMNwa1IXt7WXw8/Q/FP/s4T1P/xDPRHb0jrHg7+q
RHd1GEIsNZiTk3CHJEEWVXtsLP/QtbXtid57//1MrYdTjnoL/bieP3bLsatOxvxkiKFyz2OeB01o
oybI8N0Yk1GH8fSJgq5MUGvg27+UxBBWE8YR3yD8sxNwP6RfBGZ8/JzVV7P9HQa+3/SD5lyf1Xb1
aFm9hCR2Dm4Go8DVX0EIlDGyQclOBP3m81bc4hV2bTyNd4dgBe/0hQ1kLJbvo1wmsXxki9R6quOw
NiOBMweUBNpsDbI0q7EcdpPsJtNlfps0/S/u91l5UDbBhzea03ChJyf3pivcUbVyejRBLq8LW9ah
gYANmAmC4lvxEZCzz2t7HTYzGyX2OFwTmg0JRAudMXNu8yjqh8AhC1wM5/nLhfpz05KvEjhU4TfC
DV84j0iqquSsrYEqIePewWftKWj/hXhw2p1VOrQhgDfhCkdkbCU4vqYPsQ6RfoaLOrpilVg8zz8l
ht2SkgEWKqtSUjJFrXVYGPGoCHGkktAw50HnLgEm8qHZD9vB15rbqnUzhj19+ha+7jvwyySGBnFO
IOVMT2dzbp+PVOxU2yf3LFdFej+JvY4gDurYzKLSfk3ljHpiFEmgHVZzJBklC2I8kIOvBnoTHNmY
IHGNdaVcik34tKMJs9XnzjQf/tzTC6dRc1wGwMMko1EzfjMyM+3ppinIZ2PNvjNACS6u4Sg9Xy67
zWfquvNYHsNDOHeRDjzOTTsek5gYNwoszZxzrFSYWWNj4SdBpE83qBzZbrOB2oYxtdMpbwuArsGl
H/OnKPgwMEqRvSzM1q380cLzP+oO8lUo08HQdE4bNe3cJbdG7LYpHDKwsXKMXgY1tn4vjPzl9/zn
ADcQ59Bs5cBJhA5Jeucy3+3t8Zly67mBSOLBbo/uae3dHtXp6oIdArCIrHPi6W1mq4Sxb4nILqb7
OhKVLHcAWpjV8Xnz/jPQ9yc9A4XoVaY3eaZD1ijEdQHRPyzIIZpONqqrl7J93mZqZYqxZIDDx5Ia
O82jvuDIcXVy1CWs0G43kQUpsbRTJA6B7ueHHz2p9Id7weAGScS+U4lxpmik+Xmv3NdH+h5yKFAC
qRAh8zFkMrhBTkGq6/GWYOxFNHbaHV/MytNTJbbbC74WSOmeb0JsRJPEGAmt2Cu9rSllp0blo09Z
PyKEqfVPezV5VVqGOxqndjx/7xUmUjTDM+xgYinnI4hO9U/A3OE+3wrQnBl40jJ7hYzXi0K/dOHK
NcIPoOnu72VNJrPjC369jn2WuWN2Vp7sb92W+o+kF5tk5Em2peAZgTDXPPfkK1506aZl/xWwWtVi
76tQEzotgbI6rfGMKbfQMXk94XJ4fic0OO9CmJjeROZhaSRzvaKWlS9vy5kfoTg2WboMqqFhn3Rg
2pf8U7Xm56kfZZWSky/t9OKzEcT6WMbgifBfe5vLrdnBbFEnPPXqjoCNduMiwBEVRxuZJpUbSsQP
y2WK4Q7RExKeUojV8yIZqC4d7bfQ8ttR4QfeoiYHXrBnurWTlzRunEhxpiie2Q4x9MpHUiuzoCy2
M4rn5da7grXlgvdB6AowPqhOl9AWR+AJIVXJ8OAQqYSpJGQtQnfbytgUR85onND0RYXB6FA6+O8V
rSry9SAG8L2uHfY9RRBpsMc7oqi/V9MC8NselzPDWpW85GgEvnOv+2HHtPI0ru87ShmLo4uritlI
+wvbnDpOAR9vXbUVJ6HEq/fwxzGkTvC83zkh2uTzmZ9Bo1Wjap83TOks7ZpmdUOC3BAN4Kk4wYKp
qWO6oP8Q40O+c7zSYxppJS9xZC4T6DVw6pH4WgGZxBRXpgyVyg0cswSHnkyufFKD4d5YtNAaBSNW
zTtmVgreDDQFWU5XmPoK5JOM07BLN0hPltWs3EPxN4mzFFtqEWLnG7NujikW3hrpeHPXSS5Qv1hz
aM6t40CCI4bS+QLcMr5EUygtFfKTb3pL6w1sHN92bbu031lD+WoKRG3/PLy3Dk/86h+U3IW0rnty
CiW9q091Wtn9UfyF64fleeZGvvuuQ5l3ssxQlfmfb9gNlIIGWFNmAKwfTBE4N/0izkDskZvhFl6h
3Vm25NWBeEnbitRPCHKR39mXg8J8kHuEZi63J1NXqU3J2YnNFXdhDkwr28SP2UTj5TrYVa6oy9DG
4mZYiarc1otCul/2LGf8HUOCxSjUCR+zeGPsfW4J0AwP8EsthZYnezTVJJK5wNmIBdPgJ+W85eAU
1oqDTO4SZ+RanIFevhw0AduvxUnsAU71ermTe825OUtChRM9c4K2OIi+8oERzdiiBd5b2D3WRRzx
CpNLGpwpBIE4J0DiOx+kG6el5ukT+oTHmDlkhO1kLA7ZqRmfY6ce2Y4xjkj9GW9pWAdpGQCra83a
NoiYypOJgbtCu2H88cZQc3WyduNze+q3MFE59xX4sRIBkJWvsXhHzkV8C8tfQtmVea9rMaie8CQd
gb6H5s4V6b1fn7GlbcMwoG7OdErZtzNoqlBeQ2RHT7sHisR8JUarkQez+YsCiqYkecSoklOr4HCq
nxU7kTH/Wiq/W+jT1n1eRqT7xFd3A0dphsukZQ7VTf8xwdemEUrVWqI8G8IEsmN5IJunl5FgDgtw
XYXGB8JmTcg7iOw3ZtfZrerbfmdfSuD4dJqyp0UaBk7z7ktrwLToVkX/OQMjPirqK4k0tk5XhU2n
AN40K0UwGqyI+BpJfeubPfzEh/ilT2e3khZN/LqQoZUPVLfAlUmDYkGe9Zzs7WOOmbw4o4pSq+rr
kavMZQ6Ph1dXUEXfzsKv3dDfn/zWHRjuev7lqtYiLcX8BeCFvupmu1DQFtBU112yGEdP6TZQSDfG
i3MDh1cggazF9rVu8OPP9jlbFYMhYUZAj2KVAMX4gPTJxruKFhXZzmdGAmBJ9F64g7AJL7JBCzSt
m3nkJejc6KI4Yrm/QHjgNX7dn+9sV+N5/UV9zpczZpb8UnyEhrZX29OFwpDY2z3ExrKfHQmFMsAy
XASeiAc80bg85NuJgtXTdhRMBvPty8SLK8Yi//9BPtUd/fXa6h8pHt6VDIYpFJl2wNN21ytubflc
LMAUEc561yWaIi8tQJOfdxts7MR+dmsEjf/2JY+8/zKwi2bCBeaOyZkD+CkIT985GWn4OvY9OzNh
7SXQ9XbOZ99J8maBqIFYOQE1ZJNGGLmiVEfR8LIR2NTMqnM6dwiRohqrFygxGBxTd+icq+PuqZUr
y4yjVA3xUAlbSSM7ve1a23CiLuJoYJBhzLSESVeETuUzegfC5Y1bL/UKsOy0mEwDruY9Zujzx2OG
Q2gnswpqfMh2C7SiM7NBqgWSMd1C4gzmBCq15BSq9FaFIm3id9ySU1JE1gaxdPcUazuu4qxn81rm
4u70iRHsh8YdGKy/5dfYCV2kB09VyxGEtfccvfnwDjX2mpEKhaaY8OwHoRv/hd8rXg0w5bkQ8bVu
KU3j1Oi3LLFm9CpuebKRNKi7dY4D2HgZsheLZ6d2A9H4665n58xHmuceltGsrBTW7G3EpPOWs8BO
wq7X81BTBgktRajF9aNr1/qNpGytfcv0JS3yVFp5TqlNkxIqh4r7Fkc7Vu22TyWt8EZt3MW+dygv
mDVD4arQ7KygT+RoQb2X8ieSLVXCldD3xLIGSv330ZwbPjQCZaAj5q0RAtIxhB8QTZJbri5oKJ/n
yfWfFvnMJf28jcp0dOTiKwaSkJtK6i3GSi1vTJxe8D0rPLuK7HHJZZ84CiyZHTIMXgDxNaiFVm41
SsF/aKJ9dF9anFyeBIKqkxPfsNlUjtYvF2sfzkoD3h/OG6OjMlcbANfRKzUh+P+oJlwTkH7MrMqe
gf50j8HbgJ5qg/f49QivReCwfPA0xh8ajkvVNQ+qSo5qFALLmHugAKfgOa57iqO72SBUXutvMNiJ
TJN6LzECT5nmp/AJ2vB8k5fWmD2nDOelql3IqpXyBHGI72eHC+9u5sYIrwWxRrQOFp2fUMenWN+o
XbWOXmmlBtmKlTw58xDZMnGP1rzIbNYwQ2g7nOAOH/UlMDUB2v4mtIckiITY/2s8AM1O1UFfWqFr
NGPKI+NWxpRHEW8dGSKR3mi2oSY8xKQ2+CVqj4+glBUzWLoF3JlR49MVyy3z89xtmPSg9mZ+FB9z
0qazvamCPAKimqu9TSjte96SAd3mQ2gtuNwuCciDAybVv9DppZeGjJFVwz/M3bAdSaWs1/1YhbqS
yZKS1wFiNZ4XT4PEOD7odJp/Uj0dzpU8FzCUORRntp+0tXCPr6Gp78N4+Z5NNGzpM6MRcmjd/7+3
ZvKgrmq7bGw6BMQXo6gGHHDjsMU66iSJU5h1QrK9MSDTUe++iZJGWS6QW4SzN3CABvm9ilqj52Yl
fpPQpFyAL/7EBHutaZrj9ryzGm8I1UW3OQPPVnkT5cmBv6vhNucQRW8sGmGW2bsn0Q7++epPM+R1
2NC3kbynBuloOTbO2A3Q7vHFF8qbX7v60lo1Bsfmxs0HVtTrhI5ThvlrwRvzM1RgBoeSjplXqsFu
DSJqLdOjk9HCBC0ccrq1GakdICVz+vUHRMghUHs6A6bwXKk2cte2Vc/itkJIRO1oXyA3BaP0/P3e
b16ZxUWSr93jIGgrbMeVU8aKy2cbp5xtz35OwiPm/VbEhvVSnUmM/OnR5RaNfc4bwj88NVrT65op
a0qqaN7dONCwBuap3hr8E504QXMzxsy5/P27+eEVzn05xlDJcO/3uYYXj4fZn1wV2/io3wM8JA6M
7rHHOOClowgJEMTNeypUiZ5SRt0xsHMONxMSFBiD3a3LmYRzSXPQoMham4A88Rh845jlAnulwb8z
2Jm6QHJvx06cd1ZnLHwO0zf915jTOp1POn7j27RhCdjffGZ4WxqCKljLNccfPKe2o1/o426aZGTe
G6DpLK6/Ytfma8rwwIrYiehzNJCsf2ai4nNmfLsl6pY4xH5fYleMzh81+NHiZhq+WuaVcH85UkPM
laWJbo7lP3n/QNsXCVbfoIEJoFIshKfQ/8ndujTZ3XaGRLX6NX8THddF5EnA+HBjbfHpso8Rshur
eFX2tgAU5mnR3H/OWYtjFn7U7PTwhsIbpvk/tbTjQajlCkps41bcbw0E0IIKsoHVRo1CreHyraHD
ufwfpD1+kHqF1zBsMc/GSkKMApKM31106Zq6MAiMBgPPOuAMpIWJG1cILOdto2ZF7RapQv35GJOg
nxrzTCxCUMZqdhSbmOxIwggtSYtDIkM8OgVK2trIaa3JxwE/JbXiPAfGtukYFfmaEbFpGjOHfJsn
5bfRQ0mGXUgDD0/QZ8hUo+8N/2ZWDC5DDyElxg1xdj5ybHPVHaI38A8FJ4p68pTp5FUNbufMi/iE
IMedD8suWYoRLldtd2kgvlFHEvOoeVdojZ2tuTXeH4/jBp/zXaepFmXlxDN7Gwkdm03xbDZPhkuw
A+orwYqJfKY8MtmvxnoQ9pbgXEJz7LIw2b1PFvgZIMOOm46HwUI1FrYYGiRIarPpmtUQsPV10GtL
TYzZSOU3iTKgaipBvpQKBH7ECqjs8md4zl28uiYYeYtsgoOEMIIjVTcpv7XJrM1fegcg1js3dQr7
iNe/Ag62N/JrHew3N87PzZFsR7DtG5CDariH3KeXufJeiiW7NTX0RWXFCVhq1j+DdkeFRQZ06T4a
dYC0oUdpt2AYBB75GByaR8pJsbfbIMlCDBPRqXksO0YNbVipN/0dzBaJcDmGKTJuO2uMTKvVIegv
v3VTRmdmPnqylbWA3sKGqv3VD5prIgaAEr60HZfONJv5Utr+1hzc4ZYcEqgfLuqJRtIOLShpHFT3
O8GhM/Trcgb8g+DAHc4pG3S+DPteBZZWm3ICirbE1LYPQ7pM3TwVlkXqBHXsNtQnnl8pDspygSZE
MjOjGypggiGFvCZggfJiPz8u2lel7wcnNMXUB/wP5QGbfZbacXts/YpUCqwqXvjK7Wbf9nFqSMm8
nQ0Zvq7PxClZyn0sN7f3eE0oAgHiA0J1ot2scVvVhz85nt2+svwXZEq8hBrbeC6whHsEfYlh+sGo
eEb3au36FxwhBSpyDjv8ThWhjMS43HBBHxmi0uoPDkrulBuHUoNyQ7j4SCtvNJ+z7rNMfEEaWpZU
GQrQd153ZlSid2Q79jZefBnt9CaXws+IP9ooBEaLwgQN0SGDnGIHf0nmCkiPKvmMrVyiWjvfNVtg
VJ4qs1hsf+D6mFFsbCIl1D7/+S7ij2GonQdLI+Jmu+bEGzZd9kjvyrbciZAoRIQKqLEkWxWUMw+a
zZJ/XSh3RiOnhf12cs/EJ6GAxo/o0qraBosbUt42i3GTFZ7Qv41QrDNcJIsZW5ES5ZcKGr/Z2odF
LoO6cH0T3uGaIB7LBHvFi9ucwrgisqD8Q1tUnGdFt0nViNVY++vOVuErc6q3ez7kTWZdVU2ZNHAA
mbf2RJoKc9gxxC+iS9PMJ/oAz1h3g7IUI3nIqSRWRg4GV5Fe7+Y3RjwwwMhoXua4skGi2YnnxQZs
EYLRZTyxzE4FFMniQkcYBHusfMr7gClWS2+65wBPGh4fWWbx5no3aaFDJcHNJKj3tgO07w9vavcs
7wS3REaOMXCn98Gcrzn4+eSrdzW+D9eBWse3UCjBXI3Hrz3EAZyheeJ8SYcgqr5lWkxB1W+5nG4Q
jKRhY79CIllg1FZEdtSKsanIFGeOwpYoTkDhouEtP6TZKl2uaqqPk7LVWZ3tmxLVluqVHnis8vFC
keH1yvukf3e9Dob0aSADrirUStsqrDkYQsu+0VCX1jV5GcU0k98U6GsWl4QCedV43ktmzB32psvQ
Gu9+x0RtS4s2rsyH5ev91RDv8yVKHFCHWNnXDR5cuFPlAfL3c9xG80iw4XVSVK8pTlEBczzbc2AK
2zkfsnOKVFCdDImdRjfX7FhRyklJ3RCaTJ8hHXOJV2R1QS6Nk04x8xA2UyPcpzj8dXYsT9PCAOCo
SMYfj32jbSKg7LM83vYXLOFjj/UmyWfeoX6skItNG+yJTWiaw9yQC76eOvfCmBjAKyrOhs6x6ZvH
DhrFqxcTkAizc+wKsQ7CdeLRJIUa1ll2R/mDdETse2IaXthalNJMPuhK+mUWxgOOUc3FyfZF5rjh
p5aqpdO+O36FmIkjPccbm9f5jHG8tLjhQSBQskiz6Filuqzw+wPq85yAkxic+Od2HoZsoKyRO3Tk
PfdgCCDDT/QWc66+Bz7V0XOdGneHoBrwJI1tSoa70IG7h/E1CEPGdRXuMv7F7wwiOqe8eHAjIFm+
4ZnnzVoNCYnpB4VfWRmRzneWGTlhIgYbXOrWUp73S9tsmFnejlKUGjvI9MQb1MPMZbbCmiBdWEwk
n3/TkQvBnu8Q6VlJnIMH+Ibn8geNCgMoUPRQLKSZzNdSORlXzH6iMnMLNG2gVkOSVFLhzIemXwRd
drAonCFG1P4XN/nbpP1caynnsgXhb/J5LE0AHKGuuWWvcKViVKbzQScJy7DtY1pqjccmMEvJdmP9
7t2dMZoPlSKV2SVLgciVvQP/JG8DnMLDfGIhZDzwrnJK2E/tcKSQ2jOqNNUqMTgafxnBpW9F0vKn
MU9RlSPK3wPvTv3rSXbgePna69rsbSfbvwHEodR4P7REcaiz2pwIaKEvaivkDL3xZ0bYnLFFPCF9
YGdXb+RBchjB2i6KfqA/TRJqkLUcIb6zrqA4jGzvW7nHB85ksz07NKXb86wbv/Rmsy7XpyxB94Zu
6i1hPI2f99plKx/QZc3siD7EaSHMULqZar7s7fiEzDjL4FZd9D/NLjTGdnIqYewzzWtCtibEJU5Y
SOGNAQD0L8l7xbOHk7/avbbGR+sOmwJPbotVCkFuM3advznUuTzJCezin1T/Y8KrOsJB7ncQpT3Q
mAmtXGha69VlS2qhDXg16nir7Q1FRqUDipjzj+94D6ZC7sFMdSNIBW6Ytway6IAg1MoqyUs3nuRJ
97owacq1W/NOMlnuSe8TPbIYqFYrkplEgJZN9x5d6v2rLo+msxPn0Wr+zbqgy+AcvFyvJnAvDH4n
el1Rb1UwITbCficYtSJg91wZC7yufKJ5FbqEPCsrZe+VCpbTtZx/RRv0CSDkCfpaJTLhynTtX4Gw
WU9xg1rP8BeN7S+Z0ulbVvVJCjKkRjVz/OW2LMQGum9qeZ20WR4xWagAbqbLpUJAvBIH0sM9Begb
lnPTIDv/2tEn5jvhbfn4Tvt5NkyvywdASZk3ubAr8h0evCy1DTHhJkbTJN0LL0oeewAvtLNtIJjx
1vhraqroyRMzZNPawPuyaS4eWPbFE7bizkuzkJAjdLKnaPdPaYYumodNSMYklt09OQmlZXGSoflK
iey5v+J0iAEOXTTB1Sw7fK9BSFEe6eMHO9gaJAiOaZifWG0yNyaq/4rxpGusG5826zIicEqB543m
yHVM9zjh3v8M0bCNPYaSkXwgT9RlFVt0ORThvYmqqcGYGU2CW4DAHTZXGACd1DLQcxmMaRhQADXE
uFfVrnruRKnTp6IqecoWXgi9DbG0Ohti2vDHTRxuTFQF9h0RsOBB24F9q2Yr0QortchvpQi5HtSQ
Q1BwTCUYfTWzA7GxtUKaP+kruh4aVuYppOEjNGGfObJSPnXDCI/F0x6SIIEV9pwq7ZBf+ufpePUJ
W42I/zxHTfs77HkchGKl66Ct+sfDDGGD8ZG52N8/pjL8f1bVPjwmNvMAc0bZQmMUN5YbsXJ7volF
tVLIUaghu1wa68SuGyKdEt0cYuVi5bs17Ai2eadnDc4jRAMGWMOgYJ4A9Bxj8g5I4I2mV7gFH+1F
kTARUNGjou0RoO+DSUgiB7qRTb/E+YmTUNhPkLw6YBHbz7I02FvOWll5CHGzdqOCQk4f3ExNpxni
ldIfLmDVwTEQeb+MpIbGgHLkbgiOlMSw7TcItqzsDEsjDzdWxD1JwjYYR/IMsO1PkeckTedCYhKk
XOJcoYFSzIDUYOesJW0PRXAYC6tw7HXZbk0myVkbCsxQuJIojxnn+g11rSzmi/BH/YAzde74x+QT
NyCENo2oB0ArSAfbtYTLMf6NTlH00kDINBQXyVG09y8tPKir0eURVR3jpbsBpLMLJkuZQ13K8gNn
whyJgbGhU4QEm/0/OQHULbof0en4jq5Vf0FghJZFet4rEnEBoPXT+QGOTVNMHkAJ5ew8qjZzpelQ
xXh/wAZ9Dkxcro40bUh7ZJ5l8Md5hE3GdkLHzpJtkpTvXy2ZVIHKK4bwuDKUWt/bMUl+HbgrjVQ8
MySa51nI0mHV7vo5/Mv3tgXn7ryetw9Sph3z6gf4f2lwAaOPlfpFneAsCEbjZlw1WWByunfMpNJh
NrO5hU70aRU+hE+dkJ0MPKtCLxqBsc/CuCocpBkeB01CF+XCLtQIcafW3QSWRyeuA12NzmZTlYgW
TQH/E9E000r/z2oOsuecfJOR6ZZDq8x7TKa8WKUheuTrSAIFx9nN+/U9jr8CedDsWy5NwGIRxqU5
VCHQ6xV9jp2PQmuxDXvI0J/opC4DUNG92F9QmJnPT8yfhVRQgBiOT84olXAdRXd+ko3m9WWmFpEE
C1dMO9DJrjpaozMppL3YHDr+kycd7d5enqcKLWK0EkiGhBkpfKXh6TI7ECkJx31lxbaYTetbtdm3
MECd1Qwiw7iGKC9P4q8eZpLMo0kfzNl/+bRPDW9McJZNkVWnWGkD3DymH+f45DpacK2P1SObgz/q
vaMwEn2ZwRPs/EbaWLAaYjY4UooW1jqPT0lcaOJdc3nyeWoTT/0p+fabG6n94QynwXUn/MeUtKfk
9MnjJZnKyAgmX+WRj2MMHkbnRF9M57p69X3pVKfWCLper3eGwfed2gPAzv+7hqsbWVZtnmrUNOFr
JgmSDekx9LetUcdaJvcQhVkUS412TMivja8HFHAvLPe5LO882vkNsy/dwV3zJn7VbY22Gu0SFxQX
5ANyto/ysVCE6q9GJrmDvoMptrOAwaV87UJdo0YaC6SeoXVRDepqj2Lam3BvMOUyyXIClW5/hWwx
Ltkwgnt/wyWUEVhb3MBrDq/Oj6A1m7elsWz1HNi9topsOenNPSYc6aNsGlV29DE8i3Nb3lxPgRlq
TpV0FA4i6JiiIdgKpP9tIMRBAG/DeVuHlShopYEJMMiBCDEw9rS7byhOoR7e95vU1dCwXAKJ6gcr
MKyF6GNC20gMvIkBKWkAqnxuGpEG8O2lMaS5Op0L2EEryxnXoQMwlWs/ZcpM/wz7Xv1pYUJ36cAn
IPxuyHgZoKcyaYaqPR/PBPBvk+/YK+u7pAp4ZneO1r+ONRCqOjTXE20DvkB/JwLSDOCYOALMilkH
Pmd1mIXHv4YQp6kQmiJ6ngWk2HZKTRLc1AyMiUUJwYksVwIJEjIg/KMX1Q4fpX2jy7MzbkR+L8Hk
sSASfXOlL/bYlz+VudtjvwMNuSjig10JzsO5o3jbTmw7Bqsy4U84/zK2pdmYGiSWzNYY+BRftWOe
mCDl3J3xp9lW5CkEhRJJrQUepygPJ9GGc8pVsEUOu1tKnfgjUIGYGqsmufRfZIr86dfKNHUhESsG
vfWSL1GTMEJClUXdq0zlRHeMt6cRtQGR/biY9my4YJPh2v60vID2jf6qj9U2cJHsWCkJDhLrZxyL
kIm7tM7Ubu9+2QWHUKAttYWocDtBJXZ5q5kaecXGxia1Uo2FJd0absOt4IEjBYo6kCWbXPURI38g
UA49+l878t8KTn9WbpO1/Pmm9NHiwjKnvpsrG4qEuIEPGuHxewWCUaJ9J+URU9xT3X/UnXoSxLcD
2bqRMnSCnvug0bbDONhVuXqAeEAziAalCKkHWNR7CI9Z2hm5dNEEpanMVnPugRvzHvXATmfbhkS3
E9VBLGDdCPWg4DxWfvc+/5BmjmRw0KXBt78PgVmwljR32XldQjN5JBWx/FLgwB01VYtaT5laWlKh
gMwhpxrtamJhvGETx6MogHhhhAUASf8+eKO42RAIBPRDYJjyVNIftcT+fUf67iFVvyA+cSOhjDeb
S06N0DJFzC7gdHI+dru8VlV8SgLrYlg7+XL26EMLLkf7ZgnHdaC0OWMe3kqldxFpmfSIxNsZVYF9
HQqaupbb1zEFa5DYUGyYlpNvMku6VQS1O275z0yQZuni3AzIAy853GLmHp/ot5+P15dMlODP9wgQ
uSKy65QS7SBWMDhOQIqZSxcpK1X6tCqi7J3DHB/aUJfoXZYqUvC+wArctGlRZ/SMkoZVMxykNuNq
1+QmsKK3vN7phe0pJH89aj3IFAK1FdH0MbpRm3wEPS3lEHM94/GxrSzjUFC5fkcmwsNHvWbmNwjw
+JLFayAPLbFSJNdmdsFfoyO2zwzvVbSLk+OMctAZVyKsV4kMc/Z+SfIWhquT5n3u4X4muJMGPyPg
ktLFIoaoOk4Yf2cAB5fB9bQ0ZtMWx2wZ4sk40eJGgvzGKiJGdB2ax6SZv8VdA/3FkbE6QxLZiyNl
jIPuOMssiNGe9l7tgjwNT3m+Rq/adYxZ2tJEeCzG5i5pk7nkDX1G9VlomNtJSPhzEf0HuRQ3lQe/
l31htVuq6GpyrTiX3UrAi27ETT4nGRHJekLcy00msbKzlxbSDD+RF9O5LlkXkE3avJya/feioWeW
wo7gX6RbU48EWDJMWZFX9iUhqrlVNQHsiSKDZXE3HW0pB9wzNqg2qeXdl1Vkvcf53/pZR/sfhy1s
tRDSAqESaax77YyO9AdJpWGrUyq7J29kAdwSerPBUeKFL4SNaLKeaUcTnPNhf6C7nLyBDgSAcaRP
PTpbqCifcdIBVrJPU/0NK9F42M5AoE4Af2vFMwogrbEGt3jyL+CfNhssAHJMB3PBDwp4rAxVAOo9
8fBrNu9vOF544ZkgpPqSame932EkYqMjyNYOvXet+g27l6Tbg2M0aSk+5btbtAD21HdrhTFML48f
vNn6JgOILPPro1DRqvOV2uPxS/hc1kG6swI8G+KZfAirkbA0F0rkO/40UKSAp1bF+JOmzXApuMCI
saec+6QL6C4USCNEf69AVT5vM/fy1o+/nQX8Ma1lwujg9zdJBQoWs/Ba5tC4YsoIcbUtuZ/JEIUq
fxisbgcr7GaUv3I/h2PB9fJo7JuA/loxIZ7KLcsi9aNWiqKB16Ps38Q6S5o+2qKuYjA9YqRu5IkB
tAE/2xUcOh1W7OONEXfKkuFg2z3Lx4pnuxRX1GAEzuXXMT5dfY+qtrpzsrDmZgVKPDlnlTyd8aux
WLSftQLpbJ9MdYVzKh9t2YbS3pFuesk0M+nXFEdA3t4WtoVnN/vcE2B+geqJlciccUZsu2Otrtuc
vWhKbgF6dS87I/D7PDPK6NaJ5MOGJWKv3awsl+6bFt+jQWu2xbdgOffjHRI8enVxJTa2L0Wu5Ftt
Wam3HTTd2UwZaIolqTwPOBiBIz3vGwpqkmSSuFMGQQsw2Sc5Js45QvD/941jkc64uIpArwhd0BGj
GUVIw4g7ikMgpwjgBMj6kADKgH2wmYN+VCafVEe0B5tzbMhgJ0XQHa9Y07DrOzePW2ecM+CjizDU
DjF0vmXAfE+9LILlnCO3uDXCET/1zqlLh/D30AgeAKkBpN6rUHbC2AHh3XuJIlOqH3PXczJTGSD8
JeVZzv0MPaZtKi64RqDK+pgiikES2UvM/AsrG49NC5iZvD5ZK5FXV/XqXJyicIuLaHELJNWVMoKI
V/+83kue+xbOMXChy/Q94VNmpq7CxPtv/mFABCmbmFGHsj42AB2m5VnJukQq2F21fxi5abtRtcuo
fzoGY/iutFvfNVLgZ5T9B21/FNcu3QNbfvQzvJAlvQye9qLL14APGLwXOEPj1bA7rP3sA8dWgrL0
+v2o7//xvZj0zmBQF41aUa1Cld9RnAXCU3/k03mkHrxGq10AYyqe04LGJzkyahC/M4YLna1ZSWV8
0RxonFTTDCE4j+aP+hq10nDsodFYth0agf6Tw9C5ezcDJpYYAw9KsQG6cRzKQaWr4Uxyipqd+cZM
XeFkAlctJvl9SLsuJt5Mekqzct5QwRBxs/AcFty/ZGWud+rDkgxeaRNomV55GxEoZxiuUhJEtfEt
MuzAbqTiSylULJzR9MPpjwoY5he1GftF1UjMBioTIFTX+NlpRuxeeJzFD8cekmI7gGhDcgAvYjwY
R5o8HuzOP6V4eHQRtvaqznuY4u+dpvqDH/GLDaPYGFL3HdQCX04Qqb/WMHBhk2lH8jMzGNdaMpLK
AYrZc4GhPFNCC+Hm7ac2xt58z7sAGFC4iuRNpWkLFJV2JGUW+7DzmBkFnq5JXJtALYlXI1y9mbuM
z9IcdEk1NaQYKDu+ldQg9rrBYvVky+YBD35p/iF4huwblIE+SezotwTeOkIUlGS2bVrL8La3FLs1
xFVxl5jsvD/fpHQrwaOoYUV4kRpYviwsXYnX+33gWhZq3u9BMHJVPGzFad6bcoYJl12joqhc4/ob
4z6+XmuIur6WQff6z5DOtG1oayj/H1JHngvM6Uf7hspSaTKxA8A5G60bqYIXsNzPllFoDVRld3d+
6A4TCP4rTtHXUgVtKO/STG6AmGDQS+0LT1GIf/ZyyEc//WIpUxcklqj6QPtPNynimMsmyCGlMwUB
Y16FI6mXodcC0y3LSAXmCmKQOd0eJNbELFJd4IThhOLMpjEPrPaiRjaYyOtzoMEeU6XJ0zyNnBTS
61nGmDrrKZ8q5vlHImsbpQEnXRaFgsysXrfkNesoyH5gvXAF7X9qrEqamfgwyIe58SNl3h882BCf
6X7SgQ1OtnIK5HeLOvokYUmJl+t9y+2XSadaItLUaXkYD1QS5bryGTWwKYng92u52s2wsmcmI9Np
qdRrzly9t/imGKBZiTRK7jF6SxH3ou/DEn3IPcpzpCBq4m2nNnxAT6Loe2VZ561eHS/J4O2hUDnm
P3OmjTKkkZJhbf6RtPjSoNAdFKNeaTewZ8XIYiZ1MDefmmbfs/8xxN3dxMCouSi86i8KPfTJN+tP
Oi5upCoViXRevKDAqgx++CogfGLH5B71wf4c6pkX5IBPbdNd4b3089aqrxVgngGSVuOoesMyvzeE
yOpn1g34SiY1r46yvVg8l+JYklhOS0X7v7YveXnTv5LMR8+Fja7Rzg7+aU8ffmsvuzyJK0lNDsgt
pe7go9yX7MKdwvJWVx4g2kGl4peBOdkCPs4UO4/mzCGOfo9J6QEx5bnyb95d4mDOsObr40CxH6dm
AMLBpksrHRIriuogQu4LjjE/owfqwEq/MrfC1UtK1SJKxSdzAiSy67aCmKql22Mjhuqx/hJYQak2
+2C5BetmOJ0xeccUxQBP4S4xbSIZmGF1MC9Lpbul/4tYB2tLKYIALlQ5WjiJsQRlKBBrigVHcMtl
98oSSe1SSxXg/qDYfz/tjnxB8SHYEjXAMOWgd2ITErg+AAT45oFu+lggINk+vILtRoSloafYWhKI
GlVeGPliAgpFjxqgdIzuSvDvT0CEHVzw2iHXxfqAjM56HikClHQ63COgJ5b4DkCu+WQoL38MDkuV
ruPF1HblF++XX1s/ZcGXtWgoW9wcJoI1ic3yGxbakSrweW+PUreFydLRGez0L9uPvJn0cLGdPB6I
TsJx9iCYImwtUPbcvHpQ0O0Pu+Y1kfFdx/jU/89WJ2KWBzcjDlWI72WxcExv7rhe/3SNdWkVx/lI
7DRA+Crn9VU23nMVsexbSiJlv7EM8/3i98ctK/LV74/TwWGh9o4qosqHR3k3xnCByNa5z3eTsnwP
zJ2FQJi5McdUeB8Y9OkGq04yVzxa/PJAQEbZm+aufW+sWRvYJbI1AT/j51s3aN5PeKteFW0/MYq5
VlE7ZvPN4UL6j8k1A80PjyOz46XpIt5OAI0Y18CwKVz9U02N593rUM6z7lquMzD48VKv2zMEC3Kh
kQfF2ipjYnFGeh35der47KUS/dwQkBei2qfwAbk1unAAZIDrBAnhDKJduOMw6NYrp3tO0a7lYZXn
PzT+E9ObBiDOINrhO80heWeo7UG55FaDRNp0Ffi0xWcHPMN+mfBJjGkyryFGH2F5EroKyl9DGc+Z
NrituLjQw4NeC7OXsOMZX+EEPye3Pz6L7OWE3BAoB6+mZzg6v3oy4Kja70lqIJAQGsJp3FhaMqL/
FmJyMfW7dOjLgZFqSpZ2xOBG9SOeNf0Fhbg7T0FBzo0t2TliIK6XxCzIRuo80utbi0F/FRkwlhFF
GJ2xaVOtt7ZdRChwqz3k5mmfwd0jPJdcQctin3llr5zbYnIBBRFn890YaE5YXwDlbwC/8r/twv/u
Ld33qloSVorvnovQyZOY3elR2s1f7jGWlabQuaT2V4mFodp+OylTR0+u0Um+UGtSm1KF4xt1GEf8
33xPk2kyIsUOJpbbDfM0VINrFilaukQPPxTK2GTYwN5HWTWzXRzy64pUwTPI4dm6a3j9enbspjvn
Q1bZ6IAMLxXJNxZfsNolO8PeHLjZSq1USk05kgihCrBpT8H1RI0TcKy18oWY2QjGWULVHSGvBnk7
+zJ7cb7MNGiTs3VUlmFi3cI0jf0qaEDSVEYceeKX4nI7PB6jZ4cJgKHp1GOpPvQGd0iiGzkdFj3s
8Rr5BMjRUmTT9cLw6xH4Ujar7PV1aCjcbSjf8RAv1YbK+v9g7etAHVYiiXXAmLk528seKylyZQsO
XkjhB36lRuKBf/Xm73E5fov8GyIlq6cDr+ff2UdWP23bOmtRyF5AxZ31jV5jKQTWZdisduR+HGrE
9n+WoLu45/arSapAQRwJ8+tZfpmI0Exyf02nihfk9JLLzLB8FbE68N/U92g3abUtk4xu6h5ElLNi
DT7Sdj2rDyQDJSQ+2/mXQvoYD7OjoqmMBM00tc7wSgA/j9CpACrnKVj+sRcpEW0+y36Lj5Rn4LJw
P16esE4l1pfXZNfqBm5bhJx3Ll9SJIVrP8m6JN3IMAsgM6LfPhB4Eoy9C4l+I2CURr16lDKCkI1R
byLB4yJZ8oKthoMSCzoANe8LKusGnRmdQVBMaAxpPhUee+tQXn91Tpm59DFlpflyiCA6VVlbbnba
UoP0XU4Ghk74r1bXYqJzGfHp8IqVjKzmDaI5rDM0u2nVKudD9LEsfSt9Xd7Z9y1TdoFQNcJL+MSE
CbYtlgkHEseOp5biC3y8jYuScK84ed7b4fH4rLDmCSlolaIBNT5lNS4gULZgpM2YvBh0LlfacxfB
uPcUqoKC7dBVlMNzZ3c1X32R87p8uUsnaX9zTORUVc2qCMbxz8JGd77BJK3WMwdXHMCCV0EqYps8
GCVG86/SWrW9zws6q1RrVgABW6Z86UoiEW8ZNKIwbyIfiC1hggBnCBhLr0ybgaTb/TvR0Oq7W1EO
EYOEPcl2Q4OiVDaXm08dkCNWJ2e4KASDXcTMbFmh4HP7OA+HFQ/VJOl6XqWUKbGf/6ofWbGWvSk1
wXPZ/W4vUL7e7LVI1pfaEPD91QxOp5qsX/n4p1XJ6EN9AmA3LUzdqHpsZjcBOvOaY2H2a7kl1aNh
Rzykn86rHG+/Au2COH+HSicYeHeQwhfuAi99hmPsM+2UuDGmekG6IaIQNLbok1IfVEDHcOvSVOnR
mHHfVI1j7cuBdRA+VkWHZbadCbsMJ2KECg1EmlS5G00gwVOZoGwVhIPtDnUG7591MznSCX+GFsJ8
Tx0Lh34Ass0qby6uObeMdL5VKheQ0TrE7efpVN+X49tRB/GM+x65RbtUu+EK3cDwF3LNVTBisVYT
2tOYDToOqS/WRr//4/UnVPXOrQ63hxiT1nhrTzuczGaMtdfZSrScCxzSy2wZUOzcyaMhl/nNbdkZ
sfVUbkcGtGZzglKs/XFFwXj3C+WVMUdxCkLTePpFgl91dxemI3zoDFchSydi5uQy2o8VgfvhUcLP
r3oua4d05wWrQIRSjs+u4R1imvWFvpjDEXuAbhmYqdsFXzXnCoWu/DIgWyr+Z0zQpAcShMZXd39g
vtV0TEf1Kws+vW/ye7Lkqy/Z7eiPocub4GX135UEyosy1MTZl5NrUfqMH8lGMZQtLu5aurT+IZoo
qrq9sQ/UMAbFJxziVssMJt7q9PtRFcvia2dxqJfxlhuX4kYPVAPZcJGbKT7Qke6t+AU2tgwnbjVJ
etTf++5YwIJPoD1/NKf7VUzK6f5jGjqSPG23IcbAeBy8vqja62FyaxCwZn9jbYzdf/nUIlxjrGu3
w3uQbdNKhBQjhuVo/TYyabhTKIx1Gl41geAFAnuxmMDIfb18kzPmAbN4Xhpdc3CsVhkhwkTIvR2L
nGBW97/FKzq49l0iHlxGpuzWXHe2agsQ0JH2iI6P2edO8mAN6AMhsJb0Cc1lSDO8hIEJDXHUlvWm
C1DrNUxi3WROE9PTmFsGNLnHry5Wrq76xK9rPDZN6Wpevnc4siJgv1M8KGgfcyfwRSejvcdnh1eC
FLBjMrw/ZS/JGcjblIMmM+ZuK5PWMs3PxCtMbyXJl19+dWYo7RaWPJUCHY0StczX3WT3j9UZ33xU
izGos8G4BN+Y4pBmiDm6FvZZXKN4DjTQkbGYFk/NsJd8TKxs3zbyU8mHyLEAzwU2ERs7G+2AFnFj
dm8RcX5nfHGJgONDU6etj5LaF0b3Pc8QK7bcrVhdExgQpsU8f0uji/64YONP1QF8rs+Neib1Fmiy
/vB1pI6IOpMrAol8GchgsLugOYk+EGynhv/58oFOK+eNa0X828VAlWxzgouAHIsS6K/43On1EZh1
1sj/qSG9QifYfmKEHf6oqXTmeLyF19JLu4kOHYDUWJh1ieCk/g2ynQMEWwnb4typSV+3iIayY2Kb
talLPQPmx+V9b3Du0K0TOlxkPOk3aAJepli0iFNHYCZQOpGk1LdSFzQkHjEeIbz15CuHMSvOJSuy
w7yG/4QZppoykGw1JqetRU2Fwc8VY2c4Gakp/9ujDkvYMut0NjgsyAqHKgdrR1UxY8hRkWxUZ6O8
SIPNr+EP9cA9nwYUEWf1ZWIT7z3x+z9tFLzwoUUh46qEfM9af45Iq/GYHqg2tsCSbh12skVSn29y
cRqJmY9YkiIkF9cNp9YXK2KNZfFfRzQ1RhVICH5TEFlSYl3sXNdBy45BbMQOZrn2denVJs4o7RGV
2DenDMALsPCwa9dVpHwrrQfOEBYK7isrlUweJyocEEPKBjRLCYSPx++gjXrdcW90BYqbvV7x1hXX
MA+voggVPqxZnQEOOOtG1NCNbrfv27uY8xlP92Io8lW536XqLZIT/GNmU9KhP4//Kz6ccBGJS1Fv
xKc2QfFq4vZBXiQsPCJdCNV9nrt2rx5shgETIYq9kHKW0aENfKSAeOu9rT2Yp1nSb5PiDoJSTeyu
d4ePLnGTR7jr7u+41Qj7QT7x5MtUzygOKJlR6tdfwgExBJhcfmUeq4lhD07TftpbCcm0ljIKDM8T
eByWJ+YJNH2gwOQAGIVv4onnAp8IdtS9Oz9A3FgFz4551K8surzLTSpmpbV7qdw5lSqQYRE5XpTR
GVnRYjPawcu359vUBPnXG1AXBReMemzxPKmdcK+87vpQY9i1XdERaCvMTfR6Q13NLUrDAFi5Doxg
hUWKKp6slbVDCsP7IuFtq5bMxGoDnLFlkiznGiv8ACqDPpf5tTiN279k4rp/ZOi2uKDfj5Hi8hkp
DOK8BQuXMAOU4po3RZjR59po2OvO33usZPlHiZSUsbjCpTTArfKCs8c+F4aicxlwvZXAKsoOdJ4i
VHXfAjrhAzeFeCWj5J3BTioQMIC+l7Ero1v9f5xDRLJJGHshO8H30klI5lao0WDhwrYuoGwK1WMX
93wE52UXtvfB6zmx+MrarBEF6Z4ZuKxw/IeD5Yq15MaxhkH1RQojTm/QNwUGRxSdI9sNYphDKgzg
VWXRgpllBnOfd5ZKx+5/bpYem5pzaHsykeVunii7mwNhy70/bLIi1ZoDFGabmkXIqMn8DLZyWxup
m8ah3W5k5sEqoDsFbjFbQOCcit14gT64SWeP8AwdhwlPEMRqC1ex6b/h4uBc0lVUwBRg3PLOv4qp
jZRphE+KuLxe1+qS3sPcUKJw5e7kDScsxrO7sc5l2SjGGvPMR8m9VU1TmAQ7vWgBC6B/vL+jhgbb
GMVab+nSaAHzLaXx8KVlXGEvPGLfhVa1CFwFdKEMT4TmfCx9iGO7QKys7xp1tZSnMHQm/LP5ObKF
t/db+fQpeHxv45d6soin6PCNuqSofuCkp0tVrT3mlRTMDJ6sudTLAnkumThODLkjWvv8n68TFhew
rlv/Sb4Sk2LVQby21ZEhJx2bPF8dXqJxkOa82DW6BNmlvKmaVdoLSCDqoH7kGcZllNISlWs5nn9F
xoXOnFB9ss6zkM4R+WuYvEaM9AeVO4LxJ9McOUwPTFlkEH1fK4J/d4CG41ch9G81PsLyNxXS0l+i
xiEgmKg4sFo9Iz/OoKoPA5dBBGMZJV3QCigiIKxnKKcFxrnw1nPenfU1f1QfhXMhY4+wrPqxJBBJ
pZOYZoE/lio/LE5NYv+DKSHV/vdNDbRHJ5UoV28WzFazNnd16/JBs1QANEHxxi9tRTS3xOO5kcTY
Ub/au7cMVIUL3Qa7gY5JeNVyrZxSXtFIq06snBbpYrmLm92pwis+vtKls1eW6DlcpsaPZVbld6Dz
BcWO5AnABmXVYOF8V5SMnCjK/nKlVkCqU2RREZD4tbOh9JAfDLpomh8Doa29q4BkjqEX30jWIaZr
5rzx7UM1b1BXzapSlLazF78fkezZeIY5XliQNh/hHrDV2j+s6K3H1Gfzwm/QPOPgU+JCND05Gqjh
vZ2ZP78rgv/4cdCy+rVjxN4nypNNwQsNP3wa9dIXPjl0K90Iml8EH5e5XawfOO7IpR0Mxp8zRfrW
Lk7RpE0KzREyRYDsDUH693wT83VTBEmSJez4sgct1TUVdMU+mCIyhNc1kN1Y6yjPJk4ClyRFrYup
2hsAfHdYc/zRiOaXMkFPT5jbqQVjxXd09edat84X0mrFFQxcWAo3VigenutRWTVANprHUvpkdk9C
7Gm6Q3O6eFpg7JbT/UgeDZrEeGlLEW57Z6RXjwZHY/kC6J0FgveKmDG1UOiHay4pzDMiLzLQnxe6
loR3le5JZL6fz7Omia0fVyewZJstaPctszyf1a4l/H9RWE7Li1L6lNJ4QV2p+qLCAxuyfSFCq/CB
R0TvknYBgXgOsoPeW/PQtlXZbwfDvoKqM2PEr4NtalG34/jfkWaLmGANPpGQpBiAC43uVX6IAtZc
tgJkfNMN2rx/cR7iTIrVdFxNMCNoy5CYiNSX1SZRIKKCrj8S6qUh+XxJkcyvxXv9cTHhGN28vPD5
k8wYtCt0FtXNkIKdxNdr6jlHAOKgdbpb4K0JtjykEdjZf/6pYmPBOMf16agyZ812MVkZmJzAjsHe
/RXMKlwt3MVNRL5IClykrwBAyk1QsmCxyNEOpZDSL3aeIgPlyWCdi1CdUxzzbceyqCytNDlIsBOi
PtATVrVF0Dz5QbTBZixzm6gZlOD+WpOsOkH/KfMgqdukkYoXyyRojdTr6xnRlLFpqcow5uniUIZD
yXJXWZJ/QJI3ITEjPLSsJnHz/b8h6vGA2Dz66qphNbPMSRXK1ydLkOv3FUbkKmmURGagpl1Su4+L
uTtdotgFLA2h4y5tHrViUaLBRzNc2VfNAXYF8yr2c1VU/RKCrq3Odz3Ork+mTUOCkwIHjhtFch5Z
kBG9C6p1warOeCISBggZK2H0BTfGNF8n6XY2W43EAeSTwRhzm74oxWe9wuuFtlO02O4OlTuKtgMv
3zivSr+BSEd4R2juMnFZqomdh4cbtj/c7KtKFMF0Eld4VumD1KIGCMrAgRrsaaPRL5fhdll284XS
R1bDZtccx03+jPMwsJI2GVAbHRWT2ExA83NHIOPI5q/7Jo8cH4R9znkXex/FopzT4PIAcnaMPrcs
zLN7dfygPf+PhRcffVsk7mzC9zwY9A9+7f91Ouplm7laNr4NssZoNjeJobWIeIoSOg6iMa4QInTA
N0ShDaMDxLyGptz0jn6838Mkw86ob2LSHyMcQpvkuguZ6p3kDoSH4Dfw3cA61N5tne3Fepkqvvfe
cYoxhFwaIbfANy1NqIB0ozHKeuS4yrZYhNCbCrpgtGY+qDACfWlweFLSVFs0SQJ3LzzioXCw9B6W
wkWc3wU/+cL6SdL9TQP/0HnU4PZnNwN+FdUWkUiJjSgCXG8pY3mo7kP3Jz0ztjifBGH/EajfKMol
dqGpjsDfkjtYnhj6O5rAkLqsfXtLQaLPObAut0nrP6++76dQ9MV4tRbT/Hr3pWqqP+gck0Lid+In
Xs6KsLbDJjk9ccKWiBkRLigzxJ08ylf9sRdBKcN3FThupYEFMw8oGPcBml290U17cL3RiKgAteR7
qmcDZ2NB5IiVW46iLfeXTf5h1C7pDFBqYK9ICg/25wTFZQcvpkWS6wOiuzsCHT4sZKC3O7VjgW8D
mmO/jeufDvqrgthVpsGSHU7Zi8c9719bvCIzd4BxqTLZtgpfYjaNstnHqbfYRZxbW2l732KjGEit
e67da9m9dobgrG/uoYf60JMx/+uGO0iyGflJwHOzJErrB2M0AR4XLLFtQZF7CYA2IAwer3Ci0Y8P
22zLC00TrujXQgzeDxl6HRGkqnCKghtndAPIotXeoqxpDxbZSnFsoqnaCyz99raaWE8i6xyYpKnJ
jew0sBXZHYa/g161dLctTgOJtMOH92BGWeMZ2YK1DSrtIVRVsb+RsNaQkNTRU1S/V7SWKBbBahYp
PHYdm9atPKujVJ3NDef9V+7YOSEPDzCta+qBIj4hmjcV2hZdY16ndHk669aqtkK48IY8qnN4i6kD
3ExXSqaXvMLsVNtsPb4wopcs5Xqp1lwFs7eWhVWZGaobrOU/a1tSmVdo4k9xr4Azvt+B1IyWd1gL
F/5npjH3WWmBtY4rzPnCkinRd0MEC+6lpLm5JLSaxSGm2JScndu0YP/5qbJdDNaX2XPMK+ut5uCv
r9aVrARIzzOr3pLw8K2+h+abIKNb22apt1Xh2XpKgIr4JUxy4VszYV1F1ynDN3Ta1fIdLMdFiTrt
yBBiJI6wYotDakxt2nQDSEM/fFZLVUsFTlPKO7BTZbcxssA3UikyzyQvF5HzA4qzm5c7ufhIbnOA
l5qn6sq3xa8I70OuL3f0gTpmX7KY04wlzt3o/feJj/Wg3/DTvLDteRr/bpB92Zs2V1KQpPMB8oZb
BscnQ1/N4zXBw/Jatt57Y0QhtrfCf7lqqx99M1gSfke98QO/kOAxEQiiO+csoSD2AVl7tqBRNT5l
8MVWq+ksS/rkmi2/Ix7n4u5Lv+I69xaVcDf/keN1+ZdtkUf0wpEW9DcjhBeeZHDefCyRUBAh56MH
JYevXJuOFeipbEqlU7M8XteaRmouwBosqUusgvIZMX66jWTLYfprCtSS6Xq9Kgp6gPOX+h27X+5I
iDSWWqMS+LRB0wbgBexLrGQ2OkyJ/5cFgQThbo5PxHchM7N7dMDmF18fa/fHTzzKtHzTqBWW4EZP
oGIMoPORD6BjMxfq7FiJMtVk5/iaBbcSVznfwGEC4JvU2o8btgd6blDbsO4oWkHPnaL2G7lxw1Hp
ACTcAO5x9/B5wFmfIim2WnNncvt//ETtAID29o9kMHWIuThvi0mnJvJktMZ7Yp5vhSpfJEoHTl/z
ibNBh7xKoh289+AKd4xT+nYzU+sCmVokv/h/Etw499ErxWXz3dP9JoswdkFHQYKwM9+08O9WZmTL
nXVwocYMxHRTQ5wEbhlOe7OwZQhpPyT9N3mbWsNlmFFZKTmsEpn4ZzqLKhDMeFWvvsk5ljU+Bl+J
XFQaCTnUswz6jnM3jGBJBB3ANsbUBpD5oOw0N3zi0O1L/toKw1g3IPphDR/Dyjp3UzVXfSOUTs17
cEnG3O2qclKQlCVBLmTh2fEqXgdthadApYOp1K+eRRsZNaz5N+w8G4hCaboN5t7E/zTE3IzLtZeW
4z8q9B5gygkKiBdxRjkxTNYaVwV8mG02M2GHIWK7o8rXtCnQgjKSGnNpTPhD6mMIVd+d973Zrx6q
sT+a/VOuXUk8Q5YZcpJxxcZfw3xzSZhG5lHYvRUndVpuCeARWnMZ4wCA/93LnmtrGHl8u37rebxp
MzXNyZ80psBhcH7bpFVd3aIl6eb22+BYPQhBsVQpvfu080fBFb6ndDn93DrRH1fDu6Wq8cKxVmKG
skx+mGs1wesNJgm44iyjUhEb8bjVrtXvv/olurYn1DqeNlKk3HsK1GLp4m16FNxWPyQ09RR+7XsS
Wa/VS4Sc+fJRFt0KR5Nmwjd/U4pC4eheMnZ+jYLFBSmjQ+azYt5F49dl4McE8PyVRgMmS/7Lsr2O
T/6nGMRQzlnzo+cwnYGgOpBvBL8AbmQ4WAh6a75EyAGDo083kvdIfL1VKki2q+D0Ek/gmbmoO6Gr
mDykt+fG+7KK0e5Il78r/hEaBqpqE1SKqtXPCJD7hSpRdj4dZIuAesUuFoiCsJKgw2VifXlJzgfc
hrFFY++7+6lbqMsSbFzbRm4uYekce2X7jsSyndyp3/blsiRFJnYORva4bZx/aY7Bovf7D2EoP3xf
ocVPUyvT6XDsPHbf1sVWgJ1qMneay24k/jIY3Meo6Lsl8lmVMQCEOd/VhoN85dLwiXks7WWIbgZ/
COAL1g8gqo0wHxOfMDpqL3UxKuV/BtswDR1HTdkz6jY+UrBVJZl19LI1jegKhM3j0wbAJJQZ+Ydp
z7aRfIHCwlOkUPxXL6reJSwuaLmnCX5LFnm+1t8I9Fa+Yaa6Wr6bLzZq1GCWipiyPPTRN0N7iGqX
TsLzxskEpozpqQ3UKs0vbQi7csxRysnyZXWBbzxH4BLdlanfXuMr25JUR16ugTqxLVImmsRVO3kR
Mvaz72jh9a1wiNEokqc4+X8vwkKRf9R/PwTdZTIR7k0wLTLcafqgGTtdZaNu9fUxZ/Js68bo4qQr
YFXnbE3RUcUJ1UU/UC9G/QaYqF/TFjtld4HWAWD3w5WLbOe9aIKV0y2hYrmCBR3XquPTTIrUlZzB
73PZeXRBfh+T4DXcheYqZtVU/MjUPdsHksuj/7dkjGwl/+a2oQl519g03NI+hdk+yPCxiJ9KVXrU
4cPB6G6Yw8nsdHpnPsLfdrkM6DTEpoTR0nCNA4p4hE8q4djwkAHCniFRfwLorUcB6+BmIuNLpBTh
XAs21QCFi75uOsLi986gU/M4ippF/K7bxbSP2mDYw3C9AjP0kPTXYoVFfQFVjueQ/a8l6wTqsf1f
7JANHEYBU6qTulybEAYurgi0NzL8gYoChCx432ooiVlis5Y3V1agOKRkqPKLelEgEipoRwrE2BJP
EnoBBQmY09ZCCiCHtdnuqctTFmqfyUxa8uFR0UGtCPc8YhdZ5ERmGQS3/G8ncs/Lfh576U70H3HF
GSQJFlrGd+n4mokOrWcYRexkV6atiMXmIcQVkij504tQeo+ZhxqC0mWXWnWoKYj2PH8s1YD8AT8m
VgXsN2T271FBvAj6Sa8YX0ddCLelMDP55z4YW+XyGpkeIQYWsCs5WoLN+3vJKZssV6vOUCgHv2PF
QdTEbpWiYVwti1IN7Z7hT/cda38EsBZJt+J27wUKGsIyCSHjfYrYZP7VKXQKucscJp6MHsmqFYs4
t7ZZ9JcrSi6PbBtlao8TF1+jnWS+M0ly8KvfmmnxUjzYEgCLByVcPdOjxz8OtLootuta74y10ZNi
giRkQlIdyulHTNgtDCR9wajicHlpL3ey60HL94TpHOZGgWyYHEyVQaUIeteBzYYqXEe+x85bKveP
mcq8tExSv2OdMVsWWNmA0Ofzyp3hjNXkQscDVKPnN8ZQJRMwm1POFK/PHdJ6HADqgEH8qrfio9eL
PVBTWsnSNLe2cuAFyResaN643q3E+VmS44/iw0SUROTW0JjbnNEvsPgmGGxIn15XTvUIGY4hna33
xcS3b8G0SMen5gu18Fz0iz43iNPxOxvKmxrPreSBqiOrobk1SYPIL7dtd3xhEih3dw8I4awcn/GP
UPBmCwx7V9gahe8Uj2I1J3RgWRo11om+kbxXtLd8Bx4rDAiPY3z5wWYDh9eBazzfkXRpACJRHzoj
7G7qc8koF9D+JCeO06QYVEmSFHbB/s1HLXBw3RYKzcPCeH/xOgogdPovgLLhjZmok7A/eqLLL/Gr
b29NCR40+T09ISokfc5QeLs+97Pjrahx+GR53WnrMThJGzn6w4wH644pOB3uzZixtgJ43mfHbUeO
S2jHvrpYAxUM3gIFuxKMhdcIX/vsSVO7M4XUMno1QBgxKktcDAGyzwaiyE536afeTPETEwUW4OcM
qAVKHw0CnKc11vgY07/fc3I288cS7T54Bd7bO6vidcf4Ht78apa7o8g8wByG6r0Y4PFphOhdoDlI
na0FgiH9rukKPXHJjIr6wWVfHP6IpyvGJtuK5QMYhPQb5poAgPwPjob2jMhPsv7fUSbiDuDBSNVY
+XJ3t7AXq+ChPNMBqjW23eGUI7MMnS3t9z3baEWBOE7Hwu62X0EhNr6AD8PVbMtjbhBs/EEY39WY
8b+W62/HS2+Uc5O4EH0DHI6vb83aLU4hEL66JStfk+CGn+3Zv755mMFBnYCUWD7rXikxk/qkNk6U
RjEiEsbuz1ntICdMnwkTKnQHw9lajfxA+bsq1YXvnUnheLnMqCq/rIieONACletG429Wnw3n8H2Q
50a28dpSsz1cPuhjdhdM1E5R3GTyQJXhPQyUQOkK4yyIbwYuHf6/wfc8HiD24XAnkFgHKDBtlnnu
d8/mVQytd7z+UsEFw2goSs8TkVMqtOi5GB510KB79TmHMmZqZBanwDKjvEBpGBuusKOxfU+OTUPg
ibYrZ1o8btuwThbhBYpI0YjLQkZziT5YqeaBpAhCHdZSqRvWaOYPfIRJfXRfiOGy7XXrD6xscE42
kSZcoeQDhY7R7ZgQn828E/muzAB5kHCShlE0U1HU+WI0A1GS9BBEsmsHjOQ2FAqJX78Jqq3mI9MB
vz9IRZ31ienUIy2KXPS3rtaptNSlYuNWM053kWNZXYm+IkiqBI0JvjIfrLyN4eGbHJqpUh6NORHI
kfDK+Jpx2M8UEnX5BdH5fj4BfaqKVzLfhqFMORjuwSd2hxRoYfsdF/q7hwusTfE5RbqlRGVh9bmJ
veDd04wm9iPUnblP7Tq2hBHSGo2ObpYn9/74mWnjgGmQW0grl9hOu8uY08EVTFzJPWXQMUvqUAjS
i1V3Zj+l4ZiVwE5Db5jR6kTjjeqFizjNoWM+QN3lO2Ioy6DQl9X7bJoC3rz+ySBuXdx9vzDCIZVW
y4KczsvB5lR0y0iHKcrBL1ITSWnrDjrjrb0/m/dI/0W0n1UOLSAe1SP/qYUhNBX1c4KJbV3/XHeV
hoCQuVyTNhaNnoeQ9o1Km36lDSNupSmzbYzbVIgKJOoLOEHyO22+IxHgP8cF/QBxIecPTFeH6jWF
xM6rShTDF9xmiIzGXmRRsMfPFfZkWtpMp++3Gel850F4+6NqOUao/y4PKwSdmTfzEY8gt6tNn+5j
Kzw6NT6P134EvY2ALJrbOyhttevoidETydEp6q/UaVuMuKMwFpQbuAiw/Y3UkEa6K6zH3a0X6l8g
StAj1F2e1Nfb19j9d0F8hp8ED+awFAfNAICBhHsC4o65aQ1z25fWhP7nML9BmZ3FNcfb083nql7Z
Abz1qoliyB4fP2pKLTIQzcXS40WdpU+Y04LFRnesy2IUm0aKKOw+BowlGj7ZBV8hVdZ4eJZZCrnK
qlvnteP4M8p4rGDl+OCVa1Ua2wJ0XIGfqfnrJ7FS4IXvil6wXlNOI3y/1eyHVz/IxBM79iBm69Dj
My9wqa0D4Np9kgbtUCNC7SZICgQXVTrPuYQnIFnapiaIIhzDp733TBQ9JJexfAAG198Xwb+YsoLN
PIvR2XA8hqwT+D98v0kOgoqORlbmhM/jIzXcGOstkWQBljozB6bpqkKhbJyW16DmBonE/qVGSrwi
WTy6fIt5jcMgxhWGyUn0tOD6/gGzgR+8DsiDb3BO/WHM+uJseXbA5f4O4cuzuMKoXQ4xbForHEWB
+mGIdksOUVlqPCd8gvXGcPt1/jhXRC+XIQ0g0OFHtmHWifnuirNZkCg5SlqsiCgtCJqjeD91wY0C
+l5bBG3iZCpbd8rYLxcTtafeJ2TbiQjqtTQ0zGkY7d+C0/ezrtWy3+YFGWROOYs67ftyokrZvjg6
5QO0mv5DJCthliy2e8auqf/hdISVon165sB+leFRMyghBwJEow15u7WKR1leIbLedaOWEe0ebaAT
H+FrGNN66cslwHzQsaP4jEF6NF//DI6s521Ryv/NiPnhkZOzRiDxtKeu5cyIAyXfkoRJRqzXvxUv
OAwbJSVRAOk1XCi2LRsUwTTmdC10vWkXXNvbYWaAdJRv9y2jNlpebzOCNA4fe6EipC4wDSvgM7x8
psalElkeze5x2yQFXSuoyVTIB6XNYDw5pbtcucgHQisHXqo5fbmLQ2Si0AS6t+BLM+qe2fT9xbvj
stvXy8RSNhzU6hIhjIIFszYyeMfVv+8T8B4kb830SCTnUasf2VTcF4BHeoAGmM7k46x1hH1TkFT7
wMMptjaUEdDh0lCoTFWqPPVJOS6ACd/kSSxCm57mXcGW+bv1xhAPVGqV/ILMeUn+t3m4WsN6cl/J
4S0SayaOJ57D8a3s/SPp2JDtPoILQ5tjdunXik6pG2hsTzAlT00X5ru1VhVLM3QeHWTnMVv317a4
JXyUPfjSGXhO/eyXiBygv7fInNQV2Ow6g2nVIZkNQgjF/4hFNEOcbp2tpchhWrhaL9kRt1blZUJH
PeMsoWqsXmdogExpnsJoA3I98SCQvujrTJyrJ0g9qreiodlgYBS4hhHqRuBxFuiIO5G9sDoIr1u4
4+LnKaPOdx2cUDc+dR3ix1soHmoFFy8Sp6DAMtHpk6SMe6cC3+7fTk4nugFOdkup2GulnhpgKD0D
jpQjFQHp8zfjgXnyJMLuMkOPPKuV9l0o1h3h0mVJIJinKcXg7csusQmn3tjc1SCX0oS0FS0gMBNq
I2NwoejnB8tAoiuulZVQifxXOzotx89KNZyW9e9uLJ/UkfR80Qs5nZplVxO59bDHdBaqxTo/eocE
o8MOy65aF0EK3VbIO0pz5KRIZ6L0+QIKIhSEmeZfY9V3VocBkcikEusmn3rWhablUjOlLRKxNmsR
IB+tgM8KZRkoAef3XjoglEY478M96xWghb9rQ+iKFIC7yWwvYWbvQgGfyHG4KEdASPaH7tjDTO6Z
w8OE0m7aSOB2uQDhyrRpnCfkRzeT8hoEu9bFpmtcBjddeFc/ZhDDAB15MhWAysafJvxZAwpnIlzi
G+zaIi0Kt/mJhShBq6w0xWBwhPwpgtZkwri3/pOmrsthmaFiXvc3111E4O/qCgrwWfjcBK/g37a7
YMFiKNkl9emUnkj7iYL9NbreJG26hh5Gzah00AYTk4wfyZkspqryILGt5e7b9txmVrTX/k90WGGY
hu0hyuKQBPMckBoBlnzCMHsPWi+2kkm6JzBvkZIgN2GVaxyrob17dE3cQurED1hVxFgsv/e9atK7
WuqJHQ5eyASJm30tBfqNBvXapOBLOCtM8zjmgTaFnQRd+cWqiKvnYquIoNhvjSMlnEq3jvHeW9Og
m2v7saQNnVvs0GmTZnw6cz431Zo/ssEOXK370XGnQXLPrLzXm2yhxhOKMZXVhLcmIqvjUu37mINm
pZpfC068Uuqm4yyfbX+D8ocd0Y1skPzaTQTRthMrT1jpyPlPw2sYZAnPwNmdh3hknE0ct4RRCsY4
6mQ0o1r2ExYJRE9QyVwyeuCNllvio7fQQzdQyzq3QEEf2xv2mhWV/7rw5LySkozo4G5qtxlzWErj
smpZLtGbPRMpgXv3OMYRJyJzQ21Df/zZ7oOPqJT/6T15/f5JtT2E7r9SBAaEVsVFHRULiq0JKvwc
0b5ETlTz9H6aDFFFIf5nw897dNJbE2Nv+xnWnv/5VN19aCGcdu1lWO2LxnpwfGTLRZr3jhwjlBzU
oEk8wwBLU62CIKrexu/0Aw+43r8R/DvCxNhiob56zFb5NQon3ix7pDhfW/6Cjau5vehLyA8EgSIT
kReaNXZ/9okgbgaXUmPbDPiR2AmPobe98t/mMKZbrOnFu13pmcGo+K2MDbQHMDn9n0rYzBFW+J1x
zJaSyh1Uado/DjsH324DuZuMMCwt5XnoQSOIZDzsX5oW+1+wu6gYpz+TZUwgbz/c2ia3zUC59fH+
M4xVuCgD9Q01wAWhFqx21PZePaD1yF5/VOAo7EukmPrJ9kACjM1EkYo+e55NCF0h04cY0+BS2olu
oW9BVgCnjnoq5FiXT0INxNR1YjiZABcUBt2iP+d84pi9UklJlEhTZb2NLYSNEJlLwo8Su8t+5D4C
JWvfYJ/rJonu3dWPitfsJ2KssBkzDWV3pY1I5IpFTrKph2ssjaM3HQi2tpKCHllkHX5vgyuugyxG
XBPe1PWb2iIkeHyUWm9KPNkVfRIZ9kGODFPgSY3EO9+OGQDVNlmH7EwfOiSg7Zh4+v3/l4e+KTxh
4pCm85wa5C5b0YF1py6yEC+pXi1zDDGBdqedXZO7KyCf9buwmEo/s/nazBfd4bnRT5yfxKZjG/pJ
AqB3cJ0oNVh6xwh8yh9V5kGcuYEYd7AOZruM1hT1ryZVP4E+ejq7Z1vubtBqrxCYcYKfqKFrWpT3
14QCE+wT8mlaUZlv11nitgSHozgiKW7kHQI93tUND1qnW5jyoKfdQ4QGppZUNwg74cD5PEfvSdmZ
5TrokA9ZJ4+RP7dQ9adhodGiRfHPIaADq5HLYUtzFHil93gXtOSnYnGLASxdVQxxafxgSWyeKQHV
cBuHUisnqZ6O3oY1MfEtx9tLIPC7+I+TKWHPItvDviaJvb/gqFEXs0rlPAj3AMY7EN4zWLO8i+yP
YLlFFKWFActECMQEVJp3FGaRT6Y/Pz52awoIM6MP5T84XdhaKIXBYzeHSwmBWoGBOtRmnongXZUy
DiB+LDEhiI7FAslyI0ZDoWpr/aYltXrfXG3Y0o/NhryMp4a64GW2azy8ym/lhv5nsrsIvlTZei/C
iH++zLTwZGiXtiKoCMHyiBLB1qePFtRs8Q+QoJa3dLdaf5ipnDy5KLGdcXvgJTRR7oQUlSAn6wgg
mHCcn4QFF1gkCdAfcD+F26p7cKGu5CJLUg07JQesXK6VuHWeXjTeWp6tNiLm+yG6wGvCgfb6OapD
jJSO1srelJKPSp6lIrrLdN58aiFmqUpD9PxV+iaSOMbwLMls94tpxdPaPq88BJlQQGe3Ni3rn7mV
i2taXk2pjighKCBiNqxqlKMvmK1ic3d/sbB7wgbOeU5h+jmi3S3I1qBSZbJSoUXBBmNdMt/Mru97
vho8wbcroFPdn6J57GowJd4dOQ/ZBoeC/3HlqOfn0Z9qrsint/436cOJGGS7oqFXj7gETit9iotx
1NZjziJXZEH01BIqAhVl7zZQqz6vFBlgPz2lItwD4+ajegBrJf8wRWsYsrtFrSZQ5mWeH5L9ALIb
ZlOIoYPhgcbDwf+xIjVJOWsn78Mbr62dOKHZtb+l8PH6e4ODx4mnTn15RFJG5QmlPFJdQFZdAZG+
A06+sWlohKMB/5HFGvKKIHy1cuKiyEEMBfUbC1LZuVYlUUTEqDrvM31zHjG8aI0Jwgo+lKbEWJZ3
jmnruzkPzVcVNh5qXUIY/H20eIPkhAQxB1+DVampq/I5ddH4kCe1NTIZ+MCZSsBvIY5dpo1rNNM6
ocBhlLz9OpzFOeusbmJ2CJfndfwRx3JsH529414EShROxpXxxXG3f90/XcyVs8v/pcjq0NVS6c8U
i2DKp4Yc6MHQtNUH+4X4T83j1REnN+/CClWNv5HPjIb1d0L9QA2QP5q8u70Jp43nvZXng/GHR1Wv
ciPp36JBF8BKzmWXfX9M4aljKEphHFoi5bNUTDrn/2xnnOwjilvDzETeWCZTjqK6yXuyKt/IMZVP
MnIaUJYDpjgNTnAnTAA+XTsBCyQ9WjSarOT4NkfGutjlDozAJ9+ixWm56s40tQOF6Mor+eQHPVOa
Y7ao3bP2O8Ge8MSUg84foTFeo/yN9n82NI1c+PqZ+sPgQCBvOHebZizAJ2w8JXrKNpTx2NRFx9bs
YnjLlUWz/l3qfg1tih5gHAJNRMK1ASEFedcS8vhYVGO73u4aa2c3h2VgjU8zVYBEjFh19Cr6cORt
Uutzd5DcY1zMTft8rwWBdJ+dPrt61s7xGco1v+rEA9Ttd/l5zmZUMN+qeTyTuvXREbIBURf6Bt+V
DWs9ttM1wYvmDd9nkLIZt59zGHqRSYxEPLsPMaM8FML+MxWcmZH1zYD6TNTckIS2dg8cXYLjzc/2
Jx54u5r24NGUIyoyJmo19xXrB0aTVV/lp0+XapVz8Z+GRHUWYjL8qmFM7PN/Ygmz5WWIeMROs05H
xC1M3wvaItJ5IrqlSr7BQLMYKrBuB1QvJ/xHvoHAa5bic4SEJ7mV+mTMbMMNQynhFJ/z8UQtVIfb
WtoB22zvs3mjYOSJocAAre/CjbzpQMxBppS2rsAeDlxwGT2Ndj4JIHZhBf8ygPLgX5myNLjpze+J
7Pr6D/of6f9QVgkMnsNwjiaYRfDlhaxuRmA0DWO3dIc+uWLe759D8sbXcS8bFLy06/qAWl/b9tS9
foA6ykipUA8rcYSCBc7CjRcbPAtXEuSppYREBiIu7bNx1pujrSC/0f+faQ9pvnEd//ATlI3HcMYv
L7tkNaWcjn+iy26mL5hMvVpHbMLjJMpxwdJTJd7zOhS7fTTdRDxNc5vHhZq93H2iBpHVOPdZkj99
nN5KhYUjV2Unoy6IuQ/FcmAdfl61YTxthig/K3wt7UCCkwBEkPa8fB7oXrGX7HwSshnpbRFSqoqx
2QfHqwQQxPeIKrWv1XdLZ0HYLHBvx/vxBQtzXIWaJbtqOlnhhyl//mTqhxllex0V1id+AJqFD/MW
DS2i0JzcGy2Dp+vSnr/SqlrzmTjs70dm5tt9VWQItz+FHel/iXgF84swL0yEXeszQ7l3Sv1Z9x9w
1wCZEKRwkZz1brl/zUWTSXjUwK+66hwgm//y0ClG5Sjfri4GxvPLSY+t/UlW2xjtvZlER5puB56Z
BwpcTpg1F7qR2JvhZDKXcWP++qX9om0mQ4kRhOkhtaDW7to4g/aWOQj2a4sKn0EDKcWa5dLWxhBf
ZdgjyNRoMqdOZv8ndZyq+7aJp1cK2Mgllp8krI5kj2wdNu2sJvfpOhv0OHkDQK6rxn6ewyAz15C7
3S/j16tGOT/OHhdCzweWt0KrcsRd0VYguHkbxb+1/ThzZolfHZOp5gNyn99mVm/bOE7/22uLzJad
ThT0O0mu1G3deS2OrqU74DqhfCJ1cRYL9zpZd2vM5DWUNdtt9VeM/SxLkOuWRBuyL1d6hSyyyZ8C
p6qavK1kws1/6O9FHNvgHPy2cV7WPyfw4lFSKKgmLQguUTTprojGCiN0vq/VMCe+pXTpdjuflzLK
5cf3UhqTygYbDeNZgAIbMH+4R/t+bCT1F6ZjbJ+YKL2JTQMKS+EjerlTuvSQA/oiRm2LdnoZWU0j
OE+u6Hc6dNar4qvZLeIYHOAgfVWwML/GPbwEs4R3l1YRiWGZ8aTM8Md0zQfvMMO+ZC9wylNpW8pY
tofMYvO9BYnWvNaC4xiaWSWQOjgJwkfZCD37iXJ6k6vV517sT/RKaLPEc9uuRRAjILnLl6xyENWX
u2hIpXNNUPayhdezyLjYg7qi/0u8hYjvx3AUoEMoeJeP+KSy1AQyiK2w4fK42DarP8Y/pn8k3Jfj
3hsCuXALN7S3kM4ZWPzb/anIP+2CTNPDc8jqXYMts8RWUOgel9/ruxFnlaMESmag614Su4Ak/Ftb
etffhvdsWS32YlwzX5Fvha/YtWftbXXgiQeaDCFyXXo8KFwjtpp/zbVBocAcd8wzp/rfhb3Fscfn
V2iZt0m9HE1P7Qvj6F9AlVrMORZqamVYqNW674wOWjjnwj2lKLt+jbLMpK8/Q7wR0SHc+ZPlxKP1
C0fP2wia1OWGbWctQ38bwDAMtH8fFDBLG8zqYrEhdQuADEBzAt9vOE3Y1vjRzv2MMWOp2DCA2dff
XXgp0N48XAhLMU6i0hfC9Iyoum+8ac0KuP2GEoqC80TwmWF4Gyfx69yJjIDUNkeK1/HjIUkxo/3H
zp9P0tF+N8kCsjEE2YcMUKeGFFLXgMxW0T5wr6mRtt1CkzEgPakVAMfR4GB0NFeq1RNRSKkZoPGP
EdIhSbZycJ0gU4YJTX4XiK2BQwKNJRAOrSrpi4djbmoPWWf6s1Qc6Gg5HbNDDMwNTol7dphV1ks2
/I/l0oCu/yOmIg8yxFu1wKWQRZS4+P7TrCTg498gkHCMlVCvZCk+Yjp2ghBRLs0+SrnYiOOCqu4x
/kWQgT6TXcIy77wpAVLvQ7pw9EiX/mO1vr74CINXaPBDlxrSL7m+tabGPp90de3OqrAHtNqD2RZA
gnqrP7DqL4Bw8LcVcHUyu2BwlyHbLCN/CYUN3qVQtLvVO4rMbQ96VEMPHu6UsOuGVhFrpym6kpSb
PY9lmhNvn9e155Nafe5j6aY75Ue++A3RjabshK26MitvjkJHN+dvui54WnGwbza7nz+yCVc2y5lo
xCeguc2RhhTLi4b/Fv/3APKBD5VkjLBynRmdn6ndjwqVv/wftdx4wFVv77J4x2l31zhFDFLiLcO6
bKx2QjdqkVylOSGiyf4cc3QIerAnXC70dexl9an2mA691PXctUJNFd22PHqOUBH1TheNlZ7CbBGS
YOqDMb52+xpDxGfwg1lSLcOFOTnOZfcGcZRvNL5ri+jYsmX8FHqAT2uJmyALdVKQHIs+83r5+e4i
18YMXCc2zyK5HT91d2f7pHpjiccpU3jeIT276W+UuTHEUgFKst3g6XHwIDIpxrZQtO/DV6xalmAJ
6oci+/ogth+OSCrSCVNyGcHL7DMX+tXDyZ+IaeerNemt2+AkwYII0Ienkx+f1k7/Y2U9H9HEa2AT
OD4kSg1uFGeTDfdGtyG/BNOQ05ZzxDWxnnau3zrxtLM8WS2Ud/E9qg0P90ayWKQmOrqx1t5eun7R
i0Y7xFwi2wZhT+rmPPvEshYQd3USi/E6UQ6WJcg3sTY5DgGZKZpMd27cdacTyTVHwKhT8MVDo2/X
SPty9ClcqoELd7CYApMqQICJi8peyscBhKlDk/shdmrX9feRwypEWGX3ZEWVEw59miAbI1KlIVHv
HIiCRYOgBY9ej0iINxY9BytTAm0VrqfmNIUxwCmq7MK9uo3oAndLplK5OByCgPb6e61kURdMnVWK
V7Fa92cT6olLfD46oMdBJKJ6TO1RKQvK71a9EKdUAOuxkWTuxpADOz2jEuKeqJgm5sBHg+N2bVt2
pv1GTadgG9BVA5RNHJrEP3SsiKwcKNoUH0o9e+a44GpMph302qPnlS6XjtVfS1Hp/yiIa6amBMJm
k5SMzqJjb0ejNI4PPDet+lQoFTET4beJtv6cjtL91OSOxlu1Nl7RzBxDyHeWqtVMDuyhYE9Wwyvn
sLPa7tncqRbtGPVioBgXA9OPuDjvaUGvOqxQrCM4LlvDcTW1fb1xTOjicV9G8G89O3rGmYNe1NBy
xsaPdUYm0sVSPQO0X2NfqlcC+40MAyDDpDepRL5t1TF39rSD7dmlE8JMJIDi9CkK2zDjReEpNpub
nwNK94vtLeTRdlQl8yiqY7yHyGTj4oLPmkVJg6bobWRe8zJIMiYCgBNlgYvgQRmiqHoJ62abxWHD
+ASl/5wA46XxbvGycD9hOwmTVXNJkgis7+RG8AeKjK2hGvaL7JtLBLxGumIg8E9yHjANE2tk7B1v
ScemehvM1ZLGzSz5Xfc0hJyE9Bc2pniYGquhQ8c1aMittMYHnvsVBNRQxmYuTAI4nn8Xkrd8bwb5
sIC83lGRKG6y5x37sEuEwef/BUSHGwJAxabwzDj1Z/k/8KIk4WubrOT/NO7xywi8KG9iqsKuj8cF
dNwDF5hCpvZNqL2yu7vDApkHHla+4QOU+9UiD/YMsPRhykOay85hnPd0o7x9KrZDV/Z1qAwmlcV+
7pJh5jrxOH57mwRWEsaqL/mKHGGXTdobYgO5B2ULX2jHox5KV5QPzsU67XCNtDPZDWtSVf1Gqz2+
2w7xS6IHYI85yVtZyW8P/MxwUVBQ1PqLukXZV40xxxSVt7jpF86fIJSsJ0JIA0RUb/rz49Jkq7wa
vVxSAqXSpnlm7hSNtrqkW2in8mmes+rMFA0TnaFgnnxfAN4GeIYDH7Rt3UguWkbQW+gtb/BaBj0Z
WrYt5Mn+DonNyk9m/YtgKjwIly5DqFhPaUtOsdF0bCCRN5r8c3IW7z62DCAEGKC3b61/qw6hYu+f
ef5CsrmpNZoCXW0a7yZ46U2k99aZ5wfttecANZa67SZAFWi795PACKzAeNEEzI9An/MpaCuXquQq
/dZIjD7oio/1eZs1FNng4dwuxb3CoFL3tXs7dvlJlhvs/zcuC/26IWOB+Oyuin1ojDw23pibe7EK
cFShYP2RC83g1o7hWpTBC6xjZm6r/YCLB2BJUwrTyt76kE5Y2nqaY3FOoaKjhvPKztclf7EkRmhX
Dti3WojCGdicihO1YcuYTMqSL5RpYga29QRZMF1V1M3p1mogV23jCVnisbkUv5aqJrspDgc+Bqqq
egi6FE64E6V4I6441R5lngmZDjiisjyv3ClbCqpk3HdXpbd0yJ3q68GglzmCoZ2whszlfdTWMY2E
J3/Ml4vIvu+6LJ8EVZVZuE3XG8gVVt03isiU/DD/e/pdzPPV/YMQb9H1MdNds1HT2VjkE58mhRSR
UL7h327bd6Hb/SonqFW3AdOrQvB5rd28s1xE5mTS968Gqg66aWCFsazj1fUjs5Mrj5bw5VShYSV4
2bXf2Sn/8b8d3HogvM2FjsVf5SdCBJAKEOUR91q09FHHEbEy+CPF7/QzwaeUQi1sDmRSKgKt6MZX
xMKulrMWw8RpR+K6VNu4RZUZADfInkvfzXb6cGDiNkTLUfQUgu8hhaYzhzb8mquMniRLdjupP7J2
E5bdVNL9j48Ze83BUbmMFQkNXMeAqCiMtuJHuHKKEBRChENcxubuq9lC/poJ/ZOj4LGWhgsJ3Myq
EfKmsLvCkiNVvig3yWLUSS0O/B68tIjHWa70fRAsYl7yhIZbBYb7pbu+22YQj3vRh4g4vqgi+6hC
jNJiyu3OH/EMbTG846b9VAdZ1bwvngwkwp9ZcXjmu5YfUEy0OxwmIpLUe4qUwliUncxztIAUW5H+
u6C7NjoDrE+QgCgRcxqXiehLwCwsxmsImpeCJ99LamEAUFJ6TIq99JS5k4xZPAC8sp4585VCCrN/
6PgWpdw9Do7CHVUqoNc3vOVThFQGrFMTYaz8SDq958Flq/n/3zE6GJ4rtqsjKndO0KDO3AkMjtJb
tF7H1pzRBXL+HQ0eSH/rFEhZucSeQzb396j/+w6R1ttcahxd4yUfIVOg8B4U/RVOZSxnOCoeAFrm
/ZYxHSagYnvCsDW0c2c0Im5MiJdNNic2USARo6f0Nv0WwYfo39Ao99M56HR3nS5DCPCFFaB4z1y7
XFhRNjHcUZVvUQDxxCcVo32xTQHqC3Fd0Dug02PadjBQpw+xhfbk8fm/oNrxRTIgrF7ZN/UyTxj0
iCErdosVTqCSsXECwI9mav6LNv/0m1ehMpIFoN5ICsTXGxlQw4drL/de2KI3Z37+HV+atfljc8zz
OV8VIysNr87FpaX4Cdys78T978NhmtNxauVskvefsRs4EJra/0+24uaRtyp3HmpRCJ3Es8kJ4RVL
NM/l1fcQlR6d/yqsZYg0fsyO93ks3V9Y3mHI8FfYtax7JRJvqZpgja53rSQV7pzBdFSO4CuV0ZRs
cqZl007RaNoxwigtWde9MrI1HCZzwjf7hNy6TFhCUhS5KFMoS008tzTUL5Ue7pS2QJG/0kapvuVu
7lmaL/T+m2+9/nE755s4oN3wdVUktt7FYZ0CuCEouoM0mgPe5Kb0AcVT5T825BLRA+7cbUCDCLDU
GAlAP+z1PwkyCRSPH6LSn1R9A7Qg6yVQALO1Nm3DhKBk/1HxRjSC0z2HygYrGQKQSVkFCIJmbRsm
/K8nLrFUA479ERdC8aoJ/zWmTwjzbWrpvneFVZS1qEzaaK5b6MhesdCz4RXzbUZoT6aTcoc4ctXq
tHxlk62iPavRzkTkctMrX8/DY2e9YtBDVVdU+wnhelWs0SZt+j0LjU0jLjP8hLBUrRdXVdUJ3v3c
b9mz84BL7+qKCFwzLOcJQDNbGYH8+vrP8URorY4PE1Qvc2l68CVSSa84+NA0cxgsLARbJ/pJBZMz
6VOXc3E4GGBybK/TKCPvl98cxWf5Ir+XZefZXF0NKV2vsCcHcVzbzR5ojQoU05/OjJnHxH6/cUSh
IYtDEH5AF88roguWJ2ClCAzGomiM90qGGXSbsfXQx3tbaEk9m7KaylWOkzNbq4UcB957BtDwWrhd
KiBeS/5h5DKFZcSPc46+hBmsA/tNj4Mi1EbJkO2V3ECMktpIFfBUPJyov3f+fEpZPC0pWHXqrZG/
vDP4rsOslyUpfUd0vwL3xY4liGZoBUQoRTl69nJHfGhjQomejFg6tll8pr/aco1980s6iWRc2Jov
7Hpu1iQtOXCzUuf3gMXXhj9l3atcmUkKscTBJD4PsbIy9qIzJpkr543XlaPl4Lw5O/4bFUqNZVee
gq+jmCQenp4NkwJpNvTHWluEKfeWsRocVH3+O6Y5uvN1NjccTAhshgnkSzuQorfznxndxSJJ4jbH
tdYf1hzGtxn44ws9THnzn3LrNCJiSG7+dwof5Upr93feiX1HSauctnLtduVGpslDaeB3bmZ3bPRG
rO8cHghjNrlmth9WriAmR8P3vHeRe+dOZjNZHIl3L98m1sN/GWVkeXPSNlIC75+lS78YVYy/7XLY
1NDXi2NHu0sXC8TzYOUs+BDjF6TpLUofLSSvpHSPXWVkL8QDCcr0FP2ISD6epg5laC8XDWHtQ7NB
BYLHzn+csdJvFTuiwtFGLMiqv8KLinPSsXfBleFlqjmPG1S16jb6kTAogq2e8C8IJK8az0jkSX1k
Il2R2LP7RKM0VLEdLqaMSHbNR5ioJRdU8mTWws7lvTlBk08s3kThmlDeKyKlqYgJeolYYlIrrjSp
1FycgWkiJIZNdEuY0JhCs3SLCtQDskujJw2NDGArePncoPtanzZvvOHkruJ86AvWLH2Qxt3uhBV3
VUeJqf/0wsdfS1IcMOPiVjv9fjAVkCV4nHPJ8vdT4zVzJyRsZ10QP80OByTvvJ3PVNIrS8r15v3y
TbN70vWII9ifZVp3vzgryettYFN4sV5f5DrU5ZZQJPKDHfPwbwlOK98kNB/OhDPZ8rYv5bx9TJ9B
v29vMNZajK34C5efXRzaAFcsEB3X4mkTxgMpG/Izbs4aUh8QXUMN3juSxfegEzjFf/5IrAM7CPOl
GSKM4z+hBULdPRQI39wKK7NoT3SnCKAug2l8GCmvkppR4ST3A+xNiCqqJlT6eUFNk8INeGDD2Ot+
2fEmFkLTEgyncwmmgW+vdOo+tF9yEEM3mijbYn0xzGisvcpn7nX0KPDRaaajnN9ju7p9UFcE945s
mGfvgZFPBjIb4i5Z9/13xh6KNBoyM7Kvc9sFWK1oHUAoN+YAXj4Qnq8I1YQF7FWnTsfaXTMcZmPX
qvfriW6QjG9nvuTnqYny1ChLXWVL7up6EhXvxkSuKx5dEkiW7G2qxIf/AkWUUlVriYZj6M75qJyG
INP9tcLuK8adSr8AtmMNTcMuaOZiuU82yeOtO0s/F+97gjBnE3RzZWUw8dT18I+ngWR/k9m/A7Wx
ZIS99zTBXlxI6p6Hsvh0U71XugMSPykKq4DgmtMoz/VJvlYIMtz+sKv6kcwB8IBJ+i0dvo/pEflk
E4e8Kw3UYD+UJmhSY5abaDNTf/msMIyTsJMyzy772oT6YpwAbRk1wl0lIbo0cjLF1BS+TsHVgB/t
TmwB4OGkkL4OvcJ+GNvr4kt7fpP4RTnXRIXhtez7Dp7RLJ45KEMivL74xfqRMJcIhZBon07iW5yO
VCnhFK1CWdBXUyrvDXcfMWrw3x3Wxs+8x6H+zGnCZjMzB43rwTCupcFrHWojV/p4dxeNPmLX0cye
wdRULHdVRciEU3FrsWSV/moZubuIEr/cXs9O0kNij2ZMzjkDRXxAFFlbJMofRkXmiJggmiwz8MgH
JrqQGtn1uYtbckhq9glWI0fxdvfHJv9vUHmqihiA1txGau/XV8rSRY3ihkY8JRB01bAY7lWsBIuy
raQ7yIPezDExyLZWsHip99B1hDDkyB28PctFEner7XJ6fDPoi6LmDDW+HYhhwQM2wCO9KfmWee7B
ulYABQ+kgpIPMFcSXjsXJkISmLO8A7XfjwUwUiXY9yWfwkyDysY840nd6MzQ70IC6gBYstUFVPFb
5CvABtlDYzknPWduIp5ihJJ5EXV/1zmG2a1yhAWyU5p777xWUgl+ohRNPjpez4k2tv0QvSGsvioI
ulE/tINRw9ohLr9cUC3IYEFcb/HevQ+IkwSPPSvf2+sDHXYjPZJkqnwdgnQ/e+ARKOZv4Vw+FD5Y
cuxKomBEcdrBgmejWBYi4iVsI325dAcWntg/cJj51AAHP39OowCcWAlRNtsiaJBe69lOk5fSH1nE
oHtJGrBiQvAqLno7XpRl7S21oyVoOBEQ6+1mpvdaDJcvayMlM1yHTBplwVXjR93GYGJyU5OafKkA
rKwg5zC3y+cxs7a8l+8JGQvoiuokEe9BOS7/oHfZPC9q7RFZasVQLzMEQ1lu+XOLz8nQUs0cnqZI
Dd/RSsHGpYXemp54Y511rbncah7UGaxD8JVoLHtHMn5ZIAq4KiVDeCV2oqHVFcKQU2uff0yVAq0c
gBcTKlyiiEnKH0YhjC/UT4aqJ6XXzv4VFkheXEBmp/y061B4NEI5eItvTecaRK7IcyQr04XwJb+1
J1as/cTx+Qc+DEPq5uWTBTyWyjSB5GrnZwb1bJkn2Ge26Aym5UHlXkHaq72WRUnKzEf/c0KMrHLl
zcxELfplvtFTegDye2tuvo5QNcDEG1BCjwBkdbDsj3TV01R7mjqS0onSwGZlFYfUm4GUu2ZCcA12
jwqWsw+LZurbyhF8rNh1+LtPFAm64LiqpyW3sDUVrQaNBrPhuqGNguNfHQHU2wiWjhR1Mvesn0P2
gWxTNxzgw3FkLYrsTJ5vJ0kfN0OIGGi7KTZZFgv9peB42zwkpNENQdMLXhklc0lcHqQ5Z7R7SzDu
/6wrwkVO1n+iPmHTDWQFmalUdnDxBmc1Qo2QUetOHmFRb1PpDZicoQT3gDEGZu5BP8biwWX3JhSD
u9hLQs2sFZpkCLgKWMBCdHFATXoYUoQllHHRQ/Hpb69eLYm7NV5REnCcQ8BLKcOTqvFB9s7r2lfo
R8BFHJWdIPQ+7uW/ON3lvSOrtCJFim3RBadzxcTr3E8yqizuy4afkAc3wf8IEkQr497fkyz1RSbQ
ONYw9xuZWqS68nS8RPHbJS0OajPRFmINjaZU4VErMxO8J0q1pZkNI67jflUY2/eqRCV6HonpHLKq
6LFqnbs6BzConZC/LqDtyZqfa3hLMpk+jP+8mSmWA/9F4ibr4/xxV3oLfaLThtNIz6Nj1xYwACI7
01tIaLlLE4eJLwx8vxGskosWNauSNowy0kjp96Af4ZSz6BuCBhkjvPIWFH8f7oLcWkshal4hWRJ/
ywE6NssIoxLVeZ+ZEUct9f5YXLPasPRSenJZ4Zhe71P/3RiA3Ixzwel0VTuUCkZhn2ixvwirxwwa
Zfvlz0q4zrTnA8tmPwI+zENwWhxjDrEZLYMESasyhjEGBQOuYRKxZ5x4aMfIWOsru1bT8IC9opFd
zfwOduImAHv/70rCu5cAZ4r3MTo+G/RuxfYOaGvOL6wYYZJFDi2UxW0rC57B8hiBVEPg8rBY3GWS
7G13Grj6vdxt8jW7D/AZcH/DfZ2j94F1RtAKoUM2ilOfqltbuZy+z62QSfwmmdL9RwVt2nuL1U00
sHNqBcBH3HHQa4n8PH/hkxGF28rV/6BtLg7oj4O57vJ/6qF9BkL6OEVpWWUuXGP9vRMQxfGnWQ9J
c+91mbnPxugIGrc4eepA1XyDXXu/eklZBqzNGNEGReZAj8014bBxqZQ4maOxzBjG68rXGwZHg0Tn
AIv4DXIgzyKWj3iH1Zr5d9OiqiOWeNrI00LrVvS3wFSfB0g0kSwFX0w4tNgzXV3Slyv9PGlbjoYS
gzYLWQAnHhc/qebe4K1qjhlyGoaHSnWzEr/EyOwP2kdfeY7uejOtbCtaa5I4dsiaSFlmGc2FIkfr
aeExfI4U+aZ/okfWxCo3ZpYGSU2xQAcZz7C6mUV4jho34gexJJwxLMSnw/EK6Qs9F0Ry4GS6fyF0
fSsNe77Vy/NMBkxSwh3my8DjHjRT5i7RRZyoFfm/+ns79Lu4WAPVlFR17LE4YBM/VYcZU/OFG5fh
uLbIm1CEwfPmgbb6jPArpkCO50PsY17OOdN5R5Bj2VUf9pSPOtvIJUyX94nD4eo+axyMKtphYdwF
L0u1BZsblfSBkChuey0MrPZZ8r+QHDKXPk6v3UkilkTMxyXtEKHDZZCOoWhyb7gTCN640Ccixdji
nsV3+wyx8VN422NBMyS0wN7HR8iOzUlSm5oU4FPCUCsEC3DUUh3Q/BecHyQEH7r/O/yjogIFvUf+
M5ZRj1pUtpBhwu7sCfHkbNu2bCoX1v3Ha47A8hTjkFENSWBGfhu86EJPFZD0p6707G2UDVyVhITL
T1/Vpw9ooNZwjAzsG64catFkdrbN5+lDxH2Sz9I6KhR1iv9FXM/pA/22H2icObPXXi/Z4sGFP8Ww
pYH+nFW5b6PX7usQSth/x8qsykBa0wTCqsbJ5I3y2ogXLBO10uDdJylL/f6JTcpcq3tswNTWCcWG
aGaDsRHLlP+oKctfM5+3dMpu0QNJX1VTOT/l5iVYHRmDLcsY5FuyuQu4yYK3S9lIkdOh5+a0RVNb
yB9FmBD6+NolWXEBDlDOn3kd31cMVmh/jkuFh9WpoLOPEKxiSzXvIIiUFuucTpZbBPbzbZe9oSzz
cMzj23veLRPRBkyjmmntP+/2SOWCwtc9CbKbwiMEziTKQIbPO2lkn3uhPJTO0DJLcc2PFnr/lIAY
i5waAwz9pWla+z1t7aRXfvH2152vpg06zbqRXO8H2yoV4PPqJ18GLgIC4+x0UpGG/eBm/5leXNtG
cN5IkOuJ9/8qT3gXXpslrqHUCF6HzKAq1W7kRAXTHq5LfcMP7h6SPPA5cu5b6ibQW1+wD9Byd9M9
Emk2fQYzIXxHXv7NI9NaqZVHY8PrftKaWapp8dHWNZDifm47heB4EmYjfCuCni76GnznlfPLmwlC
BaZz7yID4CaIrfARDzJJerFzfX15LE4Ap59bzjeV2DReo2O9RUIR3BApMEGR//NycRvvHhKG6MBu
Bdibmk6NqRW0Ee4/wwzqLXgud4pMEjBvAxuCVHDySXT5el+7YYKJR3BgdRJoogEUNxoI4fzc5W5e
nDRidCHqvRB2McTINRJHbhM7V5pbY16O77wMYWbI7PGU7ozlH3vEtx4w2vj0kVIAZ3h+4O3AvLWt
YlA7mkrf80tIBANiYJbaCeLrjeqTpyXJ66xpX2v+n2hIm6RmCY6/GqRZdXo7JJSjUwWq0dv30nTR
bGBiPOBP7KdehmSlPqum9b/ZsXALvFHiptoNioRSL3FyF9b/IUpOUaTBUiE8dqEgFjPMX5FyxpwF
6jlsa6j2HY+uaIzZHOEfvHlF+1APyu3504tveeQig7w72K25I2HvEAFRf9qxb1e4zk8ZsUg+peXV
HCXSTc9kbCB3Z6hjfQ6qrPW9z5h96tQ39vSNHFIqwLPGpkipZzffW9Q2mQ9cZhSGBz8yLUubob4V
PMWNe2bl/bw5dT/a9m3aYKmyIoZvVyb7TqP9l3AFYZ/tyaOapMtKIrnmNC01jinXu2Y3xXkDQ02z
PB9Adiw7BXqZhzQSz8RcL0t8m0o1qb6wDxbwqkXwXEZx5GrlENi7b5YCAQguYyI4DSeO7j1bz3PS
K2kC6qzA+qOAQMJ9RzKtv63M8WvkYpaYb/xpzHwtXjos7qaiBeMcjcDhUjVzUZY8PVjq7sfntqLX
HkMp8RhLHs5Y1agEF62Tss9lnE1xIkxbbFD3l3MsabcBzz25eBSQxwaNfRlPT4Uj/VLH3no68GOS
cY9MTLKNgtrd/Ly9NRhQpCDrH9K/6FeQNkR59sJHcgn9vBQU/ZJHz67gTY7KwwnlbQKSISlIavn6
OsvZmI0GVd+GuMLzgSau8Um7LGRFKlerLDnzn45tUDVDLgKUK72BVIV3pJwCJ5cDNJ73He8aJxVj
NRWTFCdZukI0nRrFIjKYOJgCMaYmchX1ZNYu3CBRA+BapJ3rul5FWMVRvOzY02gVGxb6orUDIK/T
piBRYL+G2vKcF9RaGtku7KRq8ZDxhD1bakeZBQGWWNc6Rl0KgIP8gbjIQ52h0kJ4zV0DhHbe9b4j
RME/LIQXhGLRcSFY0Ej1XvIU42rA2Od3FNP+Ad3JATrUR1Z9TteMvH2ajpU7TAFNG3PCqnLM0AQ7
bSaI/tDJcNa42gCv4cpVqdW8xVjyJyEYu2vqz9trvB88woxxv/gXtp4bJ3kTSsfwBi5ANkZgvZ7S
cpULgKPwHOGTte/80+T47NTXBWKATc1YGCdGNifONSgFHUabUFZTSHDKbl9GwNImGRiCKh/iYqnc
lo6N2p+dOMjV/dCV0WSnRJBHdi7WUp5xAVPgNs5LUjrzinoJJTEZloEwQy2rai3IC6rynvLamsb/
r0msoA0ftEyiFI+aS8DQtWC2nUGeIJCDmCh06ncHLp6P1HUY2QqHA/Ce623mjCRKmmzLTIBdj4RP
QIQq21wwn6krXZBUD9LznGY/UwT8V2DMS0yzLN+FwRu2PCYGSDYA0DJDiETpP0FUFwJ2MvFvn/dQ
HlDhNG+5ggMhzVvg+qbAOxDah7sJVcOGvws7LDgTAG1MKsqov9z7Mo2AlPnA0QG6ljMb2YhcTZRf
zS2dabhXVg+VAzs19UHB+9RIVYARXJC9z6EFsq1NOFVx1rguXLUtqaNQM0sjrHLlxhZC51Idzk7J
/koM9uH/sNGl9aZOm4RB207AEy6yTjDJdzBrWeNoyb4I17yNH55XWo2UXzUvXrIZ1RnvPNo7CDUO
VvCJPW5BWg9SYRyLLiglGzgzTKiAgviTXN1bl2nIydNyRBULCFJe6DT3RCqL166GH7TMlvMLXBeK
Z/5JDrfCs8nNzXsm0cIE7pCp6uDwiW99oNvVjkA5dd/9aR16Ri45VncG6nRu18pMsxXSyzeuor+s
TA4LGKE/ENSVBgbN55cxXFqVIeFeeRSqv1ILyx9rJOaMIxo8GQqx9YMZYKG/FJoRiaSdsGOUriGy
FzsFquYNOJKdYQ3m7cHNT9HVXhFwte8wLcjvgQYAlPDX67ZJFWNEUSdbY7TpLXUUKSTiKdBRWD0m
/GmAd7KZv6Ef5Cql+GIlP1kvJfx42xBPRAOvSUAPBWbO1IVY4Rx4uVd88ekRzmqmcZxbMp3XhgH3
3Dxux2jd6VfrsM8f7lWDUc66n9ANmXZUK+GL4eV4ypM1QJT263RQyXaQ3/+1XIyWKtaHO7pLM4l6
dEiuT/WdwQcKkL9Lrik9gETBKDaOcToIpYvT+64wrWgcGUUFa9+ovsC01l8eaRC4zvUv9xhAvT9h
vOPUZbIgB+7pqBrr8QjF2uXqPsVSiHVITopzbosZg+rcjjak3Qqdjz8+uep0TZhqywyMAMJxjBgd
Y+noJDlrAMgorbzZMIjg2S+3Tu+/SDykTIZ5wtbxEPVv7CGAIbkB6k+tv8X6SiYj1S6GZ0yxudeo
ytz8/df1ZqTfHNrcKCaaTIJ+D2HauWRL7GZ9YK8WhWLQOvoWEony/YbIZG190Xsgi7LeY7GxrhBL
eAxOHc3XgiQd54xWyFnJJgOXKtFJg1JZcIZ55upAl0hJa9iQVi2tDXNEn5FdS2g30/KH4L8LfJaz
578NoYouhv17mpS5UUoLwjwkOlrVi1/3Shxcaf+H8TwgKXuuJ762JhcTRQrj0gFDpGng30lLyTRc
ofiGuWPWe62QfCm95+uvoVXxO2cYiicsF3IHyPNwrxpRQGOm9hVxBka07Juta9Klcb8Ew5WqppB4
+ZL/k4hS2YB4k7qmM481/d5w4xGxOwYwOxAzS6zSWa1i5qK4wk3Ozc3hDCdaDCukT4CUrSpVxK9o
THU0MTWTwQBK+bCcREbHbCE0bkm4EnbjFL+tMBttw7TGVekS09oLP4oLsN1gN3WLFFd4reVa4jzY
cqXOSyERIapTDJmmdYYf8zIKLZH5mvU4zAt+e5053c8JSC/lpxlYDivaQ0SAFhMzKKV9c/q6tAvo
a2N7UUzsE6Dk81G2EGRMnOz2b02JBZpjxmRbAgA5oWJSvEkpn282iT7KSIUDrhgx2M8+5n4erH+a
pluJ73kvR4w3Qc6WyjryWwf0t26S/2kEm/t2j8oS6wtb2R7njOmYSLo45xjbMiGft5AKHZp74YQg
8Ev2gQCRC0xCo7frs7IPEVn8SOCBMOaj4D7MWVjAXnfXaDQD1GewXYpDraE4ZINQOK1+/7e3T8cX
PlrjmpdU3OadatyDm9wMDObYo5GZCsUHdasxqpnvDQHoorMfiQoBQxlwifuy1V9wdcnxKUnNm2Vf
WfPzzIG4YSVr/1lZ8UtyOnQ9XDzHU+LEqDpFHjlCCqydR6EmQzxFPC4gly98NnTzFWbk0lYu0bX+
Akcn843Tx1Mjo6fWMW7dj80+T2ssNuQpjRvAaWv8Mr9YkXEAgmSIKwSramAxqZssBg6nLWQIoDGm
XCnGPbvePEtDNfoYeQqsPvhIzaGMq8/wr2yNCrr358Hk46Cs2bo/M2qPIDsfyRs2Pl2smpqHS6PX
MmKv80Bq+TmN38xz9GDMQAKUkxGFfFLiDzBjOAJUY6PJIaqfY7Spyx5P6DzvgjKEA/S8pl8VF96p
iGs218n2adI1zNyjifdHuOEgaVJ0QMRQdp7CILIGsCnpowg+vHMOYVr3GScmhe9pQUsJ7/TBdDH0
DlARpCNTB/5Lbzn4tk11FZVicDKO3IelppgeofpTi9xKbARVhomcr5GObelBV/LuCv/MpwjEVTrk
Gn3I/7WQThnkQtu0Mgs+sjfr6TYiYIoiGdRxCrDKQFhZxqWNUpf8pnWwcNMfuprTNTmWRQQWYhnu
hp8564Bbz/q0exvvOJwWeywGNuQharl2ExqMJh3dpPD60r8w6k9F8W3ogwF3jXMALDsLJVYtSx1+
ZalndpU4iMuPpXdbJAvd/pyhyeQ98nKOvyLdfKWJIT80vg2hLY+/eL6s89+moO73kXLJUAW+ZZbX
QLiI0QA8NnZ2ZROVvpaPvmoMEcg9LKxfAPMzzp8d0ID5hMQoySZsqsKlkXUF7z2zd/uvh2AHJwZ1
Sfsz/55znmA4OIXuwCQFAZuRZ+ue83iYa02jW981o0yGAvacpWB1La6CE3klv2SJ1YfmhyX2Uk5+
SVOQAug27z0GOUH8Rc4d27JO/tuYv2rTcfVxttvRL1Yo4r4GgU/nbcV//S1IL3049RuvnQ45GQQN
AHd4vdUL5vn8W+pqco2BSbt9AQkmkgBCX2Jp3sCjCQNGkLh849zPFfmsmHBPWisiIeP1wQjY+LxJ
AWBjTRSFSKZwqE8ELzuSm8uMzZVi+En45bYYGe3X1DMeqcvBPwAjCyMHtObTQRnXHoCnCPDMsFGY
0kKSIyak0dEuMFQ3h3H0d2RpFp4c1zhxiQOe3RYNX94DvsemVwx8n+dem0BVvagbeh3a3nfaxAU1
FJSctTFLmFIYqhrmW+K3Kevjv4IicjNLL1e/QkKaVNZZy+d+QIcrxqzMbvdHinaKWFniThR3RERJ
X3zuI/ojsvhxRpOGV8v1cl8bpYNueOwtCQ/xjWWiIvbggavRXJGxUDI7E/7icl1jG5tXgUHIAoe6
unuoOBPB/nF1qd1xhe+AtsKVqLdALVWz4fvwKuUVLPPqW5zTFUFeR3oEgqCotosyvcAaExCSmMAc
YzcFN/Q79hmuf/LDEpZ7ZsknuO19qu2UbjdH8gGwXWjJmxLMcMTKm0lHXvjLloFpsnOsqRXh8U4Q
l8SiOQNni56stR361naYliJExpvy9HheN1fqRHKZnAqRams+cy6rFheHnLaKVshsoFTjJs6cxnJ0
xeed93HNIpEi6TItnAKTVtIMjLkerlxgKgS76xlv0TU/gTw1SS+Sts6tXVweE2iNsWCIPKT792Zz
9lzwORt9vPqOaYE3ksCYDeK278qB1NLfCLoqavKw3JQfQ6iBh2PU7BTEqoXsMBHfXbQijtC9zjsM
ftjIY5Jh2Ya4IXMDPxLu2lrq/BR6cEePb8gSCkuxwGxnJhOYGaqjthsRPB65DGLOyNR3ILC3gkmS
ZoPO7yLHLd9P1brZ8WOiyzWNvEbPbrVKbOnzs0sJP2V9OkoLTq7lw+CQWl+l7PYpjfHY1kXedh4H
wJntn0dVWpz7I8tE5vg0c488YtK9l28Pqj0pzetrCn4V+y4dRuoxK9xpNvNwlgbFxyDOO+SJeLoV
wEGb//URE3h4iEce0oQjmyV+D1MPqgMc2SCfOeTuVDg4NZE4xDCT8vTxHvPGK3wgGIqnEDz2ZGMk
fs54CAzPZsVWYB6epewd+yl6QkJ7zk7JMpKqCxC4lOVTU0UEqXhIQWg69EdMOvQM7lPNfA+ES/Hb
hcyHYH07Q+F6RENv2CMq3KpoJRFR1zfIZa1kxpi/1EQVklqVbMTK59QCSE7tV0VqsjtfBWqhVuCW
oTEzjkHkkbwZTMBmg80lXZ9QYtgVIzKCt7jNiqcxq1OKxEQqEelp0gmkvuzTAHIpM6yiziT7uzvW
5FI+hlxPxSh2tOZEuan10jYwnKh251c8WNWZpXw6W55ZifV3YRX/DHVQquCU4tNo1DnRruH6UOuz
YDgUIxFrrxxsqPz2PusDa0S11IvStEN8q84UakL64qt3bo3D7qXQKuFNl4ine7ynHPKumCVC7r88
sIPfRqbayjTH8mNaIcVJtzsp+FmrqpKsSRhbzBb80fayPzG8bkglkHYZ8huapxiWec03CieUEGpl
wwxS8dmKdZuqdG3NLLnH+CTmTuMlFFCoUkJ2Rd1bqd0JLT4dlWDCHKO6M8thdFS89CU7tIaW6jil
pKFh1ikJ+Eav0nvzUgGZPBCzxcE1ktorxwQiqkm33d+lgVxvae95OAD1gOKezyejeMkRPeV+gZiT
M29wUndUOsHkmEd3y2Rdr2Z8CUJFtZRQc6Szz81wcXg9Y/c0iRXHZqKFkZZrt+5b0BKU5s1/tDbs
xrsCqbPHNIPuPOQkLJQ3/UsM7gXTcqnPCFIzwnZfzLQ+B59GedzRWwGvZRCq4PinDkUPvA3s+VNy
AC/9qqzamlAlMckKV0qh7EEcbvwKECn7VCRRyde7rvcaccnOY5dmDd5EO+NbJGxaKAokFpqhYW/A
8RspBNzIClkUGvwGUGbedHdBN6BqRRQ36ymZ+fgS5c8mdgvP0NVWl2fGvrixNUivou09uN44Ldbw
sDcpsiDtYfTgEP18FrNhWJvuBeq5WdK7TaDhABoqtcITSGnik9OyZnRNaJEWole/SDe+sipwAojx
kD9GE/rRG+5IAXmG6CDb07wiRCQQx2jjekCxSPge4zpmmZn1/kwXeOhRoC6bhn4e5bmS7J3whRys
ocskJnF2oFCDlYahDr0J9z8ysw9jd6Iu3h93ZaTvOnFV4XJv9+1PVINF+s9VQp1YJoW6moI0dA/B
1Cu+U4/caE/ScfTuTWC9lTAXsD40hdNuR9IwCp7M0oHw+Xfi4M4QL4XUolTYLqzEm0n6LaM+hvP8
+v5iaU3m+pOgRVa7mh1EXjnVVl+S2b3Lf4nPmyFD1x0Z0Ov6/2uA7Y+uICFIbjDIGvLz7LRrPWVg
0Gely5dSyJQMzz9ESHrPreR5b+Kp0HuD71L205v8PDmUi/7j432DnuvVFQ3adaLwvJLJQ3TwDYYs
cqui1sBRwhUptWkJ3Z7Jtds3A0EppPXibiII1B75SQVRivdYnh92YwmOZK7icSjoBb93H3Zfzdu0
oDytsIigBLaWEAF5faGTaUt3mdVJ4A+lVqdzpFQhx0u7tZCry0rxVU35vqsyDW/qsaIDuwKB+lfJ
xDVADS/9u1PJiYp8MsjWlbAZLkinEliHzUNMo86nEufjetsb2b6uC/3+EaQpAY2YsfPAzvpuHe6O
7g+9GDJEkP2pZpQ3u8N7F+hRTjkq2oFgufrU32VsWnm4Xsh57JroVC019EZbmMDwOs9H1184MLFz
2iVJFY7UoHTApfRIbN6nCYB5C37xC0KhbWwui67KEMyK7nDLJApPBa21dJwaOPKfnZIp2Fh+Kd0i
Dn8Xc201HP4aByaFDg1X4nW0xazNcX33w1+dOan/DZcZNgscW0yvLk0TwU9XHgTE49vLmOLGWGRY
G+iYFRFDNtz1/ipxaZ1LKBmN6i7v5aU4YXd5AYM0rQ97hGhngBSU+PYXU4EZdWynToqr+0IhLsIL
PGDti++DP0jr+F9+UIeK/eQVgmMuOWik1VqjvFPWlCynf7z+3TiUfV2sLnVw8/WOaubefMHQE1NE
+DOANBce5swEJrrrDst3PJrfCqeacQd0gCyA91b1+ECsao7yOUGzoma5ycyvVnOrVuAViDaaB+kI
PkuUo+vbXnGbHTSWOPYeDxWtbAAbDub8NhPPQPhv+AFqciSs+9YnFUpTNKzYjnW4zN7J3m0yan8S
eWF0w7b7UuST5emjpU53nZgH294x9tPIHUitpQMHDsNcuKOyOgk53eTC5n+eZWOo/A9Czce9uF6p
dS+Il+pZxn60P2XhZl9hLqL2zLQMpVNSCZrst3jvZSzuvlzSR0nGltQz/zrvYLTVbiHZ0k1gu0Yf
qMvmZ/WpqK8IZlX8ZSkxOPkYO68VLhKUSz3NHzRWE2COz/6RfkvsWY/E1CyqvGtqKpBF4gcaKX+K
03vX33+hHiUT61PYLHKKunUBJbqCXSed/Au+wOmR0yBI9gMmFEPL+Ad6pC6aEMhAWUnCnTKwEkhA
0SsMo+KPUh0p+0ysfJ8X+EV0/OykNc9M4Xi5z7cBjA9B0fqosghjAuPczOzeuD6zJe+7mU0oMypA
OBACsttcsljzKakptxkPezdXwcEzGnBrC82dSV/GQ5VIeiCP1Nr+W8JrJPQLRZkWapoF1tRFhAXo
yMfcTxnX1p7Hlj40Vg7ZVNNZQEWrMPeNBE8Ku4SaxQhi91r2n8P+VQEvO7Fr+VoqLL/O5n9OJAXG
zdwgt8WDLySnYCRVCip1v4bO8XTOPlhloEM1lBTPtg5ldFWoU3DFMNN+F4qO57UQyIw606ZJFncq
h+EsFnLp/+9b4oahIe8QDHSGJzORyNOcBnh06biSrRhYJm2g51wwmdbNtcXAf/TqRgvbh33u0aYD
22+sSgfevrc2r0Ac5WnDiEChAeHP29iLnChL78ieCJ1b9ho0C4DqzlJ4TjeBKbNX/q22xd6EsMHH
F6H9nH2ByG8i1K5k3O2VmWIk1vsiMbk2jkl3W27hi70qg+6T0Uk24VUckuwPcKxLwbkWj4BwwVY5
QL17JzNPx0R80h03Fkmm0oN+375iAhlkjYT2vzct1Z+gQxaDUfdict12+CxVjdNeA7bqp66sMZu0
PUzoYozoCOCL5Xm4XMSU/lQ9ih9xB394HbXJg7EF48jc99Sa5ruAxOgk1wS5SMDLQNRdjCC4XSre
t4AY9QuSGM8gA6jtJxXy6ab6CVKmLqAqtgDTua2cB8VQgIB6UpHXAsn1f5KkkkwXTpckPx87u0EU
r/9ZaKZi7EJMAY8psmEZr39d+FG1Xl2mM+40lgpvWUSwNeXvqXNm73jh6o9TSkME5jmF3bW+Adrf
wEl3dvv9rlLzifZXbuteZ7F3iQfMlPuBeGPOgnTmioAiC9BHq+JcePaCVyIecD3f3H6uDxdWDW/3
ifPec2MyAZKmBb2U2/ukpQ0WdL3VxlTz9VHpZ9Wpw2pNftEXnXs6q+we1Q2DknPKWaBbVRIpDAro
2Esy1nHoPJU1BW3k/fbuYvntZn4MvE3nXPCNvY2+3aRIDHuUOww0Cyn3zSxB2oOT4KyetpZP9J5H
3GnNDWt/gTQUSotb2cXvgA+JQw1yM/3w5MV9DxoSYbcUa8y4BgGVBtPC+NVGRusZ8H+zjMjNT62X
8vohrr/JxdpQxw0rlZJwYOMzhOcs5qqeVw3UGhIit4aIR/gGpIb2psQcak28c2HASJhd28JsIFlh
PMvterpLLhYUD7XzMR2iVZgYSNW1pByGLfVwMGuZ9jO9Yvij46VnlmdFUNeeLzyepol/jDYzQgS7
QzW9hF1Ux/ndDw3W8wwwL8H1U58MayAjd2BasO6/AYtY9exGD+ORqTn7v6C/tY/o7dLVg7M+gaqQ
NH9CF2nvD+T44Es3NpBm88HcpHkaDsLVuudMxuZL5+DR21p88dF3zupecxG5xbBVHo0B0/KtS0PV
0I8BLNzLc+N+5G703uzyTFmuMEofN0axKSLPUmv3DlcCsqTWOk9iCh4uKETcBpEs4YhG9lfSkDwv
QLD+HOhAJJlc4+F6Vo4DDCtTX1kTQu4wM5AygPU745QKtqeXHa5fHoN/aLHdmZ6n5gc3WilweZJJ
njDqEQNIcXei0QItjmvgZI2+lXIe1TbuHi5EDljRpRyHjyEvOXqkgDDFM0NZpn4Oa4XbWmWBMzKN
oSD3OamKPzNaQM5HB/YK8icvLecnzY7Tv5iTB/FhSChvZTgS5eHzbRcTAEtjMARUDzA2aHQl5EXX
iWpdEF2GBRarkn9blyalOXF3ANpSOQh+AeI537JqUvURp3NMg4GpQeFM8GosF6MYgDCm8DYYp5Ly
VUVcq4TOxL1VHMfmplZblBfO9Y/T2GywQ7+2VLkgayPsQ4Ury7bNhcBBOiJNET9BOwgvXqDNy149
oEeODX90hUHMwSskzZyc62pThRxyjtgf3ey9smwB/uS/cccXF//ENBB/hGsFrBwQ1kyLbL/0h84O
saYc1HiUBu9a6H0NngNKomK06qiEYamORwg5xRMFzJboS8SyYlJcHrJqSW8sx9TZ6uJ9JhUOK42Y
iGlz9Dw8cHT5azuFxfZuGDxtVHOtkPbWF+xMMZT4hcf3GehkGdRsEutXYcumWPuPo+MI2DlfMHTJ
hYG3qwrYqP6WfEjOhKJfzB8ksxLOYqj0ZNioSU1R0xVeWzE12Y87rVO+6C/rkFfxX6OvWzDTZvy3
lhaH/a/m7cJp7gFoK7VIBcK8M/rYztj53s/0Z67RR2HUtkzTGhZls8MTXQSPAVE427cpTDYTwwxU
viac/MqrvDsMM5IvEQnNde9RN+Jz0yVIYJk7bTZLjs8SRUIeWcmhRbOgsUp6SsICyOwU/Pp0TjyW
4hCKeFgrzE4VJ9OEFriQKc5H78MmcpbaOkyi6xg4wxyl4xtTC+A/YEsFYz/8PJ9zCqq+0771Rrkc
HZISQFwCEzr4OP3J4m78iyXYgbbUO/UJ6qNbMHWR1c5Auhq7ZvhESb3me4QrI+kFJZGQT6J95I5j
MX1zIKPlyoUDfvdFHLlr+Q8rLYSDY5FUu3pG5RC1fQt97PB1bzqxcuAwvgfPLJNofLtvwlfHLeWb
+iIuCgTR/uW/fCy/betC6uqRmqocNaRbYGfW2ef4cx+KtSi9hDX9o8PbTFQ3eB2k8CpjtQlzOXIC
uTPzzE/5eiOyplAIYriRIjRDWckzgXBZYr5e1BVHSWArQ3xYAJG6jpO/vLEqnj2zexfOqlftK8x4
g3H7PiQXnm3p4tsG99FlkCaAQqmwdXjwp2RhqnUFa0GOxwlIqvpwdgN0mBCSPFczWEkSRDlNkiyK
Q49vOh1Kga6BgDfGJyZOW7tNsh1c8YnC+ajGi46nWkB7um1HXZLm3M76Qv6JyEtepGO27ecKfZi8
1uXf3GB/7QFffeCtUx3RZ12HrZzJsC4brQverIknRdYApBpkRurb+qggt59DDrbj84/y9h3wX9gw
nBZVXrw8z4RCBfANZxk9k69NS86Yhr+hV3+n+UqHjxiYs4xhZo8xGp4JjMA2Nm6ZqmikgdiVR6tO
F6ZJfvl16i1/i8+A/v8QC3b1/Wis6y9O4kkM3ALNWpOkIlf9G1np+JiHWKZDnKb8oIUZpZSi8yod
WqHbuPcxIA92CAWKGXv7+XWXiBRUCmWgc28nbuT86uOc5a/R7l1Xrr1GahH8a1+NvETutILMM8DF
vSTa66nQnNxrTYMTz5QJO6J8YG53xltB1LhqjsZT3qBmlJOAehyuOH+/5DhTIR+khrW1ia+32g8y
ChkddChoKNbGGZojMZhgkcDqxZOqQ9WnYF1I9VS/wb4rSmftuk7QPD3/Iu8X28DR87qxT7kVNZ48
L2ltfJVVaB8RE1/rEamGi+qn+w/wW6+izdAJOhr440O9pTRy13bILhbUGI+yqOwzlS3XV3UQzd/q
KzXvrEVLNZA882ILA3m7di8KTkETuZKEE+313j4jNmvHZqOqeTcR8OQ59rrDJ/13b4WyG3dNj7yX
Kt8GEKpZsKt/O7fOKhFfeciAYDodjj5RuifNVBpfn4L34ezD8YdQ5BCZ7U5pUD7YGUsZlZ84GXoR
+L31bMdm5RkdKj9EzqIQMLyvjs+MqQsxr9G25XMj08tcr2QP4+jwJ46lysHZxkF7+8vo3J2Ae78U
jGkolGRnlkBG7kiNvxoqWrtfiXY+4l463XFTmJKQvD+w79oPcm6MW81h/0tVKErGzKb5HHfEJK/1
ojSAyPgkwB/Mt2X/ToLlzqVy5NaZBek7xKNbB2coHPyL4nhBd5R2y/gl3spqHE2c3aX9cjLr98Wq
amiCnK9RBijaZKhBfOF9pL+SM5W0rPlSXRBgyFOoleXVqe7s1RtIYZhf3B/vbRN1Lxc5xSwTZUA3
R3jFYm0mCoXvFU0SkETw2evgCz4oQW5PecG7aKM6c4ukJnoBIBxnWZgUUkRXmZjbeFjdreabKG3S
K5W32Wciria6i5qWvZg7ePKOxRSZonHtNtlr/us9tpqjfxgt3rcgKkza9yzDjfFTYXxsYJNm3TGS
5tgTb3NU3pbG/tp1HQTudm+xxH2HBe0IRStvFf0zVuCvqXemeoU3ftZ5689Cjhu74Xazw3HLdzoS
hqlc0hZ6lksYiWS5/zKpgumc0kYxvthiKvNxf9kH6IPRs21VqGk/L4n6lbxGhnobUb7gZzKEgeLw
y2n/MgMjdemeTa3N6UjmVGmz0yXQmWM5+kvrfY0M+qZIbLVgvvKZtxUCqqlkp+5iTWazOiTBTfc4
h+jzPv9mDLblvWpVpQ87MqSz9atkgSCCRB3OUyzV2eTGlAGSvJ0PanX8sGKvAq6Qefvuv66gpG6y
kQusPRULt5yBeWmQGCmVL69N6G8/JBYy+moB4aPeWxUhDExu6aaAOmGx23qMBG32EGxSAMRC+jVj
sL6umZQyYxKRimYBk6b5dRps82hvpbpBT2ry3ZgUYgYK8M3WBd6METMh2CUO5KOSsaoHtxEIaTY4
ZcavsIJTMRORKjwsqlGdAtUd/EcCVMeJJdat2xtFPdtla1QsNKhMz5SrsDnjOSbMKkjYpptd891i
dMzjuNT40J+qSEJgBeMjB9h7cEPI+TRrVXAdLLA0GXbHWREEJp9v/N3uytR3etPErtYHGDM4zOR4
fvqUruhAWkThjYrwQKXWQO80GubCBsCyLDe5TpVQt4yXYFXTSHrwKxQw58SxwfPhwpfCbaoi8yw/
d8lZROCe+PcroCIPybCpahFiUb67Wnzd3jrg+CUxAf0DEG3B8zYhEwIDaQ/JFgGX8LBwL9hmoXFY
PWzpTKWPKbk5e5rxxKyZLv3D6JnEawtorppVI0QMVJFAd3j9CA/js7sha2og7wABiPYBwz+hktNT
q0DpzQIAyvEvkmJ9X2OUCjiiaSMsuZWOhnX44sws2ScddHG9YaT7+lJBsnAgreaYBoIpT23BlOFk
TkcI+zeqcocxWOzg7buosRcRnNgSuFz1tRItxtJXo9Q1WkGjtmYLN+JAwCF5K+G1f68OwGZSQBK7
qnpEj250djg1ke2peB/g4j0RJwP9AeGAZ1YNlx6s7qh8l/+e9QuS6Ov09rbTh/t8IE5AoaTmmoVp
GRfp2HtxQClBq3ciYWRbzvodokFvfadqWuDAkxR08hfR2P6grb2wZHDskZcJqUIBju/mG5HBeG2V
CafTug0JVOsijg/cDPocg4YWgpQkrViOFsnQySRwQrboKY+uwh3ykxWrSeYlQidMpyYgMlT2oeku
BdaHQr9gmBsu/jh1x6aYJhheUi7e5mO1sO3SiOfH6flunzOVRjQRHI9yg+lODebyZAsut5eiZCH6
qzU0nEfvfUy8uct9egEuX7h49nSJEEKXuYzYo5pbhoeYECmrwYwy5G+UFntG8yZ+sm12NcpwwbJo
aJAjWJpCSUWcSYQ0K6PkXORW3BRCWmv9VrIvHQSyMCy+Tk93hbPGbfNosMVtlcUnT+uIkZtr+ejp
sJihuR3Yb7Lm9qPuw17ibsKQLrir+exW42cYhstcvsRbaYOQXddmTM56SsnfX3ikv10kjHI5u0kE
WVgq6kfDS4KL49zxEVN9dR/JJNCxktdYwX3eOgX0zJWa2RnjiHbz0qbSb3iPhiCq9HJGO18BJ1dm
TB3PSqc/CtsdsMoSEhA57O4BzmAc4HSV6o4vCtcq4qJ8qYeOkoULDHsA/hn+Opfu1bH/qN9SO4fj
tbvhPs/KzzwB38TbYxRQJOoj3Hy2oOUwIb7VQbTD9C2ON7lR8rOGzqXe7B7RoAKkgABpp8zwnyC6
0BjioQsZ7hxz01QWnLdliYYdVxHe+qjAyxzc36PmJDP//YoE3gRWX5Cxz//78JPxQL8MCcnabWh2
ZdwnLGb3VnasKujoOG6H6gTs1zJt3lBbMFX+sbgTCHuiGUp39cB5zko5zkR5WKrw3odLhLf3vgQk
byMUUU+d+qFax972Qj8MTtJacjYiMXZ6uRgWS4O60bUQicNNz3dFjiyGApbY5CnNMLW+6EC48wmI
/7EYRRkjIzOFpi3WhYZ+1+S82Onh0Z4JkTBZzngnLwdt6lrm4UYnJ0pQp8n6IdJiGvCo072Wx+5w
VuUhMxB9jCJt4dYycGi8vTEHOAStARd+gqkXFB4bTS3Fedsb1RBvHIPEE5E3WCIcabkQmyfT6TFZ
+EoJmH5/ljE+LEpI82wBenEg7c9ier7e21sLYUXLsfBv8z0u7xXHuysXTfWkFFqkJs58B67RdiyV
sifiz6gvG4li+FMGI4j0F7rSizzxBAOCeGIPtYAJtIK+2CtrT6LOC9djc4T5lh7O+DpQZuTmbw6a
aEE+qivSdqIMwbS8MwtvaLHIIsfmXExO9i3cAgieM06TGlOMg2ve8iUqgfMploYuVVS+PeDfRgKB
+sp6aQ1cvxr0B8TiqGuxIVFksBSDVpcPvmx04U7YEs9EifJwBBVBCgZkEbgxAJVC5vVJBuFeE1os
kyYgIfqtcfhu2X8veTT5eTSp5gIQbWxoyqHKniqhHmWY6K5fNRovcLs9mEiCD9Y5FKnHsiiB9Yoi
UyqbW/44VrGIrYUKT8o12Smzpc3WN9hVpwca2TWBc91rOeyRiNaLF7kOZ5eexldAQ7ohjmKOH5m1
IkMxtxwl8VWfa8JMlzvg7PMl1qG6/Z6qIp1+s/S3mmF9UGJ6Cs+mRLhjzyl2BBC9qSOK90KEjwcV
Kjwhqgo5frM1D5plydoQNDNy3jDMgT1rk83nFE1kgH1XJ3V4Bl7LtO461xvRh5OFoDjXObQNxCrY
OC6tT9q6itr/SSgf1xG1TPoyPoZnPA27Uhevh6zRtB+NOKtq37TQyozPI+QeXpkMaIVKKb42KJif
EbMDHzfsEqahbeNaiiqyFX9XPIxgDSsH6dtnWOKI91zhhDfPYqbjf+jfWL6ZXEenGc7WlSgcsoRU
344+IvBO53rkuMvLtuTEvgGm/9qcgGLBzOSZd4HsYcQqs8YCt9ew8yZIbkP2bdNC4ETlPJ+usGId
8i/rQW1p1/P9IgKsrBeNVMQ1NpbzOdFPYp+mTr4PUpkW4rD/OAn1jAaDvbl8SKHGMVIMZKK1VWTy
kd8Bt5CteUC451OtTQ870cynDOJI7Ahty/uWE3Kq2W6jXMteKfTEr7exUd7IQPTduDNRJA8bjuOi
WoUCJDaBk7o4TZCdzX5GsFubT0UTrELxFCygQ1m7SdMOjGpTEDQhjCBSTP9kczOFo8jcnFkquHLD
qi5ADoqky+8903mz7BEFRk5cx2bdgQLhfwn20Mfhq5ziSuQuuoXhGPhlP2S2ErBazFuSmNaHgKwg
5EazI2cb+2jED2lXpjX7Yis/IhCXNEW356NsieyatmVPgAUvVHgmySCJYruNFtpqtWHgwMCBn0rv
9sm7+cQ1PmNk+oUkBSfDbq+VFSnEM+x1Jj5PiscGHoXAx9oEQMe4h/LvyEzh+QfgSYeGD9DwalFS
EXw3RZa7DxKHloUkUIxeDM/gD1t8aaSE9/etdMinduVOlA+JjmEJNG/vsAjWiiFq42xpHB6tEYU2
0fzwN5bOkok1n3voY8RZLffpbSqOq8dNQB2yc5Mf/8BFX9/VbSI3bjZ5Q+cwZpwNhHgtLcTDMxfn
VGQhTTfy8uCdYqmHQzsYBLsFSdwUX8WmsqEjAhrnMrT1Eoj4z/sZLCW5TYxpm5yM89ZfIE9rg5bE
7TFmbw6Z7pIAcDxBV37UvFNGZuRZutd9nLnZ4hBnXhZ3KkprXPTrpDfop3TCDw2ickm6D+6cS8VN
TOwKkbsTGF6gE70SjHjM9Bb75HtXbBiGCQt+h1OG/K8chfV77X1F1mHMPyfRU0KEAj3KZtAU9cAs
0tmKtj3H19Mvj8+5lWDNu54H/Kh4i4RJXpHL1+i4iDt5XBkBaEE1VAeW1ZDxAopeReRS8oks5wbf
OOhvX1WKCD1YqBgaNVheZyhay/amkJd9JBIezKatuTJHiChDYuvuyxZfriSmZaVmtXN/7gGBUmvk
vJuDTylrkp4nMorUTYGU8ApqE7rwft8DUJvd3jlxjxj0eVej7Z7qwqoyAEMvthL6YrFbVpWxiYOl
Tv5XeD+RlQBLfzlD1XYJyohqEvkXPPyuISMWxbld+2yK2w6ISswuPLs25eYEPv/1njT86gywCgNA
gqOCJVYtrB8w9+9s1sDHwQ6ayF8eMgxJfNCGnYmhYM0blijSYc9JtLgrJ3sl94GYKmuLuBtMUtSc
+Xj0x2MhQgZoysSUJ6pNV0woWeapj2KUWS4KwTHyT3P9VSMWEafaQMTD0OE6VUfNRulrhEjuGP9M
gJKOk8YLIfUc/+yLFSCiX/ha7jKTXaRJT5k3D4BrMurGbp20ECkyujc03ZDHag/zdXYzYDJngH+h
wQKHSobnbfVUdJSEPiBIMIiAGu2TPPegeEwQCNMf/nX1+S9FGlG/C33zDH9b+o+e+0k390/FZfHI
vGWnSZlZ/taVYe2mHXFQZ+EftMtra3a5s7abe9a3g71MX4hTp00AXIqeXqsMXf6nmP60+65yR+9v
LaQuEOXvOsQwlchnm0JsjJjD8uyw8Fw3QowmgQG9Vni4YgYvw2W4RAfOWfcEJwzEMPdDMCXE+pZW
1V2TdDystsmOvhfU8nFkW9nrYVMAfy0zjUrNr3yzCKXqcmFZ2TqrIdW36wJPPGHW5+X2H7cA/dEC
0b1PG7eWWSsj4o8yQzui9dAltpVpUa8Cmh2zJOe1G8mkDcgOrNhvo4qxJhB6PynDa3f0rgGdwr7e
dFPARY4pNKXdLZbBnVRMfkINq6p6KOVSaHsm2SR/AjE9g7c1DG5vKuWEHE9Wk4Sqtfu3N4xNs7sF
J9zdEz6BZnp309vC5/61Z7/pXAB1eFhUxD967mkgQWHRH+FQsubRI13dAWfHITPomcXUjoUHcr6i
5ynCQMUxThU4BPiEUMfZPNGgJDShgk+YrExmcXu32CW2kGYIH9a+mTKzQQurOft3lyGXEr7pPKN9
jO7ADb0hV27xTkB97lsVHyCOjnpRoC3UJy7e+aLM/Y50P7PV9w3ne7+8hkorQqss/vmunTLEpUBO
1keXLRKvPD7d8j6WJIlEm98QuRPHZdmT3UmrPpQSVL+THcCm6kZV3d5YthuqYQXZSLXqYtrs6PcE
SLifYDtS/E28rvIDw7WXIGM7TUBv6i0nJKMIWB0MNCvcgOvE5uL3a72fc72jvKW4M6rnrHfiNGAn
7QXWhWn8BU2W4QuiiclW5wxurguG4gZt2FsMcZlPElXE26wREZLT7A2gV9twb7BKiAa7lDAyoOYs
eyUBURCdvy4Yh7qfa3bJCuhEr715z/K8twqYD1WkgV9l95ldDe4gjW9jT/cpZhObQWx3MLGE0AEM
zF+3jS0uT8SAsGELKEoXY8AkCr8PE2Vsj8ObkE2G95tyFQ1MgFcnIR1QrlCz2qNCkgtLo2RFlsxS
t+6nM0LHzPGkhmkZaU2vrMnMtbtHCEVGSf4Z+nr+ZVGQUr9AU9ScaD/XUtXtAfQIL7n4g74TujaR
88mIZJPubjJKJaiClIcuUwvMscd9PdtFzC1IezuL2gOsGBqMq0IaS1LHnmk6Te12iSy4Sw0wsFj0
CJCHPJf5Nz9Tf2xnJvEYEILI3uCyHGRG3EcVZlQEZ2XTnRnKq92bdWr+AIkeLgQNKMG52zEON3cD
mmPNVxRjKUdTr6YTUENnxK7ENoFpueAjfBcvLJawtSTSK9YZHGvKbmrwPzKbMdwEB95hWK/G4dmf
Dcu7REE4Wf7XemnWFL7L7xRMCPZDwBXscmMkdv+N7zARYkj4V2XC0QkShkPKoQmj5kuTt1BO5/kr
dzVo3180By8q+cvzJYbcapfs70WXQ/1duMewWfBd+MkXr/oR2nxIltQUISjpm2ofSZJPvF7Nshda
GcAvTApgHQ04Opu/RoJL+B1eperBq1DhhSxGgFly5AxCN3zaN2WzYziDq+GHIguJ0euFc5w9vhx7
+68XuVWTu/f/1ux+6EnJaRaXFVUjYTeoC/0gf+hCyn+pSBuCfFUZW/r5n5g+Wyuxz44mUacJ55Zg
ivQniJitah5KErjU9/OEHP5vKdDRWDePP0ipZUvedvcoS8WaMGpKiKrX87caCm0xmq+dHZv8LDm6
vROXDwETixXmNbhFNNPhr4lN8OSVm1ojSL1fOGLWBTqyWI5zgtQRdPY7U/hAgFW0Tk7dVYAnrxdX
zsrLIJ+i/tVXz3ntqBf+3UjLhAXGDgIbDIyOLic0lgNAo13cAOS1F2sX6/jemIYPk8Qjr4/jePJw
6+TBg5HcLyWmmZgpVcIKEdIJmGuOt58pNssCQeuwU7o+W1G//sFLkctSynQzGI+b1gcJCJvXYglU
9e7SeTsdBPfBC1ihUusW9oI8dTd0WAGgT9WVRr/yvMnw4PdPz2zHHMG3hhucJK2u9OCWWOwi2yQF
C6qzghN28mAK1XSVHwc0TUzj2NegLqZyWwi6U1LuWUbmTpU31sF8Kf7taPlXEzoTodUQmzpeGDRV
NtNHruId/9rDynHRySmHBZVGp+gJtD43lLFoZYPh80v+9GxDAYaOdJA81YefWrjFI9b1Jf2cm6xx
h+y+9OHBsCny0iWOfkwq2LTCYDOFM30aEtMCSMJ2+wUJcM7p9hAu7BQwHmhFWmtGAEGyJjpWVrif
7yXOY712BiInPkmhcDC+3X8BW9fD5W5Xgaj/+M9IqgI+U5vefPXjkOK5SbaL2eKbN9YXXY480I3P
GSQRdYW6Wd7i+K5EOX+zJr1/qZH0Yx3SGITH2qE9DEAezsBRssF54jNvvVOdNcU9cOQD5Zhkicza
QPOXrGpTf75Ts7JGP08nyuBuR5+hvVjpVWtyl0evPHOR1NmjGbLmG/NyPdHcxMWb+zy+NCrajjef
pOg4DEhYqJGmghzTdYmFLORrGzpeaEjoLOg2YoPuXTr8pdUt+iGhSU8SAIHLLfL23L+ZcstfszJp
uaPUO0hxYSG/E442RTWvO8KFfuhzRmdpKw9XtzcRaHgY899LiioYxWz8h1iMv1RyAH4XibNInp6D
g+pfcxpOZ5u5spA2and6Xv6Zlp1YBVmtTnXiVeAT7GissqsiOiSFIbItLyHJiWw25q6+EhXd4fDI
7xETXs8FMV2oaa4QYyi6opm1i2opXukjyDP1yKeRJ+1f72C6Rie6sJGEJbJu4EoXKuF7CP/EwtKk
yXkKC54fmYyu7Olyf47DCnwpFMnqvu5RkukA8y1qLKxlCtds8nvFhxE315WSi6aJ61LkY5CGp0KU
p+ymtO1BzDR2CpSzGfQeVuiS9CX1tWmdEmNI592jok4/4qG/dsw183qIQNcKCgz0zHthfxFyt9uB
ZzGqK6d/pcD1Z2FnzPe98+HTQ36/HZ3xl2qswjUvo7AtXIbMt47z1ZjSRc0J4Hgtf7keOyUONF8g
QGnJIjZU8Ny6mK2Mq+otZSyfc/YVLpbc4BtQJ6XEYqTqaDOIRvhxHIahtYfxUHN+niPDE7V+wHA4
F9sBML4ndrK/17B0KwyHaqCQ9m4zy+Ruf3BTAlO39rEDOOpyNXOHk+eD0jp+X+QxU9ASydDfPGNj
axYfqc3pooTtfDQonRpWJIiCou3ulYATejcLFV8hj/VSdgEHYOTU/skEBLWcmr9rggzw3mUPaIAJ
GQdyZsSN+Wsmm9AAVBUL8jQMFK3IyM7+pIPC8szdI6MlLSWArSyQayEati80DFFPg9h30IrT7Bsz
GZsS40oAWmherz6P8/JE5AzSQEDvhixdbF0dsgbeG9taWmjiOZj4bQfKcQrkfYKvZ4ukmy/bU1Su
xniWgOmkJ3XLXJa359JUoWJ8kPaivjYVg+UmE1VQGrWlnk2oXZibB8Y6NTwB3bfXU6BvQ1sVLSUA
Ds35mH3f5MsC5QPKkhONGeMlJJ0ldJDT9uZFG2BcQ3rBJz5BjklIMVM71WJjHIj6b9cC4zXRLUcf
uSMCqiYEyq+irebcwnUJFbtJ3EX3KTkgANZrSTPb5K7ONusoEvoLB6naKdZhFPZNBAZzuvQ+RdnV
AcFOjrfXnU1jcp8qmbR54YFC1dYi1/ibYuoADvYANmgQ0MUzTNQrombC9PNzro+DCfoF9BQFAHCU
Jaamu9yKe6JrSfYnokH9+McfUXS37ibOP/G98GvluTiYWRbfiZOCYXoOFuNsmGwzc+3LZi2oPs4n
S9s3UPhmOZdl6y6svljFvCPEZoMzGMv7viGoJN5J/UK759yLo55vtKH942Rr1k3TpaXDIgl8YB2l
p8pDHJqBEnNodxF2L7IYQIFt37nAYQG2sDW5KZcKS0kRjVbXxWJTK3eToSTFcw9eBAyowP2FSInM
zzUl4FuhEkHaO3m1AyevJiQcGi+UKux86KlU+T2FyOhcpC1pB+bRcsukFiAeMrtfDuSNSzaLLBAD
V8xJb+FXk3A5vBV0rYAjSZ6s1xrzRhmDWqdovlztMVSgjSlocdD7TUHhgwDxP7rA4JW9bD9agHk7
fLhJ1T6sRdZbQwegaTIy+vrtJGoZFbpZeyKhUwaVVuv1zF4MXt7X2jgVYP4labx4ZenH2KqYEoCn
XG8uircE5wf8IliRgFbjZ9TX14oAQofwVk38Qj4kwQxx6lbNlzhvx9lfVpF7IiIYc2PdXqCDQ+yb
l3jC62pFwVkY5oW5Ndhd1ApeoTxPn0DYEippExZd388r2V/tBed/1K+L+j793TeTwwOASvOCoTgq
Rc5T4bYalfB5yrXnMxV5YdiYDa0CNnLoAafFmKkrzWB7x+kSSXNZACMLbH399kbvAdb9OMY6TNGT
7tuduKv4dfVcVNEtxahrNWtRlgoZ+EdWkD82W8cyrwSz4u5CX3QoVduy71KVR3VICTE/VsgVWwD/
jHwRyT7Gz9EgPoUumyyM6fgRhfpCSyXojtheTccDvh3Qx/OT5oniFFrIyj5n2SSn0N5NJqX8V5EB
z/qOqWMoQB5MoItAOWwxB4ugxhlLG575xp5c72wa4o3e8qlO8jTO1SyfoVhT60bXtK7Sp4niTDjZ
SdC0OHDWoYJOjwCGMiwZ1n9F5/lxfjTPNLYfaWCcXRGfQ9MC/oQwL/5fVqN2ydlSU5kmsIMnIkqq
5qdZKaxJl6JLrNPlQjDRYa2NKCBiJXPGbPQ1anFak76XVL0pT0eRIev8b2yKLeR0pjO0YumUXkr6
JtFpnYK/G0A7abMuVsh6+4x49s4iaPT/F1vKXBqV7EVZv5eZAcmmH+gy0FBNiWJOrfuMIUfXGVLU
M3zWTNm2nuls1qZIq5RjZiT+vOJqVSErvW9Jbih19MFkVD1OWPMqjPW5KDICxMwMXXxfU54UZPzP
30E0qt8BJ9GJVGTfkYjdSVMiWPGz+YCh3Dq3hlTzqU6/y1iAS99191fLXuzu/11PvtG/DrOvtnCO
mG0W345XeVJyXFg4xVN6qkhkvbZzO7kJWWZlpD18C3/aqsuWHNS0ywuINhKkxhz7NINC6ExgKnX9
c+9i9BjEbxORK1aUH32dzQTBGJXXEWKQYdcQ7RsC1hqyLXbZNdXKEwwnZZHzHrMnyAb3VMGzGROy
sTYPJBECYaBcmIw7OonbkEEgH3uEnzi7DBpAm/0OsdgtRkCP57XqwmzYBM5vzAWZBDNyC5kc1y35
klUWSu/7kT3ZiS94RqyyUBZ6Y+22/WS5W4qIb92gG62RQxeudaZDP4kJCxCBTWEEmoV3+ygbuJJl
lxGrR+9QAYfIsizi9Z/v95QdDdlXng7gr2/zi4VMGA9Sa09ysFzSY8we3w2dssH5v53WdtAzL17c
q451Ei5FpRHXsMYP0u1ZKMoAMcw5i9jy/KRG4hoh//QPksxYKn4iDXuGauw1jTCmAeXv/NLnY/o6
V6q5tMmXHD2SrFBuBCmDTKkrg23NDpQ8TEo3bdBSQSX1dpRHYKKZn6HOkc8MW+HQrcaHIX5FV1q7
ZuZPYjHhOrtb4MqYh9iWeDiPqOmup/bU0MHLZ5m8utpAgM+VvcFs/IaBnPkdOjUPKB55BRASBXMy
j5TThpptW1/hH0A39nkEnIgFOeTT07Q06HCdhHgrZKAQucdFzSoUvZhw4NIgoCnJ9sGRG4kwVbUz
9IxXiql0gzbmPQTRvLm5+L+6yafJm/x/3jQHQJV38KLYVNWpePaFrTDgroC4e/CMyN0PBBeN0xci
YJMBd305YekZyRGNH9faI9pHMe5FRUFnrI5A1U/ceikW+CByGswq5WLMPMWzwPY0aZVD9agQoVOT
kcU1mhBhY6nySC3DKLCTuzQ/9SWWkKl6Bt5DJr6AdMTTVNrJaSYDrHxmmeSx5684CsahzdJOKLS9
GveAg0LYIqOz3BsR/c+BtEzQ5BYrDDI70lpqmWEbE/LLgzLiwlLTUN7g1IJM0Dv9o+jFDELwRFmU
lkwrhHdMTaBbe1yLbBDNE/ThBuaJO0T44n9Y7oIkRD5E9xgjMjbS2qSddn/zI2p/cQrTEKiNB35e
1wbUdVf7dGqFpgZ7Jbh4LQDFNZEo7oBDyq3hAWZ6YS+3rIIhOybz4jy6F4GPUkiKLTQJPZtaBcek
OWjnmXG9UeVwPNKqaac3OFGL/xki+s/7zjiAPPTuAol8PUic6+KN2BHoWFRKSF8kVaB6PeX0E8Wl
X8nMXv/GltWXn+QJtXy/fZ5SDWpKZSyEbkOIa/DAjz4ADNqL97zawmh7iaNdvFAfno1mxFzCp7Wg
duc1hi4f7KpE3c19cSLHX5zLEIgD/w8kvL25SA3TIusC5nL8BPKtZqtj8UY1F0cfD2GKPmIi0rqJ
RGcejokzeyoFE344j63xIR7hoo5e4uwtJErLe/BUCC7bZjCsqwkyW6aVudz0GKnGvxQu43lPnZUy
ANt/fwjWHpDkwGmjbT0FJJySvHGfylqcbXejq/jZe6ST3kVb13JdHJHAoivw6v1nMKUyDldXeUQW
FKFgKB27gj0WLU9G9fVvFmaKLpSz/sce8u2s8w6bwGwKbv3tKHmAYixPNNCn8TbnzH7jiVA5v+35
b5nJvwiCbWJFtUhxVaojXRzqxd6SABMgfqlpz3uAwymxjGpaE/+sHIYlwaXHdJ5qEV297QhVrAiJ
WTYeb0SpT+3TLBalzQryenG04+a8s7BF340W2QoKRvgIOEbEuHHrYviw7Kg3znzTICFeh7fpr29W
gpRHV8Hx3WwXdP562m1YHroYGB4nVpBRB3R0+p25mePZ8/5TnF2N6xGzQdMIoU6pPzNSQzmaQkxH
HVyBw/jXfvx72ia2jwPFVbPNR6T8HpDoKHWr2f/L5yvf3fFNzTx4Ep7QVDWW0vDPt6m/ooNy4JOf
TqXfUcnXP4n5F/XPgNA6DDjwZDiKqcD6suRVO0QwKCBJAL/MdT4ZYsQFXEyX4YuVlz27TKo2211q
F1HDXZNGL/Nc4jbaNuRMiEsdYeTI+5MdfVZD0zgFjrWmQhkbV3PQi2z0Arb651zvt8SVfvIDrr5N
qoxkxgxw9l6N1Ss6vLmXiBmwpdeExlCBChX/LS9QlNdyG3YjQi73Wz4YqmNkIZVIuJjWW/HCqOce
kvHoPUZEbS6IakfO416Q7nauUVfJU4jRYwgC+yPC2IjpeHkNiCBKTWvUKNvIRT63j2ediQB0Dm+A
ShijoO65VVut3t1nkz5p43CzJ04S6kpYtBm1L56O44Lo4JIyRxxzcakJsPONkCGMHxWKvLtmU/hq
/I2rF7tpqdSMbQNU1DpjfaJWgoIfiCc+qCvHMGolF8yeFXo8EG+ihh0BOOmSj+Z0/uY/BXgD/NhJ
ifD+M5jUqV77HqyABQjQ0SmoY0ZOJBg5mLuRSD76FvkxM81grpUTLEVqSlED7JF53Ze6ZoglpFr8
wwb2dBfnF6uqxa+y2Aur7yq0fWGevT3P/mHBD5ElTpign07XGzTIGxzPq4bFZeZrS8sI5XtJnlHH
TdJRUw/NTgagrS/24lYKvLOx8TCx8DiDia1MykhCtY1Wcnz/8mlGInUPUil2qP3kS2oE9Wz1TLra
CG1C2JImAxLOQd6L0mBS838qfLbtRPbaRwEryZiudrQUHuwWC2ipwAyURkATFH5Hd4u8uTlRIeqP
Z61+mi8Kh84scfD7EdGRBrSI50biPGCY13xYieUul9eDo7GO3GiLZAadWuzz3x9fHPXwmh9ZzLya
NveBuO6Hv8h02u6GqQE1EhbmsF/eBNnZR5Jnbl/7S8KbLVWp/OS5yokj7884p+8yO3rX7Rfm+6sW
wQ/VET5Y1szuiwL7jSl3JQ+0o6Ucruz8JEtbV4J5D8nr8+9Q7TCAXpfuGU7I+Qq7HBDaH47ed5vV
8dMCbRJGJ9HGK0tBf6iFRGPJZPo47F41mPICwBrDS3iHoGAbYVOEp7TVmy6LPcd2MNr4FphutS1F
MrGdOJw83aMgxKBOtIeU5CLDtL7GYwJqt4P0i0RfTrqHgCxtINDZhLayNvwgr8wR5QBd+ZDUB3Ua
KCcLlBmlURl1eXCmFO9apc8aUP0l1hZBW8+90o8zJ9cYNanNHdsA/ItaCnrsM3pk4pjywKGctVEn
KBEyuLziLZUSpnHl0jGTCcWCdJZHN8qxGUhmdkIBQzHieW5pet4ix0aYa+Q6K6KM4asbWWwxIVYI
vo2PdCXv0bDqEYSH91I6+cSxDsK8BvQCoNaVD/jiqLiiYnXF09Dp5AhZlYp9/fY8Qt/+22EZNIgv
BsWyghsxrEAeHrFXIguUyIeExV65Z7CoVNsOA4EIO9q80t3yryyezoAhlaF/0ozeWHKvPBNbekgq
wnPuP5OazIChB7GSjgJJ/jhZblTlO60nqGgC0PsUvDpNvWnStW9DfwPPxJP657aLYE5Ig/YhqyUa
bWbiz+aEXfMlou+3p/JS9IZu5I64U83FPHiIbEAE1Sr7oNZUCcHqRuHBZUgVhAP2ZUUt/ydMciNA
D9zTZzS2zzceioNovEi2hhiTvJLpDyFKEzLgMZi+m8y22rxG/64DF3X+YPI0sQ9VMjiJuQJmSmz3
KDYQy5HalHkaUyRV+vSYdR4y6akq+kzrH5Off1uGWRr9VhrgaPdG13d2ThWaRJS2BfFyMfhmMPBQ
lOdnm7zYVBgKLQigVBHdukCFDswl3NggO9MQrp1b0E0MGxfxzMl/YKEv233UXfgpxSSAvu8j9ckJ
hmcnpWZ/IHyn9rg1UNyn06Sx8WiaR5KDE1hihVeTRa4VKHVg6wo2pk/gXz5xxoBc7gTdh2qTZ1H8
zk9gBxI32hrLlcO1+SAj+a5BkBWZ3OBdEcJbowM1zKBqS3D/votmQGgj3hFj+jSSBWPQ8hUjejbB
Cl+2w4fYkBsA64iDvathPq30OjJyPD228pw0GOpJb/a/AOpEJQ9897Y1I/oEMA5Zm6hQwEW3kLQs
5q05nijHqZ0k1atCUriy6FNZ049P/2vpRzcKaSYVsLoQIhmSgk2ljHvTAQfBX4VQsQUJ2p/n/7Ha
Ei545TqErsWK7mhu34nOvua2Rypx1SjC4kiGqCS2Nm36Su627N+qvAt7URomULm0f0LozlMDF2xV
SqcUUQJGZPH2X75Y3+KzuJmkXLLT+zQO0LZWyk6/lO1yvRNSuDFXe6srYQopF5Ez4P++a87Y/ljj
m4WUGcVrLFctnO4Ib9VcuHNJ8VBK8PjI0EcjNi1hNORDt9FNdg/TC9LFXJHdn32woDsreKOJrX6i
ypXwNxUc+OU9RGoGnOQZvfATil6M4hd4AIVSLmj80bWAH8BF+aL4k7jnd6FsneXfbIu2+ASnVkag
tZ/rCFCT8ziqj7/nVIZn5bc+3dln8CTiDfxxAzM07RrbkXSBuCBwRvwFvSjEv2zrMn32JqudrnHz
w/fPCT796eRVVRvf5xVNHzlyNDj72R9K3i+xKF19nZa4HsKReC4p1cXU9loY7+CnzapjxCLPKs5/
evi6TmbrmxlNEiVGmhqoyzHjD9Y04723C4EuEkzbP4ljADRgGrgyqvUDY0TUFajBb/5RjKhO/4tm
tmL+PR3BkM6hlGsYYmLoSHl8+3DbTnTN0nhBSFjS0LCX3onOof7E8oIAxKmZ8TWszTrQ1caLYyDG
/TIfKjPw7qAXfD/znM/R4Q0diEhOy4nK+hUwB1iJHAMj3b4b/zPUM9Ec7IRPQMysdwO+fVvaHJkJ
98WJEuAGKzsYpZ4ER0CIFYsEYESxPEiubeompcd4Oj1m0tgDyxHvXJCUmCf3P0V9gb6+fEwrg1/O
mFXWxEM9wz8jomCdso2MYmaazt59+9/QkOrwTwfvCkK6bzqJZqT9mID1cLAnOTUTbw/IcHPangPD
fv0AIURVpJlaPzsUE8tznulxTWcKaxkSFZqnEbb/WzgPvfUKZ5MHK70EJZqAQENelevTFnctFdYm
NqfKK8MksIGDzYdi/5gSXlbRoDq02W8I5f5BAw4OEis18HPgd49OUuAaffI6+JqyatIlzCXC4Jjk
zulsElA8PJn2/HcPzaw2VWYtP2AogFpEO8YrFtFAPpQsqKXoTlKwQdfKvlAj2nKtW7gdIRuUuLaq
441wHgQ/Cm5WiaCUfOPRQuo0d4srK33nyLmNidcw3TpbNn5ROWWbE5SeEssXAX6kfefKtdt8wsZ3
LKD22fmIQRTyGa5iJ5G9xz36SBxPEEe3hqrLHyNRrq0NfMb73uqKjxXYQOZytRkzSSqmycSX50NY
KM9wNyUHkjLFdY4Cjkqu9HpENf6as/uNySd6p0lYq8EA5NlHHXsVBEjAFFNrVcA+JKloZxI83edB
I2632RJp1/rnBs7hGHqHKkIMaS8Cs4W/vs/Ttz5RIqUiIdv1mpZJ6421TrLSntYby3dp+RS8k1tI
ewIXOi8hHOfybzF6o6pF0ihIKVuqzB/xEP5aK+tabiiK5ucW43MeKok/d00R+4kYCJVBTMZc74Qy
JRCpjRSlr/77v29EQXkBzHBfC/RVr1w1FPiuEHfqNig2oZge1CWpGf6x8OFVfnDDMjpVO6MLPT/y
n2TcmQgkP6CA7oyUY2zv2MLyITcDN1Ko2/MjnYUniW/fnWi+ST3ZPPzBm0i1GzZv6RO0buQ3bUmg
g5WW/EpGCVCpLJGFyGFQqxLQuC241mvsNnQFkroifAGrfdc21VkaHLS1f7+iTmOXcMLD1seQqOEY
yTgw3uP2i6X5QuVHc3CRbkQehnEwrwyi92k8bFVgMi1mt/9oOros2OFH9kyOihxKeMnvWTqTSJNr
uwKaH/UmAw9mGMBxoLg8xRiOyi9wQi6+5B+en6yTVWShN2TWpsumz4QNzJLqSHS0O7I4K1R3hdf4
p/99YNY3ihix3AiAo6osAkp9LjcsMXqdd6034qm5UmztpRLwxzbr5I1nRQJY3ZzfJ+GVC9+cF64q
K2uzr/Bl4kkHzjtTIgkiROqh3bGxcSOViDONt+ehFyS6pHDwZvEzcHtyhbUC25HVhJ19UV275gKa
qdrRIH34PtrHXWx1PFb7kdnd02C5xX5Lcg5QbVHri/M8WreMmenomUVIUX2J/rcizP9uVMUn+oNN
WuoC2FkL+KMEPb88mDL2wCGhrXf+U+guZcGnZsBQS6+bp26GJTuIjWU6r+5mUqxUEN0NalTVrp8b
ZrMZ3eqle7VA5sWilMlkKftLmlFHroaFljVzLpKuC16w5C2P175oYpf1/mjRfsYDL+sQuBeaFWX7
JUhJRU39wF1tk3c6o1cEk14yowXNIGDlPuVbCMXXND+B5fJVet1PFPPctlQzN9ur9wA7wul2avHV
Pl4lTXprB6UrS/Z6+WUuS3HauL4uqkVkZnfyUIOURaKqe9BB6L+GV9K/QbZojq1LE6wOwqshbnOy
3EWi9aMQxgywKnqyfRJKlx3f0pLRNDM+DyUAAVvF4Qr9Yk3X+bwtqLmN8Nspv2TN0FEGhzJ6ABOT
62uLHqGHKW+L55Be5PAp8G4C8gacczm3QHnqk+srQrtqPnsNGkedJRrNtc4H4rwO+pIa/x0qhjgt
gyjSVs1ViHtrdYwt3QQGcOTLCThHc24yxLgCSl3oTCW62kS+rWIm7EsELTLLupLlVGhLrcTK9ly7
UDA12dHiGBSuEEXp+PjQhFbBAY7xYU1ppr0aqRbDsFW2wHU8DqLj1khz6oZnHc3nizzkrdvUQVCm
j6V5iSgsiBX21shqNpS1W6KaBQ5w5xrjeh+ZyqlifHqodAZ6EohnOiKr1vLvWkJNJGBlbODsHs0H
faT4Up3tzvVC5RVUvKjT3bnsjZhDuVStkdJ2kZEdKfbX5/TBc8Utgha2UPYv+RlrBgc+4+/90Q3i
Buvdp7KmRiQ8ME/8x9pJhiz2CSpheFiGYxMEXs+ea1DchjtsV2fDfZCxKQPXzRs/omYeu+MnVvyc
2vPUzWlOnIDaoAtaW5ukoUbFIyDPrv2zdpsuBnsf6xD/MFsn7qAIoxp9fT05esaR6rOwPqX26+SI
XyX8Tszz+pOjf0vmpu7YnALYN9GHrhQ/lSodO8OuYg3YRQVfLh8XZbFXaHO7ZejeBaJV4p+EobcZ
fkCPYWNB+KaTaHpecqhTSTxkYSCSu9jKSd2/m/l3q3r+cR3fEd7w55Keljp5npVkSrkVMOf/88K4
wkFbfqSSkhOgYsUds3SFSI1MJfn5PLPRZpGXLiPgiGi95tAuqlhAWMVW+i82nyMBTSZZnJ8Y9rrT
1N9jdIKtnNfh/CRhbNtGm9fPIYT5migKmk1CWkZ66JWRFK60Jlt9sAfQtJ1ssLjPSiu3y60tAjDt
hodx+qFXf2PMAu+3geYsOmXbIC6vCjwgutsesaNqyaf3Lilr5wPmAC3riqKhZFTLlgXzShCJ7Pqx
p5mW4fD1Xp4qbdStfhKZyAHPgkku1U4qymYyofjsX/Q7C8wmO93P/YTt2CbIG/tPA8GXedNej+p8
WuH/qOJHmZV3rIr7S7vftWCH/Svqiw/wpdffr7gr2khhgMMAgWrbj6wBXTBbIIUszv1TDI0z0HeZ
+jBZcOXl+LHg8xxz4w4s3xVz5dDqtbp4aZhXStBSA5EnLuY9LqKyiEh1OvNl8BtFkrri7BMeJuNx
T9BZSy5fswjMsaPxapBJQnZ5cp+h9snCthO6J6je+ajXXut3VYbiGL1disHU4ELs8e+CJdieR1rH
68tvQBMDpSy0ivaKXf4GWa2zvzWlOyOnPWMTBeqf3fQkqhnDleBN33xlDd4+rptLFzRneod0tXKn
sgo8IWSKW0jJac1fgjFXpwnZLARcj4qXcf6avwMBXgw3sPc+mP7cPofxfoZjYMPNzj19xNGcOQme
cROnMj0eRuuClZhtL56nYMqeImQ/7NbuLV3dDGAIBK3e/EKm99d+vGBnCzyMvdkEN5KaCVMutnUI
jly+ixiqKfOaT+sZHd0AOKIHoRHe9HQWbL84dTUNoe5mysdmRCdhAR2Ge/CyLBueGXLfMSdkEdqx
UMXvrbUGWrUVyfP58a6A6pf+PA9HxAkflo990jLBMass43Q5XokDXd8DoaXk1EHxDT1J22oe4kgC
TPDxPxTuVI5gs+2SbR6q7jIM8wJwOe5T+nsX7LQ9rsGNN7z/KVtda397VkwJeEl+xJiASSkMXDk+
3h3nO9DiciChTFbepEQqhgjlBHBdocJwkFhHmm+TMUj5rZj1yK/fJs8s6OBoC1vnIHr6/SvGSynt
0Aw59SGNdBnxqa5h5S56AgR8muOH9ehHaFKIyJcWzNW4nqAazS910nmJRPTOGMqOxjG7VlC5l6q7
UQ5mrCjCHOwwqShgsqXMSxTTy00zIaAGuiP+WOHXhlVPVbDc1dCoz1sFk5Ve+9XJU7feOSGkF698
tm577fvBfwDNI1Kmey97SqhnrBeZT85lFrQALmOR2lcye1A3ztTAHT73KcCA1mkWHsqz09FhHdL9
TnmYSWflxzw12AHjC7xrbfOiqezSO5epIQU+0CiTVDBU1cwAP/pwjbXk8+NQCEG3PAkotjrBVipi
eWkMLmblCtJmiNeXjtwQwqW23ZnSN9AJWVBvfC8g+hcz+pg9JLUHeSTTnnEIZm+hJ4Cc0/aq92WN
NTpSq+pNZsMEbzzstkhun1ysajMkcVy/m/w751cYNdorbWKSEOwf8IKoeSHrbXS5HrE23PQt9ueS
YSUC+7wfG6Poc4wLqJlwbI2tSRW4Cjd9AG4j/GShi0aM+Rbbd3/cSx/GqQKlQzZN69XFC2rQ6Jn3
kx/iuaPE/ZdC5C49m57q1KHPxV4mCP4LdFta5Qy2Hm9IBb2V6PixDYOCVOi2HesD5JcipZa2a/dc
D8pEfF9dcCTLbunZ3eDbU2FVfl9HWnkOV82v837ljMx01mGzq2K6Dh/9DvXgXLLwheHkgaDI+/on
NAPiK00qSP+C8+Aif1N2pEBQGu6EJXez96AawuOoU59msxgtYoBJg14qXdIXTPRBcaFNtb/yk3ar
Oocm6hetxos6HBexJ/Nb7Fb0KzWpuTC8vh+wO+NNvx6O/FAUH7BY9ctPThCtupAY+6kI1Ry7K9fq
YYLzI5Df132Dzb9CfMAI//djWWa6L23yWLLfcaRHWtz5eAy0NypzR4/HaScHjmilR7qEB8Xf09MB
kAdkBZlJ8epdKlGrGUoImAImfxv6UswrmWmRcy9WuhTuOKGohWa+iB6FyLWjrqJTSJVHBthXpOQ9
NWH9nCm3ubtRt2HNfrYMEHjl03XJ7WA7KL+4jtARBePHsY/l/gS7gJU0R84EHUjkScpU874ld48w
5LVPVSsT4UVLkdgywi+e7PL8DAl8k5/QUhqXNzFJQxTjvT11fivI1gkbP1YVxOPKASF6F9SKT5zB
xkG5tjI52hs2KueMs8wQQRXWGCsE85tMDAKT4lE11UAxpSIBmHix/s13/6Z4cDX05q8DFWY32ilC
gi8Ksn67gtySaikpxrKj6u6fWS1dkF8Q6TxG/nJnjijEXhVBV08grukFC4gBBBFGYxwquc13JgzB
TfYzdpCM8zyGkL7H2zRffnLGEywha5LrEKA4yG3i5dLxL9dVw63/652rAjS55a5AUydgZnEzykTv
rcJ5WpKwotQRIHmd1iOWHTzgEedbobI/YNM3yaL/18OfGYEWrJajsqV2SoAmS5O45oTc4BjEzQjI
m+d0WTTMl8jxHixdutwzeiOhVrIG6khzCqbFBZ6Sd+fyCpvS60SfX4eZGkNL3OQtIr5Dhzo0EL3g
tdLyHbnUSKmvqh+GI2z1il8UJIja/vX7fuzF7VeqKuHMHNeDurHzFs5z7F97avD2wy/7oQhKp0uJ
lQ7hGWMCceyNKiJ5ncErPydDE9vHSzGVeKR3m51XtqH4Ktc6csXmC5G5i05tyfptMuiNoAHpamU+
Pa0JZYzycm6lk9cd1oQNpc06FmLbbuCQ9XgQRjkY62kUln59ZmDy9WvW3NxSjRK5FOMn0JRuIUwX
j/fFGtUZ8m+VnXG4yfaOHT/X1RTWvGmYVq5527T1blqEXdc1KZlf6+Q1UcYXye73SNoT4hd+7x0S
dFGSIjB+OLZXFhn2H+l2gGjrf7lF/ZnDHi1RN8ufgR4DEGRwxraHYwysUEn68VmDxQw7k1aMxveU
dnl+tms9VyqKCjFex0ZMMcRRkXcvoHUoTyblTAKPcJsNZ+R1oVHvFzq/6HNcZOieCIJYYtaUZ23+
tKrJijnrzLCl5CPOAPv7pAN/10M8nImcnxKSS+0hOVG6yYznDsXEunn6Reo87jzkewf39KPupNSJ
2QC4xqVlNjTdQNyJloMQrIhPC9bfUBZc+WStpU7nOp+ltytWgyhbyPgumkz+bHUvR3O8+AECWg0h
fPMUts239o48y0+zNb6xx7Rl4HI5iTbUQ9Zwu//Gxs5YpZhVHEshIBMmk+OKXMJTeE9Ue2kpSE6n
p7KkuGhTrfDaOo1/mZUGTdIs+YSmwQxJD0Fi1Z0eX3KmHfIdLAlFmNOuE/mSuDTXyY0q0PattN3E
oXXqjDlAaWjGXZ4FYkVpnl525AckypsfYhVTL0oLB33T4kt2YkbuTr7np4tk/JOJWu4IEk46A8Hq
1gX/rDRHt91MrwPkN5xaILbgjfaEiYexx4d4MbNUgl9IpH+F+OOWCg69v5NFvfxDa9UICVY0dIXK
/0os27CvjApvshlap/aCF40q913d6cJo8ym2tgh1UMp6ggb4cB6Kwz+diibCeotwf6d8QBJEZiUD
dhcCE7VtQ+/WzxLZz5o3/NiPB1f5umefM4QOp8SmblXyF53aYJphJN+Q2iWAGrDntj/KnyoufvRC
gquAMtXG40NYPqbyqb9LEK1oloZRlolpHnXXu7OZ6grJADPttfLMxWJQzHrboczz4kwTzecFhk+u
TcUmWd3qgCpnlh0cRowoTNmUvt2gEzWHR8EpcRl1+8crXQwag34th0wI4HfHF8TNtcEUiVnWRmAl
4/rxD+/mk1h4LNs7/YMzCtEt4gGhEvNK/AxcVmTzeBKopxJGYsmNSlo7u1RfKKXw9mwNaTLChCD/
BVZKlfOtz8VDIMha6bfTrfajqb6734asehWOJY8dRJafiE77J+VgEe7Si417Y+mjUtrotS0n42wd
welvNokpUPxnAWvuvJgR8BoqUrtLDaRHDuOHCMDyzjTNYofXRGDjiKp1YaRiBasHEGE7Krsm94SK
TUtHnxPjd9twd58p6eU9Ep5dGZLMq1krfEBM/HPZSFnfDLUFOixUJa0mvdJV1BJAf5fZtr1+qnXK
zJQDtQ+MIa5rPLed98DOPBuGvC0KaVN4HvxwEFH/hRoXxGXzKOHEiXKaDBbjjdPkXkoCqL2SD1ih
6s2GtCBYr3RDN6Kh+PLncrjgZo3/pt2A0klPDpVad5ASwUCyghNNzuMUnwRNZLmMRUd1OSDJPnBh
tZShMO0lHqcnt4kV5Bi7ZBHHD1hMbUbJSB06zOcOgnFR6HGTLjNMF4dULSGZUatZUo14bMbFQgq5
wpSXtBDcQLkWIJ7v4sUkl6qkWUpVrJB+gfEIACDH6GHcFVKKE6guUnkrmUZ2jj2k1ynzpPuiHQpf
oUnkkyFo/PfAWrCUu4KWwoEVXETQKYMCFgsQz5ZkncU6uK/6Yfcbl7uXfMdSQQ8uwfMJgX8sUvw9
ZNVetDWz1ZwYKjgf5EzWX1LTRbI7Xq1IEBGBKI7+QY/qM1/kDz1/ewCWxRybQc8z/0xdhynXI7sa
qWyxfW+qy22n2dfSwTwAN1/v+T28m01D+JnXP1YS1vIypcShdFUEhCaEmjBJpGjDQh0r6Qb+/n16
xppUUIbQFyTNBMAmcu1VPnunxTqwZ3Sqzhxqh6mxSCB3EwIqu+RuaKHgp9QsREyeMeJkwMwwnlaa
d+yIaFNXbSL1aRt4VwsZ/6Cs2Czz9tBYNnJAqz3KbHhgzdWmV4LPSyapLdRtPaaKW9ccHD1RBPMv
QpNnF3Ku/33L/MmPatp4IUsmbgb1k1XqUYmJPu8AURKDffvF4mSu8b3hXWiItKWt0PkHrgYJJ82Q
ym2ZUk31uM6OZR7CwTxCkr+pmgJwnFgKpKSUwEl9e88VIqfdxTRZ1M1BuieixiL23tZGFOazcZyy
EZhg7XLH/sAlr/IHZwHRW3hj1NMrgnrBqWRVtpBFBRT1B4XgJxQuE1P8MPS5UXDBIJot3sZnt4V2
IXhHzDIdNUTzDnXphHm4nKUd70sTSOjE8f5uiuJo3tQkXC4GyRkrMCBimuL8SiJrnTRs4ZX/7OYK
l17S6JGRInDJ40lqIdTSp83faFoP7xrrufijeSoEK4huW//JhqiM/ZGrqVpe0Ba/KgKENazmbZ6O
tHpddyLGl9upjSqHnBv9htX7npu6JH5JjBIh7umpHzrjScm25dbJwYp7eVuBjP4PfVvkS0HBmOOs
Aj6jv55He/luTYIRV6uzO7WtnM5sKplyMprh7ip7ZoMnEfTVIFvX1NCqgD7NQ4lvsz+0an3KrAK5
CJlu+Wzmk6YoPwIZCnPSfRuaC526+6rtlWDFbXSN/0dbfsed+WFJr62sEUnkoPsAH9Y2Swp81YHE
LEdJVs/uo9oqCtVhJ6+HjpYqV+7nk9y1pm8EccyniuHKw57w+0gjR5gZpkFPfucOg7EwOB1IFhrx
DjuQQoDiVgMRODMqfEm1wINfJLvgN+SykHqzeZDSKFadpmNWq2IS/J7+AGI3ehouWSqS8bmdOeOr
97WU4ibbp+8FW9p5KEOMSc49FjgsEUo6vn1S+s04JGi1ggJbbq1dRbhfLrVueqsGjbZQDwIcy1DV
jMP7/EDyT98zkzpogwtCTNUXw4VzmMjy52l45vfbBAhFzWsx7Vrn966D1zAzceN3zbepVJWEGbHC
mJ9n8HacTfRJflFNIorcC5yl0g3x3Pyj22i3ApMnCbqDDXZedoobLkdEsm2YzmtdQaPrcB+daNDu
vlMc5CQMRixV/RBwHdHniTiQAkbvnXtMyMhOQ8r2eJMjH5FYFIEuHhp6/Ozjj9XpN7hgmILBdOYA
vFDgINd6yH1fbDZYEuJv+DdikrteTRT4CfuEZzmopbEbdRELi9Sha0pTgQhGsu9MA9BMV1cnMyEm
Ne9+w6bUzQbZsUVPOPjNky5eQizXpwBUbxf3bhX17m9c9d1PZYrAp1Pobi8bJdBpncpRd8O11Wis
Dlj2X3vzdjnjDyPyz9VrrT9C9vy6vHnoK/DipqQ4hqLBjOz9HmHhHSfOJV8JPsCkVtxNIXqAfT6f
rxAph9xU92ytOPecizTV/JQexf5eaXqWt0UtxVuzcHlejWmVw+84YQ/GqHCLUwzVAUpYmwJo5p94
WncuDYaErMh3FJ8wDl5qfc6TJXwgCMIHHn/+fBQL/qVFl9zAxyfwXZgJYgsxRekciLxzyzCrlct9
GzwU7z2M5bLh6YFFnFLhmo3upmMwGo3dJzJ7NnZd3zU2XrWpmkKcnEaht3E7EQLvEcJxA0DUgI2+
co54fUAe2/brtvIVKGiFlKrRPVhU7A5fE3L5osFHHBUYLdwM4HF7EGqLkvW2UbnBnY1JZtc67EAb
ferDgjbpPqhT8mz3mPJ9kWcovUeDU9ryKm52QyJGBcaT0o0AmMWiH6lrT83OQYVRL5drapmD/Z94
2YaSE4PZVfNqSKLezbY5rZYpVEFMNTVq5rSdcdV9lPw+ii+9CYcVPkBbaEiRfOSUQzCrgEZgszze
aJZ7m/zeGAlSRq1oIH9E5INKnsvs8ZUmvEe+Fw219cBwLAGzRz3sij6ggUSX3Xv+gC/hzAvc7ZzY
fY3HMmpxGjk6vfjvQ9rUgyKbIeKHAC/R7X/x6FhVSFVEeJBbLM/p8/VwxuqVAl1VgLZPTqNOWhN/
lwtwoGdGlvTqDQvubiEB0uUOstMtJ0OUgmvACE0MGmLziAtB+IpfD9L0jDLUfVUjlLLW2L1LbBtT
tcvQUYdKrXp2UfhPbXqKMMmfXuapCBdBl4L9E8AGKwQ7C2si539lfHeNLTSU7HaEY2RRCCwQu3Db
+DwFy9pMb+U+vEswK7pizD0FiWtSJ63cIbzxBVKiYLz+HVgVw8KY4zt/aiZZC/JFOQd1Vw+/UHVK
208vqBMLOFBBXnZFDCqhejX/Yi8dRx+B7MlpW/FqKEFYvFSz04PjD7J/b4O9Zx3ww+tl6UpejhBx
GxrS2Aau1hnxw48eL9zapfC99tKC++NxVqV8Trz717Z7wNOVwo13Ej05z7LcJOTQILzOSgl7EiJk
+u9OUvnFlStl76dasYlsYuN1Gd3aqfBocA8LnZApcXp0Uz79x1grNCODdybAZs7mdKi7kGvWKp8o
IzKr8L41nGupk/7WXIyZ7E2Uup7WzqN+mE8YPKQ+r3N9CJWoWegMz5q9Q75Z9iheJXgKTJpxbZzA
TJ8AghpYb6WVeSEM2tL+dpxtEi5AvQjSbDRspWg9Llw5i3bAj6/mhzZmOFWVllHSfbDiCwNE/iNv
livfZMEsp077hgu9aKz9ZkQcIqBNzUN/FFKav3LsriWudKW6BUTJvqdgRA6QrgsuxLc3orCJqAcG
sTbMjXDhN4Jp/+O8QlD5i/D/I6pvOrAA/kvgnomODOt5+jckI17rfPkialhLlmPiZEmJKM3b0hE4
gkjZy/GCnx4ldRZa5UtxvaL3+JaFlu09lcpNDJhqH/DbfJMIn1YHu3oU2qS+NDRxRHdYzCIc2WiI
0BgkVHX1TbCflmoa3Q/CstCO2ac+8CCnE1pu0fAKApxcmUqT5Sj8Ho/JWBz+dGbqTzDYP5NXvfzm
94zS1bGJCsPF5cnFtvg6LGibH4Ugg35XsvswGlXz8Bb5PiH6mZVb/dABBhUskkzvgOU7k9dH4NGW
5PLQO85vtEgbZFFF5baSJpszmsqnRjA6zhazZutLDBI9yVvcTmjItwqboJRYl79hGHBW27hwQrRj
naURBhFs/GqLyRubdF2L9h0YiE5LEKggqRthmu3lyxWi+LjQyLt0OBWmTvZx3jt8P1h70YZ1x4er
RSHZNPPvXO7SRiDvKa7WIrTj4Hwl4qePA1kxq0qQxgdAYMC6/cemzi295Y0O9sxeXArWOM1P8Spx
nNrjBSF8WLvknRKEnnGM6/zRepNm8rSe/Sunx5z9FoAKD9AaG5bRFsmfSi8Nq2HD//NzscoTi7ss
jdk/ss2K9twfjwj8rwwRgnzxzrPf8vb59NLt4Fi6WcED24HppsompVLnnKLdRaOXGUhIJREKWPzQ
sG8sAOXVaSp86BIKIddNVoVJuR8OmYbTYfw9DBceRor6hP0QSa0RyMLL2PhBb0OflPyQxWtqDCtf
/z9KjDGhN6JlKkZYuTs2tdsgS3pX7m9DSu1TzWrq6Zf0uChgM3LcpYmHtWmyMIyBQaT2cZeznheO
s6fbadfufvnoPluISrRy+IEYxWpbZG5fUnX+yw+l1guwMzk3355pOuvF3s/YnzruT/xIMBy7AOiB
uv2LJZdpxQdnKgiJ9yagM/vlNFrVI60K2P7ADJp7iWaS1h9tjy+tfMlJUJzjwUkrI/8TpwzCwtfZ
V+3jdd7Zlyk9FJXxOn19MhjJydRMvdtFSNop8VKMVgX99t8toilR4WY+5VwQRFUDNuihKUF7gnvF
bileLJ6gOzlzIxgzUggFy+mXsZm4Yy6g10n4Qq6igTfHs/Yjg88fAjrOfDI0k2PjisKLCXPuq7xV
aAXLQo5DBEbz1iGOeT2zDro95B/zxbLltMzkv5ZrhZaNEp3kl9Ljx20eijPqib2XvLZpxehG1Z+M
yDtUzJVUOVasdHu7sisLnXPwrv1gBh9x7IPL98J0cvKdysQcX57uDHjdHkNbEcrGFQuA8uPFv4OM
zPbbkfSzTArUCsn/leriRX3Wgmf1Ut2o2OykUcmsUPL60aakqOqJppCcX9DqAlUcbHFaeMWk2KCn
TRzjpdxcUK/h4jP+y3cvN4djnaOFz6oXvNLD6M312vg3z8yp9FQjjmPV92tfk/xMSXBP0C6sOCgt
+dSkkQulWHzhieXVnftihrLhejyxnDatKJDTl0cKwtrRTiuZZiq0YqcZjyM/8L2LN72RSVUn8Dbk
ycK6OHhygAnfUeB0JPTstHAonkg0bl7gwcGTD7xX82wNzmo8NItxJz+npvq7QmSkuz5+9QXiriYG
hVXzHQI1IasWLmMxFUodWsddV2fOmUJy02K93icQdcAym6LIfaCr7KprVGt+2hiQv99ceHIJGDr1
KZ0yophZudAizM8ptBzuuGlzb8d8L8zI3h9WllWNWjmAmGiXXk9TVBoakBfdUfSEXFMmYxqoPjwr
T98S8lpLnMFN7a5LFZoM235twpEIqrUwrHefdFcymS+Uw0wHYRI0mOFHZGQAcB3A86+oBvvXMJ1U
P1gM3lECJJjQqiJbNb4XyCFyNpoV9dB/sXWH/n41ZFodDkFisZRLUqJag8CdiwY3wD3cuU6gAAmI
Ap4zEwm+SwsxdF6FTVzJA5VqjGS04L2DVyz0JytOMYYIOooxHf701x0Hg2Rhutv4NJZAitOw6+vh
xIFoJz3BJn22qVvFmxhNmTO/J1H+o0bgykae3/ZXH852mfXegolrFpvTLCo+3L9LQjcldXiGPAfT
UZuHDrXb/XZ6PDlu1hHzUcoaazfnz9HngUf7Rd+0b1uaowpgA4Z57GLsCPzwWE9Z1d9bSowIF9LB
VWeuYPKV5ECtSOdGomD5K+6CZiIAkw2RDy3mVs+LNGfu+cmlCmqBkUj6wWAtepJV7hY3rLJJ2sz8
WDzNzfK4/KLBZWr0W+d100ilKd4eOAgWUVoEPlrHzGcXMdnfkkwCzGxL43wSYC5+3q/UY+TM67H+
dPttXTXedco5PO55mf4TjQLyL1fxb6lX3LuQA4KW5kpIKs3bIJs4oV+tFuJmz0tsB9GR8mkBF3yN
nnY7Ep2vSeac36WdhlAjNAU6z7P89NWxkZvEn7oqiF+obmcc34paF1+mt9iWI5aES6vM2tkP9/ls
q7BATRJSAL2fxxcc87RN+z6Ka+vFksn/8Sy5qAHdxToL1klAu7u6rcPWargeZWh72194X4haZJB4
66qG6ixK2koD1zBFxZV9SXKr+cdSbvQTSH2KYwysEENxw9GAkMHfMuyPWRy3d/EoSCMuNKvDKxaA
/bswbLkg0og7adBLuY+QXVwuurT0Bl5v89QOJe0RPZZX+dA3fcLWotV0goIa9Fv2SujG+UrRnE6h
XaJlMtsz7oKBYZI3dyp2KjIWw1n33vDPGnFHIFNFQAw5rgHTjbt3aQMvh3bGw7xluUSUFb+WDd0H
mI6Bs19iDdzD9JfaQb5sJYE0cojkT18CJzDLwLbT7qmla123TvdftD8UG90JPi6hgZJqESV0yvpb
YveZGZvPBUZY3oE9i/owyO2zJkdwIoDyQXef1eMx5lVNKWSO7FGzQswZbpDpzhyJENBscFKpi3gn
ph/y10p/PzdmcE5veksuBUgeKi2wWboR6UA5ka4ow7QCU5Qf59fdN0myJnh3WI/INcSv9XMyBnQS
yKRDlqscbZCxLm8RM/HNyC4SbeaFKP/cOP66H6/yZBJYges+XKUMFr/qnC3LDvSktQIQc3NohLRP
HM9xjLwJrIqZ2OPSDfeTaoAXttnqmLM8pCiCi/AmAnOgXF0YDABBu97xJCsMmPkuEpWmMd/JvCt3
FKOMW8b5yCqTJUAp4E+FTAGxCwM4YYepdw4UBL0AewKcYQCPXnzuh8Sk0bShIqEcquo2zxvbBaCl
9adhWWHtB8uM8aCW7jZphsE3vFdGzH8V0xF4W8bHwfgnV0uFx7bYqrQOyqG+DBvwG77zY9eBeV3y
2UACyUPtPWAdrH9+RMEVeu7wJ2GGqCVslxGTd/iYu+xRVdTJwEzaHoXlaLvc6ydhS6yaN70Rbixc
cDWvLH295AjXR+hCCZbx7PRFt8xmWbEgRiwSaJsbzUCBMJ1DGBtfpeedLqvXUEQtTeN3UzyZKqNN
FY/S/HqO3PTrurut0OZrQgNL5R2HNOGzB+ThNQaDT/99utoVX+A1opYGgQ9iuKeN3FNI7VEvC+cA
f3V/wNpjjGxoJMnORlmZt1AQyNQPbyh+eME2+xnsurZNt9HgoFA4Cfi+nC7nashkWkd7OmhJeCGF
fiZmn3ekxEtGNCOZLzmrgeKdXKczKUzb7lNTqjELjzYLt/TEHBevK3oknG1cwX/lWLrGqJGetKEb
KuuYTSpebVC+Ec5OAC6ctHmFMUkEMr1CW8DCpMXFmhRYDfGbUQ06BNQ1Ao1f/Oevc3wszVlcYjsd
EpF9/F9PXWiH7LcW6A8e0QfWQOIMw2T51pvyGKeb2qEEf1/egpaFgeKAFDE1TZJUD1BFslaxvwqI
LIc7Z0Yos31rpEU2XUC2Yt860ctJ8RQsQmp9gED6GQNCxqqn3whLGgtP5aroeBlXmaPalwpv0QqG
q1uHHF+RbqlC1XlZpZmKSQJgpvVtBXIRVu39N7W8GXb8QlLKUSF2Ns0VdSB63FB2Hgs3qVnUbnP1
Xhno6Il24Y7QiiErwgjcvnFtc6VdgZVVg1hdDHp+1KQviJ3ChWIozd9h0Vy8Lc3j2E/pPcmw+qTl
7fk14Hyk2uNP+b1iZV1lcdVG+uAVI20VYNsjSeQQejq1mM8Off6CxEqcsWNme+SnjGt6KhDXhFbx
okFeleR1UCVfDG/OA4rG2Fw7QezpIIbqtalBRvuUx5kLM6s/NT2AQ/HEssZjy5aLd/6uTMOZGm73
0zRQs8faNF0sBtftVpN/tOynBsQAdWgj5ww92t58WTneneZ86cVIJoVK9dEBGSRl7nAfv2d/ONkC
YfmYomHZ0fnyjuaB8eQ3twXo+3f7FKA7vb4RgkVqaf3GM4EkcRmJpPhKPalj3As9xMQcZ5kZIUqu
Yh8VUvRkSV27DEw4eGpKu+m1zFTYBGQxowcIV9NdmGXDnzY3qRBWSvM3U968WpNLP/2SbcuoIl80
2/lsppTDEeTLrvTaKhEk09pJjs/Tab0NEqIljHNGPJQktXo4B2VBsqTQBiIS05RWif63tbaJyLqZ
an/amWWX5Gb2b51L/boQTBHeSaZ6oI/AmXyXZepZZCoJlFEThU+zEbloI/vGVzZlLnr1adNBl6FZ
ZHn7W16vxTyY1LuN0BIN6Fjbn0Z1QDBSGYUXgmIdmHXOnX68MAXNr+zZIrfsxyo2OIQ+/rEg4Nf9
2mn2VC5y7AHUrz7QVGWi+GDdXqNHqf8QYAjI0NawiCu8YT/hQLiAXUtPR7qsHiH7EansKjBObfuA
EaCLi+JqMSpVv908slCbWdxzcQfWAH7jK4iznR9q3ZSUTHLgfi82J6gaF1n7i0hBtiKulmJMJSGl
xZwaBVtOyZyyZzO34QyT3UxfTcuBoUiCYNswm8sk06TQoWSM/BPaHNnqGEezhy2QgarasCHJLfL1
jxEoNg6L1myMCZc8HQn57NAX5F13abCnKEQPkdu1mXY55ibvhcJV+2gsM+YrjBgs4JnnlE6jg1UT
2tYgD+TETcbBDe/Nlxyf111GggM4QRWWrGLeERiiLXL5TY/sGFD1p3F1VYdT+ejFAmDdTxPh1eSW
k9bZlzFXNMJQWUMnwQtI+YT/19jALUf9Tf6X6BbQdCQhqhPwE965X5G3A/BS2dImnDTmTfM2Q5am
M6Br9ei4cKIiDX18Ehnk7HZ2ZEHFNuprD3EMPDhHZfPwptE0yN7/pOwy0tKSTncdaxzW5AGMx5nE
A1NxJZs3HTiVi/X9eniGfkl8TfAEKTa7TS+08UfC8vUn5rbgpKqD0LlNvaHtnwOJdVQ9bIVuhgfg
gHFlRGCwUiipllD54i6t1cOjfvXD0uR1IBXerVK/fcGgtGKAjY6r+jknc7Z3cULwe1CHkfwaiKKm
bKAUgw7E+iHOKlNaC0ZJ6VLNfRaSEG+3vFxbIk45Q3TIjs6CyTKC84oRbNpCAHkxcc2pIh4GUjjQ
8bDCMcYLcE+vj+Rp/CuzzMaDqDLFqyz+v8RkZSlLx9wq8A2w9Mbo6/wmYsQjz+BYAb5SOVltDMcm
sx049wYtWw4AtZRA/pw24AlrgvOrHbn28sb1LEnQHaCaqFez9ZbfLqFFxxL22cTnyJ+aE91qRyXR
i76x6To3d5RxUsyGIHmDa/qbVOarCNQpBpN+HehK18AiSMqSz6yvKB9zKNJCUAPGM/wwBXThE4x1
zZ6mzZO+0S/MNEoN7MSPeiMKvOxOsF4fmCcnam45qirmvc0VPoQRN+vBGvpqNqkBs0X5JW8Zgmmf
7qBLFk43dHSOY3NxnI5PdHkt2R4N11b42C/mAWYIIWy7c9x4rXT9vv9uCaOrs7noxhlCAAXUVN0C
1mSQ0/T6iZXYFU3i3n7X3U6FMDYG3fWPifYj1hHk16YEbl4EqlHugVNeDfwCp3Cjr3j8hiyLiI00
1wRpq/QHMHKdxJsl9ngEdKlklkEqr5l7+vk2CpmqDfnYO6jqsKGCKp5oTe4NTw5Psk3eBsv/0cz/
Lx4B9qh+DXgCKqh/tmDpOl9KKDKSflU2OpoOhly4hktFcUG0HDqFGqIQDEl4M9jCIygp14dFQyFV
zp2ciI1yHq5SfGYoChpiZ1Xoux1fmSGTIEh+a74a1qSWCjLnXXCIid2BEirbzqug5ugHrOcxfg8E
BOHyKYsyiJo1LzjPo3eyQ+su0x3LdqZoM8YctqN4oataILeUUXChPcghueZ9cSkgR0f+getgLvcQ
+mq09btUPahYngjUiPrBdbB6TxrTCwqLZ+vYP8WeGbTyCsbE7EyXvFrEg8e9t99MpuptUakhVXBg
3e3Z6SdbFmRcqoy9MzXPUNiNaLpzre54CcB2QF7A4MMC5YuI9eSd2rlucHhE6xoboqfaILBxnBKV
GqwPU9D9oRzBq33Pc3k8Yq0+q0AlXd2iGFpYUNHOfqiOjgL4pI/WqgttjxE9gjF8uUQ+eC2dZpED
bhdmvtkXqGo9Fv6HcmvGed8VaYEV06WU+Tw8p7+DYiW+RSEu9Ptwr0JvoBpSPUAISaK62VaKV/gt
HZ16uF9zDZrZZyavuQWNyJSqjm9sOY+7iqdCxVCFArt5CQ82ILNu/uJDXrG5ZE1rfq7rCS75+EMx
Y+nl+AeBeTmuxPaXmYubmaJycEtX6jnIHPhvFkhBTV3LfmFlJSQN6xslUicpLsyMypBNHRoK5fTe
9yLmmNU9l6RpVnouDJJIZvVyO/9abn5PU0O1RCnVJAB00kGe856Dhn6zd+oIW1TZXkuFzeR+ZRDG
fn+6FAyuazSwGeebNbRAWNwqKwM2r67iyTBcMu24s7nEYFutzwimC8PRKZddT6HnhOu8zeoy/i+u
0Ve7gZcACajeSwQtvIVCvnZfU+DAKFB19KUDDRbgBPa3pxQZx5w7LHnYKzEynLCx7m3pMTDeGOQD
26v0nPKGWDZzI4n8LmO+1KZPzrfm8Z4sbUzn6T0DlTcchoIsbgYIqhjhHkh48vX8+nwH7VDQZtMi
eEAYWM7LGLYHB3ES1Q8NEPgy1nfVCncd5CoJZcoY2xGan4iYnCJ1I/uqn1A4JRea3qZ/jhjRlaF2
OWsKc6c7yNVqHqTTyoOhYQKvLSSyg+7HOJTQ7zgfqhi25OepTX4sqk61jvl1ugb9oNAukEfrJkCG
E9LKmCfCbX6gazSnEiWTfq5dK5F8EYoaskGZRr7Hf1w1IbqJWglHTwWQtCkcP3gAKPxiJDDBs7mz
DtadR2g/7HabLqzTZXP1xDgd1N4pq5g6jcFGQDtoLj6jiQrFQS3nC7gaGUp4uV+Tef3IWBzz5fvh
TxV2gpqdnUnzMZTCttMtLpgWaos/AosukTbVrDc6rH4EehmWOzwVIVTepunC9ab+LmtUZiPp3Hwz
xZNgDbRptPOyl/Zp4DubD5NYYxDWGIcYE868gpYkf8v7+mJEWJi7Y3MecEZejwdI4vnVahI4lSUh
2av79zmqO5NxLOXe9EMxAto8otj0HHj6Qht5nWrrTJGMbRtqDFlBxNpqFB8mvP1OiH5cHtyj5u9+
2YvTNYNWFdIDEtLyx/XhVWCV/ivrwReHN4YhK6QgOIPuRRLR9ptsO4zwLra0QdNabX0p3/PH8xVz
Wryy2zjYfogMkVrjNg3l027VrRE6Pp7s9V7HdOpp12nv+Qp/5FbwlLIkp/WHY4rTIkVk4+Rf0wT3
dtoEIVL0Elci9+oUPev4X3v83588xj8IzPMot7+1tmV8cCUF3+HihChiIEHXodY2a+SCbUBk9HSv
9+MV9GE2+NkDPrn3LrcTvqkP06aFVCMviQG+nsnHR7fWhZrFuoxbSv1y3QxKcMjkrB1aBrsM7PvN
Of2lWQoVBtZhta1ocpPu30VHs0cQGCUWnC2y2/qoe4j03C5nk8qcFFhnZpk2pWVLT6FRD4ayeQTZ
Cfd03JcfxZ54YmdqDn471owTXeSUY5ydGP0rL8yxAW/3GKW0UnyOlq1XMpQ3uDtSwwWNMHU//XBh
83es2lPn8dWWfVnzn7H1dyBagGpKXH3FkFHXGAFrL0IifEFey69UK6URAVH0faTUhrXbDoLc5upk
3wlOg5USSuqXZdiq6qZ8tOeC7w4DclWjwlySNaaqUJcjroj4J8U4OrCKOUZmP9Ckn6LT/O528cCQ
UsONJx7dUGc8/XhadIVXMg8RWtyS4d4AbqpHtNkmYhutxJXBzZ+pNmMplrzRvu56ogj9MRqcoX8m
1LudXQmsvv696/Ufwz5LXG7wqfoFw4sGlat4kOYQ2cAsItYnQJHUU+FgUpRbdp6CMqymwLOuPpoJ
tanKCWo3WBK+oDI1uiujxsdRoRF5gTBumEC3L2Z17rAi5NcHef30xfGIVsRsI0ZjwMPWbt6R3Hbf
WMOBGN2ID26AtDjVG+XR4+nydZXwXvs9inrwJH64p3kgHUTQI/N3Jhd86biTZ1KCXNS+7mkeYy9x
Elx65is+FCyYdrRfouDKTMEolI2mY+KwxHL1TpeZHTkiOt6inXU5RKZQpmrJ0xqZaY2O7WoqTTBg
dUtGlMFMFkqysDsocRyAk6czHIFbK44X7xBRAHwLnm2bczUcBq9FpnonOEL2F2J2oCkAe/Ev7xtL
AtWH5lWuXB5dnM4BOsIT+5qGdOtzU2tXB/du1LWwTaEtEy7wQiRVGyO1rtDyWpXu+f4DhVZ2flnj
OQ/UMXW+o7Jn4vRsB6Kn9m2XIN5/2SlJWrO193mqzMioVhczji3CvlCJjE60fAg0rTNplXQmwhGf
LCUOAShpn9cos9g8HCe2MvJBOt+o3a1kMvzxkU+l/g/Le9C0PBFmvQNdpnV+LFaDJVHT96Msziwd
KvM0WWNRbFCLyuRVpVdJ0oV9YCV8ng6FSZMuCzth4y2n7LmdADhMw0L3dBvf/o+WMBvrqZGG+EmE
SEYB12k59RdcnTjv9f3pWQHZBQK5RajvkFvLsBYuwyiII1FttHaAUtjXBteXZJiE1TXWUysdfvqu
PxY1QWF7MAPTze+e8uN+aJzFDiwJZWF/QLINiGgaTH7AccM6itYRAvAoX8xNfdu41Ba3pNP2AK1C
00CIpZjSYB6L1V6aMMoBIHRHVEvfm4WRc1CvhcxUbFIvtKGNMoRlrEypPoDbtgCtx5rDEHW2/pkE
971O/0GhpfKwEgVIMYLDAtPVNYmTbld5qrd6YTz80ttWG428uTpKJ+yc51+4CuWdvr/SfDyi9Znx
dTivMvOwsF5+S9veMXC5ROtxAZvDdfKMc+Ii+5T0v3/YxnFsidngfzi62UVHG4TQLq0imKzCGksI
jKjc/PecPs33pDWxOmH3FzxarBoaBNgJoTmp0WF58T+zG7PD9TCvcVhr0JWOfmAYkkunLjYcn/OB
KEmWrRqOM8luNed4PngdFnQbsZFeE8jxaLoQ8rqD3zyYPj2okPp8cR/GM4t9X3VTz4MaJY2VtuDe
1dc22V9A+Efh9Lu0gZQTUGpYsA7NWzk7j8NBBkYkNEww6BWxjeiaD26xiW3V7Niww6ObUCvpd3s8
2kVNU4l07vMS5AgQJTpNm/gpNLl7LFx7xGSKwqC47RO+SMX9QaqsoVsev/3P0bVAZiHRcVciiEEh
qBcgDgN2HpQ4BEVKMu8pHH/cWreEOuAt1uNJu37LrMOJ+rqYLMbj0cfEovjgFlHkhxcX4jw0EvH/
2HFoWrZ9UlYxjzLZS0s0iGAOVCFFPL0978qgMdKUohAmtVq6Yx+x/o+0Kpkl8qgA5tYUmx2xQ2Zd
G6poJ4R59bVFkr8zRNvteXmYmcKA9HZWjQzVsou0UKFOdW6OnJ6cHJhd53m6LNKSemWxTjCtm/k3
ZQJVHQF/YPCYtyjezx+Us1kPfwU73puSGSFg4RfNamy5ETUuaUmAjCmu1tYkPOX45/Y3NJFNfNRC
Vk0ZxJmlqmC7XLdoS28p/ucLNrKFBH5eun6tHROiMa6ry7sbzLSllaSuLHv6T0EaGCG0lO7+KRsY
gJ46Te7Dl3NXvuLR9WMrTlRWpmvGYSJwl0yQQnJZHXqCLoiZkwI/pczHXm0vs6JI0HRUdwUq4sHM
i9ze96hXnY1QfEEdriWbSvZpoYegBMpmI55JtLZAUonMujOsZgxwMFZELMs8dFANUFNHRdC9+P39
9meRKwh2AplElFmcelQH97NiWrrjjRkjGT023aFEe08wTop6Al10RmOfv6impoB+NaUxcgHpD5xi
KBUSstjpxGCnHUC5cFKeLlAFoKXZFiONHyOcKy1v+kD4yMxaJCREskhCtTeg9fDrhqWfGRWwGpz/
pSoaEsxMCRzDzEj5MWU3QdXEX9LNuz0zp6kAgguWGxWJNdUUpGHbkMJRuPb5rFzxMwA4ksqPKGKJ
ug0MAu6dNvUnQtk54F/qVnHY6XL97VQCxnBt/EP+WbMyJsbw0egQBYYE4+AmT+QmR/o9l4INmq5K
crzCu9xY8CvVSzcLBIdvZ9qxG+jpLduRoH4SbJu9V0ik/TgaXbzuHtU4xKUF46SniTlS4iTf8QX3
Bk0I+IwdFZkIR5RWXKvAVFjrLAiD+tyd5LYYVy+Wtxi+acST2W5woBXviFlv333A1/CvFJDxRz7I
bfP0FQlLuh0ufwMcriZySd8uP9/FF7fQVESgrbTzoW+VXXbWI6Ufi7Ikj58rcpvXsXwa6coAZTdX
Jp7+IyrYIiZcjdQnkLDTHI6uzR4jYUx3YMDZmzzutjFnZaBDTkiijr85j3eJa/Ae38OWZiunqUYl
Yt7WhFV0y59j9hg2FPdfA8bNFCeiSNMigXVYgU554yG7LDb59d4PG9Ny7UzymcqHp+FQ0B63mios
lDysaqpfc6BOsKO8kD43GYyn14imADujoDy4L9IccGkIA21kpAXE4VzcK9wg1cSg9qwdeyK/BWyw
SnMTgWgo7bAs5gCS8gGWuMqrVGzDQoWq5zLpVE3uWw9r1/NMlPekV7zSwrC/pyXQceSkV2mtkb92
9QSQ8aDaOis/F2zAK36jLwDhI4yjollMj61u3+C7UPquOLKNClUACcEZRX1X5AcBL7fj9GnI1e77
DyLouE+Dse/DBdb/UbqxvtJgJeQh0w8QQqJMQOM3+KB78o15VZelgxRI3hudZwE/EucIkiaXZvt9
aPhNoigoR+NV3yFm5tIUIlWxLt3075cchZsNStgLj9Ehgf2I9FzZYuji0PsiymfQQDj6wH/eMxRg
RKwCYA36TV3X7UkurpS7znxbRTmbAeVXsxbcbtZOnf9/6HmTyOhyCkA7XKgoJOb/HYsx7jkftvi4
nkEMyaprdTVGWjwZLnEdYQIeKtWELHRIpPoCUCxXnBBh1/Utmq7LdFHiya5bEG0nD5Cf+lTvsu8I
YFK0MmcfuFE0onYe6P2JZipn5vXOk+jSuzA8RTciBvqsSu1rakREt40Iy5n/KHy1mMHqkw6b2W3m
7kQjpJxnhul/ZElnfUTUq6KO+Yx5jtFwA5bMGi9tEYrkSkTr6ZkM4a7dxrFa5wC1FMHKxn3I3S/a
tlpzwSZ/+/sFT8rua1k6Zmk++uXnRHnn6KqLKUXhW0861/H54v8syCnPbEv6JNbdTTJcB+SZu8O4
9gOTK31Wsy89jaTAqNNSIZ9lLJ9zj3tKjveWNMTqgCjdQhuHjYHGWhdhJy3dzjJHLnmJ36DD7EiT
N+vra4WrqkfvB4cKSvtywTHDDOLiZZz3LboD6Re55Q5+YEgwHodjrwWyZwEjDm9szepOsquxw0+t
WgRbUr/uqHROr6TRk4QSKIXrjLF6aFb2it11qfX0ZeX3b6tybWNXPfodJpn1owFIab0afS/Y9wFS
q9nROjO9Zstn69njFISsrJwEU+f6nnA65QRZGYYow9gmk5aSi0JyLnBnnHKOAFOweFQ1YoBu8zEh
4HzllijidCqEOjb94ItAmZLY53NZ5LuAzjFrQPTGmbr2ng+wGJZuVStLmeTnMV8b08SEolptY5nw
iqpXjQEx/qxLvvwojlY0KpIaRd9UHTGhBt57KZBZme/aZoTz90y7M6pls0iPYFvRTLLUr3XGxnBB
6nWxq0RYbiUhCHVNQSFiX5ViUFJFOnoqtD8JOdfkRPHJDtR0URTnefEFkWiMjg08H9MXhKSYTBNf
KBb2aH6qAxRE0jmDg+VS/HD0gA93/cXRW8/na72HBD/Em9EkYsyTWoTr4nf/E9ok0PFsqSgsjGMU
iFgZQrI7nd1y3O+rJF3+RseOOuC6z8vEwruVcsNAVwOyRwL3SCOcyjSK45tV2XoUFdCsfAkFeQrl
akHq6rp6EJr3ZihCOnWIVTjyuEnro7X0xW52GmMBWNIdERcDUrHC+IYqL9DDWKcMRQ5grPWU/Rg3
Orif0Rh88dL9OhHqHJc6QZFS3GGeE8eYkGrmE4u+rEcj/PqoJWuzg+HMsPLz7AA71dOzY/GtPYLT
v897JCcCJipx5QckCUJcSvhrTccoWlov86o78jsvRTxA9irzRmZu7eqzR5msDQplFhfG/84kLxgO
ykPHX6crYGpv9m9zGlyPOaohlRtO+UNqUqELtS8MEDNRt5muSjr9V1sX3BGHFVoxYOvI9qpNrdAz
z+PqEFb/6CyuIPvwFRvn4h+GjcxZyoEa1vMSbgosKgsM+oh8JD4NhfWSVmqvXAhbDhSSrBmEo7qB
u+toZ5mkj9/E2hv//w1PuWvxPUC3sd5SSckseymQ+bH+BNwrAFp80IYLVVmBTKv2pCFRlp7EJzNB
uiOeroLo0mF2wmbnuodi8LqMHTjSFPxwmBaVsQXL6PI84hxD99X2SzApXXSd8TqUNOLhtpfacvtY
5w0u2Z7ybqyiZY0T1LAm+haaKYqNDJaUAHw+kJ9hNh3ltSztwbwQUF3quHCAnirwhI70VKJoLqdL
gogHThRZgAw6JiLWvOKlpP+2efCd66mKwebYkEpvczd5sGr99tyMmqdcOXw12t1expX8CHpiUJez
seSbbEpi0LmAj2vGlmCMZfl57H0/Xr3CatUG5nqrFf+1caefozcAkhcO4TgDjuAQGSfEfu6JMUZq
D6xYz9PgmjuGEOk8n64ekCCsfQpBnFxigfu5GyC0WrgDJahTg5oR++rIDNfnwWDZdw2dFkEvyKZW
ldhFDWdiz5+S5gAgnTWI/tRZLerVrDrPKZvUwFqQY4e8P/t2cBRkN4qa6+tBA/sqgJAuEJOcJkMr
K8spOHJqJNPdEfgG3bvVYL3WfR5E/MeN3i9v7J32Ih+ZhWx70UqQE/xr1N3UXiFT6bGctoQfJKVm
graULRaitWTK8Ha4yfZN0vBpc2p5wHMFO0MjOdxXaNngQkKzgpJEquOgLZR0eQiHO+lnvaF6fP/K
sMjlYCBH5P+EwCsvdl3UKwk7mt73cf2shjGNzCI34vNA+TxsAjG7/v98944wJJlOGHNg17dk8P1o
NlfvJ9xgTLRtVOOpXTsbVQdy6y5lgou43cu62SJwRZj1QIvx9H3ABZu4RcdDwkkq+GTwOT7iMK2n
EQaka6HJLWzJCGYXi5b1VM3aqyBFr4xnXQg7A46Hob70xAJC//lTm0m9w/bK9NNQk7GECmbOSZtd
/YN4DLqaS94poMFMgGRbe8PG+eLim0aPorD7svFEF41xF0GaecWLqg+K9aYVv8BSNgCv3hkSYLrR
yVk5aPJ8v2husqYXPSl7RZgRFVnymrKZyMsD0ZRoLYKzodhDahdTJ+rS0uMJiGnYofv9Ppusqunl
koQ2pfG9PZD1rudC85kOd3PFWHsvznEY6GhyIjBsiuH7apmLyC5ZHV0npy3Y1QXMP/ENujjReBV7
7CUaa1IW5p/M5QeeONdYZr/qSLeP8VJ30sJ4GiwQPzuxVgbEA+4DO7o0GR0U5c70ln5BUjkB9fqs
KuUX9mDxJ0s70lBCX+1ln651+AWY36iBxd1W/6Q9urFDZFl83bqhdY/QNVpYChF2T1IkmHej41Yk
ERKUwTfylqfjN8zf4RVih3NMdSld0PPieECGUE/HXdaWDsIjYSiJfXQr8rdpLMLBgPCNMnZpLmqI
nkxbTxpJkuwm490f/rlymEIcBfLi/u7u5W0jwpo795aJZm+kP1n3TWidn0LnHDVYxjKB2VowVFRF
xq7LhlpmhWyBxKXsDckqVzCOK6ZQalnY7rdqh+V5knwcKDiakl0h+bTdRQy+bX+TpiOPpDviNHnn
2CQPtnaycPLw1SsWVgyFcEQc6AbpsK6QnATMavZNQAr4/ZNL+FJxWUFL95bImJwVJu83rQbQkuqa
Lgm992XQT1+U/E92KWTQ56m8wutMIco6pvJyIpybbBVhvbXR1k0bB9lHmOE3T31mVZ0ubTAa28Bo
j+D0dYvDb8CIYaJNcqhF+uBnGD2EKzms0yUVFZgSvDYWL0Bf8GV/nMWJQjgei0AnR2+dN3hxs1NT
ghn5rVyJg/oASLD6+Qt2M7CQHMYL4dUq1dsekHZHt2fPOROh1Cq5DpKuiIyr4QG3dToAWa0yU/5w
ry8npaC28T0wHCEKHSCoNH7LjfqWQirDUQvhavB1p4KrhYBTp/8ZtDasPMctXY1kbS/Z//f1xJ3S
QuRunHcdfM7UJWv5wpF1N7FT8+1xRDh5S91VSOcPcwFJfoIE17XVZyz448z8G1xxalNShgT5YcjK
hrxR/lUaPs2ibAgjxaNUFAYbAgDbvMVKe+pCexaOXnv2LiuyS+7nzEalXGgsAzKageXlcZyeVISh
umH0jOBI5DIRaGofo5VFH0AOJQMe065KcId+lTnK7e42wmw11IvHR2M+G2ll79L1aj+cFI3msAj6
d5kK7IfTwfGi1O4COnQ7AP4PdsMb5LV2Fgf/6CYR4oMCIRHN1t7NqJENIzwKKpEsS8YqVDh7baoQ
3ZOgLdTCe5XDxfIJauisC5WuKNg4hegwVjJZJZN+ifaejPVzOiynR8NFAOjVaMSrbAeQYGDlyJ8x
krxNKQ4oWykXN7PPZp81E1qikmkJLLZmRCzRiyd9d8p+W/nFSbueivZf4uoAaVV9v1J0l5Z0BXl8
AfZTAcWZxQBwV4G0/ck0yloI5qFyvBUovSH08Kr6Y2+Hw2DQvrsgUuNZdJaJcv+3hgthsjEletbz
yhDGAXoDFhHEgmQR6JEfXYRH8hL3jmq3kJX4R1GWd9IADjPnkKc+XDIake+eaMrkGiJy19LTARb2
4zDMsr4uHwLKQ02T0WZQMvZxpZSA34V2WJgPihaGE7ekHt5RyPtQG/WavPTFNyanfvjhrs6M+x0W
OeYMVhz7AM1gxE4lfXUnSXhTXuvPr7BPfcU/4PPCjgF08/Mrci08ZSvrFonanpMJTe4BESREtZpB
4aesj3ej9qGOpRvw7Uc+GLhhA65CLYJ0iiPUmE4uTtq0pJ3Xaf2KyRI9j9i6sS2i1GAb3F9h7gCx
2DGvRf5MdAILSdYJmf+QTA7HmnheECk6pTGvS6gISD6bBEZ73p8EPDMNFistXuxBg+05jPRpx75f
L8SZfT7NMTX+rEewmAeOMvWBxMGT1DjoApMewNOuA/ka9QFtFLpK0RUqqvwVP/vZz31VoHByoNeU
BDFRT3GuYGWGr6GR8MJ9zA4QZlaAu+pNsoL7SkGJrtdB36JI9byBIuPJpybFzoZ33KLO7jzHmSMo
dbRXwuSUETu78K8wFQM8T/3EDbJBSG2V+rMoA5FPM0b3sHsglyrqp7RsIxG6vi8SOuJhpOqNmt+1
gQaZX1s3avdITgn3sjWIbji3sSiNZfLO8h+IcsonjUs/LwCJ+EFMBaqpNTMP2aIxdJiE88jwj1M1
853yrk8IN/fQBj0KRTVRTkkCiyWyffugmULDqZCUDfptwnWb9lD+I0AGLwf9O6tfHqLsS/XFJzWV
+JN4NiEIJSV3Zmg+G1G7MtRBObeK3hADuXrbslyOemIMJSXYj4zZD0C/MJ5wGCgIxXcD7EQU2OfX
x3k9ScxHMhpcMjrDGLXXlcZoOgue35M/Up6Lc+8Ktu8TsBTwLkGMjLdDKDadMX/mTGHZaZz+C1VY
TqcqhHvYRM5bvSjbzPJULcFRkx4eLmqvakf8wGJXeUxOY45iDWIiSkvESIwCQVzwLtLB2QrcAke4
CtmBm9Cvv1GlXs1aTNdf7hSKTNb2By426D+OIXHEZPjVUiDsbmOPrUSuYIl1UYgF+v4csWsy2/12
kIgy5fEWJ1ztLkPac1m2jX4WqR3SA5gsEnATH/5nuF9DzzVPl03d5Cw1Y1SWkdj6GCOemwW9jz37
PMvSwwQQaRj/sq6q0jvm+9qckdZQTLswVZbRU6AXbvfkFpgSKajwj5Z4+AIHTP5tmFOYXDXegPuO
sEbVidlKI9pWEvUsod/xNVGior9x8VY75volupyIeDe12MOr1UmdoLiCo0X+RJOZOWwttxa1X7FM
wAwGEiLHvEtgMgG5InXg69+jEoXchplWFSQ9/oUUv6kBoF8pgMk71wjhnGQEZ2cOBkas441MBRvo
8hUF4kcWon73usEmUiwGBi22+Y8BoQOQMvG+cs9zdLK/AelKHpPqNczlxNwcRqtIGrhpMQbUfmK0
OblDOijm0yw2Q64rYJEjTltEnA2TzH1rxkJzkzwPXH/LFV2I8bhoYLIRumzDciDDQZtTO9/ffkAT
EUNbHzl4/Wf5RTw4QrsGSzFVhNpi/sGgkHmGkNQ1LCYJJGIjTGeUiFicZI+Mf5OV+YZihgxunQ4z
2E0vg4nAmNI9EVEMD6z1tBlxvzWA97XRh9jv1oGjJp+mg0GAEXrMae0WRLG1+IzhaZhX++WVOW3o
MDBQivi6+swjZ07jBie8UMnhJ7vGeSXV928MyTAz6OSapPZJ2cUGGADo89vD6KwgX0u83BUZVow0
eBSJ54RjqEqx6CaG9AbC6cr5ku3PE7ZUrlqzxKGQM1fmsxl2hxg4UiYecz+DGOqwgULkp3uoa7g+
ilBAbN4uN8/3B8DCApXeshltC2Thwd7iXJIpBmc6Q9od1L4w02L22ecadOaoh7AE67c3JVfYdNDb
4m8slFHj3c13VRBssXF6eWKCmAlX87JoFZtuqIQo9gJPLEDTs8ywPooYGeoAJPDmtIxdT4WtAPN4
Az7GG8XNzSZPspevWDvaYpM8SlpGg02itY1PeF05F4PZy04Wo1hEei6nmuFW9rJ2mPz48fhtRGRr
zaAYpY2s+6xalwKwot3s18Mz7lJ4vVJleTxtVO7yy8exRgVlaESbms1wxET1f47X9mir3LV4R2Ql
HTI995sxx8btWIVPjv12559fYioNY8DgFZ0Fj7iRFjngyiozIjnNLxyWomMK/CNoBS2HnJE7mEYo
QajsdEG3isqWmH+vnLg+itGRUHSEHuuJXhK6onKnvqf97tUnbZNG3e1JZSKIv1WCpU3Od2w7eO7i
Wrdv9e2srRDwjLDo+CSXwBHe/1r+fAKPMMdWkQ1x9l3NlCJ3ObBb9Cs93bfNs6b3QfBAcGGwzBeR
U5xZq3POwgGv01o8ozLny57wz+rV6WqRJjleu0YzaODUUviZJLc5XZ44xOmkOtHoGWh9eVRH5cDB
9S4r2IA7d1K07lqzpxkvZ3hgl3A3cQG4vYUKyVs/MKfzKGER38IzO9MVmF6rz36o9DF4Gn3DDRoF
1iEDeXdtCmC0x8q+9C4kHg1Kv/xT65Tmj2I+H3rbo/U6xQhcGUmLLQBzmiK2Dv9/MJF5QRhUghOd
Ad9oh91KjEivCv5U7kAkQ30GW6yBgbERC4a1yEJJ/pjVxKDPPgJ8Xii2y60GCZWvjvC9xYk2bUpc
NqStUoUJIb8YwJQCf+sbWd9NI7GvM/Xy5uGcaqPNaZtACj0DynoCWX7jP3NbkjWe+zNKeq0Hml/Q
CG54jxp42LdQ7ciw/JZeoHQZ2YDokCNL6vcEBg7HFv8VdtIVG2lmpkuVkwv6YgImo34q55ZU+IEL
81zoW98hgyF+3k0BuTzBr7UhZBaAPBjnxvrrYBYVR15IKnhbql/UWVP95IOBD3Yg5/llInrYZOy4
QVw2hNuLhpAyNNTdWiKr9C2tHD84azytonUVjMrF/qY0GQSd9ebWxrWCD2LwPaGvOv9mQ4/JDYD6
des4wF7CiUUTVPxE4MogdH+eDo75n8N32lTTqbKlR9vU0eGFmrXzJHnHCq4EHsOS/6h8ozNDqpYs
53qqdUZybXjj0Af7MBMBL7TQPvqXHD5rn74YNlowHhQoYJpV4bh12/w9OESDPqFdWU2KekUaOxwa
NU9YUTg+YCRguwGE9qcrx7Gfj/HvWp0L6LojZK59IxSJgc1+paVkzyAwkl3rpFF670Uzk7Y0XvcD
XVy+3ulmoeqkcTl6VS+9evfOS6Kl583TCqgguai0Dfwr72LHtpUn/mfUjzSfAJfnUmIzFVrbCsp5
hcuz6xMA4nc/zfgY0VGi0c01rrArKLzyzwKjetcknnbaZr11fIS0CTHrIoTyKgr6evoCDrvtIpB0
SZvR9gifozSJhgzAHZIWoqIMDQCFmR2C0f09TqDdhCm+LwVDEjX0ncUOMJC7nfR5eHkepzRYXDXn
DbqtCGT6GUEpLZZJC1UwdAkJviWJO7s+icIXmLosrsZ6lhR1qpwNo2aLCX1slcUPoVKoTkrSH0U1
xkuuZiDPJgz4bYwqWlQEf1R6THIwnQKVjnlFt8bHnefNqnVewcAqdr35aDSeu/hAYCNwmlE0x6mo
CLCZp6aN+/aY1FnnBAtlW6IEDBE6UKsoDrN5ZLg3N7pAFmhr5HTRRPKvi3ds3FW3W3ydpqM8rtLl
DU/BWp9rkwLT3uy2xbKq8josNXHCDWcZ5sHW6cbXreTYVwCCBYZKszEO+MV260KEcLnhta5Z6BYw
C2IfOzqBIbOo9ZhkrzkTSW5xJSyj79zFK+k8NQ9TvqFUDj/AHGN7pPsnnvRuZLuVBkaq3i+fZ2t9
y9P4oZ3UCXJqj1IiidDDMPfkmu4js38suJkzz8IumI91aBmT/iAIIJiS2qyHaHL3TfVRlOrhZqO0
/s8QJBAvWymjJX58U52VT26Oo1JUqr9JoByoRUu9D4Ls0SPuc/hqS0n9RvMF/D+sxpkIiyimx+CM
I5lryyVlPR2E0k+/r2IEbcKf7kv79NHXEcxTL9RVKICEi6RwMkbgPmUDY81N11MH82WzZ8MdFlxK
qD5+ziO/loFYRQbTAfBWGrs0RYRSf4tvc5T2Rih1YtQY382nNtojfoU7Qew4Pp/pZd+hdpPSgDMB
aPR9E/k4kMEjTECl9x4rkgxEoHiGIEJt58d73FtW9w4lkoHoKKK1hod1VWPWKPhUnmy9lZI1/iwC
nhEY3JK3nPJRhNExtboAF8hznWamhjmvmY7+oDubXadE7Lvtz5ykiwcjcXIB044R7clTRgROqoV+
hoHWd+mApZ4ZoaofZiVP5+gU0dziEC1FAHmeJsp3W25pYoQGlzgnXeyARDprQxVoBYoYRyj4+1yt
XT1VQ5TEnvcKhhf1IPJCiGzpln0Toow2l9Wq+qPQGaglBaDYTeSU9z90prb9Nt2OhWuLjwV6kvyw
QDQOII3m7ivSs7FCFZkNSug9u7RdVnAm2BWsaOWXwkHjv6XWnfj8y2+fhq3P0hkPfSXZ729niExy
wWa/pj0YxXBXuyhqxcOUVW3lz6AxBHZhB4ZvJzbXlGkmJtnavje2GjpLIjaPZ09RLJ6LC81gftiY
gA94PPBrEipzb4z33SuBf43EZTt0SwP4RV1zcuPP5NaDNJhzdu/fhlBPt0IIzQK54PGgL2TX064i
FlCHBckN1OqAchzegW9d3ZBKW6FkFZdztGMpV4dLtwKYKmcvYRpW1qKYNiBOMo/RhCeV5QyZ7h+4
+e+Vw+xVH7XXS77wgu7L2oRyDDBD1C1kPH94Ac5+vTNGfVaAiLLruPedqnRBk7YD6spnznSY2h4D
HP9e4AWFj80JXgCte58KldPBSesn+8ipsl/c3U+RRpbgUHl4eIIZEi9R1bDKOdu/OtHV2NUSgqVW
6m5Z4ShKVx86So8VwPZC3KgEKb3MhPJS6c6gc5/mvqpwVxWvbkHnIO9+D099ka4HeBH4RnSwPxe8
qlBQrPDVWFj6xeOhdktNPsDwCaxQhDIsgBU/noHGcT7u/lm+li+nHMsj1aWoeI4Ou7hIxOgi44jv
4a1CcfQ87JH0dVvTGd0fF1WkOLa8JpLZshdnYDw1FlmQWO/j9GaDeiDZamyYArKSvmT4f8wk+0wt
KrA1msVXQkXcaJnXy2pM06fmgYZosF2nOBPqVUOTl86Jud+3/nIl9Z8VZVKLFH+Z3qnJwzxJ+V2y
KXyfXcM7fH9Ac5yPQOLGR2nfa4XAQnwQiddn1Dy2oUXQa21qpCxtXxhtnFjb1jCoDVT3w4dOrtue
McQZjDjUG7EUnIcgi0CbBYjyhAfqUM9VroH6WG6GBmsV89d39g/TU8SWPK0gM5I4z4rmEgSEAHQm
MAU0RiJWz/Tx5pWyy10X1t/9ymTKHR+EKJsqiT+YVLE1c0uCcMdAwTbwO/jIakIbiKmtL3Docogg
PLwL1I1cxDQccwr5LnZkl6hekcg/ThVEav3ePTinekCQQ1lp50KwBhaq9wqlEsGbjkkmNYlRs31Z
GNUbWnQ9/4K/CoqrG3N9iyafd+xl3tb7r3php1t8PUGOBAI6TBuw6X96/igABLWTVXOaAI9rixw6
f5lKbSJFKhITMzX65fjKcOI5ynovCyoNb3pqLcdusp7UaKQ9p+B+niK83gdHkhKJqFRuuJTyz+0i
5LSSoohX0Vs2+qWWUWyIFQoe0qRx1IwQ1BQAF9obMWnViSzYet9r5swB8vilVLM9QykPf4uQLWjY
EL/KD1OWOACOB+eNROYDYEZ1FKfc8ev/cYbw8vxsdVzZJboLIdV6g6fnPOZKXYDXV95hpgRNS+mV
RbCQgyAbtUYLbwhe6nzM7sLplrZbmgMaXwaQ+XFKEr1EmmLlQBVbmDIO5Zuggpnq3SGZzPSJ7NLJ
aaya/lhWCMiC3oyGuLjgQx8zVZP9CRyrLuYTWdfDlxjU7gg0n5ZbI2wCuqxTNvOIm7fiTWIZebJz
T0IKviyU9t6aCSJF7YfVZJ9B0QVcpUu45Wou7IS7FdPdDc2ZJOgLZ+PaXx7q/vjInJTplsSCoF0N
5kOSaweXqa1LPyrJXN7IdjwkWMBOJpb8DgndrXPw0MAPqXMOFG5dQakACkBhLYYlcasbgr5wBfnt
yTkAC8mOHIMNWZCeOUE76F20z8oFxvuDj5hqrQnsuwVURoXnUm1HrvDKsGGpeld/iu8BhzzEK+W7
+G7R5XAu/d3WCl3P76ukjDUJAJBhsauIOBLg4MH4ZTpK1s9kktbPJRr+rMJ940T2dawyJ9K9+udy
yXwMjidpTMdD5Ok1F79mRbAf7u+gjOsWFUShp+iafV9UbHXfLsqrKR745hVXF9XdVyfVBo7k/BRW
cCQeFwv7aKufaaxEJKWOnrtsPPEIEHmR/xoetJ1OsU38XOhb4yG1OJx6QAQO+PnUCltGFRSlVSsf
Vc22v0mePcHVh1xFQ0VmgY4kTniHvqGtrOBmCbXqYXEdCxzkrLKyjDgXXlWyksDUJAxFCsCuXYBk
fzfVaKAVR1oBKiNDwrvZUwtj+LNz3+T6H9cmPDq4PsXty6tHp1RdfDyIyrLPz1VrKd5ZK53CGYR9
wUc29c6siFQiyNrNB1SrRA2Y6NkI7X7yJ6zZVGx3js67YV4G9tkZaZ+cOzx/DeE4WMJDNRhjgm7T
s0EShb5s8u59lJwRwa7ZQBk6HGsw19WUbkcnztDlh/PJdRgdbEXKiWJecOoK/4P8rsC5PMzjmez2
fuXyoAmjeh+uSobzaI6Lxp3C9D1wpQ/pmPakLEsUasWvfkOl4YycDt5aLjaLTNHx4PCobByjn/Hy
fUcNIBgbtxDsLJtlVlfEMGtqjB5NaZ8P6w8L6o5wXzK2b9XxhCww7b3FD67yPhGarxnz3uqYf/cp
KzLZYVQxAtpWslGU3bokAuqj9lYfUk4NJZgX6m3rIj8OtDXVdNIzVMc541pcceKFB6jev4+KMwC5
Gnq2j5ezthKlwYeJagTikw56GZY1NLZVP85sg/iJ6UZTjs+TUt0QqCqK1QRsJ1L1ENFWUxBRs4sC
S1fHp9CBmFBDSEOs7my9FqD1qxehxs4VfDOtpfDFozCIvO8KioZ15WrZjgGeTbsJcdRscG6gAGdo
5ZX+J/RTuCtPDnb97GgtwpX0usAfuM1a7x67l4HpqANytNhrWGFF6ARsDIey0z2NSyPjlyB7X3u5
H4sqjvJ8d+MkKBRhy9L6gCOphihjiSu78kYg0d/kqJ6HdqmPLJ5TQIDaMsP2Ijo2LmI8bM+LyLC8
fRwB+XcvNs8wJpyczE9FiuOgWoBmKPRA/KPjF6MMN/g5b5H/8eaRekqfrC92qqbcuBUsT0whvmid
sjgigZGWiMVGm9qsTQU67bEaKBxzke1qfttrGu5YJJhzZi74vO1/QjpHENlqiSm2ag1noMOQDxqR
v51Cl9LH7hKV9xBK688Cc+N44E6TZbqjWIYX9TbNrBw76HJMZ9K3puf1BmGutDAFXqE5o2ccTImt
qxb6om36OcaPi+25g2AbWz5o6HUb4MtwVH0oWqH+VqzhMqISgZa/zb2Qa5uImfftP+YaEFiQ6tA0
RxEHNjlXWlmcFPUzNeug4a2fU0/rc6FbB5jVxzKu1jQ7zhpt6cOObMozkX2meS4UKnpSXQmFonfI
8CLCaeck6DnCErQV6yLxsIcYiVY0As95nq0EFESESTj/nKyY3Si5fp64D7XHAQzi70mHgTiZQv58
H7YPh/vCmlAiq37mIWW3KcpvfEpy3MZdTbCSQkys1aDbS4VEQJEGiRrKk27E9f78S88sPdV50Fx6
E+du9J7i3iZBh/0ayxXND6U8FlZDADUX6UPxRRfSO01PLhNSnsQUTN2lv6zWGsXS6XS5hLSdKQxT
2Z6tAThycTZ6c1+4vXA9CZB+fMtR2BNxZ1JLIn9FpC9rzTvcL0cr2VjflwjeOIj7CZO4H80/wKoi
Gxe0H7usdcevTRRoTsAetZhqGtA6THQhJDdDyGAMPVLhibMfA6ecU5kmLKprJg4fkWw/jPgwq/2d
Kxi+AzNNL6LqC4fRF6m5PdEuw9cpv3tCwDWd1sCaBBQMbLcyjXhCnmAfZwiktySIR4mAYHocChb5
Zp92YZVG3GLSji6SMDVfMddnGADAe/wVBcQ0PduUQfu1P3TRQmhVQSML0Xq7lSBBRxmb0LWsX8G5
8FpKtHKTM7RzUa1JICpFRMCn5PLpwFxMaXKM6LQA5wEnPtZDnm0o6DJ6+TqW2Vl5qiae5ilo9KDO
U8co/DMIU3rqfqxjrq0SR3UcnXlkA7BTEI95hOEuNyT30IbvnqWrj3VJxx+k2fZvt8AIOpN0wVoG
Guddm6Idf4I+ckpXxitsq7VeNH0TRwRTx0VC3deLw61d425fXPlVm+28tajoFGrJ9rzGJhg3GKrX
h2zOtrobaCzFuX5b8lo0Qxhh41K2k6OqPrqzD4x6+3Llk1EbXm/VO3Qyc0OUlVUDBInYCqUlibuN
C9nQRGI+ZAaw4GVNMdXRWpgfkiyOu5iGDhqOuibL3VpHoLUynHS3NcaJ6GgATH1FuX1IZBI3diBS
nbdS/0rWax1Z8KWsh+efE+vbzR84wJ09C/hPJEJf9tA/WRnC8WaI6c2EKCbihBysW9MMCmxQoMJE
WAP5Nik+NtoJqPqbzoxxx6forVPdU5pJctY61QlhniasxWkcJ8vo3t4gwmbBWXMgHlaxJotVXB1v
FvCYBGOqe8UjTc3gXUma9Hxn137X0t0dK5i44+L8H88EGgErAltOBYbAGWDHg8g1A2vcfSKIBt1Y
l4uEQbBobF6sOdR3o/dTLBfzfvShQwBTbgFG+aNBk/GFUT2qaZxySyBL0+EgRtGzu3Hbf9YVfADA
L9KEwCWlx7W1vMa/SWIiNS+olxx3//CmXBVg4p1vhhg08E0H7UHEECM1VvVm1xXvy5GktxaOCf9b
QrOEWrKCrP2g+5QuzpPlAPFkIqzUrpeA2R6r8nTT4TsWrM80bA5PRqABVezL8fMFMxW5870sUjU5
BhJ19jWsfojO7fJ2Mr2/Jf54MHvEAa/RX9qattMerux14VyDifgLq1onu4l9bMg4Xaq+zc7sVZCF
kt5IicYW9nDvd4DAeJAPdqNqaISBl19L1SwQzQ7MkGGpKxQommSC2LsN1LSx2cOsS9ZnEpKcmFp1
WRGZ//qqpYyevrZpt4EsNSbwwTPo5R4IK0n5Nfsgn/lwmO9QXZtebwr3J9YVWXuoHkkshFrVs90X
eL42uOhdnG6QvTE4b7frb0HcTJFlRR0nrrvVr+kb7WY+dddLUAvaLHSHFu/A4LnVSk5Jyl7/jNo0
0gqELvb9Cdy/zwXuHxE5gxbp0Jq1l+ZuXRN/d/TcD1HoJxH15t/U8L0tSbO5bpd7WVir3EOzZ8a1
f/GG9KuOMx6XyV8r8lp87kqS1pkS+3GKHrz47P3sQXP+wgFBhtXp0hpPbpim0DfL/IRwNOssfDMw
J8+ao9eSuXKh499MeJrVbKRiowgnU/icqgm9CiA/WEtHfl8xs8JLLoGde591JhvLc9ZetYhFe74h
82EGYWrBsrkMOvTHP7+WGRto22le9g5irs4lkfwToTZlIXTXwpyeZnyFktyjNIB9GDgPLsxNNrws
qJFVpNQVy/u8nhiHR6t+E/glNUKOuN+8yn3QyzufuHI65vS8bR7K99NJW0SH0N+e1IvwZJgTKhd+
PrbCjPaFKKk2zU+ENglpqXFfxtueZauu9Vo8OLqsDZLZYvNsDRoQu4Hqtm89ZepUJmE1/XfeWfwg
mTUlcjS+gEIfHApULtlUPr/hdsITQuFdI0eWPpv5ECIf7OXwvCdSlEOcLH0UJk/ytNzIPkwGikBq
uLEOweCBwuJ44ViU8xel2f9ixyOYvUBGe9LmVoiBvWLog0h8CKDTSNiTCUYGp0ILpcZbhxAHr1ao
BifZiXo9IYRwgMXz5roIhdP0ZgiVbHLsa15vTwzBqD1Xk34TFoiSL/OIdUK9dfXiCGYrc8d9xPve
1WT8YdPmTZLVb759LPKf1JUQfL+SvnYsS25qkyPB+0k5+5w87DYwe3GtWucL+gjCMuvEEAa3C9xD
Gh566ZN/X1CuWJ66HUK1XvX+ButqhzDc7VNN2TRwgITzfuYPdhNhRDH5UsIfcmupYMJ4UVcbhJ4x
JxMvlZW3A30zaNAtWi2MBsn7/+OiDKOcEMxQ4nCxXEsQOCbJR2VFQj82KgwKsMeq47XTg0qLLMV9
azPUdgZPgWFNnVdDoOgiiFQj0dNIPxbhX62JmIOer92MbVUI4QDQawmd5FYcVqK5j+0BPI5J/aRe
QSzGDCZXWwaxx4TmVUmzpx+k9TL55du6io9pGSwoUpzahWdD82k4GF9Z83C3t5lxJ56tvkvLoRyE
XVELsVT/ZS3bI9Kr4tJDpOtJVsJaxw6g6S2jNZyu3ZeXGEPiAHgUTBbUEXYLs0rpPV4snyw+mXny
itWrgOJiQwv2hpXVmjfYIRH3RzXRYNHg3uEF1Xv5xpSDQ8U9MVixfPRSYQG18cFTzviSgnr0Y2Ky
qX+944rKIwV97MfdO8TpUwrEem1W0l/Bvx180GIZwdbi6RsuCurr9xWyPIJEs6RtswzCGJ0HT3Ps
AONBgMWlkbujv8JyUmzL2yJOCUYuwVOyjMR60ASqSomURd5xgywddGwpPp7HAh57cZyDzcUQePWr
sbFcre8y5cqqloyvXEw/49FuW+C+2mNcRRWytnFX/PyK649qV2B17qaOmm5qVkqnOMOAjW97v3Ef
gmAxR1AJZLWSD+4PKKK28/lptBPhXWFb/e9xba40z/FSovKAWbaFz27uo6ooGGwjhgsLcwCRPAQ3
RdLb9JbCQPZ6RHgMzPcqZaVZvCvYYtijiFBcFIsDD4Ww7f/kM9cy++YUE3ofk+ytZyGqBxtthPOo
W5IEjAYxb5r/qzX4RhNCHdpT3HHcKRLOPXe8kybl9CRCbxHrlhdxbMpjCToMd5DlxF/Zy80vkW8A
Ow7Y+QirNFwwXZD//lb0lT5rjH+sleBx4lzNY9J29z1cIQLtKTIhRUfdob6CMOfcJIczTNKyxVWv
FBe6/7BWOLVKOERY8FlpZPw+QhaV8PBHSThahUAKPlQhqSvkBaDTY0dwoY/UStpHGqx+hNR+etYy
tFKSie/8v8voKgadEvRcKBulYBEb7HM2UZaTTb8y3ZbWHd1TfkahdyaYvISUq8BL85V1MeCLrNZ1
R3950/8R2taPnJlOGkVtaNjMNhrJP61tVBSOE3y4jXLxf49uf17X0GJzR8Kuwc5RkoshUMDF7wUS
Ml1ZSnBlCV8gX8JvpF31kP9S8IE9SyVnKjif9zs5ayBJrzcbtV//K/MfkqCrZFWa5OPTqt5kpL61
hr1Ab7P1JIQ5LxEILTG10yaX57wEAEXxTy5fhW7MSNFpa3EiRuYw9UnxKihlx54CHenfjMmz64/5
cbgrWmccOlvr9PGV3PCYa9Xtp1zF/nGvplVRFtZrL7erGIKortw9v12bMbRQC4SJrQ0NnPTaj3UU
dHiWtinDd6bPCUokTJKgb5SxfjmfOb10dGy72SpptTzmgkClYVSyobMJxT+wBUZE0QHQjCEuppVC
TMwq41H3p2KiUevCI09w95Fq37VOkW3LRiza4WoBR6/C+0NKLv6vkubHCYscbUGdciUJ9WNCW584
ba4OkAGhQbZqIMv1S2tUEGibb3ncj4eEJfnpt6VSkjBDj2sHBq2UaJStT3rl/zcy6pokYf48yqO2
eWkHbmdK5Sw/jxMTEtSAu9wqCUEIWRwwd32obZaiZvVxos/0uMp54cOwb9zrmn9rsj5G8RyVRddH
0ZiAUJEKA3SUC9zhPxedLOYkE0mdzuXLJld713uMvl6bh48aWTkBsZ2Ian50ql7zn4vGqN5N3e4Z
RXIYnjv3OZXP5s9hlH/qu2w+OiTVZnxOPwAEwbD3ajBiW9dFFIvJ5rgJ0NHqbdpzfSe2VkUeoO0I
C/KT5mxHMaCPXPDyNDaFhPo7PoSA+f0nCCe8vTIJE2sJdAP8TtoVOoPJ8BEiL9RPO1T2WWimiXFz
kFxeGcF6u/QtE4QnoIvwZZghasbVKV79IenbElvrbjN0qeDjO1pBbPDSOa+9oIrow+A8FCD1iQjE
dSrM2bIG+yNiJGSMSmP1npMY3/aIzr9g9ea9as00ukTz5kgD2DqRZDTxPgLRY87ZHcL7W4xxTWzb
E3nCNN08l27/KPeZjq4TqyJumcKJrlozw1usMsD5NuTHpYDM/h6PIQ3jMfq3yOOTPujaNmGhFwgn
Bq9L8H6QkhZ7YOwFrxO9dHWISimSmGLOoBtS4R+9bk71tJ1Z3YOTzEh/mD2KM7fgkjgLapCmiRUP
6rinoCWbRYIc674jKM8yYjcgL6TtvJKg2YoBi+VK15GafflPmhvufEtvhZakAn3uhCkvWgYiSjr5
Cmy1btNbAxKRZdNw0xH+Awb9RsCw8q9+CzFFu+JaCyGPp6Ednk69CMS0kYrYRHdAT+ElRom5CX3e
Na1ZNfkKMqy+pOaRym/yQlHXHoB6wHV2eqycN1dfg1YsZogVSBintDbE2U3g1fLl5W3FcThYawHJ
g1rvjvJrcxRFiX4fiPncbtorHkQAaTRTxoNOQrAAwWNnT0nVDQ3ym2ajG+xq5fabdv2WJTPTNqFL
ORGfFIZS+yL3R3quXaXfHXQEGJ2NllKcnutiQUHhHC/URzAdr3atiHfjSAKr93jYG7ktszZQY1AO
cTPs0inwrxayBW/uG9dvYzw6OKZmY+RZnPIULfECQZuvmn3vCm1MtIbDbyOrpeNR1B6JOr/iCnej
/k7nkOoulQyTc9YNaI0MtOlO/so7rw1cd1ltH78ie0fcTy/OCvzSX1R3MAdI9B8BCojrLoN18lmm
Mm0y2DRCIIDIaGdD1vJmGeE6J1/otBs2DNz7L/eNXG5qH33xjDtL2EjKl3eWfcFcTMs+zRy6YVwr
vyDVIg1jsFQtUCYR/A8TPj1IstmZDukMOPSU9s8AguRVjgqsXf5GA/roohTHLZAYWnbWZU0M3HOn
0NNJccEB553nfsNSEL7KdJreD/6+VtMW539NdEM/8Ks1HHfUOOV7X663tCcX2xqnm4TLXrdeLN9X
M7MEFuvs+5/ke9t7owoq5MxA2jCQ64Mwyb85RT50lGKvq9cOBEEtnDhcK5XiUWLLWpdBrwXb6w9t
V6imR7MmhNFzdManS4mBnDYsU6OZOBiqb9dhWcsOePc2bjANpkMSi5oT+D2RIfkpFVuSv0vEZ865
Qu+GNyRdcjAwAxIoFaVhRzz5n45Pb97ABy/sYheF2msyOm7W/2WUxhUudAtfQaThVzQrU2xuBzsu
hIfJDLIHkDEOC6cFjexzjC+vgaR5W+TQHExb1w1Sl4IUkr/2PtWN8X6IgFqgNJyd2imBYxcN0Mqg
aFoHVyNcOKmVabeiHyzvccRYJmbIZFU9ArKaq/vusofv/B+gyAmYOyNtD93hx8VMDcv+2R13zkUO
WTPXFF8ek3VigkBiQO5QkDWghQT21GXAjNP9DR+xxxL1TEOaBus7Zxwp4XPXb1lUrcYqsudTnOMW
y5k6JNI5TZKKSC9h4QBmP3zYpKTu6v4F+JdmCehFQ3IydcJJ9h9BMdU6xZR0OiP8gUB5ywFRCi7F
LxLmY1c0ShchrnKXTYyonHl/JNeubANvF1B6p4+3UI+sBzE9DuV5cf0pmkH6+hSRfR8Z5Uh6VfHD
K7QSdeatZaledhG5FPaDTp2jqX1Un8sARzcYDRR44kji0U/RmhegrpyMFWAvhKJsxXLCzw0G5Z/h
Y4ro2plVPfe/eLjst7+zX5qRAMzQDtjMLVMjSqCVruuxMSjOdEHUIl2e0gS40mfYOc+fmaTSoA//
Jnar+JtnXmABlfZ84aCzcgbJTdPDXJ75hULB1jLLmKKA29otiUZv/UtaV2sURtoBPwhLNwYfZYPj
zMKwzY9w+U5c8TW+HLCB5RYNbVstcLcATpq6KZMBthEWLGhw8QdV3eXI1WFVq8UCqjd5CLFqqPOh
RKtEYmTHkmxpY/zYkc0hAjRJ+RzBXX74NhFx4xdRj7ADoXrLZwGTkiWF9C96x8jph5zhdqOC32jk
B0nkuar6S5uegHg5zF9waRfP6Hv1z1SCTaEa3SPk5T/YHYutojtLJGDlZ8tnx8EPsdv9+KfjZrjs
sRsh8awkfnZAUgEp56+4DgBGs3jZrD9rK3Egqb58DUREPl6DhY5JjST2OQl1WEaC0MIjHbyBEu55
J2M/KxL+Wkax7hMhFtN9IpZBK5EoTK+nrL0ziPvOgI6Y/a7vPzepr0PO97jAUOk05zLfyRXXc8Lm
QDS3nrEbTImB0r8Qo4Q/5WkoqyoFMPpF17T6eLlxV07MOEt0mjAe3uHLnz+pBXfwPCT1vwormwUx
CwpwIvpqdX32UxWpek+g6JMCn3eTUb0DX36Gjzpf2uwgfpRLi9/jroelA3WjhQQfopBs1WV6iw8e
km+KWEcgj8FNQ4UFczQLFDvmUcKflZ/rPzAZ88x1ESVX10nTjQLQEmEKtePc9gBXZ4UCIZXDbUAS
Sw5UMhjyxf7O+px4JaDyaTFZq3YyPhhvkY6ny1y9Tm53vt+7ocr5Rybg5M0W7M4iTDtiKk3OnrsD
6lfjwxg29tawbCkH3OJGD1yeeHwCC430tBNy+ee1HchpQQ180AD/S6CCtMosRRCeSDZIv+6zIi8Y
GXPRwhKjDWF1xUx68JL19tJwCVjk33DtUIQbQ8JT3f2gHYtC9U4S5+VOQQX9/Q6u2Bc/H2I5JxOc
0OhGYjs9G97r054559nzRyWogecqZ1dDLdCf9mQilF+Fw2UGuhZmjBn6xxzCVmjnHuRx8TemWMfN
LoF5FbH1BNe7a+cIljaIb9mThlkuPPLihukc/te1nU256AzfRNKlcJ434SpZofjHgPbH0n+Q3Tgr
nImJDDqgQCwNaGOD7HpIQhdFbZqVteMJeqG/xRYgEol9wJBnz8lJKdtZpPUnVcfqhRehUbIZWR2B
u1Zsx9MDJyWHBdpb7qu7OC77zlYDvapxDCh5ej9hyaHmcJ/sbMxTyFLtm0CRwdGFZFwH7oQ372c3
lCHGyqc2xIrsoSSu6DGwsKmqQ0cwg4OFlUmfGP78kTP7PDP9dZAznaFrHv/MMm5lctkWzt+OeNk2
6kD5CVU9kXEn47/MGGaIIDEKqnCVL5rpdnSHNZBOb3pFGIKJ/ypqZ6U89gvsJOWLgUAGYYJ4hJFC
P+TqoBCXZ/cM4OW7ll8EJqWq267KOYm+gshCj2IN9/on+v31kPhX8Usw9FgKp0vXIO7v46VVLbfh
42i7jqASjTyvl2vOLKxp5HksGT70YP00cIasE6Qb7v6jedmn6u/6hvUWjdAA35bG/kmEteAfIMC4
FuRtALI3BQAcAWHyMtxzArEBubfG/8ACf6PvF8XHz37bvu6AnvZ3pGlOwil2rKZYlwQIXseKZ5Jr
sutIS0bx+zLd8mMHhHeq3BCd10UTlaCB6uiM8CsbYW+Bkfhn0XTHrlYigybiZi/ryr+YDzLvDZRO
z4yiZnXEZhtxeaYsr6nIKkAmUmJ0dCq5JqfLQyBbsgObv6dPdMAmaJcM8/1iZUKm7HjlCK4N3ei4
hePSp7Chv3A6gtBsu5VTNN3lwoqaQ2PofcsV0e/FwTTiBcQZhcKJGck10K3yJNorLz1Ih3ujT6In
szR+2fIrtZZWx6yFwLWakaQiUV0y16HeLhkPXdtHKunvzYv6SvyQR0OfXv3AdE1Q8M3u6xcP68k+
N2mRLQmsAxpO3hy3g27XZy6lRHVB7V87IRUiiFx1uvqVsyUqhIhDPHBZKe3vy0QCJ4tc11XO3IMQ
tQ2iSrnXkeQp5uPN6Vz4YDhSQxMI1K4bfFJpET7V1eqacHppHNReCMRo7OfEaXBOG9JHstS2n4L0
SquarqogrcVUVp7QC1CfcA5Lxk23ufeoJBN46blPTBhDlHma9GhSMEWVACkVqmd5a7XyZUy1nSaG
sU/xIPMD5I1zAYPiOB25yZhZqLB5T8kV6MUMF6R+G0Q9oYmL2r80mVe2AJSLcY1tepwkFCRY0oXL
KkLG5G1XFPaBKWs/uCxURZeQZHleCOcmcjmF37xXHsySzdLI7lUmHEDPrmEHEsiPlvLXO0ULeeda
8V20COPC87NbU+tX6qQ0E5MNB4Ju/U6vhnhnUYDaXv1w4lTYfWthI+NKsq8j7zOXPsWp+xGgrQlE
Cf8/5nIdo/Mn5cesir8xDuQGz08SKL3ys9/aEl0a1lGohNGEvMJBF0WLI6CKHM9o+UzMZmfXEz+F
/KdIpqmKsPlTlBhrPoLq2wz3QA+GuKteZ0vkWrsNvCttPX8jFEXmF/vV7GhYQVXXc1z4NCMFQlJV
GReNgOt0M4hoXCz+s05RGZFW4c7za93IW84CFsS38W3PbpNzTOgRiFamfQGHyMToNh3gFfjkZH+P
rMIhcZ2+R1PjGCq2DmyCwlJEi0FsqZMrz7KEbrZ85qWEssHBuFeNMymPFjJTlZgAmdpo1XA2Z6DU
Tf541+DKJ30arFC2GZAkUa7BYYlfGzP4/TT4ZiCHtUgWy8iLutPf4uBWabjH90p/JwMj0w9uWIzW
SaEinQPcFABENCc7ynrjE0Ak0yfQC+2Gc3AJTgjhzWqKcQfG+2SAB+YMWsCjLWDitHCRY3B/+vY7
g7yxsaS46CdJOAKNA0RuXwgNMjudcVdg8lJ9JsxQURIFTDaACzhnRp8lDod53hMaXeQOMProMAM/
0Ai7mXVkflE4pqOFQqMkMGVgh0nCQm5mpnLgOQIF5G3tUHqlzpSqySHw5KwsnYowWy7VszcBx9vf
qwenqU2Q9mNXnCufpMUfe5/BAr8Rn7fPWWO0jYOJsjoGRuchKVWwWhxI/Jj7CssPKozfJeXIpvib
RD03iYykbHk3OxS365nhN4OBQqaBRE/omFxwEUIr8bZKQ9im+P3WRNftXPyuPIEW6B4a9/zWTCaE
NRuoXFQM/v5cgv32Q1qr30C2/zt4/ma/8Y9TnwBZC5jMNHRk3MfDCCVnlirKKx/rhNOQIw0MORcf
TO8FuCjJNccZIVaxG/eJ8EKX6BWAvYiOumreVw5gYNseQQ4M3I/+Ep6mhw55mvuFxL3WYq28dz+k
WSRERzGXQtbHWaiv/0kp7NQFY7me0INB5RCT5tsgKcuhmaRwdpcAnw9MRqjvM+0tSUDVVUzhrSQV
D2SDFxjo4YAXMmfP/XvAA35xGFVepfbKgx5QTwzO5NZm03Om5mNnuq1CtmfrMlIaED1xTpKroimT
x+sdHgsH0eRoSXcYHmlKIqnQnor+9ZznJu6KrTHyCL7pyfApzl2bXSfhCHbOCHo8Y43FYvLcYnzC
wQgR7xiz8pjzriNFdulDpEitJ5OorcvAkc+d0JQrYf+ISqvncDxf1PfkqoFKWnHBPmcF6h7HMVBK
NFet5+Z8ODbeYdJBhcpxbRsMpUu8rPJXEyMkNyS1Plfhm4wVsQPA5lxJ7+hkJp/vEt1Eejld/XKO
PsFiugmdLxpnVZMN0DAHqIb13+JK+zcnVcRiUPWWtJbjtnTOjCUgouZT+l/Ew3XZQrChIIwOQX9y
BLvotSDeEEQKk0aSJWDeFFqtkUMq5I1MkPIH9GQw7/4oO6/qxMr3rKKcsEo9i+Hk0i+BAaQfrm0g
8t1BG65Fq771qmjT/akNnJty2sJPI9sYuWjTeOR2HmvyfknLMOH5De5wd8OA36aDQhfsgy8CHTdU
XaEZl4vK5UMy2Ov1HmHc0FMINN0A6TxlKpEEQB9oDz8haC1Co4oVjGtOGMT3S0YmaAzjgQxbtagG
MLYPKX4fZACWCRUgX6htSlasTKNf5wJ8fZ0RS4Cy+qluPGYqg3tjVF8/Yp+mWf43B0zt6Bmsvh0V
qVBAgIM72xkWsTp/75exp8BSqLzXj9jQwkKRVaX+aBZ8bvlSxoDjC4j3l4dT1UsgA7eXEn4cmeCb
kzxZINqiuThbC4m8bQF2F7izXo6jaZmVR4gGQGaP/BV4ybTOENF5KR9wOwdwkx1jguA+x5u7idbj
/CNCliZVD1d68tyv3eHGJytF/9WlWFJbaT/FeT0NxdhQaH3f/NvQhG8uJ1/X5tyC2OrZy3HDyrcZ
hgkuTvLqxihQfuXkstRwSg+Rd/vFzB4EGx65cLNKq1cvVLnemZRI2cGn/wWhcd1EuEF9IZ2zgyy5
SXn+JECWfx/Ws2UXGYfPyx0o+VTyNq3hh12AukJYpP3TsbCUxGu5RwVyArLM1pcDoJ5mi0NwkgW/
sp56tTEa+/GzH5WzmLh1DRfNG4i/TLl5TsAHjoYXw6WFPkgyLuzQOPlf7NwsLXOxT9baJSpcxPSX
FcMoUS0lk7W7PA4pFzxrsE+lzFZYmXF1Iqpm1tOOHJegqDhyTBn5irokyQWQmk+Et1zUSAbjAOBi
vDHPa7GiL+GbMaQgK31J3POHiGk+egHLzGU/7TIrjJkSPRe90NdJW8aRRTeZP4lsSd/4wnyLjhnp
6cvKxuzxDKVO/8PIilG+3tUo7ydT2ETM+bwRw833bzkriXaAL1LXypXZJ8Ol+kyIyTVFj80GNygC
L3T591CmYPo5bosb05MJOY0J/xeMkFpP+aCrh7DO7bNIhF6xZpAzvVcEhyq2HzXwWLP64jEY9Hnv
vkT6oGWsqfODUe8fIAT7YRs2RTvrXTccoVfd+YEnU8bPSWRVrgOoi98FlM4dMpVNWecF+dz/XzG0
F1w8lCiodYRFMs0haJ19+/7WW/0w9Lg/pEWH6FWYs5BTk7Wsqsq9a6DMn3esevTgFLRTVxCrDrTH
H3NizoKSMDZjN0hPSm0mbiYlVUDh0gTrfvMGvQmQaqTxO5KM1lqLZeGjFd2kM6CaB8WGpKf/IxQh
g17ovbe8xCtkdiH7rVsyCZ3KXWc3DSgekzM+BPworVIa8hwt9yGdfeC4DwmLkKvXmugR2HBZrde4
daGY79B8F00bMvF9Hf+y8HX3lSaaj9JUlDtghX7R3f4+wH4RD/+SaR4C5K8anxyzEw8qBbg5DNY9
o1OsTKmz8Hlkl+RDKHIdDDlLM55d0+kSrr46cznc2gvkI3YhcYXZVeI/TRyp+6Iwj6cUDKemTM7Y
3jigCSOIzjt0frCFmZ4D/r+s8qDHAPQovFOKlkRVD9/0JADpuhLL/VVNhrS0ZX7+r+s4VqQcAzAC
wVyRDkYN75u+WrOa99JulFeOrGdcE1P6hstgTidjDevPrgp2BkKRNh0Mj6DX3mkf3ONyuS+XL5SQ
dnC8jnPNueyStI9hUd07uPqz+fUfIfPrO7VDBlSz8LJ2FuabjWfVA8MXLde0kADQAiZ3XB1+z1pV
22u03fCXL7lf+Q0F8OHx4qAaZBMlIWOvmXvwq1BUxaseR3bqPYSlH6NY4KAildHYTIMVJ3LL/y26
eZSG3aW/AInbg6zINCeeYtDh87T08ms2YUVuyxaNlWH5UwJkHP1YjWOq6UsbA68taHBhinrNOcS+
9XYfI57FGIAoaJHIb8cGNgG1Tc4ItRkUPXI7/FiLTbALyqdHtmznY9PxCtNdBTP67+PyJySAs69d
HeRvRT8E7Am1mU1ehoMNHuz40QVIXte1v3axjiqaLlq1vAjqC4fJ9vzkRYtzcO1MfWlA4wzasVWF
NRpmf/Ri4UnupcvRE7+t7PdnM/r6+4EAQXATmjWrnronmU66blWeFXS9VyHd4WWv2xNxDKNrxkqJ
Ga0tJPsul6VWdGVlw81rfxp/UUFBSZsnTlZShLLACoDWKVRKdId0XyCCS7ZXG+k8clsciLCdwamb
mHAYCd2xLFPdpdPHOhhFwbo5LhFRAemJeSeV/6EgAeZKJFYfvOdFYbkyJpEeFQYGnFG+G6uv+S2C
wMWF+zbeg5/3T5nD/gmVnYGBj7YOXyKkTxliSh0LG8rHtWBxOMRmi2rxOPbQxCPBe5JFoPQAwZAn
ySxi0pCIHOw6J9FEJoTi5WR+8HnK5cBDpX9ax56AVCc1MA9I+1ohZHk/oghiYo5I3OXPFD2LU6z0
Aejin59ndmJ5P1yvFuIwIGAOmed9lQwlJ5Dmab+gOYMWl5yXyMLPKOdX4u9HuPe5B6yIRyTiwitU
Y2m8mXoJztVHgI7lbmJZp1ZTjWvQ9YTjatbHUCjM0+oG+QSpn46HXJxRW/3qSTbYgi8lzYOg5iQN
69giaiRI20zH0olT5MgrKYtKpzXILrX47dFgtXcODzciPqv9rdr0RjYRI0dqGtcAEiW1B6n9/YXc
lm4Y6IYuez0QvPyyEuq64tqDIDZpjj0bRswmckYXk8Cg9UoUgDR2t3GOGY0L/m2gaT8X8938slwZ
kqwt7YjMY8298TsKdp445+tkRDxoNC9R1Zhj1wvhkEhnOSk7S5aoMCNxLjVhmUWEJlkwcAL6N0JC
j4snubxJ+UhyVsWZ83+Q06rlJeLnNkkR/FHcN6+HFoiwQpi3hRhbOgqr7Nkxb7gEH0NgwOWAFDlG
lubpbn4/di+A5D/7f81tUkDkwRoSr1hybogBpnYz0trgWYvqFhUhs7/lSVokxzVRyPvOKpOFQZbg
zLaHkG36/S4XYR6h8LbWsZX7OHhxyefJe3EOGgLM1XbHaydYpzHxL+hJpJCaQQiMRMuWQldIG/ER
E0Zi5LQFlUR+NXu8lf+qazDJhO+nop5ON447ox7tAi/ZuLomCERjkCUHY7jrpb/XSSuA3mROPkdX
ITrlKkm26SZ4PKFmdliw3FpuxeT9nDLSWTR8vCMxF5Xbh5bglUCSV0k5IY5KZrtVk8IJLoXwP4gT
9h7MGuAtWxotaMZMEJK0OAah4CWC1iKa9lgiR6Ey4F5j8hzWpaUHW9bghuag8q7tUosAiQGags5V
JRWJ8DcQUu3mDh8zGxBcY0u97h63EujI9tPjmd+fJY8dPE9GL73fAuCes6DichpFsCf4uFcpTLPq
NiYuSbckegkQ23b0ByzukZyQ+JxuRERPl2usv42xBB2xLDaDy6BcFFS+0sJZk5GWl2arJe+JE61m
FYEkzAYEXRBbkpTcNXV7BWMn/scEctD8vAXoz/M5KNW5hx6x26GaOF86VqdvINevzi8LtM//WPvE
oElKzR7Vlayh6ZflmUFPf8CIoyE1iPyT4YbqeVeXG7A2D0YhE7ailtpHsxFxlUcPwTlo65rrRRhn
6eYtt8bdBjGa/KPO26DARePZI1lmsWMuMZGQfB7AFJm95p6Wy5iOmJGN9l+DKqvrlksvAafQi+FL
ovPUGLmFM72FApV3Ot75shL7P74VsrvTPdAm2d2e5T4M2F4wVHHm8vKgeJMcgq0IgxgIqMPohl4C
+xLRT5kbtrUY4NuE0gbv/dsOVbGBRWvWiDnlfFzbgrREDCLvq0UcoKSEhGjNJXMtj47UYpD9znHq
EkTvnY6E9LKyQdhhzU218Ow0QY25r0njvAEKnBj+Pfo9MB50pBh0httjyp7vE5e0K/Gf2RJmVMJC
eapPJIWIPtR8diTjaizvKP5se2gOilT+bwqc1R4cYMInmJSrSLrl3GED58or+K0ymCrcpkTbN10K
3z28kiVq3qOkRGHPlPjDaPkAq2eczS3KDAP7RjvDHmctODIPnruxf32BFjxDG/krsfoneiBMdodO
n7BST8jWKnq6znruD1493jc2aFUUbycJYYuVmis90GvAn2SqvJdf5l59ZaT9fJexZLiEHZW/UND6
0y0aIsNeLKDMaGTnDGuFz0/0DJEY3OhGiCBSbC8ur7H/Rnaq67JsK4EaUeEiVlNFOxFp/7XkBS7m
lRJB+0KZR3PVPYogj7Dmaw0qjtqCux5mxick6bBePxv4sl6Yn/9jy02HDvo87pIGd9WDXbcZ/4sa
7Y0Q1FxnFK4wv0D8EKyP5x4swcCBvRXsYS77UGw0ws4riDTwZmCn7ys4kcf5lKjG5IDc2PCY5V3u
oLuBzY1RCxpzccCg4BDT9PmM1mREqOYIxM/U8g8XRsL3vpgjsdm1QJERsZ8xK4WtltKLeRYxHX4y
eoCfbzFfMheB0Ml1jUP5RV36ZucUj67skzPJ/kINi4XDrgF/l1h0WZ5Q782YyqC7hVxqnlxjIS7D
GlRkR97mXaAq2MhPf0qyZKem+SImoiuYnm0QZMo+ONcRMILTjHBQPTuP8PyaUq0aVbXgaSeKgCIh
NkQ9jcPG5dKHpbhNJPeLmTcEGWg1CGVgZ1YpiboxL9gthwpSmTai5ydTYIZug5G+RdUaLedUeK95
IpAD2JIQ4a5EtCjO1QJXuIv6eXZUGDBrTfu5OGfzYwJZSfPV66DCpn7UNPCAR2AfB9D9qv4aRe4P
ChX1lBxLVj6jotnB0YmjEZ8jmoDbpgkP4LDgIljY0sNecnIo2hYOuECjIntjkK4strMlvqbfYMZk
kN/+C9LwB2u0k81BgOEPOn9k8atRSeersct8kn5QSuwnZCagycFyf/P8/68zQ9x9wkQ+GPbAFfJF
OnYTYTnpwPs2NTGt1dYC/KNUBh404E4FtDRiTQTw0UpwEFaypxKJvZWNxlTD8MMz4qkYeuJqowYJ
Ds+k+Wk2CTTU0/vMlC0m/5Pv4W3deDQa5taGjMzwS90Ru5CMJFPhQR6mKwFvsQYOvRA0SrmTIanq
JVpdglIcxpTe0lBUoBAfC6bPtjkBIz4Q0Q33emvnrnjKFrFrl4k1jFVAeBkBPsFZ8x8OsPRFDoGf
AfxYcX1C9Uh1NDhvNEDU5Wh2gfnZTb21xIehvRKD5OB3CBYaesBIEuCTKoI1+w05DqDl4E8M3wY5
tkIBtz1Xwh9+qbxcLFWCcK7cJt8gRPj2kbvUtje49jCMIOr8oECtqCrnYkKW1q60v2khzf7nN0QQ
F6VWXTeo5aW8ZGVCUMNfY8yFeifwol4Ysc8SAK2dPoWH1tAaG2A/A6mUX3x3EG6ksfV7vZ5IgStO
3AZBEGSXZ4GAt5n4I3zY/4oG6Lgxpgr0Jca2+yLoTwvRbMRF97LPfPhmTJ8Ax/nq4Ge4e+aOyWmm
ufReUf9GNpeBkUrJHaHYbEXCdBi21R4D4b9XE7FlUQ+CHYgt3LnCqEcUmWns+c6g0VrSIDNFPtB0
M5yOfZNFH3V8GjMdfgwrTwI3fLK1NkfGlMiNIozChLAK6vI/44J/+LqgpgofNMraZYxNPl+s0m9F
OgbIdwSLNI8usNSn5DJyfQhVfHHKhUMldcFGngEMCRSWZI+0g5K8sMlhK5DYUpaHOd8I5tmaxIjc
QIw/nI6bJ63KA96Lc68fM7yMe0sHhBL520aobjxJ3TdZbzIwCXmTwS8g2ziuxaqla8wHWFUmlgGu
TnjQGunp49JKUbnfA1860RgBZBNrjoAT0qEhu81nqfTIOjSJEp1FjpLGFvJWPTrUbeB58V2nXCU+
NfcmEqGSKwPnO3qpmjOx/d7wAKq+7+qD581hCpOP1L7IGrTkdbbpxGzN5RnvWFTtG8uwj1DQb/DY
NBRUmV8J2E9RSQ7K+UtLL5toFP2wBKi+ilN2SHLUfGZUuGvucyF299wr6QjwOpuyBrgRkqLoD37x
ezUpsiT1UrDhDQhRtj2NHHqLx/TRo33sYGeKl/OYnQ/7OsfROqAizAoaCirbDrcq7LEMHraCzqiG
aUbG9hLbauQKrw1Iec1IAw/KAFRilXMc0ZkSp7Er8e4fI0CjXANGjgT9LqwyKxDknjcVcPepCjjz
lQndaYjrgEeWFhPad64LZtKNhFyBLqX9veqJd4kA26PT5ZMwfc0sgPLjiOyJWTbrAizgjOTn6dmv
GEhMt8G4M1nP6md61lT5MYukAseif4Rqt1FF6g6svWM/rfmRa6mp3n7C7N7j8oOlwPg+qleFabLY
kD/ueHswC+lBmhN7rt/T0KbNQebZAqB2FRzRXHIBS+uyxf5yX7AufwnwLFrDCEKAj5wqoE/aXJJB
jV1IpB2PwHosTzZh9H/WI4JwyYrw8tDCKQGTkG5N+aMeFzGYMmh5o+OTKVnmyyg8G6n5aGbJMKM8
rg+B/cIEOWm1Kgrotz4XJeWtry/byigGXwSeejSpteD1Wue9DU10qDdGWM6geLxiompgI9HwwbXf
ZDTwMmqoakjV1b+dBmL+PiJb2A5Bkay4ZqJCEYsTeaWpBfgPBsePkw4PqOtcrg/UQwIsgWuOSfDY
e9bAHss4OknLP05iPsNr1QknKZ8BM5c5s9De/zufsL7Et7nUBgz2iGezFz0CfEPCX2Jmi0lbJ9Q5
9npMKKtv08CRKfbc56AdWjbUOKUhVyhe/fE2iyvAP+Ufw1ER+Y3eDwOUIFjuVP8d9435cbdo+nl9
6Dl9SG7MDwbxbUzJzNlzsNL/dNLDJh1XxOBtE8+OXX3c1YM1Fr69bPJtj3/QYLH2nEbEavagTcQb
JJeY8JwD2O6Xic2I8DhaYKtlP4QaY8QZ/cvQanDtCNVXF2jXZM6vYwWLY1OBCNXZfdRbGNtUg2vI
fuWqkGG4tgRzYVfgZm0PhDM+r6cPQnWBEIdPd0xalO2a+Jp1yPD+3A7GjqsFGZw3kzYfdYpDuz20
kj0M6GAYOsyIEXXAIzG88cUavV3YbzdUzn/LMrb45X9d7/EE8p/ynT66b1Krx6yd/c/G98926PZ6
M8FlnFdKpeget755xG3Ozcnvdd9InIUzazAhXgM646cpDd8uUfZG5q+/Kai25uz5sKtt7/AFsrf7
dVk7ZKodDB4/58O5Uo8sfhy56LtNwBIaQf5S5i4n0xmvCnqKeMXkCvEwNqq4YUFh8VTQMKok/4I1
/TnEKu2baImedAKb11DvC7u38ndYMFkfDWMgdeIYGhd6ZhRn8PTKr3OLeeOUQ7UpzjSJnGhlvBQ/
lIdEHmWyUlfn6JGAxdG4z5g2TLn1tyPk39v3oLsxVrBviGwT+/Bcr3xxznPXwExVHykzDO7OUVNs
Gz4rryyqwZY5soAc9KUDQrexcJq6o7A3gUFNCH25V3hu7UgdatBtuDd8ttYyGERJDhnjhzq/d/xp
3XizNMvFU3n5l0pggK7OTtEu8DZMN3mUllu0TEqbYYOKlOjTB9OlK9WKOOXVBa6InbYb2TFBBj0t
cKA9vKCdgqVRw8ikHSraEN+AtsgujdNE0Txw8HM5jhNEJCfhpBWvrKEbrVBUQgldDeJX/IbKQlYh
rU4goka7sTfG+laeJLZ6QvejP6djP9xR59/jEOww7yaWqLYfYH0mVdh7QywZx/Kf6+TzNqH0VWRi
0/ht6Y7FDqPRpnGWPoN44JDNcx9yXT7xmXlPTRgmLdNQfK/huIPB6sqquXfPe2wY7NnAW/gQ3sqo
tAj4sHfiX5JTuLOtfQG3MvgmDynx6CNQi/vV4Kuvmq0W1FBQ1jrcc3+jbeFAZs4kx3u1JPYucymt
8mgl7jqFK6GXUNjLq1/F4ykka+IPQX5ocPoxuWM3leqLleHA0Gza8KgDYE7MtlUUwQjuC3iT8H29
gCFvDwB9Ge8TMCNJS9L+0wuzIOhFrFVsfNmqxCAffq3mzWvV5GZ3CzkiF1HlQfisozDYNtEHKBl/
z7O3xD8uvxRE8gq9eYW1wCW8S9ioIpGmtcEYKLLv4zvBLN1UOV8b/XeeA4t+x8I2e/RjYSk7889C
41emwdJFnQEdftHPYedAJ64nkbCsEf8rVwpQMTaAYSAMGD8c8z6507xd1+E/vtyHFLr6AFeFaEVk
7aBTZLXnt3B5Hd8gijwNrZIn6As6i9JVBmc6XVEuzBbKeH8F+cq+6tXBfcEtMqvrEkCnlva3t9jO
kqWPeJVHjdQJ7nTITXYHQWG9okP8WgtxPG5Q4GuCMLp66r2m/uP7fHqMMoGlsub9+pja9AUaN0Kw
SxbyGgh18xN99fwIICXgbzIZOGuZsr3nkyk7p8h8A/TZ2EEs7fmEr2SwVC7gtq6x843ZvO3qA9qR
gKLudrSPFSWMxye5mkAYZ6h1BSJVBGjXJ0XZ7adaG/wGIiP8pHCyDSDx+93od5wF/dg0RJeE4Y78
cinmg5jYT14Q9m1ZzCY9K6C/p7qiWeVYX4CDypBZE+2GV6pn6m8po+HtHaETveoj4JMWB7lJLQkb
Q4876WuIb7/zy/tIpN3o92RMOCtDnj6JmN4/SeUHLOm7oeKfwCTGh6Fj9Dh1PfgwOEVX9nnPMEdR
Hrkqqw/MqNTTnR/e5lyl73ctjKbhrvTuI3JPAmcbzPtNlregOq6Ys/ARwAP4liPT/B8imJp8bOo3
lJbuUgrKhkOu+D5Zjo+CX05I1NcuwWFbEc82dDEAO7+JV2PZ6/yNsPpRLQ0eWsB3vvPjoSLQudgR
qQ7hojM163q/pr7AC7VWJmRxoOxAcv55gxmCJtu+SXSYPC4KxNenNjQ07QYHc5mOSJBVitsuzFkP
YeQxakF+kcAeF2+RoWg1SYElksxlYOQOo/CK7S3N1zg5GBb/pMyW7kIXsM+QOHvLTNgMmfi8QqcU
fxhPz+q7FHbrFcKgpR9EmxnEArLKaDTN8xKwdoGVte6paJ1mEJfVyu0QERMGPMeCXe7kGylIBiEI
SK0SyITto69kNVPBSZdv4w67YafjUfXsdAzrRHX8ce3ZOukF6dzs6lNA12Civr0RPLhhq7Hy8naX
HIU8UED64wyDeF4ssK/xlT7djL47TdorpR5s4e1JOBWEhQNC8/aIJf2MGnbYIXNtl2rtFYpAsEZW
MNkCgDiWZL6RoN6TwqLbNeG9tC0GB9UC91EUxIBOFfs1CYadWMNQglx+hUh8kGBZao4MUw1SY5rX
0/J2jo5Vodz35QAMuhAFFQjPhzr7zVm4bZtMj9CJyCTVgGLqFwT+L0Md74ol0jws4/puIz6j1C2m
qSBv1DhHc1OiMPdu21I2eF/fHQ8lg1QBdc2MlApGQ+fwfFgWW3bzUE1W9R/pc/ZVJT9KwaZL+m70
1FHhgSmBoySYTDKlVXfJ7b7m5NmS1OVFKMoo3H6ziXuBxrbzNvP5xDTdtWdnH+1ymmmjzo/KvsFY
ha61mQBSf4/pKvsNEO3aBF4xe/EcI6GWj7EtWVHrch6M2ZugqBokVuHE8LQUlXmjDWN5JT31/oFn
tG8GANpoGbFG9U7z0AElq62zK6oQIksnVtRubNKHOFlIbrAV3PUEDg/QOqKL5MTaZgHLs6Ckdopy
VWyT4h6lfUHRpWnxX1fSZJF1Z7z1cQI46A9aclpuoaPB80peO4n/+73LyPSBdMvaPKkWdl0EWRGx
OdjbCubE9qGL62m/vwgHgz0b1gNb/t6Hm6Y5n0jptDRRWtdBMC63PGWXxsTZei8siHmviGh9wpg7
AVjA6N1EzPplZd3bVMVs+yc1xYP2bHKhjH6SOR1c49JlDqzfT6Lw4sHy9fV2souWtp85PYNVl/2J
rinXUuudYK/sZK8s1a/eoDJ7VdTVqPTDgSuMRviwrMh0Dywf96FniTsOzFOvJbxxkNE5OvK+iwKQ
yKbSiLnPNx+vqBxYOGtYT4I2oIwtj6P3XtHsog61iPGfA+9KkCwuYw5I1XQGgjcU8CWZKWZ7Jot2
gRKxH49iVZsJ2Rhd77oLv5zjNBLUr/fm51YLp7nmKsmPliQIpd8oHsVsjlB0gNSfqLGmmGhsOC6y
UIwtYj2GC+0U69kiD5T4xt4fDFRLR5k/Au9otT/TiRpmlc+rxdYgp7BlKakHoz3p6GxPcx4d6dd2
RQ33lWxo3n5NqGqiSlT68mml3w3wN2S+JNwYcXCqpuccGLPVyrtXWk+Tr3Tr08F5ZzKGBBWO7v4m
umIYgFka+48NTMSGcv0ntLNVQkTOBHQlT7qyrvYlAA8Mm7J5Lg4cbCr2SUz2t+5reoVJ9ZXXJfdc
Z70SokZDDalAMsTY4NM9jXaAv3lTFCRssJ3FVqdD/ik419stnFAcZvMW62ZV40IHit7sS2UVOVOb
aF/M1DKhlNHWLuxYY/zGuqBzEAe8/uG/zQ3Zu4AQgR+qgQ7lzPT2m/9nwo5H4qUCz8kYi9e02xD4
AlzA3Xv4qnaYDb/QE9lbPbDlNOE63sNA5j4mfntgU0OVbpUTK/FcUgn+cRYBU84IL3joxjtHsRi9
Bf/GqiW2frjf/3YzQDGmuW+zFubm5Typo2yjYHnwpip7YlwVbJkXfUoEw3WaDcQAicMgdCDUwXyW
OL75s9Oz8pqKAltZaVMl883ogZByK1MvfIwc42wZ/ILbLUxXbig3kLnF5GUg4kl33Ka78REaWeZy
767pk8q/UNgCHowXOtWNJ66lOu7OtBesrcZME4H6Y/CEyic5UFVM6G6pi0k2JG68WtGIFWlVrcOe
P0vooqVoUM3S3Ldb6VBMud+t9vkD+3nEd4FJme8nDRf+DJUKeCQgHdHgkrPONG3Tla/p8PNMf636
GH5JhbRp6PIxhHj6TZDdnP6qdWt1TLjtGtDQMhaSDxLq4sqgAPTpPbelohjN/L37VS86Amgfk4KP
q9h2LAiHUT4IugtVwKFlFXKc704j+aeOjk+Vx4TGi7Yfei5dIN/dO8tdmrkxpKo2yFpw3aa3rAbl
ZXqqIfMWiJSc4GG35xFQ1Kh12enZGuWMBCvnSFhHLGLb60Vu/Do00pCZksVNsHt4lXDlwCig5prk
o/tn4cxaVFLH6mc88wBVAGMEz5mLd5FxkZEDqRdMhjJEEdboQCqxOJUbyFKuVJlRBUPItexFCIl1
3Kt022pCAu0ZRgBF6SbPp6ySaJqQgvUblne6/mevLrZok68E6luqL7cK2KrPQmGRruiPMcmw13Oh
bgpHsJFLjH30XRet6dh+fIr8bIjo3fTIU0ccDy30hcyyit0MtxRBtqahiQWnEtdBCNL+VTaXboKn
SIEUpps4OpBG+2CSaMjJJdipcp2Z+Zt8tK2s4w4NoiK55LNKxvBb+j9U6Kh/Zvme0EhiVkN4gZjc
OChefs1/sghaRFSCsJ98EuuzNDH+kW8390xLKFFZcXugNE70pim78NhgcJUGkxfgFs6aFkeUlz2/
vwvEN5efyfyWYQcFmPNay+1RLUD+BWEkLOyRUSXAVU6q33FknVzlETve0tnUiwyEx+286xKzRlSH
80DmzPEb7cjvpNTtTu3S3ywF6B6uFhK3Y6cFsVbuMM+r3YWOmdny3pO/nXuTyG+vvCDRoKwobJj/
YeJnZGMDsBLwjpyrjVgDgqfaWAsTPyf8ZVyT4BzqcqLU9A51FzEjVgdu2TlRlklgeKWrVYvCRMsh
lk04adH2wanlAhZNMW3f7qa8DxvbRATLyeqHJnMauVQ+M/Uj4SFmJf01gS2TUBN4lS//ozdXfgdu
hFOeq2A6UnxC2mU/MPhs673Xfnttx/D1ofFWHEx2CeOkKhd5Korkat3EUC/YGb837zp5g0njKA3W
jpkJ0nN1gSNjh+pSpxVaUzHih9cTblYdEDN7ke1KAvcI4jfI7t1nMjsb8qCf5Gaw15gOpACaWJ6j
ifW9cN6P4tA67LCe8+blTCy5KRs5IFJT90ATjO3ay9Lm/NgNsWzYKuD8PiE4EDC9aRLqg5k9pJyR
vsWFF07aPLoePFUH7uMibSlkc9GgrUgPE4ODEmZcQWrZr0rz1bhYsrOw1ZTShLRsiQBEu0bS9X5G
SxL3TdPddydY9PzKDDz49Tu4uVZldETkPYQlYRqg/j2ffiIyJSgH8/cgGcUs970DfoxVbPgBVm6i
usZ2MVQsBSUeUkAWRrvg6sNuvzjo9OSM7uqJP6VRlaX5KkwuG9ezeGyhFQxGNn6pk/IciasPbvz/
HVaEVFVfSbPeRhmPGwDaRzILG0rosNvlyr6qtR0XNu89J165KMDP5wC0h3jCuH2hPYWKHUKlbpBG
phaONUjYSUDSoWep2DjNjLlp4DxbvENiPoFgHrAlSG0YD0AYP1gRnRbBCJazN6ABazDSN6Buxy6W
86gDq90R0mW7kJpsb77C75FZy9BVCII6JoUcdCcz9Ot2S6R2sYw0gYLgsjGUigcXxeLAzx6OOq7t
rOCdul6wc2GZM6OAXnNIlweKb3h/IYV91IDETjPIPg6a1fh48bLjjEU8ouQFyx9xLVvHNl6Mada/
QXzPsfPscqhpthokd4nHSd4z9HyRcUP5YbmU/+obLiHYs1p3xmXzdvRwKcyPCRg2sD0jV9ISk+3U
7jrke/ogh0N378uxFZfLULsFXS47AK5rgOtuZxhA9keLjer7nSQTer8o/IRKb4cJk2GcjlOCcl1f
Tg5a76yJZ18uJ98KzETTjE46o/p2SKR7yddWEcCBLKorUdonuTNVyCqvxNrk2wAcqRIMhrsou5ET
zgS1BzILQMozQOfg5kDYH+r0Yqa3fCAZvMuqqpQ7gSdCDEvwyHB5LXrmFTqMRDKcTRbzQIaq0zgT
69dd5lDd8Rairh6gw3fEBrU53HAYUFG+/EmQf5oltfL42Gd46HQeTmjVa2lDniMcLw7/JjizpmLR
v8WQErYyPrCHJxpavvfEai8PabdRhhmVwN8/1U6vY4t4DR+vpWZwaWq2oNOVRj/keKwhqoQFyVpc
7t9PW2YMXrvFMhPKcsyyJPrZ3RnDKleZGok74yr/RmHbNyk5JNrHzKyq5l8g4d9qy7AKjsR/nIFw
dFt2EelSgQ3/TdTvAwWiU09t529kCoJ6Mzr0VCCEjkxm5BXklh7uMz+/44Gbl2D1o8URSn8wLyWr
Z3yOWey3eszLnK1wVIY7ra6u0MbkalLgNH0iX3RAQMbD4CScqaTO8vghMaFsLnabXUngmi01Z1Di
8BuE00lXy3ZAXL4S4Iz+3kOH9hyp+h0QlM+CoKvbMttiktjDkw6ugcPQYVxXMQvjGC2rgYNPSc1l
ghYo1Qy263I8jvHcKRqe3W4dNh7aJNgw5Zqurbbf0K+2q3rC1pc6YZQEaYcWIa9xe6UGU/tJHgKi
UNaOa1oYr87iEZNtfkShsMdH89V5QQ/IzFtLDxGg6SBQDvv8g6SecsAW+tTFC/RHdrCW1H6XXoa6
a88epW4S2G7FR6nvQGaViKSLMeNv4Ld6GaEanXMM6/Atvml40u9+1WVraMMZsf/EU5mVVe5zvB7e
jWCXaSCX84HfD0i2RbVMJyleLfjZu5M8ELzKbm9QWCy3jOg4yfLoIm0OQ2FE8O0mnscKmF1UhPVl
L8CTNFCq7e4iV6DdC+48KoTKD+By4yvlMOJByuWMHl2+yal4b7NZ12qF5vBdBRjdbQ98Ch6cE+//
XWkntSKCzUbTrTPstrP5xOW9WPkeeIFlkpiIMa/CLvvpy0DCsYHWQLXyl1kGlGz+xq/gElTFgKub
pFHbJVnAA0l5PMqGoLyEgWckdFtMZoJpvDlz6xOANZJdeZhAt7h3LOAoPFO9N+dDFSSHJ5Zbr/jp
Bs/BMsloiADs3rFzo308HwrIYz/v4WF1hVd/tXascbrNNYbd8UT2559pr3Nex+m7v52E9btpNrhj
3/zWl7H8ZZcmGuBkeGvCeMr8sBWZvYNdZFXhNhUPS1rJRSDsNh55JFQTpx89A6fYwaubz/AgBLnl
MkHVxgOpvxmEr/hWk+pKu8cCqxX6aEJQxeMG3QrScAWfsNWH3tBMqFmpN2om8Y1oCzxcGyN2a6GT
fSitXJvBOc4C+8CtX2T72UyNgU6seho1SWRhIWnJqCCqpMRrU2zzDN/jp1cJcnxdCpe3mZvnoNON
j7Y1LQN/y6SH3+TVuNGpOtv46Ympo+9MqTVskaUDJHYL/f6SXWmnm0psWLccYFQx2gc3zBDUZPnH
xh80gJxEYLQRXXB7P0HZxmDEZkFTnIKwOZCTyILx4aCziwgeyChXIJYud1fSsp6mIX6bMDl4XZfN
KniSbaxWAQBW9Mbur2kNxCAP1C/nqyTiS6BL4eEqy33AVr/nfUr1Xa2JbggHiE7LVCr2BlDGv5XV
yiEctOFdcYsCOHrH9BktcF1lCGjJ0+bEFv2vNsgmtti95l3d2oL7uq7kc81YRPj0lxvq8A3EC6Ni
nAtYv0EfKQZl3FU5M8dlM73ZgeLFBPhMgOoeOloxQDeVxHgPXVxYR/CZB+YJT5gOUnwmw3KxUkdJ
pBRlhcVmOC9M7ABFb7tlq23H8RGjaIH+0rwlQh3RaJAxwP+8hmWTHkFToEk9WgoWSuK5bUrWAMRS
Ays80MgLS9tMFlkPTm4CNOZ0jIyFyzj52v4KmrccP4bRfci3YDOce0o4UU/iYoO6LpKjnx+vrR9G
0mLPT0A+sigJbJq9B1dQPJUh/r2Zu7I3kdZRY9HZcILvtHHV4vLB544x7wEydHMRf+TZh3Sl3pE2
7M57EKiW0C+9UBUE+TKkFjVvCUhxScGDgD6A8IgXFNoYr0ao2Uohxtj01tXpYaMykrGLqeRdr3TG
Hbh7M2zFNQIzmtUaYm6Kt0rqLHE7anBhd4zSYlXGoGFDZxmj61pXCaYha7LsuSX07sCA8Nlcppce
k96Lk0/QZTQAC+jwObbTcWa8b8RKfiKHhjXr16pP4Kjaf82l+Xq8uQCE4vb/uqSgUlXFjrMa/U7b
u5rAgwA4Jyoo+150DiGhtpvM1qOhne1VILwpvYzOfQjNFpxVpVsSi48TZOWmAiGf/VH8QJBdoA+k
2GZX2W1JTPKXaVMX+EQgR1Qx6eeeb9VT/23WMnfiLIti83i2lDgsA9+7WBXAp5BoskYnJMCQ/mEw
Zk4dFbfLjJ2v7WtQIyvMetAi+jpXyhLRvmkR4dyE/OiH5txgd18EnzGpBYuo/MFIKcZ+97KCNm7e
PHWrMJYTvu7f6rdZ/P1CWe4hZA+32jQt4vGC+gfBqBSaWYlRo7Xe+iEWeW7s4tKOYuoJepTE8QDc
HOGUq/DS+c0Hgy8y3JDcdW/MyoVfUoXNzjY9x0UAk62sBAilzZ7riNE1t6R8E+7HGbs7nKQZ57D/
e42SYbJzDs/KmLDWjwHPoXfrUzf6Q5P9twJPr4CSwsiaehm/elHESldxc3tG6bYA07VCfoj11+Oo
BdZ+ZnaGVyRJuvVF5TreUzeG04ZvuYxiqkWN8QI8JXHoWeUXZhZn6am+cEBBmW3crAFHeCp5sbau
wcGGAqpj2lehUlLzWHNO7OhHVDKi8of5kZZ1cCRAqkiDXRjJzQOLU/K03w9xQ7FemgCpKwsCYSqj
zPzKkD0UwbfV5cOIWZJwF1EP+7XA6BzvBRKEF4XnmByJxgieCOd2hQezoTH4KF+Up9ezS9cu0a2f
TIvDMAPKo8TUEizJEtWA9TKAf0G9YCVp3ms70xtwfCR1pG2K9hhpx0PugtVbXgGIHrTRLHtx9tK2
1SjMumzjw/t9GP59KqZzUQfZdybCGsO9Fi1oNjb1SKLJytKKCLOr+YzRTISCdhelCsPAMfTJJFmT
rbzFDwKHLIAmOb1wBuMbphYEjlJQ3rV3CXc8dy3PyUxrU1zaq5QXNnpMm8hYXDGMdACWC2szyavD
3VdsqOJ1UNb8hUImiCuIIgivQOYoiuxvxNcre2YcMTY0DqeTNcfgV8h//R3ONY86weHiFnu4mG9r
CAd/gUIUotqgspByJUJ3CGh8YLVLcUts7kFabvXhBnzep78aTedHd+KJNI1w1F0zEPp6SCp4Wuad
NZP9DmS4xxGrTI+MT0kvG98oeVcJmxgYpB+8K/ivlylu19DNHda57c9YSfXvqnuEKGNOGh3w06ig
StUSAFL6j8iY5wZOuXXr54DW5L8yvh4WgFA3+kN0BbV0yY3IHA//35rCKBQYjFRAeQK/NLTo6G26
XNinz106Rl5RgRleJAeW25cUNA6ww4+I9CpqUpksIvMUFdFuXQCMaIJxM9Y+HOuKb5otFvIeoAeE
ZDFBhdyZ1PIOhanE/BQflvWGE+lIwpBHFedLoF7mA3qP8p/bzi8gOYsKCy6MspdjUd922q9/4JTe
4LYt8dlPqkDg5EGHtg7AtzbVT7iIRPchxJAU+nsPiwawYEeQRSpQ+Jab3Ejed+pIonvco4SR/pRN
jB+F1QWubJ/jpm1vo6jBmJIt+gDngxI6sShppYsglsWLqL5GyRMXfJbHrVnj/GBoVpJqvVJhJpVx
WkWA+wzzOWF1mw/W4PiRm/jJ9/caV922+Hgj30AZRwDEdP7LPPnfIFJIgpEPNDNmE+Jzdqrfuxx9
8gmPJb0tKgpHWq4KNDwF3tVzTXlp++mpYrr0SIJX4fJPPkMYMAGo4VOcSrYqkAbrl3h+1GaGeSF5
IT7xq5U/M8apm9lGK5baNXO8l3TYTre1UWUln8Q2kQwugS/qiM6OT96EDzZTaNL9iMbaKpFgTeX6
cvNmNKrNGPsgyRf+SfK1LYDZGT6mxF41HNWEgLOF5Jy5J9P1tod68Q/M6VW8PgIvLiKj9a7QiKNl
U2+muZ5jvnl68jb77aYrH+pwy6yvb7E/SyPnkpGwURmepixGBpK9Sb8RL5KqP1bC+1dFGvHGEY7s
JBo0eZbt9Zjig3jXZkfdCbtmInQMhbjh8laH0340Vrm29xgLIYpu2FNE77pK7G6o8FDBL5DAoKJX
3mzF9JCPJqYmdJ7l4MAYRiwAiNWNLNxY008RDnAQAnpV5yzsKn+fm36D5vF1Qryr9fqKcIpVzKKi
oUWmK5uTJ+ZOfLQd39GDX0MY2CfQLGyLBciVagV9agWRYeHsD9+Eje19H5muCDyqll8dnkb2waBY
ALGol2VecQttn3oTz74MIp0GVCsanwf/YhDiwyXj8j8qcl0tOVvt0P1vvhokGO9r8G2maA3PLJs5
Dbj8Alyp860aGipO4pZubK8cCDprtV5jLAilMH2QtCKHQ9iDdGGQJlQiMp6wi5p+hTHBYgvtu4g/
HxA0Hz9MHnKAYouTJaxXo29OYD8n0zZj4++r9/2AKDPfaDm7YMex4IMGD/hdjI+/MA+ULpXlIKMw
i9niXZVXRiZsokS/Xai4U4KlqfLWKzt09L0mtCFDbzYCrZnkbJCWpXf19XwTEz1P58okxWRRoN0o
OSsV5HEAjgk5oIJT3qe4WiD+rnONpQxksxWMqtZ1l5iT7wu4LhDdLDxJkAx2uZw6pv0K6o3467dQ
9mzitBqK3iYU6EuoLcB7UsDhK7arK9j6wBZkhGnr6XMS62mBkfBq1ATnPEhw4lq9faO4N+T9aHsF
mOEi9a+/vpAnlWbyVbWhPAEmZq/i8qq29/pFrkI8x3WlgM0Dc9a6XbLwtmqm6iZmkivimel7hzyr
IgK21twKbKauQ9GcliB/jz1dGT9vpe5lerMmUqQmkBXvctVJaZiBS3O4++QX5YjjWHfA0ubviuCH
z+jr69/z065QFJnFDtiJIaVw73d3X36+QocyixUOlqn6/wdgZUFPmxgi5JhQZWmf6DmJ1tJydrJq
h/N91LaykKR3FAL1+TlwirxtXD3SzR6YecbtUpoAI4og864idNh0ZSvWT4Z/pIOUncu1Ov4YQPlS
yCgHO0uqy+K8tDJkjEI/sV1t44qMgkos/m/x3LUyloS82shuuLpRX1dykLcfNol+XeoLMpKlymCn
qRdKH7gVM23cdCLPchq/OlKFzhTvYFByIbuR5HNFWJ+cKavdGoeiJeO7cdEG9SDf9+wm7mL0lG3P
NiZI4U/10k8vOWXcsqHH5ug4eP9+m52miMktgAPS7lF/Pgv6Nfb9Ql5dDFyETf+W6vxloc/bB1nH
hVd9YkQIktjTSg7bejCf/XtREvkGkJEHpud+q7X7lHz4178FbohYqTRvBNQSiaLMjikQph7oEW5z
98E6ckREsN6f+vWpr/17IorDoThq0fAz+AWDQMtJIR+8AQF1PBj40Fm0BUkiOwCYBJfyrktBTfh9
fuaATQngOwrpBJ/4WjQOeFlLEP1cy/jbIvX4QvsRljILP5NlV0I24YyYchmjAAgZN5RW3C75vBSp
j/Bdj448MXTkwFW99egC203IJX/GY57mk5pPFxYJPFbRdc9psdLtF7bGK2vGkjP/jJQfVsAjuJq7
LmoJPK9TJJ5zAgffiIzACtPIFbIHrPZPw2X7JLAExpJ/nAzTMOkSWlHr/3WX5j5CvLlm7GiBRHee
HWJrsEgWZDh69RrAalODGUfJgThtjkIUK7nxRGAFi5HVL+svysIaNjLelnn7pRa3AwMdkGQZToHH
Llq9cJIty21m4skA4yuyqVInGBBmPEWw2FfvBZ2+u0LAfPly8is6ba9rozwn2sH06XEN8GUNYj3k
B0zm6tWIM3oCKfq6DsTG1/tNMJfPLBG0aWkBoung3wVlqnGKKjiTmJr5hrMDdbeRlsfU6PquSKsN
vuYil3XeY0KvDVAV+rCIUq9s2U4DKPvM8G2C43lApIYYVvCfIo2IT0QYXJbODm/mOz4INJuL1AHv
mc+8DG7bQWuCGaz2lEPQrzl9FuT91fUggB4DtODAtxj2SYtKHKs/szMm0rtvqEQPKrGv1sPsbcIx
e4e2pXj/LBWCzB7gmeq20Av/0DYpbybh0XDZt8uWOnX106lxpGDZE7mm7SkvJRT3xIrAX4qMKbNv
op0ui9mitqRpuAgCbCxyBPpBQcl6rylxheraaU83T8SX4Fx/OwnNE6NYZm4xCAlTLhB20iqNWv77
Uhc5j9RCbau3OBbTBdHuDF7tcQMTG1Nv0jdxH3vbuzgFxUDoxr7b4vzd0bZXsFmuuX/iI11W3HFw
0GH8F3ItoMlO1zCDtt+eofOytuBbPh2bHHB2bvXMtndkzqxIK8dpZbwGrpHIlHXnFqdmJMkICdZl
vj1CONC4P8a0Wj1o+oFHv8khsxPSmFnk5QODdSFjlQWr4Y/JFBis2DQ40gqirAOiPEqgligweJUS
v9hAMwxauxz9zqhYWfneNibvKG+ZbRO3oRAEOl5qvfnwwNLQ0lRmwh5AS2w1mj8cw3kILNVDM5m5
PyK1YVivtea4Q+nA6FFBA8aLhH8aO5I/9kqm8K1AIQqeKqjjbfM61q2qbKDCfHBVvSSgU7VHpPTG
2zUSj2qTJNdv707In4GTaROgYU3Ip7AmSF63Phys0pMEO87HqnbEBO9WVR9BmTtP91ysLDKr9Ae7
VztQg1NDOQh+Zau9/dSzU+BVB2ocplsBFHJ2tD33UVgBa3XRMuPLDYiDLgumyLB13Qwl/SVsej3G
XTdcGzx9eqCm8uI4jquQ7LhDIdHZTKZ4EZ3wvLkKxunFGYpHpwR4ahNcgi4pmpCnydqkq5ZljFM7
udB7pE5X7rSF8/dH7FITSQzc/PovTmH9SWnbUYDcbQCAcLy0PKVxqOAwx8yzqkWAtDNWsVvqEP5f
ZBaLOtgiaMenzi5HCSAQd2D7esx1rEjYAtYsdVphWwmHiTzcsirpAnorJYJuj4Rjz86GV4pq625K
2c7OBUhwyLFt2L0MajZWfgJC7/hRdKpTaUuVJKMTVwy3dvbEiU2iaGpOC8vUiw6vn4GYMCavuXyH
Pe94u7h0IB4BxJ1R6LhDnLPOqqbHbDFTG4LuDnLheuC0rguJCgKICR+uOPcs0A73WB+AYU8nLdWf
iApcSKWweWFKkwujWIH1Ud45JU0feFOwmRQJYJHUsbedMQQ36ifSfFVnRcgRvSJKmki4SyWNV6kU
Y9mgQPubAZ4Z+Gbn2dFTXsPlMrN+xcMjdkyh6HD1eQcMcQt4pQEdod5+atDzr75SElz+6nTrM7Z3
Uf7dvbNGCqQmKOdRAeR9z1NAjFtbJNsRwWdvkBu+lGi40rHmNVnveOhnWF6iSEqZrFq9ae97B7V1
2RCiwekaI6kUNXPo4KO7U9ReCe/FvxzV5/yJCuoZ39NvjX4hw1Dm/eD6x2CJLzVZlRw+IUQf4on7
lu/d0nvpdl5MlyW9ZBUX3RaUvf6rgjTJ93dhPn4nxdFKAWbWguriw/YaCoYtTbjPfaDgxpnBegaB
jSdFcUp8iD7EDwvw4WS2FPzAIOcaFMAhlNVI1t8a6VHBFBlk/fmOwpmv+X76qF1IdNuOMq2grq2P
vguB4cu+/u/Hn4ugBuVF0eLYVPWhSi59x+abFh75UOiWNzAQEAQOKGhsSgp+ZIQ1EyoJiEX1bTB3
9sjCGeIGzJ7i5pEpYIhgwNyr8rxWuKEVAiAzTzR3DgVPz1lI9vOei+f5AcZpJpMUfnM4JzzXiTVh
+uk+yc74614R2GhUzyR/kwrJhgvkM02iF2gG/5zBRHJXCLEBZUHZRg3Fc8Hwi4ETFy+Ar5wzs4LE
8OJovh5fnqbXKCyWl8QwoExtlr/cZJVuMQQQih5IQCNYCSnr9DZw89cqP1ptdF4gDaHX1vhxIyNv
/W4MATNSpfVJs35HTgB878fmqM6eQHZFzJpfibN1a7bNOF4FWNNVaKTJxfOAgpTUYkZFTQaToanc
Ay9HDFFpFrCGGjQ47el3CizQcNc1mxQw6U3lZe0T+gCFCcOotRkAs63NqHKg20MZdVMmDal2wPhA
QjUPxntbCFPo/NLR5kjrGMcXQx/9kIfdBjXU4eSWT+vlHYB3xXI8+MTkAFrL6WBYkv5NtLhO/bOO
/AVg7p+wVB098Zfn/IFMYGmtx0gZjdQl7OhX+v2VUfI3jRoOstTU9uvuyktqOZ9S3u7S7HTHiYQP
i6N1Skizcxw6gM4B9fBlbxqD/whwzXXDMRbD9Snr/1A22ZBOY5sMqrGuiLwGZv1K2WbX7HKq/eq2
zrRM17q7wB6QkQ9FNXZ/U48SOQusbW+NhZtyQl0d5KEku5vf8wpDYtHA4Hyniax52L4lkw0qW/Qm
HlY9mnoHymAtdd/N3LYjFjTNQ7Uva8tlEkgThvbQRsQBSPp6g1wVPT6ChTrqV8icROXC1oWtQLI/
PtQ/vgpOKNXjHTnDPXtjF0+g0/CgJYzUVYTCjiwBhGtdW4k2F5U+Vpyh6JnWjXteA2B6qm4QSGGX
NlE3KB7m9RI7Kl/im8hN0jIJotk9+zXD8dQkdr+2+xM3TDNnot8G189OROyR55Z6rZPdGZzJaZ5b
khIb5k2DtJX50HthtKiqaOyrytBtwH3Lv/ey1iIG399jiQVyKQNtMApm8b+DLMWRm+oNCXl47yND
T2zJYdFY8Bb1oP1n8DVBg+i+tsyrmVyD7lcDf28Wuz7rQRn+vQbr/wPedsge3fCTBkGJeuEL7pfd
icO3PZfz7bLFz2kJ0BE7NrUQvFAKNBOPxhi1o3JWFQb/bW/8auAU/wkb2+j0qVmGMZyIsFWtcZa7
iopluugKrdRDrTLlzpfkt4Ky64i4mfpwtcFWJtcqblWy8f+WoIyXtGtcFDCvCkZ5SakJv4k9Pj0p
IM5xLwvRHKjUSabs2M+4cgu4Emg0/AppfuylkB+lkCaQtcBocZpDRVEQAsarCmBlFJ1KfwVnuWLn
YkJkVaesdwPBhOuAvb9uHl4XC+jZrOj0AjmlalmTen+iWqjhhRzvyIv8QK8I7WEnciaHbBAmeUie
pe75SRDX8eHYV3TDQJbko3tOgfZtSCzXl5ACkJS2Pf/tEJk618blL9rfz60sp4CjQEXogypwL0m3
OkPPzTCzskr193aaYFRkqxDSHTh/zFXLvu7iWRGZD9P4kuucuGFNJk93wl9gxeyoUb0jMhYNzEuw
L3nlG7f7FiA8OW+x7V1DcnyEY7zWJgzDM5jh3ujprRvAkJS924vfDpT0sUsSnhVF5WrCXzxlX5HO
WZ1lpofIkvHoyrFiVxC2j0WmwAItpKiQEC4gDoLmvikN0lYz0TUkCVdZFqo2ezELbX/FpdUIh0mr
kVtEUpiqxvEynpNdcLJJYqsJq8PjLhSlfCBkkX6hZXLRVdKHjY9j3puCi68Sju0akLcPMvB0HoUv
5KsJsRtJWsrLmJzY+8kxSBi+gLjr18ndojytAnS1pbCLaWKOX2JTjcME4k7rdUVSrSXCaoFafCIt
IN1CN+FMkVdplYfxVZ2ymye6AdRBmM6pFonlULiI30kAOcsE2VwTTxhst49QFxXmipodkJkpVnXA
esu8gHPxrbL5SSD4swkWVMmJpPts883IrbQnL5VGDgpeMdkShlXyYrOVdlE0Fq5AyEAPoPQqyjnq
m2GOEEUs7YkQBtDGLzfPKdbOqk9WkXPSxZ8cbqo+6Ha/CnFRnHS/qtpaV3N8GiOxsBx1wN1pLltE
3EXImkJ810Fsic1xqJ1CaxiIdJ1jKK0tjE5rcCkNWTT1N/OONBBDdZPJcOepXCh0/2BE/PZJ3mwb
2RgOuI5Ey0fxhEvtXlN0P35VmpAccfzN/UuRzu1JOpg7QnKVFINiUl7IcKfsoF4tn/q4NcsiODj7
vwoXgkSemzr63717ggVKZETbocXI0TgQySwheh86qNzd0o9cL+tQT1Vrhp+AynzzfWcfj4Z3HoR5
jLvN0cgYDPv2YJUVUwt/Pad6tu9SVNVRiD6oQss5bgpxJQeLGcWNcc7jUc5/0hHykXwd8V+gONV8
VKPkLHCJ7eodu370hUu1Iz0IdrNsvfTuEXOcAOYxEQvCxKF6SIG5S9vlDQzXqpTatETNkOXA6edM
wyRV4O+wObY8nPd9U02hxGcwPn7ICTX3pvnXYtxnSs5DkOKSPi0cHt/2jW89Ds+3ZGGKdnwRfM1t
e9xbqQg/1I8HyXiZxolP2gahrrjfeAQgcbxYzoM64Qw8ajDVbuV0Ilh3TUyO6Ib75NxwiH59hXja
iuKDmJvzbmreAKogTnLNhO7t9dU+neGWw+7IHfglYT1S4YwIzNr9e1lUSKJSkBzU+lm3TDU9e3tV
z5ntjU2bhbr+qP5EsjP497h4AM34zF1JEeQqqExbnBG9PZIZrDc8I3rU4R33GLFgua29sWxPEeJR
e6JCumb1zAo/oYp8DVhONGyyvMV0es7Ku4BAiTPJiYYMkxnJ9gYk+hwidQJtd75bqYZ7/BcInVL5
yStkS/ICVD25N9N3hlCFAHQ+e9jSFlrzSiVXh4lwm1nxz/QkSsEZCbDTNVHz8vKoCVTXLVIYr/vW
jRSGHzz2AYWAeItrl1V35OrFfBi+s/rmLtUvkx+wZdkPzoacTyQjS4zSU/EO+hRXpTSEhKw69G/Y
AzYpJVnOL5ukzojaxF0i5w1w84XLu4ZyALhzumd5VsKsHhzGdHt9abdBVTihoAL8fHbZU+V9h4M/
4zjC6wAGxZ1+BI4/jua8+ay/AtxlQa4QJPOB4C5AvZZXHZy/ZN0jEgqClaP5XEjg3RwDqpcovqcE
NBkymDoB224mVxGbVvtnup9anmy1HGz+OhHjvq++oG4xAocvh+ODKngvh2Dk7J+6cwvuoTc74O77
I+x0jlArrM5IBGn4B65vTrS7uMLvjQuRSkMgjI5uCBBVgeAda0QyfRypfBmwVE+1n4prg3hajZ2a
N4v0O8MvhBTVY5mR3iDESkekHcl8arwHwECQ5ZfXq08mUMt7Mp94eHXC01poj1h3/5JN99WaRa2f
H6AgikBvnP8qXHiyZt8uOpI2auWY9eLIh7WWle29Tjh3gQaS6aY57P7g/P9fwUmbt+eJQ3ZBgWJ0
owiytw4vlDYttmNFFTwY5i4c3/0nzo3rmiDQWt9FbDFJ/X4IaMI/kv9CYUjaU5henJJFp3B1tPZo
EYv6GcFrdQAkPiOXAknNMqMe8zK+T2oocZXJ1UaF5MF+xhCSPn3ErMO2xBgNWgt/dQmptWltivv1
PVfFb5jKJvUU23ic+CKNvpKyAKich2Hv0ltNfwcR7jiBX9JVTo6fChBvPi20kTrIZkXdKvkJRIzC
v5l3ANOs9NKavx+W6qVESOt032tJjqsRl+x2t7CPbox4wIMksn494KgWaTtRnDDVNkIIqjUuJ7ts
Lb084GwTzH9ItAsbLqh4r234/wO3oNPULfWydJtwyGimLCobeaK8TOR6LUDb0mwbJe0mdNgh2LJ9
oGwxcffY351A6/8pf+AKThjM/PuHjApXlMrXj2sfTaD8xrQC6S5ktomBr79ziQHjWc52f8d9vkVM
RL73XDh1Dza8EJw4eQgez+qhdYUrVl7/b7TPAbJTcsHLAOTb34Vjh12HIBWG1laYQE1juLa5jrOU
Pp9TS4A26f5gO2mjmOZgbwS/32kon6SlMeRVvfKx41JCnBcGTtuR4+Yq++7nfL/rJhLlSzp78Q+P
qPlOsm6jJIvcoD1JLCLsLJBKSZs6Y5T3l+iqyjLZIQKJAK7IQKCbuic1XiBWq1IUWWwPlLR87jfa
pa4+RouLOi83a9mqym5wCD0tdjfYrA36g+LR8W1EjMDrnyH8kN+omlgWWMoAP4p5llyhjLganjd1
t5O2vJwlzKOYrSrwb/A9TadCo6aE6ZNvZjUeWiPBmLqHY3pWd+18Tolg08Rl99cUc+qwozWwb3R0
hFURwholaqkcc7MwzgJ2KcBoQDjXGWKXEZz6ruO+7ZFF6CSJoeVUYMrwO/GFE5+ervVRKvdOQGUu
jWwLERg1mTAaKADA3I65kFKTKYHPbcVpbJwhP2YEDaL6v1SZoB+sQPbQLCj4LGb69gcW/YkzdeaH
dCr4VJIBmVaHWsuD2qpFwFJAIuVtKqxg2ha+8Ly1NPS88k6Vv8y6gJYpvW2D7+F0j34EfnIkKMPZ
q1AcMWxWa7TO+zBkA153xBjAyiZ2MppHtB/vWDx2tpqsIogutbqGTC6Akr6s7Yt7sLwBhjKKY3M2
jp1sJar0hoWtNqKKT9b3u7Q+fQ06B9HSdN1jhm3jr1AoTKjfkhp2odDHhaMYnt9UYYeRljHzpeEp
SuaBkXumnjePRCC7FNm1gfLZaMe6mK82+dGol9h/NHMzq3sTIsdKzTMUhi7Huf1MaytHgHa7rxvG
HCjt0CZY38mCjk2GnwJmtvLiEbhnIMvfaqzzLP7u5JQwEIJUkbRv9OW9fwk9qGk2CUxGWR/kRFyn
EoN+TdgylfIebVjYfuTaAwHBE+JECE14Nv2ZEyGCh/fyNIZDhwRcayKXA5LY19enNtIkr3CfAUeC
CgbcKqiT1jK5OGapC+9DAgOcpgn9tiYC/JvU6BIvSGiMciDcSoJ1upk+iOhicVjvYMXlim4ICB+E
yz/zZqlQqKodY1Hut6l09WOl2HWDUiuyZRm5M4A8+bKghg5+sVl3hqGp2jkUZjx5bJZg8UkVGL9n
07UN5bnE0unxWeyvLkQlUiP0ygEa55/obg7DbAKT2uSYwA5uIZNrT0kiNIGAnbpqOLcuf9rvTk75
435i1lk0tpBUV9CMWlZymjKSr5YpndgSvXwW22mW57VHlTY7xXA7xkgF7+Wn2hTHiOWv60RC6cxy
4sUI9wHd+LMADv/5kstWfTG16jA+LPxSn+06w2EPy4KxQApWfGBJfveq6walYQW1RsIB+uEheK9Q
DafcWJNFAgWvdDxSSoJfFfS9uXoTCr9Y5i4wwN4S7EFwl837CpKKDjCZaY6bM20WZOtVgMvuMw5X
nQeUk4nH7j+h/MRB+1O+tkOsmUX9EoD2APGxbvQmI/AWKZandkY1COW90yUh4NYv8xiHa9sqYGne
xnU7A3n4QTI+/hOItmcveb1SmxSGDe/dOLe1IZJSfy6UzCHod6SvVAnxxUQhPFLl9I3XPLBQ4zw/
fEv8cS3jgmmEKyZPzXuO3ehfp1+SysUdqmA1D92hW6kVop2u1Kz8cpsfWdcUmTrVaL/qcL1kbcwF
wjDhsAWL8jUwtkgruzTAAGERJ/CTJRWd9EUgt/AUpOEEQ4yETavYsb+/6rt4V/H4k3rRxNOODAfe
7DRl7oIU8O4ebRtCbIdX51VHpMzOtgq8SIqwbM8hEsQ01WFSXtGv8eesEDDX+PZjs6dZ3qEGdMAA
C2LGV+j1kSkjNoUp8N6pHM8gfD1VW8YJc+n/Z+rvbhZNOaJ/EZEz0TFdlPBb5giBrsu9RNJKnODH
JdBz150i/Lu1+ZA2rZ4w1whGPmXYdagbb8ehXO+P+J1N7kcCUxq0D/XdrV6BbYSQMBLQEyW59uVm
6J8nf8wDJ1/B89yUHJ8JAVTlpjj2Kk9SlwxbKfcNcac8emGMsJvABJf8e0XW8aJQ1bzehNhn+9Z3
1RSIm7WurdsJm5qpXE04htMn3cF0pc2/+dLN4+xys8vP/STZYjwNPRXzhyt537U2/aHtY7OSIJse
YY0h4X0zoZZsycvDPtlEkWZrzKwajIZI3d5x2/vwYHNUWp3NpvK4OxJIn0kTTRmEzgfHQP4S/YgR
vnrCZpmbCrWlF9expDyZ4DYt8cx4K/D2ddYehI/e1cZ+SAIhUy1mppollLcIyv3NBUuKmeOMGj0D
eaKwnqOtIPTr6ISv18PLW+/KQOe6dgPpIlk2AadsYtBL0VwaI5zwS7AaDV0F5598kvT88abpo5PO
RkfD4igPLpcHDhn0WhwjPOIx6qazVEs+iaHxOw/yxhMOMfD/HXDzPr2KnYUU5+pe5Bvl+KH4YXXy
z/4T5LBrSQ5ZtZSidhEbI4jJeri+ZTygLpKj3fVB+rJgpWBmsbUaEc9B5Xa0c4iyilug+8/EhBDd
Ol7jJXH7UIxA/HfIaH0Fsic0YySRHYPPJyfjXa74qrsU9IeQ+5UirrcrcoRv8F3VC5COB7yY2iy6
AubxdgaWJL5CCoAllrlo90AePKVkStsdnkN5xqs2Pa/GtMH1jaBF8Xk+tAnCN3ntTr1D+OIyIqyF
aSDoKfGwsF2lwI6YQBdtnNjsrRvFgyr2vWklyyt/Hne1p/Jw4dtMotpvVVkEXp77owhsS5Lxh0lN
RXqzXNwnGSmVtIOCprmzfSVykh0o/LYcoVi0vVZxjIW/qiFZf9tRHJxMxNyusYaJHZSr9ogFAKuq
pgv8AhBqguGRLeH9IjfR1NtqTShiwzQnn2441EIT8f99qbsz1EhhjxjdiTeBRxGy3T6t8AC9FTJt
0feT45Cdv/BrHLtomkrLebFKYTdp7qGF/HbZkih/Yvovy3qkEKHE/X2WnnSzwOoAcXzWVff9jnLX
DPxLUELkE6nPNCEiiMl/QR7X9eftHYDyUsUS2OalO/AhECv+GkCxQQjqS/e9WJr0JuE6h8CJvOEt
+F2RoiMMzfqJ23nHPjoFWl4V+UTwv4xgdb5fbmj76ISeaybZx8fQkf/p23iTqaKFx8XqWndM2ilJ
6RlbJI6JaB6YdgcfLex94qOvqOh4xOc4YVF8QyexsmfrZqSE/TNOYNyBXXvwz6JPrCAsHULt2sc4
N4AL/adlDzav8AKoN1bSwRGSKA6oVdmrmNRHjXNFDW2D0a6nxT6SahLEjIISJZikwjM0kZQBbIC7
IdE8IYri2R3nbmcu8jzix/m1ATmFUrk2WNpctjSNYQvRR+5RXii+5sWT6n538YqVkfL7jUCxTkb+
FABMkErH4aP/zSgFUFeQ8XY4iR8X9TP8hvfTbqeG56wTPq9UrNswD0GUaee98riEHtsoZ1zIEiPF
pHwPjxrN3WT+/jyGiqfcX0/nyaLBWVBVDPxRgtDuVIp7RJnx65AIFUzyW/DbY15ZUsWmnwHIwtVI
/bIBxN6gxYC/UP8GEWM3IvOsVP3ROXM6hq+qxGgECato/VXZn8zLlJrADvZqw6EOkzpWb0YEupZP
K7NWSqGGSvadMVp0xn+KXhBbkyspBgDvQmYKloDqROIaV2rgrer7PU7/ybzo2noY14qfRaFih9ds
TPPEdeJOrUQo8xwn6f75awnsjbK+SAPEqdNQyk+As6y1EmKU9/0Xv0jGOzYOn9u8+WAz9/SABQ1T
aE1NEB/2tGoy0/SMcbTkL/5R4CF6m6ZIUS2nHbX8yBI+ywYcwH8TQWEBF/xMN02yq2SebU9JWi+O
YcoZHTWYL/o9o41PagUPuruYAm9WLqTegVLiyuZrhx5VgMicYILgCFRemIaBT8E6VIMfZf+kpoLK
lgqa4T3Z5NK0CEpySCaNCfMoqD4AMfcjhHrBrTRgrHuQt/mRwV3ZJOiPSQX0ePI+EgOn/vLyevVl
pvhjZNpJB9oI4/KBrIRsbTDpru2n4Yak2q6hyJiZSVimQgIojaj33ftfwMRr7F3XkpaOrq7qmvA6
UZPkmdyUA7CEbJumyXmD0XNuLg1lIQLKcHlCsLWKmzxiUjBbnR0pddja+pimZvAHjQJRrqUfSBjH
AIhVuslO+iFeDZPGMmpsxd3Ojf65L5cyw/Oe7Q7D7vWeIF9Rn/9+nrZLpFdZkd3caHArN8qwy9iN
W3Bl0EklctsWVipDbUvC8XNVlCBvQ5QQQSH7z9/Mt6AJ/NLsN8js4RnV8tO3TDQqv5uUwsNqAmVK
px9mIyoAA6aPDSC0KnzA82wswpt/P3UPkwe6tptQRJ+jbQi+aJ6TkxGOC2JH9BX9mkFQvT1pHSqz
tJU2vj92DQdfHnVAROVPv0cl8Wo3x/7Bn7tfiQZ4Hflym8Qq80UxPeTncPOYUwLT34LLQcgTZ34N
0saiUr/coUsPvhdMoGLKfPl7ZFF16XCgkls57sUAP3iAc0Ex/MtIt/NcMJLvRRTsPin/zOxBBkp7
4ymKIFyTgDk62TqUnkyaMhz8RNni+Mh6oCCztWehmvXUSOqdm4764uKIC7qzl2NlPVyTOfeGn07J
orw45/0BZjzxgmqfAZyCgZj6721gjZWP1g8ihKLg+V9XfcE2j2Er/QC4fCBc5+BjYZqQh05Xd+zb
az2AmDouuS6yjVSpgiB21Ou5j7MM2cBqTw9n9ljmRGrlpDlcdQZ+djNC2+MWRmBfchMWrM9HHEyy
oNe9h7f3HvghF7ZFS42qefZos7g5iM+AcaCuZHTjsVcTN91Jh3rpguuztMqBgxmAXt/NK8k5/N4o
4NXNV3L8AkdZR6wK2oBdKblpvGaU0nKQ9waFGhyE5A8XoXszjTzozHifYq0FK0ojLiMB5Yyx3Ja0
A4NXQMLm1/jSyn2aOb2UiuZ7z9g2nL4DcmyiH2y3j/pZnrrP0pBdqc6BfLS68nNk+BBTVCxs8pOC
Gc/Poej9lYVaP/rXe/S8SIWe6ZcD8fvbjecfUDr4kUSo/UEqqNkcpWR1tpHp9fdaHnoXJvlAYlaI
7PzUWFdh6845PFp/Lcike7BIBS1WtQLIqhvHOmayHtbnpGFcARq7pTR+klSOKJ+GxpfQ5sdQI68W
hVVirDTgfiAAYnEsyNugTSM6T8i99pq9PpFr+FvOYcXFZf7W39D9GlZK008ukbgpj350wzsWMTre
C5DYk4Y62IxArMiGP7g50ZlqYHK/lIxVByK0fHfk96TO4kXlQZn545LrWwgU9WHEwCK4hZvC7j8O
w+3HQhI1UQcTnio6hKW/gaIvlIpctExIc0jCQYvIlh/c+PjyrZmjN6YDoIhqakNqaw/7xbvxaXfg
F6hQC4o1pDrtXMNOrfBEWwXhCC4iDYMKv7j3We98PUmSgtdX/7CJZ1J9JGHOIDS6LRudYNExw2Wp
IdQqNYrm8sM6QjP4SMbiQ8LJlNcxpazcHXUsOkDxgD01MWo2f29QrtBbbi14PF1sIpz/2yROKlTQ
nuYjhvvwwvoqjQ/5tx4Di77/iX+FrZborbLfM8VGlfhzNiaqZQUuJBVzq4SmBKJYU2Dtn2MiTGOl
5moRvrAzdI2hmTAPFJLU5cBYwRxfYfBA49HJ6AN8qL2FTs4400YzvwJR5/tbOjy5UGyqcEQOnE8E
M/vRX0jLNe3K5ECT0k9CzMCoeJoS5fuuCNpgxiR9qWWiCzi0Z6Ka7BEayI5odiGqbxV6BMLszW2d
ovw1iyFjci/ndvbGRm2kBAeXfFlfwugNJVl44WAgUD45Oy3yMNeoE6e/SPxbFoTYax4IGJTwNnr+
4POCqcTvjGY+rOe5ekJAzdQv+PaeyirlsdgIRO+AvbcPOiUZ+acL260V2AdRZCFoaicjbvkMMJs/
bXk73j0nDJAXxL5YmkinpItfUGVNlrNdjoIcXEjQvkyXyW8sE4oEmK5AyHpViDvp7pvhJ89oh7uh
Szdj8vuWqLbZpcVKOPkqU+gjr7Y2Rl3fxCrxl8TlmW1jimjbg96HIcCdn07/DoXveQ4olYs/TOYQ
FgXtgKsdQUlEOKCv85qY5jCNB+AvmGgAFpR8OwFVoLNDKOJPz9xIqKz9Pxz7S48K7TBClV9A4bbF
8qTNfwNOmbxifORjAIvxsU9ikOAhjLtrWrmquzxXvl+2WaBkrcRC0zi1qjkiTAYUllU/X6iBklNL
QOU0d5d7/qEzh/LEXAO0ETkdpDHOcuV/TAFKfk1C73Fj20PTuzbbrd3lsdaijieZ3GUzJ7362M1W
9VTq2n6KOR9s3/HPa/1u5+7XUa+9w8+eTEVN+Q8u+IaHcvHDPsUM9lffkfbE8l1SCSogKMr+N2cv
N7pHj1mH5KTNBQ/2dCUiwYBEhvrMzKbPuJa5wW1FdhRd+JDxYZkxHEhw3Ld7XV4iWguAhEZdg8hw
NhHv9iux80CARIvqYku2mfj207KAXEide+WUApa7ui5Dfu3wsxL9nsHsSMmnmCtsVeZ03yGO5Xkr
FZsdwXi4R6wIr2BhqjVEcjBgdqXXsZlnKMwna02JEbw1X70hwPcf3hOUivarWSDyciwW1GQWHF4V
p7WciQHZ5eJv/b674PTv7yTV8lPCBNsCNvsyI+DqiauMrLg5MjAlkgBoSWFxWyLuNf8S7+41lTZg
4o1YCp58zb+izpRcfg8r2KDB5VEWhZ+997FpRFdB5NarcFM/38kQCkByO0BqM6Ay8kbTPzvi7UGq
GuVHBZAzS6LGX6bXuC9jubW1y40qtVmWe9AqGsH/+YFSwXHiE02O/M5pMmQ1Vf6wj1LLztlZy1QM
rGSL55vBMohffQJXrNRpvZu19atuasCptoUonpmFHH03QLimMvdf6nC9yf91lnKS6bBBy8kCAoek
Q2mm9oydZaUZhMmJRkFaCyPGLcpTmQXlVJk+zI3biUbXikae98DDZQcMztivwGjNLEKfV6T32Gig
d3CywXhUubzTDbXDVzlScjojixvH4UK15O6q2qUFZMZZ+TEJ7zo1kVv5w/gASGkvYls3Z6fBfSth
ZSGSlNlreXTfAGfxOun3SnzHrvQYV2msXhxv+e7JHuOjgJ24nymAOZNPkHXo4vl9VItFQlpUSZxA
lfAbuPImAZHklsTxlJPHs9n3jZzWhe1vS5aEfIqF0N4jwfMz6oLBHlK/1/2siHj0U5WfhwtJt2Ua
QZGu0YBMxYTmqdL+DaoXgQfsbeSbMh/NAoy0/5p4r/mUQnFm6Z8hCHZ/26dZAHmFD7428+jt6KwM
xAqGHoI70qAsbLeg4i/Hhy8uAdyQXZ8a6n4kcKdACzDQA2MnkpE+oWvVQGqZ8YKxUQB7gqGXj006
wclnR8yUyLrAufACJFrRxLjNa9QQnB4SwyWByadt0DVAbgLeSxGgUAVJArTXMzCTRh0jz+MrMahr
VJdWmX0KW5Fh7s1vJ0O1zmijW3QVwBTkpm7F48jfYUYnwUYtG3BUvYMkY9rREg7UaNCAzjWUcoJD
io7jblcZaZbtGBYYk025HyOiVdSXmw+rM572ViD4DweQYjbHDG7KOaaARgNdy3FSSvFAlKD94zh3
nCzu9gRdqTMRS7QK6SB5870EVdIdeO4pwBO406ITTU6KJFDgPdDi3qVxxe4EpZSbhGKKBbo/FA8Y
QxLbL+luumABAWzv9kbmSkezzl7r/dFg9wIfE3TGT0V0SJUIGmNOtv0I5fD0PhclUketme54ewim
fo49ExdRfWt2DRG/DVftbzoG77wPqn2rCRRnRBzfGbqm2aE3Y8WXLqf5ivxtOzjhb/oMnakN+K++
AewsqTfLymDETdTaP60Q8CfEgQO6oE/9NvaCPmXul959uEfmnEWlPV3/kHgdKpnYtrcuhwaiKsA3
8NHamjhWy1xo7lPc85wivTEcQv7ZVziF4F2ihDcpxTxVp8sE8EFp7nSJaIO8sIhQoJ0N048epY49
59OCuL2yOwp/Of1MR10ncKgwYP1PaDWXXezm4/OmCY9z5eILXA94z6mcG5koiIjC22UAVsm62QCN
+7S9cgUkSYKxb2GFnxOSgygqKX7c1GrMR5IqaDiRF00sVN6zNtmBJtA6D3EzTnlAe6Pie8QuoisF
Mzs1UZPoNoSH93wchSxB497bNx9IHtfhAZlustGGwRjMa3NHfIcNJjhEAF84uucnVsm+Bu1JE8lt
O1FEYQlFgvptgF7VEPuKTpSImrB06opMetUt6jytC9eOZTwbppfkJtFTxEVt5gDQrXVci86dSgtH
Ydm86QMqYToDRGqzXYnJoDF3KvMPrkdL0XNdFM+xTFtFdPmwdjJQ8UtCpxEYNshg3mloTFGwWGBk
bCyYF+js+HDyGnCRLjIST+Kq2e5uI0MVV/l4MMHl1+tBJ1L71jtv0PtjYgcdEU0sGuIyG1f4Hum8
t5dgl2TjQStXB4MPJphRGooIUaj68GoxT4HKESFSsh+etQ3aHQ7pNhU3DCM1NLDdj+kDSQPNvQRJ
8IJDZdmLqTHOoKdo+yRX/ggfnIdJbXFiN5+T+qKK8ubS4gQnCh0Q8va+WC1ulPS9/4YVM6YISVQ5
sKtyP/UcuVvz/GXLRT4HTzkgzI4sACgVZzj/Jd4ZjdlZ+vT2VMXGqwavsny7w7S+S+S4e9jCGRjp
eOci0OWZEBRKc6nakJHlAGUtPRf+qFUdtZ8Ul2aDezzp4Lv+mbbzFeKimySWllIlYvl7RRVflcje
tK9OYI+svPXWwWsP6UHU9peaYMAWj24/1PK1nVcSdxo2H2QgRTQ08MzzBneP24nbWiS/Zl0MgTQV
4OJo+ZY4pBWgRB6oSKgDXMGXB/rqMdqOu554yv7gqPggh/UUtIle7QDmQMa9/RccKaooMon9fi+0
LgLXrZFZgnSDcc34PgqZ4FGhLLmp1z2mBKlXsOUj5Acb6SONIeZ6/ft5HdXt4fNHvS8Z08NE2EyJ
uB9CsyYzcT38NyJP7tvkY7ctfuvKkBseMB09pOde7e7vXJ/Ecs5ADXpFmv3fA/AedvpqNp33WFa7
ZR8wY3cMic1V2oGP6IA1Xhmoi0mvbx6NIWVpLIg9W3j9QTW2CqLadsyDl9jHksUS1c5mKYHP5uL3
MkSiou+3vXnDqCQEQbsJZw2V0UvXTb1WYi/12di4sqthSCCtcTOTBZTjV465tm4PmBKTjdCOolvZ
CqDCLKDYk8RQ5MLpuhYxRL5hv5HaR1FGkibHuTLXTfumvZaknkBJuLbGeSNTuRJBSoGIMeyIX3mS
S+qJXHHaB/Gla+Nt/M44XwG+ycDsOEn/OJzXIPbTRy0hIBZKDgmDzoaBqAc47vZeC/J+gzuUOIaH
oCqYBd0Y2dds+YmcGDlWlCmEMGgxUdrGbsHF9Mtp0HJ/nwvsdWcwzCm1FXrUsMNPo6YwlpbR/5nb
lTQNYzn5+x/FK4u8rmwTtCX3QT+WMk+yuQ9e1zgR6YLKCXtcOuo4EFtGZ0l+lrqWroOveS1sm0Kz
qOWTxoEbKov7jJeXbYVqsD4bwdtixwhvXudQrwvPp4TW41QaATiaczg4fdcDStKy2JfJqBcIlJjR
UOeQ2CLpMLTNtQ7hmAoUt1TQ8qwKNQfnor9548loQcr0oAgxn4MYEkuQgzsrvFAc6dntNSofU6sF
35z5mmz6zU6z5x9QrZe98mqrs+wXU4CX9QHMngxjD0I84KkV/toZInwRJbg2JdUpyk8eziCpY6qy
LycPbLeJYpnsWL7p3dFVVRHumGEsr/3esrMO9ZZPyEZ3IiiWV0IQJs5s96OldYNhkyqu57aIQRXJ
gNVQyoCieB+74S8LFuJIVERy6A0Tmk8e7iSdvZs255rQZ2SQYy5mAH3HIMZiJWFgzkhMYP90Q8ba
SVxvDnnefhnyJqQ8zxgEFD2hEWrRoMM+/Auovqz1mejhpLxLq7F6SF+lurBgS4KbcHOXqMUoDs5B
jIat6sA8UTtzLFy1xPgu7M67ESiKyMys2YL+PnWfUEc4O2FtoC9w+OMEanfYyqECm5+1zfAnsyd1
oSXt8cyDMkDRBjOX60RAcInYXYJpADMVDO2SfQacAjbFJXkjlqpomTa3UZH2DhvIurlWFT6gChYR
cvW7lLmfyWLBCDG1gTDBx0hfY6XnD3+v41/6HIWIYeNVrAnkLnQsg9W1atKvKbWgnRaITKNYFnSo
OLyrCNmXyXxyISbbPyq0U25GEcwdTtKebSqiv+13Mlu3IhSYUWf1yDCkqRQrjFEy+dX3u97txJDC
ArBct893+pK2Ql4PE6ncYpFRHq+sRlmGijoYVJqZ1ybbL9jPLGbgPhXpZKvPq1HO6y2CHGiS2Oz3
vsOmfcznaTcPYhbTskVptfWto2/0KZzApDe58ddL8qxf/LeZGZiAq9a2KOLxoMILOyJFzlFCl8xS
ZZmRaksPK6zEiHiKcM1V20szctP1i1AXgdGJz/sxldbSk2rESFFLLxjP1VvJoLq/bI61BAvZKAUf
EGI9BvIFDu8qqAxuLC0Byy+MAXBOP46AKeBeHR6h+89GwolOHSdhNoz1EE+TubBJjwpuHS1Ma22U
OyU8Eq02SXXTzd3OJFbKKcOTt6IxYSpWEPd9NyKKRmh/qUeTtvqK6/30oiRAiq/mN6rgesnB7NS4
sG1cnfvcRdSpje5iDh9q4YYqnwA0mNaa7wjrp+anuaxpNwg7mJtS4fqCaXpcwNwWQrNwjxLHndsD
tBoHGBgh+cHdB1Lvd7tdVOy49mGV+90yklfmBjsgx9v7pIko45q4vTbm4b37I6rQ13HbcBEQz1Xh
96LJiU4TEhhN4pCwcuHkVoGnTDHbUKaMUmYQCYTxYMi9LWuOy99NrJVj1ireWhlVi1LMp6iHh0jb
dXI6/0LsgnW/UBBFO95kSQRQjTe2x9eUDYUyHHqTyB2bOHrWLIQUCq8rFWQP5FjtI0Iv09pBPCbZ
bXlCbvifOr2UUIHjzUqBYO+MsL7HbuGe1mGcXgabCGYYX6MgO3pEE8YSMsLIG/uL4FoJg56kgTK8
ZnJ51gnY21kuzZw0BoU+YBIZ7ulb/7dWEzd9VD0lR4ueT58SaGZXxsRs/9WlObTsLPPIM3J+A6ZQ
NUZyXo4mHSmnTBZjDYvVkAO1CjC9Rk6msSQQWycv9xoIvfjTRU0SSiwl9Bbi+EOTvMbPHI+sw81U
UU4gz/KE7UuKLcx/rgKoI0MXW/7mHld3kWWKY+uXqGrPdKIJK+wgioJRSMPR7ZXLdjQ5gAgOTdjv
S6DeWp5CM1cMymHyzDJBdrPfoqPwmI+ezVjFuQqOGOdNzy395cOQf/yTV4WXEmgrIvV1jbsf1N3b
HA8z+634IhlM5fg4ObutbaF6arY/yx2B9Z7CBSwD92yd+DBDC0nEI4QUzbeR0un0bd2MMeafcOvi
G4LsIUPIdfIiITAjYzTkV4phCYDp21A6bQSw+Hz3BIM5yJzf9dVEVQooTpITmN2rrNwwZ508KmaW
qULG817sgtO7Tj5zKiZxB24WslJd9bIiFS4O5uDckRVlN2BqPNIKrFElqnGHuPt2YnCEvwgEvEAg
SrIs893a7Xjg14oF2FlNF2aZMyYB1tc73thGUASRLWNjh04qvlXC5RicyoppnrHhjLgtANG1pGYc
9ZxBnsoUNujXCSkWs7NocGYqkvmRQqL87CJQqxNbIztVZMKTvrepryPd2DbndTZ0UXJ7pzzzzf0i
USPKz+TN69Z0M3mTJgNPDCnjiBBs7KX3QuwHnRRbV1pts/qF8ghA4RoSbMFOrx/l6nRY1QiY8VUf
15Ul78+uEUwqsC8JYqkXPJOCFxuDQMgZrcYABcDcSiuv8OBXL26BboaCKIHvmt0Zw1mXT9N1vSxu
RdGzWsGDX12akD6zdhFtCyKt5oQ3aTZebGlMmffDdjVRbJpXlET9LtvEtnUNFubizOEyUJW8U/J4
6ctDtEHEJuMQZ0aQmyTSsEPDWas22V36WIXk0ofSRWjv1f0zJBWqnKJ/cHiw9V52RM1/7+lVZGzp
5otEXTPlS06iCj++21owrE1Q67FwZtyvH5C0ROuTJvvhKp7aanGEhF/sf1lj6evKM8HqloJXoCkQ
64rfj+Bkg8zAgWbTZlyvw/WLTQcMxGVPiqgjeAVNfa9cpq8tRkCywU0jbhgl18ZZbykMQGFwXB8e
g8CxmnMpPXQGUw9s8vNB49wsrEjJH4Fz8QiYNNRHXRLWptfLgxpYVIPt2rjKgD2SNwZmEn3rFnny
MWhKrRlgwRjPTT9BnRv9dD5gD2vI6uDIZ3rVONwo7HjdKsl2NugfUJLJ+46Neehx+tOHYEK9hC5L
AKxD8ZwM5qM6wwhAQEpCcNciKUAk3agNRsSAt2MnMCneA/BOFAvXNVI+89JhJ/KAPiK5ykAeGgIq
WloOXzSXXdPVvTa1KwOUeCs2+MjQRnJsr/mo6MUZYmdyZksjabNd8/03n6OTQL3jrdjA0cpUDN6Y
9pmeQLELSgL/eugYDY8OYFs1l9h+nt5naS+zDO4G5A8nLETtWT5TUl2k2UalD0575TGTVg+Jv5eL
KsnefM+kjTE/Cu5wZ18TmcQbslVlp7QAZD/6yH+r0P0qN6n1DV6wor59vg6gG8w7lnYJmGUuoaPS
vzaoeVVVTBq+QWOY8iDWJAfXmHa89xl7tgWYA9rMKMBAlDJiwuK0H+zKTNxvK5F7FIgw+8vb/5Ee
tgtW+uX9xz7mbrRP3w8LbbygUnwDt7yHe+GX8qzQnSalFr0rlmFZ5J2WetP7qk/fn0DUcE6TdTf0
PuIJmsLwfSaUXywoTMTHcwPf3z5AhYcr6+adtIk0WdDr8W8ivXQZcSNHChhMiGc/gwES2QC8aFRY
CgGGuONTgl010weG7CSQeL/7F+paUzN7RLVlFDIZ44PEnAgCfKuJcp8yHSB6W5v/kS0uScs/vpL0
L90Sb+OHLNFRaNlXEhslJW+2TVL4PUHK0l2L1G5JjXlRXjK8ZWViuHPCTkCvtuPbLLdh+gXLtT88
StOkXtla6py3cQVUF/JkCgoq9McrYhTo5nUU199CQUIxbV42XPER11Qr2xLMRKgk+ZVa8lMTqEJH
S8/ZyoajRkleGttZV1dwg5axpC5xxqlXC9q7xq48bb8dWTXGHRGKE/6YbLllHsVG5Gl9gey2WBRv
WgMHZxbchVj6x2RANeNBZfTiS+wRx+VByHYTGd8BlQhQGNehrpoD3QMj05YMY9f1B/zf2fSESINx
Cg2pa2AiI0gDt2tDWENQka7wVyz5GNp0QZednfQC6IJv5XsEZ0hWPJLgGU8LUXtVpr0ksL0arKmx
2k1z5KRn2YqrcnswsC0vQvYCQzxeUV/phmI2unl5DOXvTNChYk4bzXPIQZJ1anMVrgZic2giEF7N
h+Dtm0eDEPEgtcaqWaiBEo4SL6fUzJ6QJcNb11IsGxyJchh733X8nUT+BULJdYKENUACIZPOfR0J
obfBxu6D1jYxjxByDDtjLn2kf7dF3cC2VrYUmhDst7IoAav8YALX1CfPaCkCI4T8Scc2bVH3UW7L
3OrJ0neKEgI7Ua3ts6OrNjxGg8r2mqkCykl3F0GzlVC90il/9LO5EnmeFhYYlz2ErVkOOBlE/htu
f39faXUxEoAS+zF8ibD3SLlyqqxEHYNBP5ZlvK9unZuuUISjWFVPyAzxUVqpp7vfqqt9skTx42HI
91KKEsk3ICXnjPfLCBfTxxo6+4iVZVfmWN0XOMApWJ39zN5d4YusDwhB/LNhlEvkQ7V87JilNJ8T
hAhPRrLv3vblyr9dhLX5BV2FpcxQLL4LtHoYYq1s0a+T1mtWUCPxVzCnxFSVy5mey81cn0/1mx0o
nrR6frpcol3dGcyKJFMLEQlqvB9zpbqWaUIFpEKwBqIw9Sv8CMJ+yOga+rHqirFqy6LWqudC3mu6
s8Isk5hqLMp5mg+jOKsivwz+v3eubFs1MyB3d3pAd8q7V7oUBFFKfhZH3R2Ei8EpiLsN119s0pRZ
mRh4tyMaSl/Dnl+1HI/7TSf2CKn9FafL9Tf9RT/u/Wzoz+I9GoeDKATTbOhAM0pr5NPKokDOdZ9W
d82rISgPp5eNrjEeovdgxhh3X9sHJpPIVEoF2MjNWXlOrOwEQdgNne61HpcH1YqAYzzk9SpKQrRI
ClPBZDk6sllqjV39wqs3IcqcGvk3IhPiSbbg69Zl6VBSSeJl5Cs6HK7aqODOUU0F1cqlDTdvpuSb
EFfRfrk9hM159+MqeNtUVVjupRxnvIJcnQSs0e0S2+oIqVfOP54tMKjBNkXAAJzYw3PkioMQzHlN
b/2zsPlPF2piW+mURx2PWNqHFXydh+9ZDck0t0/bom++C4FcRsUO4slCgT+9v+d0mWoU9UmtcTcp
Kpgi0luZ0+ayvq/dfDzroVxPLAtIndjEqmMQee43aZ/VpkZ12+z8dSh4YYBvbYA81GvmixF6wGAU
y3y5u317OIXk7O/InQk99gsVvMLtC2CmyATGxpMooVp6C3TtPMSX+aDANhyiVcH03h5yGPwj3vCN
3itqztSe4Hc2tdwEKxA7bLluHxpov9Zmdl0ucwY6jrMt0oBYkbSyQn9wT1iXM0MdtEz9fn9JXYwj
gV0l5irH4Wb9LXefaR1/DTSijH0jwmrpp4nUzp/PzbWgtuOalZE3UUob9L9EF+emC0+4ApTAdhAW
HmPeWCH3NabqZ8qXtrzNgT6zoNfVInWTwxIvYEq/1GUiVKope8ImRIoNcCOl0ERGT8uE1AX4LcJI
aCFRCswd1v/dRzahbGvFgV6d+W1mHNCKFBHbKPnZfSQkio84Q1a3aK/xAUPiWxUPomJdah16GqZY
aBqYi+Rend8t+86ZxVArSKxPfx0STq+CPzfgvGZfJhE6xN/dtN452Xm3bqBxVBaB1rPHfiO/dOzt
UwfKwc5MWoIkzweiBJ8uz0ZzX26mSM3y/R6M+7oPfVgDRMwRQDA5wBDXo+rAfxjTAyg/jcjKWNrf
Ruhq6fAINnCIxjEFW8DoWaRrmXaAAK69C193gr026nj2Y/51qAQtZtoFxfQ1okcJC4wTaNEli9yp
jJJx5WXzHMRA4hCrduRVVcEDnE/Co3zQZmbLEXy3Kjs9iSQeokubiHM+VtMSAcVezXY88Qk6uW2g
DzfcESXyJE9c+WyVzPVHGTJqOHIpLko3xtfypJ3MP4dVCBMTny1XMTIgR0kM/rwntGUQfwCCtP43
dtVIsqfSuabk4JGR7ZEn/4j2f+4X+JjRwLV/hfxuU4IK3ic4s6c17eT7nqjoMsjUvHe8tf/aB0uz
ZN5vix4HMDOcj7Za1fOAmja4OIX82SY2M5nP/9cm5xuyIcVRksGuAcu8tjQqpB154v5bFqItXqLg
HhJiLlRJKXAVS2/2l5pzX40nx198I6kNGkcHij40Yz3adxP3ZPQ8GKfRFKvmI3nl4Ju0rbFj0z1t
SEByzITFmh+ovW646vuSjIxKbkfcYx+ubG8QSvN+RPMW8/E0NZP676R6hwWEmZeFW61BMwP5PWRt
Xrqz/m41iSqFjnr0CRqLOZaBp/c4qkpjsr2Yyo3ZEfwThuoPW5XSdaldIIGS+aA3vWmanLXUVEtB
xskHnj5fgM1elOs30NsZ8f6qx7LSGt5kRLGsHmGjfshW73RgEsMyDgchatr5Hfqi7kBdBvSstJDa
p5YAR/DI3lXDm7FYgCv5mQDXPrWJc8Gz49ptSgT4eT0XncNTJb4Sf3nxE39wDs7Iwv6uxnY5BWuL
5XOGyUejMcef4kEMap8FO0FbwYXd2dbpZCeZQ2aQ/7gyOtmvy9oo5qz34/vcOTW9RnOJ8fpc55QS
HxsIGMC2+3iU+HHrZvRN86g4c+xLhIzHi6Q2wpvb29dM4LHv2xN5tbcR2jP9EoYxv8E5B2mM8hNz
IknM+4d4KAfALXBomraib2Tk5vAbXwy0tO0qkhlHaL4gJszbSxUYcT93/HPgue3Kv/iCJJz7uZLt
m+GUmLG1UFef7HbvsoVTk2ohwCp9xWIrA0H8QNAiAAVz8ObOl2DegpeYmHSD3GOnIPDcVEKJirij
bLIBcLU1nB3X613sZxJPFNNhrBujDgkx1ONmBJXovIMuKe2MZjrTImQepzkwZzD9Fe7/K7NtOvTx
nRH2jM1AHy/cFJMSkcu+jQovNzRBZLt4zFYHm1lI0FhqttteiZNf55RmzTp+j/yHckXzMlzmwhCm
vWe6gO4+6ij7hGHNXFbzol4A3Nn0vSG2XafS6Cqz/1KsO4LkWM/Rbs7VkQEpbyiYflLRWpltbGiJ
FBgkOFD/vn0R03ysgH+8pPnBVp2REo4UtKLawl7qvtzNgrVop0rlbkS6/NVwPJFk/xXRZ9SC6e+b
Exf1ETxXgMxGnUxps/jSbuHBmIDVIil5yjUiK6184xrnMwEZtfnRc7kEdUTZqIO3qivNcvTixduP
jhz/5IIviPGngG/M0sWjwj/ywFY+xKmhhQCnrYO/yjIQU+WYHTN92MAns8o+oJXiVLRlpL4mjZkQ
nnI3PbLl2yxEsE9IwhxKu4A15qOFU0c2qvfU2R10D/fHA9mFPfHKlBI5v6sgl5/Fl+n0qgRO0kd/
AigLAKidoI5ILJkp2JESIKZNxujqkNxa3MlrYtv2Ut/P4a7jV3QN94cY82kHAqHxNbxls/XITuhc
DUCN9Au5387snEZDCaNPDxxvitm13rPj16UazWn0b4xZJWFKf95JxAkihUtNa8PFgZCblKjRpgDf
L96Z0cji2msTdV6H+uENISff0JLT7BRrMdGJ/g9B6DNvNMd8n2AYTJ7fyYMWqQLjo5p1ALfkxWHV
1C1S3NfPYM7s//HpL2Mm6BVBeuXvxefuy1KNkU5hA01KiRfhU8pJv2P5oGMucCnx5U9LtcRWrMbd
ZmQ6xmZ0DN3c8ba1l53y0VyQuUxuJ7q2LebDP0s8rB2pvEQQiJbnMDi3xYZQ9UOZ4oERpGXl//aM
Pc5kPAbLVzRvc5reY1P6beIbJZjPzActD77uCh6hfNJ63UZ+Ak39iWPHR4r1nF6UPeMYJAcMHah+
fHg/Uh1ra7uAIcRqkC5IFLLnDf9NvrKOGtKRz7h8CWyf/YB9ZGJ2jrjBHRiSAJiBveGNT3LJVtsb
JaH3yvcnZ0UJ3fPb+Y+iULbmBiyqBrXmXq7avxpYvFmP+QHOwWGutedaKrCyqcCIX63exzjmBbJS
DAR1SSX+NV/7b+qOpB1S5T0VhJoRZZFI3iOCutoo8hMMY8oklr6bcRATY+B9lxTNk68Q6Xz+FYCj
cu8oWFeyrtnPpoLqdRmbQ/yiL9KbS1ksNNR0UODRAHOT1RVGUaTLm+GChYOzkvJjDf9ourcR3XJU
3WrSh8l9j+wUuJCKrHk6ozEFZ4geEPLzfozP4OSPsMKzmCRFvK/NtEZY0EBOW1jmYdzt99icN4FX
+zwalaGY3Yh74Pa7Mggv3KxjvKLunNKYKDfPPHi3Pe3rEhyzd7L7u6jLP2321zrQXhi3BiKOhqYi
m1mIzkmpJDPYsUXkk8/z9b1Cxs71sYqJkuOrlGIAdr9RcJcmRfE7/rKM8efH1daUGZrVtR7oml7P
vLvojwKiDXETctRqMt5Y8SbTnqZpAAStYTB3nWfrA+bZULRCw29ze0GckilplZTHy5LD7X+R/Cay
4XPCKB64rHyzbvXi9DADF94yNnoIIPU6I9Ns0hpGil9ZxLZePxgRRwxChu2BkphIQ5CITblibM1k
M8jCu0GxIDYT3SRc6UYvyxT7W9MZPvqV0jobrOFsPKKgbepwY320402jMiuEFM5o/fpBtKGEt3Jq
qfEq5rj2JeEPS4xwq80cJfz5sLEaVmF2Q3vcxG1C21RXUqLYqsiFgc+MVnSK+b0e2j5Ba4CEa3q2
w504CuV8WIIdi5SfC9ty4zws1LAfwxTTwDdVc7KSy1esB6kikM5+dc9xKX0iYUPC8/40Bw8DlVGV
G4XV88FAhmNKXWaxt4vS5VY3y52votLxaYOT8QhizC/do8BV2P0hfDNZqlvAlORdeTbpxEqVlT9d
+XAlU8PPGA7cYeIZwb2F8DVonO2wjtXatgK2udYRsOBgituShPPyT+JgsFGEk0jzQ259ORshNRH0
V0mHm7VeCVnmGWLplmh5MhS2Kl7FXsKe+RX67QWQuF3Eq5NXOyiufyG95j7WuJCGcdJYm+/BynUd
daIx6bNpWxHZTEXL/1krBMNtRfM/QSy4fpmXTgBz3jZnYxOODmuetXvjL8JbKOidjTaB8QD3D7Jr
JmRQ0jAwO1zH0sdsOPSgeqgO1MJnzk+k4QqWN6l4MWWx2955fmJNTKvphMN25nnQB9I8KSt0aRgE
t/v9RwRzJPSyJAbRvughNfsMhW0clyKwpl3FhLsZh+eHbK4mflEBSPp0Dup+W6s1+Q12eVEj3j14
UYId6NtQtpYll0Z+7tG9BJNUizgch0Yn8isPjtIfd3K5BCpxRLPdeDTJE2W+a7Sr8o5TGE5k3UW0
VgQVK+FwwtmINotPvhTEVP68O5aom1vKhoJsZ8eK1WevgPIJMyeAnN9syrYUADLtSET5mREm1kH3
1r7rl2KjIIx31LU/VVc5U3zLUshWGnXZjOxWzeXHUMy2E20R39RnixOvwl/SCeOPV+uiyJOzBqBF
w07HCHCCWso1787FUM9VFhAVtfAcg5UwRTxgq7g7PReDtHC2hngc/rcqPGVhQVAdPfvSK0g/x2fb
wVKtZlXwnXX5ePyYFMotMyKJKTM32bvN5e2zqEviS0pWjic3aBeuSr6smkCj6jQ/K3nIHf6S/ikU
/NwdZxRidH0reS3nJJUFloIs9WP8wXlGGgmr25V62js1WInHlEf/uqCjbNuzyHX1JHyQPjtHr+WI
AMfk4OlyaMtnsasGTqF85yO0+YmW3tjfc92rdGY0/QFaGUfajxT7SHeFhinJFY2OW2q8tJZvKwdR
pUdvBUMnwevVtmh0enegIMwP4D4DoYejHQDOq8bGzbJ091OvOmyT675CLuW6ZkQUhr0UsQjZrzOo
JEku0nqp5ou8d2AOl6osggMPqdbY5oJ3EyvCGRuqz130ql3G0XwQioyzK4wVfOWNEwHt+i4jOD5F
rBMu9L0ztONHfLTLj7p4G7m+GYvEKTfrv7gH3SUL455NcJWqj2ygXCfz15kNklLEoasv/iCWxNj/
5BKdo4Vs2OnVYXTP4qfI5yP86EtcK7xrh7G1ma5jNq2zu9lOVq1mUn/+i/2BH8sO4ZD1RbT1NYEp
12Jdgrwxeyppe//yzcj6QgVNdtTqsemsTFzpUwN1EoRZzTwCCOZ1xkq/DihZS1CMA73WbbvSRiKa
dFGo6S85XQN7u+/VYwvIhnxgpaf+d+E+kQK4LU1/z51dITLmv0uR2nKk6OydQxiVHHOJ7mpX5JJp
o78Qe97ubYGfoYQ1B9+lVYscs7KwxNJf6pPpfaJ773lU/se6zbN5iDBIhMlimGxGqW9Oro2MiB5D
dwjcXyg5dZIm6r9pWjzEYvS6lqK+6sdueaqH9hhyDUzSYhYsenNvC82W8JvFIjVQNXuzZHnDz6eh
G/etubAnpKqjEFkUB4d/g0CsYSJtsiRidUbcd0lZBGC90RcHvnmiifrQdaVBvUDafzc1ribWT8Pf
V3wLAQuOGPuJaBVM9BfBsyo1QMz9YP8C7I+yP6F8CTule4NO+f92Tj2BO7BOoLnqhqY0145m25wB
PSMyhRTQtpdVBFouSFHdfhvrTdnGk51c+J+ca8s7M7Wk+2nCvoO9l0VXZkLAXAdA+vCH2aUcQ/Yj
jScmk3OJh3n+IWHqYUu6tnMwXNoVO0+kAVNHmmJxN3zbh+ij0mqK2n3x5cr9amgLybA+XG0T4y4B
aHl7Tf5OvEiHEitBQxHMljMURHIPx1h/KtFfYGeoI8SnUf+iuzSxhgydQoZrKB4CUnNp896o+MgB
pF9/C6UAls6EWllPGBkshs4qv1F7YDQF/vXn+hbfOJQohcqDOSjmOIGmIIGM5e0KgWlJIRCTruij
cB4WoTtvIPn2AFFY8tqBqrZKEAPs44TI5n/GPIHC4vGnl3nma8cNlnfjhTjF0PRYanLllh8PhoD9
nf0jP/C9rWIvXwML2P1x/1kucGQ7LzC1FcM8Roj5cF4cVZyeFzUcg/jiWsBP5jztLUeUxEbf9ld3
aPRnXVVq/nFyEBb0k660IyCsdQ272FsVQB+6q+3QhlGHghJzDppYLzCPdg5kY3Hu1c3EbWAWRx4s
jKmbScpPCFcsW9jGlGw0pNs6b4QI9TUVbGai7PmJSzp8mSd4fkVj6axx4C4RhN/IcvM4SULSfvTS
JNUo8hSR6o8TLHnn/vYaQfNzijkjIbs27fIe4AdsU0AlHneAY1os8rAH/LwW1GNh2HntEaDoRp72
YuJjR14Ny1QG95byScgm0Q+oM+DlDvOyrF2vrf9SxOxUeqpFi6VtmwUh9zY0NnbxfUPlerUSxP0W
QM7d4SwLNWc7UHMDPwV8LWEBfa0LVWGM3AUosqMbKIstbgDIwuCQS+QpgD9gumUXNhHYz/CkKx8r
ccUp4zDRgjRM1j0hQKKXqydsjJJvl0WiwBVvTYBO1P9eTmBk7ynw8y+7hnWgVpO0oerHOkEQlX8v
Ax3MU0TonIwLOMOhg5DGxRMkWWmoDrXZUbpcFjb6GUEdJJ2FIp1CMIK0/1Mkau2iWP1n5i+8oxJY
6SaHzKIUgVLN4wANZlyJRckB/v7njk8o5niGNVtK4IwuaBAaLNBc6Z775NFzhoMdurdpyuLqxlcO
t9vyQXEU8/O5jl53YSkHYi8RyMtWwmf6J/ypVVFb45ZYONE88md9eS7ksn44NRc1yODijxD4IqXd
GdFFN7qyFuQVBbjKAwL3eBauMiodeekCuRbv/gcf8tm2lAr1vKew7wxkpUyrZ+2arljlP5vzeNOl
8rnLE21MHIKy2XIsyXYMhmCtmPpnQiWcect00aBCnsQI6z/FEFBNJSnqcM7AUJSQlixY8seTXOU1
6PLCD/pm/bhJKhAKj+PjKDkOHycX5CMmFz7GyQnqtRVkYV0V5PDIEMxVrR+K27i1h5YeR+Uv0rnB
4C2Rys7rJR99zAKDOlLrQdZ4HEz2h/w2zzNJ6ZLfm9liXqfx8ZuFhaa6zfYgP3gNW/fve+Rmqsbs
EwrYH56IR953WC9GjA3N6Iv9pXLeTExGWDgEYPDxPJ4McdlNaao8PhUcHaX19D0JlPUi2nCQn5QW
hYUSomKJfnSOBhV5wi1739dLNIhPQphmWveer/0drNFDepX1XbpkE/7KibLiqFVIumZ1t6VAiRNw
0N1smw7sonuhkqxKPOOrOHpv3nXkS3YZ7O0vaZQl4dCHHzuRAJv5xFigIyHeak645gipmIruUp0+
nIldRyrcZVid9f6zBNcwYKFkPxMPy2BbmqN/dJP1b9CJtvZEBEihvUaJFj9WMYhSxy1wCn/eU6yY
/5LWIJTCybMiiMb3xht/GuTpus9QYnenPvvyPURLs6KSvOnlYoL/UJp1g5Si/O2rxIH9bE8rg85N
KQ3xQdgA44MenvMEUU6cA1hfXiMbxlIUsN8q8DGf0ov99/bPZmVRNIttkNiMtp8+pf1c2iV1Av+3
RwJKsCEtrFvCmsjt3njeP/5vjxk/sQPhebuy8f6AV1LMJ2+r8t3BAiyy8Y/wZpuv9XMqGXzyKsQ7
VDOx8v3Zyq+ZfwhXyhCjYxVkm1v2QX2byVbJeXTzHLJaDo8JSNOWoWhXCy6KCf9peN4bOdJHh9UR
BwHt+KU6JAVSpmsn2GVepkU7Zd74DxbDVqW+LY2dyJoVD3J+aEZJ1YiRnnWAe4as10kyiJMdg98f
2373T6sKhM+34kpPSQvqcMLvAFyKsPQXOlYBVpJKwhlBP5N5RW2pUmXu9zwuz2SUIrxe7EAi4cEM
UHIWO7qQ4BTEXecpcOHrnYZfv038k/agEnkHYll5C2gLUfte2hI3EGHB1zy+SNBZwS1zeYQAwABI
Bn0sDRNekuMoNeAvzNVnLx5L7xDycR1JENYKay4rNUkHxn4keTCJe/Mth/10PDNdNcMly7jOEwVg
ZpasWFKnbqufZ9FbzmZyB0tLXXgLBSGCA0WrLizPkcjRZCB1hMxlqRPQaz8NfIAtFI5p5ZPAs0Il
ZMgsLFWbYn8dwfxAYuvqM8NRM6njS6Bb/hc4/engkReWOaRDjpc5W0Bx5eNlppn+h0/03kLV2NKm
cGEV7xy2cGjRhO/KPKOa/dOQ/oExrkG0bmcUxHYYgLIzIOhbQpO8G9EW23LsTXnNMbmgSLxxXaEv
7/nHW5MHIJ2Dbl77/xk+tWdCOC1IrwCv2Nzd/jn9sqE7OvnWxQRFZLpf0e/hZlFVl/ebdFMbnyHu
SJLlUP+x1llfW2roRdSo277eBaGMu+mRXTgtRi/6RO8BoLeDMpqhtrLRtlsmcHuhIZBcFayeWcwT
mIELQ+eIUrxGlcKnq5sjNAmmB8kyYkTGHyeZ81i87WuFwLSmSI8AWf5vd9GAEtOcWNTeBugX07IS
vGcJd9bwjkenA8BcaN7z7fQksm36/6XheIB8i3/bT4eGoOX+/sCf2vBIQSnuBRvIOC/t5f71zHvy
Z+f455TWBPO6eGEjfC792o9C9Qd5QFnIecAIXQbNF3b/ymFnTgXpv2VC3IVXMhtBvC5YV3DmzALk
jTMtWQ7ddtfuv+cua2LOEwE6C+9OzKRo1x6bi+F19Dsu4V2jGpqqFk0DtuU3jNdBSxo2z2mXKq9U
9A8LmC6O6VvTuPVfxJEQhnZhjZ+jOoWynJaWvmsPaNNmC6ljOgAdSERJyYGo+7LgIuwH8VCWo3l9
cAhgnYyHkh0Yte7rvFN6tyn4JV0hFmMEa1z5m2rU+bqwQcJ9aip79HGUg85X+d0IVA+BurAefowN
ZyZAyZfr8SCB6AzELoVbFcWe41gfQn99rFWa9ETrDa+dDBAUBhPlZexCKqK8sbQrb90LnN777PBD
B73bLSeQJSUE80d7Xokltm5S5e6q/lfqDJHl9wH/zSKrv/XKv5t1hxRVsW5A6S+S6R78gsyHO9du
PI7EKXvQKd2UhvZLHCU+TAGJJpKcqg3dInYrfODIRk8vMzpj5US+fIK2ZaYN0blfOa+9KQ6YUsJE
IbDPafadm2pJWuNGhLJE/4u8gKTgjqcTiWEBmF/tdTvtEVkFT/Tl8vykqgU/cdUoS6C6nqh98eAA
JUxIt9iemwVxbnTMaj19V/JnM6APdWz50LA6G6nxEaA+9sMmi4IszT9TsCvZNwpKtISSkUs8L6gV
nJFo/tLP9qP8ajBXMAV8G+2P8pqibVIO+re0SDzk/nzYq1r9KN+GHuM7MxOtURH9PiAd5nR5+AAO
7+vto2BrsOMg5OXbHlsdNVXfX6/XsBScUPEW3ycMBY9WN0U0Gt3+qRlB7qOd+FSIb6KDYwFMa0qe
hTWrJ0FUwWTMwoSuYc4OVgL57ScdEy/o2wn77jSxeyDUmCwxLqTv+Ji6jsPr0wtzj1hyFXIS6mW1
k/gEfZdhYnQCjaqBzBveE+ygMy0mPqwAPSgFHYTsfa++uN3RQfCEwGqEq/p62iIPQ1Z5ffxNpNQ8
b8LZYlbOjMJZyK9yAbQjAJAYlVI70hRUch7sIh+M+ltT+HB/mK4ByhJ9J0B0fRwvaJkAoMRX27V8
cpfiPp0AN1BNy8k7HDmjgrZ+QgTzKOhVSPTZn+74IZ7necAIAqxaj40ID2T9DRLgEa1JLjcn6jBG
aD4Ey+sw1tzerJnfl8ysrmTRNW1WwP7qRXJYcUzV26Wf4p8vD+Lx6hJa+3kZfkTdrD8F4YiQW0FN
iMhakMZEjHcKMMVT3W+5p2NKJN0xviHovRsAItNcWd+/cp/r6/kbqAXy/GKLWNd7ct1OOwCR4rHk
QPggQnupRkqw1SrDB62UMXyUc3cpQXHxRtqBrPap28NCwoMSxF+Z83lOa5rNfwSZR9RW3J7w9zu1
4Tczih6qH6dWVn8WkkAvRgbUgL60uCJObvtYzQFzgQWt/l9KFjbK38DWLcwGqzrmSJUaQmCHZzsH
vsezp21BBk4+P0zWccY0IfOfwQwj2Qfia82rxTCd1r4AshTIIyvcS7CRfsOI5817AkOBlJ05R7/h
XWePJCOrNPhq65mfebabVfeotViVngCn/M5kTTPqs+jkxgstXGgM/+htrTZZy3QjG55fBUCL1i4b
7p3i0HCvx/IQY6uGhMVltBa7enjW99dJX7/kT3D9auuhuFUF5/MEoHOCbUmOwRLob8WAnDZhjGgO
4ejvteIT0ZK9iIKgwHaIjV5QIM62nVA7TL4/wIjL+idX+qOTuV5aclSwS37QNwmZAaWs+DXLSx/D
YohliddLXrfpVgSnA5GKyCMH+X+tqp7N2HVFFuTYMmA8TqwAiooasNagvsZzhbhul3hBNQ8fYhdG
LCcEERcLyHhbCgSk4BMRdNUrgkI6u5bGIXkym3XhwsMmzKKtxubgyHJJk3pgk1blqffN/NAe6QhC
LB4wUoedV8HWb+pDyE2HJKImBsBfl7RZzoDKlPd2cFPiuX5jOJ4/bigDutzrtU0e5orGatEzflOg
dSAD2YLZewbIVo2Dys2OwoltWCryNBvV703JUIZQX6ac/vwBY9Tl7oUGygBsUXByOC5biJGXQKAf
BycBwLV1PROWAi2wGrd8chBS80t0IcijcvjRwX9FzEsf6Yf1dBqeIYkEOdFmBEOgoLaMDj3wZNr+
kJ+AhJSlNnKLpBgbp7jmvL72yAEGW4iTaycdFd7abT9n4mmxRUCAElu6T7Db6AAmpn8+Mo2PfIqB
qKKmZwwXka/REVisvcs7f55votNuYIYYDPW0PWlzbGKcBSL8mIP0OhxuwI5WcwpNy2vE0F1j0b4G
S1dWCLqcp2kLeLwjGWfGUWxkA3Te7p1oeoaBTftYwKJUE3TSfO9svREQdwOK/9CPZlmoV5rSWKl+
BFTHdCCDowJtT2uGL609fvG3BaOrNsKbmCiGDDgPIBkoqHWb2AO6CffznjpGATudfu6jwmkMz3QG
yyUMCAoPWNZLM/GBIbDz2Z55b34R2S4Fsjn8XtM8o4FQpcRgktRQuNf6Gk5TD5rAzQPRv6m5NUXF
T5j2xFAGjzuUtY/xgNmEe3atbLf5x7SY2xckmBb8CakTtAr/2JbA3MYcI+KyYdAyAZ4x46xoDZ6j
ZjrvGDQF/1s2rjrI2dmGH09pydbnYP7DtFbczMR31gSbO0DqvGAX9JfamnM5PSG0KYUNZUpxB1iD
guaWVUwQQyY27w5RtaO21XT12PUdugjqefu2ro7OAOIvbgE3ku29Fe5VmCJ8+sUBAIJ+bRhY7KTI
fLb1ryBMIKDiUNf+7HmcZ5tWE9u3A/nOKJV6QUdvzWZaVu7QUQaDpy/vYRfMHl69DZU0/8Qg3cvO
0I9fvXIfT57MR0lMjj+dY8ZPZPMAe7fbrQxXb9y1EAyBnHJLMmBkx4uMfruc8IFf5YP+yy+ZpRcR
Q1zK42d0ggoMGQH7bQLnLz5adbW2XUGPfVxEkSOHAs1lHA/upeHZbvTznalUMx9fkmnY4Am96+jQ
NNPpbx+8I7sDvE4lnCxca86VNS5GEb8LrdtH9TGCWO2e7HRObvA2WuF4KCcve84tzXVC+kFGonve
Xz52Ek0l5B5bV8V30WrIV/lbXJleTuvpu+QoTdkyhA6OvViovXXd3hF9EybedW3umHW93glPPL35
ux4/y7wp3hIrUoh54QjHbJUeDzs6URMk2QqiKEZHZHzIehwSviXgTuOBXW9RE3ckUul7cIN58RfM
bShPqpiNNzhu5EmLGqHgxDIl7ymBTrrTSvqGD+W99PdDxHr9+O/C+VVOgjpxS3MhyOfVRbONRo/z
pK6CIzNJpmwXwQBn4lrIEXooeb7qQdwUVejSBUaYy0njfCtA5sITjf/5eXLIhbBPa+J5NfecweB5
YABhzef1GbqBqM2uvycFCFd6xkLqa7kmYrRXHEOnwMOCnstYMNbCaxKs8t9Uv/6axOYJWKEjHcy2
51frh/vDsvcPgKm8Fek+gk9XlyQlc9z8cOwXWqUkA4Rp3aiDqjzknoFDbHemCB8L2F448YANx2Qo
FeJH+igk+SjilfAU/4i2B7sk2INsEp9FB5Rv74ysJ16AcxPFonNy7rCV52eMfFUiTwxMSnlYJZ8J
XAovlUTjsupFTdn+l3wyBXzFBaNzrgdgu1juenZZi18Y4tqZ3FtxCSitLExy+RG8xmnkjyXPI3xJ
v5lKamu5n6NpcBPLqja3IGAax90GFIEw3y2GF6ZcVJ7VTY8xL1EHG58FtGA1oZs4JtHgD8QBwJfl
GhmIKDK+UHsn4z3mQcyjxU4sEizhfEz5+L1goxmlICwEqafD1hOhTT17Cj5kRaCftB/eSpPOZBQI
gqrv8Ijaj9orsPRhXqeNksn58z0ygL+KN1sofXhtlieBn38eLIDgDsUmeguE9loMpKa6L2geKUeJ
7sT1eEomtjH8csVEpAJHVLuNoYRgDIMAvecVUKATq6PXgdoN0SCPw6oDJYD9ISpo3UQONvuUeOB0
SxoBWJN3g30N4YNDfrlfFFMz31N9QjHbRFvEewmufz4+2grsF2H+GqMN0/YLBaHo+S5tlAP+GIvz
ysqiDbLpRGM7rMsCiEb6QDuDcgoX34MP3FNRCtu0ClP2EVvW1SopR3OZFHXWiWL74F/xjtdVe37U
5S3NV/nF0K+28LgIKN3AhWYUa7I44Okq+A2nsLV6eX+exv1LYOSsXJ6b/t62vJ6/uNrzTe56gepi
Eyzs6WXti6tzSmHi7H5mM/VcdpKUg7GdSFYxNPqF2L0JG9Q9L5h5vLmfJPoIcYh+BC8cVxkWEpdv
RxyXaxaj4JKscBbafnsZQ3YG8zrfv91dkcXgX98itgklQ34Ej8JsdHlIRbKlfCZpZXFNfGjg1i9t
JyVaLNkKgytkX7+tCbzp3OJO2JEDIkvz1jMHIrCPEDQ3JwW4MJ4myHN+Y2vEPT8uevPg9YB6VnET
J+8+ZCOEcTQFKAmIuntESfnz8C33+YIYdxH1oxou5DfCbaiCByTde7e/zIHqNZVRSdsY7Pylj/iW
CcWS82nEj4sWZG5ypxA/wkvd8/bS67Ffcc6oNNv2vHhu8wZtfWOhM/1zI9z+Z9JARsB3xgJDlCVj
h4qYj1CbzTtDxu9obTbubx1hAZj123bbu9Dj4M+NlaMPxTVk1xjovJVqVrhRWBzAJN1NMoJqPYXO
ixDGF65iXIArp6rkzWmYnbtzWVhPPuvhPW3a6FG1X5OyhV1IuUg/jHaWCJPh0DOBvDXjjSwLvDhR
mPdATQoKMD04VE2T1XdXJOBNZFhcmywX19MdciHybNqAAnGnJmXlqJ47IFgYb/aSE2Mq9Cd40EHo
RhIja+IwZZVZvIpF3WdSjqgAUa5NIhA+J6aNSKij01cGqNNy8DQFD6oMWZ6X6+uaVGIyZ4G4kYAz
50qjxDdw0klBtBqv2ekKEWCQEHvoZXkxUuvCwIr8nwpo4iPB7bt6A+pBCwAbxQsSmFSFOJPMoWEy
eodK936Wt4l20d+gt19pwjdm5oe8v5gHEANvVBoUrx1ccptVJuSVvHAH63mH0tFd/YMAoQ6294hj
LasrafXNfBTnE01yyqHootXjqoC8RK2YMhaBdhiMVYF5Rb2kTpFDwf1Zw+mcnrtTLucAF0Hc+utE
MTMyc2Itn814olHvkBWshLUb3Nhua6x4m3E5sN8sCWeKpW+cbJlTYV4YwNAMG/CrNBvdcdp1UH1d
Kl2yXpMitnj/KBh6U/mHK25yvhMuyOJc2uq3blkfG41N/+5+qzg5lY2ytIjhp0eDLvKauyuXlkFt
Wmokb3XqNzy5dXFySKRpY6AZpOXZTLqSsVbPnRMYdBre2608DLL1n2iwgodqk/ZfEaKZsrruznAy
ZO0O+XSEhcni4gGWFSX6/UX99GFn58VHJOyw3yDgJvdsWIxFfekMTaTNJ3FEsjW6RrqOeoeGPbhM
FVTOB90Zz7aB/VI3m/eqlOIg4hEgX7jpfjNnkRWh79XWUjY4XiyGzCczXpstDmVsR+IaRTdWixcp
nFqE0q++I7Uq2bmfEJxHUZnzgQF4ODZGu/XN7nuDd6+ebdbbFuKZpLWXFwEbf3bBWJ+K0zDgmJW1
Mew2FFVrPxJOIL1D04nQRH3I1J3zBK1DbCL+mYnxhuwwvEWPUNO4CtRbp958G4OEASj5jzblVry9
z6U6P+A+FFEQ4wflpi5PnfxxeUNjoKQ1lv78k+0N9mynwy8iRCvAdWsgFyILwvu2TrrE/pBsUJZV
JsIdbkQ9Rxw+IKccJKOBkdJqyj18nPunQj2NtrLx6t2ACcpPoO8VaRO1fNwXldxGfRs0DO8Hl5ly
eQqhDYCLF7RM+lX+e6mOfe/FJGLqFNgMDMq1nrt0WEPb0q1iCnKwRhbHfO7Zd4Ytb48qBmPTKVeW
RrppMYqH5TDk+AwEYXz2aAG8HXh7HMglSdCu46ygTKtdwtwyFjiPVWYtiGG3LNLs4q+PPtwVx7OS
B6f4dl2TaD7ho37hzfcuxPoiGIMyTDboPFGpkG9PDHF1Y3a/DTQWUrTHdSloSoSQX6/vE5YO0zJM
bz6gGYvvgXoi0zqGZCmHLPCUdSK0nARuQnxnQ0/TKnDIA7M2vgv20E8VoOyRVUIXE5nA0rjBMS3s
XnjWqVE0DfmZAd3uO4G8oku0iFnZRsiD0A/v2ZpM6NXOD49fuJM3d3DOAnrnq01alZ3V5nGxvNQj
YjIecYxCYM9RxI+co7hewk/7Vfo1Q0mgll7Jc8mIKdF95rOA5aDIYqChpCzopjHeEtLuxRSVdo3T
gqWoM/3QC9C/RCoq6i4TbCEgVoCalJRlpSLz/PmCs3pLebgr9TdkNrBissq9lQ1Nk0uzgTogLFkB
P9O2f/Nr6IGUXPRXqgUbj7S6XCWdrMogIWqxosWpOlnc8Y9K9rRhKuJcZ05Oto1CGpj72mcqUsbA
4SodGCaBAV/bUzT6EXMeIDMVvbKsamQuONWprKyNnsxCFcCq5tH/gA8JHewEO83hQiArFyvzY7X8
1r/QPK8pxClmwhvkOukgW/uAiJyEXG6kJoFzRJNDm46ik3JvW9RYzNNiMKDsG/mLEivkAM9q0zCR
X1AEfw5n0EJTj+DiUmAwBXDlRaXSar/ZW7WyDZq2xrMqCh91lrQB3NG9/8QWLn7+UieAqn5Xda9o
Ut6AtQLFaexh11CkRAPztyRgFs3h5tR+R/FuZv5PGk1Cau9hD7thRA4ASaF3/TqHqiAiURMxCCz6
NypEe8oAb3kC33i8vWbZlWEZb3Nfhc6hBawoFsVzxx8gNxkcmfU4qP1dqdUfQym3qbyQBiAr4jEc
99XliKDln/eDZf3ON97h45uzT0zmBX7qp51BZOkwHUv0GBndaM58ejbKz8wDU7AA9m8LqYPJF9gG
PyTnLEfEt1jkYQapUDd9/gT121Qb1fVdjIhdpjVeQBr22teQjKiGxIlhK3HtvUPIAlo0b9qM//Oy
Gekk3wJ9R/Wz0BUIK+IxV7VtpQ2jIC77loPuJYqYUEnjMURBpWtoDdaFtqGaolyv9lTdPb9Rr0uX
zz3ZVSDkn1XVz12u9NpZoKDyxzu81WcHzqyjNo/IhI1rsv3vJGvfVHX3VvHRH6wxJyirfClQsxDz
PHq5lecEUQagoVOuT4Hhoa6Ar6uTcRitcLLJCh1DcKtEEkJLSqjEqAyp7+qOe+xC1k4IohYkCupc
Movkim22Gzw/L2M6e1HhLuHB0FH3xaYtKPxhV94gVe389y76n3RUwhhziUsHSsNjZypnc/CZB6LZ
r8wkWLtWZ65LzTQdHYU1Vnm2Qg8JeVwCc6U4eAVQ3KyQv4y06/dIP7IOAE14PwDoCluEtUcw0Z8J
YYCvFwxd457gPpUnK93vLK+b8njGBntK903lgcynlasKkOCg3/gDqbLfMI/0LT8rdrAanYrvtT4t
fiwssk1urd3zTN9jltitEG9X6p9rICEz36N3v+jH8N80nio7O1KPGIKRp28N5sKUV14+XzaUB8gU
XW5mmGMbgw47TSusiwIdrX96NXFOI8kBMCXIawhEFEogBSz9C07+0cjQOVIJ40tihGXmf0smlG8h
GdBivn3C7u8rjeKd/aB/ThYJOZCLTtPmexgCG5xGJhysG8YuziqgwTaYGHNRnTbIdPSUr5p7r1mK
ansGa/i+p+/J9WdOlZMh2Ue3+0nqEpgS0oBkFJ3EtIk6ViaG3uErSjjS8nMQg1LvO8NwvGZzlMK5
iiBSS/AkrR1hDNmfd6FyQyOLfHeadJw3Cdm3X8i0KAU7Ko2Qicjpc5sP61wvVjTx5NB99JxNsNSB
qJxWFdtLGyAeCvXqauAEhp2+tDT0Yr8zewLv7nZLlz0/OUuvYQP1hlNZD3a7V9PDh57hxkyhEKtc
/FQfJaF7eY67hcPm2wGN08JeWbBS61oKqPyIR2+0rE+bcCV4uaPOP9m3POtdNmE0Kc2RILeN2oge
7ZjVrksoIBUIMGdHXpDYYWvFHkkz2CYDm4ajGOgK37v2FgssyzaQIhZ3xOkCAvHWNaaprlkjVOu4
7a8uGORvKun3sdJRQHYOoTU5E1m1pagZOk0vwI4YbJzAkLaTKYWKgMHRXLI8VIu/3MJQ0xiHv2SO
BYePS2gc0t6wiKI4RlodZjnjuW/EMgQToToFUqcFIerShqkk6YMwyVs2gzEyJVhUpMWMAVGfoWF3
GdUc/7H9SxAFjfzyqhVjDQN0R1XeW8GHD5Z+zDrQkI61hy0YaQ8gPu4oupyi+/SOFjYuBXvVjEhP
4qbf/qJr3fKJpQ3qlubA2LOLOMz09Su6yA/+CzdfTrVKt9Txc7U07Cuq0U1Ddz5xZ2s35d9faHRE
zac520rx3UrwAzGdGe1GGeTp+5KQDLAU1DDwFWMBAfYQIPcz/E78yjy+DUo5nnE1pz6SMCz8XnOW
GD93nKRZ7w4Kj2aAaOJQjlLxzithdpeytaTC5OyGv+btYvF0XLkNbQqUlahxFQKbjkb/HO4x5RjX
DCJ8xZivpvW8Ep/GuI/Attzhi8yk3F+dVGjaKQgORmTNEhEphbsoNpYFnPsDHlU1x/v9jVq/WO7W
B0OsvU+iTXYbd2w6VwfZqU5q7jCD80Hfw5LqkCpFxeQG2EyRMBysQY+0Pvhi7ri9YG/Mi2sS8dsR
dpKas4saBe5G0DsTHm9+/SqSNiGgyJrc6xFepIIAP9e53tTZPETxiPM0u5LxNHMFgKh+ACDL2oJa
nRx2Bx1Zjsjjjcs4a5bW7EQMTeMpn8wA1ZbwTzZN/Wrk/59Ep9yY/vqzjBwCw5xSgpBK1ZW6Rkv+
jWWU//NpodCbLRhtOtpU7WEo/GcOOrYl0VACzNTN64AnpjJYL9LLX+8SM/4BbD61BNKUNrlhRMER
5DVCb20fALmXzJ9YIp5CpEgKxyElDI3TfLpLOpEDXkO5gUihY2yCyaBE/2aU99GAF9hGMVU0ssHO
voKhwg5FqrRTNf4cMRfalklngL/GJ5psuMd5QJSW01KkeBILn1jO68TTER+ld0C6w/7nZyXW+xHc
+O3kgXrWSsoA8wIX9siz96wpvp5oQU6TrQuW+a7HQgbD9V2Brszbj2/ONOT5Oh2D6iW58rHzRpNS
VfhORSeOCml/eDBGP/nxK7hwto8omnIqqJeZexCT+KFp8i6Gs+V6Ysj6ZXbt93uQIzz5/9wSZVtG
/TsodBdxxpw179hzn6JLC/6VQTSQmVSSgagEOFJBMx9flYqlbvWh02LvBRMbsQL/ATxcwTIwREQF
28rmGCcmQAY5/YX8Lpaz+Lg6mX7p0E7TxsID+m2seCuAKr1DLZ1zKb1vCAf7ZCebedHt+gajsYkL
FoB+KOQpjBj2octwc5lDqaUUdEpf3dCWNuAk4khYsO6nj1PKr15fPDGh3zr/XR9OtPSQQni/sHIL
UbEHGaEalaJuvY2ewQiJlUCbD3TiJaaxHpCEXwgyyk+jn65KIiI72d3ia94NhAxCOL4IJlEWsX8+
7YarLw9mVGJyJU71lLJUjjlNm2ItfV13L6Mu9wtyXS+msSEH5B01TsBgIOYeBM2CWbuj9phpyEif
aP0FaGH/r3PIuhtI/tpsxJlogzhvUnR0D/QiOJ35D+KVi9KazHoOdif0smvlthJvHXuhIyNweeoG
JpCKrTmwvd87KHqRlIHUCvxnopv5m8jSOB3k/p8w7uHbwNF50ql4aBUQOtjUGYTswnhC0Awpv6sg
vnhJGU4tQ+D18GlHR5fGoY034ozigaIGZD2NrigEb13MIau42DR3uXK07FB5cp2/33DxALcnt9QM
XKxUAfkW9QEo4z26ONXmx6Zrp9m/TKvbPATgjcAM0YkeNXH0bPgl8GzSdOYGosyG7i5sPtIHIwJO
5jPG8x0+bjoW0FKaVGcx46jYhup3jmKPYjcM22U7fMq5kXxLZdjhsUef6a/DjENAh1HsmjeZdpmr
08FKknLUMDZ8X69YNx8t8jOWVPOGMV1s1XSo1yv1Ngg9ailIMwGp3Pi0RgGcnPYrgBGq2b+37QNT
6sI+JVZBmmRiK0etNBK/vHeaLCHFeAte5YJpb57m2f7DrTWxuaRf3YQJsUKm+g6/dxuoPFrTEgmv
UmS6yPty44KFozfhmycmUdjPKkI/9sn/tMqtktUyeWoKI1i3sDwiJ50xrLCbev7v33b12EosmIT8
rF1Kno6cWvUQJgzW9wP8aDDvZAbbzHnhnyjDu4ZBOm3j/p8vgdqajbvLXMAbxjr9d858Mkzi1srz
o2Nid/Mj3oRmFtfaWjDuoF88Jm07TtF8ETK8HzCFvwhVga/2lPa6vzHF/qS8+vQfJiYXloJT90xo
rXT9Vw1jckiesX2mmsLeYJjOviWEesJ4qTmoJEX+r3UWAvlH30vFLnhev4SxtJ0BKnd88mFa+o3g
7U7zpIWnT51/So1Dx8hNZKoVkQReJG3H0x4zPj53ENFJtCG+xT3asO+rArPBHql4w0zUN7+P8EX8
tPQcfPmfFgBf/LT3crNn/OarFzkSgqG3RhUrg3Wk3Af3pL1VPULd8aMpxQtr4E46UDNnPU0c45Z8
I1UOj5+WI0nvDOdZp9H/kONEg6dDXA2Qut3ZiB1GFOgOKmUB5HgmTmzXn/50m27LVMi9dmgHc7a4
fmEJ4U6i/mN+ElHLRXQDbpWceeaK82pbTnP1vRsMC4q0p9pO2tMklVrdTmOYNbW3nJ/ekBhS0qZU
Ys094MU3qbn7xdn1XqpozuxjcRy7I8fmWz4QeA59uzrly4HcKdJLKop1n0IvB6r3F7Tzygb2mD0P
0fdrRh3mHfdO2/BTFsDv8BsoxFf8FjaQRefdpygipc//c+u1XzL5owITQeF9Xyai43m8IG455ggA
+Y+Y3CbTlzoa9KIVkFqTUb46OPqRFLC6ANkj52fkP0wykCpud8DJICDjSjQFycMK5A779rmw88Mi
Yg2qVkOuUemNGmXdp4sEWj690TX51QFdY2M1g+LeHZWNhzqiDJm+1NHvgaj05wpwjv+KdNjUHG+W
9XQi+7EDPoKJGmJKOu6SK9wNxC+DKqsaZxD5nkZbuEmS3txqY+H45uHj6aq/BUIo0MNEwD2r4mks
3LOfG4bQfFSicojnzdyNTFVe52r0R+KpOwMnstlhJlRZB3GwZtba4bj4FuwL7HcSVV6apJV1JQWj
AZu39Zd7L/MYlTi/IdLqOF6QTPgrjzfRrgHOT6RkM/2p9k1h7LzIMvWiJawE8RoG8D3g36Yj9vSS
0aJAp/WhT65C0yVP6cspaF2o/5P8Kjj/Kr6U3E2nDt55TJ7V+JdrCZcd8TiC3M/psEfhMlwnQGe1
pKPny+c8icPELtzI7q2ST/cX4bLBhzcWbr8+GsmomKoq9o09300O13p8LdiWOZCDQ4/ouPcdRl7z
B2YnK22WSM28u2CdabyRxdg8kC2UKq/X6kLu7xsqJbbw8PC7s0gdEp/We2ij/kZ+yGlQoScKXEn2
zoJyVcnlrks8asJK+dJbjdxuaLWzkMny/bZAgqTbRZ4ciXz0pUOdsQbnQV5akya1lk3xNzZezJyr
fLB+6rRIdwm0Cyc23AU1YMjpKmPSEbnaHJECQoj2Y5OIE/EdPJqUKR6MQWoGJq9AvoARhhTcyUk3
psAWS5emOVw4YS4AvsImqfvn8ko6nsYslxiwPAvh+FVDxeKjg+OZAJ503uiwFX7LjpNd3BTwfujx
g1sRvZoRJcYWD9Y9/tO0G+VsknFM0GYnmhBWFB74jFgLYsFmRvRdumvRRlizA7Eq1kSe+gmzMcPu
vtuhT3C5CmOhQgkqqphQk5Qe2O6AZz89R6gE+6GC6zIUp21qfn16edOJQrFtiJCDVJM2B3/OPF8P
P7wyDNbS5ZJgEFCCcJ0QfU5vkQo/6bPmwQMYBQd2RxlEccKbC5iTxL4gqJOiwaSrnuReMr4HcRxn
HNUpMmJEi/WbXLjeP+qkheS0q4iaVWj65GOPcMSfc/mOKCwJVGP1zqyx+I2FLfjU09atSO1gp3At
AOgIWOpD08g5DJVEgeYX2+YAyCyraluZSg1TGs9X75mkM+/LLVg8g/v45sjC7U2NI0DQqFzIUyzh
1Q0TCZQ2M5XfizMNcSZ7Gok+1AvJWRmkTvwXc/yMarik0BwPfk1IuYAznL8KCsl7nw/bE84FXmNJ
eSj2eYRAK4JLQ6teqd/AQ49tgjWPAJnPXMS6oQFdrSjgCF+jgLiJ2LHfJQGOFtYrG8kBdZJwjtLi
t/cgOBoBs46VOq1g/HVtCemqAPcFDSKsqFpW0FI1GtLPr1GKHYDyXwnUHQ1D98d9LosNxT37cPF1
6PGYAj6kDqGnohHQj+j7TFaL7P5pVb3kgTtTC1JUxeuq3MZLS/if2fgcl9YbCb/67GHN5dScsWly
BoP8Xw6h9cuoFE/tq6GySRn/EtDd3B6J4UjVuFaghjT4f3Xt3xYr7PhSqd63HhtzVZRp2V6xtHer
M/UgfgjeMBsDSZkACPVEoERs5QkywPkJ4oK82qJXJxEBKD/DAZSc3dYjQFc8dTFC02FFgXA7MCH9
9W1m6UkNyZXwhSw6SDyVpn2viN899mp9G97F2SaU3Gi6iiUIaba0L99FxV3zewoYy5xRfPz15CAD
PnXZ6OXsmqIiLwdnJnDPf0Djx5QHdKGhtM8MOEGvbGuxE/Os4N5LDF55YGhZZNVgmxRWzYbc4mQs
KWYrEfKghFduWcSYmAFlo+m4P2n8dupccQGew2TK94OV4I36bAU6i0MipbnH6cmqo+YCqJvpQ3kQ
MKNztvNIf0Lu7PNvmkX4tsgP5ajehvgR/QRo7PrMfCkgVPxfvdfe2U2wOd0B4nytxa0+g5Uwt6C6
lDmfpHuNfW6A1Xh9MKz3c7pm4B0MFgjQJbuBwjHLKFaL5j/sfXNQyJnOFUD5FHIE3AX6UhE0HWEH
+ZJRAEuTkeVMAIypGe75YW6z3LSIfHipcWTUd0T1kL7Agf1Gkfv3KFTCaYv3gLHxz1XreCsEXqsm
KX/p1waG+TxslSEPuWD6O+bo3lKWjT5TR59b4g0e/xIbqupP2QvR0kAYJcvtxqqqwcz/nuryogJW
NNYlNOavzObilUSRaGukOIo3rgGp/CJjYh0OPprgn5Z6kTbRxXM7I7fWpd9C0HzD+fbfu9ciMqY3
kb3wj8u1tdVJjqiPG59TMR5h+dRtVr29U3FuyjOwzTV+gXNTDa0UyEnzRAOX/as++45aHoXUhEw+
uiypOM1q0etA8T6IsS5CoQTbNf0xSGNqOJvVZygJl1kp98RDeev4q575oNXRPrFyj2m3iH7rowwW
LtqUKqJaCpAFu66s3sYfIJpHEoj7k/WVbOYn3qjoXY6tt/KUvM+KkV97MEKCbIYCnvYJXwQXsSqN
iS21IZmarSPEH38E6IKGzDxyxwkfAsSrybh2oENwSJxI6POsjhKzovXlvoj83fCk/WiZyCRvyCd4
FMRg6mYcVi8r4tjGWZvTNWtNRLdVdCRaFfCzVkBvzQsouFROVa8lOTcgv+hiiyJVkSddP6hd1t9b
mbH8aLeB/8S8Ezkacfa/ZEixCVS/kPnghJ7KABDOkNFM0rVO/WWZ526lcJWqfe7q1N4R2YEjFYqk
sEX55aRMr+uMW68Bm2JsIbVEyXwIODK9/IC/ja/yRjQw7PihljCe1P9eVYOZG0DUrlRB2naiLvg2
lGoxWF3C1Old7peUaEjSgJsZA9FgPipAwEu70O+c+uWPUGd8qsQSMsq+J9GuaDiZOTi5JYIz9jbw
zUm10aZEwaaZLRsBjY8UETTlb9h9H9GpQs6CtOqAOCiJgRCtI0T9sq1C3HIO1wTubOJeDjcCQuqE
VzgjZohJLCx2DAPsGG6hgO/3DOM6rahMawPXWHSQV/FKS12hn76JiClKz3fRdXfRqyB+O3yZhvkL
GsGjHmUS+B5MruSrcrgAJGNnWUMrOqW6M5N2HmpPuPQFAOCrk9qEBLFiUPxgvq3lPZADxu4+nN48
NVUbOR/9i02hvd85FO94orP7p37XsBpIZZ9wlfkkAaCCNsiqqjzyXSAnGiNbaERTLPEIV6oKJ4yK
ZMp7ML0qwkhl1A3k/JdWrsnzma33h6aRGqzrqs8Lwye2S+HGMwBkoreBMz3yj8IBuLelzrnnV/cU
A4K98nWz2+Akcdh18gqB183TVC3uOpyC+YShvWK/aFBh8GxBIuGEajU/hjlMhrf9BzMVbP5pzP9h
cStQQjXdOx9zKaUCLeyS7pokPv0m+yiWI9V/ZYOp7Phlkk+xEwscBJdbHXlDok4MEHFIPx8+INEI
/sSqhlPsev0n3wg09VldYc+c7sp8bpOWeJczna/W7m7x22n/slvFV8mEEFFbqoF3ocLpHdomhNxr
UwBLEDFADh3beOljIfHPY3FqCNeAqQshYDCD48JMvFhQrVxNOf26IwU0fDTUDuAl0wdhPauiU/Ay
SO6srg4ltMjkfh6C0g4YBVjmrzU2iuyr9EwsZflVH04GQzT3RTEKaM9kWcxncbswBNPJDHMrCu1Z
nW9mYDhw+FAbUO4C8W9SqVoNYz/9YSFyWfKxCLnEiyLnT/S01c63QCCu33fNAUz9jCbhAUcNa3L0
KTNRlJRF/wljGee+PMSH+h9hgOTk4Q08Izf3Yh1x4axMxR83f323JW24BenZvvu+ndwf966KsRK0
dQiG95ske4TtReQX24FMmBmJFVCrEbzN8GdhOOL8aqwZR5Q+VP4DOD2RmdlJKycb4TXxNDMrz+/x
nqdtH7y5SdN1rp+ycXZ3x0fRozePkV2+k8wWLZp+cPQ5QOCcig0qHzTymgpRL/LCbDp2c56YWSXv
kNxPkbrkBMPV6MQndlEnOv7L0ne5pxpmu8Wiso8dvCwchQTJHbzl/uWURO4/1ikRSwE7WyCMtnBP
mUL5LHqj300fatMnFj89oZpUtEi3ZpPvQOfFPrRnulAtwAC48ASC4zgDAOMkK6usaOl09h6Esrw0
bBh62zFFNHOgl6xHChqb9zcgyNrRfrKyHwG/oNKbwSCntrvVReDlPhSEcyiTj9H+7aTwnXf8bASw
GQEYXqXPwHpCFCGp4LVqOPyrJEkLWRfEtJc9owEoZNMVkznhQqHQlpplFZ99tHSGoej3kW9t8gt2
bWmJf4DZkbCmW/G7DMjsTTBMs5L9ueaC80F2v7uCI19cI8a/21KTpfSfM3k8GMa6j6B4+ycefBpL
2qWbqkmGMXLfilhatzZbaW3w/8gBIt7yKabSL8jL8/nXWpMQoP2jByA31FDlge+wkOfdC8Bvd774
EpsHlspzHo1MqUXQ/BJVIuSqUWYjtFIsTWCyqpO13Nt4tny7MomyrTNuYqochoLa3cUkfea2QUZg
aL9b6k3fT8Hy6LvxLc90I12DXNOiQNxVRzAyez9UwpzxFSHhH1uANHXFCjDGkASCltEsYnmX2u/J
y1ZgL7ttFtvxyb05OXgURtxp0fGOs9Ywq/3Ygc45h9C8yRCDTemRuAWTz+yFKyRFKR2mdatl95rk
cq7x79Dzl5pPJgyqku2/YYOs9UrZ2mln+zjcmzTcAOVZLCyZ5fD/KPvE5AWDHZoRJ7JfqLEB4XOe
yFCVn60r6rfQtXahLMWbhMNBrVSAvq/og9VQAWmg2YEusxXgj6IPMLUnRmaLXL7qiIO865EVXf3/
2eHaPMsxm6El6W7RLl32XlWpZz0Ho9z1KcaSc5iBLKO51KBpy3rFc8Iogiwkdem0aWfnIqX/ZkdZ
3idWLFuib0AjHAwZWEQgprJOjo/h95aqmafHqUC9/CIlQNrsTM7SkHiPJOVePaOPOc5pKvDxVM9M
y4kBNkEhi0ZYxf/ZjQjLWKWThax4ND02fdq6zSSTzrUQponI9LV30zGbhuyh5n1mKwaKoqkEBtOr
B9jdOevkrL0pptFOybCVCe520wKKmOECspzTLOTZ40JTRYB/A5+3JoCDflHJvmQV2tn5FKiPaFRv
NZy0sH44AUmSyPS5Sa2Y70x6frCsSkd1KSi9Nas/+y0wiVXckm2qi6akvquxK+4ytjnoX/9ZTZSy
n6QYNfN/zNpfVMP8DTyogWCiiop4h34wtT156c0JbPEeh5ctSEj54BQ1qF+EVqtN4yHBDwnZX41Z
xFBnmyrDAKRcV57UyEK59FuiG4dGLijWJoqgOtMg3Oc2SaZ32QCCbdTxKGAv3GdLr+GklPyK46h7
rjhrwU5oAL3pnJvjs2gfa+1A5nYhVtAg5G8+eVlskW/HqHPjbgaUsWpX/eHiXI07d9UELeEFzEqh
DFDL8QWPywKn9Lsj8tBFo1hzHmeFw5NloO2g2hnIfFXN7yuCiBgYuUKyMuDVZPWL5xgfFFdTqb2s
MzWmG8DhVKi4RY8MI5jPyMPZ4q47bUUce5G+p28OmK5l9hpzH13EBkJlNmSrjTgXEIoKriPRZfQ1
JyeUPqMxfkC7GvBF1gRVTX6F3KNqDetCFiYjEwaw1RNvrFVGbzLGDHc/R0wWbV70j7ne4HGpOpax
M/l7RIiwPhiji4DZ/MtVtIs8JMEXIIHtq2TNJUM2HSfxIdHdZ+V8ZCbmqjh8teda4kQKOuK01hPx
/YTd3mQ6oZyBAVw0Lkfr+03MuoBdLxT4NQ91WhH5eH5tWal3jJNEVcpCI+eUfJ3AwIeUOb3Sfwao
iruxwWXpu7431NczFemCwU/sM1XPy2ozcbX2stGNGCppoScRYZ3HsB0JkXbwovgLB+Omf18v5299
ucS3+usuh/FzyBosRj3bplBNGFru7FnCkwfo1FXqQQl3HD/PWx/IOMFBeNbtsV6GVLlaZn6FRkeZ
0rYYTikLoO3+HlJ+EeJT0ozwOUpTQ/O7CqgNTJWOfhi/8meFccZ9qPwxu8PNfl59TEQWNK+sZwnb
BVdxjJRE3VFt7cjQx3KioBE2z3VUlm1wP3347OwpH6PnhD8rBb7wh6KYa/Hmxn7SwM+E4kw9aDMc
VW3pEhTLFgnZms0JVZyAQsUuvUT+w5k9IKOZ1UhnOhlcmV6uzdUMWzsXbIq2WNEJjJbzgQYxYAQk
VRJbtI9IJY8+uFxqywNy3R7E7TtvwXYxFstpuPTbLwVaY1K1/uHW38eCdDRPBk51ZpjyFBBltb9Q
EbnKbCsBoozJtzM1cvWlQMgfQAxmQLXdfYiMHvz0HWSeVCoSqI9Vz8EwIsPuH+PNPYfgjGXgfI1S
xuve8q7AIfst2oUHU2H2xHoNBylJ184niXqjLHPRCwndG0FCbRTbxZ9sWhdXdYS/5HfiIMdkmlk4
Y5Fr028MBuCW8m+19FT+/EmvTjj93Gi+AhQH11H4XBvbYiGk7idbeUFBjpKm5vUO6V4qOGlIeCGZ
K3c9ZDua7LzsFQQqk4D1ybKKXgF9tyi7hgJeP91KE6xywkO6I46uoy2f1aEbWAWJSn4dLhYLD+p8
K3i+V37YQwTTQdK9zqvvZ3128FuZWNqd8Fib3ei6g1IO8osVvRbFrxEo9UpfnfXRMsqc1l6Hg8CA
N0gbkUkEOn4KB2Ewu4x34p4SQ4fsmnW3tzTCp/lV4WnlCGROLycXlnSACtkezB6A46HkxSWpMZeP
xGuBouJJzG3IYg9+N3aDr34HfyqIMjIYP7v6MRYc0dwPegesTSIsMVhoD4QFsIfoY2P07McEDChS
8KA84AJ36lvE4M8gL1OybcWQlLpSJOVbM0GmkM1hMEAXt+4W3LFx1yjXnE+7+Jes+K1vAb03r8wm
rPpBldJt2HeCNPgHRpDjFWOnQWkogYPWbu403jfcUv9tHmU8yIrzjvOsiRQZTnnsjz/OZyWrC2EW
2HYj71wRSaJ3UUIZ06CE7N2ZqujGcpjqCxjP6PwZ0vnsQy3x0SM5IpUBeCn8Iv+yJD/DCMPEwCHs
MXJZA/nsCq+0BwY2Sd7x89Fvh1BkDsuMExU3MOnHJRVZ5LUzc6QfNbOl6H56I2TaqW7cKC2Uy4cX
es/XeD814Sl4EnCQRV42mMRilr9YLT5gGvOyID/ddB7mAA3cS41mRvCOylz34qS1NeITl8VRQTGB
rSf1inn4RYqfxWGpWK1RGZOdSiss+7MkERX0KkahrKrJAkkv7+0fz22jPUa54/BDM8nFALG1+Bc6
PzvFQvZ9mcJXghMy7dME+VUoCdowJKKJ+XQH4jDvCePaekEhLcTXA7LU6S8CyBP/lchm0k4SuC97
d0d1jh/nVLSwq0pS80bc9f0zmoM/FtxtlkFObyWRLjdG35jGvdLnFDllDOSuvyCIqQY1yb0o0Cr7
9uHJCXXjHO+8MdY2BFZFPYN+xESZG4FSXWqiQzMHTgjwI93hougTlrfbnjFUPISCYqqDBRdJqgfj
0O6e8y5/lfDOAIkDIjWRFxYGHahdHDMil7VAp6rfaeCrraopyyjCBD1/r39OjlfE3dILWau4MGfE
wi4qUZek9yIHKFo6xuvYb/yEgqa9dMUcpggazTpW13o3hrFSXWdNnoIvOwRp43DrWpjOTbEIgged
ziDiWktbIJ9n7izDJXy5UqoA0pmklu2I+pqA0XU3fmNzXdQ5VJInteadrQBI/4yVwdzRoyUQhFu5
oML3ey2UKyHCBZHZnQ211MOZ8qFbFCZRZEidjePY9YsITGLP27njo19GMra6bQem0hG22mwqVcHY
iUD7FyziKmL2sGLj2XvnYQ7FhnzOWbIARJnRn/fPiKJnxCIXQ3q/stFDZ6qr8kKV4urUbOR3LPbJ
LF6uNNIcioYfqc41Ue2wDflYuIphYTkVZuKoxGPlYFOXRvg22xMEetCEEuOcA05WNRHx43Suiawn
EHBSd9VICOW9r/3tSZk1YcwMuM1qGPvz2EQghKW8PCR+NjAjRydsLUQlR37aOnW4vxzhU+UaW8z1
U3ei9tyhJU76GzLung1W5pD+2A3R6GD67Alr4iuuQJxSbJaNqLu5Ibn10q49mh3pw9Yyz62C01hl
wWPf2z3JQrffhSjzwkBW7GAC7q7b/xv3l3wVAXro2M+mVrngDt8tqcybMTI8hxIBo5V6/sLZYw1P
jklqhYvS4BVp2+qDObkZ0E+olc2boUmy1r9qMg64O6CUHPbp0AfAmdpImFC58KWLIB1PjoXwwSGi
9OAYYPKW1WFYCxPH+KhwGxJj0HSq/IASU8qEx0EdUAThII4Jesqbsjrlyoi5/lWkIUqXVUlw0Zmf
RB3H3LMpdYmLQheGoUsXEMpAtIULqsyqkFT3ap1lyAltDnDxskes6Olp7T5Nd4MIeDDGq0ubZ1dW
UcFUYHeavT6lrSqc7kDTIHwEyAwQM93+Ga9uQlrtc/3vHQb3JBK1VNV6oDS5FeZR6Xu91vOs3CzU
fBGZrPUE0D2rwR4n3saFZQEw0WzntlJ4/fHFj19FizOxG6EmoP1fcII8yONQ8JHGAT6M2qXtHxlk
B/ZfxIHWiogN7Bri+up5aglkiZQxQkrqi5a+5ZbIG9WMtTbtIdGCh73v/i8Qv/XWiBrDyKKtJM0Q
+Aa+qUSwxcPgjAF5Vmg9cmrx3hL4FZu6mgQ5eKCj42W2Xaz3OU4RdrwZgDxATiT8UJo611/O+rCQ
n5OeCmAwJ7dh9AQL25c83U3mG77yu77feAmkI7x+ZakWsw2m7AzhV+Dk5BB/b3F/vclIKwTXvFHA
hC8f61cYLdAPDfO1raAkI+4uxHVBncrMTYaaPzCL3ca65AxyRmn4Eg7kVn7ESD72ldbOqTUZqFzx
3jJ0ktinfMg3poStSNiEHgEQG/nDHQpK7oK+JIwH9Z72/IHfBmhrU9lj110cbBnrIkmc73Hiz+mq
EeShQ81R7FkGpO2b0wyNkHcph/f5Ib9/YD+7lrDuezspae+LuKTKaNNH8HQyq0HLiR3LxviLtC6s
JbtFyuXFM5qwL/hEE7cEuKk1bxKfmCck178xQ8xuu0Y+MtS1dPo5gIwV3Yu/KnGihxB8DOpvrNgI
QkWlx2+9KkUxdsPkkAaPxhZcgfIcvx8xOAIoHUytvLEiGeCpmmvP0NmdD7nb1sY0wO+veqtQX78I
LvbnveVREcEWGmFrF8N6ok5TZyXZl7AmlJOQrv599bjKAeB3ono1MhFCDxIwUeYznCAnmk658Two
pejfkJiCFm9YYYPBJn5JP8swGYpgooTMWZ8BBMZSIn631jNDl6Z+kHKS6KYRIZc4Ur04P0t6JCNN
ADtlG7rqqR2qS1cDJxunWyZjb2Isjhsvgqp6+Euqx8I+zDoo/3iW9cSW5ZG9m7R6nnAxom51lET9
V7PzBHujERzd/7G5W+h4gEhxfDhLZae6ULuCBS/TjZ205zenRAmTAFDWqv2hEkAnZgg9GFiasPcl
rQiIvkZ9RUavn8dNjYsECtOCaRGgRIpHR2LQEPsF9GD96drVUNbblvCiRqLFVMvAxB6HtMptvT1a
9AyCu15qvHwIeGgbciMl9JrvL3iC5TfIQrmZhuUYLeH6tNbwFFmF/TOkLyJ74xX9SUj/bLEuNXfX
gKXG9+yk098V9Vp11MknO446Pm3n5mKbxr60Xos5m4XjOEqVY2uZ0RsM8YF/XkPEE0iX2Up3ekZN
jz4Dr6r04fgYLASH20C3iT1OnY/RtVYikzEbfjF9QNdjnu05wkRwxWBmPmwfpeGbAfVVYutw+5Ol
+QrteA/zJJHRfZLfUFeoBVaZAMzvkH4Sopk5lFm1/jmTweQH+xELuBXbGUIcVyRr/ZPaFXSUQmMZ
nsuq1op8CWcNKBFclsZai3Jya36yHCOUdlLJUvE6NOdQidziaqdhGxgzNxMAduEfR78ujeMDCFKJ
/YHSmqTLZKVIYs/oDSaJAyKCkY/FW7FYg7G2cs4y1xWN4vbj54JVSw8shnAGehVYuoe3bWXArtMZ
2LLxKJ46Ob3lEJpy5iN0r/vsAMUnS+9K9B0KS6rmAGmpPjUfcOlRKO+B4K8sCNgy7Qm1Zg5RBW+g
fC3veX4ju/BC07A9yi5MRoLAZwQE5GFxAYRNLzBRRIjfMpY/v/OHEcXasgB1SQHPD3DLLykRxspy
Vl86F3Iq6e2B/Ou9WwiM+RQkMjYpOHbAJuuafWvpOMRd85JYDxuoxF0mu2xAXxL1xY+BpXfgzh5e
D7DW6RaKBs2F/5abwS1klWowkj5Z+gDTFmIQ4kk5FoanpN2A+QOkad8+wGVGH6SUT9NOllohoUej
qWyyJde4Mq1ywwxx/Ak5FjvULunELMR5v7ZKbgFtXQ8D0QhAZAdIhPppiiZR5t9KuT+Y33x2WtnO
t8LO5lAGlfzfE2HWV4odhb6Ac4RxvHasS6n0lvtStRPc7WsEQRGLsaBybXNZN9iPHcXBa1YQuI68
/0V6ipGMIqR6ozBSj0lBQ/YwhJcEYpGuJimt/kuUjj8Y4iMoLBhPSDuaOfcFZolNWmuTybETKOjE
HMwldICpbfyTXCkdhjcsNkM1kycC7rFj+8i3YFDdZRZbQqJeNW3+jhLDKPchOnDLS+dzViZQLi/a
JgSV253OSTS4L2nxPAc3rcSfs270OJfQlqaylo2jh1r/3/ijV1DxcWvuPFalwUipOBU70q4VIDCR
6Cv+bKZmHLQhZ0cDZVZUBggVcid8u+lzhFEpx9/deD8V34woOXFp8fCVP+pgqtgyGDNmPUWKp9l7
NKC3/RFEZizPSZGZTTbWlISYndkRcfQNQ9SbO2vloSJRP3zWzzIQw0+q0njj7NgLXZlWbbjjD9ZK
04C6YrpZ9Z+C2oP28PuryJ9AfQSns0U4S/YX0JyI6URusA1viEvnly368B7uSDkhascnABKssTfJ
WDE+vzP2tkTaE4tIoTRDjVU/UJbZfzX23zBZyhuEaCSulBcsMSkRj1mxGGOxbeg/ke78i+5Tb1mr
/7u4TTAwnXAc4XZoARqH/Xfrinl3LAEOisvEC7P874/R3+vzY5/6ybjt/ROP+0s0xZ/hoIjofiCU
3T4xapLG1Y8ZMM23RzJecCE/T9tNYMVaLaQ2lUY2CLeGeL85nOphTRTB7z4o8nshnQ8Y4FeGfr9h
pUSzw6TR4OfFUW+/PlN4yzbG4EEqsMDKO8czcH8Yc/awavxzICNilGIBB5TI081RTMhwCKMNgvoH
LXLbPM4uaAneCkR2oGy7kGM9smh6YE+kroayC/UkpBFzpHmxfHam5Ss5MJ2hknjfilZpDlAisBzH
+u2dBbyUZ6Gj1NwOE041F1e9oZbyDWKJZr1IUMTYn8t1xpbowZHHocYb27kASWTe5yNsNMkW5nG7
bh+x8qw5uD9icYAB82ldrknod/yT385fQCOGzpFWZkH+zrVuUULTHOf6fg915tt+ckTijzt+v0hM
x+Rl4oD2khpl7iswWX+yejnyBegnMyOzs/EIWvvV5pZme9SeAuIpjlyaH9vcA7LH4FLoeaIQ8euX
P1YgwnxqI9WTbOW6wj9djy14RboiMNALTjbk9X+1pABcaCow3kIOwNhtiof89byVTPEaa2Drn5wV
DgHaXbbarpxpks5CDZTkfL9rm0+INaXKmRHOsXal5hcMvFnAIAU034YZDHkWL7Q4w3sygmsUMdwM
phk0waFhXOtXiGd8qEyGMaDsypNOJc+/gR+8TgtZRyBO1jPRjYdXOGDdwBJnqMX+mzg1vGGN+q2i
BgqP9t2OSfXG3oRV/AFx56J+4tnMTbTlMfjrlgv53yKLUl0Q3D0w1ZSdYuq4wmJQA89o6fD/k36i
HTzqu/eytNU2IOTAXSTttDXkhFNagFRVNTGYP7BBV8K6xVMf1UZIxaTqS1XoGlubzuWyXi3LFaCc
qrLIPtaxZ+q5LMc20pGCcxRH9avPzxJz629812TDqswApJxwQm4Zx3Ph5x7qnqqfsc8qNKQfLBRV
g6imjJUef8ltI7ikPqzs2yT+wNgjpvnTDULbJ4xXX8lWlkzUx2SyBcKWv0wHLOJdO/ZoYiHHLhkA
oOW2oR/jXq00uQyi6qk9sYWutMKnOrwdJeIQ6HvD4Nn7Vwr4DYxXT1nbVdz3LYGEw0E8Dd6cI8Xw
WljUlQ7mKKHaDqjf0DFdjhVpHTxiyxyE33nQXp8AA3QDnD4JyTo2gW7ZDyzSCvsQP/Bxvd/MU980
w1pBhgeHPoLOjQcIL4nkYQ0ewYP1vltYfG/VJOTxOiaOMF9nQYO3qpiFlUDLTkMHDDnRclb3uQt7
Ec5xeByAsRZnYzIvB5Pw3Bd2rApBPO2falYhJA3oZ2bEl5vjBl8Ts3bFf4n94Lv8Yosj1TundyPS
3hwez9Y35dbvV10lUW6MoWEIkKZymB1BDreMkJgtPvvGfxHAE4ZsOoqTG3hra5ZSSUqKLjo7P5q9
7pa2eWxS3QmVmkYiwLK3ORn9vb1axuYru0C70f1bwpetBDIl9ZMc4tEdfqq48c1tpc1OJYY/Wwyz
kAyPINFlP9n6mkEsTZKx6i2Yt9fkITZlvINvUQrdYLD3k7nn9ZQTTbBvQZ9frLZEOnfQcXXJUbb2
+6MHsjyzLOyNgqB9RJgn8r9eIxo49xdWAe4XVIR9TGba/hH1+36x3YkyU7tqoe8K9+IwgB2VazWW
ClhTRTIlVe2G6FxyKmCeS0XJ6OKCdZ+6MyrXKPkEmJECEFcyQesv4C1gWPpuiZ6B8gvozJ2eib3s
6qPxuz2K470enx7qAYamCDyKVhYcmuaygOtBf0mKofUWnvCoTL6g3KjgX1g7eNucFzaH9relInxq
+Cr415WYAwOHceLy/85zcrX7hLrH1A5ZTXd2CNPrGZWLtcFTwXLEFC7F6LWrEc1yd+k4b3vsRd4U
ZUonHtocgObrzytiVndwE4by+s44VqqdacVXojthID60QmCXtigeF4h49p3oDx7A41YoLuvHpKwh
a0kDcSMAdyxRuqHp03uq9aosGCQycnU6hgS+08L/5/5lMCtvdSv+WHjKxBFu1XIjNnT+fuKBE3Ir
QDMzyw1SqMw6ZrWdZSVbySUikzWOQqjjzXuTjIFkVqgNrlrowLwcwFiVLNStErMLT7mr5HkaPVKr
F0cpMNQpQAbJ1Mkc7u+ofehsWYSVtXExycHVWc5nJWbAy+t3kCmAVx5a6zGs1MFRvpX7A0vI4xy+
QTXQujjuIQcFGnaxjHB16JwklZxSM5Hw3clJ2epXJpqE5yX4Et/SJHEjvmZkANM0E7Qm3CHGdjtR
NLWPWCGLAXGbaCTDNJm7K9Q0ENZp1oNeDSLRhUTOE2z3RnhrKIpfC1em1QZodhkh9DwWt8S3iYxI
c0xGlo1A5NvupQ/3xDbckMdFmKkex/gr6drb0LJTf2lDIJeigiXdKDLrA7HeG1mfvqhArN6BvwNF
izYdNAzV2OqG/ulO9BIHReTgCpqK51/8XGbt0l5qBS06Qyi/OTzURGKINUgVUtUV+tAIGu4u3m47
ll6Vw2pGNXsEJnxN/Wimv40AbCz2wUWqqPVc1+U9lg+/NCqlpbDiKL3Yec/VqVQCwf/H61N86E0P
9E7nGtVs8prmXWsfy8FfmS2UnTuBjYJD/d08f0d+IT4qx9wBhCTNntZECK+qMZRecjrabtw49Q8p
Z8yRiBR2wgaBdcWz5RS3QBYzwqqLShnyqNCXZ6gg1xNf67AQphd+iuIDnotKZX8FSCaPfBciSm+p
FoqmdKRcwUJeTMuK9p8NHoLawKY8M2Zh5uSMCMGUMxj39Rva3IV+iqPDCdThSS1/vqnM63fbFYO4
PccWn8bq15bvAAwGC3M+c32aoQjT6CtFAO8/DRUwoPc4DXL9Gnh7GpNCjmIAIovQEsj6RMjJmIik
MihhTGrTOfzLRdJGouUePzRyoMGA4WMKGNgwA/jrDLwNxbHTo2vsxMb8idCzjxdB88erqmkGvIvD
uSmjbgs5WihDjxCUEY2RqRb66XuvV2f03+SKVP33sd3lKwrYmNPuB3QUPIwo83odoZTSrC/KFnik
/NXSy2CLvuWcnzAu8+iobP55Xtz6N9umYn5kqaXUHh2aBcN+nPU38d1fy1fmFZqUY6faQkRmZ5tu
01IczineejM+4FGyff2N/uGipPztbbN0ZTjCEzzkY5Wg2/JorlxmXjZxdjsna+zG5NYOmWBkMu1b
uOhkhONelO241WYaVJv0xISAa83PFNzc6nakInNgK/21NFCylGOG5GDF58OBAe/lcgFW8A0Kc5Ll
RlIZHWzgmX/aa13jKDlUGhLBkPHwjixeuFbv9PCCV9S7SM4d0uxcczoiO7ZFPvby3/fND0pIOrjo
9PQ/4LeibnS97IDwTO5+K0ken6TOD3AVlrCcfgo31pV2WBxbRquKkYAzsIsQ5ysIZpDpKXSuYOoe
koH/dKCLWY1vVm984awXTYugBCqqY5SgKlRs9ETxedPVAIrtbhrgdNoeoEkuoJyvuZVHTLa7iykZ
ksL1XMq4O7uQrv8Vk9Rqr0Hz6COyCsqW4wiAplxsAn2ny5SUACBsVKpYqkfIV5qG32h8n0E9+kRP
mdNgxFXQGYHcnEEotP1UvUcEcS6uptvX9hPtVIU7Cjmqn7qAYmuxgV8vSUI3du2ebp6xISCWiiYv
v5XmqrlwpCjuwW9Ec90ogEEwrmtS5PNV66s1ysZUuYwhG5ySsxPaABL4Gtir57vhw5Q7GVFLWAZl
yTX7AtDj/InPUhid1+PX4LYFHuckS4wifiK2WhnTCyLc/t56WGnhYf0b4T1mLcPV+EaZoL8rcHpi
DxBL+YdmkGRRkxnLSG6rgO9kAG56a4lMnjR+F2AcG7EHmLGh9BYRQeu1PjfMRhvYEZpdUlzy8oJR
L77tEHOyUlhDbv4Opb+hC+KuqCo4FIQEQpx8ky7+OPELXvbbrK5eWj0jR8Iud/l76Fx3iI4RHz3C
ieptfJe5yf+6KnyjBDhg26KLl9HWHJmioQFgEC3Lf1NXGAD9zzgGkJ4K7JiUZFq48pymRVN98jMA
o558LDDMGS7XIBFYP57BiFww/R1vXULYcEXVY0ty11GLWpvDlKz7pBjISzBBj1ulDtX6OXIGBOsQ
Q5Twel7QzaB/MXBDBQsHNLXnmtYzpdumuU+M4SbkW8/vhegPynGyWI+U76layz+4pkO1aew/uHEA
QQOnqKrVrYCWTqhlL/4TxWWVBSx/bZFpuwayLdBQKWUpFTF37TIJWhGGV2T5gy4eth5PzuM62S/j
agm1RjJWOvN9RW5bQFto/MnBUc1TNzoBYLw76RKntwvQLmzIghcRHbrh+OFJBwIrGeHoVs63B1k8
kc4Iu+q0YerXEFl2WizAFrPX10QM8Hpx0Y4it9fQDjZUY6Iqla6jfHGiLlLZD9Yvlg2QhPXFZY3R
uKLK7oddvHsmJK2WOojxv9y6Yph2DR5dZMkLMDlSFA2QdpOx2HyaVRiKC/u0caijqLwT/qmXYvA9
Zqpv1vKks6nIcuraGsFABn9FxVBIcC4EM1qVMbU0k2GrSHfrgsQedTA59266qLwwZJSTPyhtaDqv
LhAimBSTu3pZd7ggU2l8tdIRe8w6wR0jwqg0clQv2s4O51MB1hqI6iuYneuKnCIfAaqgtWzjgDr7
ProOT6+nXz+AF5eUv33NtZ8dZkPuCc2fU1gLHWqL/aQnpt9ttjqnoDuuAmMJqqbDxT5MQMPF0Eyp
601X6wewd7byb1puGGl/IYvs22vHwyRtZZAsAJBvtkKK2NO2vRQX9+MCednGVHAJRVTMt1ebj9Dp
KfOSQd5az55+gQS12dnCyE5YzSRTkm/PBSjoz/jJHOsKHRasDnKkJr9lLgvqjAKj+DE8UwIRowLh
J5/aKZBorLcc5hw4fBxhHaKVA/aQyft+EsbmICLC/yXfKnVU3n136jN3VILq2GKQBTX9t908/2B8
HfcL/JOVlSrztVsoAY4b5ZKJdh/kWqnBuG7r2z+Jp0I1JBI4E2N2NREg5IXs21VtNAOrQJi6RrI0
VT/9iV425MmpdLWhh1ykeJGzrcNjo8Ni/J+gzVBZCM7LaFg1dIF6h4FgqrhaF6s8MymLyze8VWME
wtd3pou/8ZiPZTNBjxzUtnj9GDz06GrnUkl7y4NYqR0rUBGm6xAJmeaW6hpLI7WnVfTSk9aqEGHN
eIn04iqzfL29qwur1xjwPHNGjx0hjSpfS7Q9plnH4Yzm4SXhe9fw4pJkxquyUcJnf8GBlrFjXFRi
JdFOwbUdatvojgdhfQNFXY1XYCvChG7kKlOYN+rKYxA165PZccKAc7YjAFk6gxyZgFuo080XghPu
cg77/YR1YXGIzB9UuwmDeyF2Bz+eBh1R49M8v14EurgJmDYo01rWyXwrtf0LzqkJBuaueRCqZh04
edo74J/T8yneFvRPaeAREu2PQvcCo8wIsqZYFpnLN7TRn1Ng9SW/wc0ng1MUvITK8ya5VhOSG53i
7iGrldaP6qZKvuDEJywz/m/slwlvA2MyDhsRd/xN4iKbtASE+6GlFVTIgQzXfGZH6hxYIb8urQIc
gZN51ROUfZ7Yich76Jp+db/00ZwyveJiDIvb4e/ZXpE5oSTf4FTikfSk4RJeKxkxjwiN649YJbJc
hI+MFf1oEsv+hbE8qSkynkrk/Z9umIupdjNO+dQEl7x6bfyeF1SAALOybG2TpZCXk/H5S3UFlgg/
0IpLXnKuvpf4zV+BbALfuB/pEUwvxOd3sq5IJTQLveUbGhfCwd2g1Rv5gqGok0ZGFi24m6QPUZaM
TsNh+TKzCOBgnlWPW3CGZUBLEyjNZWmVR0SX7KvN3LpfEF6ZCByqyHKPBW2uHzZKSD4TNEacBfHt
UQ8h96DId6XjqLpsOP2Ludy8aGsWzlCteTrYHvKZm4HiyXmzFWCEIwzfvJyKbmCrkNz4AIfBAl/9
vxvCelW7cQX5AvKG2uqDgpt17sW93SY3qCY46tvVwUS7XeKyf1IHGNgkpr1LZQ83vPoA8G1fLSkR
+6nssNHQZHR0EQnvZIqqHXtCnr6DjDZlZH9mZDNYln9jONZo/JqM+8h6onji/bQ1Xa/dFAa4XZ7O
5NjUamuxvcUQAGc6Ce+pkQl9o0e6KWnhpP8+85oYSeUvCmyaXzHQ2y3WfAraNbDC3R5WrKHmSvSu
yms0GGa1pGky/hWqbhJwophuA9JCAbPdxUJlDAG83352qZTsCSxnFrAlGole+Ts9lI+k+OTp6C6H
FxlG512qc0m1r71Zd41T9FToO7HDJVZBAFhTFL6KRktuhIii/tOmhg9EB3AZe0tZNB5xNGZgsiAu
G9+mF2k1c7HPIyiOuaLnHMoRzggEamuXcDsbf5jxH3B6+0KYDK69EojnbeFreDKB+YdPvEAhq9DN
nn6p62ySZbiTsNkxWSr3/sYhZoznh8b+JCDOtUD0VD2zNPec81VHJ81AFa2FNXlaj5/ZchIK3dWD
cffAcwGsCnY1cYJhtGH5VP94U/77Zj9RR0UW4RQoj5gqJNad1ptjXC6Szz7jR2wL/p6Br7xI9zdP
fjIc511cfmFOtKYmRedS9xlTeAImrfjvBI2iH61NWjtp2XcLjFEcHLeBW1gbBxji4gAAFBLYarb2
z5zgCek99wOR+BfWMkW5NmHLhAtIuxCVmfNLStL9aBYDGGMHKegxdBcrrqgJrXNy6cCrXuaM5ztH
5Br0gpih6wjes24d7/RlargJwAHpiNjFFkeXiSOzCcBuwDXPQH3kbRXgdIdp5WyplmWuTJMYPyqj
lJU4Ql8OoVnS9JEYRdVX4sGHqdrOYrgBxXwYeTd3e8MSlpuU6gOeF9rkMvMmtlNDhJ4gN3z6hHdW
4yQTnqL9RHL33t5SHx0iocfrBpizBF7853jJ1Z+slk5Ci4+BdR4sHLo2IyHh6EL2KiLLmkgS2ezA
o6NxAW3AzR2mMMLU0Ey37n6vzLn9D4suEMZUpg5jgKEE9416y5U+CmTHsYKTpPgTLTIX/gENjEVv
sFpASuCE/3/IZZ16nVeJ1VJtNkZuB3fIh+p795S0I/eQfEA7NtWHJjWasQcD1LxkLKQgOzcLXXJw
gzQGkchhs2LGYQiLAxmWpMNi6cJrmgzFKIIiS72RQO1TH2/J2hyzqsCZjX+ZF4KBkeEw68jWMJMg
02s4R9rdaqONrL5mxiGWDs0ImTMOm+88ms2Y+y3EErNklPSMPdpgudFGc0erN6okdlPappNufTw+
Y0c5IIREhjzL2Uxg0PCGF3GCaDq/DbyL6J2slhuxiMm0WUtg/h4D/clGLkLVrM+aN9X2rj4IigDC
LF7vbZqOXNAOx9RwqzxsftWcanehBul0ECKtmlrVAlUVf/IrCJ4jNz/q7s1eUYKZ+dqL7kXLiKJB
gYsgMVA2JXnItWUBkF1+phSnk9PiwyWkrPk8H97br80xs97GT9P7PxZMc7+xl/E1YOPAj6B5u7CQ
Sm9puq0QTUhvrTWE9RAJsAKVC74nTXyNnCPeT1eUGYz7y3K9vOkM6fvRMeTRkh6HcXTVVsBr9vR6
B+yj/6Ug52AtrIA5S37fmN4gnOlYnghCnLwgqaEESNsuGoKzVcu2oy56OXS3JlhwVBHpmqOsMD+N
7Zy0HzAHPGgQboS7uoGe+CBh3z4yMgGKKaPfcNhmeu4lG4EHNrBpkEAA9YLON4WrqA18XdC/oTtS
XU+/cYkmKbF9qMI+ugnU9eSKnexH95k2w6eJv673Kv2cD0/Rt16b+9Tsugrs7I8JO9QmrLgeAUkd
wzezCz02S5XRk5iU7wWmlLbckm7fX3FH+nT83kRh2hnq7ybHSt2kW5GBvy0ZSVzVL2nsb1FBt4Sq
z5TResPY2ol/JdCh7olDk/7mXDEjdnQqLfr5XME4yiirs7Fq0bvBXweP6I2BRsc4xL2tEJsbJRlJ
TTydullDzqR/ZuUA43Y26dkGBou6R0dC5K99F/j76l31Dc+oJ2PXgnDTwDYwwJf6xALeb3X2zfs1
5B/+xxbsKuYIFmdqNmIXtGVFj04tmBi924+2p/pM616AWEwchLOVePGK50xQE7a2+3vF1iD7mjwm
wUGHI5p3/D4QjFgIWEtZtc0Nbpwc18+vmRltpLUIKTZIbB9HGe62TBzL+auB1HQjLEVBoAwJ9J1I
jCe4vAgnynKD9CmKMSzv37Fn4cipPsAxJPfCmQNW5a4ISEcX6igVSa0/CEHF9QnbOMwNVL0j9HzC
zz4CiPztcNPrDPeskg3Z9CBMEQQgGz211RoeBZhAP50Mv7yntUvvXX2YMjXXF4D0ZoLllDHBUMS7
F08ebnWsz0beVLJ6d+Q8JTFVEuVOanNb9H30t4ZsYt5sWnkXNk8gl3sKVxtGDuohwU7s8waDpfgD
9/rGmfZLEvELj1LZgilPfc/C6i9uXejBYuCpY2tryTuCKSmykpDjXH/f2i1uI/RwJlwQ44SSyjo0
t+fpDjbSPO1biYByumbd7nWLZWHj3b43RpjHfeB0c6Yzg6l4uU8ZU5HRzs+s6iYlksrNJghCxFfB
ohWCPXMlB9mnHEfVTrHSPyavwmVuH/RQii8QBz5K2MbDGBKQD24m4+zDZhBOjWM5FQl4QzslvTFx
M4p0xStNvIs+DovSwr7Wvlq/k+EKlj1ipJKI7I8B1wXq+Tz4fviQAb+bUDHR27WY7nyp7MhXSy8M
7lsqwipDuu5NRDO/Tq/tHMLlo+RRvyGx4R5U/+3UfzJKqhVr/lE+IdqRQK2ZR0I8nUk3TKei6iDG
tVaVtbNk2cDSYBJ31EEcKEY8SJU70kH5cN/0bOAVEQXTDPR/Lo+QxYjsGnuYg5NMxrMvL8X4Aozz
Yxd19Oewlfz2451H0rtuMDbOzOWEXAYkxhIwlP4AXuHPxakdTr1AppE3KexyWp5G9MUE23A59ToT
UzKBg1uo9LXsXCoH4Qr05SiYxfDKeoPrAFedlSPaMDvxIqO8AkZM3q7GLSPx+wvgyi9atSMLqbkr
4OF63scIhFlrbBGgUHJx6npeAN7cnvq6SAWPVIQEMgUgvJiryQwXM2kx5lQVaB/V9iu9OMK3yQky
pKgoEpOxrQ94R1lGvPAfH4JDWx3uLgayU8HdcGFvj/By8x+yg4w3zB/4uFC8xVGuCw88Ay5cKKgq
eEqe8cbkmUNUK18+EZqTlugUiAHosR3wupjianwW0LHhRgII2y/LvnJulfIb0hrMVdBAm5a+ldvr
bkkY7d/nYD7rFLRPh10Dn4EsXO88w1UxH+A5RdoBg3uIuGLnYExaCOvtK6Xa53PNyhkubePe1JLc
HBNr87GytMQovHdVh+BHeN3o0qThTniOwrQJYBmNCxbwHUkV+/w3WcWS281Diqz76Fn7bOx5f3Wt
daxvLT+wtGNxgegt4YVUpz+qiiLdWd1iRmf5u3y8DcgIjdPttmsSidoB4oqrsv4N1DlVCz5sggo3
Fgd3V2l6sr4PWam8T0oPk4d0WYlFlWCQwv2fQPbMs8tbJLvyYUY85/Vr2C/KdywYXDH+nzafy1R6
zgWEvNU2DzN+udWrKlMfMl+rsp5L26DHmcFt4TUPPwVj8eq7tZQoCOt0O1QsMN4c9YorNcIwpbX0
gqKQW4k1VxporBUmuIBYlPV0Nr84rgw+AIUlZTWnCJX5xNSeqviJHo6AyM0Aqzrm5r9MxvEsaaj+
hwooOH/HOLLQYrqX7xGP9SIPugA+TTAtu0fWcbCJ9IMK7p2wRFS+1qg8v3gl1Kh9agPh/Cq4sBoG
7DrXWQjN3HNk0KV0EFIDFGVwIg3d2lHupt+FhS7j/UMo8lqI51PO2LhBthCe0w6MQpqfCLngKdqJ
zlIIO+h+hzz+YHjjSkL03mwI4p5i//Ud85EexG1b/lNdZxk0xogXIcpZJ3XmXs4k9t2FTx6mWcee
M//6nPakuZ2nYovbsOeYSG9fLI9oqCbhNGLf9lr8D4zEaelgM/pB7Ww3mkcs+sGFSkkY20MXZy03
fRZWvv6lS4Fyn/x+Y3et1NrTcATMqcwaHWjelqqI5/fGBSHhV6b8fDSBuq513/+/JCBDmjW6lQO3
PcZuBt7IOSd8Goe00oLKt0SRguXfpWzrTtlwXgl2lyPK6JexdXyUVWxUxhOkJk99lHJTtkZ4JUT4
hOl3nOcJAKWCV4/7cALoZ+ZkDfr/KAQTrDynFopOwCUf/IT/DR7JFD5NlBaloNBk2sq48R6O6TPN
rsJ+G31TcdXaZb9y1pYpIWGs7iTAxrxqdUuQ/SXKpTugyQ0+/ki1oWnwiy/R8V5zFe/ScI82rlTq
+QxB8GibDmEU5q4zS/RziIkJNznpE1WDmLt73cCBjnxlHo2OX+HpKXPw3U/w+4DG3D+w4Qid+E35
bwQE3qgQEut0iU03otQxiRzC+x++9TxGCvYVPtx03P63AsdDnzJb681kpD8+/AE58BEWKeMKab+v
NflJxQx8iZfCLVQpZAIaK+vG5wtBYk1wzNjA0HZvQaKfgZlrZO1wbO9g7AEAjFIbBtEGuE2yX6ut
nXinRFHxOHGcoiyb5DBkwAY9qAijaCGO77eppPPNhjIxq8Wl2hqzGdUYe4VBI6A6n1sLNlGIaRYR
wjrPNTqfHkNzxR6qztxiEXGJpoMSBgeKUUhXengAMlpfTh5WyOPM+W20k8lx2W2wjKUwrKlCwWDM
mbycQab1UWlh7mW/6wwudZMgNrpM0C8Of6LSe620fldm31LdTU79USJz84DjcofRbUrnaRoinxq5
lnzVCgAFqLi0m34iwWeMEuq8dBSE4mgp+5jwdo2BRdVPfjPHWi+rRLiN7Sx14i6RKmK6ElwZTEB+
ECiYhQrPerabnGw6Uys5gvzXs03DznH4elLmpyirRqC9JfTTUtT5H0cXcZPFNzkJN/9S4MFP3MFN
sWGCWpPhZhQdMy5cTRq+T7llyhJC9Kdh2jWgwFa2yJ3plE2INh57EHCH9tcsyYD2RXZl+svEm/Xb
zZqjOxCAfLPfUDDivRaSJmmqR4oPdWO0Sl5EN7aQlTI7Z2P8L4RsxMge/22DOC3ZgOqfrfRTJuAf
iLpv/17Zvl2zpeCo6idfx+shJEQdmCp9LVxwR+Ojd+kuOCPYoHT1yJF9gVB4u72tCa8sOnYW60Sn
1l4xbl6FGFCzRFWmEiFwRDRoJ3Ak1l6YFXuHV828UcLHuQhgSCnuEZDfHbEe6+n9StHyqeL7dQcc
h3AumoyW67uFPNLpnavtU0lYg1ETYgbGICGs3wV4+iTrl2ZGTvU2eMzjyGNAlF0BrzZ8teOYp3D5
a+bga42JCCw3Wb1aFg3X8beAlS6k0eZsTlnIYEkFCtrflKH7G+yJ9Uh9oPT4G1ti5SzCCO5BAjEw
qd0o5usS2IM77Dw/qPcwSAIbLBqlwk9XJhjsp79tu9mC/TVqR34bCb4/34myKQ822fvfsr/zF34R
GjMoPwMdpOPhz6fzpK0SldEBgAtqufnGtckLwAKh9s1Kams3pgNSLMM0uaCeGeAKFMJ2//OCCluZ
si60eTeyJQwIYoIXlit7LL7Yew0w3VbUTVRERJ9HlBIxzRzzD7Qxs5L/Rj3ug+9qS0lXzpsbEFAT
4umZcZm1XjUKhkfl/s55ffvaEogsXOBHJoVc0B9q15eb940J7iX5mxEl4FRmLDcsw2gv3PoD2U/p
GwqYwGFbW/ze1/kW1n2sqK3wQd+WdmJDbBIJUI+ezWxFcvLiZN/c40Bs8VwrTa8JkoIfsmwEglON
F5+ozzdACUv3scpPFlKRSpz0WaIqSQG5KkjQfv9wJCP2PUBuo0V4+TP2tS563FaGVh5I0Un0ELG2
HcmKhRK2by2ITDu1LwjpYaAUJL+e3jGcwH1iHakR5MkjE2f5JBNaUff5Yw2MynVlYuRg0rULQTdO
JhpgEgy8zgPpMnqZ05glEsjAkGNec1W5g000XvZdMaPcIg2cyNl1wcNTNZTDHMj/QPDP2Tc9Ozh+
yWG6X7opsSEucW0rZJqSVoNe5lUtOBfYPBzFYujCgrhc1/odKN9N/tSLAsDBjyRj1NTbCoX9i63d
WVXTHXQcXj+2ZuqauLN+gigZ7dxdZE5CDm89XFRgTwejsidBdLPahUQawIjiXwru0knyaYnwUA4H
iul/TPXouxpqp4rtmS1w4pAqQi0ZTZwb8ZXLWdV6sE/GuWlxmFAwm6NpuAwtksirA5tAgN6hY6id
WEKduwmgbixyPdOCgXXrkrHRH1ouDLelOeJxieusRAU+dVc9gmeMWkarWSXYYZKtMBD5mau7iS8l
hWWeKYMZuhAe7hKGpikn1YMj/uDth1pmpII5XP3TmdZiNFVWN2qKhUVqim8/m4mNmlLXLMZwRkZ+
9gZRmn4GxvAHwuwib9ZwuntXjPT2HOmIuKkgK7BT52d/Jk0Ijy421fwNpcVHKlv4v7FOJKEgTHeC
dZUwKBBngMuPbmkHp59SEhBL3alWCNqHzGgaU6kOlU9NKbZhl4H7EfXugsvkkvdd9JFyIir1G9y0
YBV3Q5pvyJHm0vgQhC6El1rkOJ4lejDGwmMmoyt9DFDNe4pokcVcyygvIyLYAtNR8EKQgB/j5YTg
90k8+HYs375D4YITDvprIn3Ld683RNPZi1dnHBLBwZMUcYUkTTbz7qdAyApJZTuU3KZqlkEjMp06
MHK+waDJihlxXOvlFOTPaDvCWTD8A1Q4ovgBj8Bqq0togG/4z5U2aNytqnk19M/wPEq0DX7I4Vup
3Cp3jwEkoZKWol9/yoSv+QPci8ic7C8t/2pLLZ579Gy2SdWcJYj2jABtHYZhpphAAAOyxzVsXeHv
NDCscnA/3xn38iwhrUFKrpflGOPPHYO3fHETkxXS1gDONew5HrBlTgZ2eragPilP/nxDrKIY/M0+
0Jve/YE0DfIdzFwq/t92W8tMc8h/2DH128OaI10NFzwhjMsuPqcIpoYOOhO2pDvryvrx/CNW7Nfa
SC4r0toGfQ9GSGMvG4fJRecsqLs5yFWVrcR43KCWj4enrOZE9TM1TNy6ZjH9XSNfl4BbN/35z8PV
GT5A+cphAMs08Y04sWogH9+XkFAVp6JXMbto/98cZzLPDX5jlNiDgy3cgdh+0iKIKbLSTV52SQCB
ILNB8CtWS7smumQZWMEnb6y5Rvn9QVY7OZqjO+nRn8H52duCspMumws2lkc5K6XR7cPxL7oGhx6+
+gPICZk6HtK1mzFLw+23IIhdBDKsZkua/7FvA43RKsxB4Xzdui5N9u8Pvzk2Zx8n9v5An2+N/4JZ
7eY9M2EPM/DCbd/WmZ8sJ4ek2JeCE1xKex9UzA7MMzMOHI95oafrQ8OwM03k+5JaOBGMexqsm5S8
egEeZvFNDlBGh/jaoc/VHdeDYs0hytE5cK/4Eh9aZ2JdiZG72RvKWd0Hn8fbSEFntSX6xukvRFBL
7rvufH61TWp9ogiDO6M3/rJFdEahtchgF+MZ6QedPyf5R6nBiFjp9A1ji4SucazAToQ9uyezBcYf
v9LZm1S+Jdhkj+Znq27eHBQY/FMCkkmxRAxghzujOgyjSNRUh99/XWCREbg3rhoiyGio961nkKAj
9dVV3oD5p9wVZHxvxZzHDJDqprR/xtOEK7FafVkh3E4+iaZL33uc+2pgUaU4+ULLplAlColhm3s0
264XdAVecgNVR1PJOEgPGRSi6tBAcFoU8NkuXIQ0E+4Uvq0CYSDBzKsQnjl7CTa05ig6AIuyZ6bd
ma+mZzpeZai5tRE6r+Yh5v22gNUYfIKxe4Gv+hHqJCaT0obSACJARmxwy/QeA8n07HLkuzEfuSCF
TBvM5yYIQSthmzkEYdK1XdYH5OS0AxK9Y9po2TTqAtn4Zd4CDmEP5eYmiM6Y5O7jFbvQ5yE7RYM3
lxsJueAicD/D04oG3rEz9p5d/oWy/lW/ivUI13U6p6ws1hOJsbaRr2SfI4rgx3ZM9x/wnSL30iH+
c7Zksy+v9a/0jsyg490rUYZp8A3e+e6Pl20qksVkW6pTf4Tid5aWrSlLMcgfRdToZvJnb+CFWv0X
3wla10kglc94XtA55Q3NLkwAIaGQDMYSQOKV+fZEdfi0/uDA5huwv3LYCofzqMVI8ckrfZCe6BCl
yHKplyVD2xJix5pTG9cisRghpe9ZKZi5UAhAtPO/y51lEJy3CbZnR9qRQX7EXdAdPPbBaKrex1E5
7dJ2mBZJwiYdghwpFxlZoBXypIZ/1dfllI/PkFx08EV9S0CfM+Mp1VDwfuTIFLR6fYtyHLQM94c8
5rpSEyOHCgUBP6Om8TSEhcXT7mgsagMwIoekJT2a7SsIUt6eqFEPSGtAIgIk+hltXL5CorpKvUMg
KXAHzuMQ/4aisj9qvDRU1ilr0X9wp58t5syNGEOpEhJZuHXESWd6HjfcLZ+F+qRXwyoGXOmKfw0e
wTOfQ1Hf6uoq8hFbDVmXZxAWNyL1WTbNndB+N1NA+Ooq3xd4DdXkxyqIAO0otFoqA/jJFkBweJfj
7cjekwQjuJM2Xxoscnc7oL9iKZ0MDR6wq0FmDNoSft+ZiloMqhZibz9dnYZQlzUkcZ/EmvwaiFJw
7YkjUpkh0qBMgQ0GMN/E2liFFLAHu8569AWBiqhLL2bI0LnyFlA7GzYgyAETbi8SYchGNCJKvz+B
0vQ4DFSs54s1chpjtkoYk/aZ+SY8MeNrLRj6V3RVvHgPOVrSQ4nQi8ULRX19v2PBFh8I7HSv6DuI
nXVWhuVnqYm6yayKsBWEllt5jiElYyXZHm2uLFoZMZjJnhha0mRu3YAbalFhM/YGV6zdR91vQBxm
D2OkOEK9LwkUXSlUWcOXnx/GkBqWB2IfER1SIuo5hKYwrKpuHhHS7zO7fs8V9ho0zCAgks4N2RSz
F6PXHz8ruTKVv7qPuy8whUbTRYqqA5ZZTs4o2ZkEudGem2wvjtCvOdGIKWpLTHHU18OONrFaHk92
Qpi83UQVkf5NiuweYB0d56WFQeFtJQMpgsuLAib4waPxRCXMSD2mt3uVZK6mCEtrJCggSc8+GaPF
bZYosxLYV8hz7SjIyUyM35RtIc1PxI0Aat2xn+2AJJv0q6IdnbpPbbTBz9QeZnqNSdj2jRQj5brj
Qm/GcJpGTpkLsmzbQ29WjPcez7jn7+EP47RUJo103SsxDP4gRSLdIVgVluj/NyXyqJaTiFsrigVf
AWJMOM37ZZ07vXqqSzOZpUxm71uZaFe/9vz+APQWPZXr55/qj9EhGB39RXxk1/UpffXBFnyw48bh
7vkb1hui2crMUWDC5VrMFPyNrEpFUW7k7EjXe+9pfuDp2QMKGn2W399UHys7UibaZ9JqiroHgQ+K
wOdNXklxTaWj4qovyWV18F7hEhHjRcm/vlIyc5haO5o9QB5WPn5HlqK3f57F8BrgUnIG5QEogVh8
2BrYu1i9Va0HUzXCMz7stkg9Etou1aYKt5S5CSd1JOa7ZGvEJkmWcJWsHQjQrUN/jZiwu/8lf9bT
zYGYyxsL2GkAzptEQ+TsyMTthxfyWhd7LRSp6LeNXA3GFf84QtXFGhry3APP5Ee5IDWveaPAcMyM
EHBYgv43nzVEeqGpVuY8RyBxLtwnspDz/k6RFjr3udn5+btY9/RDFvsTiTi9fDa5izbFqM7Zbuw2
MYGWFm1aZ0nB1Dl/3AkW/tv7o6Py80uzKO5fikqaLHyHXv38av0WarMJOF+FmkOKc3yA5YxSElkx
0KDaUuphSYzFEB+Y1b/w61x+pQdbJaxvJ9cGmoG8rKCsYcACNYrdQz+mvDMF2frr3K2qWgt5D/QN
3Ts2mV3K0quKbLmDGue8v8/f29pb5fvGWl3lM8mru4FT7eA9SO2HVnCivtx0bsilzkqx/fnfXKv5
RJmOwAuC7nQwMa/M0Cv2pDdK0Xk166dhoIgvtArYBIlfiWxBem5az3nmk1XT5e/dd6QQbpY72qMk
EKhNtJ6OpNwW1vAFIQKWAXjC3bP0FSzh5CKW/qH2MlsTH4OYD6Zhca2qBZkxM0BZEdGBEID0c2wK
RRJC3PNk927DKzhg9X0657MJAjTsC/jTsu5G0w/JpfmwSTqr4L7b7rP7PFwO/BqKeyAnhURciIsU
R5+vjtRDtAfTPvTM1q6wh/EncN9jGJTsYPTN883XklCzbZRQKWEnzfb/0doO7Zb8Ey04p0ChVMXQ
PHA6mJkMMBfvsdUQeTxWHfz1sNj84pbLDGxrd6Zu7eryvI9DI8vMyaO1wi65eqeguXQhEJ2Y85fv
SvL64WO3RmcXhC60ELKpYESGgEmROMANayYsnQov2N934KxU08l7OIm3m1AyaeXNwATYT9ivGb4Q
faqMdvxbJ57KdUAv2vIkIdA6s+3ur8wBFyXA8+S1s0F+yihNpMC8n3iKEbk5K+VwQzjY5ZFEsMj5
qzBJ2EDo+3qVIccMM/coHmddPss7QJP0yVWhkt5FAK6qPCYsaFZDEqbSwtV0Bv2X0ycvCmcbs+lN
bcpI0o0w+WKI06mwO09EVZjrk6aJeD0y7ODyRWJP1pMVaNLK+xxzJKZKHon+YR77fVPSSRxlFssX
MgAS9zFYhbgbecNI9omeeOnSA7h5HfSnSjM2LaS/sQQaTZbBAoK2UkcUb/2PkkTB83oP/twIaXHP
cAXl+hiMyh2sINXHyLKAG5xhHG83u3mxsdMfRPwng55p81o2M+XUu47IbuRiKAUGfa1PASupwPUm
e3/jBZbxEeU+qSrX9ZSejr0FBnSx9jcN7rSqISRvJPAsBHdNSMtBRaj0SDYlomFH9S7tny/1v2nI
pMJk+RdWIL9rNq0mrhM95MFA38JVhDGCGEhQwuxH4sE/JSFEaceFLuhQzD6+TptuHANeJ4C/6UDX
omc3Tz3/KHjxhd2YzxW3sQQPMrbweMH7/dyD0LrZjexsDKKr8XRBDtpszonKwRofU74mKyQfWPNR
2FOgWQn1LCF1ezs2hEcdIAspNlFxUkGDbc93TF1HcnJQ+rpnBKOvi8s/6rKx8OVBI5m9nydbNqX3
oU/K6NJjW2YR0JWlIi/yDB6enujnWYCIY3ubgPHlLSd1BN4RQUeGUzJpDW1os2Gruq2fQTcsWah0
9iu1xq7yL8fkQxlv98oF7sC8ebzwsfP876hqnfu1mo+n9AFc584/N7fXZTUfS5rUL9egtrP2OB4I
BeD8bMWjDUkn9lrMZpCnHQs+ukBHiAj5s93mzx2122BhkHbtHfxV90/diEfOcmGPUV/szQTub5To
Nqdja2fh2EZskff1iXZV6R/t7Q9HYtQt1wpYLw0ujUrbqnCtOV5A/o2M4JMQQjdI2duS+nu2fdBf
AvkxHLc0TrzGJ+hHllXiRxaycrg2e+mJ96CWB4zSHp5GGlFLOAVtnU9mh5iwFk1vlyURfYuk2n1F
PqBQQlVMtFBbPSOiK/3EuaVacXWljnqgTgs+nO5P6/dAMap0rjEZVqbhAGBy5ywvZghG2by5o9xC
GTL21C/zpHQO2Q7l+cYGRCtZbILuOuA7B6l79dw3mUIKqaTkpDzE5qwXcYX/+JvFTOZLhLX62oFF
8XO7s8k8Rz9oovqmIy8xzqIEUa/KZ3ZWwZvw4AJ39QHxHSfmoJDsk4qTsClPP1JjOOHcWeh6b6gS
rSeEXnorA2JRMTUJQ+g2ReVAgK6V9a/GaEAZX3b+1+xlI+x85ebZD+LI8crX1oNFDahyu3Gb5ybY
EyrjO77YUVlxOG4RqYLBd52rCVO2326bx/za68a1VlfFOlbpv3TDXcjXiMM7L7wEQUDB6fcg5s8h
nLgsnk9t+HtcIOxqUjma96Pd3VbD07kPTbPYsJK1DRRU2WjdOutjOoY2utlQt7h083Uv5yG82C8o
SmnbrG/Zyps9cQCx+Nlok+9fG6Cpr2vMQZJMJ98gQZyqpz09//I4nxITOZyo9N+toBRGSIN8jMLk
561MjHsn2XiBC8/Sxl9UoSKtdvZoqwqLqpGyoKxklpSpNoO23hNpCZDNwGxLpuBgXOHA1mM1vtnR
JOcoRD18jRr0IFBCi7nUXPRQrc+Ph6bttLhespgU9hh0dbMFkjhifTOscQQDXGLSIJh+5lju9t3t
MsNCo/A2Kek5u9EhRw+7b5yEHNFbpB1i9XSkq1LjX3rjLwKjxpaSKSN8c4EBJ/TQhDDIT62JAf3G
nNwVSRJ4ob7Wo8WVAf2GBT0MKW9OOriAtn2F3ZqwCj9jvZmIYDQ0Ly1puVhPNQ/4iSOtnfM9bVT1
LAn3e4rLiCn84d6Qg79jF9bYXQkxxshDAEH99Qh4Zs6gdREhQbyPYCmZJJ2ADqe9B0Ye1mhTdyBE
EX1xB2kbXXTo1xsTG3b0ddtYUGiHGGplkr4wTyweucVeMzKNyv1DMh0CMC8eK7O4y3HDtQNW1udE
z6SeIAE8Yyub6vy4XTieOueVRjq3/prDhAVsysMv9mNrzIoD/p/f/ar8/WmHZ+MvGExhCEhDm5ed
0TyvW2tUKZoj5+tZPeAc46X6KnsDC0UtCQNrEdmHZXvpBNO3eDpFK67CZDQ/vcD75XOaGQjRGfIc
V54PTJ+kfvX9wqRzhtUVH0dCAmBqXZIxrRKIszMqm+/c6xFdBr573Vw+RaL6oKSQmczZENNCzTHw
nlTST1mR2K1BpqHo4Hd9QrN8fpSdQ9agEFZIrPz/ghky9tIDMBYso/llLlzZsW55M4dy+j0PZR7y
cN5ltjMt+ZLz5tjGcV32MgQrhZwPKWj/mALglZbYbrMmB5ELXcx429Bdtmltqi2VLWAxkiX/fbaq
+Lr1J5kKdW4f7XmZ2NrNEhar6LRvt5a26YgfuqmT8ywAAAV4wI1uSbfl6j0E7+bINR3vAzUYbeq9
xjuRhJzI0t5II0V77WM/9fN4MqWc2k5IpwGHea6lVZDv/rMWRG1s/RIOnyXosZVzxb1KkZ3qjoRI
kMY8S+p79vy2UC0XUUSCLKW2+gZPnfVZmyczk7XCItHtpzP52V4Vcfz/puUJdw6n+CMbSru2TVVC
8T+0DE6gSCny+UsrXN22fih4RdygQaFdc8VFO/EVbI3eNxfLYb1uRKi2953wQXZ7Pufi8ldsa6Pu
3KSy4xJF1dmTf2Y75QWkyRipNaEbKS5CaW02SK2RG5Anttla7hb8XANuNcK6q90WRucqRr9XmyGA
azG9+INxaHyxQI3WKYRijGU4GeQEn3YYI7oliVPbaGNWnUY+GXEmy4UWLbto4r4hps92JRtbTNd1
oWUKE6wRyuMZyOVSuhozpAqjDk3xjq5qs1y2YYJRNm8iAJi7pHUgMH9tqi2NSt1rTwwLa/fTPner
9Jioo902v945Fgv3AimMaEczF5saz3eaksuM9BlWkpl+i8hVfIa1Bh9pNb4wAw7rBaVOsiAyK+L8
MaeD1DA0gUQ0zP8rnJqD9+jBm5OidibBzeTkmvOzZZz+bcih1BzzuwdIT1sIk5qwOmpzoSJfOHGq
v/4ZfgWl0+Ln5PeqGRZ68ZmvjgcYAJxi5frId4jtzwM/B0VUbVr559IhQr8QWVIEHntPCnCpz3iE
wH1go+J8vZHC86A5F2MT7NehlutIuk4Xc5q9U7NbGNan2JcEX28v8pOP7V2UsLe7ZvoPC6t8A7fi
5nvuziqOdIR32xe/eU/4uu6O/PMTxCR3QA9LJwUYeYzz64qwZArhjwHYD+ihwNio4CuEsqd5yaKX
NupFVlWb9DSgxfxygAS7f72DRvjb3xqazEHxOnPZUhcv2aYtJ+7Hqxe1H/BQj/TyeHrsEK7JxKJ9
MaMcz60UGAPfV4iYpqbRdTD/T2RbYrAp3K/YeSmOxLuBE9YeOGYRGAUKX767/cRdG2PVm5d0W9UX
eRND43Unat6Xy5fV90GZObq8DxUokhZilSS6PVALfqfYEg5S7lw4bMW/CU6tpArdYx2tHHcznD2n
CyW5HwHtwf1GHuqwd8tug/I88YxHFSZnycufwWEsNR04PT2QLzDbqUoZwZi8MICz0V58p0/EbWoe
dm6xkhtAXifRlyxmbrccL+wIdwxR88nwCoL3k2PRLtjYjNYYSXd4bHcCxUlFuy5HWmAU1jlRB1xL
Yi/tVi12p5tblqPi5iNwu3GAtJqao02+zXbo1co9uVPlXNmyfdjQe4EzwJfMply9yQ69Tg0H7RMK
uIqEpSMnQ36SsarKOVA8n4HDvFfInlHVEcfwhYuTPAfOc0zk+yizfhYiouZJ9q1JB+Glv0dguLMJ
yQ3P0PcSyTXL5q9evCEFlKG6uZJEGdmp25q916lnqYj038VlE4KTaZJ9gU68OwJf/GCaGsfDgjVY
YH+/vqYUPJFWL22nxC/LtNmaZiY/wZoR3AteByeJ1r+LdaJci/kXfPhp/WNlxVL8Q7q3hIdzpDOH
+CROy9DERGRaxqyZFmmnNgTq1E0kFuXlncCIk+EA1cknPdMqV5BNKVWvmJUdWj80oke1dlLpUehw
LQxw9cKom/VJqTQBaBAT4OuZ1+iwMGGTfdQpBTaqrL7Dhls678j/eBdxCfACXhwLSefLyNULIRgG
BG3pHavts/ThqZ8JDFn8lhj8XCoRk80beBuFSN37ncF5a0IvktdZFFsWMA4H0Hi+ukt2Td4HFg3m
i00t7OSdqsRRZwxK1EGq63wd6fdMif++6h4OePu1wAIf5+nHvNxtLEBQO5+6s6+mUpQiYmgZZ+V0
Ohatchy5dSGeL0Yoiu595nisa6EJO7acCq+TZB5407ybrY8QAwsHfXJe1PzKs5BbAUbNAUaXcEHK
/QO+dxX+cBLfp7kPADSGkpXAlIVHW48czp28PpipdskM6L8eMfe388icMN1jWFjxDZeSX0uEtBYd
KU8XssTIQM2E2fTibaxk8nFm+D9Rk++iLNHNer+QaK5Y5ZA5mFFdEaalhRgxE0S+DEn2heu1qnn2
HxsjVClyxuaRJkcTTx/onsTx2awfw90jn1RWcWuk0Hm9aWAdWIusEeHEw+ErefeHYuBlHAwmTBrP
um2swJxejfeu7sFAea9R+7neKk6LqYf6cMWDJfZFSGo0zKchm0lBEXZOwcjfLGZKhbQ0cZuDvqMo
xkTXSNnRkgc0x+0ZsBX+HxO43bFh1njF8Jpz8CmMvkrrFrDawfC1SFdbMJXxFVbj2Z6XGIgzpdPP
eK2Id/NHzLEQPhqgpVFCzS2+cbm+WdSuASh5w75TL1O6MqXXupiEBLQ5TUknx6OLuSeGvNYhJM2b
9tH0SnvI30jQCrbMhPFk4ObEte2L4pisHKRZwEErnpRfsbC40H3bRxTQpy+/uOXsR7V3YwdmLcOE
9h+bBp1732kIlLGjyFN51fpHxGFdICgiAWHTosmr4khzdBh7iJZS+kssVE7ARV3fAzem7WHrfcGG
1EM0IX3Q9o3+0OnnFYGuWIY/TE66zBYwpFoRVDMFqNU5JCF3+wk2GuuAorBkAosepJ7NAvInHP7+
Pka8vSi7Xkhri0T2hw4qjdvcY7acnNzrSbk6S1cE3TR2B2yB+0vRuZsIaPNyhswQKz+vH/L5SKBI
KLsRg1jPAT3KcoF1Suf5ttt4n1cmGXMOV8ywBKAdBhRjUX1PR0xLJvj+Ve6B22qYdSrzmLNVjghY
yJ+cZiR25dcyOFN5PpivhhIRshvQoluuduthZyWzFYB4Ir4w8ST343+aq033ylFoo/vBZ89Unkup
FnUTlFBpOg3ttERVrvtM9eS3mpQFj+xCrejyyOWx8Sxh7M24lfpv8kgCg6AdowyY8bJ5YcAhV3Oa
yihG8d8JDJis40Ov5C32mL5WxvhEYBAgbDONjJK68EgMa2BOcPQDO9X5jdyQhkupmjPpXtxEbYDy
NeiMFl9edKQywtrDbIBFgxK9NzCvKq5Z59uybi00+Qs3Ujpwk8GRlUU1jz5SGZt0IX1P4e5Ahfnb
0URgLfLC0HPJCOumXVVHNdRymOgfhzjrrjC6s4lTpOb2eZQB6C4HhV39q327YrYhktuW2iKX0CEH
e76PwKm6IQ5/AEke7euAdZim6HF9rV2UQL2+nR2i2Soi2JPfYkvhRbSmLTrp/j50asC57MrQJPho
/JAjo0GACqMwcoeRdQ7RWtUY7VFlff3Z0sAr3XsMotCe9zyXIbF0jYzNMc6tFf6BCd/U8sDoBoSA
GCWslemYi4xXdxe7f7jrz8SQE+lQGszmsOrb+Kb42kT6OzZ+Dq9sJhgYt+qoRIGRpGIml8Rez732
p9/nvWfAUwCUZ8uWoyJS0rtOuwanJVm8UG9gAc5BwrfVbJ31gPVGyE5ON0ckRVceIYJ2NTJNdMeg
ROtWveKH2dJdvKyfRnr2vK9hsd6LM549lKe/4CtxAdy35+GnKee1E/F0bXAk6ItQ2CcE6/g7KStM
e7i5ElBumFyamp8VHHDvQXeqoSGjzacub4vheTIJmdtvJh2lFZcQXHV3SVzpJ7Gp1HW0fsEQJoTv
LNz8k+vWtQCCgKhF6PvJa3G69qsrgsGfvMyHKQxrCta3S8QyflMsD+PbqsErsxoP24PhJIfQTWlF
gzeq86GnAKeCGqgx9JppR68X12H4ldB5l9tQ66dCruxzf5lVRY4Qj7RbMSeKVu0w6gJXDDeFqS+G
G2OhQ4JE1v6bWQ8zsTciRgnAGtcz7VGs5cYOf1r7Mf5xW1Pa1lAUguMoOYg7CdPWFGpOU+e1eF1a
//ilX1u3DavqM2UKoLDIBPlLL6kTxvLBYTXZ1WOtRp+ZFC83ueKGjfvF0Bx1MSNbeabwp2QmWesb
LQTVxVEaTIlmX3lOxCcsU62ByryNtWooNifH0IPfC6jWYRk+aDnNVUt7g/YMdzfE3hT8NGIbaEXr
neaPL5Vj1QIySMNJEowgkFASd4ApZLPYpQ9F9eF8Qoe2L7SM0rKr7d5jdzYkDb68V8KcKzMa5ISQ
5ImR/DztEB1uXptXvqAseEdriBywJj9j69yueovqXilW2YoIjag+3VesyX6x8nLY3uwsujKGPcdj
3v6PIMBLry3MQ2TbYEPzKL/6u4ZhHYRnPW2V06Pf2GaFnSyzGadPLwKEVWKvmzgSWHeb1uWPSjHR
lUDJzIJDJLDXIQK9gzbzQ73BcWgKCYytcvYLqjSEdHqzjoJrosF+Je5vl/0MKERD5ecqdizfKBSh
4oxvH3C15VX0UHiAgMBU44llqFBeueMwXray2FoP3C3jGUwL1wuRvxg0cK6AK/7YZMHWzLVQ9vq2
X+lZSspHtCkL157Cf9uF6kzYzwDdUgpdgOLFIGng5sSxBqxLlZDMshYSWpfWrc1COkwR9q10soOn
u306Qx5oqvhdpknIml3FHBNFJMRVWhttLBxiSGWk8H2j9TXMiQDBbWp/2QGencgecoyvljYqFXIY
ChofAO0z8zmrEXsB2nhBqLSGhTFfl19BOlbKwH2I9C4Y4LfkNz4uh2eYNi+e2W7Btd/CQdgR+IJq
HcKPAsizRbeu3yeg+PU99ahZ3IEEdPmJLDVP04FFPRe4oRIn55o1aXd/JrrLJ7w8xuBwIEaSDPh3
HMz/nlyqFNAoEH1+vLLJ9Yc3KSuYtiD5t2MkBmV3WC1VdYMaTadFgA5cEGgUKpeSwurU20m8HS31
x+IwNmpoCjZ41zwJPu6k7yg9DEFbxFe4kI5QtSwqgWO0dZmQ8IcWZgSmcroGW6oJIDwLQIhuIRKh
XEs6697obfrQUCrzIB536LeCEGu0Dxi1tnTccBPBIrc5o3FGT+9DCW0HntZegiqDJw9SE2n8H4CB
vsD/Pj7kXNiQOFQk9fZqu/Etz9n66a9BzmyKhujohtMgUIXjaFq5Blj30v7l4oHqTJMdqBEEEZHB
xQBeQ2IB+pEKuxgpli/7KCb8HLOAUThwtQvtsz9E/8hYxZoyGbFc3rgCKgvejqk259e/qcVaYrIx
4UysvAWHXlConSeS/w42BPi/MhAJL9hiqJUpLcsXTo/KNvDxfpg/5O+Vsy9i3S1/xDIui1ylFaV5
RaAvkdNKrqKKGFsuNBLFpCqxYdsdKoASOXEhnw8s70w5W5YUpR6TwmXXYGgepFVTCUCb0x54ebpP
r/2viCI3j4ey+dDvvlALjIrVfhlfxNjsQku5FX+bGPzRfdvcUAnA9rrsqkwyCJdQV0Vz6bOPawH0
lp9Xmzlstl1GA+TbFVtxQR8LCB4KACYH5gwcIlWfsZ3Vcc2kkoVSNsAhJRjXVXJsunmGt2Jk0gQM
pKEAIw08NGqIQGSrr0zWRqWWSToq5ieMb84yre25S0JTbi+l/BTGz5AmM90jmNnWzHki7J1uiCYY
89EDaMtgxJQ2sp1/TMYMhDJDrP77LkhDUJrQE0hMu1qLBBCGpbja2vTbof9ArvTUV+lJFJJS0bRg
L1IqNYqXJgN/PwoqYDNpzv539hi8ZO+3dyGb6Bk3MAAFFrX4qnGY29qKMrpWCe3TFJZVpeTsE78N
61fzOzPNYJMZcbIt1WbdZJ0yf/bor5DLrIlGDa8FwIKOkEr4MB3Wuv+STr29xiO85EyxSL3uiKAY
ceTAGDeVTU5rV5B3/YuFJkvBP7CyaA+rtHKpdID+HDPEEW9f9hod/81ap/KTXN+uT0mWsWO6cFXu
mGWfQrbJkjMPUABn9uH4USXxzW0Iw17z+Ll6KY95bVceye1TRWs/6KXTd611GrirQJjKOYIIvhxu
iS0hu3qU3x6oUwqGBFGKtL+KIdtbvFUUZKAWGw+pCv2Pvduui9/mmXDqq9RlewA6p8sVAeq9dsxN
jiRgd/0jXoF/w7TR7fVt6psxCwfGwD4iJXaghD4SZmf9/0SZ0IKSyODrQCiXJX3WvqGwce+PBHsE
qnPivOjDHAVo1H0KpEzfm2F6CLJnBOz1Ze+D20oC52NqF3dOJ/6gfBA0IFOhaZeYJ3lCoilpJ/Iz
EVbLdqIGpKwktFMRePP34hHVbgcE98s0Da4niDFYDExgdnwXSThvdC6YRSyQ+h1pfghPk6fnqSQB
/FVHL13PvK/niL3kuLRbICni6QDalnKsa+s5or2zunNdu8Ox/fE+pOOikp60PdwMG5eRJ1lFZpwX
P216HdTeJMKcrvWNcfnp5/bmpDxhqY33aaw7CaJjd1jj0+ViGj9hSP8ilReMPSkCo9pJghJHFeCP
3nERipa5Ob0MzgSuxDxGs9ECSsaFOE/IQFkacqRatkfPvXrCnL6RQuxRXbekQ0by+cHhmcXcROo1
zF8fFp5Z76yarbCMbVAA6CdbZnLrRmMx1YJRW+KV3ywZYZRRWhcKwCvMEwG/nYH2GMJgKJNYFKXZ
q6g4H12q6VyV7SDBumle0X99f9LQfDm4t8jnazrRzyUlmTMOCXZtUq95+3eR12ovSgBxwjx/8Fq4
BVLSZ9XRgawE/B0ghjDVAnUTCI4BBbiBRHiN+e/2ZvWYg79LGlU99+hXcXsaGyggM0gpGD5Fuaql
5PPgfSlAwE0c/vYFXwZHtjXchFWvEO5di7+qnMOdElyiuHZ6lV3wUaYRWJEMnmieRt/4SxOKYHWl
pTeK3H8Epq4izwoQzcKk58r6i7DLuGQDkssGs2hID8LS71HJ569rhMEdBJ216LL2sI3otM2qNMA6
/TPZR9lya3BmZsMfploEln2nF+KuSBMj/737GuYYOq5H0eUPtoVdgXhsubWY8E2pzBH9y5kKSIqp
2mhdFywMXLBYwEm0Cc349Bl6CrK6RMErRq1MFhHhnKFpLYcMqBg9dhqILJqVhy4jTPZqLvjdH8BR
BsaxwNFBhOyp0rSJQmSdkhglS3xm3+4QT16tXc5tLqMM6BzK1LX4T9BwybUOortIuzoX/OXXvuW/
vNO5wDIWDJMj6ZgQzapP6RJqmTqofzDKwPvuq9HMv8V3BO3ufgoVZTPQ0BQKvd8jwPQKI5l0TD/7
V/lbYHyOWosFCm8nU797Aw9Z06WzO1vmIScundJAeCsVqgF+nLtz/rImRkfGOf43VtTxesfykEHg
pH8iaV30DOXCCumlWuMyoXZ13crpPtnUtBYVibZKjAMeA9dzAsCy3iTVUAW5hjNN8uOthIJXZes9
M4BPbnI6BtRD2khqzQerPdux32epabtDNoZo9+U+hHCdPgxyrcR796cL8wlxfNehXJKCAYhpjt+o
CRpTa/IVkaYDcYz98uWSyDumVDnhnyvSqvqxrhStQYRltVnd5y8BLHVskkFzl3OPLmtuij+qa3XY
QZwGdmEii+Ugfo15e79OXSf9SkWCdOSLJTGtJGEG4OlPIEU2WN9suicbQOErM0wtuO6LUaFFpHBB
iwK0CKzO0ez24wZh1lZiWvetO+iflq130O1RsXpMjqS+jcaO6LG2KcV6s/S+ta6MQf3mtGacdYMn
lJNRJNfxnD0zWd5/13TBn1cLaYaqiS6oCeNS0szeerd3/AVS9Tg8DuGuvh1wqTHquVp3OB7Cg9Lt
qS9Ym6jyXcJ6oieek84/HZmTZYpUjMQtrn0Ht4AVWG3eayjDJ4cdYXf3/AJ+uBt9Y/bp+XFpiqrv
cVROIAmjdHw6s/+USF64GpwndppBbrTjsPw1B7/7vry8+IyUxJo36b6rbNkHw1aOOQMgxVcka7pt
DpRt5/mQUOc3ezBrjIfq+UoJDFoxjQ0c1CpCyQ5IDMpHNpi4FyyFoPzTKMZIjiFBJO3mI1LkxvkK
zgJpX+eXIo9I8OZNbMHBYCYaiRx8U0tMKZfaD1oIpYgKpLDnHJh7cufILK/MQX2BzNi+LHbubPcW
JFY5RTjmD8h6DoUPZ8SseLgQPfHi5ZhlA7PsdhVMtc129kcdK4us542nOU2AyrSuCFcpUHJRQjs6
pF7ER/UGJ+JiJ7UJlWKNfZeP32PEGzqUlKyf0XzAwxCeX1qjDMHD9AyMOz+YwCY8CGZQfDQfyoBX
RiklwjwUvtv7olH6bmjcGhhhtkqbNYXUu7H0ixWVjMFqXMaA6BVKBXq5QBmSbVcuFcvOSIhWkVI6
Aq340Ch2qVclz2SBztmUchnGRPXfWiYWE3u8OVV7eNm5TSMiVMzlPOpKT9XlP0G6n5smxYtowasb
mmL1XG7HlSSi/nLKLKP++yHOXP+EsmzGr3HlLBN7xkFuNAP2tpiffLtqxF/yBhu9BbalUOG+Y4pN
N4g6Rf+2C/z2E8dQUsLseAEjyHcPuJD83xHzLRUncaEShGk8O4r+h8JypvOWYJ3WL9hB0Cc4syER
hXnT+9apQjPi8UG2eHEWK6hEkOz3hYvkoSlDlNCoSltgWBIuJ4lhlJYjOs4fx+wrkzUUs5bXxG0w
jO5UdBP0x1PCtqaxYyPn3LtzzneYBF+4sPi6dgZRPwa5gF6Foqx5lpQbKfBCImbfvh9ldqC0f8Pr
dmgoSLedz4q6PZzPUXVOA/YtN8WGsfnZOlW7U+vmS8YfYyd+6a2mCJTZ4NkSYNPt/DLHKK2IHPnG
S9sdFb0wzs5d1f35jBF/wDH/j76ZHNCRgRuuyy7aREpqVPvMD4qsygcFa4NFAmJ1d8EIcLsnAYGD
y1+Ai8uhzPFZKeaJqhtkyKH8bY5D3MqW1qwyzseypQ4/OCLxvt9iLD2C+Gcws89EtPqW9qqCdPv2
00u0uY3iYDGCW3N7wwY/IWM9Zih4fTohAWYeAZ1O0d/awAoYXMy69LFvQo8X7/ORcNfECEHQonCT
HWjYVO88kIeV7b1JbaDvafoSHGSdc1WDpbhZchOvcoHyPBGwNP5eUTskLu/Tej3lbdWTvo+zGHa6
Qh1lFd7FkhZjbhOjm+zUKAKkKm/MuqjsVWx1F7PZ2KadaO7eW+ztDmkLx39TPwLAedCDGy9soF1r
xu5ju+NVtSoacbEl5t23Pp29pUcxflgPkP+kHBjJZ5isY28Wqw/1cXhZZSpZcPoIlVI5Tc60GAz/
HK+3tRZJkFpNxRWd24FjXP1NR3Ll5p2Kx3qra1pOM9udDefe05fqroH94x99gsTppMYnW3KnAyHv
Y2Mz4OUgI5HBCzXEDIKBAhLZBDGJ6c7abbAnDQsZ026awqPyGOdG/38GSfeTvV89aQ2DMSwGszZ7
EGF57ZfBMpLz8wsKl2KgXiZagErf1uQfGA1h7hMst9yXMaT4tP95N4ZSLsMmvDIriV5BWGB/tXGo
Pw3c+8sPq7Cl5o7GJjfJ4I8QSAo6UKuDLAyQp+zHB1zFrzFiJr4gJepIYll27vvH48uquavKCArz
6xn3Wr5I0ofQ+3syj9VE4+4MHRpVgziHArvxyWIFZVte9vI9foSc10+g+q6ySMabanzNAaJKGuZF
MUp8IBcCkEPPQX9fJ6AR4AATUOCk7gTMm+UPtk7jXORbyFJUl2oHGXiozCWEt/2BpUODVop6ESUt
ppH3VwP/H7Ud5Rn6WjAlX3E/gVCVU2NEz1iE3PI9C/qPC2RbCak65sUHjS/2o0KNI1dqU2vt2DyH
WH4v4oqiSXtg3NBG5O6Omjh6lC7QcFIyuY7ylZuBqxPbAVoTUmRmcklB13Lce40WSN7w10latD/n
QAZ6YCeVOrCwKkYGkuWhOakodEJI4c6pT0SyHeNsa+B7xR9Q2D+awvxM4PhkBstH5sIxSLE1UeTH
q38LyJvqQRirdLs1GJwxdvlpYjAP/+1+nH8Eb12J57Irf1eApx8tqAPz3O2Ip0M4TcmoVyjUIXS1
Ja5UFdvso3pdtKh41klVq+1YafpTTT+9+ep0IXieNwCm796BhlkvX2HlrUOBU4FAIsnwu2lkB2KT
g5a4/lPVCD/XOi5H4RbBdlWPunqPxUSbDQCVFOmKG2lt1MozbF/Xmwz4E652JN3AKA6a12OgqSj0
FqQlC8Mw9DXTZXgPwMVUCvhRVreO+yBK8p/oT7xduZDS0UHjiMKHKFM4aJ0NgcXKqZvJoNJGGMqk
5+/7pVnJGLEDfoFWmCOQYWFxrf9dP++bUJvB+g/crf9NVsD9+aPOgl5LbCa9n7vG7o+kDVLTLLru
jTLUBKD37GKPW59XC3xH4l+LnhQdPQ2cPU2umkNZVSA7o0YIwwYhqD2FXp5XT/qEcZ+Pedl5660M
++hA5g/jabj6E1aIb91yiesIUi6wGpQJ3Gg34XGRVYnMawfH1rU98Oh/B7MiHxA5JJwW83ZdeShE
tAI2Qk1CWmZoNALIlXBPARTespWCEZIFZlNCv4siwdrS+WVJylt/donx7CdZRP2QjVey7BgnaWEz
KbOZzLGksLhHj0t2kZm3/YfWY4eijob3NXWCOa0QvIl4AGNnvWdwpoBLPK7S3Hp4yUiGbyZnVJHG
kok3FSprw/BfcKXtEy5Hcj7lrcxK8AUwMkN9hBbufdom/RLzSS4EQHbUZZ8EuGllHn/i1b+7i60H
xtKQB8APm98ub0mfRvkHOOw34rsd8Mk0BS6EBmc0+leR+nmgFfFFOqvQSwVELYEKBYHlrvCItxys
gCNP2FtrOXasonNwT+9ofBvPXa4W6L6r3yC9pnqnLpn8VJDqQMyQPmH/TyhRoEnP5ObNXBkT99cb
LZUvt/xqpIK1YrebOO/VspSY1IjTPevJOWXkY7NuWTi0kXsxMv09IYNJU6/2rStJWDHvCw/eup/g
Yu1AaMt6wwQDE6cw19D3M8YrRtYIHxA0XfXuaSbhmBrEIEz8i1yDkwscyW/hJmECZf8mPU2SK3Nj
VVXokmkuzAzuUumkkkVsAbPLiXBBaQwv6DT2YNxI4bv9deUBHFEbEdtUUhib4qjWNIJaoHKv+lKc
6IRa0aQ+5izZM7kA55eb9N2ZjmmtascTLRo17Zmwg5DEMgvmPsgvSrW076C5oKn5JZLKTSw0Dsem
ZPHmbwS4XqMoaAgr/ysu3o/YQSS/VXfcJCwyNEE5tn9ft3BNxfqzhSKIquWB/Fqb6JoLfAQ4iiDj
GFFxYZYtzFLlaVV3Teuf/kV8JEuiEaJXCwtEGdQ3Y8uj+5EbdvSc9Klh4SoTwzf2S8heoFev6QdL
Ca8LImgetGvg9ewrLd6VSW+21i4EKTWW8TCBOIkr1ue4GKiW/+GztHLNva1B4t5rVM+r2PUCWYwa
chinuJqFIBxER0oQdYV8sKDDVGyJI5fQLJu1mZl1GCPzaD0nr3m4+ZjZRqzdC4pdzGiUdGSoA6MT
4zpepA7CQ0+f1pUvA9f9lGdUCQd34vSJC0DZSGo2alNl1dTmR4efd4DIFOvxYX6YeOwQEIzIeaog
JtDG7XP1jCCskOxU+9wBlG2Roj8kxjOtrZN4Vcbsau7zHsLok/Hl7esZm5F30o3mVqIElCzyDDME
3Uqlaat4dLWldV0G9ILF+PqiH+AbGFD7uKYF2EvJ0gj9ajvpWLNnvIe/8M5JJa2MGw79wQ5TM2j0
sszXRsXjFa95rKCVAhc7qT0v5KTujloD0Of+texL2bcqhHfflzMpBEo1DrYbfRE2P6MWkldYj2mS
qfylP9Fou8JfzCIPhJ2Vps/2ftiEBFi0y6Hr99+YLIF7WWNu0uPz/nQ59hL3gVkrwTCkDG5jggcz
FDhvXUOM+MlcjemuNwWySh+bpyiQg1qr6qd4RpOiT7v34aHl9bJfIcZfBNRu0RIr+GWlLR6a1jsQ
HyO/dWu822QGhCg9c92EHTB30vyZFW9WrmHHe+u6mv8lFBMLE52Oue0t/8VP0nhFBBUMA4QpK58G
LgUgsARENKa3nIu1UVcn0ZaajJaf6XAp0My2+AhJJABoA4EMR8fLUKdFV4uL7CNNVcxDS6GBGV0q
i27O39/uyN0egNWvAi5h5MyQGNvxNiz7QoJhm+D6PSCbZuRZRxhXt4iidbVQYKk9cRfdxo1vjr88
gkvY93DAYN3vsPUuj4I5EVJwXHxfqpm9LhUQw4TAj7P+k2nN60OcqR+RcPQpaQWHINCQC3y4/s7s
IZokQVRoM1zCwUs6rebzEx/jrkG/bmaaGkwOjJBDeVGps8sXiTQ3g3EAdEnhtF0gGi+BF1vOISkl
TRacbKF5rZlSovCEk5/pDs9zjMUpvvrbPaH+W1GDfD0HpD2v9FDeAZ2nZ8Lez3iCnfiq/7qxWRIK
J04JksgmmV+kGoqYOZjbr6L2HeZHXE8dG+Ox8T3PUX+g77p23RNJyaVh06s9x/UIZCwC8N6hLGqZ
BiOdOMGrevqrxWnQQAlo7gGXm+5xZEYBzJtyyPs6781aPCrHuvARzXbsEZ4lGLj9KU17ioX+LMrV
X+8fmsnFNgXoNmlMOBiK/JKLtwYBUHG3LqxiP6mERrK3tKJ9UFG0epeiBXW2Zq782/qAKHX1uoSL
R7mi+I3MsY4EU1UmDWxJA06frgmjyZU8PU7vVm+wt+kiII3cnd/x3RS5qr5TRB5eMcjCFe70gQAx
Wu8sG5fo1c6pFr3kvDtFOI2vRc/tKFy7xOb9v71czD5oS8hV4fMXDIAHYkANRoUd0dY3qN+RGMou
4Xo88GKvdRFFA2qDj+bXtrqeMFoiz/Pso1IFczF9I9VTtP/mcvpLfSONe7TfuD9Qo1SM+pSl3J54
+vyELeAJYxDSwijzaFbf1WQ/Rlyopfjne/ZHrKw/edsMYe/zNlhNvqCGkry5SNZ0sODW6TNw9eu0
6Z5K3um+DoJAufI/ApCuQHxG5UVSvMNRwQ9HzYzmdO/LqywYis1jnA/Rwrhmu2h4Ci9MmH30CVph
JMjez02zOntpx8RPsVKzDZ9fd4OoAGxLgNZsh0N0G2fjnSotj5Qz/MWHuoXNLAnuk8TgiXmHe0eq
TApI0gvZStJVGoBHznz7eWDtac3TVl5TKILe8O0wlDxVxMgt/Chr4DmAfZ+uDpBK9xQqIR9FLDHf
rBqQ5IZQujMiz9obHY78JIvE92tlZO4lnPyUS/R0E3kdkM/CwRro3jqd0X5JGe9gmbyjsbzGDCuR
CvdpokJButXdjAOwVa9Liw35e3r1++WkRX4n0Oh+KHml2bnNKuuihy8TcjcHctVXatUaKxLvr1d2
WAFRPrPXxT4bSwMvo1nrkbbCmAMdt4LZd1XRKsw6vZoxMQpxWTFhrgWHS3SVhCj5oTWGmEDSXKJu
3qY8rgdQFbIdrG7DHj+HkeOgiOkiyRo9J+rR9TZvQxDmiOn0p3Oi+juM4QaUmrOjva4Rnj51Kg4f
zcNZQc+4Wcwx9m6pMd70BGCjLwvVXmxBIjjkaTGtPmDmakyUvyDDcwWs1vn2d6GR1Q52pauhTZea
PMCGiGtAGHrBrTc3+Glc4R5TZNbUr5eLsT+0fmZl+hJE9RhiwxDWOLfKDwJtd4pZhPYErVQZa9g8
WLzdVzIwjZwYw51LPqGFL1n5NP5psM2uWH+0WVCmdWTvNdSHfK4h5iC1j0+X4LpyuUzYXJZV75W7
iODIziKQ6+kFkbtWSa2pzE8YzFlaSCeEFBz71DqJd494s24Tv3829zy4/mBVO4mIj+Rqg4Uhotfc
/PX3thTIaKrsQwLhhWVuWsmrdn6p3XoQNL3lI7s8LSU2x+5lG1kc5LhcKnv+3h33pJHRxVIZR9bZ
Qw+OEk69aTPfKa2ohZIvlQtb4WTmijdGd2oxirfAY8e07dH4olO6nrEzdBBAcOtyU2w0k5cEvhar
VRHLNWFPG4JKY4K381wBMsgRpRxDIePwH4+TxT9NiBiVzIDB7JhFYz9vApPx7zkd7Bm3qDbOlA/+
MxtFMz4puxsXyPxweKGnT+5XuM7dAh73VxiN9nTy/Haq82/S01YL1rO1ilxOoG6mbXTytRwGI0Xx
iyfsD3aeIlCxQmk2+D35QHRl3I7yA1DSZM6TXYHFWKrwMH9esYoELUOUXz+mDbqlzqdGoNnwbquE
Ey3qmLcCtRtCp/bvnMqalG6VIMj4Fs5DpR0IZS+gizSJj9WJ0NjR4nE7KCfFvC0xIhyXVpFhAwdU
RvhosREfOd9v+pDxr3b4LIcXYYFylkIo04Srvx+hjAM4KcoCpCiRaBnWT29Vu4W8ZgaePL8rDVde
qxBdKAq6E2430oHkri+mC1O1oO3bNFqdZOrOpT4aq4KpsQnL1/T0dbCF8MTY4YEK4R/BBU62POhz
kDOedF3WUAhzRtE10LPSNjYF+M8NsDF51XWMk6/+n1BQSsmz7gqi5f65FMlejXPreekJMUGCRmrw
i8ODtQl9kGNJu9lM/33N0gfqLIvvTqfI6/BpyyAOEUFuWrlh8WBvRogD7hcKiMJkMH3TdRjE+5KE
gMsovApN37vpiOwelOAHtRZRJcIS65YKpUgpjcmd0k/OAJ+l1Uj/tVRQitmFbPhl+stlVWtMbzMO
ya0qKppkCda5SKNDYAMXN5Z07flutBPbsuqwVphV8utzffQFY4EJkmr5Bd1sGUdGEU/Wf6TiccAu
iNsUvnuL5d/iRtygxeKsjnb+dyuENT2wk5DC5z8968hGqwhp+7WxlOfjX10hRqO/uL1tuiMK+eej
E7Qg0Xj8WGYmVhaTpS0i9zdgYg274+/gqFJ8EcCewPTmcBs8XQ1rfhI0Svu8ClKu1UX4W+Fh3xRx
hLwbHBYT7MG/1Ra3Br1MJ6TAdwjUhR3vM99o9kG5lKcvRUTfA9/3DLxfV/6Lv2AFpMT9HLpZR9a3
Gx8hXOSPmL3xnjhoktfY5Otxoj9HmD1aPBFlr8IIE9H9ELfW84cN52x4Hb0mqo/z+9tk9cGNehC+
Rjrv3FCOrxdeyINaYLH989wVlaw8stv27rNdTL+74LLcM9t5eJWpdPEQLY9CLQEp//GWAoaNCoED
37MWdutEfXyfXXE8K3qYWmOuDDtLlbIFmgZ/LsSRLbUQPyhpPjJQ+c9y3ohmSPoOB4O+sLWDxe3A
ZGhdqb0J37snKEWSwzORDRwAjKm2xUzHEjHQQg1hjsDIT0YbqGZsZLsZ9A5/XUjupN81EIdQoS/+
Mt7hGUj72/jAblg6EUDe2ozY2xtBe2iNPGHW94smIeDZBpex+GYzkKlaxqW42ZcrhwVF1Rx/jtL+
Yu1U1PIEg1PtYsOHEuea/L0WXuEhhvheTagMTNiri60mHo0bKzdd6/obF7WmVC0I+hmNDSEw4CtB
CJFFMJC+pwLjESAhD3bQ3AFp/ebkin2loT1ZAzSoh3ZNE2Tws34uUnT89QneehY5fcQOIlKqOVGe
pnUP1UwgFEmR+VniqEiDkaLYbl6QwyKWFS/dxHy7Z/yrbYMVcL6UbWfKpA+sUjfPkljJJxdCI7xq
yPWspK9MMH5A58Jq28honlPseMBn8CbWb15bxtGC0gH0v1+hsCafVKz/6lYIW0KyFuieiSsUiFz5
AV3N2uep7PnErsfbjnWQIujdLKG3a8gB8hYJI+m3sXe5AGKuIeWdz1Hf6/F7DOp88cdKmxZVMvt/
kLIrOllZPB0c38eizYu8oVu4YyOTMJvOrtX55ZwkpreBd97wGNYwVxemYn4v6U0HL0dvNO5R7C2q
0R2+NEux59Eq3nyxmMzjlYGX8O+BWmyaoCYKk3r980w/5abRmLBsPZabsTLLxpnQ6md1DHZGQhiL
3OFtE+uBqXiyzZ6FrtinzxSt4Wy2Dz/8WokuhaPdCEa8OwoMwvnKTLlZH7AP/gtIWXXSctyBY83D
I0i7OUVmJq2KdlX6H6ThDsOaMlszUwGJRgu1Y2Cy6NPNbwFL+gw67VOhTFPfIe+JJYSyZZ2W4efi
VYqJzZcO5HCXrxXZy6Zi0JTZoRHMNvlgX8Q5CROYcKzAyGvEbCBCpttW6rYJ1cx6NKwDIV35XNf/
2SQIjvZE6uZiE/1XqB7+ynwra3kYOMuQBfGjJeARzdFRlrCCO+CjtWmBNeVJi61dOb/cfcWOxZCg
uEvu4tOEYBNSL/lntQ1LulJwuZtMbqH8NbPJ7b328Qnh9mUdB2hai80NGZ5R9aXTbFiuu0c9iY3K
94whmOjR/Y/x3Nl0qMSgTTXPL/FO8GkmF9+fRtjF5KOCnPOEWkyPhK4/qvS+HvUctHf+eHfdpYvR
HKRrpm91ZDuF5EP3P4RA+vFnN5XzPmxB7LkBaDDayljDtRVlL+Oo9Wbo0IJxrOQqnOpCRUt+OMI9
3MHgv88Dudkno4r/+OIaYT+5DdVZcu0QeEJa8tNMBRqm0pvxU8WUw/YSU0eKMFcoD2jaZHvCCgtp
ZBbbiEMu+NBTpB4ppre6i0q4MyVQf2LZ858aYqf1YMFzCFW9bj6ZDoGCsvejryqdjYmhyWeUTW+f
ncpmCp/plYowJru/5J/Px21jOyj7yJCwG6h0V8hRblxAFZMJ8jFtzlEzYaj6jImZF1O7FNfth9cm
lHDM1uTYhmSBsgt4OdBo7GZhEXeIbZUdUL5w9xDdnHvS8rn8CQA7tytktXWyaptCZnawueKbNj/o
HM45QC1ZjM1TOcYxmjH86m8iFXviRV1VoBZ/4CsaqjG2lATQ+t5SPRJ9upZARHND+SkUfGYAVLZw
JnVU5O8l5lpfc0Wb9qmceae95ZmIdZVFnuJvf2E7n8CwyVTD2mKPebM4FHAyNS1gj+PuYIgtJxeb
x9uFgJ7u8iW3siK0r8/QAwlTWth8BT3DuTv+y+tKSOuaEi4erVMWwlRXpFJU/fw8gxhyP5doMbaK
xx8cTk7UL+ydNavfswtVJ8RR9fvEzA0CM5y/QmcL6HQXzsYkJO8hqEWfyd8nuJDDp/sZrrpTpgnI
hYJkxheJPYiLo1LS1lhioo3VJuApoACtUP6DfoGh5IMCyJQfU+yCOwLWkHYGbcQKY/uLrha2HE4Z
GWMf1xrTP1tkW7dBk/5Cq8x4QJSnL4fXKWXDyigacqRGHQn57/hbG8mtbEJmpj1JX+HImocFzlJe
qFt9vB3Pd32iFCCIn77GsaYJv2QnUyiB4W9W4MjMNZpQBfDzig1idjTmOu5YtM/MrdoY7sTvynsy
KgGhAnjcWMQqY0IBK9YhY3jYEPRpXDVg2enlE9KacMxl0d5FX9fcT0UjxqC8cMg11Lm9Y+DjMI3s
1+sWXN+r4rRxXuW+qpW+kQFsWeqXs9baaM9ZfuACT0Nas5h0QU3LcV+0rbNqXphD4Sqn9kx7XLwr
deJ+5aomif57G0u19GCkHUEQGjjx74kuveF6FLMwip6Y4T0LjlQLbZCfeNA7qTkFKwCr5DflcEHy
OyQ6zAbVgTtqcMuy8K4JNyqCnU1LrZeGbZgYKcDLbKRUWjs+Bi0ynLiwulcqE1WVMpmeLV0E7//v
oMY+jxfdNVRVkMnvfovw8EaNmVbkPEoru5Oh4XeEarkQLZx77BZQNnUclqsflQIDXlU7/yYwbCpO
ISH4F0CbOh7qrs9nfkBdKlKRq4qMJANdcLVJnzwvqOXEp9OP1wITwSsopsr7SiPVAzdinhUCw/T/
mSDSC6lEZijazCSJo31+4Dv7hqU7348PhRD95EB3TtGKQGBZ6EFkCuWxkX95bbSA4LSrLylfOpn9
1pO5Xz60P9nAfPJ9WzIU/y6U3B/MAvdaJndVLuKgdxYA6owulBza1P6iJoe6sTFNJnIRgh8xz92c
6fI1zEvjc6Z4ncbrYp8tPflcitCW1NmY5tKO+3HLB5Ct/o2nHvi287UiXtni1h1/ae95VIRK7lX6
nhzkYSNIMnumOQlRDrR+HZnK7Pj+DOuRuf928sQl/XhjbDgbzgFlx+I9xWpOuXJmuSEAzNDCs2q+
dC428ycMDPeKdZ+P274Z4kQQyHxXZdxAyKAmkEv5S/Asx7SW5+jpyPfmDO+h46nA2anmUnXVzvvT
aDmO6Zt3rsqA+1pf1MbaCoTc9KDU1/ZX5jf7ZKdzt9uHWgTaD+9k3qKtUVVwXgKmlCBIY3YAeXMj
YtC1KCvBXpXYW54xaQA21+Psnw4WrDklqYoKKS7ePaDdXtDCjY2jvrkYdcS1XFflYPlUVCbaqdhk
zzKv8liQ3AGAFiMbDnsP+IMw9BN/+ouEe8h2eCGlHgY5AJolKZ9Q6pxLvUaosJvxmO8x7Lbfz1kB
LGD/F3X0o4zge4w4GjZ1+NOYctzOKaWm7CNWsqB1k/k1KZOp0mYtLl7cNwhV+2hwQnO8pE6Kbq8Y
yqlv3ldWbql0QDR0yoGM+SXfDjZWInWvaHYXps68vbwviALMZX71luvr2btlx+1t0m3IxtaFK2E+
ayn42UPior6AXlNbDxGmTTGIjw7/IFFkzFFfXebvTyPiW6TUc5GKz9VB6IxKj2rtPB1VacB4tafQ
1g0w29Gj0nAs+PDz+QvvrNyp+pX0EjJJaJseVtY/CGD7DHygdhWbV7Ojdx/EzqgJP3JSXNDuJz1T
AeesDK5rVBlnHgEIQxBz2VPTgYMfz9UKz1R7CrmtlSJXXk+wEr8Ifu8bM6agQvLP8uwZFei/S0di
sC+tpo8COGzZrTkbeNQZz5Nw7DgL/fSf9kHsK2sEeiJnB5mQCrCFKPV2Hl39XvOzcwHIsWxsAdsF
fuVZiK7SixOuND4N03NWLhK3JZDzopwNSjm/Wv5eLuQArUU7CdZgb32VYxgKiijdT8fqB8pYFxox
kWMQOmb1IFJ44SQ/NXVYarKkh6ORHeUQANFk9e+cOCOJWqoU1II7R2hva73PMfmzfIbzX7+LX+3A
VWV0nsRuCyKcqyw+MfN+PW+rTqPwmeyqi/0Gp8xZ6rAkAuoJ9j4psX5tCZu5aaYihZvvERhv3AJU
SXSPmM9pAUQbnXVp1DquAARnycGCNKmS/8iVT2vpmsGuzpB2V7Cxfc+Eu/+UDzqnrW6/M+Pf7WbM
YJBdmMWZmGnR5qPCPQg58aAmJx/pxq1xejShCerd9/DGzq97ZaYZkAG2bkxRCFbVJVVTd4F59dEE
As5TpRS5phde19qXncYwRCLXKOEJc0FaIim4wqYd4BPIjh5bsxY+xl3+jOLER4ZWUgKw5S+ln0Nv
VFXpMEBWXCHT4UzoKEifJ90LpqvWbm4M9mG2FQSiYwaAHHHUSoCD37HZMYinl9ItKRXhzmK5EOru
l4llTCnNJ6q51woTm9xDFpsZJiYswXwykWrhDdW2MGx30Iiuw5xEVouX9TngHHkMx5GZclvfiUFD
DIhVFS/3HtZMmW0zIFoKstouY3nwQNCqX14tkAYxv0OnO/JlBJ3BsYG+GZFUVpNG1DzUNgWhKJk9
/6mmRrzA2/+rWeut7JsKp3OjQ+bjPXa4KyIQetvRvw8snNFTFqpWfm2gVD3btx3ekVMfMheDT7sl
I0pP8t0wrFXCJ5ruYRKZm19wek9Hcen0YUqnDnDR84Pe+ue3GQB9ZN6/AzlfhjGvyMPzd73UqWxl
glnoiwWZSUaN+5kO9QRlTqOn7xtgnO7PIMa0gpOdm9Ln0uKExMnvlZ1MBQjtpAvtsO19GlIYTP5q
3b7WRh8e5VUVsUA0hNHi4RzvCRAe8Z+gzez8MjorgTs9/8C9DpzbkxWh9Wp7BB+k4lO0qhZ8vQnA
9xigDZcpDer5zIfS8xjSlsI2TgAAMYqOnUUypf8leMYlBPx7/xLnH6ffKZChazqbHxko0Cb1Cme/
01hgjsUt2GXKIXh2W9MuPLMrY3H8a5KbfeHjj+S4iDcmSpEaUrt16y4/lM4KYOQwuV0n/3Nsb+J+
072Z+OlUAeeNgQ3PGlnhiBrjdhzBbFGbuWj6dJzl+298r2GQliRXc/8vjSEAqbXo5fP50yoKHjcf
PMazboqXXepflqBFc25GrgkNH6rpPNLsRUJNyO3r1X4A8OvHYCDQxib2ubNJwTevLbI+FeML/vuv
Xz9o2S5psUJuoidQ84SCk8HQ0LkxyzbyeUZMX4c/yhbSfAieryiGEFHFi2TvuyFO3NpL4rlrfmkC
6meQen9xFJ79RDuYpJSW4eOxWIczq+G7vJGytH9EAsNmmI61NFYm/h2blsaH5W3RDf63yXaJMW6X
mEEmzIB1OrO+BuATcuHOLNfllczJM0u42RVL70osJlYanUUl1fCGV5BKThdQ77FKRxDHBpVPy1In
K8NCD9p+cL+vo68Nlc3E7n2BgiuWxuIl7coRbhHfqdnHd5DZRUWXJkoFd79zO/FUq3BMnxWs1Sxs
oILExaPiTAUSFskTrmRh4Rglh0/XEsW0RPRWo4gaJvoaLQOfE4nvhEXUzgM/AB1HPx0HNjzj7l8F
qvb2xjtkhMV488NBiQLlqQfuMoY3lcC6nJoHRf2/tJnD2pnK/mmB+Jgcru0+U2Qtf7DDfFyC4khX
mwTTE7EhbpWRqc7OtIMgwpXzeSmp+eJQ1xb+qsN9w1lcVazO27LADGOwyIYMu2nEW3Q5zUvYo5/X
N0NVkYRbd7U++6QvCIJdAjbL3exEJEeSwz6Sva2TMLnb1pOdO2LKZzNxeo1t4mY579ijaIg7R7hi
Eo0lQRZpnxwgkxzl0wtdX2/YZJPJzFk1BZIRBGm3/id0kVc0JEHAd6+dqQFFuQ3JkBoUhukAhhHw
lg3YkizR+s/6rORKS6/OuJm41B+GI8rUS995lc5HgRWcZeX4/pJlpRgp9WWQaZ4a5Sq8XWRZsoU3
2DQSTb2HF/Vo+odthL+28nFaVcArnofH+eMShG089or3+okGFNI//sJZHn0jbiZQK8JVNzREti4/
ZBfFdHi0grnGCdLkXT3nOYYBdyC45ZTyGBdv0xDv+8zkmvspdDVeW7sRDjSMfzctCqSNmaDWMDVP
9nvCmEm8WONoX1XL22l4SR4MGrXj4lrGFF5dwV6rw849mLbO2P7VffHUE5BzRCzMuSb09t6N7bYa
a0Bu0vGeCTD2zuM0PU775rro5RvuUGRlSATlMl7cMCyIPxTk4DzsEvNUZ/PQ2G8aSe+VNHatZmhr
UBOCQY8cpgoGDCtCb0kcwUaq2tJdUUsPOxsMxTNkMhQYkHW1Qlz0GSNCIgMLckXG35WzZRLoMcvq
6N7dVxZ1k3EugZ2pi1bjuqivWcFJ0v5fuNHFxmFxiWWxE3KtKd2cdY73SCZ265OfUB7gezQwrl3i
YUFaIhyXWjnmn1/k28GThA0CkfXB2jYziZrECaMUxphA625dtJuGB3MPc+rBp8ZBc2krsqLqObzO
GHv3JNXtI12h1IYJfrtM561fIUMi+QU3N5QtGbFDRljT5k98qVr/Oqdeuynm3kxlnUFbgtNmHatF
mE/UJdKyfifxagiFoa98UEG3FTRldjw2E8wjlDgXLnxn2LAOjmhEgAkmEJsKxeJb7WUCVyz3zzPl
c+3aTr3XgnDCdi1ULjDC/WWjYk8xHVBtxJBQQAQ+ujpoPeosKxXYwI/Q14M42NlcyTMRJ9+UbpPs
+0cV6hvyP1VU/LdDCVqW+xEfn9XC9ZZ4DrTrcBsAXYpSObkCpPMymZoBrOx011fP+LFlV54qxdv4
3WfdARJlDZTIDvUIG4t0ajxLMhG8rnhrxbSYumEcViA0AjvOeaeeC/KyiaEsIEq07FYse4Lw89WH
8yH5ChOgEuQ1L/DuxbpMQ400Jj5avUg7B7MYdoIx0cMK2INSZiapV5M9JR6phVa1WpTBzntOWOea
g3D/LYrBO5tAwZXgmdCtvr+LIr20GH6jGTjAtocugDOu0SAeQc429sNIe7NJAYnWEZzTUEWewZQZ
rNUmO+X1uuKu3jxyEKyMLvC430BINdZKRl/MWWVW6tSqef+hPWo1sPsyGPyD37CAnj6K0I8fN+8r
mLsws+cp2z/tCcoXfF1IN/femu10At2WbepFkUyzDnf6OpIZfpswmxZxnIkDSvOcAfRJ41jDgyBQ
IDIk/klpODNwmjYC59GP4zd5qp+8qYA4MV2Q3abQDmK7TwhN4vfXR2vppqXp2L/sx2Pkh/GrsfbK
tnRQSfBbOXZvq6xXt2hLpOARmwabXxTitUagcWV05DQDerj5NbpmptR7ciHnzK6LfOz43mkH6Zhs
eJpSifZE8rtffX/LodzBVcekrAK6b6EE58mJ01yVry9KAejpLGiFO/I2ze6m4qnPbT+sQofAnyM+
XrwJ62s/e5aQiq9h4o3QNF2mvO4Yyo92/PTOGIOkxdHtzNUIw/FBmvKIk57SJ0HRJsr8BrrWmnnD
cUJ1vJi3XAc0/fxm/DmEcrreIePJjDMOofMrFEWPh7D55Ywfe1JupoD5gDJGv3qJvH6TBfS3blU1
i4Lyac0TWpG1qGYjPQkqfNlmqkaJ+AGhYVH5IcRhsojWbCDS3o73fw1e0eYeRtUv6wXO53DBjZlB
tEIrbVtooitVx86BEZ7Nf8+Cheh33TWqM88svTg1U3rbmPWTGjr0nu5MxJIAZVDv3lVwpFVkrGDD
O9MF4jKrtWv85wMAA5vDJexPhWXJCI5tTS/IfTSyhZ3uW7QITB0o0jyiylkKwhybDeT5hdGL3VjY
bX6tuEcAS31kvDCSYLDtsIohL7o4HGcQ7ffSf9jVl/RXXFX0rgkZnWKFTjVRAQGCMD97M84KamkR
nmF+p/fFTJ1mahRhCTDnYBjxA7Fh7Lb/rnOWxb2v8FDic3yY+vnmE724s1rt89OxHlM5MiG7kwQI
uLxAE4OuXzQAILNEedq5qQCVviX4e/qZSCyVZfbVcXK/p+I7sbAhhI/g6kbZ0qugLyX3SewnpIOt
K4bLMTIQdaDKtAy4ulqmwrZt8iWeJf/Znt3yH/fiRf8mVhfy+ws1ZrGapeUOA0i7EcISKiX5vYlC
t9i/EB5UVSoQKL0IDDRSrrwbUe7Cs/rUpSkdenUOSZ/OoQ6K8fxOO4kq+DvJAm64Kk/GxcSRDMyR
SANLxXrMLrajc0re9quvEvGEeht9w4V6jjkGnUEvE8AGBZTeysnvl3Cam00/5QjKJmYqQUNcsrsa
YfxnVGU0vjSgaDW8/g4O+VLvSrMKiqtwsFgGfmehMSZiHbyTlxr/VUlsq8dWWB2RoRc/lpGKU6WQ
DWPTcfI3oQwGLELuX0Qu1V73NPh+IkGEtI+FxKht9Pqh2BTL8CpYxFRKZSKznQ8qmUi3xDc3QNKK
D8u1aUEbrUvwJmZ0OGEoOFpu69gUSgLU+Dh1+vETfzrMRDI8mMTj/SAUcGZdDcPwJxrhYatAzvQ+
d9S/kUKXx1Ux+dvA0j2Pbsor65n7fV8oD04F2RPiPw89fuVqNfiQdJZ+j5GhX+H5M09JWrNkpUuS
qUKOPyTJmNckjbsODMC6P+ALvQcgjzQBkqau3Rc3DpSj2XtfQ9AymWGVre/9uxje9WWs3nUmLhqT
9BaQVwGA3+ooQKjTioVyZxRSqT8xuFJSqz0fNR/oHLYSspxwJjrPUWUe929bZokserx/i+Q2uqZk
Zt6XV/RZBiIBl8kq6ABpbJpTPww3nv83pM31b7QRCg1YCISvt+b1lt/TTZ8lBz84eQGgeZiCtJAM
5088/jXFwGQNH3/0PBfSGCeOHhLMgNf4Y+i10t4Cp4judmRFw1Ce4iS0DNWXZzGRbeBlokgZLpki
PB0Dsa0CpRyz6899MXZczPMCwD2sJkDBb2d/vGHnupOkIk4ZM3yqFWve+1bAnX22T8RQb1D+gG1p
GtAQVucyg0+bMNdVILP6UL9i7ak9znpHGtN8QaV3xGg+imCA2BV0Rgu/DoG76E5cokcN03HoyRGj
KjzuW/MFrnTAT97XMtv8M83dNhUgFuOlrRCIQF/Y6qYtgcgTvI35N34vZcVDvXtwAxqRXcR4/46Y
5nCbgpazH9DXkMF87WTTMP8BC7jwCL8V4RyHWReHrEpsu/XHmIGdUQb63exF/KAQEFQlurTytVV0
z4qI3ZYXMpfIYcTKDddMfDMGJcjjpimIlFZpTQqdGZbczfl93Cqe2fbxH0Yws7QfnZY1nS1o7oLK
Ve6QTb5d05L1/QK+BC4yvE7XuAryPNPP/Gg9WQXUlpQp4CSAZScEqSPaY7wsOHQAybfrrg2QZ8TL
s03hnKsONtmbDGQT5gpr3OTVybdErnwlrCFPK7GR0y5e4tkjo81SPR1PKocJDsKnH5rvKx42fAZ4
pArUgQnmqzV46lyA87MqSn7S1OCos09puumBSAMR+fcSG45nS7A+G41fByCMjBd3n6GHLkQcRxP1
5Pyy0BO4QfqZq7uXUh/XgaAFbWv1x5jqaHjfBsQVsbXR+tG+xUnYPQvtLQfUxo+y9uUgOVRsXh/C
W3R5mkFlQxyDFAL/g7/ak0oZ/l86kZ0ieGSBdqnffUzziKU0sYliTZXoOGjshOG5sOI8ZOWV6RLN
4/jXh05mDccL/KIa96FB4GWva8c1HL0f1J6qeTEhNvD2oXbkr6AaBkp1ZkgaWTrp+l2E3th5Omr2
BaQVutta7dkKRI1+7jUYfEBvGHkN64geStpEzaf9J2L6WZjQ0r2INEhYDGk3seWzIPtRwRGTU6am
IADW5FwGDk1qRJbplBcnEMYILgOk9yNbpp6EZEvLCZ0NRKiMkaSszmedtMvHFZQsUexm4WUwILo2
7OXQb6wm87yEg4E/B3LTlBI89M3NMDz27tA0rT61CFOvWGzhoOR0tmgF/s+zIkyVE028z7aH/HPe
hOeT01+PWIeZoEZ8DyA43NXvDT3lq8kDMwRoNVbXdbk1RL+0RBR2G+efPJ3lgUY+xkSzHoJ7Qb5g
+XZ3HaIy4JQ0QxV1DBgYaHu5MtbZZ/AnO1tcqhaZsy5QnSAs7DOVNZTDYndnGtkcIQ5SI3LHMrBC
vOBbhApRDDBO7CYakWEeN9Av1Mp3B4dB1Yqb7JP27BHa3juWrSokE1MXX9sH7Lqq7dRkfWiFm8EP
MeiNQcKCUu/7TOXLQehgv08ZVD0GGyCKLt+thR4JBHSaJLiXDsfsJqPFCxhRXPsE5AQs0mDoY2j1
W1l/3otdqFKmn1y7KEHjvswk5W1awScs3OfGe2+/sZhiaAcT/OQ/2xyDEa92EP+EanSE+vA56DpK
siPVPIxtd+XDgqHMojqSl/KvqTxQBmCJTg6JWPZ32YUx63Sm977lggEMfXl1Cg5A/x9MXdD4AX+E
n3YWzBLO077E59qP888vt1igZFP6ARU6wKIaXXYWt3bndj0heSMxwGVFu3LNSKPt4l+y7UU/3T31
wZHQwH7M17LwE+3Ehyj03j0iillQSfSYJ+es3dJk3vR39ju0P3V18yKCUDTpYTXk9o9PvJ+64sVZ
CpeJc6U9Y86b4PUPunOfA1m2iDLKpzBTf3jO3pxmpbQS90oc2jwQxspbFmm1pBioH2AXUqfKm+MO
ba0TsxkqpG2yI3Hy21lLP5fG45+8IRxxclS5ckvMZMBstxFQmjN/Ms2SsZjK4PKqJtlDQX/fpoX3
kPJhiG3T2ayTky5+6JD9V+objUruhcuE2fSs62LTtgFHBBIeJWEwfKNfFM32z7WfaMcPFN2j5YiS
ahwC2ZPSJUJYI9xQcWKPOEClhUwP2K3ycRFdUKp9MgucHNWen0MRLb0UxlX0jzMK1AVw4UVA0KoO
deU+63D+4gXtNpwDHJfQMB/d5Hl1/cOh0PTXA3R+5XC6rJARIvcvdFZ3A5vt5978P+yNmVlBJBgr
ARnXwKAB/rsWUE4qQTZnKqjuRRqvTOygvEFFCVQ6aHUvuSnSlDI1IZNW+Cn0crc3eWEXd/I66MLs
9F1DnGaaEjup64MhzF2MEU6THRnAadoS5JMz5Xc0VyWrx8hgULMjLH9v77CViBGpO2qkr/U8ZauZ
d8pMJA720s7NjZH9RB/15KkvmEOUcpiu+bUzK5SJZJhCoVqJL4B/cPOiOtC9Yh/39d8jB5KRcccR
QWqMduJOsgNwBd+dMQzshd50ZllISNyti8IxEth0xRJF3X13j6f3q1aY3kD/QIcizFD6VbjbBPnw
MkJM40NP5xu4P5AsP/XEJzsld1J9NBFfdYUkdu09s0x+f+j33gkWChntGk8xczYa5j+7qtTounFc
SgDwrKL9NuFYyLYBjfqmliy91Urg6P2KVF76BoTNEuq2okfLzxhwg+UQUiSnod9QpR29IhPNzXDl
zbb5H96/XmKyiYSPgas+pZ9Q57KRjai4uNUsabFGvgd0gWuYZGNGEi+grRwfo32awwgK4P6y0hFD
WuQleP0txs5BuQr1Bt4fMiK2DCEokwgS8IWp/TwX+tQD0ryBjuBgO/DEsoP8+7+W0U0p5cPwuC4J
pazp/hJRMdxos2PFI9xYOR+8sDHdZkq/ix9VtviQGF6g7ehRIrDaKDahINd8o25XcSYSVchIBN/P
tbJAGddsE2XS4dN8I40nfd5n0UT/F44hI2kCfG0kv1NFI1qwtBKVMp97BQJakmJOILpwxf1bhKTp
Ub+QOjwpsb+KNcnuW1IOgw4F3rTAroWhUscosXglgenL6WtLdn1fqnq/FSih3TBqRdqJV+CjO1BU
jpD3+gZMmHA4Rh0yFLvK3xyOS8AIVKYNxo5mg5C1glP1uy4u4FZIKR94ORB5X1Q2sX0V4wKhPzSS
fhZigHh6R+t9WlO7YVk/7hjEzzCFp3YK/uorJDFRkN7Xo59kEi5zFDowQaQVfi0zoMXHahXo+t7L
IXC9G54gkHvD7HKemxRUmQIf+HYOjuwzyG3j5YllOt2IrKcoNU2Dm/pyPOt8Mg7D/39QS+vmYFMh
fhzCZhOa3lyOpkZwptpAIf3Lh29y3VxT2MEBKAqJiZQ8f53yygYYCIvuscxKSLyj1NylLmDKJDau
zY0UTZobI0cKlLbLrrPko0xPNVAcj6cMqjSDzqydep7n8p3Lyyti0tbjGexdouzSKAIKT5lUebTE
PRkQQ7mJ/al7sv2v+YoIGmOGmoHTDVZioIlOOfDGM05yqibZuj+OS9KEolL50ojamD4Y7oAGO47Q
TVXtUXuLNd4D0Bt59A+/g8pIinw5kyX9MRckgh7lxMp5lkUTeyfm7vZqq3BeBekqFI7ybfi6SBGe
ehr3oQgy3I8optJwrdss26T/pSq8w75O0JVJJUkBBHjglSt75SnwTTLExJ6PYoRYevgvTjOwxiJY
A8WaWTjFSLF5SjXhBy2N+oQE/IGgDpAE86vInEMCyZFCW+wnyrJf911GQgjRifI64P2Lf2WBk9gY
UJ7q8kCqLCW3yoGobT2NbMWBKT9TUnThvts3LViEKU5ngIrZo89ne46pkFN5zX6hF55xofBL+cT6
+CvVg2wv45+jSELmPUl9dmdCdP/7E8jveQBYvsOl6prG8NS4qvIn4Mn6Bz8O5NKwLOc67gkunTDe
prknLQ7ArUgt/GSPMzZQZQey3kL3K8x6nNk75YkePo84ht+iDlzNqvy6h4IpdlEkMkERBIJdaeFk
dzkedZ5dzaBmJgvUN5AcAV+eiGnvXKgST0dEk/Z+85vkGJWtM7im+Bp6TGGKouzlRi4DFQVCXHG1
PF3S72nwHHl4WskpTcmfr5S6pyndNh/9nlugYFWzI85fZw43AkEDRKVRxxTcSdIp6Jev9CWy6HNM
tx95N/wRb0s8Qrd9GMOn0JQG5BodtjWTWtR1xSwlRqlHHJJYl/7wuyp6ghM1CytPcziLwjZwTHxu
p4YyerJ1TfQKr+R9OCyGESaXZmnVodH4SzNlO9K/EOekwfv092DIaFDhIqqsGynlPeACmtrKWKkQ
z1GCkR8XYQWcqjpuzJ2YdKo6ocUlrr2oGINhpaKQ+5C5CRt9QxZmrTrhh6c+NSL5/fnjaE/RM4Om
rK1/51qfTHlxm0bIPfuIcA5cIh0uM6tTsDFoxipbwPSSqOpDIMSfHbonjr1879qc1VZzaK+CWslK
JhXf3ETJ32troO9elGgthK0oApVC2vxZEsDRzoQCdRdGK9wgjskIZvMYx6vK7CdseL2YWW4XNMBQ
sBJ1dIr+6XFPc8uhqPrsnfVq3oCuUvWHyFQ/czoAOibAvybyzqgej0YCmJCo5gIxkiHmbkAYzqfu
ENNwL9ItYOoFDDPiZth2ovOulNgFbIZ7pLr9qlVowNi+PoM4i03cF3EwHzh4G1yuM/2BcQh7/J/Z
gOazh8S58Al3M4XTifnxiOhxg+jb4PrlutCLVnM41BcodJIBRY6gqxnFAdcNS8crWxjnD+Cn+m2g
zCsKdUq1JdhHvRF9YE7T9666BVRUknM8+Dskxh2eVmfjQ/x4wRRuP0+9/2fdHXdG9EbS+nhAb7H2
6y3hU6qfnScN5z7l45Duz7jevZnVkj1JJjD3Jkp3IhGX7rAkt0zjvGU0sdx59yx1gmSttHOVXsU1
ezSssLRrp8oewFOahoL6LN+2HTaoB0cl0R8NqobWA9nsFLm82Qme3kdPomsXDBZywQm5MK1vzFpc
TKTEQ3+XH8TleiLBTUgVk8Cgq4jjL1srdUUgY2X5XkXCaeMTEWg0SgYILO/0/NHhNU1Myusw0o81
YMylU8+T9JJp0LxMKSkJztS6b6KVwKl6NsskM83MqeVjUaPtI4boyEB2y9TvT7k8QyJn9ba+xQW0
tx9VFtqoRm8p2Htr0+1CYnKsRu9+b41xygHcrLTpcFWkQicZB72znLHPC/mDnNTWqPrzA+TtFBoU
Z3M0n1Hj4vc4dMl7BMDj4ZPivbKJKBpKaaTGPjQimINaqn2kPWC7T4BJMs9Xi07ekl8upCwWUTS4
mDOF/Jj5MDZ5oW+T6KctkeY/K2G9nT1FV26Mg39iZexa2+ZbDySv4ROsC/p6JbNEbhaQJ62U7RoQ
+lgUayw+SR5W+guUVho6q/nNtQQQHpuycqcyXLxXwZrAfJO0cdA8A25kzxtjXPwIp/nf0w4iSzJU
MSuArbSBTS0n5vIZLPLJzLyQiidfncAQlx7Kxa8jXHgDiQUyJ+fqep6XaMbXolcXRI6VunKtA6En
kHt8m9QlgtLk/+30oUJBenXVyZz41QkhBpL3+6yBcb2AgRDt7q6gL0NV51DXaJBThqfg/JS41Kd9
HJ/ygziwllnafK2d08zDndQM8B4+JHLCcHHz/dNLm5aJJSID8HJk9m9Agz7dF1OCUapV0CvhD4Fo
2eahQkI00WAS1ZPq+pr8J3JX2zsH9mO0/Mjv20O17XrexYBn77S0clpQp5Fg0J8E3OXzMdJn57tZ
mwDGB5+d128yzaX/9OtuKrWIbyElzy5Nsu0gBnJrOUnBhyHBHjwMBeTJTbtnXZzgcJeQitrkn3RC
03LH2Qt4IT1yxh9hJy8GQcfw8iok1aWjvzp43EDWVnlGioo189V8o+asJ9DqePtOabyp0kNOQsdj
rlV3AwCr6kwebZvqTbpkUYEoXOxjB0nOLbseh8a/1z/ezISMg6gEdynF4bVP1/sCz88dV8RiBV+Q
32v2ZAxniCxdgef2kF8SxtEFih8hElVU1mWxSsUUFq5/K58m2ll52o+d/ucvEWgEOsTaNKaw3YNw
VuT1TvezI2VLDIZOFJOKfPalo7F5Wv7DX8EmCbS9g2PzmAC4FNNB4kUas61nNNfHelxcsNq45J0Z
T5piEXZI/cDQ/LSvucCcjeP0iiMketbwSNaLg/E06CPArE2G76kvqRu5B+fOU11qYhHE6U2MkxKb
cvrWaeIiyZC9oOn+vQwVQKyvHs9oFveVOLntepYoGKSnugnEIvwdsakLWMpRfTzt4klUUB2qNcHY
XV6e1KvgGpX9CxT5MB8yRN6asYD3BxRBJtUXvHRrlL1axkWRQqPGTcT/gD1ogkwQ+6S90OwEFRa2
FYCM+w3IHWI0RzZ7AeQy7pKihE2xFyOARjpo3oIgodI1HTZPVwJ41lEYbnk+vZYeKzMKlKDWeCOo
CuZkJE9pRLsOthYuZAasJlcrLxubWBEG0Dwac2yXHTRuM7aOLBE41gs4LjQn3jMB5769SBJJi/IB
MGdDf3NJ/w9Qhr3VPiETdRH96xsPYYC4DKx8XdlluMF0CFzoxUrZ4o1PhdguP7qCzq7WsgPiwz6Z
a2dRxHcyJW79Yw/hUmItyRTgtk3qPAhjRTRDPI8I764M/NKMRW0424mJQOCC4AolkfHCkP+QFKAI
RzyDpvpC1wZM6P1b+hlvSMf8R1AlMA1HbSGWRjoYec+D4p2/C33qyCL9ukUvJCWMACwoK6mwjyl1
fOYSferkHoiec91y6sZq1kuYVXmOVodnY0mGvYnAQu6UTdbYd8cGGRyfG78nwRk+hmvmmTWmbc93
ch5LZy/W+K0HI5vEMMdDKXhNXeR4NhATsVvSMqFGPAMzJF+QgI2rpDECrTf6m6LRP+Hvc06cTlvt
7TEyezjpQrz7Os9uGoyjpzy9PGGEt1JQ2FwvqD9OwwXT2x0vsPlstKMDCCU8tKtXmXsWVJKBfx00
Tm/QH09u2i8WU8Ue5wSZdRQo0hObZhWhNc1Bz7mIn3/G9NiTfc8rRrBEY9QUK6PkKxGf6ZuBwVIX
tHCTDGvZLe/qUjaVSHf085DQ2aWB89gj2+X9FAQE/fJQpbS99YMuWsTL/Udq41V9EKLo1mHyvsYt
tZtoaYhhQuirSW2yVH1+P/VMb+/kE4I4n+VmKhu/OuQ/3/5gphz1CweAX4YXaoMkU2IPbMJR7Q/g
cpc9HD7ZBff1QqFZprS2MTGDzjPYEh4XxBoUNrzTT5hvGcocXo5drk9x0WNEyvNs3dIf27mbOCpq
MulSfS2VOQQRjqdkboprB7KqwDecQ36OeEOeFgl7KkXKu6yCOUWPw7BclBSO0O91uehXQ8fxodwm
XQvpoeeek+MEL4EulthoQQe2mC5oIA6w8mkf6fjMcS1G1AO1968fdFtB+6qLNWq/W8xHbwbi5bbL
4qFttNXrBzRTDTELtXkeYtI+6/DtoC/9W22jfY+vagpDGmXjk7jf/yUss4/y75FidNbRCevIkKLV
6JFHQy31EClIrNC/zr2Z+lFG6mMbkzm7/jHPVUkk/NfITDnA+70xpO2qiueB5Dvz671aPJ257Mlg
FSDQDM4ci1yKnt7y+JN09AJknT7N3s/BvAZ/HxiPrA6tJkIb/Fk3JDjG1/rFOWkWvOkwaIJZX4Eo
snYWKMC++6unwPPRmP1PMQlZC9ORftohZ1PSO+W9AqrJQuIl7RB+ZdIgcAHK8Zj3CXFv52sh9hds
ALAt0t1n6JAWQmXpFaJG5Sm7fLqvKUG+A+Ghzm7EbhP3lkhcJ28ZI0eEI0t3HwvPr580UoIrUvdI
ehip2J7mS66oju1fLQJZ9l/bmZQfsJUMmvYuw9IHmAEwMrW5H7L0CVfJVr39ruIZhBD1Ql3lwjDL
vblZqP0Frgdd+LJKqRhOV3XqqUCCh93ihB/PGBEPW2MLB+qGTUea2okoh5gLDC4ZF3Oh11SKnHqM
pMhDZTEhfRT90Trd0MC0yzytNlJzyNVN01P8R94Im/h6fSz5fs1kRqZ5nVSBIAVouJ4ShxMI3dTR
H6NH35V7GmtpSFTkrRE3z/VsL8IXzp2wJGZNPihq5VYFy5BfrwqtDjJtamRCVY6lJL0G7oPn8IE7
W7gWNRv9iM3C3UghzcqJsvyjC1CJW7PCOJI1Sxiyc8TVM1mZ/55W36UV0y2VHeTA/kyaMg7/6hCz
h+dtv4VXQ20gJIVoIkDfQi/7uHegbevVbiiEAIXglnqFNYUvbVXgyhalklUGwLsDkR0AqolN3Z97
9fpPolfN9O5qooTdXIOvL4RzEIlBQspDsNMUGvlljEMSZYqVDjKVJZp4ZezvMrryKPDCVlDC3FO5
pUXPupBTZeQK0KKZR7Aw1D3/b6pNVrJ1EI3UAquTI9psw0Yl1yhbYR+Fn+ZDB55pYU1jEDSMk/PG
pQHCn5UdOSM3IXSRJM63FzusZYWqAS17tfpa9krXg+co72T9F3WJqXn6NEfFtI1DfNl31uQ7ndpk
+CXwzuVNWKtpi4q0ECGCGoYgBT5Xi1+Sm9WCbuXtwLEDc9KsuDLa8TOwcUEggcWRmgjuI7ZAPcXD
miaPatsa4YZLtd6SKZb9vBnQWhlH404aX/yPtKcPUl4ZAcYoLuRDJxKOOtBZpoprlzDos1L9tzLX
AVj3eNoO7TZuKuPe9tstJc7pi5xYPFhwSa60jfYUCFQ2RBpkI+ei1OEaFdw3ff5CuzfgWpQOZmVI
Sf7Wq++Bn6ALvl1mn0kt740niWVewa/LQp61S+WTUs/fpRhuIgkpG6quI+tBqdu0OxWAh9hVx7Uw
BD0lFMMGg2OnUWk0KSgV7JVv1UHusGzn/ZZGmmXB4fk1T9yHJ835jjjS7Ccezz78JOoxCbt2qr9s
mn6vu+zMUpwXVLa194tHTPBhoUW9ChN9z2adr4aJwRvU0XCd5uQIvl8dksbtyd//EJYkH5P1eDw6
jpJqZle41HwY9V8BUmYNw2l7D4tNNEMLp+B2t1ohfasRSSlIJA+GNW/VqklXaI0rdQWsVmEp0ob2
CrbyspbewH88odA2w3CtytFuUXTXmguCl8jsk1zfpXNbRAE2B5G8P0cd1rgY0G+VJDwj3TA4tPIk
R636EqDtrTRBUc4if0PFKoe/JbNLuZcrM+h86bR6qEbX5tnBqOhFTfeA3yNNDtidgD9wBLewkCGp
xKIyMqAjZR4tEMUfS435lDsEjngdweusgxn1Z5bL1aJtC7w3798qa5l1mQ7ON9HGqdwzR6UVNxas
JmameyD9rYsmY2hZKIfvqg+bS0Mk9IHQCPpHxV6kxXEl6Z75kkM9ZHFIXBYnVhinutNKIqwPlfrT
xg7SN1lkD0rkNWrB6FMFOh/i0yEUMaYj+hn8IFbTmMB01lJHcu4L7wvFn7W7aVMeaoyuEVv3ajDl
ClKMkpg5rQOyulK/lPkgmHTA8rNNLPk8gcy5ZoUo90uBPRHhu7hn0VJtTjp1Xd9J+15Q7revsibV
p7w2/wWVTsbfaa2ishcPwdyBBjlhsxzgpDzMoIS8Mgu7fkPWb6q8xivjP++Euekn0x1ezJ7QqRFE
beX8nPOHEa0CqIQmPlf1+sz8C9XpbC9AGOwg16o7BO3XxMhQxCJqT/AFwogJwq7EUQe5+WF7xcYj
UbVPHV4RiNyOzhxAEc8IY/PyA3qGof3r/C7prtn2KY1OOxrtpWNqE/laiAC1h5X1e5f+mfb5slYG
ggBOoE4vBKjsY7Zp8B0mseoF3kJyBpeH1AXKHkpVsJXfgIsKQqDWU6omuhnYWdqRU1KAsYJsUty2
tDnljCnnZS4HOM89quSFSac4+D6DXF98H0yu3qge2lN6HQxaEgz1QXnDwEfU+b0BFqsfE/bFi3Id
QQkalV/Gx/Zs5DptT2AqRI2uvONZNsEQSDyoKtQ1kijMHW1a4HNMPhT0mZP7zp7divYb0AQZOavs
NHnieC0TuViiSz/I7Je5upBehOP0jBC2T5hJgU595b9T0GetwtsUMoYhUq2KiYK7UQE64YTJCi15
wgSJVgZ0FmacSXuXfutV6cTY3lunxxMaGnobQN1nGiY++5A9vgqfbmzovuQTgpACWVS2HibZjRAw
bOB5QZHg1YA+Bqx//vYCUeexg1mMF1Cx1afQfIqh1+288/xZ4dBUXsdfiCFbpdvR1eWxFlzLzXQ5
z+1VQqUdHk4u+El9KBKG4DsJAJ7FPnS3ITLlt21YWblxnczHGHoUJLzTT4fGpGB1F6kwT0L9uBap
0HqbLNqUHjgqXuWyhjf0xu09FEUV/Qv6Uu5DKYY/Ns+qiopKEy2NSXP4BopLj45uIas9sD1ZxU73
DbbZmYzj/i+IMa0l6UtHW2hX2HtKRIJIsuQbBrjbEoQZ+by/1CiT9MFUfsDMG2v2E4Z+FFXxf323
uZiSS/OulYGG3HwEIuuJTNh3ncFCbaN6GJvZz4fuWIyjTX/G3cARf/Y7p4bnfSrLLx9ytykQM23l
jttQdHqSLE+XUVygzamJijYGHqjGR+0h+F+RhgtwSkSviUJJNkFi4woO/uGM1YK68gP4SjP/dqaF
7EL4eStdub3RjQvIfkH1u0lbky+L8oZn8n9vaGbgqUoSqvQglO1K31FcfkBnJuFN58IJzl24ljWC
NlPVOzm41uqatGJ9TNusLFT761zUMVlIeZeTzs9/GN/dwMICv48c6Y8WfWCwpS7kQ/kuxrRt0fKK
1+F61sLsxbv7Zl6jtX5F118odEwboywrxkAzO2bHwPS0K3h4xXzyFjbzopZGqtXB1BOPVNIJYBTY
z4NoL6sdv4iVArKOabuqEVEyxt32BDoCUAmefyFnSDnWcRe+tmipwIoNecibHHkL27EbZmoFVqjm
RGWKqOLn9J1QLtf71xnHYKfBj4xm2hPW0j0UkgTcHta0b5QaBu3RbC/rL0Jb3Cc5I0uUuivfqm6p
2JvR8lbCZZH/Q0K4EPEdSFrXyWIsSYt7t69Fb/+wPrP5ozxsMZUr8coV2xwVCs+svGXoODYcFJLo
mA/lFGLRxSgYcUTkBarzIDVi4sQY44rh0QM4WFUd/d4PpaSWSIDd3JoFHsLgZdBSRt+/ziFevyxD
9RtM6oOz0/e3/8oLjLbyDQ/95nGlNsxV16Nv9yYHSVFVFpVdXrECkuZvMogVVDQcK+qu4pyU6/an
hRnIH+w22q9ydk+YjuJWUInLW6CrP3rXK2owO5e1UjkXLnq2AR1ViRfBwMc7cXs0/WR99AAYTYan
qUAHwJhjEZfSyG/3j2JZbr3qdqvBhsrLmCRi0+GHWJLrWv7Q70FLEtwCSPLEFDHMGCmncMrFNpq6
MtL3W0k2JZXq7KIqtIXVimWQIv0aRPx/9hzyuOnHZ48WH9cH1/PxjzNDSqkIFF4xvn4fn+58cHFY
JZwEqia5hBT9BOaZYJ3Sme2/0bgCLLJjnsKy14FO9SLwh/WAc3pvyFq2NkLp6zBhuKlQVEaDI/wK
Wiss3tCCzTs0NXKiyLRg7VbYy+pszKwto78mKbdxK/EeDZRxYUZW/zWN+PvwLJ6jzJbRJBqS/3AJ
vbKkXjrvWeDLK5lxi2biikKz+hlLT7kW1JFhCYu0qUG2wL6uLP+5s5Lx571WAilU8e2ab6/R6V8V
xBEGitCREXABgEZcCUYctWzU/baUbDA9npM/xdPCkxU/f4r9se9Cf3bqyzBBA2Wg1e01tYX87zW9
qTX7kuttrUQ6XyCIWRvsy+csRV5gJJif1CaxMB+u5Yi+NGQUI7ObGeZgUytXjADs69Y1Q2aCw5/z
QIvzSivGiQSduM07rYAl8WkQTtAUk9EifEXbvIxlMRn0CWWrkcmxk1+boonnETFSH9D7xbpcvL+h
TT/77NpI0irVD1P3sMFKrAw1Q6hvp/8LE4aL5ZBc56nfXPLrYfahncY9624PFC3bU4sGr/JeN14F
otKsxY8QXQOTdNDdINXZN9GqPjB3tuobusWUi9qurEMCGC2VlPhbdrbdmtSuLW8FPEGyrIy8dNpU
C+vj8iC8bLT3CDSo4j/fdwJ5ZDFGClnPrsqa4eh+37ESALRyEo5630bxgMPL6tC9DvTt5E0wgeYl
x2yKjXj07KQEDsMiXzilmoS7zogVlMKqE+hJkyWVFyIfkHW+2P8eMHwBvRbbEaK600yXxdRHp4W0
2o2LSVXj7VNkRMHPHxb8vvlEfLZsQOc+YR0KH1rbxvn/9TDcnyNDqLsOXd860xsMgesDeF0D/NbS
HCplF8T4zjTYeGWy/XT/qDO6x0s97/GGBkmf5EQgrUeDFs0um8upkrAsBPkKx2u2UVCoxNuTgND5
D1uiE1p2jpZd4dxrjNAMZ0vhEY07lmIqjAfezlYXY5toGVnqP4jywylz5abiWNdahQLjaA2kRHX9
Q8yKJfL4d7k77D2hyuBgf7V7J7QBN3gxEu9RXM0NdSrO7I7s95WM44yCCEIJ5RxhK3rGArm0EMXI
7sKMsF8won8o7WHjSy+//phGkXI3T58fWv6L0nP1uMUGrTCFtIaLw30HVVV+qEqkGohQAU05JheI
0Jx0s7IV3JSpVOeOqXPo5s9vs8fxoFKiwssQ619FqgYnAmzKbn0IL6Yk4rygi690RTVXeI4nmUOw
qVj66CMTazxkthblppDvVlmtcQxnMfIf/mGKloH1Ab2PtRP4f3fExHo8WG1qO/Ud55T1ebxjWNJX
2Nh64z+n93h+UgGGWue+rI+287NI25pmDvADbgPnIlXxNR7/bOkY3CeWiD2U2vpwx+OoQ0wwM2Wk
mtNqEOAD53N/3lqsCVo220YcKzoOZPaq/83rERtlRfznFjZNwtfBNPasdKuoWKgqHFg6YLVA6IM+
pTAsn9OROBS/+xqPAwx1dnoLiLgTNXzvX+q3K9iHwDOdBe4Szg+Kpv79dqBCvD6IEqFmH8dXVrnr
cbOU6Zl49lJnCpanrKcXndq5aoRiWqG0H1PhVU0xEDuIy1AKllnrilUvQCkq4Qzr3GHHuvIEv7ut
X3hb73NpB4zK9TZUAc/UOyoXFlgVJT2qnzPnuaTHAbJgL4NpKOAxMgeqJl/EH44uCSphbhm6jQRZ
rJxWjIAyMPS/vcvxiscifDWUfO8QrQ/NAQgpr7pjSuT7c4MNebR6JxTRloDI5N1DWm+rfjXDcVZN
C7EiNHbbSeygKiVkksjWwK9naRem38NaTmyM8BOGnD2YKdTfVLssJlGbqnqigeXQDiFg/UX2B59w
NjjlLSLPJFkT5RSE7ZNmlHTexJ8bA0ugRmMg2My5LYoEVW5wE8W0xQ6nPXkFzp4DNR7wdf0BW2IF
s7fzR0RxzZysT7oHe1qpzGgiZSdSBPYdPn8tT5yyEX2j535iwn/BBd8vmEMucgVI0Jhukjm6sUBl
icCVYj7lKVCSd2EUyi6KeKyRlhuXMIxhL13xFc+I+bh22rxlNIQg1g6iZxowRdoSJoQDSSg2k21k
badVzTAwGeE+NRmW16JT2ztLmDXJDuWYjPcZgOOiTaJWVZCugkclSkkpZxJ0utw2FnEE8NdIlDJh
zSTZwF/fWsD3zhJ5985NDMG+1QbYj5d9K18SqwgdY+yE6MNCasRwIinxCvejGAyb6mV8KsPrupto
nqg+ns8YPI2xhLZ+2GsO4JID98Uj6RVSeiW3f5DAiFBO70L+/d9Job1l2alX0IC6dw/0dJe0b7lv
3ySN0u99x6jLc+u/BrAl3HjdfQbr7J6n/NtR51nH3eYFTEME3E+ArewNm38g0IpQnEmyo+/zhViM
oKYo0kHFWcB1xNBE5zcxPKmF2nerfWy+Q6/hniPuwyHqTSALkOqqzlCEVkVApOtsCjDrmLWyPFND
pz6ADmCNaSZdfnVjJt5bDv7QrLu08v2fWDg7146H9gDloKyIsahRdRJDyAur35LqQgc4Mx+j+idT
XFd8UrSA7BjYqGgjpyU3T1IDrE71nHC4zNGUJPPdXKD6lLudjY/Vq1yJEIliys938gOggmDp97nC
NwRT+QTMC2ciToxNLSQWw/mCYgPp/RqDAqYR7R0R635qufqpNFsLwilcz2VE/ot/ITKcKfnV3hWU
tR4RU0xxfr+uD6B5CfVFVpOTUuZBhLbrd89K0aQmVloNOV1x5eZvR/GZ9UrKezCut9yZFmfQRdem
bn1F6Vf8ZB7VFyjLXLcgA3LbiT9yXgngKdkgEpiX7fQsDoljiErY1wXK3VOFZPwr+HAImsyGBZqU
7km/kzxxCXI4dNIvd0BPUTuiWTzkeLkO2VkC0faDB3/XjmWGVEQgIyBPzhsDP+2U4EjtHScHDjeW
KuwgDIm03F8vPWs4J49rdvCWY1dBMdyXPw/92CtLfEJNzTIV2/76EM3vSIuvIc1SctXqTFrJ+1j2
H6WFuOmEhFjipAz3FOUG2vEJc0/xdVUgcUF0wRk4LzrWPecFEWk5qFLsAQ44iNYiZNeR8Oa4mEXx
ygYVbXYP4CIGbPWRpzwAYBytN5ThP5LYks/t66S/HYQFHU8mOyMOsoxRRCcLzY5zfb+HmhRyJF8k
7VREP9jquEPiW9J4viW5sQUFnWlucr9AgcadmZIPM4EdoS1cTnfzoAZ5g3LG7qfREj8LszMcu1bm
zwL9QhYQHrFXixYwHf7fKpFUEzwV2rS7gALdWVlXtuBCePSRq6utoxedRnMD6wRZJ74xrs12+Jcp
B49Qx0dMYBvF8uZhCKbSyO+mvKLIad8vv3arhxBCE64l2GNHnZn3QPv4U+LEnv9ROTV9RlKwRjGW
96mXmmE6Ipjbt175Rum9tNUzqqxA+B9G+QqzxpfoJ9Xvclyy9D5K7B3T4Dbys0+Fdt9eI90jVIZV
jjOuRxK35A5zIKs4wftp905XxkZY6X2B7kpq8z8zI8OEA2+zuD4o+vRbdyjYv2PwXW6uqmaQ5424
C3Y2DuvMKXptWtzKTaNjNA83WUcDwK+bUBXeT0aVZGu1Z8bHfWxyvDTcbgCZ0IqZjVjeLSlFYGA9
E6gLtabD97RCxhnelnmqP1zD2yilRttAo2LleRTRulOV59dZ3iXeK0p51mJe+UduPcZxehX/nchd
aiL916mXykEmw4Jw5SvH0OveWVAclzAaNj1k8y0RuLTX+KB40QYggQT7l28klq+9OTr3SFZBHOda
gy5QULAaXFPg72X6ShFN8zDExYhL36DIe4LJWkhYyrSmb6Xs0yOWgFkRaSisitgri5IOEicH6xt7
UD2D5EObmfLZSw9kj/lGNes+xGwi/SmtO3VjFCI8ZM+eW1wOIJBDZySrGjQOgtK2zY7WLSXG5OmK
sK4QGKDoswm5ajLWrAWsp6MCvuwu+1kMjIwhI+nuzm8ZlImualOgzBvFy71WfwrGKrve/g4UqBjJ
pY9Kct3VJcryno7mp/2KymR5IajLWPIaUw7CSlwhb3nQ49u3l0FOUyltTiRnm/vx2gFL/DSYTP1G
0xGCeiAlwMJo/q9ErMYsFBpkAiFzwlr+QF1B8NPcYYTiRwtLZn/AgFaJ83o61ZpliSo+5BbLCu5o
Pm3aXFjCetoDLOXM4Sqhzvm61Un1yvm2rNFstW3H2vR7XevR9nMqUXEditBswt7AvON31S459QPe
80VBGYkgAUoc4V/iPPip9gBwRCx6C4n39sM0TUSCJLY2sSaG0ccRk4Ldeyx4VcEyb0LQXMVNE3HA
Wy8rompZ87yMh0rkBIuQ49UcEQPq9FRB4oKrrZgDb+bEf7nWyoGZxhUvYSFCPkljYNJtp9F34hWY
eSMIwHgB+p90JVa/CrIyFvYMXgndbMXLDf+fNx1z/Gl0m3R++h+UckeFsoeKc2O/Vj9BbfwRX/Gu
dXG7TfZsY7779FGGe91losMEBBDTc8FZ3ZFawiNQ2y7lRmRLUh48+bqtHIgm8Pm7rOAnGha46O2k
UEyYYs8IOvTOh5Y4c+qy6X3yBuQKG2afbXCWXqAP390UrhKB+4j6pyQlinV2+f9nq645xwvBIYpH
u9AiSJMrA+GgeIEnSj1fOo123O5WBWpsRYTKwZp2LbXO0Ge8LFIfn3VQKbNhKBpo91In2lLf+pqK
Zp+gjpTobhFAC5RxQXeN6Ly+c/wpdL2hvpxLY1gHQiL2DFqdO9MxKroI3CvDCfNhSHUJLj3lRN8p
CzF87ZhVDOL+K0lQsFXXbw9TmU/4YXuNC4aRD8IfjuXlBq3eSZYcSgHRp1oQIHceornn1ClxIYLg
34XZdDN89GTfnHfGhCnqFMSXCLZf8JrZaz7fHAP7BVo6U1d7M9oRvPldOvZs7rpMnbd0syzR9Ei5
1wTnbNVWBwnGnN2KcRt0Nr2KB/GWYJ2dWV8U/pcw317Utd99VaBHNCnuyq1nDsyTF07CrFxDwwE3
iv4tL/0p0WqyVyJyqmdYeR5OLW65Bg4FsUopcs9PwhacB1EvXgNQgvddEW8aUplkF9Qd7xk6MrS2
hDw/h4z85XAbMCLchXzXEOh1ls9U2RXNBJ5lpUecwTiPIp5rtk7bhOb2B9BE8LmIdQtka69Hrs7D
aQm57fbWOMvwoGkkLEr3L7UbknGjet8dXAJO5E8KNF2U3w5WBLju0tb4fl8Q3iR/dsXXg9x5DRZs
EQTQSgDjYHbMbdtk6NpME3TIEg54wIZrwAcXK9KlkKEJUobGhJFx2ndp7oDsXNuMbIgI+8Kg6rH6
73TyKu32QqeEagkbWneOf3xBInduUNLy/poiztziNjgmmyFRQKm46+CeztdCc08fUhQT0qzKwKwx
juUvjkM5ucQxGr9rKBMxj0XJ/7nKJN4kVG4BMOPfzKaW4VKjAQ1F6lwNpxC4cZRu4+4IJ+s0jUXV
qiZZtLb80lA06Ad15E3oyn8ucTWPFrfoZVFCs+El0P4yoiF1Inw+4txz1mpgjQ6alcoQrje71RY1
r11af/7hqE96xKp8LmujiFUc4AaKj5ddpLflb1OL1DkOd75yjm+Rmk41/lQdwHaJoGXsLriLumU9
q+OCEmioYwN5Qaj69lgceWBqqvWy619zWcTGzKMT/lrR+D2l+RxaM166ZKqp83ztO+HaKUAUepk3
hRi4nO3NR79tIEpONjiR0dugq8H5Qx17PAAuEYUvugqbQoSMQ99lgjIZXaWw0q286cCH5Oj4HyMh
wY9SgkMma+W79AD7pLAUgMdhYMQ9zLr6H2JXDenMmP7qVNRlH1+ks62bOnbmsa8r6liQoe6hWjH7
+NRrykkKEcyINcxytk7hWWEh0Vw5ZQk23UFGRMfJ7ZCRQxe9HnN2L7i1GUCCTgpFysQXLWk6Y/TS
I+6yqd6u1ddI1+DVOUgHgqSlkAaBzTewiiYopQPowiZ5QueFxykk7rt8NAEenuTwoCQ/Pa9WAQNU
KwB7he640MX06Cick4UGsK/9GDFkFmPrsy7DmpFFs1Ow08nOE/IYjadFzp81boyurxmr7+Cj43tG
1m0CdJP/46A9XfFkai8Zp7Xrd80lglpAsZMc+9NJAZuMXJb4f8cD+ZS+HZmaqwyuWT855+Z0etVR
dIUlq1Q6txS2BarKH1roUP8RHdNudO0MHiMU28NWIJ8SZBahH5bvF1mGsid2mq/GvKK3BavWwkFS
48k6T7rTpeAsO5NAdWgQcwpIdEuXFjpVyPMR7LITGph3oGsIYB53rSNkqeRBIIPmjPZ3tSiyfhrJ
GH3HwbnZyABoruZtOF6S1njuH5uo8gMObnRLUPzT3f47p99kGR09/DKtqk43wu+2YEb7lMCkfbuA
dAAs69ZcgV5Qq3gEAL1zfyP10OEKxwBT9U1HhcSiSS8lOanHfgYrVN2CdldkQ+FVFh2fciezuhTz
GvusEfU2LP7S0kdVYoB/+VBflzDvuA2VRvHAYGf0NVg/tPukSAr1Yumz0LMGBtZwH4kFrjEZrGQ0
kF8ftOeTPwTDnpOnIp+iJkFPRcrRCVs8hl6FpPlaao6IGMxpD/qU9PpaQyNp8litGHC/Bx2i4s1P
aspxxzhIziiimjFpurO7reh9HQz9IrKjBP/t/JGzQq4l829AGl7trVkDd0tUy7VRx6Uhzf2c2etR
A2SVQ6/UXo+9RLuWEKX3xjbzQMi76dEeTlFyAtKLMjYQwR0iyEkspQZG/m9Cetx3u/EAsD9u2uY2
AuE1Bhj43GWqJ30bX7KPFx8dfFYUWioHLtuidRtGseHUz8YKesf/mGh+UEFCbdx7gyxHX/EujhZP
7A26vRD4KPKyUdsaT7DbqCHewd0MqPV04AnflR2sQZB/XEXGIW2VHKZsd5mFieXBrryC2vgGtfGd
gRfPx/pbmgS0+fPeShIY4GCkDTuq3bFnybArPhNLhFm8CemuGa5flYTTQVWzV2Vw7Ljsm2uyN/fv
BJ4upF9UkwvU+awculDPW0/FuYNUk2YflBzroKTYeUz1k67d8+6WUNhtyTfjv8kNXLsHEp9Czrl2
THup0aGci10X4Y8puQZYIDCD3pBION2OQBoZL5HDdKLAuZNNBZQkSwvabHG9TqVEBHozC1b+V0ki
MPe87GVuxqltdb9lklISyVuqgEXTGpANuEe+Y2pA1TyIOZn77xa0pGrqpklCE0FXpJLprLLM/ciU
aPG29/UXTxETk+fOxiumBBTm87ZtYq5XIZAY//q1HWHDDqgJ2iioXwH99PJVVHD7H3pLVrt8ZMoG
J92xW2lkYRGTUhpCvEDAfrB5013XEqwHVxOZYpdIy9tlRXSh4llU/HQn8ozr9mYuFFaux3Q4xZxf
5QfgQySiLJ4Q28P6Yf8c+KnBhYfTo5hpdrv3rpbiaj3YvDryYoY1RoAIgM6yMkkldUopS+1qEVbD
djkQRWO0YNuBFvdBDQn248Hig6g08XTHw44/J/JZqVCf+MxVbTRP8UXSxWFtLgNgtT26ShqOqbwj
C9q7zG7cwfFOZKLyzWPrGU0FJblcMBsewpoyofsCFsZ1dIp+asRyjJOp+13r85qpVyz0p//v45Zh
z6dQMwDPYfRO5thonfDjQtYKLh9RfMFDfMgfGWz5TBzNvPnonlhgAO3vYZaJ19KVYR3robk38wOb
nYQXDGaS49qAvmiE839eGTwNJoZUVidmV9EGHxVmMhQ3Oo20KuVxf/BE+ERRJrG6sYRsyHGGJI+s
rvy/YZGxqD8U2WYxfWnvHnxZzYRt1CgFjyrY2FVU1+iKlYMoICy5vYXFiT81BuGqdBX7v7xLwqBZ
FD0EEtSsq85nwI+ofGCw3IWpgl0BZD/U3q6+lz34/t5LeVLLfOj2fiHOkTTzevFmPtAnzX7KfCWD
aooeNjnSoV+P1qp0/MXP/qWBS0V6OSshm5pJQotehbMqqHNMY+VMj/A1ThC48+SGBGuYObyEiPwB
sJIDT1iCpeoPE51pcnxlpohhcH3vIsxXu6yPhTasWzSikbi1/2SJ9KOhGrgLfMhTcEU04JuWe6/O
Dk4TDf9o6B4CNdbzoKg4UBqZFA9KnFeQ3k0GfpSbemN47sumWbBbUta32AmYQrxDOhtVcCAmaLWe
nfAe7gjJ5eoDJwKqDQX914zcwx02iFm8cIZQdqcZ/wgxz5ETWNBercZg56QPbUaKRPunHV4qQ25E
tx4bsxm12fxcXdWzTwy18Gd0ty6b7T+K0/j40fL7d/6CTdD35JPdfoO1jday6lOWrSWXoUcQ/baV
kx+egKn+KA/yhMGmJ3preWW8ijGa8QqbpSvrZ7/Isojvjp1XQpdBKpK2QMrdT8mMuLUNTIE3QcSU
vw6fJ95PonR8Ye0uvq+eUdvLRAiQN2vm44UpJChx47ecdWL9T4ZmfoHM9YXoOx/RpzeRA4PtdpOc
n1XJXIhegcPMjFQVKIiE0P+rsokRUA3j609FG65YqUHrZM8BRZUhPScZ8nje0uwh9AF0Eyej6WRw
iOmChEh9+fkwoHmcGwOeXjbe6avF59Hob5s97PVCOv7IYtelIwinVpyb21ZA4Jn22XFF4sWLzr4d
CzR4SisdglxkT7MPVjDN/6PdCVbCQrCZ+JooUgPphnj60X+AdrfWKF7+ehjK5DOKz4ovOVm6W7E9
0nImvdWsty9hJ+ivzFV9Zpd0C9QUSArlZh0rofe9lp1vP0Dz/Jyehs12Owkuh3q0rwyAsUu48yCn
QXlyxKZA6unTRw8HqIDnoM1Osxy8yJXh8mT3EALQr+fCmph8HcWDp/TXzPcLuYLEU4UUqD0H5zMR
duPHNL55Bz544D5ihA7Jh+5Oa+SNxuBSaIB6M1HJpvvOtg0BfdVBZXKeR9bsud4y+zHPOWIZf6s8
4rDq0cTKzKf5aRsn9yBAPEn1TYuTCQaN+GwIzh5tU74nI/8bxO7rjBZH+q1BIz+kN8ctDTJIRw6b
ebG/qMoGMO2OqY86ecbdo9/2LMRmE6SfiVjFSrem5OYQv6CGQoH1nG3Sni42QItuk1SDZCou6LQD
TtPTqASPl3SkDFgJYkuoS/qv/c8ftlEQuEILRWiMFyyPHNGAYkrz9RgUFumg8M7bZFcAg9SN++3p
5POdY4P2Nllg6z+5inM3r5+fEpyYLSSvth2foMz/5ngcVL0lsgBjGvtMuLhHXP5VUjWkMeFlFYKB
wjiGYHEbrtXjdum2tYgIA40aw2+8M1lNMce5xL7ewYBQxd+mLSLJtz54vFMBTnaxh5BJbrIsjf+7
wQaeaKA+DzYl+d8ZPJBBzQvTm5Ye4OC2AkkxHB5ffusbt2zbudAGzIOono/l7kB95lnRX51ie0hU
x+cHxQqFMkv5c0e6qD/WdGjnJwcQgCDhkqhNTiWnEhXHhujckrWH4PZYqjK+9nYeoXSFZJOypbwp
8jkMloP+IbhSf8TjbhGy01/Gidb3JT8OQr1GwNu6pC4ySx0N4t5vy9qQzEHEEeV9eZNvJjvcN4NR
V6GWSo+B1Cn/rQOsylu5MTS7f7eaLEIbgebKM0DJdd2pQO+9f9jcirLtVU3hEQFdg2A+cVv6FYCU
Vhoxj1d5tnqT9Ish1Y7dd4iidgTjvY7gdkhaT6JMdPYmRBfhCGAdK8cabReFBQNRsHXJJ0A5Zg9H
5aqiz6VvGIjMRQ6/5Oe32Rjwud4ROdjpp/igV8NJTSKLDfHiT4WGlQAIcX2AINCDYGglKVoWGd2U
25jxWESZMXmZuPpmFvC7lPX+6s87gkHbrBrUNBlgXwc61uaZMZOz8Elf/XRS/Nf8za3sIcqQXTNa
GBSfh1nb/K1M+5XIEaWWGX6mrcplXaz6PgfzOqQVEecGWuBtsa/WfcLr0RahvWZXOkXXvBnONvjV
5q7XAEY2wnulx7EO3CxIsSUWwyR8rwZiQRyusjIXZKRnYGUS1vw2qGVTOhbrtR6mCE8sz8sa5dBZ
EO5/lJNIqygkdGdgKQG0Q05s/u/L1nJLhE+DLfB3BiHuW8VrFQXztVA3bNmCWitvOcjZT37wH6QO
hcYW2QxZ/YfWrBFLUdll294/KXEUs7YxNJvCtril7mGyAS28jahldTEWm50v+wiZR8Lie4SMk7Yg
glrsoQ+I8cqYVMjDeBPZ3+g2YnfT8dQgZcKExsebC7bgDgcDGbSTLis39zHsLhimXylyzJHapjwP
U8WPiK0PbUhIlXMtCKprs669SlPFAaWz5wdduvQbK9XdHD8SVimX+Oj/1xju/LFl+sZnRDiOtQOk
yScXezJw/+aMRC8FyeBdiGoJMdeX9C52gm6954zjp2PoNxK1rBdymV3lDrrOagRzCayFbFE3TlPs
XhbDwVSZc37xc5unRWTug6pFk3YihZhp5crr9+A0lTXDCyiTHXLYcij9hulSGAwPiZIoMnn/aaNJ
PrUJxncDijBBL0nKjp7xbYFWlCGLDDwxs5WiwIFe1iTTjM67NntOc2BBFuLntBcCLta+JCVK+i6r
AUT4tW/spwiWUzIjU4Idv5QD6vOt5VvcW2Dgj1/Ma+EHnJncX2aVv1kASHYe2nPJ97d/+EyTfcWy
ufSCQ/8X9l6+OCC3ZzEc9aRepGQXWubvgj17RsmZHF1349y4I12fpdEkP3X/4JivS+kcmJPrK/g3
F88x3dAZBWdQliBdbqrExRjSlwLARHzq41tSqmcvhuL4iLVEm+OL0fFR0cjk0x6+fYKdIlOonBKO
xY3NHn2ccLD3TubIbCo0OBYJsnIzuSBDFfBzag9Dytrfrct6PPbTb1L11ZPZ1p018tDoxEI4lmtY
MsXgy5R7kQHfeMo7rr92H/kzMMwO8pqds2AiYrMtg4QaRWuMiV+mFFXlSOxP9l0ro77V7aUCR/+V
Mz3C+FSjxPk0S1GsAq6xPVrMYZ5aOhlFTBfBwXYhgB0K2RLeJcMRDH8W5DsjekxP4UMDXwliy0ZE
h3gioTj+js0AnhPDhLPu1unn5WiTXBCoxUzVJml+322qJFCN+ERMXuLmeZH+eNBPWSfYHXe17u/A
gqHp51iS2T8OuPYIq4IfxzghLj/yGvntlXZZbVBk7lceyiszoou7HtqL9OINmkatgtM4O1383eu1
7wWr3KlnRdkFdIIpyb7iBXrGvZHoj7U5NbwgiUzUOReohBGQBXBSawa+G9dJSV6PYq3AWc2Ehc95
RE0xao9AfR5YJ6dk2JYdAthRA1h1jyLacXOMku1f5rGV09W2Dlfx2/pImZvfqcJhQVc0wwroV6Z6
AXApB7TZ0XZ05Ju3v9uCnEDiBnt3g5E9auz6/p6DqJzSUjP8sD0ELezQoZq4+M+59VvTG5v7ajgy
WB4yCwcXu9gbK6yy1NvkF9ENSwrUboyPOShW4LL5rED12QfzjB0jgnED2FCvwFc56cQhGI3bMfWr
dqvs5pCWzqyFy+ByDX8sucH6wKXMWXBIOwWerN25x8jcGc47vTnlARcjZaCFa8Rvtd2As7aNdbpQ
11eV43n7j5forYD7vc+PmT1mBu4ZWJ3OFNaIkT4xYguG/wSpk8rA6omnysSvtCW0qy+XtS5W1wLZ
YrBoAr7+6n1krMngpCX60OANqwf9vTuFjkFWTShZ5dRI1HrKD+LKPYH9PE6KVS47o1o4n7x+gy9l
CWSDnGZeGWGpRyo5Ybli5J5Ph7cL63rMZtn4lhTXBdDlpAbuxuvy3NoUoeK+gzhByu/h768jTm/3
TMYiYmGHH52siVT+gjRkLjsMnLqN+bR08hGlii8DU/AuxiHcrw0rBe4s33IaDtCbYfkG3x4684zz
y0Z3p1AyCUW6GvZXMlMdAPjUBamIEGPtY61ogSuR7Xhz44kUIBW6hCnQn5wqTpoq1opmpDuYNsuN
mLC9cMLfSkSzVgS5TEXZies9I1Vm35Bciz/1worep8ER9Sk/O4XorDzrQH/i2Zjos/5IR03gtCi6
Gd5pnskcgv0sNTYoTyNh230nlPe5bG8v8+NwgJ3Li3kkgmBGFuh/Qs/QHujiGAs1uZiCHak851bw
RK9vWR1o10I/HBlG6RedE6Yb50edLz3ip/6MpkhsOjcAgHe21QBWuE51nO2z92wA9/0Kdkajt3Bm
bo2lrUMo7BVvtMFwAvEtTnzqUMSuP16Z8N4cp5EDE+lJKPXY39pmrZT1OfA3Sg5+Ml8ufJtH8Nuk
UwIdkTjHLKETlR0FTP+yiKcHAYk9A4pCcy+sAA24m0L37mlQeByj86Ofy3XhnazinljwDQ2/+NSE
AeUFEuUSbKlf+IuIf25jn8l4L+N/pqfXHW3rkBd6WYdO6MU1IKrcXCuieHS1jM9swY9/nLLWC6WO
AHop1ekbQI5KQFGVNcmDLWSkrDxjRtlb+THTBbNAxns9BPNIWc0bHjxP6/Z18hjT5AkduSOsw9T+
V8mAqUwwUP6qrWjjg6drJ2mqASR+phPRLuztZXYx1njuf/HtXObPy6EHJ63oqCvEvMyATEjWrORE
BgwORrM5SBcY4p+v+a1VzE5hq8h8l8bKVH/cZcCSKj2b2DbhHykakvXz7t3N+BW7KiD6ElAUQhpo
rWYKKbPl2xOWFp3+9T1SXYU3/A6+hfSqoOmfzCP0NvsAdcW4o1E1Y32j4bFqnw/Owd8SimsvL1wr
eLZMDYftd+h+9VW4Zm4fPeDW+mVNeE/X4N1Dn8gu/+gl2h+apLkKtRR9raNCvWael9NiUtSAiMtF
C+lE8jmckGRpSSnZg2XrAfSi9AwON0MWq6T06XnC0gQkyN/0B3ck9866O1k6w856iAyPw0sSJtvj
MAXWDVIlcqGqesudTgIe0kzyxRiZEbNWlQDd1J4f4Se3OSHdO8oyH1k3oAiifv4zL0PnGjF9UVGZ
/wbVCyTLfmVGEdrEV22JAzXOE5FN6IP2krXKbVtvnz4K823AyZGXv/yWjm7yGjOfDWDBd0J90d3C
zeSD/wsY2gYeyruDsZmRNl7u84Si03SSxQ4HjTC//3q5rWfHRK68p7PQZlTKJkHf1tErK5Kh+efe
dMScq1wHv/04raxODFG/nCJgcIJeOjdtFYHVnezcaqh3Al4vkNLeNvifAmx7/EaKax/Jnlnsg1rt
dlSJgg6mPZ7fKKzV2xR8JThOicx7xUV6vo1K7/acEjlZMscVhoAYzP6tlGZEszBhSWkQHWDOwB18
JEPVVRd/xAiV4b7NZ3O3Xahunl7CdoQH0Omz5tup6ib7CgcUK+7WyqWnIe3ATONCwo1yrrPzAkmj
rDONrCWKsoBmFxyqGKeLpZ/YRP4nzsJD6hxjfkO2gYqiKjkl7FmDyyGIo7X4HCd3uSSBe864OsGX
heajhCZcpbC1hN+eaAbXmzZhmcPmjsgkHwoKRzqpClIsZQutJW1naPqP5JknCZ5PuHAy+awv3hes
CXCL4lyt/dPN7Y3r3Im3Au3TvLVKQW7Jly7KmPRKak5c3zbLhgswVJelgJfs2/tRXY/WwS5uzxiY
mzbb25CUrOavfJDHaMmetgfyQDpzr6kN5A1IB1niEdIb9Ou9+Oj0KbruVMziZshsQgRJLhNsRRaH
oj7YD3gFVS1OZGx08LNXzZjJUGBWFjoFt0WoXZ8MlMlVDK3imF3V4s7N6Ik/hp+hdobX9GuJ+gtp
32C5LvEeQ7Vgk1o4Yd3jIjOC9LITJ7uxEEZVjij0FVowzh+f2HCn/NHi2opY2RWfAHPWO4cQXHGC
/wU8bqXmbBWtAGyYKUczOeez2PBXl9Y0hHR+pn5v+kIJUiTnawsOm4q5eH7id7qj6gpIRVDGCLOi
w1oMigueCLuZd5JhtJiK7PBVNxhT/me7BAS1i5+NBWn1cpcfuRkCFhcA1V8+gc+TqzcpnrGkUswb
Xx2tuS1kkwd8WSiHduFiKRFZx+t0qrud19xDXov9bhnG9iUmBT/lAQpE/oCMIfWgOZ2jlNrvPcsf
ZEu6etQorileyglzKThUNIVW4hUa1/g61wtcl8r+O0sz2fuDhbqOA+tIC9+QLHamLPRSGiQMUmgv
mr0Jb0qF2jsu5bg44imLZirD85QliEDXWtY8EBK5WlYSEnWNbr3vS3WBMBZc5ndpK3ux4q9zlV95
sUruK6oJAc8bK5E2ev77rXvOgrAocoqBYdtmGOb5rByN/jdOe1w91WH0nsw6lKt73HKFI+XW47Tj
sTfqF1A7sI2IltYuiM5jklzY7oR9iCFSH5Y7m+yizavMB96hsmSlowB6XRcocwJ/b1u7iowEmjac
0bW/2fP4i373vLV0EZoogFhmz3ItEBSdw0LSdatWdxMztAsRfKHTbbz6GrukKoURDvIinU48LYLi
myybzFTvJnS/tm7H5dRocMAaSC1/UOyjl6Q9k3Ddvw1pTEP/npEEh8W/NBan4yD3slBXPvUmsVMy
pTAC0+kPgc/Ue8X5zywZhqw+TQynzJuMcFJRK3Vf3X7jgUHyQl6m8JcMJvhZD9TTeoMJQrq05r1V
QxxtbLXlYn1n8TFnizspo88Qri/nUWRLGSOJxra21GEmzDYSQkAk8UecjUMqlefD5Go3jcghtJGL
qEjIKlbQrST1eNUd+KP5pIDCHeTYgJDzRGLnf+T0FCe563XDHdASJKt14KY6LmWs0//P4ue3/hVL
3NfZttdlqPnOV4G8V6A3UkRybK1s0PB29kFnPZHzEg+dn17bs5mKoEwlmGuK8pU85zqpUOIo1MPl
1/DAvuVHfqbqGVGfcZe4e1hTbafPZfTkqsuwgMpcJyjIkvi+OLHTqD+oHshDp20Zvtnm/1RQS8Ki
DHFRb6oZxckeS+1EvVYKuCEfY6VtM50jRF0mHIpHFPhGIRJP050hoNo4CGSlMgWmoEFqfo3hREN4
3Q3zNWHp0bN/ZivtmR7MsLNKcBVFkAZ6G3qykcHgcvmrlZa8fImwcOCnhcfsfRRNSWIyafcYROfh
fKV1T9dCi0eysW7+dR2gkmKVEujHHsUSOvncBGTv2Mxk80x47Jkn9KM/7FdThuMe58t3QLD1SwzE
0liN1B8Xzegf5xrZriRf4KxIgu/0JN4GhW/NyYdxKsf1Ziio5YLWZxJpoGzlhI4jiAMvhxJrO+1U
+TMYlEnd1/tYNgOdqMFbodFdIS+HKzjRzzzuVoWIj0RNQ2BFpCWani/L/t3mMTjqRP7zpr0p4vyI
6uETY9cwhpn6gou2zSU6WKuQ2CzukiEQZGhBlZDs8Gh+kXT8zrb7FsD2e73Wo5ZOAK4Kmztt59d9
hwNd9piycLw6HjguRq4u1/NeXY8jvCbgBx8P+hI6I4Oou1WnicDWammeu6sdo5jSl8CUOXMmGuH3
bNdEyDjmPmKZW9hkdYZPd5DFqUDJ27aHn4zLxk2hzDd7Pr86qyn5NonVUaEYr2ST1jXPu5mrXPEP
nVNs0SlsnrsPb5M8B2E4ytcVEBDqjmRx1DHwndFTEw1xzCCX17lTZJmVn//LB9QPjg70pbSbCsIp
J+ndqjnK2tPlmoXYIOVaxPd1+94dSl3lgOKtim4+z2l654TPEaKey8SJaRpd51hEPD/6Wf02N6IA
kSnxm23fl0FfkSKIv481dURz1urJPc4yaqyEmigfpTFLcVt2UyHegSRz9C2xRI/vOgG710U443aU
AqOedXZnuBRpGSpB7Ro9hCY+Rb/e7oL81EHiDQEgekjGxYy1LJCV1PteiBX9983l3G3nGQJ++Z1P
ckExxZI/Qc6ch3q7fShiE80K8t9lSmnP0fMlICUxZExFmD9v27XlJB3RTatyY3kE4YYOCAyPjpR3
oz+6ulWcO1QusoQjWBF2M1n850/bjLb19ED5sZA0jtW5T7wsHAnSqGQHkCJcivROeW5xtp5vxZ1I
FxFo8j+s2m8JW63D5wUTCuUPcz7pPeB8FHhWjcBFt7d5fHXgyBQoak1+s3mAuhcnLKT6sizFU+2o
YADdCAf/ZfZigM303kmipl4AiSqtpHuXaohLAf9hDghKEimrSDECVZ3r9+MOR7LopL6eZ+55jUcv
4xd2ZuOiW1Pu+Jwc9LUtQiD/+ciY31KO69a9TPfGopkDDbRJngPy2MEUyBvAnRwgtVorEWF7m7x3
5hLGEPX5tctdYfstAua2thv3a+TuD0QRS1kzH5JJ0WERgL8662pKl7x2FRlwE8G4VbbHPv3INUWJ
fkWTSlOomSsFXfGRv/oI00vlH66wJICk6+MZtcWTbSVPiP9LgslGLl6BISuGNyYdz0+g47sTZjtL
C+FzP21lk4iAFQpm93et0RDuKCPLCg947Ka4PO2KpK827wiIAil4akSMFQFeqWTuMepifRoLCqZh
04BFGPqPO/ZJV1rUE+fEK6Uv082urKOqkPnWAS0P0j85q1kimIvYo4m7b1z+aCV+WcaDU4vmvG27
6b6RC18+1jTQW/1vqSb/XvtZIqqt4NbQEp9gelzE2amWHFWb1ZJWra62dK5NoDXi0U0Glnlzmjeh
u0GQhRzIIyoiDJFkL3gTfViNxm9wyWOObkQBw9WXUcLEto3p0mquIUbyp38i+2lk2J2bKsRBgtGr
LpUta/X8ydXAzRbYn2JwmcHb8fl65CHJ8BBy1iK0tgj1uOQsj2eSYJQKW2448MOCjVH/XNCnupca
aJK6QYon/KncfeM3JWD9aUMKpWd3/rPNlup5zccE918dMIko9CO3F/C5wlZMoD9oGpXJrqfgrTuk
v1vpYb1T0D9tKmf83UBtBSGsgXRYUFLs5zkQcmvsdmd0IWzG9ytrIGVSezMKKPVbi/tuKe8AzTaq
lSRKlxfNdlx1JqtZBYVBqGQ/yfDO5K8N9X4XVuJKxkLZuOfhA9hPXw+Dfci9yIy1pYF64rHMs64X
zNGHRQRQm/i3yqN1mz3rLKDtgW23OmKqyRXbf6bsigssDn7rRWUZYWEagZXv9f76Dc0TGW8OewgF
OJaNdLdHeR/+hGQJiP8yQHUSE7aJHBWdTMHQ0R+sldYJ9Lp0DV5IAxdnzQGYiRL+FMAUqA/oyZ+1
RyeuoEoI71CwDPTnnoq9tLJvMuvCNosM58oBczFTJTpSTOYDLKdRkVotPDNlT+xXjYVkewFbT81r
b35/Os4Lqf1y6j1Ut1o9zcGXzII7y6/xWyOXYGZHUpMuRM4Q0m0b7ml0ttnSu0i++T7gN9IW/Bw7
t6nP5YShl8+GHVdRTJaA+uulUMKObLDQ1i/CCe2WuyLlZyxJzB+1MjS1H5ZbtfvdNzz5MrQ/1Nac
R2/gyGniNG9Ke1snKc1L5F+mB+uqE1lhyUak2Hohn8BNnRC2HIKbLCChy7VD7vXXxizWLNhNu1lc
08Z+5sddjCIixjAizZn5tzy28ZdYasK33lDOt3Ah13xtoVogNv/yVGD0l3S4M3UFQ/xDUniRBHbr
CVW8POiQkpfjYh6sIWDUNj0VhkBWfvNpEGBX2w4JzoRiu8Gnk9HIeQfqinAcsgyh+EeWVE7LdXIN
kIHCzAEcx/kO1QxBisH329Dtg51DLy++XNWQ+LDTz7f0NDsbME78Ab9rssQ820AB5zrGZRos3HwR
WADOEsAdz1Hcl2aN2xj73CG8IPDXX3lUEct9fQUhsKoxExSvwZ6kKZLTxifY9LQQuQ6nTDSP/Fne
/cGBa7TmgMYaPJLNPhugiy6HduArBYhfwYi/a/oSJoWfx+cHZiCQaXDgGW2r+vNofYKCUrmB1CmN
swpHNCv9jW3znN6FOtUPPyAhSnshtAxBDAdZNlFOjn1vsbfZ5i510JsmNnrdGyApfKwdMOZ64V6f
kjBphL5jnaUrpsi0272OymVvxSqL3bh2AYu1JJBLcpqdT0XRhlO4VkVA4nuEf3fJdpXnLX2C+oVu
X2yvAk5mI2BseNN+cO5oChe7M8USqmkmEkMECjtlDmxNGNlNME1vKKxur0bmiUWEwGG+h1ZQ3/BK
vlL+eJv4FEW7MYaUzaNDyCgG42BHTmEYPzsmVzOXxHcIA2INrI46vRAxUBk5ZR/siQPhYmzeubHT
FaAQwdrZUvlqFlY/RJ5Bs5aIm6erpDz+IJKiI9iK/r1z3t8fM66y7FCC0J5zrzq6jXyWgv9+2sPp
NERCRpeWPIIVc9CQYr3SHyrYRtaKK6/WtLBEfVOa10qoawTWsllQEDI8unfmYomkGn9qRwK04Lc+
lgaIXyajY+FdJR3BYedZ8+S1kvz3yPOO9osJZB9M6V2uQ3RE/PLcgJR4JVR7kWxaVzNWcqFK2usp
Q5voyMFG0vQn9P8YTzlDTQwF1fkugcfIFEMxGQBuM3hoFOgs3DMI1WrqHxOkduaMKGguCu1rEmxw
h0qgaOlJ3/ZwmvtSP2u7cqA97ynlnkIYHG9OgBQmPnQXQ4tzyUtFT7dbif6fPZKPq+O0AeY2xgS9
2Dk8r1+ZfjxXtfjz2Xvbhz+QEUiwqjr7s/Wsp9evsDXoa39vYfdLSJft99nYfV9MsaHXyApqwvnY
6CHbxNIaeX0kvx5HgFmNJUMjIiEIIysXh1fG2T7Pz1B13epKrvqb8agv5hatzu3OQnqHPujWru7o
R7Alp2fBFZO7jayHJpfR2c1RLmm4xkwqLEENZfp5kfX6hX3ziZNKpIgXYQdc/VPl1oWyJizNyE1I
eGPppFqFRMOTIM7bbyAeDD/3p1cizpATxc03HluEiX5DncEcs6+2YpqB+sO36PmFianAs9rE2lLf
xDTHRW2SeMZH+I0v8EiuGJyV9r1Eb/pZrea5adLtZncHQitt3FYlEoFcLfZm3/FrjVW6CHzQ/9pf
gPA45aFtHMdDIO4w0SUkZHIapY74HjMMFfVOBuSuhwjhJIYWAoKDqvE2vqVlK06BMc1pfE+cpDVW
DJcu0y7MBBkCKErZDC432XDiZANOKto8Zo5YPUgJvUtX8FHVirfDQzohUWpQAB9pTg4ZoNHUcAIc
krHYfEalDGs22/tm96xhJAhX+6IGbE0xnymhV5lCdagf95+2ybiye07LFuzI9wmWjDVGclQ6k2BM
YmwisZsFKpGa7LkgZpYfrALvl1RqcePQbE7vsfT7hcApTyItrOd+7FKIkPIWnCYO6DmSc0ZaK4wl
vpZ0s457JljZRpa8N8VKojRwVRgWxEKS5ArWB1GFmBC+BviNzd0AQU3v8aR3fWfJrNIUpZBDXipn
DITldMwaBkhzYAYuO9A56sC/XF0fcVpriMhqf1g9uxF4LLlU8qjX1twEF8FbJyIXaf8EryVAkWx8
Im38rMOmYkjnj5DG+QWRFiOu8criMEMVwUVhgwK+WuQ2HvFlYJFbvYAfXhk6WCaakAk++9D6oq4u
GRgO375ur5riShVU2b+S3cdSYSdjwClsIJg+Un7iDAFh5dxrNGtNNaNKKfcPZ6AmOR7m95ojfchu
/kau1tcEvYMRINVfq1G1rpgXKOTTS7lQfZWn/LtfCB8fjDbB+OsqOLkCSSCTn6ik/q0sSq5f/p6j
APZhG5oqwYrc4j2TuBn4Nue4d027YZn0m8N0jCtSFgO8NiSyfQ1TNZDR4Ofa/7xodEimwLkXsqB1
m4T2gASJnYiLvTR1JQQjzOfRblvzP7qnNNamhVqwepyNkmTexmu+ghNCPHG/O/RCdAcAu46w4zAp
zY0oiqgJjyS0zKlHC7aH2t/levIIx3npSv9EeACESANYEkdmXVB2CON33s4Hot6S2pHiWIXAoF3I
7ENvi/juJ5rg/D0FAkokoZPJhXvDPLqxvHokZ5igToHiaEPycJ0fkLykTO+IDv2JyDSU0Qn0Hxed
0AfeveykZKcWj5JRrIk+Twk6q2hJgjCKWy1O9+DvgJig8TrLOpgaXuqFEW++sEi/2e2v8ql/7Sag
k8jTKLZXjxugrSLLvUHlgzzBB8Nhh58MoLU2z8BGCeKdtnwVs9Ncb/oHClENt3nK0wLUNHmYSaBE
5MelvL6vQkJDTVkEVI7cCL97ufRwfFOSVX9Z3NUw8FhvfBIqWVR3pgjSh9WdF5Lc3OLf4CDayfZp
V/LWVRle+4XzETh/0AGnPPFzWjc3rDcNaYVDWOYIS3m59zFac5wUdAq0nEXF7qBpfcAsk4U40IgP
SfFrIZOfiBjjsSMQA7NRHEruqN8PtljWH+MloI7vewzTNVE7gd1q9CP3bEq/BCdIm4JP0jxSgw5t
FYDyCtYXZjV5lfE2/yL6TaO61aflwCJqgtiM0fKQlE+h12rI2gg1yzYCPTpaXbivaoaEZBnaTnK1
z6bKXlv+dPOeWddixgRHzzqYqQlTwcrcfsk7csYDCZCqLzDvhmM+aRqhq4+SipoX6O7OXWqZ2w3v
69Vs/z7pVwuNIQ2A7VpeTGqO+Z+tkUqjpTzr8l9LPy9PLni76UoB/lUKap1c0cb7J59CwB1DS4JS
xhDCJqlRFxyKqb/A+tjtwbIWGBRMdNk6oUiZbIp4YRD3+SrteGmskqbnEhw5Urg8Hu6jKaXArogm
lnawxCwyTFaiNSRcg8qrXC5CcK1i4XoUdj/MlsIshJd6aJj1ZVA5zccyqSNx1CctwyNpzvziE6jL
RDiVZU1LLhHVIra0DrXxTAszj86ZGPiQKsW/mEoWEmPidWjuWfCF3pnhnzDBQIDi9wkppgbqihwa
3W9ZOyFzy+8vGAnqvjUk9RuUJRJCZkQlBrPgJFBGGKMkpJdE2crQuYaPkH1vij1Hm4hDMVDG+dyt
4KV57U5jxPLfWpL1f5s+AMUz2uuMQoNTDgrZHtTh0urjVqoodBEFGD1XBFuxiIkDOV9oKeEB2jCY
vBzKTogVBlBS9BfdvgdBbaTqfjizKEGrZDodv4h/92pwt3QgBnnEDr+TCYmd647mWtYvt+ujUZVN
fzesKznXRcPFFb/AJ3MqGlTCYi8e5Nd9gR6FUId4N/D0Ov95824eUAEFFHvnJjnqZkpebFQvyyvL
UphSmhRzpktN1yg6grphkgo2mdvN+eXr6GeYeV/WESr8KjqVD1OhBUj3Bd23QeL+6/DLs2taaOsh
Lzfvr+F8ddLHn854SWDFmJdhIDcZD5dxU1jIFMsStH/AAGpwFKSNOI6L0LyulYOwiV7D0byQtCS+
02vLoz8j4MNPwyo8V9Ghs/xiftjlqq8Yr7NtFlb08q1ufvJlIXUZnur4Y4UkNOnE7eWbsHbpZ7HH
/crgFW9vc35P1OA+xmvyEUVfWKpf+IfPgJhKp9Y+IYbHP8h/LcnpXOTMttc9CwRbi8jsWFCiehuC
vE/zIWXi3fjVQameItjiN47ln7RxvPGeEwQt6w0dAXioAUqDiHLWMzBewuE2WV4VklDIyhFt5p7E
t8o1d1bE55fkW3f/Cmf5koDXJffwArKtjEaZftpVGrk9SOw6CPQaTBfo1R7H6dPYnUAN/Xr85rBh
Er3rfHiXBlWEzLzcdk5wUTF9SgKV3apSYA6U3PUHCf1gpg0pMPZ+WeetE0Liu5ngshnuUYI34/kO
dwgiUyqcsvNSAbS3QBTlLD7W4pocSoD38BjA/vDnOqZz8t9bdbIMAWl05hvcX+WJAjkpj045G6P8
s13E5OE/+oXe3mcg5SaeqHIia6EVxAuMjqx6Bd9A1fyihxNAW8qmvQoNjsQjjX1vV2FcvuvTr364
aUVFWanYyGJDOzDkLivQ/oGdwbabt3uLPtgy5yVATqPrf3cYALrMnzqHnYmKj/aZiYvEkMxoqt6M
QLNhlCMXDj1Cl+kc3eLODx1qUZ4m7TP41ieLjCF/7vE84Rw8BC2zmuA/kigXgeuo2NyYKaIYUnNj
nqcaobpSYVw7CotDUJ4hyve1Tj/aMQnnJqz9EPgknd7gF02d4hugWui1rQ53WNEG7WH30wMUV84m
8+Rf/obeKEXx9AjTz0s5wCkFe8owpP9irWZrqxb+mPawyl5mrhbufKFQdyYr8qfm4F+MESBSF4B4
lYcvD1VcGKmYzfx4JhvTo5UdFMf0qNdW7moAcLdO4gI4/EHk67+MrmdQxMghFGLp67yl+VaMNTpy
XDnZDh2TWo9jFS0joWmzNywTu6H7jYuGoSyM1CPTn1qXSrkXk39ruP1cIxbFTCW3gz77PObY61Eq
w4oymonyvUT3XFWfW99sBKhUNfZ9bwwee6hacAoaDE5s0zIC5KARPAGu4193jLPsrhhcPGFpuLxO
S6i5ayqUl4Hx1TDIH0Dtrb0BNJvTv04MfFL9Ls+ET4L2CU2TYXhBF0rQCDgdBlE7EVar5n9HCDIE
Pk6E7wFDmVXl67khVqSE1qB9Wz0n8VaVpFsa0P6G4e/BI8n6bTVI9L+GtRXRMY4fyFZOZGhi3Qul
Qrr45yJTla5Kg0uUBwVVysjH6l3RmA7fgtN334G6OglsTn6hp6bRK0VEV07t1KXLbrcRzOZQaJ6r
FIafwxhEQij+s0bPv1FyVPEamF9K3Xm1vwtKqF1SKuL+038iazGWqVQyZ1dHI7wPpPpwZRwJtQ++
7y0jX+VQ3K6x9qZdVd3MH/VfJH6vDx9oXYsO4oB8Ix/PUivE2sj6WfCu2iMiDlgXxQO/7CmfejvB
33xNPjeIX9cH2YT1VYiZ1SPcQHd4cxvhC2W6YNdCe/98OW6bkVd3tgE73eyoTfkMP2wwI/NNF1bI
zEu0orCpNZ5xfDAKTu6XiPGSX6+fkWlgo3JS8G8q/Yh4OoVLmrot83+CexE2G7nn34cNryC1UvFy
IbhXPKGAg4mDru83jpgHqkQferY1FxaTXwe2LW29VSiL0ZDJdSbYT4u/IkzY6rPS/B8C3bB39kxp
/bp4lPFFLOKkLoOT52kRs1OafIe9lGCGdD51Uj8789cR4rc/hnitexXmPEkCkQZjIFqnvofadQ9j
5jNDQHkxEmRo2CWRDigqKq2EHatrjKF6zp1ccLnI4iB7qGYuvtUferSoHD4Pzr3JXtNX2PJy8Twc
LfA15FJ4fmrYezijG0xAIaUpWntwteexR3sofCgnOjM8QXvmYlpaOwJcgmoX5pGt+xDgF1SpdSoW
YJmt6mZhg/8MabE4A7Nk8EPytsCaP7VLFSZTFZ318hfoOXS+WA488bwQRUNfDQHjqnsm2v8Y1B8n
Ar26vvYhPv5I1rV0bVd+ydNYpVzJmFn/sniW7r8RWNSIG/xCeB/FBFLItFmcVXD6I5gZstFDz1R4
SukiBUVHakL75EIDo3yPzetDkG2X3gSQocxoXKngRcSu8omzQNokIcs41L30vzKCIOhlSzmhjySV
qeOkYubNV5trKIeCgRax/9YdZs4i8GAVT71JpLi4JgKR/x/To/HTMnBJX0UHP4d+lhKMUDIxcMV0
yrNPKPphwFzi6f+sFpcVpXRaWgShbCHt3n1kdbS/HUyYzHqNNn+k92uzE83pN5GrgWsutp+WjeYb
r3Jz5AdxUDBbydITKxkVBt15QJY4Qn/hz+cV0MwNZ4pw2p20GETQyThm5df0da503+ieaEpP0W8L
FBeL0irB94NaWKW73AmJddQfmBcdk9gMwy1ZR/hBv+driOLwdq3Iu2npTMQphlBUROkrsbHWnJuw
xDBC/9+qkVdmj0CsFcZSx13Jdovxnlu187KO0em3dacdXWn7Zu8hA2XURAWas/jhOf1mMDTbsHrO
c6+dB4a23fEJTOnVTdbQ84Xpkb2Dpw6TeUCkw8QV7JDtT0Nf/R80l3MIH8z/bSzl0v977KfIS5Ft
YzK+wwr+DsikvbzLfZURegJmWor5mZ8khn7jPx4g60OddmG6tJnFW7/cvouaMy4JIehjY634YjZv
xD+Oepbg27PlXwhPVY4s15oyehUqlkVz7L8ZhXBbmGsA0x7tiKxVfYhEJJIckdPC+/2NiEHxWn0d
xCaTwj71G/uMTcp2AdRQTGAI0XQnJz8s5ZYXzBmcNS77qk47Nnv9UgsUF7qarM3pBZ55eAN1AXsv
F1qsZRBCeFqqoeoKNI/jL5JhrSGzVLVkKSCBz1lyotv3ZiPwtGqtBx0z9T4Zmi2kOva/6h7SLvfc
i2Y5mUhJFdjMJgGG/pMDblfLEst/vq9swr5kmvWJhw3W4zPiF+s3mHU/vN9HJcK4/8L3RWVvpx2k
tMVDHmhKX//2ffudGyHWNTR2qXcMW3tQoqk/Umzib2TXO2PWMxoeF6y19SDkrizEXHn0PpYe4STG
NUNxfRWWpaOedOO6C36qm6cAU8bVXN9HpboN57QQhRpU5yEMrorlaMswcJJmhWLUGZNwooG/jrJP
BledN7Iou66RpzvY53Jala3IoJoH9JfWRXxuGBeE0amjj90qiie6Ql6pEIR7l4Oi3FneakKykNk2
PUqV/2/7BpvNkhg0KsXNReq9eIpWjhD8LV2CqlW1aw/JQQ7pWtaMxS/gnQjJf1cfXtsSHRCzbWGO
T7uWQqB3m3kfhq3JDygmVj9TJG7JG2NYZp1R0PCzVi9/HutXQn9IEnUylaQQQTRDZdcJ/20oTq13
lYqRDCi7kd4DXqpq3MsBaJkNcpLpQZ4GBKlz8hddfKCzhLHgKtAkLiydfyqrUt/w5+8Hcku8f7XJ
I6Qbd9btquh+U+iAzDYAnZav5x1Tnz+ci2fStks0my+hgCEcJlFiM37qdG2FD/fgs02Q2Q15SUxb
BkHQFX6cGkQcx2YaNh08gi+luTSdxx3eDG1tz0gy15HKhWP17U3ACIWKk6/F2ZL121CypOThfA5r
sD9KzJvOC8Z4DvZ2HvKVl0JaPB1EBgePJoQYt261RNex1itJxgxa+5tBV9/mXH/0VgGjDBZsZ6od
MDnSRqbD1vL5UmkeI43Byn8CH1DfNyr4U2IZ1v+l4/kRQZ6InExXsHCohOjKD2V/q42NN7YAtJEh
UErABT3zIOqTcp3XmG4bHlCGiP21/feivPaUjBUjmJl4RTp8wJtkI/c8G3o/EpbmnPTnYOD4Broq
qDMp4LEWnuyhe0Kf5ySvWw5KPQuX2txekQbgRM+fvggX9VwqiYj4KEexBpV58Brrd8BGJt08ZDch
opBK4zEptM0sM4qDireq7SI/YLlGWZhhuBhk9Fkk0esn9YWfp4V7KWancO1/v6I+sTO7VXD6GWQ/
CDbIO6HME+zNEQSV7KZFOVKH1+gKO05NlIfdqyK1PiRdlx0+41Gk/Iyf6X8x+E4w3dE74EBoqlsh
oYQkkkYXLKQGoxkJSLYU9tnJuAlaDT43Hw81VXtcNxkrmjUnfbp6F6v8mi8LiRJIOAtIcVjksqW6
z7mAvUsn95fdYgL/q7U+zgvy8YSk0vX7eBOZ15WuHW0QrLd3p6Qwma5mAUQlWjGCfUsoCFtvACEt
CAxL0ZKt9qqG8roJWmkHpfHOECHhvR95wtxVlJuReGoa8gsZRRLqbU1AqEXnJxA6uaLZCrd+VdEa
QLFAuzzbAARGafLQlmOT5SQl8eO4RwqahOZszi/y4gelyr8ifWbTTJRVO+Cttbs586n6Jp+jAWHZ
X5SwsFpEF3G5+FWmOZDHik/szsLUjlhqgtx6SjVkteP7k0GXFfOfDVUulQBaH7LUPkRdfp5ldawG
5bT9GtWBj9ohK3RdrxQy/IXx0/zlhsjLQEEtBArKPnpYyXXaQmL3v4r5fPKiQKpUXIPMerBWz1Hq
f1rHinPk9itYR01bjIIpvLCmJz1aPJ4NWbSETBiRVka7D7m1lItbK2u4cjyOM676VsDqEQnyXLWF
3AiEAGxMaxec7B+yMKHUtx3NKT93fQ0qUphfBvCu6Za8l4Jwk+XmYfNEGOWVsVovOx+GagiSHlMu
OBYvMBBJpR/ndTnJCe/W9H1c9rYY7XJQvIYTJFBV6VxTlXUiT3vG3qotWBFSW9Bw5WAsJL+24vOx
J8poG6biuOGkyYEQqAsguiWMqaHQ7USM7q3bFuJIXGRYwxbVORYyJw8L44vh3vpd8hUr0tpQIA8M
3scEkSiJ0SzhSitQ0zU0zb6k0c/OeVVtPAJycbJaJofLCjkRb2QCq2o3qeiJ6BWT1cIt47HQiVR2
Ku/It1hOQC9w4/cp159psSmgokPdExWJVT56zjyOuh8r6ZTN0v4JeKH4ZmJgzwbzRw7uuHAiU8sV
mReuL5IU1yMsPOysONANtDSQaBdSmsckTH/KRxO2KiysorOmEoiqahDkvaw/F8VoC3p1ov3DoLVx
3JENrMmxDq/c2HDQi7X/lRYbr1IyxX5Uy8MkFIertD1aWTg9EYz/gFpCCQAAAWhY03iC+tHb4pJe
sTqJrIhC9Qn1AjGq+EkqGMenewqg6ez51i0VqlPar0JY9H0rM3gJZP3ibZru0Mmpn1bAGzd92UOj
GJDgE7qbbEhjgJ7f5DWXvnE1qeH+jpdwVBKHkzgAKIWK5Iw17SVRhwWjjCDzIlFhffbQ+DuqDGKb
ihlVc9V2HK7PvSXGlui0IYfOzZkXBY0wae0OtxqNhJUnyugpPlVyKQCRx3Xaf7NDf0rdddK0AUQY
+Rjah5P2yDInmukhh+wVSV2DIM61R+WtTWJu5OCxF44hfO8K+r0u9YRdGTmnWhQz0Km8JTkNx1Cl
cYiBe47Gb9lwaP+aY53lE2Z2IoQyoOnYqEUqt24QpLUPGLdx4sA+yCHmM5uBB3d8p9VzSjNpU6JP
a3pujAf02rfwBVo8waWbsdLj6T6JNVbvOPvd/FVv0pO0ZjeVp81mh3/OUfZSPKJ1DCOkQ33i6g0x
yI1BGW43sUkkmoLLWR6QkBf6uXoU0ZRa4MJEVGk5eUhRli6FOYmksHLxvChCC9iT7s3f+h3KbBBp
DczbB5Y57998dqmHlcLDwyKWFCb4tLfFKsQKdVnzdRIHq4X2KUDPI41M2EMEbwS1qu6uf6G5MYFb
WWSFlHpwJQX+TiauMY61KNB5+QGGhg1jrqm2b98v5zMN/ymBsuTdfBZGHIxMcvFa5fksB4xHZctN
+++T5W+6k6Xskt8EoNgSaUdvKjZXfNG3WxfbjMFkSbIb4YvKpUF8IqzZqawZHuIH5UBEe3OlYWaf
B+ditB12GOv6SspbQlUYpwFK1voSP6DZqAwsDasJ3BTN6frQfhENfYCUz3Jf4lDK4mK98fj/eW1x
2AW4z6soVf9vn8+CnW5IK6xD+KFEhTjT5KuLI7zDGmBHvOrp+JVkg64SHnXhJVSdVaH7ikyLM4is
+kwKXVD5air+iS3O7oHshw2ErbOd6NGTb+DS//ImxMHOeH6IjI+gLaZbkuJmvSdTkz13DGggGDOk
KcCwrg2z8WFLUVYThdGAjCNvcMaWizAhCcREU+pbz60FJ4RY09oM1kLELHPaB3ZTzXJUBPNbJRXU
ehmjvHvdnsOxw0cevU9N2PvxTRRYLnZrC3ZvQFxECX89DoOU8yusxvLhBwbTjoO4nRemAJoJSdIe
59Uu+7bwwwupVNif+v6hGPZskIzEFCBh8Ms6CJXCwiJdw/gKkac3cWBb8wPJAxzx/rZ6yPVKm5sG
45sRi5CObtDI4IXU+ndB88bjr5oO+Mpd5D/yExx6SKTAz7C5LZEDiWNHocZyAbcwNsfxLDUwAAdY
8VYzzLm+Rii1OKv65SlRNum9dNz6idjaabVva4rjDevFwm8wqF8XmjojgOV5O3KykHUaAjyXb6vV
y80GpLcfJRAXvxE1be6VPE/exA/bunrFiCwmvnuKL4/rjFm0MM4vIxOa1auA2CUnsXgZ1Dh9Br7N
FfWe4I9Lmj3Asr4exulLHrl5yuer2EUColCxsvjPYEKA7ucon6LzqeUa90rR91RdnQSSUCACwlv+
FUoG9b8EptxD59JI9wflt7KV5li0vMJojrOFflr6DO48Gy1763rcn5QnpQviwxFCAPym2wFvpmVD
WSnGGr1ag1yXbwVBSi8IrYfALeanggIHhY2pRdvTuMMLrkpUh8t3FL4pfXRRQyEk2sNCVG4YLGEF
E3182bj87KoQ5T3SPCFay1tw0IfWUncASq0+BuBcAR1Rt8MlbFO7U6TjVAyI99ingzOBMKxzRaMO
cQY39OwaW17cYJKlVnW5dvL8D05BXGzGQO3cG2LX45SscMILNp19R3PuYqUWMnvEadX6xhmYMt4t
oJBYVED//vX/4PbwIJaGe0IdmwRtNtIn4NqZQpqaCL/n8wD8apawvkVL9Klbt0bd03ssBFHKPOSR
EWLOo/vdwSFAldHEpZM6dM8cp4frpEzKKB9KvrjatSNZ2VabFWy1pv5kN8TUGdeALBE2b/ZpEFgE
ExXcruGgMkgtUJrxE0rn/sHkCBSMgkTY4RsHypFUBgtPzNdgbGIHBV98xCy1ruxUq/UcBnAfBuJt
i906RbiW8YIJgca2kZbb2BIAmejqvnnIPjTa797o6dOTVCxLl4m1TnflF32g/5c3OkI5sURUrDZB
cApJCycVzTYmOk4NzNYyBBc1Unad7i8G6LgZ7+YIUXtv/AGMig2QD3aHp22WKHj13lmOq3Q77nRg
I+dtKDzgoDKupVFHCbX2YtH7shJn7rc9/YUYHVjh/dhoou/AIbJRH1PF1d8AxWHUnVNWv+cxuM9f
99av8LKTwxekihGPvoeD3hmuXlK0a6K5akLVtoDOu5v8OPVax6+26Rv79HKGI/T2UsJMjqgpXiTh
ZfV82fBW3FCB3Q29Ohit5XjLaPtgDorPoRS85Y12YLQN44vyfF/EES341lHBJL11+zGKGD4IHuCt
OuxvAZZVoG2I+bu4DS36kAht5MdtiEEf0JP/BXi5PMj7+TDGM9frQ/09+aGKyuDtitIfZ1dnxWiP
TJo2zNHwxdEghPTJoj/ukFi13D0FWrO8DVAdx+HYCDXzgwBh/DFUrB7+YVtUvrX+3wdkk6VAFWb4
vdSeKWXwgyt7eyevYYhFcjaDagf8JWxprCwqEL3JSWxj6RL+DiPx2yDmOqBBFCi+gkHwGGCBuuCj
ElWn11dXSjxdipjYCaxma2PbG4iqbhbPq3aFRz9HzVul0Lt13HQIo7IvvcZzVhYRYInZKB95gQ2J
Je55C1sOHauY3ip8MPTcqzh5AqICwsxqNF30Z0m8CPPOAFQV5KvVC8Yc4taIgVyhHMKC+0FIL1v5
uD32Z/TL5ZHpvnmAdUHcC/tUu+qAf+mQ082ManVQqbm+4mwOxZ8cu9Lg3KjKERcKdGGujmV+uV5B
66BWJ+TuFEFfFG9K0DR6UfldeSHhwJ1gVoYGmYBak0FqvKNFjm1t7nVHTPIlLBfNxOvk42ugmVZt
X0ctjBWPPjAi4wNR8qK9PJgLj13nqOLhIc3NF3BPjKh0GD2FHzYaxY3hWAkkxvf1o0M88ag1jOBq
J+yIG/DFD0KYNXkKsTGA91WTMsEaw8NZ7In6ltHR7BlCTDLSiJKGH1a5YivLptI1Rh6pcL7oAxqR
XwkJD7DcQk9zXqKmo5Uzkuyws4C9BUElQsVzJxMd72pGeNv0cZdgvKb8j6QLkBgLtjZME+r6f/Xm
KUT4bXjYw845qP5knLArqZdOCbkppapHV+TZL++I6SP3oBGXFDMOMSaP7W8RFazffVn0xqiQyCH6
NbIE5V2OSSsPCIAr1DBENFBNBZTp3hUBRYkO8uCY49RQNa7BRUuhkPdy76oMfNa0xOCCcoWj96ob
IcnPgqsdg5sp5KPczTBy8bWFbZkuh8oDbeqLpoTBoz7ZHbo5ML97v4WMp0bgJzcPfVGSUM553vK2
Oi2J42njnNMtGJk1tRsb2w+wvJePVC+g0yAaNv5HuKetilICoBP6w+1vhbvsgwgcGpLpD6WxIePC
8qTjOjr/qQ/lOGGZbXhZiXeX2DDRv6jQWJPLzgPm7ThslC7gNwFiCjkFerUj6hrhpWJRwfZRJ8kY
qlIFZUhhLUx324zTy51b0YL8G8+miaoxiIsifwJt83EAosN5zIRMRCgSKFN60OPBJaa/x/5hXC0Q
yfPwWTC+VnC4zkQIRhDTOwtK6Pv3srGdJDULuCOewo0zB5ZuU3/UeZbn4D1Dh5LxznAYKJwwWlMN
GOpHHa3Ovtkb2WTugrSdfgzzNAnW2bBw4cMjL474IzXM19hjnK9RirMlcsdx8d0fJTRPOQwfyJE+
gL88DGYFRRdAm0J7oJiezVidmA2ZTDaKnOfxqq5cqiE9LBqfju4ogZwvvlaCMK3KS4e1s6tRTpTT
juh9hJD3S7cHCx+JmGf1myLunhTUqBGwWi2XsqYOGTG4cN+vMLQFgQh2JPXDUZtU2a7NNPNzuRuA
iU5nwFnJ0cb622TXsjBDJbmfzRYDri/uRYtGQi0IwzMT0UBd3YFfv9Fn/0rnCjc0o2NNv4anKnXo
th6h3wyjr8f7PgY851kjGAtBVHY20yubszDnoRLfE/Rtpo3Ng6x0sF1PNucvTWmZ6FgL5Q/JbK5W
T6aRNESazzklc4OLf9NGrvc6ZZYDoyTUC/Wqu5BRzjpJsJuT0s1Zv8QJxQ2u5z/QnvC5wUVOU6Bo
mZZHfvVTXBQrlLyr5iaMxzEz2q1N9z3PPIdMSbISLxlRhzW+V3LVWJ0C/J4dhAMOsAymUQkdU2In
gbJaelNWQfqrnQUxHRUGP9gDySY0Byf9eLQqXqLOUDaWIxq2mB/WJryRGGRa7464CYsRZsqZqzT4
/NSm720FPpnFE37hP/Pmr3f/vZAK9qdLkQ3/oJLN1p/7hpPIlYSBUMAQWnPtKMaMMeALMQNeRFZe
aLnLYhto1Yo7CYpjHc05FPO0jpaZbGD0bKqPntEyIzgpQmSkIklr65fk2PYaHS96hIiMC6BmMYZC
mOABlgRyiCQCMqgeDBECeL3buLwkdcy7BjALGF5YVIK/H+L8s8PpjYUmUT5H6cgisBnkpGxNLAgR
qiOid4scCcCSOgtJm2d++jcQrEpHofM7I4VxCVEFkI7sXme8+C6YfcA+KHOaY8mXYR642f1+Xs3/
bKVdmycn+nU+fYtT2W3OeXmIKfE4RKJwhnRZj5udQNK45uSRzawlFOJz6hMAeaBgSjfwi5dml4Gl
T0DWIyW+blSu4UsiZA4BqFm/lc+cEsTMFhmGjLOxbKgVoAInRK6Gjl1L/Y9y5MEC1I3HT8LM1MTh
PDrP71/NoDNPBZoif6gC201vx/Dgqs5vEZ4N2WwcE6kagEdrZOU49INx88wQTdvi848LZ2ZwpkH9
Z05c3a7jxn1fYzhje2Eb72u9j439ET0WSIriyjnOY4EvsiTXh03NgH48mI0QuW29TycBMZAGnlBw
86MqDCRPdMWa4zWtPijN4blsQbbduPh2IVVq0shUORn/jnH2pfK4i8SiTV3plyn1zrum51gl1eov
ttuEFdFfW33X8IHwPOGMwUXDtx/imCXTlhsaHbATHrdErgL4ch07jCb94YMgMUsl0Db/0nbVQMPS
4wwuU/LqeqAO8r/MYXhXxje65bBHToeefsm0tXXSEjk0Li39IusiOgjp4BujR3nTXxmtYIJegvCv
1WEqf3kPEn/93tj/X+lP1UEPd4phF9gcraN+hp3OdUuzqWOrGBo4rKHa+QJwcUe5Q8+WuKkCLFPT
WgDECpemNe5J99EwJ1WBsvN4c3kro+Lf8a3c/xw9jJf+ZLcEFJPMro4DgS1j1TNisU0iK7oPSquF
crgT9h3pNQmLn0Uo8sfkQl3ms6myAgUGHbW6JntGs2B/EdhHZ7QbzeBAXVnlXhFaq29LOHWg2E9E
JLF9BZIfx147K7ZjFCwzChHmjTutGtKAZOpUz9xehkjdfoneWXN94CUqoAMeng386n4sWNhEDwzF
uRLWD9K3H3pB3TQC2AhY+kjyhhbPh8GDi2UIoxrdIWdFVPOCNQY8npqTH5v+ELmMz7wNSWu9FVfB
fwQHr2p+JHlDxgv29gtqjlx0zTk5KH43hrmqxH7XCSZX5/WQDyUU85EgTIfZ6cpvPhIbsJ144Lzm
NRYzoDvpyWJI4903uVCcjVr2C8INOu42ZQOsZvs6E69agNJwzrNJxOph6ZWr3qVRNzYJU1jlU/TZ
t5FPcbStEWymhl5zvu8raCQNcpk+kI5TKGH4/X7Vv4Yt4qFrhEnActpfLfYdAHDDuP56PkdXR69M
u7IzjPSBY9u+ikuGBDZ4d4FhfyLSieyTOmrxPXqZNeVGmJtQGC5oDseZfF9E+hMW2lNUx+7A5nJh
MozhS/y30QwwYAyRXrIIMEuDNm9OXtS4p8cxotCz/C6DRp8rnQ7az9P9H77+SBZbGvtLUDm6c049
LyMgBxhmzh92k5hdq2RQsPz8J/yVzxreLMJ2NpR0lIzasNP77KYChGBOb4CME7UCZ2fY7zoVsuUs
sCpXY8aZ97JUpwV+IDc8Hau9twU8LQbEkcndqcZjBgsP5XEmdJerKRfLNZZFMMf9XnxqSGC8xFj7
UsJbYp9lBJGdY0G1hbLE4DisaVgTId4TEfLxtvON7vjbSaLzZRJQc7oOOh2m2n5EXiS3FPmg2EqM
NtqOdTTeaxgbEsBFVc+2JajIayoYxa1Gsu4uG93PPdcmmi70u4Bh6goe4AyPptVsRzgc8cY2CFiR
5VG4BmLU+8JBkwOEMovAbunethW6GhgOG/CXRZcXAkkG56AFPmeTSGUKaqq/vUunVfVHi7hpDjmp
E7b/4h4/LJp07wtBpi7zDUL3v6WpD72m2waaCdBtK9no0Yr/a8MJRfhuEdpIx3vCdYAJ29bviPoD
Uxcp4aiI9SJeRIqkBjIkXKDE8SDaz1xmXiNFgzDKMvwxgGSaRSKdnMSstfiWuu6txc4xKHLXd/sa
CSLdJtrBRxRWIFry5F9avnP/5c/hO+D43peO6CGowa/dWGBYXLi8lLd13T3q2579Bjlwris50DBL
l4vOVBZQS3T0xxcHueb8qub2T4PkQwQRydDAANb38IKv5bOOr7PzcI9y2fmOxSDsVkbfNBzOwV8A
UNvi8dqekvs8lgLJ07dCw1jSGhw3jo1ba5bu1YqwSUcbLda3/gk9Vz0qHg4Ve4ZaX0uMEJx13QEa
y9TO7RFm3n6rfXafYhiHKGVwIYDvdEQWTEu8AlZhMX89untwnGszlRjdvpHpNtLm5QMq7o6ZNG5/
tyNrKEsv8zM6BNDhlSI8RbYRFq8ArKm6c/lq/ivqce5792G7nm4BguRg9HGAeIo3BC9sn05tbOw5
43hmLkX2Mp2iQe64m9O8hMP5ZKiFz87uheGGL/V1NkBGiVXcJIED2I3evBNhIuncBEGQRABSyKFn
q4UEwo3pEq8Nxad6agRnjm8K7V4q3bolDTWs7cfkpVcBOMWeXDz5eH4hqJtYHFeHDghoD6diI6wG
bxPvt+vqduy+xWUQo9QMWEW1COKGqwfrYctcEq6fy2xrL/I0ya10DYqN7asZM/L4NLuClDqEvVFj
xtwRKZ3dBDCFnzl9CFKqTJW7JXyU2wp3qF9B4kFYRSHjs76gtp5hPMZxfV8/lgKRtyOfarZHyewz
UhtzCeX8cF0/hiYNbsp4t+GXFn0+Dab3DwuJzjC09i/dXOUwl5XgZi4IdZB30kxZUpfY/8Cl85li
WpDB6HEK1UP4J0dRIvEHIqqcgmrJtIuxZ92lpCV72I8/ORgSwOH/PEqfPECsPk6dQN5hQuvElQg5
KeXrpOeJmvl7ZPg0br01fdPqKV7/IT8WO3JOOmn5RWsrJfWFC5i8GQdW78U55MMiS6QpVPW0OPqv
kICPWEbLfTd33FsJsOzakYQha/6KzIhXx6uTJ+3I0Ih0MoOoKCa5O4ZYLuRaq1HKBcWlDg6c1FF9
EnNSNZ2nLJs/5qb1izYkaf2hgjfUe/+sAKZ27XrskPLmqAtlI28SNSpapbc7ZFi1PR9bBm4gr/1G
aH5OJhBi2h0JYpUkbsCgxrnAyOcqQFYMKK2MeiQvQbDzqKlbvUApU78glegjW6r2+rgk8luum072
NEkwY1p4a9bgNn7a4ACi0TLpeQKQpaKb8AGy88Tvnrcx0aC4BIR/PqgIe7+wWuLU2k4TOjk8nzKs
HBSWb6KaBwxz9UrilYwpcxr8H9lgqVgyrWQYg7YFyydsCs8V+l1tCACwaCcqdvEXBqUuQSi9buC+
gO5GeKouDttFRN288R00PstVl/kk9SQwUQOtMqAjgVH4Rpy4pNICGg44VcDVwBCqhI9+Z26L8uP2
4KxAWpjTb986BlxBtz6EeL2Sf+8IXniGX3WI1AYtV2Ix9G0/HSQmiH4sERt3OUeDkAYxN5GcjJwE
w3OKxsuDj/YRj2GORUDdKVhcAOrABXhrefBM+/oKGMR225v+ozxmPKJyRQWmAepgqeBapHF9MbXJ
r4NmZpX97ULcwu4mVLw97ItjMjBTqpCBh1uDUEIH9bqI3ldyV+lCW+4bJBv8B9dolXqIbWa0/sdz
ltw8QNZDZcnIuGGv+ZNTj8JDj1u8fr3q+Mee7eER7YqLcNcwBIIjxb31tPIHVvacC+kRe9uBz8C+
arJnoq02KZpusgtmSY8FBZbA3JCezUCAqklBTWH+7r1SSdOPgib7k5+7XgfR9jTK9uPbhLlVIKjd
aSe1q1M0UqGQnSckzcV5vWpS/pbM8fP9vDGAurVs2cSpNQwwaVZETcYaWO90BO5VP7Vpxpnlz0OE
fFUx1SYuHWChCRxvI+9Ca8cXwcIpmX2JfiBtY2lAsx+275G1QFfPkzR4cND2Fgj4Qx0s66EkUMTK
kHyf7Ueuz+902Msk+l8YjuwxsjGtUma3nCTvUPI1+/234i17Yi3ku5huSct15mwzf3MlY8x/UmYk
pGH+8zssGKEns+6mza/suoVsAKxNI4s+E5uiz6DWPDsqXdxN9q35GgfsauI4VDyn/1IZj01TIQx6
tYYNbHwQc9UI/dLJ7tfLNN8wVXAE2kL2EOTGMIk3dMOBL8WAuh4IqM7vLx7pZrtIFjyHfP5szMQf
cORzR6/XZ9GNJkIPmld4pkpalzO/WzssA84F+3zbIegzHUxoB3/BttfXxu7Csjora9hCJhdRbGHi
Fh4gDcPK4kY8tXL7E+IzRbTXk9FhyoaRfpVJQt+hgQIc5YQ7+A2JT5g341rsm12l74W/YmiYzdsi
sVVBgGGAmiHTM4hx9S/PmP7RREqGc5Ci5k7iJzLYN4/idBfgbJ6mcLz45gY1qSYvEtbOMR23rMEY
lqlqTGkkmnZBJB3kzSLfs84q7U4TxY6LDuFS3NB6Yon9Tu5/dAajCP/4IZgqKHdHcltsuPJvZQdi
7lmQRynYGAVd+2Ow4ahLEYwgjBc+DOsU+C1yLANwJYi8TGJlr41ErT0gqU+G3I+sguUHqTioBw+g
ErRrQJjwfK0PgqltPYCY66gKfa0rciM3avCWBAnCTlAyoOXVM2CKmvvC21sBhWsFZvU9U7NcFAbW
rsPo67/w1Dh79Vatm9uNi0S94EtHLHjISzJQf4va4b9axD8twltC+AphATcc1I/MeerPeLYNH6/2
Hfs9UCLOl5MQ4ffJi0wKiMZW5fZvjjq430nTSBnCa4gk/ig5Dlr7nI7GktCMeMB9s40jddHrDP0s
Mww9TEEhT8ncWqdQ8yIEUl87uOdKIjnHTVH3/lu2No5tD2PuLyZdtRHs0KTXTJWDv/Tp2SZVUgkJ
irJIbz91MotmndZuo0psKk5dn9VmNSaFfUONB7rk8x/7boZDO2wdy8xvn0hYuy4kFsc3Ox4B/Qpc
AIVPWVAoMaS3/hV/5iwYV3NtOWI9faR0HiaNSpRmhISMKKGw1xUeZ+DkX80bkObUE81JQd/3QES/
tjgHMU5+rtmIPWNlF3q0Ac5XYmisI2+GW12qDITSgCWEnhouENvyjUwLWQe69Wor6MiCad08pKAv
N9fCFURM603HXfMNfDnk1qnAZKf6hzTb1NzL9bWW9064cuWn3PwO4XwTBXiVMPoVFGtTDT2Qk84U
vlXCSzuo6ezIRwGY67QVS1V5O8YEMyAQu+ULTE/8AmQJ1RwyfVs+bDrRq9O0pSqHwDl1B/LRgTgN
dK+SZmfqVJON/5+sRXRfrbYKgP0WmGk4gTrk0XstTXzCfx+LSVNhy5wcTasEj3koIweM3gvMmOEy
3BKfE9kNrjgrrOQsLFJGsGLXyTXx2OlfUi0TLWN1gR2fGJbOqfX5RqrKg7WTYluW1Fqthgt+1VZj
w0xfp+d/lU6qVLEABuly0r+DphodTiXZs8dUkn0sMbyFR2pepXFRip2Mop4h1JgESSpx3Oeid4Oc
fmlAHGUDK844oBeBLXRxuD8JjyHtQeXOMxKqPBpBPsvXh7rF6FsjazgkSb6zZgQ8zAzJsZhdgOPV
P+SyX2+10eJWLeuobFKi+xX9pQ3Dl2q/Lr8n8QoZIlcyYpvWMyOVsoGXh3L8UZXVPWanuwMzWjXe
aqoxgd6t7hLKMHoMjD0LF9FgsFb0hNRDfMdxfSiCauRRyg1YKKieYjKmjPML6WHAEbvybf1mPCjE
h6PkueNbQU/XtebVbiCkWTRGny02nVsI3n2s8LLJ1J+9HigrjIifa53QiCBujywtJDIP+U7+UxgT
aSIetQEgWFzBcWCdeY5rE5MHl7NYtInuZ1f5lAFYKuJt0UDQpWml/UuTWO7ZITELM6jkrqcEnif1
fYw6AsW+XIO2ZzvGYrwty2KV/aSelNbV/ihVGRMMhVaRD7On8/gd3YyEBIJoPDW8BykG+sLsRKjA
Y+upuYfBzqetsPIYTMI38musvxDaULci/y/HYciYsp2WwiHJkrLhJTGw7kN4cVDrOPwhjqdaqakd
LNl5nczyGdKtcpL7hozit1lGH8/pzEEndHCNv5Tnw+Z3vEv5kJU22qrsKIgMvZ6krSd8a3jJzLWe
91hlQn5HxBK4d+gk2c7e5kYvaiA2e39wHczKT1PiIZ09zc+YsXfTDiBo35t7vAUHlwbcOkoY6uMb
O73bikJfhh6vCkZRInd3jWdDThyM9RvALDy3sIHaWd346tJWdEKLrXefwovF1qs/+XJTap+PmlTt
hbMeXffoQ/g/62TNpX3uT6nvg2XsNOslsbVpCqLPqiFuxwH7KguE87Y36voenrm4GaXjYW+Ds7D/
dpUQo3ypFFfSPU3rTVT4mldbOZfPLxSHCqyadTV2fezfdnx95zrS9rXo3znWofduC4TLd7wPyDaa
e7/Xd/dA5DGp7Y4CpbSNeOr1983NcNyv1JOCDswdnuiNyFjdM+MDEi9phSmho5NB8onXdMw3zNKI
HNwsUVZ7mp2nUdQWMLG2F+jOyZhUYO6TZB8qqJ4ctld4q2nLfYWd6o8/z/Syp3GeavgKdicUqRAT
Ffm2fddOjXa6kThBSSKu4TgGHz9VYXoa4BkzBA6Tm/rT575844BZEbCKg7pIxoklSteDf4WnC92C
rehLp7YXsPWHx2akIcPoEKEObpbjYE3+fOFtag1acw2NApnzbuXn/O8414MUS5kvtA6FhUuuSnhv
71Mo5z6sYLnSIecs+moDajAgG7bjldSPfbXOZIHBFtukkggtCAaSdEBqqbcYmtA6foxfjQkmSSUZ
gR5EVIP4CXaEydlxvTlXOSKSpX0p66uzceUETR5L27+LlgMVIhe2Q/6qe94TOw7rdipVJQ3qYzel
i8wEfA6bgHXJiVjSQBM4iDyGT4il40du62W1xSfBADf+1dqLP+nPstKyGdgwoZ+1B+QDBYg+DEbh
cNMSgERX4aBbnAwfr6SRK/3X85IM5fieY9GMuFjcXyg93RlOzAnI4oE+b1tJg6PhBUwcsxKD0dMw
ABV3XkrgMCvaxEhH9qW4rFt7FNBLsX4wTWaM5ZxvALipY+FNZQcoO5tGs1OU/0+My38zIDUos3Jy
vsCtX5pFbr0GrVIgvgwCI61xTV3EDoeCn7DDz/N/7Tz9NQ6CaLpavtJzaxjIJ23isA6rkavj2gLA
ta1/t2A2YdQiEFCL/ayNTSpsfmuOh1fPQKKjOV2T8OmypkQIhaaivNxmjP+AHUdLAAE9sFoHYFVn
3OaZITLaRt2cjXdTp8StIihzuvUAmuOxd9R6HZ3waQr/8Quum4hGkVp88W+hlwTowXYXc5pCKmSc
P2BJXDQQ+HBqan9YSFH7BNZ/4j/1wfRRCAtv9TeCgGr2GiHsURKnilFhGlUnMAwe9a87ciFq6Jq1
ED0dhcPcMpvqvlAebmktRIezOo3+2qIPE43aP4XTZOQZGtEFS70GcP74oFv0OYPV9fZEHu0Hy5Ij
eY8LY8p5KMQALu22eBS7i1elvu933LOAw+zWDNiHDhWFatKb+lTU8NOAGfPPMFi/VPveHWM1owWA
Gx7ZZzDYJt6xmVx8Ax8KppCb6CEMh2CC38c5FeT+vOWbyDU0D+wf8Ez28wPWPsA7nusCuYAzxtnr
Ju9R5wYg7pvMph5o2Du5cJDEWTjFEd5zfzkA+xL/jG+JRzMfFJ8xp8lI8QUbZIKRgEZypq8hbuDo
dpBOfbdXxiRuspTXxI9h5vo2OZcYqcxDrYpDiIw8lfa8NM1HdxkNBQG1+OlZcrwEmqHZJMot+H3J
hJWFQ4DaZ9cW2WGIUpZBAgKy+ZVqT4jOIm5AUKQCfrFxhZtCvwCK8fzmgXLyp7Fl+/sIHLN2q8ky
44Yk5vaPMcUua9K3ItU+m+7nYMZ4U18H4IkqsHqG/XQCkQaHLcPJ1y7AUfEe6ENUeqQFAKL7SMRx
a0I/oW8wZzslcb6vzHnI5S21EyzwbcqqovuSjYZfwI8dxfljfZW0DU2fx9rRmmx/g5BhG/LZZlQj
TWTBBw+stIEtx2jpPxgZ5gWQLTxvqBO+XqojEDL2jzYvnV1RBgeFymdZvmTmRpXlsq11A701eyFV
2ErwYveylLeRoOGyriTQ2Cx52j8mBE1ABGZ3NXE3CHpCj4gyFcW9T37NlF4SlBouvTp8CfXTrYgM
Xy9wsnPx9/fQLHi6+H8O74fXS4D8joXaTT8jGum61EqO/aVYoHttfu2ZEQX7iqV7j5DZaRYISKjq
0NLuz80ZCixrRj7t+9tEBrflGk68pj1dkj1gQskDtJwsqwFn9pmlZFBij0yP/slYkRNNDqiA/zVs
IaaBlZF5iVqq+APCvJn8uaRrO3abCzUVSpkrAiuV2ZwEBOuuybgvdoTORL5qeb5uAkz4PnsV9xZq
zN541E1GO1EMBirxhVHFZZG4GqTIrOLq5ozAI4aogjpzHOaNL73Wk42jiE3WifKSPWed02Y6cu7P
93wFJq4iyDghBZT0AHbPOPbbl4prb88DzVOfyiKlP3/O1L0ToLAZGtTjwbrDQX51hmj6v0cMu2bF
0EooH29pEAxydh3pf+/NQjPOjcaT7iomLcK9v/PREaU1E7zRkGLQMTr6kSJMghGrJKojVsCwBNKm
1lQT6zZBr9oawWmwFIH9tqqNboSFO/0+CHrcjOiOUtGrXCZnPrVZax+G2ZZv75eTNqpIrJz03ALv
fNgI4ZckqQ3jwblAo+T4Tb3b3IWcf+TCQqbjEOlPNotTu7wwCvr6uPoGapeJg8ABDiXf5YMjFw9Q
r4PPFtqDZwIM5Yri/LXj5mxRTbY3Q7xh8HvHb0KMrOKBftC2KwI+nvKjBQ6e45hmfrr0EFjB6RTd
VTDInD+vv8HYZJMPCB4l0bW5ZQhr9q80cfdOzRNIwzMcOkssri2LjStwp0bfR/3at+0Gx2jmkiby
kULZxmfF/ZQ1ZVqzd3SmO5ErjRHpnXakZZHInbW1gpWRB8yLgFxMBUwOVoCBbhJqKBLjlj3xEVyG
I0sKHltzQlAh2+S8N41XOu8fnAV9dxHEn6PhZewgLMg2AYaJ60aKUdt0OwkiKGHChWf1tKNuacWP
E/lyavlHVdIHp9GjEQ886ZNDwMAzIKilOioXGhg/clfvutPklwYMXalP6hncyO2syMQL2jpRdWEJ
iTZbc7O4nCoMfDr2o6xTtshtNTToMRzjxjDRXO+nGD7fdmgFsC1x5veCya4DqQn7qK1IlR8OxED2
DNgAMAvB44HVHj+p0iCmZGIDlx7sSYgcLYavstzbiHP1BA3epDlZU+8dJFM/wAq95zDSne9yi6b4
SY/YL+G/Gbui6tip6GUj2pOo5VTNR9OfmIDKxAPNc5ct2N0Tr2Lp63QkH+jpohV+InOzTVslpaCQ
WtkQZGv9iUOG/VBmrjU5I54Vz3tpdzeePWsWb0ErPkgZYxb2efzz0d04UiwC8ug7ftIStAImc5yk
Pp/olubavAl9BgLNvba76WBlL4MGYFBMj2HYKp/I9wUi+EqAJIhrpBYt4ruBGzqfp0VYqIZUdT0w
8ZGg7ogHVJTzW/yMA8Nv4ozgdKMYkte4N1W59IWvFFfuaSAhi1oR9OMwZd4NZN7oKZEgZMGsxNpM
kYzIqpwbUSlTm4wZLBkIfZ2csWOHiq2Ilt88JZuBCgZCxkd98OFDjJFFMazhA8LPV8WL0APhodiG
Arzq2Eg8zjw0dHW4DtDOdrMYa2jAkZ2VPBRt/8qdxAnAY4ZONd9LXnLmuQ/CIDnWZQZzr7jdrosN
awIjLPQmze+4pU4U2yL2uohl3sUb6r6Vur+cdw9nbbJNNPfJBOEUY0NV7v/mpV+lvfHEeEJZtR4r
x//nn80KSPVWiWeIOzMN6BIWMCFJivwVSzNnS543Ce2Z6ngYY4JCXvqFhM76gdDhVOztXjzPhoOh
CxUS2XV2j0wbKx3y7EhJNgbh0lAIOIWmfoX4cuVORbFeAFRnFcOfkQ9NBLFjw/oVCvxk1YOTIHnv
DvEymG/nK90a4bzududQ9Ws7WtrQcfDJ9aAxhpUouA++QzSeZyPyPdmu2wNv/W3neW+70nZBKFbM
v83887IsqBDTXWd5ZC4nqmB1s0Orsca57nL8pMGOSRARJHuscUYA5aM93bKoN4JXBfE0Cm7RxTnO
TfWhSu/5uFsbjEyK0E+KLAEuxmwEEU3H0OXOkdtOorA2Y4ZUZin7ArO1muinRDhi4McLFnalgMCn
LEvlADATpmz/MsFw/qKatSR08Pe5/Y78IAKxNHIs9PXgfTBS8Q31H2rastigvj+zCeSEIolwtmO3
oNlDTjx1VHaP6lLNkGmBceoUNqc3OADoTR68vH7OCYGoNx7yYOoJUwDGC4EICmfgRQRZmHqnRs2s
hYkF+gCSNN4ahTjAXu2nuXS553GbPfNH2gqLPOz9qTVsndOe1SFivE937s4cPsJPNJunSCdHdE6Y
bPOLhLbNqJ1kJ4C+g+PZ05gHEnIr3Q8tWuVlcVBEtwtV2S8KDihL+K5jiFGW1yM1vsh5Dbv5tcRE
9hJmK+bfSfvkl/zl10t+JyvjmpZ5eeQVBru5Xge/YQ/5AHBM+XWnqueMQlJ2vYf8hNnR/B7ICe7i
bPWlELNW8LoGsub4Q2TyD+5kWBSogjmGqHTSh9XNTeTtdVtZKqe9QC4gkrDYVzUCaAVVQ+1kwjnB
1ju/NSaW6HdR+no2JSpVB9zh6OoXZwYWrtq2/quKdlD47t6/NBG0atMJzkyEZeNLJKub707xSDFn
x2vP2WcE+dffYBSijvgzqa+sQIhFgX0o7AnO+6UC4unjGEaLoyUXPj2cBAIira8DKlSjXo1n6I66
ZJCZjZJQ4q5vwRXfGihCFq3uJqbI3sgSPkiaFJ3CrtwuSUK1TdfQ6TggUbrZhENJNhFmwFC8fFH7
J+gGa3iRvk3Lek+139EfE6W9F2b2rXzK8WquAPTZR1wXY7S/ikDMdPqZSqHwiIfuKlPXLoX05zp+
iqdbzeKbxnEVNOwa1UnobtiaU5ITyk7ddCS63NTSMuMsjjbOb8JL/EiQi2fqdwysOWvowXEAOSVY
sQkI8i3vcqjiG8/jrUEzXvmUeQEvCl8S0JdH7KYTh1BZYJpKqEIr2LmV+nXFmlavUISs6UgFFf9J
r121AFYKLf7xQLAZTYh7r5ANC2dxlyw/9LM+XtvFmwySzBap8ZtBy/LkUYonutDDimeki6ksI9vy
tVfy16QugyZdC+BXlYF5DRnSpYxi3njMLaTqAOlMwhDJrdtAarv/wznqfHdV/Gqv7oFzgPfkufn8
Gkr7KkkTGVplYzuejTD19rp/VDwI+VGO6E9zYePnwYfTM5/MVG0i+UhqfgcuoIYqUH/jzyWPPyBf
9N7oMoWsENQsu9sHyO1OHBFlKs3/iDGkiF6z9ELe4ffUytiWhuR7yESWMim0g06XiAGLslPbzxWd
dzWhUBFKYpWoCw5KbPp3C543EcLqR4gBmDJNZEUj29bEngi0KkbrG5ZBlWI1gB361zl3LoByj8Ec
El24XCCJJfSKB7hk7jpLVmfJowefW0C7gqm//908UYJDIxUWwzEJ3lxOryKFd7tqKNIbCk7dpQlE
jjGq+mc0zOYzRL+ykKrnE3mozeygTT7OlwxAu0ztD7tmow6HLdLRpsFPcwUrvynRiUm386tzzHv1
+6BKVC+RFMQtdqAO+YLWQgtkmAqMkl0KdW7PUI3D+A5zhNsCV2fpqnaFTC4wFGT84gFxEmKJXPiC
K7/jt+nNL7Fy9f40oADHFtg/mJaThXntpuPwukdOFj1y38f5I/SV6/FL5IaxfFaNlWW4u2KsxUOz
0luEVNM6n4nJmBdIL7RKqw/MzG2uDysmFgp8Aiv6LX/2TpAH+ISCCugkEF5z824jutzFxVaLvQM7
vWztlUPporCCE5wTFSFHdV0jhEs0VgQhtn6/7RoIbxgMjgJ2lwlzIVSVNSavqa7nOHcaonTCzMl8
LnN/Tfw0XncqxOhNzz3TOhg+P8Ej4myjCffhxv402YYue7CgONk3f5WvPvTzSF3pxT/4z4zcykPu
dluq1T8pzZIrBMOJISh1//sUfOyun/ixENh58Sv+Q+li780zndaJe4gRIpX57GO277YK2mnnqL/F
hrzbsv7mnh1szVu3JhAJxpYmOZapYj25tioZVr2BVGvJXk9sIFBXGR4me1kLXA2g273LBysbfXV/
LANR3IgXZao0O/aFpeD9gP8ZweAFXd0eZAvwvkaE/GSckS5O0dp+4kN/x0TB05KAQllaodF229Ke
vTsMOpwyFcw/BMme8U+eDUGpYKhXJfjp2Pw/NP3V5pe7XJJLX9QHtn+Nuc7FryckUZlOtqDx1jaP
U/K5oA6u7OQQxAkrfpNDGFkb1lkfxqMpX+9LpbT+CtmI2NPCHJu28dnXG9SGHqMnmdLHxYvu2CXq
ViWDTiAv9zV8Qn10Syd5DqM9x9rW0RgK3pkArM/w0yzam2TWgwttO9QsGH9V4fSWW8qdOZ7x9ajO
lpQvfPjKljYfTpN1zYRqiHeQl015yEI0ARt3hhf8gIFkprwfwUIHd7zoOnhq/OchxAuwrSvsKsNq
GOwyNI+6SlxXEZgIfFXUOQnd16dcYJhtHxxaQC+vh3rvF2FEsiYt/lLYn4S732JEIuPM0NPzvEIc
4kViySKuI2Un9qxr7JBphfdRZK+edvXaXgXq++fcf8flJVvi+TwAWdOYre1PvZmgmtbS+Tt/c6BE
ucRDDZ3AMXblCGpG74CGORZXD983FmDdmPbYfx/QCMUDTKuCWrpEenY0LSmyQ6pSFoFiM692kmB/
/jyQU4LMO1LNcEfT+WxVDfM2lt+2pbvzCxJrse2TW7oqsi7GIcJZbrqzzw5HCeI832Cx/qNRGiCA
hyl3unVCuxU3RqIe+M/cojP1bIu4JS//v8X7TI1BcEC3C2j0EpGXzPThzlKwwfAphkvIVw6AM6vw
CNSIgChE3//IEu0l5z7+zAebRVkRGyKavQbPHK3Wrk6NmlJM9HiVyDiVca2t/zfA9weJJPwII6yB
iEcx+NDC80FN9WFThIzekt4VCbLXu3G3Srpew4mUNVev5K83xeGQNVol6q17ILV/MPdTdLLm4f+v
lpZBEr7vXtptG5mPtJHqhOAApKwbvl/NVdSM3VTToNzyukLXv8TlRYfgptZllm0ZkU6NgeflgVsK
GBSHl9VtkbQYQIpEmLpKEKvlB+6HIMAu/+nfDd/g1oGF7NXfBTo0dVPbPK4FTZzLW15baMW7k07q
22jWZmAMaUnnqxkH9k90zftU8O5QlQ0LV6Hmh0abzY7nBd7YdFbYuADTHhjeqYcU7xDlROZd80lJ
A9Kk5JEG46W39f0pDD4D3+IXb97HvSuHdvVQMHrjN6sGTyhrob1ymmt128e9J9c3zC5QG9KEX/yW
/Cio7kjC9dz8PY8SSV/LwACzPdfYAJ6kcBh3oMR4GHQqlXrK0nGJH2IyxI1PJCXALGECpb9LlIRx
PDP/eSg0I0KjvW5v5H76avglBx35JwJUVWAULw3f81ODJpFr5t7h3VZ3+1j8FO2DlGQS6IjhSaRZ
GXHnz+2qUt7364BUk9CEKBt6rwEqyteIfwVrLpQzxo2knlatOTS4UmoZ90dDDUPh7NpN06SiAoFH
LezGFNXNcALVCp7pWjCzLy590f3t6uvESQSOqtGD2PBfqEGPauwwIPWJgsjmKQtwbRxaeWTJWSae
56dktNQwKD88fFO4pFwP1oQyuuvUeYplXAUXjc9n+XwdKHwCASlQzUkF6Ga7c4Q3FAqS7B9unXGs
FxIEsVGtLCUyiLgc8/VdxvD3Re0PCdvjgUOzBDXtdmVbTuzuQckm+GmIAa84UFe9AD6CXC8HovuP
PafAhwnH1tqa1Tw6NsrGQkzA5lMfeEz3ogEBtDSbYezUQ3bi41Hy7+tQJ/oP/77vCZO2gcqXCkjy
2U5gfomriEgUXb8i59SS6NCgL76XDNJya+ARz6Rnq6EodsPXSMDo5BfwkO5aBaTlyX9TYvscWNgc
d8HBopgmoPoOL8UGzHOqj43A34pXSza49qAbchoifXCpfTRDqkVIc+QNDMGBALf9abAoPeVW2+y/
5+Z/qUw6Yd5AqK56YEsVdsh6dBsm/BqlMrWletzSN4Nm+XMPZPWq+RR/sjYJA3ltdlyWlLlZtG7M
qwC3Tx3Gz+vRHPHfpRYjP5C+TCddbh+4eA60H4dvhN0ukoVorjVGn6jqgNFP+gzSl9hBoInqRbBG
A6zXjGXcLVbJrnoxQQRfaFpwCTJHYw3jw/Iq2YErJwENF1oGdRURG7sY9GkxRBCwXzwuaQRQtNKJ
/alwNXSr6pEy8xYqVb5Xq4JBIRKZ3MBESEPuTy8gf2X1B9a4ffxgJUfk4CCxV2Q2ZbVQHPulsPBj
zbX3xfNf5iMFrwKwpCE3xsZy/RIhez+CAOdtI03+hqbyKvp4ZXGplMiXy4EKr0N2y3u7xKgMWASR
vJmFAY5Wu4Dy9wv93nbz7rte5gcfIckXravr/nzva/U7TigX/GpFiSAufrFEUJi/SneqaPMIGoBD
B4r9zhp4JRkZwot8cRvorCp0VuNFEgEOrLX5oM7NEZHz2uahRjTWn1FqGIBBM9Okj4svVbB3l007
qUdiSxTNHaGPXpw7XRRIcw2nbZrOER8CrESpcS25QFXDZAx0A7F3AVJJybo15a5p6Qx3Si2O+Q5u
KqO9+y00gB2oLs7SGiyh6+YtPELiGqOK6jz+zEqbmom8TaYFxNTIqf8zJhNQr3TflY6EkDO9HuaD
nb/URaWvH83iHyJcub/YqlIo1L61d1Iw16FPe3Ldk64sgK7FQZLrPch6vGr2bHqrj393CBsB7xaY
EETLDxf/XiY8PxF0AAT8r8ba4xKfp+O2d0WrzbT4x69JyGNFctO3kMxDoL/tiNyO332fYwsCBpuJ
WCggaUqdnrY7d6N/rCkwwEnOczgcwrM9VZOKgIHgwe0q7t7vMixX7P3ZMOjsBXoK5NKJCNEEA/qo
r39dsmj3Su5UFKmDwOBisqUqT8DocQrdHxuF+Wd68Mrx4g355Aht+azVJ3m5pwAqyJ6cdyR+MC8b
me1L33ke9Rcop/j14oIrVAA0s4URjK5e7XtAhzjIX6cY9tV0uPwlgfvw1pz9UuJ6FRCJuILw7Bj/
Kvv2+rrBmygujiC90iwjoJgbEbkr1wD1eO5diznrw6dVl4yManGEEIzszcTwfjHSvNIfo9WkegLF
CIY4CStH1gq+wDA4E90x34tJVxl+avy3pqH9AjQlvgYRHgLGDY/y7xAYjYmVLlCvByy0fLCjo7YQ
Nbj//Cpq0xhbnuz8Z3Ot9KSnQ9RQaDpTgQys7Bm/9FaPMsEH/T+20YOJkNCkYY1P+t6d7+d9c3Qv
mFOeQKBlFEM7INZJ7icskhbA+vLfLamOlSuyMmN1/gWmMJdCDo8qIeBTfzYN02iy0t/XbTrF9+Hj
jzjavm61IWYx7CnoQpQjLyL1vwcegGwzPHh47r5F7KG0YfEGtc6hADQdA1y/kYlLthJfAo01vdfs
aCGHKKg5dVIDK6PmgLAN/aiJ2uaWeQrwwhtQs+ABs+jrI3Un/d8bKhRaJVIXoRpCFGo/brIWtCAM
2myO9wyZQtRS42YJaHY+pJpLRCRd8dPBcv2aPBqXkBB6XvahnURXPBXlwgGW3PgF06AzXStHvJRT
01rmqgNBcDhO+AdalNjAxJvrbz44S/mEa22XWSQkxjDN8Rxy3sXxQ61Wtk3Fe4eMpmJnxA0xe2Oo
OYW3GAmKxR88HO5BrtBleDkrne6xVac++q/lTxIozmsZ+/XyeQFQY/q8vaO+NUDSeuzzoRdsdu6g
OJbRbmvjntu33eF6an9355PN7xld0D1CKb8RajNIqTuqV5MWs3/osDlJI3Jq8PgyKQ6/f+8VZ40l
bsDFY/rcrjK0OEEe9Qdo8YdC7jmG3+/UzM1YG7pXbuoL4Io0v5CLMwb5H52jk4vhnLqpUvzEShA2
17Fgcd4Q+1U20jphZOvxWS0LzDKWkUCLyYEbsIiNxgUFzRhVnaLZS1FJhS+ZzxIAF0FTW94+FJ2H
lwIwz7gDHRdz4EzUG9xtn1u+aSOxL/jtKfoHSB/U3Y5AbyNLbHmIZt2am74NoHIaAyCq0wQIrLID
qKx3DyWQBqLY+vDYo2sE/ougmPpllwjX3VnpNCeLHXUo+D4J64A8r2zbxUtvPDcAYVH2yqj5Hds1
GqF7Tz4TzEmVl/axL3iu54dTAVJgiWPTQ5pIQVVkNM0t1b5KoE9/AtoP37aVZ95qnApuIuo5kg+V
7hoUk5lqim93T/d/2AacviIvgKRaOxIhy8Rz9M+9UQQeCep5rBx+lKEmiDA4rOPECGP93nnkV25B
FV04lHntEdwm9+m0+Ndvo+T4pjWLz9u/Y7mbSSzlPPqbk0ukoS/RTlX9lDVHfzEbtscvX9hJWHvt
zdkSzdSimuvg6AM1b5G8HX9dAULJhFkztvyVW7CwEDY9Yc6msUP/VAVgMBvA3cPx8YPYEQJwFCKQ
U8Ydw3SxOw/ZsFdHkAVKwvCWdEblgaNSZltoDnuxTm3+WtKZobRrBNi1es/OADTmTT57ZqAJUOjx
O1HyvmETb7JXGfQD4I1TzUsNUnLhj19gsz8nrIB9pF2GpkTDKtU8uA27cyZFhO4cUANz4VBQ8BDr
17f8HSzJgNCswwRC3gz8xeY0lNX5AwVoqPSVRbNNEVnuIvQNlW2+e+wKW2JdJSF0AWuFEOhPhrEu
+P2aURuObsUISl0DuyZamY9yhN7JhyEWKJjvvLW35l4fP0bOBLqkTi2gIoLySgb9XJO81XK5zrHL
RcLNJOWPquGS/bWiEkYVCZwDgBCJpx5dgekayIX5JbSS9Ui0ez03cYw+qrK9/QsuLKUvukzIsloa
bhC+HB7HyvBE0S0NYABgNOM1bGOry0vNKeGWhYURnNM3jtGh58ZHCcSv7l0g1Sg+Xo7Okwe5EG18
Y6htV8Z7WS3AGyPXYz5kjVkbiMelDI0ctHFTr6DEgi4AvWyuFEETePmbQwIMBKonfETSZM1Rv4oJ
YNSpdnG6umBp+GCkKhCTnrlRh/FW0uegU1O7Ka+oE5dundCISifC96yevAuQMEWQz6IBBjUEpwTS
IaZgyyGiKsNgC1+T8Kxlc6UK//X9rnpUiNq/9jcBWykIItLxVVDHkk6hXEVg3uh7rSq8TsGyUQi3
s3Q+xaD52yq0IoC8PPLILEU//jcltwemeIam7Akgzr5FtGP/BFhEoA3CFGoV/hmYmOpakws6BC+o
1nsXMbki87dYcP5MZBn9gn84bSZUSUo7v19sxtTWNH0Q9Xy4UkP2PY2QdZ5cBxcO7szWEeJY6bfV
6eyKp+QkkRVDk7h9HeBeUlcNbDAq9eNthLOUFia71y4btGUnD0CtM3SuOdEF3+esTfOq1RrWKvaD
1/gM6hM2T9sZY1u5rnKHO7tm29+uh3M1HX1fgH4KIjuekxaui7bLSWwwFCbAJ2Ifeh/UYwX82e5p
45S/VbYCpzO5gL2tgzsJZZCo9Iuo41TdRpDe0ouJmU5fuNkcZkZAAZGG1UqjCY6lMVn7a1Cww4JW
ZFelOSOv6py7Lp8bsdCBJRDCa80bJHzdwAtBhpLjejuO3hLfvPSHzVXq6HC0S9WuzlMCar3AppHl
6eC7LKSWOT5/jv2hmRcsP1mjbqr6R2TiQNWTokRnpL8KEAlkYau4iNI+ceJpIETXmRWO9PsqpE5I
+W+oTl8KPDUa/ykqjYeQ2qLYHI1sgDLfvU32DYjaw7MTKWON/8V5OqGqxh1BL3T0wClP4ubet89c
l9DXxGusQGB8/st+tzHzAtC4/fgwweFJj+bL2LSTRMfMdlHSSuxzERYme2L7UQOEZeAyDKWeI//p
2Z3Ftc60RcxNv9ffjOmnr+bQToitj3SeMl5Dik+grzh5Clbz0q3eXGjyYX8KBGtVvcPSz/5MTDqJ
WiYS4CleQcQ/VDd12xiBp/a2fCkGmlH1qg2J+AGyKStT7GN/HtYwCd///j4JlEEZ2p3vWV/nXCTk
s7X9XPJMADiRlxSuFwaNdqX5bf3hhp8qDnjQ16/8+esioLOW17VYiDtmxwsmD65tTdRa3DS+smey
3ViQrhR/rG1CZAopU8ghtvMsg77xtRlzyxT3+PD8verve5e4oOugAzezyPuXPCoW9UPVMCXC4LTa
MxvDS61VNmxslORgotxn9ImbDPd6AVZUVY8IFf4SLByLLuZ77JxP+jfbLIr1pmFqufr4+5wUQe11
hHIsd7Ae0HtzT3SSByG6aCoLdt+A8Ih8pRk9Xl2EOstFzED4RM7DwO3IZI+HWrZzFcf+uMUngY23
KFnqCQ3DqnwBDwjCcC7bbjVrG/KBeHTgS5pMPtcr4o8xG+sHKj56mvy/PY3pZKwJlnx+4o/VPHDH
iqvYRpuZfQipQ1Z9pzgqLPenGHr7BLk/T50aq0/FzX4l9yDoWSvmnFu69aY8kRa0zcapR6dpM6Kw
ahoHMNRfBFh9m0X1W55/kCjWc58SPboTxsbazUwD1yEAkDI9fBOTPwUokTKCOABPPWtptd3sjv/l
W2bu3jkZJ/SLe/0vPK+9KQEUX3yTQ06G8RLusPV/Tk9ILDAokCQEPh3hzi7VGyLi1g2YSojeOIFd
vJZt+HVmNsHwm0sZ6H88iH7i73i3qurSgkwj82GQ9PkS/aPe+VcfknJRBv9Heu0U1iFc0zCCPFip
sEP95KkkbLKrkghPoReTGx388vqkCPskDSXLe10DfL8m79JCZ49L94pSRJtRBoYgRBMlBwRtiDWS
EFATFhJGkOzQteyy87zBgpnHgwmQVspsDX7biok/08ZQJdWRTeOFttSXhIhCga7R6Fke/y16mFKq
f/AEQUKEGmH7v2JrCurK0yo8MEQmoOQ8t2/KGaU8n1xjA1TaQBSuej+7UQU3woknkU8WsV1myw58
TO09MsObVXhB0xSW5iQYODOrfuXss8zHxP3tZEq1KBBAmFdDdR932XE/KBnm1ZP+Q4FcRMJ1rCzh
FOtNzhefF1VJJxmqsAgPduUO+kKDXZzH50BO0NVuBuBlMRwhxxOYq8Pmw7xOsqopQbTZNs0nvzxV
X9/tEM2Vi2dvR89HfmBIm38xXp/iXGRW6EH/lrO+UwDQUZYnZ8LEQkgYB0951yj5kI1UY0Qp+xi9
ZUvjgusxjrw8VQh5ab2bQJPF4e4Bz93nLrusLTOHkxiPkV5tq3+apHalT5cVjpZP44y1C2H+ftbO
pzmDPSokM8q7RBXAe6UdGelFWh+OK1ZGwGAlMNjuZiu60PuZvlAPJb2DnNxlU7kaHvq9LxIIAAgd
yPRi7OfnCMSgdHsKNUvPLqZOQ6Guk4La05pt+78RBHd5tIG2sMwio/8zxZrkWQtjaOsuIyBSTJmM
WRu+WxQ6lHUDtLJGlt6L1u1PiLyYqQj0xFcNy6nj3ZpYz0nbTfTzxVPOGrXEPJMlb9IdMGjlEh9O
AnmaNjSoPpF29xh9yvqWDWNYaVlMnJDsVexeP+szF+qWyr0P9XrGypUUF5YNla9L7zXUyjWCSx1z
vXQWrMFtIRnuoUGCu56+hNj6kWKCgAcjvIB4Z11IO1+MuEAxB4+AVlYKak3e3CvjWVAJ6GGgZbVP
skm0TXLf01Mz3bhbJTB7uwmf91LJ4r2qTJUBSJrirn3jhg+EvuaWWxI/UqWMszMlNWLSvNr8EzlN
4Gi6ac0x4usXEmpIBq51KQw/WQeu+A29xfjM3sxdqnQDE4qT5X4GkzHa6PumgBwhDItHBPK8cQMw
LRlvdFjXS9xNvLLC7XBJTIyZM32QRMZunS4SBitHl6ADR0bqwMLB2UPoIoh22X2eyuEAji2aMPfu
cTb0D1B0miwRoa7eMQBnoXfZ7Mo9eKiwGdK/M6RC+/HQWSbI030cmqc5R/Fmui/o2rKng8wri8SB
EsqC90z9qYxbSRbbh54wh57qYgrnrQzcdxNok9ekrgchv5Dmn/qG5tMU281J91t85RQG5fmN3ddO
AkY9TSXsUJZ6hakBFxduAxRQTELtQekPppd7NBCQv8i48Q7QAtzbpdOG8wODFHcqVempbd/+aHLP
EsUEw/KQKwEdBRvBvexWwcCFpFkN23cgKeOObCOpugvT9kCktNCFJ2ZU5ixFPivc7z5jXu+m9pI0
CSEnwwd0sVT6ezjyRsQNJaFZ7bMK13Gl97iGQEfEjUg3VuiPXMzt6T15nEd7oA3P7bkCBVPJRaxS
RZlSdoX+zxmecv/TodEAHVfVn9AZHrhZI9/IMN0P0sO/wXLYUM6qIyLl0mwfxcGLA1/cC1uB/IQ4
daMf8OJICbiWhfCzKMuqBu0BY+KJ2a5YCU5Jg/9c4hWUjzipeVDWQesq+vQBJS+bmsjM9L0tdBnP
JAcSd54BY9B58/iz7R0mSELn3aUP1VmhtRDH/sUuDRLFsWlHMRDLaz8ezrGIAuy1L52720IgeR0w
BDtlLHHoWfLTj1gumkIyFwxtcYU5VDDKOd8bgZgJd/PbpzzzGo/l0/lkr1EI7yB2Tzke1L6eQvd9
hAIKAQrDbBdxkj36Hz+y8NGK1C3XBEgm1U/tZrQHVMWNXwbJ1ahOo9TMWiX8P5u3jrJRAaS9FHQQ
8Gs8k2dNYPerTGPRDxMbiFijpMPzkOr86Li/35EEK/PgpPRlYOBew0KSbdyR8OOjxwPyDhIjZi2O
RmO1zpjvIH4OwyZvxhwxe9UTw6bv8dm2VIOnc6Q08U4qsb8gZaNEikAaqYSjN9OeIELUpc53xm+q
Vs5JRmIgDK5D611QoMvtQYrNcSjXUGToLyOjkMJZJ4MXTmWLGu08Xed6X58VVGD5Jdcx2KbMI7q9
YlKffRrh/f1ZDU45hFS8r/qG0vUCiRqLH7VSadUTZ7d75hSi7yPWt5NbeLZiEmGV0gxYv7aMYRUn
kDj+tME+w+u4zAPm1YC10Qe2MsKDZ/h3ZzwC4EKpYv9u/fJYZz1nNqG9XncSFaVO9Ok5yjCOeWZM
a5MaPXyYXWv5/yGH4qdlHdIitfIqPix5qsCCta/1Ts/VBAXXQuEbuSJd8KfJJbJ0YNzMZnMBfU7Y
GrKST9zVCoA1KaT4HNw733oyEqDMrCOc6NXMlkA4lPbeTLOTJ61Gi0sDYEScFszFgNlh4J+62MCu
tEOKpuc2E+g8QXhblGJYMsYCu4NdDyXKsyph7Z9Y89LmT+8mLdnntKSFLmU8UppnbCbwXw3L8lqH
DbBWShuc8JpQwuBThf82F9XeZUnROtunsDOTKJO60eC2jmQChzYwLOMI5KcHCNj/iWbPS5IG7ss1
fgpFGhmsS7IUsnCrC299W62zHGlsMIwPJ5DRmnlkmfszP/URmLPHVgL/umOlIMOxpqtj1RL8sckX
B9HWyXmmgXb5NH8IS6CCa4nTh58KnvuUT/IQRL8C2lhqI0phCWHoIL5EfD3Mz0WkGCevawFKhGCI
Tyt5lP893hZ/xvZUe2eOjF+7lQEBdSfSQPpSHfpR2kuks6UZ3pwpb5IQt9FxP1NNZnii03jtbx/6
984jEP0c4wjBQb5TjBwVxm5C6de9WiV6MhRL+NqnDsGDp1mXDBUD2HsgmMy/Rc/BbHAj1ozVap/V
WDmmwoXT2tHskm9M/EXR1iRCnm5+rv+MQQ4UIHvKnGERbVnzDu4Ew5RU0YuG6RInmwkcE928+9XL
i8DHkGC5XnXnUnGfbodDr25MsjeUqsRXXfzNeHgcA+NHsT62ha9uIJTcp6cAxaH7t7SPI3Yycg8o
hAmSUml9skcI+LseaYAXuxVId2cX3xT3Ldyx0o6I1bO7IfZPQ8/A2uC9OLEGebU7V5g0yRWu7vSO
JEK9ORgaiTlr9GHGwmUtsYw/3MFWh7rYeVcUFQjrP+o3LJcR82Chod5gmsQJv5Xmiwl1o9Hu37hy
zTHjzZ4lyH4rJ9y/eTYFdlfjp2H24xNwSxamcLy7dUvRd9S3g9IRqHY2cuGsXoc1xlbBV4GWRy9G
zrhe5TMEHEEAJiRFdlLJhdp12NqnDKJEnWjgc57aO12Pqwt2Ycxk0ebnXUKwHupWyuue1uaD8d9r
Q1dTj75GTjmVimJwfIIZGGpMbm5/VC7Bkyv3rk0dV0sRX2nIpmk2Ja0rD6cIuWlqpZ+2ki/kMTx8
IcUhFiazBPMvv4Bl2WNPlSoBZTyZxzmR3gR2oY70PTJnhKOaaGPwMye8Uwn35e7rUaMAd8idqZ5X
cEr5oDzUSWk7bLBYVgygKZuus2H6TqI1xly5RMIg8JXwIMfu8aO5P9ulicxM9L2DNebWWDE1inG2
Qot9903LAjBW5yl8hWV4wdXsI3kWLkV4PY/G0G2+CW7SArLUs84w4LMM8fTUagbHdycIP+3DTEa8
S+zWrEIkQXcxCWAUBWBYCdCx0n+k4YVL6+u0i4VXoPpcQUeTBlv2sSMMEyBUU4rQ5pYrIhUgf7eY
VVIe64eCNu44P1heEc89+jBe293EyjFR73Qp8DKMD5NZKSY9LaAnGY0vuZMj9j5eDjjn6KI9Zt4b
Z1z/8wKcOxLifAWaXovOTb3cj5RjhRKCCicnGhmT3gP/gz4K7ZFOSq17bO5l5kr2QwJf8e+6yf4Q
GuhISTVqo7+gzKgnuXFleJKMVqsgGxBOSOCnwKaRWcc1CYbG3yA2jG387GC/cp7tLqcYvI8Td8Y2
iIUVgAeJ6TveqDZ6efgXhT5uivuJSejzhJPga2MsQgJXmUBamqQByp36ergmCmfRjBcVkxmQai/4
YpqI705OShLnDSjA/qkZ0k9sFyoc0OKM1ytCt21lzJptiundxJM99sp4ARegneEIFwLCefOdgcTM
ud5Q9QL5B1RT6zcGypw00J5G+b/3JnuAZj7fMd7qAQE9C8w4ONg0pDUBI4h/xn0rY6y9PueEHfgg
0xKKwWhn+MxI8eC32f0giQisBBUjpWqSTMxHBRyez4VEApdOVWRbaT2nhww1qZzk/CIXNbtVbRLt
IJ5ymc+d+s5KYTvWDQ3Ww3ZIo6s0FOzAmAtz3keEk/twylpaXjupZx7takcuyysgdJXwiLpKc6NF
ybD0ppD/JuNV+bvLPp7pIoW0QvVQ2DRDT/rCQ0MBX14LkOvYQhHL/hKV5mnRlhCwm59/zkZRZ5fH
jMINCiFuf64+M9WC57WndVHg+wXkArwy5+F+7EatXugJJ2kvOYyWgOTnAGEjd6RK1DUJTpi9oBc3
ac3CxYvXE4mQTkMXtK57aUDiQZ6FXnbLJ3YjGqo8VdnkoU73UjZYc0pkFsP8d2Lsosj3225OenNe
qBoh+dc2jU3mcM025LynKIKlo3sbgZf1/lk2TgsL4GcYq+Ow4VCg7ciOBdYMicYfOuE3nZPbjbC4
NisSV3ycNWMWRpztlJEMQjyxf0qCZFZEqTbPr4Zzw4iOSA5jL5rZZC3V5iXA4jEU1pmIWc8hhS3V
+1/8rXTjrs/hZcawq0RhXXFIorzqC3MDcSS44GInJG/Kf7JBO3EPyG4BZ3nw3rYUEd8D7P7FOMOT
CitU+MZMFTsiKqTnxyg2vp12VkUF5yQ3nwYTx2kS7xjB83jTIcWlaGb0KwzbxEbCCSdVEzAXEEMt
1JEMbkRlDfeO0GlAYOFdo3+S9bcITGwivt7/ux6LlR54ajjeRs2duFxdeVARn5/ocXVxKcaI1NRe
STnU/rR7FkRjQu5C48FDALKiJJ2P4RonyhdD0AUvt9UCJ+XSzoYkzibSmCaE7O8NC/oMn9kEtVkS
/xlkghdlbuSXEIBg0HSe+iXUZjJDChhr2FxeXKw8XvbrTtuw0gnv0R3H76FalBELLWWY3IyF1odZ
xw2jcuJofiz6DgO+YE2KaaAjxKuGfqerklzFgdyWZqHVKDWldJwpIoBItpbSG8vTNI3ANgvDJ/IV
MI8uGSQChvWXSZHBVM7JGGlNvA9C78Hn/Y9Jx7AW7pwxUs1w3aoAD/eKfkqzR3sy2H/yhM40Lf+r
0NmG4fpaMd9DDf3X0tMtBK2iFlSWeVUh01avvHrneybktBuqA65Hz8pdbbTgsMgLcjeWmhlDVN8L
RcXiuB/zpXzWBSRkrxzHpMfXZs2Ycr76uxcnM3gkQ/Bxu2BQ2lo2U2Qm2tRqMZFtIFzRwIYdMHil
JuCjtlOUBpo6yBwsrpf8Z3nPvGWxtTZ2M9P4qidqZJ1E1n63KOoDBaEmxhOvyXpqthkH+G3gV/+x
sTSBtsW5QQOv4T/RB6NhtVaaVqXJ5w3Scubhi6mdz22B4utTc/hJewS3e5boNP+GMlooAm0pUU64
lrjNmI9eAOW8o9MM4X3tk07COeMAZZVsFxor7UfPV0T10vXPoNqxF7En1USCZeeCK3ZrDCKUZLm+
s1517TUO/V1obdp+RR44XKSRRxCUJXrqrbCrF5TPw9BW/aqN7Fpi+3iC68JaA9BbAZigbbsFgCI4
Na+faGtbWntbtzU0l8ppkBcu+tSRh9dn6eio69hz8j2QCBDV35/5Z+e6hmAV3DgorO691Dl0Q4tF
seZlGEzfWLFLqmsdqK9gLGFfMgoUgnx3/EU8nV74BlNxzJF6cIxh+Q6Ojx9QVM89GrbnIAeNmxdY
F0I7q8mgy8V6A+rPwtz1xHNAUIsD2fqI6aH5vjkhMn0dRmaJDHQgekQTAxQ1pPfnpyLl6pofLc1N
Y8j0qLjZk+K68r+oRrlmjEOCLnYKVVrjAUtTvEMzjMJS144Mfh4GHMIKS7AD4h8Pfk1AY0+ryVy/
kEM+Wk1lyRh+QgIsJ6kzlqzqw2/+opj/tFzLpcW3PJ/Ircm5gGll7VLwH5ECHUB+z5sLVv0+hRq9
5+Sz6O4OxdHEkEyqjykjf8Dyb9OPvmDGxZA7LqoWO/xKjXSkdmcAxoDHBrmE6vhQuPVBsZLYtM4A
jdH++RP9aM9woOw3uuECxzsM2mzJdbVW1rMfA6EckKTGWIFWBl4zPHP4w+Dd2l3bCXVus2FhgOhq
xGNgIyzi/Pl92Zg/Npk6bGHoTF1hF+nMg+SBEJik2Si+yBwvlH5JzSRx6E+8CooRlSvPZHeyKcqF
dVcSTtBUVLSPZizomHGx/ThyMtIf6VJ+uQz1j6ozhGZYc6dZOGN2VRA9KW6NViBt9gwBk5h3gHbM
C+MkukGlYgEq+m59hxVt1xur/eL6Z2uW7nx4VoR9ajlr9yKuWOAJsaIt3wd4RzCbTw5vVzyobKQR
HKlDfi4W1x7FInwYDdZ1SDxNkqCuKzSMLTjg/I2ySmtLK1LtQJ22CKFP0wSwSvGSlFuprCeKUZyq
+0ZPAZRzM46PEA6h6xxhJvcNpYNGPNy/onM6m3ah+JuR3rd1mUKIYrEQFrpnSDTsiQY0DvcewaLJ
KIIAGhKBBlhB/ykZw+lRwxLIq6IE9/0cXoJsKhb3/pxWUGZn7opHptiRljsHCUAdW0w3lyyKATZC
92sTmB71Hdp0NigHSRm4KwrzEbWPEwx9e+vHze4ZmaDNb7AvMJiJsLQAqVmKw45cnbUBhir3HlXM
ACKX9CnFXIj9uba0OVv7EaDG/pWKBh/eo2ljrjp4C/jYt85XK0/fiiBg7XdctsyQrXW5AoLO5l9N
1rO6iQvU7MxinikOjX91GrhxU+AEZe6ZwGFXfgf7DIRgOIhE4O6eNwcq8ySheY5cmHZoDSCzb4lL
PhkLUPQM9dMmUbByjRneO0VlDys53WKutskeQNGbNFj8peJtod7NBobpgqGHKsOUwJazEowcUiqJ
qNiITQpHQwnp4XvuKexCBL/UihPQSY3Tu/SlP6QQ9cxP+JmfvMN0QVpOyk15Zb2BEaKMv8w4bQTP
Qg/16SAfYbmZEPMuVyriNBrS5w7rtVqWANQ2wjQWa9eQG/rWxvCiKcxwkztbTTdhbrrDHmjoWOHU
UuSkJJxlUZynBpA6kF+RlE6aUfji7cYUdbSRzqBlo4etSlWQ6Kl3FKnHEwpD4tSawcT5fuvna8iQ
l64JS11zBiEhdHhGAFmRI4M22Cwvsv6Nvc50ovscImErAT3NYvYQS2aNUTFM64JDbA0/PhjT5NMI
JJKJ+jfVsAr3PNkZn5oxJI7PkkOsbYjjSSYhXSfrP2XmnLOBGUyGUGJSQFaOIWgs6J4gulj11PHR
J7SkizfsccMmqBtGBu7kbARDPVWrQ+k1Aj1RbTcEuWvhLwtSz/TOd0pNX5BUrT93w6faRspuUQbu
5anTEYRpbAlEl3mzzwDJeCFFs0s0MK1blj2oew7eCq0ZA6HtLgePFpeL8/bHbjJBQd3oN7FRE0OO
xFhVpHiZvsm9F/WsJvawL/l3KasLgzZm7TMgmW0UAI80uyaTQPtBUy8si6J4txK5snHuoAhwoufy
EJrq8HT6zbBy4abDXtK1jeQ8roAipJ80hGk1lVFZV8xzUkxZn8XlGHN0ppjGJAuUZWGseO5NUGnw
ojpp23oQPod4wQt+vJguOsLhiHvZ8aDJzDYWFwHrMOZ6i48GZvVqaPHtqCgD9fPC0W31hE9qRjaM
+bRgS8p/lcwbyoV2efxZKPbNDD78lAJBQP1rSyNuTrHGE8obLqezFrkpycciNdadwPAOSLxg65dH
prLK0nqpyPW7TZzO6wumSlI2AoE7J37vVaJtZo/uMXCx/WNromAFezpC5682uQwy9IJDCnBLmLfS
LHnOic5UD9e/suuE0QJlt5hS1cg+GDM+qIhgQ7+hiLmEEZanVGhhz3J1kHfJFKkJH30CcDNkg0IX
st9TVa9zp/0fNUzCEFkXNoCRGA8WLAnG/IiIsiKoN4SQ/mCrp/g9eHR1I2De9ISyVHWpSBGPKFa4
FxYcshl2XbOA/rA6JHROArz7kUI8asfefhLra0mzEWbEm1qqAGP0JE9snepelWSq3vCu2Sgx7QG1
X1avGQAF3SpJjGW09JYwtJEwz/wLngk4uXR7Ovja72E9PdMB4PxeS4YjNTCrGMp5GpY/9AOt+6Qo
4Pki6RZvxu8nxg8742t4TSLs4O+KOcLOkbnt83wLNEduEFuZFzjvNNoyB+q+9AWZKl/iWmXnors0
5pWSbjVp7v+IKZWuydtuQaeu2ptKmTcJr/oS9fPFKIKg9MPQIVV0/Gx2Pm6GHEOZOikssk1CdQ1k
6c0PAz6r3uV1zApjk/XmOYAETwE4ihIXpLpPzSsQv67AkIw8sh7ZSBB2wAO0zAnTfg/8i2YKcjFJ
IKAxLfPZILFnOdbR3+1SXu2WyNC0T0Y6TxkxCHGZL+6sJqZHAHpF5XAhJ+Nlpcx10UIz7w/4QgKA
imCorHKFWvlfyRUbJWCCkqKYH3Wae6LSCse0MDC8UkKS65tRrjA4Gc3DPrb2+jD931b5Mk3Af6gl
Bwk8djOI6UvcccAomcAFlN+mL6evEIxuyKeHodI4VWAhvGUl4kgskzn4nwHk+iAR1H3AIX5ZD/RS
aqmcBgARTMjdDszAf2rRrFJCXHGlrNqy9fXSUKAXpJwuf0gwYOcGWCbPwHbKh2SKlNwIi11VLyyI
SWiBhKaeZ1yRyxWBx8gqgo0hZ1XZUB6Ithhqe+gQNGFVnkPbjpulqxbVWTFajCj/cWrGk6kqhCji
ODw3EsVShWnBV4qyiQRKCz0J8mma6KLlNW5blRysytS7eaMQl4+2GpfWWwcXJYZK7TT792gppSpu
y21vHJ24Xj+15v5lTq0Cafy2SJi8DAAoyyM0L0cBtR71On4WftFZqRvYMwy3Cplawvfaf145V4WO
dMKvgopNW3AJ4rg2oK9qmQahCPFTszVqZSqTJ70i0taLLgW7yntU9hIw9oYhPpvw2sivFEN5Oiif
sfgItnEMm/GgFyb68v2uK2Z6nww3eFNX0zbBOHysm60nO9iekitrDpzKQ5Zk55KYw1+Jw4K4+zYC
3CVZVRXKVCXTRyt4m7ZrdmktW0KFUdFGRb9L0cJJZNLJhIHqaJIySMLKD7MBFldrfl/yvupLsayO
vqieE9C/BNVDhtDeM0Z7eltr6CWCfeXNvD7e5BN73oWuukQzbJ2R78sk3v+hDDipjrsdiu+1Cnt1
ey49D30qmL1bMyiVE+7q+TyNxh+I9dh95cLxGTZ91/OCGaJFOSq38Qd6hw805qhlpLfa3dr94P4K
Ef8yEJbc9Fa64psRivZOqphzAzwPDAc1pqitKdslRRwRUtL1LKHMnXxIv7SSNYikiOI0rdwT62m7
bBbh0C6uZs+WuIzcekgMqh1EM4f99DDg92U0NPNmo4N4l+77T/IbeCKYvAv6uMHkJ45Qm217Rjnc
0M49BfesapW5FS9qRRhgnOe5/7ugdti1ZHuaMSU/Co2C6gSH8RwS4YbFg+/mPapHwg7xBMNY8DBu
+pYDLpcz95f8ZhsOQBrE4Ieui9u//bHD5gPIU7ru29VsuQ+OAgQ08JdiTNmBG5sDsKMCy6sUB8Wl
1g1ajYuven94O4xqame4R72MULVuST+RxLZymwSCWbYOtGi6hGXGQ2NDXxordYRwo81aFk/ekVPs
bQzEEQTP9Fpt/rwEKKHMpDhVijukCmUJW38db7/OqevHPGUo0wfva0YR1lf/QIe1z3FnBJKbSs/x
JPXh5PouGefMah3ivoPjK88ijawRv3JQhGA2rR1hHH3EM+JsGzgEXDmGfVsqTPfTUvYmuM/hWcMI
f/5caW8LKqvDBj/DTSpnL4cyFHSfHN4vDfKhrvpnEwCjEkDipuSqLWIlyKWHG9hizFmcIaAWOZxw
7wmdU4Krn8h9D3PoBhVg5kckL2iVVYjwFQxaSdRkW1hzQ5O85fD3/9VnLLnrKuBQnaU+fXll0MoB
UOp+uDqWinomE2/o5Wfymz3Mac6YNdmXtciPikoLMsfpFYco9q+SCrSWsiCvKcqwBymNMPhFaY1k
pDqnHrTyVMduylWzi79pE/BEd3HqqasAFrXjwGoNAS4URdkg3nrva7eLDA06OrwHkljWAlemi3e0
RRBce0ynY2YdhfTvrrLW/C6TGbDTqTNpgAKkGPYY2RQ4CyJ/zizgI5Gx+Uyr64ymq5A7Tsq0u2HN
nJlcc2cQguobfSTcMFW6FAn+v9z3xKoGryzd4WbJ3vKxg8fAta6MO6n3yOMNXUmljvuxV4vBNYI6
ztpv1Wr3VaJI9xbUMg2CmftK7HRx//bSGW/sAafkJk2UUl8T9jipRektoxj7e1j5rWt8Bh353fn+
MJTHtpxK9tdydrqHQFK9lKXYoo7QKIN0fvRV3Jbrfx6hVpuwF82vy0w5F+AQINKYpMgTJtiuUG8f
PUvD/fSDQIp7sXU5HgKkFY3a9W422o3Xf7aZF2ghLTGc1cAfMem/PlcWOF2dZv2NgYsW06O56V85
mDpqOSnI1153Dudm2Pe67glr7WZurXtHzuapLqdsOe544mADrD3sHS4/JVt9M4a4jPLMil9D4uBc
de826VZqFVn+DEitG+RD8w+DXJjznsg4IJHXM129ub9wzECJV07vKEquW0nXB6vk55jwTOXCjs+b
34475x/PCkI3vj2RYnN15Q3ek3QjyY9+2X/FIzC5RCALFJQ2mundm6uAFvzXLFSLgI4uEGOBW0z0
wFxGmInoCuZvhgnh/XDu3kF/Dtli0ubyNPatZcsnPvo0WqGy2v1AF7pmHpXuGVXIod6IAh81CY6J
t4fIMmgKz3nk8D7ZDjXMxlsQeZeMM79YE7x/M7p2765dGvEOazBZZDw53xZESmyPe1Pc4zEZC3Lr
1SmElHXKB+vo3/S9uQO2e2qtwsEqL7gY+PVtyRHWfp1eXr984x5CpSikuHQR5ZbbY7T7WmwHpvUw
8fLj2sle5tREJwS3XGXgFJIT17+aHlPo98PeZmoOWSm90I8Ii+pUkRHJWt4Rs6kHPP6pUEY/hqRq
YkPzu/4mmyNOYsyK2NkBjdfUZZSkIpLOgf8YPMjntmAprvvqZaBCa7qVEWQzSTF8jmDc6llrcFjD
aorCXuaqe+bRDBdgGBf5yhOZ1Clo42ADhaX1wsBlyWNnMt0Kl+NrGwZVweRqiuQfeZWKE1itRYcm
6ZMtemY7M/CY0V26/zW3KAuMsIPCefMkDQKQzzhGLSmEqPptXvaww60Vvp3ba5ZAZqf3e2lDrOwn
xuE2aqLyLoLnXOOoHiJhJYPmI54IP0x4DjISAUf8LV4XFoiUbSy/ECxbazP08nSHhJKiB3xoZWqy
63Qd59RkiSgKshhbaV6PkhknnSWD1AIoPQaBToBDj6+CBrbjFr93WtHdVPkOZ0s6IPUzG9fzxba6
zDua4ZbLqVjvFnYDE2kmN1gua9YCSd02SsjYTUje1TmZXfd0uGsZv2j70aqWSbqVQvanylQPYifQ
ruAamtjDG3bAv2YRc10ZNK8HMqLbfNPiAqh0OvXISz8ko0S23arfiUXqw02RsUZlgzPg3dJuh43C
IOUAqzhoF9RAhVR5akKxK8diuUvoRH4Ti4M1cBH4gyMCDIkt1bAHCW5feyP/T4qXyQujcBfG8O8g
i82YJMQRkcrza+nNLR3SlIq1PmkSOFClxrLWCjel29moZmk9PVRLqob3SKH8MQgFjN3ygxeoa/sv
f1sdlgCEz4NsGaX7I25CafrJOyBQeKfxvGDUHBVGIIxSQb16tbW5uD0aRK6mwtM7/i694MaXK2ZX
xW8DSBKL/V4pTscGgT0NnU5KeLJYdNt2FdXF1qcXaTIr4ZEg9nNNkTnEdpa0Bc/nOXK1Wkui3bbC
RRWGTlDrmZIu97gCgRjwchUcoqIQf2/FgpTrZ1nmheArn2bdVrlLw01+o5IhQZcPJU+ah5A1x7hB
Pr6hngBjqimaMMu5ALGZg04clf2UIT0ZC/xhu6jTqapo7xx6HKUSzhGyS/6V4U0rS9KwJgZ0S+vX
1nW5oeY0KcV7xlckRgiAm36AVjfaCYwPDLENGT4nf7C0odKL3aYMQbEBtNJGwOFIkyfw9s3dEVU4
y/JCtcHBmDYxvkKGHyLgjQXQTZAYNUVLYNUGjI5cQkMcVue78afduy25HUkRbQs6sRidqM+2kNCo
x/+8SdHYiJcGx1sRsAFG/8lpNumyVPKdwlkhaDgZxf+GZel7QGwzLAmiPpIoIC88hdOIQkgDTIZ+
ZnPwY9WmrO7YDS1o6+mqKJYqtbh66NSVxSK8Yg72icXgkK55l8F7M7sybPvfo9j1RFT4MuaTZ0Hl
cxWbgO2D4aYf0IYdJz3UYD1BFgnuJWA3bHpj491BXK0IiEzQ3FthBMq+Zqju8YKKOi0gJb8cHMcn
zLtfLHejEAPlqexBAiXUy6/WiXt3PFNaxxZXv3Zq+GMiHEf+NGPHUAfPTEnem6gk0IgSoMN6TwDF
vB1k4/ZHWhRU2pu0DA6cmTyu6F8jFwB6o6xf47gEIS75rE9D+AVaPVPFNE4TBZwZFMuxV0PuPAKl
5sQCW4QBuMyy9GPz6RybeOXVeiFPqqm86LSG2Zl32XkqQlyTc/g9q9Uzt8NqFd5mFauEXv6LbvUS
0QFP1a9KZmiv0D25XwKD2g6++iOs3uoX4k9HOcQRPfp+kVjUfh22J7MacZ019txVuTSYAy80XF8a
wyrNGp1WGvhsRc99VSl40LtmF2Rj1+85Kvjh1LstwKZ3t0BM11AXbWOOo0LzrgPB5WIsyzoAVAp9
ON6bk48h2tTFi16r++97q+smDHQTLEyfpMD6juRx7P2mwFAbxtfARuVlLsy4maqTC7iwsVhuW8y0
dEocsV5GUyzbqYQ1q4vSFtfaiquZZWFg0QQSOPmI1dJezZGbdCeA1wALqUasfP66kpfa9QmLwqBL
UcO0vtDoQ77pHUHZYAYANod28PqspIgLIoInki21tPGID6BsnCDUql0ZcZ6Bb4ZBEmtsfg7cWrYy
bkD8U25nEYYm0N/oow9uFcya/KXq7BWDxf1acnjifIV3UhXBb2q+kFhFsWSlrJ6CdHp4iBu5Wqwd
oAfvQD1ejoVcxlUu2NjDZeikAa2+1VlpifBfgqtB6+ngtMJ/rUZ1OB4fCQ8AN+kBLeXfiMEocnjH
j7rXNZQA3OGxecAZSXiLTlodYMt/OtSBnzJKYiOYUaMt46rYhS+u2yZdCFS8Suq7rvTp4W0CbI23
Qpav0lyWnUSUXamVdi2YHYT87PMs6snqwpExpXJSBH+Z8wDwA1hIJZWoY374DGHZ5TWHKg/5pPsL
wjGZ3RPsLYO0fw10mAClOa57xHZp/v69I/HejF8uDt2LKMsomHAH1HcoNaYUQBhsWArg2m3x9fio
WHtuIEpj7JXS4f4C8kORYX44j35Tsk0zWCn4r6P5DGWagTCrAscTmuI6fbFCYKzDnSy5eluB1ujA
QrRqEpEKlTXTZScgjjGgQ9lGBITWAqUp1d2kyHaBvj+CoMTTVQB9ocKQFrJUpu5HwNKwpT0hTFUt
yixP6rqbNqFr9D7F08Qh1O/r951OpihpBZhYMzMbof63uH+129pNDZ0VesuL6aX/aV1YTZC+npRx
RGEAKJLI4CMiH8gDmfip42H8ymHPwEncjFsja+2ELfXE8l5ga2QXvNmfZTftS6/uMdioshHM4y2v
O1REV7kGN97pJiHtmZGt5Ml7xuo7dx7OGYIL7C3NjKeDOmjxtt+rD6iEDGyl7tVQpuLbymYvj0Mv
SOU9d56Ans61A0aZvo2oh9cwxEB+o2T65OBkY7OORyzP1T8NKnS8cDOyzMB5+rclame5eF1dde+J
rpUxGuLpEkQg0ZKPB7ihwEYR+rAIDwy9LsKtZv3K5uNYO9ToKAZmdNZ/EcGbAVCr5Mu/afX6cL9f
GBCbxXIdVt7D20kcTRvZ/6oTf3keSyvd059LgPp0QBrRu5FXJ2FdJ81igud/F1e12ypR6I7FUUJF
z7OevY9j9WoS7i7olXY5NSZRLXp0KU6sdBHbJORvFT+vVgyJGJ/Gqhq0A+AUr3FqF504Bud08npf
Wm7cJ+Ho0jfM8D3/S/mnyeojs8x3Zm/a/4MNgeI6Hcx3RDacnEMzmVrPymFPNNkDzRvJfdfNWhED
eqH5X8sJQ6r43Bif8/tvw2LfWWWFN4sTRN4Q/x8xl6hmyr/8klEaYbAIPkr9GgiTtRQ1k+U8Sz6n
N0dU1Om0mkVd5R0Sq8xIKL4ZZMAyTiyeWW95e4dG4MlRM/qGTksZzYVNM8Y8nQBwPFFliE7pfx0C
ctgK9f63nMYQPP7d6DMRES66lJzECvC6gHpzpJU23zClNIA0OHLQOUFCA88x1nTNGnLenqmZmHas
mKVMkl8ZuhRWEiKGbwlc8javaA8PzQF1FCWs5FHaGAEd1Vzx2flkOEzVmaZFQgez79LN8GOl0065
OIppX7p8jhrvu8d/EwCjVP7W2EODY6WLtMm45qkSFzknbKRzrFg+Ssi3JMEUnIHIc/cpSd4TGq+t
TQ4OKjYIYq/3moDBtJbRudtZks6kXz9zLb50RVpxW4BiZV4c2xunU5YKGpHyyGwsJPJpfo3VNeRL
KDqaWkNLD0cst9UhGSyy7lSDp+UHrt2BzlR5uMpoe0ciQIriCO+uXPzCN10Ovb1Ms+jNdcZoWjuu
WKZw4+bM/mxj06RSJ6dcFetq87P0CEoCJ2J6ocTsHymlmaieSBtf/bR0B6wthjaPZeBfQs6/ndk5
rwjRiUuK2R2uhdv2L2vm7FaHtngfy1rKUkb5Qa2/0yvrAAfevG2g0URW/kKkoGdf/Nkouls8+F4w
ypWm3HTLdDa4ZtZumbNNvltJSaC4b2bcdNkOmlbYG7gebjF+/qwsYAPa9Yfx0klG4VrwH9jqn+3G
gqHiU4NjlkUTHdfT62IdDYAnPsTymmfpA1jlv+7UHeFHaLx4cF0YMZS+5HQHcfFpS/fnoXQmBB8n
wNxyfXyBjlInjI1cdRpKUuzEUIBqdNyMFFbdI+KAxkVdKghIqKcebnsyc72uFfEmAWhOssqZRDe7
eMI1BD60DCjRifD9OU22ZXrSoPn1QpBkr6dKS1mSQNM/n8puqjYzixI2qRxTVqIBiZ478wDpQWE+
u1yIfI9dScJjXrZPGaS/ISdE2yIsQyEvmEbv4lWetHLDK4yry+jp77cFx7kkS49efYrw47rLSFNl
qhfO+MSdZK+v5yEFkaYswXAvYVS+ruDSsOYUKk6A8bFjAcwOQakz6XSm6dBgMfqwB9zRLHuwBU4/
ktmgdOfxDxfRvofxeKZTBqUZcv7zRjUQ+icZWY+HaK7B2q2YIIR2RK02UH5/O+wPxiWMN0V4ho40
7AnjwYZofXDlkPPhHzfjnIRymhz5QDs1E2rGYXtt6yXO/KwR9ZQIGR55dR4nJuS7Lm6p8QrwWigZ
UmHRikL+DTY28FPUtpdxrquqJ2wq7tiM4GXSfv+FZXGBSdz5hLbZVjHOIOcLxE+JUtWtQMtqGqsd
VPB6r2fek+SrE2yFwhnrU1x/2JxML85h8KQ2o62Bd6XIlJZCUeMkTR7nncriM1Lfh60SsmXUUl9U
JegaC8rg8l6PghDefFsGlXCkSpFIyWtSv0InBiuSw950dU+MkqziBUeX1CdiEkRHEgKdlTMPRCg+
8eJj26LwZ617DbeNsMBcIwLW/JR+RtIYKQ2UVeL/kmjmV6iBEpcSs6B9TV/l588UdL6m3gotJ58j
o+HLFBH1EFm58aZDoDrO53430zGjYbTwJtk69wfWWF6pDjzCr819fH2jtj2GYsoSvE6j+zMoEkzp
nIrlP48a4QVHXtvnTdbzcQFhjpHtFez2SzWyDmH5EP33RIpmSsvGg+4wmkXVQUKh9yYhLhkaUDXV
DZpW5nzLB4C7dwbdYpT7gc9ErfGWzCcHd78ToB42+FbUKSwp6RJU+UVaXFoJV1dVkQf/Zi/U9a7D
JnQ2F7UpGKwKRsInoQEULlRlJA0FnTArHIFrU4nhUffz17XLqdfLSx7YOzJOehG5Z41L3JwVF17h
mnmyTh7M6Wlt3gidjv66ky8/MSzRB8N9eKlPA2A/yb3QD63d8ZuL4u5l37ggj6PB6WOhfGHKf0FT
8khLuLigZu5gq3zlKmuT5UQSB0nD1jm3Etg/tI2fc3s7v13YHrmh/6s0xYHGXjoaxCGcl6yxlgru
arL6zyS+2YoDfmjmbSe0r98c4ex7ijw2psAmEhcfEiUaxtTTg1mbCFkZlbM8o1HNmBlIA7A2YPJl
0zMXCsHBRbKHlhbYf4IvFxGkwyT4Lwg9zhlmMdHLhV1lLlQ0sQpQxP7v3aP8/SI1LrLD/6aD7Vf7
zQ5db+bw1VKq3FZA1AGsmy5QcQ9pPqrEV4htejT3+0imSBvXxkcyNewB/y3kCEr82/+AWClF3nt3
nMtSJQw26+T4M1cPz95Ckgh9g4GGjtt40Sj6yZeo+9UA6+T4hD5gyDiJAD9e6tZM5zJ+GnccfbHf
ytBUBHT9dhgB9IC5stF13niVU5419n9DfTohAMPzJkDd4/1N88V4hQBa+D/1A/+Hd6F+7EhzRjmb
/egddtDpfUrZW1lgZ/mgO4nkZeLaolR1DUYZ984vLZOkXf1Vz+uurA8G/bsROgLLRX5AnVS8vmU6
ytZYvg8jJOHNvydgicbZtMiGkWtB9q7EIvkbjK3oJsph68S5s+rUfveCU61IepJAwjF+g/rPC/XA
wClF+bUiTh4IjONcLtQsxck6N3ytuCz/Q+CQKj4cgxfbh01UI+nZ163wTAv6l5Q1hZ6Q4j4HK11h
A3T/dZX6xfn62Oacy7vilDBpaaxkA1fBaJ8pKIHLGs35EwosXSgv57KA+5ZQgl2QqcnnZsyBGO9z
MBcHyugJu2xoneT8cJbJ8iA00s+DitvQrsBXCqvtsvD5c07JSihE8JMO95l3N53ugIXV4T2kiTiI
2mNfk2E0b1mrIee2EZcNg5Pl9X1F9m9nE65LDm1jhKVuyPxv1mp/FNCDq7blMm2gpXvSZmq6Hs1W
FYC1FMs3I2Nqj3nltd8ZQbyuLnmxhUrfF4gbAJQSBBe0QAHoF+ht5EQd3C0G2DAZEoCm8hBRvJs9
2GWFwpIMRaoXi6xGt2vTilwSTGcYfZ+BB16fQT2qcTF6D2fLTHy+MEMzz0DcgSHdA99/VtypaU//
YLE0WNNrJYP0qcXhwmwLwRuOvYGUvM00fdSTAHuqzV6L9C4wW2tJ1jHlZNw2jdZR2OfgM4Qvwbhx
Y8LNwFf0FBczxl2VxEzJZeEVcJTlRPI+qpjyx7WEd50dUcbEQcdse+2ujJ7nWZpwrC8YKaJu6vyx
CMCZC5xpR67AbI0nN5RZoc8Ve2q+bKfv86H3eloscqnZ1+go9prIaln/hSR/3VqB3nysdEwnRV77
LGasBmYgrnulPQhwXI5qYt2ctlyAi3RUDOMK2TqUIad/tqw/8Zq/+OJvD808pZO62qCODh5KZH6N
VKS+qQ55BQa/86wdbcETlHuSy2MNZhuKvWMuLnGp+2ndo+fRJvDq/YDzv3lBvUfriu01bHGJHOVu
Wh1tIpFd56OrestnSlFmXLXqVhOslL7rEjGXoGUMf3hogP+KPhPCWd3B3p+GaSRN3J4zXolSSbGG
723dCOcRvZyFbYQJw/y83tstBbJtyw2v2iRD+JCcUlWzPmxzMUW98vnWnGb6L6epIY++XZOF0I3r
NVA/WK8B2xX3j0+Ndn/ZAprPUihERmXHxg+GRFTgASLI+6+t+0dv2bv3riz+A4ILO5f6+8VbP0Zl
y4DSxbzuSY2CkvlN0hgsGZ013oW+vGT56IoFNNuEEF/O3GefJpyNPnVYgACUxzrxN/57EoiS8fgm
/mdR92IY07wk/PnbSTOG3yzZT5ZqZPc8DJ3tVpIAAlua6RLvMGlFV2qSKInzEggodMz0tktHZuKw
4/TlR067FHL3OA+Q9tIVY63HYx+/Rfq+lwe22tJPr8u17evG/lVgfScdlKfqbC+p1O+TZAgZHXC8
Xwla7zO10V2jBGM8b8yu5c1ZimxtUl+cIrj6UYpK4obYT2ebYdP+YZRiaGni6a2WBwbmhGcEZVdL
OuvQBL+C84u6ZWAI+5qb0wussq+2baJG95ll5lpWvbAQyQvcPC6z1IqXHooo6SE+Zf4E1wFy/2Hy
Tn+sRc2S8QnnvYFw6KWmz4sGzys+rx56NtBzt1UBlBvUXATjFGdo7FVqzaMCkmJUV6LTXvP10xJn
vb9rCEI0yt7NKQ2U1M2783uJPwMhgGLCrtYGngeZKsos93zKYs8xZ8SUzpd66Q8rRsVHq63MkaxR
GTEpsHeOJMrnFfOl1BPkUe9iuYGfMDa7B5lbuw1tccZhBjoq1ax75Fxs+qy8O7BIb8XF/KXV5+kH
cj60uAZp+yF2NS0d9QnWHD6IwFFDxZipC8OwKVooA8636tPRd0TS7B8gAcjbd9tv0Mh4stLz74+j
N+UwhibADaNEnOyxbLTxCmOMPoJ9bpwtTThFcqW8dxVp8reIcS0tGmgUeixGAwwfyQ/2WMVbfOot
wJGwPwLTfuepoexp4PrZWwEKb7AhkzVZMksRYoLtaPUxVKMo9TBLBWr4cfEcd9bB5fcqkhdehMKs
F7jMK8jYQIWFFkMvWhBD3aWpFO9Vi4EnwsMRa5tyuvu4vT21+kqqHgrvnlA8GYwLEF9vUdLmzMHo
fTAZJQ2R8uR5BfJsue3zwfHjZ+vypPEY3fVGTVy2ImgdrxeOynBwUItIsFEsEHXhppyB4HTHaejH
t0e5uC6l0c7toHZMKrEVCejCzh3uVLiJh1/UZnn5rIuYanQq/Yk4AagtO/MT3A+JSwZNLvx8bdiC
xuv3Sf8VRn4XM0q097nMBU5McAPCM0W2drPjBjDIPKxD0dvOSnoW04SM5JXSxjsEFShXWquuuS1g
g94IZ3cbOqMohwop2mrIfY7r1mrtjwtbdR+WrDGGG3TFt1GVHzn1ishbnKZ91ws0DISO+UtJkG+T
oLhoIfffVVFSdRisvHPqYJONrURvRcdYksa/V2U3yQrshjdsZ2Dnb/eBhhk1ZXAS+YAMaXZJOYBb
CHmNu+ui3xdUN6xxWfU0cOLNbqGRuWtKBaTrnMoSrO/hkUUSfvXssr37dZzCvQ8jXDbRVz9h86yw
w/hNcrJ6PKZ7W/VI9fEpJHi0JkGik1SFxJDgTOaXBZkR10HE7cuszBc5za8qGaAF32EwG1UaNXO3
uf3y4FdlBM4mN2uhXhyJYalvKivWfbskTseXNQuiBhGao3j6rvmj0foyUZgaVm6UYwgK585SWCWz
8a3XW7fN2WZxRTLaqsOr0TJqI+uL8IgVHnCXCUq30yFlR3bZgo/wz5Ze3TVJLZl5oDxGGZFJtLQH
HPOZ3y5i5vqynXe/mJT7cVAYPm9pAH0KF7Dlz2gGZrH7jS7KWvljFTaB/0n4J02NWLzMhmPsU3cC
LXShBMLgQV+UXKFFMcBanf8oPvISp1cuWIp4PqVbYk0ttAFpRopobAqZeG5rncf+Hc2vNBDdql1g
kXzftMzIn+XIp5KouNwrQsqj7W4SDM6y38renCLBplPSS36qDwAcJz4iSpZEMJAurHoTh1HkfHLg
N9S2vRoGOV8TiKGQwFSazawXoEFrEK894tlgcmk2XHy3UXP7ZXbpsnJcvbgAZZ2JU2EuzorTP7bL
QUoWfIOYkVXW8pQX9N5c2bu5vnvWwzLbFPiC3k1g9wOu1WJfUMe3/qLkMo08VEGMZGPWtRpyby1+
+wu4yriUqEuDfc5PfngliLaQVU3jx0rePPoLMVA76/ZSOP5NsMvn5YBQLHEhO+rmj3/2SHSTnNHA
0h1uDucE2SGWZUekFug4+B8jD2YDoJQ0mp6mUl7kHK2+TTyxd3TFp5iUUJzBNkDH0xo6YhllC6H3
jRQ9mRjIxTJHzpsaFMvOnxS8djNinxh//b0Z5ki28I/++VWSUwuHhOdKKJRVBuhfTV/flBlcq7rO
PrZbo3JR5SXMhcSEUJuFn2KXXzQAIYds/V5BYvi2GgbR7AWissMrBp/pyO0hiloWL3XJWw87WfJ+
qYNljN9jvZ91MiduGKNWeFb1p7H0mKCne/KaZQjImaVpLgi6TOHppbVk+ROcqpyhdkegyx4pN9RQ
TUwYhEYHwtOeqvTOiyAuFLmZqW7181iRqYuAFx2ruB1+9nxoRtoqTTp+vM1h9lunhykaW7RaCNVy
n6iehAU2sBXnV/6dfaCjTtSyF5c3A47vLCZBMqdxacMKjP4TJeZgpo0xMe6bQ3IBL/0iz/uHg+fv
w/OEDdFmuU/FLojmJCa5wCNKhQ5krkJf98270HWP42D4ymOFiWrQuYCkpL8YMidrKOhRFywghmK7
oy/LarPsPntvQTg1iG8jQXLt8yGQZE3dunuhOv49gMX9DFykZTtb9BGUJav4XYZoWgtVwE2xljHj
HV4up0neo6Hnp/1IjmS8EhvyS9Tb0kLede+sT9Fzq6ofe1dtNGwpjtFscypmYoq9Hdemn6q/qutv
tAUiqbrH/tErIMqLTb7M3dy2csc8M+eSFH6RYFgKTVIuUU1dnxKm4c12T28zl2h2SSaa8TN77/O6
8GDOTMkNC+PYTp9GzcRpqsCN7A1+mMaGd1zq28rgCHnlv3boUAWKIYNEkTr6nUCBQpengpyas8rv
QpVT3W5Vc4UIllW8I1RdxmDlf16nNtxUtt0pFTv7fAyyQN3XMloTFJTCvazublOs2pcG/pqQPsFH
4F8X76KbQOSIpS789oWM4YFgqlnmq1uBLF26G4gws2eAFPGIVq7z+MKGcItqhkcDemwQP4MZg2m9
OgHBZb4piTDWwTQgT4ALXrvPbS1Hp2vnd7YllM8sGrzWuedf9Vjk+50HrIvff2aM9GyxbjJifbwO
r5xALPwUL+US5TSmNbS3JWDBInS8Tz3CVUumyQFPh3e7bVoZ0Q80RrGVVgCCWFCtARrhLCr5li/t
dUAi4fQbGsajI64T5vlBq1SqN4N7Hy1gQJ55cgEreOcxaBpq+8mpfcq1ZMxyDS+3LJ3h5MHGF6S/
pAhIUobNpYIm62V641N8InK6OECor0vKAvFG4LB5SonA6cUBJsFBKw7UtkKntajMvm0bNxRzFLiV
dFQKdq7dnbisAjr0t9EDmI7CcjRcjreQBZWJDEePji5worvNpffRd1aP4lbt7Iq43u1ZEsHQLzvH
1QKZ1n4ZQnt7pxKWgxMOiqdMHP7rt/wKtd1VZDMEjktFtf3wTdxkueowP/1lVYAMMNC24aTHXuRC
Hn0i+EOv1qLZ0jvNfEkhZ6LApSOPu/TO6k2k7ZraCR9co5GIFFosp+gYyz6b5KJxdFi4k+xyIqmF
eyyvmMStWuK1ZaOjxBwMXrZIx/h/x35pl1nejDlcqnrX2D1DkNS0eMJvzX4hcqNkTkUw7VaOzVRp
8KRG9X2AZcDF6KQppYGzCFLYQI9NIDB15fwO6YQF3npHnxTzPZygE/Pc2iuVrTvBbuwCxzoPPXlp
a1OHRplwIX3iWTYnfjbNg3nSRcWocMPV4G5JV7MUWpLYVTgnHWevP2BN/LjgT54YZPUc2T86G2Ml
YE/3NRJmpxc7cJvghoIUNErPZ/U5z/ojs3XRRj1MMf9zmMqbIvWiDfnhSxF0JegLgXZQcE4TCscc
/E34tetjL0Co35eDRXZdTKs3L2JSjr0PO0nLCpMY+iTb+PYHOp3LA3dqEwjw8BvJNFzFuRYVILfH
bLjmycp2ceAxYJDlpMaXUM0FMxYcQCEvdHFubX4VaU6kISoLZMH57pZQLRU5k9yKhm4+BJRSKUyl
BC6/QYELjU0BXI4R22PWcqiD2UUujNWOmRQFWv7VSf80fYkF9mb4K8UEOyY5CphqqcfEgcjfe/mK
NArE9nD1ZM0NVGJSEpOEc8h9nQ/CPcq1345PQkH4J5cVkWNcGWFyNuYnd7qwfemwj/s8AmCuCz5/
UbWzaptcN0+ts+IImh4NNx9CbnqFvDVJYmj10ks/FyTz8Ql8f5otZSWP2/gkMfrjxxr3Djzo6Ven
rE3RDyAiObyG4+OuRxbaojTtTI7S0PYWOTTAvizqQzBOlN+z0rl3HlY3v60EyVl+ZMmKdwou1WUy
4owj6kke7GaBsj5PvQ3gvqzCJPVmpulUeM5WsGEWDAbCIugoBZ2xrX6uZ0/6SBfxmIYygn5GLXeB
uEkVCuyYiBajPYfBXp1b6mEeWQiprYd7TWMX7D4YQvBz62JHAV+ojn/73QVji2FfIX5Kyl8yCsXK
RzaWUkHgFAfqHSoWoLq1Sw4IBFGEOJzqpYUVxPCj9g0J8FqtzcLgmIlpYjdQNr5Qb4KwYu/zMk+9
GLt/pxdp5JURI76ZkZ3wN5e/QSTTcuKPv6mLzR+WNY1JBD0GVEfO0HkYPojO0XgVG8nPOHCN5vAI
pR8DmyIzwOgVR+SGjEDHgPPL6wGtEKxx2riuZoeTcSVzgTrrKWspedv9eqHtCLPICc9g5FtoEJ8r
Cp7kT26ikEDQVNRVWezM3SNm918cXlBI40qwcpxHprOlk+ah/3vUO4fQ507V+6i0kiFhgUXKvp7Y
zEFsq6FiXaYyk15yJnZWzyF5OXaQG/fL8pIDrfnWOHEMjdk+ORBr+zZBAstRTcmHGcjgPKEBU2Mt
2QvOK2/RAqDSjSzpmOKMjXwiVVuJkbjD+NnXJhFmWt3Oca5WPP1CU7AjBR7HcNAr135fQgZHTUdr
spN6uVAdzujg8HG8zpZVNkgQktZABEovTDF7Ld3vpPE+71LNuXaFdIuzy3+Y6MbuZol/S67hCuFT
kVKZo0X78ljMECJYoegXv8K/vdBpC5KnzoIYNPP2gTHvbQFDxo2oW9wxre5Zsw/WIjLphRKo/iND
VWhpXTh0oJvO19N7F0k0/+PwSBBys17I5MW5zNfcUWSnit9JGqywIkP5tLCRFVGAXcizVaL/QABW
7Y5TwXXWYrNLZdG/hepRpBGMycUMhDaM21sZYcqZYTHvgj6kAR7xjHQMgSQBLTMSYdGgQN/k53Ao
xnOifzSlrGygaWLgLz6K+DdoHIrltQsTvCEsSUcCo+QjP36RYePrT94gAvGGcszRagrOLdBVl54i
FJYyduUe8xgdsTJ+SKIppubXkidxoyQA68NDBB+p6mMPv2mjhkJkohzWMYQ0BipveChpbEXye329
GEJgXvEXCzK+p67Eqi2p2JELYRgk0xpHgpJeVyybgsPAtkjT+E3idniDYJMUkor1pSTSQARLEPry
SFTZ+Hew3qZBZ+3IZ8sjHOAhSfU0J5dIPRt/Q0mTV8Jz0Q2vGfUiDqb6jR4KgNwnWm0ElpT5wUlA
GOHF9MClAeqgidfYXn1DBIQtS0FytLdZgb2tpxWg3WM3oROeZ7iVEEoqvsIe9naMLuHjYr1qv9v+
G4B33IXEIJ8BLeHCdCSEW9XJLZEjM+tqjYo1+/tm8cOMEjTez+hdWSZXoHj8XYYHnkCp/JYtzNaO
qWHU/IAo0JBFl9M6OdZaDmci2qOgLZ6dL/x1tgTZc3JrbAOJagZWrQm3Dy4O2OPjJ/R2hiqOpShT
PbCdN+yIYESRMrED36Xy5GH2RnoarFzCgd6CTAT18qVoXSRCx2+NzhZX4DcVKjJNU+VwW/FapE1l
+7cKdXEZFnjW9o+UxNWrjmZGIbMXVDyEd9CBSKOWZ4n1oZg7oZFvyZkCcAc8O906AztZy1vAGdjQ
mvECgZV5Kf1kkuGQ1kNmENVxgrZZiQVugS0eoKF8XXge72TCv/CmZDW0msQo7n0luq0X680oZS2o
RzHjAgo29IVYnBHb1UrUEMSygT2omPv6TcT3BMuIjsVMSu2MOltgtoQOeJqgzUM4hqMkody1gGFL
cVF2zy/wA36QyrpAjyNz388awevoIgki1v9PkzYA9UAI1//EQ473aaGVkWi/+a11xTX5nRxC0gz6
SxIQDfoSF+blz2MWNG6bZwlRg+oJ3btz9+8IFbcI92E3yCC6Z9klo2YheA2mWEozIjDFPTvV0Je2
HeUGVx0LJXrF1irPm7xSG4crhhk5v/CEoW/Sxmf1Yxnfr5qin7x9zOqxN0yrorXU3ZIh+zdoWkKu
MzaFhz8RBmNbDwwI7Ja7UwAYqHwjmJi0/e2CSkpTSC8UGRR39oiC6xafckuVo+2xLrmJzHOfSlUG
wfD6cMePZ9omW0219ShnHQk3y1Yv6H4jXg7ZwYFnLLzYynz9yzsyBZaGjo6pHwGQOwfdaBHCej3e
YID2wVefknmFPDmsHCGm3ILkDMRF0/6mkD3qHARdvzGBhNAcFrTqzQSKqMpi/sgvZtswHZiyyfUz
uB2jwoB7hPASVsSoZ3KjEgtCaGIcBm5s3V1EQXzCd7EzEgrqP0sjbq4CgF0XTKL/sNe3/QmYBdpa
6Co5t1RTW3LhBv+O2kyPPsH8ECR90ewKGIiar9az04hs4PRY9nGXmHSFZyGfCnhjyRfoyiQXaSuf
HsuDZIw/4ydPd8eD2GFNntlJSyM+51uefV09bkfuP38OZdPofy63aEZu5LN+EdFWG8xFry7eGxis
kueZ+WOhP3okOVcTUJ4YJRsYoKtQIdEYpC5a2USld+lGIMGSPozGAY+EqZQsiYTFn9TtrcAryRD8
ZdX5NZg97YGni6EK0RA44I0kSjPFvVAWHZY99cOQQMu2u79KVjh2cvEX7/FfkaSLawN3GWDfhaCa
Lqchq+fX4zw2yxhfZ8Oxxy5lUHItk/4+S0TpLLZatgIJrtM7LnI6sln29TAO6e5QZvh0GHzQemJv
U3TFajCRoc4tKWEC0rHRxe5QE1h0EgJUc1YIF83jplgt3f0Aox4YIgbUbq9AhVQwtQVUZlkQUv/e
4QtpYTATUr2o1kJ6G8764gFycVxPEOSUP7J4VHW+70jyhvAZTwY9Z+7NwSrq9G5ldI5OKyVoMj5v
S1BFq9o8F0h6k0liCLxe3vnVv90sYkf8+IKmGK8bURfhJk6zeXSdUzdfzujOT6vKRUopTOPKEKnB
g/BR6jzma1i2KR1yXWVnzS0olLpyRaYOEuqm/YcT/X00UB/uhYG5EkDCWfMpYDpeBI+liUv20SbF
YGaC0AUMtUuO8BtDJGxEVR8psB3jEqVs72iIH3siJ57y/uoYN6AB/W7yZ5AqvDmDwKUmhzx0rvWD
lIxCZIq6yx93Np17/hMCDuGK+57VHepfW566JqQcJfamy+prDxcurMwDR8Y6EmahdhZTSxLc6iOs
qua/9mkEVa9D3+LI4UxrSdYTGXT4XdBcvUFMGJ7uFTEjxjEmuSXT/rzrb9i3bocwwLEOsi1ZwJzE
5t6V6IEEpDqOBX3+NgBCYPSgqDWxld8DKc3dt1NROpXLNLbj410Y/FnwSEBILq3bY0sfy9t+87/B
pgHEqGvESICd9ScsJaaZ0XA+YpywMg70nH4jiNLh8IwPlccyhgLe3+e5a8vkRpVEOYmAFxRiGtcL
XCCZWH5L1xNm9w+SACJfnwrSXbZcdRDdhNLyqRvIZExBpzOtMSp7d+0lINpC0mFmuwKr/Ju+7nwt
6fXYHAy29v9eExCx3vpm2mffpc9hw6xBSPoc6xVuDey9uLq6fLT2nGxulgQzE8HZDeath0OCAZr9
gbtmAkyGiYspPhczvs7aBT7zgIcRHS2vPsdSuCyZrsDhgXkcB7B4lT6YZhoNojW5d3Fh8AkzLbUt
cr5C7UPQAnSVSDT/fvzWZD8oB2qHuZW5BsP7od1bpJVeaxDYjE8P/JNgiK0AWgY1x7zFxx60tgIT
U+ICiYyD8qOtMooWuFDJ48CbIkqgfMuiUU9BGnR6YkLgQyFAiRAuDFNiw4lre+UK6AIZpF3DpHdU
oafExeeUZecmIpWPB84EGShvizAFIZTbp6VXg/NAcZZEr21nwZmkFkvqYS6/AENzJgRctIWItEH2
5OAK7mYCVAN7Z0OYKSN0dEzEl7f+cSezM69lAUWSlQn3qxZdD5FgEqd4+fQvPoYpvchwUNsaqEpa
amKeJZdrKDvrw6otFBHMaTJi8XY027mjUN1tLgnI+8Bg+r10E/MYknTecXIuNpLn1LVQ0VKSqxHo
TmIhJS5Gq0Xx7pMFQSDtXXdQzoVks1F6M9Te0BmdOzlHrn/ck+QSqgo81WKJ2O5elzzzUY+ZYxrB
pBbIb9N9A6npWZvOyQJdfgChYc+xYZ298KksSKXl1S2d1qEhaIvwlt/3mgRFZnZDBTMVIbzoDpXO
3aRp0B3KImrsSM+0qS5MRxaIKXCPALbJhHFEpWjwCNvE4P2QDzw0gMWoquiufO/nk5WghCbjb7i/
35IkM7NN8wVEQT1Heqap8b+ZT8nz1zrwdNgbQ3X+ATPYdMGGFuo0qIu47ewOPsCdcq+iQYYzQDar
lTpbdZPXZGESgVI6E8mJhFXqWoauGviLgjNwjgLaf/KArot3QA5+A81Wv59GNcO+TL3u5GRmYgtP
DKh0WPK/3EKHjL/Q5xtIXBk1pgaQm8gr6mIbjW3mO2OlTk4GSdRR4LUAVI/MIAq2cDd24JgMzQD+
aap96OqcnaNKB0WcPg498ZE9VD+KHuyJiuOkesPy3sV+MmxEXHMEJNFlvau9o676yaiklVQn51JU
VYba6kEuWssxULthpl0g8rAKgixn9q6LRqBqkwAtsn6ELoBxNehaec1GuLPWpmdN6IFHT08AaS1y
45qSeVFNugrG1CEEnvODCiCumsm6eQugPr819rKuTPL5FIfegD9k5zdLM00GRaXISoUd0Rn76PIh
9YKyr5i905x67w0KKfsZ+HXDyAmQL7ry6NUb+faFdKpBiTaisoIa9pdm4g2Z8lkLMPjpBhMWsVbv
VFd19vDhRFQ1MUPEq2gthZNWaYizW8ISTHrdtep0HOW1OxmSastl1AwbL79SdSHxILnb9zbQLOyW
MbRb3xMoYljhN9SVxDAXcSSg52Zy3Oh3UuvhCpE8Dl87IxGhwty+F/rfwYNcXlbjCWCyG8TeyBFk
BNV6GHNpTSLEFM2fRXMiOwzc7FcvceBiztLLUlZ1Ugrt1vV/JcEsC0aMEpObNri1Nr/Hll5m0BTp
hooXoFIQuvoB7Ye+hBMMenEZ1C42UVwUnKC5+9OBdTI7/LrgTLQuywPh0lVCfxL/c/OrCdrQ14g9
+0oEA42ZF/sEQ/pk9w7BavHj4bXx3E8aYp2jMyhDUqulqeZUrPqMrCERLU+f3LCY76XKC6hB43Yh
sWrp3Jy424SXwGnnLXaJwlhDfjjBnazd4mDG+H1wTZl4lBAJsjqFTdwzYpdXGyv4sxuZyne9GwUd
Fnc+nLQQUmQj9a1d74EueDtLZzW0jvgacrXwHWGH9En442gqIcOGFdCyiWPrCQ0g2g/niqKa3fkk
/5PI4idVOzy5nxjK9TZyzAf5m/uo41u8SWNDBw+iui+1Yxz+0uCJ/jZZIwEZoiw6aSqp2Mg6tNDI
z/ozkaFPcO43Ujy/4b6LpVuF7yHCWMPI+NRWdtL7+qdTmK8Cs7FmOMJcLXXkUkwjWSecbmctIciD
i6SRQRy+liJPrezeN+oRZBYLZL6I1euqnH0jfr3SUSRL68Uj+98xKzzHcZNH/DdQO+ePwAwgnUI+
aWwySy1woZGgQ0EP5vgDIrHwT08WlS/jhXlgv1MjYD0wg5NFXmQAZnR0HPMgC8oAbUYlE/hKsTPX
ON4Qz0yRTFFXJHdgE3cyJHsl/+NG14g9k9eO8n1mnoxTvxTSsIswGMY9LBG4sJaRLjrdsYa+YCYu
VfZ5vvNpMEVjEYGB+1lMXtoE5CsUCbWU7bTOTxVwIQlOGFDSeAku4NH2Yov8XhnhNhNscDMuxFzh
V6hrBi2TXnBVjRrNMRTLYaJrnMMyk1nkGa0wZJZdoLEF5gHMl/3xe/TqUUdiyH5WONvN3SwSjbPc
9X6yPpbGNGvFHbQ3tHyDd/3x9yQJcv2c6UtRXTrgmiX390RdNweq1Lgc/sGgIRbLiO23aJp3qNmr
iFhes/xbfE2OtXMrbdQkwgp77UVeAMIisT9jEBXtYKU/XdVYFeHPZjJs505iLAqQWD0dXm8AFOQP
k36nQdZXcN1q6hPh4SpS3o0btPDp1y0HR0tMY0LjKpGeukYdFT03JOQwDEho9jtqRoBXCCpCuaYL
JJfvMocgSErXtnsRDdgJTomZTsCVh1mhaEmNPKbF9xeZo+syrniKNT5LjJOmed/m7g9c2b3FCdtP
jBYdJYr0L4GfMccqwqxTeGVwJyyXKTXJNZWFH1mBYITMXLlLaPtCkjw6vu9Rc9WUq4/2MpMg7QGO
IBd+4ljNR8GI1LvFit6FNLNnfgjh9bc7Qn4a3GpNoxn6xXKBgksWW4nd0oao5LTI5cyAJcmWjeUv
ChoiBWoqsJMGVp5EPgHxoffxlkNJLwrGL5r57cAQEzXdsPZkSYfqBE5EZD6FkZcOLB9oFYAZCdCL
8OovtSUUy5ZXitAvT+Mvbfgpw95nUnLLmSk+Ewanbz3lXmC01gDsMlxoXvkyJ1ihAQVXV3R3/wqH
/GT2bD0dYD0cN1SPaCw15wM/X/3PYfBF+wmICtbfhY8bb3AYWSRfEfuFSp3gkR7yQSG2Y796zDKo
sIK2U3Aqr7r2oyL+pJdY228j8xwBBLwn3n9iTGmjGPBm2YDr4o8/681HOt7QB9X0t9Lpq4YdNtk6
G1O/bCHJdW7rrXbXh1hZlr9NVkgvt2lOuKFq47NvUshTJEV4fJRmssHrSUI14bgIkSwjhvuP+aS0
22w7Y/uVjhCWwRQGwAaWli4T3Wz4AdWK8JEb+fON3V9pmQQnEQPb9PMnRdxV2gBKktyHxN2CHXzm
KpgMxHkIW9GJ1qBp85Zr47c3OqZJtEQYL6egmPRhS5cUbn/3ZaEmXlZDoftvnpbKzBY/7Mmz9zje
igH5gxxH4P7ZlULHjWpDXZqKuk+WQNEaTl2yAG52GkDITnShsFmrmVUadxVjFfEe4QiXdOOiVl8b
609eiRsCnnJGhgM7pbNsWWJt7fm/SUGsHmgloPs3FdeW+pnzs+66aEp/kawRaMOHUO15buIDeAcx
Jie9gIGUauA1s6iZ5jlHgTcFGGkaGW4J7h/VWtAdwTIaXMmHW85c5sWPPMDZrXyH97bBb9igVpqJ
Bz/c7ptNcz4oOekQF90Hn1wR2t/mRfknqGbVGZoKZa/P+XaygfZjyeAVcmVhRwk94kJTGGvjrZiP
Wc3yS+0aFlHiPhE+tpq3aUHu1N1dCDfYEX0ZrK48w9U6ER3xONlkQg9bcU0nID/oeWWljorWhGI2
hGWlr9TKuTdiIvoeNZ7yXH3LivlkCaJC9RvUStfDicob6am57r22KdbAJSEmuz88tjdii7s7nFUe
N8yseW36HhRF+Fk0YVmMzjA/IjEKBlb9vxF/4Ybl9BrvIFOMyzzBFm7KYF+m2jcSUJu7Mp8mYP7N
gREkMvL5CVj060/9IRQu9IQM/ZWxV38QWpkyJYKeGemIE8X8ymW+J7C9NrO8fSN+PWn85X7JGMgo
XvD/LrtkOaQpnnh+Z3EmtJdJq3uhP4vxlWB270yM9qJ/RhHCARR+91O6Q5U11IQkawOsUbVtHpzx
a6YkDO8FpJzwu/G6forUYBfHHjck/RdjVBzQ4/qTKpKOmxc02Kt88PsYI/YnEnJDYmcCs35LAupc
aslUsB4hdmYaFgZo2d4PehcZ+QEW5szzECvtJuE+9xJN+nodaBy+wQO0dCDcO3R9MtpBCwU7SqR+
mjkGRLvd5XGQn/tGn5tMZs9BSVi1RPI5g26dVQ1luIG8Kf84olCzXuxPgIAFxS/+ot4jWk+VnKS+
3NXoe7GaixQY1pkf4CUXSDOSEt2FfS9WJzj2XVBhqzqMPtkiacbjLh5nc3FGm7Fur4hKr393iwQn
rFWyIqrjQBa1FGmahtZJm+YvsSaC/x02raBjX62bZ6KaMZ6Qq3P3oGbLGZs6h4jbXh/QMPIcDYDh
LopAZVBf6+RBEZ4a9ErIT5GwSZGnXUm2gerNOXjdC4a4GnLZrqUTMGSwH2bDFKGJKpzsvI3ZYW9A
rVLX4XQdhzH8CkXh5w209PaP7uTKTAqTyhEI8vvmJ7UqQOH4bynXepwqfy8sti898Aq0HxeAR87i
VUoXCU06lgBG6kxm0eE1g0sXshgjuvF0iVW+H1ic+68oJqutNFgWJ7dYD7dVo9YlmDbpmgWzntTo
qjYrybcP8R3PisJw4Bzr8GkrY9DQQllOoXQQnx2eQffTHz5OCzwHOAphkzqfm8od0GAs2whofXQx
XoJt7RmvvDQHAN0qi08sC2QnNa28rnlAaGi/rJmm3iwa93at3PM3zOl/TVsewMTgpraq0XpTOurv
GMTwoXicf2hU531kX6qI95xWeFiaQ6EuQg3uMN5ckJFn/AFV+gytTObxzcB5aDMGzQdqGGV63eAX
gp9MX3AaMU8AB8ahRJ9gfvrOSG9PIWTUs8+B2yKdUrBlCcOQc2mHkBxvCHNbbYeADShXf1s1GGKT
QIm6G9d0+X0TLIMk+oumA97iFYzCFBSnw2hCMgZxM6p6XuvJatsTyzeu5Alqh6VFeVX5CPhr4+Ad
sw/LfYHPvtuARdKOh81qJlvjGzCsof2XKe/WEfaHC/7qza9E1h9ty2I+RjYxAQrfrrJ1/UkeMqTF
WjYNrUJ4wO45cp8eqoFYM6Xo7U3/uaiKAWc7gl+xYNms92hvs147t0r4PQXrjp9rb7jJSNvB5uup
MG2YBoGmbzAGzkW9FmNtGMWVoL2o5gniqe3+PylAKYhCrXelwGq+SK8X35XYwiUZ8ZECzJua072P
79NPgB2dudr1LwOkPX0Fk/ufiQyvj0ziO6owWROFfzIeBpXtAYXNa2EGu1WJ8gz5Gm2UJq+KdRBa
kbwjXTXG+eJ3z6L6ePPFsw89myEq30J7P0jedrdWMARXqUqpdQ3QF3cNWjrHV5B36foqnHOhq22f
kmr0l2srq52KCkpnzeazN1/euP0BXLJeQ954/v6MqdAFQlEF4ktxoe0W3PmGdJvqOE1HJ4c979zl
fYKvtUK+pK4PYKWgjYmwWIZZxZgd4NFF7oej0rLj+1DVmkTMnKXpvwhkpnXd8tOvYj8jyBU3/N9e
fEXVD6hI/GwAm3EOdQPatRbsQYcav8qxa9J0y0rcP4CD5N1dYOzzOhybdR+r7OJS4OZIix61eA+/
ue87t4ohqq2xUgvT8+BYJOFfUIBy0TLl1Yt3wN+LLvhuVN878dPIMN5JVD8mkBytmGv8DG8SmHq5
kcxUxf9Yqj0/ynPi8uveQpdptgJy+Qf69LQfDOfWPB7ydRus9gsGbqZklbd2eYEdukSzfq0+uv2F
ZSH2l51ohUA+KZWGetoPVVaDNBqqLKUN+uz6Mq1R4nVNbsD/NbQrV2sTNALHLrKpsSt+xtTPdyXM
Z/Lt9ND/bEpaPgbea8+m3aDXg4ZMrdB7bWBtDpWTFPkGyk5uTJ1I3wNQPNRcDGDiMBglMY/VXsiK
GRBH/WA2iuutlLMv9N1N3cK9L1sc8cRch7mo1lpQ6Ep5QY4i7SiAIb1xJChi6LuGHUalurCp/ps3
XgABwFFtYEWWQhCmLQ9ZnyuCg9SSeuL97Y470ZCO0gbV88v0RgmhYMlnMKDXl0ftPaka6YlxBi+d
u6q5GP1r3CHQGeK+eRGgJRA3GqgWArT+xVyJ6f6C4l5byz5oiPAOmfIdDcP18s/hymN6l9o2D45l
eDFeum9fKk/W/btXYwwmdjXJUfc984cEojMz3PHoBaSV9D3o9rX9pbzjmSwJ/v9ByvvndZS4p03A
Q5/FzSHJU5F+oIta3krL31Ho95Oy4oiG85QPmkBvCTOLhEgt07FeXHLRWP5/CuVlTRwj2BJ/h/2+
LMzO2BkpvrwwO4FvFxbDjgx4rWSpL8ue68Xffgyzuxf4OaZX5Fhdjh2ye4Uzz2CkDinYwE7A+GP5
R4KNukVaQhAPdAcgY/L7X4VERY8aCbLS+FMlS+B7XtJaYrBLTfAujA+jZNzYpS3mKIR/SUPt1wKI
RqBd5h+g9Q2pZEO7iIEJyDLKM/hjB52DGgq+tdPORuE29SHuiiaaDK0bH/iLM2/FqilyQ5Uyo1vb
eWo9HdqLBCbhrNcCJJ+xngSJDX/a+moHRRbtQjUpmxj/xVFJZ/ZGRE5jOeKpyUI00N5Zy08zdY5z
ngXAXEw1P+YNLssffg0AYwqdYiWnCXId5HWdW3R65zMEKWrrCwXtFdqFOV7450C4NlVPGgP1h7Md
BU96RJ74IW862Q1TbNQfFmf4VwTWIsLtC9FbuvthLkKLm9O9xX2qV8GNOVaeqtluuYe+nCazgKtX
/8SfMnEJ2s1MGMEYyots1gNsHKdfnHUYK1px8LJomxqR5V5MJVVoNFA6PRJJpGG7R25m/SC+XYnH
nGimrBLqbnhfox2VEc7VRd2nP9/9Ok847UlHFLql9rSYPVrE8Y4XfPtBqRdj7V3kNZ4dFXbH+Eoy
k8qmhpeIvrCaknJKdE7TkjHF/GnMPPVj6N4dsu8FRMOEMDoyq1swLYlqLmMaPjtosvrl1k6+Mol3
SrC1LcMV9MxiW8g5U+KztzxaJTEAxhoCShIVFJdXkY2n8LgPcK9MiDZEyomKcJhWOPCtPrC5XluS
TVyeVQxuNUB4anhDRkg4SjOgzjPRjGaPzN8tOqUBRxI69NbWUpMfCsxi8ioTFZWeDq+vusERf0Dr
+pBVdYVNx3FUVMHO3hU02AXhNchZxAbonVXVPtWj9kD/fhn8QACjuiCSsKXezxOLSP5EBTRhSxml
UGkYHP1qqS79U8I3DrCn/dl4VXOMKlpczJQIuZANIIKCnVfuh8NIKHtcU2Y9ycCkhPne+lSrvaOS
Frr7QXRwu3TywTtcp3biRDnagTsRhoriAzFrwwe6KkVHuEQeO/9OiJYEVD+VIwSeKNk4EFd17l5I
G3xu+LxRz2e9pQzS9ULazlRaNfHuN3WSOHk+9/EhPdNaXC2+GSXwRZBg/nSadaJ9nWEbkeW7xuuu
0ZzsIMhVrHvorCdDlMBLFkOr/y/GIxcwD7bEdixGX1xaWxUKAbqOy03wLnMgJYV44GZJRwFR2P3n
7L0bHuU1+Dh4yzvhB7UWr7QIl9sNfd7sDGTz7lF2i0ABPLVmdmXJvLVSIso/pX6oLLw8GQPVBR5N
4qkuRgzEvrXYNHpn6aRNfFL0pKW0SDzSpAX3BrJmvXTDJPOrE8ZG0ot43XWOQshv+rL7eicrf3uG
e5dbCbuVmTHTeH/5xcHrNfOeTaarVLHovdGTnNA3U9ZA+hdEQL42mcJsV7qYz0jizWLmMtuDdMbP
lis/AWoUyiMjDOu/WIsVvqXr+EijaAwXu3UkmCh7qs7feH6Wjry/fQES1TQNIfJrXD6/jWoyBWTD
htdsgJmmhWUPe1MDLOZJf/MtAs7COWwChZM0YqePgUP73a92pOtGqEA0jW5JzYy88+DsMSJzRt5Z
ra+epXDRqsyOySCgz3WQqsRU1L+dfApnn9ReIn0suGe9UwZ8XoiKbXnQzB7tr937+2C4YefJocZ9
OHojuvcpK77f6KeHB4xgvH2DIuvUFujwmhUiiqcbkMdL+RNlUmR7tJY1SzfjbG31XMtO4zbaNZwn
w77M2cXS2RRx8DiJC7sGZKze4xkn2euAVZNNCPW1aeeT62DVeyyEVf5nurzPUKM4FzNIs4mCknfU
CUcXl4Z/F9mb9bmm71WzvMBxBs7Q1s/gl1zAxQQiIQC3xq0AwxY18jzt0X/QkyQiz6QCjGtbi7ss
xNDQfBJBLFLMr/jxf2eJq//wclbOnL5ixgJGAXCyyMQzzwimIH02mPpWbpOicENIJq0VfRa91v/L
yqbglHJ6f0HaV5apL0iNTTDhdzQW01MUryhqOtHDitYnOxEAM5TSyBBQcr7mlWXaKEfRsFsA15+X
SZzBEpSN31+KGSu3Dg8ylaSe5ficSiUcPVCDPA98QKH0GFc4UD6u9lgyZ3f6t7oJDGcRxMriFNsa
eUWYKLt3z0q7agEAuO9WXRsIeuXTtyE2OkEUM8KIGwPwTuY0T+eofkgycftYz61BrfoWbXia9Aa6
sd2F2n/4Zl85tmsJPM6lJtxCZrjCmsyk5vhL/xn6XA8YRV+QYkZPWxPfAeqdtoIOyG+z6b+GZNHB
g6iyO32H8Fao7L+wO17QMVuW9hd0Q8GIRp9GRxUKgB9qd1q3ZEocB1goK19+PHq5OYRNFYSlucDb
7waIeUeYwAigNS1/gqRfvaiPlkBUL40tmt3+9hrChE0HKXge5Wt3jGNTMFYLT+nqE74C2a1Klou2
SWwb7dkZOficFHq/4oKXY+wQ9RpssejiN/fwhCD5cxJLDefEJlfxR5AWIl+0WtVJ/iGuH47kgVpe
eWZD6/Y2nsS0e6WbxJnEdL83yQIX4R5IyhYXAzq0kTUjf30Dd5MGZEbQaIO6CiGmNkBjnuQybl/x
RA1VuNUDTiGh17LmqVx9qcoF2LCIS4LZS9ISM36T5RIZviGEc5ftiR/SZfLUnvKBOlx0uYqWQVLE
iNIi79L0LSh8y3Zhqw9Is2zwfRGODYf0bar89sFMOakHc/c9aJWCqmJ2KNEjEN3gMOGjQJFit01R
thuhxTMIlax0PokInGoWq2MReXTcUfVs83f8QgHH4e3SD0sKFjWhyIOIyXCm9uprsZvLUYnlsMcJ
vlj4OIlp+80qLcTDKdyAL2ZrfDT951E93RvQRGPgfUt2CoJvvbDPcPitH8nhEIiVILb7IDVr8px+
HphcXnl5fkgB3HYTsrChZc59a9P9xx+LusLjFWkahSUDNJXQcmT8+wL/S0GsSBpIOyyTYrN/O+l5
HACTG3+udv3y8mCjnXt8OCmdf6QHTomdJtom7268deovaJZUCTQ8UPX0DEKAA4EpA5Nvr2kj5LX2
g07lD9Qq7nZ7xOTIF/QIU/9wG8zadGO48/S8FKlYp8j235PO2hhpVuiQbUHTbMTVjrQupcpaIPT3
lCWDCMx8xAWnD8wZ4a6arNXrGYrYJODsIHZg10rPg1gxfjSm/uXUl0r1VRTOOPIOyy6j6U/ojGvv
ivK5DYDsjVyQ1kdrPh3Y2YXk5zpK73RKP6gSwYIuNaEi5EDTkxIAgAF0Q7fckgwndsudPVBAhVKL
DYgChapQ/Kq/XS4UcM4wCakzT/lhliTQt6qojbc3UBDEgAgISCEvjKB9IWtxv9oiP74L6WvfBIhs
N3qg9SlJw6o5pw6E2+6r8/4WVSSowLQpxnMWZRApJQz5XJwCveynqEbVUw1xZYSiSdQsfXAkBfUr
38NDexX2R5hn+ijR49mBP45pczsfDUVVm0zlQrsnLgGGzfSZwURVr+7IA3U+wwhAnyDMuM1qJDrg
bnXUU92dYsWP9MJEeJuauIHo4kQnr8E6zp6nIljN2V2VsZ7qdIsIFzOerzmxIO3EByPdw7dD6xAE
50etOb/RCMUohcx+AGRQZc9bbB2X/Oh5/CCwkF/G5JdbNsV3cf020bti3Vk52sWpPRlnvONxTZP5
6vvdOGOGfz2nGJ1j2olrKpE0TDzYp1B66z6qwkB/YMqbx+IJ6i22c70G3j40XaJPOnpzXuYxTDbX
T+gTQuq2rEf/2z86xfJWlydtwqYOhcUNS69a+jVVsnDSY7zVemA8AzTmNwblefv7F1UGXMRpWEfO
8vwZVcvEkEtuxjWtoM19ZI9J/qkx7RfNwHgjnYDbmjstnS0eWz0WrTl2ECy+zYOAMosVMQal5DLw
YpYncaHkQCXySp0y0CTRQp23jGLLVrMZa1MpiB0nrIsc+kX/PrbZsabA7KPkQ0TmfBhu1CN+2V99
9b7DeOMs8kfVgKg1GAl1GxfcOm1BJuemwMa04f2z2bRCoGyt8NAUsQvud2mlsOQofvLTmymlmR8I
calM8d2Ks8BrQ+ii4ll3rLaP9YrQ47KcVfuUhkFjiUITu2Le7TIbtT21f2+1ASixFN3rp+Q7P7OK
FnveZjtFE8fbXmyGaLCMp0yJ2XOpxqh17xheCeHz9UIUeZNEvtrxbU+lMLY/pFaxFukf9xwtAEzu
x0UdZdraZc14x2slmNhtYnCVDUx7MJ0uwS2b9aDvwR+dxKORo0mQxnFLtslwxkCRCYfSHZIulT+e
N5OmHkSvY8lU+3CR0F+9GHdSyaapFSZ3o1CYtfPcoD7/AEJtWVKbXliHovkiPBFSeQxxpaGE3KfI
0rFK8NjpPzDJhAqIu36g21fSNpozAQdur57kf8UbXh5cvaTxilSzaI5ZaW0iZ+lborfbtXZ4b9s/
ApVwJEI72fykqlY1N15V6+froGIet2UKyLzQVkEbEJUwwmMuIf1OzMDUCezSjhbLoJ7IxUGUxUWy
6S1ogD+CjPHFYadwcPtF/oOSTv+lFmcP2yZzrgbbqLYf0PdwhtaQ18+2AGRnZ0zAFRM49f4lApSU
Ay/SX+IvpLRybtXTH3u51Tb9rD6rbumH/BtjOiQBkeqiEbSbnimXNUVXIyN+SSaHUQky4PQA5YFm
VlZ6rC++k9JmNNm3YC0sYxczclmqpFXYlg+QuvpeY9vqnaeTre5XVW0ODMUPjirgnuT2NLiXuZ7+
nD0cJE8E1dUYswH2v/vqB3GYynZ4/UrJKQ8urXpeODgy3JOI1flGc9xt82Dnj7J92GWHmU0KbqwB
At+DotU6SOg0pRaSnGoTWLOiW1mMylmkeZAI8PH5tlx9qgZuv+fF8+F3wv6fiic5NBzfq8Uzz9KP
4gI/CYiwEsRi8gNsHwWQuN4NwEHRIcPFUzMAnuF/GpIG1vfN302fd9u0XDyUhMP263F6ltV1NhDA
JwK6L0hKgURpLLeyYToLL1az10sgUQ6c6xtEicwGymHizeaRqIDYnWlR6D4qAce7ZT8wLmhYH68j
28yrXpgrZhnuQCbjOZXwL+2nbWipViBYYOxhB8p9sd1z7D4kzu+UgCuDQExD5DTLdBngYDkDrEQY
fFrl1vNB+fUpZKTGHuRQXn0y14NsKllot+exUR3VB9JxAepElGuHYB/8+SkJih3z7rd22/XftEFO
e1dWFGm7jUaCmRZOaN9e2Z/1EiKi6cl4S+NpOmhBYRQ5nYmt4YpcgQKm11EiDmVb16jKl0dICdA2
VE2zJ8LFFrsOZdnCTyi8D8GSYPXc53Khr4sIdTXYPOZbFq/J7tIRiRBJy9TNV0I/gikjLGexCKO8
uPRc2MBVlkNj9OVE6TfJGwynt+HD8C920lX0K7DNUZHyUdku8tlrUKPVV+ivc6kQHrXKC1FiKO0F
Ac2XkIAH4xTu3dVcpeiPeO1aYwyZ49yWjMHTqHN+r1ZpcYPaKiSf80pNWEneYTYitNM1hD1EOEfL
2UW/PKWG+n/0qQZ22iiagM5lVla/3a5YvdjEzmzHvAXjlg8NiVlH9lpYHAnCIyseESJI1tm3VZxM
9GEWxpevhWBysrHq/VnFb6KuDvb9g1txI7usbETTNxYi9M6dvfwLDdyuA7fKcJP7Xk77gt2pnxB7
AubdnSl9j+NkubzDmVbRUK4pk8FnjxiqH+H5hCHGKNisUOiNZnp9g3ISKGdxWoRjSY3xRL2GFRRX
Mbv93AwHLwV3fwfAxBZwgctgw8DHx7ZtKrHLZiv5HjF5+9HSckTPSgHUOZCF1RYeJMuy6nmuFfs1
xDkydrtgAtDJLqawASCxcOatVMABFXZDW5oJcuAftclVBLAqDV1fVqm9mStl6mPv/WK/dapoJcuR
aMuFG7mePZCzPpWjgOvB1hi9h6Otxbskubegdw/+g6t6B+GVYtzW4QL4q5k/Y398xhHomf7t7ZRL
x2RIf58y92Hgbm9kTmkz+0VyUJ4hJiAa8VTNeMSALRNHka3w2iqpYCpkN838YhDFMNH1NZ2A5806
H/RK44WuKdWyAaRZlD2B236wOikKEt/m4yJsBh7IFntCR0damcm8Q2/OIFMYIjQa5pDEWfjba3Ye
nXobBobrHImpYaEAUzpFxSqcA61JbOA2GG4SCUkHMHc7Pc0H9hw9dstODVrrntJLTw3KNgnwLTKV
+ZG2WbvoUsO4OyFFxjodWbJtwW8UN20QCXfoEcSoBCu774OrOyeq4pHzMEXRSOrpeQN+uD5f/flO
UMO31mwjkSaPMFfeeBrzH6jlZAyOZx8/jwsz2l4/PbJuHO90rR7N6dVWJnzek6xFyAlCiN8dQW6/
L73U90zG1e69NEi4PRVp8AHjz+LuPI/TLcMaAh0i9SJFlx3iqZQmbW5sGsM4WQQ3Q6TTxOsaxdd9
/Q3ExngoBrloxr5PvrAOyaLoe8CA982O7rgGCj73YviKJVo4J80OJZ7wxeqMtEl55ZccbfNagiNH
utxdOWAg463kklYS97bpr/MR5VBrGs82LTcw2tMl1rDVtn2NKj2g5fX/N9VCRjzQ9mWwW7AwfVB5
z9kDe6cMSHXYL31kyESoYYJ3StXp/5glisOQreeipQt1LtLrDHwe4BF2OkpJ7pV+1dsLdS4B1MEg
yDW29aZl7FNN46Q+ToZ+XDnvtoH6mpEcJHFeCGTQ1I+D7PA8D7liTDTo9eh9PrAKlTPyJSHpmXyR
MKBmklqeJU4Y98gX/Zu9KEoF6COfZPvT7KNt1F/0sQpkgA74DI/ST8k46JhU5BAUsM6ILUdc4Clv
yI8/O/2Apkz1VCCfj5L96+wNdt7PhC09sEYrWeDDO/VcRXxIqVrCl9GM/t0VQhtUxyJFOeYA1cE7
cZUCsrzbXtpJxldrR3V9KFTPMRXdY922gVzcHKRB+jB/WX5spEUpAUYqnT7Xs2upa8+hfFBpVeDL
klfO7TqEJE1J/bQq9qqZlf4FG2Z3zWxwpxtx+BTHwqwp9MxDIk6gPhu3jvlTDi1DaslAtnaduT/a
waTNO5T9jSEcWQHPg+QsMS+Tu+xLLA1Edy4r9ZrjkseA2kb4Ka15T4tMPfnvo5Q6f2j7QQ/V9ag3
6AaNPu9Al3M5mxKG4P8IgGr5zx1ztRAEUL/y5FKObD6hXZmdopG0wBx/2fswVUjjjlDl0K/zbb7Q
iEiLrhfeUCfKOZVR6JbNxc2bRcoLPYOLScCXOsSfpgCX7GpIhlBzz44z1ZoVh/5gHsuXXPM2lAU8
Oby4sMK/T0DftyXH8Gnt9qHlN8jlxQ6WDUyLJIkYowxrCq4BACiUgUL7+lEt2e6LugWNLLfD8ia6
sECrtpa7foWYlAWxuHK/G9CUOFLMYBjtRrHjZsw+7pXpKVgMbtpybwrARLf54hApLK9H1BlPtbv2
yORzOXNZ3aH2Uat/vJ4mpVnM1pFsi1lgNHrhnHwA1Q2Med6XRpB5N88DOH6T6G2fkXMbB2wMxuAp
fC7VBvx1oLd5BTzdFUaaUaO3KHobmJKwuPtcEhocwIjiuYsflvmmooXSgqvF8URttOUEqQoX47yZ
SRN6pf4kYnlK2fBZKiabgLDbt5M0XzHpBTMu8KBapmGP1CWtY/+e/MbRpGxfUe6cKaHU+VjIKx1u
cX5nMH7snjJG3vLhhs3Xho2qoYIwKE63FUlRbLrcf2vuQyYxGuRWWzE2egjgpxMTg4jxpqGmxVu2
/u85LNvfUqlYNDD2IhcZz6BrYXelv14db4HXReD8SItrTT8Q6vqha2jU17XXZA2ukX8yseLO1jvy
9sVXsBBao7+0fTMhnvYz7RLPYbN8Arbzaq9AcE5Z4KltxJF7dgGqT8dB9+Qd8M1kwucClbjwge1E
d9QirDnFPXxjQsZDbHUJg7DU0KB3hWchB0fkmqX14boQgCMovSdMNVx8s6tLkz/j/+VbaGHhvwIt
Lyed5WhoewyVH6o8ZSsD8DS4apqAJl+6JOeAfaNnGIR6Q792PaXlkiv8MODpxgXIICq7b+WvR5WV
/s6091gWXwwnMVIi0JMV56gXmFbG/l4WM+vOxb84Kr6vKpXT8EhUX3y443shfZv5soliXiM05yZb
FeO2wVJEJUDU7AtOByJvuAO2Ik+x7z9/F7s+sYLvDDmomaDMBg4PJbFrs3oeI8Rb6wk3AK2fbHwr
TuKfBWSRMRrYr/0R5ayxg03m3KYYYt6Ae/xRSzENrl9KCrw4z5ToNc9949odWuoOp49r8Kq0BswD
rNmHQnGNqpYVHVx4dccuhzzDn8GUrw+00IigZ4x6cpvZxBt5XfZlClFXtGxIeDtML5Cqhpz4XSJO
mVCiCtk1tN34oS237EVstQSQ/mVk3vZDgug1h2GgvXkyfih4T4dl7SQaHwarLMbQyY5/xmAF7EHf
MoqSvVOYvREpieJKAlcNAdCZn1JUt2I9x3qCZQJBkeVznZkbJEz16aGCT8fMgdMMzOuAX82m1u1o
7iTEGO5tNnLA9IwnH+OcrdAwYVTPIi5ihGvb2XWnkwPo+LmlWcr6yhGUIghyV6m02y8r6D2raAa8
oPAvzguov3Yfha8KR1TfQWhRPrPAAa9jMbay1irWa2FZN1R8k1XGILyJe+WmlAXE1V+4fJZ/PFXp
dAleHRzgdEw5QAjnPd2T/LTsF6eAivUTEEvQthYO6vdibZPWQEGQ/SIFVdkgIRaEAHKH5WTbLMYM
bw5JF9h2/ChEXzZbJc7BGtFkgIO9otesa1W8iuwnsM2ZAoCztvTK8eCh7HZNg5arj2Q5qEg2v6OW
xqBoe8nfB0TP6Hwn1Zt3ZHROZNC54vyfIKAmNQ8kHkaQ0tYtXghkWJ5NcljNqa3J+IM1WAEmmplH
ZCHRT+O/ZZgVu4h05StIdl90NA+ngcbtQMYe+tK+mzih66W56pZ/HgSXdNxcGTCoqPJuYv8DjRba
stgJFr0bUdt/zuM6fc6/DKRLd/AV5shoAiPcjxCVdAMrxqGz5Pkdg8GCh6p0fBDFoFhLIwSRhm54
XuwHBrqa+vuvekiC+QXDAsKbCnKeKj2TUNLgYsc2WERVTWLc3QU1miCNb/bUUX+MsH53soVcqrtr
d9+PecQvcWhkcYrfSJ8ps16GHWCsiZYlaaoEvaAeDXQls4Xp0mdnU1ESFqTmOvUKvtiv0CXQO7UB
cy+7gZAEctbnujBzUxangdqt0lyqQy/7/NpDnhX9nvEEjhmr/npJ7qhryegYnnGHgOdUzUdJrkW2
AqTfX94NQeBhSEtN/6u75UzcYHKEYXtT+FsSD9dq8CdPw3iAXOKIC7n6mK0k3ix81KpGo9hYNsoi
+CYWfyTDDT1fUC5xZJcAGQxjosbx7bNKxlAZCFoUbvVS6EtS0ShRpbt9TkiD+2VZgiyNn4mF2PY7
+NbZiG868iRpgXEUeCwazYzAL7XEsFOYeW3mJ7/pMt82Sy4+aGmrzlwoLyco1kWF29mnyD9qrJM5
2JF6FW5Z7BfREO8dz27/viVeQsC09S6PR8/joRafZJ5dOwNmBM1394gEHI2pzI7ywzAQBJQxTSpH
LXfXA/mMH2Sm16bAUALzQxLC8AxBBOpoW5Rk2Fd5g544P8wF3S2Y7jJAr56MSEuaePwngHE1zvsi
wbhjWBzwg5fLy+bkQMiZ7cK95qav626iE/P/IrW8ttCobQtASwl3BEOcp/zOQgFR9v+yLVnNTlm1
e1hzWn8rVUhcapy0u11V0QvwtLkF4wsyXtWvLK3uvWblm0VTryp9ngwjy426lta53PwTiZGA7h3R
gXE0Nl1YmAFg5OsTAbLSWxt+4NtObX8veNCeF5UM9t9V9VsXEvD105pAepheXYwreywHUqwdG8ME
EdLGrLG/Hp/etie3CQW5vn2vU1E1vovteEJLFSNunoMYmizShWTE6y4zvgPXz7iwrhHLZzkTaEo+
DHiBQThOitHKXLKb8pn/m2pW/tsj2JO3ylEzmkRq048l7qlDirIzNpZ0XfTTGeUgu6sGX95PriDz
friONtbiXiPSM5lnH/N8coEACuIz0TTB5ZaJ0r3YfXP8Kha0pcr9lbiPNgabPgyfKvP8KZ98wFwp
DhzebH8FV16rfPfHlkiGLJM86qdXD/bEawGwXDygsQYMwOKVMZqxIvkhiGPYz5ySJgphBkuYHgdh
NpWe2GZ2IY3Sb34MKKAUicpBJwAYjqpLCf8ACj1dXcht+wlIdao+37KgdJRAp6QjTw3yrN3WUhSq
3LCOQHIq+wLSmcLwiXzHX5g005NPj58uDOPzQQskuwdDLOWWjP66pBZeSZrHQ8CTuEL868k1n4oH
wifu9Tygk56pmJQbLRgXvEHx0zgyDjGvDySqm1pvrc18ZQiwfQUolkd2W8ymJ8qgWsot/7cygvhg
MpV9fsMMH+fc6jBk+rWwsIefiAg5nL7X4gflk15RI+NuSQeAyCs6CDIOkdGrEDFRqjt5uxgyu6LB
bVYZVti+w66QPjsQa/J0Z6XlN7UFaRQzJgrVRWJZY+YnY40/xnbMrIwMFz3w1Qnx4FM8vXItmGzv
7SL3sCOmXicJorJTC6U791QrVht8+35CQ8EC5WfhK8ULOkhVSsxFVvfjpui/KCEBYlTZscnBHLuj
5tF+MFc+jRCQ2Y/9L+gCTlxpCVZCBjhitOV58vLafp/lSCE2jHr5FjR1wH8a95m2SrD+237NubAe
/EngcjF8ydlxQuk/tKCABlTucuRwS7kR/SaC7OgCK5DKIrcHd/AZG+AvKGT2Uae5GRrCqJ2DOUOk
HNd3wS/rG1PjXqAfQy3PZLplujNX9pqZav3qz8TrCxALOtLzxlHTSjVRJmerajpzPuJj2nFD74+2
NxMGwEad+aOi6NBoYib9/S1tjwhlqLySu61eFOGKOVS11sd/tYNcpjCiWlpeC95VWjMtDbK4xfQN
HPNm2J2b63jdjtXcnzspLN9kU0hC3RIiXqG+a3+n+MttqvVl8hQPbS5/xcudtsAm+rCmBevO4LfA
K2suoJE5p+yEQfRO6Nz1vEVqWf16fo45Kr+nNaR4IHwCkeLbVn3xKSI9hdK5oUhQcFTVoHrw0rbA
EfixP4H2SzeSJLzOh/83FuPgFllHUIPCx66GLLhIYhqIfb0jXUMHs/OmgpVTPCuAiTFDStl0LfZw
dVHI8ceLocRPkSOpwIp1meiP1NUkChisfEg0kybUkF7FabblMdcXMQ5+rKzslcz+qqqKTN4RhlJG
D3E3eTlUxu+/xqyk7vmXsCt+bSVz6a47bWw5lGSIoiHLku9UQC0q3M7Ts7uRRwI80RgRgaIwz8a7
7LPF2/vcAn+DBxEJjWZnxOi9bC64vx9Cm0Z4kactSu8lf+X0GSLdqdhotW9VHZt1qEEulSUqa9dq
TAVz/h3kUZnW6qiCphjpbldwpA1+435ZrjaS94cRySNh8c6wbmOXwrWnNSpj7bHSqE0LzT6+J4t0
Vt6sWFMuaSZd1+hHhUYlpQW1Crc+LzDlP43qGnvgbOtpa4nuME4ysQD4NtmKq8gceTQOsLToJgWj
rqVVT9HcB1doABGDSi+tMd3BqtkN1/YeW7K4gUne9ldCFztorAH2rIQ9dAnW/wWZ3c4SIhIK0KvK
TSC33ZlX3P71t4xd5rbQvfZZkXiJiAVhIn8FI8JVt5U/m5PAXKraIa2KO22//IGzgGNzBZRlqOBP
MydyfF68J8VzkkZhhrSUMkJ05XP50fT57hKqdPD6tGAzeu1qD5m80MvYjzzqfo0c5teuAlhZHdzv
tK6FDlVQuatjWZ4w3dP6wTEKu6Gwd4rCnhh2sL65lm0W/V6Q7n1SAl8yHmBkNE1i0jgQ086MxAv4
kzjOdh/QNWDIG2t2iPGv0nRqIdyRAyeOAy6hHZGl4cti3sx4Q/LvJOAymxGbhR7ZWpu2mky4pMEq
0U2oes6YwJXAWR3MxFAZzs7aOEqDhET4xzGtucE4fdgA487ey1Lu1JlXLGzO5CA55W50kj8GsDQ3
P5zIQGD5ROIcbP4G0pAe0FOnn4XA8fkBnNOrKBOokds0YeLTSuHrJwrOadErtPMAgPGl74NaP4P8
73oXfwnZ4wbNEqDuUbgRbMP4UlCoQQZh2XGSYK+1fQZGwMVScNNng/ry6zfXQdlIZzWkGxlxV5HN
eKi4nIK9S8zyBzbwUfnNI0sQF8YStpDVtClr9/81SzSRmTo2Sdw5xENZXIAvXVg58bt073p2Sxle
+nyx01IpOq3F9pIeUfcJVYO9tMd0dat28yGMWh982rYm+n0DvaGUh7Au0Tp1hzZOLv4v4wzxuppb
+n18cJvt6CpKTnyHkt4bWvVax+H8CjG2GzYVJ+qICWAXdEdLS2JIZtJmNECfEFeTu6SHA6OEtI6K
oclzwkqxWJ2Qgl5BET8ExC95pXfTjWn/2zAbc2ZQpCWbTEyLd6MsveNBfgLg6bMyxs5meFWnKnuN
w9k9LtIo33CmqnuaTkIrEq4sxA1raTQSyMYJUalAQptIpYac83BtUjQzByUPG2JZrRHeh7aQL0GX
pZbtY3P8wlveFGRJ3P6Y571bwAa2DwUMKBS5wvXrW3PWKV8PYoBaR5EP4VD+rLE4z8pACzNocWij
f7U+SbjeSNfBqDn5RnvOW38XlWTj6wUK0R7RZugaVirFooRyyYc3/8093dNQwV3rNANTsFzy8Qfh
oLKFdFoOJNJm0YNSVT0XhSZU4ulSMNDVKPGKu14YO/b6tPc/JcJwIkuk5RjVNQVJlDNiDSb9wR14
8fEBAsGE6hldeoHzH74qTDGlEoKgN4iK+GPsEGOinoX7UOLmV50vnsT2oznHr/NMhGQFcRA2pz78
FMYdADrkcHKndd/7C+KiC7u8JevOHyEF5hld3sxM7s5cMXCkFqZZiKZCH0m5ayP5nfGwoVw9FG1c
bZ1hQdbfF5+weVvNtD18xEzUJUzs0FCq7tZDKedVLqum+8mtWzZUFjF1J2JqEBj97sEV8bknNcrJ
53vGG8fIHkFvZB4xZXQjqPmEfAxrIVaIVb6HQr8UtPETq1BCq6w9shVfM71uoRFD9V3J2miORgEa
ca+tqvKo4jmuNBX2YMUp936k+PIQewxkaVRgzatSJAJy8SfVevUPqo3yLXjtkIVFRMMhP9GCz1cw
QPHkBE3pdwXDSU4BwCs9BgmcV7aiICsLtymbcnTu7PlPpum2Sjddc9JJ0PVusBIq940T/9Q7MXN/
mT9FrAXVeELpy5J9fOtR6byjZ0eKgs0qHhyLjKL6sry2FMoyHALIs13oiPjdJzh9jSC8cJ+mgGXN
qSZ2c4XKcdvVNbkMOEnku/4AafmHeuLTQhSxxF54NBP1FQQk4Bhe35ys/jO4K2Txftgw7UexjTbX
EnP3yGy44HoVlCf2w5ckAKyhafclUXam/KK6u68WTenIJEbko4OMSQNgPELdcEvOYkR4pIpLijdy
C53RuA6pl5mVze4j3pX8dZGILuu6yk94MFVNjigNV6FF83o1TDwiN6MkfnY7t4nA6cAJUGMRXQi0
jqqMM7MUXosrZkiadkA0paDsPXyCgpRrYhzkl6uBjvcYK6cVVZJtAB0827uDiJDn7+28mU1n593Z
55uDS7EGZzsM2cC7qINUJ/XS5A7mJ90Dzn3cOYf9cRcfaHo4roTp7hgx3MT/mEa8yCKQfWH7bpkP
asozh/FlGovr5FQn+5u7Al5iomo7jNvLvVtN3yJ1Cd5/tNs5ZuqI9Eq9kBBesw5Uu2/meQDh5EIJ
DCwNnTMNNle1S5AmYkKmn15YloTn45nlzCqguWTWYUPeX7EmQyGvX+0bWv+AjDnN/dPcn4bvDu0W
pLgXuYvz19AUBCaMDj7sdyzfqhqGft4uf8qreMUtPQpHPFS2AogbD6hghxHuALGsTigLR+0bZg5D
KsL0ZTbXQEX5zDkFiWTNXYoag9+COMhG66feP+qIZNx7cP/8JZnuKLUHrIpE0KWx/aKvC4oOB1hV
sKvCkuEoDHOp2F7cOUMnU8KovR5m+E+rJ8vsfqUoL9cCPcCfB/100a3RlOiklPHwH9z2r5qh/xCl
X32o3dGSZfOCMCKJyJWFBpZIz8QwzUqsQjXpUd0CJhHHMU03U7qznAXZvfm8xvJUv/0pBl5Tz9CG
mU5+GBG8QwhtkJBTou8RqaZFBOV3xdvVPdPlRde1Vnh1WZyD55W39qvJJdnXyw2tJFQcvyvdrvhr
TPbo6gZPTHgDFaoudrk0bseC7WXLVybzykzOqgAL61l27ms2tXOFLCuElJqU6pChCdzyZsRZzkUc
Tm3oexjThM1so2zXW+6ZZvjTNwI5iurpw/+Po6O+BRl5tFEZTWqpZ9jGxbYjT+F2CgSGx1ciTJn6
xOFJHQzf1LqebuGV0urCF7NV609oA5LNVVfV92jao2dYRQJRGKqYeBMFEdYRsFa2elQOvIlzm1Zp
ejW3+WUusvb8A4NTehps4lgTNtWN/aGDxzuXoLZHxxS1mrLQXHmYR3ufdbyTzpW8YlVkSBaK7Zz8
38UNqmly6aKd73sd9H8YxxGVj5/Apoy2NaJd+mi5sTauRoj8Z2ah8gK68WX67YdMlHMgmdojTvpQ
NI920Pp7lNtgFRxCxQzeh03kvrpMPjuJIbSwc8iv91ULFu3EqAYXjbca4dXNnZLOl6aoJ553DZ0F
LccGkf3ZX/niyGtJ6b6hNYbt/ip7wveq/88iHhdv566EY2LWLA7Rp5z3CqVEFbhW28O1DBY4w/k/
7gpuVDBcP3qZMBVk8WJjqYR8MBRtF13oTNFf6mYFCp8faJDgcd9J08Wv0DV+ApmgD8m2byVbJn2v
guTOueepFTS5VQN5cDC+RDHDqOEmc+DMUA0bqGByde3RYl2tc3vIWNe5biPEdYanMR7J5/HjTf/m
exfpdx4cJdVQzexMUDC0tOyFARCwHexDx+yrchUSMySmJnZTI1lYPFmQ4aRIAgq3IWUrjnzrmowP
H0/ZYLzc+hF6RXGksRvwFhUhSptNAcOJy+ylnxdTl5UGpC6vGAwg+KLf9cHC8UoTpBlfLCL+PDqD
nLoGSVZSfyj5t23QXD/3NBkPSBnBJmHCOHv4ZZQSDO8daXg+Kxx9WLo7PjzzN3Lz/eNRpfyUnK7w
9U37oNebDREahTCE1i5EcT/KEEF7jKgXYfTqU+8w/bLBrgeRiXZpW6YK3CAAH4NHsNm9cbk1qvxT
uTjSBSnm/BnewCt93fLJVjwLRM6KT4LSkyBATyXKrDWbAxivhEGyRVd1KclN7+YctbpjQG3fyu1G
7tXoZ4wz3DiwI5XIGkofBUcOwt5RV2ZSVDLXabR7hYXTjYbsKoLEKStB9wC2wXAoRqvZC2pPXq5Q
Lvz3PkJpr9L5IYIvoOP5ITLeU+5rSTArb+JTkWXdixTMAtUsXfUiJFQntipaex/Q5Q4Q6Ddiu+Y0
ZssilM3t7I0Aue9kqWyJHJZYTLwPGlHo2u5He8iFGcyvABdnhP+u7KMrhR4QhFM4n++OsiqzZCek
1W0anJicc0kmpc9sHdfPd4LmZM1PGG2vfHm2XCjy4H9FqfkPNb68uAejqyHp8Yy4aA06nz3lPj52
puJ9wEGzla9gR0+70kstoZI18UPQpUXRBYgSWeJ3gT3WegW5Z9eRVZOVIgwbo4WVnJ7q0t+zUecq
uuuQr98c4tt4rtcpo8L7drNbxpr/7zm6ktPkJ2SVp+xsjfr3R6aZDWzlsr1dLcpiOTeRNUxhxj62
Ng8NewkOzJluE863RkfgJwoIFn5KOUJsBVDiiHLf3GwuxDqLGg/KgiBOkPfgClxxZiNmVVUDqZSO
+vBNp2IN8/Geqim7HGxnquXBQ/GIezUGCwUiiBSYSQYGR+lg+vb694JVO7Ux4qfU1tGXS076kFAE
Vbyn/ORTCAUd62ZpvH1OcHwC8jZrumN6fNpnSfyk2Gi7SIvUgQUb0XW1Frahy7hrY6uWF8Cj+RoP
EhRP7A7fxCoLnWnOZUXwGWjAr2DwQR+C5GpSKEanebBBix/d15uQroEAWD3rL6S3VC/AVXfdF5kh
+Uho1lNQsdjqiJvuX9dMwLw6/bJLpV+amUpfePFkVwyTwJuWLynUUVFtvaICrfe0LR/WTx8mBFJk
Jrzebf+cXCPp21vAmygCfodIZ70Q99nGAEueU1+hr0cinQz3WOpBY1tiXlH3b67brrHbMKUf1xDF
U1o40kEngK3Rk4oeAuVEc0vpVhHqjUcERtB4pHhrssfdFzG5kyasrKAU9liRh31XbcXaULTMVg+e
NZNrcaFYybzXZRngwJCdojILeOTyUsVhvtGqm0aBTFESWbVWkzINZ8B7CCBMRg5Bz/POXVtAKxNP
/h/RrAT9Vmrvv2R/a5UGsbkk9ml7u74RXlLX+8B9Gfw4cUoP+OFZnGq782T8ndWCp06e5S+cr8rj
89qnkTqFXR7NTciJRNyAsIeDPACtgKPz7MR8R5eUYkRfxb5DU66XS1IBpk6EIyNecKSEls9zxsO5
tL+MlRRXtUOzVV6NTy6y4HcLoNGoM/4dcfo3ereqmI9dZZn4E3gVAnVKG3GM84hhWEzKEG0w3vvi
8RuzT3/uYmKKxlnH98QAqz9qC3PNrRNYQfihqNv+3SsNOrIhyEDhxaNzHGrfky0imug8vSBEUvzs
K0mt0Fk5HxDO+BVEp9aYdQc15xsWHHciEgs7VsT1/eKBt8GetP7rUYaLzHdHKmF44RrFkr/L+ySl
sK4FVbVu/v2XDfbW+8oxv3k973jC+iRLmoSCcxGhYE8iZreUyKn/OpP0NCKIhqRK9sOomn8vxO7y
OMb8wOQhDptZ6nyE27gwLaETQK/P8QorVVxmnFWC7URPJfOJZtMYIvaCbA63ScoFp/jJzwzwTfGH
aXd6K9BQnFytJJJfza091/4NruyS/H4OQ881D5iNwwBe3XDV5Wx7sDXp0CB8TIBn0JjwGUGvmmeP
E4PTkkIDfjCDJ2AEv388wLoKgOHtLB46BneDCOqlSO2giBgpOOgkgpwnWx+c2vb6KVAQtUrCGjJk
IwsVCDXLnG6BDZKpeU+IFZdF+qkT0RFuHgKNErcIozj3fCGCqeE2tyWZ9nTpzrvOsFzh7WKB2qCF
J8367wkYil5k0u2P2Az+5IpxaLO3AVo4g9yxMlTdx/9luA4FhiZfj6OsJgnlXd+/hZ3J1R3JTOSS
0cSw7RWLjbXplw6t9dlnKZGgH+zG7Rt5dM1WQTz8RrujW5KDfTp+DwVTb0t1hrGZjQNnEwAh5REo
gfyd1ytT7OXiPgXkKyYhp67W26jWidh/PvFhAxaU4hibVVC4OW22adFtwEZe1BuAH3ynDIm5Nvg3
B5jRUDqlz2LqlV4jMF6UUhgU6DFwITwlmZd/Sa4l/NGG0pHtrzUsd01Wk1BihChTDfoatfyRlaJM
xNEYwG8YMhhDb1Xg78q2gtq7IxArXD918urhAQNJTTO4i68QdoXRmE/oKLJQsLf3jEjUrruh1ASK
VALnO7MRV3VkSAxycA80kAppCt68H675n2Ip+9jTSYmIgFWzw4IpoWrcu+x+amDUhOXCc5lYHewE
Pbaap2NmqSre9Ux9gD2cXSUR+h/C36fsRcWFUfmv0q4BLr/DfNmk9kaHdCIZJgGLO8oApGpHupG3
N6qtYKdFJJxXGrAWLH2RoE8ghxar8oIJPsxCTIZeHLRXjR+vMrXNoXIVFVfzi9/DUbLJ4WJW9SZe
CshFdfUjWviHOroW1sl5COi2Cx/D2WVoqsfagocSHjaasy94h3NSYVHPSB5qqb7yN/n9r7M6o1yh
AEnC7SvwJL/62zgiBxSdPKs1B90nLxToZhIInBnbgMsNLenKmaeihYgIX2fuvFAlAIo2c1xpNeK4
D28niRq8ZjFl9vZBi4XOOTDIT+aoH9DD2vGMdlDwqNGrrkaOJmcgKIXTc3nrBZXWsqI2BinWBk7B
gsSkQ4I2Yc+oEtV/syY81tqRh1RjsjpT/opeCc4rmPXf6VRF5eZOaMBaljg0FAE/3/vnfQor9mLo
dm4d8SQjVjHCir/jRxs0lBNj914E2fqOR4iTDAZkEZcIUXPcctgy/f8KS9jkgiIVQ0KQ9umbi8mG
fq59A/jbROrwywBmKJBmM6/rKSVAiQKscJvmPCufYspKD/vMUvfjEKAzg5ZQepDVjInziGurOEBv
hDFSGm2xQmQ3IKsxM1LumRIkMo3cVzVKBml0z30Ml4EgfQz2AsuIlpaA6UrHW32bgVyV1eVC+5kF
ldn89OGjRRowSjUs11Cm388RE9Z/prTSfJPSm6c3AfQ5oN5hJzFb8qmT8KEThgkvAjlx15t1sZKp
sN6Hh6kNp/jsRnFlEoxocVXdRSL9FGxWYZcEMdDubK2Q9NW8Ax2yPPKIRBzXBvQ692e/2UhB8cs/
SmH9mFMNGQGAmQ8o4oUU6rMD5fQTeRzC3Y+2be14BXAg9sZrhiXq5hCYmIGDGuEE9JNzeVk6Qykg
O7XZoSGf52voklpjadTdONu45EXc+X5EG049vVJd6EPW2ZUNir312CgLHX5xD6Xg4qaekWVGPo+u
OaNkgg91eb4RDjqAXU0mOJZsHwwX9EsNVyCPKPj8cj2W3eeWtjZf/Bd2ooEbziq8mo5OXnGW3yx7
GKimWn0m3U3dx6N4EX2m6aUWoqtPHGRbPIxXBkAszu3n7w6kpphxVqoNeBZwMch/aU5XCQpc3DLf
LRonMXgVd+B5e2+7i+lAKORA68+gCOywnde5uVIecjxiKg81wDQAEtBZAX1De6qECKnEyzFSFi9M
74mkByryauxz52izLs6gcgeuME9MulmZKVjRMHo1Of3EpgTIlCiO3fg0HTawGjPYRcfs+0tLw5uG
5xVBuxH7vRxFr37NgrTpnOn+RkaEC0lg1mayLdx13QA188q69FoyrL0i+xgCw0LepimqGt6o79NR
zjfXYuQYSYuOZNPlqOFnTmrXlTe4/LTieiW8nDdwhjld+lYqC0SUCgqRvHIg/zkynuR9pg8LYL25
rwN9FtY9zGKaDCmX9MbiItXCsxnQdcmkBWHqMSEs1/GBXmftGV7GfzH7pa974JlOiXfff7fQ0V3G
8AMyh8/22PFCYQW9HsPTLBf/gjSr4xpCRFP2g2tAMvcvNxKLNqiYqAWw7nRkWK3Kb/kvRbTOkq8L
TATWPWJ2IIMHQylc5Av98p8QUXvxJhwtMrlg6nwgOZ298oSNmz4JKPMkdShjTgk5iWXNcORv+mzb
ztJ2OmDaw9UKpXsHYF9XB3zFN7YcGWl4bVEBqccJKKEdbwcy4hRZ6EpQKtbAhO0oVIuclV7dDwxD
/jBS+WKyuHGWp0S+qOCX9zANnXY4VDBfnRkn3WgRThYkrU9ZCpvkRk3tfQgzNzLT+wUVrPmOa9SR
m6HjL4aKW2tpAWjSCTSNXEHmrtGXkwBo2op8i36snDk8dOO92IhY7HxkT5zE57kOlYsJROOdI1vb
z3YSe9icMT15ZcINE4UdCT8qfGfQI7WslgbefpTLdRA20LV1wJcH5fiMRAqjgdAzw4HsFHt+OceK
hqFmjOsMlLMMG0y+3FUIdH3ewFDSMhWG5bZikdlXL0FaCApt/gekabiCgA1Azs9dtZiApWzPCg0I
m4OCcaVMMSYHfyf3jMzUxF19G+ar+LKOhMiYN5BL0uniAzNJCdU6f3q1Hxa6fxmtBM81JYbeI5Bi
uFp4euafHw7b1I1rCZeycZplPU76j2bHuQkG4uFF9iI8B+VwESmQOlbdj8LuXwy3MtGxlOBGXeqt
VvjkT/RXKHSuLYIEFoGeBr3uKa24Ck97pXX4wUHPusbUNIZvyZxk1FUBKk9ERCNXcULed+90i4am
u0/GlyhS/5Fvi+uNULGWeiwBH2HyiN81G5g94KCFgm8pEqVKz/elcv2t1fxcdCA9LWxBbT6XW0YV
w19TljLEbVS4b2jpSz3uES8W6rvjBQSf0UFg58Oon4YMAEpLvT7/FfAotb1G1wR/zmrGLNgJUVbU
WgX0CA/TOnOocA+9BXgCu1hC+IboANV+AyUtVGo9AoWFJnU1zuOUVCLUQAMJYNIDuK4WwETGAtsx
Y3RWVUtYpKXAxKSeVingFe5b/X9RJwa8SXq/eS1gN9OlDrQe7GYaj16TRiMRUtwKpwos7MChyVB5
w+AHv4RvJS4eCWu26ojnEqhE16FdArMs950wViYvrbgtfsLvunZ3yg1Iy1yZmFPaGv/mujsW4VGy
P5z9GB2N1BVJ661OKvNTT6qyrQqqUaGCMXsr3f9cwgQjquR5wCEI8B6SKwPamx2Vs2snztmWzWXm
1HWZWRDPo9bCUwo4AT7qisn+G41eUuFegs2h9culyQg4zn2f2DcGDCz8Jn2x0lkAc0G/EmnW5TSx
X//lUbjAoKBxI0JVvk7IlspUgwGnWJQY5Epd9q1D4UiVFHg020bvHEZhHWnE5B/FNX5BWaU5Bi02
+oI0c2mfl6yv84olqrJP6pLtHmXZogCTh6n4aKgo71HIQJtSOK/ps9TEeK9rCvf+EVfnHpBoWbZE
Rc69zEBEc4pRTyn1PvfhmYrKlEvs4kbEIGDagqKBAQjmG6bxnq3ZFPfnrXDb4tq1rtieZPCBj6mJ
QQozkJdeDoQnkIn0mtKCs39PBofTfBxX4mvskzk6zbQaYau6W8yfy8qPHBsLu975IqR5gVFtU6Rx
7NC+aB0ZiX8earDO+/+Eanbm7MLumGKmUrErOGcjQGE2qerHRT6OLZIAyzj6KgBMpD6yiOdPVdP0
ezgIYlBjaqvGNA0e64dwD5DTV7YEZK+Z6yjowuvfpJz9WmABgh+KRTS8Q48B6xCHfmBU41RdQihT
IJlXWxenjEs481bPdeT4TC6L104qklQ/rGnXnJcYRA6+6ldpvylHRJr8YwVITDgHup9i+crzg/Ut
fsyl9NJKa+14RatiPlW4f05bS9WA+6XZJu2V/ULI2FhKWz8FXOjXpayibw3mQJGsVEbQr6Yk8WUX
RmZSCdTrZiQc4D0YzthqjYFMSjFXp+8mufxHBvsmVj3z9X6I+xUNriv2L+fLFddgIsRQFULWhKUL
cB0NIfNDnokc5AQaTKb6ocYKLQKtRdJ2/0PiMHkA+4BWXdZMgslEyntgwNA9qzszGbhGiQWItYJK
8XMjaJdXpUP6tiBmSv0n7HhGagb32fbazMtPrNNkDdLkfUmbJueFNvGSspmNLJH6BgvPO/WMTusl
tc/qsNIgOGVr8SMgZ6EAFB5C4TpOJzaWy01AEYjdAayvI09Un1dsAS2qKRMCbTC7HHXEzIaCEluW
9mDQOK/UZgcO127YqDQ95ORaZEC0LcyoUiQTH/yJXcUpAhZf1XZqxe2f7wmiNN0OnSP6qNr8hJzx
YrNik06dQh/C6UecVuiAQub728VK4C7cDD/sXn6W1R8uJ02DDP4Nvjmtf9Sco7Bk+etBlZok/bWf
k6nLcEK4Cu9ou3KK1SvhfrnynCUct4rPotUCxRLf/e7tZTGKMcl9WXeU2rw6Qbh1k5ERHYEgqmmq
f8DU73h7ezpcfmw1ftsRR1aRBIyBkR7yYFl6/bDDnp/2iq5vmp7oHNuHgqZhS4KpA56qq+mtuZh/
R0HuyVqb0e2sCOAIJU6XFhyrWeS6xLZ5QjaTbA8P94sYbmpeY79ScjG/iuBPibpyYGputNwuayS8
E0Jnso+wwQvxIQkVjfzq8MQFrY+4T7KHxvxwrgJfF0PmAXk+yLsDLgTmZurKGzDjO1yrvl7hyhyQ
WNeQVEoeB01Quo0LOPLWjT7TSTt9GMt7O9LDIgs+eyYu3C/7CZuG6kwVeI+W46PUu4B02pZHF1Bd
DLy4WIu/09r79uuZGXDIYxoZEs+dvFACLf7anfcxh9+INzoLCu/S2b3blVmU1eN3RV2kLdKPW66j
2ddjo571/MpBDgVo4phGwa7k9XIeKWJTBHdEamNmYOFLJ8bd+tiot2rrfgZvYKK3YW2jQu4+ys44
w6eRtcMedivLoYt65+6Gm4N6F8tlp1cIPLURMv4vQ/+mS0U+C920fU6Q1pTACJlw9r6NjscDnFfn
Ji86j5PbbTVsLvTSF7/HMzbkLntqnGe3pF+Cvn13t1YycHGKe4hwQaXIRmX+Dda275BGGP+eKtPP
Y/Ak2pkJDHaHV9apOtU+nYpmlAKPaxOlLvWM4n7dJHst2jQ1nc3HHqreA5UqKgQS0SqPEb/oM4F0
2Ex+YkOk0RIzoyfozONqKYtSih2QABJEJDNJUPW3MNCOhqdhydYJHRzhZ507/+V4R++iGPgf2L7Y
8a3bIbtD6laU7IZuy/SzjWto9GiIkH/1yE3NHmtXDwAPY+UF4b0iDMU+4ZlG9UKiZamuCtdO9GUT
x3VhuDMHEhP4+6u5cwmWhyqrSPaigxitJD395S7JGWv9LLPiXPYlr2CADfy/t23GmIaPt3+g4//N
6Kwa60tWjlPheK9iFGW/yoWTIBkOJtIvkGTDwUcGJcIrvYoLCTrVuCjcr94kM9CF7Qr4bHs98J0/
+S/lVeSUKg13QxFwr4ajKMuMOcgWv5RA3uEg8YudQxx51vqILV71xGr8SqrKGebNeJ12Ro52ptE0
HfvilpzgFMpQ/7MImfNk21q3is+dvKF8rpY9vAJ/YthXw9sody/135Z7IN8JE2/ARFmxBwPuEi8R
IgdYVFfdJ4UAwRA9mYda6yXfkt16PcnD18qjX49MTTMsEHu1hSt5JVC1Kr5dyaOfTXlPHBwUW2ue
4Pr6yYvIEnhpo/9LDiM2Rv+QTsVBitjVUf5Y3470d7svuYgETL5om6fT73sqTenBfSxz6M7BlwYs
G0yvVUVCpY4jhs4sO9KbfeSTnArZcW8FYdR1hPXrqKnAouDz6U1QrsKZoJjLtJdtNlRqksDPqNsX
h+uBIOV7tHamPoHMfj8xc4V04mAHZar/tYObLBOs8ZC2Iz5lVsueKRcU8B6n37sr0VUNQyDHsx+M
98mCGQAzYoRAPRjVCfvNdz+YGeefyflS5Hj3OiiB7cDapiZo3EQGFxHb/UJvrhJbHABhKNd5g4k5
lOgiVlJM+qt/+riARjHmJuatmvqN0e1EeLeZmNbj2V3RDvux1MoCr3HYfoAcMGD/MgNR39OVHHkq
L51iwJs0Zrsccpp8L0uzKH1ZmKAwQPgDwq19U7nyPgx3EdQLZnfFdETX7X38Qmv6euF83Zr8jbIz
ZNXMIn7S0v7sGxtSt1dODx+5EKkVhUhlHqLcK/C+phwUAtrAKN2xEL57kb8qBZnVX6cM/uVuVxqP
A8xmfCy1oClFuNxA4QDqlktNQLcR4MejMboAp+atpod3nqLi3X/1rISEYeJGHzd6/HFnhT8b4lz2
7POui0Cy0sZYMJ2lismwGR47UQCijwjptbO+PyadaWjCdNxzFM0FDE5XOSgybqiC9hyjr8Wn5Jev
ocmxWsLm92TCFNeRZeDzt++QmmaTvGkCb9e70k4F0alPwB0eRLpwZ6uyLGN5IlXBl9/834jxmDHI
YYHCI9A0Obomvbv//CelrExQWu184KeaiBiiihZQVw1c6sf5KTd1Gpx10s0b3UnKt/t1xFLkR1AL
3zuHOSRZtYO/1M2jq15ZHhTB+Bsma/Pj5no1UkNCzv/da+LzDMwRFtlxqRxWoCFnDXH5xj29fHIB
1FW3bfRPAmWje3dt6yCYHnE8mBCLyaDcISpI6rS4dqRut1xHL/z/dC12ZmAwF+HO6zbVh9NBKYhZ
wewttDOIFoFEFW0Ai0S449519eq4XsPj6dtSl2FLQcUpqUw8hDQWPhBAScUYGUwgtpU9YpOrHpf9
QJeQihXTe8zFClxGvna07IY/ww0MyDYc2koHybMMo6pSJw3r03dohNXUlloOyJRrh8Mwd4hVcuqn
g9XkGllFIGP+Y0uT3E5urBpAhz6qA0cT/V5R/4G8er4xX8a9NxfMFHSnxCFDWKjx+JQnIGQ6Yi/X
Lup4sQqFTv7Q1md3PAZ08n6/DWLVNtMvOv46GRbMoXLNyHuTMaUspJL9DqcjF0uQ6u9UySzReL1J
k8ae9a0Qt2NJXWO6r21yxqKChcFh7jDqyXbaOYYeN05Z718NzGjutBFscPvyMI1K++w7POnOGI1V
z5E+YS1mbX394YuUjtqyCtyy71fiCzysOOjZCtz1wMkPS+iqWoaiKUjQkLGx+hdzgnyUQHQbemOs
oTNnjHRrpIkNDMZNSNfWZgfIu63WJwt5k+U/eoayCsgIK+QY0oG5awSLLiTliFK3AiLTIFtl3yT1
ArmdTSYu+hDXESL/3EM9kkSwmFs1OO3gvJUeBjGxWNstKZpbskiCzXMp5IZeHxupOr74axEnaP9s
xiFT78NHI7mNZvvlYGXdckJTO08QY8GHUCAqw9IJzOjWX3FaB615GHvxBnNNGUI93A0t3Cm9+X/q
3p1qoLUUvZEgCQPiZtpHufRgPNA+vXTOPbhsMpeTnwl9peSwD4RTIA+IafWMTD8PyX/SPlGyWzCv
kCGc2t6oiONSwwgoMDu9IV/uc+a3htu/l6FNYcI7bihKjdi3Ujpqe3UW+oIPA40TEjdCKKFKS8fp
QecXsULY7keg/QbGFec232k+GWle7oGrDqqYLR3XJNgoHsRTaeE1WAnXkBLjj8js4Eoas8vc2hWl
or1yrq/fxb5E14FOHLYLk82baUHGUNwe5fRgM/vBXuhV7QXtUEosqWS6OxKocQReHd2pEmS4e+an
n80K9yaeCrfKqbbc2NZt7ADcASkcPzzLTOIM7klYuobuIAW1mFKRfmEqhiJpdmueYJIhKDnu3l65
Q3XBA0mKLAz7l3BjjJbFjON6fl7EPnYrtCo+UMZ+Z7Bs6DiodObvMIKqCieQrZV94QBDCepVw/Kq
BsWINIWmsgxKFZam1ONDMKHRrfyidNb8fRmoRt8a8JULVb2FBNzweHC1eoU8a9+FapQVOmHTaNrx
T+bQfXbcItpWf/3uWW3DLHsl/rR8o6MtsNtuuwzqZjEWYgLf1GdUi92IueVIqcyCqI+hMS/WdeOe
ymcX5Lke7+PdXCbkS69i/92JsogxBGRJJFCJ/tKQSwSfnMLcKVwKNt6AJxN481ckvLmaKhrXgn9s
bclSa9IwPIazIRznmclBNOR+6LYWD3uZM8EaNm57MFd0hb1q+zIN5EUTIInWK7MFvethPJ1Z8Zhr
pdZLkbybWF9PzYVzYtRZuEVrR2BJR6H6rOMx/QzKX56LH7ELeYhSFALLxQVLu23J202eaOG9BC7A
+8s349OQQ4Y8QZfRh4Nz/SoD9bj3Y7d/wzDwp6iGdxxLuvOvzwPKjKqCBTa7FrTF6hPji9NV8Qa9
2g5EluyfjXXismEkjasVqawHuAHVIja69uqVMoy7ephNR4duUtgJfzOh05zmvNRJeG0gtZya764O
wSmvuEXxRbn4hzQxchc4319aPGhrqlifwPcpKMKHvWdDAWQH7mLwp8NZ6AK5qWDtPddUzZt6gziL
srk8JXXVaqE7V0qIJ7irD+lMQ+RBLTCgVo0xLej0IlsuYW3+mfUViU07vmW6XvkXtol3YLefuAS9
GarsR+KnZ9KR71zk5DQVRt3YROTfqSS/sS/cimnHgwt8NzJJImXqxFo3k+JiNM1Mw/kTGFxm/TAd
I023tPbLq/AQIkm24k2Vd92WMqdeiJjzVHS+vas/vERuKRzxylUJOy0e0lIkZiE0j11Xrf2Fp3+U
b34mlu/uS5lS3rGVNJJd1nhTglrjsnf84A/2kW1AmDMdFPfmsnIx0Y9SW6ctPhvuMIU4G31ywrQZ
zGrpDcmHZamPgNI8l8ME5RbBp1QFqkHetcTu+ld97fJqWu53UAlliUovVL4+42+Zsk5l7YEap7uZ
W+ov3o7b9KEPCKmAWwnxGBfphi3EIerPqeJKtz2xqoFiuqVKa0dkUZ6Bgj4rzYAWlq3HuKR5Se53
OqyfmDimExAQdIUhkWYaFY7/mHnrKLss28aXeuWu0jjjaCO/uumudPKMs48HVbM3rP/RWU6CH09D
Th6aPglHt/QFqoZC5bTWWClb8gyvCPRyP5SLg7OLR0q6iqG8tWd6XJPccj3I1RRWOeYMFPQe8dtV
YeOjNaiRzc5PT9KLZnlwQZn5RhTb0IcYpwRYC/39Iw6Si5gRatlofqFmM1eR0E28iDF80h2aQi13
imYgm74rPKMeTz3kpm6j8qlgUV0vObw3GmMEqB3V4D//PCWLhSa4/7ZXX6FevtUSxNSj6LRb0zrb
ifH4/piPK3Uxo0jUXY3GrWl0vhp0/WYEYzVqRWxItWUU+qe5FvPCngQW590b85GQRSgBfTyV/o5X
RVV1dyZqAbrDRlTetVWtHJ/2sARYCWfWNIPeozm8hMDxZ+FrS5ZKfJuTHyvtYM2d6i3TqKKjIOwu
qxjOramlhygwZrqF3lbSqD4uRcw5oSwsyrVgpLNlB+nMiLGXH/FhP35ApoIyvmVyEOM1R6HF49+M
aEYrkgfBn8LkHh79Oxf3Y5/iKf98TmBHxdgmX2l2XxWgdGOsWNJSpnPNVChbHi8+IlwLy7ds1Ehs
jascWdsOUx3+twZUx5dLVL8j5KKa/aHUFHfdR5mdgK+anJAoHock2TpOBs+A/ThbS9heeZw5whwr
f0Z2Gg+q2u00n3blj0UPjnk86qieE685/MBnpH5YaQ9gm7Mko5kgfcq2kZ9CXJtb7Jw47G5pdpsA
s2okn+fGlEjDjbaDnjCRFXQsyneFXPWeVsxa7mgORcRKV6wBHHbWXrfTZupk/ZzTnukZUH1NGuDx
1iJMXuYj8bpVgsALFt+l5aSm6CayVzUs+OcOXGUsFJ2SxxG8RgTOqSfZae0+oQ3DPVPSI3t3eVL4
6qWjKwOQsh4BVHZCBLuSt1Z6qQpae5o7a0p3oh8te5KKAu97q33gsuHitvyevWIxgEsnBCkbhQBG
Xl/XJR4vPvG8587XUJyIse/2MDwWzk6G5Tbo2mfc+lH5w7XcebOHjAhJdkPQ3fTOUWhKcpLcYsz9
7l+uZQNw7/4LHAJLyoRMUomq9cccB3NZSO70PHDU5aZW0VCPegItwJNVSOWVcZJQ03LvN+p5YeJ+
AABy34U4anRINSgyhnkP3QmVX5Uf8V3tP+OijhaemKk4yvl+GXHBnBj0Nzhp1r1OXbRh6Zbex8Zh
EcgDfcCygIj7vBjT3QXwWehj1Ux9dwgD93H1k+bTvWxadCUdOMKDXWBfVdum8+sI4MdS7Uv27HAz
FJAtLbNbex1goAJVX5XC/lGEF8o75vgQh9mGP47BTvfXYAc9vp5WwRRQxhxZmUPLSwB41ft5vL9E
1i3/Vn8rsBWAqwcxZSre0Q6DqKpRCGZrS00te5DQs/+v2DRg3+48gybNahLDfZotn9OAyDbgda0S
TJZ48DVE22wUslFK1hSp6y22769NKEmbtlIzFfedVdrhlD8NF0vCmYvHJUbTI9WmDnmtjRV0nA8G
I4l+3Ejpv5p0lo1EOiTqyo+E/cvgWaQPxJsZSA+cqTWsKtIZrpzlnFcLCMNhtYOgVqw39QTJ6i/y
g4stp2pUPUJlrDwTovVn9XrpTBomMRpKTGQchdtlVuze/gUv+ulXe4XOdEo8yA69uGwdx1IOOI5J
srZKcgdwrU2znJQQrDUvg3MTWSUv5TbAkfvktV7mmYK++LFFEA8DK4iyAFtQkD7Y44vLKM+BRL2Y
5N2SfwPQtnDr6HTL+8ub1CgZUpeMvsrLH1dHfUBAB8faCTg2+nZdGDtWnzVtW+/YwWStkCGNkdwz
CDgdjakGub7bHDrNfZ1a9l0J52TC5wseTPPkBq5dBvdsNiMGm9A5RWTMqDzSl+8v4W7TFqAECXSd
J9uREeQaxgwNigllZ4asQv1ghnBLtelpGBO8Nn7lxh0kc8FY+lWM6UJmlLTrwtDN+e3IqzpClu5v
eJqBr61X8mDn2VUOXNApkT2NR0Em1zZFIU3Sxp2OG4d5wYil+nxytdgHwOfinCorKZtQaGsL0j5J
ztO6b2oJKsVU28Vn5S0w+d62QMKlQkoFtrJ8mp2swrjNHhIya6rK2T1xGADxSZD/q8TYGL3PShHq
JcSUZeDIDkW1LwvatgYaaPjg2uUYhZUi9wrW4k0fD+iFe+47TBXDPA3fBAAE7M1/P84bh0IAAhKX
KbrOl0Ric7z27bdXeLGinH6W7h/c+59QBk5b3PUdtDoLNS8OCi/mBljVePnr/l8LuA+yymhpDAoU
3Ygu2R4xfM2ydA0hA2sEGrCi0Rzm+DRQxvFJP9xI3OaYuFz9PUJNLcmkqH2cXFR86kA8LugLnhtM
35/bSj498adwh/kws6Xh05azAFccauo6TQXXwJWBYnm5fyxjQpIOSFDF9Jc/9f+YrfZYLr41t3g6
Bm+CdpaJjsn+f7FXnkMTYDRWZgTg/8T3enUEGacn8hURs6Em5G21VtPoGVvGEY24GuxaxusGKFMQ
EhCoEOZe4Jxmdh4oCJRmg7Xjb3heVfxbvrNa4gKLlDC3f56mHf8WT+010+vcXAhTT3+lU10WOhZD
3Vwn2ZnkCV4jeg7Uztlv1IRr75+JLlyBHPvH1ZHgj7qwmrUk7jwcGCvXNkHgkjwhdfXsWPY4hy3S
BvX//ILfgq7tzPvFh92yjCqO0fbT6UdHxuQDS7pXU8TXUeMND0WDAq/mqr2GyH3k/q37BVXV2bdl
G1AYP5D3W3o2501AwIN4T3Zia4H+/eRzi6FNOtlui4rukdmh8GZS8yQzYThZZ38XU2j5DZslv5Z5
ggjlm2zxcw1hJAFbtIjYknU/VVJJ/Jcl8inkYYo6xLKNlGWnK37V0AKBLWx/rcX0HwEY2INl8Zjc
Hvpy+V5FDetnkWXle9O32MsKeBobQzBnx0fcWci2ZQ97uIazMTh2xLRubgSJeAcbBa2FI45eV/t7
mIdcjFQN7PuhYheAvuZ/5Hq0yz64OxCBfaQFxb5xu8qa+0p6ViWscWBz/tWzd+K6vANBokOwFpmi
0Z9/Z5EYsOHlYRt9uIxsHrVWWdj0tOoCUYawwG8KHBNg4GuQTyv/O1n4JEzTl7KPGtJl2fsuXAI6
/LMcz+hrzBBJaGSoV+QYYkeiWj182MfV8YKQyBAyC/U9/nyjtYGvaxY3svmX0iSm1O9eQv3YS3te
np5CWydjHJqRj2eGVQhnbAoyX1E3fguZT5fpHqZuVdlQw3CLiyrRZd2vFtjsPE6SD/1tJL1ZkcjQ
PM7uxfGJxj1EI9JK7v7tQemCHACAqIcppXFhna8+HzfNyRY288P8cFX7HIBuV9tLOO6YPrgXJ8LK
BZztK8cthXu/7udELd8Y/D4cPYut6ASbha/7g3PBtd3DalelyuUHcs+eogaEwSdSsYutsDqQk7Ly
KKha0kA1mT54Ga6xrG/VAuwtO+VHqXoQK2qWGMjUnNXpm9lrnSmg2zKaORcty0k6pqGjVKBrLUJN
IqrJTVw4TIg+HjYG/TRhpekA57NL8Fy4M7kuGaUBSyllciO2H4p1cj7HHJHS9uRMCzBX485nvr/1
3LsTqXMdM/RSL8NlofWo0/op1KoH+y79FJv11D7mFMY1URovKU5m5/gOH/mUvZ/ZC6StMB5WA6NW
vWRRXbfNTqE7e//7nLQl3rZBV7nt0+Vi3aljlnnC5a3kWLiazAkRqAfHlqYAgH3bHhyBzjtJvnaC
XWffe+2m5iWQj2YRL427apIh1LL8Sp0ve17UrUAj+lFVDeOmMWfQAtTfOHKy8tpX/0WnuIFYwrg1
uDHrzUvgcKOtFJZVd/MaAZohOoReWEOsqKeXwKmW0gmuHO86mjFQ38d/ugXOK5YYZHITL8V5JVCh
O7qVPu4D4d0Mn+KtBXSMwgSsSM73YamnYMueyuURVeD28qU4KOXcnHGhlkzY7yC0ZIJNmiYXwrxJ
DT9qHKbNpDrLLWK15QtZiISM59Nx8lG8sK/Kt5Q50xTjlkXjELwB/+I6ijsY4DIEDDzbC61kasDG
//hhZGVQ+eXGkmD0dtMYbIfQMzHkA0OqFLmJJbZZlR1clIjYjwIsx7WwQsDhk+F/StWROtzIkDaV
c0fej7fuut1NOavNcbg1PFxUoZQObops6J3MpDUU7OSme9COdGgawBVQ8Kr2gzCwTfAROS8RdZ+z
vk+lMU6D/h9YFKxme0v9gPc5/KP4fDc4I9w0OSPcE0rfZoXPIrtScQhGLcCJkHWq5Vi0aD3saT3V
APxxxHSg7Rhssq1K6fC1Vz3ihGm4i3fExFHCrEt8WTE1seSBYea6J8BPlcdd+WVczME9JxQ/Pzjj
VNMz/olQRci1xqQjxOwDLB4a04qQpzZBZ9jWZnmCXFeck1OMlLDSPr5kQODMmxP+CFThOglKSp7P
3tmelBdLUFE6HNuiEa60nS/19/GCVtiavmWGAmuT/nwQB6lX/eYOLMOKunBq2R6K+M/pnAQMeY8w
/PXK2cal+ePlnFoaoZ/R0P+b5Mmn9OX5RvMH2wSLfvUJM1aywKfema+adEfVfxZNqXuYgLX4dnUb
+vw1bSkWPC9qDlewXuwT+dV6oKJk2DzrdcMOmUkIrqqvE1Qjwy0XEbiMn1/uGCvr+utvvSiafrN7
AdzgyUt/FuAIFqWsXDWB8uvD+pe6gNUuyeSOiAVDUT9c9KniLLzfgQPvJqd7okvxo2geKdvjsXQH
B0B4wR/DCRQPlmC841ZIaiJwn9w8yaY1bdX5gcpYMUyrbsoYga4ZnERLTIDsasW45e40oxX9oATk
CFV80ZDMHSpubuJ0yV+VJQIJzfw2F1J129RHhPZGoweS3qj8GtEQeEqwcHvblpZTdk1eg48GlU/x
ljU1Jhf+VBk+LzW9+nkVxNziY6774W1SfjNILOry3qhfgKnfuv8/2SZSmhHM6GInaus/ZRhm/7AN
xtU2odCYj5k4X7udS7AMhuF8bV+vgVGMNCCqOkT9ES3M6Qk09Z4rolPFq9kBBboZBMXK3Q+8yxFl
okOc4XoIkXnBrPBdBDXey3f7YC/C703L02YKBXjOrWe/irzZxGtrGVQMRFkLWAjhCtRveDH9qQzv
DNNbcRpf+XK8Tdj271QxiW1DhjwDO09U4F0lt5+nGyIbBdl3Zggia8f1TnSSbqrSM3tH6Zng8mA1
7xbZN6LFTSfdxQbc8ycg8VbTLQZxSF+SRSn7jvMwIXEg2cWKm5vT1bcYzTKlwEX0jQtNEbQXhD/v
kUnkhWTKtVfQExnvKokdc05hpFDijVUK1NdJpVmj03xRygMu+an3HnyAQtVmP34Isptt4J0726m6
qFQF7SbQ2xI7j+VOsZKLvIU87fQC/uJNrc6xVLUV5wmsZd8g63LIjCJnkikE0KVx33YjI3rcK1Nz
F3R5jY/xfHZJkUTjZkL2mVeHqI6uTIZuiu0OuqgfhYnKjNsEW21eAplSIBM4tqbWTRLFoDROZoUR
EHEVCLkz1ZHL8Wgy0WSv6cdo1xEas7ucifWTX2Xd6i6ZfsYf9WmFKnsJ/FRh/FbCnZAdm+btf7xP
u7CfydAwzHfvlkoMW+Smr7ctXKK2T0Y4C+4Bo1b5gfpuHAyk+VZdpAg+SANalpf2Tf4GYzt525kz
Qrkji8t1na7Ju94nIM2N1oMmKTvOK8pSkl9/Iadnfw0uT1L1XLy8VxcWKUjaNe+sq0aA5CKDawqF
4hjcEAorS9xz2txnMtr/iGgIWx8RnS1vC4PIDawMfBtvw2uP2/OqEZ23Uf87QGCFOfsAHwUoBPOu
UWHLbGSoB49o/ivXT9aeAYPVOWW5mCO/T1Py5FgRNSA5D2kooaFNFdMVTK8piKD79nu7+JERqDEw
CLfAl80WOiEYL6/Lytm2FcjH4SnIMVKDIzVALK+IjE92KG4IRLChdXqEpjz6OTKEzFPgJIbXkUeK
ScHUFFeCWO2IvQLmIARUjWNIIlEbEvKnQat1PHVH1MeJWB+Btp40t6XWAlIEDyGR8Oe9p1vjbsLH
t5Sc6mgx5YUuUx8WXhysjkLDSh6UwsilOrl4Yt5Cf1TKQbOF3BffK3sOvDeejS1r53vUjqOMlPQX
AUq1nlTD5OGHolH3iS+S3aK94X/Mpz0whaLtQFnmmY0rV0CeNFz/Z7yJXwjzIjl0Ycv9iyxqnF6+
YryvQDuvk/AwLiMq9/AS+3DuHanBpE6F4Uw7Z5IdUlXYWwnSX/6UTFLVwQOrDX2LDvNuTOlMPXoY
rujOdUS1jM9oocxwwOp8bL2StCfUYKpQNjte6yS9p6iWGwFGaI0QyFdoBdh2B2YJiGkxqJUWYxZb
IhiLzQd6dYm5GAHx1Cws+0I1rZ6ged0MncRbBg3rTEBZDFYNelY03Y7kaBOX7DY0QM1wWvq31O4g
RMo21FI/F1/gByBOpn4wii6mCJQorXU8tu7ne1WbtSiqhIECaH3YjQcBowdc2eNJ5uovZR7blaqv
0CSpObbaAzJL+WWcj2/DiD2LywFqZ1g+vmb8485NIKla7rXGMQkYoX5xfXa2mUPi2Ltot6wpbZ3k
YLRVHErpN/JInA8IbS3gpvOcQBlSQvdBaikzb3EwmHrIoZ6requXyNBFYGcyLlP0NMngCL2eNVHT
uJSS90qR2wBzDhwufWGE/B1d2LxvYfrbq8YOS0nMlDLUYDh057c7sdJ+0EkLzhYFvVgxhw++kFeU
dFpk551tXn+UmJf72lGqAkycYSUXwgcF16OBBrfUZxSWqiaKGv1XOF7VHZiCndFk01ET61YSzgLL
QgNCYP8AYjWQ6J1Ds81mdKAAoxq/IizIYQcF/eayE0XN2YlC+3hQNimIe6x49YvwZu9pNRv253Oq
WDylqQVoVfXuE/ZGUC3Qr8CEG3zxIcHZ3g5sAXpIIi6wtEhXxqrC7MVV7nuTIbpKU4LPnWz+2uAD
uR3BALB3MkR20DUjAQuuB3EydXr18SD6vNnCn5CaD7fWGy7G7VialaaZEOZUAAISKPPOKQXtF6lg
kZ/SdAZD5CJLgPRCpkJkoJ8S0Kk/z/tEw8OyPwCga+dcZk8u3cvezX6iGZ5HTCApMVA2+8c93FRz
6dUq8ggKNuAwLnGsWP4Je5cB6tbALwtW/SoHUh9WW60rqgHKed8xUfuJ9Pwqt9xdn0qKP+GzC/Ay
pXsksAK6mw/Ow2B+36eAYPmuPlYVHHhaxTtiKETlKy9JqmPMY5IN97C0NCWl93qgZZG/dSqrUWZ5
oNfhaqEacJ2X7T3IgK+UltmNlYF89tbVH55G9WIIvDi2Pw2B35fKgfqIP77uo9156JOSNB1xJP5P
GRXgUppfopI+Ni7q1OwIG1C6303AKHD2dLYr2USdAENfF5HEAloCePsMmsgUHA9PJ/aHtTNS5wQ6
okDuhw+JofFTeih41DwMFswyiMZu/fxeiOxXeM3LvQJyyfQIudzmtLwz08H+EiCOmj6Xt3lZhszu
DWVqWaj7GP8edSPN1wK9OkJMIZEJwMDlNOnq6fF7gStLQUoCWKhKOqDp9usgf1GyFJKVfsZnxPhg
p40GnjJAvx28xXqaDjOJPOv/YwT/fK1rRSuA0t5umu5nii/JjIfueacbT/jIoTPWzFKv9nq3OB+A
y9CHf15/Ag+4TgGZhWLfSW85YkcxNSOi7k/cwN8VjXAybj5LvHtorrB9LCI6NKay+1aAZ0MLA00k
19NcEQtYWniY3Ge0Z/QbtsVnTB4NdHEf6L77rThxWpzaHeLgia0g2keCeQTLewgo+cTu2sG26T2f
JNF7muMzJZEZ7iKhalIH4/YnhULqpwHAfcMqo/A8dhIIKutyHagToR90VQmilEWdMkbJdHZQyNIF
FiYoLso0r/NxE9TezxnpINpLvJl9l6jP2VTwMT/z8B+9+J/T4RWVPjLwwKeDWFG4KU/ZVGwKRBMY
K+jY+TAxKHYiASigE3mxI54FiDw3Q6LBw+PclH54An+5WUUjx6Lfrpt955BHdNBoZz+w7feBSGqB
dSueuyGO4ugWod6uKdZ+miiGU0cLLO/Z4eN+Y5AILBFWTs10LtGIASb5/APPPFdFK5k9eSAvnSUH
nvNiEfK9GHmJkoisbwCC97bNiF8h5nWEgx22gkNY/WGDB7X+qh6llk+sFiY9BPyqWvaHi3SkzNGY
53bJXwns6HHZgU9XKWIDi3+qbNnI9bUcFTwPOPHKZxlMY5GS5rlFwxxZu05eiBZdLI5/X8KEi4RJ
RhhIY2ZJLlypLFCFgeoy6bV9mykdvODB1unNXoQPW3TQvHoqRyR/LKJKwbBfJlnmQUXkqdjan+bs
F2tAweIYDr+VnpQKKBTwvmpZ+8InQ6BtCpWgDhvmNaDehRNsS57CBZHJN4/SnaDZndIRUOt0ovAE
z+iNmc8Aq9uIR+F6Mv1A9wLeoKX16vMc4xb7ekahH9mKeAAHKgGM0fWPQylX9x612Ak8vpXNphhY
q2bztjZoS+iJVzaNWfEfsnnQBqzLF81q5dpCBGGmb6VcNzVDkFrfROS6+5F+86+n2/Zi6xepdgOO
V0v/u7BhwPkOAOfVJ2MzVTcNNgCt3Ep4TmPFjZCCK5cwDVpBO9Uj/rj0SKui1JgMNQtikwTDNVDp
3vCucpAToUxe1FcyvZjvMLFDkbMTPBmSc2OaNxxEBmL2yP53wuWtrbHrdEUyidui5gC8RNAD2oix
tpQkvQLyGc6PeiO4pzv/IIS2F8GWfkJ+t1i7EhVrrJM4VGHoU++OdqwZC3BWXL9fV+kMnJoVZLsQ
YJtidu/QOuR+nOsqzS6lqPaB5s3xuw47V3xY466PMz7esPV6BQiSd95QATWe01FfxIucVtHMATAO
ES7OnS5NCIbOcF6TFKFkyvXEMKcZBGTpTSZc5rzGS4F6D6zaTMRAA7Ne53XHUUWE+KuF2mjGuSu/
3ha0+xpfE5Rlxk7KnNpS2zTp5BanJPLwTjLnhqyYVZM7eeaytgwZoiv7ukfcAoELGjmybSi1q5jr
hF2JFhil71xOWgVtMAeYg0s1G5ZjYWAWS0r4gm47WZbR0ZsCpmU63eGPkCTBSE8R+ilO49qfvnWm
T+KxFE3M7BXorsq2Ft1SBVAgsmObdkBL6fG3EGBdHghsb/YpgK7bOpqlFByKP8iJL2QryCXGWGqM
c3xjUzSB/8D9PNqNYBLMKnExHsp0FwAjX19wYj0qE0wGW2ftUrOJjoql2ey8D6xXskkon7mMYPJv
VmecDdLXLLXFbIdPCiN42EOdc6KAWMM+xSxgPYXQBD0tcJWFoPxbS0Qotma1G7Wr1/1+nH3ATJjt
NtgiQN3coQUl1BJlXcWAkYmfhYNZcgpuG9rX0lMh05FTmNFKI35WxpyTjfcAey9nCLgdanWP/bXA
9sGMJ4ok64OZfmHSkRbY2J4L8BCvuvKWwhAoJSSYp5QY2gINCkhytYn/HZp8dQmEE0k+ceOCGU4y
Snj71enqQT38JKPj7h34csayBI6LT2e75wVxKAwww5DAIri5xsPF87DlLSW1vMzQ9HboeACN9lLD
uxeyGVZuOWcHQFrCyalmce+E198cffbpDfdkoZYTRzDDjqAk9qOlnRzboQ9Onk0tRWOMb4tzacQM
kGj44rmwf4V6/g2EtqYrD6TRKJMmb5FMfRPGJJv5GwMQ+rvAsU39sCI2oDvSBWUuZREuUFs5wch6
HmpdBtN9fbh44SuZTorjP7yXAu7COfNs2QzbRBbJY1pOBRlBSBubTd4jAK78la5D3vZDxXBH3jQQ
JXhuEM8007Z4j95aQwusLQE+3TqQElv8zOO2qXdL1mGZG/7drjGf0L//JBBTTOvxG8VBSMbOsF+5
M8lSgjFm3wJRZbBgdnd+QzNdXFBdTLzwdIsHqAkqNAg8y9pROubo8UKPzUw4NpRpdB+F+tHGrxDa
+ktpytCfHvaqRiG9/yfLP+q6Gc2uuB57wPnWT8KH4DT4Byeaqez40z1VkrqmndOlRb7dPJWoD5pz
2MqjPzFMczRBok47vA9OVoKdXk3VI8rceuM1zLLjSAGpo915Vh0mEr9Ascq2ev0B8T3y7sB+BJ/m
X7Y2UeZY9EcArphoDR+0s90MTj+J2kNDY2vlg/Ch5g1dYlTXVoPa+nRZARE7nYIiuAOshaa0wk5O
0kQ5fl39iJYGJbz444q1KYoxxR0dJ5tAmY2QksvHFbKWevl2A6a0/cZoBNWzVb8qsurLBlIJ0PHK
KtGrgd6Xe/gkKEdk4KkvXGyZDcsqTr/SIqTUFbTPXTYhnpQpSFjSlkiP+U8egwUrggqo6L8EH+u+
RR/Sh6mcn2dmTtxJVznjUK2X7qaNrvG4n1fNa0C1gUnIMuYrcXd+ASXObgwcOOOR3OUdW3gn9Nwq
lkx8CaQ/19anUXeT+UJXcaZUs8zQxMcEbcqbfSxFHEHyTJOTjkR+0ZYNADRaa5/BDF8OkdngX0N8
b/MstGCwZyCUGQCH0uruOLrL++DtITY0Kk1n5cdt/Jwv67zvbl2fS8zvoM8zEBHgOsxava2HGKbF
sfIdYcuTL7WB3pXaHuc2dA/1d7iQ6i0EVkEjEr1xnB3GSeXG8GIrZIOoZuQPcNrNeJEtKx85/SF9
rzObpCASzwRfqUgxQGF16EFQiBj3cdXuIG4RrcOcXGQ6ZgWD0prwGNj5NVPzJenTiXx2835cK2Sf
eRCE3H7/f+pbvDsHT9uLIsJg2jTwyfRc4ny0uxphcLY5VdbFZ5pgFYM1+c9MG9SJ3x3Qh+gqYZQH
xxXA9LgjZb5Kp7phHBPgtzJKyo/p1lrcSF3mnhR6vriglLEfY3oo5q8o/QIqiitBVfB0ugNNp+SL
mHo6aHdkwMLzC0wxCxeMk1EhOWyB6GtdFt4zfa6Rf861hKrqeRHp4kWQQ+k6dPFmUjMeCcbg0tIR
M7qZseCzbtHKRnjYn5sLDLi7R2221lGcxO3S1t154WDU7+ttiSx6gZwaUOPn9qk5Zb6Tw+zE/B2n
GF5yhIl2Xm9jsnUcc5xmQBkHL3CxNSzOVFiS22VRjViNdA/Pa9IknAG+JW7oDNyJVbp1bdcXwSOw
lMr7dXENgKiQw6XZ8n1Ukt+IMgaML1ekEswtW4+I461QYg9X0HGOsYTmZp2q1fMK/CGmggdO2uql
we4d7IvSobSLzgAYpsTKESi8uU+RCf1P/Bu1lUMtk4em/Ilkszw2+tak8YLD+AMCGnN4PhRB7oF2
2jpKESIDU8zrs/Sv1pwo2Qr8kgzNhW/XQ/FPRmwF2EmcWr/ortFSN1ecftiqx62O/h605Gixj4rh
/IxNozLgPMFoAlpQkWaCENzFJsKuVB2XWyMM01VGUL0qPu6AdMUqwp43uiqqavooageZA1JU4e7x
g2yk+JXwOZoFzewmKzASiJDJx5/0Evw76lZ3DPk9awSJudsFfkI0EDqIZGw6DduFJy/WZYbFxF7m
0lpsiUt75HvzIcCztKbj0Lo6rz8XARnSkWp+iPVdZuOlM0IPhW4hJRAzMeKqSijFLJJy19fHUdXs
+09JeGL9BMKf2JYBzX9WFvgggiEvA+TWDHhGX5EV54VHOAChshSZRpY0HAsAnmgeqTY6TfnNjtBc
lh2KakB7hB2upYQ1Uw3uWKrq79ziwtk7yeHJRLgFulllLRqVqe7wspi1g92eRzJaidNqd0qYbQRu
17REnSZYUoM3joh8edCxS8ZJFwuDL8/9Ko+52kOvw/eyTLQXG8YhGogdp6AbM7WMA/mV8OzPKlxF
YPujM+d3a/ke+lxreM0ATpucl8I8UOTn/C8iNKNUqUhh/I/pC+r2R60jnnM+yWLMZtVURBToyGkA
0fa1c7DIKsqCE8NYXp9eW4mGnci4ZWTtdxSF34eznxMnr3P0L8Q3Gs6wtaHRA7djyTHxNQPmJWjz
FjQM+lF3ajCYWcsQq+KFtPyNiI4P6UzOCx8FTyiFu47kE9PZFHTvpd01uKDDwZ7Du6fRm0d2Vj1f
uXydOZKUVnZ+6ACb7YfK5ZFEZTRrHYsHx64rdhcr8jw6Y/p9V6x8Md6FXojLKpH/wfJHL7TqYXQJ
D5dx364bXgkfuenA4IMIYE3HL6Xo6sSViyzmX7TvnHwlfVrfPiNS3y+qqwmjFzqh6mw+Z0DAsvX/
Kq3XnaeX3s890Yt/Ys59EYD33t7zA0eIABJCJXu8i+ch+PvJw3ImFzglpsXAMyYp1Z2y/CnV65DL
0o3X6adFmDMrRDzw8XGB23QFsBv10letgL3QBnR3gdLthyOMjTtViHaP6zwROvXfe/sXeHoUWWOp
Z3MIWBG36LmDJ0n+7FXTIuppS+rUcZUXWVG3rJooBGDtKWqlnyZXvAUqt/tFeOOSJcop+ofTozJA
E3hYctVQXtL6nl+tyrjoEOr2I6FdIq6YbAKt03pVz+8NLHcjRWXJiGvoC7AwJDT/b1W56l9itgpZ
LvTtTKOz/lNtRMmYPuQoaaLj+j0wRB23OyWUXiTnOhpLOSI+/MDBweeBIn+KBBZFQfmj7rVNx916
IeSVdmJMlRmv20zDiOOpcSTECoc3jp0hWebgDGomTUeHBV28eWpT8pPW9eIfTNUxTFtx1defrPnU
vgnb19hu8RVZw4/Zx70DKWtGHCOf4Plcb+Il7ZJBoI34HLGAMW6SnSaMIBY7eXu7XXA3vmnmZX8m
sLgRsNfJy9NCTKlEhTGrXhvYfjl0Aah6PEQo0So9iWGhd/pChzpdz+dPAMp/BrrbkLphfTryAFl7
BMcGYFLU5eqJCI72+BabUrFjRlao8CFjql9oWL68MMoO5VqLeFgGR5Ka39zdAq3OX38z8bMqERYV
9jqeynWA9oWV6Gq+Nyvt5aW8jJaxOQabobg3R3/5cHjn3PNMhIMQZaO+PHZ1+02ko4owjO8i39U2
Sp24mtdhpPXviWkUeTI5ffjmQRAILZJvlkGBkrVeV/qCFshxbjhHrIvt6oxUi1Qav/YJxPDlm87D
+3Lehi7VLxPcGRXhekUjVNcZ+/Mx3Mdp+JfcX6NrjT0JHuQlkQ7z7S+WKDLf+SEpnJj7W3MeYwLw
0+WNDUFQ5f5MXsIA3wBckymrJd5EzAD2M+E3dIKlWyHniZKXuuXVXNNRYuO3hiZhJDyKhg5+0NS4
l/yCGJ0avc3tm9M0ao8yrdh0At82Sc3CAzOB4PdFe+yQQnvQr5Pa0I8b9sLC1HgJWk9zR7Fmwi0J
bpO6Muey6O294i4+sbZ8ZMMIdoXI45WuNfgyS08aqn0jXiaHQaMTrRc9GViZP31fHNSp2A3sQj+3
WKtuGMwHHtWBrpbBuT4YEUaVs+wTqhqOMX2CCo9MWnQdJSCokGcF3SkQGKxyy27G9J4FuAehoQTI
ABlREP/JKpz1d7/05TwlqewujMLvIkbn1dasTgDuCguPDbDlJElV7S6E3SUCiqH9ibysoNVy0g66
vAwb4VZQKpgIMG1kvflisM6zo6h+fGWOfneJkT4TgoBjMOe+YqKbgpqnqLNAx6uy6I7hTMBjrsMi
ZbbHNO/EXulMq9hMNynfAYi07DI3jCS4IrVkMblSt7IeyWXFO12eVv70voOLRFLTNiETN2dLuKpO
z2LIBhrEUZIn1WDOiQ3L48UV7L7NZPrAqaghESgAxcuPYeuA4G+mjIVBcSASZ6R4+e2KxVUonK5H
/GVbXQ4SVfc5J9bO4Lf7z7xRebFhjSXxJ3d26WzQeA9gnWcmcarneqoy+FZzOooAPj8zY32bpWIz
3DcHCLX0oaT9bZdD0BMV0pUsDzq4pWlemJmC1NvWl4J8m2m6Vonc74XBEnScStomZph7qKMs6sZs
1AHuHJICW96qVj+G06+rU+neDY9rqMabuyF61cjjfm5fhWU/jrLHji7X8c7sz47cf7xAr2HMgpiI
F5rYRewqkvR7Gg3pdZQahvD5ABczxZwKJ4GBVKHQrum90U9Zve6UKIgCjjbVNccW1ZqWI3rQ+/iB
V0ru1yZNZvXEB6357b/OiNDFtRdmmntVHic0JlidZfVjtfVFm8jAsi4IkRLSkaXXxDs9UDE55XXF
zSVF4fqjKzX26qoeirKvwHTe7x64YM6H8g1cqWZUjSP9RN9IvMg3HzTcW4/PBPNCLIrbxdHwwyfy
OcPrECuR2rE3irvSWL645nsDctSmyWPMmHVRv/uOXSRDueJjFgzUg8WqK7tiJA7cKX2Eo9ZTfBno
e2hJyeM3KTj4NK9X68hXAcL1hYXpX1vvuckuasHkw3rrUh60EqomM0Mxjmsb+mvofGo3Ulyp+Y1P
3A16iS2ZSDsC6DgNdCG5hh8QxBmmCPe0StT1nTwya8Eviz9QD8m9RqhmA/zKMNQVIs5GaawEcmXc
QtscBpoSJ/SAsr31MpqL78nThA60LijlwbMMhKC4FHUJ49WgtXLVtkHXdE0Gv9qJLnqMa0ixmhF+
PK4DBwobmf7UtFslSaolQ5wB/UpLXmiubGXmEaaG5x+dVMNpj8DRARl0ej8VjgnehKYP3f10UUVu
ucnVbl8wjfu2I55ljHkA1M2J3HSQdjbLDsNcTDHzljs1+2WxLkBcJZiPEJN256U7ZskXwKPNeUXY
GJ+At3gu1jUEaT8pylCwQ2t+i8zJftokJ5LKPxypV426BRWPbauVaR35ieebG+GEpCkUmVajcR1r
rgyXeEyOuv7fga1j1TWj0ER6xeZVH2QTZiMPbSmHjESMugfAncE8AOfBdbdB7QVFrJyfJTM3BXSq
BVL79Eg8ECCqCSCUND9Hu4cAdsEOEbwSy1avKYnBpwpwSuL8Ugtj6zWeqlMxVFu3XLdQ7YcUFMrS
LhkqqseXB/GgiHWNvFVTMLhi4CTFCX2ZfpjOP7HELnkBu9ERemo2M/5jP8vfcVyMHTAniJcBjJ4I
QWwkDcdEYEK3NCELX7v0PQHJVFB/CDl6UqwEwNAyiz9tpOfSbjWd3RkF6LdUvbkaSjUm8YSoLsPf
LDrxXNlxbrQr8VYPUjT8gviDarguHTu9Pd8PDCGGaNr/HbDlMsSRd5diPzce499j2/Nl2E94eQZW
/gPHgoVN3Ne0iFVx+QaiiFEIcKCmPrsaaqj56/Y+jaGKX51Vx7YFiCUGSl1xn3IW7R2kuSdrkXXH
AjNI8BoQQbbUL/VYctLthb13szAu3HzzkuHUQQgFx6NA30vDJCoPvrJGYsK/uoyth7gs1OY1qzx5
DmEyBe9q0wd4XRJKPSpF0K+dM9wlBxMuYxzPDoNUG/ANqieVE/pnmzzr33vPnRrU55pIAdNLzBuA
W0E3gBXKq7kzxXcixiVgHC9reZMGKzzJy5QEOoWiHCmxtNfSes3PtPoDgCcybuBOjFzIPlmTsNYO
QGJPDdeutMWKhQRnca7sH4vNdBIDHPYNvy2AtUUvztDV7D+TYZARV4ApLqIjp9TuMs3ry6te14TT
y3hEtb0DDDA4QrCuaY7/JCbXy6GliLNRROvPFpoeJ/xURI002XBfJCbEIQnew6W0xZdngO0MQVAq
ID9cmYTLmXvBpGYRi1th2DHK1puhUcgadGjH3JkPDsKi6oM7aIZAiwYeCdKRKzTPe/GIH2ujWXqn
CC0ioYdGAeDXrn3XQKcEK2pNQvfmk6+98zRAHywboSIExVFRHdu8qVaeMHT2er4/Ch7gAzwh5TjB
LmAAZlKI/sd8hPIMvQHOG0yl7/sE5DHfeFc4zawqXy7xqd/YOzXCEVw9bI3RDInyA+r6QvS1rATM
1FnNfa6y7Hb+NmfKZvdGxTkuNtbSpHew3DArPEKvIEIAQnzW/ziG8Bvs72+7FVV93Lr6wbS5cAXO
+0TKIDd8i7aiK5WR4P1sPZ8tuOth3CDQXa3n1AXbmzhiKcNJISuAPXnvFAGVw4sDf6Gut0UAXN8H
1Wial/97P7IeEDbb3vWMBGgjI9DaSNsXb+NiWdvAQybS3KbSra2uvLHYB0UMEqSpX5udh8/eYNq7
WB2wF4RvL58X4rhNlgK69qKv4OvocY4LXy6DQTfIkz6RuYCAib2DKBZvHaE66YzhjePp3d6veYjj
HjOcuqfDhjRGw/B09dIYGl9G+TH7Xn+UiB7SM8o564GQNNHlaBOIVMsI8+oS2mnxAYt6vUjCKtqr
jiRvHQQaBQpCPi5z5DM398Uq8AeqcDWI9vl/Fj9yiikmflBdUwDYJ+Vq34IzyT5kGye++VsGJW2N
aI8iqBLjscD9vWL+UKvQc8GVAAATMMtOoYLi7FlyDPIIZKluBjwfdFbHBDlJCEjx8RWQBlTy3L4Q
nH1ZkKqVd5wAT8ZiVoNO1EmWWu4254j/TXyRs8CctBa3ZKfrWAUeEBIw7dE605aeGfEwAjwVc1uX
9w1MQeMEcXr8+qGl9ojS7mQsRX70K6SCsQWO+S8zphlmT6+72gnC9auUtOi5PEqnbw2LvVdWZW/4
G7HdUrUsTztJaOWNzDO4YSp/hAjeE3oivD0cveYV0e5s3P9C8OYouSu7coJlvcc1zKXed43Ioxyv
htDaplHl7lRlVvE7VbPc0StCL9mQ2UDcY+4ezTibSeZ4zhz5v+p4JJUAqv4zqF+54fx7KtGp9Dlg
N8+rjimzzxp1wH9JHkVV/AInD4Q+Q/KWZP/ygCuvOyfgvCvxfS7613/Y8lSQQI48wmi6O3H/DcTE
Coj/v3DHpnfwtTOhOjDM3lDJpfHwbRL9RkfnQ4S+1JI0a087YhGLxbPwbAw2CMt7qDWdyszMv6cm
4DWf4DL/xalVnfYgyqjpIu+FecEoeI2XdTLMzG68S1iGN0wK42nfuufH8v5XjtthEl8EGuL+cC8u
p7EnXqT5I2UfQ0leP/QZuboa7ldiCMmkigZqahBgpsUzvcLfALgv1unfmlgoWEuOwbU8mucII5pd
tWwM+bH9DoDrLDSlIwwBN/jNZqZgqW8sF26m0LINu+dSaROQJ6X0ym3ylT66vdXQFKKXKyCyU8cM
gFzXsdS9aTT6UPUtna+tzLA1PhDj6l647hQ4GN5Za8eIF2/nIFgheaxcSWicCGi5FGwVxNjiwqyY
qpFvp43dp9MK2k3vzPTTtfzLsirH3N+RR2jYPw+eLlwb2U/+SyVqyw/di31Amx6ElVJzI7msn/Ys
H/Ike8/YfiGj4qx94a/utqdSNU0SUA3xWE/oSqUmfSjaIPgzHSwl7kchtbvRp/3kvo9IEDyAbbah
agdgyeWh1pZAvex5mp9lsdZJ/FwG7N5q7ZowejFTCLbaC7Ta2onZjqIntcvHTKbUR3pIYWr3NdnF
AnKBPvUUHKMDUy19Bk3PPdiYt8V3lGohIBCHQjqSLeixGKxJTRpTo3mXD4XQ27Clg9LZR2AEhO36
16woG7bWdZe5T+F5G1nsCRwKUhiukCOvCJ8NhBf1RQjoQaEtwUlVHBZf+H+TrJ3ihwwnMReFPtzS
klQ2i3HdGQKX819q+1kaiS+43YqD/JPE5xKANADGkNKisgn9RsUzOiS+yQKwayH2JuNWzYt0Yba9
0BE205qqb/Gynfv2dvTmqE+rgBzJD3KwtCuhkaeVcXX+1HQ5jC2Mx9lWxwiBqD9BpQORej3XCczf
rdeGBtGkaKWACREDbTLTL2X/OqzJnRCr5IDHRRMO0cz5wsxFcQA2AcgRMRxwZu0HGRcbDLseO38W
FZFRS340G6cVLJOV+PVQ9Fp1E+unUDpbw7o2uni4DlWrQCVxZDihJhTuGIOn9qkth/8HpXzNXpKn
QH7i9lea7uTCXgXvE8f1VoQi36XSA2cMgqH5BXpdDgVehT2j3NV+yh59iXTUl/x/o/hSM6NSSC3h
xUHbs+sEmyKFZOwcWqgyXmDCWe1kqdIBwPQV9J5aVAjiHTkMO3DETnST6b2gT3a0FmjCYiRrU/PA
8SqaFg2CXE6/ddmfzqbKam5EtVoB6hEJURADfpGXEdzu6W/ENC7zUq5VqB2ITCmDFsf3zKRo5toc
HRSr+5fA1bL/7SoQMnGnqt4eDIb6/sNaB+c/cYxH7eyrgL2GQ4bnmEHdbwp6X7pdJMSW7I8YD0W+
1CPIP9pMXeRj/9k/++WFG1HLC3HznkaYC6hrwVF+s3+G5/zRnmWaSDZXCqd/C3qfaAFBD0oan8pg
HMB1NQtMAN25yoPJQGcBtbe44cwFBEeGidC59mFgKOsuCMRejsDzjII6KUnMSHM9PLctXhnxdanB
9jYmbBbHpknowfuzL3t09Fv/LCplyr1AMvJ3ROk+Pm9khnZOxi4hfiSGBGzOVDKUwKzm1OXQXNZq
n3/lPGNqteyjmHbrBTgbflvkFwz4knc/ymWf6C1RSrjbsEOzpA2o6+6IzeIYBP7jMWOBygRX07pE
rMsDUKkPAscRRC0rG7zX7j36+Mx7QiB1qIgKgKVMg/GBu3GKrV9p1cH4/wAOlKrEDr017m1WmqF+
lCsv8tDlR15w3RfWbnYDu26bAEeFolvIk9nkjrNbRwFRaMH1cgtmTEC6gZRo+nz9MPc81TxqhfrI
MnagOKCkT66D0yTVp+nL/S0pFTzkb/ZigXzUNWzhVfxFgWb2y8yRxw6T2NmGZ9Er3XUXz0QABRyD
NyFbb9WQBUrkP76R9PsVsfugaVn5x8xdWI0+1J0lworthQyl36sgQk1Evl5d0NK7iiqDU+oEPQi1
NDacgn59ywnsrTBTV+150LU4MMvmCows3p9qb/8gDFijHPgFmbiBT4hIuWAXGF7V4h6JoSFVSVp4
uGtv3yPvpsfqP9mF+R87Qct8P7vkGiMswWVWUJdJ7MG/w/fxkMc4beYmKPvYZIi1nzbhlohQaeCe
nsv1UPbDAHkJPOlTv9muU6CW81FOHDo4S5AVI2m9AWP1lbT8+U5ZVcETL+GfzehWyNcXYxdMd1vD
7q6GIYYE5+V5bs8sqTM2er4m4A0CNuh+7h/dzDnZwywWrmwJ4+Ui1qV1XIw2ljgdZxg5r5NMVFYT
05R5DTBWiHv/1BjG4gtVhW61u1Q+yYgXgv8v3vUp2NezYmsw5kEZz55XHJIG2yGW/4Dv7JAXDK8n
rivXcmn28cGYaPrc5I3eP0Vx6YS5LFBjmqUjgBUSqVmwrwouSP5Gb2iTN0LoJOYfdC20Mvg3jr0X
bTuQW9vTo4pfo0gvfQoMiLqO1ObOW/Vfa0nTSRkHkGDGZhIv5iiVCL2X9CquN1s2eElnwFrf2bH7
9VAT2KHXwA68v2D7g6X7g820Y/Tfr79RSREo3rraZoZgpXrDSKpQSxtnFn+RJYTHMI2zr/yMKTL2
Zq7qHjLvP4lgs0br8zimZM0GO7U/qlIhKPBqNBDeZiLE/WNhcaUdCj1WU4jkkLqzv2haAxXwoc5e
QILkRPzcko1CWPLGcFMyKR+M0bDyBAEemDmcGOxxI6de0dCHGe3BANUrUgWTOKb9NmQrjHcfT+go
J0ZrTZor5EGEhr50rIxfNVIBAstj9pDbAuI2NQ95ZhSVn5q9ppnDSLG6CJk/O2+v85Cl6LWeDMU+
1H2Hw15zc2pwZNy6tSan/Y4H1wR36RtOo4rtOMDXqPDRRC90gmmTxailYRIv5SMEW9ovv0M5Eb2W
Bewcrdv7WGPfOKUj2/Rmb1VzcCcmWQSFPHJVIIT015+lgasMSA0OFJj24t/o2F/ju0WoefJ2wCD3
8FLWmEb8Zt1CFWg9kTr1ABZghc/NLS+Yd0Ds8ewbLdVkoU/qQkGBI9/fmpxhvxolvcwSJB839baK
oy8PL7RVR5lkKEw0cx49zi7ntshF3Z1sV3CSErUHxK9tmlIg2xyviVCy25/KKysxGqv3KfWa8hcL
hxWy9g9ZTCdf3t5HBfo2D5SZXbK2XnsIG7MijmWrf+8572XiZpmRFXnOPh8gJC7QqKW5ZAHAzLVU
LtYmkGkanxV3NhaEG1yvL2fBmKTqr6xQh6f7xtUjhS1nZcqYLZdcVprEU6xRvDGfZopAemKi0HDh
nrllGh5wKqILGJ9EFOt6JUvvfC2KV1er8gpZjfLF7a9HVHpsHzt91xdUOeAuwb9LL5Ionxg+HPU4
FmNkSi43OjD0wtGIXOvk2L+d8k7G3gAKLc9JmmVrcdjXAUE0K5zvXjro0Pm5xTRy1QeRQ+PNbJNZ
fQ/ydDEAdpc8IWUWEtI0FrqMEXhW/SKj/4fA9b1nAjeRUcukyxkh3NKE3GUPLfpNxEe8HEVYqR+Y
LJNoZwRC0AcEtsuRqAFjUhNQgFpA0b4IHCwMhhGvppYDlt3v2BUB/68h3J1N/TptrnjaMmlFmlDR
8JY9TVRv/9yN84s6YjBmcEx2pC9TpNPhs/imcCdb5SICEhTN+BUZV0qNLvYsBlKsDe8JNmIYMYWx
lfEeOvjMzI7TFoFwpwf63PdrdJK/uS+Kts4TqeYaAlZMf23P0ZqwOnjAyODqtbBT2qgxLchaOy3e
wuqDUNxUejyw+Ylra9JQksSD79snK9RpuPlVpoQS3aEJFZKTFQCjiUV3sCWdyyU6nnfGo3EAUPQ+
cwIycIp/ivfGw2ykFRGPcSI700xcNkjyv6Oxch9S9YyBLmH8Rwig846hv/lOAQ0GWMiN+te1L5Ll
c0HV0tzRO997cHZjFKvJtmxCdSxo4oKE77wJN0p5oG4bUfUUZTB8DpNlVXd1vuZf+KWvwo6gCQ+Z
mKMmPQUG3jIR4thEohtGbT/aLsZvHxa9rVqnx5XMk3kPKZGKhTxpTvCYM05edKv1Uyf4L5aj9x3T
pBhOEXRvR7N8zMHICCn36QjdMpFEoDzry6UYR4MnoZXdBgAVoW74/Fh+Itnr5s4tnKu7LWS5vuHM
NjG5elLI96Q8SEnR2FkOWvfr7ESPgqRJ1S7oaCxz04B14y530IzqGR2Xf2uu6HqNJ7gvZ/oOwE8l
BHGqYfKsF8vBNldbm7S+fOPiL/8Oe/+l7KpucOehwixNNgnXNF9wofvrLlY5W/654K3ldM4YBV0S
DDfE8hQCM0iXXPDJ4me+gWppu+XxXqcbYPPzSMsfX0UIrmHgLs94vY4QdHb0SumGbTxtMehN692L
kJWl8aooJnPcWoF2edzKM7pacYgrFU+tp2y5ZeCI7OzR6U4aE4v88LeEQTXmrZV7wZwPVv1w3RfS
51H/Vp9vERxigJuMDoz4oDIS9G3dkc1sqLo6/KDl3qwY01un3fgk02bg7NSIzaYViKP6BC8HSVCN
ZtqLAYVlzkef06aoYE50WbLTviy7p8ZoZyw6tvGPocAtNl7exQsRNR8sn7XYVBQafijuDonEy3Ao
f8aOC/GAIlnVSjtJ71O9Im3aTxeTHUACWMGTklYyGrFL5998TFxjXlODHSLRzktErln6MO3Ka9Kw
CJ7Mvf1zqIN0ewIBBUxw7GzH5/zZklBeucSBQe2ty5sFchEZn/3K6WQvz8DoAXUBIwdxkaLopSJo
9NHPSRIIYZ/qr1BNkSDHGyegLSqRTdUfrQ05r0RojDBsdXuHP7feRMdCBR2pzyixiwgNnl4AXY9r
oEt784cYgVcBCzIZhj1oEAVDVo7YzaEjvs0dLuruDUGdmGPmYZ1lk07XCLTKPsCOz7FOciFJPjuz
SpTuEmIbsBCxlwZtvaYnaiNCXT7v+0FZ1M6rkT3Bk/ZZUPntvpbPo0J+vmenQrbYEuVVjjG00Jyt
Y97aApSv2zO6KJgrXj2SE5GeS9buC4f16ymzu1AfLuTaGiQ3l3yMw/3T1UCk86yvnY8bf4HqtUiQ
GbZph7Vj1npJZy0Cbmem+i8wCW69X+rz1UiEhB5LdUlDJdXFN9Zi8vSKNS6Mmeaq5PMnPamnaXPF
kH6PDje0HKYqo8LTAWJvR+RM9H1umiJRjEwZ+7LwahZ/g+w5wK9ADL8V1T+3uSkYO137jefsP8RE
57Js2tdcX5eMr5mgcK2xymccRvQFJHKLF3aALXYjlifNmsNuD0OAoHfcDXJX1GWmLRYSduKmHyIq
XnPVvl7yOa8IYxDAxq9nTgFEnc9UrdV9+c2UXdMuEBlbyPujG+L+SlSBLGEI29uXDpS4zrQY9mds
vGvWuZQec8gDqoSGlcqiERaRjEOjTikmDNhJK/kk7Z4Uq/AP8TvHnK/7CAHKRcQYkp0Lfb+i+jzH
N3Hot3Bb/40uG2MBuPRyNCvug8DHiks7mtdNxd46hzzXulfPCNPpeE2bGWJlv+h5pFqzAo8jqI1u
nwkIhjvQVb0WjENg9vrfuvGI/8y/9uw2f2e9mpBc5CQiE5nGppQyiOuVbI++lmXoj4TaZMBbY9xN
q0Y/EdOS2eHg0+VWrv+fTNay2COqPqGhU8mJXXqnXevDFOOX5EVFUJ7WB4LpUJt4KyaZ6HPbYLWM
V3TIhviQcT6tLjXMvdgeIJyTyVd6EKEEb6fQJYhS4pHuIeXxeeeCpYGwL7UnsvyQVvMldnVlCaEb
HLgh740nF7/u4Hwi8SPpTm3aXR4+t/bXk0ghSO4c3j+yiNM7WDs9zLPPb4EwGTRTAQupE8Z9CRvm
j1EVziekA6UJQ9+BipNLbga26BMdvS/pm9NoTbT79o7EhUrt1UzfLlg+fetBxKmUwJcoPngoWgSL
0U04X71ZBAp3km8L+ZkSCb0eEM1+WtYDo0r1L0jttWIl34t5Zs0de3UxQfsovPldDU4/Xze9ihwd
f1SOqKuLw5cwVWNDFdUc7aDaWcv4zm9wyrbOoM2Eh8rotm9YNgxEM9AqDvOF1orfVBBmYFbKyJ8T
Rp2xnFw+aGxuvRTGp1PqMzxSqZPAd4a3jSlggzvFSAWoS23k/zaTqmVhnpFiwrwZokArWuyiY2Jc
bD+BQnI/QMzDWvfmuMFzrBkL4x35703JH559UPzFJCvMXIOWXSNYZJZPzk5DkNTcH95oR5eGUs0t
XuLrESYdqUo4bokzWxKLDwYLRkNb7TU2ie8GpqcGHDzmqEmZ8Z/kNtz7qMRqLDgoQvNtP7WUqDcx
IkU1GOS/5R/gIF8bLVx2e4BXnYRi7k+3Rdr46/amSz5rvyrd20xo6qCoZ/APT/O54EXR8A1gK1iF
dlSfgQZY4BymG0lWtaxCIzvIvHs3Nea70E9lA/pG4wn6g5k7T/qU/0oNwH0ZhX3Uiwasjy/MVsoP
fR2//ugQq3DP3wfOWvdXjCKdF+PrHugFa8+T/bWs3pzWskxDh6zj5ysU8PkVgMTOgI/hqO3prxKn
PQ3GbmT2bSCaZ1/0Za6NYhVxiYj1Fggv9aAApZh8TZSZV67oVmlExgrgT/t7Tthk4LZJeI2zZJxq
aKxJ4HAINxDpc1d6EdAgXDV31ADTpLSGYCnVb/8n2Z0k+PzsspfLl9Vvb/gWBucRnKPByJNC/EHS
TB4DZ37QSNA5SYfpsED5cE22ojitvX+euL/J1PKm58ItHiUeDAbUhmr5f9J8CDWhN58DldboyJ4E
eMZmF5Hmstzq0RfphuZjwXBuWBjoWpMF4g0LFay/8o9xIt3h/Q892hZKKYAaXi6upQBcAfRD1i5u
i3DWQUutroatlq+FmAntRWznf87mazjIB/zPL7q/nqy/UGBIKcG9/bmiAg+RGxTeR0aWtf+NeO7u
pRUit1JMOCD6hgMAjVWl1YFj3OBmjIv1cGxRH4VIWQVxC3hNAHqOshncwg6CImjadb6Dv5f/lnt5
wQA7RSZuO8ZBNtKmClIX8EzM7oTkbX+xdJNq0hkgIE5TxQyTCf2wkvMXb3fM2GaMSVW8YYoq6ok/
Ze1mCRXB5BSH/ODFmLj8KadO84ah3MVeynUha4QfyJ7cIxvyWCV1EIRvkFgkPREz6552riaHCZgw
eFNkcB3NCDnpTte2Ji1leTHcCtZrRuC0+N4PPVZpwPv89JodfAydGiTu3pOd7/C3spqrcLIB8uOY
uBF8dGv3YbLrjxylTB7dDuuAN+WmUXBPWHQatO2w+nqB95raloTo/JsXz2sTPQQxh0x99oxiiutd
h0Kss8n+XdJ/uIHQ4XFmFb9UY0SNaNGAsbmEtjUkp8QTYA01Cep4BGv41Dc0tuyC3oYIpH3qMdW2
uttp1EkDVCEk5SHbGLOoHOIHWtRJoARHdIO0BVFVR67929/WzfJ3lCvOqwb3sWKwpQtQIVY9AOdf
hVxI9DerleGeA6TRBLC+uifL7YnAmoWG22USatUgdxK4ZlyXE2S4nnEb/kAu+2B0OYqC54Vm0N1O
fiO2ETkMeWhosBO9Yz0AEfwGFLwK8bem//yiB1nxbh1cZnQfbMg7xP4dI3vTsSIvVZB1vg/i7p61
TIDIttZtgg4827naJTlHfk50QFTFEzAC4y14iwzpTCPlYd6kuL0qQeEhFkRukKHdYUUjm0gCjldN
+LK174jf0/DG6UB5NGS5FW9To8Zd96TpzML7zAUaRyny01ScIV29kQ+NC3I2fMvTBvmysTI6bAwa
ttoxeRNlM4363mqxHGuEvB0OCQ3HJefhZoyl3n3B8RI1s9C1zmnuGAerL9LOG4TciW2zMcdR5i0E
nKQ6z1WvDD7CjEjRfX0SMKF9uS+VgenOg6GfoLAruzvVipEXmuJ7+ElGVQ6vhpvEWIxUu0W81hWz
xVsiC00e/5KtjPKvjpdainUAV0h9OxXjSchUfUNz+y0rX7xPAInIgAXdjfuzkBjhPDYcINeH/7mn
pQaq91nc9IMH526JgdfNeKjYJdjUux/P6nobcJ2Awcpm4853+i2M3s4WtwWSg5JX1nnYVljDS9FL
ZHkZ28mPfG/I4gwB3w3Vo5V0ohkKf6l5mPKeiSHAGU7g1LerkrqmbUZSX1Cx8i1y2wEfHQphcopS
4SblT82UfVE3Y8sxmNAT0wjlQqy0yKaNptMUJTtWY38RzEskTafDtVE0klsfpwkAHA/1ZkOUy4Is
a9wXkdSKrsAd6UpxCpzo4/qS122T+c1wjEHLYWqQZqrpfK017PQrz+G1jqDWs1GHsrER1ulAo/aU
oCP4UfViUFJBEadg07vptfHy/J7snFhLBhg7VOYE9M6Jtutezr5vFpQjQDz/yx4XWOsf0CGLQrcV
tvIJWdkhZ4MMou5VPzEtua2LHHjRelIOrH5AXSCoFxHv4+eVGGQu1rqAdEzl9eCT2QGb1IOqmqzx
XPOlO+TX2WSkqUWSu4LtFkpVfUQke8x2/Za7/4ZiFC5ht9hFznJ5DpBMQPhUUQYT6TIXzcu3t14K
3j9w/9KwvZ36P97CkdE9+MY7w4Th7fdnI4tZ5D3DLJAKS+1fUr9Gd3TjHwDIY5iZXw7beQkv9l/V
mTFL3M3m2MM8q6XO5j6znhWHIgtSnidFPOdxgCH8AgjOkvs3RcXuqSI7rpy+yjVn16V6qIKfavv2
U4PZnfhc4JecNWuZZ0vtZ+i7figrrq7y2hfjmWPiJhEgV8z9u0VANaw5ALDFMIS41gGPCFA/5mc5
x5IGl85vhaRZJTh3fswMl48GX6cHErOT6CFJG/NU229XNjUxyiP+chTFy1Hod8jPhyIwz3meKtbd
NTN+OSuf7y0at9C3fb9zCywMr1+C7jzli8r8SnaaM0mLSlLYXyW7mKXCFDUH998GOx0icHP+HLFl
7o4hDtqy7V+30Olb8Ic6IVvXwxKIMNz69SxMPmIOBFKqGjLFphfZzelKEGdOkKGJQavSQ56b+/aQ
baKzCHLCOK1gO5MSOMSmsYsBbIXEydopb+DUvHTBM6PgxXcIclIoWxhZiHG+D2vGfTa725/+DnU1
AU+e5CKwZGzva7Z+6pRdRbVnI5q7DEu5PZIRTYO7eG3kFNmHXgDiPlPgsu9BldCY0Pw9a4AXsMQP
/mtUMXYph7Hzc/rbP1dkF2vcp23WyjJIOp80wcymYxQNz5sjTNHOlB8g7Qazvj6ab2DULSjBlF63
wDbvWOnFR7Ut4BjfcGYCw2CF2q0Z1utyXNxqv72xfXHGjHahqGo8FFYD+jU0JocxYV53NHCfCMQG
07iLTR+3NaLoQcS78ddWRuKiQOhlxac2iswSrzQeMu5k6teQR8V+3+cvw0LHACOZD2O/LJTafPzX
nPdoGbfV2rnr7JY4OWTMdkdE+9xGxD/YvsZa7tFRjt7sPEhA5SeIaZAMtErWx7x4YNX3RZHlRfsK
yMgQoIztAePaZXdf7RGmtr9Z6FeGgTadRH16/ekOqCsFutm9zMyjhgpnk3Z7zCVkLnFh6k5qNnm/
L/VDxAhQSAuN+/JrJBP0YnD0Whh6qcCZWhxTjjMQ/AYebWmplkfUmW47WEoSz0oLE7yrWBFQ8Vh8
TC3zSZykP0R2DLOjnJcsMWLAH5c/irYzmEOH2HleGcMgzrPNwA77ZpXXQ+C1uKGMVzTt+EbO9ZHz
XhDybwQ0SNnJ5fKD2HchNLtjAekTaG4GMcfkLdcu5lQu4FzFqgPmBMW9AU19DJX95++ccv+AbNwt
W41zRAun92/NSL8GnW5qlXn1gdPHM2WlYK6G7VG2aftx9bjbjSoUDoUyRZDYUTZHgBrGbPCCHQFY
nuRdO9aTZwh6AP40YwjwSI4rp+4cj7+uVLoUmtW5jhN0PNoolI34lw4qVzJjcEvC06tV19pHzvMH
WqY4s7XdBEG+2rif3vGUlL4o2tX8LCHglazTUCjZWUVrBR4qAu/bnDWK5w+98IsqKAc/CtoJVSc+
TiSelOVSwCR689pJvWdsWPzb+dG/j3FHCYxeoJWpz/btD90Q8XV1K+I71KbGiQexEJHT6TXp18wL
qmxFKaAhf8mHFQnyiuLRkplZBvhWXXXDp9Gr6VWiOiXjtPAb0mNUACP1VR4usYURloRamSP4Z4Ks
qLQNGoNn896Lj5OrFfdAc0nRkzNqcjkoQDdTF8fLZHlyhgrh6vj02HRoaLtNUs7D5Al5jPxSfcoX
/IzdE2sCysw+MbVN11rmN4mwt3qn1s8Sa2Ip6nyu0e8aVktsKo28OWmduiTz8EWKG35zwlRcaUVv
Ipky007lfYw8e1K70RSGb0x3wceSYHb4fkAPq969ovme7yyouSxSNfGWna4M2cFo5dWOnXali1iz
6zYx0G0Syj93ly/Yo5bt6zwNtYAYia7nOh03jgYAVTcEjNypgMmhiLJ0EZJAwPXTDaxJvrg+3V1g
R5u9mf1TkX4bmPjrTHJuM71ddehYkUsje/4qLYXYIgd6dC5ARSsHDOoaUpjPy75tuHhXQVRy/dUv
Qfr+7N7Fdi4Je+JI6nzATeGp6fFywF0GmIdmCsxedViMa11AqeBQ5sdRKo9spgS0XxCi+b2UY2LQ
tRPE5akqwS6rhy78T233UjkMqxUFCaN7AIbh2Ug0GQyDPd4iz/yu7s/C5y0LrHusYmkNdVOx/0eY
ks8I+2g8fph073zYASjVIF0Hl8AlQ05i3TGiyQRWJoSYXOgfDuEyxu3cf9I9DJIXWog7PJRgHgxd
fkJszjAAJW6JDENKqVS4yRB9GGWcigTfyLQ4nyHWjfWiG43Z1DXCQ+61K29euNUes7gLcZw9h4NC
iajfe9usBI8ibngJseMSilprQkQf3RvnaKq/qC7JeCGzUBTkoUhrf6ViMYGbjCxDjopdpDWk1OCk
AlQ++mKKuc3tPrydTNIN8fcIheY1NRyxbVpnoXlfiOSwH26ibnZqfPS54wW0A5IpNGWqNlHKkLGy
p07qFWRlSBw8twzQ/Uv3ial5+u732Cly0SlcV9Up5xchGw80jpWbIy4USkZutNa8M65KZDm/qHpa
3el1AY/NTzGn/0EH4B3iKu3cBWD51m4JWDSFrPh22J4nBfR4s/bVVAwhDVnPlvqxKTbBwDkpyXok
ZOaGsi9xblb1ZJfUNmQEs0BeTWmZ9nY+qJzVoQcl1dxweeCCYRXAZ136r/njisoKbnk1tqPNGNLZ
NyqRnxr/M/IVhlgg5GLA2hihotILlAPS1fh+3JbF7RBLteIPvYwkS0/nQ+3LbF0YhKFU0zVsZpWy
5J2fVcSzOcl0hlWqr71/KVwzkXULV52ItcbO4wjFOqKP9bxvxKkENFfMSbcU+LuVtQhckkI6AmRv
BDLM5vuRzinCgCd+VFSuw5SVeU66irGMeN9nLlKxS2iOc0vj/g3Ow+MOjDBgX0ighb87at+xoawR
cZYYOkgRZndUpgRHw+uWo6C2wpBzlCE3/mba7+vHe0umhmWcgAVlNeN33Fd7459DLP/dmRu6THif
Xy5lSspZOfiCo9XUhZLq0ikhzTuOfXhe71gsWVuOVmC0WcNX8N5pk7edJ5cUxnh7Ik4m65tzxb0Z
1ucXW4VehBWmDUkMvKAG40st5w1RVOYl4judC4rADvAMthNftMaOPpuxi5482t0oOmGmxt6GViJD
4QlTSnFF4cKxNBA8lwzwDoyaGDF3oKnHKpoh8sLZSrgoVgdym518MKhPY3JD7uGvNvNFkX0KVQjX
eBZiILLNzlp0auqCAW4biSc9ow/1OUco1toJoty6E9Rq6t1Avo6NugPPPY19NLNcVhO2VMgubuyh
Db2gFFcM7BeuZsiMw8JSrDoFfFeJxwAqQitbaDlgPnRnqjZ/m3QR1+jOYZGx/ArXXQ9J2Hg5RHtK
mmfDV0zVMlJ74OrhW9PkaC0rvz8riYumsVp1gOZTtF70kqTjdMQRwmkjI+aKElqW30Hz1pT6aEPB
j/z9vex14BriKgkP1cLXQMLSOQGrDHQlMJJaK8jf5mLIj4WxYwniRhzp+8ThYtfaFEpT1c0Ytku1
PFAX9M7do+qAPWKvfIoQXDrEaeTL8275/D4AVpN6jBWYeZ5prZYOdBe5SrbmI9pPk4GG7x4zAElp
snI1OOabQjGlCHC8zkelo9x7B5QNKB+hVudbvwJkAFDcwKVstup/Gg1ROZTFlDQ6aP/AnimtFe7J
oMhGdWMahGnkZzNeqoQi2eh79AT8jAbgC+Ir0taOVqElZC9eem1XQ/gtGGp6ICD73ecU4QGTu48x
6ZOr3TjSZKGi45V22szVdAIhvnp4Pc8NcMMy9aHCefZqO3BHsYunQsjRm6T+cn4ZAq/C7Sy7RoLj
yT6e8j4IYr5JoPKJtQE+Mf2HeIq6XD+59uiVYArn10PTzCowi+6FFR31gjGO29GW6Xj2JIj8X95d
1r+fDgophR3UEVGHbDztqElQlTPHmPcGAerkMHBDiL1XswGcKlcHLVr5gx5oSAlviipneMfcQbE4
BFZ1uaR1BeiX29XbuvAvYF3YlP0k7qGjmbbZsKUy+Mz3v0YlLGZn4rXz6mxJu1BcS5gwvQ+6dsOQ
KCMZIZzxq29dSdxldR5pNrdRUx0YfPVQsU2VSkQzIUaOHPOzWPo2RNsXjkZviedMyGkkfQCDxsFP
JhgGMH+Gy8SwbnhBQ/1UZh8/OXH524DUWjEGnPu2vnZvIAYCGywkkhrlz6kNOX+7Ntsj57ujNIQL
FVGB92d0Jv7LtLkHpXlzDHOQyBxup5GsdMDHQpGdMfIqCJsLsFBtFjoWYGjzgPWtT04RYeSe7NM0
aHLIJ76SfsKdEXbfHHd0bTK+Bs0J4SRMqikPAc3Udc2LOtUSElrGH1qf26/Wrxf9eUUaIGVHRptp
XnFzgbIuO4jwnDQTJ8mqAP7Z1rQ2jbrlZSfjaZgL9Fa2Rh7dW8PsMMvxkYM8DsbUl+RW5ktKV4iE
nb8ET/3sF/kqaUUI5oC0uPbPWvckQG+rixZSTRPY9aUuyxjwtcUEzKD0sYR6KdE8iO9ASAA4W7EA
DwFa5Led/gD61hKwc2Z9vr//5fyixGeAujATCTkUoL7PldM2dBCqoCePM7XV4kWLkCiKm2lu1/GA
JmtiAoCEXQgzIhjrnO9VRAkRNu77+39yC54RrgITP4DSLBhf8YnOKS6lpjSTcTBUMWESFcnyk1va
yZPJy3GDaVSqU1fmC4Ds+iW+0f7Gd93BwBA1HAHTLzcw0bci7H862u1vNN5SU96TslaM/Wvetgqs
V2vR+AKzPq+al01PK7DW9wKQ5TNFBCjV6BvC8QTRX4Njym+Bs65Dl0FExd40FNpDuWfru2i33H2V
FBNYiK7ezJUwHyAjmcz7eBS0SMHtZDbOlMUnPjDiIeVKMB8SEqzIIPQn2t+t2xOrfOeFYftbT8vv
TiayDZJgwHWly94wgglSXJq3V1jQb9IVRfFTUijJsqL7Ve6aCfsPQrTWTLiQ9v1scTapycPCGe0a
xKl9JVkVxtO/pIVKi14+OB0uUzqu1LT3BC0mOfzQu9avKIZ30U2I+Pk8QAEIVJnXDoI4Fs/77Hnf
R1iZEfah7IMl5LevutohBf0htlvhMu8aAjIT65m3Yy91hdbeaoW6AvHH44GXJOQ6X4G46dBjdQPe
py7X1ydp/1JP/HGDJFVCo76iEzPjmPTwQInVaGH0IxnzGJwiHuKUgvm8cH5GlGdG9JcDnYicvrhh
Nmaz5QVTFguIR2nV9YBkZkzmGkKtdR/OCAAspELom5C2OWgBJ3lZWc23yeK43PuQV3cgxTaJI4Pw
IYHG7tkr88ozxgm4Vf+CsDUU4Zze1yPPwe+gigLrj6FeMmITbfIShIW10Hk0uZv34sReblGK8dfc
DkdqZEt3yJFnigfyrvg/FHf5kRUJwgCwZUitoD+ya07bmFt0B3JzDdPorAmEvXMk2ouw4K+7YWO0
Zrcd+BTGw6NBrPj2qW9Sk6zMj6XHyQ/kj6h66/YZYn+UDzhtUFnWiEheB3B+SJa77QKz9CYtachY
mxg1a8J5rnDkdJlkeX5NZkQj/IMeMN5kaqsDBKHulF3vGwC9QnIVsNWSLvyJ/nTy6oyojRoKy3Zj
B7QbQB2qFn4kMfcKonEGgo/x2rK/ZRAzaWY441ePxVfI8HBUlLurgPP8brtcbF6SrAJNhHtaz2pj
fj4yqmAH/qRBMoZG6HzavJJQ+iqysZyIIQp7k3AUOs6ApndUv7bTUHkjOko4TdogToAR4TUoNhD9
jaKk8ldW47417uC3Y+bIcGBcNFXyNO49fBsiZaxcRvOqYEcv4pK6EnxdBecO0UO8wPWCMmRqol/W
KGGfDjcdQMmMG1n4XBaZ8YmFT5yYpmMAH5uWwO94iNgJy3S13in2wgGUtEGCaB4KrZg24EhMdq8l
MPaCqno1RoasvtxCnjCKlRnYmSIBc2+ppu8I/ReHHE8KY9JDMEyAuJDlGDhw3TnMeihAt8QvO1Gd
KzXJOyPH8vvPfuClwYnUVEgEy5RlxZUVp6oevRYlpjbwHa6rqrvWWxw69osoWy494NQFpJvuejfO
XN8y/gq0y6GRydR1aSuT+yc1YG1ZtU39g+PSXJl4tGyujmWoPNs6PR+i2T8FWC5ofWlH14U9Q7pj
z9Tavj7Zucmj30/TOdNXSFc2wUp64Mwi2DjCYlb09k/CC33lQ0CH36Dr1GSoF3J6yvMLurFVmO/Y
ht/UiQEhJNqrNm8PZ/dYKe0gHpD+O2TJfWuKiwaHcclqwq6jNwdCzQhHjCi2RpQBWklJ6fTAhs93
rixe6sDXJFgVdgyBSxdrFNSLbzojfwODNbP/eMQ6bbDKpAwiSmbriVbse2KnLbQK3ySCfUjNa2h/
PhFJS2xNDKWtVcs2yVWZzWcIH0U5lpBZEiDu/vS/lYKO3q5efZj6hBSu1G//FKgKewYbTj1ooMj7
u/7wJzqA/9kSwWCJEEp6WjX3hN6SEl1yxywSgvDHSh9jxeczwngjsv/AlMIeXaX858zJeg2jBa79
25jxl6FstXOMT/Rjf80geggmao8X3IPalW6sFOOYXDz7u9Ux6ve5lyFPP/HfkWD0Zsh++6R92uRF
fPsLqcLS87v3c60AxPUdsei+NUNIfygsbwTZ2TFcWen4CBR7LYyZY8Ut7iaiTTuj2BRMf2I+IEe6
NuuDtLHftHOvAzcI+pGIp7qOMaLpJbpvm0XJluePbuS1nIoDI+ILNOpEe5vtuWTS4stXimVjVt5y
n/bUlLPpGikam6zW9/6jPe/602HbbEP5BCW44WRfWonWpvbhtG23YGgxxi4B7K8lNT6PGk0s8PwO
MgZPINS2WVVtkE46TEDAyldhOQEtN1hKMk8YG9JNkwPTJhFpsEJ4skTc1SPhkFdJLPoNntfPTTc/
dycwc2n1aW8iZtHL2ZrTjvxCIQ5z/G6IxmqopC5Z94BFw/cttENyBfycgzQaQaNtDxj7MZz873St
v9if9FRKODGlsNBuBnKPx7o3RMHSRrxOvQxebU8wK3zB3zwPMKBlLbuBvkgtEGGbZcULR5BgQsXq
cgYvVXdlKRY+ZLDg7vGyd5MzE86t/DGq1q/6sOxT9HjeIy+gCScLZvaFPlwiq3t/llmKLgiqZK9o
5jI/+w6LXtEbhPrUsBDy/vliwt8E/a/ABRDjj4bKXjLb9rBe/StkF2f5g3ZeISE6Pgpxccb9nULw
V/HBL5ULyo01O95JWSUbPng1ntYJRzMma0ZKOtigZ7rNocl9jfctxQcYB/2/pTCysTpF9a0RJhFv
kpQ60bBoUOWSBV7MDIPVv8o0zRJFZ8xoELuZgzugzfOrPdUs6esnOoYrppa5piwirS5ZN5fgpZ4K
zsXtOEjqtGjInBfAUjYwEqE+2mcQ0rWHXfEkUopJYNvbH/BGSlo78rVehfdY0jC0CtBJpsNqw4aO
/fllykCHeHEhAvlxL2CTUKojGrJbi7Ue+0cJ6NgvJIdaOCOGfFURioF+pYTSodyVgh0QeuM5tDMz
NrRVLEBZRFCUWuoYs1PBpunyKldo+rHhdMR3BoegEVwOvQ9/45piWoX7dkIMII2Aa6nASThRH2iS
FkHN8EJyxPegKOi9Qafr3fVHREJ18zGk+k9Nf9EjgiI6ClK80lMf43o9FT/9exilKj1vEn6hwLKg
pt7MDRYE1SN3Je20Q+Z42M9nT8ao6YfN1Sy+Uf2CpGtedE7phUGT6VQKApBSoXj6EsGM2g2IiciO
rHTcLR2EsWWaXCIsSuxZ221EsA/Q9FHs84edvrFw3qjqpzS2ydNyFsQsv4poM4DdRpf7nKgGxSek
DzL6kUUBRUbUNWMzxjBs1v6wTOr26WssdEbo6CK7Xk7qwLFlkL3WHBPV+ijOspcZl7noygaSn2Gu
EYu4LEeJHA1I8QdihjmRmLoXIAmDhgGbvPTxzCpH8y6Ml2QS5O9A7UvC9P5bD5aUIiLv671kdtv5
tb60f9p2VanLTP5/Pb2VvmwI1we3NH79fS6LrZjPM1byak7bWVZQJ0Z9hVXVH+0I3ayWqe/2KEUn
y1XOEm0T71fg/3YIw02O8dcN8rf0RzmXglaaRzE7rw2f7E+pD3H9RViSZB4Rr2keeC5UFnaiv0M7
jkkOJlA4pUhLrQ4oPw8gRPHvntZdaJbOfu/dOCmsgJnZvUhzIKaULNtCsEwAxSPz4L3mYfNwGX9e
l4muTIu43W9/UkKWOVWkdrYE/VVqRbUbCrEnPtHycHL1o7Ba6ufUoomQFBSlKGjiNkSI535rvZcB
2UOxGViO8Xkj0Jd2lxqmCFL6g6sB6IcG3KxPVIarN3u9nz/X3K55vPkcKdBBGEjAvaofqI3WyP/T
UVXHr6G75i/CZ70nV6vJX98s404tNvmec1vjC9Temf5gIvqH1nOcBLa+BrnQDaqF+VKDxjA5LOfg
a6k2bcRAkwcP0k18DhwJoUqbLFAmhLrtU4Lq6FPMEkDrSl9Qkb+MK+EbWM2Gxtj6w/E/xRPj8ZYQ
io97FPFAZR2BJJnPN+UCoNREd8h6fiHxwntVkO56r5LdJJbwPzOmJoBdWcRmm7AQl0Jg8h2TG8qh
7+juNVOf1hS51TgN99qo+FaHdphttw86zr5rkcCp4MQ98kKn31Kiap/ZV+Q0U88FQ0f3tEpM16vY
xRky/bStqv+KRoyAqVwu5l4sfxshK5qwS0uLwpkkKPPrTrKuRa4yDeXzI+NmNlmQ9qqaHWI8ZmOa
pyxTQr8btmlqBNa6AdjxE4r2gVSX7LaL7oOGycwER2RgsiV9m84VS5FKv3jp1xBWijG98LXHLTWG
DVRm34dN/zqfcqhigEVNLL0aHe6Wl8jU7MJAbQmCAzJEqVLS4Xkt3XHHgPp//zfOU92WUH/f5tlL
2BP8N9VAMa686Qf9JwPlfyPfchPLialFuEKJOyA3I2yTiYFddGrgNUkyoin/w2a2fhhLydcDCW3w
+fmlvWpankx5hOoqC5a368ui7UN5WC57KEmJUDkwK/golKsV2tl6QjKDfBkppJar7lcFOMoIJHR9
0pBe9GW6N5fNv5ztzHiZRa37klYTeQtHO+xcNCeklMduQnlY6fiz4esoVTRa4jg1uonBqlTTEZhh
kMfKkj9kwWDzkGpIw0k7Hj6vW0+vXLokt22jG1fJlW3RfpIUb+NLxjBsYCnriMnmSodtP6LgZtXt
ZhSyLbH1NgJiQUYIhY955NAlMWa2f34h5XC08JW5FAgMWEEd3pg5rFbHVNSjbUh3W6+Jj+SBQsqQ
BBFf1fIvGTYZNYuXw00s1bikTiHe2oGHoSb1aFjc9tgjamRrBS2qW/E9htEja8J7YACYX2ptMIcw
jpx5s6Gd1kgCBEjq9/JiLN4bSl+DK2hUdfmtXWvJREDiin+6+9gSa7atVp1KkXeP2S6niba3pE3h
q1gJfaZTlVRkvVJwEP/3JpEyN4J521om2L919P0/JwrnKPE43p6m+9zAYswTkpJhOk78cVyyZNwZ
wMz70Nfk33rZoEE9qSYtw1GGsMWAuQuMmSGe8RFBdTsEVkQ6QN1X/e8i9yq/HaFVQLSvEH70A4Pl
22uaujq/ff316kdAV6MDbdq2tEu+DQm45e+B2VfbUxeMVIu+KDoBlBpJ6bEVNTHRKZBkUdyeqoTE
EZCEgTLSgvDOauhvmhLO3RDhM88h19/wiX2ber89Jpz2dH5InJeoriPwh5ZQpPa66U7JJD1PRahV
VGlRiazHhbJ3R5vREPe4Mz97t39fEuwMihmz3et08PNyHsnHUiGNN5gfmMJFT+RYZATJCwYH72CK
HQEZWm4CCiPi/uUGd2AgsOfSwcdJ/zsUMe5n3bKWbxM2xos4gqWgU2MjjMh6w1h6zeIrcFpxk1HX
YtYRszW9aHFbk19krBYDwfXWdWpiTI2n9Rw2ON1qWnhukuTA2ukSBsCK57GMazleIdlrzfOqQqSa
OSUh0UFeeGdPdgrhWr8juFA7fSy6sGcxAm2Q9Oo98dzETVAmAQfOqiSpeUjU345xjZzPnMAHtoti
x4o3RwJAVB3Ppi01qQ7HxdCWUnBVefdcW9S5AcZHhxiv1lIm97FGPHQS0x+mHgzfyu6itBud9aEL
5FzHiezt5Kxn8vkpySVMXHUoxYheP2N2hT5GhDp3ZRnQE3ZUVyT3Q07HdoI0U/56GcrD1+U/1OjJ
84FlEwh6Sk1E2KZ3Pz5RCbHNqcmK63QtxWNW2AFs4xytMYycYrlOgLr2sN0LSIHFYpq8+D2HWNfL
Aa35UHY/OttojhKi7V4sEHuVxRmFzTCK4bfmNMJnyWZ06hmwAG1aam0J10DDzCRcEDOvAQ+7VpXX
HpDquzJrc0NcE8gzLpb2n3KfeJJo3W/SBR6TIJIn6Fzh9t7UFqbXE+UzYLZn5c0xlbjE7DAGqPDY
UmjLUicxzaimuIpu9MkC8lYSnZf+d5lh8K4jiEtfLv+j4b7OGTFmUvSQep8ifUO4/+6/d0M8aK1e
uD0jvbbwCLjji4+tAhwV8aEoJiHHfJoftj+NVdPvHTJ7pqafwL3ASadahvR/fYu21LIcnwkP3HLM
rxJ9m3gE9sNUQ28W7PYSF8WT2gYs2JSXmXvhtQvV/NFWj+x5j06wEYgOl89zdRqFjfU65Xu1YGXk
dv/KQKj+SC/KWJRsI4NmflNo3uYtWXeslfOEnuZqPOHUGro5pcdJ7wTbOrz5SpgcbZbdDloZN/+W
Ss16CcwKUC9xU+HCWPF+MzK6l7LYopRpZII03xi8HzJBMART1clUUtTWsqxvBG1yPekVn/UGo6X2
Aq1h4SWoSbLEzStFUGqxmb9npywrhaRq44rtPRK2Q5/rqXPP4vfwSMN5wkX1H0Sz2vtpLLIliu9a
J5OzpGObN8iNhs7DVR+mEzmwAEBxDp+R3f/qFsuzMIgAxYIPPu6cyckqF16A8AE9OEuOgCDawK35
axBll7G3Szo4ZUsWxAPCgF8d3sF6u08IeWEU58jZdD4lwgQnBR6CYE+qIQDsSrYupBBeBlacX2BB
arg3/8aMpVB5WS2YRrRf/3+xmtAbnKqUeXKSS0irrFkDfWqYO5bywiKWmC5al+jsp3d0XTb97h2S
EhA68LU0qPGoIPfoze5To9WzWAbtmpjz5jv3cTP5YPBNy/Px8MluaN+O5kOtgNZk/7Wi1SlHt0/T
Inwc9SAi2LPhNfGnCAMZ3Pv1SC7AwDAtNDabpSir6YH9ir1U7mJw0zyRxUlFRqQ9jfM0a5C3MQNF
VSzTUDT27pbv6ymZFye8ZteXFJgNZcj60yLwYTZgnngU+Dp1G1i2Ta+tirXIGWjjMfqIuJzP7t2e
++cgTstBs+MliI41Z2SxP/j/CToZNk/znWcZ/poeGTF1WEiXowuWSuuj10eWZRDqNOOZNfZH8sLT
aRAfvxGxTo7y+fsrpfQnDgBIB2aCTZNcu5H7RR8MEJLnQ37elUYAZr1hAlr2wZ/rX8dk+igS62CG
aQelJ9Wym+bjJ5iFdZn34piJgVv4041CNfz6NerywcgMEWMo8owvMne5//XsUpImdb8ANGbGlIPi
jueHAJ3rS+zoEcWFUgPpKy9RC4Cr8luwwwqsNT1yoC2g8nbj1i667j6y3Rx98HmqlJs27NxzVCaV
d/xhcAoKrN6dls7mnOrMQgv5oSYHGnq4QndsBFkNo7TsatKvx/96uNr0WXPnj/c3ASj/rZVnpkYQ
js5uA05luKhq6G8okqUse9gNttb0HipgKHsAMKDHjBXaY1V1hAoe4w4uVDHdmIT11ZO9pe6LH0pP
eFSNv9Ea7tG/CxRtaSaTnmk7XNQAYlxBUcdka9U4LRP+we0QdiyBlcFJ6lIHRutZ4q92SAQS+3Dw
+N8bIJVwXQuwR7KGVb4JjaWlVAKhx17HoKrOjDXTke/UaHg8FyvRXMJAgTmk35/2q8N65g8gyWIx
UD3/py16HqyH73gJJckR3e3DNNtDdPUChPZ8zYxzDLTIo3dB/mFyCnKLhsgNiUeLdMlDV0S1s9Kf
sN+8EFV7MFbIBwu50EqRc+WBMgagZbzFQpnUzB3rdZYgm4aPsOPe8Wq4F7bWXTundaPrsDiWNnnu
78VQ1TE4Trv38iW2SZt0kqu7LRDlm0FdqioJqq8ebS7u3Yz8kzH78rFK+er/NZUxmMWfcqlhQ5GX
qB4k5J3FhitSQB50vIW9Jeqx0ks6SmD0LiQ/b+jPkAQLUIfOAr9GeRW/yFTXkgQ4n2b5dt/OYPEH
ujz9wCjJe22DnnmtZMyyx5FPKUng7Yr/9ahZxH/Ho+yEsi6dGG5b3ID0E967LlW6zZUXU+fnKdGY
8PNWrLyFMgw4zlvY0kJhlMU/Ja1VtkINhDFqtbgipMH/4VyCElkZfH58+j/cBiSmXXzDNiOmOmWR
Utsu+x+UZqsrP2+JbA1Cdbvcoy3UgDzEJP0z/iTqmcV9SQqyKo5/GAYhoV+xoSihTXmJa1xNLaTN
bIz68xjDqQxOLzlj9+gzN3uTSwpS4n2eiHP0PUk0hVX7DEO1NLdqP+3fB7A5cn0ot6FyNi28klfz
oe8rhtkZpiS+DypL+Mn5j1kI9EXy8spPzrMJ73YLZ6v7J/kSMZ162C5ckxxZtadefztLUTVZVFjz
3+rMG7E1yG7LNYjwKM6782cEFycXvgOEH9raOgsIDGGq0PiND6fejgu16xggHuvyKedFnyD7I7E6
za/wFCIhNRPNxq5nsYmwH7KHMUR28PMl5fjgE4EkecuM4sT2KHIe/4oerMzR9yXRTeDljalvsqlE
JrNNL14zcuPvLMUhrvNRef7drSre0LQVFlO6MmTxsZCW78R0k6zHfgph6v1jlgc5Y3eHc4wkfVOh
vW4tbMudavTMvMXWmjbX1fXSUmvauiP1f/IJVe+Q8aO23qVREfwgu/K3GYwaryu+iv9jzQaiGNA8
xiGjwupGKXPXpYxGBR2iuB1M1Q3KVsfblpYzm7FkbNtQngvbbHDpCdfmm5+w+v3NPVS/erI+Iiqx
LeSZ9NNtZ+jO/P2MS29w1tKQj1423oJlBwMDUM7+Fxa4HnzFxXcaV2v0t885/8m+rwwitYGMHCWL
EikXAaZGxxOlelxaFzIK0IJw2fsNa8kv9o5oYbORsbuydDe/BHRl61v8rruNSUV/MWNMiTNZbiC/
PnK5sEJ3MIj4Qc+4qNU+DFriC93o7U/F87PFDzzYlkPw0/ee8L6/ffUua6ZjVMMgjT4av8ySigpC
Zg7YjVMjuj/yclBHYeevp9nX+FA8OGMEvJtGoSC3XXWsiZllgr/JHUkoTCIbYIeuudIe1w23BaZ4
cAYoZJ3Zqw5HZDpo43nw/1OoBvk4ou2gIYZ15fSQWakOfNVHy55gNZxVCxJcnjl1tmVmevk4Sxju
oyaZvJ8Ed26KKd1qMhVpj+nQDNunEhIPFSQdcnwg86b1UDTBxxWlzju2NMo2KaLlLUcqAOoEQa9b
hH2fdbzytT99mBvpdpLBsCH6umc1FJb63B0UD8DErbZCcKhbUp3MJra79IqZLA4VqxavGl0hCV6l
lUxPo4NfurScBJ3IEZVxBd3mmEzesQOAWzbDUHvHD32cRmvB9SU/vqFZsYOfs/q++aHLa9HLYl/m
rexADw38PWuHbke3JCDBPZBOCu1QZHx5GMpgvGTwetHglJRhs1rZXbIorM59jOIaaVrH2yPSnZuQ
7ZJ24DeGv5RoDucNYmgyJqbO3TmSC8jb6tupjcZ0433KiagbwRUnBaIuEf07L2FtJ86wssKEAMAq
13In1DyL14KmknaILEaVGpytqCFuPEL6CAa1mZtIZmXhnQAfMqhBmW4vj27fvxeonPNZR11/AU8K
Piy3MhD7x6+FxZ9srf8+i6Vi7dzJ9Uz5voEi176QsfP0WE6JLPDCPqTlMuZ7f+cbsUvvXpmgDT4w
mbSbV67yKhP4HrkKSpxg3ksAGTLG1AabiuMf1oNMeQEeVp2WUwmx3luTbmXdmbLt2utazY/u3M3m
NpkeYy7U0vNhm0bRpmQDnV2EqQeo19DUwJAjjb6y1WToMdQHIYcKJ60CpJmJK28lmOMA7koJc4v0
mj7TOeHfFhwzXk3TrdHWl+P4Ulrpro2wiNABnhQIMzW+oQQ0xxDPxsIhpzWmiO0WxOAbYpM62tYe
Ns47Q1mmW5hcRnUzw0iYGeRCtM+yF5+gMDe/Zliar9rBrDsqK6pNq9M4EYRougN8U6ASvB4i+LNL
yAcC+Ko+rn7XXWfijwUEng+GTGhYRWWgz34YezAwtJHsH/cRZ6umTTcTaHrY2SNFxbCvKC3Fd37g
OWFVUG6zu493xFpvF7u4wRFjaFz06Z63Gfr50W59Mi1Ua7J6YNWzTR6K0/Ah+obyrtkUGR3DnoIM
sQa+m9ZFOPYuCecQnpkwMz7pEAHlkbGqPRWPZW54RDLN/9J0/ti6CqqtN3j/CIuu5chHmRoZmiCX
dxMY2PL859QkEnehYet3CQ4pR6CdBnN5DweFV3jENYhfWap+9/3UWsPbNhF+JGmwsTjgidd2ddfU
JuDMjLw0uFwHzdirwrcVeNKGfjXtzy13h6MzsJyxM9LpdrHwI2IZXGQOOuKnq3eaQGVUP7qDk53o
6GAFJoupBPKBV0z73bLyj22cH549CPtPw2O7czxDp0yQejeGgI+Waab1Ts+EM5Wxqe+rvnENOTrM
PMO2QzZiYW3HbrPz/P+azq1QDuqJ3gEpGKz7xBgZJvYD9JzDR58bigVkgOcEf4nmVEzqwbajEuab
2S3rf2ED0C0RoJc/W+8PhWmk/j17omXGp+WIOuhzgW13aSLTjizVPUjrOsPEI8X5xocltqOuevRP
X+1wmJfn3OiJ22Lrukw9QNPiHAB2xFbzik4qflK8faz3B3oJKJgGfVUjp9EArsr5btPWReIpfOvL
8I3Onn7M5wYUv5tP/EOZdVyH901w/pcAZ5H9rjQnaTTJv4bqk+GUWjiDZJrOgI+GSxK5W6UBe+qF
0OjYANI3xPZHSCAjPsSN1t4uOrnzL4fVGujwMOuwBMWaXKegxnFW+bC8JsY3Gne6TEbWng7O/SuI
cD3aT06mDs+NtwHiFfy19V9KfNMXLgXs0Y5vAPsqAdWq9/PlBoWYGBiKeBny9ZyuddtHKbB7L75I
VBKT6VHIEj0DwAGiK2BYC1b+Dv6O02+f18kd4gpA7hdFipQMGoNO0UQWM+HNg71vvdCzUa2tL3rm
Y6pm0D71kk0rDnLuj3XLvWdpJwj1KRxyeduYsWN9e9YW0Cxkteg2a8FJExTiqDwi1rKTvLcoZ+F+
33gWmbZb/4gV53FX8Fy1zJIC4Fb4BkQ43Zc7q5ScafWqzkDdvTVDPGlaws+YbYn5mdw93UG7A0Zs
T3egFgaAGezwRPSJ5zFdyiDhjcLCMEIowIVqMoofCPydPcic++RJh8YzQP1rmXdaWtZIVRt9xl3V
ZtyCiC3G6I0HnZ0/tdkp3qw1jf6BTEMCKpzU4r0qH1YkNnGKqy02Lqk2ZLdg+f9vlc9eCqEi+kEk
m2tEvJrLfwz0rm/JsCC/pRNPIM13c3y8EMSDIdeSbRwr+zBidlmzqth6E5eKyFxgTAlnOl9G/WGK
A1AH5NN18BpY0v9UZ27YIPAJelBGCXN1pe93Bs77G8nw42fxjoViBOqsTbVvJ11uftcNAtLLY8vU
MCvaKetHSw9yu4WGmJQ8SaOH7k1v56+/En75oU5Xn78NTot784o8Ti+sreL33BtXukJf+K6BkVax
vk6r7jDvGEXT8ve+b0YKTJP6wCC8mSdJKFkdLy5ETt3AhOCpdNIt/NNMQYGCAA+vER5xwHsVciNf
6D1F2L5vzB/QDZFR8kJ15/jS8cpwlusvnOi95WpCpwAIGCZaah3hPlbcV5sngcz/7l0lUL0UdIkw
r2LLThLAGL8ZayaOVkuf0l5IRxsx0RPi4N6ZGwZWxBNtKENCR0C7pNtXhjuwYPvvM9xrKqwnCmE3
PvAaY0xP4eZAgX2giukYe1MiKkeTMS7bG17UaFYNO143vDwJx/VzzoYqvmLTMLGvDUPabdZ9FVoU
Y9ZMQMpqn1dx3vzJM7Tg7l3ldOHh47lGH2JePIA+1sjES//iHqz+y8lHnnyurojTMWDypQCRZ1UE
16n9sxVmPXqiwDcfzE2LQ0LgcLbaWv5skqtFg4LZmdtMltN/i1PhIFCC1FlOtLgL0NU47QQJ/8XQ
PMKDW83W8m2FDwEHL3adMLMQmn0mFOIgmfILdjzxHDm8UmFBpZoQISw60pHbSHFsJgP5hhXtPlbc
qQlcw7txhRJCrVuE4RZkWZQLnoCvETv98nbdhL9RBv5/PTXvlDJ1dAJi7WmyeaY0FYAPc5uUM04y
7k9aCY56r+fnhmQhj6iSVs+oE8ELMBpGY2wx8Fih456g/9G1C/RKx4RmSurrQkMjJzYceZ1FhO/J
qPvwkRrJuHuo8hnu+APzXKzFCkPi3Weij+L/LoG/VLNXUBuXe9IrqldbCNMgwpE+xnPx8Iu9NitH
DRjoun5sbRaDgdfwp5y0f3Br71fBw2LFM8F5/vAwRK81G6EupJQ1xP+ux9PE2ZqQ0RfqZOia+32L
yZZDh+FDrgRvTr4uZPib0K9Xb/nkJDksZLuD9oWEGT7mLEtuYnXfbYthSXp9rJj8W2k/sBhnJWzz
GXER0f/DX3bLpsM6246A9dA9EpnfLQyQjzjxkXXH14jMz2YtmAvw3D6j3s7+QZLCIV2FVg4fU800
LWBLEiTX8j431rG9MUbUJbB7BKxcFMnPk/1nR+jyeqLA/KVRcaE8OXx+BnSZjw1BdwUns/zGXBXF
oW4wDwbiPDERagvGiNU/6ccZ/ADeRcShg6dtLdiN5rTB1Xy3ezlsiC69OZuUCadQk5SFlJyCfCdS
NpCUkhbXo4j5BRxFHsYXdSMcyHPZE1WCuiP56qfyN3hogRsG+R1x3UkyROSIQCtAFblGalkEUpqe
ypNiDzEjX9EwSA4CB6TgtnfVi3SGxc9QSVVo9HNhkO5W9lym7XNIytcdX/U2pFk70zZ4Q7g57MTM
MQikySxXuvoNoeJKBx8AHOV2YqdMbqFUd1V7dKWILwKM+HTOOrVTE2zRfLBsbzKPyNG9FYimff/h
Rr4hkTC1T8RiUUrRV8wN7vJhUoMl8xh0Rd/PTEf/P/6crR0mjSbwLR7qRRHZIseQoczCoOOoL2UT
6tYhPuB58LvIP2hZYi4I+syD/yN5tq36qbkbsIZ5akkIhgUaXOPVVMyyW9bc8Knwl3LMQ6cIyuUs
DWbMOowqxyu+q6Vm+BW1FNS52wrrrk1o0xGQYpAPALn4oT8iK+dtHGZJ3HhYkPo7FhcOwqJIq2xL
6QzqdD5Yw4qozShc+0WkCuY3CKhnmIFOc00JBY6g5QYBkpdMeGKumtm1caroTDyG5lF/oBENB4oU
mXYMgHLAqjPfadCaX6F6DepuabuQPUaUdnFRNK8j3+ZxRX+mO/F2wgHKpQDLlwD9paVx8rtb+TeC
I/9ZXEYgW7iAnOR9IVNb87sFUPxGryxAul6Rdto2wFnDyGF4MTMRw29szooZ/55FBn8xCoUcFCzv
ObDKD503zlEIg+2BwUVuT3qB47fIzQK+ShBFcKGLk1htEvMLTF7jHk0c6/vfQdGvq9NOBa9hX99X
NHnt86omvakABF12HA6nfTHDK/StZZfv0QkLgOK02ujM+h2aDC9QJKoWgHUiru/HxM6Augr/YbyJ
5Qz/qtn39CQzsnvP7dNMapVynK1KDDX8g22RIOTd2TMAuTy5KgfzuO1MtNc0AvaM7P8kiLTjlD8L
aIWlcmBUQOcFi8a/E2hAys0l2pBGleOVYB2ohCsShY45MxrC3P8AVUNVevu3Xuq/fvdQpgSE8kDP
y1oATMhCwdOPJgxhg4pCwBo9LgzMcAN0dV1lRUQG7l/rt/C0y/FZJqZ6dlPZploBBKzF6eJg7MXE
CFn41qpyFxdqVnJpBWe4of3ePKefUTlov627z9kslBeNGEa5xudmaQg1iOP7ZH13Bl5gBtBGGeII
UJKac3KKKOTPHvk7xgMztHm2cJLYbVFfFxrjQDknPbJP1u9iso5s00Edg2YN6k1nftoFyXmC3a8D
3LqZG1xjVHSV2SWBZcNTdhwssPiefriBhYkwS91qDT3oMs2gI4957HE5HI/gMVGiT4i/jrdhdTyE
CwCBnaINzqrt4X6dc2bhOWknyDMAQ6n45otAlelIRb1lQrbZ7sqzIb8AabWaBkjEi1xoFhoOLyHu
BS7DPLWPFBe4+zBsP2rcAq5eg4oZp6OH1F00wJRcaegBjiFbJYECOQ9a6G8K7h5w+vN+U/lpi03p
LDxC/tULhZU5rOPFoEpU+ZDN1pfgV2CRMokZDTkz6e0YoLp4zOaeWOmHjCXZXuc7xdQ9qxkqFTmA
UKm4WObFtJMcilBGUWH+EZykkQmaFqv8JY6RrsSMaoeXz5OW5yl3MOu7x5IyW0Oz2DK93mhAqJS2
bt1HnU0r4f6D1FHfceHyCGfSVVwMqM2579SQEYU/xVpJwdbq2OKRcYoLzXwt6TDl2fcX2x/sOHhP
0ULjahNa1DxxWd+LTfAbO5TfL/wgyk6uffms5ad1Vj6CWX5QfXpfZO7BD1I7bl+lS25ii0htfyV2
UHcCaf/yuFqbagyvH+C1K+tuB57Wy24wWLs95PEDjuK/2q14tymgNZR2ohk3UhGawaUGGqqO7dQ6
3utGSZRJ/GxWh/qfU/TBv6ttooq1/uwL+6JmxzdaTh1lB/M86DQSSXRAXsF/TZ/EXcKBhX5AYzKl
1N9zqD2xuPuzVd4V0/ZiIMUb/jw+SD0eb/N9knV2grRK0MLzV2vk02yhPb+rvdZN/jCHscFPpZpx
VntxeVdA9fW3iO09cTy/5Rewc4e3VWd9fRgwl5BLCsLFH8JdDKHJ+mkFt4jOipjZviTGBfKw1L8y
VABKnr+IOxIEUaCnW/6NuFksyOHbVOvMN1kEWqkQ0hTgBUa6SSNcUs+ouuM7IRuXJDgQZ/8P+BDg
eCpl49OpxEx63BPWWVW0Lf9KknA37+qJl5GtpsYdL85tZD9Yld9SEFbxmY2Mo7hNxgWkVHOSYWlE
chAp6wVBtwH98f3OyvVYU3mtiwJHjNgtpPXgPcLiBuarEcMclhUQLlUInzF3KnnsdyEChZYHen7Z
SY8mIUfg30Khkn/AoWw5iNh+pbBCnFLfjOAKaK+tFBnAkoZcJvWnwgjJR1StRoNVqxlbU7J8SF3c
doVrApgVMTivGKtLA4EVFQJ/QuZXA9QN9+OPzA6OzbY21VfcyHujbFnwKSEHtSwyvxCDajSYU9j5
tSnMBzvf3+EwdEx73HNNeFpSg7Nu5nABLd2a0sRU2berjqOV9y2Go8urrPr/WRgBWl2ATLVg00ec
kkTvE4tfMqeSYPVquwGNOKdn7inOZThB2H3DiUdrQGWBMcnORFV4VdrfNa78HCpsmOPBBWf+69pk
5RSXdClNeu+XlwaIQ+n1PP/KQWwF5/qHSFo9Lv7VBfC6VMXijYRnPGM+/lIBReNAvo4h5YeoyFdb
zyU385MTLOmDhqzVY4YgtXgyba4GzxDoDUsXPahDsfeC/6PwTlyWEcfBmnUGxaNVChzzTJF5yDve
7AJsk2tzL9vb3ylrezxtt/dA54S8cOOO8XpBtZiCqK/+YAo7CRDtcw+VwqCRC6w0DUz4BmhYgXJj
Vxv+CqUSdE9/JuqZVJ/Sv4kwNlZlR2Wnc2zBsa2qq2aje16xBdrO+ejXua6aUfF+fD+xConvaTNP
U+Sz0t9mzgiaJhmo/d3jHoJAkdfau4dc68ym3MCuxNBaawsREyRJ6l3458gPRk5eewwWmsb3AL7z
RmwpYSDZlp34/MBchCiWkQ3Ug/pKnayL+UzN2ZbxfnhcsDoQhv0SlzzZuWTvtlfLKzKh1SFdqluk
41CnJhlFJMEa7NJTLRZ4skaGEEzouB5PPfUGfxaBezivGWlyzRvVk1IWYK+IH8IccqBSVYrrJCmu
Tb6aXU0FekuHndJUK6mxXYdA+BQJPefVRENmMts24mrQmeDD1Rm/UvAwtfHE2G4Bs80ygyNbzEuN
NikJBROY6gDj/3LNuyO6E2fkG9rG3+NfVdIw+f3H/Du90lY6W/eS8GmHTCyk7eSzeNcqUr0xgeYd
bSmdL2FsX7qJAB59pV8AqXiEoTUkVx6UNFgEOZ5pZ+sXu49F/I7tYQnPddKhv6RNdc++Z6IjOtx/
JelD/jystNz7rIc4+Mxd5oYF34Hs4HuC+GeiSJJ1F1IrmozqvjsufQIu6TAl3yCM9mkJSLTDsZsK
5T9+7lYMDYfN/4sLknHmnqXRMNKVw/RGNAEWbG+xzvBeuO+Wuot0PF42OUe0e3i7ZXBY4jkLfWyK
fgOABKWlrt0Inkdlzt1Z3Fz8UImuWADoL7zEZ4OmSeQNr3nYx4iSGTwBMHrSP7o8IYMNuBkZ6hRv
TyPOOE7aQFFqhKcXgwqUUHPmjplYOwaAAwBvrpmfCVB7LsMQXrnos1D8dkpbVYf44CgPA71WhQkE
x2fr1JhYPoEN8tftRMFLpglreCpljwkR3CueZIi5y1wAixxMEkGu3RYR+uSwRyHmk63R9QCizYJT
fAKzJMhw+GwFQaA5DN5ufbeHnykJKqpneum2TVtetDGWDWKsLBM/h5KH6QCV++0D1y7mERm6CFBS
MJ7EW9nb0d6lZSdJKqa20fMBAI9cW+Zisr6sB+mA8KZqasaNZebiZEEYFwDV+Ass86wGQifbTaLi
lW7b3fz9SOzn625gBH7quEIXYVAc0BoV+CXdhAv9IfAUBt3bCz1VSfGQ+GgHqwE4rXT3b/F/UXzA
ypen2UgZb5DV+YxGI5G4zPdUuyfA9/n9eIvODlRpyAoaoQ5d04T6u3Lzq7FkmRtWYjoWvq/fK5qr
nYqPJKJ0B+Gjj8FBSM8vwRXW/WIUPfOoI+d8LW/uvGuz39ctgoi2+eRGQrwGqtCwpzFMK9jC/WK7
xUaD28NZPFObtaF3HmrMEx5uZBVrEuYiu6EXc9ts3aroEcz+I9X029/h4eIBZeUvo9LzybnFsMQ7
Pf/ptnoMQV1ExCjvXrI0wHtI3V0cxhIBlNBhJFyeEVKjMmpCqNs/9YlsjvouBCwYdA1xScumSC3f
DjhCEdxYPQfNCkIS2DT0zIVFndDlGTkRFO73zPyDGsGonr2DxSwW302msq95qcbUitArRQd782sh
mAZD9soCG+6xhpOmLxS9shaBM+9Wy44iJj1UHOkikQHnAJpFOKoE0dw7+DOIfohLXBkWXX12Te2h
htK0aj7j0/NW9tF2bELmGGTrDfHpbIxnWd4OeCHqygZPbxfx77AeKvDgPyCE5/HaJhnnMHEP44yW
V6ZPh4FWtYEyUmiMGrM2sQGZaFPwp5QZ+Tf4TRvIoTcPrER8kRpF8Nlyt7JXnuX4il3CnDSHh8Oh
o451V30JaKfVt/5yDl9b3FNppL7/03VkqUzav+EsDY5iiQWAaDIMvI0VVQH4Pfz7KifFUvlpugEJ
ucdNUpNHuXd+FRhfS35Q32Yn7iyDV3XZgeug6lpwxhUB2QsKNRhx/cRB1zh7Cev8ab3s6Su7xFP3
EH6TCtjxJd8Emx/o/uJyIduJhZJb5vR+XAAqR1fEDrxc1XESmKYouDBtx7zqHTkwmNc4xXITz27N
85ibW20CnWZ7C3MDjqNjhAx4h5SJwAn+iO0vqXKK4Ed8+VHWleA6b7z9kNxiTrdzEs428YkjqpA+
bPnqCTno+10ItltQ0ygtKRXMsxGyclpVR9875z5XMBXKvrgsMHP3q2AgqIFQmodt1/drKqbUGnPD
Wj0Y2Kxv+XcAPdJd/FLRWPomCg43yu6O/EqQu7mXfUlnlAqw5QtPtyzw+TChA4NyFSip7W0ClVHm
FgJpD22IP+YEmtCqjvpJFajOxPEcyMYd8i93Wv72AXXWQNYIfCsT2G1F8Qd0eXST4t92Gxd/UhXl
TJWu2jjpACJHw+HrtSOz/8YLYNC9AYZNlO1Oajgz8sb3hcwayJEQJBI/iP/8EkbV8x37cbJ1BLYI
vX7V3Xpntxc1cCPibMU0f2lipR2RfnGeJ/1i7zxTO+Z7e/EzPxLvw0b6GP0jWDAJtuMWO7hgNqk6
tDYwctS9/GnOCS8E+8+c3n/nwwtMfKJJBg+MRErT0l3Jl+eXxuSO+mKSkoqfa5VdbK+syul4GfUn
L992UKMbwruX02J0uGxeaSEW4igs1/i1VI2R7JY8l2P17sVWAKqi9uoDV+j0GUupMmAz6T7wSfeg
XnADJitFSrEKb/sCvkvkZ6OFgEr9pD43K3YpJYVllxKHQV3Cux2MOmackD39+rkPWqOd4s+bUdnj
tlcK61VjP7khKk2h09MqRCZ65MACZHbX4gVVbZDBwKWBhyElUANdQqAtzJfRAZ9ywbpP448Q0slK
Hv5ml3M5bUBgp3YZV8FJAEbvTBLJQjq6EcAUg7SzUOSsxwjylFUI7UhLdgfqzt5dKAIk2YcV144V
12W+EY2AMsyVf2NL9Kp+8zCGNON+8SEE1/zyU9jsdMMGzZAb9g+VAFwm/WIUWRa+fL675UM/ed2g
hZyLrtGWKLjmWyS3P1zykiBjK4Agl4XNqD/m8Z0aYF9b772xA949C+yawFmI1VPk1tikQaetD9Mi
0iNvEOUWg6P1KvQf5aBwj9mn1sNDzYs0Gg3C1xfBqdNkq5lXGGvDeV9de5LFjbHT5AjqB7iAtC0P
i/jMVzL63s3PHE3uIBxJV0t3dLDKmLqTU+/yTMkA/0OshdPlAhdhAeu8plbi3fRV6KErwJ+BKYyR
W5VtY+G/64a3/VkGtds6337ZBStT2MZ/PI9gu8iSpTgGiftkaotSuXVkvYRN3Lf6Kvbh9gIWOXBT
KmCLCkB/csagFuj/tUBw5aIz/txchR95XUDw1evYBOXl48Eaqfv7LhoqXxbOYBKx9Mt6it3yXFWh
vxVPuTmT7ImsAwDJMiJFlmm6lczGE1MRW2nXjBvnc5zOeT9dmQN7vh3uEcJtc+vso5zmcw5iJvID
70ilHezPoR1BcvAYK/DFO//75U+LxEKdjsUI63BAzz+mAe81wmJZP1x10ID1dUbdj20mxYK99Dmb
ks3knPjk5NRsKEPFxsDnWTXyOjbLGcxZ5QG9LZ6npIJbGIwIJNr6/geceF+AiQehI/t2YXBJGb1v
PySx4oop7wAoE6bG+UwBkX3VlscNOWD6XXbypsnUr4Idi8biDvrrNd66DCfucF8RBDKbjecNQjLL
OpSRIP9rQtTNYo+IAvkzpbZCpVk8HIiTqQsjcUTfYifTlTWuq/skIpVLiSnbtqPtHqvUnU7PRoNl
DU9KDXeF+Bh9d/qLZrycGTM8XAl/6TQruzcNAJczbqHoxv2v7vi5fylqMJVJcjU5EqE0yZBVMBy0
tpmpciuE0FbnuyUDSuPAhZMx8ViGzr9aUGZk4jqDgnCaBHDSjvCyK5BFjbyMzOeYe1VvPsYFn13s
rK8Q9xDhXwxw9OGBMAGdXK53pNIk84L/+mTmWqDZskpZCfvmvbBfB0wl64kJVHjugU1P/RFAzwYS
ci6hXh5IsCUHgzIccuYj2Odwe5DhkOBnsK6vtSqgwrvTfs1wap9bbQecc59IYJvUSn8PzZnhKp3k
ztMVETMQHRt/UzjSq+z3PrPBxhjR0B6bGxnYxloeZnijeBI2l5dlQ5Kd6jomuqXD4aSPVItkfZ4e
lnTryo+BP54TzU7Cbe09cfKWZs0guwnnyrtc4uqi4VOTLEBvFw4a4ssGREsXcaW3umQ5zuFUTLWp
OJ1shScwKtRYPBGJ84bX59c430bVNkp4O/wusrlCxyQq5hzjIJ3SZHg2R2cDpDtCHmiGgCWFZNTN
YiuR3u8VKVeTcQjJsKE4K3QuBrFmD6/3gky5XBZ/yUn2F8Rz39vZB2RuyH95wuB6K6dtwM+pT47q
gZAxG1moYZbZtrHkJmvgHnVaF1tDuJKS8a368lNNB94BVdKdD+zHwhFjBLGOgNbD9kPYueN2kWSH
U33ImYjEfcx8gTJvEB/lNRkflv2NX2VPraRKhArIsH6PCZIEhNVuY4w3vKygPMCt2bUEQEkWQdu5
M3StFqDs+zORbQNpx6GcXfSBYDvN5lDfZcyELp23irXmrrj4a51ZF9qji2i5iuMoX+DNpxfA6T21
WIa6VWaBQJN37t9ZxUNetcKit5n/DILazB1+YFUIJ7rGd3E4oiY7GLKG2C1Cv8ke5uHOsrj18dmU
H+Er53w1EdmQGYCHMvmmT5K9i4vz2fFgkq4x5YTkRPAUj6w7n1bJEIbx17x4p7wjx4oE2SbGAOgI
WOPXg6RXtypPiGnfCr6/4xRydb7LF4KDgpNBYv3V5BlWeYzlEC1IG8sHkMruJ5JHBM4AlBqx8yuj
nsNrKgKTM7ZLFU2//T/70ViFUrBbUM+BXClUG9ZKhxeQA/7GhUN3LyJwkZx0J93xMqua19c/nPNN
Y9gqxoPt56l5BMFq4xyCWi0doRzuC9K2NqpBnvoHh0sdBKt3jnVnuxIAfyciFSgKFKbeO+JgAHv8
QUYkdEh+WNLY9SWV/t5t7SgytnESDx6w40hrQo2HEw9GlQyNV3yL3s2Oe+g2MCuCmqAetkxcQnLV
PXbpPnSySRjUjais13m14Gp5aJmeq+aubKFh6HaBV3Pb4AOYPQ6mDHLMsMknu7PeUcGqWaGtf/Zr
B+mPqMEFZfN2IeFx72I3BZuuzrFE2WF+swj6oqXjfQ6EMsbTMkWAbLddZpSSq/X2wc4uRH5vRXJW
IPvJww/9qWOrjgs9ii7olmLGBRo7t814YyQ4BER1i7cXfpVj+FI9j2eltYsn1HP3PgWHHoSf+Ajt
b4PFT5fNVRoHV/YkfYsaJ/hq/UME5G9H2Y9agyCT+u6DM9pVsS5QMURAvlhyE4qvYmU7+MP5cC+4
TvUa2A3+W9KB3NzDuMXoeV/bIbQPgE2iDoBq3Z/TzSCinjpUxFP6BgOvO4wXoC0cukElgdD5KZFJ
8TjSIgUD57PT7TUfxIAb8ntOcj7M11Mi49Ebp3bQe5SsR8h3p9FoK6/PLohHeeEsf6TC2ItK1Ota
LSUUhZWcLxnrRvb81qW4TaE4Qr/+eITfZeLE3j9NLP1EaLB3bmB73OE3FyeNf0sZmuVJSaapJpCr
4jjBhLRRiQb3ZQeFPjceAzuuKOax1iry2fahc2B5XvXnG33ab8W5dmaOVGAyam55M/xx3zrmfpXE
hAZ6nAjbXfjzZVpGxbvcSYMgsscj0o/I/OR4fJIn2oubqqYchoioRcsueeHUC5/Om6D4/1dGrUhW
mOOS3ycmXDFr5eBnPNemQIglVB4fMbm18dcFF0rxTpkndTk31SYex53a7GtUaSJboiDS2g0COMhT
HFL3/09WyEbljQPDsHQBA/9dCMGpT6bFALiFXv/REIYa2reCo3Vx8D9T2hhRr/s36YUnULmYdA4O
Fu7aFHASeW4MzLIakBAdEfT8Mlx9cjOhLq60inN8/JbLVOvQ2bLUBOxP9e9orc4SVf6jEtvX1Asd
bZS9vaCwWSiwWINIDTZ0QQTPhXIj38Io1MX9VivX7t4QdyiIqvzjcWoMAE61pMcYQ9PzgGARyw8g
4LKOzK8qoqwKvsjFHItBqh/gBhsQSXGHh2/HMtJJbix9JN7qHUFpa1AojG/CQZbgTYCe0fUmvRWb
oqeELLemyH/jf9PmxAjfQdFOuTvwte3ZTzcJLNITSLvZ7bGxwJVZjuhcIEPORD31xLMoDUfKVJww
s9ZphinabT7okCF5bXaJBr03o6srHiFbK5l/xYBddmrgTmY0eeZWUa2NVXl/gr/GFP5X1HwHmn33
uXvMBvt8AsFuHvjASLLcyB/rYoj1LCvH4CyZp43dhYtCA10yXdrEeC5rsikit0MqfNLXfv0ekyqp
xeTwJBUhP3rMc92Rge9k9kGvvdCo1bxr/a9MHpQHkImjLZnY+r5RvShNj5ECESMgtbrvZVq/W4qd
JNRBaSR1gYLsOcqlcMIjAooTmeJOz2dG/8ggxGWFvOBvvysC1tPyNdgFindTokN4TcUAIXJ5+24l
6cSY+Atr9PAK71nmZoIttTaHbcB22Td44D9U5+WVB15kapxTiIeKYO4HyOsF13BBXGBvtTyUcIv/
kkeW5x23qZANkrA2kIbd/e56DP2yhg+FccEBV7I5c/khpJzobQ9LSM8THnQQzBck3zJeVlNOVJF5
kRMz/Aj/SjpGv4is3fmLW1TR006C7FTltGE8TJqHG1jU+J4O3GRCIt0Fj2shtYUQqAHr9iXGhABz
liBKMSE0ivI4nPQe2WgQ04oO489kLO+tn+C//ItrjFzn351hIQ+EFBIbn63jqj0iCLpuPqTXH0jV
Ckzi3+zcFeIJN3TydZCBig8KPKvTEXAFDcmJlCjN4NOxXynpRmKxj23y7KXmjWPpAUn+TfpqB0kP
3F6O8go43vq4gNQ5nvBDvK+icLT1i/V4fvhG66Gq3k4A82By6Lku7lKx+wSgdsO0xOvp0AiGKJt5
LXCl3+fqhyxUv5ITW5ekHDdk/WTvMtRqmnFhPnikVsYzoyYHWaC4bcTnT+rlde/69G5oLUbEepD/
hdsD1XF0iVKTA7rNVVyfkn/PB55+RXCFWsLPWonHMWG2995oVzVdnTwp5k3c1fV9u9PdYLc4t2Nv
tvn11Ohr0yvLkGRjbW20acHScRSQbM0DyTR26Ba+J3L+YP9LPwmFherDy3Y/J35tNAwERREJb363
ijyq6kq6on9IPr6ZYlblViLfMcGlHJwYaU/Bfd5i5K4bQRlpIZEiQlMt7dMts0xKhb8CBrBi9jKc
h4W1mWANaJZ31w+K0hAT9uXcHko/6eU9PrzI9MJhbO1ekgy3mymKjo5YZFighD3f/Un0eSKYCxfR
sam97xVM/9IG6hmuQGIwead95qf6nQash0fCWa+Y+JwS0BDTsZWvKMYpudMlzBzhQ+tRFrMe8ZfY
41DMPVIP3ed+JowF3YcmRWd/MHDrSZuXJcXT4V+rPmg2jeb0Qq2WXBQxvYEIkPMTPi4fHjPq8yDX
ist9efUu60YIUTO2xTahIv24U02PPOzs0gnoDrpERionJ7MtqM7yxf4v8Eti6uHNp4at0tazWKfh
uTZuw/L9GmoN5A21xouz4dBT/LEvESuqyasVnvQAzjeq+5uSD32uduxEY7k/QcqFbppamCyGgZIR
HfO++yQIpiNwZ4x9jcUNlOELVWHBrGaKofR+FHXbplhdA27Yh5GoFgyfcczSU75OiVZmm/XxnqxZ
SzbHhFOm0R9NPeTexWXwNASJMGoZej/xnK9RZqvPqNYb9jfxLC1KOgfPV04Zn6c14PonQBLgMy4T
Q300h7GBx6icz4eVBB4v1D3OfqK3FdO2irmd0rpavURS28CzIDYwSxAk71GqhRE4wBevXUDJw3K9
bL1oYs7sgy4RF584VRttLxHcuMD3EyD+GgryHjb7+oidwAqSCg6oPwrEhccCCSjtxJI7qMxNb4pw
SohdnD4k6LI3BWl0T2wkzy0xcv8z1XfllkHGzkphqFcWtb/okFrnp8LXR2pQ/HMs9Hv3tlmqUZKU
lrQ1qBzychYgvcrci7TyxPZqtLvBNfjKZ2SUK0cTijaeHHwUdY24hsXwLlyZ4AwRpEf7uQBHqTGK
BJA6gpM7O43ZrpBFIuiB6JB4/Qd0jWsIC7Ufs/TYDZ3rQjQHx27M3JYf6+LCvWXjoSj/B+/YjQ8w
X9qtI4AH7b/qwM0SnHrDaK2rAYFCjUyIN+bs1rIHiJMqqMamrQgHYlW6Yxc7apJNC+Nqu2JL5rQf
cVimV5pF0MHMpbpOFw7Mx44rHUXLQaE9kx/63FzFIxBhlAKjWwwaDTjhf9g4qARB2JPvPlZNrAgO
FXR9mcKXNe+OLwaozaKbUq7ywycyjmxly5+7+RvvnGpEqqwzk7TQxec4ZvPjELd9EWbCCp1JA1WN
Avus7A9O7opWV4cinNSpVICJOU8q5je+c3EqpgYk+AxgppjidLiRMVH0wsxgOFCib6hBDx+8m3EE
ZpNIlihAnZkINS9pXhXYvJRPX+IO9lOMn454y/lIF2WtyKppJlpZvJsAM945UX8monIZVmVFzRoi
yFxDK+0s6lsvA3njjSgIuDc//G6yYZYNFhYy1rwg59Fk7yaIwXd2Ep25K0lpDlRBAgUHDoOH6wQh
IRnuqipzP3PhYIA4ZdcU5Wnld9C00Lxtp5G+tCAktNUGhG7pUn4TAaUah7zDhzkp3VKZDiSUR4J1
r2oVHoRcpCDX2IvSKdfY36AQQui1GxjzT5y6mT90xkXuPkMybvs5aJ11xvFqRljIDo+z7mffwJHB
SRXwaSTt0FnTcDDmMXr6b81WFY6GGag9QGQfCKuPiIbYtMy9AbeD1P4aE7T2cYz9a7ajDfAdfzBc
4pD/e16rVDjt9dMH0DlK1JUXKAdodQ6fXlF0snvAFIPMm7LsZ18dPEuHiI7ufbLixGrRHyUUu0U2
fLycCD4z41eFkCPkQzw0iOC4x7lv+DDrRbfps4vXDs5Jk7Ywmoj146DfxfVImQGScvILbymJKa2c
fhkcZnvItVqYPwSLQz8H/Kfe2W0CBcbBsH6byIe7upLEk8M8HxDHqy6wu9eaq9aS+XbTPLVf22dA
VR7zH8gA0rxiIzHKZA3pVr9bSCi9YT0OGkMVTdvOAcptuMRHSxlncscXzbu8Ma3Zoxpbo7yM/892
fVUbw+G1mvJwCYyNe2K0QyEjALLZp1D/fr4m/TnS9vhqsRg1fQO6I0GdfQ1FojQ1ctnpFBsVUgYb
Dxof1ovvXCWwVBDk9slpPorLD4tguIUJmhagvHagOXRoiXmATbQGu64VO3ye0qsBBDFr06uPh2oy
4r18GIMb68Ql7/f342ld5bmY2VB3hGnTFIEotL5g30fpVRo8qNJ7y/SsokL+RZNj2KolDCrmLhde
6V6GeM1yntsgDKdKAWUAywJub11mHgT97coB0/hAT7OwymXu2LFO6BnNsZW8fbp5+HxrXee9iy1P
C8akfAax/D048o1vvQCSH5IJJgG79ijiKgfwQyHLrjqqBw40i4cKQxu178u42RziEoRLQvmZ4drV
4uYZqhkgQOzgtp0FNl3lNKrtwPI802y4g+tFGenN98AY+3hhZo6b1asTee0GNwQHX0kCODFsSesk
ozmpkvg1JIYpEfmjukQ+4y80ud2FwKxCwGhopJskGJc38Cxz1OjWL+ssZGkF9UeUo2/Y/Br3eQmj
giIacdcVsfg7ZKDk2yoPBEL9HIg6lo+pRGZk86jkIM0ogXl1t1hbbNA24RpFwYxeKBkfK/VkxD/p
JThJFqamYmG27pjo70jgmM6A/r0vBjod/8GOYruzUx67QCnWC3/sI8B0qRZFIiubOe8fpsYHPLdq
craap3enXrPVD+6akFjtYGTJn+trAO5jJrsCBshnO5e/wOuGfvx7neDVS/3F+PeaW7jc3DbjZdg8
o4D30umzMz6NojzGFp/sF1aPcO6DAEne7shIdQXezts3Wo7tfItiqkcOTkBqrEcCYKDl+WQdtSDW
NZzEBaviNLFdoAm075JW/5ggF8behSbLoKfQwjdavXlF2dQm110q5xeEgDket5q4p7B8vD0rfbGM
NPiCANL/hC2oYRWnTBR6ZKw3+n0aw3KciuZKDWmmW3ds4hRfLlDmrnQn2BscAs2jQs+zkY5riZ5J
RJr3U47CW3x/XsZZJROcWIMWzacvYYvPSVDYyLnAjqDIWW9kOCxRPIFHvv/S5vMGS7813fCyY1cq
oEHTgvZNeqPWuPbXeVosSE1emaNQCxophIPiwKNuKZWxvrdJ4OcmROcap5iWR7oGbhSOBw9FH/pb
cUtZlPZsttHdZAxizpChsCQ1x4K9MxDD7rUZSpvFVSmD9oJvLdnRI/ZGh86oFA2yo2iHm5rWdV1H
wTjFPeEE8MWAXO62DV1LyMEEHDQgP2EQgrcOemer9PSaiVQHEdjwaUNIzmL1T9Sc/Pq4HTiTT/1R
Ox/SErpIAcnHOKMPHe8xyE+fhHIP+zN5NS9NVsSBSWs/eVg0k02yTdob+9wH5bKENPfba6bdcrId
1GG7mDzHEyvV6IK/ihYGu+54nYgvmlhupDkZGR85v7iXanGe1JTLvWgIFgt0ANywx6jKswni9I9s
06MTQQk/AgW/jydh1U3W1JIYkXriR1gM6l0jYA+TKupqTRa5/QHnwAN2m5qTm8tE1gb6F9xsFTa4
ngs/c8Bm4LuVM9XcHlEh2CS8OmqWxyvKr8hNl4chjj7VFykIlY2cWyL9lkiLEj6JuU7Dzi3YkFwo
XtGJGLr7cUyHZLcvvQWSOviNnRs3CoMUkcmLV8EZiYyCr1tImaE/3FaVuaqZBsb15LTzdYEXUBW1
CX4Ng4MJchdFULTdrHEwTDZ/v/rcvtJFc4feMyVaOKrBmidky5ERR+A88EQpfqSXhUMmNOron0jc
8ZqjddzQOQ2IoMBrmgP5Gicgz/5p79iO1KlY1/SSbSwifj+pRbUZR7701gidXIfaLQTaB7rHpdVa
bYlTtQj3twP+w7KHjjfwZvs8bJ/MjGbLM1Dol+y/dlJoJGgwjeVhyc37aRhNBCWv2HZy8YqkEDHy
Xy2aSTTbzLUnnt2oLXu9p6rGcER3SMqV6Bs74pM9LhQhPLzS5tlTxJif6OpN0H+NRFyWNHDLkolR
KCu49xgns8Ifxsj/Q1+RY9mg/mXYs1cLEzqWbbP5XJsAgSk/T0QO/6OWJU/z74Wp8ChcwkFF+Qts
td9q707US0de9iczmphMLH5i/ZS4Nzhn5QY2iMoZmW9pW81aLW/C+cLol1dyXUK/Jff0F4/vxYe4
DXgszVxNfvgMkcndSJtByMw053cRD335LuviyPP2L54z+G2OELekatnwxij3F7hdGuMRgjO4ZbbK
/DLET9ew9Ntv3ZK+TEAN5GUc7n6OgvyFpx6VSbr3+JJn96fq28btkXsM/GxsKpG0fisYy+vqCqdF
AX59aR5kzDEvg8yJ3TSFiV6um0qD6vUciYfCzXSc6YNXkYxzK3g4AJvoujSSEtpVfdV99/An98qM
trdioMHLrPEqZe8RTCK78z3f/Hiefk9U9uA4divhkXue9+ml0HppHl46Kaef3yiArQNLKiTTjVEh
OkRLqAOfleXHrjmcujECXDq1LVkbOZcn8l4m84GUgsbBySMM+Ud+gVGPYvZwBVcw/s5/rjUMQ6Ue
uDPZ8VaY46zRFcyHbFvcuXmMfE6exM2erjevH1q6X4G/n9rFVFCkxjh6inAvmx7ZaXMzQ5AafgVn
SiDuUxi3vsa1rCcNbzV7s+6+nbVeFzMuOVCcCGVvmszePyin26gDbg+KxMv0OeqdYcMmnjPgrz94
9DVIUdEDoLZzQIr1tKLVWRTmD9OZay//TC7AxsQEvGQCMNvCP0FiavXLbEMbQi3q1ndKQGqjiKrK
A7l1NbgNNFnqcvTEHyWA4SwT2nFraWdAsQi4CYbw192nTA1uT2xeyVOE2Zp7RriasP/sK2cHgSON
dmP5wkElXN7uHKmDUv2aLWMYaeUp4bF5tKaksEmhd74kqXRxdOs0QNU58N8KMhrD6yc2f1HJ7b1Y
ud5f/WFoEQqCph8Z5ATll/hr3aqHwWayylO6dolRzP8w27v8bDtuik2JRtuZJPkyNiwW/ozbr7ck
8f3zfdPlEzLKgx5h7yvq86fyd6F1ZwjxUe+VafKuNtJNLOcYMOalIE3eT1hPMU9N/GQqcLt7RAmk
rgYZFwi2YE9anStiOKzETmLgvDgNbTzOboj++ufs+j+5BVLEifnGegSxnKQdZWRAlKFpL9mzqBTV
SkqLbrAvWLyxuvcHEmDnyABar6Fs+vwo9H+IuCO6cFMXegEVOfy+rdzwPNrWN0lFNweX53G9uYhB
7YvDlCyzYslCBIwdCNG/jshSFfx9ZAG2Ny/ZgWyiG+X6lgShGt+ijw61qZ2f98pvBkFtdPGQ3hdk
J0NzH1DSfbftQJot57Ip3Ey/F/Wb4zgH46f9sPHztV/UF1ddq0pNOev44/ip2i4n3WtZJhDk2MVd
2npey3Egi8wlhuVkm1zWZPaDf35LcYWg5Gw6TLsUd9sZbj6mCevliqtkQQ7IO2K8oGx5ot+Sw8W8
xNssHHudL9MdHxNlkAgeykz/UR0ghJGw25L29BN7ynNWitSZKZ9SsPszkxv6vu7WX2SRmfp7VOLZ
Lq5fdm2f4BUXXMMWStOoeBZ7J15+mAX1kDofBRNp4/hmajsslmeFIga+NucuSqSMTJQtcSYy+dph
FpPn8Rx4XYJqrr55COxIHhNaJcJVLkTmORMUe7edqFfg/P9TkNjcLWXoRYRX84EvRW+ODNRUi+Cg
5CO8g7j2rZ3QAxNq9T5dxyupB80qV8abSrRbIotMAJogvWl3448fE5OFH+2hUlfDKDK+YiQZcPSF
gCfE4+xu02XAElIVKbnoT1Lz2kywLJxggWnK9rM/xoYCIlB0mz00vdQgY97FuHmfXHjyB6VogKJA
E1UIKh5lNue57T+fych+6oDINvLSwrt3crPJTXBDV/AmascGF7t1c+WGK2r/qWeFyYDwAS5zdHTf
ouYKZUOT5KKVK9w/bsG/gguMOR5e8cv6oeDZCRZe7dgKU5pm/awHPTy/0iHRgbtUEdc9flbsAhKi
MVjD1NT5LXrgL0L0yBD8v4PGuTAsM2qfiFkdxpjnLBtuD3ajsAspY7ZLRQVMQSEHuw+Sp2v/bjCF
sO/3kI176x+pYy0Cwi5bHoZ/0EC85d8AilynfV3e3PdDPgZ+C98wcyDp5itW1F/7GeKqMgTKwp9J
gVUaTRClDM/WbVZFECW3M3STQYyWssz88cnTqaVvTChHIYLRQewN65V+Y9vy1q3aS4W0K8sh8c8r
wcHUDwPsJuDgD6Fu3YKAZwN5O1os1PffwwqtVtl3a2pcOoMAKNipTxLMr1B2zk5kNTnzTVgcthZr
BOIMCFdXhsCS9yj4yh/fIKEpW3BmgaEtMulN2YKjBHG17KzvUGR5nEBDyZSEkLiBmaYMP1Bo5aMJ
Bro/hb0+Cl9c1p1/JoloYW78vcktnKCStqV2WbD5YPJ02ch5nVus5IcL9J29KnVcWEodJC7y/DcW
TtV22hiDSpRIw1F8BeSbxLuPV/lLIZn2m7iNMqh9pWfEEoRGy3e7wl44gzfV+HdpjWdfh98NiiVW
jgFSXwkkRKV1LVbj4hMsxcsIRZozdpbn9x1LPN5SFE3GUmPwr18lT9kUMO1Lt7QnJaIraH3AqOkN
Pla0QSxY7B9sqisSXJAM7zvnysrdD56OracbYpcY8m8pBedMw4b6Gn7eEZghxtj6ckvSw05+VmNv
T7O2v00tMoDVdsEruvy7c5T+zDu+Jq1fDuiRvepeskvgcLafuai4iaD0m3EpcXMOLIMCa9hBcoFJ
3RCQG7r7DI0FwAvgiqiUJHCwVI47qDbpM8WujFF7g5FA5hxQoqxQJdgUgwYz8MwIEAg8cvtD0/Bx
RBLmW73I2Mf/Th1F7sgx7eg0nu6p2z70oGNRECmALOhKEKUqjaHRqebphWN0Cv3YB/GwwuaMbwVT
fOaGAI4JCS6Vgq70ZmMhmdjR5I9v7hnDqECGk4du8V0Ft/yA/RMgyb8TjOvo1/V17OLBSjJ+zc8c
grs3UAuEB3zbKR5+Y6a9je36nNt4sHstgDgPmuFvLv+zu6JCpEcIyYBYd1LdU1ALwkuWF5DYM5fT
GdMDUqsIE91VW99oQMIDiezBxLnuQ/FkDRgAQLq4uQQliiFEsKA/mmxe5JRoXCRfVvpHa6Ox+SNg
cUEE4dsZpgx+W/M3SSSS0+tAFM/2D0UNkF5v+2+L+aeHYxbvLw9KbTtXhYGGRYfwfErDymDqGCh3
hX5UZq1B59LvgE3aO8iSfnjVl0IfLbzrMq0EWXcOCcXhV/HbcVdf1JlPJlItpeBO/9n7qmBxlpmh
mVXYDEAWsJKzLU8SL7E1gQaffGV758yUZJGFaMQu8qvIfIXt/e0Z3f94HEWohchkqliZJmqiq2UX
SW/+VWmJ4SeXEbDn/BFQPur2dcyb+Jt1caoUhv3+HKUF9a15focJGUCEaNnME43JOnmwskpB4mVF
eOOS2uK5GOc5NWxylKvHI7WtZ5s/vHArk9MSn9ESn6HHx/4L92jeaHZnTfHEAvyUZc0Mg+YIBXt1
JsBTKDmIcQoajlA90wQFv15B597EhVxqAKiw4gZ7U6lXi8JdJk8EVDMcENTrTMNCYBaYt09BDXP1
MKYCHJBHgNozTj+vF9tuDfaU72jf9sxL6BLT7Je2nt38ysSmPTv3V2pSkLESAurMrk/90PxCX4Od
M8G80T+OuSU1MO5BBpgsBXvktparn9Pol7u8mP6UFaiItO5JqQPI8GDGOq8zjHxQ+M7sutY0TALF
DlI8Db239mKlgeA0k4kmsJUx953x5iP5uXx9Es9IJVo/LHHlEtrB+41zPwEyoehfD3cO0s3JxzbQ
GzY0JHBOyRKHGF+PlCUnTj8Fj1NceI8MljYMIx/+d0Z/YKk1u1qR9+K9P5CC4rtbgV6UnfebnlLe
NKhUlVHzbXNyWgjwd+Jv2SMvxiEyB9kYA9IKI0MX+PMo1HVIwJnEAMoXgddopdZQLo0h1LoF8wu3
Y4/KSP1KPCN2tV3d6PoCo7CRowa9CTSTCtw90h7nIasXHSKRGy4rETfG5oEVbR1J9Ewh6WHGS+Y/
1P3bH+dwNj0dRj72WIykt00aIAkNKLJlquUcXGfn/SQKgj+5K3iIBRLvZBPvgeIAUukko0pO3Gv3
zXQMZqfMD2vnSMrx/swojDmtWf/NmIuVN12wqXIU/ph6y0XL4kgOGlZer6L2FDCdnOgV77X0I1Y4
byWo2xzMZm29nzWQ33+CZvPZfh4KEEaooTefDeNZYRKMXCy/PZNnI8eoUCZh4Oht8WNVJqh9s3h4
SCqMlHxUWS+QVYo2lrBquH+22EmNLqonKbWRPssaU5ZCzB6fW1+kHYTpQeQzIf8YWRqSXDmcq8m/
YpKlGxTpShPbSeVRgOoj4ktw8O1RhJxOJkuvIMsVZ8/pvhq0KTCTcJWVdmeeyMdO430vrAhUNEEa
OCKriw1M/8g2W9nUZ+5+tPsKyfVv+5o06i/FEZo14D7lPAP4T3P8x5dPQiImySoIDkXoTvtO+x3j
3+VR5oh5wXbquoXp1/JU1N0ae+atMXQfBksE8o6xMzO9W+CgGCjJmF5w5WNvA0d5JZl0V6C3167V
Fg7zO6NX45xMntmlWETgoZVbSlIlh1JtAnDUfULokj0yHQenxOqePkQWC8AqI5E50OWRo5p8b2C3
/KYITPd74txY00vKKUFlBsreP+QOfg6wX7dqNtLZSV7msfdtUT336KFU/5HgMKZFO3CE6ev75sYV
OS+a6NX1aD9AHFDcsSDs4qruH8u/FEwbjQ3tNwsvcAHRU6BPbhgjSlVBeE8YM85wRgvlSoVsXtze
MN1ZyqvP00TX4zpDt8YgEhbPoRu1O3nDErxs4R/te6kJn47bpXUTcNwG8CyzFjeaNaAwSEz6ZXhg
VmhJE+bgvTDDuqGS86ZKyskR1Jc3rElXyfyLd26k6x4pTGUnzrQNn/xrlqNnz0gJa3ohKi8DHJrQ
htaEK17GLIiIU/PjhLyKyeRrE8Bb3eAkxHWptb5jWimXilRllsitiIlsTIQLAJ50q+sTkeLtjhvX
QNTR9fwJRS+QwbQjF79Ykq3nHJRfREwQrpTIicu/77US+aLuSsqm5mSYmijhPLu95XDAJBpYOctH
a746CqICsht0HUDKLJZrPNXiwunX1vaweiiYxetgRBBjKJqEyYuvA8iQNN9UyosRV2B3vCRHvaMU
i8IxEdyJLcxj0UyBjQYZ3tGmZtHWVrvh4hMqfoZJjGc03cjAO1axkrcuC5TWtajocAPceMj2Kv04
y+tReLt2joE4Gtq+dGFnGp4zCAMxOKQ2AC/Tpd60qYoRlCQn6hxv28+6N12lTpFCzIt8t7D67yfZ
8PyHkFEQJ1QBnz8UFGqw5Mk1vj4CKVBIv+/3cSYw1D+/0HXMqPjddOa/1OZoyRlPkcN51fsCN3gW
E7HOCa7pcrDn/N/KzWcLx9efYKhdwwffraR+H5X/35QLQZeBDal10ySAW73m2+FDjvqiotBBf+vS
Ng05ldcWmKvXnNqVT1U5nxwCImC4dlljGkQNm8In81st2ML8GOxqy06i87nLpMOox14fYYS1SXGp
P/zXZ43FDsIMXarHWU6irrFBFyGYJxjKdQhrZ8Y9GhbBxjee1dIyGsdjq0vpk2bpDGLzHaaWH8oD
A3IMPBVpDIZmkPMqFO5xlFJ5oSNnL38Ouc94vsfAc6SrppaV2jwigPRm5Voky8HcODX6Mpmt43sf
l/U4nzUqPO2/c5vK49eVezAsSS5JRUvS7PZPbKFxD5vYgtduDtp36sFMYFd97RSuJ+xVIevxWX06
DlGoGco6NXIojHj33roaE5/a9liqwND3zk/WKopViqbK2bLnNCORujSntQ+aiDjGSMvdSRF7gnKm
FTVvRGfFmNCQdfKaIozahQK5edy1299ml8pHuWuMaO+PTF/ohMAHW6ZWXCqdql86m2btFXqeagE2
hOGaYvmj41Fyyui4fxZ2f9svSu1gNIGSrXy6KbpW0CsEYaDkUGRfLHoHWULdrnXUfkKF0vBzXDiP
BjZ5hdTrQUo4btXostpFy0YYBJldyW0iqPQEL2LcYKRvLvI6qmE4jgU5CdcrZh63fXW0FlDaX7J6
iIrTrpm/hVK1ybldeq0Mcz0chxvBFRibKhZElEzAkVzTjPp7BRKUW8qoDqtmLBGiWur+9M4VAN9O
/8VKeudE3jdxiHd5nF8AGl7XuKS+fl40ZOrXCjs5DMrNcl9a42KaAsyW+ro98ZCAfH2eEHpu6IRy
e8sLHEhaiOqDuwNU09cZUFttB4SohM3z2T12/9x7u+AelLCOiXz8s0yvm5eH4Q7gBB2pEyXRaDIW
J44p1LbQHSnFI9YGTcJtu7VvHVl02LyhFjwmfOSObSyKo7CwhIfxSSlyuffulse/cIJsUi78eUCC
MFZ1ELawL6Zc7O/X6Vt/mXSgn53pS/LJIwVeFaoKVz9ixVLPszbl/vDcdbXvPaoVjxxw03Bn8Lr7
/T5uy5Ni5FkzEVvmf/XjKBAq/ZKbI1EvVndxxMR1a/IR/vwVy06KFDlZag/uqI2dkYdL9eb421zi
2D7qbuiM8aqiS+Odh/netRFvjeqjIytNOf6zszn/SlRLgS1yrCJpiBMtPdDYvdZWJOtssmQSe7Fn
p0Z0k9IJDydRBw4vpzswiEjoVKrkO/iKNuTXeR6nLZ0HZm3qsbY0m9S8WBdE8l5xu7wzDrhzNnx4
7MjQu0YzA4XEnB3oygrqCtOlkmOcPu1SK2x3uBvc0GTx+OiILcBV4h2UUVtUoZvGkf4GDjoNrK5B
6FM8c03rtDy7qacl1SkKpzPT9hpT/LFAyKXVeVZcSNmGUbrUC69oJ9UBM8gDP6iPela7d1Yv7QYu
jPgtFOUr62/UDThPyXQOTeyLd76SSbIP3kUOP3yq++g84NPriF+42+x5OoV5CGycD94dLu8qaAPW
Um+nxLsoO/L6uHYyKPlR0eafOX2OosAS3GS3a5wg6zkYVSqG4ZJh9S35z2z07eQv62pXuMv7aia8
i4MHh+toslYwyKsREF1YyTbYlhof5ncuESrYbuM8bpYB9Xvn1uov1C/zYRh7eR1+W07m3M8Im2yU
XrUiZXBt1BQ0o4x0w00LNwunwNaqmmUD+AbroCNlln+mN8Q1UoAXJpJ8qcHD6styG+i15CHiMWOQ
VvqjxUlUhV2kCBaFUf3LyU5SLZMzNfzLXsn5vyvoQPGBNrBJ8TS0wdByB1aP3PvKi8/UsdIQ8rmt
Uvp6QJpY6klkUgzuCd7j0q9ZCNuoyLaoa6llT6ChYBzIwUJ4/+8xwvZh7pGNxr3AhYA91wE9Cm/R
Gddt9MExayIDLBQ2JEm1SQgrlvamd8iwnq3PVnc4o0ih9IaalAB9kVv/qWHFAhO+pS08dfN8alUf
gWCNFoYU7507CnpzJN8LJ45dcmvuar/bnDqxw/f8wZ6KDs2NwNyMLwedUkncdMNH2J4h8WS4Qamz
zSv5K1xARNg5V/cX+jWm10KQJA5D7UatSLngLaEgOJd99k9VpkgwLUqy3hFAFq2spsyRL6DJM6mY
mJcFE7rg6rxjS8xt6BgT9DR+tgp0FefEGWTmo6CgbpR1HSsBrXPT6B2MGL1MS9wWXDOqBWr3y6CL
jFwTop3q2+157o3qzn3KF1/zzaU6nnHe40Chedp/5bntjSHSfu6mvQPpNU+fqFut6zmYh8InHccP
+V0FHn1DSX51n/GN9BXLevL9c2PcC2uT5msxfbR/01InmqjkMjUC01ZsO49m5SF71pgoqmffvqMY
DUs97KSLSLVDk2Ccrjf6INpw+QR/j1qmXGhx/ZMGtTC5egsUuZVfDTNES5ogasYYVySFa6e8tvwe
hUkU8tvdiSogsW4CzoVhNgKnlvkV1tbTWKbQaMsuuTOSAk6nDvn8yncat/J4bkKq6YbUR9dBmKqU
NAIZCMOH/gOWOFaFKYH/lB2NITMqvuJnq15wNHGUaYSasnC3vxR2FHTPWHeF0WMk2jm7qvAluzg6
o79JzakK2BwCrcll/xH+I7jMYmIAp3tp53g4/Rhi1waLHpBmTvtDq6mu6O836klLuzMYWzPOBrVd
ADw5AtuKv7vekfOCjqoT0z7+YsxPbTioedG1UByMXc3sY1PYC6aGn3OLV4lCM+hs9w2c59chcgyq
UKm9Wuqz4A1S7a+wgGVa+8hxtt7YcfK22wJSv5P8aIRcRXJ2svC7viSYGpQ2+9YVkLL6pn/Z72XM
OlaONRiCR/Nshwi5CoxqXIo9zZ6tRiVMMr6zx/ej7uV60Ffrjsui9moMt8buiyUCDpI4ilIlR2nm
JKBS8PhiIloCRuafeFnRFE13zynPkICz6BXQmnoukbTFT04xJHoUGV4Kley1fN2vC8G2eEjR9H/f
CvQqPgyCGUIjJ64cioRfkKThCLAHmFdgk9kDhu+BqhVRZmB2ZmmEBE5j/mnnGnsF5ykgLEQxi9Zi
i4XBQ0FjHUJGHpYqA7ansK55UrnUdc6jSuIJFMnQqX9CNXkdeDTK72s1YrtGz8ZjQ8dZKk2cubWK
jn5H3AE0+s7grRzBrhQmE4/7Zpg1lpcqJWgj7XIQL1erjc5Hz+kv+zA3it91xYGb27MrbSMRucUO
5XjeTOdMLmYVHWTsHjJOPZ5IBf1gOphFr+eQv3caiYT2tJsF4iZtBWElJFsBrKUKh8NFy+6IZkWg
Z05GhalEWtb1JVqTJ2iJjaA0/r3OKTYZHAo5EF8O1pb3YJxjvU+3nbAqH+1c9YPgV5xZjJAfOlr9
MxR/JOuHWPS0FEW/NrVywLoiUOeFVET+5pF9fK1zOmE7OKtg/D9ejTRRdU7G4julY9QDIz1u4SoV
7G2oKOm7WrE97k+FuoInAln1mhBhm70jrkV0PGzDPS3S4BDKWEr/yGZDRdGvIgIzPVX4Owv/Kymz
y5iDOb52qm906iSdaxM90bFMtmfL1usbnxj5AEZPMBfo3cmyXZz04UnSQ2FKMXE1T50VNXfPOG+7
SKCUqUqafNB+xU5FE9cnARgx6SVPpmJMaMtiqEgPCv0H0NwmIkz0RR3hBZUWZqBjZZ1bbiWoVC8+
eJ/ezo7BWEQ+OUnIHX3lewUVMk7UxA6bx3iC+SyLLfQuh4ic4bcNt0HAOWLdYQ0UXPHSJ6HTkYeQ
37VTnmNjMKXq6PzFe2FHj7ZSPaPKZi/wyFP2yluaFn5fGC3VLB2NBnphSWIkyL/moNhoH1/nrtxb
dQ9apX1w/VVn840jptacUYaSA2EM1ZCRxvoS02POxwUKYPvfOYP+9CZPkQj9m9w15SBSGg6p4pEb
4bbU3mpqYcV+2CASQo+ghjKdGiSh7OBN39tl3HH+Pf4a7aTo008NK9/qk9UnRsTybj/SjfMbffoQ
IgnEsFKyXQWZY/Zx0qU+GXMD9K8KJPEQPnEBTtWoyqoU3k4NAGrkmGnF3JF16f5vksJ8ofdA/b83
94hZwGhOXwZj7sOg15kqQ7Wxrj7S8tgg03QLvgNTn8cq75V7W/hTG77WoNBOFeX1kFe2E7wV3jGW
IoVshgE9LgRPNegIWxVtTzDCX+9tTCLNMAOIRJgipjG+9tI7XW7o9qW6LTAC7BwpOZAaNORy80YP
M/zzFinS3OaH5K/8rzC5wT4KLJ4UC0DXfNo8kZJhS8Jpah9z/lg9x3g2g65fZVkH4jTs1RibVOVe
n1fYP+a3Ht4WpX0dpmmu9Dp578Su4CG/1D0pIWJNmFY9OSb8wqJDQSy0A7K0vze7mCgNziQRfYS6
4VQhoobO4VHQVFGbTDk1rXsUynNuP36R2ZidcG8q2fpsjeCfAVdNmxDpThEjxGxjGyVaEho6TNTF
X7gdM8zoyNAyooDejKYD9Iz8Izn7seNxhAKC9DKm14gNf3C6t4IAHNVxafoTv5++blch15MWRRk5
/i+3pa02JHx7mKfc1ddS1W32QeBtOaE/M+qQal3uAmrnnEypyWXwgIYGT7JfiNkQdZLEL3a/NQOb
1nT2avhudQWTKVjwZAnOZKIwWFS+ldJk97Xo6HQtywlhti4PG5iXZnfTduNavV4/TqnHZuzHBLuR
hzR4EHxTU/U5etgxef6ciTwxd7hKeSf0/4AfIK85BMyC/tmUHW4uu2iRljRjwwh3RoRh3P+1SwvS
PS6yTs944+0SgdpmKcnQDIewxsPiindRVva8dbELhLNWNTJFJqmx9dG3p93Yb+Au4wfHWjyxvlrs
YFXy6MfzI5VgzA4p5CR4hywkbUKd9gGXW3SLJ/FUf+3BCO7pmUB0S8S8fcGTPXtBtIIQtad8bdAY
DznI1xbyK+qC+zAayzaHD2p4vmHlpO8lpWXn0jPynviHMy8SpWNVeuCI8NOIj4oQR18bo0qsDvrJ
kAl/PsfHpFVyVYbWHG/T8ahaCMdovW3Pnh0m7y3ro5WKgJCuwDK/442xU6FUKXXymHVCOUr2wDGf
IUvkF/VahkCrijFfZMpqd7UrB/FaMyVCjSf1e7sCyU7LHgMi/mHsa+IIXtH31blr3QN04Lg7rH6+
PG07txVvSS7S0czaBONg9TJdiFmNsztrB8IhGpockJNEQolLFLm5BIcUX4eZv04SLKvvYxXfheVQ
sU0mmuY4u1515R2ngTa+qMsaz3gpYylMg/keq4Q18qGmQMkZSrTlV2chadba4f5gPbKg5Lf6FP/d
+uQIVwcziD5Kd1FviaW19pJEfGZGDthf9I4XsaD32drksIYLsn67inzO8LwaKPfiqAnig8qKzk/+
nFY8DdQD/icfXkhZvYR/FsdBGUoAYQJL+hK/BDAcKrBXIYq1LLNhw39Qzn1/qXIJ+CPKFfvvSIWQ
JXe4r49dkK437DIha8p7Zy2a9H/bgB6GLbGNvQx7/Z8BDuGxFlAFRC8mUKIm7zNIJ2UcxjY5lxIQ
76PwhFTDV7NLBlI9fLKvxylewa2a4BNHm8OHi3zxhFjb+6XiskZsy3wVA/09vpBcieeEnX9RHGm0
7VqanDHId2lox7ek5kO89l8Zl7OH2UAKJ/PqDe/TqQlDrSHOnmU6tXb2CkDUYVdFgkwekjw1bXW2
tRL45SAyHe7B1Y880gJu3nCGcHlRfUwgEDc7R+jFNeRCDFiGH29cAODcJCOHg0vC3+iRt864QzQi
J7G7FzP/wtPXCvJoeFAyGgphq69+I6IPon2qciyxq7wu4P2kjUBw365R1D4CK4IdDnGLytYRHYJ7
mmuOBz2El8C8D6dDLyNGLkwu82GuBRf62CBueOLkWpw5JNJutLasEeycVC2CuWjHxPdr+H+vSnAR
+i2NgHtRQVo+D3q2uHqh6EByc1oiEXG2KPxK8I1SWUiabkMjnvt/YxKfMX45KIREvl3QSdEn6sRn
4Q9wloDpdKHNADv29+6QasOT/7s0vpi6XuM9XrrMwACDpWiJ3Pafhc6ojz+3eveUrVfwMoFoODQA
XXzi8y1SzNSvMxOnHuzZZ+jhMNBClTScNkMtiVDdG/E4Id/dxrzWbZcpw0kxqPpbK69xqzDrKjuD
U4vKV4gZk5Tc4QpDyHimRkK9LTyt4+HNA5aabta3WImsi7hcr4yNBenxJAIZsrLQeVViV2abvDWE
vkGm4N+byiYlF+LImw0QcuFcdK0q4RWrp0KWyj0FEuHMKwKGpA++xuCLKz/UvpQYIKzyx/TF1bTQ
EnaXCFVNI2lI5F5gvV6pkZqtVNxBEUOu5kEdx7NHIfg9XLKBLxzdtXXffvi0yB/uivJqgyBXmogj
zkFASjuu9DVSKo/2IftdHTyeJny3YOPmyvWK8Lcprml2APN+0tQE6JsBonGemSgBs8fSoVBi72Az
r8R4nSaZbekXZGWKhXOE1kMpLsLO1CQs7bO3h6hHa+C+76fJZpURScpdoGBOjryl3Y5SLoTvA0WG
mWwbXFgxxG0lHTQtBkbCxTnWIPc1nYTDcwqf2B3qPQg5cf5WZ/1+mzJA0CUtNVXUrrjOHS3WIPUx
jHe6URf+kbElL/Jyyy23AkrEwoFEFMrV0xmJMJhRNiM0jMT0yRJTkM2CfBPpdDtGQPDwGZrKV6WL
RR72r3FqWh/9/DO06ULxiuVp0jbVIwYpBE1tRdwFLqDzO87tpGtfK1hdOUudksXMruqSlt4ndv7J
FxQTqzNNtHMJNlLhxhy81NnTMmWKWkD7qTu+Y6ELGHQRJnNnJoTdqrRb2ABbtVW2MvR/ruJWb3Aw
1X5gTxKJR4ZybOcUbOpqkUMaOk7GVCRVmhkCszB/6/laV2dVcfFIgIFIhKcIXnjbCQep98byqdAL
bSAiB8pLRBU23rZjF42ugMPJvq7cKc4Yoj56wXPGOXwmnnaqi/aRhAgxrI5HK5Su4oTiiSlDhZto
zpxEW3lgyDFVrwTWn9W3+sNuSVdNsrg3pgkV/HfA0hIGARv9nB5ZziS9W0EjdVQb5lem9ViYxpas
gBeW0iWVwf+vyuRYLKUtYtS+Bpo/lRaWsWaNR5UpVgFuemwlqcA4TrujRlR+HsYzFHCb/y7oND/r
dXtAODo7QNKTVLiJTpkI6DUfeejdAPU4wJTu364YiATtt9S7uye9HoGVgyt+mOz0lWCWwlUTs+h4
AxHEaXhYQo8t9pbc2YNURM/nLMtNyn91WRN1KOBn5tppoNoIRB6KZis/Pnt0Aem/AUhLbIG3ZvTP
abNLYfqYQVnEJS6VAMCznQ8FfDwD6ZjWNmHtwtKd0fssi05nS975MkBoeEjBZ0Om+5FZgpS6rxFt
4qAYqmf9mPg3l8/OVHJIPSboSOw0pCoKyQn2N7hnQOBulWX6ardQXv1v+tFQIdB9rq0lrSLIVlvA
ZkLLfTLPq7g/rfjrhfz6VDsTlxOrI4HmOYQDcEQtv4mJ1HD1jcyUhWncfVS0UQ4fs+yLp11l0B3v
HIGCHLG0fQVnBuiIPPkkcvwdt5w/CK+Nc3G15K3dp+HWdpt4ukByz0ZltS6GwYtiIRvNAlBpcuTk
G1I9RMBJM6ejjuGL4P2/DFpuz/BWWRpilkI/RrLIOLlvqTbQxTJQKrzyrO8i5WBjVJFjwV2nBXdJ
kO1WFg/eSNh1gI/giD+q56gQgPtqC7k9l/s70ilMoAcJmIjx9mjfP9AX7Q4LcKCD9w5g8laUdMxw
Ly5wM5q21gb1ohTV7g7Upw6pOQoSrepdjxrd2Fl3vklMxz6oqMvTik6R2thJOtZ+lWcjTA26AXzq
xRlQle8o8dYiXYHu3zM8parKZ1fT7KsGRv17OmvmID/COxk8cy9+AsQd1iCpcaDonAOmy81Nt5oA
vi4rGIQsyRYaLo6xMb55A9AOS6FLcVnOzV8rIexSBd0A4nbZ7HPqahz0IfefTbu4GdWm5Puydo4l
AAi+lCkHEgnlsJw0XClptK6jEX9XEdFkFxaziE71EazHIELBSsciynhLuZgOP/yDuqi33IsBZczy
/moV8xWSQWZNGsLmOfdf9oss3Lpn0gcsWvVo9VLQjlFKvYCybh6rq4/yW6iU1A44Q76B+7HtVeAv
WkbArqyd2C4cymv3hNytv2av/Uc9W+lqnNUn7nbUv/rwVSzn6YDPFlH434QeUhbRDgcQvGXYqXZ3
MdDi7jHsO+WBgtYT9QVJU2TrNdO2GcrHcSdJ3un2WKZBTLyaw3FBNSW8WfmozZfRyD3xYSQ6Nt+f
T9xVEhNdymdPPxRFjDm7fDH88BZhl+JkQILB4a4oUICA0ptuQaUBC6V++iXxw9BkqmPN062ouZTC
wYBTJY8wd5sZiAplMGt44LZaLZhZnrxZV6FhwQeoyWwZZZoE2kWhHbtSYoF5wjMEoFJ/m/jxP9dE
BO8QpmOL8wmjhrBpaTF1oHqWu/YnS79711IhHDY5R+c3FXc1CGjK9w/X8QitfTmtvl3Ou2IaO+KD
E1hsdgpFtI3KuHZHyygSbc0wOjSHOJaM90zEHGbCaigZXFTO15iu/RLNaJu3q1cBSgVHZTqDOr1P
WsAy/ivkmef9Mj4XHazJbOD/rqC7Ouo+zxqxEbut39upnY4GV9qBQ3O6K69T3YDXquyUObVUOIYp
H1vcOclQ2/DSA6w+ni+mpKlZjCfOTtOSeY1EQ9XZLiL3yS+e4QABRN4PWCQg4cz+40EsuhtrDvak
fCNH+Q5+kUvQEXCIUK2zRnVSA5LKFgyGpV37bsSa5d00luKRC8ERaq460d54j3tMN4cC1GfnFUsT
WHRu7GoGh2PPMmd03n7GOPqAuQOFdEjSOCAvUlkbPISLGR/2WCXlBVMhMFg71lFZFV3wKqpjC8Zv
RpiMvc9HAPPGNO2Vu2kgWN5asCj6EMtCL/3h/XYl5prEmXJVXuMwoLYQ+mSDOPV5f/4dLJzLbwc3
uA+vdF5Yzxvfw6Nx3IuINpZeDzg4+XO/783LgTvbG8Ru51WkXuMD0eBmiJR868JU3k/TeWRmssFD
f3gSLPxAEXLnFPgvWxYWOvaZU87frsWWmogpP4RL8RRULyleA5v9M8oaFgT6ZuPpF3VuxdTVd3aV
4TlrL8tPDxcNcix5sBYCcYMp8fbreh6kk2lBieNQ2/H6vJn8EjoyOisH0HdWbGk0H+GB4fTt8NXY
83d7AOne5JUIU/cVFFC1yMV1z1T0s63jllv7p9THsalBQvqB3VLMb2GElPmZfxX83SU63m/K046O
OaG/tnFZrM4fpNsiyyfJWzca6qTc/5HXdYRLNnMLzzehuFf+CLvtj6zLkU4rMCxL70uMHbA83Ito
VGM5cDMC7+PxRF5bjENC+94DhCaEGd4yybI+NvewbfTalVt+JtRf1Xbm4jzu/v0EYhqj35Ejpgp4
tRbDPzZ3f1MywTglQ/vSw5eaQHXOMNuyy8WTqV1EZQUtXT2Cn6kMldaTqASfoMx2Wcj3yWNR1nRh
60rbA8KpJm9HEhEab1d8KgCw1FdYPK/jA774xzP9e7DgkvunkQ7ndIta4DvAz34pAPc0ta3qenIx
hHh9Iel5IVETAkqurev6xhJdqo8hd84PwuWMyVzfj/5fWq4d++4jkz0DkLvflZy8j6J8ftMR1K/o
Av5ZmG5dsQs+JNsJ/9yKkJEFQvLJguaciA25VUrVbqm2gEQH65Fyt3nflDWjVwvpQXk0y1y6TaQy
rju+qVvyhfeD3s9ya5eOsN3Yv+0N9w+hz65g+g+gbU4fhMp9dMI4kZDJeV0aVA1Umbpn3MrcIM7f
ZRD6LZpskHpsd0aRJy+1StznXh5lu3TvjY9KpDG4T6bslwUk7rNib32EQMFIzCOROP7LSJriIO3l
pcuznOEdSpoiacIBSpPfub+raxf2x99gpN3lK32hHvv3xTjgJ5cUW+xO+9k1shBRVIQZTiL15/xM
4JsCO5qkiins4ErKTDmPsrJf65RE4qtqXB6Nymd5fih/bvFuj1B2NtZyKNcdlGHuTBgSkPnuP+Uk
0f02ayiNg9G60eVYJ2EiwL4Ijbx6u+XkcFjHc+U65ekSNbmxUjKvEYIcieNR4PwSbfrEABPsMU41
F6qs1uHFOzWqvX9tyBhASENOIiUq3qegHMn2+4I5FHD47vnmVijDSIQxca6i2fFkxnGA2P7Xdimw
sw3zP8AkEZ9DL1kWpRTyCIxD1VxBLZ7YSeD0MIEYG9AYzF4spjQ7mPtMwIjodenVqYpUnq5djlbx
kaUeTcmvO0Tjzot83MVe47Yyl4xqITqVi1T81lz1hbvHY3DDfPcndppoTu8UNBgEHPeq7Vxg75rQ
bChpw6fiKwiCbFncpjFXdhqj8R+JVhsOWn/vCFl4yeGmhHzEeoci5or4ZdCn5kOZQCkloT7KUbbz
SfJD7y17Qp/JUIY4/dopGCMtEK9Pm2UkfsIWf/bMX8xhx8W5FgWaJK6/nnnvFvsUs2qGOf0AGMGL
NBKoz5j9l4aU0mfhV75NR7hGxQ+xyuSA8x72sG65KSVOk+MKS3LtWzMaGy2ciokBxVEtnUbzSQMU
UlrHCynxtlO0TocOMp3CiLxvTyRaXCuV+hNHFuKDtVAhdwNmVJ8opvCYrL7qXjmFuV+JkNtODpR3
Jo0FEA9qSiYR5tf3VIj/xwM3q7J/1btmCBYdHUdiFlpCh4pkCXf1fu1gCbf0iPTLdDoTNPWEv2qx
eFhHYtV9kv70UxCuLPMfmwPxgZnXfQcl5DMhTZcxMrrRvXJtwfnvaqR8rj999KU3yu7ULUjERa1A
i+64G9jN0r9f55r+GcwoQG4vNg6kfl7PNKz06DcExWnI0arpdW8VK+E3P1s7GCVEhYmAcUMEr3R1
KwGdrgHPOlOH7ua7c110kvAsc/tdHaHuoCh86RC/MI1yJpRH5POYmXkzHWCizIii80GUQUGVsNtd
xy/nG7TLZfVfKdlt3mcxV6s6xbv23Tc5CUt+Qz8OK3wS0z9NgudVSIL9ZkihRZoCVxN472xqg/gG
oimJENacN8N+dn6BPYa6c4jw6EMtlX0JrS5loi/7eEf4Ib1zB/BLEnAaRAvasvwGiGRtw0/KfboI
L0a7ATpbriTiQ9ib9TUY6XoYuexCdYwOlausNk9tYz0LmQUcg55U0kE0DUzEQ4rOE68EXegbOBUp
XJp2gYt82m4SK5o3flCjiN3CEXQSNKl8gTxz7GKAMMv9wW+sdWTLz1hNCxnx2E51E4EaoIWRmXPC
Xo+II+0+ndzvYOBHSycwctqc5fImV0AGbW6no7r/HsZlGbHuzAfeyHpFrJ3ShL3IOj8zIFHCciXz
Sm5t+uxIRDRSPkGqfdp4nPEf3UdFDOWObBxsSrNeQrhDQRpccUha3n6s/8pNgRYT3iOmCkn2syoE
Iyqrx0P1ZB7zLQJvKNFHFF3hhQiZ9ZAHSExMYmypOt5qZR5Id9PzgXsKBBASstddyh3HHiFkRQo7
Fto9e61Kpr7ePUyRrbUhdB3wW8dgMzw2dsVG5yThj9wyKQXCEcRssAKA8irNI2ZDnphuyFKbqLr8
KsXNjiEI/qx5fxW8IwFqwHF0QBjHIIZPf4DtY7pXeBmQ8slersaEQ0yb9Y4RCyVWaO8rr7Ey8Hmo
NN+p9H3DOdqt09xbzpj5FM9ay827L9KLUNupD00DdOQvWfEK7fGkbc2HK0qCfCUuWX1i1UTWI8Bm
afOUDfI2sx+H8TrGcyeuUjdE9Sdtfn95wRq4d16WTV9ftFvQ8Jss3Oz8dwgmANQvKK355f8cI4ot
Yk2ceFHh1LiTym+a0oDOO1qY3f/1wAvd1w4Gw5PQkuTMcjhEmKTrv18Cpc7yR68/g9nPp7DWTgYn
moPQ98AlpUkiAtPDvFZYFyLlpyy+7UkaHXmOPyO2l6N0/5P6fQK1xbHCQ/n1ijd/a7N+ccCd4NT3
N25K0RrxFkVXjROmEpwCAgsWysNsrICt111VPyFADZfd5jfBtHi1n1BWv7H3gYUhtpUHToCUAmpw
U4ByM1FPo5UmO1jM4Q5uUBSFLbAt1mYdE1t0WvtBZ6o2x6UWqJQPu1PpFmT8x2uU3XwzRPCyHq19
3pPBJI1Yksywtob0RtgDTi+yEF5gK7b4RkxHK5DWEWJ5XnCY/vhEtSGxqcGJJ+zgzcrAolZhIYi7
jbJu2pcrIKeRF6qv1+AgpljVEMf5QGMird3RfxnF5Ij488MoJDWFt3HsDACxmV0xYe2M+6b4b6eL
WTBBnpGPElMDXIM4BePd2dg7kVOMFp/Dqrz2How39GAsgQQikCqfWyMvCtGzgPahfevQLUTcuXpb
QpWxeFqzoWPSDs6fq1XCkf3tPN7C104rV9N2r1lHWhXzax5KM7lqXfN3iHmlAOi31jIUOtKC8m1G
4C7xLR2k8IdNffuuNfR9XxHSb17M6qxl7XqAF0yycjEaevRZYyZ7R6t8fIEIzY8J9bII0DKX+LK1
u4VEyQ8f5U00gUIEyhQU4rJoPbO7yn0F5TLGF8EztR11LsME+PTrorM11WmlrnsGmJ+w9dJbrWVz
pu+LO/YZNaBB/dcVY/qpZuFJs6cIm2AVaWQMVYrSeuIPq3whWKikzucZwYLMRlf7WUHZK+Lz4qm4
9fkQucm7JKoj6rVLgs0BconriRz7eajcOD6JCfHmgq6VpjSVtO1hgDEBYlJac9dsQKYZurMD6hVF
HvHLNRxUd8r5ruLVUUIVgay+BCcMhdyIKxE6Oa8QNRdsVB7/rfjSYMvrymbpbL9FvYZ4U3IjMw1T
IJA2n9mD9V9eEfmBWPa/V6vSJJ/yenUzjjoRJN1MKG4VmZCLTYU4w0DqlBx+U7sJ99FYd6DjOFEj
b+nLDd5B1j6AOUPnt2jbLgnpzVYmALhobIvLUscSo7m8AnDA+VvZ8gVzXEwIoDrX5ujx1HF2B7KF
53a3veCxovX+5tin1iIK+7FVTC3u5cq5nFqC/ETcAqSHqsXgm/VGZPDjBgAlyry3hQJl29TosODM
9rRecgGK8KlQEtSlCPtzRnZX/mGtiWKYK25No2+IttvN5SQQO65ZG4oDUus+vWdRFq3nU6OlGUbO
l+rR8sX+Caf9JLTEal4W7O3aTvJmskKCqmMeBMVdmDfRrfH8Yq0TsiW0HZVNLB7lICAv3JKES9xS
S672UdNp3C3KymN7ClFqYycGte+IdlLjXpWsmJBaZMjkIsOZ+N4xCmPGLpNlOFRzIC8uRYxy3RRE
sbwcngtVBVl8yXtiCgabK+1IDBd0zrCfz1w3I+SxFDNvSyt8oJ55Y0S2CrcSQNpEwo0/VsMJQzuk
yCDXP15nkclgRwoDARzDMAsW0PeX9gVEBj/UR+EFO7rgImIUapb7yvj7mvZkeGqY6jl1WfOxHdWJ
O+tPqCjYeA3/60TK1WTnxiVus4oV/p1+3MkoLtrm7Z6zIRT0LcNZ602l9VGegytxf+kvhnDk2im1
v/FyXsWWLLjNZ4yyESGp/fdzFk9CVRbFTQ255/77t7b6j/732IgmThVgATRpmD6juMpXMHGrB/3C
bLhiet/DYoBQ++ys8dv9QglcNduGToY7vucmLGJnBhVJ/A2XFuqAiktHNX4isZfLGsmxlmBzODkT
0ITP8JGIHiQlCp20+AWLghZQnei3A1/5VH55zfX1wvS7UcNHp/vRwjjthvU5FNi8/834+mTfN/rv
wKEO/OWZ++hrs3enu4wqQR8toFbIXNuHRczEuHUwRglqtocRDpz7vbV8WyqoHbiDQEl8P6xr3jGG
bYBEu6y7QIDyvGCvGDINg6PdJveydTYSXCtRU5aZE5Czp+moipDErCvENaf1Lny9X0n8gTaLDuMy
2FQauv/CN2iwNkwThAKXuNTqDFKsw0rkCZebj1sP2QjOXhuYosFSy2x3xv9o9uRWN99Tm9Tenikh
Uu1cjD/3ATSV/AqXxpYlV39KxyXc+6XVSWupUt9MKF7w/cLOmnjTeiJQOJv2fgdduo5ml8oZqXO+
yACbEvbMa+qh03t7xLyGD2SNJyfqlS+9MyTtjO/XK2mwWEpMCIn090RSbLyahBgTdu1FlJzNwBQS
6wCNhu31WrdgqFm+6h+Nj11A6pkTrljpEwQ+SLuYs1tGyDpsPIw5jq/qmYWEDHtkzgQ36nEt+TDp
hPPZv6zsDGD2n3WSClsvWGmHUoJVluMDOmC9W7dAOtSzNZ9aDulgeCcW6Pedmn1CzuDN5xR6xctV
pb16pmb8U6N9sqDAeey/sUb4gTK+Ea6216G0k0P/UFzZTKUuhOjzu2OjpntoZJFJUxFyxt0N26m2
E1OCn3aOOnEo0eRJdSPG9GfXZfUNvc+WRrl6xPlvRVuMbUnrxZbwAqx3Tw3667Qpq42vb3BN+RWp
9iw5vFjaQjaUj+uRxtt0SRZ+ptKJjeJayW6vI+5KhVaArAnBPztcsPr2usfPkixPTrmczM0P9xcm
Yw5tZcUY/bAkkfEqL5C60yjzx1lmj3RGnM3ZtOswcIklFbal8igV6uhfs3+kVhrYcu47iZVqdKhg
F+4FWHib8aR6vG8WUzjpsUmKqZhsAJSTyX4Dzk8b94BeFfwdyFPlutXs+6OuCCmKfShLPhIA+jNI
0R18hMvWLEvDxyv63T723BOqEOvjR+fi0c8NseptA2p2B+EVP88u8MvbEKKizcK3dqkpVJDvTYgN
vYruK3DZ45756Ogx9c4cPpry9tJpZHWSqGYYbmWNeBo+bYORV6WSr0nZCqIP5RZPJFRKRSShLJa8
fpIQnJdGLxbkNPLe6x0xIB6jGmDnbxAG7PeIVjl2Fa6HW9cW9l2WCT2lds1QPLlLoRuTwBbmwyrO
D1M4OFLyQOfySUQGFAmitfv1b71qDNHavBhattL1wY+F+xBqQ+pAthmgvFeP4XCxtaA/JJQ4k4WT
Uf/RpCBssvW2cAgY+oeMUtw0x2aCnRFjzXlJEzWaNhdA4OZiivfQZ4QsiBvCU/fhpv+WycHWRd+s
IovPVXtrByKEI2jQwtXx0MIGUxNf5zskwVDXCYyP4VAIO6w9Yz0sa9V3xPoRwf1UnMTDp1O4rb//
m9ol85kOASmRZZ6aenIo7ISft7oDkKIK1aylDH/7+F8SUUvJeV9Pwrbh7Kvs1SWVRV/GS3bkUeF2
zZAlqjDGqcbsFeVvkDe3vYeLVxJIWaEvvp+Jm5yvFunMLxxt8Am8BXHR+Hkpq3Updzidki+KWOJG
ngqhDJSid38QgUa4uuBdPo+0WsfSyMuyAcQxcuIq/8H/yyYqpqQCGZxaip1sc2523Gad72t0uS+F
F/wwXFt+F4GRINNr0+bftTTp/mikdg8itnFUX3G/NYsKEMEAm2bxJAQSDa59yakhsTh4YLIXMvy3
tA8L7BRLV3BfOB5tq6mucRW4h3xNumYdI6hKimE/XKpY8CY9GzdU+8QrOsLtT4gY15caPtgQT4ZD
ptzOZQ9NTfL71zQVpKkj2WqHIIAI4qJxXlbM5vHBjfXFZd1EvzkhDv+eJkGNtdfz/efAYPakArV8
hc+SISmI5qLy/NRklJIBTP80efpOQiUmJpJV8I+nOEBwK1TjYb6SJa1RHJrZMDy2cb9Ti9ebYkP8
+rBXUs96kTgW4IBPER+pEegyiHjm5QNHCm9WBQOYOOGiHdvsUzMp4cTlVQjdgHXJRSaqsJ3h41Gb
6CSYyv5/CxvSO+VNE7q0q9YFToW83x/eOpaga70zBU/jHh9hpX5sthfpcHL/vYb7qGFxDqOFP7xY
QjCWdNhaU4YjbjGbDw+K5yR8rNuogcWpGFuytZVF84+369cr3UVP08Bw2/7RNh4dyT4XfY6b8PJH
Vd2M3f04HSR9GWz9o9OFPPSUxJruLb92KIC2moLRH9I1cHwkB0o+2YqPEcvqRu4O7ZDv/zieCvMM
g4Rmn3pvOPkK2og17gVH8+5eBsWQ7lB8SUYbEZ7efd0Vi518TrTE73GSdxDDa8WhLUWRcMGwwbri
UyZ6TeLeG13akmJz/AsBZs/uEyU6BA18+OkpA+tzGMcElhQKe4mSCLkMMWe5T+bzVavf/DDzvRym
BIHsz8qGgLDcbupqchU9nAgKtMNyuMUV+BwAIy0/LwLk1R6T8XStkrDIccIXZBg6GZinR5NJzHxi
rgV5udJKkhfvrP3oLX0o7WC6nWM+XwF28x77ibOJaRU6q3Vc6Hlrj/KQBGvD+EEFLWvujsTy7LOh
8ns/yZc4fpyYVZj3m4yXmnB+QO5hsb19TEP/AIbpS5X2jKrJxzTntAzhPnQruRdiaCTMERO7aCHI
30oU+tQoGJivtzztTzJU50L7YzRrwKwLKbbd5bd9CXSFpXFTYSH6zqCF1EZdjKnN5ANgy4OCMYv3
HcMmjt+noVmnWIR01ZwdZkqrpNc9WMeFfEKPKQcloNknLmAAF0iGCJlu8Z/YqKgydwsCtrF6itEN
l9mHNNqsVyu2+OJ97PXccPmONPVwpmm9CivX0MmwuHKU5wgmkvD5YJb2cIUFg05mmKNgGVqIKK3B
nL3FWi33tALrUPELR1SIgLhB/oJGuY4LjtQqBWTQY5iQfqE/Do/y6lAT4I5DIvBQd/SYXeKKLftL
4y9+SKBzj2rmuJCcQlIU+n2o189PLNFJoFBspnPFbyu23TxjyEnAOwoP5nriixDLw2MTIsW/sVGN
W+Bej7PvB9dzMMrRgUG4WT66fHxsjeVgCnJH/buG9nYkKd1DlzhPB9VILG1QO0+4QfNf+V2uYKJg
CDlwbOjR3za9IZWsX3vrIq1V87uY9XePZC7zt51PFDIDBQVhKXCLmpBhwxHUdGbVl6Bq2ZN+zibH
MCI8+SwrPftJALA8mlNJymrWUFiEZc4zm47ibhHbmXFQPDZ0B/XJTTKMYcGhD06AmRI1Qg4/Wwv+
/YiZT11THvIswjpf/TvybXIFlNrR+j3bBfzNjAOKwjjaEF1BugM8RozEO0asrDTixMRSkMXNS1az
roqOBRf9AzwqA3ZSFe17qmFIQ6c1/fCLH/HSf1ziY1Nw6HHT3wJ5N8CAc1ZlYsqxot25knua8Ktg
H28SHWEnG54sqgUe2SIDtnlI3vnwXX/a/s80JPqlkZjFHig4GrAa5wAfL+9b77PsLYRbD47iJj0G
0ZyefvUhem1jfUHmFA/amlAACSn8xIeHCz0dGM6r6u1/Ar6n8IqAxKUgen45KpQO3OmO1jMPAedj
tuoxghAaTvJ20pfvOn2oTFvUl3H/zfsSBdDC56JA/APIwcxCl01QJqhxx+AH18I21ipxYDJRjAeT
52SvET4CLNRnIzVm4ilUKods2rl94IrSKIyDR+gbRSDAiDi1S7ifHom5Y7HHYARupV/pNJKo35+0
bccEHVOts5R1oej8Zfl0zNdzbRoCEeJrOnPUsUaJ0DS1J9bhRQ4pj4O6QZf9yPz/vPziMf6MMYXH
hfjYrr4qCH2AnBPn/NYuFJo7XB5gLOmuZFnrcPpkHhyz3mTPjHSWoUMsxKkzZQxJoR+Jh6NqRWFw
BSGoeUB8egq3LFMFQAAlRAtFAtxt8Z/Cl4ne2v0ycFwO1z70Nd3sW6D6QzyrzwF26/b7j8urDytH
2Edz8eWZ17U+lQnw055nn5ZNRGyxQEyLICA4kFEL6EEpwbZsNPuimSi17yWXCReS/GjNQW/sPAOk
yRx74VzL2RAuvXAG+ugDwGpK4bvA0acWrJFSvrFYBpis5SP3CiT35r1eujGAuNJwDheJ7nkT4nWM
Xvxdcv88wRcn8nqFKL5ywDerQ1eB+wHjQB2eFH10FQQZNUw64Ec2IKh8a7534rVyZ/BIKTiyu12z
/lY5daUfKYE6vIN4DAG71CGHTyUaFxAPvl2tNXh5JM3eeO3odPNXx2T02TE2OQj8EeQ4XHKTCavo
x6HQWRvIxxXBHmDs2sH32SeHnTW5VJjohOwJZS5NkwUP3Mef1hV1vcJZ8BQ53Wo8CNntjD96E8tV
Bci3MkOpRAArgCwMIVAakMwFMtFJpxwAGS2eolhDEnD+QeyPcs2qnK4vkh4De8lcbueXWMFpSL9Z
+o6t6tPTF8MauW+fpoR/4fx354GNX7Kd6Rfri+f42vRIdxYw3o0Q1EMgv9L0MJsp+telGX1facjb
2rLj7NVeiwppNnTs/r4MZ+2/1OBcOE3Bk8KvYJ2YGCQDDpjt9SJMAsUrmFZGoqRJdCUtBO/KQ6xV
4BJnwq9gxqlfZOeoogd9SXx4vEyiMIPDmoTJqCMtgYT9QDxAiW9035y/H+i22kyt3Qc1D6dWCLWr
R2m+TCtQXEZDSKVUVoF/kBFL4Ct34IPSHiEf0ZfwSDArxgJ7FjMTsARM92vX0bBp9umzjjdYxF3J
8mEwhGCZClFWMbpDFRhnAWg/D20m3RMq/+EKJmw6iD8rQ18qdAp0eCEordF9d0Wrz+WffPfd9Fw+
5SJ0gVQ6F8mNBH/iSw9Blho2dek9a0UwdFGjPv4587L0tjhVyK2q4k06mOSE4VkhTFkGyWgdANm4
mpZjz78ON7aBJmi4U8HhT0NIJ/mMMaOasT+iKsau2WNJvFqIEBQ9dEA8ouDF94wjikH4Te1Zl241
S8hwv3yJphu3gRWtk09mQzhgLQQnJJ/DNPJu043QOXkMLncefaPI/yfeaS3RR//xFhiuSTjXtG8y
7RH91AgaYohepIdyfbJVsVXXD1XEzOCM283LEUId53avrjO+nqNzcSBRfmNnJ5c+OrCPa+Fxg0Cc
2A+qpCZ/kqI/cibbuGLcuGMij9ejHbolwwBy4MuipB4/lyZC4GqukeKqAm2xFHJJI0WeUQEX5wkw
MxXvZUkliqJySqHIEm+584mTQRmDc/IO4IZi/aWWHNtsblBG33nbzoSFX4IMFyoFZQp/pihL5rD6
r95ugb9l8ADKJOSEV2VT0tkwWmeHkAwsqDZ4jmBLZfy+AtP3j8QRfLiZx/daQA5o+DfSrvAL13Em
U4K4lyzPohotmH1gDPl9jsLUZHqh+W6sKrkMOLdT1jdvE1PBhWqL6yB6ohri776dwN9/UAa+RnwZ
+0IUqOBkL1QseDZjCtiuxOWep4LWA5jTcAjVR6uCnQuGNYUsmvVE4Vio24NcPmYyBhnKHOXZmP/9
To9CuSEsBxvsEMmF7xL8dtmOY5oRzH1oHB1BYm8jSi0Tz51fK0kKzDuwAWG0u+eE7aZYyvSqIcsK
qathuqfmg6DavwdcN3J0/0Hyrn2mewzM7h67Zg56JaQscXvvYiciCUczxcpPtUJYoTakXN5CM8ec
9k8td6XKDOlRv57pLkwo+VZhB9ELYeHCsc/oo3H/bYqvMRczZ6VK6ljiJMvl4um0/7NdE6HXhGuz
VsjfgfCzpnQBGvBaBuLGrKH8mPyJXyc7S/rcEd3JQV9g5BHEwy71I5XwNqhcrw2WC7VJdPNKF3xa
ZEl04UveKc2Sofwy4I7UVmaFhM3sPnfCQ3c3AjWVmm2sbdKtuEIukmUJlR9qvCKvaKO1KYA5j6uo
tgh2ywbaJ4GdZYABpalXEFDUlDYa6YfVsTTTWNRoEZBL+rqBmzV4xipytrzfHSabdu3feigL8jhN
2/U3jA5vQvjsuEtUXthM7CgnQmeStKBHLkUchFPIHGHfC7WtjmkO88jkJ1HTeC20/B7xyERC6uEU
GhOXSZMKnuoA4GgwSdbE4MYnn9Cs4wxRRj2tt5/bLoWuSP1qpU9d017PCfcCRu7v8ZPci3RMkm5K
RwZeFrb4YIH7SzaCeRjhUNyxz46zg2oZynRQu08k9F8u/xEFJk08RkUrCNuJsboMMHAaVMBilfqN
BUt7tk2z4ZTOad8mJpmMcpZ0pfdNdO64YPZoKWgFhlrIdbub3wGuJduhzdsQWEmoc1j+DtUaygRv
4vii+WI7zWF1F+z4SWaNx90gvJTsOgzBkqlRFgbeAhvE6GUhgo7BeTizgE4RCMX+r0uWfPZADRkL
49ocJesoUs38Qq1jo6leLh1ooaliENq3mJjOTOTKx353tvh+W2NU2pdVssRVlXGnpSrnV9vB5Iis
0dO2TpL2t/fbeCVrOIPqvKFRw3jUaN02aHgqU3/Z5oOp9wL6XCSWpk1cUAc07teFKCmwQxdw1/rY
5puT6/rtjrCNk5LcJbN+uy3BB3wsOcQoRFxww+XnL9XzGO4rHADGMi+ofVdbq43NEKVTi5yqB9Up
agPShRKw5cIn9LW0xCKYF2rlyFqiX0dtPUWGrjHi5EcqPnIXzZgkokGeVhteL8BLmgubptQAN6bp
N4loBTwwdCYqtsW/YhfAO2JabipUlJdFlIi0tLWFyQWH2gG4T8Xlx62Ca+7FhnHvX8WpERrniS3e
IPb3BYuZ1WRW3LWmtezBWXg+gSvPXiOvqdmXXUyLTLI2Lrc+r6UCjC5AO8NHjOoarzDGuW9YtcO0
s0EHiWMfA+Rr2uHCB6KyBdznr/Uv06J++5deWY1BFo+0iadaZaXFqmz3u1t2pO5Ge3f7R0F17hRp
Sa4jHM7N6R224wAPQhpPXHQJo6zwOPn1/InZAidLnP2gpTivYGw3lA2jC3yYE5LGx8LSmljc/oBF
R/p7sYbUfLMP3PnZPBLS6ulk2xMtVLx4XJkkyDvTZ5SqwZMFEmQNkcYa70y1/lfZn1RfdDgvnDSH
GuO18BndjGHj+6Tbjl+mRnTxqMREqgMWAGacyucL1oqxW6WZWZFeI25BSNHZlEoTReoehYY2M8Cv
eLvA7CfIi8gkvE1sdHoPrZKg9sF0yefli4MdFNUp5R7fPKeGDyRedmUiE8LrUiPsIzBXDZUDxh5B
eEYB5LndO5ZxLuAevjBHXTtyAUayLuA5PSM7C8eyVBO4l6unABoB/NqDnDsAwbMGX7363XqtNVz4
gzWywSH9JqMPAAFoIfB7Y9faf/CyyO69YjodIDASO3p79vkjWn9ZYQ7VLseHuxjw48NO3mNjv75d
10DS4+A6GAEZ7neBvmPYyGwZLqtpJN92Kd3P0XHFDOBVNKfCtfkclk00oaOKlE11SO9eeIEbt4Zn
UiJHKqKzaAXmatfH8EeJrD3v5FmXuNab9r4fcLo6wxLJKc9y4cV7BD1/HZZKnk6NNQJ8YAH34hOz
N/Rs01vGv5sltD1Z7JXvwXPA89/k5JXcf9qsUFLE7u+FMwi8B1/6RgoBaVdOCDis6rJNOkmeBVWH
ASmha7U4wroEJrwM12zFwmF0kijcKqyKIgHvNiGfXHgGCqCTQnB6yTp2E6EhknAc2HkLy+6/Bva2
yBUwfwSlmZBMHRAlJ4vc5VExQb9jEe7E4lRz3Z7XGh4TRcHmXSP2roEkLxjv2SQPgJdTIYxukDf3
rcTJDDN7xv8ZWeSjE2S6X56qIwN6cwyYvfAIb+ozeqWETPJhqnTZwfSWvL8sDAP5TNLUPZN4gyN2
IQQHMjlTz3VIuMd9NkjUuBw3tQ5iOnwzhquNp2RUUM6EhnsLprzWux3ulC7bYIUq2CV8s4Quh3+y
c6rabwVGILbN3J9SbOIVBTquH/2gLj7icKvWM+DkYHw9PAOGVTEt3g6sOrv+zQQbSUmAZddSy0sh
e9fMw1UKCIQ3JdjVdhZ65idd7fKICWRqTxolEG9vppsouoeqfZEsx/AH/C7AOaXO/t/IDqLhInay
30B8/OJ1Ocxkhg09TE+XXxDESCtSn+xIVJpxftDQJqhYHx8K+a4Dsqbf4hdTepqxjiBMxax31skd
XUQrYqMOA9B3ScMRHd+11Jnj8JoYtCggxAFKWZtcKSZWxZlyTmUI8GCVMhSNGnVj0A7wm/zn+yQt
gSaMwR9P6pmbIeu+ONGY6MAxhMSha9XxGnnbY1OEq2hK6UyACZBLKhSjfOAoqggV0cEFRbsRM2w6
TY2A5S2wITP4svh43deBZSlbFKfIoMT1tRFPVwbDIiwQx7i34hllIVjBoRTH6CPkq2/QoXxyd8rx
UuNH2REfz2SLp5fhmXfGMIFDPCtEzKXCHc8qlPIt8jR2FhTh7OuIo+6iEvXIQG7WiDU8sdr2kTi0
DWPMX8QnG045CtOy0L96XynjH0ffVE9tMT7I72FCqyYYfdvnaG1dO1qwpQ7gjipWBhhr433Er+qa
zptrUwFEzrlz8FgLDmMvH2rYWRuQlp6rm124K/c9r8eiAzkhqV8ES8AOOaI2GE3/Q87Ya7kR++NL
v9ZmhCw0F2+Uplq1rwV40DQcERmE/nrdA0I3F3JGnIAYVxF9ST0bB9QC3PCz2su/HGicAw0Zg7IF
I6y+J21K+/uKmeiZ8FnyTjRsAZwvwpuRoQlOCueHXy+/HximDaxpeXVSBSIDkHkwVM0P5I4en97s
uKjHgeiV/6kDt6m4mb69b0OGk+gezdpWZ5fakQ1038GUr8NQCJC1I9ThbNoZHZuur9wxYVVPdddU
sisn/UIaoAy/E99gHTfBwteGvrwnPTeNQeobQwlNN4SKZeSvSN9UWUMz2Ymx3+60rG/9h1LJiYPq
yDBN+YWuGOd8fxtQex5POQXHLGTnv++njrwwlsX+PaVkqa/pwKhfu5vWN/XooX7CvRfpf5Uu8Cku
DBPTtTeTYsl/7qRW70IkK4ZNlFQjqkOrU1mHAkQbl7utt7rjimIgae+zwKtcTVeLRS2EnsFZ0+Gs
HbDLjRvW12nBt8RSr3R5k246YVDOxQof5KxN4LIi1mTTpxAPh125e6+mqOtDpFbW/Kv+LCBKfcNC
EhG5XsTH/osCY/wUyHY20RjImBf9RKdFiNYXOHCfNhZIrvY9pC1Blp76b9nZwaMMvtF7syRjyT10
jn3GgoMkZlPXAmh22S7pKI9sVKyDlDlhyvu1r/CeoE2ozg+S36CCWfegQ0H3kUTZwJABk44rxqKP
penqhfsl09A05zitxak6YkSnyFfAm2u+0N0uDNEJKRsQDbT1PLx4lnTz7lvBNZEarWbMPTlzwrW7
KUNWyK5NcsJgEkHE3n5p+B+wS5ymFeVQYh4Az5klCcjZrOKxXU+BQcOsxaeLLKfnujMm/bBXSPKS
ekpB+cmc2elxqiZPYSB8VnCMux1rQnsjeHPNnj3sxkTHPCQE/CyglmfITL5hr/pmojKM2lQZVU+q
wxtiM5sw4gHMlYKUB7mXFjXZeFefe0grQOoCRQ6CMKf8wwsVnhyjWrT7ARNnqxH4X8lQnhNuzZ36
r3rx0jrDD8mO6zrORuypYRohdzjprApH6lmkpGegylSkDXnkRm/nrT72RTctgjgWdGeQTEdoc4Pn
TIw7/OBmj9x8IAMXpfcjoGXC/R2hHnG22mg7gLcQLqqzi39NTDn7ojsmCv/mseInSjN+VEo2LROI
stdo/izH/pjrsekIGXctMNtSJwW4GgEqIB/4trp3PuonD5Z4Wztuu/dCVQW0HCgi6lVWb34D97Z0
ClS+RKX0aw5AUj9Tobcm7X5Do5rMvEubtxqtMth6aTrzRkxomQSEm7UlS4emrEr5/K0+2vg0yPOH
KCyetdQGz1hO2WcrkQA55KBR3DrVTVX4CSkAEk4jYG4xhpy+rBhBP8E420azmjeK7rHRNj53DgQ0
ZCenUgDfGY1DLWXZuGQ3GKtXPyVwTivBY6hpdkTInUmRD4mbmOhHDhgnl88H5+es1spaWM7EQuOD
QNQmylRRxZInVFu45rSc4U16akZSIROfDI9Ze07kP4xBi9dmstyA2623s5MFF9/QUEYFUGp5tw8T
sJmZ1HVnlTf0sJ2sZY1KIQ4345cPCCqWPaBI8kdS4r5pwPpSUQ+/AZnXH9lw6hpVgG+CcKiD+7q6
4nXBkDItstmukVY3O/885TanLjEEFiNoZzJ4QgOdbkml08XEx714MZfqotejXkOFuIYoS8A1Q4m8
M39ctKkAfZZkuEM1/voJzviJq2OQc+Y4mDi7JksXYd5qo5mIPWgV9PJ8l5PMQfwK1s47BniXFZap
cFex5e3ZZzXWyt2DA0GbhyJ33rXeHMpuSVneAH1SCokMh9Zjrk2XmIvkSSxApaifhHVpuNFRSlOm
rsz8vQucMfh5Gudzsht6/KdbQu7YDlzK/JZ3u7AF8Efu84OXq1AMWThjdiEwvc8CILcs4zCtOo/k
OgGWq1XMo8fOO5Fo8vmYrB1wqi5kE6osWmehLPYPGdHLZH5fW0PsK0zylB6l9qXailmTPe/ypsdM
Q1nZt2eqwXz9hL2/Qfq1lex9nZl8E9ozuHp1A7wELQUWcEJbpw+PK7sicVtwtLLrWvKKFqvu03Hd
gzr1kEGMDDGVLRtJBVurue9VcBRpIOP3v2Ul/0oolCS2GRND/Ns+QbsWCDh1cdV5b34Ss8gBRZD5
Ksz5jksCwlmwIxUI+SI0X9CXSZ8uwsckom5Bw3+DNjRuv1/BAD9BS+daLB4w9sd8kT2cKuDNhkno
RKc9YY6/LYK7350oPNuRgVhyLr9tyJ2sa2r3m+T67HyoOHg0BImFzy0pmBblZogUtZ5r7ueIZCGC
IV9kYc6mjfOADxsUGcrz0PcgRehLFxm+9nDcFIJ8dwahTs9U6vUvLPyU9eLQbOmu0EdfSFISKIXr
djBFCePGUqvFOA4+NGI/mbR6m9BZMRFPmVWDZ9V9QZDNK/GNTXFU9IxQ+FN8CgUiJuX6bBLcNMur
LREacEmaDUqOTQzIwWdBB7LapJv3jcv/n3Spa34fuelXDuDdi1rZzoFQ8LHL+oy7RNLOYVbMPj/u
5kXbW4PWwZJ9uMfZKlAIkKaB2y+jM7jUyGdbfr9ovmJ4ldssG7sMQpdIlzhG+gnpTbMKUOB4pAPc
Hm/U2ZV1SVT1Cml38p13vlFAiQZv54ZNnigsF+qfkSK8KIUS9caIm/XI4JCzIHnWRe07AUVsiQ4e
xgxd3ZSoB33iNoN8RT/69TKXUd3AVn00zecc4JBw/Q0F/45Typy40DCQNgJ0xnNMFfwpfFetOP/n
ByU3q6y6olJRN37ZCRvc907jD8cH42p9pIKHZmY9nLNPd693+ahmZ6ZHI8UORJZjr/ubC/KI6XUr
hEBemFzvhu7hqnxt4hmdRa4r+uk+m3ZdtUrs5GtC5neaCSOYgNGN/zB//4zJsxu16ut4/7RyVtnS
18cgQmdNVGSkpBgdPZ/WCukImeT/ciULE6OolMnaDIr+eVhSWYcnHG8CtjDysuQU8cTWF6zqSeTS
N5zCxWZZu2QTSVqp+hKbFvCVMtRt8V2Y5riUvsq+jsQahUCmvSpXf0BuquAsCTftWDQSoYQzFGoC
csehn+T7owCIEWn0V6e2dj7FN/Q0NZtyq0L7HgcRorvc6JHyIhdaOYKlFeeUChheQecXmFNZTIMW
q5UvamvhweEMEatjyW3IyYmEboKvcUoSnadHHN1xOW7np0Pusg29t6za0lT7ECglV7hpMc2IwAgg
3+ZNx8g44Zl/zBmK/SRNYr7Z4CoTH+srV3NJSrGvMrB2OLq5TUKzutCo+GvdBbobarmzi8I8aX9S
sNUNio0Pes+B0u+HUU8/PK4Z4y9CWj3vLSJT9PO253DJJCKmNyWJUzOakOWGALmpKA4etxecw70U
Ed3xVzjVpAqqNg9xuGMxOJAdZpngisze0oHO9loVj+/b2XsSkPGWb/y36JdNC39579UXunZZXr0f
bEVTQM0f/5Tr+Kmhqki6YGzHsRSQOaTwKZsvZZT2EiT3vKPTqX+JEPBrK9qzfcWV9IBinWRsCBvB
sJ1fhw7eXTF/lWnffyynSUn9rOGbAoh5l8rOkHTxFcSS40mxk8eJi8fHexYnVUtcdmtKQilQX0i8
XG9Sm8WCqenn+KCVoc1m8DOt2Ye8LgzXGzYVaX0TiYXFv708SL6OLUJMSjHnZdFAzwL5cdg7ARdj
sLCnoQs9E/X2Z8TdWuQZHpe/7FKUPc2HEuWtmW1xW2iBaWErf3tEOdo1gFHxOI2b/SOlS7ie2kx3
cb7sNxCI8lWaC3lv+V0bYbT9CM1hZJLGfzgyKXwxBSAWsw37er4gEdmCwPduNBtmP6Qgc9UejXop
RdgKqKFn45CKiZyipgKE221FOzmh2eDhEiccxzByAmHSfeufiTdp8k7uQPike3t3hevuhcJAIP2F
i/g3wIUwZ6bxUpOfZRk2rA8ySTt86x5iijuRtsRyNxS2tPJNsM4/OTyfprA9pBX9Dp+/HvZjOM+x
ZqqcueXpd6RnxpRaRiI25rI4gP/YYLhF/eQYhkwr4104ZCGq5ZIQ8zyIH4bn1ImPcuqKJJrHT7C9
rzR5T7qGlZKvJ8YhpYw3kZFSwlP3/GgWOOyZPvbZeXiTw0OBdkNNBSd4dyzbGJWfkFccgfvxGxUs
+N/zzOB5oQ8MsTmZ+8xtE4efc/SXNIPRgvNHGO9odM1X06b/d9ucvYgANhp+P6Vq3neFBPc0VXgS
oAb5sK+/jbFoUqHDbCFhkS0i3kaGZj+BKRORnXGkYZf7pY4mNWx0E+nNDEPIXZ4tgZpidL76x6XA
K0FWv+qhdVSd4p1PiuFPBrOkuSyg9AUh5zprOwisKDWpwsA26kfhh3LnfELqnoBKA+wtCmJ0amsO
zTcobhT0Z6jn4VgQw8bGiX9Ab2kLDP4uJe/AG6C8iV9ucKpvuERFF4fSiBClKWdEcN6WFWm3mhfU
GWjJlHzjliSf8eE5RsI/5nSOSIk3VYcJETh0yjaUdLVSp6p+6WP3/zFBq57tuCeSuBqGwGTNdcyU
hS/yUxHdvXzGRh1vMNM6X2OVmbHFMYYMs/Z0gpm3FRnRH9l2cKn596GcoXIhyoyCwu27+LQJf2TR
VMnl+AhV+HbGsqsP1/IJKqa6VrcTV5RvnTaaz0xw2znIp5X8jrCYnBjV4vAC1St+nJm317vVCXPV
CvX/ZvrxqvGVnJ1K5QXtmWbf6ckBFeFo8y/iRg7jQeLtnO4DW8hDJ+1G2kiIeNlyQB55sciFrXx8
HvkaMUK5E54KnvPhC4Fu5EPX9IdrHqa8qwwmPRpO/+l/9Es0znizFhL6e7C9AmcUEimiJd5nUhes
md18TcLcdfb40ty/hN2l4HebLOEo7NP8rUQkrDUfJBD5MkuKzxle3YVsuz5TIWy2AGFujZv2uRSx
ss2cmPK0odsdg7S8GMh7iMT8LVMZkT1r/635mT5Ta1ns5GW8dolVSMIeYBzaaGh72flKzPX2agSL
uMt5bO/gkSq0+4hLLn2CRDPJPyxsbky3gYJOja4G0a/06eWs9yuJdKTWYTO1w4zLfRDKFtU+dLOB
2ZlMZ+pYrnH9obdV5NTrVZHmx0P8Ne3D0/zRpPunCtyKUm4dNyJEPpw3DAJr2cecqXfY19Uoo8Hi
G8f9g/G/p8eC0xyGczsgUBWJpEaNVmesGGBKNVtqPdgsAUOiSMF1Ue2IKeffflFOOk9xy0GH0R/T
1DJpRs7u3l7bjwqmXfi294TcmlF1JSEkpLG7vzK+L7RQqO4fdcF/ncgcBm1W4bXxT1wO+tK2s7yY
4eVAvY1wrOi+nnmTPf9DDyqcgltpPu+SG29W4AOg6hjtAv2rdcHbRnDclMwhW2ubiopxwFTrIAec
di60OsW/7b5If6rGYi+H6ZaK7+YPfsVV2GVsK+WA2NHK9/eoNxE7RgkiXwIrpAb1nOQc0Xz2zfQA
5B0v5vFb702TLVOAdOQx9IlKvXq4vNca/E//cqPmutMkwdBiHbQbzTUfBlS7t345ZIfj/+kUmnkx
MBN1Enkhg0g7GO8yeVzWE50DOp928+4y6ZCnVAMF+7/PnrocKeE8eDgfjNSGwjF2ZaijG2O/6+L8
iLOKhXXx5lvQh3OkMCwNdn7LHTh7DAJNYUdLvscJay/m8l4xB9cmricmhyfyA4YQLRI1n7UrhBt2
vd6SC4pibi/WkIKQ85atmyq85QekoALkyGUBnAQihVSx6bnbvc1aTiPQIDY/HIjXB4Uxb3Hjc9tD
C2YP8R4JqrxpeS+LefAy6/sGuW7CPo9an4K5vvRhXO1EihSSuANbWWCSkxoLLnYRMBV3Rkkstiy3
lQWz0bnAmZFB4D5TTMQ6QSskyDPvT50d/kukYgRMjaAKRJ0r6dbGteBg4fDN2+KrlDvTIsFg3F2u
ebp0hSO+eoWmd5EgdF0aRoErsA/BAuHakAzOrV4KNQp+cxvL1fIVUS3L9pWJiSo1q9coay8mPFqz
R4PX++Kf7KWhGIu1THuvDlhOEzwUb1XZt3kmrvrIANZsq7HXBxs4VZBLiehAPYvlRNrDF0u88uF9
jbTysypt+zF3CCFTqWtI6q9Ah4VByDKyLpWh3R0xvykDmKFtWip4435rNwAmegoPaI0RBlikx0GK
eUSdv/SPCDp7Et/fVE/TtAufvgGwgHhIiykMjO85gMLriECxvU0GYYhtvkFGq2cdPqzmMP3jWklH
7Z1/8Xd6CY+nvMLiJkeevweiORWW7bIQLi8GOg1JjExHfwqpLXcF1qVjqN34H+vE+UkA5mdxGZ4c
6lMSMWoSKpu04YwV7BBTFNOt7jMHXVkQg/XK8SQWa6Nlh6UfflO7A0kFPKekvF3wjq5oFMKroSFJ
Yam0voJJRTHjfUTxLjgSnolqNZdA8nzvbKQzM+MNtXaKg3qiaGOf5k7J8Rn0VBLu0Bapn1PT4JC4
I5KX0XUTGaPqF8LmUu9wgm+EBRIvCSxOmvknCrGSXI6RjcnnliDqILyfAoJPf+l04NyagcJB/QeI
vUI6Capu6Nwkr8Va68Z2ih1y0Tb+uLy9gUT+KOnit6/TuMUwfrAwX/gd/lkkuaOMePnUqyzURUqW
QaEe09gGUFJwQHReOf2g7/vUpif1KWO5C4C6JqPGyFD/ERR18XefMavVAgI2e3mPKk9lXyL3Sro7
oza0BqeF94rS2cE52jhhWwoPQ8JiLReLSNgxTCf0rYy4U1VXTYHF12SLEtv3hf3GlKB58MQAagQ0
AKgbvuVuRZktUzxDyNIAEvVMcti/gSCSvYqWoxMi3724lTH2dWE6sEJALRmYaQHGm3cVBBTLaBmr
+GyRUsQr+GLnOdqcILFI7j7NG0+ZiPg8r7mu3nYvmk/h+CDF3TzFHaLf5wYpw+BSR718ASqAtgWp
ChKEog7W6fvmmoXT7VMKQOMpmuWxaF6jNKmDK1iWLE9qyUvd5dWkAkqDqNPHJPl8FH7/eWQZiTSd
JM3PzDrFm75iC7WCJvszM0UpymVJRhWmIG824IFiYmOC60wSQifTVQhxgH6hnXSnmXuh4nKD4fSP
mXWh7vrsoDbwyqzlT5m7DR8w+LbPk2uOKXfIHPhmLm3+mJ6RsJdcx1gbQBIJfcBPSqOgXhrqQD6h
Yqtnr5TTKt+LWDaqA+JvuDO1GLfat8mEvirwMvZUxKv7G1B94gSslxCKyWmgGZz1v38tw/vGuUwq
5IrT9uoBRW3ez+HRaFb7/pI4WUn1sXZu+cTDsqWPSEfsiltral30QkxsFC4unWTFeuGI7d3X57Dm
74grhPNTnAmzS4eWM1PwTsvLSWabQOHmJQCooYu8bCpyy0a5EzqjRA1FmGY/SjlbigBchLC82KKd
5G7y+AxgTF3Qr5plhF435h3d+GG+saIqaV/CNjt+4rVLOetTyEgQlrC+jW1Ak2iIZviKnA/odvw6
zpV3RCnzNmWusMAaGtJEmaNAMXEvwEHrSqiwRlOiilvQxq683i4L+sezd8SnM37JkmNScqbAoZ/c
ArEToQVF55eKOQdy/ZjcTBeZ3eDnhYzTbWnPgiCxrcr+0wBgSh5GcJAaDmZqzRyRTe/Ddg0ObvBe
ptRGNmr5MF0Z4TGLm+13ftIHgC512AEU8+ReaLL6/gPkKW0xnYWycyZtTN1zcrFOd1ibQLgIdAho
p0K9pgZFeSqMVZhbZvUhY6uz8sW629OCQmlwRHfuZmF3qXRbbxyj3RUXpj2DpqYDkCMpBGQqt8dZ
1zzNKO2pMLfGh1ukMJkyOiV3kuHEJO0CHAbNtznirJLXGoUjIEbVFvTqeS0VN1qCrUumkSNR0Qud
xAoVYnl0MXXyVfsR5/+gw409kHArl4THD4PNArQj3lf6B5t1fsKxaNb4kHPgEwmZwRFWFl3LfKqL
elgfWiTKoTBwIrEeOOg58mWdECw5UGJ8RAD9uy8A8kx3agVbAHLMQiZYy2yoYZYyW/W3kVuaCcYJ
7oaWXcOeShMvHahkj2iPT7ZK/mNgzpkPFkJtqWHgGSAyzwcMrlm+ErEZOhO5ojoj9r+/jIi6/MBb
MnXOdD6u4YD8MB6EI69X15tLVgGuh06hGn4zDJ0oaqZ8Xc13dYF52+NXhox2c5I/r3DZMbouWaQi
dKJXGdrAtC6ZVy216T1dUJCLYx9+/5Xaf173THTObIj8ZNtsNKvoSutBmBDpvo9yz6eUAqNGyTU5
S3TpaAGpxA5rRR+VxH0VkRqBdU3iko//AnsTqCF8GXyqUunf4sIp+ZwsJAnizjC2cFmgeNxrOysJ
l8WigpFO1PsN8QUAw8nLl7rdeL8xaeYtEFlTeYTUYD33n+hDUKybQ21wIaDANx1qoMLCPBWPa4pg
aYuwHRvdkgd4zcLgF5ppDz3E3I4DxfzHZJWkZ1QvrcM3CMJ1k4KLbo/xv1YtRNNaqFC3LobDtawj
CW6NvDcjBtFR8XOjBtm6IUezF1DsO2yq/GekFUOHQmFRH8PXaTzxhg1o7n85Ed9wHOr4MftE7oCI
UqCE9Jbh/bhJ0BglTGI0tXSOe9FQEikp1cPLLPu3Ca2iiMyN2yXVl2VbEonyPgj12M0DDRldhR4K
yNgBdfDi+tpn6i9CWWdf2A2lZttqFnL0cuhxJgdclIooaH7vYMR17qfENPTGGcCMEHPlBsyurMzd
uoJHnwXXHh7QJdmwbYV9GcPF601XnU9f910kUWzFUrAptZRAbgmlnxfKXeTxvU0rA/dGo4CvX6pI
25NXVPoeX1fufvuo81klduWpZq8ywhks6Cii/O2/gsFKhRH0UzchoydZB8Uk2D7Wo18AugkSkR+B
/ZTZD1t3nULcwoSm7r2iEMyT/NSocjXa/kf5Y7GGOsA4hEWGQE3JWC49vSOI3e3JFJxLUbSA1oLg
j2tinkEJ4506ywh+m+QaFWa6VA23ECtrF4gR0uobow5Ta/hKMVuXizTRcGDIxlZLKTtQS1YkaHpm
wXC62mmfn0FK+vndW03+noH6erC0V+B5S2dR/x7gzbAmSgzz2OU1repfgYNjrifNhmYWxS3v5/Fi
IvT3QyfLOv878bq1UjouucD1tZ4siLDwO+7OREeUZz4xdkF29abjxdPwZbgUX+pmehXK2Id7LnaT
UrIKeW1EJQ9ilFOcMFlUToNoHyECSrBbYExf/cWAnXuILoJt0BLd+bYsWbzyKBp6tT3fthHK1ArT
oUmKhC1PNlNWOkdES67AVP0OJQqZB5o+N5u5TiY4Rhn9R62TVEViLixkkc0QwRH30gzxVBhi2GXO
RbRDkJpeERBjX8FLcx+CPh0zqS8srvbrC9cHg0q3poBRUmo5JIqjBTJYvZPd17To4SBi3jKiUIGI
m3PEx5ncSOVjGmRit9SdMJrZNxKDPL9uz/Zrj0bBQwzDret8Xi3PmzCCi5UZlUd7kY8D0XuACybK
zivSjHTAJwE8P4I339qlqhHa8LUOCqIWBmKwlOaexLFUg0v5bqwUU8nW8us0k21yqFWhIZLUUmbG
W0YCK4whzL2VKSlMkFXH7oeH8ibgqmwsD5bzGnT6siSEsoilesTxEDeGkdUBvin+qlQK2fhryhRi
mAnPURTz845MGCqCV6ef58HdeNSrp4GtsNXjcV4k0Jriy4gq/tJ8Yz4qgT+c5y4gSRYGQM5sJL3q
EzlfucjxL1EDjC7K2HbXEepmeeQzHv7Qx+ey/K7U6o/Oug3Soa3Rqpf5rb7UKC3MC/DqzibGLeo5
8uiqQEQ4zXNv89VgwgGoZ31qsLdc3l3xqSDKdCmaVVGeIwDu93XCwZZHIlZgOXu2DI+tbBIo8y38
X4sO0vRbyvH4hG14qWB+FYyNPISzScjtkJRd6eZ8Upf4FPbQTtLzDeRcMSehZXTFR2ELN0zOav04
8Jo9mt32vtduQjIp3tvy9kpe9KEFYPEUcQOfDhJgguykX6Gr2xfb43RsPjloWC529kYPd9dsX9ut
ePMEuddlOhwm4osZ9k+c3ItWNyjOpF7lKl3GDvaaGKP4ibMDXE+WvUsCrmJnDJI4ZFH5R5scbYWi
TZRUBR8AnFVhVKjJqsuwzzPtIqNWZKlulvafmVzP9pXkPDrQ3EYaGQDkKK9diPqP6Ge5efohJ1BZ
RBDRnE+CSPo8NyAF1Ov4Cdt5oflV5hH2SiDrgJX2k6iL0TnRNCUkre0l6O6ikuMmSJ0uVboQmFcl
oLcisqzV3pwrlwpietwMAy/TkCqndxc+o50UNqsWxDpLyiH1UuWs4b57osqwuYbLkMM1WSUSX/17
iD6LA5xFR5+z/Vfs9/HLdnS+d0K9+d+HDAC9mUngfY31uQe4TKVZuN2yqIpvyLIbEVzBES5whRaH
omhTxPOWCufBNrEIbHv+73ZizQjiRpFx//doOgoyHIzIIz8rfzsFjtZpY+ab9vNLbUtFMsdF2qZL
IrVf3cIk5iynxhW6JxVVctcVjBKfdm4+4HtxNgcIeEedJ1nrh2N0gsFErUDrZIJKfVBFvbU214gc
YGOfi1qgEzmeuG6UjruKcG624EiH/kChvDglrAXZ4kcobarxN6fCvmTihzC4oUW7y3M5VbOV21Qc
JdjVAS/XUn+y18e39gUaHSW1b0e3I8h8jQhAqDvKh4mx8SMuwLrALOeRwy4gF/PGVMv6QJkTYOlL
9yEO4mkx4K3IKYbsmuIaCaNllpUZNkF5AwOhRe8cpj3EzkYvTfaAKPYpBTZ/xxEJSxxDNNAi/dem
LNtUg/9He3JBZcJ51I4jRQW1QuN2KXmZP0EaLDxQWWYeqSAWCK+TqRRV41M+XhpMHGuLND0EgPPl
Zrew32mkXiVK+3RNwP57Kx46nJt+huOYoVU1TIxTBHsFOj/tf9muzNPRySMyT4JOBNeq/5O9jpwX
0uSbLE9rTlUjhgGlW/qzHmjFNRSncORx3HrD0a8OH99F8w0MA13R1IofM4SthaDCAk1dnIx5K5ce
sf785xDRNdwxv5bX78wklVGeWjk5f4JUeFeGtod56OjH3RBCeNWRj2bgBya/4eGORiOteWNXhX00
PuzRjJGRl7LmXT0houv6nGDP96ZyNNSHPdirHl+X/tExK0rAC/16wgxYebeC8jebQacFB6Ene/PP
earJLhV/Lau9MT63GUXtm3AiqMwbFJYPrtyZFUYXdE/kRDQefamBlqGBLru0wTxPVyvcS5zYpjtE
LHTgn+GnNFX7ERYBrJ6bs/iqOqY0Af8nIVeDXTn0rduJMhEPPYxXEhubX/oZAhuTPF5GhSqu51dY
7TO6bMNRMKooVnOc/wqBOMag2wb8mmHrCDHQTkGU39s6OZPTpHPFZvB3T0FxKodgH6uIbIom6jyj
Rc79rd9l3I/QXstO03OVifDMYcHniC1GzA4xbb/8ygGEbFKWT7E8BY37YPAWcph00XSTXnO8h85h
aXJqOYsxlrsh1BgbO1WOWjlEdVHLGbZMJNyCWNDnWYjf6LbTUjLs8+S/X27T9+XdyGAEHqH4cOPP
YAnp2dUnFosUEf2TyN3z/8OUjjOGr8kGDuWSxd/nZvIPSTgP/mTIrYvlihrk2JgdtMmWGig3kfK+
lH20DW+UdPkrHzL57FVO1674MoCuRt+xdPauINhMYszPRYs9+mZpQWZO5Scsmi6gIHEeOORfgyF/
XhT5kL76avaFnRAsgASUf/Rdq8NyujbXSnXwEXHpm6uOqV9Jmk6+N880daAwt7rsQQNTnGrD1ViF
lLdQU/RabypcmMF02RdN3+5mEUL9HMma8zSEB3V8GvJmcF8SWCnbLxPOMD4+Ov62rHnnvPCYB0pH
kK4+UmGlqKrQxLbR+iEwApozX9bNSsK5bMqmvru9GgXwd6vEMWRRwS1VfvQaIgQ6Fo8/iXzKu/fd
ffDZ2KdFeO1mB4Jd0gDadolZJuJsGX1o7RQ6hY1Lv01+APqEdPjBdaSun6bdX5FHAHncOhQwAAjb
YOZMJaje6MO5iUVWxOI+KEP4Di+U9UG1ak90QesCsepf56Au1b7OQgBL7nMWdAzb+0WwlYaeMVMS
h6Da4Daul+Z0lm9Yawg/MujW05jv+7ImH4z26spOWMY4TokcfEtTzHO1swqwdiL3z5/Bmb0B2MU7
ze9XF/iRU59pGGjMSpconMfBvb00dBTgeWHviG1sODHHzJcIS5R3lCpoVwJW6fctdIgbUdweGDwP
whi0jaNMVPv3XJX4NfQywAj38IrI7Y/tWI0FAG74kMS6zKoL6JDjRgyOxbYhmE6THGKiARKUFofQ
luhAdhDSGyILma5QLvAhDqPLLy3lAHGPQPlAkwONZ4wHzgv2iGVyhJJ+J/4OHvyxSbM2EheYviPa
lFXe2mCqPOkUYoiW7pAdysVckg2qOcXxvPOn2cSyaqkbrrr+7gySjEuou5F5Y40nk/unj8wVDEyb
3AzTwnJPLBuTF+FGjzefbsOx8PkO5k8QveAGM7R8D7W9r5GyE5O5F+VestJ2UkMS37GugED5TzFw
dmRNDxS76nBN914+dx52nb+7pNkwpVfJwLxWc0Dg9MnB0Z6wMgAYrgsyb6fL5V4PYXMLhjs57XuZ
6W+EMXSfBTd5xh2XrBy5oiDGAP4XShrICf66lVHa2VYA14oemYUWReqFteeAlupGcuZXduu5a8M6
+llaZkxDPNCnUgclr9VHq3uYyN4xPdqJBDx3RehDkbNKUXcD5LboI6R7ege+2lcjxRg5ixCbe7cF
/IMMquxhYEqQoBnITzidVIDcNjEj85hWJGatgIV4zCXU09H8CrhMhUFRM+NPvvCZ/MQeQfhp7E9a
9tokPGJdJSMXR3Aml5IjXixvG1Cc67vdRNxVqv+37/k/H1z2arjIikrI+j/4VHjGRbtERugvPrny
Crhuv8gisEDUrL6IQrcJ47YCzb5VIo2Wf+Kyz8PeK0TFpzEXTjYh0ySqvVNybaEv7A9jp9ThA+3N
jJUyfsg3doiYR+f2pJ1736AQI/aKIrgs4u4VeUJP0aS1i2BIYYTXH+VJKvQ0+XDvPfdYV9fEZLx/
68kvQBdpxEAsLC1GPsWPW1S7O602xFe6fIOW/Mn4dTnyvj8Vz/UvFzW60tCZ74Qk3BFDNTYC28Am
6kmaCAmy5freUyD3yIOQ0axL0qkZ7kW+rIVqwUrlT9vAPdLLONhBWkgkJrkLbhUZ2oBqtweAxcFi
LKCr1XP/CCN7XzkYs2IUAKuAhsUF1Arl9lJUvauj1xoXngRUlYML9RQCa26QvGep3L3egtiYIfjb
VgCEDVpMO3Nw9/Kyqf6nlqIzfNU0itTCHQg83F+hUtrCyrKBKlG3jEKOe+PK+2C/wq2B4FiDrUHt
Y9s7jH9jb3R+OpVldGRMHG80C8LOKUpC/ot8iJvhr7SCs0ksq9wUwLY9gAkk9nZA2zSnH8O71vcW
Qnse/14wHfdXVnaTXMeWmprWWTsRgZDZme+3nJFg+HkjNndBdHV0tI2Z7BBGZKkEKTM4U0y795WE
t5prFvNZTFr40mRM9UwtMk9iz9wLc7FONU/LGuhRJIKVqGXXs3SxNG4ZwnIlgOqTlhftpQysy/Wv
A1Rx/PQthZa4wKrR3t5q6L+Y7Kn0MXtSb4ee8kjhLpy1tDQYU/EkCLe2u4aI6FP+/0iG8OlJA/8H
IbVcKiV5XWt2tVhpAofo5qyWUM/exqvmCPvfvzo3xk8An13aWaWLP83eakOuDrGp29cgNlYxoQ2A
+Ess/SJolFfeuAzG72ZWudA746vH0VzM3HyL/KhMfUkcPNCZg1nX1GQgqtd3cY1Fj4GtmZR5dxG+
YVUOAk4Jy0dIXT5LlTgjuNvGtxZdi06Lejodc2pD55vqfOSf/5if3Zt0Ae1icx1/jzp2gHJyl7aM
xw5U7kA9ZHtwkbWGHtzrTG+KCrm7s0Ff02wqnVbXdp5VMYDa9EkxfWWcEsXRJaVEB0Yh8+aOEbMF
rUILOwoY3bJX8IwJ1UFfoq7U0s4qqp3EfZt7Op8Ee43zVefD6lUdySGRTvCy4U0xcSpuIxghRuGD
QShdmctZOEjHwuIlmcoSxJfkwNgdu4J6t+5I606N4PwjioJ+PZeC5m5FoIJokIuKOaxCMpsAl1rb
xWAgP2VldRCywD4DUJIsaDGhZVTraV8cY4IPFO5ySuyGDMjCMvrF6VIbs9tCPk5EUybB2KWiW0MQ
pHBrbnRPLI1LORBd8+gevUto4nyuwQk4l+yAn+pClmsB2jEQM6Gk4bGTcNqd/+fzildMw0Zmknt1
or/1yEOuC380mPD2bUhKLqsOx1jZX2016/nkh18lUwTS4JQhkefmv2XquewMftcUVskUiwW0l6j2
O7DLAczcQ79eQ0oDo8LF1u2+3W4OlRHB3Wd+b0Oe+ovWVi2bdptmQ5sMB72SRjlEq/eGQzNeIrob
LWQ4S9hjerBSj4PTtAqJow3wHRiYhTaV+3t7nGO0MZOxTj/nnDfD4Vs84MYi5m/aItQDTRqhvekf
Vd3lXJqDej5Uss+ikXYFtTL4Nl6mywNvRzXaAI5uQGOL2J8b1U+mKEhixmYuYqF03pZ1fZBBdh1t
0WSGk+k/jnImtrPoV13qv9/3vRV2i0dGLhawwLXGtxl71oGmB5vvml1d+kHsLqQtSF6N6V2MjRLw
vniVs/AMO+KMU9h/2CpqGc1yu4nn6xtfroFcIuohJdMHHTHwB27fU1TL2/BjoYr3JiKCREyRpi/a
EofrwIZPGSGxI/ZM46NEJe8eoA1tVRn20LnzsWhJDqOxyK+tlEegHQEuIKpho9kyE+mEnbfDiU4T
BeRrDJz6mrlUzlZuNmI7WM/GJADE55xqmvqsmfPIOAzpM4XfxNL7qlcm1BC6xuphV5bjJMYyYPGg
+okH7h6OHHH2AnlTyUTA0EbNWhe+7YcrOdTS9+xxGvMLaG7AykantDi0LnPYR+yOzWfye93V6bTX
W2xM3WgDaZ0G8Gl3rfruklvYb7ZYWNo+QuVKG/GO1AK2ESLUlHfdnIW0kcQqW1cUVgX7PTT+COAb
7JQKwa3u3d7g2n8vnEsROz/mp9hj86FH78DSo6REXnMC/vHIImo84zj8ANt9HUp1JN6UuEQh2AAP
dJhrERwZEGfjThYbltrKQN0mie6CQH3/PnkJ4sNqbfnDSkgTSeq3uhO28pAKCo69M8iQ2Ge+YPX9
+O3Rve1uHZDRQ4z5sVpGoXpdW81kG7ctxQ2eSIng0har2NVA7xHYf+T24LCrKrLl5f/i5XEU1BqM
6gS3sYOIwA0tO4bQCe+Cw8z/zQ107/N8FPCl7c2yEuWhdxPah3FbuweOmoStneTGzs+dZf7aqQ31
QU9einIDFIIROTVZ/Zi5/oQHQjK/rdZQD7L0aJHsc6BLIoI1AhFPD5Sb8vj5+ClUWFgbR3M3lFAX
jjnjhbz3ojEThkFjcj5ZKzar+ycOsQSGfRzVYwefaiDW2ggyAmUTVVafzhsh3jrT0IrwKz3RUhzw
whVNa/5kO43mQ89wIq+huqwBK8wG4xbHwiYWSQKzeIR/vo7Q+8mR2vRnM3nM/0tW47zQJPIeArKO
YzeSpBWQY+HlKU6/3cg8QlMhCP/o5ORpAqIJERcK2jNXHCSwOZJpnapDWtIQbTMV/YmIPu2yUQav
bjplP0GXoBHDw0noq3KrzLKMGwNoUbvCgtqMw/+8zRWq3aYZh+BhExipihFOBP3y1/31LGTSSidr
4dOLmsPwFluETHYGWXwko1RIwrdUHewMdjMbUPQ1I6hjWMrK3VqRfoK+bDWtgfXq+uzUzMlTYSAy
DSNgaZJ6N1pKvyUQncVz3AXLuBTpT+IWfmZpWqAiVvHDoIHhHFFfuj1DziCZb33mDL7Pa1j9ASCJ
rfMHfmZmw/L60uHGbn/IAoBUZYsKy3/PiNilJC46Hdly2Yj3z8Xnhmq6HDLvzsnu09oPwJp6nWFG
urR7e6MyLob/pvmgkzrSYoZ8VgcdNGKnLtlig9lmTwCUuIF2C4Ik5BmttWTI6rxIjYWIQBtLktNx
nyCf+olloTr9WazteBgLqjFHSjt1mtbIXmSoZITtrGmF6rivg4ap9V0YTNZBTHKFOljYHnZlTUbt
OCAglv3YOoajAdh5It3SLDTor4MH6HtVFRjUUOe/tzAjsfdNEwawn5NRQA7IsOGVRm9SWtDuilUM
37bi8pJ62UGldt9fz8IxJQVbdPF2RF1ehesWK2fYLW7M2jGopYVCvpHySPrWvf5fw0Q9u6gJ4OVD
K2RRb/eR8owGNfNCc1kcGJaxo6mODbmQM9hOU3/jmnqw19i/yhYmoB2G7LvA3IxVt+nLZP8+xk/z
CUN9IHTKvhy8sb/GD0C0G1ZdF8YwXeR2Qk8FNVsQRELGF4fW77DTcq9p9w+VG5FMOAWV1vfAkxgB
4facobJK8io8oeqhFbxttHwI6FiD9mk4Pq+pV9dBVe5o3+kZL/BYAkk+0n+6rOuBwcptS27czp2K
iH9L3FNO1JILNbwN9A63Rv3Yt4nSii59lX5YTxhozglbFlZoDsXQp8Xn64VBneeexXH53Mrv2MMT
WFdcorEOJJ/p1FeNtNcV/CaYxvKiz8h5gJ41FAVtysYNIzUVSr7sEBGgme7yifuYJGWn6syfOFYd
SD4mBVKnRFOBkAo/TehyldtN1BWEvMPKuYoPPAe79lM/iBOrPdgb3C+uqqHNjuVk6SQWNJa8OBNK
tRqRnZlgHhoY+nO0JcajN+zt8MH6B5SHU1QBTscQ4iSzrlHXktfxB/FULBZrolSW0WmbZrjtQpTV
cF38A4nzQ8wrZdt2IAd6GAQrOn0yfb1mVjJEtMxvGlCPsUdxLqB5EY6hlFvjcEBTdsexEvdGONcZ
uc7QY6F/hieurJczD+hzGOyRz+sUOCbcchASp4drSpNyBFIprQVPeBq64ZTvqMDEUk9M/8javjuB
0Ys5LPJmCt4X8KWkh2v7lIxvTnM5/MKTOw8T9dpWhhCGX4w2F07SzY3vAcxJ8N5au+qrLA1LkuLw
C+lg2b8g8BAvKCeOcsI4NyphEYv4rKT/HE1MuFaUpiQ3+67pXJJuu+xQRovkgt0ULIUvbxLdoZLH
o6bz6Bhtu33Ae6KeDgrZinQInFcGMkhrYqgr8zse7s+bxBJsxHaAAc9gkm6GBwsGy7ERZIb6OsLF
61dHnW9MncjCZ2M1zBpsvHrTt6Gh9DUDTIQCBInJ4kjILykcw2wd7kr0KGmVNgCGO81MK86eY21T
J1lCTJhpAmtyznU7SC4zm/LChmjqS/qJlFuGpDWj8P21KswpfXvdKvGF5o0IZWk7Ap+D3nqAXA4f
NJwFvOp3qaI3fciDocPUZDCBkdZTVOdR8t+Lf95pnOG6usV+GPO8q7Ku4SuwhCOLN/476XuFFdhE
HQacLt2RZsjZRMrMsWpDYC+IZ09NXfzTAesfDTHk7PittDwDWeZID41q5pJZ7jOrtVPZHygjXLef
ZWb49pVOKInnZS8Mg4T0y+tJaif8yyc1p2+y4+W5e3hNASzISPnFDXH60iKdx0UNERKCz8NzUnrT
HveBAb8wD/36GbNQxB+IVd1bb0NdgWzWB6mgenHwHJmSUSRpwWvDFexEJeDnsA8sLCtwj51RT+9r
R4W+ZnmlIY3x8OIgUl5FVwZVQy7UiEsXRoYCMBjHtqv4U9KfsBKsAoEVsp0B2uxF47E7jyn2QwP1
r8dwMaqcASXgfC7j8rluCduh5EARkhBU/D+d7/hxuMc4IX5bdwEvyS6n18CcJwxZT0pdTJgciYYe
FbAQxhv8Fh/93RKU5lnJ0vpwi/fCu4WIss2H3dYfZjWZEOOGV3a5u2Acol1HR/YBKz2v2ZhrzUh/
wod6nu7kPmgJMteS7TAowWvtj4KpNXKdU8WSxj9DirCKMoc2S7VDWQ7WJc8qEwBs7TO0DmtkqlMY
a9hCVUR6E/6Uom1LxcN16cND39trpIx0Lha8u3sQnmlJ3nU31q1WI+LEJesUuP4FeJ6B7ASlr+qs
jOCXfrlArkC9dTupNP7YhZhpEOxOCTr2Dan1SA2I4JHeNpR08pYqx3A/q/bDDdi7DkRqWZJMXrfq
Rb2DAMdW/11w3RC4jpqmgRga002GOKTD/PiqunERAT0CxEBKxdr7SZpHnRYmu26d6nfv+wrGzoAw
pMsMhOeuG7uN8temAyv2P6SUHwMDBO4QjWsJvopBXJXjgNuQtTbupnk2iYfpNb6s3uf2oVFpfemv
olDAj1XbrkM3EO58DQrQpwNBpgo/K/ak6yiOHtWs4ijs2WJ5B1ckp1pnSi0YvH84nJwFKQZHjH6W
/QCBiOF75RbT8Dk7B+I1Vioc3n25jMssve5wBelb2I3MNPWHzf1TXszW83qnXVqH/emLy1QJmh2C
PZ9yCeVDqhfg3RV8u4AHadot+itWOk6dovhE+bg5v0QNzxxBaGLymOJdAKhEpHKl4K45KrqsAIzb
Eb5cc7aue08JzVAg0AVw4yVyVDuC6RBhFVr/99AAWvwoKAouY74Hi+MFh6CtEW6ISyDyDh3iuy2T
DbkXR6Bcq8wbbDDerkLQOXyQ+3rsc44LK0+j18EVt6xf2T6OLWa7Csl4rPqP13AmVqEeO1LqHpk5
sZ8pQSdHk5mHf5nfq+UpbKtcIgenZ37n4mPZjoeaWyG7aeC1vbFYkzatJN627XxT7PTXkQO/YJUO
2Dd6EySJOWvSWo2LtDcuf3vXNuiPyb2Y1EU4cKlgggxYAVM7LHukX7NJhFMBPY1cbbnBa7aaOMOR
rU2XmRHmUwR4n5SvZpsRE5czMPLXsrDuZV8rngsjmDOezaTj6NJvMS79/KR9aDqgQ2Bnl8dhEDCe
q3gAL2v64YjAwOpOF2ytFrnSEfrKqkgckpLTrr3wi6lWqwn1/QY4LIs+WPOHXqVlhpCq7djVh/P2
u00qHma7ZPNnWtW0zXcDikJkQKwoL/omAN6AlmwR8eNGkBBPjfpAOY1S3jI9JAFo1SRMvL0rv2hk
1I9t0kZ41xYkMsxnfDCljV4OozGoEgZYokQ9C/aEZm1bwMyvXYotpGzQmY7+CPrEUZCd2PWtooaL
NP+SRAdSjY0qOpi7QzWBrxVm30X7iYKhpQSo13YwVrMNZ3VUsQL7Hsrm3Q8+tL8mtrrzrZNy6jMf
FRRqEXCpIOnmZxU5h/bR32U+E9BnG/JTE50LUmjpsf0mlNV1pVbnwIKB9UMY3XgVyX5K/5lYBN3P
1y8scPissIMxSoOmp75MzMi4HiVdkLFT1n2Im235uTUfXTKWuatFB1bKfvJxO+PseTXoQ2+M119a
AScuII7nvOngtx11bEBLnOEA4RDAXX4d+7RlJlmOecFYy6HKyrwqan7nNAAcvwaSVgXQJRXGizLR
wo6MM7+5iaKPeWceqFNpeOrT3YTviyP7YHvS0dXEg+YZoKHY7ZlAMJyTGmqElqhuIcVZCk+0gxRa
CICk6mNA7kLmMvHlzgehmnZ7sR3MkLQWoBd7Ujx2cQqDelp7JRzaz2FhVSRcCbpMaDcGfS61hl4T
QhHWzk4Y7DUp28lphix5UCkyaAMsJhKBN+yEOr1WuNgV568wSKLCL81lWFx8sSrEJZuOL6W74EuX
vnWaRFz2GLP6UVdk803mMgmWn5myto9Yy4qDujr3cexuIJf+IjZkYjFhWOKJG4ZuHEuq/aMcZBGT
FiABpVTz0pwQ6vBMXPbSsFBo+QgKBW0Kv1+7KuRwqi8b0CqwS0nM9QwY72XqM4ggm4+WL//cIRRv
X/5AE9g0ZzxyQwkDzFCh9gbt8oel6ZmqO385Efyc+hkX/zabjWoFsR2i2L3DKQhjh4kn92YbQMy8
KV2Uqy17EVXdlAlHALMAuwVZ3pyyl9gPJhzsvdT4pUaJIcodcvYmvwVnmCiEY76HrptjQ3OFv6pV
LtUS9bPirqsYuO6XaEsw3/mE3NINwzoxzXH7QV/Yq/zAsu1smD6opv3d5k41Ir12YgdjHWmtDozF
bT5auwXxmYvMKUY14eUvIK2CMst3HJ2+D2/iy9Z/tm1mP714+eEkHHHY+DAjoyK9FIGiWM9rQtD9
iUAXwye077OUaP2KJyc+SW5LU6SxPUar9A4B/L/TjhHDNpVHLmkSplCo8mcLlGw4nN30ZzBpcGyi
x6c52AHIlSvj43i1BYlhYONz3p8If0U2Vm3fpeFpCHotw1R15QkpLl5sqeUKM7J7Z0AwXJMCc848
uwjA8gUPpYuhGmJ/q1JNLKwb/9glqgSXZnyDI99qshxRj4QrJsP7druA2gDzKu8CR10YSC4kUYlu
nKfu47rPfoY/8wIBsNY3nR4IDtoSjVwtWHm5p1kZt6tLpV2h1mCcLwM3BidTL78sQfX2jcUprTKg
bl18XnpblcRy0eXPlCAadlG5l+mcji25pH5Fc+x/u1413M3LqGzI5hC/TECCmp8T8U+oMSPtEBbh
HTqE+IATbl/T9P52kbnhdx+pRD8qzrlw46Zq9lBsmHFMBy0gjmhoua4L7xQbEoYHlPGu2uRnIo5a
1wTq63H1HgALGG4zQD2z3oPnPBl0oLdWWUAIegwcd3fpftofVkkv5zExPKcTxr/FpaypNd+XYqoB
7bOQS36J0Kej0ZD3dvpgiTU+oTjBell+jWpZjZJ9NmaUb/xjLxApLD2TIjoiVAIan1+O6l2UACTx
IKcHRMyNLORdRpqUYriCSMGxXWn3n4+KQTipz5lZpHq1ihXE/1tJrwjrNUbGOdz8pRaFZr0maf8g
ZUBj8r+HAybXQoSKmOVgKEEElIvsThjBsKJbooxm8KbdgDNCzXZSzOD7IWoKWVnipR4lkiBpw6hv
MGdUzomRaU0Y+5IxYCNGo/9FU+3ZmbM1Hr3w8BNQVjFHC2BnUpAObvNF1hJMCVDaKNInYiOZ0cOh
yl7dt0CRjSNJfYHo1nMq0fdotXDXKeu6hKQYMrDg3O+5J/FVma9hHfHGL9PP01QH/rjONEwH6qS1
PKTApetqjjPta0KsbTYb4wEAgQDNfsCfi9Vm15iNyK6Fpn6QPEeoFMMpfdje6lvW2YAUnVemBPVW
ED9uBw2omJ0VGtv2/eUQJdZ/M3L7bjtqxequ4+37rI4GaCHc+o0/z8l9Cyl5A3G/uz0IeF+I8IRR
v7IUtAJSOgFC0b4IvF5wAGXWMtmLUndQrI2swnsF9F8/3Apf1hiQ8vXhEcK/PcVhlfFORwAzpVfi
Wl+k5VLsySUJBCuMjhfMeJ/yp/kkdxMw5jt+e28BJuHyY2W1S0cNd7FOG4VySCaLrRiW+G0aZv6a
Nan4LcFudWM4oLfemIdI5CEl0g2oaxLqfEDaW9A44qWd6smGhedvkQUxKao0X7G6ty7gyPRM6qkR
H4zbLYN6ON+lRwWsSOK61W6MCQUmqhI8uk9Vlg6fLnt/sEOEkaLT7v56tW2xQMo3Ats0kfhQIya9
N68NUxrquGXNtaI1TtV9PyGQ9B28dVCHvzojNLEqQnenV46S3D3fqo35lxGtLq0RDb4irCozdmDg
kiwd7B6xL71VISorV3BvG6SWioosTeDqnMKaA/wEIKgZdV4XEExCMwAhtXB1qI7HXBvYj2uFB6Mj
lSFMj+FAqfP8eF0bgcrvRkkN5K/33sKU3Rka6ulzg+Q5hWxbPUtvfUao6Nn8/dLCv+91OtEVET/I
vvbRUqqHNI5MPcsiEHrNt4a67f+YRVrhkTBfOeLJnyzlBlfGeHr23YYsJGVPRDYsNawFAlsDpCNd
15SoBEB8mE9vsFSwU6tNODKbUYDQEcGIX5GMm1jKQiYV9HL9Uvce8kMk/OkVLISuT1ZySFvfoUSl
bbwTQZ4vLPlqqx9JuQIdIX3SXUy5f78uu6qpuF1GCXVewx7GeD286hBMVtTU5+cJtplR9IzQ/Dp+
Atg/ug4TVFqR18mWtegLzMSwZdUMKyWWYjwKgoU/+OdC/f6/2SsG43BqR+cDko9cqTkpy9DkjWc8
xDE+SD+C+wgWb70wfJ+3HWS8H0x5o4GnGQ65SW32iVxXu0ODJnkRffuzQNgofs6S/907tCEmUJWC
mUVBoDu4lPj4DbmxEE1QBOt2cWWQT4TsXTPxEnQnBaA9dE4Bk6GV/fmbOwtiHp4FJ4HJoRDQPaGi
flhIj1OAm5BR5E6npke9EbOK6hgGJrmXF1d+nV8YySnI8SC/PV3VJM3p2wqwlThNK7ZMzWmdiNop
jG8MoYhHHjVp3VEV+Gtz4gS/bHrqKjXQH776HRA22GXI6mtZYOl+4phmYeR+AyxzL1tkXOlB/4Kh
XiJFAwzf5LaEGxIiePNtt32q2QQzo0+Krm79rnRq/MGlXmE1EE75tcvh0N7WMu/VGdAoI4iyqccZ
B/Qq2R443Fu4JvwzEqx9C0XicknNvs51gPZ+GqBpxcCnQO5L55c8jkE9SU25/Vzthd3Ksd8huCN0
pGagwN/5mw+o74zenaO2WkSx6S49HvzZNYpnRFxNJESR1ivfKEZvcQ1TczwTRWxSjw5HGmm5VK6d
09Js5KgRLnhe+A0WS7HtzCe0gYdI5nTJPku2pEwBllWhdsKP/NPo3jZ3jCNDNNs/f1VtL4RvYc4C
5FveOGQ13V4BdHrb6E4FXv5oA47nImDNOSOTzMblBmH0x+Wum+QsPkX8OQJyDkknokOqgL1Nku2q
gTeEi2KBsMmIeljqRxRiAyG23+M7oGZd/S71pcVk+3MO0X4t21mWTJrq2SMVd1qNHSO5qXE0doyo
hXzOmqhFD5hJmvIc4GHwuENeZnGtCEXknLftPptSZyLc/TyGISJ7kWGiBWDsyE+AceTxLspucuAd
wmCzNw223dywxfc8kMqwecN8roO8JgDbpA3aoYLYmfLJawgPUjt3BtQrtt1i4PCEEjEnoOoAqx09
5jXwJ8LYaH5nHWR9j6QbsZWA7bMTeE3RDNv+2bgF8+rcQN/T4W/oGgctQ78mv0uyZ/GQl8YQIN1j
5ZutRw27CIO3O9I6FtImCLN9vUV1fw8WiwzUd3voYKavgp5gN6cB7aDeZj9XwhiFClUAwl6va85I
6h/h7F4XUE+lHiJn6NUMxszhFXkg8khuDxPSZhkrKvziUISzuKxVeeecOguUPm14LD6chsYcT+/L
hpH/WR9vxiRwMoX72euOcY7QznrlNTMZt4jIwmpXbXV2/om4tspVmsh7KiSG4HeqSQ8xPu8qpTtI
uMOQ3Oy7V+luArxaNLRvMwpxAbMm761ACWqNhDrsBEW3Dzgfd5zXCzNhEFn0fXDeQNSFa+N3QAbR
dz6FWKSbG/2EOxGT1cvJ9KgYCLxCvgw0oa7BE9Gm2xcMZgoAnfmr/T6IYUe7flOpZ3RHowUDNuOD
Avlg8X/HqiEiBYPeYKRkgYRsHedafvT1W/qHaQ+rF2yREgYTz59aJsceAzEP/sXg7pJ7j6qNTwWU
/D9KHXTx40qAd82Sfygp0TTdchoKCpGe8p3QlfUPfdl3tU4U3OwFw4sP0theYig0KNPFB8951ny3
iws/kIIKSROrSK4kZhgQbMX7G8UE1agIlFoIYR3zAaKMr2VaYbydlRtT3dddihBAO4g5kQIgX6YH
bbdsz7BywuJo4sUF1K3FdiXKKPJEF6fXppQyD7mgPYM/7gI4K/fH6p4y93UdCBqmJ3i0AAU3YeSh
QUxViDMnYclNLi3OENv9xCd6f6dfJ+jSV9KIo2u+jcMz2m49NSZRvJMwd4tQ8ypei23Hxv4a5sGv
AbFfEfl3Qyg9IFAqohWwaskEJO5e9aaDpFZwAyxgoprK8vbgY0vmf4b4C+PHGcJt+jm8gw5P1X87
AvnEkzkCDvruj1gILHHsjb60rOctPheyUOC2er0f+6/ARczmQi8tCZyxmgxF+FTxmRfyCCGnou9w
Cth5vWRKk2PzaCAGu144o3HkJLgg8IpEUqAkqrSQDaQsLqq6MeVNjCGxrKEWTG7jqJUJqDJ3DlR6
nAeJUbrqst4AxprPGmAEqIYX+u2DCny2mV+iXMpBHeBFVulZ7c/NT0gljOGKR7WcvuSURBWE9DHP
SpLw22WXA57pv2uREUxnQjvV+G5HO/lLhN8nb95KOxBKp20+ohl4BROi4f5I0D79TWOPXeHRcb8y
pFmYxSdtURzRd3BrqtH1xqEJAWY/UHcs0JBX9sVjrryt50P2Ijs8o2GUJ9+icA/o21kRNuKq+6Ws
4Ciez8Uplb3sieOVBNY6BVmpJC3vA1RmTN5n0GMUM1kwNyh8RdNtRDKnvPQkLrXNh9lX739w8zYL
/eXzHGrh882LGSqKiy0t/HjkrBaJlwh6NEiOifi0PMLlrP2NaFemTyt0tXqFAgippkles7nT2LRV
rbZI/BXgYLG4Vv3bE4324F6K+rS+QWlZjx5ShBa6DhaST5xoaT5mPXy4UH2mQHYaAS+TKEaYPmKa
CEL9/Ew5StztCOQOFd36cnG3Y+egNZNtraJWqwxI4AIDkZn/qrPY1ihL2TaLF6qLpmpO5SFx2/Da
ApOb5i4kbKTH6pboqVKLVrKtwgvUMpZW21qVKYDDZqaDZiLg9lDJdDcOw7+5a7anV4VKRUAWHOMK
9EzQMqcCtv4/h+zyIudO8iKYYKTDNSEnPgZlUQbjJHwy9tZskQ6dDX9igsHTr6ERNVERJL+C9iQM
cCf2qXzMPC4FHwwcAeegzGMxKe3UU+HHXIaUraqz/7fbi2+B20T2cLc7BwaZ2+9uq5VWu0ji189J
HGvcB6qUzrit364fsIhE5BVcnp2dC4bnvdcFBamn7NQdMk3cnuH3aTJqdZhP6zWA0xRZUoy36Joo
zEnePWkv2NTWDxnldnwbmuwaK37g3O0GWlhtBHM3zgNdqxNrAl/y5Hc434EQ42NHAEexfrMJ0gIP
EnTMP5SKk26puoRrDPQVUDTYRQ5ABEBRqc4szEJ4ekUZkm4FQVvg9EWC1AFMl/DjNOhqBKzNq3Jg
V+dmplCuvDZR0sAhRZSQ6RaFiKyD5zOM6k6QpVtakHDAZE9etd4smnIfp57Qs7I6j2YwVuJl8IBf
3KYuK4WofIfKwKvUcxSM4XJLYCT3jIOMKze7Z2Yf6U5DtcBURqrvi27nA+dIA4dc3rYvO2z631BG
KimNJuN8k9GIRCgSHXIK06We5gBz+rCMk8CD81Vz9BWTxgElnXyvzAnDe8XJL58sLAKgluh0T+X+
akCsS10NAFsUOLdDMobmDb/pfZYJntUgNdaVV0vDSo1o2NEUQYevq+ixBVMqgejFk/yBjttHvOo3
492olsXjoUT5e1h1B+GMNj5W+QFFAQD/eXT/xyQB+ZuLzMPBWY+pBalkHXxFRKVjcGFwnCbtmA2k
jNnDR1/LQr0sYTIlLazLKRjT3NICLdWodvZuakB+FVReOSJk7sJAUbMPbqgEglyWPQZNwBeM++gR
dyGxjm+ksAULmnpoDAF5bAZ+fTTaVD3jlCiJYtqNhMV2ilr3w5FIGpWHDEoaWXltbOMvWHcrVBEE
pan5pGqjSYRr5d4sAC1my6YEFb3+Klap3SsglQUzsj87pkc6vkynluceiBTnpdLxIyO0CTdPHUNG
K9iejuytHbVN30XpngntFXjlmJUHFDmZlDfvyDoHNzrTUW+3MrAMptzsDPIIt5qspnYw2QDcm1Wx
mHcbXs+qXDweCrLcfEsv7xIn/wn+K63LLKRslYLzWPMYRDxfi2r5IIrtvzCX2VptjydyVlXQT9Nx
Li+WVHIW3KF+PsfsVA3I6gURMZLTOREi+v1JItC2NSLkZy/qX3PSBJHlbF/Aubf2Ihr1HR1QrHqB
x0nBLnZ83nTDt/IpPVCY3Bsw661L1lFuPYnKZCADWUThk/9QyOxatvX8Lpc91W3ewEf//6208t+B
qfk5nKbFVDJFqf1oMSu4YWCCQGmhNzF2N3T1GVuK4e/blLkZE/xHofrpDkRM9aqE4CCjXLTrS6+i
2s7I9m30Irv1ec2p5vUdZdMXr61bENj6Iy5KYb+CW+6UE4Hzfa/HX7NgZNgxYgqtVHKBsYY46UKj
ZU1tmeYRvU4aPIOv1RBxf1pPfEfD14JvZVKSe7dGB+nJ94NRjuGVIpNy1qJ0Rik21s4QRJpgzHmi
Ce4xhZfuzh9d6L3VqOB9C95iQbO2r0Lr1xmh/IpHRgxcjZ4HDHEJTF+gTa4N2h4gMvBKv8bqqxlc
zrcBln9zZ8cn6noF7uZe+5Mzw6QfkPcHlAs8FgFkYdzlckB4oSHiUfOm7T6v3Zorvd2jStgCTbpu
/Wl0Hm0eEtENpvI6jaE0MATNk1d5bkfgZjgbpT+xo3bWaQLC9+U6O1PFDtPIof1HY4Snmv8UaUvx
YrU2/M3MxOxruz8PISLePZcMLYzxeYFZ3jlQ8EPpQGgc24Tl/X67m4i7snrM8YgZbuBGJ8+Jr37b
Ir22LYJrKx2XvGnFFGN30lAX7oMExBS0Y4AUm6mFRyQzBZJMHuwgwj0KPAICHMR4g8G1nXIwN2D9
ucb0EbzuFU25XrvA82nrEBMXIa4F7bqrUN26rt9keUIPFsho7sLWcHZmv3lcm1PBhdemLSTMncgN
/mW+5n5M2gIlqFrFdZiXTvmIZC0Byl5IwkZbGEIYw+C/auxq5zt63/kzAah4w2rJeEVFpFlQDd6f
mpm+BfQkAdHYBsDW3kPhAd+DrcMms0YOSprGbNPku7w4UNm7WQAK8oskRk9F1uE1MrzNjCO01AIQ
wkMeMPq67jjkRwNG1ih+ArPfiz9+5MVCzLZzoRp1tU9aybwgdxJOJomIpahYJ5qdSkTirqEmuaTD
fvuOEMWV02goWJMsdXfjCrN/kbNGmd90yjl6lKNxpKkKNdFgb+Fa+OjsZMsmxkVh92hNtSGI4mwJ
kTIFZrFoiRuhyi9QoU7tsfWHy8UPhPxUlbSOIY+GvBQ/ONtYUu2t/JpU2q8NT3CJM/wwNHzWGzTb
KosxHEJDhVx2tZnjkLlnx8zW+FjjMtnahQ==
`protect end_protected
