`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
p8A8b09Ra0o1o1KBqnstYxn3Wxme5JrWvR0+B3bRTycm87GwR0cQSCmwGgaNHYhcqK8MENCyANAP
9de+O/RI/g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hHlcX7YOsoX57YsohrVUVPvRPUUS+AObuTWv/MS6aIrwW8e3k2bbkBh10qkAlXOxiZ0o1jf16hCC
F8080L1d2hdwEXf/C7Radh4xEw9hKkYZtzK9SUQiIH7XpIQI/z/cggbx1xvUaiuZ41cmhYtJcHQP
g511bYFnhhuhHrFVBjI=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DnamHuxmY0qTmWsmxojooz1TTTsfuLef1uX6jDyUSFysvlV9VQNpQ3xYg5QgqwM9nt6wgRjDCncR
zg38n5e1dc8l3DJfYjoxthd1emWfCXNIDZOf1q0Q+180ymUTXjtijRD7Kv93WSihuecylMGuqqyV
YLlGG1EYUPkFDFldrwFockL2c/MOWI5MO7298cte7f3xYx2fHDFMLoGv1WqKlfUKTMvodsxljrPP
jUQWeis/TlsqWW4ERkcuX0LDyc9EZGSdk1MVuftNzZGndMAneK55nJjBR4vKuS0wNfFsprGdysge
AvZP155o933YHV3tFlnQYFsJPwqbHKbAdEf6sA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
2UHg6YmJcyzM/mdtPgeb3g9MbF3T/oPPltbSXo0rbrNLXEOauGM5IGyAHKL2JV6ZNrsaMgLxMqn4
nptShxuBGV0V2jQrXtVGGopPqBBEJoz5Oq0pnmAIUoYko5yGS/hdRX5Dx6WFHDX9kdPk0j/OYTel
fNfCQj8MMkn0vr4lpY8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
PBYcqLJZ2g51jHpz7H7EHcP9A7s3UvicMGjCmsKazeZLfNmO40rFpVjaiBjHUlu566E9sHy1IkNm
hKtC54tNVI5ZpzqCyyxZ250vWugB8TPvc2zNLxmBzUp7eb3fUJcH/Akc+rcnvB4BD08YjFIoOiCC
NKjwtv+ev/UHZ3LNRpo9UhDJoAmTCnQLNnVCwqS4JOfV++QciIpzp2kQAxXjBsWIcp3FdfRz/MUy
9YO+OpflOqBr4XZGVxtJlwGqRoC0DzaixrFBmCxdxUW5qD7Raqlzyhw3i2vEl6Xa8PYQbRY+VOY+
s3myYWlI5bCRvDRuFU8FIij8hnwslsK5yTbsKA==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
E+LzsRu8E46Ob5yD44bBcg8CkEaYZF2uIqYOTOdvPDdYuFGaCJryCUQK5gy9JjKqjExq1u1VfMWK
88sDiz26jyftK4sOWuM6GGTXFZDxAnPKab9BsCcLNUkymfQgKo07H97bC/iZl6SCxH6pwtK6oGTs
PHxRBRokVghpHoKv69saziKFaW+6FsRvlpVKZl3BSAJAcqCoNorRAqOlLPswrHQXDj0AFO5A96ig
onNQVsUoAFAXwP80bJWHYP9kGhvnRvA2FI5sfPA41+lAoQIYHZmevTMbiURBBA6hMDprmENsSW1C
VDN2OilXO4q1OipnCjNhuLoi8Xa/1aZ+ob5u/g==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12640)
`protect data_block
ojoeTBXwI5NuUed+LNpw317gVUoqOPvIG58oGWkxTW6p4z03G/50SrR2gMDS+7QIj9hrE0Pxq2s3
YSyujdQqapvudTWpCvGoBGbKkkTtcLMlE2sSTxcEoWhxp2QFB4VjAzFPGETaszIki59SILnJqnIc
MWbJzc9PWG4PJwh9fUlmwkYvRCewcNxJLSlQAMWDOOjFbMqirvoyGabCRgZ3KbXFWDoFnj//hDg4
LY7rfSA54WEuMvjvjcYVZvv5wlDgukreDDgBBzEkbZ+LfV8xo1mHSjNFU5CTPv2PT2sSYKyn+nQP
yqa0A2G35ASqzkBJU5rTv7z2M2k9i86vgZ28VB6ZbgxYR7hnfRU4+zy6fciO7wl7LduelaclH6DN
hFKHvRGp3tws1zWUpdxca+Qg64XLnUI3ceRpTDC2aGoyfOOV5DbnsbEB3L7PpXA9xmAKNU6J2YIQ
xSyGDo+2XBqqJUR3KKZGyx/hUBsLDvKIFqP784eJ7ALc2orw0HrMxkOlj6Hc7wtioU15SYYWxDq9
lN9jYOLoZJokAS2+9NGlxnA04FlT5eBW/Xws7Lhs18m5IlgPPc5yCTVnAlpz1i3MWvTEiMR8avov
pxg2ChbO/ukULaSGAWm7SnwxA/fnCBSW0MyyMaQD4JQ9nPkG1ZC5WSDEQpv0R5uMo8QjWXbfTtK3
3PrKnyukdl/lmobwMnrl46fWjXVykkvpAh3QzHPkSZfAyHbDbop0wajGgad8Lo1WttdS0ktx++Vn
unlS2130FbHLccYYD1ccBGSM1v5OswoaAddPv0THFJJeD7TM15GMDqD1KDSz2EDq+I6LDtX/4jL9
6lkf1WllQT5JF+2y7mKieUe3hoOAh7vuTR2jf+330szECY2xZgxudZe7+mxMwLqIaK90YaHQCkIF
stfB9lLHFG25Medlx6GaDZOvIsmHyKG6WvUjAoOga5fSxGHFBseCK82nbz1jdsQSruf1YJnhqDX2
0CkXSuLS9WE53rqH34XzJQP/trOLVUvPL4it/erLOAGb6hqjvl0hCIPRmLT3mSPZenDg1EyH5RyY
+6osGhoyBAewyNvvFLzlEDah49d0GRigjG/bHd0fVqknohShv6V46QraHQ5/wMWLusO8JHQ3B6E+
4qIllvBqZI1GCv/tq2SuhdIoukH5YHzoPYDRVPBi8SogFZ4ThQ/6IyF+f4c1NOeEYvfu6OjdGsGm
2FX8vKNQOk+jAzZaWsqzKaFXsoIfZois2upuUXZhbWDL5RfJdc9tZJCndfDqG18L5JHdiGbv5Hlu
5U8T54HvSOmC54gkiu7RnyYfcFKQzzmm+6Q+fucE1WgIvgxeyOs4juwLx1xIPf2p8o8LDejpNtQC
QrEfq/smk0nenkIbMkYxBQrwkP8O9NlmdlICNeyWFz5lFXMu3T0SiMUxSbGCMmtV6gIryHaAxYmg
WODW/f8ext8ttfIJbvi2+OlNtwtZyHIlQp64xCzdd0paiadRsEjWsRSSdxSViS/jAZdtzxLBTIs2
Yfwp36HsvEogTdud66sTGqvs6vRfhJxO2paW3yHwvKgAoEx3CUlYqAQ9BqJF3/ehpJ9BfVVQq674
YerxzdSkNGH9tqWR1EfO9gItjt5PrNwKfyKgtPLnNqT8wiKmX+o203xRa2lNt+DjEd7g7FtaW6Rk
fpkhrLDEIqjqXRA32BVoPIRxSPMuSqRsK6eaLh7XCAyuYB2z6XURmT9yKdtocWqLOZRbqJuGRuam
T84kV/JugwyuGaZ1lIIvC9P5JEllCbSckZ7clI/VhqmLsYfqAmJLeXMeVMbmnZM6h8oFcLzJu5x2
s3wkiWeHzmbhNMEFzptntxPpiR7g1GwmAZtTYpget3wA3avjXfdz/pGJmUBOCn+tO15vEZEAX8PI
TAi+dzWU2N+aiaD02T50hqdTUtkgALDd7GcuvR3dDFH7G/tQGTfAggh3YZ2Mf+6Wx3fMRW302/T9
M/H3c5JZ8nygZBWbeCfUIaZOgBre60T9CjeH6SsF2o+owVa+nZ1fT5FMa0240NUTfiabSZO3sNoc
700Xn+++Q0CRGZZkv7jnWf7Rno/1lzoC+m1hdWd3IsBx7YK1XmsPFpidX1gnIStvgDpVC1p0y0Xh
GwWvnojeR05SOPcJzW90m7NQp9mkV+OfFr986ys+U+QCD6zUGEOUxjRgI8oYOCXFREOkASM0fUlm
QAF8HZFj142tVinwrjR4QJ6GGEferKnYswsPuKS7gGhPaIeg6lmS1PKllyBWTKCllPAOLMkMdxVf
YFLGOkwR3WEaiDJPNJjUv/1oDoBm4YAaAGR9swyGB1GzAQ4JjqBuxoRcPaqVr29/ukmDTlaTLIA+
xRREdgrpZFvYUGruagKJKgx/j3koUG2FYESa4YklXeyF9kobUGk3wZJcMhsXBBBKdpFoLXaH5h29
4+z+Gqh7z9M5zpzlGNkP6pk0X+noiOcLsbLmZfd5dKb1l+Oi7BMRLdts0ARB486GIjNbvPNVrBH/
3n6VoOHXDSIJddxEADRZ0cQCBOd2uVXAGKZSDa0b2WAlHGn/LCL3HFOfhymV0hZjxQe3WUf+dm38
uvW7IaofTRnsCeGL80rq/b4k86LedgCOPyO4Bqs69yJ5nlct4PELFn4ePUYvtw3JIyR5ETTKjbgL
k9QeVg2KyPsnZ/cMKmfmNKXaHAKIbHb61171QUzodv7h1UzJ8YGPvZM712Mjwin5ZeMrNNqlj7ui
CwvtHUgRd7HZDuHGt/snWe5fKPfu1l3R4tpwSUsPzzqj1iLhLCp8lgc9h0ONz8Svk+qHK4aWT8cU
sdrLxWwniYMXH7e79rijCH92rIOHes28I0bRUQH+Of9UipoqnM2EI2THBt+X2BZwOoxe7JjPTQNx
lwS2UtXi7hpPaA9iYB3nCOtyFgelklzaHCAmTePq5lpaFPJwufD0JPaHPnjGH2mXaqmqcPZcEgw3
x8lBu5JvJjpXDmSVLi2kuL1iuPclAp5nnnDryRE0RBkL5yQQsZvRJS+SKujsl1weG+GSPwx6D9BB
r6C0L+Bfnqaj9BLSu8zfNXN4udzpJfUy3I/D6LFyro7K8nU+sNULCZbGnfL+jGDur4wFOC/audR9
+168gF4f9qytU7O5/Szlm4mFUhvC55yOEEn4I6sbJeF6fhmoqW2E0qUaEqQimkDO6uZciouMIlvL
q8kAZCAF2Fsg/BrecNOSlWkJbuzurYcZh2Ykig9TCU5Bre2X9u42tG8XDWjuoFYfXhgV/PGlvs8X
UqFLIr8rZqqebNUUi7sK1Na28Vf1jqGsJxn6J7Z5cilgKVozNv5yNh2oJnNx/EPZqj2lPNzPMquw
Gx3N8uAi1YwEViV/WODhyado1c8Tj4Eh+tNezaH3Aae0VYTiwui/NDiZ6rJRo9i0Ydrahgr6JZzD
sD+iPk7Atr2DT+/0V7SJH0z6j53KOWZemjXHr7xN7o9nxo+juNObYUeN3u8P25R34MFEf+4rICID
0orXug7orpKHQWfk7rs1G9frO0H5kk4A5J+GeS7Hzj0GmlJzjR2wvnzBHaVXJ7UEt9rGJhm8Yb5b
uMB27zR5VRK7vqbVKF5toOQ7LUXi32qFw037eyBdTFtHxomgTMe99bq0sMyhPSWh/+Bze9sE8Pl7
TSTmfUWVdhl3EQocf0J907sTluGOjOgUQQm+8hu8HpT3fk5RxE8S5WD1iLl7jR/Frmx1ZPdchZrn
AimxHYt5qYQT9/boTkK+bRdlOAMf8Iu4qxEvIVal9rUumCq/sZXm3KxF7alJth5aK2NgmV5HEZYO
/AVo9mnBEE+ne5LDDe+xFcJMLNZsTI+0rC1tGdCBS9fU2QiwqolQP3K9VaBhhqYdmT0n9BDMRdXB
kKSlucExkHFExEgLAMXZcwlRgvE/em94iypjOq7Sh24dZHgjZzbzyTI3pqma6xzBMCoSPyGZVfE+
BmtagvKEpnEytffmPCqReVJQpW5rVn8EAHJaq1CCynhBzoCj9l+szXAVTHzDXLJ9Q9y/KANYlnEk
Sx2we2eB6RrQbKwi9Si6ybt3VU4GKS3njhpUgmUP6mnSls2x0pK3nl1h80eeuDoj3z4+x/kQ18Dt
/EptvygiyjuBBMCFSGAKeqEITHB3Zo1S2UAYxRNCbBJxpBy2EwIlHyJxLqPb7FdhivHhbHCwRdDN
uflACAlvoI8gkXKQtjG4Cb1as0XUSsACiR93Uj5JkbyP4rU/FhTyoTmbYxkBtk5kk+AK8DC5Ji6b
XKYaiR42JwcZyT7cRFTddi8dzjM0jq1B//B1MwsBext3x3GEgCkUhljzKxF791fxpR0lEroSlbyC
txtjlpsWnG9oHAwklWXON4PRl+vML4AiMz5Rx7IyVggjj3M94eeMCkrl/VizPL5+5pRFJRHx0Law
fEDm9t2WWsPYLHZzRuVMZnXb0ooxo7abamC8poct0KhhMyAye27aMT2ycLxrXb67+PlYIAveSKcd
8IYOdia1//wkZFFiaCU7AS9ZnJaAKhNHmIF5R+NZzJKos0iYt0SQ/PxGGivFdQNTAPOsUm7Yh7Rc
nDFP/c0/bk7ZiVgRF16ExcwzQmA8Liuc/b7fJgWuIsLMhxeY90YZpOgtNWHBPlPL4fEraNoAx7Yw
q6C18QBakVzR1ryP1SZUp0ldSVxaMboiIaAOZrulhiyJqoVtmOGhQ/q/Xw5CFzkrKjUQd///639D
icngftR4qK3WapeCpGq00cJSP9SffTjq0kmq8lLGdmr0UXljt4XYXlB0Cb6PpR5LfyLYnJkpOvUG
9N4uVc7pKcGuIYDhFDqJ9tVyv7h95LmocTe6wA8/Lrzzyz9wuFhwBkB6rWOhjLcgikkE1fh46B3P
E63yDY+F53M9zMRh2E0tSa9gmPJ/Hz3F1bOSLq5Zd6IO+83vYqDuTvv8ZnX5wirV8wVezQBbhIpT
k3R97j0tSDxH4lOontCeevbKGv+rACnnRY2M5VRApisty7vBamfsHZheJe3UJWlGgC0mUzrzujmE
Ugcmi5A31s8Tw0YHYEl48ttZQ71kg8iKi4iDIdr0AjdyKE5qjt86Optgwh67M7iCy27KGGwKkgda
ubeY3VRNEczx+j5yDHRUUcXD1saXJjI6kvu14k2VNZTg2miOMc4hZyI8fGLc5H+7Laj7eYZIf2S2
CPkpNyU+wsTUKHljbch905CoNwdzZdhY/gHhbKouNaG1zUU71m5AoYgmdJ3k3pA1HV+zS9Umq831
ufGqTQ6jlFaop1zrpMvP3ePkl/COfwdLlT9fV7lAS64sWewMzvgDnkUky7iGg5mRuyS1epsNrgsZ
doSXi3uf3AybN7/XhcxETKFm8k/N/s+F/9nd1eZz/fa/dhdg6wA/41/cKPUKyIOa+FHanrzzzV6m
RBYgRibX26h3Ub10dwVRJoHrHyyo2Kub8BvOaBeAAYFbM+Jklf2je/cbpZDGPlk7YSDjHTIlRYJi
S5gB2BxBVhmdykGfkGpgf/2kgiwR9NMXyqPaVISUNmAp/Dzcl0O4dmt+k4BPpc/JpMdPJuSbUca3
sNEPo7lR4Xx53hHo+HZISm0AwGhgSyHA7ypIk32Yb6ThTGqZsF+GFxNoysIw95mYsEY+uvnB61Q/
GenuMTMiZ9uumM9Vs451Xlml+djNtkm/qlzmOfRPmzDsWKrBfU1QwsOZ7y0IY7ruQWZoolC977l4
uOud28UwFVg6F08PrboZeIYLUBkYtzY6+0y+qfTKXlh9zZ9X8UOMfiucv/j6tHQkkVgHDP0tNI6u
9gbnHgnaJYbchZO8q0lay9DuZ4fmsog/uI7HcwM7iVfNg8as4oHAtI4HQAPzXbDx6BRws+e1lsXF
OkerrQ3pfcCDQlr2C5UVxRy55CXn2k7gDda5HvlGru6vhms1Gu0Odd3TC/K38XBy9sxhy1Rg6ibK
c2r2Pnb7z7TfaWUyAu6jg6mJV5aOqOHjW8NAOnG4k+lasTGJ+l2K61YxvTul/PMsZ464eQO4brbk
Qism83SKY9wC3R5KvWKKxv7aRueEA7FRQ9cv2cf0qbc3J1AC1XHwuohd4cTXWcPZaIuK8s+eXKzQ
s9AhFkIl0Mw1cur6ZEBfqF0oiDcIC2O6ayFaRsO541uWXkwcvPKupNQ8/+Vp7gN12vVxlZC9gCuS
mIrBcf6zUC3HtlHET2kiBp5KHT5J605kzOJ1SnPcr50Czx7pB9mjfEHEc8c+SspptVggVNAp9Tol
1P+fnu5qYUiLqcGvXFJLea7eT99QlYQB4zGR/TcV6DD/haICnieB7BtqQmg1m1DatYX/eHUn5UhR
qcH928aVEn7gBwD/HtUmP9OSwYZHBnm2XGTfa3DaVInrUGy/WOBLcVHu9m4e4TZge9dEDAxDgVAU
s59WfFUTDJ4q4AXfI10PXChsER1txi/+L6C0A44fgc5CzuJEfIToo7eTkHB6Z3j+QUD9JHJr6j5P
XPo4s4a7j5q3/IPlmJotBQafo/5vCcU1ekYA2Lh8CqG6Igfn+mS9w2hiLgJ378mDLp7q12Qduj/P
VAQjUlXbpZu+fPkQnXHtRBeHySQ5fpmKq+gvdj6DPoHca+VNxbCD5cdVNX2sr3zK+3yFpWYhiriV
o97lftxyx7zt8Q01QuhH5sb3n1FmoWxIEAWmyAmWDwJVaJVPE/319ddJhnqaPCicmbEaZfY6vDXn
hcX31DWlO1h8buWPdk2pwG03ADx4thvfyzrmkMVxXIkpVUTCYa4HeMG9FKZHrgEIgnGrAkNz9AUl
/3ZBSwLCDkmArDYhG69srHTFX3HcLr2j8QCGe8oE2LDXk0cG7hbbWTdTt4Xpdj1b6wO32nXTIcsW
QJgnVD/tLjWMnZBoc1TQ81tFKV6mj7DCNFtD6VXXmaRAw9535BXt6FLvoksltkJrwwIlWtx+i/ck
oUPKUers4YhFZzTx3tdwo6AeVz58tyoOUy5Z4O7gtQRan0HXmtFbWQp1hV/qjkxTlT4AqD/PlYD5
5SsPv1D7Agh2cDb+SCbrBL7D4cXfQ4QZG6Mwqc5w7zzZ8ougyi4rK+N7yXFDPpJ5rh+AHpjo4fRe
nUAaAwola0XXcN6UHwX9m/sBU/I2Dfr1rXQ5mZLufYbw0fBnYY6Yq3x64xLxRt8RgLt1nPOL4l94
+Rfju8GTEmBCV18qNrHjZctsRgMCZ+znkcu35bDukA86MaCYfr49e3icAIgwLkouL0+PAvo+iwBx
6a7ulocqqty9Sl/7pUhsfscyZMG1hfuV3lQeXoZ+VaAL3LA/GnpE/jjKpFJPDpf2o/EctCScHtGi
vsaj0TiCex/6UQQi0om8Q8Ui2I87XSbasyRKCCymO4zWUF/NvaPLEVslWJl1hh8jV4eCC+jwntsp
m+B1ulh3ARZ2QMrXXWj1D0A+aWTmALtBz5d9SJzc2PUGjVNyM6GFMiSm/SIDy9qkDPA52twgPxgv
xgucd10jlQCQUncbGy6y2AIJLMwZ9k3SNH21m44vL+OenEDx26zh6/ZtKQzizPn3nxOXzOmsXOMp
5kb+J3Pl0I1/fI03Ayjgx7rhdn9+k7tm7jD18oBT6Nfu0NSJp2ZLiuCYigPIY0S9IStRKiDMbaop
T76WnjFqwcgfykoq4D5GwQ0ZCaOKAZSXiBxZG/Tv4JO34MY3mgoh3eWu4sAEbb/Ilhb9Ma1ofkEm
t5NNDs/Cz+Mnvuk6TnGVW/J8UV9Lns0Z6RbuFn1R2CGzLzLTZHgyWwkKaoAi3vE1zyT1oB9yVRJo
ru70gsGrqriOMpi7W1zJGyVIdForGzFrB92qA4cxhDWke+apzgBO5G0nO89vgVSUpzTNDMu9IfLM
MEwflsj8HESYsoj3ngO3XAabXSWMaeR3ooOEsdhC70X85UNwSHDwXorYwwydEFm/w5oYxQw8cGW0
oL9gTwlQh/VcEmxonxmf4iXmY1c36n/jKzZR98hzAvXjcII0lHvEV8v+eNiyIyP2p8MLdGrp7r++
3YXE98kWbDzd5x8PXg3Wl43d5s9sS0+vfKORXoL+MEPm4UMpII04EoJg/b+Q8heaZ6VXqyUoIkjE
XgODNQQfWHb5qBlhJcxKyYvMHYkKSOA7ixZT2DTKFkdw0mscUNb6GiFaIPaEn5ONvjJsVBTEsLVU
GmqzTlAPk/nsrFglKpfVjmG8tMFscYLalyPCKZasY4DgMbngw0YbfOdfg0n2udy26+o2ezCjGBnW
rpq/GKnRGzc+dA36Hec455cihicGSHJE3VJ6/AOzGicFGYtktuk3g6djFJM7v48oHUDB0TlulBOP
vpyCFFV3UExjG5Wh0l9q8h39Cj1VkRkOMFNQqLPotr2ob3vGK8djJQWAaeBNVLeWUcb2Q9+eZr6c
miNajtKYmF6E1FgOzic8oKfMQi8OUKCDNY9Sm+BjAysS2GS59Oa0U7BQCgC2gmyoknU8W5RznVJf
SsOAmS3XICF0oUUPx8iAjhOvdX8KQpvGU7XzI0DQFE51gHmZnHJLndxkV43OS/yVau0IWD3uV8Ia
eyY5qdh0d1s5veZLuzisCf7ekZmzqtJpx+avjPyaOsCQR3E5jkUot3KTnqF2E5iVUB+Qmm2eTxu0
dZiCmtJr5u28QOpP1HQGuNfX2H5MKjwDAtFrrIgN+BvzB2lWEB3A22UJ7TwfZSgDTWJAJL18L/KR
0F0ZWiPvlhHbIrAZrgfSiTYdO7nzXup6cDaMbgTR4aAPNNzUuAuxlXnR1RGSbRkv+V5nFBNvhA5g
NG6fq9bmDxpQnArXy6eCmpr2zD+ZRGpjj4eqODg5M64yCYmi2TWf645i9Yy60KMmj7kTAnudeuPj
JEvBfaGtYxf8hQhnCf6oN9Nz2qwqG6gEttQmTZgagvQKt/MHmYASnEk15wAPmiCMM92kRjLIMDDs
uO0mIUv+QbdasqNYbuI6/Ft3dCaqxyfxYqqjuxa0+F9Q92yw6qzyoQ4KUR16PT0eYJ/cUhQkz9iD
F3mGuzINe9U/g3K0IF+uRDnN+ye5JQaAi3n4SZVSX2xCQ57vneZGCB2lhtsaNiP+5YCyyyH7tGpS
zdaZfoTjXYKG66fjH3QObH0+zlRH9xvIbn1MxGfWZJ0LVA5Se6U6zFdDvxbUDPKF44SehpeCy8e3
yAb4gYJQ/o9VhHgmt0mqdHi5oMfjewBHwFADnTnRUdvSnlUvzyfAjDWoEp6omBrI31Dd+6CMAbQW
qznILrsfV/AVAEVq7IqWJKCJJvxZ6+eF9jGLWRoic5oNGgPJMkECBWq4qQpy2CRFFSaZlVLY4UTP
3P4tL8p/IU1EbvX1z4ZuVYZzF/De2meG21RpEmRNvsK2U/RDzAbGYJJlKOVlF+hHbZN1NJlL6YMU
WxQFWDyh2hF+sAg0NUyr4Gj3CqI+vKcGAt2FrgQwwWJh/V814S7GNTiQV6gdOcR3PcdXbCDxT/x9
/uaHX6ecWp9/nM/TawA8Fly32uIw+jQHzZvFTEWkosmiARr/Gfrkdb6Xhu7MtjcVnlShR6t3G8Fo
ZHf7JuyLCrSkZVcAmv2ulU1jkxtxbQyAgrJWnvkFakYkJqQ2wIqABM53sCLSFQNOoIPkJtNScWuL
e0zHHTJ3hoaFv69LneQAHbeH4GjK/Qrr6GB4joU5+/nvWwxdC+5YDxMK3etAA7dGBgxTyTWfuoaq
ELe4M/Vx92r/69t6U2qJQBSZZebSgJaT848g/llSygjk0fRw1Zs+bW2KIejDebD3zbYeDeNPmvWI
NIxJXOJalXlfsyXH57Ocr+X4+ZbNytvAaxv3IO4hXhCjE1lVfQrGrBDe/q407Y3sZGAMNrEN3R+6
v7AKa2VvWcG3sNGJEVqZNwW+W+5qDJAcxpDQZhIHt+JnBnk59kb8I7oSgP4EkKGJ501npuUaH6bW
QY7H3U4TpX+uJ2El9Wecq/ONwJ4WaaqgZ81xITTzU1voh7gh+Ib00SnLBldrI5f+id+jVYuYnP3Y
tjanXIkELGDbhLauk5IhZWQnsGu5LUuVgpVrjk94bQtZ6XCKr5nwr7fVorzrkSZbUIH77Atxtrs+
KlS6epaSnm8I5Upqsk/tmGVY4Yz6A0SqnLpc9KlDk3Mb2W8P4/szRFoUe/GDFCOpdZWNJOJzbewm
z7iOTsI9ScaqA7Xx826r0sD7fEyBqNsDksTk5iYJJyKOF4VaMbN6DxlJUQI+8UJp1zE9O0yJVuDl
CxvrqAIAhOcwTFn9AWCCR8IxYuQ8vfmEhNcovLKij/1N1ov4yJJ4gXrSA2QVEDg7IcdhHdMXLiSw
sI9FuXtBTSXIzlzs0TQhW7R2aKO+aF/IxojRDB1c6vqYsDcuCG2rs9/NmglrTm0G4OyXF6DJ4DCF
XZN+tLAz/CIbR6MmgudaIZ83UsUxh5bxWfPt+XI74m6T4n3zZeh4/nXrPbaoER7w8Y++jXl1dCLx
6ZJdbxWFrfF1i+x4NkX1TEFwyZXcyTp+aXxk70EBWH/lBwPOR6m3nNg9iXgdmroviSeJkHbVOfHU
O/Hnj3PfXQ3r5BHR/p7BAM/Dlkk0KD7I1gBpHWQPuU/OogqqzCQjR6bDgiLPgZcM/Y5Ae28twdMX
zYME0b1Fwq26dlD8VWXUepDugnwysfRlZgi+4awT8WdGquLstejOnbdaAN0mz3ExfFRZleiREdgh
8y9kqKC1dh95AG+b2VtbJ8TthPm+lXfbR1Ryl+vGE5ocVQ3va0ktGJExRGFEs4FHcAIvewKkQV7p
NOyKCmSMl5AF5oC5ouHhaeLSMbdSeWETBeZeIgAp9SR4Ee8M3g0jvFdVcHWe8PVSD6TkEN4Z2M1F
HCNpW3IPNxu4e0bmlRsfmfpYmxdhwf/aMnweaIz87dZMp8lTgwVHfIluBXNoPOEOaFEHyOQSwuJO
JeFAKwmKt59C7IUbVyEzLWjzY2oAHdlg+qgebgpMPv80UhZ7zyKYB3Mgk1NpNQ9t2g5MRewXobeM
xI6/mwa8P2K0BRgTQhnXnhvhQAagv0adePeCoQd40ypJKNg2zsAKNwBpoEsdbSbLqy8SE9FAnfn0
6mFIETJa2j7SJgsJaGn7k9BZwSN5f24LpYhRodMEuqW8FGjv6oeZoW0z965p/+EVaGRO60SicHI1
8HC3gSN5lpNFSIDkpq5vqMrQaFyxlYSRANrHUIBEWacLAIBTdUgLB+8xSSzQOrrWky5AybBYoiIH
kGJ7O4sxmC2qyQi+jMJTvynSilvbcbD3WUe2KKgvv+SCz/sYEmdhSXXP+yRIPK0o+iQhBjSC4JrE
5+3qnlKJuOrDvCMEYUX8eTqqbMdFEoZFo2QBwafhI6MHL0zKb4f35O2Nln96+rvqOJ7u8J9v2cRy
863f+38EpkozHVGgFIsNOcPmirR1dj/bsLxdYuvCMR6tiCKZRDxYOdZUwGovjhZOlIR5XY3xQ/x6
UMqMkjOr9urWRInOwJtWan29bV3xyCgODsn5B6Kr5L8/Ya05NYS+i16cnABCf6xdEklAHrqikpHf
NKZ0pv4z3Iptzfn6F7vRLo/J7CZ9lTnE8glS+hnP0/gRawmY4jECYYHhT+KYkHOIMHeD3YxtpVwu
9bhCfekoZryR6NE3UqMWpVvxA6F3zjjxsc56NhKqQgp9reHkwlFc654Fbw4rVRAhxdMp2sCYpAOl
mo19mVdgTiKJzmLKcD/VMVQ8mktQluVh5xqkZq+pf1VoQBm/uCpfvWFSk8CGtVLC7NBoOmvJC50D
jkdlP43KR93cN/233ydOjoVg9PXl/oM3EtZ4LexeEx14PsTWxK4Xwg80nDiG4CD6O0WYBD0fz4Mm
3raGduOmDsZUXCr36yZgLbYiw/ucRXYdt29M314v0gdPCnI/9D58CqeSp/00wgADKI04yePXFbQI
bWxsSaQOSjdT0LCB41YBuhmr0syz95HNDk3bIYOJZ8lSKVG/jBdKOlvDjPapyGnsDQ0kjNloymZ8
8A6OViZgiESbX2cSopsRsDGpM+QzYIz+0PPP8kjDMquQBOc76d/b1rrIx6daah37yALmoK0C0BGI
o3iy0e3u613EhIfsbGFF4O6OjiBePK7Htpy6ccf97jM2380B4iozjJzyIVsjq0NNK0yhWQwh2fnC
ZLNliCRgmBpHE2ikTdp2HK3OSLulscMI11lYI40ku4K2+EJrP5uh1MoXRamF6rYo+8baWjl01RrQ
WpA+oAAqhapmssYPji9+vmvoLoVetfuSDMLy6wqUVBoqGhgAFiB0JI9stz0t9N3pUSSrIgqPurLb
Prh0X/E241eHJRcg+VIvJqtG447JCJZKJsFwKxR5NauEj6d8vEHWTKkHDDFNzL0/9BHE2UUr4DkZ
2dM2JLGd+xUOdzqlgp8PZKybB0jM460UAWnT2sjbyoMbgPMtq65/zXexmtAHxjJj2AmSZGOKRVtR
I+itSokNa2NH5eSi89G0NBQKd3shOOdSvIjH8eFgoQgJIk0vvQwAro3ZANGLAmRDS53T2cqgSpxT
zvMHSkZ2FpSm2iFLtogz3mUQSUlHgPfmUQ5EAL04hyWrkuIb57L1y8MCpgwaZp1goHmz8ZI5Vu9q
XM5X6szBkJrVt7oKF/CxOWEyra0VqULKkxzIlGiV5xU0Bk/jwnYs/c3nm4c6GntvPaV/VMc5cTHX
bPMH0mEQtOxzvJEZXQxn7aesHv9WM8YCsO9a4yYBMWOncuTADh/M6ToBJj7BKAvPzPNuRGnRp0rN
9g5sldeZWeo838zQDv5MPn2ciijNncJFC4pohtGNdteffw09vBqAmPofDvqaWVnwY4WIogRh30S+
ddEPr9yVA7Y9+NsL708Czz9u8U4n8Z/zJ5rhlrvNKbmnQAiwK1KwPnTR1heCk0aGuU8FYa9zx2Dz
loTrD+CIosQtAF0g28HGoF2lqYEYd/EuFP3h2lRgSDDFYaX6xfuZEDoTvvzJds2MMgwjhxCDSN8t
uKFjx9Nup+6V5us5xDJtBUutea5+vPAbMBA+xUMPAShgIff9Ka+XUgRp2zc2WF4aGEYfNpVaoLiP
fZDIahQuKNYOrRkt4FdbWHBOxetKb8qcdomZqbO3xwEyoj7xhItdtK0IZYeBZeLjfwvsAl6GWZMY
NQjhOJBqRZKxVvWNLk18JbmbiUV5gisclSbGZEG33wflDeWcADzanGoIg03xBXMMz2d5UR84ist/
KOqrg1Jz0g0lF5FzA9AjAy1ap0BeiiCzkTWKuOuURM+iX32FGy80UYF2d25PIFnd03iiUJPBDCja
w+gmpt+JdOMJXxSauWQGpw+Xr0hJw5d+L2ciAuYhYPPLL3/tLA7Ma01UFFuMRWo2u2SOUpbZirMt
22vBH4yGZ1Lw+2TEkK8E0PqqvH+lo7nH/3mLm+3xKYykvvbDwUSIS+ldQkPG0XAtUevfoGnUU729
gSs5EoMrtPhvEn9Z0n4n/wzhZRMWIOM2DawOxoY+t5Yu+L4yr6l6LYcL2eZPqx6Ymq7ctD3Iys9U
gywIOURPOat4r3DNPRRIj5L/0xUUICbWRGEJ2mZcicZpTXK2n9w96r+vp/j+LPbx4dbl1QYxi/0p
DxAibDswjVgdHY783bCW6l/J9b0TauFL7f2bM2PQfypUsgxzDcCEf1UAl8TljzuNfdAkbkNMJ4wn
/YV/E4fIcZdctajzW6eJqhx3yOxTJSfJpfiSkRCVHu37DmZO9cPicVnHU20WHBrJmDfFr1htU8kv
9NmKO3WKsd/f9Z+8njnkJQMyk85J7zbqQZS6r+dL/2GfU8FcPOZgrAwYPVaGakdBrH8a1Gfq8Ole
TabCtGuty0x9ach569PbIuKZdZHQ3oGHkDUqgvUBL4EuvMfhIPmXenHKLfgtFNPOUMpigxtZKuQw
sTkGS+eroj/VCTYe8HnaHxDwWxitnoSu5tnkqBq/hohOL3Vdb2UnZbJSG4AIpIdMaNe+9zVw4+zG
9cb79ql3R3GuWHkvEf+ElCg/sQlnUGx0ho00fb+z2ejdIL1Z1Y9yPl0kz5XtuoPqccC7mTcETOUW
SeCArACqUT73j02pcxYy71dBUmUGwiVK3ZbMuPZfXUUDZQZb3hgPp9jK/emQ9ReXiHIPX6egZGkc
r/IV5WG2lfjyJhQaCLHeMBlfyfzOqzEXFQ/Y1wri60fUBZozEi+vTCYpjdFVKniZQR6eMFMBisQy
5tnJGx40AUAS0X+J7QRbpQYyN7LckD/FOJFROvI9qJoCIoApIq7vLKa+7md3vYKeYOs19uvAR+nV
htz3Lois5yUrgPr5WzGJsUdLLGl56/q9DP0VcSG/upLCFes3v6CFSdVi7crTS0kmxJxDOvK6jGUT
Jad1IFcg8g3gUQLnf9cy16IYzoQujETA4CqcrPoUm9XfcVo2MgGBUeoz5l8yqQEieQSSzGpH4ZWt
VHbo8BwvUlqGdj9Ls3uBM2rGgB57EYvbkWT9utvc0g9bZo527HyAcNczLA8uCcI7r6ZvzEqcjZaV
EplmJwSlZ/G2kYXc876QGt3vzvc2iTFOpC1QARTSVHArYAXvTF+p+QUTq2g5ApT6WeXUgDATV6y+
0PICKI+agRE8s1Yf4QgR/h6oUudrgHZTtPlUUBhEtuxs4MEV9gLZKaVaxQqpfPRPAaY8RetUvOWx
5JlYx0pPvPV/K6DkTNuE1m8VEKStkPtmK2TI4t5MQQgx2XzbcTweBFuC9wmYr6fXmI6uckYHx7/V
V36cahSm88s7I3A9kgt81SUI6mVsQLbMg9PvSMjZ/kB23CyaQOgQd1sxrLgMpiRiF6kLF9vtc3UC
puE9COoKXbYTGJ08AZJKg9Xv5XEc0pBpB7nLZ9xG7zIUMwM+jYJSQbJxW6ue2Mx2vjSEkdS6692E
3h7uDmzQUqcFneSvPCaYfllMtzddXVO80a3TAUfLspHs51MlFowV/8OEDi4DJ5t8LMJf8Vsu8Czj
8x3ZUWtxN8xk5MdovtYgeEvvPt3bKPXnsihCwoVu5ihHZj43zJR56quKM/WFCwUsrQsntX6k7Nyp
53rlPw4Oe7Z4oKpWLomCHTN8A0dfDwhaDplyL6SuSIIAncMGNmSlupqgOaF/56mNJ9pxtMk/I9Mn
OzYvD0dgjhNbwWYepmM4iuPtc0EUdVgPnV4gKnxM/KL5JL2IRShE841ZkG0lv03OjC5jhFNGwZTQ
+Q53i9+UwBMUpAKeRLelSG5rQQk3qb2j1rve5vcjSNPv/4RTmIkU1MoIY5b4rRcNiMx7TWRt+Ae2
/WZyN12CQC0gCu+LQsK1rr/S5+w7Fju0ahrRhRZ48gsw37ExOgHPkk+Ra8NtOQrw/B5oM6XItMwU
78UOMEcUmXMK5Ngf4LPliWR0wnFuBtjTVeRPeFRVSLbZSF34glLkTk6f1jDeoMqTTXo7DtkmUNEc
T3Jnab/yTtNxS6TYM7jWGEFuyy57U2HDt6LgID/pigNfQrTvOWOqEU70/nSJj4HtCi8xD5hS+hOo
Xw03RO9xvqG8XUUYbxHjEySSNH0QDOiDaFmtWk4eFSqGq7ej2QMQtXjMg8cXRoBhaLRsa75ylkyT
wz5hmrwqD1DJybQ3OH0HHSiV+wOGGmBtTHe9U0uFotry/9Awkb5IwOE3VMIfcB/NxlJ8GwbFxwrs
GWlQSI4m1Ja5Uteog60yJa23V8DxzIXe/wOm72lsPo1gr7us7zrZND2Zqr/t3VPtbgsDpByoXBVE
30/9H4ukijqdP/3hvCFBgAQeekCnfodK3w8iH6+YozHL8zoygFLum49h0B1GMureWSNMSfUfm5YP
3CE1PtMZ1TPy0fvFuYXrh5SUWWQXbtq8qrnA7m9Y4G9jQkUwrKY+1KUH2JFJCkBPue5M3fFCgjfX
8KpjenN4jKSKJ+6fgZ4r+h2pNHCUhU8hgJJRiK21TKNpkBrpTdK3Bf7xc+mNTCfGo87uGZCpC/CN
Cw1UMdMEw8jUiCq755JJwoyjrnl5OnK+RR/WF7mnXePCqNyD7XXON7CcLmy6UFU/lUDprcYgsS50
/ui1fAOcUYQLB6v3cyVskQO1rg3robunXBvhnnEvsxnkUWAAqP48qZXhIwQnC8j+IDvPYyjUIVRg
oIpx4cj2YxcoEbnd2c8vSprt2aIQCYaW0H2KxamKt7UK1y/As6NAj1V9eaylflDIHvIPPt1omxeJ
bbwLq/8ys+bBfcueyoOngQk8J518ElF7s9qtS6ysSTiEA6vou4XbWxLRbcGG3Sx0PT0vFemR9WZ8
JtqGq0tezuC27BcvX+9L924amZSMLQ0xAkhqp8PMB4S7SZYeLJk5od9pl8SPHu0BTcnJnQ/etdgl
n/Tu5aUhXQYriL4+gR6z+ZCZiItI641LPxRvdC66gLS7EJQEbD5qJcCUo2GZuk4ZEoL1WOufaEcw
SNQGHXTLpB/gs2eIDt2epUCFkj4FGe2QZXVKfDVoVIjL2ds3hS1tvLlYQFuYtnkpC8FdMl7PikTo
C2lZ06OOmJYz7HQYXN5qHpFIIDThXte0s3Y79hZ0H8uztBaW8i503faqA11+hhgNV8BGpWBxUHmS
ydEpBaVhLqRKqAww9fQvKrWMwf6VCBWlMzlauACNVgSKPSMWWJeSfx0MTB4fTGzWm9yzHeTK17rI
LvAeWaiRn2Z+LXenWD1mbOxVoJNJFaQlKDnvEPW71sYMAXRIZ/q+6tcfaYLmTcA+S1mMGKrMFWS2
+wraJSg6M6UxspNdxYXT/ZSIm+1vIXXYA+29KaJIi+zfSgsVW/PKb9+CZ0IPMMEhTGSI+vN5FxPS
aaxmyKmswg57dpjqR8C/2+SH9GT8MIZXZO4urPxgY5TjdDISTsdbf/vI7uHbO2eqK4yhlf78uEo/
aadgeb7EyH1zDK9JY2RcWm/m+pyCE+F/C0yJ/gHM9a1Nnd2t/AiI4n2CMw==
`protect end_protected
