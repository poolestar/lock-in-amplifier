`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
FWJUwQjBjmpS5fzHVnupSDdqmhC2OFCDg+mGSU08WuN+lNcAeoJYKUUQnaRbuv2FH+Sea8YzbrTv
KaWZZFlusw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FtX9k+Nhr04u1xwEhivd/iYo7UzwiRWTKKkDUDMzXTfSnQa3202aN7pNreKwDtl86B2aeUD9uhoB
uyqh1uV/vjvdtALRZfaugrlTApN+HCnk+zGLSYvoHxa8JSj3xG/GUae2C2DK9/DU0tO6r2Rr854O
RjsemBgkTRdtQNEFOrY=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lN6RxOt4Q9lkXDV1w2WOP4ecEiJbRxkZrxzD277j5dJHu2HqHEP2yB9kJ7DZqiaO/sNnqSJOAxLR
9MF7loAm7dO8RZN7KYbrp8qgED8IHsYzlfwaIQT+CRPripdqe5noccULLbeqQ+9snazw7uNWdMb+
mI4OVjgTh6MUvUKhulo=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
zNd88nG6vyShPZz1xT3YuldJFZngkUv6WDSwHyfJr/r1ZLWP6fVqJiMls8mabWQfq71S5lrhKx1e
+o6ver213W7V7sCmOdLfbpHYB5JtqcOIA4WW9k0EHz4RiY7mOxKZGLdrstpLZv4lRs1HM0hAB1dL
s1zREsNpPZqUxWkzZhPtjHD4HOUuh0wGZPmPkvbFU3e2q+Jp+nrDMvOj7DJHnAp1HqiFmN7WwogO
da2/VPgL9vVF5qQvTVGRa5NkHg/XbyRX442hRT3ozJm1tNBZD9uOaRuoU0F3RVqEtjQPFS3jp7eO
gRKtaFU2KIhDAcyYk/LufyEQiOFao08Ea+735Q==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DTIVm3D2Qg2CJm4w4QG4loWB9rWRWi2FI34aM44klha2tzHLFHO/meqhDD1lvLjCqOJTLU2M8Pma
8zlu5SCg9/gwkaxnYv5mkYWytplbO0H1kr01H1RznP6MEp5DoUGyMpK199edCkwksrPmNULxzehX
ky8Ma7RNyOs79sdLwbpKFsa6XfNLZzxP7X5xhIJxcAZZnFFNZumYa0OykUZgtwKuPz3lcKdMo+zc
HY3p7u971tIRBpwxb0FLmBRiBsEmFO4YoUsHGNrWFmehQwXP6wANiFPSayNMPBCH/5hETYi6op1s
nqwwYDcYawr9/A+xGHOb71RqpqtVtWgonq3bpQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Sx5PmlDPJ1RXJSuT6bfbdeQftlN4hz5c8JsYQ/QbhvUbJ40vuDYLpROJVUIYcSEbeX6IH3O18J3E
j3vbfDu/NBXjozPV9IQPyxVz/2wQV/VSf8xQnqFFQFoj3HEAB8Jwq9mM2C/eNWrigp7i8lhdPS+n
RHl+JlINqid6t5hw44UiKqWYZ4QHz9FNP8XlBPPsE2LfTx+vNn6WfVUySiPz2j+QpxMpd46CpsKe
mWIKt+aiaIgVGz2HrsxswXrbZzLX7yueyv6kErZBxbndlDXPVIf/1P77iCaF8g+Za/vI0HfTYQKq
HHlEHnUZpeq1j49KLB5KljK35qYeXyNgBxfcyA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 122928)
`protect data_block
d7H7VE9x2rIvg3A8GUNQ6vl543opZmeaTf2hEbRRo59b0SMk9kDOmireMfFdoHtqFe1uO0SAMfsr
QSbuQa35IK2nEpiOCA+SbthThygCnlU/jTFR6S/tS1iGfOshdflRQ3ktS23wWcYsz9h6tDtLITvA
xXblSEcduhoYBEWLl9JOfnx/+AUR0mAPcEMaW/G7mNPU9d7ZshRxhxy2SJZZcVLHwuBaJNtzurMh
Bwti9Ssx0dMyU85qqTFOIkjhFvK6Wgyl7d+2EHNF8EklRyK9wShlLFzTA/UpBLMTkdYtT16nNM8q
BkE512Wf6tIvYOnEf9T/q9hFYlHano5x35a3UJuE/tcB3S2xhY8ogYTNHLjXLivJWw/zhk3vsT/E
aiWGVjS41cM0SAGg4B/qzum9E/SBL660C9D3sU7i9bRpl9/7hV6ZRmfMQvU9ARpXGZ7/32/ULDcC
DnnVpyw09ZVWhQelwjcITk5jaAN4ISnKAoErxeEzF9OuChacz+oQmHHcKqIC1oOuWG/1bdg61dh3
zgRBgIfLXCTYCYO+w+PZuhZurgWcojmERcoNkKua2C0o7QkVRK+mkSfG7xhgKzTGjQIxiohOBrxl
4ND1WkSPO++WNlXzh26suFxuqIzIWiJ3yL5wPsMFxgPLDHsAAwS42ju3OVKs2o6b7JcWAc5LXoy0
GccycVypCMAlpXojKUBLBsJoTlD4KqBE7bq7wCyqVz44cnG+qY3U1sS1AGnly9z0kb+BaE265DfN
Dom9dnSeYLuHrLfW8tvU9+Fp7s3RQ28eVeju4TvcpODctuMZU3Q+Gq7N5DHkBOWvGdFsuR+ZKOqz
Etdjqvs63gO8xurrmyOYqdbylHfoRAlixWetBZCcISiZEECCHrGnhiEXt0M2hWFwf0PeySdpUDSo
xva1+HCPCkFk2MDmY1DNAJzeceAiHs0eM8ddB3eSgLzu5CCv0UmOeV2lE9ifdDV5kbUs2H0f1P/z
WmRXnqIIVLxpuSJwI/2dR0IcgLhu00OH+Os2cF89b5RTewiwJEBXdwTB3RKIrkt6arVnrCJ+HY9S
1SNHpwunR/U7iEWh3t4N92Jo4CHogYs+5ncIHceBMavqYBuK94mK7pQKg9OAUBlC++u2PUWvF9+w
5+seCkhA4Qnqs9dtmOGtsCgjrv701TFce0jYykPjDWDHUJuqWb3luiSguNPsjNbNKmB9rTg8+K50
IdwAVeItHcwmQAmkIWs5AhMze16SAsVd5bYYGUzFbNjd7o742fsYF5uHzv1+76xENqrfA/S/E8v8
JeFxVAymhl1ydVkCQKrCK2vPxCiErIX2GdAl2/eo9hPzptFAdeBiS9iZ5uf+4IdUmY5TykXqamJG
4H9fClDc+Rnjdmpg7bv91VIoLR2/IsJ/IDeCIDI0KUPGYQWO9KGt4IKgavF0zPrDJf7/otwhKfA9
yN/x5rWzfFblP+6GWI4DLr82+T3sWspzOlU6+U0Iw4rlxFdhvleDVlLNB3o40ra0OsWEfEaNQvm5
gEkd49uvUhu+2OcD+qLWUQkXfSPH9y5cljXmS4BhcVET+YQE7+puLxyOhpsbhRcZjIc4/iYuaLD1
8ERdvlHBF9a3CNlldTqqn9ds6j9Y8FnCGwYPYmRPyJF8PBK4p8jtnZf3uR9BR4B+FUhavira1DnL
ALNLSutVFptEQPxKEmc6Y2CJlAgZt/g0/efBpZnZzvt/TNgHip1QRI91MMPh+NvwCxfM7e5mmg4O
wT21r/AwfzxFu4k2WrVw+BPp+vEPi5deRhAAZ47KjgijKJZkctVkaMGcDeoh5UoNtN0UIe6h23JW
anEwolQgrRSbNMOhPdms+LEtzFiP/qK/yygryvAJUm8Q/VUI6MLTVIaT4RzDmqz0Twxg+xQ6g1tP
XTfDZLJ2yLWzO6JRQ4wOLzKeTt0WZtmbwBZyOOrBKlw60V348N4cIdJlVfU3/tPlivGr92tWbtkK
YzXV6zCHcHquEvHnxewd5Sh7ecrDBkOgS4Tx7PN7cQpAKA05+CvCgwR7jZOZs1Jcyb3kCBUtoRdr
MPwnfJgUaEd3D3vezdgMaAygGQcrs24rNTNjzZIPxMZw1f/pGw7tC4G2dbJAeLNeieuz68qSb98W
Bib2dhW8dluizepHkD0s27f6OE2CI+9ZwdGxDPm5mQe8spmpcsqGY975KWojKEzbiauzXj0BsKfQ
qkdyC67xRCwtFasO0/tzqmC9mGV/zlya8tMVAAPOn01zmMKUFoSta8BHspF7s0DF1ySGaOhMiKf3
mzNch+MYdusg73dkIK0RAfuiF9Nx1VCuvY2djVlvssSkw0902BPXgGZyNicFD0qJ2AisjYql/MNw
LZap1Y/mbbQddhFKMEk78LpMjdWjJJahqURYf5vT5LDjtng3wFUOb9plz5paWNJa05voesmArsYX
eVNKn0vwJGlKtpMlafFaocUg7ZzRoQnVjvMCJA3H+pZjG3MbYqO6I2iICPT08ZVPWlugvyQvCaJS
3Z5YJCMX3yRw5hJD3aol0wyKAeu7R8ItvwZL3HDkZU6HWHiseiQmY5dVT9fy1KzwU4Y5HjG7Zt44
ufWLMKFou/qTldx0tnfzQEYFOE6xd2exn/AGSm4E+jLDZIp0IawKWShA00ZYfR3I58lESS6QSP5I
VqK/wzkXerWSGUJht4+eG5qVEVqipq6WRaAk4ao4PZoI2hBs9QxBeLWX4QMutcM8Gkp8lTDH+ttE
z0mLPY+faDRT2e9icazIsqlEW5BxPBd7GTH17yK0i/X7RrIenT1iAeB7Hl4im7iAknWXLAIpSE2O
yW3oEoPnNKU9U96uXeFYL14/OH9puXdor9j1m9ThtLJFsFhkrZVu0UbA65y3v82H+A1OLnmfM1ow
Brj1JnwkmA3O9xdDxPkc2TiJZYt+xHOVxTZM0xzYvmF5Qj9NNuyiRN7I89ZNBO5UIuKh4y5nXcXh
CaV5AYbHlbZeWEXG13ZhgISq2z4bQLBc2sgEQQGLaQ+fySjPJABMLlhKXBlgESvZ5Dt6FIVsNlW4
oQCp0ouZIUaPs6f3PeFeKkjhvXgiLy1WEl/3K0ybxUR+0RhPUWxV0aYqEk7JRzX6csv+DSpai7jX
GwWv/5O8Yg1E5QVE3NMSPYFR5HBfAqgi0oBv4vqSEdExfMPgUBVTIzdKXP+++UuQ3ZrVulBaCKTA
RtmNaMUu372eD8BN32sPM4tjBiKzA0xuAfFS5gLGogL4PdBGJWXv7OUugohcO4jnNIX8lYFy04rD
hu0+XWVAG/2fKcoqyHv2mySxGyj98nYQ/3Aj8tynAWV01/DUu2KFVj30h4vg7PGikZWGN+k8PQv3
4ILF299yM2JCkvyPZoa2LEAQkzeEY7NJNN2TxO0ZrNae0xpSy0Q2K/pDhEqyZLy4Aeb0uTIuOMUp
NGrQvgEhSli438b02uw6QUcno1sS5UtxnHx0KmE6/JN7mgnKE0zN+VXJogNJPqI2s5tp+xkbB/DW
CwyQFExG+GuxVWocMl8+z3NNzvAY24tRbly9ewJQw+G9XL+RKJ/AYX8N4hkJPAopJ4wz0S4UIM+A
JDNcGXV1r7YWpBEm05pQ12bswY3WZuIvlVCTsQr+ySY4h9tpxfKzS2ES30eZM9Z66SV3tSbTWAnL
ccHG15Mn/JtR5leQAlsGutZ0Dl/U68e5I+hw+TUXFj/POinE1S6T3y7k6pk46MQzksFoSTSrzaMy
dsq40gi1RKJ7wLZN+Angdd4J2LSZXxYlUTwOuiB7zNooMO9vLvp2q++mSP9XEJDzxPPD3fhRMhr4
HiLlIEWe8savtdbHFf7NR8Tp4NiwbPoyNwd8a+/iEYGt9g1cvIVO2kkcsk8m74j0dSrLGvjBvXr+
XRI0MGqTCbpPAS1tMlVmE/BZrCsg7Zh5eadoogDGj9BWdCGJhMsywHrfT01m+19fRsXpcfWde4ub
U8n4uYmoMHVilqjWFu2fr80/DEVCjWA4+Q3Ptp68Baoi2LuO87jH+iAomYvZbwYLXMgQx7h0139J
5PYqQgXNs+bL0v3pEbZgQBrcZFWSEVny0T3mJZWFmdjC1bWjwmLvqyyKUyw89jw2Ni0jTfREQj03
fa5yzoVtN8AN4Dhu6mCr8tkG1w5qJPYq64pKWgi6+dQR0otOa8ROAHcW3YC8op1GZGnl27oylv/i
dC1lYoOHmyyAAtzVJn1HoZ6Q5OCrqnALUz8gvc46GgCaKer8QbYnLywGRpwhA9sSleHf7YvZ9sXH
RZHSRr83gMqkW1Kz6pgcKEsUpDY1p1HOZv+Jlw8wQH7GmCBJmOgR8sXWHW/aKuZ09ptQNGY4ldUg
IlJl0ThvF0LXw7o5n6vhJCU9RJUrdTLU5l5N1whqO8SmvGr8/gBfHw/Ohkfm2Vien4NMmYs9GP7f
3kBalNLIa7IPU3BrZM8dNazLgTTO7ds7uzI7ccXSBuC9rk3PV2BlO1gXXqvCYaC2pNqsd7Y5OiwJ
ppdjPnsZM0D5QduvuNJ9DINm/wU+gZXH5AB+JZiByWPpl1eiDNpUmOz1d/dVwV3y0IxplRhL+OXq
Y0qojq2cegJ9dZcyldWRF3l9nZeDKAwSR+RRj7YYmhTDnnhMkvtu6Mlx3eKcPafYrLP9tQFT4w/t
AUkyyGbbutwL4tCTUBU55YUS5USETCeNgxe8uqo8ESLsCs5MbO7XokWMByE7Kq9ZwoaU0Q3saE0I
yA96INCRb1bg35OyXDcRGsVwEjI68EybIrhdEVDFRlC8KjEKQfxvzb31HYbt7PRp7U7iLTtKvdgj
ugpNO+4Xyc2vCpM6NeEHyV2ZzLx8hsFQNiaCUS0MghirPcPk1Z+Rs5ZNoty6867OdH/jFTChldyz
HiYCgwEshbUn7jq/kdih2CRwq4uXl9V5O7hsZUjJwjbkaQs4e/YoxZDqLns1wjJrD9VlNbwgd+EL
JrGG2vvVLMe/XZ+JjIM2j/dyPvNAa3+af7b8X6sS5iCVAF07PxXeRcymB5mYexMm2/zsLpuuqkDo
z10sPdj/8T1udulpjM81yhUC0Rj+wyyL1Gv6JwyFGp9jO8Q8g+9YhegNwjXioA3Oaxa0WCs19XBr
k4E5l0UTARjL6rQYDWoflvzgGigiyqD6zTHdOW9/fPDYqYrBL3R/Xfb65r97+gFi0JKo5cYa/Lxo
MeJk10g/iYxAkOWqa8TRPJxo3HtLMpfhsBmiqw3RYWxc09eNZCghYH5fcZy6wKv3h+PrFkBlsDC4
QeNJfVYub5SQEv9DTNrhMu0vhPIX2pyLyFoHRbj3uxa4aR+GKwotUDwEk0DZWxsUr2b0fFX9ZTG7
e/H0CeuitdpadD1du5qUMZVwjgfLJ8M3GyHF6h4sBwNXDSXaJM8pErRKSLUozUTSADDpt5yALGJF
5/wezKGSO6SFkvsAZHTI+2+sMByI7iKFI91sOAGQ3mMvzLuYS9xLv/nlKHsZ7FdDTuyO2KXz5WMq
uuBERRICm+ObwZ8DdLcvcxzaWHwQJREteE6WH1Fy2qXXRhMJJNpGIW82EJwDC53Jt+lJPwhSF/a8
xZMAXDBiWkntGPKk7/takTASvyfIK+U/RddVTyUsUR7cZO3zHJb4mNxn3RKPFND3wKzANSCyRb8c
+NT/qjf3JfKSDbvYjTjXCbW+kqvYZcNGRPMtokbUyVGTKC0VvJ0b2NapV2HgBWnuD8eyVh1pZe4a
7epQAdVq6suZ4oKEnld2ISTXkibBWT63DJZRvqRbaSyVzFTGqVjaORfiBfE/JcDGEwe/qfi5cQF7
Fh9MhbEtPmm3Jl+fc6SAyrzIWBGYujA24ldNNmFLTdUb9MeCytFnWvhPQVxtxZ7VwUG2VlKq7Aoc
hDCne2Yr5OD3BbTARmY/3sXLD0RzUHLITJYLQodL61h+RacKhbxcjQWtxZqYmakKezNvpgrZIpDA
TFps7OILnYvTfIvaXkZT4HST9yu9gdtbXlo7YS4ohBEZNL1ASiShCJsxHc+/XYm97vSBkkrDBFN0
KcIuPMkNM44z7uE+d1an6spe3df/cRP7y1ui6N3ZG+1H1ZnAlW6FZG01d+zzLDLsillwA1PbjiAJ
AvpFX+MqBeYwEVuJ2O6Aqmu+Lzizo4Uw9niLoCQ+HtgjuRGWaUFJHWfw2TP1DQRbZiJx9mDKxYkz
7ObN/zUEOXkXLfHXHmI/ombMrCcdJ9rbLEG4dq5XIRHGpg+2oZdhlJ0nHFdfnHkn2tO7HCpuQ8c6
6/tG+T4O4ywA+OPM0BNs4VG5XA9MJyLtn8C4Z09yDpHTsNFB2Ss6c9MwdQtkklkSym0+qyHthWL+
S7SoblRt/RbDrl0vzl5Y5YckzGEdOKdIf3g455W4wBJxUwTNXu83S2eLjftvEsXU4IZgJFdIvnO2
Viy1jDmpg7YFoU3DvpBIaQPjxPlAC5eZdw3Y7TAaiXkYVywIeMJw9LJeQZZpnzrKnfl55+YCbEfg
6Cv2OW065AsRZgfOxeu58sezcKmaCgoJ68B7LTqCF/dZSP80b5WeQ0imCg+VuObiHQ1nc+hg3BQ6
e6ezGTxE61RuO1yEc+sKUjvZNJCXOgtuSa7qx+1RfkXYu8iugVh2a6vwnMVRNbF3P9JwKLWCcDlR
/128G0tJwRZ/naI21K4iVfedPird4yoRgIxEu5fb4R7KYi8NZeRcycUJ09UaONTNbwG7ljDT0Me6
338/Y/gCCGs8NZ4be+FlmoGKWZ3AssT/NfwSlrKNMb2W7fyaAErhUun69KblzR5zS9oadBdE3GIY
MZkzXUpszZ3TK5Cpj/MnvF1vvBtfGQEHJkvnZ3/ksZPtODJH3sA5GNCG7jI4ikcJZHAdxC+lbzeV
uphvzMIwnYqorSu5gMmhRmKfNQBvkp2qUXPdlYjqA/yh4HfEu0DavtuPCHebVJIBnTe8cWFDgVVY
mpsxHpeUML5ugqJ5NxvdNFAkVIVKE+RKRJPdCUmylx7gzjcD74hcG2B30h3kEp+BqmtrE0XxLt49
vq0T2BI1rMz8CsRDFkcZOZ5ugQnQZCxv3nDk9HGiVgVqMQV3wsReongui5Vxw0I7Ch/jxaqarbe0
0St2C88Yk2XJSB1hoadcCZfJf1B8vfMHngv/xjVIGUSlCUcHVqLWiBUTIrpVhNmT7QG5qnWNEj0s
dmVD7j4QlSw6xs7k10mTB9iVbgiS4Tq2j0CJMU4vskXRoiDZVFF2yl3FCdhnvXJlqKllzzxypte7
Bhi6aNA1JWIynQdjOgclvdOkJSiH3tC/BXLVt6s4IIasRykQQIs3O3UupFE4lQFJX75EXPV5ZYFC
2LixkgQN/QPjYn3GCkk5rTfofVW4dhIBwnG97OnWENIYpEEp3EEHTHm5BvdfPbMsw6HesAxghuev
23beN0ny4ZyrhoTbaz4CU0OYpw1dBlIyPy/907Bcw8eqw9J8bzs0CbejjcVlmboJzmaiu7VWR+wo
Fs0Iy/CvaxkaETd4UvkTTgxHe4A9WHg6cCAGbwD1ya3+nUbioymwHbbOq3ef6n+NWrykm+6G7NpO
ETUc+C09NNT7IQbKBZ2ZjQpXhmp1sazbJu7wBZA8nZzEllK5m0z8V+lnLqXGAvHoNFI3s36msvCU
1cn2DnUdNMA6YOWYbcn+FM507mzGwnhAF/MkCIx8kpnx6X6b0uZS+PozggkDwObscc3lYg97wYWp
oJ6EAZndpSbnvhBqOX6hZtqcTsotBcI2Gqqihrmx8b5TAsZ9j//uh1eSrO8kfTye1numO0rYoWnT
wxmw9AcJmPpbnFz06LzZE6GBVpbgolUcxyZc8twG0GuPlNO7MolcckNDK9u1LdMH5Kio5lDj0tXx
v1gpJrYzQNhDAg+zuso624EvkCCYI3BCymoDeDEifgFOPLLMeR0ENuHZqf+1BF7+ZAzjuLKfrvWb
1ZKYZBF3K4wI4MoL87hsNZnQLDq3PTj3CHqQM/aZ5uB3Yc6mH0FJiD+4COl4lINTqo8qf6zrTL0t
S0Ag28XP2t3PGdTA8LTO1kvKgemyhIbyo2ub2fWl6kjcpUk1z2XT0ZrBYCPPkUEjopXCniCYfstB
UNqVFIj4q/YHEXFyku98zOhtARc3kN8NIp4pEm3l+kl6C6B3hLs84HUU6ATkZSyo2Xf8Q9RyFyHa
Yr57dMsnbrdYRfn14QHaYNNaTCoIeXPT+qETHTi0TC/2hJCEW9RlAtXaMQMxxtN8q/kXfqAmPwFW
k6ApuVR7kLfYEeyq4h5cwTbxN1l6duwFtaAa00TKiu+W3CHUfmdCmcuTDAuqQjis/VOEhjtXgN8+
KcXrFwfKCkmvkug0yonQWTAFJSXVDCDqQRXnuxfGV4owB3ti2BcuYjlZaDbXPRu1e8Vy2U5AjrSq
G3L67nHmhy3EU3dYtRQn8gqJJ2Em5mooCsB9HXoTqz2Vr/Q301HnXtJORUpqOZJuAeXNzLAZPS8B
NdBT+1HQTOpfQ4omdbud3nGngsHKuTYxAGES9qzq1OIEzlz1IVd1ppe0ViHTh/pawncWxn+O6klu
F7Z9ZDjdlsldKNTnaPcCOBjeXcfPvlJVJMv2+mW+WoBJttU+nCauTwTvlNKGBmBmMx2E4DNfzcq/
4tmXzj9JOWWJfKKZnXJascFM7yce6RzyqMUvmzf2Il2w9HplqJIuOY6mKOVzefuJms287wPzGEDv
UsaWO6sQSbaaeU9LT8G9v1nzdI8oGm0KxCQN8E8EP8JvGfTnp4Mv6e7P+80AFonM3pfYieYryQxU
M0sYQsJuM02MjwzY8SIVuLvk3aF9qDt4iPjiHhaveHX2fHQHfkrXUwEt9vvJZElaY1zIdVOwdgXN
ibLF1djSaVTzryCyypLR20zdNkjDy7Ru/pNbMx3buToUKwHWqTiroIHYyKucxS57luhKtDznYRsH
CewKg2+K4hVhdtCqRjk8fmmtiTyxKhl1YUTEXqMkGGl8jVirFd8mjFT4lHiFSmXiaziJBuktZ+dh
S0nUx5A12Dk3rOX8Wrb5EyIF2DxtXR/UkMpUiO71YfcjMAIiJyrSBGuINc1xzzybb/tdDB2Moyn4
8zErIhpe2i46P7SDtuhrruvyhQRK8+dLFZI0Jf0j6VM5XcrpeZuSZi9Wa/lVZMdN0ntyx43CjuWF
hMjIt/MjyByU4yJYR8xc4AeWeRrdrvrdLaxeXOc1iGCP9Kmno0+QiwxTIa3RjqGsDREJR2HhXwMT
AEf/ZuCPOR+ydAQ3FxubcLXpjX4cYnRiRkN+TTXsdV6Mucm2yuLeZfSblBcbtIakRqoqeaWGW8p2
QEhIj6bpmxGjrSaZ0arkkkvblz7ng/31GnAgHtFBbIIlGVRB9a8w5ARpfHtITdYzhc6ga9gcl21k
SvUSuRXau0gsM0YSrtnwhyXad7xyiifIHROY6cWCgWW8TbYARGSPtxiEa4erYUPYaEMZBWTxL8uQ
zcFnzFJOWUFGtQu7IwNZD5hdsfyTfJhuwgbeev4Tc7633ZtHHfekPlKvYGrjGBzgAID1Ba+j1ffc
FeGj+diPoPmvd8yU9eH8iJNBHYWWKaYbQ+KpQ2aPQEamklGBdjhIHOsJql6DLu3AZDadYvv/DCYJ
9Zkgd12yDvgU4dRYR3Qc8THG94Ovp/N9SMY7K66+h/2PXQIJagNoJ7+pZIkFBNWqRhabG0EBfCPE
bR569K+0qXJV3ps4qkfFIhOta7606Lvp25fhAeEH9WF/WQsx+VpaXKkozzxkWTM3DQr3W5azg6H+
ubOln5pEtXaVZKTDueCDL5AjEQaj/yaZ4Wl5Y5Y8jCLrNTg7DWrhEhjN5ezVNL3KLD+1JBXRfArm
8u2zmvkgXIvR6UDEbBH/nZqCnZZQ8aHGtRDa1B7yYVrCBBIc6cSXyZMxMwKpI5Q0hdvAmS8VRmU/
Iw4r/uLjzoiLOWhXa50OuaFsYN7DV8dAuIZ9LowCq6Qo26aoUobObu5fbsGv6O+B1rHmcAlWepMR
cVfwngB+vaysshrk2/iWu6eD6huDXo07SNlDR09cMGlvG8i2GV68g2h6Fn/IqwsWpiA/ZZo1si0c
elrWBlSZJ9eNCC19D3EByrt5NvPUaB3bpRKTMfCdQmkshjCOZakNTYAaNqEkZKzeRxYUhi3BZRLL
7tWMlMcqsHQquXi5lqSTd+CemT7VR42BSKc2g4Ol+3QJ27AXGuSt3WY7Sm6lLC/4co5RX/IWtiQz
3ZnTnbVLRX0duET8g4IeW5hCcCshap5sa7/cj23DwiANP3eJD6zFRGHCLkC2VoHwI9Gk1wGVNafE
Z5iyl1yGR+mKd/sF5yN6iDY66PxsOEgwRvO4FI7PC/4BRTnfSik04tpH61Y+pP2kgdCOrBhE8RU1
DRnBHSh/5deWyIz6TxvHDh5Dm3r7KvfQCdKrLoypcl5Jjz0Wg0Xu0QMAWQ0udS+wyV5UGnAi/ZCN
p42HKnd8IKTj9jHokoHPU3SA/3hdDm8js8vG3zykRIEM/8Om3e3agxsRgAJnx2pBHixWUCB+jelb
BGXxSp34B8a0cW7T8QkVdDXkj8S/DEHRoi+qJgwARDE4G1ULc2CcSz/X0ghANYqpK+NSzAYQgcex
1mQJwyo66X3yRwteHAAAQzJAC8OsDlsKg7d/Zi5cynn8GoUulYrTbbxlgc+QToCZP0DQ4BteypDR
DkqBs7dSeRAzo5avBi+br7e2aKxSdOBYmmIofXtyvz6pC4ytziCeKE29zUjqnjCpyiVjLKyEA/bK
+DmVH0jo/BDJdEIge50hkneE02QAm2eD1phundiNr4e60Q2N9/b0rRakzSeKxLOnGh84DjUgrpiT
n553pNW6qO2r/SZjyzlrzo20jLy45OQS86+0b2zslL94E1myji1WZODpXCOxIU0z9IAi9/OYg+x7
r3/x34kxS5S2DHyW6GSM+uSJfbBzXHwabcEC860oYYq0qL7cOQJXhNujJw3jFMRqgUuSe+DYSsj1
8CUdvyOP+Bk0JReK2GTxCbxW1NXtVzh9JCpwypxfbMTrmNYC7tZb+2Rk0bvNVQ2OqvNBdpvAg0Al
WLNmk5lKo+tKfDb2RasC57awgOfXWXCdKJbqRUtqXF64M5s+6rGeIcj0czsrdxN1fpCMGwhc+nF7
rdEjF4oJW0BRBuRtCc+5kYYbNGUsh2utUmctQph24l2gJGYit2gM9RC+PiTpitUTei3MM6Li9MuD
Tj6pXRGPKqrVe53K2bbpEMfWuDQCLPpgzw1vhM4c261LjlHWYldxtHjEtlDKuMrSlPWeYbiO5PQI
fPLYuK76BB1naKNgbaOmYVlLOVWrCfJWX9ZwMtfLhJe9uTM6R2lKoxOq5gLt37UYLDBOphk0Ft/F
q0XbMx7SNwQEdkxbnoGtECKfZyq8QqNxuTsgY0vwDEEfoLXof86w2HEwNuH2WegURCTine78xnJy
f1h+FAKEf3R0QIZTngmgahjT+mxnSODG+e6vEkc7DSdFtAfnfiTFlhDztqqjZ6VoSTljrrUxiOLN
coTnxH80DfVuQkULDp512WSgzxMhh9f2mBGDuOmX2xynV1K3iCpGSpqkYUlKH+oD175J8d8NERxA
LJ4nkwqRFOpErbkfVbsoLr9hX95+QJMMN3jcu7uL8A7KX1crcOJr/XQ74p2loh7q88nk/5M0dch/
CFIVTpIm1X32hwARvj5NxDJ9U5pSBGnjTCc1FiqrwSFMLrKvrvqjtnxBqg2kJs2KEmPH1UZ89mdi
+3yplrMgqogMG7PSZJYK8Nr1TPkdTcSrv8avxByn8wS+GCxEAIOezSczuDvna/AeolAgCuiZkgP7
UL0XYNb9abSALjs4nnd1tD79ztN6JcVh17Yxl3OVcpUS8xpQcfPfEHSKuhumH0gyCkqy3q81KJ7t
EhwGrHYeUkQwl7jnocbnRs7S3J6CWST59/HwAwnbemEk7eHkJDkC/BJE4KlRwbWeoR30f/PqDFdN
4vaF/RDBnn9DT4TFtFq2rvIC13EiXQFPa+oofOBAF5CMWpDsoGR6bUejXisxMHInVMM0cTpk7f28
zCID2Cc4cL/3lB9P9EdSsNKIvtU3HnGGydR1y9TuvzEpCgwI3+htNGvQx8/MEDNH95ADc2C31HSB
1l9p/2duz0gn+Q7A1JPhG+wouSmWS9AIJy4LvtfCnIfXywHYCC726uJ9e3WGzBHQjZR16cply6Vh
8hsPQr5W+hhr3NGBkiuGlCUWsb9+XhqmPr+7UOwNkGrodHoOrFB2YL/B5PlPZ375haaw8IJYBfYz
5k6eP7gQRUrjrme6VsTygfNSFH3pPuD5QJvoulG7Lc6UJt3ib2smrl+69XY1Qx/raWzY9SSiIbce
bpB+/4r52FBUjUmeTnzkugscmS6G8Z2ZpV9W4nbxqj92iVAjzlDg/WtQDppuuGd+DaTmZXsCPOsH
BO+YvAyreUd2og9WpL8nx2RlKguPgoqSOxtMs9yElgYJJuI/R3ZVo0LZIscvetNTQu2DbJIaAnrX
4XvTIVRWcqDJjPYMzUhQPu1/UYfIXPMyY8XlpKA78dfG7exxSSvZlW6RYGS5djHNpJHUYt/JDJed
EzDrJvJffwAgr1oObtB+Nw/V8US6LbUOj2nXeEmS767JZjr+Mtl0gouoEr2l+awVyOx0DfyI5uqt
+IYfNBchyYZW00Zw9fykmsdZcIlxOwrrMZ+aXN9Z3rjyVfL2loUZVijmX5CklYhe4/MPW+gCD2Th
VSCBWI9QazU/fuLst2y14LWlAbCH1u6Om+fFN1nsJNGatHcxxhQ3xk2lUrcZiDb8URkdXrnwTSQ3
xzKgfIOUm9rjZfIsifS3YLJgmv2lfWZlbG7WxAXhSsKHUal6bWak0yutfEib3GPRqAoXgu/dGuf5
sr/pNW53chwf4N4VaSfF4JPOx3quMXHLlBslneIdvrvxGSFCXOK/pdzrGexcqTe7SauseNz0nhpA
X8eg+Xdhg8OYMYF7mW0A72rwiECCNCQA1NoOYCWzmspf2/0VQ1MLU8pQtuIwbjwLft7eoztGBD/v
xPWWqTZlDRLa2RjwRVlMlLp1SEx/pCHvqvz2CQMJ8g4tiV9uNRW3DNzw/T2h73bAtQF5csmQqogA
PQ2SSgqrX4Q/W0p58VucqS/f87TojDUIElLFI73jTLGiVJc+otg+YMyPoUTn9g6iMJ7dFyqktGUu
0syeta0d2I9Yr4oKKSV0xDdzHjHk9+ZmEw9Uv75yj4LH+5w+NBGvDsYUpnCeNoZWf1+20/RwhTHA
pJggdoAMfBAtOR9IpVPmfHOru5xXB7xRjcgGs1YcyKPt9frkm8EYQShKkBahGtqshvMxa/YnUVpD
82HmoRnJ7mHkYTlQsHCcZdyoskCXwd3D6/jd6ql17+WlMJIH6BAaLB+tXEN6wzYZj3k24ded0pfh
po6xhIdy4u8LdpsxhRFQ8NT5WGyfp5bfpmw9keOx5wRIuV2zIhjlxkcSZE2IgpKteKbiKRYbXhuf
n9tJ7DmKlCnjrH0E/p8nkPbJmh3QWYhKGu43e0KPCF0XRkjk2Qq8gDCgWRjrtJw1WxK7EbM3wsSj
atOY5YN/UrzdXTZurQxExMBNHx61Xtj403e39MzP6aaiZV1BHW6ZN4/PUtWOBnN+ksOCj3f8fEU3
0g1wHmEraMtw6emtbNiF00Ry8H/LEwy0ZdVdmiHNdzPi2/tvx0Da9pt8+xWoneZ7p84uKPoaK36G
NkdWcF+S8exZ2K9gdvFChhD/OFfQ8QyPZqwkokzROK7XMnf2NfzH7pBIQl7Tf7luT+1bIw7bbt8z
UYHsdkiMFF0qw6ORz8kfAp1kT2cPFe++2u1VXt3upvHTEimIihg+3gnKUCT0gkxrF86OFMjMG7XN
Dp+rPpfSx7g6txyE3NpNW/C+oeMBfcb9uFVv7DDm8l80c6Yz4Sp69EFPs96ubBK5+8sF08GFFSpK
HQsuQ0mE+XSVGzyBw84Hu+mscCJP5eNbCZCy9nnO0f3PzHtpQj3PVaMi6aFecFyK3Nm3n5rPSaTV
h3Z/Q8V1MB9M+1NRdG83DIUf4TiCCBCd43Q3CJenuw2DuwtZL66WHGjb5MPPuVbhKRGSTdy3Mhb3
1+sPhUR81r53rxxEf/9EqAyxLUtQrJ47ZPtU5ksAsgs7KfA6H27MKoP/WvueKR1y24ccnoZd7NJY
qjtrHbMTde8vDdRLs38Vcmb4KGr10DkMut3bTm9A9/6wP8Qj+2KNOMdYerxek520nj/7X+4tsohe
BgmXp8ZwvbHOF7gVaSzAUxG+jRc9pMLmXJSMNnFPAxJLim/7z+f8sRavi91dB0JQreGTiyRmFKJI
gbYfVCNt7UZVUnigUkRYB1PG5iKNl1bSf/6fc6tqDROZzuxuztwJylFP0U9IdWkFk2HRngcTiSoH
WL5LhY09gxJ6gmZ8DCBwi3eHaeLHH7qRYN/wR2EuvffBkA/xLnul0vMagxdPEVMUT8oSL4sEJZRc
p6J9JHGOfEHtVinifBsOu+b9AxeRexG9pbALfYtTjQU7aq1zAuORfTmPn1h+VgXTvPpI/5jPjTgW
zRrvz/zPFBMeZJKdsAcXagkSBqiZChj5PJidk038Oh5B3c3HsJLCOT4875CxeX4Jximfgb6k8Joo
oyJQmha3pYvNOd5h4UNMZ111KLiH3hAdbPP4/F7I5fDLS0LFYysh7pHsBYWhOkjDcnvNFhvCuX+/
4g9djwRMO08jxsZEELX7VokR9iGPuD3HPphCUSEG+8uc5lYYEkm7hyIPmOsrDMTmES6LWBnKe0+j
itClIPr2jWDOjVYmwMZQOcpDdB1Wch7UnlXdNQMFziW/IwJSMO9OmbaT6DvtOFiRiCl2QTTB6Xl6
Ozj1OYQl8vz/e721DpbbsyTjM+A7Q8hc3HQ30fR252sIBLseSz/+dw1LLif2iiSPCbHutgI02yEU
cUeLLBF82+68j8MhaEqIrYucPsvqfxDZ3mU0iMFpPjiLXBA8pV/EZwsiIT5xVyknvVF290DE8NP8
TWO3hJDEmeFJy6n5ju3pZayQQA8xYZyK5JXpAAmJ3t/dUpD9Z+aEXJFVjBBesiius1xGN3uf3yd+
N/5i2lpeUhlR1abklIeSe69HOQjWj8JNqZJhppQSNq2czEMV/bd2IhxZbvwB/KvlRZVKTFWAz7lO
Yk7c4Sm6D9p9az7/vscdX8Pa9Tdk4AZRGj9OflQgoU5lEhSB1k+kJzSl95FcrFBQx0sK/17DMeGi
ZneO7Js+AazGUSLBYHAe6GuCIvHYkWsbCi3osyWrzPYVQvQ3XID8moGEdSZjS7tnzT28vTcVQX2r
oPRiZK5iWB9WB2HnkTWrDPvFoKuEtTT/gvSXaoAsKOkXhqk2i/2OpuDz7rx+gy/6eNtfWt1EZN+2
k8Z1nE2XTqrw5iDKqq1OZb3XDLjfMCDgR2K+9tfbgjyTQ4TJu8kWiPG+3V0bahCoThaMYGwwbsI/
nsVscG/86Cycml0JhumeWWsnIXeoDYzLVnEwh7xKkJR1P6QGYiam11xdl1hBR/EBTucvsO4ZOSGj
yvCt6bwO+VMgKCeAUG/ny+/IZ7S09fbHMEZsugvGD3FwEDgHmtYLpolurw/7xCo1BQiIRwom9KxD
PSRzn3aiCT520djvE3/xig0Y7bbaWfZNyo/PvnuOiDZpk4nAtttFhBQAQQ2bbYUz4+YgCYEgEx0I
wwunBjOOG7aXLmvP+1XQkkGBFgzGsMo1VT8m1tupGynPQMTolLgxpOMFgjgz892pENYqNis1yNu2
JGtXENB6LBr5NgRDSPYeTv48nIg8HGlgdnuip0bXx8bGWYn46WKmgYp05pvqtyhnik4djcGwOFqs
V3twhdfnWwK721Dx3aAii1oawnEMNDQLuMoPvnCjMN2QUNfniMXhAho4itvn3LKLroyK97zV5HZL
4BoivCJSMAIGLxdb7gS1lQNozzcPsmpQtHND207VacJlNK8n9+sdC4nwx3e2TfceKt7ODJKDb9FY
V/ymvxfddJ8zs0VhJXuULGEAdWdgVSRoUMbTdXv6bujYIJfWCBoG8hezeTe6o8YPn2WF4VTtS2jR
iaFmZGwOE0SHpNGeqSLAGfZaOW/ZaFDoYnBPJ/vzM9lmm5IIeMPo14DzhGA9KRrdxqlQzYevbT7e
Z4lbupdIuyqXQwURuAq59D9+JKAKJe5dEbLB+n7pi4KPFOMZghMOgPQztCRHKhKg+ujk86+kYm+B
APe2v2/Wqtjs6s3AgevGyrN4ZJPZ2tjk4vbj1fJWsNvNS84F9awsN9GESxg2humBowVNdDtEc8pI
u3U+YQYuBdc8WRrPKiwSbejEF4f1AwJol1dVWPGncOTBblJ3mPB62+sPlsRtN3BEJ5ujY7uCDiw4
Kh4z/gEVBM4/JErwretHWQ5kPc2SP3Gc3wpUUSCq0lwdKTyC0Cz7K6nToGmrmrb2honZnrTQ6V2F
G3uu54A8Sj/FWT9j10L9NBkXkZ2+yqax79G8tf2BUusl4Any47VrOEPLBT9BhyzI1SrRwonBl/A0
FQILX/5dT9KNlzBMbtCPThsyBK1v+LFqNqT8GBu5Hdky2YiW4GjxyzrziV7g3DQrGJA8TAKhYOGw
lx6YwhWGZprpAUV8qFQth9ftsi5U1NbJnXDlWfkfBsbP/2uIdapxVHRw9vxNUGxu68fR7GvcEpdJ
3a+M7RQbp8+W9Tqp7dzOKZcY5cykVHjeX9tyfNY3ZZbzkesyjyf1NkYo06lCVihsMCcMywzqeiWB
DY4LVo/L/HJmR6fXlaTpsEfzqQWksQPUBhgRJp9WV3OnwBR/4Liy5M6iSYbRtC1TYdnle9HYiX0Q
DGHWqaHL4RJPGT9ikaJLIYRP5RT0R/sT461gxsPcZXdWCideCltu+Is1BYRFg/bD9U3yI7LaLsdl
z46+1Gw+6mPoBMkRbER+jRLN7C14IU66atBPzgjjOU2BGQSjiJ9PrGYtvC553KApadFuisqWimHh
WNvrGYkoqn9GaYNC4kcInznzmXE8AkaAbz7RkZo6R2PYgYhVPLQkaVpRteXdmRIJf0upOT3LAI65
o/J8sqhJiSE0tucL3fF1gU5jjNBEzBwUDs4vvyshYCC9XbEIGV2vuYDkmuamrVyWcCkSPT17RdJQ
+Z79jWtEdbptrqyVnIO9xqGTC3IC46uIVCeJ/mQiJq9SwdTBH0cLPqloo2k5OL/LXwWGQACyJiBV
dYXf69UeCz33kcRuavIsHxCVp32rnBY0N1HcWcrTz8u56eBiiHOGmkaXr6uVBiUrD42D66JqGlIw
1qYf7Ir4r1q2QrMIOZ4EB+toqtX801ECBoyrVk4DMO0xNx/wlaT6QD2Fi4pg+okJ9J7ZjXJOWHHx
8B0FkL734m83yK0bkxCFGhx1Uh/Izy3OtNpPdITMO3biEIlQTRlpS1tiIkK1eIWmQpLQBlYDoaE8
cSeh2dl0ybpDm3OH7+2gsQhB1a0SE1zpsvCHElZW9HvBifYpdEc90xBcR0Qsfh4v4WPG5Foc+u6W
AyqyMGxh+aKp7YYL4HSvzF6V6UwWQ2R5l83nw1YmSPFs6KeMJxWvTaA2NPrEF92JfltxHVoiQVJj
x84za06X+cOFnixbLj80wSjWefaF5ioFRJJaIS4uNBHE5JCHZgVGSF3UxRvQ9InTVtnIfV5T/6PR
HSiYrBeDGB3SUcqGuKk/wrDEKDC8RWjDjbxdR3uH/hOb5vWw0S+4umk7NzwzdzqY3I+uUYW3i8W8
XarPLgHHrUrxMNHIOBADqLTu4UZB9nYrgSEU7AjqJ8C6hzOuLBp61kaoY9Bmg0r6k6gC2rzn2sxu
CgWLCWBfNHAf0rJAvKJfQfXwSWt0bI907HirMAaP6UYXUUL6C+3MDNzNsJVC40RtuMbqmClG9E45
u3sET9ESUsmTuUtRh+WpggzCFYGGD3h30vwXvFu2pt9WZ/1U/0xbxLk4izUKfYvjfdLGdC1WQQeg
J+FOiPJjXc5BOVj+wZgeVzpzSer+LoRB606Mal5H/qetS4nk1lCA+oL0YI04yRh82HGwn/BXX2oS
Ay6KslQOY1G/bAQT5bl+//ldrg8YQl4MNwNasOD6jhBy84ZW2PP6mpnVFv3e2ldsVK3Jmaf4o04K
5DhIIQOhnjszH4+G8QZxARraYQCVPD7ybseFZ5AR9ADKuBSR34GOakOrfCJwW2x3rkRSkyezEXAk
PUAGEz98/2xxGRg5rVj5Pb5KeN9jc3X82QSd/zYbmckBi2+2R2lherVdV2z4H6fMH2n5ajV5V0m3
7zN6Ftnye28FELjPaEB/hsmJ2CGLG72UUMDBFuwT6TY3p+lPFRAi3VxmwxP69A4CN9dKx9E24Ipk
n79T+40OifmOHl2uPkTZrBCA9rB6SLAWSsyFqD07LULwGwB+gLyQrx+hSGXu7zN67fpll72goUAE
7M9mS1cpvbRozDQNpjW1Ha/PrPLtox5zoldzPIPCTlady3KUQ8+4sl/yXm7SWrU8i2/P4mLr9Utc
XJxWwKQ2oU6pvkUf7DNSaqNmo5c3Dl2stzySOP4xm+tiw8/GJ2w/dZUuK88WhZhMqYKax0mMZIPc
rZz/90wArsLrzJLd0LrDvscvwbMbkS5J3K4wPZ7byrmD3d77IB7vFPlaKVZOk0ihGWKBHjJ95j5n
dWcJF4CjlUDMCEm2+2jyB9ngjFByeNkS0xzjGucrO2/lEAQt/AAKa3BYa4ft8A0EkcWHTNJM2U/r
Vu2iMjJjBVLRUHRZBO3i+Bm22NQYbVgtdvV095D4xKgPxJv9U8aTilPk0otPkkSdQy/N9KYDfWUl
2jM5WTA/eQOXhq98NQe9uN2JseLmas9gZrpMoyYgX6xkPuBDJ8UotdaNlNHrZjKf3Svfj8ZnaU+T
oC5veB3XIoNbmbUDG9AqqdDIldxw+q27fOzQEzjgKCFaP8iQa/Xp9XYl9KQBRJLgBMU/5iuZ8Bjf
EZXz48IR959Zrr+awMqHpWcy8Qi+iEoTZ2AEkW3B0lFuaC9Ny3uSKD/jp9fsrXq/nIzAIPiQklKA
JK3JF4rKQB4ozzOj9S03bPbrB+g9l9LUoplkKXOMerM7h9smMQermYwLrKy4OaR3ZsTNLII13mb3
OV3PTrW4utXfvgHTDLN8YTCg4BE7x93l6lCQQvAlqdQnrbRHQ/j2V1X6OnWymfYow+LibZ24RX49
oD2U2zXtSOco9JCHBS2g8MtZX4LPg+9Lhi863F6rPYbA4oYBqV+GXNEBauB0kJzU7HQTe4WGnTUc
lPWRURqIKPS5hwc/pmCaanZXbqxbCOZgSG6Lot4uTUm/Bng5eud5olAMhurV+VJmMYEjO5uXxTDa
ZocBzcg3883kax6dhgIHDGaMT1IOte6RRlbjX9K1n22xnVlJ2JAFjralDhKapDA6jW7gL8OcWdwx
ojG+OM9QpA6epWnMZIgEf4D9p4Z9aN+CgStlnO83RmQjLIiTb2MPwykSbG4SqkXtZ01BufoSYyPn
DJngAts3gl3/KHaj4aqaMQsHYouyp93Mpc/TkO6I2sCMLyT8WVygRVs10HXTJ3br3XIuUdiT+OsD
IQ6+kOqmhmkK7uDhQPqzcaVa8xI0tJjWaYqjtSPmSPJx3R3Z0NRtdCRV3SkZ+DvE/E7Ml4Sb0cLU
S7CyA2gIU8eFYrd0SR8gt31PBNlkmtUE3aGNu9+Jmej9NilmM1D1WZTL9Vmy5ciiFxWfYkX/cOHH
IlIdkpD5F7ZzSxKHpT7Hyjk0TEqFSSdWge7+Kq3PQedrQQaA4NQM0orI/8rds2UsDnp413GwSTUW
wj+SUI9oXk2MIxUZgSIwxaWZuLiIZn9X06lOBWn5D2xuvOzRpul998zXekSDImprF2GTceGUwraV
ZbLvKPPkRy5FGSPHpH7+6HgRbYuwvau1scICGZKZusDpD2sSRVAMNOvGKwl4jexdyFR1qOOmINxP
dE0xNHV2dpQ9b7EZz9gi7I7h5sMTSNzV9FZ+6TNUViY859ntVHUI84YLXgRoLpsPnjXPbc2Qo22r
Al7NyAffz0p6xWwdLjHexMeiISd0yk9bEnPOs5P0RSR+dZvAH0TnlygooXMn53IWO2M6jqS0E3qz
EkB+1Gz1P3ChERsXVG0Ks7Gg4BDuAHI6Od7cQs0/2lNVfBgFJe+SU+at7T+gSs1x36SJ3gnTPSHV
+9CVoWfORt5fl4mYUhA6ev7i/9C5uhmVl2u2+Lu3NcuwiwyPh+CiYKqJrxYSR9w9B5I6Ggh9eJVA
vLGBUCi9VAEfrXLd1a5rtlOPegJYm+F4XEFRXCP34IO3FJw3uNwXG2TYPNPJdFcG2BuDQq93NJ4O
EayqAveynfN5NSEwQc99xHbkUlaypxm3pLxaYY7eeDAb1S0NNkfEXE8frtoxLvr+dLbuzBf9weoa
wgPR04tFeCK4aOvHO4plJbC4qhrE/mThwGmqhOtjmysg1S9mNr5uTYp79E0xm6qRl5gh+pN148SM
n1GA657in5jGfGM/gVbTQT5jJng6dRvsgo0I7DuRf4rJy/p9Kt2gp4DfNPCEtt+Jt8IbX9UZuvkQ
Ip4ICHwRQ3Lu/DrSn2MNgZp+0vSLy3iaIYqlvTvvyOCxPZ2IWtqyGOhMg4zV8sQif/j0yezQr+3u
KU7Ykxrbbrm04WpwjXy7zb6M0eaK0dGhC2DV9Na8LTw53Mv/sfiuvmE7MgeA0Wort0AQUyo0q05h
p2dx3vBYdFJX+G7SFXki3Zc8yB0iXJnuXY29xCxGbI+XcVTbcgeoK5CL944d9z/KPmSXjU2/37Qu
94Zv9OBKxRObWQ8FSWsQDd0wv/+mVHLWqbAxnsvfJLQJmOjAlAoIRWvJ7UtEab5pjDd6Dc7inFZM
n9lcnJ46SY5CZrKvMmsVdzTYeiBvn8WB3uaLmS9KuVTh8zbPWCcLafMps1ReW6a3g+UpimhbMB66
FQxS0b8BK8GHkyG0ypTwXAARLoflufm3aJKVaDhENmEOkernyCn5OeSUpWfojpUY6m4bmK948NaN
XgzOw37Ql9tDyKM8zjyPdvsSiDa9IOdWGxiRWsULtTvWfvu0mXPUCbYBaXXcC7uMrmQQ4/8wDhlx
tAzjMJ6WaFQXNRJaEgRcvIEfPtFlmNoOh4vY+thrnJC3wH9+mt08of1IKEv24zkxgV5s4vMF7IVe
BuuYXazFcn7mfdK810/Z2Ah5CKR/09wMr/ZDzq85uAIv7rrzmr+Pl0p/I7qqP41UYkHhQKuBHYoL
d0vYwxg+arFO5Lihkv4bEh85b1KHdaWk3tvEIxXSLRAGKZniFBiKOmr6/l+wkKKFTc+6FQDB2MU/
NhhKwSdtPH0Js4AxvR8zt5T87iTD7sadTgP3XdRIn+SHRn98eqxDUbTxtMTQ0FigBvNzOaXgr1yo
VBplX9qcZl6W9NgeGgWum8q/iPpMACE3IWMTfYwjocSFVSm0ReJ1w939kWugeSWeiHrmCTe8rRgg
7ZCYaYzTZjVxe3O4Ao1wKJgAic7ZdKwZxlQSbL8NPOOw6kKG+oRXN/hU4j/uEYd1YizGFbC4KrbP
SQjMPwa5xp+7PxmzFf6ryiD356LDMPfZXr6XANjLLTrZ9X0u1SA27azjNeLmDcVkdNUvJBYbjVcf
BJj5Wmt8iAxfNhf5n3yiI8NquXSU1zApvTgVFP1AW4zS6yghWrT20pnsIEaZD6qFdKNrf3MlcfHH
OgDHG4TujQflrXbot+UhdEZrnD+7h0tUweqVW35CwDAHOTReFmXhDp1S75zoFkmH8cj/mxlnIQqd
MD1JCOfq4qnGKZZGkaO8gLnYbUA/Lzd6LNpiPvGczlc9Kxgkq/S1as3BX2GETdx8QRq6Anvcs2xv
ZNdJyrSIYSgwdF+K+kTTV+r9cmqZjqq89eYSxJTweqCHu8YtqywT41/EdpKSWNwSYQ9tZUPwEQUu
IVV1R0IiX6CxLib4HpgZ5mAlVlmG5tye/kt0F7McPM/1EQpkJl+0yWN6rUskbVT2jTO9sNYWKIdt
pErj71ixRDLpMHNPP+jyXLsYSvo8nX9xm9KK1dBf7z1jqoLhYn1UrEWl9PdbdcN+OBybIrV+vpe+
BQpswX15r/yphl1QiS/X1ejQuVkJH8o3D7BedxwytEY4uLi/Q8rl1WH8qcrlBXTAkRN9sWxAwZyX
KKsb1cuPELuDO8B6WKZkPaUad0dNw3SxQ68cFLPEOHqtVFDD/g+mEsGU+rlQVzsYsVqWpWF3qPPM
QMOKyy7lGtR3OT2FhzIRDdcgFdWJgzMrAFRAOkYQdoYzuWmYEnKFWpxYLLe666I66cAjfT0evrpv
j+lGTjb+ZJrCqnM5TEjS7WKxtq/jRq0hM8nejj1X0G96U/3FF3RIENWIkONTuLpPAeKrknrHmVbT
nEDGPytw3DgDYUUbq2gCYz1AsGCtlL0FZxYLuFe6bi/muCzgQDZ/i8DRG2krQXaV2Imb38FaKTSw
zXgtSKW0rdKyhy1T+gyBbKtRAK1wIty47IqWtDIVd3bQ7hBY3b8l/VdPxtPMVvM1ifnaVzZwT9KQ
hwEvKcMLWkHVe4q38QYRYD81fpHG2WKo0e+SezubVcKOBwrcecNhBZ/joQv93j//dv1AwquwEQGJ
SxedqoREvO+PR7IEzBo3MKB6njGVSJXXwkd8dzS/1aAd9JD4xE9urGtXBfrKCTOBuK8l7Q/Ghfks
wLn0kNUTJZ5qMdMC8jn2ep2u7lpi8a8umTGNl3PD6o6p3KQCrQX47AbqwTa9cLXzNTOR/5qPC/FK
Zcn9F8uqbJ/5p9rB9IZgXHxO8c0OgFwEzty421+XXBF89DdABRPt8JLb37SMlLjuaCOZkTOdML2i
iURr07rVxhxAXlKFAqdImt+KH71aaFnjbBxH6yHuS9/YHc//t3cu/K9dotybOgHtIAU0P56iegv+
mhFxSJXDoly8JIohXx2rRI8UB+vxe8g0WLV2AFjXGtPUNPluftfDrrwtbGTOIcgg0zBzNQUBkXDb
pXARsdcOqABRVtBeLgpuoMKPWcEFD2h7VqsgaWEHquHKEkW46Yl1SJtFBvDUM72K+ttx0Dtn7SKo
UEiiNovICMqZ4dxYUMHjf55KqTilfNne7jZpXYe7LyrMvzoQ7HP8qmjadnrfeSlbEhrfHlB9pxaY
P8vwWOYHN6K8EGu14vZx8NTI4Hcglta7tMMgfc6Kjuz1joba6AWnYjE8L65QaE8wGBajk5gvSwqn
ZlYSvZnoQ7Wjnxt/qS4cFZleSDuJ+uUOUnQLjlIuU7yQ4PNnGgHSk2gYTj8T8lmWyAGywVKTEXVD
Iti8JAlVnHm/XR//y4TiMpvLKcrX2Cle28brUs1nHSebEKf0hKzdgJKjlRmWu5FQyBP2IRGlDqK9
dY/MQlQhGTiTYvyu6TE4/G2NVvUFYX5BYleOEPsA4/P/tNLR5zd9fl8ppG9DHdcb16jy/qBFMJG+
NxjqtRoCI/myKG6xP92f96pZejwBE7N5/5Eq77xNk4JDA5L+d3jUtlhlSN6cYWrcOWrvhfwxw520
c1RwQU7sZTS0h93Ep4b7VuMfFjxQaqHWrIpzvKFIHQNmRYScvOMyKmROBdscvgO9Bahe+DAC0BqT
bqkK0gg0xI0kN+CULjnHusEpisM3r1kwWMt111dr8bspw+r/M1vnl2OSbD56taEFtFwrag+IbpXJ
vTBdViNkWxn8zHlgJNzKAlsCZRdOUqnBeHdGxPCA85AdNLU9FIvtFzxn/U2XhVYNb/4WSakSOAOP
GhbvXv2o0og7FScPkP3iMa9BRkzNHDF7yyzIDlCRO+IQdvPdRxvPRkLEDakzDXK7zNgLjySSTdPg
I/EZ7puaWFAttNaBOK1XCt6bGpCF6CuIO/j9EciUqaAA9GHZtLxDkSHKfew7nhqUPgPHvQwDvMq1
fym/+hePOTHdKwOr4zd1Dt+dOaIt+hoqbYHJ5AQFSgOE7e0bvAh5plcGsbA0/yR+QkNdpk479KDU
EIPewGpz2SmDGTfe9c1G1vb3X0UKdMy4KkIODBV7NJydz/cOEM88pvSU7uEu4NSu68ktERWSz+UT
wepygLdiNFQvr5qYqyS2oWjIq/K2atTwVAaUeABIgFCYqpCNsSo8By6wvcR/O6Ol4xPbPzFdbYOK
FbDvOL7IsGK36v5cmC2SOaL7lITSK0/8xmjiQq2m0LwIVMOfvugNuOvc4NDuEHg/3uO6pQGo4bCZ
HEpZIFwX1pikeEcnVnBPQTwBtb+Zm+6c/+YdwuXXuCenAxoYAQPMUjyoqjPgQqQSrSHZC6YokhLf
HCmCJsD6PgtjsaTGSqFFMDg8SLYFHiEAi+bJpXbrEFcDWLNpCYrliJrprKtdBUz8Xv9zgqexpxUl
n9RKI+HJn1HIf9jcghtJocwxRNrTO7HiN9zX4CBAdgnEZo08YmCfDWzo0m2/MJOq6xgPi8N0qno8
OGBjKrtk+VXl0UOf7jY1aSJmbgE6G/Jg9BWvaXG1ggpVFfqNre5Q8O9Et9tS/PTfACXbP3xjAfis
l5Q+AY96V9NbOU4ehKkF9szE+VHHNgtkhA41MKIHC8BMGnP9eA8u9lXfR1kQGfIMWxG++G0AECPH
5vg257PJKlrI1VAP1UQFJDEKUu1G5b+JSeUwdpOJm9UWFgOAXOyMMeiXMQhVQUA3xrWXA/MqioV0
dDBcxb7w9AVhp/I2ffxfhwfyH2w3NEUzZjdPuOZtBJbE1b6Jb0C5tMSvoY1JAy0zQ+6D3FGMNWHR
lDWvzSsilUoY3b9cuZCrrdB20MdkpaQonc9rk8xOt8Sfb2U2FebZKUnn48qRTtO++AL561tJY5Bd
m4BTtS5qsv+NN8aOvvBNVMsem+cBIoa1+vxwxnbuqtZggeXspHA2bOan3253VFUJ/wx83TDM9R44
n8O0CCY9qjN/IYXc7s6flqvFsd9FeJExLvr9ojyMTSe5A8kzuyEXeelqrYDf5B6gN/Wew7lzc1vm
V/EHsE2TELMt9lmSkB2VXa9VzsLfFHU58aG41a7Ay/lNn8yxMVdfBw6kiVBYKNKAdPlQj6wUn1Mf
ZCSbMl+G3kuGeLXg+I3SVoJimFxnL7QGZ9VoQ6xHrRoHEh3K4BcBVMcFLQoCLC8SG4ZhycKGO+Et
oebvxGPllQkybGZSfGpK66sdeshqbjIp0jATezeIQbt6OGnq/IZyjxQbilTWYvRtnU8MeKW9cbGN
n4sBufHqiTvb3xan9nDQ71ezWd1eELAls24oG+wY40bu91GX7wRtgyd7E36SxrTMn/jJ2DXtE1FB
aKR13JFGvGhjSEaWHbzA1EBuovpyQr2AESCGT/2OCUhmimt60T05luTibNW7kIme9SXO++2Nxq36
iKr8ZeKitHNjA+eusROCWNarQRXKZ8dF4gXaCiTAuAC9UNNDZvTTJJRA9UeZmKlaf6E4nCm+5cET
Ob8HWkXwhPcpGZOQvRGM7q+X2ikqHeYFYk9yndC2XSVo42sSLqO58XgCl5opoyJ9S81Iq3lq/lFi
ZE/ijbMU6Iprz2qnLgeZwPPTYlJOCulcyB+IiSAabZdTG6lMElKdwzmdJbXoUX9poUNw8L6dZXaG
v8rB0VkZn1oMA9KsoKD5AQsJMnlAPluLcxl766vtGB5ewI8NvazmnQ2IkPwyslwLDQyT3fKrTJDQ
5a/3XjHLuJKeeOkLFEFirUc6wbFc5hvSU9Rz6dmLLUMIc79OA4lByMOOOPo1lPmu7oOX1WXM30qs
zRAFnzBaTOVytgvYXFNNqew9fH+YWUDjVlfWjgQSj5NJcceXLvQjpPpvvnWweWKeNNGFZllTqIXF
89FRzoWxuwE1W6U2otTxAC1vvd2rwBU9VKioLRVj7/+h/eqGth1XEdcHRIg2TFM60i23NM/LkN7O
l+TFhDxxCKUlYzsmsTnGrgv9ArtWm1BOfUPSIb2bfYFCpfTpW+eZsmG2CeUrHnNWpHbdwwTw85kd
BU7s31B4dPHYdKnAUf4aw6hxFgKVIOxOMj609jWIpm6rEq+fPMGgbMeu+Vo+oATB6do1zIfUVkoc
ZFbPoJL92101WHylVzh/ZN7iOPS9lZEunGKrsjPsOBrglc412V+9Uv6BxP9He1xDNqa4XEbBk7iz
KAHLbV5EHEMxVlka6zmhQkKerbuL865LqUop9/gwPSa8MADFg/S8PfuQk3LnIxGPLvVWHrCKxwCV
2Nsxsef9SzIQWEpkMa24sCM+5Id74GPZ74d8Dw8ELfYzYKffBqgi0Z3mElpgvv7SagB0L+UCgI3F
ocjbZSiTgYd0AgibpwMg3MkxJ6Fkjzrm6g4teT/yzQXxqi2QSZKT1jY6roW04AP0cpsYtkoEX7ld
SuXVdjLh3e3jXdIW8k//zdZNj/y9WFcK9FEZIfioR8w3GnzmIwC1JTJ919wSuu+/t6FccMRRvW6o
ThI8RH8Av2iID33NrHutgvlyHPHY99GBPWN8YQKCOC8iZ1gQAvXVkZYk5yiIbNr3QtEtaH5wZVgJ
qeLI6T5Pp66W+C1aNPfD34G/teTvnxbsZZARUpMZpDCHcogyAZkUOzgADvEThqj52/ubE20xCj8g
x+xQuBDi7peTjgsiEOvyv3RBMmSS/b5+pBI4uu0QBIFUhQYZrh+iHItgJjPWlozcxn1h6gK8vMNe
oOeejkxH1qPW4K1d/AEqumQOAYj6+78n/a49iRQjY7P032Qiw/bb4xni50NnIJ6Fj/IEbc66IKPw
tzhK0q1jTGVcCtJUztD+c08SWuqS47+eem7zsZc47d1p8JeaVSwDd/cavOOWXs3cxlVZTDUMXxk0
IvFFelNE2qX0wB9n3ST4Nizky7eftqb9ghvI5Dz3wXU87hvxLwjuW4UsQhzVlTA55VIExFdz3FyC
gZUVoWbxGLCiHYldDyzZIBrYQc8uTiLANNk0UzNFoaVoxvlUo4anfwbtOBBmLuAJELoJPsUIEHxt
s5XZeE/+Mob08Tt6LgwM/KDTHl6B0hklzhBKUwVPVJRzrfqxiRcbpV1NW2/5muD04jELJFL1WWHv
VxIzjyVP7aWzCYtRQjYltT65Bsx/NL15DSo+FwmsSHm9g8R/4CtERUc9SjCce5WC652CWfK0AFn/
TMYgOddo+cROYq0+HT6+N/MJuDRJyvQaAMCLmsWo9wdTWOg4MN3CfUJehgAVWbueWzqCm0oabQJs
JZ/m8LrdAMEcxa7WENbRbZ84ePa/jFYbfRjGvAYIqPBdS82lD38m80hMVPsZDt1DqzZZWqpLX8uP
vBZcPgna5iQYoDk/HbWV9NY4spzHpnClaDMb6VZb38Zbwc9IX6zjDa/ET+kbGpSm4TlayNAgO9Yc
YO62mf6E4aiZ0wJhFvAttr0qcWYgIRrjkr7dUaYEs5Bg34NxfFJfrG+PWKEeBdKQqiWUcnncn1R6
3B2GtfcopmTQEBxFLw1V/YtiCKz77bggZ2s9RnqtZ1OAWt6Jdxax3GkV7poFqiBr5yz7vzqmfxlx
pvgt2L5Mimtc6HnIugD3Jr831Bd5w1ZxOu6tZIzZB7AzQMmF4xTPrOXZkYUmuVHm37inoepu0Hps
7zv7NwZqmkHm/bZPST6wKp/DEa+x8nBswF+G/95/flORBTEVESPS07fZJ5KO/N2ER90XDC3VeA6D
qNMgs4rdd9vPP+jYCJudk2Ey48IxJDWLYOzP08VPgRsrsCzP8FoBnTYb1W5ysy+u4Ujc88CW/XE3
r1QGyKkuBNW6LyznhHdd/o3UHA1BTzyYAAKPm1JsZVwPMlUba679GgTFu64kLJeLldl0/TVNjv+M
Ss1h8keNDHZpVr+ZWEZzxwl9PnrPabtyCLkP1JJxpq4wj3Xh7YdPsRkxp531dPUjLZ2TJIpN+uYL
vTJU6bLQ/J+AwLO1o5HnPUUVU4+xpUE0WYhj2yHiBt5m52vH1UpQrR1XTH9/8aBPFm0OTT8E8MId
OlziiSNOFQ0s1keuHTZqwoGlX65K5cOHqMDL7E9i5nqp/LEY1v6ff05GZmDdcRAAveALKwsmhUGj
3Pg0AhR8be2AAeHiELJV57rBsi5kUN2fQR0hebIuWdoSVpYSutZ7wCaxD+ZQjTWbP6wuz47MZuRM
Bs5w93vSSaBCqXOEYGlEZANz+VhcHusj+N74YnbX7Pw8pEZqzJXPUp0j4pLk1B7fjoHWOL2jRaPT
Fs1n/xh7UDVgfk/KL2i+uB/vBpvV40z5b5cNDJnbj63pmTn4JVZmXl3oDkhlqQoMobAvF2QCAWOA
fJ9C25GZ4Q+MC29628Px0RPGaJ9eqKvEWkpO+lt1nD3De76ZP4acHDX/PCl69C2tMP4jnA9qq6Kr
DGLd2Wde0KwXFuxNbLsd9lyDxqu09vWEzk54xNvj0NWVXP34ee6Fhg//ok4fVKdOzWnHjW32m9VJ
yIVI3/LWRG+DzLlfGuTv6TmcllCSmeER53Z5MNZYTe1MxlfZv07uCFHRYL1iLOmwNTYa55SrODps
kf1qlAsqfAfZTHhf3XYuoHx0aCZ8P0GzxEuh60kSMyUbwGV2xoO5SU2wc03d9oPNarzUFuTHalFH
ZymN0fLLdJYKnSPfk/1pBRYAVbU+8qr1bVfoxgN9BUAIN3VIR5N7baL8MPcuAZlY82xkshBQEm7t
02nl81nqOlNCO0j62Zd0pKhCEYsiokejqyWrMPFLNTZ9PPv9NDO6YeKGaU0jfEtqYOt/WAZ3EIhf
aOSOnfwVI3ISE+uhCpN1nAZQ5bNCPPspP6LGh9VHnAgM6oIol0Bz14mBzmzVdpDWxEaK09eSygP5
vJv6P4Dt0iBBWaPW9iPkOKkZQTy03SsgXN3iNvLqikllXyVoIqEaeAt+6OlHSFdblOKjqLn+6X35
/xnL1H+0OAOqzkCtbiwjdxnUMkI4vcQN5icK/2SAsHQ4APQuV3rn7AYbHh/2L0faJnZyrBGSDhNX
woJw7+zdktmH7Fa7bJQswus38sznKKjM51wn2lrMTHXxlmQwhtjkRDTYGx3h46d9SvRRjj4MWI5e
qWKRvFxLOhvL4OOHCuOkFJRaJ6OYEePYLJ8b+2eHO1QDSKUAsnFcuwoFV8umHs5gOHjZplqVcJzG
rk2CKJetjPA/fupOcfWulN2FahgmLmWxNdIfID2W5hin5eqD1M7yE4XqSIZazWNdkUAQ1sM0ceE7
lX5eNbmjJZUWaAmlep9NZetf/gMBwg6IrCKLVFpqYGEPkRBfNFnPbTU+n8ZU8Cja/q9HvT7Cz4nP
bEHN9N6NK3GZWmxengb9urqt7EFu6vRM9qjHwzLb5UvNFHHXn3QoE0t721wlcWKyrP6Hf3O3QLat
AkeYUq/4oI3kgBIt7qSLnaWolEPSG0Knj0nqC7aMnt650E8HEGUEOeFGd6lJq0JUu+aqUeAANQZ9
Z/Xb5XtSTGHhgmh1d3Zu+qQwavH6TrN6PYYrA6A22eLvm9VlrwcEhFICIX/CC9eKnDWM35gxJgya
xmc3ofKVYUyUrcjU25JYS7A1OcQYtM2CSc3F8++W3Uvhbr6bagmKOJnHC4Pf0L9xtZojNLG5BMjr
UreI+XUG4Xp8HSFa/DbAzgFNdvohAhL+NC/4pp2FMmY4Qp3+aFPQr8i6Nh/moSvczhaEpAJAhVGG
uOyiowILlRmaLo9lwATVhMGYdiRrIxMLgnoeYjIazSTdst+TvAikBuK6JakaNDv90tgir4Hqzbhz
oZxEvkBrW7SNkZKEovcQ1RrsOFScPZgJ+6CPxN6TbMPLWUL0bd/UGfioij+xzAiKvCCYGBoLtN2s
9xK47wdr/UuPLVGkWZ54YFNEcS6B8X1ZaYhF/CL4UfFbKfsB0Miwr5zdxDi9k2sI85APBH1Wr0lr
rTL7UnYrnvDbulyag5xKANJ4JEP+MzB24RrbFqWXhS35w8eez3LzASVolxbfWXDPHOz90EL7ZuVJ
AUvf6p4sEzaQ6GNIHtfMr1OAxa/sYCWYGLAwqkT0I8xy6Rm5dHuDMkTTlW2vB9Uh9xIszF6SBYT2
14SQHqH6CPiGr5wjyd+a6i/YyZNOzHSLTnPwQQg2QQtU7J9FXf7CCMinV00FlB3v7HpYoc8CpY5B
qJ4aEysB9mnkX90+gTx/sJ0myUzs4CrGjAnZVNf548gkN1NLJ3bNRL6OZSxHHVaX6DAqOufKe/0+
LiZ1nZW9FQiXdLYZWmqtr58wAHl8pLn2/nfPT2K+PoTwWm+y8z8nUA0BxbTw2VDd8QoMN2jKGfg/
GtbqFXFk52kdbjZuscFIPlUxi7whfXxsilbHiZV2pLvWCM20ebw6c1SngwY6AP0qfcSCh1fkhTIB
9ogmVseF1SQJyJVY2Io2kErhI5ZL/UZFnbLi5OnXFt9ogRL65znj9HPa+FXQQwHxLZAScvy/YFDq
Am2IvJalhdlo+fA9P0FgERvSsR/5y4s+xJ6XVLa0iYXPz1yN4uI0sKjt8b0GJm3pte5tJjk8e8S2
5vOxuIjotuqOc71c2bFuvNqphwQE+jmFAOXKIJpKD0j/2epTL02ZYa2WcJkohsv5UWc3uSjggvAv
Z1Yt8UUU9dKpZvex7FOxEP/egPiSz8oszmYPW+g1S60Ixiji5ZsaV1yIOCdBWa260ulzgBW4RL+B
HzTVyY5u+9yK1fluptzjLpgc5PSOHm39BEdjF0A/bx+HCiXXXAGdxYVFFfpakH/InMUEIgY/deXx
o+KeEIaVt/E00uMyARGm72XOdIbsXwDORyO6ofwlopuy2sMPTl1/SQPuKsOL7VjqcFO/1CevWSWK
Xurj4kISVmJz5G/twPwzugw/9G4wf3CU97tEXhZSseZ8fUUlsAEJwiyvdlqONOmX3FUj3ud0XUaV
9XWmgQQyITZ7/HkAIF6jjCdDx2whb8kLNgAKqxHcXkQIlZ/6DZ3oRPk23Hz2QC/KTT/pploIYlJ4
8eFIu27yVgl2N7w29T7CGZ1R1g3qXbd0FGpPQGlHwbooMgNyVKYzTn1AWujAtnZgnynfJU55uplz
Xs2z9PLSYN5me8myEF8NMTnir1wngyzsKR9sv4hygZONB/Ev/07/OP+QAiaN4+gcSBuJFRekJZYR
JR2d+4+piYMXblxJ7bBbh6lfcKMw2gUZo+tzFvDp2vi4Kvvz1iRSXToVdpw+vFWKKSLV79MGzphS
ONZw8WKIeyFOrMF2e+lrcX7r5c/wJQBc7w3j3ISaVKXixp/5LVeK5Z3veqzg/ZEFBvZTuzUEQCuI
lBS8iIyJNYhCEMRNCfnwn0xPB2QRTiAO5RAgkpsRCvM7WcR96sMEFbV06QqOkjGdUAQy/yxCfsXj
Rn8aPZB+HUUcjVvdUHGWfu64IckdrMiweYW2OnOtnsfojLllBT9GJ4H2+4F1CZ4kwG6u+NworojD
jB25uKTn9xGhVFwUEziDUK+w2y6PNFnvhy7DBu0TsdFjrn0LIVviu5da/KQtDeY0jpCy414Bqhk4
fdGlwJPE2o55EDK05ttpf+YvPaJsOs3uNq9d0oL2nQyvVYJSjfu0zDsn44dtV6YYy/6CkM8SZfTv
t6Ywr5mdIaq05iLexmvDxqkNWc7YUB2kil5K/2ek3CXlDputIdaJyaJKqBx3qf8Ru1Qk1WcYV5ag
BvH7cxhZCbYBGHdLVaCDRIFIwMOk+v9HfUc9I4klI4aWmJjI1hJencIvQY+WkQ8VnXdX147GxIEn
obYGaOr7n2LlWYUUtH5uSwLuEPTIDByAeGmO+/pvhF9L/vPh1Uok8Ff+K+iY9GbqENewLJuzS4BU
hCfzpDvrvJeJS7WzM+aw7nCffvlCeTY+yTlmgKMizTQN/Zm3huab0HmkLrd+cnaQwCl5PebQc/OT
Vt7P3i4du/osyD9xINRF7t+wDpFZ/K6fb6XI/EVSMAuqvy6f6JfhLKdrtfXpjmtel5ue0uhP0Tdh
E9GFYqL8s7BCLUwLBSe5Cvz4eCK6U+TqgJC1BqEXZZUoYKUSUX2nYjLQ44qvROm+2NBOZS6ZuuzC
h7ljQotdj1eiIle5NIeQV+VhlFYyX2hRoLodjdKKVK2Lj/ri8qwb9uz0zTM8tCidI0KdB46g204x
RLTgq3tP4ZUGmb56grr5xBeDEvvouRYGVlk2E4yjS5azwmM/vHcpFkVQo+Ia/VmazK2JMQ1+XtjD
HYZDJRLyQKGGeRdAmZ/2A/ll5b+OSxxWIb3HAnIra3Xqvd/JOGVRALr5LbXQUFmH77JIIOTjl66n
m2VuwO8pvDFVm8ALwxoFWD+9OYG+N4bvAs4Fi7WbfX82YpG4pWKrtdQT1NMA3KZpj7WgU7ONOILI
itE8atIDktTi31LRcZmU662dnQgOp0BCATZCXMPdKBwAAkAcGxTdQkyv4UnaL5OOpUv2KVMi/cSg
tf5/1PKDvF0SvudoUVtNo/Uz3KTlkFpmgV/mkzRoX+T4cAC86PbeZ41a3euNc2/yF1w2M26e/S/U
jJ0IC7s2ZPTPQR7W+fB9BzUj5IFjMt0OuXkbxvnHVzmTOVmCFSt/qbVIZJy37Auaf0OMVVxlhq/M
luHM6TLU2wk+63pnz28L6yqKauEeVFTU4sSid+ULSwJ6epGb5u2ropuLEh8Fa8DRo+d/r1WbidaB
n0wZ+a7q2TGxspIwFSd30QZthmJ6rJnvzVdvwvdh6ujhX7WZ3mQZ38zHBsIdXT92RIegJj+bJgOp
xNhb96NE47fdZVjKs65+5hC9aigdiFLkzlRijGSdax4yv+TItffaVGZVs2LQBmEa56Yc2+rYzeMX
xawqa1QEqG3XA/1gUhVkqbdoAULPOegkL1uxKw48Rx97mLyrqKq1Bvj3Y7poCO2goN+WqS5NbREY
HndpSW0QyNHE9stETmG9onkWKMDmUW5rviHWKwSNp6JjRzOKIodJXhbPBAystbYXc7BopfrLUAF/
4YXL/vF8W00MYgVHrELhh0zWFaKNhHgMST7dNNIWpn4GzzuFEPJoGsn/tK4O7kyoQQVnqtPNvmBZ
DuDeNoZY1dIRD96rB/GSreBVuKO4V6ecB8p4FgGiK8lRvo+fySYnA41WVxE3DHROiGywYZVWF5fU
/I0Z/rXp+0MOEV7BGtp9zMOFsg47/DaBsUJFbSuDKs72eeblQxK3RbXaxcbUSfPs7+0wh+ZkPq6T
Gf//xzRdahTBbqDYzALwX1yAvEZCE2rWmu805rt2hF4xZfUMhnj6YXHXx2bteUkQDp0qFsg9hyCp
yHoXlc94CDrkRFpimXog8vlBvhjdVZWQy9orVdV1D1SyA9xoAMPPRJ4R+Oy5Kk16OlTJLqON83CI
iz3WxWMndrvj5iPoI7rjHb+RX2yUMfpM9+/dgjJq2y9PDxcCyXUu0Z78ridoXcWNc1g8J5FWb3fz
h+TeEImMj2YF8A9Y8K6EJPrN7+NjFXummKjjo+h1jHKMzJrJgJ/O70KuSIX/UygHaR0bSx9I5QEb
wtKEAbuH/e+4PH7L419x8qdcnB5N7/0H9hd2ZdTITg2AjksY4BiDpOpaeQRUNd0ev0m5liOq7GZE
TfUQIyI/Z+KEF1wI8WdomD5bgYMKa3gBnicWTUi9UflVgzFUCOj5c0nEFMuHDoLqkRyiH2LanSJn
dizMrXRGGB46elDY/cNlzNA/SwZVFOsuTRcyg+0S2UivdEH2o22M1DfUCLY2H8J0oKMQCv3uhViE
XFVDbGvZsJB/BhQWpkXMdHE9lw7MGArhCIiVm/Tz02QQhEOBjChmWLLJ8QcqfOsOKrVFhJrS94j2
rKTK+uCskkocJ1/r8XEFvC3wsDi4mHG1PcZEFCnfmfhTrrX/Ex/6LUZ1RMdoK7kMyiT1jvclyt8X
Xmm2ok+hPPXxbL2frvaCkyEDRz5v23+BHXApfOkHktIXdGIcfjp9rD852frAWpQMdYkDK0TNK3Iq
SCrCOKpsqnChxi0skFAbNLnVyvzQaxD3Utfopyyc52jO82+5oZpj9qN5JLwUOVN3x9q8DMp9qYk2
yzudb49P1ydk9D2ckkZ4qcgw+96JM2s0ZzMT9+McPurRqxJN4eGpvXkyhIgGbd7PQtqpqfASWWPq
QWR7eQSDfrnsLSvPyE0jnBvnCuL/gJC1yrOkfhfOJpnY42MHwUKmn0f8bHpyspnwjEa8bBrwHnwd
QmEeSdn8etl64hjZEtzOFTUycbssFuAxMs10pNsvCG4Yq1OlL5s96a/fDXkclp9LToZ5F6qO9tzS
aIEwzvTYdNfSJ7ySG5m/h2pi+uQV7+y+frwyJkUV7wylAgYbFkYdyWituUsyOR2fa8XeE6VFSdh6
qJ//aE57MCmBrjgt0CiwTjg4tundlWb3bxhue0sA5tTHiFR4l030MbKh/O3HR63TyT6/QUPH3VGp
GaY7V0hjfY+h18EuSTmLoGUiyjDWHCaXEB6SxxQYX2BCcG89C+iCX4z8/IKdySox/LRJyOnxG30k
aD+Vx40M5Uc4eM/A9KbkBpA924ouqJKS1lUnu+hCs+fkCSyXfvgjbukljq92xNn38ivoN5PT3bRn
rcyS49ZWomPu9kevt8ciM26wtMJte0qQ9jLYocr1coqon5CCpl0FewNAStm78sz0JAoaozCciPUw
IeJxyvV9zgnr6eGb+NJyXMwmAUZn+JJTY730bF2PqQq7Shv8kglvTnRpKueuQOk2YzOYjC39zN0w
1h4ROHvyIO1T3yNNgT4UsbSnvucv8oHqn7jNzBV8jqlJ6d5DsvTSS4qK8ixhwde/O8oB12XznBvz
FCpqrbnhbDq+LCMwHJKIsPXleoBRpwMV5cvIJNjSIq5iO/nRjlL8yRBP10xGKVCevp2x0GlDrf64
I81VuCsQVB6e6/4tvIC1pyyh+pnItJqvBpaemw3+8Tw8LmC6gDtsDybtbWNqEZ1czb0FpRMTp4LL
azBEsfdOQIyaRhi84pox/MfAB+e7CJ+tyGsDWR73wB1qexEdOp/h6NPekZUAfFGUwcm4+ACC1CIU
mtp7Q73Ey+brkl/Ylsy8XP5esFTX8pADtY6gobhxstTfbXXTGN8SES7pSsBcDjA8lnRQRL+37UMq
9oiZJ1IV4wx9JSahXUPT0helvd7UuQN+CgKwjrdOeAP3QLqosAveoLtwnaiB0wqrd88n7Z/m4Vom
lXhulbqwGIb5TcU9b3y3zivKihmqT9e4e4MJt/2oFXSwJcuERjH3omPYvArfCt7GMm2pHKDFOz1w
it01o/TgROtG9GL1OfH4T8UNRoPGTNU/44/TF6aWl3DplYZziN4t7ZbnPt8uFfkeM73m5CszExLW
Zy9M50AFJnb8YATcWN2guBh4SOfykzy9bYhVPg/vlllt/JgOlL+HQ1bpOsq4fjc72dvKnWp366q3
WeY1Dx67D4mKgWeHJK8uJwtyl8fzBVTnQXeDj4mbeLJ9Vxi1yGjQ3JnDNMv0v7q5DxnUCCVdMLhP
FhJ2J/Zh3RAqN4iQvaDO057Lv+7jIln9+1pHcQhE1ACGx+AmMdlUuyZDsnEOkPEuPEX6lERuHkJH
Og7omKrwxx3PerWx+r+YS5+uMvb1XbqRX7l5TDrXYT6RDq1ZU5xYvjfDcGI6TcDGyagUAPNVHva2
h+ntc4d50cj/SChx8SiSa0lT6eZ1U50S3LhEvER+F+B6SK5hulWTbv06gEyBCG+qNPtRyqrNvowt
JHVeCky4M7g+SpAB7e9dLvhaQaHIiFiL9XcPfTTyA7fBp+vemniCflUJyDmLGakVyqAKaSwOOiZs
BhgC5V5aOG2ZM3WuLY9g+a9wYiFIukUwgic88XvyU6sSItuvxzt8zklbvtKEtF/77Jx128molFnK
GZGMC+ynvCivW6UaXggac78NXtSzwDzcUitc5Qu/0zgjFF/gW2ITGBj4Q8W3ci7kY+HhR0YGALVx
zrqdT+BLxEGHnRqfXLyovOiOQkmgAGrHx9FcDuMC+esxK34ukX7Phe01ESRr5+2Rj7RvRjZfT/xL
+m7A+FRjUoyJfbUmctiv6E4/fkMoiV6rWcNT7dMHPnzQ33/A7drcCgYLqyXcQDtnG8dfPv9TM5Wh
jT8+mqG4J0w85sfN2CrvomLQOW1RqM3TnCi1KzkJpfPZzr0qFWkEsWMt0FPvb0nGbXkYmutaKgla
qF4KC2OFOn2Rp5+TRZQdjcTNPkNSGy+d6ycBC1GNxJV0Q26hqP9E+WglPS/r/OsQJukQyuNNuDap
hVeNrpLZgnrTBOrsCjsDa/htVdkHfRUR64aEK+t7IKEiSzJS9zP/NSywRjWOu6sFcHuqLdJvIqrs
NvdFKvRYMBnIhZ0BVxx6NGrgFBUEWKd2vBVPtAxtAQzfi9Lzg0/tl+dd820A10MnYRYz3TniRCQX
h2hRj9QwGnlkbI0pxmIAkGahgruudfihlsYVwxgABkadEcXNctLsOcTFeQD8nDcJf7QIzTBCECxn
Ir9Zv+rBMz/1LL+OmsPhAeoSNutNmrFTzvQ9SC9a6K4lGkIt8Y0UqLoZMXWGfo8R4DXu2NDCCo24
VRo3JQRSPPjVp1OhLxA0dL0XldcNMLo0p2oaVm0sFWPc6C0XSUP1rk45jza8FygfPxQu4+I51cP+
QYLwLI+KsuRp5nyhGOgse94xasqF5HVEVc95rak2+x3b14Jne+nPu6NYI+CanZtVe3FHaHYdD0qt
nqFF1luPxas5JEiQtumtvO7KwSBnYPp/NTElYATFd2wq3oGPMcsBZaXceajtY6MD8F1aHzUk/N4a
pYjDNJZ4/AGl9okqHLSuvwrh3W6DsnMaN2CmPH/OW0Vt26H5Eos8KI1dHLZ2aVqpc7XUOwPUveV2
hYNDvYVmsOSJVIyu2OUtTgMqxDtkiFeP6x+DV0GFw7vJ8uP3jfZRQUjVqZvffN8tiMRmSLNcNcVy
l0AkCGXB5luUTl4tUGqoX3OWBZsNpm8cQe0cCWJqIzn+Dy0aiauWv6DiNCwZ0o9bW0qo0e4YGwoi
1otoEI+JNZLcKu+jb7iHRkSc2CC79/f7epihTxbVq5mxuMCzmQgS8L13+GUcJukkYpQHNECsLdQc
WwVv1B9dvDJkkT63Z7pQM21eZKcmg2bB8J/Oi7H7ALV1joSX//2uLnYPujzw/w+nxzZ2FNqjTAMO
K9pUE/HLtUFFSCB5rMjnxkvwwhn4Q6fcs0ptXSJrzq2TfPPzSAsSCg7VNHTCVIa9Xu/EcCrLkqsV
tuRpPfGgZ9juO7aPDolZMJOEWLYIlZM1OHx+J29+h1ag3ZEI3G0G/cnkd9VA0FTwtJVgaLzpAAuz
DvlTp3aLRx6nm4cv+scXEn2TFrazbNqwCDWLu/TmN+Yq/GfvQ0WvrO2jV1DZUc4bUTgJgB36h0Wh
bmNKf0R6fVajTfW1oI5DDIn6cGHgAZZvsORamxHNMODqPx8An+xn2hD7rAhc2pSHWE55VA4/LsoQ
vuPJy1rKxADpOMU/wVqr7tFpKLPHYmyaQi2hPtpnJ9iQqGhBkJAA/rgplDMUqWLk/Zdho/c/mzxI
oHcLEhLARyhNbRhlxCAqybokc/zNbK4bSq90YZ/Z0kwQNGMHvBDnLMidFa+nSx7KUSLRvUy5xD6T
j0OCJh99tI8BH+e/J3SrnCGGyIBFkYMEBepO71/pkP5bb5b1+cG1q5Br1CAA7du9ldjZBqFOl2Qy
RuR02Rapcc1lJNXfaTHORAR6nbedvBy6xZUw9YPqyDZc2C/xNTenOEvpAxMnv3KDj7cA3cIu6zWC
hMVU+WxNB/5qOxkctRuSNM/p7ta5q8ZTF0jlsgyy0NtN7TqMS34+cLKnT/+RShJb2TjfRIJqKlCb
A3pJIDQOvOcrlUg/ogGqv2oMSe0VPmqjnwJJFnBMQeEHvm3YgvZTw74T0IRxswYCefkB4oHqLI6s
rmTB4lJwnhYcaCxxrbG0QYszUreyEjrYWTSaAzbWbAbSFDd2mrOuS1Dhulzq5h1z3HblC6TxIl7F
YvOHuT95r7JMKNoUdgGRhn3h8/x6Dc1LUauTF4tReGn7B6JtGNjyjQiNMaZ4M1ybcuGix8p535f1
6kvqGArG9tW+7PlkSt9yv/RiEaYreQi3/wFENIFWDiLYGhIozyvqTDWpH0yhphyLkJ/Bv8adKzPy
bF1YzI95Uw0gtqCTR1WZrDFcY+oZ9fJZFQJM11/xrp42wX9lFSbPCk9essdWlng1DnMvf4IUtdAm
6y+BEVOmw1i70+PHuwwDt8q0qSsn4jj0gJBXMKfrahGkgwAG9mzr2p6SzuwjX+T2oO9H7Ejho6wT
Tf5ypeECsI/d1LozOEdxW/xo4VXkspZ+acn02vLrGo8bUr5+5o1XX2lWhFIszU8477bJ2uHy7Pea
zol8aLO9Ofm8SosxGiekUb5LvsTBgskKUDK8hefWBYvIyS/foGrBnfuT6jJGw5U0AhP4wQbG/FgU
w0wu27ZFczgSolhgs67TIyE8AuHl/zUqhvh+Z/sgnZD9/iN6n9UOcG616pki+dIydLt6xdk8aBa6
QbU79pMIVlkbV8aikZoBndx7ILXcNYJ1vJ8j7DAwQmmXldYKriVxbBCJQcpV5alh+a6tZlZYnK7k
dVcZd/wl1mZaHNyBpgfC7xsFMrAArskuAsZyEkSdqz9e+XG0GXUn9mOa3I1VR3BPmt+WXnoDyKQ8
aQtjjfI0ln7Ob4ZmkANVIefrQmsIdyCfdj3HA62DiKRNET6L1zR1JfmDWi05SLeAW9/Ajh+7Vfl/
VopQRO4NoSTU/DRQsQR7LdqybBcVDnzQAy4XC2NsZzzhQoQfq3hCfvHx6WyyvQ7VaHnmmtEL6mY9
Gnb4zW+oCZGEzTpW37SKu/I03Rqc4LRRCxYKX/bviQvM9ycav4TYpIxRPrr2qIQkar2gUcM0Vapf
ewj0QXcs+nDG3zE88ZRggnZMtSIQjqwgvOzno7GoILgv0/3z0Dp4xwo3eaO+mfucY9u3evQ0C+W6
XFIKcdLWEizYYlMbHBGTIWpn5HQZDC4piLqi9VkEzNsYUsF+dlp/AWSKctZ/FwUqTHphUbbE5mF6
pl/38LIPAot2SWrcBB5xNkp3w8+7sW/DceLiX5D3Ssv7urshmd8QV6o0PI3tiG8iCLaXgPwp0zqV
XZRw4QSy3aS69HT3L/vpxa607+wM8zBSYcU8xUfw39QKYf+pc1bp/t4lYmX+tmNYQyG93swk39Fu
kwrtZ6PTcT/q2lyePP6Gc7kv2zPaiH+HudduTjMgkIKf440KyJZIvGaZHIUcGqfnJ69enwF/EuFf
wJ7ImKkC81Rwk9JOZm8f240ZXG4IwzshRh8WS62D3LFnBVUarjWCeNecL2eigHPHxZubC615zFvg
dT/qj9TOFm1ch1It7Vg/nxnPBqIwUN9cGGp0JEvU9yHyC4WyF1xaeyqWyMLnpurKkY720u0JnGfN
gdKhQyDJ5p5N2lsi0+gN76j8E5VLZfqdDcIpCtB0U8PZaT6PCrLibffewdn+B0epTxaKxQsCrObz
Mapvt9ACHz4WhT7ftEhDSJjocAHJH0xGXWZ2MJoj/OjVilLYrhQul/1LWJ50sDHDHQNS4e71LyR/
liSbUzfm8OqbF9MFnm89e+S0P7LIKatAWHDRyYAtag1jt2raI/ZY7TzlG6bsBwQa9xTUvLWSF5aX
E2LXko9dBDzxd2tcAk+//vifGJasFCg1frfs3jSWg//kOBE4TnN9huODD0S1uEKiQ59JYzaemYRo
ZM2D1BgJIVtyrSX8O4U6ZMt1yetzBbZDM/RZ3Bk2vQAEb0tFbdiYBLKvSSCXvGdN7pgqiGlPV0Ol
4HNwHEe81iicDN5royFgQgeJX66A3FtcHuxRClm4GfMpcoqhRrI6Vpcw3aFKDV1H1P1UyAiDcT61
X+5E8VzlfszbKOvTCS8m7/rYmOhEsXHZykGwdAI+I9KEWjWVPaZO5UcTJQGuekzL6KErunpD00OS
+Zv3BZZsS8uG2KZ22USOYUIJZylpblcDK/+YUOKULLmmP8eJRRaQ2vVjVKQ87orhwA63Pu6YlMpI
hTWgqbsHD1mmjtgcnkBzfoc0GUhwfG0bWxSJB8zkCgbEsRA39lesBD3B5yftJGHjsyX0xw6+XzTK
IXxQy+dshxpdCSgkO5wAfHDo5WZIfziPVQVTvib/EXbd+3knBz1dUAcUFfeNBAUfzsvkYC7QGS5l
vokZCk8n9jRGBkbeAbaYO2GmrUZgVhk9lBpopVQd5fEqW1E2vm/nKwbuZYaCGL9LR1wEzPu1K9yd
FFKb16nQocjXsE9xiY1mp64XuTBoudSpPyIy8yZJ5rcrLcUgw9t1FKEiyR31pb6+gW8Ux6coD5+i
V3Uhbz81/vxL1zZF90g9pMDeuguEy/cYnK/gb9CuFS2kuxRG7YM3BR6guPwXmfFTpp6BBIl/oqBU
wGqdAlfQ9eXwJ6a22IkpC1y+5Teg8UDZBY03dCC7Ex/1qTKgjRhSzfoK2YJX41C5N1FoU+NbZyHW
QtCQ0GLvmj4ESuAO7yr9RFbHz8vPZ6dlrkHH5mIzzhDbWFXI6pldvVsJHBaz+h8O5Poo0EE2v116
SaT/t1rpnWxrGbFECSVwVodW6ZP9KmWPREs8Q2sD9mo0SIxfFZfKnh8xuReIeUicQr2c3IBRhESm
6frhbGAH7j+Ol7yjX0wGRseW0l9NsjNeSWX8F4MjLFMMIQ5g+Qvn2BbrxNH3khop8NZ4fjSU1yQa
BrLkc4G5yXbqUONM1oY+pjnm2zObqGFgKqv1HQkuiBNawICdSt7U5k3EdTgRV3U/3MlN8HwDA8Um
Aa7/0OzQRIDy0+Pc8SbMIDQXw52hQyBfSK0btwDfShkvN70OoHUTKoqztk0ZaVRVE5UWwXR4fFwo
OF9GKfkkoUZs3fR9cscSYWKkoCF3eG4ZA/wcY2CT/acap1pbj4XbGF4mMyZOKOHZyym4A75omMTL
vxJd8yf9ZXRB7+bnPxbYEDtcgQ+ne8kfd1CvM0EVCyVT9v/aaitmQZ62VTuthlNfpUnbqOAN7e3D
rfTztJjNw+JkUBfiapXnMameZ6TJYzzMZMnjGw3mHF8pg12k9ULUKl4yZbiJJDDNMf+nhlEiiByu
4gKPO+up1xSd5kjWxgdjVr7R7RBXdA7HxJds98GO5tPJ0wC+FhWbYe3mbk/PVwiW5bgRUhx0jDdz
DGeHdHHoOLCqozMgFXsCA+es56AAPUHgPC1g3xaGkucL114zxGyZRIsciPL9iUUqntzciCgyqupF
6wuTZe+vYSVBJVUlu/OBjq25WCOD92dqix7n5YDtymuxFtuvWdVjvGbMN4EkdFhdwVDJSLxvY9RN
KlK4iJyvbDHcPGqCt9ZW6eVep/pMAkTxwmvdi9cLJWp+mVFEXNwRBI3d1rBW9EMq0o+SuEeZXrQT
UIGhYUnJvtw3VoyGD/tTBt1vQid29DKpHN2knSymksg8y5hHcNxMzgS6ah7oMBknF9MqmPuSsNW+
NNJ5uFy6zQkHX8LgA2FFzDJ1tRB6Xc1e5jvn8go2h+HW1rfWoR2uYzDGf+o/i5MlGXZlv8ucZHCh
bqtIvlPGAUptk9wBHBxOF68FuUFgha9hOep7QR+7+f8GKGzZoR4LcM/10z3e6NqJ1K6faeWYcRcx
Scm0yDtcS2bKi3j+eQhimfmwt6hA//cYp9VQQw+ApzUzYEy91ycqtJIvECfvdsBjqL2UuaKGi2Fs
o3shHqJbc/P9itZwXC6ULMAKhbNelKCMWyXIAu8eJVVCRwBufFvN1EEt+yu14ZfXEgE6dWgVkapL
UYijxCQ62+1gM3pcLpDsmJKDoMhPKTalq+IC8Npg1YHoCkQGSH+uRaeHb2eKAticc1yKdgIRIB6d
uVQ3w8fOlXPB/T8qon6K9bUZk2AbzpM1u3extArNRgHdQxfmIKjXrwL6Z4atLL5Zs8lBNc1r5lm3
WzHpSsmF48Uuty/84aC9Ehf7f6T6hBVKYY1SbyJy8491vfhJZY1AhtGjrWb1x4wX+U9WuvvruUnt
iIjM4fr6SqrktAu9RA/YIMtb5JD5YJpEwz41E8WA7IwwRbOehPmOKMb0UZnwsXgbmYXZWgfAL+GQ
DGjGuTlN5xkzuCu7IaAKefLDS6zWNE+zFrI5XWTqQklYIfIq6HyU2bTh6l48Ei1fy8epb9+W5jJt
A4m24OaCSL9AKT9YhbiXS+pfHJ0eky220FFHi27UHBz3LiUrMzoDmdljWW9tkv94509RfBoVT5BS
JnDzrdMFohMx9TSsD2vg/PGlFER3ag7TOcz1w1OB4SL6uYLTJCTNKLBWVhwutAJwaWs5i4Zz2Rv/
dG9M9wNeAYMRiuDjYv3vcqo6Im8HUCkKAbzxn4hhTrYPghktQo5TF85x9hkM9JRiCyKSOmba8TDO
iy5ZPkRzGIbTlZP4RthZkcZRU3f4OfkrMxN9dnCeoNng8EvyUQsyopSfg5wHSFMwXx8OIK6q8ctc
k7RuzpGcHq4m3+6bG5HsqcuRL2vMiHv38om7iWTFxmxd5OJ7WCfL8iDzpcTN0QgWeFIRZsVlgVmC
udmmHfMsF2NeafoYt6pOB5lzzxWnejPGx5f32KO7TLA9DDSwokRUMkx/znpI/qCBU3EOSPU2QgmY
T1+qXXoD0ivoDiYSVm23Dun1IEExuvDDwAFVZzpcWlTj/vzPMcQWyAgFFdoOqC/gsMcE8W1H8/c/
6gicelCnefigs329JNukHyNbNws/27Maf9dt+RX1MvUMQpGEEV9dZimeb7D4JH/ETs8FU742fWZM
pxFvqXH0D6ZpqceosQszUhK13bu0ylGMIBAZfYohicMtd7vs9wys0oNMqD/p2l0GigdU7hzXPEv0
tUXTUmHlNLVc+fm/YPlaveIWsrtbbK/6yb7HwkSES1rzRzBS7k3TvVl2CRxyyN4qESU1KsM19U3j
Mwmk7J8u7llSevW/vlSdhDG4rFHkLC/Jnia0yUyVWu1wkSn42NoSb+ypMFJcV0hfI1vnEB7rr54x
Wadnjj3j93ILhzzFlJaCbKKlcUFl3QU0UB99UOJP24ilfygbNHOBVtVNowz2yLucZD/TzLSHNdTU
0tjKYqGvQatWZ24bVuk/Tye+pAhL+K6L0zUaOWcof47u0UJ1Q2s9gke1FjwJRygpxCb2PY7fLuVy
QGUluZbGIIlvvPabPd1k//0BzDgFdiGD35RXX83Q8pm7F8Z4cxjlwuwMH5P39LTDZ1eDowKcO/v5
eyyUSPASt1Rmg8oLnn564xTmtbpHAdho56i+3BBcoi/sfFIol3LI3367cr8DF7N/LEyf1fi9qGIh
y/psly5w+/DIeMy/mwbaHODkWoHz+aoePtnha9nKHU319m2WFzK2w/k1LS4H+MPccvgd+WkARXRt
NIaIhfcPWLeRryHN9nwWpeL3ylcCxiDPSeYLy0FMFZ6E84jMHsfSAw6rn8VE0iN80ifs9keI86NN
oZeHZ0RH0sUnsNHJdsDTyxY05qw46qqlE/R9rztB6UC6ToQ7/gqdRD7o0FwnCKqQRNuCFzLe+OAs
z3WmS0dCr0zMS8yw1w+FBU84Ub5KVVP6qUDGPnjcr7luoPGpxVeEmWtIJbfCDPSwg8kzC0CSTFVD
Ikx1YvKwsROzXoziYZPq2aOITaluGVD6w161KrqrqxdtLn3o59Ax7AHBS87Zi3GseNuhXvfstpWQ
ehFoobibixwl+BMmuPKPFF/CBCJ3xUiE4DuIHhouaxRkfh3o+ogDK+fwUL9uqRRHPdKBR17vjRSc
nACU/exdjqBbtI5Rus/E9VuFwin4JM3dp7nXn4UB02BKHQE+w/qYtrCjHK7yAdHCCmUk4z64f12q
BXfmKKviRPTBxwn1Hftn1n6RMLlh9BmsNZzKemo5H5HNUoHCApfQDIqfh9dZHoHX/pVLDGsWnqKj
8zPK6a7lAT7UH+aj33obeaJ+ZaxCFWXAI6oXStPXv/jmU7u8o69Ij+YmQsHXgJ2WDlzmAPgCi2z8
168XsJNLb3UBqcKd28QeR60CX4+rHtopeZV1LhyKy2vWgHYX3QYhXl7+2VUndwOKcp16zQcX6uL+
nbRMi0kfc2BIxYfL6pM+tgLpSs35LuMtn5l4x5TqojJO8yTpXGbW5Ghz1RJ6M1tD73J/uDXNFMQ2
zVWSuJKAaP0Ym1Dtdnar/r+2SlwkAU4waxA4HCmJcs4lkKKVsQAE4MYlybrPdcuA7m5TFrz4M12H
+g1nylMNPsD87b2Kq02f3Z/aZMRqnTn/gjRsZtgYiV/ALNIC2qiw5pd4eZWFHSNvm+es9AWRPE6n
ISp5curorQS8gZbtyVJNNU46P8iQPs5oTV8gOWQuLTgMqXRRJESdsaeQQIGzSG5YgcTxwVJA9ooc
gvcWTQW1YEJLJN3Nkb7UqOPaQNpcX7FdfpRbgyCR2ErcbDOdofn43HJYjA+75FI5qTrzLJwwX+zL
WZZN28Xb1BPOuXbsFJ+zXqEJ3jG/8QjDNYdAuP19aVzPeJqrIRXygGc2XrqhIVcVEf6uwpQrhjkY
MKPOjreDAtE0+kOmEqym/lC8vtPAr2asfMz53L4YfgVxznglM8GR15AGldJJQ8/RX4bJyblQpHbC
m1hZ1eDgiN98v+JUVKUUz+v2Dmvap34SM7FRs7hhHFzgRzvYjHX7H/G8ARc0JyVVKXhBsYA8jOok
raYL4xyZqxgOqPcz8si/scCT1D7biPHRYgqqhXitaskTeM5Gmv6GVgWvBHGCmB3Lu2o1sBElVBi+
RPEo1Vipy+S2hAr8dkmoZ7Y5/VaxSDDS+TSL5IpKDIrs4vZNQHi9SU9g2sHEa65Ob6mxnTaaCwEp
l1qJpo1Ub9bTmkCmTzIzNzc/AtmHOg5q5ImSaknp4HvBi4wJFg7Ukzvk5w3o3quy5XiYB6dWu8m8
6WIBWcJzNurXxsGnjPyQN20Y69QEkSRsz0ARXs3C2Uo71D0Y1OenAtkf6E4N/jKANIjwM1zYEvm9
PKznuAP0pQxjpjCWiCPEHIZ+zrMprx2371e7LJ65QCNQB1/U/tJuLrhMLRGtOR/f75Q3pYE4JRb8
ugGtptU5nSBBzXIgCsCQtWf+syULRh2vR5N7wpjpyjUJ+UcoVgjxrcrlDSnpWCxfJ11m1J9hgPRo
Ukli4BD4Ek6BaE5UtSuDtPVBasLmHoIQGzOfvG7mnhAt3cT0cPsdVv+EjkPd9UdyWNL8sjRWsXK9
NWmikkrIDrHDOQMhRugiz9dkVGweQE5DwMLBPm+JwxWFC+WF7JYEczSih1rw+Us9KColZJCDV/qi
Q+rImUw45UFSdbR3zGIgQH1WbZ3OV+ho7pXlBUIZXHh8PPhQYPniADkst2jTyzZ9m1Si7YdDBweD
A/1Zrhg44NPfGN029vtHyXcpzbhzmflAZLkpcf3nHIG4EMV+TFXUyCx4Vl5cYKrTYJpZmK7sJVeJ
G8GQmPjghRHAlh8/2YQEpRiUMnFghue5cJdNdJoYQSZsSskIhtg2exwRh+rzuQLA2sl/cCAXVcun
TpuUmJnnnsDAipOKdBn5O+SpzAXSYzBNu80jzuw0siwd2e2fsWg3SMMLelFbQd3yVlDWWvGGe9UD
g8vxEPqHO16gJ0jhyNW+JWqbsKlw62XsqJQjkJ6v4f0ZqiBqBfLgo0Lpib0jKNX4tAiUjG0/T6u4
BgIL4XwaG8Jop+5YtM0p3tothyrPiFjkU1LcHj+SbCaNq4pEbusy1c0u08zibf80/zhJ33bPjfvD
hvCpxchfjX4ZaL5KOPcKDkHhtuqnDPckGv4s0uhTDDMHAg5W3TgxtgiY8jH7MUD2GOkC69HUashZ
inzuDjgILjuIgGZlvm67RYgPmSCFevmdJbX8COzG8ajNB1JF8rlLLxFPMlWsUd9+7TgCGYGTOiF8
sVRAlybrx28XRkHJ4Ah6afBmKsb4whEd/qwcY+Eoug84+fowFGVJJmBeDJo9GmDYGh1Qt+EsV8dx
vIr50wNRx3DHkT+Lc4ABdhEdrEmDpKe/NiAIOxfsmNiODeg0lw1IhxKvauPvcUo8Mhy7GWiignVL
5izZyaoYfw6A6kD6TFDAvVuOOxX0peObh0+DP2thW2xtXMCTNlNToJht0WXj/+BbhRv+RwcIMIMY
pnVbVEkfxzHZ1WvGCdss50BuQptYRsn1mewRta7xdZpcRwlTZ5ybSv0AbpXlgomhTg2Dhm84z6KO
hQm9S77fz7DSIDLDBHTrpG0V3McO9qdOwt5ylik/adAfRjqUGGanXhQb2ghTSSQ0dvUuP7u0lGBG
1qvRXqW5+Ut7l+xiqBVM40o0FNQpaB4KU8akiB4b2VpKYHgAXkK5FMxGziTW4AS1Dt0HNXtjWoWN
69TlVberbLzAEwLHPLRBQdZgWShhy6Ss+aQF92QfHcrlg/5yES3+d3CL/X+hYJPoDWmKjDk5lAR9
mjRNGnj7ZvwZcqXlJsP2aoeW1wysT+CSNN4C64cUGJOdvEw0CTz3jZSN2kAoaH15vigydc36NSft
IySk8DUX51MOzOqXzaax4obCzZkwknNEN4Cd2Y/R1YgupW8ZKk/M8R0H82IuCstDj63IMwr2RQEF
UvbHFidAfDwg1tGQfBpi5gQzI2R+b7nI0Tszxdxz824jUgyCMiL4p7lAGvcwG+1S+1Cou1T7T9aF
7zgUosYV2azRR9Hahz3EBvueyVww3O2TOkxiNZoHXyhxH9vUdchPLHnSD4NvSU6a/Wbp6ag6psw/
EMhTqz7PD0j0MdFSlFADuL9mthYfwYOEPbGkWJKfUKjbC7OUcgo3BdtMIY5SUoFciz8WqJzdAqF4
Ax1trUssxBGzt+l9fs2jl2LhDJpWIL2F4e2NeNkBWtOkq84y4IuMIKdHt7ZM1ufkF4tCuaMlToOi
INWablsPz2jijajTP256Gs7kPyVAGI+VncIP6Ty56OOxXN0bVrbwahPaZM9l6GmLTblwnKRYrIRD
8V3ucRtr2ScDVvplYeCSv5NmETiDiWGq893DfQdnD7xjVsqSY2yni+RM1/T95P4HBCtYXhTdlTR2
FShGQSuQvHV3fnuRt6gzp8pfOGyDEufeYKtzePASh2pkJ4rqW5V1SgP53Xq1KqyBisjfHe0f0zme
3n//fZVnidfE90i5id0A5s613eHxpv4GlsfQA5NAn6ip6/RvYV1jE4rxbu7zMzKtQAK63V2CunmU
eFa93xJaIqpmOSZHtJ9KZIke2hFSqnlO0FZBZPxYdo0Thnkobm7aFu1Li69+/QwtP6/Rlf33W2f3
n0xW4Hk+vsvr3IOSSCI1Y3USnIiSGoK/Zr20+rMx+jRTWZ2tNKHJZibyHEm7RK6Wd1Cd/2kXhSkB
Dj0oF44Ll7DzRChS4lYFw3TBcL1a2vC0FyEf5OMacqicgW1BzikKnKKUzwN6WzwZ9HUnnDH8BfAu
beH2RBFJNx6iXIAUIWSIcZizapGpu6qZyomiazJDMDsiK2O6ZZ5PRx+R9iMRvRyEV9XfPKzJ/bag
HAEFH1l3US0I2hZZd2kN7C1OPGMO5YUPytILgbMtu6A5zItn8WMVoazgg6RujNIVcJEy4mMg3I6A
J29dzzK1QDJx3n5HCMuuRc0JY/3nQHYZfahXNoBwzapQxpAwvfFf3oqSGP8Tb++bF5y1m56nZkxh
/EsVZyKt4qjQwQKUug78zH6eGM657wum4qdhcTtb3zfMWUL2B+K76pyG/HmR5tlirMd4h1Lr4tHm
fLBs3FMA++bjvr5kfP/kW3YxgNp7o4RFyNY5j+PJwsEwvsMJjpHOOi63iTFQX1gPchF6gYXMCGNV
qQwYyjRRS+D3e5cUFUBrWt/j4qA76edKUnHLWD9KBGNMGHRMo4NvkejNzc2NDuummA2rS2bxqEhm
uabLRZtEG7PKxg2GyHWCAswTSi50W/B+neFcUaq+QeO83Fs9Itpzf+kSOrjA7KLBal9GWlNqMwUN
1qnJxkQ6PQtl9lT94MxlTmQjoZi8FnCW5QLZuNazwByQj9jnxrngaXW3J26tJQ+ikeolCui2yZmo
O4J1V6+PW07gH7oA+Hp6mZmAOw6NKXwut0zGhKQDbDn9c73heqAeYdjZMfWXfT7Zs1nGbh4vj+Tx
zlH4R/h/0D+E4my4H4r8RA2pIRv64dZxc4xmOaL+BoVOZfGDW1JLyel4Yu8UapLEwOf/yuao0znq
hcsfJWeKJmjqegzQhVWo2PPqa2Dfd6MrEjkFzyrqdbPr9tZ1dguPQkdOSmiGbX8KusB26LHLCRiK
zuiuoshELx/Vq9rSpUy+NVYhFp7zp8EwePyBq29Mbb+/Fgab436ATxfb0TldvRwkz2pPREgX8QnU
iaZTMuqcTDfZ784PnU47oCgXgBkJKECTzK4v2b0X0B0cx739/Pi/vM0NCKNXt1GlnaBw3lm8Qiu3
KpcZR8MRMXU8WnC6CUL1Dp4Xn1hlxp+eIskpO4VG0wgzzfuIpzViEPhq+80k1AMMjpkV+lpQWsBj
7qRrsd6MydHDiyNzWg0VZ0kDeju9elnQ87vJ4MBOSw0Z8Gg0svGZOAmbJt161V42f3Ds/cQdpfYl
cTELY9RVMEZCDNxd5x4wXtbExWpntY1Mv99HFtIni6g1dM/6gh8Ou9/7Ordcpjoeqw8y8TRGzw1+
BCCxjr9r9GGHj5nq5IrAofnPTchYKRbeV7d60NaL/TXUcWJZMQQMs52QvhM42yQPf+9ORjpz1gOR
o9miU07xI21jCXvqw3LRM260tYQWxLfYLyJHxCYZ9yJy9JEHXDAgcPmzzy/ZyuUUwxv3rAqiQDoU
5DXQIazplrSXGawNzEvYShAMcsrPSafL47OB8ZRvNAMQ5ixPnUglYOqMweeDr5ZEhU+xhwtguB+r
SOSEBb8jF4gBuVosNfWzvqDIbkbEY7PDCldhd0rhngl8KJQKdwchwS5OeYYiV4LPNtFUAktTf35S
Zs6MQwROz4VzW6klqCpomwLNIdOLvrNsMBYTyci47gNUW8DXRtIkdKuLsKguGkyWk6wNoC3ygqxf
6yy4Dkpx4GTvNpoKR026+/V+AnUQicTn/l0GPYTxbSkzjCAnoLrTLiplo2A1jZBCDahQKTfbxM5I
Md5Nhg+V/QdapA7ZoznsOjZlXHA5Byiu32kuoC/poVlbuDT0K8sIr9MMECaEW4CzpJB3qAikwJaw
z6/hHl3BHpdqdZAG0zEp/f3hKkWHw+MiP3i69rqs/1JtMSZN5jkFopQLOr9Sa/5AKrwbA9siy44E
YEf2paodJ6QZVWuvdeWJEnI65wP5BQNTNpzsN9q9X26tNOzKhbNUe8HL3bz++GGb0xwJDWCFan9L
tm2HETJS49bbSMvNFioApwpkBeN3g/4lyVAg5aeG5ufeA3AcHr18LLOFB8sivPAikT2VpStm88rS
vmJNybe+Q6XO7qOwMaNs/stWdTdw1if3+c3lDPvI6PkX5smv+aO3jyGYAZvv/TR5td9Tz7IZgapx
dwdgB1vLXeoxRLIc+3f+tp+fi/uO+QRxIUuURTxcj9sd5ouFqLGXach7gzOdgWg394aSFVSUQfqK
fPnL8HOw5YF93UfVROHisUT2k23xyjrQaBGppWxmRY0QLUNbzvCQ9+bRsEok3L3KbHsuhEXstp7E
Wm8sCtJA3EwDpqnv3bMbdMxkV5VCo1DIjnPU9MW4pJABytBFebGGG8SGiIWnRf5EK40M5/EdVHSO
cxNL9aRVSEKmLPfdXWUOv9ZfBFj5unAxTqAJTPdm5IxvGkyFHATv3GOJmyIpqClXbtxUeg0hz+lr
eIEQR2GbCJyJBGTayryZm9Y15G8IsUqvKojqeEqRQVCGADylVG5vF3DgfRSeqbZHWtq7Ubv1dyIe
vou1v0bFI1V2922FYRwqhG2G66H/wJhM2+J3ornJnaYnwqZ7YdHe2kgoQGX5oENZCFaxFUwvC6NC
xNA9uar1rBu03hSbRKnLLdxqFaSgo5eIPuAcXJ+oiEg0EsHjUJCsj8/BFLT1qS0lKfqPmTwFE3wn
a6b070pseYQdYAvwEIaP5/6iZWF9n0lVoYz6qe4xKUhOrlWvR9O2jJhR4Jsq0PBXSYNmWB4CJ+pq
nxCEDgKKSNtjAku0BBMMp5wr6O/5X+4WxzhqOuOb+/KhZ/MTw40UsVWg1S1kC/44Iuqp8Yc5lFwZ
qlQ55wrVVIWF9GyAV6IZo3AUgGBLkfObziB4GGshrNDwI6FDb11x4eJ24/HNy+Du1ZEFEnO3x6iH
+tsTkfl3bZE447+4vZ9rtS4NCi4ObLAY6fmwyeWjjG5y2gJqFNwuPJT/+B5UNO08OjogbTj5k58h
7kMTOwCbdcoL7ZhZuo6yw4ELu0s2AOV+gQhwwK9RilmW+CYQRzxIJsqSQUDob0w5NPtAfXtT+RLA
jSlHcIC/Zwp5wf9J/S4DXY/7t7XCBmAl9kOr6xtnyKiKwqeKAW8j4Bsvt5lqQx8Pgs2zGlk132Yf
QKoVl7ewZoX4BsI7hO/0TAt3R3f9t1tBOqxycHPtAVKSHd/ja58ldagChGgZOPwMvMCXRsXdsbby
Qrp+jR1M5lOVitxgDt82s5dwKBFDOWgGkmTp0TY+lXVxAGFQqVRgnbFICz0wlyPVAP1BBwwqu8a9
JoZGwsaP4oVFsPAJVXkJJinbwNr4woBhUUZTgDGkOmY/CgZKiNahTjJtoKNOx2S8nzS39QxDKs56
5Chx5D0UJVKttOabHyvNeIhb3pyUwMVBBWMjabP6diUvNx3JhVhZeFTZyDXcn4AJgDhlGsSyGx9L
yt4vieiEa/opoqgTaD/Dh4+ljMcJBrw+TkuhzrBnCLIDadjXL6cjyI4jmRP0WpuIcTC4CchVWafM
wqLPVhGjp+a9MBxzKNcjqDgn9mCQabFqnMmnO+NEYvSqI1hBMV7PKeNmlYuW2ZfqSh11CU4hlTmA
Q1mehcXxYT3syb3hRpqeJ6OrivESTPze8lGXtC9dLzkh04t/RnNTaLVMFlekO0NfFpnnGvLY9zpF
zPJgHZ+/PjQvjdQm0PHnLkzushWKMCaGkRQCWrZazJybeEvf2befRBV914Yk7Xjvl3G6Yykgf7dI
4meSHdn3F684/d+4zxpVChbTdww70YbZgeW3j2tnqQsdelX/7tlIg3mD68N8IDUS92Dks8/+ujpk
C4GhQ9NyEZ2nyLXdDJ7KBFK+oG770tI5T1NRNd2fWuOD6prKMkpjtuNQlL6Bg8rEjbc5cB15ua4K
HAcD8haQTsUj7NIqq55so6IY+Aegw09DTSQl8a/SHFOfAxX8yVABsDyfMVS6jWzGgrfUFjeNtxy3
8DMpyxM4Xs4LuvCvlXbGVbPOW4TVYboRgaubIfJmHeNkql8qbzRu4P9t2lUiv1ws4CQ8bl5K0sMi
Acfggwt9ejJM7v7kzkJn307km1Ub2lWF8WXXSJshV7TA2t55X8EqvgGcCCD4Lg7QLpTP5hNHBWsI
iHPjHicEwr91rGDovKGmtXioaacGp9qSha7B5GMntkEnZ/2Ecq6zZ6STJSQqlDvmaOEiYrYV09Va
lS5uZleSZRjnY4qdXGxLlJo1J7UvPWT4Tn4kep3RbdnR3/tGt2xC5pCBIJeuz4lUhr8AZlqEow1Z
Srodlfqgfg7ZVROD9vIgJHqU7A8tjHJ3SeYvABglQ8PE0NKmCu+v2tqfBJt1ecDJANGGMqt9yjxp
3CpD9ZKxA10CuW+vMj6C0faMEQZr1lEN4diAztvHqU2ll2woGo8Ii7Go06jbQmrwZagUYk3tPEAU
nS8izcMvOTVk16JYu84CjOQXmuZvcCm9KQXS9BHpmwgxRiHWI2cd8PM3Spf00saxn1BDBkCkGCGT
AAAVKfOtbkK45B90HZuWUxVTOCrNMaLNS4Ad2YLAtmvN9lSMxg1TrDZjNFsbcnYxK8ZlZ06wwj6C
1ceg73Oy5p1Xxq1gbHNTKr5QJy/clHdU0ii5McVrFy4G63EE/6erfe8VmuUdq8HquI0KvslrQbwB
TrfCUuhPJViWIuZVAA7iHbxvQuMqc1gSd3+j/caRbtseQZk6xi6342xwO/q/n60VRXdKTk0voL+c
MMPI5UGO+4BL6pkOFlUEdPZNmwQ+A66VoVNdFSTFjqgmi3sQPxWh2kG92L+rIBfT1E6hdUaulCZ3
l/dOmoZNv2cGMYOT9OOEcKIiMfzoyBkGp1TPHYjWsbh4pKpt/QOv1sSYjxo3G6Egh1bkmTLc1/Yj
6p1ETDtYo4FPbW0dPqvD0Odu7t1bHGoPEis4nvz5i1zb4syaZHXYECWfee33CUHfgYNT9iM8qaU9
uIgLYj8MfJfquldT7twchUFoThzdTvyPbDmFQ42nbYih/Cyl35m9xRKZTvI3XyZuGw9as4amfGb7
pTVb2HBEVyxkSZ0ABREefyHpdMX2YnfyQou4I+OblG+bMNkKt34JInwZAVkaUzfO35NkSFbr5cau
9SXJZlQ62/NSWANFAbSIskOHWoU+zTsOBT0911+SVkzvLBhnDKn9+osbTHeIYigNLjtjXDP+ZDua
U0hKCuYKj8Hc2X+PKa4SEqiO8hs0IQ6ESB4IZvl/S73fHENbvt70WWgrNu9xyt6LVV3gm9fVhFNw
2l1HAS2jqhFR/T7u1Hw1BA1R1bYevcNDTLLTHaSnqDURWfB445DyCX+rQqX4Pm+c62PW3cQ/A7hK
O2fdeM4EQQI97PMCrUcQT8XZBuqibzuQDHPUETuuStdQNsWoGvrTVboAo2ndIiC+uYzcICu/kiII
6VTh44sqdcWq0DSWMdg//yinmGNlPwnw4ZaFqtHC3MRiHnFqKy6GDPu2azyidsbyRnqRengE2GCb
SFlqvslTnzKlkL4vjJ6OnybeahwOVXVDofgl7+wUleVjmod0heqqHIuy3vBoG1C4sYyQV14991dQ
OuoRDsRiwew5YJ9qyW7M8DAKlAfLx8CZL5f6wqHq1ZtCFa3/2ZikxfiuIn4faQEgrEx5Jc5pHtDd
e8w88XjzncVwZJUT8s5SRM6C4XHaUb0wdv/iqlxJ+u2OEbNyuWVG+RV7dcHycIPjnMOnNnTP0QHa
iXINdTsjNgi90J6rqMv66aOd1dr3b98ffqr3CbFI4EiUYeLblKCeh41yXsNjY40dgGCF6CVVC0Uu
lSjl8AhsALxjrB6N+aDcHCSoIJf3QzytaF0ZPDvbnkqfIQGW4RHM/RLGn9Mv50Q44bTfUfpEignq
n1nCjap7D+Qb00bRdVvkNgthb/yYbASXHWthxNvuFWjQtOC2HF+9w/9z3fZyeAiCBtE8hwWysJrv
pWxWC5yxtRjwms+0Xhp8Et0xwMeaylPvglNVLezak2N7kAt684QCewBQXSFPSvyi4WdIqLBXJU09
4TojNYPwheZSnpswQj6ze2Py7rS5V7OYpFW354B4kdBhEgM8w9RecpmPXSQrlL5eB123sp018HMt
3AcL1p3FRHMDUtwyEiGpElJvyZMpSbny/mw59BT5rMELy9DfHCifombfuEoM/JHUbFndbFzN+4Yu
pyN9KCRZkBuXhegfKEcq52xXwdnWQzfcwyDkXRKcfU4OvEGSrR3lsEIvJGKPo6PeuQsMfaCtyJmZ
u9IwumoS7/8ASsxh/+zRzU65KIWTB7HDwwM5MCXKn/KMPeyCFZJ9O4NX0aCBSQIF0x5Ql+0l7nDd
3dH2VUCHz1IIyNMuS5OWRO1UheO3f2Y8AF9mPBytbuccXxM5pcz44C5Dr12WdUnJ4u2xXhHhY35U
Kiat3acoO0D+v163sEeR+j9rSQ5QU4rgcLUZNuBpZVCCjCd/REHqASKoj64/g+NqkAUKDYc9dG8M
306Rna5VCjh8+qDeAl/0ABbxfLngSY/X/bnB+uPKiEk3M18dbLwTDS/9zFzl5iYJeKPYw/GNSB01
wCG4dvlR4Lh3bpj0k9TXhVSwPrFzWB/UNUZZ01/cTcrkywHUT94yMGeEmeNVlrx2xm2X/cmbzgwD
t8PPvCyzoqruHCDNskFjKwBObWnhjbxa0CNjC2sScwKtEUquoiZlau7KfytoTJus2hxQ6IYqXqsx
LbdTMMML9rzqTkNKllaeqU8AmH2eaRH8+vOnHxgz3Ub9ddPAKo0OjSwgrj8GJWsSZLl4iMEaf69d
gudvTHoyPjGVYNse4GIQbqtBoWM5zfhlTa0r/RJxjj9LprxWhzo8KD638yiPM6VPGCg1k+CS4hY3
jiKzVUGe1qo2z+r4X2B5mQR+pTF2yBG7jdlLtgHRXSduvrRmorf+/sIGz/8OEO/M1dSnW0QngDQj
QlstdK8G0UVFZzT6TMPY11poqs6iTDEgJy1lRvkF7WTBlfiTWMbNuvTydUU8v3iBT7gnoNffokDy
kHn+CMprzyls6HxGzx0k5xWLYoLIhd+VPGmXmIvfAcL9C7U4yr5uZKEGGcMzhHd3FJ9aCfiMgABu
twAarOt5l5d5HpaIW64C83VXS3ZB97td3OfZNcNWbPbzmenXv/tm87BttOBa5RC4Re0qiPUL/IJT
Ot8XS9igauEdNWgtx9Vn4SzayxxveUiOJsyZ1smqfKxD7TAusnCBMh0zR+4UxjKg6Rmj1ouPlk27
05l5Ks0WTCUT7jDabJX5PAi3dOsAnEapeq71jhsJitdk78g4vWPGX2qQ8NezOGRDn9adHZUg60tY
9LlrIwd71FxOUus6q6Wl4vhxd/t5AMOxrJEPCC3NAkTj9kk/e0YWc+8Q4NCk27tM1ctSYpJcVPHz
0lQEpDvFD3M3rSzs/raZGf2YDgfRX1O7HXkfe1JN7qfh3JO7ognPRLuEPuOmYTRbd9ZiC/6sgLVY
lyj/Zn3IW0h/dPgs7xU4L9hzTWQhdJNuh9aZQRHrPEwOhBWBpehjU9XWSEFdP/PtzGygawfylK/L
PL3gerX1MKtfmJEjbMKeqBpoVOqkeYuQpVLu1ANn2LDeo0K10SJKlVLLRD1aTxkxZgw0y7bg0vTg
AnFbqOIkQbc0YFS6uU5bGOpCZojJJiJGpx7SZ9kVrp3nDLaPYBts/XeQwKD7y0g3Y4Q0bsVLB7kX
R/7vqXRos+JW4/c8ZcQohDGvgI6F9YwevAyaU0VkbC+g+QA9GEzeekUXH2wy/WyRqBTuXCH7m+9K
9MVhtwhlh4NEfe7FV+lRbh6bkDgASp6HNF5JI6NYx3Ywe+gGrRaygYQTJW8ax7NDozTB6T6rUzgX
e1mQd7l12zCz2Z76IMrmO5Yeae/+ruI7MKdngMW+FmKxpjigIm75dibyghpINPiIp985G1gaIJ48
CFPjyVp3t8vGJnbe7gsz/zaJT1u5SUzsUf6g1HzXLS2mCJpBV7p07IHUTYVL0+UTuw/5fR6Icl0H
xnWrJgdJMv62oWgalr80CgsJC0xT0Ssg0HT4+qbcKNADFC2Wz/0Xy5UtdxIaak4AuFj0EKO1iOpR
5IDKafeHGcjGMPKeqrVzuGmWu2uHqEFTDMbb5RGmw9TJxYv+qUdi7hK322NJfqSOdD9xulqNINsh
P8LLSGklh0j5+TbsI3yzIEdKd7+0WefDsdnM0K6gSUXzTITCMRC7+0dBI978DPfNXQsjq5wGiG3W
y6zAL1SNqhEe7i5Ss0y2XgVyuipSXOAslsRjHFGfzH5IqtAFrafz++F9QJowCTAYqcBBAdG5tw3W
MnDccwhW34mY/87/EGK3nVOyTyfIOUNNe1LFS9fJydlcCdvssTvlcXcsw4CrJ5YZzVADyuoNrQL0
FNu9wtSjIeTL8mpRb+uqNueJzLSis6ELFG5mRq10QhXlrrP9UDhD4UOrNarXDGXyEG3KS+Rvwblx
sBrYwzpEHQX02jJjg3PB/rwdn6scVx6Dw4OqrrA5dxSy2HZvkQPowL3/uq1awISnqZS7QH3EBDA1
yT1vQnzYgyBesIvQrjX0k/cmB9mGwoP2BufqGOBTI0ksTcA5VQ7nDtz6dis7kgv0nxJPo3KB0eOE
wNc+uyEqIm1aBGvYqPk0h4cG/j6Yey9oDEnejxetnDyDAd5LlvNaM3YyS0rCiEyqRxpWZsfFm1JT
GTON2e9g5HI2L/F29HiOqwjIQ0fiTX1ORznsLfsIqItk5TElt9+8prWd5EasxGe9bS0eBifb9zEk
om2SN/Qpt4mVydiNlavk85eBZ278T4nfdEOLqBArb5j4ZKox9vv9eq92zpmiAzzuRCeosZdum0cO
0CwgQXvDj1mfiupr43iYmHZPU7iXd4NdRti9L66HcPm2WWByHlfIODkdqPMQ9volsBO614iS0ZPw
8JQuxQ8kSoAgGKWnJ9BBoB+oWQp18HHVQuFBF/FBab9ACN6xov9gfPKyQ3tTIM301F6WW4eJEhnb
KPbngSZNQIpmH+IK0IUtxkLjmx/A/C110teZ9T1b2K1womSwKdpzc3I1xHhmvcsFEig84FX09VDp
ZRwxyNzZPFWf4H8/rOykLSn2U03a/YA3Ut6v6tagv0DaVSjs2sBQTooLf4JVLx9/uRZrgqIgTK2X
efazAKBcAdVkWBtNx/HeETA4xfCpuAKMb+1YxTK3H3a63/0dk1+XmX/bcKecdAlVBcsEDoBPOQ5w
lKZ0IvHWqLXmyLbwK4bZGYc9D4PkjV+30Sk5VKom0QY3/z4s3E5CzC4I1Qons+bnVDG5+jv3k38V
Ap0CzyI/FTT7F9i5W5dnSdzHlL7Lftv7Bj0S0t5HpIIFoQZ6p4Iff+XqL9Fo9t2kWbNEZANpJ1/N
tBf5TKfElOn88hRaq6oXlTflm/cVG9TyL11sSQPa3tXN5IL9CmMnNVly7jbX+gtS2R/e3PogJ0KI
mUzKdlyqc/XBkkFq22IuQf7VMQauGFlue8zEmWr+sRw1JPZHbUBkyLRgRGNaV2b/Fjxh2SR+PlaZ
aqKPzM+uymb9opzCDkuxGiDZcHnJ2zH6mnYLVsnF8fl1emleYQJaYmRghU39p4lQNOnhbG7o0dPe
1TjEzwtElZpW2NDd7p4NOzl1osedf6kQ3L5QFIdMx4ZakN/Of78vCXxYCyzKhTkc/ogb+15WLVEo
wgkvKfWjUJ8L6Kg24/4CEPVCYTbyLiHXI7eT+Nd8KQ5ph8JmAQsMpQt/PTCH1h0Eq4s6TSrkf6XQ
GytIoqGoqbyt4YSUupxRImg0ZzKougIiOSYZM9TDHx+NgEvl/aUDuZ5eawALjKLXnJRQbNgaVurE
rc6McQzhkbPxqY863HeJZ0BhpLrpQnYY8NNIlspkcRCC1zm9RBrOvNF7JUAGgjkkibdJrxHDa/yP
0xlU2vRp5NZCfSbIoCzH1OxGO5zEMfNX0lINgm9hAwCisY6bo1hg6qGXAdf21dKvTtfkzbsIkhuW
/MQ7Urzgk8NDK1quhAWuRxLpa2F+a8iIKBYWpAIwByV3i1OycCzXLA3vQ2ji0OW82rtqbgcne/5d
buK9YsoCgXR+MCTghy/6C2j4sgTS2ofpfBej7ulH+Nd0cFd6yrM2c8MOUUwJfwKIZkwfpGzObtGl
LRZBiBRgimHkichMdB9E3G43vyFy7hp85GjPIChWRIpiJwrgfRQR2/TE4ZarQuU4b9RSECP2PLBL
cGl5CT6Z5fHKSPqRtnyoRJsh94xYuq7/RyvGPeIx8QA4+FWsn/B1WSyuRxfYU0TamHHRcfVKAMkb
iGh8fFN3HOE+SDy5dQsqOzWKeeCSCgDcilqBZQ1ZmDKiky0P5qe4XLfFPEHmlQySpsc/HiNIDTiP
NMBN5fUykSDmgPBPq8Fngn8EfyOJkD/QdwwfaoqS1Wt4o4TluiJqoXzWkjprsqRM5Y8GEH0Z1p7S
1g8Z2YNYzV+ALk0ZppASBhlg31Jtqbbpmk7Kq5jXDwJaZEfFmsYiPumK+Ykm3UDM6wRfLIeLpXHB
dQxa5Q/qvsEhYCf91xBiRIKLdYYpLICYoF9zvCStV6Gp5LY2IrOMuLeIFr9xazSxdSVlaiZyyLSa
e6F51wBI9lU2gIe36o00xWKV/VT2hIRzTBqopktimlPw1fDzzjYTkubY5FEhDEm9G8XaO18mjlbm
02dasfLFqZlf0L8fPKY0E0rfyiWcV5znrB+Jw7a93RYyH27PGykKnYho3JZ0HrbLFhGnB0vQqHcs
QtWkExhkFM4Ic6WxtTiqG2/LSjEG+Zr4kCZII+jHjTF4S0KeITy7nlRWke+294eHhGnmXjSlyOyF
jZoqm7XU1pSRCTWSU5Sra1kqOWIOzC8Lj7HFIX6KMddce3OOegqhg8rQDZhlCFpU0Vu7eOM8Ngba
MwykmIYqUW0OB2WeAIc0E64ViPvf/tOlVo/b3dQzt/Rx2VQtHOZFqjzqJQro0lMq6Phvh6tSdi5F
EqI+O8a5HlG/OB4oN21WEaUCLOwld6NBfJMCTMBZ6ocGEaFWE6+iDrUuPQWSjXE4rxu1JyBCwT9/
WDaVxK3Wfjs7Ugs4VlngUltQS6phEnMkcF5ITetiXZYdxtUGopkt9NgWnhO7rY1q/mljokeG9NQU
9dtGlfSuLloZXaaHR9kRuX8/PaiARBHGh2qN+aYoO8fE/Ug8v0Xk8osdXkLLGmvOOMik3CZs0wSa
KQcindpQte4nK8+4yIwUd4wCNecfIF4PMf1Nu2avC43TFzgzzSTTMO5ohCJ1VUXVqaoJeSVbNbPN
bltjDpx7SaDpLYMpJBFuDmtDdEitGseNzSxNVQoKygR4IGSmj2dB8vWPtkZwkkoLf/pdibcFyxEw
YzefE08vn0Sfm65NJ4UYb8JEXGVtMXZNcV2lpsIuT+oY/6Vg44fISVIQyIPfKuAEIfJL+bBFtfcb
JTX2xCl1UCzCvhqY+Hgtcyw82jKBbyIJ6aj4ta4Iw1qUI1BqeCbTV4BkYAkG+w+3jvo2oZso5faE
O+gfOXKJsiXXvedL/4IK4MkpwZzdGFPZCdlZw1lJID46vnyQImTsl0jtmsZbImlz9huwam+ytz70
UhrRhyiAucUTKTuaEfQcm4IkY5QuNtj5spuBXOEfd56Sim8TvJqRJsqULf2kCcJhRkmKL5630nAo
vX8ghCUMg/D265wVeXHBfDn1Be8xrXrzl0HhGwVsg6xWJSwxPSFWVxib76bX008SxS9rmTuiAkkY
V7718TmoV0KwCsr0IpJtlcf876kIP8CJSbo1YH3o5VdwMd7chduZaKcxiapOBu7eQ+T6qgQ3H6IG
C+3tgF+quTq1ucztP5lF4UNEBARqC1ASybjrEOzDdjjLblZluCau2wfmidfeIZnKmP5LiGN0gt6N
lVKs/LW0T0Z6fufL5BXMrRfJtGJupyyfGmr48K4LDs/dDqRTkkApVhLjLM6OUmCTAQvG95wAdBIb
URTVVjAU0G/BO8hAu5nschwKNlIfNhxpwrtK1qnsVIbkAtL9hMSGRCZFtK0jJWn8RrpVJWs9/YXj
6iwuZcurD0hjInvh5f4w/HLXfvroWrGNxYEUcP+lykLysMQDqygvueYnB2cMfT7WWy+XrnL5vvT7
y36ffMED52ZZodzih68NDTwOFZgmRSU9W6QI3rh39IRB37ivY1EouYU5NYTGFpxI1bHmuDvoSsOl
DzsVdckZ7Cj4qMqS9KOIbBN8QBAZX762ecXAbHthX1hZaF9XxfdJgHu8curCqhTszo5SPI5LEJBH
KUbYZHRhpGlby4/M0LOU3VnzuoJbJeNpAcSqwHrwlVI4G9tbUm5uSxc2Eyk9dKg3L7Dku4CYXixH
5M8aGWetd+4aXjai9atE4T0YeWx1s3pM78JygSrHgG0/YUJWeVvc6w/iq24GhVgGIhWrbtkofQ1j
kMYfd5EpAQ4INPv9qMQWUwyF0HPA4ZgfcUZ3Y6W76PfTiMKurI8Z9WxAgA+GXYMcOUyaUZ2xHsy9
hM8kbuVFCJePlyosEuA7m728FA36W6O0LLRz7L75yLZAJCjxv+ypgey6pZpJVYSPUcyuzqnSlkm1
ICh9w5i2XefxgXWTu4tb02BG7MkmZ8/qmegISaf+DlzLjVIXOTkL8Zbial+3wujdjgv85hXlsF/1
9maMwBBhAjs4UWQToImzyJhWTeVDi0usLdJHv8z93xeqPnJUJCMkfQnLsMLVvHmwweZehsr8Rzz8
Qtb8g2OY5AA40U/dbNq2HbvUfsTz7ZZAZc1I85iD6HCeFWfV5UJNnClAyQuWE+LjdjDJW3j7mADA
AE2189hPRDGOC5bdGqADLj9yqvcaq/iJH90wOtDgqlfDbHs0pyY679J3ser7vHMiWHq2v9A4DU5U
MIaF+SWCNc/uxu2aZlTXcyT9tqEmkgZObNnqQH2XMAJ5sKQMfpH4us+DoVnzPDKc5/0JUxflGllx
Wroky1xvv+yEVvZw5OzCaVbxDsZ9d14/EWaXQO7FQVZlBiTmcfuFFvWq4zexolHVi9bcik3/jHsu
u+HfXJc25UVOhj12wgDFuwHl+aMRZMuO9IhoHB1U6V53u0vICsOeN1tFVayqyzH49OhZjB5FCKNV
uAZIneUh1+qTJoEf1qd50Nxjgm+G3ozY5T2t6mZRHmi3sf5vrViwMERsuUuOHM9bBohPCTaYTXVr
+3TkFL0chjAe6mLaJnadM4gbDjMuDH7fZj4q2Xl+pYCyjC5NLe5ip8AlU60IgkMBYmuoLto/kkjO
c8a26FKOmG/aPT8Tp+NNBYzbm5NTVQqL1ISPyxqlnOp4Wc2W65tnLfujbVaFm0OlpKc95FxOoKbO
0mIeZupUO27smw9x7eFmD2oyDQgjKmsSCHTR6YqMCmsVdhXXwIpIbV7tsy7y7z6YM8F8K9s3RRUC
tH+PHYXbWD6VTlIRNzg4C1SVIAMOh/Kmr6i2udcbi3JqM40HtQi6LIRpg2JLDc6xg/N393nfCAtn
Ory7+YfJ0D3zMC9yilezVL1OANQgmj/3zgjbkxRMjwrVW82/eIqxTqN6a9ne12C7QNuFe7TZ0onM
xFiJqDxAMzGvcg2qCabMcIC5tVv39MhdaeKZ76SdTF+bPG2csFJUBXxizITP+Yp7ixhMxrseP71d
DHZnVCx+uDyJWrfJ+/LpzlAe+MxfHBpQsSaiofbsn3fov49abeVCF/enZVbn0MGhoPD8T+mz/5CA
dw4g8KiVUa6E51xFWVS2UCjoRcEf92X6gi+vAxtu7pKi3sAj3CWxSNsJh4OvQsrPynHa0++DtM8U
usbVOSViVJ/1govMCOwQJ7RcnIyx1FHsTqOUyekixIi5ucu5TxTHsW2khvxTa04h/5hN9s9FY+Om
XLHQMgYuw13RNeo4htIWRK//QN1kWXIh7L6emgFlqOBO4VMo36TOWMtVcnbCj3RY1HGJYjgt3N/F
1udLI0Xy/e6gCKF1A3eoLxfBAokANGEEeEp/EsLrIF9SZ3uGInwgh3hjpzKMFpTb5yLYQEicWLQ1
+rRs/pMTAgeMG1mYxEOVefosxCnmFgHssAifKRTGo5u9zgto4CmSGp2gAxhhuAVx8syc2aYADki0
PTspmJWG+XnW/D3x7UTs2FaqJAxZLDIj0FCWyJYt1Y3fztc5RssGTkf0Y6qS+nLVUJkbQ8/4oieH
45bTw2JueDkJhY29NSx9vBCCfmV0dC585dm5245UKu21pJ33D+kpHpgowmF5niuNezC6dZCbwBBd
nkYUxsSCJ9EmWuNghnto/fi04g7B88QB0BFRpbeeiWQQ7N0uSMRw/ek42EE93GEDUvuMHU04f3rF
uVIb9SJw8Aji3EoO4twBL7nyw09mdpZ/zFIHpSecMuQJGm5aFK1WbX5biM7QJ0Vyn/zWeWdhOGfd
pPDIkYM9OLNHQPruRUqZfWRDL2IF3hCtYnw+HRCQvsaPuGj/MYwxu5tu9UpHq8TxnBYcS6P7Ox9a
eO2PP7MuO97l5Tdl0o2YZoExMplNmAtP7dWB9XmEM2AM0+898l59wrwxkgP1iVczvjROQgpDzIGW
Q5F4taK/CXNqTfAKbmbFWnEQfUYG7TPlvoNO7ij5TnLPv0N+shKey6Lgy3RP/mTWgCGZLbHqCpGt
mv1F9wysGR9y2xJ0X5OcDpFtRog3lAZ4LvVqg3s5vEkO4qIuOHl4MN0W8+JezrlOPDZWm1lf35/T
fJt/qd5IMukPHxeABb0M4+3nsGRQ4QjOYa4YxwMbYFxbrNLGUuMkeNCr/o4dgML/0IcOCCRXuZqA
8g/7LCx896yrbQs2MHS2Sp0zqAGVHhqyjrsDQyB4jUnlGga8rGLvCjlcejWhEw5xWC94geXSqPAC
Iv4ZWHDXn9lj0DDUaGKN08hD0BZ+9nn9/HRffwtAr/9lTR+VoXqkPBD5TXZM8yrJ2Lozv23rvcvt
kZCrRKpzHm2vaYNIFwwC6kRUyb3VkFSd8If+RWetm+kC+5wmCztwdNVYgFn/NweCcDnu93Cw3A6+
PJPIiBzFiHbTd9f29Iodr9bHBqe3+lW/wSwJbZbVIVb3KWnVJiU2U9DfJMjhcRDhEO+zTFTY9D09
I23W+t6LDfjk0ZeWC/GDoujG1InV9PThwLZxnaZwiH4i++WirF1++D7jW29CNf+khnkL5YKKtfRw
A6xp48C3ViS49THuohVNbpuCGfhE1VGdw73skahsi0ywUVcNqSTFeFhbyrpWqhK0ex1L65MIDsM0
KETCxdX+PkvVINnpDpwyPO5lkecAZ/6HQeBUYZXqeS7z13WAAO6GgWW1PlLrNMtpgu3vz5PyMae9
kcAsZtwpmhuRJyC3KtEWjHrjhVskO2KVsR5WG1IxiIFpsEm6F4CZUwL6x07oNQMeQGv8oUc+bR5W
fqOODnBoWE+DJ8KnV3wvRn5St4V4syRUo0VSbjFXj1A2gny8gVQpJB63AZZ1vv2DaPw0au/UtTE1
gc5sk178MN5EYFcKOM6zPgBstxkhQS7PTl9RH8GejyfwPJWn7T0rtboHhPYT5uURoLJFE28/IIJO
+popSb6SSC9/Xt9XzuRgwSRl83D2qZtVlbcI3vogK4qXPh/gDT40byNuv/P348e2b+WlUbLvxym7
8F2/sVByvcO92BT7mRfBfkKLc43NOapr1RVWT60CGkfD0lRP5+i4HGycIdGVWdNfwDH2dKBxLY5c
zhBB5nASPlmg5f0Z31FXiwnqHDXP1gXnV+bsgJUgu23wbq7H0uzjSMcR7vbO3y382bXLlePnqd6k
aLmVSn1gBmpjHJsflxi5DwoStvQZ2wHq5D/QMwZoRixnBvdDPktT4qpRiKDki8jwpVxLVoJmgZys
WGRz2kIeEs7ISpwuM9mPXsi5X3GBaqVOmXJObTOR30FyRNvN6joFXasGK17IaWifcCedL7SaVYe2
tQDhr4s/u611xubZfpHyzkVMh6k6j1MJAV6b3O2W6Ed4oJ39b29Tv7e9RPikA1TGLAJsBDpTUfht
spWNv2gLyetBiguq2Bf91P+IYyOk3qkUWPRIhG4qV37/UBhds3ANMUBm5WPvBVwgqX6/7+byT49M
uIfBo9f4Q5VW+QDO3jqFWDE6niyRPqfYfs6z0cK/03isGzYtV+G9o7HMNK1Fi9YaJ2Ds5R/j49Dq
NAyRYWj/kEGgNcXOZ9VsWkvKfoEq9U0s6J9v5GDHyZ1VtFgPbTjbKRsdnEqTCsYLAhdpbG70g3Lx
T7ZhCLQ0LqnCumqunGED1XqQ38Yln9zcAe/KCd6eSi2yvMfmnM7++js3DOHAcJ604J6FnAe8oSCC
xhpNt4kMbqZqCkwypJss0uCuS+VEsrYX9uCJGmwod03+5LIqEtoSueQq9NMBumdluUQTSy2M7Zb7
neQYPk+DmpqWpnYyIU+QPyQ8Fg1oxgpWF3JUQWMfapvig+SunLZ2ODmgWzLknp0szZQ8RGBzoojK
B4dBfqwjaekI8JZ34vwsA/h2FsDWENcQ9iu3MCGVfgjYIYJjNO1D5RGX8cPwFZgGaEhv3znPYSDl
llGiZxOiKNTFhlD57GygZh8jYmQWTp6q5sAu8NUxdbYUugWwrUtKFBQAQdbd6UFQztfM2nHT375X
7ooAuWpeO/1XkngcuZ9PK5imoLLTDeUL4sdQJ1GVxKV0UGESmrF7oogzuzuKlmmj3lHA+RbtfquX
hXHWwDe1q/ONcmv+BmocAKPc6IFDA2chE6a7aXGtLb4dXmWgLG7x7DlO5sCmRjouszCgrFDQFgI7
t0TDJSoAtrncedvtQup/gril2+A0ZAj0zm5vbFob9b2ciU2eI1h5xlBCs/L1YrGSquh2YNIu3e6w
dWVfjlICrCFpcdEr7uu2tNNzO6c2xWtMpuhaJr2900g3+xumcDbooTE1OC3DShv/+lz9YG1GTDDR
f9mfpFnK/DyVw1sd3vVXhxgI2U1+0tL85kEiof7K0aXoNUUOAL5AVPATUiIcIM92kF7CHfhupE09
AErO19CzP1Hbu7x5EOfCD7LtPrIFrotN9H6MN9i2p57bFyafAXY16VBCblk6H9c47DCQyfmDxzxY
kqDAl4Rv9UIzSjbg/gMDUeGMr8HOg95gzConQiWnoSe4tFwiKQsruqlhTz6gImTzy7Y1IL0yrD9l
DoSvOk3ZZOXuuqeXoEZStE+3F0Y8R0XSPVJMQP/Y5CU4x57bVlq4A1Xp6WYzIjDnXreuSdSG4/Ma
CItyZTeDHXFHn6pchUsoodUVi9/ItvfCaEy9ypEXRlitQW9c8HgpFZ3hveuVwC8x7a19I4GTHCBb
N/fkqlG5YRtMm3PSASgWyBReH+5mbLwQdLFxK38R2zhz1d6b6lcHuM0f1NxGPFxkoHFRDGa7tqoz
k1U7P2G1a9IXU4sXmt6oEINxeJO3sA/Zf0wWzp3F015y7jM4/As4fc31LkMNuXbDQodMrE+UXXW0
vzomlibsLHDjPHp35m/9ckf2bc985EmSAvZa4QQBh6O3jaygYE7SU5pFfkVS5/UcC0pDPbC/3z2+
JhWVhz8IHgonsINvafzuHR7vhMYpR4ty7okhAQVz270ZeuS6P2loqantrzqcWzFON+7eyLR7ZcgY
Gyq02yCWixyh4YtAJtcpcvFB0cqhhiIOt+COu7kvOzqmDKivvutWfY1Ubvegjoxy1gZAsKJQOeTo
r+D857HHrVCBBf94tVfZ5f+HSn576K6RAHWZpEDqoZkslFYVurd3Dzo7Uam5NG6QyUWqFuD2xm8I
Dr0qcxZ5eWMdaKbDFe7PK/M+MpDFoHh91IKdkrVyaTePKoPSH5mRO5QZg0qPBHUHpEBJCwqzznkh
+uyVxbdbqXlhLeHrMlCRZ9HLHjZ4KzZFB9L9azpebJ1wAi1KOFC/Q8kq69BgCAr8qkUOkDXN9yFQ
WAElr+AjBqxCDv3zclHZivIKik0WWI4t7jddlG+aHwZ0w/Tv+091uzJMwQJKyTtLXXgFC5nLoy8J
dEFCAyOFZymyDXVPaXsw6mjIR4m/n/OnZpTNqZv9DQTHf1w7G6NHgB1x21IN/qAqGwtC5iTpAFro
pEfDOXJTCZFwXplAvHo0tSl3Ij0u2Vq2sRvIL1Ah95GZuNAwmFN64lQG+zeiJlfIXzR5MfyYlqXo
xsnj2Y0/9eHGlFiA++cnK8uCfS474jl+3YH2ascOEmAgFo6/nlNu/734y3f/1nORLb0svHhqgTYp
T2jaK2dY7fGBNx4QwK9I35KszhyixX10lx7w02zy+wz4MhKVban/iWEjRwyXWowrnjM+Q4V6g2Bb
y8ieteRbVzddoZK5DLt48byJR9P30CvaWbkg3SjyKt/gXM6O1BM4MyDcJ0Y1ckmujHf0pNFEvlyP
PSScKy8L7tr85uCvIYqyFuyXzKnh0BaTaV56NONlUWPDpvQU4vTkIdK0Atrsl08AyCme7ZlvqFpM
G34L7llPjMPHkw/mkL1FjxcGWf7wlx3OLQ0L2C32c0gB+U+i1efB4ArKkmGTIGe50plXXNwWYv/w
3Lg+QlK4jY2jOe+j/CJSGQrWxYSnokIXBFv3r14qMHMJi2rshiy5EOBtTO8QEF0r/4zPMvHVi14w
pNOaDE/0GoYV/j7UxwroaPMGuSmywlx7eQOrKnV9kQOdU8YKJ1L2JJyV2BIaRsUDh2H1Bu++RWsX
wEfZNDB73I573ITXfcux+tsexozFJXqIbUoVWFvMtGwtjKOvFrYBX3JwhhI+xSfh8WcG2O4Gd3Vb
pTkJFEXZ4v26akdQ/RN1r4avM5MTUuyH2OZ9QegEatiSe7fEGcyJykNxVa7uVhXzxxa56Jwm0Rjs
KYzi8kq1j1mbJuaFIg+ugc4CNIG8jyzc6Q+WZ6VmCXYBu2PGu7quT0QL7q/dLrCHjaQGnUTQ5OeN
73oiksuuVyEjd0tdR7Am7Y7kcJMcSrD7+wMO1MJo87Wf5WsCfToa6Yn9fnqilWK5B96NozyInn6N
Jjpt/JV9kEKpr6UvbqgFGaRGOlXqf5RRxhNZLZR9+WsKMhTQz+QZHRucJ9uR0xeWPJRT62jZXuMc
shzRe8YOQSwOXMkiSE7XpcQCWW+A5F2zzLJslHQs99sI1P4J57ZLdNCSgetPfqjUkVfvoFJRye5G
NLxvzew+/gXdqIlSeVWAk2PC3Oqa7iQofi9+0oLj/qZ420lM9pvjHBpLDS78dWjt81sgBhQdhlGO
TReIa28Fzb6XbDKfCPm7xoP+9luCWWTCjI9KmBVlzoVHKj1xzUEhuD759nr/g9WAt0DBqI1OTaZE
nVI8kKfLO7+uJ5o3azvt+B42UZoxortzWeBsntk6oWYjYa3F36ASvpFhnsqBLn/jVB7oe2AOje0/
Qb+N3Awq50lCr06cPmAFScwlRejGyOZUVUpwlCuaVlwi4ort3I4j0RjD/8+FrJx2eLpVkJN9fOuv
F/NEX4fRdjSU4BP4to/b9go6sxUL7wuVlJ/WMEOfY75BVVB5IppYDJ4ID9KY3WRxaG/XXXWuNSL7
QrxwwfqN+IjWxUwgSY2pSTx+gf6CoxjZ+BucPfg1sNzdeAK9GLasjh5PmSf+GREpXc5gsqUZPBsi
JoTjj2rRGW0rmDIjNsUOlEYoVA90UgdRWS7iDFrEb7NA96ketyxXh8o/K+w9PGj6U4ty/UbKZoTz
4uNajswuE/o2A3sBzbqA18zCKh5ECdIrDdVdja9LLCUR+0rEimu5rB1nqZKwbDZWjyzsoYiqCkyR
E1aapTkS1U0FgkL5u50F/Io4ANjesR2L9dYYwITrJ4YAoGzHRYX9Agicfl2kqRo+Zm0KsMStxJ62
chiJEttlkQgXXyvqnVEH1/bwDCzE/RfpLJX6Nq76fuBcqvRRDImC4t44Or+x+qXaISWD/oORs1mY
IuhRQqXv3SuINKbe9rbhxHcOAbYThfI8J+0n8EA5r33WCalwdHQccg9u3LZa1EwSM7lqFvecmzM3
iJk3Pzf758i7+LnBD3LFlWCgGEJoqdOgLeCMsD3QXgd/EtX3aj7IsRE2y6I7H/dPYRHQATa6WfK5
NQ3uDy6UbPX9Ta6aZMm/vNjAUGn/T1nZbBlCDFMsK4p6wY5RLIsl7WUifJ/y85/a7F8mod4s0w7X
gSj0xueGY41XDrh+c4eX5MiIkaTgToITvxdQySp2H+wLA07ZXI+e72HqXWGYJVvwp8LJhXlw/2rb
J3KgSfbBs0rrsesppAieFCUsNx8DyrSGRZB9hQaYCydapWxUQnnEHMfSYWqf+7WMBPox3MjyMS6C
peXqP+n55UdDv7KM7zxqgecAkLKUmJJh4GPJK+zuQ8AOCet+Hm8aYva+vvqu1ZSkS/6H55/k1bpB
iBY7ga7rq6ZVVSx/FAQUhtZwXDdH9YmK20MD8mCfRjtTW6w5XH7TC/191W6dn8DnIFnrgXGWC72W
ZrQz92lrHqWUbmWSoUmfknCgg9nSN+RZk5/NYmD+nuDSmWlzbDg70R9auXNmwF8p893viYtMo+vM
/u3yWLitVL072XrIDKC8E/yKK19TeJaZ6U3rxVThb/SUbmzruFLE4Rq5QHes09lI/3BxZhN+QSwc
aHuI0lnCWGSAxJ2kPht5Ww0Ldd6sBFoNFgQvmmqMPdw0reOhhsdypFUwsb+rhd0ZYR+6GZt0FFxx
LpnVJHxDP0QCHhHcnEtEGADpJlJEdqnFXJ4HtmzsaeOjG8CWqCaKMhdXfjDDs51VLGYawu0UsacV
7j8C9mfdyWKFykYirUog2XaPsO0K1X/ImtY076T5NvcgohIPeIa/gZcsTk+cQEolmETMDjmIGHKK
TKZO8JkHzJ8Zy7MIXk4PAyQESF1WGE/ogXzaU0NJCs8MXCR558LM5tINkH91bkZXwxl/oKcSwxiG
cGb5/TTO4Df3UY5ElgpwPgXnq2trZQHke01t7FtgzRonVUVU9aFZZFRzmPJf2jRolcjBQb1hnHr5
GemXc4X4fEY5xz4YvX+aclc1hwGpL0AuWHLH49gqgb9rgTVBvBWQEjwFbaO+LySffFw5HTQzE0b8
NcMzTpYbMllS9FJIQiWBUBxDVf6L58Tnz5L6fonl93p7oP7R/fYsmgiEZ/D5DByFvcA9T2EzhhfG
1j26cqZOB3Fo1eORwi8OBcjbH1nWxz7ZrAVxDnEIOIRL1lwLfRchY7XSYTuNHgFwkMdRCWCPQPCT
vCayE+R8C1U/pe72cBvqAFj0IK00AP8tY5mEToUaAoAv8I3+ul5Dn350WgJwPcfMWinW90TbkvFq
reBRab6e0GYBA2B8VNawP412pYmOIj2wUbQUUIAw9h2Kas4/NvjyRctEI4OT1GI7gDZH/fPEgCb0
vMOuZx4HqTXKycmaRZVaeUBOMQFa2qql1PEoGhAe+F+oC7PtVTt3Jomkxbo/YQzFjUTKKAP6Neey
BOYzBmNgYHq+afUKCu+Xcxg+5aTIAQkdjWm+YT5O30bLPdIBJYJ7qY4bEQz3hu8+y4afrK/LQEtA
xWDzXa6wjpzmeWT4SlhjAEsCe8s1E1/CEpcUo3yGU/fCB5R4/jLj8IHkWR36/dkMjgwE4bZYECF6
RofA1YpTtKiJqwNvunLGiMSiqHY/5FgMQX31YkTO2R5Z6no2hgs9b/4L/Ueotf459OmZZbPmodOQ
Ke660dDOzGblLu9Y5hpJLkzxvRIHWXD3yq6D9hb33ZZZPfpTsNNnuDlIzkaOp8sphWkprWZQ3h+M
SZRzp0alcXCwsE/FP6cMfPfXrZJrKtK3pX8AJQuzzUSKheguUCFDQp7qHedroqVMPcMFKLGBz4PA
8YYg6mRjPJnu0X/7pDrPY0IUtnJafPjHSWL/4CbqwtGoTbRwDv3IA0on7q3X1wmD/ZWw4TJXB7si
WD9eNlxAnFzYesYRVwAGs+NjHyY5KMz7IdkioYg7psYXCWY5y+puDxtJZQwCtuduiUOoGUu1cNi5
HiY2qX4fUYlHlwTWhYpjD4+CWO+Sn0+78hi7f0YvA01O8NstQ4eLpCO20lI84Xrdc4RHaJtPQN+e
MMGqEGk83Gjbap1zYzaBwMZPv5i/sMPDZZJXO7hu9uwnSPddmc5h+sc1P8SyhexUw5swL4Y30APp
0iJT9lUXk2H3xUzYvA7gv36oFlK4YX451rSI1ZFykcrB1NnqezyXkhg06qfveoqFz8nRME/JDkWj
gbUdp2BxmVL3lQIL3uPVtcm8pwRKbXwno/cj3nMyKuGFdbqSmV6Rydj/nL+jrjhDJOdEskRZpLgo
ORkRDPTnJ7M8YnXe86rbppBIeYllAvuuzTKJNJLOJmZOjnTynYD08npsmC7lONLymbKCXGr8zQX1
PSJVyhVfs+FpMvxO++A6jDJ8mzVFi6unHjPPsM2+jGpYvcSui9gOJlMfaKIN02WaEm2Ph+6urrFf
w918N5+qWfPVXyspWY0b1tk+YOdPSeYDwUnuUD2hTr9nuv2lp152YxwZud+QxFSu1jVI7pI5b9Sy
FQph1byCRCcnd4iOw+AzAbQ49mj+z/8p4fv9ps3OB5kLqts8+l0XfPoLbVwGPd/p8FdpYBQpGp9i
AAqE/oPKGFfdTyfblUENdFJUFVFoMRmsbKeC5acCUtvHVqksqw4csRhubNrpSeEvTG8G3iF0eu9+
tAAGTbFfRtXgYUEtWxbHRgAhgBVZ8rdQofYJKFlCUEF1NQOyOCEuOoYtC3jD64jqudhckEhS1Jcz
5UOz6LUlusYtDDNR/SryIEZXF/q1KZgevvKevGOEVaHT3e6gYLSl5YCtpFgY/EczVlupHjgXaoBU
Z19jYs+rQ7S62Bh6jE/zV0xCro/cbBYBAm5MN9rpYoGa/D5PJxsJ7KNLCoGKvoipTc67ybXFv3gy
LQvRKazzcODUMNv6cXzy1N2j+GUvRw9mArFrzPDG/Ab8XQEt7OcGOraqzVSBisg6QGYWPyNvjVl3
PGqxWEP0aYSKsHoADVtLUCvMLFgluAduDq8PMueIyO7d1OrzseQiu6eyDWknDMTGRKu70JfnEKi+
SEIWDLvKz/sWcYmCE7U+aO/IN/hdu4WYGc5vuBWKrq9E8GArcZLrEnORntw/YZ0QrsKI9SjsSDKg
eVgufCEsh3Lapa8jBQIeNqMMSSpQJreyDnNIGAQzu2GYYIKGDFbI65w+O+wz5MZGMxzWwLb+F+kZ
NOxEY864EUTgP5EQIONn+aFrkOON6/e82T4Z8LMBAwkIQhQu4GvBISCHmJpJy/nR/OLya7qekso0
f9PZfeSj4L1H+IOW35MMdVrK8wWCeSbZGaJbfB5tll/FpZU9atsvPz8PS7m+3MMsmSt0c7BWnLtU
BjyQSO3I4SCZHEiNpcztkVS/YV+EbOBkaSb4wy9+4+f3OMEUYKYLysv7gneFau+bC3as3LTliQus
tcAIgFpPQGDgbVJwj3tFnNbsGHKHY1B66gtD6f8ntYGVqxaMkrHYryr+grIkKkOgYbdL0a2CbF0g
l2JyfWshhMUzOd9ku77BxJsZ34a8++Dn/C9nbZb1q5xkXVHuGACmbdCttFzm6TM93naFSW3rdJuF
0DkA2GV9Bt/Naz2sy2pqB6x2KMxBTc7r18ZvKHlUtKMA5J6EtlMJH59h6ISZCEWLJzKNpKJsGDWo
iEJjwwtkamwedkGn6npM06Ygup16sRstX5XPw0HvOUQWDcz9NJbwNwWZ3FyNLtnh/T00bQ1K9sKZ
XpZCGUNPrtPZS/O3uwSzX4lNfE4KHdqtbX+/X/1ElyUkdpXT41gE7aGJnUD28bnbpRbj1YE6QeHV
d0Q+xXOua4vTqvr6IiiaCXYb869xS5kZZnuA7GAqP1aLkV6ne+QxDFqQrXHfdAI1VH5u6KsAjhVc
AQrDl5yRlYbPxMpMN4ZgB3k7aGQNqczYstBlosu6+F2/ILGZLwKf7lXIr/rJjsj7cAoyAQl4D4gl
k7paqP+oVNhFSez8Q13FWwYxgBPmBmEEBAWu+enXOjcJrLHkQAxFEF2rWFo2RzyDE5ZjCDiga++D
aTRRvhvDlLrCZi8UTF5TSG0FRgS+Aa5kg079b0y3GZOqcji/xDR/Rdv7PjSNFGSlvfX6ZgTDqzgJ
3y51HgDhAOKAUT3obDIf070YfqRMNZZZJO24+TmiwaAQY/mbrb1U+BOVCTpzhjYzu+vNstbJrGO/
HSxtZs6ufVx0qXIZfisO+0HbaJOagBkHthvRwcyvzV4scHjkX7ePSC8B+CRSU2kL7eiubgee4q8R
bi3I3es/y67masApHXvDeAAzaHlwpkpaTysJlAe2Mhn4MsoVscIGUQSC2t9eUQZ12J5nOF8AROjg
ys2tt6IxTn2KlLALfuxxfwzdMBSyY7lcnwnNma6Dbw+EwFQ3pproEFj1FPQUp1/wLxKc6mYlnjM3
/owBvssyQtzG0C4SsZjTl9ch+9XrvOAz9IaEkVn1gXY25MWQ9R6/jARUaA43QEzpq8/pcxzdTMZB
C2OfbtHR0vOCjBwcP7GZBMxQZklPjy2E8qjrIhsLQ/t1RPugGCE5FWCJeVj0HQNE6swM0uaRZ6ao
pF4YqadBgUaOaX1M6ssxHbLp+U0XMourcC6Q681UszVbMn4fjFqiCYXqaCMzDdA2gtNCdPVvGdFR
2BoXEcR5j4wJ0qQGG+CvzmneHeRddRvYVq3oNgGaIkwHLz13pPNgZMmsN7KTjC/8xzofleJ0VTa9
1Pce/yUxQpZpP/RmIaO2ZHs9SzygsEE+wseFv8pCgkpEvQ3ZMy0SQbR3N88z3ND/GO0ssSeDz/mE
Nxdty68IEOsigNXI+b0hvZpIUTzfy/20+RbUZsIbsmQXq+PeTJ0mFg/ifCzhWJ0rmcQIQ7ub4BUV
hZtrmW1zHEaWxmTVtvQVNdSGsY25BJy4eVhm0s2hChJJs6tc/9p891vTbp8Eo0ClQzxXxJpkGQCc
/OC62GwBJDnYp2d+hm8Vil18tEXHxEwYDgI4ejzb8pnMpFrcXTCw+T07zLursOGsJ96Tr1OvJu1J
xJFCa0eVyn1mdggTxAB7MMZlvTBWJepxK4z5fng0lBlOXn2wk6IB5BYRi9AhknHG5IkVhNfv2g/v
gdI/jf0EAgIXA0vsFGpcqrx6XZyqIG/3MJaBYxrKkrx3tUJ0WQavUFek7GYW8bBr0Ti3IfBeZKXJ
0+IG88XzCxagYT3n8XYtd7psipxLpGnv770IH/vKCCuLla7lmgIY9GhX3bC+WDWUhZPE7KSRNDgT
q0Z0mjioDcJUdUt5Y/q2TfCXCA1gTtwslSpXw1S8dznfLEqtPF23iLLAI3Hir9Ts3Xe1hWn4DTwr
RU3psl7aiBGZ54/5xU7Xj2/8nmHIV2Q6K5aQElr05KnjBGjSFXYnSojNVgM8h/FCYr4sdqa+ZF6M
Kovzw99WQaPbMGYRF8VZqzNYEzVEEC040XC1jX0i+7GC6fqTfT8zNMkTPjH/7IJLMNdWqm34oSoB
dYHLb2aodKeTpq4QOKQGG+FrcJ9DvsGUr6kfkl/D9O0yRwsyLYKJHAkxRJzgCkzWSntZkqPOJttX
1R2PX2PjBEGr1eEEecL7NaaA+Yj0yR0aCMgse7JfuxAN6g6WpC8801UHDPa9BbeNx8d11II9+1T6
SR6pOgx7MUgOv+Qnqvc7bAjyaMP2n02lhibyh3NZguppAUjqqCIC8ro/T7eyRSxv+BKdDOAS7/zP
YFlxSdO1DGP+MPKsLXjZukA+lbfr4d4SoGHrXzybrzP8MrVZecyHVnsf+9V/C3nfH/80Us5uCNJQ
BHonmhIsOqV5WsFjE5fEH0O3VQAjnOzGL4AtUPOsof17vO3Me7CL5acm/8roKDYHLMqlObng6dpW
dz4ltdxr0qPZ20dlEllWkXbSWD/5ItCSNFJ1gcyE0c0ZlNcHpAn9XoAkk0TnDRfMTEWvFWfw+SLG
nU+uE3GxvnfsMMFBRiJ7AzPKKDiZj8w0kwWO2JeJ5fw2l3GRQvPjikgRYx3iycPOGQvnq0j9GhE8
tKL7BjleVDKGuTEpF4yI762UxmJk1hcm0aAMQga954W7wwmd5Du5JfGGb6dOTNWUhk32UIe4lkK6
zGCGq8Ha7JzyOyW9SnBje/dUEt6J9dRv9O3VMNoCTCCPGrBfdIeEMIDbqejJdxGOIDquze7j7n9Z
0iRO1BSNuLtXMSfmmkf11Q66PmhLlIss/HKMmqeKspvRZp8VgyGT7j8hFwh7OU+zleA2Y0nRcdd2
uua0JUc8xVBiImJxrPZ5e+qOz4HnwJYrUG1SNJmCPu6yAAKqSqBGR1EFcr/n33D380nJlmt/UZfa
wZ/TsUc+QANt6UNxJeHptbavNnSfDmerKz/INO91LqFN8+zlFhnH1JCLRbhDS+aP4lPcnggPCXU0
IXfeyWBSprqNxLCfdBBnmFdRr7eDWuE3TQDOuLR9W9dxk6mGVRjPtdeTmIf1l4CysBv9T+XqGFKJ
zZsYJXKFBCrnj6zVCJFNtCFRyv81GDupLJLgDEtMjrt1yCntS0i4qn6t38codPTyuEYXZIpO/Tc8
j+bGNmJYPqvlsXDHqpk3CXd0ybn3Fo01wa/sNlWaQxQVhRw1ZOWzc1QI/0AqNmwb8i5LzF5GB+sS
3BYhWbb2RNNRZsuRsdF6poOy4wXpQ40gAXt9s/UL9m2t8E48AkZeiE1AbQe93SFr9fiejNRojS1T
D66ut+WBuHZ+b2NiRFNgl36vuNyQNnXxbYEmcCEV9oIYfMT3L68sDuEufKb6BP5JYEL5wqjOgghV
u37VYa8eyIfHgRcut2BkxAnTvxhxQjbDKhyO0O1VWVAIFG9ho8wLyKlL67nRwsGgxltk9Ayreqr4
jydonBTc9Wa3w8unWhyrW31QkyrRsN0neYT4QnCklKb1K7eo1yxxmDyyKoSUinpZy902Laz4Dg3Q
3kVGZDPucBWsuhKpUDgNc3JVE7f14lysx6+MCeyT9s+XrbN7gLQKt2ksmgVHIk535k38U4JQu2ch
iZC2cbEdXf/O+1msiS3IIUQSNbAqWXgswAqgkyRAW3ZxbLk4mjmaoh+ozBnnlCbFX19xYI7Lk6r8
h8M6s5nlbHXkBQZBZxylQE+j9Wd+XskKFNsF3IVCWEoERK5Q1ckL632Dn9Hm/xUB62qTkluEliub
wW53041E+DPduI9LShkNSrNM1or5ax6ygFiveUmBC6i1ceXUOqD8DJ/XpJ/wnYowMcFwKSDm+76R
kMhLTHH1Bl2PpVb5xHTj24Z4GqgiRaHKFGcq2/KZ8aRI/aObyu7EpuhCQDUnqz6J3Yy2qrSBeos2
s3Y4orgWrtrgr1p44h6XfLLYZyue26krDyaSrbh/Y4oyspFHQouhzNwG0H8fIRSrMPs3sZtVTiSv
9Ldd9kWRckLMONIhKdynG1j7LIXzsaa3zabWzQpkxFXAQuXb3djbs0RP2BzrCHIiehfXO5/yfCvb
A/6uHt5B3IuqPzk/3xtwoXxZz+eozU3c1cdMiGlZVkKbUoO92bHxG0N9oP6To8HBeiCeZcTNPmc5
afXhSMO1VicZ0euNVw4+PEQPo53n5CrKKFCPnMmw+1LNgCvGdol1DhOi/MUKY3DocPKCRmQICqDH
FGOSqlTWUgj/bvh/a5VceE9E3bY2DJkKlXqpFGi4xL2hp4yHGDzFSTrpYHBipr6TkHgLuNFgO5SB
vSGxaDIkYEeALxgz7aB2lQo0QySxdY5D1UsdByZ5ZCFfwn5KbIBI9ZA7P8SJMo2I+8ifs7eA1427
TvPECq+N9EZEhdy/3w4ng23QBK4lk+GCPO1Im5lCSDZty00DMWK6I5tnbGDlA0bTaUWuiXuUvJ9f
Qiir/ZdtcwmGHSx3FyyJwyB7Mw1751a7aRsE8rCKhhG3ctyWP7Wx8h96UM29r5AgHF1Jhm5Pf5W2
LPXBxdwL8pSpLarLqdbtFju77Byl4wzvcyuaVluOBA/QPp+B21reE7aDCFQbLS6Cm3/Z1/VjkDKq
3DPjeKvxvZwmBOwsu5G5NCH3xfgIykD8kKyYxlkVupFxL8UNS9IyMsKXpgLfx0yL3fOQaO1v8cfG
m7xUhnHeQeo1OAxz/J+UdL6AVwi9XFFwRN/vGVNwhcOPg65CXjmVr0Pyv0tQvBjR5oVnv5dhR5yM
jp0HKJObS7Zn/FJFNM7D/AsFGzA9q5x1Bc8mRkdLfyjrHNMQwza6cYaIFkXq71l5eOtSBe7TLGWr
hyg6L0XJz+VeQzIB2BRJSKrNamIDpa5W1zY14Rx/n84/zKYNBENL+vlSk1+QaUDKO/Pkl2Zh7zFO
s9sCcNPGyjQ/uRZgxiisXKNAxMtK9ovDbMQrtJ2SNPTuSyrRIP72iAmZBwDSNrBAZ3MLPKgO+xKc
hTO7xMW2viPy1H2EnSGxdCG/kXvcyi7SJOyvogvoGYG00YqVnybCdaPEahGu6H7i04RBJXYm/Oq6
ZH+GPcDU91+f9parPYqCF9zgoaSI2WTDRD5EdEM8CixAfIQaVwU70f7fzP3P8RxV1Pmw6Cp9xpfy
apV2mwCaLZr06VJWaPMDh/OKdpsClPtICUBWcTSavBthaDHj5upWiDdSCxwx7XqIoJJ40gimsVa/
tYx0evz5Ra7UXGtTKbK14OPeybO0geDP5BSQJ1C+ytWJ/KmDN4Lu8sLIFmd2byLYFdhK5AuKv302
SmNgY8gSd8WP/xOGO16FM2SZ3a3IdetEvJ7Kn5wYSdKDPlM5CWusnZqbg0ntCVubF2EQ3IwHkQrs
BMtjNZGE9xm1t7TM/HXwKhhNsmYl22zXxk0ewzC+8Y+yAd/T7R46GCNGwTtDZfLND5Elkuc4bM/Z
KHdutcR12CkLpQSw7jPWQqZD2HBkZ0EQc2/4JlG/hIRgz/ISU0XR8HuysqIxnBEzVGd7d+SefDv8
Ol7HoWoqDwCFrSMUA/lWjgyev2EWyK3USmh++YJ2QdWhWytDZi7OUlaPthRvQz2B5EjPZeJ1DVg8
WyUKZKT4a6O2QU0x5+tNbeQgRCu0YdkOP0JJ5RqMM7WAJJxmurPGDRxoVFYqzj54CHgrSS+Fafij
U0DccvnOwR30bWYdIrKzjqocvTYHd8t219aWP0r9iFU5/flDzlvJlzH1Gqq3+V8PldmyfUfT9CPS
hbPKdG7kfp0JDXJS2DbqqSuidE7Rt3RWvJR1VlsUB7bWk4ShBFsuBAKOLjId4PwR4LTX338wD/h1
ofGmMe5Jj3CBC6r8s7Pgt4bc7efEmiLxymtCxz8WEXjTDDulp/eSEyVuBEGJPQ9GQwNwPua0n/kl
ucu1lGzQnnDqQCdIYn6/NnCoJ/0HsL2Wp7RL2fic8HK9O8M8UQkObs507KpqPeol7JmNGTX13Y2K
0QS057ZPmGZaonymAphWLcAyGuEHydenCDbQUim/atL1NSj4Z05V2Pq6LyLer8o/aekaYCuEWox2
c+jvNK0Nqo0P+nkZaYkLXmMwBqscG+00lrDDaYIdHI3/IrbIkpHsUDxDmNk6G88bA45g4PVa5BGt
0haxkfksMtyjcSttpoPcym2odgVkiRvgZGs2Fg6LravHO3sFUbYq0Dkc4Z9zJn/zNZPwX6MueaXC
u35gQUGLjTowv9DNrbRPiY//azop0DC7ZPK5IXIApn+zZo7j9YdYHXLIWjNotFq0eGPz5rJ1WkvP
BotlcemeZMJLYVsUnc6AAT4oW3NR/SwIH8Tibi3eG9NEc++RlMdUHQvWpKOPA1Inmnx0tZe/EPiQ
+JeuOnSS+Xlm7iYXypPMbIg0dwgnbaTlS0JHPb+dAmQY10TZ5/Gr3tfc+6hUVsFDWoBj0ldMzn5s
wY/0E59cURAyUTo6/JKXbzsa+lT1xpIzQgK24G8K82m02FLBB4EuWIFZXFUXv0xuyo757++MkhZY
Au+21/1JYkxAoPQh18jowDCVgOgEr0DFadhpDjKJlTOijlxy4hXidu27IVLpYqvQKuYa1wsmL4Iv
5dSwEE300EO2mZwIaeKNf6eUiQdrmODX0uXIpIoFI5hT/HtQMiULaaS26b4hNB/WHKpAa8Sp4Bzd
240qcbvXCljpPyCwsagmQtCidNK/i9Nqg/NIKEaSC6qnE21JRjx+anxgE/spemRBiXAtGOsMnY6A
qPXIzPpvJV3mSBtrxjTHsUTkEPBh4n3M3dvo/8Ivk/h6Jdi7MYOE8EekpkXZTwl7rEW2yZvlOkoH
EkIJvLZoMDsC0t2hws+eErvkFryos7tIPfJWV4qQwdYw4/YFf3ht3KunJ3XqYIpZtsFiA9C0A0rH
M5t3+wCM+CA4CXz9WjOwApr2al2+PtV6JYBNvmrtnK9mBEC7m+alVxPVZyXAqeQyIIs48suS21vR
NE+tiV7JPCQrlrK9Ryi9JOMe9voPXgP3C6GVl6AU35hfuceDq+d9nl0nILj6vYke7s01q4VweFgP
evT/K6BED2AJ/oD8oZ5e6iYROL2nyLPxFvoyZ0Zn5v/wXuVduS2CHs1LsRKs9dLduu7qgsGiSBYp
hLDnw2UF8W8s56R2M5UW7s3Rz8/UVdN6LiIRkzCiQIqTzJOOMuOaH32zA1KflrDnz7wDWKpdKqxM
fmdEzzGtauMd0nla1F9s19EziqqJZ6NCIOxDTE2qec6slQ3pKgXZj6WhFds0E4ZVv4nyaAnCoFgZ
aKX3PAhqhisounqhxWNnOFun4gDh3P0yex/1nESUhhkyYUUr1Y9MFqhn0FiBJSz9J3oeVBmpvWp8
vi0/7AThZcWkr9mOew35txsVaiZ7pjy1ejlHSXyQbomKGNMrxaIxzd2zfSQzYlPOD45Jd8QhicT/
eXatXHe7SvLiXpAET9LlzsFnnptI+5M6VuMkIYWtg2F4kJnlegYjv2mwX0wVEjZPpNzVcNO0QbNa
an6lI2pETG9S9UOrKkOlIKrojD2kGnBitVaIiGUCElhPLzIAXh673FeZrX0+yfW6lx29QsuyCmsf
DzFcJNanygwjLIQbHvQirx7lGpZh65tXXrHMmH9puo2aYIuJ6czSBM3TZAQv9m8xHl8DnOBbfmyF
XF66OSCXTvBSr87iAJWSlSM03BkCs9h6STh01jgmz9dqeJcPI2QXeB+5UUWJDT7Fp6lS7SgfWslH
d8Yrxm4MXG4b6frUNQS+lpVmg/jQ/XXDYU196t+isqCEaMZ81gO00W+A2gclxWSM38iN0X8tGMsw
fwGnpYk4PJPxf4N6dN32Itk0UR69fDolmfNqaBlwOu3I325CnG97EFr4aZ+nbyFnqqtQaW0cEFXt
CiLKanvPg/kNk442yA2Efr3hY+FFiOBQfQlt6VQwbMTM9Zxnr1aj7oWslPRPIYBN3ej6611D5dec
2Bv0uKWlpiT485Ybqlya1ulAA4DMlWJeQ5pnJ9pg1bkIOvlfrheXYtYuT8wB/ZDRADYRJ7d37Dfk
dTbCxRsPNTyfH2R+fICLzdNlVlkJR0SD5aF+DyH5Olqki/Yk4W+ar7r4FPR3BwQwRCodCktMFJ5V
Gu5QWCyDomsQ8fgclfFchyy2Njl/rS9U3rQGkgYYHV1ZA4jWnQZ4fjxtuG3WNRZl8xPHuSeImOo3
lNTj3Glr3JGSAMuxipU3fmjqUr0rjBTbjm1+snof6VHON2LV7PGL0YIrDDf2dHw2HXfMxBLtEbha
S2emrq6U8aozGfSZKGbNX5+qw0rc41r0QtuDMiGfLA5uBHCLxZ0oI54WQbw029XraqN9PnTbalvx
TQtbGsgtnvXL+HJi4AMFMIJBdlJdBHUugiLBGl9bsm8+BlpFMT/8ZXwjin8cGP8dWb8wczaDw3e1
R1aPbq9an+f1p1OKDfk3wRNHiWF+Bl0u4MF0T918fHA4Q006wVhpzlUMLu1qXSPFXRQmGgun26Cv
/wABzW4xFZxMgq6/drCzIsWu+rzw+941TJ8O0YkfJ9GET3HVLRl3Ut5rnui0IEnp3EqrcR17G3EI
bMnpHMoJhleHBy3ilpsqK6eb9qAZ6atPv4GGUwIBgWLW/XHwTUlerSgnqjUa8aX2hAdlkWOv/7Pc
QxD1yfMa7pAcAC26pkSVb6Pz0pseYTbwjDalBchDueRbZ0Kldf/S2uh3rzXqhgBa7GEoTVz23OHB
Mpk82WYioYwYXQyeJNR1Koij5DuzeHfB9d0GF5BR9wtMwfnWAmZ+TMDPJIBizCrYXNgXBXoQqP+1
7n7/4RZXyvTFFhAwVLTlxpweT5ee1D2gDxgcdjV7iJpG817NL+iJ4TV+d+FmPdcKggHW2Ig7HxuL
XKq2tXboDJgbf3+2zA11QhO3ifutGCNDMX4zov9QSFPMYuBnj1oSloBcrpc7mXFtTE9bQ0CoHrTV
gau3+kk7mzakALCqjwAKMig3wBYDho8ZCeKqL2IDqikvTn46hpQd0PFmX04xCvTov7WJ1FObcCIX
j0bs1pexeYu62d83TlOFDUkECRV8cpEhGk+6BDKwTmdX6AyU6dIUcEG0uUeW+VlX4sMTHUu29wNT
HApaWkvK7e4Fh/KQo+Nt223nrj4sjjXZtULwrpPmB2sfYu/TYIvhgpLj/cX2NYb3T07ucTlpJkRv
QRjgpvWichbQp46kCB8AoBfBui5voCBdPxUiyKQozstN3sZihMZAOp8LfN5gah+hKfpyoqTeQubi
Kln3FDZyWu8Ht7ZF0T/9pkP9A/Q2X6/5YO5vafswlQYMpWTjWCvZY45BctQM406tYmHghNfHKlDB
rCyrBPrnyCnPeRH1NWoZSXvZFvVht3gvRyTsSLyAw6ePQlYjYZHbRZiePOFHZp4K9G42Dim4wlNa
7bE5mpjZcupNY+shl3JGdQYMMqCwNp7P2BBrqnbfQ0v24VBsSHKzuObyQMVgCvJvcyOVF7fVxYl+
Zys8ReetHzcy9C+XZONJe69qcIw/iwS3vDDZ2jc9WixxXXuig5WXkvBW2R1kk+L6LewAWX9a4RPN
7XFmr1OaxJi+IWHXp8ew2Y9vACOf2VrGHtw+yJz9jzswXKq949bXmhLaEIC1mgWdFCZAWq9D/Xkm
Yupv8hREHDA+EFjbDVMzudrtE667aV5WE9QHX98m9KNLjBnnPEgNCgbCM/kJmRFBvx0RRwvLoBEE
D6dArfQVwsx/IkB77ygT6C5XhRVEwDPWiyJy0675dkvnefq2Kr1K0f3bm5lDek/4hskHGzhVnoUM
0O1W3pFRP/Krq2q+l+Yadbyblxaip9ob1GEQtgBV2/unUzscHh0FdTm1QMpDAQjwCfyMvf8G12Yd
NG10bktzFHk6nFCo1gLsMRWRFkFULjbkgr5TswDdMdRoNpVGOKD6ypdCYqK0Fm8nWmweYTrwU5Ux
Ti+28imaaf4xO/Zq+XWJKVmtFLi0MRRTruVH5i3sIpMPuf57RMzse7bmft71LCh3JyM2FbD4G6Bg
dEO+QkNaR420Q2PzeT+Ol6wk1CmRQ4ytAxNtjblrP5QrzWjNIgPgk65H+7CjVyGXahTCCXkYGjZ1
Dw905ACnel/1P+UkV/dVzIZEdhREHzMEMDdvKMW+apgzIiNGRItVI1mUxTOoSCXxf5xcCVt1ZmgW
0Zpcf8qr+mAv6RluzR1AQiIo47SEXoOfsijVHbDQWqiMYfcOy0kkBgm6Agm1bv9O4RKXn8zXNCNK
m12CPGNIaR8oj71C50eCnAikJ/c0TfNxS7Xz95QedeMQt5ftBJjBMwYXbA6g9JTkC4st7entzmky
3qJYyZAGktRD7ETJq8WkqNAZ9GwxFTEOhHPtgOF6KsrrBBxKfW/RCxoxK/OIChhrsNJPx81NgY5F
jF3bH+uqssJxQIZkT/XjRl/5ZR3M+W/Zy2Tl+z5VjDRXSiJ7EBcQPA8OpLUXDtz+nzhrMxTx9fst
A0e7Jsl8RUn6wEH3iWVLQ11s2sLNcU6pmqOL4+qYbr91Ti9feSDA96EPud7gFRC3Q5ImmH2G6PNi
Dn7lw6/pW3WZ8I36QlZBmvMNjnaEFr08R7xUrcMY/M2DOCJWmQ2o7HlpM8ScljNtQfg9Sf4iv+r/
pT6fjFWEDU0zW6zRyzT5IKlFzMff+M9I/5IY9xHXPc4biYPIcO12IKM15yG5IFY+Z5k1upn8HMj/
SgdrH3Yc3hvgWOpDJk7szlBngvCeh2SnEZF9eaqt2mN4HtZBDyWkieop18X41z+CmAXOv6VqfNhs
zunkkHdNhxkZbo0aixqqBRQHknBqq1ygSNd+fC0MZ8kMkaHUee98YhyX7wbLd01Rdq0qzbBIXUFD
GgY6bhFSUYjoevxLob2UmVwNabTrcHMTg89d5I4YByvqttFdk2+3c7DzGCBuULpOFhBRut57uzQf
rPgGjE7tS+Eb73OC4ula7HNk0frsb1uXJxViNu1tHeHNbJi3rt97Ak5nboM22y6YwnPhHPU733uR
hshpKnVPkZsGziLxqPt5GTK6WoR0cEEsRJxpDhFna/bOFhO/iBodxqh94TJojqOW5zVTnz1bpFXs
t6b3U5v5Mgsp4Crg0GMYVdOgtL/aOaRnLa1BGyGcJIZG5d8F5uMcwWrSryafVF70euQt54gD87e9
1VuqAISsub2lnez+r8g+Dr0MeahkJNkoWnokXhxukFIf9wcKIZgAp82W5R90aY1GD3R47jA8CIfc
pY6H5TcstDJNMjwYgrdUMxNF9hN+4fSgP3D2418addxgYErYclm+P2UvRp7v+Nd87EPYwWh0XISL
yBa/YTenqPWKWKUNNitwvIXDhslc3N5bQ890/GzRgIEUfWSoAiRkRxkIQPtvbhuw+wqJuOtYBO0Z
J2xFxRPCrDdcfXLeIuLIWIX0nI94GFE7QHQYgGlXa+W/hsNd4K6yegfMtXHLiGT0dYtkoetGv3r0
iAe0Gc1CQoqKHVdqQbZFW7OwrBUrHk5ZrTSZ5Q+5O7XFbvbNhQSRFwAhU2tAZ/07xRMrofihtnzS
64xNQ2d4jnK6rm3jlig3jGWg3duyiC+aTOgdafp8F43gbmE8gMN4/H/SMEfgO2sM9NJKteLwElNY
g2TGbK0ePidN5wzKwa4+5LEpWRfVYd8Ai7TebjS1D36JbVOlufwoSf6O7UNr7xVe4KcOl5iUZFX8
u+1lYnEMxSzw6z2WEc+AZ2e+faPz+iFUNhDSESp4yVSOPCiN1SXhZXupLgLYNyn+2i3dPiBZx44D
Z0GsnuLokJVc8doj6q/cQwzL4g1GJh18kXXrf4SaBlPj3EezyExDcei7xTiGeFVobn6NgkLsPiXB
d5jmY0JniwaO3TDF9Vdnrd0VILbnna8buPwrN6D1pLmvXy7sk8mu3zHSI364UPCesZyfFMuu9Jmt
NtvNhdVKJpN761x1ih59Y4L7kFFUUbyf3CKZMqUUdpkXpNHFCbrazw+0oV1eVdcZuz1v0kx1rw9d
/DvI2Mmekpq8eNt5Xv/JUkUg7IqdtbaRfhPtUz3BRTIMbgyvVvEdOwQ9SiXe/XZJFHHRKx4pJOvw
Aws3Fc2SU6EMobvXbzHIAbfj2/NpY2bL9x9pGta8CrUFpUj0DZ3x2/snnLPXdAZ48dp1s2pUn4+1
M4BMLnLP8hGoJQG/gpB+thDY3/40XK7pFPujJbZnCX5yiRZ1eS7iQhCoyXvg75TmcCcfX5adlyOn
W0jCrBYBd5WuItY2Fz7f9yAx3wAFhedaIC1v6jBGRD5PzFMM9GnhvPvvcPfrm2djSoOl2OFnRP3g
YXddpoQZXFkO0Vk0pcniYeaw6QDKV9xxXwEosZhS55yXuujRxt/7GPeddaA6WrrPX1SbC7p9Or2D
X6sfcbZMJU2hiCxbsqjz1DB7uyPCPzN+3Ds+2ErdNrovuMABVm1k8xxqMvBx3OLS88P7VU06obhq
yUKAjwA1wYX8Ml4mZHtc5K7yRZNgZJk9jS3ycFZpdapuIB+QxuLmYWCw3BUk5Xkblp5HHeldDng/
Ji/NDeyxsY1RFgnvyiitgLULHEE5dlhUEGgOX7P+XydS0sW6ExeXNzoEt0/3GYHHfIUTBmjK+LES
rHyKBQkE9VY0Fs2Rf1PMRcNlkdKemFJF6HHQsKh9MifGWpY5qne3dXz3eMqup2yWgWdMWCm45ZuA
I0rJjqV3QG8qWkG3WnNyfa37ce4Kqyfa8rWpMPk09XNg5IbFo4XqhVlW+22WuvBotEF0ej8sGgD1
hc8yX/KVRGqgRZcZWuP0M5OckxlOW9ton+rTpL0cYLQdVI1QGESXenHOEXiMJmj3nivKqNBjBbIR
0xBe+9h3fPtfZ2oDzca/EURjeexVt19npM2BSTldg/UcNIy3dbaLvjFJCAZNpY9wuX5bYi6PAC8t
pl91X3w5X2tts8z6ezflAstcH3n5CmPAAwsTl6WJmj+iOTRTUPAXhCNvvzLP1niXXKUOvvwlZ+Uc
mxdMMnLApYKVvIjqR3bTsydH81MEmLaTlSQqt7rpgBdTBSB7mNFRRH1v+EYqgpLfQhDmWLj1mfpJ
DeOAHT3mmpu0Cj1ZWQ8svcBYVJt/XbAILDOnyWFASietvEa4Thqk22jCD7mdp1uGmLkkAW0zPEas
tU7Z5TdlqO2f2cHfRW8oD4U9P8zuAiBZ3Ti14yf2TIec80OdpITisNL/r6XjH1gcXX8qrJ8IQ7Nu
rCavpL6cGmP+ggkdQYcgst49XWiXo/XE43HcdhqJgFKu6U0m1eR4nHZtpkqlKrB25e7N+P4rFyHk
f8bwzaYszM7vXZz3pLtPWvgx/vSvCb9MmeR5x3TyhLsqTBS1MjHFtF+95jFFYa6J0zs4qW1D9XNZ
N8V86DLsdlctAzZovFxSdyA7R9PnEI3IN4kBpJa8enGCGwyMBcXI4uXPr37jgMz0SS46Hp5xVAVL
5eRtytaOP4svERoYMGRiddW3DGrgKFAzupdFBdBK8JCGGi0MJfOe9lORMAl7WWvuCEchny+cN1cN
T/1GOn4xkDQQgAxlot+33WqDoTGvGiX9IYPe48mOjxqAyaOC/l/saG90+YJ8cYP9HAbSKqM3WD2e
El5uVAUZepmwDJyZhB3Q5nMVgj9a1wDbpS3clt+XNI1Xf91s+BH7gjuMD2i+1f7vU/OIECkoaHDN
Kn6lB2kuiLFOQoFuYlNkMBAqtX+DxM/XzcXj8M4ukUOeNLF7HkmDoc5TVgEOLg5IZcTkAPLmVgDS
FHpcOLWTG/LmNeFZoEdd9FWinTOGvygns/B98coMdDAhQ0qZEg7Qnj2dbcww7wGyCWJzhP0UlzHr
uzv0sQVOGnIl9cgvBOTIS5FY9/OTeS7rNYn5ffguvkFG2bmXWFvcHv4zVMGHGA0iSwrOs+RidHuD
Ri0E6MbP2qxXzh2I7/NOVUQR1Mq99brU3SEO9nfk5Xrt5FoMRO8ZO4l37ET/8xIll4lBk3oEHv0v
imc+MJ749+iTpA+nGfCCuaEPgSGTDeSDLrcbJQTAxtdWJ9ZUBJBvd4nkl7Ld4nlvlR+hxeelTYon
kBjxUD7e/En2sIYs7OoUoTNoNAxxb22kDDbyCfu4l/Yxj24g1gTnjwzfzdWWyeHrL/uqK/El9SuV
lULodIcvBTdkaaLKiKcQ/Hu01edwDm+Ae1ffWmnXcj82w/G519CudyvP7vDT0OENDQtZyMeD2Mnx
sQvZX8ZYbDI3w6dFuZ+Lp1ntNIdJCf5+hRebJbyIpfZEljsM34Q3hqCp+eTnb5RRTTY8E6jb1vsc
OVej0/pPyfgeug1xVo4XzRdAYmH77VxEJ+judmO+ycEgC6/OFAOcewkEtPHqfBzjTxFt16yGJB/l
2r1J0bPVQUO3OkecS7ku5la1rjFsHNcvms7hJAo8V09GaFLqy/SJDhdxkR0EfjFDn4qOIwBBVnu1
coZILFQzXMDDI2jpPZ/wrtfxGSy3GL7voFlIvRuIE7cvs1nguN839A47hI9DQdmfhd3HJIZs4FTy
/ln1sO/jGAfH2T93Sms9bgszQbH0j57/YhtmmnmPof0KjbjSzmlpe37pIw1mecDF2VYF1mLE/oLD
Ki4P+gzu6/XnSrrmzjhFXAlE2bB3wIzRDhUNCofM+RNNywNdo12dspmq+FVkHzQcpDXAKpIW88eo
bhUNiYm0N55VPvJOQ/Fh/G/1ZkAnMi1owyPCnPJR7aURsp9C5TXAUuGojcfAGJrdY906etWJvREp
dKwoaro9/f+uCxBbChe5gi386HzwGh+j4paBzcFBGqIod81MR+vpFOTNQuSEPIKkRftZkp0m/9wA
3TVCBBcOO+bqctAuY6gkeATp9YZbLkn8UNJw9a4zApTV06KMBn6N7XYIf81umFdF0ggxHpaqpxdl
MOMx0tNHsYIc8N1/OlMZkHr8rRouPrZ0JEd1zyflb4fCNiEwMP+i8w/RoVY7kqhlJsJACxg3UB3J
fCVH0egNY39r6C+p1C82hDtCdwJ1dtFPam0wryOUxltyTlgdOWKfHS2gFsfRCtIyNHWcU/xHjUQ6
J1/4avGy3MzQSUJGWZaUijSEcFaAQ2HeDI3NEzL6jSlZmMpHLmg8Dg1y92aVqSrRLJJ9Mr0k+4aY
RuieNv1TRNt6F4+lrOopBAGArXy8YiInuBiw10O83D7txtS79zFwzdT3jb3FBVM54gNov9sxRws2
Oe3GLtvkqrJMEtpbp5pkkKu5c/0q39lYkE55NULGxjGhpviMtQXFl2jTy66q/UzA2e7VgWKQRjP/
w35XRx3msB2pUaYFd5POdl7gOuNhSrPDgLJznNcsagQDVD/qfQt+imrBsqUbq4URuTQ4DTi7HdSf
aXuruOGzuDeZImAAhvzGNo/fPgRyaqGzVCWqLK8xW9hNAAfsh5uaTdXDGjD9xCxYysNJJ4kY9x3P
EQnZhNSy3mJ7KdIPFSt8Rph4q/dLSikNLn2+96w18mY2wexC8AQZ4pqo7keKWkbRlyQDUFYyejSs
y07LjkwppqK8eaXwPGZSRX2Qes1yOHENZKry5WssTSB/UgX8yfeACmwiyBp1Tssdk2PFMG2rQ/WM
bMb7NhDeGmtl0hpAyCX7Izj5nOZuSDkVMVLK7650/PXBhCLt6q4m+iTce6m5WkAiAtT2EX2Frr3P
UV9igR7i5xYtjTiOIhIPoUZ9uuB4smXQ3ex2jZGRxPF6qQ4M8YNORNgVQS/tJqR3c7Gm6dIde16h
X/arhimutV1T7z4NxZstMMIVEl30tCdMkFW4VTTy2WG2J0Yf1oc9SyzY+KmnLeCZqGpXkqBzNWx1
LOkckoOOGfIK/+mIe/2ypO3Xx3phiyR7GJSCllyg4h+HiDN5AIKlfdpC5OvnZOU4jmZj5HE4CPAi
YPG7owIPDO3A62XLxufVNqP32IcitCW6jaseWNoY6e+w3gcwzNhJYPuOA4XZe6ITqv5VomnhLDyY
HvP4sVJsh+/jQWwwKwlsSuuSR0QgAetwhKYDo3/RMlUgPA9mBjvE4Lqi0uVvIbKHiBg5ijcP0R6G
J6h/ECC694kxJKWnw2RFpGG2EIvpvvrsLbALyOBAVdCn8cJBv3h3UKvlDoiszEFlJ4m6d8KjOvOJ
dmzKraTy1fDGI01id+O3RpD8cxd8SHKTLN7T3s/tPXxWdgjviMRuYY+WL1C/s4+2UCKbaXAgYsnX
3W/qLtVHkYOIIJ+QzkGVE31x+naOAN/t2NV3TrD8vPvHBohMlx3tE0uSsmQhDprLs4oQrA9mzzVP
QDllp2Fb0+BjWmNwK1TbzlnuWPB7/BpoZmaOIOZPtE5lEz9RWuQDXC3nfKAG/puTcPbX04p2gu/E
mRu/j4wlz5BVpz54xi3n3SBPJ81q2/Fa9GDtnhtqhMEbgrajNiWOnxSkAJgB9ZIkxHnWl9VzWhFX
GEgXJu6Jsv0HUb63AHlFqGkF7BquXrPXMZsMRwWK/x3o38G0Xl6KT4qvhDjKyaKMyKXhKSvQ/5V8
Lf4AwjgQ6z517mmUjQcscjDzSMwbydg2IlV1QhqQE6mrwa69MVAOFOLL+4AkRQwuk1Tdm/PX3pKG
p46Lb4pVw8zvCwwZgscrI6Ye7Q/iu9stSEsxEoyTHx+SOZi8N+V44tsdY/jXKU8XoVqBlTzwV0XK
I0BbDDCDM03kVmCkj00XCnrD6/mWB0AkNmYn3IJBaJDkx7LlNzTMyT8BSqbDLOESBZRxp4bB89r/
JlS6mNO/qzr3TzCAcWsxZnZDi5/iIokDVcSnyS3UKUfAZVH4Y9X9Yaa/pE0Bn7ZVuITwpWs2gSAt
8Onee3M00v35RsthYFnyg3Wv8duD4NjajWFwHJsexsZqLtWIK8iYx12B3pzdkYcmiqjirwiZalvI
p9WIxEkZZuzluzJYPNWaFRykjNB7rT4xSvjBfysy/JPY12kVVwIl4AVjMVk0sPsC9GvbT/Wsfb8i
syV+xgAqB6u6ss6MqFiZ1rqKgSL4z51ZPARCZxrEebAfFZjEpr+tMm/jOq/V+C0Be7EAPg39rT2k
GrnJg15d4Vh9df8tFswHTjNOAGH3lg4Ix70pyPXJ5fdqDrsai+U5RDmWG+cG7VDr2R0ZFQ9rLLlQ
h+y3mP/exmo9nKfb1tc4k4fJBziDlWehK2D+icf7TNvu/q+Gd5uLaBwWf+HaBROnirboGZuWaIcy
pbSCH+PO8D6swuOP3dN28KrZjTmnSPNcPgUsS7mVcEZRubX+xsFVdBdOUpXooO3RH6DaomU7Lp8v
zSVxVmpP/zBYz7++oN0F5LWbXcsD/MX4FEtwv02ZjrlSzGgIaGX0eu7VQJ+A2/wGmtnnn9BCeWCP
n7n4f42+3/GFqrhwn9alNQlaMMe9x8uyq43pdu7S6UE8W3Bq0RMZrT04i7LnCEQvdneIxHR/z6dc
/CF9ll2DJVyFvV/c+of/P+1DvtdWSvWlg3JLhO46ezeGmffy0HKqb0r6Q3JCyGZ3qzoG3kxkgZnJ
4cHD/cEX4U2rPv2TACZNHgCoTDyvOV56pZpZLWqYLNM3Rr4hljDhIBKsV/rIJnQaTopilIKCmO3B
IGAYw/kUM5LrVLN5Lpqtf9gLwju1+myNowGPWSUGkY9yqcboT2t789yP/rwu4/huN0hncueouurP
sNUgEuVgp8y4FPxMNUPHdp0CnJvfYIO8eJ9mE8f7b8f5+JgOUI5+9WnftAtQL+gcDEjN6GiiROSa
vsJWeDvuhArFBacxdI1dxUSXTPKCdhHmVWDTK/H+uHdUW7SBkehUVxWUQVyNnDjpT/Te0S3/QaHR
N85ax0UIkC1ups7C3mcCTtU4iiihuZp026nx18C7y5ZWakHczjC8ytQR9EtKy7eVtjLLILK53rDj
ZQlNjj53yAM4X4GS8r2AMlry2Cp0Xfr83BARbqIbZkMuj13P9+WeuX5KgvLpjxL9MT25MTO36852
vPCaWbSQ9fJ81woEobb9iNFxWakD0SNfA8qXrjNweu6uTk1INyB6r8vUTo3JU+ClUIf6zPtazYfC
L7bGdkBKRMCnQ3ewEbjsyusOddT37U0nw0p/TqOeGH5U+++GY1SL92aty2ck3oguHCHb1sgDTnGf
2L7Z5RZ7W/bIeJqty1xpm6epS5Afy6pL7q7kv+K2AKTCol4HmtxMFyaFUoL2YtFT0WQlVw4LkYQQ
Wk00zkX8KT5tigDOk44Bc8toB+FVMxkQTjyKekokrpRVbEA3paABmswFwN+kgeb050OdSZ6rFFwJ
UtSBlZLG402A1fVuYy9vwzqPzWNfiPfto2LwF5A7/Xg7+IvfRahXANuYGvGc7UueCOuGlCfGgwT7
WC6SySmKLXWW0fAxuDLYSqI18ql4z6OUbjtIIp8xb0OTIVLp2IVqJJ4JEygwEdwIneamxUu8UuQv
FPz0TxDCNZvffNo3++gYhrp2V2alAH28hvZ1Sbre/IpcZ+Id69ffcwIVH/wVgsEK/l9WL6364BBo
KEDwkeBvBbtVuir831QfoNayNxhgfeJ37TXqPM0IunRIjwYCXlFDh6P6OftQNiWwpZVD0pxpe5BT
uUrAxCflamjJkAyc3+CcviDa717+6z2dgLbTzslZBJHLEsjg/YtmJteH56QGCRzo9wTJEhsuM0j+
lToVIvX6BPTA4t5a/82iS/WJvEdWSGvXSHm/jcOGgXXp5s3g3/tqzk/DY/WW6ODX91zL5fsVOjLl
WM31asJjDJ4sBfL3k4ltBoXwuMAUiHCUeGmcr9drD7d8gygIckknEwLWGOJjQifpQzJypAKovYBc
ypNKS2eXYCjY6Bzio4yJOM73HUfmTA0b1JXInN5x6A8Gq06/+I/d4DNjrqVf3nN1Egyi0+hYpZDu
dbmjD8VQKtt3F94cOWcgbc94kGN4ZNCQaFYSI8JbZ/Q46tgGCglsbbSunpwr5Ty/wciMdO+7dZJY
O/enGLCJFUj7FV/9C1l14N2bwGOVh3hP3oiMdJdiWdn4LUYccLk7AcqyFMqsJHPmE1ZkdEY/u3ka
c+nq+sXA9nZRBUqt+VGQJIGmOAeEk+eJ9WYPOfki9zylp2jrhMA9jW1M3K9Q6dUZidFpBksF/JKL
ilFGBQAu1z8vbgYsXbK9Wil9je7JLUGO928LN+08LOJA2VBxUSoqLABV9jc7j68e0JV8zOReLPys
jWP67wWYMKOmmiURU7GLNOvYftLiJ4Ez0q5auD6f4HnWoxtARjqhsC2/uKY8qHWK+NWbVtn1cPXz
eSDpjAwOvjA3U9AqFWbrc2VHsmdbXj4OVKvpxBIJfe6sY8LIYiIr9NYiiyq3OOHo524ddrvxQyLp
mD0Z8NoakJxxUrvbmJ0hFz3jk4q46fPM8mSqlkQM2CZM4O8h8QIAC6NKPTqaKCgckn+I6kXib7sf
BxpWeyzRXDu17w7Hj1oL6tR6MeydSGZTV26zsXps0fm+4kzoslvkeujbG4tTyoATmZdAITKwpuSE
HSb7FaiUA/45jbqM7xt8EDlnmMmxoG+mMIJAnO5jsw2r+lc+Qf6ugtLUZhnyot8+lDOKFWTXfbQ9
WBhZlCMsDk1RIky9y39nrRHc/LosRxWZxwxNetb09mnzHZlm5Mxlin0d7K683TTf4a1tPOLMJ/tw
BfoHfriS27sA2eqn4dkUyJCr+TTI6kXBvFuXIzMvVnla3HCf1MFjCizF55BIKHeY0W3G2k00QUwS
ksUm07UFICO3Ow4Vdy/EFyFuCNt0zrZqXZsAs08amcAVO8NcNIsie2o96pjWWTRN15Bcj5BmI0NK
eCJqByWQGaiA7xP8+Z5zk6j2GRx7LusgLcy+Pb4IPxOsxyGFHouDWdnpVYf6nydHbMYzixOyo0Z8
AJNDOjKrcdBtMqZ1Hgc1gXJCw9MbarLQ5M4MVUKx8C+9byS0J/F3Fo3UuvMetjY6QHNJmGJx2SDK
FZXAg5kfzDVMHmtxtDrgCb1+OPyxA9tikmbHEGz6FQ2P2zYrPross+banLRx2TJj3ipf0/A5oFDW
2Uheyxvz0r7FvA4nI+gW11qj+fY56UIVarCQTyj7aSzggevdcQUCYTG5HJV/Q8EJ4gatFar6BeNl
ujqVDVsWkmTf8HIV1ZteLyMGQ5kNfhe8dWf7+6gDPC8X3kZ84egUawyXtR6ANs4ddl0x/DBclagm
eoYPChSYm9PmzYFM1pzglZh23LvqkWr1IOeA2B1fPcxfdvyAvqD9ASSJGkFnMSwBIqcqU6PjFzqp
A6XgDvq3PmgargCkG0ExNLdPVhdh25MyCrt0rf4bkVPgdSdWrgNupduQvgJTIyYC9bxWydhfFvIS
h6oRqinRySQqnCNpUorgVg0FkSmzJyokYSBdnLJoN4Cdb5Y4sxG5eor77+Qvqm1IXof7JRpBE2f7
uVUJ3uEpQu34kZRrpQb1vlx3TMIZDqM11GoR86r0IKcz4QD62KWJPNMLTvYhP+ION0+957GCcA8N
fs29N/6CnO/znfRS8j5pGo7YdGAB6M2z1AfjYlhXQV/Oi3ltqaGB12XLjnSFmRrxiH1BTWs4KtXy
c7qPP89pKIvj/EDf2HJA8rq13H8TW0cFxbS0tB1ltWt9rMOo1YYOs/iwHVb7OTXO69ChEygj8AIG
r+a4+fq7bgUAbbOmwRr3+djzlnMuZsh2YZeWGc1sGADUAy6IOiKHE4NTwoOVegdaQAnc34d53HGR
myN3arBziWtRoHhytsrgl2ekF3WH3YwOH7xYnrU8e6U+5VOCcFr/xqxKtDQe9umJwWJX72NlIyrr
SKSFNU86C72oyXhjALOQ6Ui7nBWXJ5N9biMVg/xAUTn/8za0KJt84Nt9+nY4vFAhinCKIu4BF88J
dxPynJio6BjYbGi0SP+VKghJglYzqxWbEgGBbU8N7teJvMiRCxY1tOb7rrL65LfqPvleH6tj52uM
s96n/HhTmWw82tapLq4MV/TrE+azwQhQFzZkEIWy6ZBy/INBPo/yTHThcW7ocvXbjMrJE4/QsF9c
6hjOQXdnwHQ5kxbPYoeTlrsH8Mx+oqLYTjMftybS6HxxR0Yn29ikTF0JfUPC8sByDfYWBbOS/brX
pr57W2BKjtWYss5bHq+zKJMFrBBh4C0JErRjE+JWrYngfe25RJmjaeD2SESzi2FJd4mZ4gG9YvK1
BoFZYnqkc0f0/ZVzf1hup0AIOKaCC2JGGH+9t3087Db33ck9uitRvcQuDiT2usXxI0XcC2ACbRfT
9NEacy700kLfma+w5DeCeeoj17LIN62u4ohbThQYhBWvhQK9oHZVN1+5h9QvWyBzW9O5C27yV5iN
Rmqub6oXO0jovEixZIYMR1zvyqj8ab4Fu+3rg0PeqQS2JQbAH5DDm5Plc5eN2UFYiuZ5E3rACJwd
EJoBDvhcEmKORVOHwsZ81gKyaG7MG4SxEkaUoWPyzcUFH1IctENNh7C/A9KQwMgijm2ovCnvlHp0
snql9Gm/JshdWeWWykp3Pn2usIV2XzW63VetNuKe5xeB4N0BkH3gMkfuRhSOwy08IfdcZaqQjbKD
P3Cxv4tsKMHCtBfiN52ZuLBpuIVfBlbewB1v4irAWgvWHi5KUbR3izwIEdtmzE3XSsnD8r/kP3LA
HeU9IphAIdNGUqFvhD1hzvA+WPlMTrSWpB/0pqhfmFVQPOZg3NBBxvYgxWEEHNDbxdQbM+zsDuoI
tZ5owxofHTt9qMZq54i3poaf+ISOJGmb0fcOtdJdVl1UWVDWiKqhRjPdA6qU0jfZM5VGmhBSDzxa
pz4AsdEUlIur7FU6U8XxCw1nFAGbiW9tEkxnuDFHhHHOoQ3s3JoPFBaZ1PHAASh+Hk+JMP4kSfS7
A60N9mQK5fBDKmkNIPYfN86H5gCuw68cAF2Au98MTwb2xiTaNbvCtzFuoPbNJszi85WeRPu1f8N5
XUu4IQmbpR+yPO3SZhLngAaJqS9P52YSvkgc5F+Y6nNdcMZoT1IX7GIH5Bh6M0Pe30kTFX196eug
AiZon7w74ueziUp3d5IKcc9oSf6B6J/qIcv5+K9+9O55o1KLNleI3f5qEdtlFtW5N0Mdk9i9wU5l
1m+uxOvFKPjBLQGxX/WuEQv+7VGe663t8RBUP3d+GraBn05Yt6qmYtulo3R9PjHK/YSUSPm7fdpq
dUI4+jpaBpgR2k5kk1M4DsCM99BaIQdpbQIjT1bQo0CGZ4s1f9n53svvVzJ03sKjt3UdXMk1Of6+
IVock2MYxzH056Y1gHoH/cJUSt2nK0wUjt8Ah3r1RiaDIijRFR/i57CZ/WFoOKKbX+vULVU912fU
8AUZJdZ/S655Sc89jnjRuGe9ZtIUuT/AJ8Ue7ecJ200xXRHfOo3NDN4r/5h6mklcl40VLveE449p
WbQKJlllLZ3JU0o27FGAEChnlKC/xVXtGqUDcGjvWFX7vf2tYKN92j0vQDkM+ZCRVzJr3DIJa7yF
xk/F/TV3xY+5fHhI+9Y7dT+SixF5T4tpcI9e5417wHHp2HDkHyCVcy0r6iIDDZCvUcmQYwftwkn4
oU3rlS7SdWM5kic/XureFxPltUaNF+ZUTG6vCD2ng/2yF9WsJBggG/u6B9Dmj9YVA6ptGRilf2lS
ErVj33l/+NiQWkXBbLVjeejFU9U0iumueWIxfQ6gX/iVgqiwSuK6kWYYgEi/TaQfvxE4YaNUqZ1L
8MLGiEyg9g5/hzscWqtLFPWlMH4cdysZtOnIQUiS7yEOxXMBHgCEXM1vWKAg9eWFQUGYyCqMBuzh
DsTfZzhUgJ8G+dhrKQVtiVdWpPrWWdv+A0VBSKfopVs62zORtR1chJ9zTlRCkR+onx4j4Va5Icwl
jNUo+FU3E6jHX9g2r2/gfvuBUK/xGWa91zvD0hpOD7gjVTHz4do5tZt5UgZ05PUKuYYkmZ3dSSQ1
pJwb9okxiJIAXHhcthZu54KWRv7G3jpe+qtWjaTiKB+XQdbX9ZG8rzAn4bmD+jTVAeml0xGzCw3O
g1woMrf0lx7IZsOv0IEcXGZ1iYVmdQTrzYxWGzJqpypT1Bafpy4up8y4sPRLFg+DylxCkfzlXVtw
nc8L9hMTXtAJ73h573LxZ6x73I4R4H4f82w694T33Q1McpynqB5O1HzgdOFqeZd/u5YY58it3oEy
BLBgwEbY350tgdily+ItuKduMlMYCT+DeA5yJwIegIsqeNNFoPiR60Djknj0OYLMBO1Chie+ikiq
2yCHOOB85+V0Faor2eMBfDZ2igeN3XAy6bpd40Pirh83UuC4XCgXcIEM9lExi8wSEPKTkvH5PDFJ
ouHBKIkdTS0o5ydC1beedNhtR90ALrMSjW7Lgzsjxxf114UT2OOt5bzDczwMnuYMfNqzntQ9B5mb
cBOnYrxJncBwusuNObJwTHx8TNhMabgb2rC4pBVJW7sGksWI2Z9eYNoypEXQng8bN/h1nLTXQeTd
xNy7XWFbHLRGGFgwhJ4AQgFpToqVTzqbt+yD6FXARzXiM2w4NEHbZhdlCT8MKBFmcV1T8sTFdGml
d8fa7GgPBKVF4oGc02XrLbeY/8ddpzzDta611sMede8US3X7FkS/JYfyS16XVJOMfwmGIZ0zAy/Z
zU3/zWqe4gD7AvNxHtoRohdCExmcU7M07c/oIXehbSQSI3NnTDYy2CFfuF9AMmzvWXLSbG8yy8jz
S32f1Tidy1FykzB+SrHvGZphrY04F67OuuJzOn9DageIwhpzJ8e8z6MDCvqhmHOhSfZy7T49hzvS
eYleFjx6ut6fQ8qYL8p/kYWxdEasE+Qy71EJshW4GLWJZ1G9JkfBFnRU+s0sJNGdeiWsK1DkMeuZ
68Tum4Ob3FoHdfedMvlu1JipEWybgFwSvjas4BKB5aG0F8AkcP/EHcOLShs873kXhfs8xWjqDElw
2xsjvdcNhL2R1X84jSBdR1Ia4UD5VvvjdFGX7XbC1w6AS/d+r92ri+a/vDGAc782qgWryNFjWmxr
qV4rGU4kC1EYUG+xxt5DqQt6KHY50mLoo0jjacvFg0ZOVMgqJZ+MX+8BMNwvOY/VI1M1a6z5AR4n
IHkNvh83SW9h4yHkPq5VLSJDzTeNY8de2YHWXDxk+8k/YsKR80XReRHGqeY3RFvfuAu6J5rXvh1u
sGtypNOobRLmau3T4sfQQj/pVqbnpIk24xT2c33LrS+XGevP0DchKF3lGhEWqLBFJtxrl5He5c3O
8SiTNY1IWlmjFsfinnnYgem5FPU0EPWXvb3qF9YzcMG7QGccv6V44gS3Zw1FfBfpWg+srWYncmXL
/9RAVGdsWRqQmz06mWzjUQ3M/Ck3qk1yQLkFMVl6Vxm8VJlhjMDWv3DhWqWB4LU4I2OCK7zVp9of
nR4zMbeidFgGA1E/eYZaecR+FsB/B5Hd5RsHg2yGAWkoXAugRDwnDin4O3bvvCNfTzNUHp/GPfnX
JFpZAfThXW1JNAU1nPPfyKDAUs22gZYCPfXfTR5zZiicYF1FSBgF2Ov7G6DfxfRPxURFN5KsoQC5
pv9rhCEwaa1T+GETDfuQL7wMyThb1sKBDP6f17JjkljVlG2CrB4RCr87seTetSeOyyqi/WGC2DMS
4Xx9fzAEjGGrFSmEYMwZFx+CWUjCvQChyJY09OFPFnVRX5jwUeZiz56xUvPBs72k/KDzjrDien+8
aq93x7D+s3WXuMdtYcXwAIaeatPRXnobK2tE7Rk/6X6cPLCvTFFkxjOwGCZQpHG+czPTXT+AM6eo
1GHFzrVScMyeh9Fr/h8l1PTfm0LOtnI+fWHV4kIGZ3hpqHv11TfmXqu/j2FRhaHt4PEzb8tK7fLY
/H1/XTYY0E8HwQ6yU5Pup/EPuPdOeGRkHtXcai85EFj710P8pvnLyKOBlS+E6r1AYZ24FU0YgE1k
E7UOMsvRtv/JU6SrZQ96I8KW//Dofqei25D3htmUw4s5qzNdihemCiYj7IbCElE7xZhFQYt4DS/K
xAyb2xf2XBuz38piaIAvAlAECZsdJCUYX6CiTBop1jLVZKBR+kEKWFMJ8ZdfiJOn4wNeeNqWEdcp
5+qpt0HQzrfk4KZCR15gYPRqQRI6Qgcrii+QDeLzcbRKPSIsbH+N4jSvmM91rgHt+WfLGdUfKtU9
VMZehfMDHtY3Bkcl3xIECnJgzlofRHczaCF1ecgavoFRTY7eS3n6YEfwO+qNSCxIhie1T6XxYZ2z
ZP7TCUnrWz5CrRnKaBD5bYrBrm+Ev9Xla3g2sN/2vwAkqrwKiXc9m9JqoTLuu4LhsqZSco3YMlvR
GLEuTXvgWmLZrKXX6ZtKFV2pVm+PS+IWCM81XEVdLdrZ4LI0a2DhnGJXbWGy2setV6K769QUVbgu
LyinXBS8yTdONwUXt9dbBtePwIdIf9srC1rrAVexTqmHbV2sXgDKAnMTqVLs2+/EhY4zWVJtnX2v
NMHiMVTQQpGZ4ZLnnLd5Dueq2/1AdcGjcJHix0NVxffh45azE4jF5PvmB/f8AXpAtafayCZrNfkm
r6uQt+MqfimTHmd+PUtIu19FuY6pdBNs+5DkfB30giojZBo1uMRjocD5J/9L5NRPMbEkAtL9DvRI
A64Zb0f2UyqrTb5izICrXUf42Rf7XvqKxQ8KMwPZF013zx6iZn+E2Nn/5AaSw+usArehxUcrdbnw
3GWAPKwFDmalGDf64qCSFnf7EOCFr78N3kUcNKX5h9uxl9XBhgK5iC41Hkwlj0hBbQtfj8egzT61
qh7eaMoF1VhkRXoRtEbXF5ElGOYhAQ1q4nB8BOlp4Fh+AntXQeBQWhcOHps/4joUGqxrrLYohJNP
fbu1GFF7AXdj01KloLvZ53jldq64WThdvts0xphqjmDy9sAcwbBZOGJ0krNmfcDp2aBTnmxloKeQ
Eegs2KG1tptkPheu8VL9DfTKg1UFqHLn3jpTIhpcXCdatuUdCmBkTKRGtdteohDdJIIEjkrD26LO
bCjBWM6VJ4KD4IYbBzbqyyv1wn5wVGMvv9cuEDAb6kL09bm4uMZ3SYATX1OqRPDUcYt94Wp7AO1S
T8EcF46d7mnRCa8z6TJVMeuKp74AgWou2XoN4WqWudWa+XyJslOxUy1NIaTm7YUl8GpunYLy7s2v
oB5spOmkOyubwG2nWa1TV0IWgpDsgGbh1P3IPZh+g3HQPBVHHiSxvKPUFt1ECIJARqHaMcy3FsBN
UP6Lp7vamp1uLOYde+kuTIMxZB5rMu1JpDiFqfzxO0o8gBZHnqeoOQV4CCTKaL0bRBL55cGfUJQn
GnZb+uUp/h3Hb7802FNJwThcRXcXjD7Me6Npidzc4sDPE/7SOa5S4M/Kzia/erbuwBVoayZm/cdT
c5xW/LOv960A73saOysoRX9Ko9vPj9+9f/9lSQICwTNIoXPWBRgB9KW06oQJTSTe797973psmO5B
hVhlHj8KN5WzK6E/GD7mvJuvsbnFvFzY4QEah811XGRK8s3huY/G+mcNHtdMOYIV6Lun6Qs58HGC
tpSrVUBKOCia0ao63bJMuIUv3SnMd5sSoAE8uSkO0Gltgt9QpDTMou14/ajYnsg1BQ5N0nzCLiW1
24Gqvinnzu0PZ0JJu60dfEeRv7THTBp2a4ztyDDl3qtO2rYjb1EDwqQ85vTBmnSo2VTJ3QBlYWpu
nNQTMhmdf6RY/8CeBqtuUmo4SjlaZ1glv2vBPgI0QQh9g/ZfbQ/t0G7Ki1F8YKissTkVOkwjUbim
XQ8437y2MLR25wtvMIZuBu6At0Fa7KyEyauBWGCZO6wtSJZ2PuUG/aGoHccU9s8up3nYKcvzQfx/
upYdib4bVi/k9SR6H8r0+GGqedy5c1s8eyytRnCuF6DaFqJRr3sOdJ5TAOHDKrlo3CXuGTIXxKrz
Xy6y613v2jpMo6LfSGrt0GwM7CtLgvCaHM785GJkGhLwO8MNVE0lVCEE65F62FxiZ3XB0LuLsE4z
SwTwdr1S52p0TDr3LGTj2cfyMrYGImgUuTCTEnCoy8UPZJjhZOMP7DcnBt17pxIYkXUo5HGthuJD
ZTjLf+S7adN6CFzmqC2pT6B93cWMJvdOTyg78Wpt7pxa7KoNaStIVIO9bY0NHVcwXgWQyp+M4Swd
m7xVTlwgGxBYNp/kaKPPGdh9bZI3Z4TwajLwmmTvT1Wc4vFuCs4DMB06GdKU2k9BkaxONoXUFePc
uRwAselr7btcQdgiQkCNoWtF9lywaLocMEEC+jXKnOoJk18B/H0Q3chvaz3fBSoBQDC68Y/kEsDj
1daW1QQuJgLdc3ZbwJUviY43wzJxOTX5ludGqc35baoMutIFdRtsnvLo2ijRrHfbWwAKicaeFBuQ
qGHK3e36FrBLiQAw4NaZOcqGuTo0sAUvZXjs432qUHWHrVOaSbBMvYcs3PVnc2O2JvUvNhGeIfWY
XJKZLjTAAqOT8JPjJPDjS73KXJ5MCBRtuY4Bdj2loY08AVwz1UnA2Z623/rWpi67OFBQ0GizBXSe
Z02B8d9TeFmnF2QDdwLPyVYLOzFybwuqdQcbPSn9SpzqPzGrM86PuVMSkYrJxv+Cj0PdYiB0PjFi
Zz4ossTkeqs1HBPHQsadw5vJVRYY6LJ1BnZ09L2vz7KTp3t3sM6yi/v45GQ6M0l/7AMzOypXSgzc
oXTRV6pkKZwPO0GDi51ULk+2HmMzhsnopdc1A9iTrpBuai3WKNuGuDtZcaPA0H8gciiU9DF8C1tL
fHDSQZu0zZpnezBydyF/AgWeuNtJ8U6qoVbNYpaBASvnW1wBqKu57mW/LPMYRyCVus7xXB4pJfu6
5fxGDhrIMVC2IC4LGgCWyczE0VOWUczCR377f/H1T8sThEXZUitlBR5KoaD0rQZT9GfK9PGVlmDf
E2fQuEuny/a2kVD/4v9LY1iEHxb4vLFXwaYgI4a/MGbEF/i8c42VcGE2Ix+MiyL2zACdZ4chdwIt
Ov5iuN7H73yoEW0pE5X2dApq5b2KUotK8jXs3s5B3RNPZrYDVyqE1zaQUXH8pFDk1i9cWkTJ/NbG
ah/57NJqDjJDAD9LAleTGk6Eso4sulIIdg1u94LU0LsL+9BDx7ueLq93lhWJN8wYSW3oqamLebug
VkruJa13v5d1CxqlITnulG6xnbDAGzl2qzq9uPf1X1nSWXyE0mzL+LDBI8DhOS9eGHT/jC6T/Jg1
Pikymp8KvXO54xkzRdssWSTs+k4g6hgQxBKqxoPHSTgi725dnvyhpO57IBoaQLKDuHrvbvXgYSLI
X9WtX0+WVev7e8YfkxN9cCCFsz6k+AVOX8wZhlLHBf9m7LWgmvmJgJ3DLScUkQ0v27KGyxN8BBw5
S2XxH90Zye5L2B/Ki6CKo0KQZ4KsMYaQszHw5LeKTGv6pnP6fYM3/Qo3eUCC0tCH/9Xgw6sajzYy
1ZyejpkuDXVGCLBnt2VchinemablsIVF/tlTig7pWdB9//uC4uaPXpHi/itkdYQ2q7TfinOVf/yA
2mXDdGAb6Fx8zpMZ3K1ic4W+b66iVVm/5sItLiqonapazKz6fo94mprBiYTMLbyUAc4PBaK2Spyg
bXz50euZOGcF248SiybSD46/1jLONM+H543XM/WYodBA5KP/5ES08aDyayrJSheO0qjr4R9YqPw/
OQGpe7Re8Gpn0QzUyOT3mqJvLuzKCeW8BDUhyqc6VUtWcUCKivthzXwnyw13jKL8NW3ylgnnzyJK
BHRHNN058nSeYsqh1jxHDSXaYGjKhI7r4eVCPjE+JsQGa4zAaN7ziJZuCarLeb+9PLJUjusmCruC
lJuq22H/F+ULeLNQ2xKjRiR7pvKOPMpmt0j0HNPIvbWQe4V/cnRYQzRkT5W3mECV8IetJ71jv3t/
aC2FD/DRKRZgMxLUe5JlHowiM1E0KmaEPT1P9bMj481V051QxrRUX0KPHzlMjyPTAl3aOVuUcB3n
mq0X1ABnc/QBnKMTmBN2v8b6zB2MHofEd9F5U5SZ8DMgdoWEU3P+7akcR3dsgfyIpGKX8Gp078DA
cFTtQk2DchzcybVgsORJ9BijbzaidtlpaHB9e+actcA0vlgbyZ6CvGn5hu9bJwKlxGq9QxmkTb0J
AGtOReO2XcsHqX7CW8p3Ll5PcZVRC7DlZ8lAmeWSeLIg+Ti+P5YZIzOYB9vXziVTKb3w5NsxyxmK
abtes4uQAXSkNuM9oADzr7P6Uq7fGfJTDPD1b03NOafVe449BvtWRivM8wJXeKlCoZWvol9GgtLR
/O+PcrEpe2QdQ0tNM0h4v/jmRrjn0v8NGTFmbKiV38oXXieksyCIo6PZ3s+5OaTCQ3agDmy8ZAKO
TiP/FWR4SFs+fhIHaZDAQgRh9V6Xokiz5nXdPKtSi8JVOM9HoAnmWKIINGakwvehpaWNkNnQaE9f
Zc9UbGj67rtNWLhL7yUEzicIvg9uB2VfMOgz66P8stP6UtnT1AO8MLSSoI+7pqIG9n572vx5EHj/
Y5BsTr1OfFwCV3UwJ2DkrapQxaPKTo4n/erie+HIJqxdTwkMmpT6QHmNgxbP7eWHZze8V70GIeZV
jX7JjJP7NFkcf+52/yKmjFMhsaSGJ0pVghyyZ839EKlTdKRFmnywKAyIpNWx+ecp8oko3wfgg9yE
XuqE+IAlGLxJ0JmXvB7ntc2i0CWyFv5ctioEK+Ti3UrB9+IwG1RsnHMN1PABAvYZxtODV4DW3+nF
E0evpb+GyLOdhm+mNYsTn0SPZKZvvijkou71VMmVX8+GkhQ81jPjhLFOjIyIuZjjryMEyvQ51v80
+G1RSz9cKLmqAzKyjKEZeT60q5J1qgUBAtE6316xQhXRChRAUaN3op2d515nxmLNyy7zsZungGI+
yhiYxZBg/Aq/B0UnLNiIs/h6t5+jI0H8zbHfTiNoKknCJ5KzRYm4Br4Lp2VcurUVleqi6yw7cxXx
chGOCyYJ0yLZRBVYM4NrDdTdWAag3oFWLYgiFPttMF3q9wkwvPQ/xJpNxBBO+O5toKz/f0Gqh3bQ
r82gkS/QePT/IAqVWUtYjhPT5w+2XuR9oBSNEDC166vhOufT+WKqs28C4GF1mczFaaeNpvKtfEhC
gg6qPp52jR6JTSpN5110gvjfT2WXaGq3H9Qj5julV/wRO+lmSljrAYI0xf9pMZIRPSv5beF3V9aD
rjrqlXZdn0v8rqrEsDEfDoTrDYnj5PnzEqjC40MhfHgFrQ5ArGgYKJmTZiVGa/1VAD+ENTz/V9pf
87X2OivpUOZ7b3kEauEwINSlOHvOTaKyK5+vAJbd5JJTFE961QEbloAO/crdcjd8ZG97nLfOxuT1
TQTbql2MCCpJAzmV6PyTRG2UEEKb5iZxh0b9rKLaxev/0/64HritTwO7T8Hq1XUPl2+eiQveERlE
oxq59yr2mHRQyh5IAHkaFbfVvXzcYhaYInMbydEMUCUA4opPELw4ya+4xVbVo7OhqbwyOwcpFfiZ
rsBd++7llEcDXjVXOgkfLAeE2pke4Y58o5DL3VnlSxTNP4MMexsUfdUgKxsm2yzUIto5pc+KUwtA
ZyCtDJ+CEAb1Jx9KfJsJs8CnfY8vH3/YB8RRADl8P9K40TW4zCCRvW9/5bPKLgZCKZT3VSmdHP8J
49I5iE/d9xcJIecB9POoGirc9MFSYbd3QfvI9MbRLV4PDedmQ+FT+CgUYUqzs2ne5Dna1KZghbUb
gRxU71WaVl4SgIcEDLIPTaJhEe1+alzVaBm/98/hoP8TSWqJlfpEOAdspZdfsrZx1oKais75rAsE
Wimm+5limJwhE3KPQ1a4ZIUu1YO6VrE8U7Tv6A2yVdLQc8JYuPaBm9f6/8871wxqPWdnP7WsxUbE
h5bLP+eQ43I6fJbnHxm7ZTn5G2cKmvc+3oMSS0vY490Bp7R2HsjRXi12r1Vdqp7zzGpZnE3BP09J
fteWVHyDXECoSqu05rQ/cUhgeklbwvAhgTSgEWwm25+YrQ0CAsOfHnKVZQEPqTQq5Zxoy0DbAABX
hbT2joGuf4pO5ThOg2JCpfRGOorveb54VLcFtwrYIgasUP4AmjgJ1wfqGDyqBZC7dlHn0xDL+n5P
G5dk+LxytvKRVe6rytefjovFo9R0xeUjtVWflEkW+zEcM440yhYBTs1qWfnUci5kSXBDhCKtjBeI
Dq5jtdoKXeWtRjWOODZkD2cBWGLFgTeVlFo5igLQBLCfk1vXpSFTFLu5OaDk26o5En16qbBmo1uI
1+ayC3moOtG5iaa2Z5eTw5FwXuYrCecWCJQO3ptNMNrUo69bg2PSIv+jyMsBSLFwcyLEDwkrQgT5
CuVLARf7M0gIXLQ/4nNHFC988P5NrPbRsvAr5HL4zOtqDYkjpUekZYeGGOHlV6SfbuXu3uEQLFBf
TwsAvbPmwh4QniDzE64H6AyHz7SvNxGSykoPUGgxHDHBgZljI/1Z8LdMboia0DOctpyLxRjR/hTH
+eMKxudVldAhSFNSxItofKx8oiztnfOWBmKvXXirNbrj5PPqtQNyEtbhklQ/IG7lnyt6wWNxGgkm
IgD2/7HRcg0HNp788spe57R+m8YcZJ9uWG+d2uE7ylQ+LlDbu++V+ui7YKiM0wtCVldXS5tI0i7T
xe/KDSuCyIAFn8zZ2KjAecPx514d9YZyQUY6nPXKyr7MmcTwtR5Y0CduE0xnSXjFwoO5TIaUNiTY
w5q32MNdjGCsWPJKhqsqEylxU6ljyxrC0ZZAgavXHdwZC5pFiUMQ/iXKSILV4Ui7HOEaHBd07bJu
TUmw42gfNgBUYnLv30gdFi9pZaCVSfLTHMQjLD3pukEPP3aWaOIxTOzAxrWu5VfFMyWsvG+b+8SO
A562wGeHAsb5SilFHl+iM9hrExjxkIIXqABuu8Iq4zB0CUtTof97+JRsavaTYJrRlHrVVanbBhU5
Pr0NlDriaS3+oCiF+jOiK5fQHsJTGd4ooTYW93PcwncFNygXC6XSWlIBWy+vailB+5IA2JrSBQbN
lrtILkzhf4DYCi3pm9CQH4NChw8+Gn1KrZmSuAyXJJcMN96ILYcKDK2nwhdm0maJ4QmvmDoEEZlw
V6scvrzbbrcCM2oBt58pPdrdbbWa/0UGionT6UDpZTOKOQdDQti3vjVSRORzL8MNth2T1DN3KiG4
uVpgIiteyDdKMr38S3uscj94hFafxRSroMcnOGlhSqtjtGiZH2wtsnjhhVUzZDo7i6Df7bUoqsRT
0XoGS0OtT4b3QIKpM+ZgQNlPYy5Qmi+XefjF1mRl3Uy3REf5gMdibipcmWVFpa/O9YZcV+XhAZJ3
g7oxOD3jYuRX3ztDzx6fPYF9a16PgDaIZCyyuDVpJNjMirmV7dXYg2EgiJ7UyUd7K9VZW7ALg4wG
HitGH6ro9Zab9+K+bhdGFMme3g9dEXG5wZnAxysJqEbtVzKAUGEyUpoEAmz8jFGLfBMZV2xyRYcD
ydHTKEz2rtdI0QiSY6g4smMo6x3p7MnGt7dPz2wzFoV5Timf3kF1RCtGZJjqdbtWbAOp7y/lB1U8
25piFUP23FV8C3cVS9xn/5f4+DXT0qXLgCfMIGmrvCOCYnsUhS8bAYGIChd0X5kTxspwdwqe/D+N
UQ9X7y5jfIeQMPP6K2anmICys83PwMBbSywzML7B2ln5RGw2eGIXVVGokFEn6S/5onR4avU+WGT7
g+06Zm9rvLUOB/TmOyCQmEYRt/82SZdvPgqkIHf4tmP09kxZvm//5U1HXLMTppVSFonRyd+XIhmH
f/S8SxPhFbGQ/kX+vRJsfnPZMehesVWPVPRor8UxJjH3e7OZS+EeAlcgejA7MawqocwL1KiRbkpE
Hrf2wLoEYJWYCmP5OxijtfAszdM4H32vIv81fAun8GifpU1kITtDZ1u8HqF6RJEOv11PEf75Sq2g
BZgSNO7kO08WOGCZLTwCCxgm03bK6fZl2LialN4sJQPEo+DQM9a35cl9LenvVhkpYifCthfTD+T9
VfbQk0W/Wefr27cJRvZ1NIXnckPBgk1HRW2keAK1tCrMld/YYjQhR+KlEVokURHmOoO9SSxfsFsV
ZifUvR5G/chTIedmWu5+ACTHbW8pnMGf6/ozTUFcSoHqrG1MBAAWtOlKsRlt46Z2fTtQlhZBM9bf
0hAJ7WoLQ4LG4iiKKVWTiViGY7Uy15TEDP1MkcTXO/dWRjkyc4Emj+wWotCZHEMNOwJFPVuUFotK
vv7kV56tRGTJh9PkHj21Xu0LWDXSCCoRWOX9VGSndwnvbrII/l+fHMZIYctIMw5rRx6cFx3rwGAf
Y9W4JRFsajG7X8utSpFs2gojOuKlYzipdTfwIrER3L6ssK/5pj8f6MvhhtOwh0gqfVHAyuX2GSz/
iTQQJrdpk+Uea9cefqtcyYiuMIdRxDu416XCk1LHzdKvW7dLHN7HMG01q3qeYW36iowYo5T8N/Dy
LTRLur++3FJ8C1TrvHzPQzLSucvWeH7yOdKKr4aY7746hVQ6gI6z6CroW6xPhvin6chNdmlB/brP
ScP3yz5ronFXhQQjrPnzkE8fZPEGP22rEdL7OPyDroDlZdgVk7XXZQDKHgOeo+llSWMInJ0uoztK
W8PgZqmwczrpouIV3QbNvhyGMacLPCp1S14eaNrYf9/ne4hi9fWdRF7lXZNmoit2ZYBAi+YdCqwq
pa6SMqFoHCYA/j5vpzX026po6W88WyP4wjijpYB9AJfKSeLzAugexrueiVEUQF9w6MCG3u0xR7b2
vbFz0zYu65YTlB1g9JKx4MFgcJmf3PWsgfFB4a/vf38PqpNSmSJ40vJ+xa92+19DnTpPRkMQ2a4c
Q5zSbqazlwdmxhCZHIUqafpV2aQ3h4amTEKoFs6qWtWTtQzysXyuukWWgLVB5xXxAUP9wPoHd0KL
bSzHzBEyB3C9appkKtc5fG2Czk6dNjBs/26YJKpVU3HJMJ99IX3bvnj7FQCNT/vgG98UOPoTePI3
SETl+P5/sGVzTrFmtO3Tcsm9aG3jIDHcK/z+Gb6T3f1RIgZ3D8en+Ci/H4vXRZQJpzmPdlysgdDS
Tp1ZifhYZY1LQc3ovilV1yJ5vKxt61PekGhuizQqDpFCz548aQy56Dvh7P2iAqni4b4lBn7nUt3h
DKm+xzdhsxWu0y10ZCKuS14y9HKpV31OZJqZ2Ys+d/PKvwfZ2jG7ALCW1e56x2TURNcckBfZRBlq
sOHkH+FCVHX0EVmnZih1g6vLeSwcnZl5egs+4uariOQrcIqpQtborv5oSsl+S5A7L8RuiN07EvEr
wbW/N2UKfo7lXnuDMAGXMBIK3noflb8PbplcjrW2lvBDAoxJqJRecWL8VhHYCPjlN0OMKi4j/zfp
NAwaCIRVhz39I6drE0c4T4MmweDqypFNvuwW5n8ookDp4BTKuU8Xujuu1/o5oEQnKIMOse6xqras
iEpAtEf+6eYhju+v/9YzPIvsI/WARkgb7q7rIFKqlYB66bCFzz2q3vAAXbtgXzTq/5y8ixm++I4Z
mRoWJ9T7ccHLOjh0uXi/OVtEKRDBDl3TWCZkg+NwbnToms+extlTEVKPr/ud2yQ7MZohVeybLejB
LY+y8flFYbL/x/OF85FGnRrmQqn4rSi89p0O5mPCocC1bZ1SaQ/4QguI4e3uL0/7CJi6eeQ1fAH4
kEqr5B0EJTfjMsYB8NzHUJrGd+wTYTTpNfQSJoEAbki1KD6vsxEaz0sLAUB1Kfy2Wovd1bS7W6YC
IMwh/2cYlr30Y6EKoqhsVwdXw3scWk6CsxipuvVJ4dsumT7BMpSnlzxkx4tU075gpEue1zbwLlhY
AyQLgAP41JMwl02uCXmXgtglcuGzhz4a4AGafPn8t774TzQH7qiPfG+3/Jy9i+DJ9NFDSfB/CH8g
UsC1XvS569ICV3whWYEf9VB5qkPSjPHIGHmElQZyLkFXgf1qhznEW3wquihgeEZ6ZwkEXtzcHPVk
hgMwYASizH3I+vBdsKJ8/4CB044wErjMAXbFWr622xYFyDDL3jd4iE6lCRUUwkiIVGhgFTxc+9kU
8Bulbj7uIOLmyEIVMsNQK29Q7p15zzskCJg1En+GzjQho57hcDWXbMXpkLjYWczfg/egUfg9yc6O
WJWmj26kVwFB2J/SBAhXxiLu/CnAcjDvFVXo+Uoc5Ui6SZRp2+4LRQlBy3ed8AP3gSRzFqjQ9MjC
RxycgGOtB7fc9AHbO0MK59/7xn1F5NHbpmZRoRKjjp13RJje61Jt5N+rOXwptdp49zBV5WRJUmQF
RrOWY/9tV/M9GJ31fJxDl/rY6x8jxu9y6ZUwQTqwGO1dM2U8WN7ypK/Sr3U8FdVWhUMf5Zu3ZLSg
Iog5VV256xAfiUJ1KW6+qVb1tMSUgJ0oV2pTD/abrJfe6Qr/Zhk6+TD28e+zelrgpGgJ00cSsC0G
brjxeGXM/FLjW0fzleJvPSK6acD3NxwvJoloH5TZUoiXQjGXfYhn8agYqZSfXfrLE9F+Q2uByeTb
y8I9RgG8CmG112rNJk+2SaEH8rCgCNUh8GCIu6WQmJ3y7jIPkiBkFiCocMuk5OaTR6QGA7LeRToe
2NmNqHfebv8yR5UQYAQEZqI1KR36CtFqvx+beLOODAbTUVAGA+LsA1U181sSaeRPjvoFOYTgKdHM
fO0OPGQWH2IcwfIBLJ0s10bAPhTCb0tc1AnHzaUwTX/SrqFHPwsdCq5QsFWgmEtlXJpnSjOHOvDW
xCy0tiAW5jFfTPuBU9HaCEopKMQhVxsloVgDmgPYITAk68hDL4Kh7DR8Qh0fSW3dvkdFNTXIl1Ld
2his8YGLBFHItMsYARWUDv4f/EfTHAbG0B1WLVBJ/Wi2CilhnkQISHxcWpzeum6JRAWv99CQhJ63
J/WvsBS3Mr3+cfQcm2X8UFqHiJ7rM3vTcdBI52UWZBHF9CWZSGpLcpNwp4GrNhR38NPLWuhg+VUg
GgE5vFj9HpGRcaSctKnEWbgYnfx0hPSdxpP7maZFa5uXCDj2exITRhtz5x2bm5IQ0hddEJArbR1m
ecMX3SNUu9K1nIsK5Q+Yrbepafj5OPGszgDykNjiyh9437vhzTK3zGDEo7DPqxZyHXvsb8o5k9fx
CYFmFCJirNtYx6dt2l//Y+3VYz+cLmE5pW/V9pPIpyJuoMhF3w/f9Kj/jM9c3kMEByL8VqNwgkjN
ynrK/MrMl7aPOeKQSECSnOc5ByPWdexoEWGPZ6Yr9ooxV1F8kaVMcTYK5UImg8pjtI7atoGnsUqs
9/FNy9YWWwqYS+CeBsBo1kMnzpqEIzviwH78F/Ul9IsqdMBIlS/RBrgWQ3QFOSAnAukNaTCCdYBP
ScYzeohR5dF9gWjuhyp6Gc7xucfc6v/n8ixf8Rbdchtjiy3QuFd291ilnKPr2WgTPEjhdHygkVn+
J1Np8LpXHfs1xL4oAtJPfvawDmzyx1arFFjPDcj873U9U+S4vw/HrNLUiibXqW+ImCcCPugL5GnY
kZrHdmjhKXrRo/Wtc/mcBMTsoWSqkxl6QnPR9zmiVvO3q5YPkpSX0fjDZksnG05XGN9OfbisoXWS
NVJgK4mEWfbmqakzv7uKsRvm/cdb0qqHnMYpH4EECeTQTVYlwD9uXKTNATBq9iGLbytlOTCZeSV1
rYVjW5CnOTxsl8e09s+VfjHivuSJy+wtgDR58QHncR1XVgMFhDit+e/Kpk3JLyYNVl6iUB43PdhT
VTmwY9iRDGMt0sdlPZLpAuNbd9KqKW8acVW4hkxA2sJi00jpHn0E3o+NIFGUSmnQNEueluq4K0C/
RnbtqKC83URcE1vTU9wVuaVjJV8i4WXVhLmTH6jVZfXnJEYYa+cWysMrECYMFYs50HRbVhx9cuL9
qagWdHFbP5iuKRbvBLHICzomC6tuwaHVllpPYT2gkSGEHRwayl8TihB7LbINfLKR2yz1ZZotgP0e
L268UZ0aT0OiXVyV2ZDC3Xy15uTtL4H4pmybK4K2CzGUc1ecB9BanpMbYVdNMxJ2rXT1HtlojJKt
RhmqexsPoxpexPs9rMwkNwapmesnB1vJ1nJ1LkZd6yOQnwrRMNSeqrWQ+x8A1tn8LetLdV1bm5FR
LK/8l8HNNN4GC7l1opSO8423ewP3qGSL+qVua6cCgNae+LEtZ+OmMoL2uG6Fvqx55xYgEitI2x/b
JTiIe+wFza1e0784pNobFXvc7M/6w1OR6oYxZTpZ94VjSUJpvpbFh3T55Kpfq3AINIKtgb5P1r2S
i3r9VSM6KSnTc/pV9hXa05PKRoLbacvf8cYPeQWWLGIvAP0Lcl/DOkZN/+QVEVWuamGUnooUiXJ2
40LreU6d8RBjVmkZwp9VQk0l1QS/gZO9j4/fVobtJdhvcOEJvLyL3gm0pYHPZfTG4+yFo2IEAWIK
bQLTkn/e1J8Y7gAodjBxUcaXnUsVBWof5rn6s56r0reCM6XlWBqCWKx4tNmohve4NwC+my13pjAC
NHd8NYTVMKpwQavXFupUhWdFq/IW9gTg1YarLCZi/W2D1CZRHMwIiJ/y8h+yHbccj41yIBTJYbmw
n5jtUbNG+4TA71Ymy1hkMWk9U5o6laEHNmG+cnXhqBzefloMJygs1ywWHa7PM+eHhB1AfD862YgK
xssbAPBzw1WOyHX2xLjrjPlj4ATTh1LDHx0DEQmCtRR9lSq643bCSJp4vhARVFACgnx19+DnZXvG
ExMe7OO1DS1x/+rc5RnwyHDqki/OATqZsyGJPEz6IPZn8kYZvhwuBQdZtJmDJarEpgFIexo7bMK/
QLFQADbtK8jxiyRxJbbr2KM9WUpFcbS35FRAfRkUM5Vri5789/7poABmCIGlaFy+AAMALoR65zRk
N0cGInqg7gEFH0moND1n8ZO51zX3Y6gjYXozQgSAGxkhbqovPNiitfQ/KXc19Vxkzxc2FXEa3JBw
NTF2FUk7mTbOMJRRWorE9TbTRzMhFNiRJvvLPbBsVJIsCsq+Hrd7xRKvFdxO/V15phG7OUqA/eOy
N4S6b6KwXthTvL5IrpRacnSl7L/H305GccjaVU+5/PbX/NK0EmlHE9qKW3jgPt/Y+6aITN0RiB2G
1Wdux1DeyUEdLmOjaDscBSUaLvfiKbgthLTESmefz6ljquROX+SrzqKm4ZDUfrqpXXJbHEJ7kc+X
XnAxbG3C5r8PET+AoDeLKbjtH3bGYq/AgoYmVHXcS01YxisectQIFewlxr4LOb+I+JkZVmSJ9lZk
5JylYzW8lA7ZPwkpI2dUCBIZlwoKubJJpnC3PsFaJqnyejPfzkfNlwd6Cq4u94ViY3WpYRavc2vo
GMHzImGKKqzwyHa+sDKKG1Yr5Kc3DKKRTPXyfwIq2Ky5v6YL7z4QzFDXTeX4vXPsNfnhnNa0bi4T
XjG+wTXpu2DsQoQ34YCWePRoRyMT42zNrgk0/Eo28z46EzXxv2Y5YdtVGJ0sI+Ik8vAERYkDlZpm
qeD0jFLdThjvyr/21/jTRPFKu9ov5V52AeaBQELBusrLF6ZaVskSanuBBYMmm3ncrCwW3bZgyGEU
WOKeUf1e4/O85lNnvLBVFejPwFpXW2bpEd9BORE1Jrfh0WvrGtG3u8z42HLlo5TM6uO8b1fLIdOS
mFdlHcm2ZRQEN0HAZfZgWdmEQblRxLhYj+GnpSRy9E078ynOO2fLoMgLqESjm3jfW0cNtb2Am5xw
597OE5YLQcpexl7uRy7xH5Awviksiz16/Cm55MqRFfim28TU8mbgjDgWi4xjYT7vNL+HAn+FCZUG
QKzVhykC+H7wiaEPxNhatRMhnqKwgSBXy8xESIbTwsq9/HIL/f/rsUrWxgRwfEPqQk2wLgwzPmJx
JyFOuGKJ2OdyZk0YCz0DF+NzE3200vQMsg8+O+FhDEdAPtpIaOOlcEIFcK5QzOykQpwu+6tRKYjM
MtsYfL0JX/zZB4ujkaJQuOBU1GZ9ht4V025qGApE2lYq9W26ZocV5JMfpDl8I1oCemcuTg6w0UKv
3F+F+k17P+C1wIxky6hFW464ubHvHfWu4zJuQ6VjTK3o+kn06zjgzmJMedcWs5x8k/IcpgLBX7Wc
A7B1e5CAHKEagOJ8PETap3Vr6NvS0ktFOcMy7GSncw+YzRIvVZCBSMzQ/iYbtqYcfgCLMnw85p2Q
HbLRRMAhyP1/BjNab6juAUNOfIMYQ+xgn9vy2j2SD82lGlQwrFyfqpp6y3xPq4CH0Xfl+Ymw3CPs
AVXvq3H+wmcFo1iMBXWzytihN3pmIAkSq2VVGZOmjvwgkNw3mSedglzQExXUQ/hhdYUCVCehzCkA
AoWVUHrF/96thXLmVUwtLuXnvWh9fOVslZ1LXxOWX8Ae2XpgxBD55ijBhFxBx1/KLnyKuppMCDsa
SG1YHWaJ230BOjQrjcx3exQD55lRuNBU1LP/LBNhDhlnexSlgzyKwrUVgVye8HfkxtESx46Pj9mo
oc1eOPEA+Kt0FDWMvQbxmW0TAQpTC0PUJS+j5EgMRtsIvMyymIyuslK3bbATk/XCyPC1pKv8lF6V
WHq4D6FAIx80PfK9N/gu0xAuhzmjU70qbyvb6n6cD3Po7aMXNrLwYojaXWyhdR9sZrlTn7ONhLAw
sUU3KN6uA8ONp6gaOtEWUJeKop04mYaBpA8Me7didzUoB/pMlVukOaXNp8b62RNL4uB2k0ky5IQL
qTbqCKVB08RMcEocplhtN+UzS1AFhnSkKShVVObkhrSGxAOf+tpI3dTlvZN9fpJRsQG/mO/YUrlA
jrEQL3uSwtgYbOJtHOE19kKRNM53465FLUremFZIzzaS02ENNK/jtLBm2JVfHcIpoNlmyRB4gbO/
+vo/sA0+mkBKVTrd+31cVjJm10vC+thglGG/Tx2jV8zXS6DCQiOTvX3sQthRVhWzVX1PuTP+tVd5
hPiFPfY9cYfGctFO19bbxZXglRBPyZpQkTxiFDY9CSpUle0T55FWGtmnR4jXEUDk3/s5LVG4z2/f
kfxsolHVOykSIm+Fff3zFA+sykyFIIAud8SCzqlLeiX+hhR3EttkxloR/rxkfg72fEEpyn1Z3pPl
kmRUHJgUz40+7ARbLDwbLmS0PqoHki/eddVmdJVxWuW8DxxgLGArcleW9QInmF++SO8sT2qhzsaJ
jF8/DxxvOz/TIoVB4ZbdxGD9gDIWUVYNrVZIfOpBksqUGPY6EDbilaoiALcGf7IT49GrSphFeYUC
nM5TljsB4S2jx6gI6N+lZjxz2WRXAqWm8VMX/un9Y8otkKp4v+ufFkZ+k8tX16dsZ2TGWMrO3y9/
zCXio3QcB7ckUncU5iNZ0E+CGcXGxbKyPi/YDF1/3AyezpgUG3UkJNhzBwJHabxDigUCM9PpIKTg
EiTlpoQJMUY4LEPRltM5w0INo4oUBgE6S8XQYvnRQDpVYUWwDrPyD0YJNTSFJSN60wVI58C9tM6v
MrZZdy8I25mGP/gjPxp3S62yWuxYO1iwxnQWzTtXceS12Ws5zvQV7eSf+CLrxaKKfpmReLZa4QzB
Dl/O9VAuIFCKb+qgbBhc9RcGI81/oQ0RjSIoIwUiTZgiFPrL4ojtQFviZL+fNpsWL+UmEEpJDkBR
nhw2x38baNR5irD03YPvZGAL6OxLMhvzFUl+jUpDnwDICKH7lYtqC1++4Sg4svFJsP+L5usmYCIV
l9sn/HIr45ilUU+VHK2RWcm0uKy6+Cg6iUMrRMQV5mSyZvTXrlTPt2gF2BbO2MyRl3kZVOF1XVaf
QIqqE+3/ADpDIhev+miYLQ/Parw5ksXSDvBT23Z4KMU0TPrS4ozFQBH6bVafOooJh46dZQR1VfOO
DUmXnJaOoi3FxIB3TLHWNMKvwn5kj4l2xguiqR94gc3mEZPmEgFsyH2/TOB+ILz34Y49C99Wggc3
kpp1UIR/b4Nm0DaW9KKOBBfcDxBWw37ARXGkTctm/snx8UdAqTZiw6uYZ5M5VJn52DgMwOBxklha
hQdAzxeiJOVUlWXjjCH0+aBbV5iXfZhrD/HR6zvRC2L0qkzOT5SMfSzSYZxefR04fc13WpmcwpMw
whCWKm8b5wYa/OX0wIQAWWXsZEVRaC3j29cqXZinF/GvJYQcAE6rdbnoUYPaqhfEa21lFwNSn1fm
Zw1nmHjrb5jkYnmhWK+9vtttoJuWrS9NA6SFerILzaoR1IJAPfnSUXYS0wNMcE6jp8xfrRHIQVvD
3fs5JZO6Lh3NmjCqhQJP2hA3L62r7y7iuK1Q6cgBoUrjh1yz9cprawBSL9S2/7ircDgoZNg7scZv
WC8vZV/aGSV3QNFE1gWQbEeYu699V2ydPMVMid7bh1JyH+yAT+jaEQAAR2S94+zFohnsRnys/ur4
nkMVad68e2sHRQ1qPH95sIg/1qDSFEYwKrudpkQRQ7sGw+WxyhDo7XHArB5aAooqHtaj0dBM8SEv
z/Je40ZMtzNVnnSHyil6Yfs2mJFvNKvMP2rFYNwDCDVNaaJnqAiRu5bsay2Oe1QFPdPQgCdj5oMl
jTB7S9iyIGJccsmzZfVI5yk0CPLkZi4tr/UZ+MkIItkRoS0ALZ4xag3cOfANppKOyHZDrzNe9n7h
sSDFefhAD5dNDbmwGirol57i/OQq7SaI4WtfaJUahJwJ0cIs17sN6txEnf4Bb2eP1l2NPlQE9C89
tnoV7Rb7jOj2OjJhi+ryRJQfg6zkW19ypGqh7R2wP9CHx5LmOv82TCMcYcuHzAfji0JLJtage55K
5omymDuKPmH353v0jgnmPRudWzOoF75bZKn7XqidS0pOLD1FUwnvbBPRZjK9ouOGLeBpzrUvSIQi
g+8F82zzOX7OtjeHVwf94feRWbuVy0bteIZWfnvgBMZBuEsoQVvMmxOaYFaTGjGfgL+DmVLt5doj
1rV7ymxmFwUUu90cGZ8Zm00b2K05H2JfTDepnlhKPjwIqF2vWNzIMNKRbcmCmLb+ocHtZ4b/BQEH
LxJnTQVWWHQVxXCN83bMh2TamDOaZRc5YuYVgp5mOaXOVDtGq8mGOkJ4g7dK4SfPgoVhywz0TtAt
51vMYMC4IJjot9f+xdwPjaNFTA217DfnLEze3TayJGwDNPJUid7iX3sr1bQ2eSihMSCOHa3nvmIM
MXUYH8ohPXUZWS5KMR/izVQzsSCuI/eLEAYC+y2F3LF1CgK+YCdvYII7RdgXd7jUTBk3qmulgW7u
8URw+DGxPwWYLu2bscsUIippyZ4J62l4Vu4WJdLqtj6uA1oE9Exuj137tL07JVlU27caTVgbvKrJ
En3zbiQdGBBQufABJShOAUD9oN8cGYbsjohZEz1JxiL2zRWnRsh58hJP4NO5wT7HbRRU6HEkrt2r
R2maNMcm8TC6uvESgPMCwhuzObGr6e+edLkRAH3mwyGrCw0EP15wgkad9efwEf8+7rnyDsuIEtDx
iTsvPEITpvvKV6M1Z3jFhbnDGr+pzAVAB3hoUuFGN99rkMDnY+sMVuVMBnYyG4OF+TeIoNB8D1kx
CWOoegUC8i+kF4DPYdKmSw5c9fEO32SMUQ0eF3ssobjG7hL7gMPdemKRspNutKWzZtH/+zX11PkR
Lr25wEGRkTUVBKyg4JVQH89+zSHhfSEAiMrcBWlG78thysXyzoVHjn4sFRmRaP4AA88t/Rq4/hWZ
eHDjCkBpfll9QqJTmYeiSLRw74zYnfG6XaT5SnP7EDS8VI/U8HSl67szlhSpHtmrQN0yqFm/VS7E
a6LmIQHkPbJ0BnhiOtHP6/YbAWXvszV4TZk9p5jWgKjYlxnW944krKWwj5vnBd+xPjL56pQ2Iy1+
+6Wj7Ze1cpWS8hLHyFmEt6V0C5gxIPws5AQEJSf+jP/WEzKe/tLsQInD+hkO/of7JAIdh/c16B1r
kS/38XtAvkumPM0X4WY1AQG7k/APs3yOb8Zt5HjqZS8rLDfY2zZbsqDMoLnQBBEVaB8je1D8racW
5QBSp/Mkt2Sln3o5F/sK5DjvD6yH+QS09gua5mQRDju+ZHeoqujObPGVkd+XA94mBdUXG3FO22l+
sjHn3UteAeQQxU2cWF/Y1OD+d3mPYqBklcu9RHQQymoQFo/Rkc7Uyqao0Rh74yLf8c12G9UFHhlT
vqxQOrNd7yfGNKqJicudD3ubiGfnB0a84Gkxa0lwCc+lGqRYO+ys/cG/Zg6JaOkOF9vKriKbMAcF
mbBZwKBOhXRlxPDO7z3kLNclseAjY8NkkEkIejHcMfRd3ggU9+WNXfsQ1jAdmc65N/MjMxUEFGVQ
4aVGd6GrwksifrL+2SviueupJLG+P6wM1T+GbQnngALNdVrUVlgiGHti7vVuOWmGa1okCe9V6QX3
13qe3T7riPRgFccB8zm5TzgJhTijBe9kjcSI2Ei+ZD+s6dvjoq3Eo8pSgM/yL6xeTgb/skHMuzUp
PBbtDEuYkBo1vX1u6hWdwPB77lBdCyy5OAh4n3UeXQdjqE7okIiN/8WVQD+7jQ86oBmCkY8GV/Zo
koRyYWtEAbJ5jWS/jzgMdasAU29tRbcqgXK7h78kjWZXPMgsvlCqQP2+F/csJkVERiXFVBQLJEZF
93aT2o4B9YY4J7LBKG0Mhi1JW2CibYbKS6PvdOnWr1fmsboi/znLJY7egjXyNWGJFu94yoibtNXV
X/2AVI5Vm7CbL3xLxrDz6XjRwDydwUd+YtxCKtUC173znw9TTZGOdgnl2D2bR9WdNuzSNNtok6uS
KW+xjBozfpDq/MSQpSg07V8WUUjPOeqxafUybs7zSuRdBU82p6LDSKmMq61HvQu9RL/PlAXdb7dz
7590KCSllbCUQrab4XBoP9FNRY2pbhT3TgxiUp8kOiir9YuveRBanYZ7wyRBrTgI8DJGjQBLSzeF
vDeGcyv9bPC/AZuwo0ZyS11i7FTqcUkj/CIOoknfuwgDPCRC5DSs50FmkKmsiKoc3FwcYgbkX9UE
yqI8DGkESrfIRD3WJ453Yz9HErl6bkJCO9zwIV4TasCueFV88ICaXHG1LFv7JLiGkrbVZQCegjxQ
kPYy/+Wtpf0XY9BfPfdPxSwmcRtZA4OGKoEVJsjjlSemgbeO4ZCgPDpVQerjk+nWdbZTfX8YVx7j
eUF+DpmY5cOG9W9oYBzvakNyBiac32J/puKoi2d5l8LmR3/VgYbh/0HpVHFOJWMW7hxR2B7siBpT
+iEQpoV0VqI9W93Zfvup0zrt+ePId3pjpTMyb/2XZYYCt0DfNMuYaUiS620KcS9pevE/d7Dgrh7E
WRRYnazdUctwJ8VPBOoNf/kwrcFsruMiKl3/YB5AqtMUQd2HkRQl4Eo5b5IQeqjOBkVuNS5j4t1/
bydaiF6LmdcxZT2uNhc54WnR6Q47QcYzzjxUGM3NZJ9uQaF4cZG2+VcmQpQuAa0XSJAzINdlg5Ds
aLW4s6mHcEaiyxEHxmlLfKVj6V7JWL3Y8uj1XPXcy5RMBX7c+7nCzQ8tFSQvl0EYtl2lMAvF/qfJ
pE/hleaNWk/sEErMxeWRVEwFnOIid2bvCK2ZdNEY5h9nOaCzneZhjSC5UWnACUMm/vqKXMrplvIu
hd6vvri2T1OgSsUkP6XdGT0Ql/+0h/Wxu8aXATyxVNHdIT1mafwO7OlIBWhwcSEmd61/hA9uRL5U
9msbiuQCTYS951uLSkRVKD4ET72+wba321l7Ew6g773+O4pInihLe0PcWs2GMLZ9pqX7sN1TphZr
lB4qoVynoyFEzjiWN1AjCtMBEuv2Gy1YhdbU+yvGaf//+wCf2w/8DQH57eXGXfY3I0b2ChZ9g/9D
QuibL7LrYTgQb9pTMLuAVPNQ0iHhc34srptVpyZHSvjHMBRFOqe+GwuG+FSvZe521cXCYfHempgw
YuTD5ROEjy1T+/WEjxvIxpmwb8NjiLQeRnzSPeX+e59ZPvTB+VIxl54CBebkCi2bG7G7aymFz8Jm
lUDMIyYT7Pt9Wx/TzQYp3dCMJ/BdroddEByOgy+Dzj4hCzolNqIT3iV8246xlO7emJBqQlw4orMN
C0lJygiym7d+RNvUu/cta+f7vLoD/CanL/7JYQgfvYWORgE1wBpmTxEI5gLDn6mTsQUOtdZUSZnJ
wyWrJ9fgcny/gLbHpczAwVXFZOCG2BzzYGSpG5KMzISmsi8gkERkZo9wxIxgsrWaxpR/hGK03G9L
dVP4DlE9o7RLRTfBXI/zuIemYQ/BJXhd3oysnjh/Ty8nyoOqN52jxTkyy1HKyNInfX6AV3v4tzD7
X5DpsvjDinZzILNR9JsmeKKOXlEIDflb//+4LgkenbAyJWt0ndVdQj2VQ8uZrZUt1JBgm8Jvv6fX
YzTV797sQfAyomAla8eZkUVYxZlmuvXxfThzA9LhbjBbYCZg4mgkN0fR/BvLKXkgyofZFsirHOWI
DSH5ZB1H8+SV/AJ7yzn/zVDwXXxi1BLJbe7Y18hin4WKhAIYBsXLX7iudxnjizUe2oF2kGRcNNaC
MyKV3lC7k1i+zdTWLA2j6P2iLGDk4qJLyyyeOAfs7L1WqpMmcX65F6Pnr7tUED2B6DoWb0JcqBSh
Dv9b8cPS2DtK0IgukEmPPFlui/ouZmMow28Q7Efq2fRcGNkfWQmIFOdUix5jp76xn5aYSzc4DnGA
Ls85h46xId0iQgWoUVyvUmxw38UdCtS5MnZ29Hfsg0K5h0ZK1ZqAPZEuM1Xn6YpAycAl9ebukhNb
ZBgyPLwrceIOZdmAxknI4wDth3+cl3zMVYMK6+b7/BNHoljixaBPSULSet1OpHtVFpyZz1hLRvjU
a2MvNxWQnZ+vWgYmde+Osm1OnH1tmHZOxUAnsncsvGAm71bg8rzTXwOrGKtuPPV+X9dA+/7eWMhy
1WOI+JVrF9oGSpWpbxLHUOxta6F8jkorsJyqrXRhKF+dwItTPVGm2MLg84vlUFndemJ9jOfmIJGt
KBKt9oZ+tUEgTufx0HGkvW5VFPPH9aot3igGzqmePDyJsT5ApE2MupZ4Ogn+DxJ2es4kqL05mKkj
iHepNjJpbVRIEBzEqq5J4ckVV8od+Gwv4RY1Eb76+HeP6Z57okGnUkSqHXWXhmwpxArErrCBeM7i
G82tRmnC4jSmdRbKN7jqhbIeyU5/KTFtH8SNnatKe7fM4NaEDy/+GhEbc1mrIrva3kwTjqqta6/u
nk2Ni+Ul7NjtSqg2OCn3ar8wpYVbBe3l3FZ6nA2dS0nXFUHo9ORAXj52XgK+h8Ty++OgQhjo4diL
7K/J0nJ/4Mtu6gSA76LAcL7QVs4GJv91GE8fjaDzoJIXeg+c4l6/aYAwW7kxINykm5KbE1wA4mxB
aNRk8k07AIr95HS/CuY1ETGUZZD7cDdl1IAB6XVN9NznyIqijmPPDm+Kh7WTHyXSx0itrwvdxH9H
xaTKX7VlLHGd0kuPGOiONBf7t7qwYHqBPxjj71D2E9eWQA4FleR1LenYE/E2lkvRGVmsQGps4lhw
dXKTks+ZXo99iUBqbWCBS4cCeFRZt4jK1OddiZmGjI9Q3IE5C+T3epk0QveAVa3+7srFzuu2mfWT
opPacg9UM7oSnCPKUIw7l2wkL3qfEvbSD7sOG1VokENtqjK3NGqbjPhYf9MBdGYQUVSdh8hpMCOI
bSJV6KH7UmLMvu9Jymmft4SKwJud1LtslQ2PZDgtXVqZYdqh164LXjLwmWjtfn/dXEGgTZ8bD9y/
QvN+aOIIvMDQjyKo8nfADKxXaKMumepGQWxyCYStG/yJuLhS+Y7NpNz2uIukEMEoRHTWtYJGBFxw
L45v1xAbae1K1YeM0gsKyWIm4QGw1KsFSNWIfTdkOMzIC3WbDH/FKJh99t3pFOm7NYD+BBAzknxz
nEH47CfmQFHOwwkW+5bhn+HglAp2Txq8HZr7r/AWLAROsTZ1FK38tuldFtpjKSYgeQE3HCsRJ+3L
zYvHcdOVmZ4yTJq4VF1gtTHIust4KN512DIvwzgBd6EiAfMwUEAVS4QjlnhH47yJJzkqij7/ZmN1
YaPTZbX/gz0HRZSuWNfMoEaoMRRaF/IHUMQbfRla6slnXbvHVfh0ei5h/WmBUb0VVhjxVzP/Diai
Bm2RqTqNopz1smYZDHZVnSIQz76QRMFUhhMN4jmYvAf9SsoZOu8QLCJgLubNU6G1AGurcY1eoGcZ
Lo1HYZ77WIaE9cUzQuqJQouhQHbYqXlFWJeqvYFKy0hKYtrtiXvBcS6nd+g5Tb6kI9v5FNfU4Vuy
v8K6YQV5+pXn7fL7KUPPIgYa92YJ6IepAMNjiX03hnuA88mpGLGKHr/9xQImwhktbG+VRaAIkjIx
4RaanmXRiBkOn4V2oqlhK8wSbs3OcX1c85SDcd+mF29xbLSkGrh9ipJQLNlAjMJ+5o8EwiSDzsCs
WTWEgwzkIOjkcg20OnzPCUehhghlkTmLvJUyj5mKurHqZJVEgujLM+KIVegUFKNuvTB9f0WGHyfk
FxkO2zRvLtr1mk7t9Tm+ps93nVp/t8w6kaRuE5+DJ5goBmC2E6ODUkARM+QzJSl8E0PnaTOydDxd
7YcJWiCeBfPf4o9uKZY7CXpEHU+P+F2vI9gVydywofp6nr+PF6I0grYBuOvTVXN6aiyrQpcP6ZST
nfmX4bAAAep25L3IIjfwu08puZ8csSuNeO5yqqnLSxDYSvYHk0c6XpqazgS4YzWlrXl389JJykBF
yRjynM0Y+EMJ5F5A9tqzdejjYIbSoYS0WMu7JGzcDzeyuV2GkwU9WiA5dJ9tcV22wTRAY64i4qjV
yzRFiTuzNqdorRtLsAwTR600wYjhtthu/FdGpWi5VnvOYpFjHskJaAuhe5yOkMOqxlILH4716UTr
V24kUhH/JuZ4Zujjq0ni897gfzMluhwt8nZDpFuErp4lOjsvR3uirtPk+Dg+LLA1PU1LpL/xt8EP
K1303cucOjp/P1LLukzZ0od3Nv7g88XsBnsfIY5eZiiqvk4Uga70bx1XlZxMXUAujg86texa4hci
YUOG7KNY5hDg32bkpZS40up2IQsOBXunX1LdvRq2KH1/w/DogIeUBGOOKocmT6ccjNWKPgaKCrGs
sqJQ+uLiNE0thdXhBUXmadSOFtaQko1JSfM8tBkN9jybQg++aDt065UqNdphoHqK0UZyOxd3+F2W
CHWdb+mTYPvx3tYskUIViNMQPJOzdeqmxcI2pZkZZigu742vFOgeXc9RHY5H0MKl+6bikHvtha5o
cmiayj7KaHhy6P0c1z9Ju+civ4QRM9ahgUNDqsd00GHmDQ5hnT0CyruS6PVUcalb761qAFvpcoaY
aRJY2hArvtkJLiwwEOVFod+edJcuTNcrdsQSiw4wvM3qiweoz81NqkhVJPAsOumGI4vhmDCrH4GG
+Ah/0Jk1G/PHnqvDY4LM21CAke63QFPWLJwhFlvpy7k95bMH567Khdc69Z68Sc8RQi+4yPcTVBIJ
WytGK5xAWMbAWD8q2HdadEC3Oo6CGRDCyHrVNlX/4VoN0kikwlopWKmRtU0H4Z0Fy0abLKAPelDK
k6poL+auiOMhoHtF+W8r8XCigSxcDN6hal7S3kR8sH7we+FcFxpcgAV0kzkEQZI/b4ht7iMTV8sk
JPKGwbQ4mgZux5Q5KcwMyvDTmaRtsyUzhiIFDbWAARPqE5qvbl7d5de1530rzMXpm/wokAJweGuH
djJ+sdi/oPyvyWw3Jvzmv7ukxrFfbZebSR57CPajmx31KYTLpb9Z2GZvcxiUOg3BnB6GwmIq5U/5
9eMVcK/Xc2WpOC4yCYwGWENbtYXL4G5lHqX0yl1I/KhIljw8+SWJqEqklr1siRPUkykqwDdi7Z8a
Vqf4A8RGWuY40DGcnTBvTisvf2mUjusn+GBuHPpA1Ta5LPOv7wrjnsjhKW6nTv1nSZq69/3pO7KT
NbxAuFbChysgkcg5XVWBMN6iYzEqoIU35Q7opNwQ0Gj3EQ/zQleqvH7wbqVfYBib9n3/Y2X8QKuM
2dNiENW0zHHZ16PZrntt17CTsN3RkXEDC3J9EnqIYDED8cZWwcN95iR6SmuwWoZQXTyoZ9qOUGqC
mMUhKeVEl4MGKJbgy552DU+yp5D9gQbiGm4+09rVrCR1DA7Grv1CwkFUxk3rdoCheVBxIAT5hV/d
rPZFEhch//cCTp2nMf3eIYh2GERl7mQ7yrvNZauzOZOyQQL2ICOZTacqSNS6i90GZHaDKw7/dl6o
dSazlTpbHVxuh0/szSx1/9Zr4ZCXXbtedatA6JUk+ZHbLPxAHn5W9YgJsMV9pARPCwMS9wISAECa
2IU3JBGXjDwEad480JhB06jAZ7VgODg/e+ppElQmcjQ53B0iJorfaTSZDl9wO3W/gz2lZKiJ6tCF
WFZT2nxkUaUoeBRe2/FQ26pmwEn1qWK9X0lRZSyfdHqcF+7D7biYyUj8KUoz59JFE+N0FKObVcUo
7AqmYTm3S1tPvnASeyLIyPFcmBMC6WIWvwtXu2fngrUHQ2fnA8bIAzNVusZmsBVlRtQLZT1sy7d6
sHJs4Hg3NV8+lA0W5xLsClSsTXJvvucBnzCaKNdy8IU8620Izu6v0B85/FNeU/+0PGiOiEUtm0/J
HnIQUS1/xV7b0UdI4wqBVrYYBxSn4g+bz/4pw2osKl373AWb6AWWu+YCajPXNrlxDD6N/jo+fPK+
1AtHOasAESB1tDNrLCwExbAVrHecR1TUDQp4UWuclbfO6nvyCnjG4mtjswsrrAlMdpw7/2K/U2Rz
QTkyIKBYwgHn0lSVS9cH2CWPiyMoNi7O19OkTq3N6FOzzncSYc0vlTw2d9T0I+Q3x5DXdBD3v3a1
LYRDyzTJEUjbcjfSdR5A5bZsSx9cMTpUQnm8tZ9GwGd7V/qLtvHjgK+2GRyNaUpezpVPicoe6YhL
+lkszmI+dERJMrRe1ndAyMWeY67QzzqWB45oxaorj/jZOZ7JEvncEui4V2pd9X1KDPwwc+Lsj8HN
KQi+Gvhk+iTZU3cJADeZJJQHOQk7iqDCyZa7+RsOEHtgNA8kZMg8YOnwyEjK2h0EOEPcAXjHW/Kh
6CaJi7tea2oFLgpwuJBXEnJs4sr0gpw9JSoH57LYA5lpCREk8D65Hg3ekbEntUzl14DwuqLHnEQQ
TOnbuaoiB6WkyW/9EBAZf9OqSwvnIOfb5epePFxFeEqf5JmG2rrVT1X6q5r9pvzHr3JM/Fd4YOq7
vG3xS1iYDr68cibeQKSsa4l4KetjIlHO5tJxCGk+0qDrlbkylLcX0Z/2+JHHULJwOvgVFj7+ayQH
DZuQfYxiA4dTjGFU6Df2QxOycL83jbdqURe+bk1NLZ5n8BEnAJqYWs8NW+GrsXaj82QE4fCp8Tbn
MZm6RbBETjvCC75HpSDcWThFUHdw6gdyBpeh4slHQAEajltih9vNqHM+sZIw4yRMUVWKX+Ad6ZK/
3sFoipzIZgkYIWFJ4pBDrXY1HV6rPRaeXJybUohG6uhcqpbXa5wA0N9kFm7ajxR9MRhnI/3mNnGk
Y8RW/WRHD0dNy6tgGchzgKaVSL/RqchcWndwmjj8idU0o1Kso2cnj+r77vn99SQDACzYLhjfRGxi
neEhmf/KFtrk9XcOvejztLrt10YvJ8m0OJ9MUgZuWMm0rHuYDnYk+agzlNTGqZ+/jyaPzJELilE+
8BWhRBPlTIXzFEcf53DAexJQqkYtm9TooN/ojWbfBucsc7JSVq2ACIK0BkEh/exNsa37CTIHQIx8
Pu2porURDNf966Yy2ZfuDYl8uTGkLnFeOJ8+xmnu1gISY/budYVv9EN5vm+OQiAhKy/S4+8pp2vy
LRXMPPj0WArL43XGXz5kxIdQJ/Hh/6RIPm0V5bKZW/hNHS8soCxFymXE1M9GxwfocjhqophSy7z8
Z9xM5ECkJB5LUCe/7/09R7Q3tX0+IXBo6zMj/mtOWnTgkaRS9DKMaK3wJ+J2x8bS9FZT7KHvggCY
fJU17uL21o7XtmJP+Ax+kgolEalAu7EFUe/A1/ECs2lyF4hS/Q8HjuCcxUZbjiqRWC5NzytTvjhm
iRy5jfdHll1Z8l4mw29U0egtUn7WeSVeBOUAG3tyU9PGRiiOsJvQe8IDvrfzhrhv8rvKHe8ou6z5
3S+n+UErgYGz2DGX3zzDB5NifLbVHaBzIo82V69U4qp56dM9U9VtXXONdAQtn2caRzU4V6fXXKZY
jvbjASCp507r+M3GolX18S8qCNTtJbr++PWO7Uyxgpzqxt8yLsCsKa9id55nLZXbbWPUO/67pNv9
I2aLVKsMQrjQHM2SP2BTy8Gc3fq6P6PTCRMNon5T6g6lZky6q1nNyfa8NddUDpnL6oSYw5YXdlVK
oatfcjqgqbCkD7jP1/oBBUsACkxfU9EDIut1JTJu+Phl6Wz5bEU/IH5ajxu/uQwhpBTrgvGqrJDv
AQpCdxKE5CZvfOKm5+cSWSlQ5kn0Z241n37NlxQ8yIAyv2hXwM/ATFvNh8CJxu7muIikcAJzZQOC
MpzFqokChklu4aBeuv1TsLu4+nuRS4K9Jeh29ijmlxB9olmCMhpzpNQYly6ElaCNeoCnNZPbF3jp
W+jR982A9R8HqlZCKfZAVfx9hwgq1wEUjpmrK7AjfUzjyC9qVT6x2LA3F/2mrKRY9XKKnJbJMQoB
vXJWYIMS/YKBg3JJI48lBWTF4x7rEUn52JUinzT+RnyAMxFSOub7u/Soyk/zCblTnmv40epnyA2z
T4aQmYbq1rjlhZYgWULCRtrukRq+hRDsy5EVRJfMA2Knurdq09ZQmT7vb0s6mnK8PSgOO8sliElq
LNwfjLkX/w5vFs1y3WD0FlYIjVIoryqPXvsHYeyba1F8HJm1IzhB5RAlh1MQVrVRlQhT0IoqtJaH
aN0XkgpbI1W0TKYDp41zV1AbzAkfel2P/55LDeKu1fFSqXwszsk/Y/Bs1NwL7sNninLFyws7lWFM
xpPOvJBTI20Wbl2+daVqaIzqmBhmlZAE9jp3pJarhEJMh/nznccRnVWoIc9yK8yEO7pAVkm0WAzf
e8pyyUdhLcrLEClhi2rOpqqXXW8yXfZTCaz59BlRrDNhfLvRBGXcZns451N2s224ALwTGJJKUV7y
VvsryRjpVHQI4euVjsD/L0h2gRi2RiuPn6FBt5mH8mL2srPSPhhvNxQy+G/72pDv/YkIiQW14XVf
Iz1uYkob+K3zw3s5jIVkF7itKy2IWbpzmT+c5rrI0iO9I4/w9wjd7sYUY/7cTlBBxRwzj+AkhgKe
0le/0g7fKmjOHqKSae9bQmNz8DvkzZ0hw167FI7NjDqeaRyOWAjP6ZFOcO57luWxjGux+R7m5zCm
cG1pZ55KC5cdK5nx1vWfnPwh/bAWYfUoJ95EhYTDXaGbFGXn85K4OkTCFJ1sqqucMZ4z86Zjbel5
2f+y8cqw2B4dMdOcwn5B7HUl++wh0JbyEuTaLlpz6LekS2JMcIIlOpFoHY2G7wVHWPDb8ejTWHtK
E4NZuFCR/1kKDfO5v9MjnXi+eDnj/6Hy0aTtok2D16OJWdknggwBy84RN94pTrpuWOLiuJOt+PGa
p+XKD4sw9/iphs1/Q4cQQD4N39IlYB2ozQNTNrI2HpHiBkanTPcmHKIf4WzcsoPiEBLJGWEW52VY
8t+ZoUxpcKJVDHwotuE16Hnpmq5EwJKmhXTkpfWR4VPQI+xl6co26jhrJe8O0PoymZeFK1jq29Zj
BS4QAKxv/Rz4VfhxLHooXF4l7GofiZAUgGty5Ur9uVzQmb+O4Wf6X4nwx6Xh8g4DZs329A8giMDA
WfZ6wTSaSg7SjmwaXVpLvBqbb4KDG0evnqeuwjTYGkjSWUCbLTyDuTAZgkXAQmEPIy/IC38ID9Wj
QGq1PMyA2uay8TqMkxBKYUJxJ0zUc+yCCAhoxtm13COf9Dsptd9zFgDi0XE7ea3tiZ6DV4g9lWHY
tTbfGAaAEETzE7EOXRO/ddNeF6U+/Iu7XVYpV8CFPCWeVW5Mj7gFYr25cgMgBVv9m4ed3fp84VWD
AKlTmQSVjUnE3tHVxWhTEz1wOZXbjch9LHjFvvSOkz1ZJcgV7yHuLBOH+QIgWTqYJpZLYcnaQ8z/
FyumJqPvpiCu0b8osEdko1UJF1QExfS7IYRVu8qPs0nodY24d88U4HYX+5JXmmHO9Rw+qNHbhA95
0RXeLzuGSy5AfYPKKjWDLqrNbTS0Gvq18IPiov5fLW2FCVgnK+68QluzQcMGQWkev5cW9K5xSjp1
1EILR/QFp1x3FFNL7QUMXgrJ8EJG/k3Qat9bmtOnF3wlUHMlL9lgyA+VApzcuLpLkJry7vzlT9Hs
Scs8oaNRCg6AzGKgs+jV+0pkvQrBr6Wer8MEN3y81ZvYZdRP1kA23YjAaSJKNt/hsTQ6+cUi6AvG
tMZxv7VHbodryPi9MCh9DSUYL8Y2VTr8Qgg2id1w4bk71ETFb8PR0WL/By7YygnPon702kMSnBei
fof8lsIZ2i0EET3WC9UI8Z06UlZDRrlajOFgzDIIHbXHUpKIGiPWAHo73YcDTwVd5yjPD75chlJ4
Ee29pGrFnze2Wcydj3Z/R1JV61QjL9w3/MZ0+EfCBKKYNj40fhW3ydDmBysY66MF8I/X1O4zl4N8
20B3KHbo9kYF1DAGOlfmtIiuOSW0aGsQwfWrFJIMBiA2cfd3eUWBnzYMYj1jEOlsixK4fRJwOIjz
ssvUPpeXOpEG03yTt5Dcn9O1jO+s/b4e9KkTWhR1gS0lH3sX6xR6SoGttYfdpj+sZWYOkEZFkU6Y
gdg5J8WQDlx1kG8QiMFLecEXEhs534aHVy5ksYx7K25cFBT5z3WG3WDGfNd41O9cm76bJyIBgR7e
3APW2Y8R0tE5XBDJL77UVqwqbofugSKGpQeCDoyaMhvcGxhIX484uoQKtNixsuFikBDHkoG24rWc
Zw1Pn/by2MGJi8Em1/jiCqoq2mAmNyKXjTbUmhpIgob660ddklhcxQXT1eUGYmAYKI6dIkpAJBL6
oF+OKzpWGb/xp+jq3tMENKVDBkHLLVHpPaJtgTMIGGdO6TwLPWPZ57ZMqxbTcRfh7AP8QCnMIo73
92IO0wb5zc5njSmMF7Gh37Tkoop8Knqsf7OdWRZ62CVQ+srVGAGRe39GHaCq34ldTiJNFb2oM72J
2YzqPo89yDt+GDdrMxrHxpVUqKZ8/oZi3bdwLv6haJ/kCrPyaJiG5b28WJ08quW2aiRQq9Rk0Odo
eZTQ8HtVSjJUdquIeZ6Vbg0ojNFXoO0dZWP6SxNYF9EI9qGKH+oB5m+VfHLJ+RhxFM5FPRAtT7cm
2kTYm4T7BM85z4hdzH6Va2lCdgwvV3wiQZcNTDyrnXk8hcz5H8uVUF4pt8+3k2OnyZDz7X8wNzyI
NiB1pWUPHMVvmcfuEqxJmA+NsdWezwrFs6XEU546hc+veKXGGl9d/jrpEOnGV1livU8fjGvWe5As
dPJvbQgOCFuBwFIGSP3WGiGH2QCzYdQGitp8j17lY2BOQGMIXRC+H/d6X7hwNc0lNr3jxVPqwY/E
tkKjt92RMXtLmPNVu5GnZN5IjRYEkkFK24MSXnOXcILRKlVFhu5vJwBI4NKDvrDqz+B5JI90pS8+
I7mbLSsuFikaXnX2Ub+87i1WzhYvXFqJDYG3YU+LJroTugzUownKkEaOjpTDfCt7kpDQIlDS5sQu
NCZXw2+lGBce/zCBxOUp6VxXUsWrKBN8can4WGMi83TYF0XMMqbkRl0qYE2T4St1yf5/KJ3GTQ8o
vAwpznUcj0TMSCP/cOj6tSSE2Ke9sSwkUg61e74nMalTykAn4utH/XYBGC5WPWVLyT5sfbW2590K
JjdyrxQzx6GsvwlybfrHO/3QkPszPHwqG4piMKel8YT4Vvn1rknsSTqQoJ5kccLjv7zZyr65NlAF
xDQFFX8bzUViR1WoWqc4U69+DNgtiaVaYQPxtAdgOZyUQr6Pxt8Y2hD67F/RLCDhUtT0GLhiNm5n
8fkSmZ6n1YYqdkW7Xo7z1eWkM/rji34kUXT57hwZNAZ+duEU9y4IK7mYe947/MNsQeyolHuuUGU6
D+uA81vNpXXYV52fAmoENEVsARGlCUZQXrEwKtiFo4fpAFMGydzayA/20/n/Toz4aCFTHgigIqKB
JMUk2aD1qu7Hc6XHq7VGkOWoTK+vwPYucDzXC/GuMlIAVT8vyzmoL9WhzNZFFerPxcheqWW7u83O
EP3QvNkKt2lsQM5bCIHRruxI9FULfM5IJucVGx8CGRkFXi9pSVGq8g+IG2T6NVuixgGpHvt/5DXe
SXE80qj0QmSjfE/QW0pYaQGs+2idTKtafVlvWUVv9y6BLV6McKrZ/W07rgCCjLthYpjtWy85PZAX
ExdJzDiiGn2ES3fBPVCblZpnwgLxUdzTh5vCu5mWUcZS+dN+AFysVhe86umfronppQKJLg124G7Y
2prqn+SNllmOJioXejtLHJyoROjc5Q1nIofPN0SAaD1E7N2yzJ2faTiZ93Y6XkIfj1D21vnhyXdq
+iHjaBfqASEPKO1/ZrH0ruQW0RMcwv1M7YB8ScJLBog6YnC8mDp3m2XlnFMIv/x50EfDhNOwItzM
zsyANsav+j5JD38M/iiAuP7APP+X+mSrleg3bwZyXOvvvGQlEd1ZehsvrRqGSc6sOPIbK8aTDxX7
buf+hZ4ChFdQReHp4kRstbMh/CF7ZLash1Jsw3a1QKvDYg05mBENkUSgxTBjhQFLrfhwjZdfFsEB
j+n+vlFPEu2pOs9Eggza60zlkoZA08KAYURhu/441mtBoav/Ysh/e3RkVv5OrMdw4cY8LrIylNOc
va3Pb0QRMldgSlqjs9Bmt0Ju1ne2Vilh10cHioHSRMTlY8Lw8MpT8e+kszfJwQQVIB/HMLBQKIVp
ul6FM3VhpxhIqxXDJwpr5JwZJodcwFDb0rI86lh/lE7TEAHdiZvDanNA8IQKNaKbknBDsy2OzUGC
70pQCShbBmx4rtwACN0ugnQdYB0L/jUMYgjdv1Q2Q/m+0k6BMohymKORvC0+rNzbeultR8PZCkuV
12gToc7dBuBRIda++MKK8nROVG3SeNvfM0oEP0fMHwkLYd0D543Wex822UzhFo8FnYdEEK5N+Zbu
hin2oAkKvF1asH0QpEE7bPUD65SyJ5FAwY0+4VPKEXhCvCwEmBjMGM3/U5sch9gY7di6VW7pbJ23
ddgopYQxKUB0wNqZlIiCT+Pej073/MGphfk2a/tRmSaAf3gYGfLH+B0gSsrYgvkIZ0JTFXb6esK7
o2vliMMG2agPkRlSSylzIT6h9y6rEvbNJrs2o/O/Eunp0PH/WwjYCcUwrey2vd8hMn8HxTHz9KTD
lAdm0k1/1saQ5hCAwscX3/Q5W2tIrneuB3/70ai06IoCH/Sw5xeB+7z4M7X6we51RLuUz/VEVDDp
jvWWYqd0Jx9iT8zhltE/4WwBBZrXWqGep+EsSZYxnty8frchEEV7nGA5/7rgbrOxmptM2AeuhWeL
nlEOB4TI1yX6Yq8zTRyKgTH2g7Sl/+1TYd7wCtQpjaGshly+HE9dN51pUCugdxvtkGK5uDYh03bb
FkLnVLxNgrEk82vpZSUAszn8L/jQ+W6SF0vtxGgBXWOMe0BF1z9p/ayoS53DFjb778WYYHDsUgJt
uMFhbOuGSqAV001OPsEXP4S/0SIFuurPN8JuilRGvEllo5PsWJg+HXLjFAjTMFvLh6GPNfcUijwy
2jtR1yvzkNOHvOzr6aNFfmCA6kzicFreAmTJJiKpCz9NkBa6BFdwr5hJXVDQAEfI6t7Yb59UAdSP
jVg/EGtIkbn04xskluLkuJSNvF1EHHDbUhdQgp65iv4Rz3izCJBbyOYmDBBC8EpSXliHOVl9yKkx
e0WbTkgJxnx9+DGdjd9UdQ83GZq7LclNhhX8R9f/35Y/iWsOVELSPYK5FPC1lttNgnPEf5uBHtom
0c5D70auBv1FB6lAj6AwWBQhoG6Ul4MEpAHGaMMjJ4i5l1duUkMk5IVljYaC3cNbJeWqsxJBnjOO
nLloiqK6FuKBX1YsYATJh9BauJC4zP1JlfjmFekpj0JXj61gs29KJ1C8in6vmR30/HhXkkL9WSO/
vOl+xDmiwb0Sa1KsBs6CUaifpRTiqTkhhp6s6xRQSKdzhVrffGDEj0g87E6HnlSgUoLkQAv/9YoK
av5rbGQULtuxTlvFxLWeS/vmyX9eiJPsocGJYHYLJIDgvXh8q5iPNOLHyy2EJ98InHlTRpB1wdsi
3buVsefuIVggJXspJiD+BtfYcVIXhNei9K3KCEDITNLziKw8FrZIGVCT4L1BKTsNMNimWxVs+WvQ
VEQMuBcMviZgdn2xKuarhqhQy7KxYHyskXHkfGEvYQV0UHHTS4UUM5sAnAcObJGKaZ1Hn8R6OVm7
hcYC73RfMFPPZTkkX/QQD8HKAXZhb5jcOC/GyI54JO3Y6CWsLmSC7JdtMrGadD9CeEB4+Z9MfJk3
0l/t37W287WNb2hN9OCvvgjItngd4CjbNK3mvMvb9SdAoJFDsTHZqyOv1TR7FRRFpXH9fdOr+LAN
57XaoRUox9R5JCeGg6yckMiR86KhzglNTE4w8icEs0xsu9qTK3dV1rPK9UKgiGQ+EQmvfuKDEkgb
/dTFVe4lvL4EtdJKSjMSEdAvrzbOmV6c9sG+vq1aKYxzgxkWTWcn/rTRZttZCmywl/I1oxCYbr2V
khuwH1rtZtwCvIQGmBEQnTxKHS/2R5cH4OVGS2eyxsAvQ06GEiFH3ti4nnh/h4Q9oOZoneqh0OsQ
74IQbiQXPM6YusiobMftPtmMJNymRdJ1MleyUceZVKWTmfRGas10fqYH82h+Qjv4tNzW9ievseoh
CP4DrsjJvwjLgbgDYMziNKIdIuHwcIWeCCQ5ajqlBQdULDHWX7/Udy8PAwpX5FVHpm2FssEbi6X0
Q9u4HSoR9cvwfaA0+Ewo5ovrifCr9wVwwetw7ZGL7b2Uqgk/COgN7CvD7TvYpaS1R7tdpnEPsVp1
+zj5wbqfJQRmi58qOAf81i8O/ztNR6TBJCOVKNt3+aB8IBe+xbXxNMwyXMjl9hd0u6QH8vbPipmN
UuzrAm/3ejiisOJNMMN40iEC3T9M7pLh8hFzWer0+CfJYQS6syHCl4hchwGh6I+BxCbZuepNzqyV
YHr0wbz2LiwWG+/vzwf7RCZRTfF88aPDgmrMUgksRwhQWZKJxvJLGEyOmuxDZZoAgYZSSKT2HKnw
p7GOF/RfZUFQpbWoVwv9o2Cz2ama+AzsJqfUOIhhvXiIazq4n/Uu3uLfFgGNg4PdenKXMwEnokb5
LYYyRi8UpgEzdUcnLTSi3bHFhqPBj8+tJY+X68lJ9K2WUxHESIMCjvo2GXUietCIgfAQSPAvqHDN
6DAt/4M7JVgKyLd+8VYQgo9WYqtocvawmFyHPqq1O4LPKgu/tcR+Fop+RxPyS/LuNSzyhnviX2gZ
30H6oAbqfBrHoVRbIXVNOgRZ7FaTyCoApkHAWj63Eaofz6jigDfLxvaNyg9cM94CXYRbMKhZe6yR
wFloTrNGdlahuoSUtfBWxa9bXBFve0uyIsW1S0f25ByobXvjHwPQiCaG//+BXKzHkohLem7nusBB
1PezEpHZYEKen4woOee2yYRWdiPpHsAVhgIdVhEt0uCCzi6xnvmEKKiISIxGns8K7oR047kVniL4
sTt/588dyqx1Tbf1C9G5dmKfDb40Z9pzlIPPwnQAjHvCl7ymOkY0/zF91BovV8eS3K72XSfq07Nm
CfoF28q0RPoFM+XDTwvhmXug5F/H3uiJG0LZ+6Mw2goFJHnSzhbZG+eHy3/S7ZWVoZPXl5k1v7U+
bZDXXLfafNuMIPofka+ozkjwXaaiB+uwOwfp4bmbS5tZBlZe2X/nCbsR6PEbo1b8+uzBz9PXz5AY
S0trxfvazAzEUYnkJ+7LpjbrUqKjniKmlFF52oH+B8yytxhN1dRe2I42qC2o/toqOP2SMfxfvrrc
dfc2fqB10UsqPoSNh/lwOEN9lkCbcnltgeNJv6i29AXTHA4WGgybXl8SuoGrCOsF+Z3PpRf0GxgA
nZih6ZVOuhohxW0WEoDZV3qW5/qjNHelDaJRBUDhLyJIvuCyzlJo380MrC4GrOSOY9pBD659suHx
FoXpz/gt9Vw9C76UdZIlLbG76ZSo1SX0JpPeGMlToOYxMakcy04yzT3k6FS4/dymSHD3J2eU3yvq
tbgghrG58I2FtBFDX+e/WSYTpsTPT8vE2CcHjTRQtSENms1zAQf2latsdOhyfCv+hEB4napGBopj
T1U46dhCinS8GkHbUZIjhdy4c4PECjZQoN4ayHqO4TIIPIpE9fnmWJvjP7ZcFyIRerQ1mKWHjYp7
/6HGTN8r1gSil0/9qxvIXPjMIsvJsjAHMiWzpCLV3Vyr8azJbvX2DU/qQbjbHHDJm9RPZLRSkP68
q3qWYoV0EfhTupikQMQ5wMskOuswTNnH2N9+LhvDxhMsms1JI47cttqpSEfX4sVaZqnTV/e9nwHt
yRHLy32tPt55RBsKw0nRk7+8NVx19LGP+3Zi6xRZqVZH0XnkFkYBxRncd7EVxKG3COAevNtEyHhg
msuSju8Cya+NAB84uM5wCnm+xOdhlDFiStRU43eVDK0SAtRpXx1wjH6NjTJ0nHDJTGZIYGFICoI1
DB4O8X5qddgGy1m1OlvxdbDUo14xcniMN94FmFX3yNlsqSa4cW3jELj5j6Rt6y5QFFFlG1XWOH0n
xU5VrsZpSB9oCQOHOkZpFFvbLCnjHvypfLPlEPSaVKsi7OxvLjJPbPi92+IQzMmWfUuFxjMi4rWx
10IGnSKcE/sKerSgYOFreAzPhUaZ1YyfgFe/mjmxNt/sP14RlZo+Emz7CxJTVq+CeptVDZqBdz+w
gZtxXIPugngFm39itEun0xExmqG3R9anlcqojnVI9n/YaAWY3TX78AqUZ80PZTJDK5gOIfK/BlIc
+IbuCx4nJOElbn62F1VhhXgPlYpBqbutLE0u/0UAXatKYz8edt5TsJAIduy7ECTr9HJwZiV5cGyS
mwOUwioqMarh1hpuDON7MD4cJoPswbBwDwppgI9f3Jkh8vqOITgpRA/BgpH3NSg5+lcpvgu/KQCR
+2WycdSXX300qFtTzWaUCRFmSxe2I4ARgrggJVbpZb8vAPvjRI3csTrTFRRGFoH/SsICO8nyR1rL
XQD4sZYBGTnmyMn+sGRPO24xiN4EUQ1gdP1tQJHcd+azySvkr4kkAKUZjSEWsvOqetpaxO7zqTna
Zg8B/V3OZDKHugnvPXeGKqgwboomVK7VPfgBQ51z/rtktu0Jy5MkgKT2pRBbosfWOWYRlK+TUXfq
mpShKBHpnybbpX92BR5P+7RWzpIowXrb0Of95Bq+6s60jL8+s9bAYHVoyK3MRmmUXa1+7FndfM1H
rJ854oftK/wRNCHFbanRzH7W4BtTrErG8IlhIwY4DvJa10XuWfoxrZdoLGzTOnUlqYP7Tpz7rHVE
ho7oroa8rgZQE6S0w65wsmlANlZKmhj7gRQgeSq+1O4BeMiu3OwUinKf+YK31vcMXLDz55BNF2Gp
6np+ims0fIUaWArLPCgT1Xojj0U94hio+3LnLo3Zr3HjzkhVdRuRvrXc+Y9JMdBVn/wKsJZDJ6JR
uk2TDZLYPGu8ESj8ftYDxHYzHAozyHJbJzIF47tKAqZ89K7uqRiqBSukVtKGM5djr1smmR1yjykL
Y0E4bu+OX2Dcu44I3XwRCc5X1YVzviojlRNS2qYlKqP2tL6OkA4qkQBF1jMvtwQc/8nudgmwQem+
ZCJmPm+uB+k+gTRGHTMEOaojBdx2Yjk55P5kbZwSYvWTZZSiME2HIKdnD6jF/jbIDMGTUSTUFyKI
/f+SGsIBZboM/vVlyXLkjgde3NPuXh5j1MKlvho3oWdqurt1liatD9yYAXB23fn6mduaKz5+YsGY
QI5mkqJpQI5Bl2b5MEcVh9npvdUjUruccj/l6vNK6pNVaqn3F03OqsErAAy1Hm9zY1aYekZQO/0U
KZ+YLqJ0bcbi0bAK36XUmhqGF9I24N5bSqCV88BJQtGN/hCSCTFR1/rFuJ8e0l77gxGDqio7A1CI
SAQPKaHY+3uCUgAgU0C0mKS/am516vRS/ouasSdahKcu8fTi4OrfMp/h9awiwcoC2xsPwqYgu8iv
zd3h/T6KAY+CWBbHRDS25bGPWuaZ5zmgSg+ludnwXwOP9Rr/gpzKQaAotN2l2mxk7UWdZDBlkfp4
MAj7h+Q/vYj5LF+LPykpUiMBfl3jkwbXuylcSzGESMUORJ12dzWC2o4DOdGJlRcp3IkjuWNaCkAD
pMi+U3XQiZbBZu75DIzjrxbtYTUIzv0henS5PG4YGwg4cx8fqjDOtdOWnYlAawvAKqyc2TZ606kP
XacyDmRSqYZM45tb2nLswzQ6HKubM8rxH3FpxLeR1Ky4L2fIOsuz/TfNzUlL/GT2iajtgmFXGc5P
/i1BEZERkn+5z50+oL66PmeY845Kdr4LvnB/W5Ozk8m8/jvbM15z9eniqzGtT6wfPhvhpqovrS2c
jczGk8vi3+8+O+cGn0aDysgTsW+t9V0OPE0D7pCbAkpE0zHLFviymY2Y2os71vkVEGPT4RHwk+fr
Gk7dljlFFEitNWl4+oWKtE5h7/8wp9FsDQXKghOs4LriFKx8Uz+c6U82B9CSU7HvqrZcor/n8rtr
9oulTdZ24kNQZdm9wAb04tjOZuwrXpJT7t/kxpBipVh5DkCwRsTf/EpJdG01dv/U5Wsm/aZusedB
0Ot9ewLLWtISSIx6uuThsVWyyFu9rbZaAhXNI940B1WvCk4B7gLJNhDmzEatP9yERuUczR6x1pdk
l2lGsS0K3lFzqDPENbkAUocJQs0KbXv/H+hNS6EuGj+lDMEfQCu4wbLhNN4t+Wtk7+DDhzD7BKD/
rGraN6Aygfduo5LCAC9O/elOrU6EXVuB+Iyzuy4QKtj43vovVUvUFq4g4EAPLzbmOHprKUUH+LzM
jrlsNc+FxAO6E5PAdm31LAipcNTOyyGDIesTxkwGVTA/UX+CNDGjAAcdRS+62d9ymUllE1PnQtPs
w2YFq5q7NdtCs+tYPEx6djWu5o1XiAjpAjLlrrkdvvQDTZIewogNKLhtc/7mIgCdN0lmB+2lnuVT
qLs6zAZfTVmpiMDSHe1SrPNiApCEbYkmXOG6ryaqGU8Jpg89n28A10kvvPGAZdPNkSfgReb9RquE
dHjf0tCEKuHoX2MXj1klEd0Gvb/eHOHIbxCR3JdZem5qPo4KI7tWTOFREtsg9lE0APnot4qqu9bJ
PElAIykPC1MVt3vWACa8cVM+k8/PmgU08mmET8C4/3CDnS1XMdroipWwOQ+LZYeUPVn+oWVvFd/g
6X/ZWkBloWqW1f/l8WRXeheS2QdxH/iOxPs8NXfJAJjfqlzd5/75WvRPD8ET9fs901FvX1qJs7lv
hnaHf93EB+ST8LAMobqLQG2jMRrrr8mUmCkb0ZIFT+ekjroGRX6gDRPlRyFF8Bl2H79DoRxuswGc
stEZ7dNEOVjsJVYyaoVEnH33qAZLJnRYoOVfRemqP50i/P25x0uYd2tiiMB+xC6ONj2dyy3IptXC
2pn8V5z+NGDS2JCdHgwwnJxFYE9b1edGzGYSoNFdSBxVfNOFBM2gTw9Gp+mipMNez4upoWknA7Bp
q15nS65FL96FSRQ+4TTbG/L6Ys1xFRETSKQtEEADVWVqQHY4A38xz68J9eB5jnci0wy11Y8gbdtU
9vz5ctaFEU+Lua4MI6FUsqT2K+ZmfWTwheo+Adi7BiOF9xJaQtqSw0q7G7NzV83fO37uAKQevXwh
W6sdxysdKR/i75WYa0dKw0weqB8GqyayhvhODz6OaERwsGB+jWX0YoxDFqLE6ven6xMdY8H9B2Zm
XwgvXSjKiEsKTpwnEDACZyi+B7aNi7makONWRYQGyK+4DCnlqNzLK/IZ/IOszdyckDk7aleHFCXo
gtnEHuPy/4Kg6oPVl9YXz3ywGlOk5kXrtzqSgRz8n1/6c79Rn2pvEfYK7QzeQJisBdCRMBG46/J7
9m5tebsMbm6WZ+L1n3P2qPb7f7xuDbjXQEbjOp5k2IHiNOESO/hRiZe2SnYwYod7MubbF2IP5yEV
QMhy+PrWXgRIZF7JqLNhQvwnh5sWRpO0wKHNivQf8LHWOBCLRWhoarn/Kr7N5GpddRANoHz3lbnO
rLsaGdOdM/fD24+8qw3K4gm40OgvjGpbrGpXY1OrhQg4x0wD7W8B2PN53cy7acQNjZ6aM4G0CS7x
DKbP1n+Azt0KvclzK1+ZUnUPn2OI5HN57r7hOCLaYe1liUueHXOiM+Hfim/Ji+cqcPjepmbSyhvq
pAhk6NT2jLUNB7C98SVEgWkulX54n7tXwPtsR6584cnqHpZzwVsLuj8SM+KvIfp5MsipoNDXHAIY
aT/caeK7cC/CX3Ev598uNvfD1Bfdbpaq3FV7rhkxQH0NlSzDOEOfs+KZR3O3XlqIcDohfDS7GCJd
X3/3YvW1c7pxSKooArmN7tcWkAeSxLgfNd9/4/s0N3QZZ+0VzMJfXWC+9YPxL4eReKkPnkYNPS1G
fAz2O6OieSpJyyY8QpF+6EXU68WZbHb7W5M0KX+xVqwcM4Fn0eEALsxu/zZdDqJcplXsiDPPKTbw
gl52XQf/t0bAgS5wg+3n3/WdZ2ZC3LJcCPNi1a8f0HutWJaJBlxbG4JDQk4l+RBscAKkfFiCAlHq
QiRswHcRNJ8uUcMvEpmjV0ufUP2yA8R8CTeN4MQLnhQREcTrBfb4NZLVbRqKcIkZivoj2BNPIHOv
ApCPVLc4h09GWD7BadpwV4NWtHPe9zQeJA+3Yh8kbGBEn4hbsd4LiRlx99e5ywQsFU40jYd9KO0M
iBoD4M6Ax6c3oPsP/J58UfCQLSqJs8k97h4H6O0du9erGxyfqP9Wgd67omHVkf7yG9W0f2zEv7Fg
BTCFQheIuicsgXjwILahcm01yngIGfOB4OXn02x9p9f2FMrQZnFONTlOxhTvA1v21UvJFpAm/D6q
MvdIWM1xA9DVOB6UvJW7xyUoIdfeF8ir46BFYKyrXDEBppCUETqMaiK7cV6Z/ZEJP4FeJqp5+Ncs
GSscO7picDXTVm6vCh+KSr6JzYXKCXAFzYJ5KtqXw6vAqa2tgTNj/jUYqyPYHuwbdq4NQB4+NBgj
lNAz2/OQ+MoGELRMxswA9rVdriKhANJmnW5GduzXVl/FUS5HgNafO5UxiTIPgP1RwrWY58OCnGER
JnhGn+6e01X69hSjUBTTMtRxAfSdTpy1nCSdPuHSsUNfwdXgU7lQPUvTDNxaVYq1K7gsoPv6ufV8
RhlnU+/IqWzMrs4V5ApZR/wotfndb0mKv8phrKXvoitNPm5Z7/LISXjzYq7Ft+ooHFESqB2tNg1E
lOR1R8LjosggaKab8wL0ljV+qI79xV/K1bwfetrD7ocBDhnKOn9G9B41MWmq2hh47nh5+jtGWVqB
Trt/uy3Oc0+JLiXrs1X6s1yOPQaWtJokTWQayryVotskuHkYZRuQilHSgI5+cOyJvNjRYoIWFuXK
U9a1kXgVplwvtukj3ag/fQgfgpyzDeOgi35Hq3PU46WPXdO8VXCCJNzy0qR3pQF3p8FPLSXX4/7h
1TUV8f3UuMpGPLSOOSwsQ+NjunIsflntwP2XcwJ5VyNm7/0r6XW9/NZU4xGgUQt/BwpqrNuAQdrx
2BVRz322RQ3zXkbT9YNZ7k5ssVgNdaED/UbMGXhfn4wOx40bW4KXpSYm43o7DNI7RQ1DYNDa8xt9
hwgt0pe73Wr+1OKzDB8+5mK+dzNwnBIm2H6hHv4VTtrsjP1gQHm/2fcL/wUnSOontTA61mZhdfOj
eM6xBXSTfYcAF7VsJtWKgytACA08VfAlRkO8iRCjFGcXuDS4uFNnECWTwB9fo2duPrXslKELMLro
kUmUJWqjD6J/9djuEDlv3VlH5cZfpNI+Us/AYRLKPsRS3jTqFColJoSMBT3d/HfbVABxaGkec6Cr
QtCtghHOfaFurLR/J+OQvUU3gjrw9E79ybqyuLu1EY4PTUmctOV4WpugAhv3bv3VSoNvbrxz8PUF
asTUIV4HoS252G1viVMD4bo46l4UYi4ni5q1usQBEPADUQ+gthMjaAkcNl4f8rMakpqYwKF1cB0z
ST0zAeWZN2fV1XF17hWoAJlWQc1NQhqr7eTnRbapPFdWY5JVT4VTYDcZPOPbzJjIfZ8AJZOZnvxZ
wHlayzvnZhU9IQ2hVtHG5cr+FgZ91ijh2WMgqbKox/JYApr0IiC3XEz389xbYRcYa1njl1AYO6ws
T5eiCBo/8JgpIzYA4PNFoWYEpbY4srkEBF6KQ+CR1Ff2grZ5pb4SZ+VXtLeSytKPf1Fhn7reM2QA
jg67GSamjcWgOPMwMZCadxl9eyTyCp9Yq/5mv58/MVMX/zFjJi6S/528HRwUZ8hKOoEqMQ+YbTUK
HBQtq5zq6iPk4VhmcGLYmkQJlzeUpW4UToMLY5cPOvWiy1M66DAqmO8M8e9lrVNO2+QfmQ7Qqjwq
jPAFAEl/48a7FmdbNl2IX9gNir0crmlqpVK1ANrvn4O3U6ME6cHLdCk0soqgigPC5hrutSHlwCiX
GUokAETCq5ApTtRIPaudcpDiALeEA1SFzE4lpFk4etrsmuoj+Nafhfq+w7nv04o8qyqlL3w8s/9d
uTu13sSa1RK5Lf3L8ds/l8kChiaiVUn7/qC7Kn+kPYIUvzRDEKDsc/ldjR+JDcNXTjUaBWyeMxlJ
deaMO5RnSqvDcKBZAO3lHCUAu7G/vK2tJy2MEUrF3RwxvpJdvZETp4slfpzZjGhhBS86OdWPUBPH
XyHzmTzIXrFMaC/QaTPft4S7B31IHIVzA/A+X/ppNR564kYnvHKUP1HFXhaMTCPGbUuxJgqY2VjK
pWllCVPjDt34uiKyn+9wg3Pki4n9mzLBqSPWXoSWqoS3Z5v20n2fWiCcTo0h4RKs0hX5e+OeL+80
65R/Nbnlkw03xvGLmm43/+QkjqUKA/Mu8JPwCxQRWDyBhQwEarf8OLF5/cj/KdSnr4eq/3JH/teJ
Fxe1pKwkvoJ31prhaGh4wTW4LiFh1NsRZ3C4sfFTFK/91sUxH0xV4wyNFckAI+w0I3c051mzvGPu
RaBYZAQoM/UKw1oZkpPDzGOvsYXuNzPmVheT9Ck69TGlUId7cLqQ9mNtuQqwqDYOVVDH/ziwlTp4
b09Xfy58TQb+m4y7mWylWaDsFm42wWKAFaBMXsvLyraIfJ0scerVVtdLnYHxzv/BFfI/ouS8FuJt
wGuKjsEbdsvnbDfCvANJWPcVjlHdMMqc5J4L8dq1yrRQ0m91nH7kx/4BYkBRnhMTT0pgKhFl9wRM
/OQvjlZyBHERT9G/g7OGRYKJzeSkQshJUKmfYd6Th79opMgKZKoxDhis8IiHrtOWP+sFJ3vIc4F7
WF0A4NOg+7NzE5uxAVW0hQTBMljm9pScjNusEGzdQjWk71b0kPT7k+4h2IFCT2pL8fvMtUQ64Zjp
4X0Bf2VxB5qsY1f5i+eRS5fobddiJS6vVcQ5pHKRgun1ef85iyMJdiJD25tTDjQvfpEHoScvwnaC
LBdam6EjICKAlHjl5u7YhbjjmirqnACB5DxSAA2BTUSHsnMC2kuga71t/aG4NlC3Hx+xs8259cpK
BJ5qlxdGYwvPaGhDuGLqhOcMcrhLJCS8/d1qn99GjtUmJLZpSbEt4q/tUEupj4Gimf9lpzv5S/sj
GmQ64QLo0QwvwFH1PMfJP5qYNgXWg1m2RZP87a2efl3TVtCAX6wsv215u1mIXylRxDGS0V+A7SQR
OD/K29jRO9OyWWIw0RMtDYYJvYFPUJz74JJ93Ap5z/MuQgzTqfYAMQd/WVaxBlomCoYJNC23gy8L
zybls/JIHIOt0bR1TFtHEdVqYesNPNY+hVMu1XK6qyal2hLozagPRZ91Axf7hgsbov2E07MEomfm
Ez1/IyvV8kGW0e0qCgG9KRSpdFDYkS+SxfbQL9sFbDtNTBz+NRld1QfOLxR0XNPWxLMxwCL0gwOu
Nye38XeD949Gxzx85HjhyImvykeDlSG3aj+/izT0rTwetBchxnpVVcFMW2n+iYm2elKtsxzOCREY
P04f43e9zQiuYyDlo8xcYLmRicZgIde8Z1XWl4Be8fzwjUFRecRLdH6ydN5MXk8/Q63d3W8vlIAq
O9tzQqHNDVJl3FaxaiE4E8p/4TdZVQMKCQObKMPEC0KhXiPTlNHp39RuOqp2E0Vx3QGSEcmRQBlG
SfjWS36+XxrE/c0Q5xduusfNYwfj16VWfA/OOfpq/Wp8U7EHCIVoQzumMwRr18OIHnbb46AkVm9z
Hp+NGDZL6WtdgVN5gfKxqyER0C8h7t6t6o4ThXxzU62a5rdZSkuBmvA6lP954TfbwocgswmnJjj0
MLoCMGibzQralg9ZpsN3WWnh3wtfsUjLfFkJfAqsj7G9ffo0bgTbFCZtyJj6pCA7WhAAyAKBbVpP
5oZ/tPJpSoG94iUdYmS5dHt4SfDtjQy/nE5XijdeZGN39i5H5z3kP3xDQVCUCyArXg9IE8UXOhn7
tpSh4+Ptnue6UExnbGVyW4B9HARRP5lNb92EtFdQwrLeDDMN/FQka9dbbOofiaeQ1s56QtIaKuoX
BLBPbJEZhPKmV9xV53gD97B8lfBr2rJRDD+hqJmkZ3CEohzOhPiyg1ZNDftTCdlp/pVbz+o6cTmT
fUf4ZSnIRVb3dXJCYKxPhtNTftkGkN6L7yfVJAo0Or/AKWMwmP3B2PSmAaAT7JmnEgUx2ViQPVBI
rsul34UGGrb8znPsDp16+epexizoP9sI62NTcdHwQ66ofrMRdk7HevK/YgsU1dpF4IZ+EK95GQ+h
Icra2ZIDmbri9LIL3HszJ02FsgjPWnZc2FKgdqabDNy4hSlTMjnwAAAnpf+zLqc/STXZNBaKxk41
eZd6vUBHHlv1xDkBUvq31PhtKyaLaNpGFhflupRKFjgsrfOHSzhIgji7n+6Z1sDXjysZdfIFRAe7
bP1IUNd2tMbbQxq5Cefos+/rZaWvTbEqnIGb0dygqUNbNRVfQbBv52maZaW+e/sUy0UYA7Yuagoz
WNzdNVXrq36GHObDRbkNLIZiSiU6mhTFXb/mhumsTtcDJEMRrMZj2dUpH6YRcDtvh7MJ/j/whTms
YwUUn0Uu6qadn/VrW+CFf1IGA7ympiYozN1Aa4zcLGk1dlQGTUMcbHnvRIoBnbeHAqZvK2VNq998
axxI2IVK5Pzo9xAkGy9oqg9oQLrKCCGJl9afgGAic/lYGE/m2Ceh4e5ipyX8MzMT6kVwJ7ISOX3N
qW6b7l9G97sf27SoYs3Tj2ZyjSudT/+ATymrAhLqO2dlbNFCXq6himOS80rAvGTamBHB6OEZbZTO
uPOuaQYzYsZ55JziUDK4Pq0RtAD7A2gdTAgrPhAGPP4bdogjlvetUVyaiP7fELH4CpawMXqV9PHg
bYvT6WHk2tKugyNu1gjWnzBa5elpQG6Bi5LdKE+uViF5myH6qHknTJT7S3TpTB/FyNu/jksU+/xf
MbVGdJwNTdgi5Bb+4i4dXRPtnGInnJ7piv1fwx+LRTRgUBD5+A1BnC6/ax+3q1QE3LZ3YsjgWBap
bV3iSmarIPt7xCboHce2kSQdZRytaXXKE22LrsL0Vt3KLAmViAO73SbfOLe5D06lhAFPNz/A09tw
vPdLTNHS9g7s938I4cvYIWvAlSg/8XZnpBnPYyL5zmXwkvFLWpT8zSVbQ0JN9FOAON/xeaUFTbrr
b+F19o/SVumkKJshxoV8mlBUDFr6arSEnhiEerrPgnJM6p6vwOuoeatv9jTfYL2+ehFtB1QOzhCq
eNOOGZSQlNlOOwzCkB6GTbVrlMJL0X+4FsCf/PbSW/Q9fJHIRBMeAG+kyGxpXqT7Rkc8Pt0Jk4ZG
5we20psgo0eqc27LVE75j6pdQUMwbxZaWqt9SPTFmBc3PjUTiq6slSUH4sZ8r91k0DKrLCWzE+Vi
nU9Eq0WgWH6ZkKbvA6Ydez7CfNmVJ2XzmeG29vM+0Libh9Lpq88Y4o5FFYOeayp0CBhYcDTw57oE
0vaNd4hDj4aJaDoF70yX3HZpRb5t2rY7kSeMMJlhokpxkQsSDPoHVxFajl8QPeE9r46sriqGigLR
1+5vPoBvEnok59gYvwLQkOFgDcweZdYB+4WUshG3K5Op6ah5rkdZCnSa2Ne/G1qRIdi001ed7/Ih
wU9segBpEClJhkjJUaOtRKOQvAYzNjRg9ApiA+AnctmAC+BjL8cH6gy9Th/chlWonpZ2lo4vVEsI
LVCBNHCSc+bvtmOZjQcqmzI9QyjhPAtoMeSx+K17v/QWNTqGyDRyY+J5+RRwThij8ys+Vd7Ii0+h
uvBVNl5zeh1ELEP7JXt5JJn9E0tWbyBC3wCnpYDTls0HB33EIdm2g2QJIqyNv2CFtsHbpi+JP23j
EDYZNzhnxstz74yRxq2r2dpmJhbxYcBh0z1eCJwQ8zCo1PIVTkPt7+ADf11598urZAtdWpPMhVzl
2OJ4AiMXMHkFhHvHsyAwSNMeUBG9XPoGPuELtJtQ1QmE7lJeb7dLWQRIgnEaoTBESldJVdDZMrg7
HN3OmigPr9/1CRcPxtKYVl8eOd4Mzpzm0pMOsINanLpUGEuOYDiNV8X59M9klWxWX3Zl15piDaxp
9d43cjCwMTDF9LQSNch8zylwhjfgGIGuLYXABxuP6AAYI3M2zaIl9HvYFFRP85bEyJheVyYfShJA
MVTjYmI3rNJDdJdYBzKRb1+WeM7nXKe6K9AbFHqCeWuzMBah2vpgaWuik2Gqczt2A0vAJT8uY8Ii
p9pdOaVd2jahYGZGBUWOzPUncq8ykYqo4FTCl9nwrY+ZwoK1fgJbr7frg9BgyXfY9cMYYT+ZSl+W
8rA6i48j5OqGCkUXN6nE8X8LTF7PhjiOO43eYgOUx0oQykyHbKfsN2etfNn+s81GQs3ItayRCh0m
hnycW1NpAfOE2KltYyHjpW5WNZd7e8Y0OauQGYW0cYCb1SPWwOVPHrbPhC2D72asC9TjVjUyAz26
Hx6Fx4Ou0Rp7wQQZ3c44FFXARACa7qC0GOHUrcAhfK9WbtRzVGbpbkuU2txQYmvSVn6LL+JpLM+Y
SUheJNVFgUVzKi78ljyTJqMM6IBo0qgXYT2tAaKaVP5xKwicb2N1fxf0qMTrQB18fTzd2i/hAezC
nJBxvqtJ873vn4llHB/6KPWT7Mh5i5XtsfVmd0y2vDP5opWkdg8NeD4H/Vk9jSXdn8ZEAzfDMr5K
XFgDbJh5t1b05azLmCFRq2noH0W6PjGbs3TFEuIImhmn1TCMmel0hsUMt6UlmI9X2kiXyol14Y/O
CO1yPlRXfmENC7yollb8q7qyDaWZ2r2Ia03MikU3l+k2r/madlKqscw5ecZELb+6X+FBfcM6ZK4V
53IYAPS7apiZde0hOIK3+wc9oO7IVcKASir6hXOD3N/fUl7NLDykO/fZCt3VgxlnJNLszLwW4Oxp
yn6ft65/WjT0xF0Uo461bfG4147s+iy3nOy79Tt/gSmGmRRKb3aoq8Q0tveuU3aCjKyp2vlvPAHp
jy7rR8x1n39Uhzn8WhyYFUqsqliuxMffgYAEfu0hehO4jPGF0UAanmAHmTgE3ZRUr9S3eYkQBEmV
wRqbZCp27/ZV6yQ+rcEsKlanyEuS+lGAl45skvRcJnoGG65HMVreQOhc7eDGLEQkf6SBTIfFTmyt
UwfD9EYzcAMDSdLkAgL19O/zvqRRHYqrqe8R8cQGUz/I+GfxWPTs9mbJ5P6hy+s4VGnYm1ogPTwH
cIJd/gxXoyB2sjPg659ssFvnIYMBQs+7UK1CpBdXBf9CWW5pGLogklRVWbICcq7lmxsvFeNQisTJ
5uZIdLdaTaABah7XgdVe/DMrI2ADu0o2J9yMIF3o+cHd58xX1UMtWi1MDUAAmzF8cq8YiUOT4Zor
Coqkvtenvhddono7158OPzv0g1Mm6aQL+OA/HmSDg3wHWtyuIpl6auCipMfhDonB/oloZt/P8Sw0
8L9TfTEW4tiwHkOiYTxhQi7XzLW4XzYQ+aZNKtOOLf4VsE8sq5uxwil4kF2XWWcU2aPTfwB97ht4
49ej1K7QoEIR62muOAAtZgiYCfz4czpi2tlmBXMuY+TsK8QRRxm5SR6rMr4bsO47gPbK6nS5wqHx
zRxBr1wR+6BOMR16ndXoVUJwmISpZBOo+Qpp9HQjqbbKvysKbBQxu/0eac3Oj7nAfMFHgvf3sxHo
RvDeCaHXSXftYqyDSHll5W7lMarizddlQ5l+0Q0e7W+YG2YajgJPLyvfkFBEPOCH8SqJMvBGgR94
SO+oOct7QKLSTztPdq3b9Hv4m7SeHzJKJ1zqit0jr7x2/+A7ciCEtZm1AV0QGYPlWp4Z0F3T24Ol
1AagSB1LSkeOQ4AcAZNNmdwQA9UJL/4OjAWIEkt8lJS9ykUiuWC+t5Jf9IfYdSWBseqnGDsfosVz
jm4MuYzY69rH9dk15yFsZT/969N8k1LY49qGdwtaUapU2wVa8bbBNx9iK6Q1jlkBEJK/4cRh2t+u
DC3RrSgael5ID8qZxfgLVHaQknB1gk3kt9665irXEkfABjkqwH2x4SxMPkl1DqxyX2RW7f8j7ryS
hyGUWl8p0Q0Tr+neqwS14d+wgZVOkXxn5eSaDNbVAes6iHxXEGhfNMVyE79beKk2DY9YqGaCk7Pq
oIubc4QP+W3f7H/VFoZzDIDbzOiRpX7IX7tsS424SldaMOG6wqsWgZjQk0MzZYQDSDHH7+xEPULV
aSOmWPA5OQFXyNjewP37iXeKZ9LDkvRwtQ/AXjRUp3BV8YWx3S2fY3RjwHWuFsNsk5XKIiXJQTTk
/AYU9POhuKd09bGgg4OKxjrboSygmOVUdug8Lfv2RvJUPgIhsCyTY0MiYqWLCo0SdamKQsloT9Bc
pq11ib8khtn4zb+iaqsGnqq2mHgDVV8m0mssq0TxgjZo++QFrSm1Dn5hRg8iWDLcJZB6pmnUhnu/
0gPee1QGNSVbgeUnaeK57k6oraohjibFOaiQ7ra64GyfwTjfEq7MOcaHw0/RgyFFe+ShbrMO8/Ue
SDqhTPuStTDW/IHReMBUaTDEXY+ANnxAhQnEm1V4TPwaM2vGcWPQDTa8DC4Vm/37gQ2WyG9xFsrg
iqR+tkKJZ93cH23o4bWgzpEmRo+W/MHbhNbj8xbapmZDuKmJfjKFdvDvkphv7LnDW7E/b4Qxoacf
qvJk64e52O8tY8dGkUHoIp5MpwUzZ7p5yHgoIRjhjWntUw4uhn3UXwHB6bcsNiPsP57fwfxqVCh4
2SihnisC0RXN0BmR+J/tiX82Elolqt+/3IONFb0CSf+jOZapoVw7TdHSBKj9RxsbkzzrY6rXGY79
TOGyWvjR0rL8/ie8iMj/ztVk1LNkf86FA2U+Iiu6zWf7lAOoDLWXvlsSlt3vWJeNqwGtA94xa+Jl
ua9Ng21NN/7JHX2LIjrucCLX4Ko5KNJ01PoqRiXrpR8pOJhTAZ5Ey6lIdCpMgYbKkZbLUx7rnuev
7RBtHeq31MhBap548NmDKQaYzWtyUsIq8FWTBSAkA4UowgDeHxewvr5j2r7UDg4bz3Q06SzzLEST
AckG0wXWWZe0ZixinQA1O8U0xyBrmyWzqMJZjx56F1+cQThQMlVI0n9YgvkYZcpUUBkC0g65HXFj
04QzMxxOJbJ6mbG7LVRWcULINt9a8Iq/bQ/rR1Dpw/2q9K0Pv78kgHhMBjT5vbRYk+U9YVPeslv6
bRkcINWVDAIGb+x7kBGpVR7cJGvH+Od9q67fxFW/Ao+7YyNB5yIwTxZfLeYUR/eMPTyw9fp0fUFn
E4HrlaYsGyXPk6YRdgb6W58X5L1tjRr7DDh9E5T4xogzaRFemawPj/s0Zk6QJT0h/6LBtUvu2OzG
9vfR36zEcmwE52xO6Ruld1K2ye9IyOeyItfgIuIuNe1tVXjSARiDNtOORQA62KgprVC9lvHaEKY8
f8K2jkQZKCfZr9UNgGoEVLd1fcrPZZcnPq13GwlmuxwFYY13BkSxqMuGA0sbjbKynEC01oYKm4Z5
BksKfvXSi6qRH7H90AJrQgmRSqN56U6NEGldFwTUXiI3KFDP2LDXkd37ArfWEgT7yo9pApPTVUnw
CLkTMAiPCDpB3xxlTQgKv9YqHegsU0ZwEpfrM/XlzRWgZlyoy0EJd/0sK4FvnaxZ3gQnJhkl3Wg+
FYCC+ouIf3yoVmLj1QgZX+BXlwtz19Ir80b5rsVImn5X67L0l4REd1FiGfiuiRKKe6XVYQXt+nqo
9qDQ7MnlCbzKKAEskwh/3ecWL5nNFe0EVMXimlDDMaJ6M2yVmYKhoQOkS4EoBNaMXR9vOxDqpmg7
fVpMAoMUJdYwDyrrJODUFkdH31U0bU445zZ+EM6f/HvuCUrBKgfkuf0V9n0yQDzPxA444PuYogMV
40ZcVrymGq5UT2HOmZJmYLvRmSmgAbgVShiygRQp+KRUOkTV/kHOgFFM6XnexAjdtsSf24SojcBS
rsDA6g7+qZTdUJnidlUwzoouZUrD5m4jwdE8GiIm/vDmXSi7NWnbBrmyP0ON1lQi8PslaDH0FGfB
xHSXMu3AVN7YkKq3hajAxGmUUCODd13M1yV7QUWr8pHS+Xt2yOH5nC0cA4NqauJ09kv9rCcxXchP
XHBsqaN5OnCLnT0l6DICrcxmv6VknnRTTDgBvdjvbqPo/+/uiHB4RUzZCquJz9tpXc0Na7Dxt18P
ATNA2MrCuJSYNMdooR8j6DN0zB7NjVpvYQCvitpphM7fA+9VYWCSQVn1w5zJv8GSTHk/WmG07Gz8
vGZ2F+mgpl7MrJKI/k9Yu9z/aRKhBBUras9kX0L222ikGJ/nx3fJ9wtGvxKajM94hdyNkmeHB1cE
y09dDS+/IQRXIreAgLC8quGXlPkORRXBARlDW53UK1XcRF8rT/oXR9463sH3L/ox3L2AhYSpC8nF
lXOU8yj7sIbkrg9ZQoQLXFt0AoDf1iPQ7I1TspKMzQYqaw8ctdJhPaDf4WYDvz65hlG1S0UvctLA
yr5EoLSxyivibkiYYKtfysN+3Fs2H8vIr8kGoLqv5WqkmwD22ohAcqPWWWdZMkwN49wODi9wTSl5
hURk8frn4nrBTZsttkdGkKGvYhndfdrX2qsabCXH0cMz3E1rReLLMevbzxroMoSQwaPU7IPboa6I
bPAkkiywGfrpiL0onZAZgAqOOcLKgn+m4y6GTgXo5aaYyrnlWwE3CNE2IF6esQDl6Hu3zI+bGelU
3W3jnVch7RzzQ0LKNLf+AhSV6GUxHPKjJGbm8qurO1pSuyFDd4GZBUj84VRbZ5UobpnjwAEp69f7
XhoGqky+TjWTWU36giR+l0t8rTuS1HWvQGCHBPtsNGbhYlSIxE/nTTnq9FrgLISTXH6wtk3loVsM
bdUG9OSMJzQrI+ldTI01WeAqiSA2vSPTYLm2b09n9agwiJMNaxWrh6He8yNYl8QrojXFm/F9Dx1a
a6QbSUT7OldCjerXDjUdFXfoswjuUT7Xjpbj8FZ6nQiqiPs5fOlqXBgfVMGI4qK4gIWx8mcu2p6X
0928r8wHq0lMCwecKhhuSapWUTB627KrZDddsZAZ6n89oQi8g4J3ePiRUetpUrXaulTFLylJWulk
bAOtgkvWMZNl6GRcOj5HbCgsqJIh6hdot6T2j0JWiZWzTcO5Gs9WKYaXQ8+FwzeY3qrvM7d/mKyk
n9jBDgrju/7/rHVQ1Vkja5yeoTV//yAI/wmVJDZr+v38jFi20yO4XZUFsmIedi+n5Y4kfXGl3qzG
t7CjVMbYnKTaR5jgMMoyD9IkXHIKg7qZGFpxG+xzGEiLLVYyj1KeI63XrHcrz5WvVMfclXUTlC+v
kXcxLTsUnfHVuZLA7Mdt8u/DlyhuMaBc/5j40PTT6IgxGch5mXBfKTeQ3Qf83XJZaBEj7shwKcny
wqoikBvdk1Xoc11R3TLb8YnI3AJ49lWL8RkWFncA/hebfTI2ypotiv6pUvvIyL0nRDrcPTTRiM0P
ZBQbaqIqyQTq96G5JZzWmPyg8q58tLdNuA1ZRcTBxaxVwgwzuGSofVSx7VxmJSLaXF6MPoQ6DdlV
GdALn3ZlYb3/dl/AWrDsM3PJCA4rf95t34sk3XF+kKTmB6a/9qlXqlRbcB+lze+/Nz9PlS/WQqBn
2r8tpRQ+87Td2l3yNQPw10uOWrmsshTd7a/svSgN2RSTDeqsqKnSrlI+98FbJCZCdjS92A8Mqdsb
+RYG/ZriZSAq23qr0NikmL564P+5R6ogsB3QNl0W3o4+FGF3c5vx8ETTvuh2C6gzRSGMJaEcuVMX
nExQkQafryBATn7y8SDyGv3qzkGvJwOar8GC2n/XCHwGPdsrWqEquS2x9o+mwZDtAJvJNt0L5TM0
Z6ESiYPFWIRd7VmMGeb5Gu4bNxAZPKNgGS9mM13oQBnpL8Bf8PuVMb9ymxFSZ2CH0m4grxCcsahW
ELTSPxUtGK1OgMfmhaxcBC1/beJv7K1g/phclXMmMPcmFA2cL2BGzW9TGB/eln/5/2zvgSirPa20
9lO0vH2p9xfj17ZD0hKlVAxzjZAjRHJCL95lzM1GPr8oSfb2QcP+qcK5QKc23yXDFFRtWB2yOu5s
YLUrp+MCL2obgtyPvAeytSmb53+xvuU+bcNg9ek03Cc9GAtX7TFCc5TXKH+O6gTjgxa4IcwmMT5k
aNlHM6onTIzXtZFewlwHNcU2VmZ8NPpQzQObhcXrcUGAWDlrVH8yUCPNpknXWjNFDLQLiluyvoky
188YdcxDqY8OG/1JX2/JVwNy5dfVe+fqudiW2/PjZtOTEZxQq+TiswKUAPUZSOaZjqz77eln8xqF
InWMA8RUQDltTr2iLhzcejmx5cfuSv0sPUMppCfvTZ/6azDCmLs5o2mERtOlC6FbLfdTwLzc1g4x
diOIMH5Yp1U6YFd5mVuca3/lkD5klhkE4FM4FbtqhdPZDrIZU6kiIYFII0v/6xCwTn4BPk9wsdaI
0+ior3q18cl9H9f4Sd7JVPXsya0mUKwNCat2M26ZIXHXKZFoYCSrRPVpjQPLXuc2asyOy1YIgHUF
hU+CB7hUBZHiriDR7RpOm6bZjrXbE8zrNGS2zQ+HcK6i9gp8KU9MJXzB/HVJCjnZcAvkUW9iKEtt
3uWgc7440QD6iOcbPssUg9FICU/O9kY3lkm1S123Si7MF6Jyv9Xqr4NgE0nfn5WC+lg8WMHOazJo
wWmBz6BB2MliJP6x10YaxrvnYhTHbS72LLzjvvJdy6pTDQ28EdBAagOLdtM1HuSDu9m+X0jvImwk
NQtJ184sZZKq5Hf6Y01nnFLYqyV2JkGKkWMKWqFzCx4E2J8/wFPAGBurv8l+EJFjGoZ6JewwWmPI
/p+Stz2ZArT/NyscOLICsIgqOmct0rV1G/nwvHQ94oQk61Itl4QiaZ5+qJ5t39tfUlUnnQTUMnpA
cpBL36gypE7HiQ/blYEgNzVWb9bokvG7J7LYcGk+MLqe2uu0Qd/OSPQOzLUPjV5GKvPCkt8r/+H1
cCWTYLVEfpGYQCfN1R8T/XXYB6U8gr/8YvpT44123unnEKT8M3IuBVtMmiAt5tAUij7Mf859duR0
LiTQbXwT//au19lHmRH3JVJzI1pdle1APBmBsAMdhUcfOFbvdaE6aQgqExsdsq4AEWI1DR9dp6wC
vo2LP0HmzfJyvwug2KjfZTrjIZ7gIIvEfaLR4GjW9IAW4qg8ITlR+IWwVaYJK/q6LEGcgg6VcOKl
G3US/EqaqyW8BiXogS6YXLg/u8HPZUV1MTrmRTJz4V8/aM8Qtlvb+H4GeZYvFvWB0tgrkjLnCXqm
5Gs6rMJL7hBmAA1SHJvzdZHPtF7jC4UlJutswAuEy2YF7ek99rqXZbTT1DVsUaM4zL5mO17V/RkH
LaBlP6I/YgRtxxmUlC7zoIn36i2YtCNjFI0rcmdCiF2WDO+xTM1Uz870DEKRYQ/aqrI98ORZwHSF
6uVGzwhrrwMh29B76o11PkV8053kcBoqiPcORbUDtF3bhp087MnDnrrTRLoeLRbIlgyxycbs6xzB
b8kjGv5PHoeiIWG62W+3mVVFcPff8kJ3rha+uB8SDTpP164+d97VuUx4IL3pBZhFlNFCu62I7VUc
tEWmne4T3d1TT2pUDaXhLHCA9hz9JkeHjrCKZNKduWBubDTVo+5TQO9zIkuIt5SuJCUtyKfg2SIQ
mmU8iebeBgJpwIATWS4fsYkwuEQCmtz+VVpOWgb/UOi8KvUpnZLqvNZ/hkqURZsoct+8PxLnZ4jk
hRjQyVjA1C9gYv4KhMjaeton7xXDV/UY0z2ZD5HXwSDjWri/5pB48bPrZtJqg/qWsvAFqtZP4/30
E7Jj2io0rtLI78icAJfCmaGtIPlH7PL7wqTlcgS1n2xeXzbl8JROIdqmNl2qE2NHoLhJm0ENhC0O
dvp5Vr+teDqQDIhVl3iDxH0h/Kafhbj9XLjsB1SJ5EpdjfTDrNtmzfo5IGlE4e86EMcsS++L5qLO
gEOLupFiQ+sBgWRKErsvqlIV2+tLSAvdcTnVDjAb2QCalRzkug/RM/Ap6Px0YQUecDsh2in+pejf
C9MNbfwjpBju/BEdbL04wddPvwYJiLRF3T3rbSD6k3RQeQ9zjouPr7uTc2og3qBArTlBGsizTtuC
PiOPlC1zMeKNIB99K/TZDOg6FgsFFZeCqOTz8F8H3+PYk85kmr7si54YpWRN3Tgf9X8lYma7jUy4
LrjsCn91OVRTdVe9VfPvpSBzSdaWhftyO9CRVLPdn9PAKRZYVXHRmwmr9uxqhlcAfts5ieWszjYK
r7oQG+HES5xb/ihyF/qwS2fzxecOpPgau4BQyFCJBNC+xU2DNtM7eq14hd6ULMh94Gp3Zp73wC8R
lsxQ6q6q52GiT2dYuzhr8CmqsM0GBZ/Yroj7NskTAPc+7QByi5Qstr+qO7J1EcUa9E7ICDLLZfg9
sYFcO5F9XmCSbiXXc3U67LYaPNMuVY49EdtPtvHIbtMqQ92L7c9UcwqlS9j+aJ2hViUi1x2eXrRf
u4vl8gn2uuLuRtIi/fGBfrxNNNewUs/75H6LvEkojzCjcQ8IvxoHbDf2mqDPMC9r+4o4Se8WojG/
KAY8gd4qPe7u1WrrbW4cQF6IsGubwAWhRNPO503PN/alnjDjmnync3wrNyOUBZ+qKvrLWPCm/3MT
4ZR6J9SyB9FIxozSQIYOt7p5iUcvEflRJtbuIzksMHitOrENWJNj7gMFldy9OUONnKTZJ4BGTnJ/
FaCSZt2AQoQpnVe/fL6qpPMS+3+cBdtZKW2ZuYbdNOPMHNKPs0pKCznErA2+18rq00DOggs1CKpd
EWN8UvWJrdgGion8CuwBh3v52e0tEFGVQmVgNu3ji5PhrHlVLxfTNGZnZTIA2uvt4zraNUoNzSiS
dthwz6AJuW1GImX957k0qXALuxBlXCucdDFX/4LKM8FV1oLaEbeId0QFiI49RGtfqHRk9mBDrwAf
gAWil9kwWN3Lxc/HD5byftC7/lSs8LpNhABwzlOazsJZseTIbGE9cvVEnf5b10EEjR6pN+ZADjIB
r0hnDtIyTwXDISK/G9mHSZq6Yhhlu2XJFcRuV+OGtWOZMQLi18Vrr2LU578w+k8KgZ1LoZgf3KIN
Rvf/BuIcqr7zi3whio6/3C/uEnH8XWsuuZRHLyLujhKcJcrWYDp3ZQNnS/VpWvAsHJZhXepI/dOe
cqKXt3HItnROqsfT4rRk/Cwu8Svf75EQNrX4GbvFkYffmAMv8KANfJPp19YZmilnuyUcNIR61Laa
uzZmkKwxqIaIBs7faJkCRT8MulGgo/YFad3z3OTo+o6yIE2AWTgPaSbMTFKWMv6t5bJw8v9SS6+s
5JEatMHt8XXHdYwzdZaItEApTKBdZ7cXIS8xJ4vtC36hYwyOdURfz4nqeL5q16lyM5IZH8zBuqin
F0dO1zODpGuryocLinRjvIVB5e2UB8eRQM9qYik14cL3Aag2vQkivcW69K2tnmfojbeLLC+RKgT7
DYEc32+DHFu1rU/+p7mojWUf/XuTZVsusACfOFRZiD0SSIJBpofhLCugGvgIwbGAsETkfgF8PlhU
lBNdWST4XCzvSteSgLWvvjli9L/zEqwG+xBLTyuD1ZUoczdCyRL+xOegvA34izBmk9iChWD0Kugh
hyi8tMCr3nhZSbQyM8ZN4x/YyCaOPa5Mbys8jp+zFgO96zvbMJfYvLI/5Ek2BAxybngPoESZM362
PFazw6fV2Vsp/lyajhmmR/1qv/Y2HHJONYkYeRmLY6N2z9wrFSBqven1iJw3nqeKfZQxnquIxkSy
LIBV4APh2MtQotznUGTbrrePpRHY/aFQCBbSvsDnUl04ZrBdPHq5Edneh5CJVauHu+BzkiLSNqAL
9q1DQf9B66bED3tr62OALl67jfUhj5P/xcWAn+3RdAUOhtx+z6S4WiOdTk235Bn58THQC6peHh0x
MdM11u3JWBUatgCjj6gFd3wL+ezIiRyPE1jkEb4y6UI99ltH9c2YVvTDxeCQ+lRydK1Hyh5OYbt5
xfcTM6Z+xIP9HRDskr0nEWFN07vLS1eaT2BT7I9ZtoRg9Ydt6NTtuKkfmAcwXo5SvnC1HjLjycQq
FSpQyWwTbgyvpX72Ni7YQVUCofmeqcUfodXx88nu//v6yH+dEPXZ4grBnUSD/dhens8WjdwM7d9u
OrJWHJIkkRr9Qq7+G8VqJa6fmtQ6kCU1UpGHtcW+GAm1EW6Sj1L4g5De4ypMHMtmqsYV/8AQLk+z
wMJaoytNjbHymLvrc7epCod9hPMEV1Ee+yPSzeQ7J8kJwfB7JzQikdGlxb+uK+yqfDbr9H3XmEtb
EhBnRRLiGKGKsm7Cd4VPezUCwSTu1cP2E1qJDL6Va3r9YMyr3/QY87vhIDo/rFDMYhgGFgrS4zb7
OM7KcoTvO7WnDLHK3kBBsa0ABgiOsPYf+ZZOh5hHl568fn+PkGq2blYdhGXbZo4xDjjwQvETOCYv
o7NVtZrcFin2uk8/bsZw4a1p5KyohTjZ5Wa6RrOmnCM3wnH/qnNNI7r7yKJ5llljl0qu/akJrC3Y
qJdnUa8dsKWN1TR+4IXiAZT18A8xZSj2dMl2j9QvwgwJHzIH8JKXCDPgQmFYjrSQS6TQKDR4dA02
jZEWdAD/GvR8FbrCPExIg0jTbTJBmePFnTSBWN+vt3zQT3/mcG4YGv2UrCDFhu140Npu+4Q3ZE8T
lH086MfQg4SLKpKpL7OVwjr0Vr5vkYa8gQvk/fR7fug+2Eu4BQVrnX5nPPM9SvnJSyD3jdcv97ty
3ZQ6B0UWbGTxhpzPqUro2RW4YdrTwX9rmWShHGolZAR/vvZIuydcXNf5XATOZVIonZGhk1bcrgix
uwXXfCGcuijkWzZqwrNR7388ih2r1cJzzKK/mcyxe1sRYbOzQNmVqcZC2UkI+gAwMz+qVu1VJ9hy
9g9yTQJUSjJyRstEpxg2Qrb3rHHcrkiIKGcbDhuL2mnl4wWpeHL/L8c2H3qX/MQuUkdZ8/pw1h+k
Uz1B4cTXvZ0bPuBI8WPquVSsx3E8L+YQfspzZSimHDCnj01CUw5uFrUS9nyVbBCfva5VRDttazKf
NGQvgc+kM3xtmHVCJqP0UtQsbpFokRWxnKY6ktuAiKi50ZDsyia3fiCAvPYQIQB3qz1pnsySExNw
TmaPHKOsV8qKv02XOFsK5niC9ccXVExCyhGKo9K86chxLSD9MVxQbAkgQgUBN6Lk1BVm1feXJxNX
az79qYhMe5S3qQOFLsBZj6dl5zkdskeujrnzTNgC/YfZDV4K9/E64RTUghSAjNXFuumQoqJWYxHj
YFE+p9rs4KFhlgCdgNxG1roe0VVS79ef9M7hf4Se8QwY2p8TGvv2HEncIhrcUScrgl7ckdAj2LVH
nHTDudKA9DCTNGWDPUP5/GWxnwO5I3F7nAovE0zJjZDEfl9aNmsApNUMY5WNNKn5oSp3ZvrzNbR4
4fSC/HFBvJdOyQXqeJh4B14X/+3uiXkFwhRqYM50+vN+MVRcHb/U+XVmVfm/lU6/P5brutkhtcfj
UHxZTnn5r7l99wxsy2u6tbmcXX9RrSuemMM/mW36CCbTk9o/IUFIj2YvkUE4q03hZfrZxoiiLh1+
lusHX3WUAs90UZnhLOuPvOFb3GyNcQxvg1nqaHxSniHT/kLhK3IgAIw53myFhNP2RZR1BJZkEHRu
h7OthT6GR9+kzDsA/0lUYsM6ZjqCJjOf8KlRR4UciXyGxFYMP/Z3YdsroGJihCYeLywe/fPDjjpN
1EESZPIwPYDP9p95C9xRQixibfnuXuImEQ2R9aBWQUoxUgkb4mDNffoNKMu4V97pGeL4SsAfksjZ
eYhAxnEFUJXLYPcPpyOfbv+8SwA9yqVnj3h4F3ZJwY70TMV+Brn0hVAcGD1gj58H5TiDQa94DE1B
3oXTWu+vAe4HfIJZ471xVbfQGSIZM9esmttPUvJEyCnnb3qnQRxA+AcM4gSLggq7X2XowLQ4+uhJ
gvAfXUWK0MkshD269wHREZg/ON7gp9WcWScPYeoh827OdmFIAzI5W/PmJVWLWIgwKwj+Xa5zhocx
EwCwSMZ0wwIjJTL5ilR/tJJoV/rB+AzGFentGzbhaTE9O7Ha2rFtasraALX/lHhBB4Ry+kMrbkXN
zMniOpzCAWlYy7SeB8rHqqwpnpuBxuR4dLJ3u3FX+xA0XLrxLHfF27lm5KBCDjh5QWzytEv+OTxm
exX3L33tNC8AC18QtmLZi3sy0KDsP7XkXw1t6s05jr/UoxaEgAnQqNedFHYow2oJtisPpTZuIBIF
JALdS2nCkKSRG18VnVwPzKTy35AUHtvPco9Wo3XzJLAtJFdckjm7FEro+H//bTyvGW4l4kTT7+Of
i1qyeK5Vlby54LX45Xk7t4AoSpaZuez8ecMndsNh0VDQ68zI8+I/q/a+NWelKQrp6Ztxju1eRw+/
gXyAHr81vTmP4dg+agtUz0QhVfNR5cIOuScQ8eH2v7Wd57tYzX1j1Pca6R/wW/qec2FWETYcljJ3
G3ESOUj99G3b4YgCH4OwkGi5StaRaYwTA8GKZ7hR++r/wgCXfV5jCSPjs96PQWLQ/SrCoAxX1/bb
ag0DZbHf4HAiQ80h2kOw0ZIChzup4mVhlUKi68oyIsW9ZOpNwbD4EGWFvK1MGJuroBIVdtL2D2e/
vtYomrZNNpVVM3sEJy9lpW1R1UErP2QXWmJpyvMGQVhuXwgES+X6NC7/o84VGCyKhymPlVhDHcc/
5ljz+M8uWva+Y+xRIYq1ON2YunIR0bK9xOsbySHFbax+n2zguC1do1eO47h0tsAFzmZhnXrG31uA
8oJ0XXSQbSEYTk9UNx1oRIV/IQIWQ8OvP449vGZwShZDgVhVdoT5IK3wpmczc6AqGbx18mxXgeWZ
EDwIv8NB/oaHUgpDimx/TT3Ghhc0NN7DPXPaD4dNuvZ4rciT2XpUglHd3SM9apILcOoY1r/YBFIz
7F0O/SMj6YQd1/miuevSiSKHs5qo4dSD1Nek1SZQo+6162IZOZ7Mf0MI/vl9s5/oBk6siqP56nIR
Rcy20wA7BwKhivzOaje9+rSnrpbclTaNImDWXlQROcciXAU416C0RJdHpzXikK+12q/M7OPLHijd
aObwThGpXtA3P1PYn0GuSQ9MlH7XHaWfcLTgJMF2q8IxmSuhU257qv6LC9Sw2gsUh+wb7aiG4Kxj
Ze5jZCoQFE55SKPClMlvE9yD8e93qOegYnmPYqEmjaiyoGAoHS/dPA8Dlekv8DkW8qCL0mRw5hcU
lBXzRTlFPj9fsB1rShdNDWe8ONhHxr//YXU0xxvWdr+fbIdUVXLnrFsTvT2a0kEeC5XDb5Nlsv2d
ZPUwY6f358s7H/atPSnhM+3fKFh0prxxk+yfzdZUak2jyUMv/AwjacLOQ9gWHoQ7cf4CQcrGnWRe
SsrF4inq3amM7KDhGzkwg9AVXB4Ex9mOr77fjLNYgJ9pbrvLT/xUNF+hVkMTSDEKEA7AKhCEsaty
jUo5qf9QxF8N8p4FG2qB2q86lkIdBmTPOG0vJ9e67h8vsaEB5oB3nLPhDXW78GdLjddG8YkwKlSD
GffCxJ6WyiBxYjjEEMB5ta67HlYi87nC8jJj4u/Y/eNN1kwEE3yZh7psP/us2OuW3vyNB7Q2YtwX
wZWjxhnq13lN+C4SDAw1883bU6BFrG/MQm+Ol3ez2I1PNuuLc9ZO5wHHUPtHJJSQflygcsTdYnXt
MDd9VTNrDm4FZN4iWHmqXSUVR2ApQAgvChXchK59jADiPEvHQBKRbSpfSWuMZVwNl7aEi24VKyQ6
aQfPNJ+wo6jnwHRj/cV0u1+uiaQtYo5MnIEbOqOdI18O+Pq0zVJSaQgeZzAYLUp2fA8MHuLyojLj
0HGakgfAPUY2dnNjitQJC7CJMaj6kyDdorbr1g0lG1vhMkLlTvqhpWmBkvEObMOOa6sc+IQcWAAj
KyPi1n7ZmS65I+McBtsvdjqEIGspNtOpqC8m89xYEoOVO9884aGXPBNy+GMMu7QwxQqMWgQ7WMkj
+sbAN/R71I/iTITcQ2lw++VVaIEgzoBguClxRSf0tOaMbORGp0toSivLLGBh4sOqVrYcFBWR1hmL
XAsL2whJXZil4J2LGeLdrmtbvzntEazF4ZOa1LDQp4tSenWMfCXNAEZBnYrf+oaQwDqWWkMclsf6
uCQxzm5KSQwkNh0TaxXXs984eT1NAGqrlbMsoZf04mULXMu+U8ODTGFTBSosneIcxFF4NwLwx4Xz
s1ILsIqQOOOO/xCUJG7P1VpCbdWPGFOBEzn5vcXqs4rDOgLtEFpJNYY4bE85HdHhXSTS+CwQ6Vii
rr5nt0CrvnQe+2FRLA8zB7nsBPxSGYrXk3HAYRhb9hEwIroh4YBG7tLcvkfgGetZPoncqrJNQUM+
xPl5H0XeVnOCaOosXQ4GNQ9nHwwPZUBfmQ4ERLO/ZqneTWjLjOsdBiKT6F2qWUbmQbzImFV8YBsV
381YG+s+iu9dg0Lz/TeuHohbyGZ5MTcQZRWfJkvO0Inoc+ff8XzvyndmTBlnFyTjAgTq7/fh/7F7
JqrPjoIsAihgrUAcqmEr/Sdb7X0R2yIoYLNrICxP71/1FQvJnNY1NVloBnxFzMOPKtYvZ8lsJrQ4
6zLxEerg30J1UIImAhcm1a4bboEhHAUSRjezxgPIOXsde5rtU+nqhMI4wQIdOUkIfHygm2Yk521Y
50gRE6HoVFbk9motDSr+dS7FhmJJ7ONUKJibkRERI95xEFGFrRcK8SUBgHFoTVDizDSq5FwyGQht
7Yqcxuxyl6oiQ9a+hJefm1+8urO6hT3SXThJ9VnH0EdA1kE7W8wFGWVqZsjghSvdzFBU32EKLTgd
xcqzazSXn5shJXYiTmKI4nZAI0it/QdTyEh0ptRal6St1EZTBrtcPtZEGEmGiyssEcofev92yrSF
4i0WHt4/8EJQulaOWF9Z4r6pNzkEMniAYHMoJGS/O1OClufU4Dv6y1FB5rFRY6yBP195hgGbzZdW
XCfJjYY/M4ekUZIQeI+hCzX8pHAU6tLUP+lq+V3Njs3Klhx7m1OsXbPnOJ25EzjauTkp8ILSWqSx
dPBB3bpGHZE8R31ftM8y6IgkAK/gsB1qU+5lkq95E5m3npyH+ejeFi1dZEKA+mOO1oq+ttw74HoI
/0Z4cmQ6vazAcTksIaeWt1/rtIPMcNFukl30IcwZYDpPtON6QD1tCAiOMGBSQ5DL0R81LX53aAJT
EFuwSzVLwtBOO683u0GUHCsSEIxo8Q7APouM/sz4/SmAcQCuTiL2L8f0n7ujTsOWjilyu48zd9jk
hwJ3dVyUzBbbaPSBTtTvVjFE44gNUWPh+4E9TAbgK8adJabVVihag8xAQUFpmLvdfXIi2AOiK1DI
i85ffHYF5FqzU9lHgEE0Qpl4sDcuI+v4+IwoVNqzrNmi8Ek1TaWpJDdhkw+QwbMFM2uEIa6SV6rs
B05/aDNJeW1QkDw4qWyWcV4oz37GkLYPUwTriLx4Wlb0yuDK+GwVIjTG0QTpsK+/d5ONOuyKhrFw
PXj6z80qNLU5UBLmUI+33QJICdq0pLsEp5kR4mid4KvOkcGJ4wQ3Mk2Y56fCDVCbsw3cHcjmvUtk
dviFtj8ScSCMRMD2jPE/+H8nVF11u+ULTF4InRlfGTpw1fFA15dJwa6fzQ82WuC72AG0qGp1FJuO
jUweopNQSCzr3Tn+/TL6sS1Ig7SuWNmbyAVdxmn1RWaUxiOGOMtH1LQE6kjV9+GcG2XaGuIx4k/J
iOx37tM6hRL91G6AwI7Yhssbs460xbHGt2ZLHsyQ8zDu64z7cPXYi7bDkLVAff00qiOOpTVEkpnq
6x77Qpge2rlyihceLRyTbIdIYmB5InHHMraZrEaFFgOb4+9OJmNu6eIlZI2WQNdO2w+DYjFHuwA7
5qBBXKiGHPA1B7b9RDJhRPEXntTVsU06onV+Sjq2nk1a2SHHL7d7xRz+rU7IUMJgiRHZ+0VbwXma
keJrgN8XoN2JRGlT1NWFKZIkBd8hAKwzxA8/xEYum6yDuOZnf17mfQueMYRH/A6i3jM3pQ+GNLW2
XGJ6EhYdmvE6qqpyKKsZUFFYQkrWhiBH8CNiWXlEZzQOQ2dxHP6IMXXPy0AUIpir0S0PjH+1Ga+S
zrPpgI85rw7C568MS9ehM6NNpf6tifPdEUx76E11i5YFgbVr1brAQ4WOcBKywyVZNkWuJuzHmza9
ZasDALQyu9SpymDSKMr7BNEyTB5hmuJGU3sNcldw0As9CaTaiu74v4Uh0c8Afdpy6tekOyaQBeUg
M+YtQlqS+FqUgdPslNoyifqvDg2nIhb5gCqrwVF+3jJ/5KInH1PDN8CqJHlfXm92tb+d0DGNe48D
2a054WjVPa53kvndlxHjXz6HCCVfrfImMDMCFJsnaH+KEtgqgGlCRI2WrJzQIDpEexcPP36xxP3C
wu2DwE7iTE0CeCnQBb/WxPxKkc8XSIRAHEJjWW5BMlN99XjQSAJOJWV6zX/oBKm3GGOpwDnfzW+c
i9nLhfQLjLaPjNN7uiJ+DFoUr/iwu+yJ2lR6lpy7bv1C/Y3Hev1YfT+MHZMRITwrMvmfLI/bHd+g
IyDdFQxd3pslo8yf6FQouqEYMNQ8FRv6AutkaJk2HyK4/TztoIVsYEzty2zLRvhr3HNcBOt7DVQX
VYvEiX0Gbh+K7wyrc0VkrmcSu0GVgQTLNmlJ+Bh0popgyOWRTKRrGzWaFzISGMUuD4CbyLeBtQ/7
9HGrfjBVpNejeNGKIgL2U5Z48k5n+un6WA51CHckjqWXcVIyT10H/VnRMTQj8MO1JpdFxPWF/eZb
+G6ijdUB1crh75I2lrLdIjOl4pFKka6U4MQZQaYVuis835Q/JLuXSsAISmUsyzAbpvhfJHGfiHZV
QXFs2WbVHxXEdlr+uuFp/mJQd/to3LX0p4xxrlVAG+abucyM+XGKFlLOczs2wrCDaAxuB5JW9Aoj
kosxgA8sU14+34dth7HoPuR1+95EwYhtbtqZ8Lz+IbTLUC/iWZdRih3UZqr7GrMDkxR4fKH7vYBa
/y6v+Fqw0fGjlRQnvkV7Dmr/G0wMrGBYYh3uPwZRKqH9ato/fEcYJ0Ll56FtRnkUt547BwyM//97
VPY//H+PGd+DFNNIiY9kyEOWhGW4hDTyCWTPVM5R9b83bLEbKL4MXpjlBVjnRZsG+xg4GOh2I3D5
QbUPBnSchlzOjXQAOnbxGYDZCXNtQEyVEDkYmxFIwHuoZtOEnzf74jhpDq+oDbjJJEsgIJH1ZGak
70bpLI07rh25aBG0+bKBOPpdrOq4CRGFHONxzbiYD6TRW5lR5T09mU1YQ1fXt3DDKshAHMmgkEqf
YTVY74D6LcFUq/d49/7JF4lubNdxZxgx1W7WnVdD31E2a+2RXLrXXwoV2iHraeAdN6B6OVr4K2wN
M5aK8RYwIjq5R96mEtY5//3CdlC51Y/LIHIVYbSe3bEZY4+CHzrtYNac+gpw6d+nP+8qUq+nPOhw
NwpIYlnd9IImJA8Nb/QUDaOQDgq29SVLyK84R5ht6VHb2QPE4NMXvju0zRqW+k7IJbya+1Iyg8mN
v/YOJZ//YV7Echh3DaDymRlFAT9oSr+ohT/z5L16q1nwovaznoI3sDMUEwhRVFANLLRjmjVq07Uy
Mbh2QcUoZly9V7mM7635xypqZUES5ABTIKjfQy621vQqsOGTfFhC8Kjdyu4aWYd1ILZ3fRvunhT6
M5wi97Pfqw5tYJv03jkbA4v1W53fEDPZC1dbYouNagA/MXagnwPQ299UtZ2/2OASGzCagJ6pMIw7
klJUs20ZT4DgXjZqsKVNpeDsZV0Z/6Rblw/PZMRArPriL/YMH2W0J+TqBT0qUNYPwqVhE6bUP1xs
9o6d15fvoyk1A6q2y/SICx1sTc9UDtumJj1PjYBnlCYQ0EWf2tTyQlnEq21Sa0D7EfMMqwSmMTyC
46G7jLvB6PEFk9MyaNNdi7riqgvss1K7Q6fZY/6XHQkWfSufTqSaojFsVXz9moh0OYYvWYWlc2yI
+GC2EtTrZO6M+KivtEZ8M95VzgsvH2xdRrJGk/Wp+Hrbiv+yV18kldkxjOK7ukZUF6PrYRY+Tsw1
1EZFOLUbS0AKYtyoGXJzLc0H/kV4LDdDywrd2MbMRg+gTqNAUmxfNkjvMWTvUbJNRcNTUjP7wg4I
InZlBR+Is1OcT2akuclARMaTcfRDZVcNRtX8sqFbCviwweXP9nOHvekbxzXsoZZNl+FXXEYZt5gd
a/aKwLzeyiI8Lpg1OeTv0Rcs8IvuMgR8CO8RfwHDIqVhGgVzO9ZU4EB5NURtsuHJAc90d4nZaVR9
mksRh7+XxpkpmR3WNKpvMyABLK9q/tAAxn2eB0v1YZKbOxlbM05oEk4/Aw99OaO4CrwDNYfEumbk
OuqbMvLMYJMshsEPg/ZRDzYoDRPSw9G2n7tHRvWZ6j2j2kqM3tLwrhsVjbe3nSX8AfZxeAu4/6tN
bV79Yg9ocjCnPuxDTbOTddvD0xDAjYtHxT7JeWmdXcBoRwmmkRhJGXUw4Xvu4JUTOyjefjcHNpmB
pBfz+EpAb1Xs/lFWUnjkGO+679SENNQFUedm6FCk5AbvALWxETAF9VOqEkl9JPAGQSLdepQZaxGt
vPerUGsY9Jk7iyn1Dm1M+7kRMWm3PiNKmInQN4QOXNupuNr/bfCQm+Oq4grePDRDVtYtNQmz5Wdk
udq48o8dwIdEIrWs24zf05Z2fkfQxExwoVIWSdzlUSPMJAKXMhtu/Dm28pee4LAholiWAlkMdjG4
nWNod0esYhaFdBc4LUpt81K4eqeNUtomAxwsg7NtsOnN9N8QhUjxyM7V0nnvDqdGCWIfqGS/TN5L
ANb/8QmS7km1M7TnKYHUjzGJdYNpvowJhegSDF9Ga5E+v67ld/lqdDr3OcoHAZl2UF/vfhqFw//l
UpIDhNGYWCPzOHPYu6jQa9DckxYkEsJCo5wInIKKfS6Lx19l00TNpjukiuHZ58mg8XAhDVZLuKpO
sPNsCsJZ8ulLTn/4JINmfmwN62ZgNZIPVLaX407QGvu90uJQpnQkEQ6Jh7mRvZ1ra4gLrfdkcX9q
3PDYdCcm+cCAHRd5gbhxBzxeOaIlcdf36m96TIW/Sd93zTAwz42tfCtgI/5e6A01+yfEqwFZEeST
fua6MbKh0Wpsd+Duhnve90xcbnPVGtwQLYpSVrnXRi7Rcm9mqZKrjtVSa4uCQ2P96qRggwtHtXKw
4P28o0xTYOXie8MlaN9R380zluGexCBnGcbdUOoDZGFTyf6jQf6v9ACSLKUKeRI0hNlcRcS3GYOI
acz6fR+1YI/As6QD/n//20oL36j9NCPmaauv36ce0FZvc8DCFygeWn28/hTJS0guW5yArzUNk0mQ
MbPRsEZIhLSsvXVmPtC3DyIInnLRt/bnoVTuk10X9mbU5tc8182reqlbrwp7Im4qC2wPXffeNNsI
uXekhFZsuIwo4kpAjRzqulxxWYyYw5MquHwfBNY14zx+WR/EgY2JtvzDId2hz5M0IasPay4O8xTJ
zW2mmimLoBUH+GfVVBdw8o8XTB/yzmkus1xJuv+wCBuxt+1Lkmz8zUlOXqBgWVlmUw2fa0r97SU5
yyaW/zzvlrgM9D9TSgOWpKkt9hD20nm1KFeTWXTJQkh3csevslWCIystwNRK32JNpCU+Hklj9Tig
LGnebbg3oKzYKGruf+tlGAAcqazfoprqcvfYNes0pvWfcXl/JQkzOJiXiSJvbM+G2C9/NL8dYRWB
mD2An5Vkmi2Efx9FOCmPIdobqEOqG+L4SQlkAPDzslLZZHlE5lUG+/42IFk6a+3FWtjkL6weKA2p
TbQOyxnLMcudWQ+1r80skMykv7U8OFPW9tSMdXQTZcKx97tgYmbrmpnE8miiaskJZ+0ctAsQE66i
M/7Ux8y+jj0FNicUXiW0yrPnnPuiDrrlvgUX/bwxRvrwnvrNx+05ip/T7Hkl9cwFO3cdISqGZ3Ip
fbhsRdZRpKrZq1+dFeROjVVsSnWTaEb3LP9l1oDAiZItiMPu9i3L06+5fJ6d7yvSutvheBVHRJDI
16+5NHkRilXrXq0+WkEJwr5DMPnb5P7vsBoX/DJiTuDwJh8jQ3TcYTF++DK+mlsPCxX4V7rNIywN
rdB3kXeFqAiRx09GT12hLXqppFr3t4AzX8hLsoMY9fjUBwX9uS3emlrXsTK0DCVTX+W7Ofb2TuyC
O3nUrftgCOCXms5EGc6vTRnff7LYfqXI/Vh+Fr6G5mmit7KV8hnSrbRLlE/dovaqBX0fS1g4TeMb
LR3SYZPWX0JiZeXKL5WM5MYAt9V0fcfPY0MMYPmnGwCMyn54KHX5ibLehU3eY1TXkd/NDsZtvJv2
k9ViUe932SsersnNNezVSLsASGP5A3VjVdqZaRpPyA68v0pcBLBI1H91uT1s5naNbhimaCIzx+Lz
z4DMzZ8g0NTzjuDhI31Ie09RRF9WwQ3kt29KZbNjN/3Zrp84njxg2SD8C18FBpY3LTQtwp8p7ubP
stHxsaZ7B8UL5JAOy6LmrFs1zcMb4wjpTORWDQN/P49Vcmu9bwDtMgVZj2eDvqqz7MkIp/5cw18+
NRjWSSrWT5qQspgzusuksdHX1fiU8oCY0DhtlnB4gvgTvjQjhxS3E+OcVjxxsp0MPwDgZ0hStpmn
GBXB/P/DQmCtG72/Ah9HigPmTGzh4b4ZkAWZBjQOK14SXyofvVgD9Iu3Tr1+YhDLnOXqm0kTWWQv
Z2ojv4ZN8BcMDS3LragDvtIsfO7i9/ENcJoUbZ92Z69d+b1Fa30Qb3hT4civ8bKeMFj0eS458OR1
adsNxqeFhE45DGeeg38WaSsonKb209uw4E80V/2tCTd6lCsKeB/vxWwK0i0hWF0TwItsTrM/Ag2X
oqyxyuV2FiKuI4OGLYJiOgYWa641HydLBw995/NKy9+5yQUqLqh/qrHE/+nS10/14J0zhx7GbE38
XiIipJLWZxSWuptvzUHiEpLJjzLWdlRcllaWBewGBXnvHizOsuk3h4U9bvNbJY1CjB0UZOqOfBcy
wHRjihCengAWGDrQrVSityLFwh3l1nES3P5TzrazkRMwSiF797+KV27HOXXPD9BE8TVp4upJ1M99
eUAC/4Wh/GAJVDtr02r1cnduO/0Z9Adoz7/nrsKXpifROw6HaZvHLGEPvtPO+l16g5YLYwwb1wMT
EYl8bULaWlDG5fbjdGKBgRUeNX7ldY/ADNirOmmEA6GAuLGV/YDsyWzXRR7/CEEfYAEbXrlAt9Gw
oM3N6Q6v/xA4gGxBjHZT4vto71wHn+nEoEfV8Sy/WIV8f/NjIF62Gy77xk7MEfpESd6VihOZCQd4
aMNm3CRtpWpWA2uU8LrkzXsCtGAUDppGgBpjYaDOqIKu/RqGr00gv2CbsMPxaUk5spSvphY2GkbV
r2WvNEKf8ZduOhm0srSjSCLlFILccIDmGhpb7bxCDZIqS98BQlG9mA6k05pVEPgwPqY+G4WlIpY2
zmfr+r9Bco/udZ5jyop84Bo2sT4Uzo/S7kNii5e5tk0EA7jusbpf9k/Wbd2Lk75IZea+lIeUi86H
IHfXDw2nCxP3327Ni1vGynLnF37oQcMeoqVSTOu88pOPDchWUxCPpKt/cUy3yodJM9YCdSAehdMn
O81RxwHMsffA164r4SXuN8XCqTpilRwTSrEk+8uG5RigeP/5Dp3rP58Sa6VrPEGBlt2oqSZgrBoC
e/RrHQqdS10qyKDoVnDp3qFSiirgSPxDh5jvqUo8p8/sDHbex+a0PSWSI3sPoZT0Nl7EShFVFXsO
570kEMj3+d1aFU/+1SmYUfIbmqHekLsvY/1Khlyd3M3qniFY6wWSd3eyjgSn/EEtdN3nToQ2YEBc
qLnP5W9rKrpQ2IYc+PxjccflpvOuDoUX27zzdVrkT4ruDa07V9qCXIeQEE7B8osPgTuNWgJRUwTo
pYWYS/i8KlmNbakCrUt3PD858MDS9wJOS0ORO6XFrMcjIdiSqwkaTkuVXnyNTcnMxLp0KDeUphT3
Z1iY27qq+uXNFScszWKzFvAZlGkbftDDIZXxuGOizt+zi35+P3lLGfcurJm0neKWpmjQ5IRQ7fya
lxmUpKJLvnk4rj51bXuvqC+kxWHczynSxmNdVQqleyNC+X30pUq59WZGSyymXYczQwWfqhRDZHq2
RiK2MxEa3ta/myEDi6yFNdssSdIhjhle2JGUA07vSZJqmXcD5Xhh/Zqe4c87PaXc3GWgV24XZi1K
MPOa2CCDiJ/Cn0b4Py2o1iZeHvHWybaxyl5m3ThjEOdcrN/alfyGrTmIyLb8iSCmXLgdKhNQvNU2
o5GAKL2++akaW9SGC4h3unZKZ1yhhD/m4YYkqH7l9vTQqYj9wrzMZc2dNr7LVYCtasXJApfy14Zy
kUi9QaDjBHUIkiKhqE/dDQIgsyja/riz7W1qK+VdFsORaGoP3Ir8ldmS21dqz4n1aCW09svu3Ea7
g04wBeRnpxFlGUbFVak/6YYHdlM05JocOcwO5XId/zn9lZXHoz58vqdJQ9Pk3k1LmY95Lr0zhQsL
3tBMLHabSuXu4Ayqrs9SSVzNLmVGQ3WZKolpqXnYJvJuM96nECPQgH84S9Yorgn5OqJRCKZSNysb
8wcQIvtCTyBiZuGqTx/Ql/qT7GxOpV1yUDZVOZB/IuM2X32uvCJowsI15qeU/888EUlwpUZm6wyq
V2Is92b/p2kfZpsNApIOMt2MLAOaSkeb05lLdBTHQ7YDC9Momn1YEzusos2YqYrB9UOCNV8lpoXr
7Zlx5rXYxNB2tZ+tiCjK5FFbBHKzoJ9HnEx9BZQBxTgmQtgUIl8zDjzIbSwZmDoIdrygFlEcj03J
pBUIfoe/oqNHMInOS7o2PPtzdV3fV80Gf2WOCCnUeuCCnk6eF9FZ5W5YcgwsT01ZnjoFjHVFilpr
AXxoWvj55VP03Dm2rkDF5xZQOUrybwEBGvAXGqTknJ9QO0qZ7CmDfT9paxqCU/pdSg0xq6jv8o7P
rU1HBx8m0zR9Czu5dwuNsMMo3bypLBHfFx6GTAOEXIyW/wZJqF80j5hawig/QNYPJlLM1IegrQl3
fmZsSsHbrZWnVEM8ys75YMzqLwmUob56xeW0lKsEmVeMhRt/jfGE9bF67ovet38vied6+VzWWz42
2vy6GGs6uOKXMJjU6+kp6AohCVLORHvIskGIwSdYEmdDIUMv+rhPlh14wSx/Ou1/IE99fVCSSDxY
00WTawuMPKEZUJyDpcDP+4ZzfMHVSrnqnFflpiFHDu5QhVtKeHD13TVaCu3ii+2qrhaRkXAS//C6
Q5VmypocWVp/Q5zOGGPnuufoSg+AQ6EpAFVGTetnXhXLFzW82nQZbYZkRmbr791U9mrvzH00bHVQ
5Inzf/6P7aecMXvuwZBSeoN9CG1aqD/DEK1PC7KS4gWrk0yW6pzXHSrpb/OtFrJg2cdJWctDtDCp
G+G17SxVHGmeKtvots9pQ9S24xqD4hxKOw9qcO/SY78Ee/U6UxiotfkZWCibYJSCHiaDNslsO6RE
ppQed2mYrbEaGzTZOwKz42NTp5GDzj5uAGRbEebvMpEorZroBNvXiQEtHLKmRZyrccfFs0ufkSKE
ubhBZoepm+kQEFzGGG/5g5todaSEpNDN69fNi7LymPseDqRguTfkaep92wfKtaJxUw9VK6FYSOtE
qpmw8E6vfbuirM5kvllpjtoNkQ8SDOQ1vdB92kwCmV5suQbd
`protect end_protected
