`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
VuMqHrS/xayS0NiRMUADTngebRTMa20uGoJ2x568TTodUM+4Xj8dbIVBgaFt8zKLsbW/KzVw2dDN
8gRsioW1Ug==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UmttAWTAeIeyI2E4omE2H1fojD7i1LJuxYxoqrIenLDK7GrToBE9ZQbyxGOOSm6o0st5sDPZoMV+
H9VT5ab1PhXyxpglLSScoQgMQpYHZ0RT/bqtWYI9S33rXKErdm17MfnWTSdBRAu7Ix7eBp6GxHI5
rH4otpYVFqXtk8wk8+M=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hyvJ5Mo++nomOEV79YebXV6OeFhphscP30m3xI6gx5/d9CnNbGTNCcm1TqO309b9bbk8iiZzgacC
6S52jtPn3KfhWRj9AibzeCSCYXoohsiOJ23FkaCk+mwEkKlJ3mDjcZy26GLjwcjbScJNTsm/UHWK
PfIh8HPiCUpa3bg23lV5ulKM4YGRj2sBTa3W3JHs9lKcUGiQk9bOc/u28OTs135SpVlqZdnYASTc
tFBfJN2JCW/4L17BBDrKeCBGTYwLhUnmFIdUzMWbvQ+mjBjMFto9Rb5EwjveEvWs87csNxKyyZuU
4BylbByYGAIJOeAfXEyNVDuYfcxYVsz83GQjVg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
apAayz/ZFVHW8QiTkiDBE53TYOOUM27cyrpNlZPLylxG4talg9Gs1bWtQMhuv92kudZyfmMDM5E+
uVJJL9tgf7BUEr1+4j+Bs5mj/5T30ttdVw7NZtOBJlm+hnyis7VgW4moDk40uVRcWGvW2grm95C2
yN1pqt0YyFxA5XTvaQk=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
T3f2toNxNbI/z4gSmTtpZtoPSBtD1LYAig8ZJobiZAfaKcWJhPBPy0uESvxqT1tSULTyfOYXy71/
VHSw/hyQjbeWrnnypABG1W2vNN59SDdPFmNmIFh9Rasz7Gx3MAGlOml71nz0dK+sRawYp7dZ1/vg
irvlz57fdoEcM7tFi/NkE33tR52W8KfEwJz0lzGQ04cPC+ZwPWiro+BHMU7qo4tuCuwfFx93rrVB
uKWgxmZH7z85MxGlI28jxFE/WYFBcSr3yneidiPyAV7MwfJzHAARt7LcOsFb6vQ/mpIu/r8ImUmi
vu0EWLSfp4vLOhHmrc+hpFewJYHknRAcDik5FQ==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
obcug/Z4bGoLdEFnwbW2QJ9Ih1MzA12XZ+BHpOFzikBdXImU2p6kx/taVMG8aKD0fb9peqKJkrfl
+78bTc016wuX4T2h0OeVEOKMNfDZxJ3sXpS1Rk8YFBIk1Z06HvCCospfy8NSG2wnZIXaB2JHOSAl
tliuIAfzuoMjmeW8+tGymXm/tGg4TJX7PJjXFGALfRYEPd063CVaTkxVCG+3y5pm2OjjWlvsdebP
syQUjBCH4s+4D6dFlMH+C9gj+3lClfX9TaajeeXZgA295mNzShkA/e+hiwdPFRhACK6efYDTvX/H
UCY78gKh+fLozqDExWHfwXLODd4LMyNvc25qgQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9200)
`protect data_block
9sP0Vazx6v/wYVI7D/hLnIVvMifBeEf/hZn67w3J7Nvj17sM9IvX4IwXTpr4JZGCxZu1ubDbIk+t
K9b6fTF0SRFjIUoYUv9y+roip3FcbkNd8lyhf/ophfWp+W2XlC0Wb6Ni8Zw/kLFfnfr2cbAbxZnL
LJNOyo6YamRssfGm75s0h4k1BX0YamzGo3AWOJf2SbGoF6EQvQZw6g/btd3PxuAM24O1bcZdL4Ri
hpDXv21xka3e59HpMjwb6hyLTWLkzbAQbYAnpUqiwNeCe7cJtnq4byRe7kyJQzkKcEIqknHtsti5
6S1PaX66IMYg2rN9CrwuA73s7mWTI+fcObsh23Uw/XThpVfXJYgbYpIeFlTNL4Il+yiGkk6AGDYS
/kuuC3JknEvl8mKWzpLyteRwKQ1htzK2BvPbBKLyHXNOfXUz/DUxtm/0EuILFfpQE0sz/tmQUUXh
CD44jOb/J///d+p3ALjPXzFODr03ZrOe0M9SI4buqCODIxX7AHjtog5RD0erbt+W68751jUWptmG
sQr0RR2tcGX0111YolDVzzINd0t311kNQsQ6appLH1T7bFpNWIcigihDFN0jBqAB+26ZEHnKz+9d
pxs6inJAH9ZzOYakzZlLqmNND+u5AAEfiH8csYJoAWqv9GDftWHXsqAlDpl+PCSCOrLyM6S0vnQ8
Br9A5XybxblA8ztoARWeVDAHX7LQPBUbDOfsoNFdYI+MFUDjrKxhJAYwlfGU9apZr67Dsno/YnXz
QVBjeywaiv1spqK30TGlpEK3VSufOyyDmGLcLrRVK+l/XYARilH9YvwN8qA21l/zH7jyGF23UOV3
u1vd3j41gRA9f4GoVlieySoeGgUfYbEKLgq0IEhu7wpARKYxKXrYOgIbrZ9L4S6wM1hXvbP9Wfwb
h4g9cNXztVnCFe0u4C/HhBAMgOk5ArRqIIV6rd3WZFqLJnf5SXLVZrLx7/kT2FAU1ws0CLHl6x7o
EoZCcAy1njH+LGywmhlZ/7iFB3yZiT/JeDnxjwLciPOfjNt8eD8Iq9RIdzPDRO/0r9ADanIWPjDO
UM7uWs5wFT2MfEl+tDiGvDqPa72qCh63fw6ut20VQ64bvZoAlHXh1FXjmK5J6t5i+CRR/+jokMWc
TjqIqQHBhIWc4iJaWIMoQdsa2ngPk9+zsICq75tqlzgK4jYk1Tgj3Y50r0GpiYHDbwwL43jMzuqP
kvj53eAmc53RYLaeC09Oy3oSSTfO0hHgt9Tmes34hboaghSxl++VzJiKPniIoL05EumAfTfSYP0G
3P6SkshBtD9WJefWeL9VSi/AR+qLvrPQbtAz4vJTtDciiTGyQmuKhLqRfGfsFeTc2lJUmO7QqjCU
jn1ZgR/UcfYOzfV0+GhrRkidkBX2G25ioxQX99FuIiw1+4NIDwnIUf3o4ZkGsMomyMq+NfTNy5MX
1ipjMtji7gpMx5nVR1oJiR/DPdxWgQdj1MAY1xU1xVNRUA8bvYPdl6xS4ZuN/QRv+zkqY5mbz1OE
Fh5Hz3sZ0xZgY2EmzXeRb8cNAw6vFNbsHFA70EpbNlFa8nSD/8TP6A/F+TnWuYhd/zKeC/x/P5YS
dRtGnnIKWVZmVXQgN1ciEzHsjK5bGlGNFiFozfE2zTr6qgPH4jPe7HuCg+aJAbD+vBnKDHfjNrBo
lZAM54PxWmM+Op8+wOYdxCwzlY9zOIRvNesnCDq7RayP8wOaCumCY7WfpQRGuV1BLwlsok8OMFBj
2rpGcRgJwDtxz8u9Fk2UK+wkiLG/5WTgQXfxshecaXKqzeh36YSa/CITvxq8FAtijHciLw6tYyso
xxJpiJANoe1/sYtn4wxufBPawnNJynrTegI0tEw2FjBzi6KTUUAqam0TsuOc0IB76O3prZeVIOv3
Cw9dOUuN73nVfJdJHcWFDKCT9dQWyB/5aI/B7As2IegtSiZiWrU5+MH7JBPivxSCKbx4KB+7WXVG
MNHDjNSiqRtaSzJnNepWj+Z35zAKPCKJTsyxo1++iQoDTrFsC3O4OaVdXFX/q38qf3y2/GYX6Nix
wRecjRCJcwXTJhWehpkbIrAa/sErThOfql2j0Rq8bzGuADnSYQtLP5wE4dnkbTg2KIjLJ+yDVRRK
NnPWt/fkA3XjtwoO++wmQ2C+WjGi1RCd+IJ4EUvj2JRhIsZFcyFIA9qpLXU/cy2IeSp4YfLwTx2/
BijgEoK922pBgJPji6O4+x0/muKZLAe0dDCtU4yaII6f5XOCICr93jNoTTcqf7SpM4XsvBcvL39C
1FvRnQrdH7+rQMMUJk30G5pPF7lRUVk4vizYyAKaqsv+OuaJ/KSoSCrIU7+zCr6yCBahLCKXsNVO
IrSLjO6Mkc5MVab3obv1nXdl7Lncv8EioX+OXZTPs+CAaSTsIqcREc8QYrQpn2do3oXlWfPunLso
E9BlqkK/H+xQQsIRb1t8sN6oIMSy6VAfFU43S7yBNVGcGpHMHLJkT3h8f3r6C4rExjk05jHmXlp3
lk0gC+Xf6r8ZjQUYGjx4q9tuAL3axgFDI3k8622jI4X5FqP8xQkuV56Rgs6kYrWlZM1bMtFisYp+
GLQZ/sftymnV+375n5H/WFCvQkt7pKtMFkh+PLF74nfmtmAi1b9NxrWx+wc8mUSU9PeEgGapGedv
FMgqH3ls9DQbjpfHoHmjkIfkW95AkgZ8yQ+IxlOmseVC/vgO953sd+hkSbErokD7ixEUFLbItpX8
+Qh7s+gHIOOEYuKXjYtzTKtAulQljPNjY63fyRAfd0gUklvoXmWiGlhrkz0N1CSUhA7jRg0Gn3S6
ao7CjhlAqZlfAjl4EMgncJ+JUyr5HOk7S7N5RKpHiHKREdxY+rqyLLnv7batFv3+MVZd57D5pGJw
Kq/6RW4Vv9d71UTad7DaYtMhzfmt5FT4GXAixBGRsxmf4Ot0dpzpBx9b7JlPOl0tCpebOBVKlAIT
qVSImSciSzXL4Bze4vZC8VxjFKn+Mh5p+Z68brOmsC9ojfId+yNvHt0UxGNiz9UDdHBx7CClmqhn
PBK709ooe3b+5KKDJfx5GowqWicEQcK0e3hxb1Evw6pUVXxu4ONyJYKw7ronDtI1rgaubHFcQd8Q
ayRj3p+q6uCklWaxUR43QDN+U3I6gTS0ILfKoRwtPH5Y1hnHs1oECyThJsOJhCV7qdAku4gSQzcD
JGdtPN6uuIKzsnTi19AarVtlCmWyR8xUxz+5s8Y5eHpIImdXcXaU1K7PJeAw6qQTqgIoPRP4PwdF
0QgNH64dzYCYG3bnAVp9V64YX2CeqCWQqZd/9I3axRVqZPSUv93lNuPjwuN7B5gfXaH6vI3+391Z
J8wD6AZ9MjQDfnpQwQQjVgl4+zAiAv/Qn6yn5Va4NWApwL6bJLWi6MXS17J60FuW6COp218S7fua
1uOBfFNvw/Qd5m1uTQvAtKlh86ZkBmuc2PrOPoa0oYjVX5cXWxVSvBkEAXfuXK4jemQNlLcNPqV9
zZjXPZ80c9G8OLfsZFLAK4kGdcKO9579eW0qkf3EeRP7kdARTFiyf6lCbblIdN5ypPYJt43KJJ+1
gH4cJo6qDM5DvDG+0VwO4nYLXEx4cK3+A19yvJnyzjmjXz7i4ReIM/zRyV8PtGXqEd3Vc3I3nFNo
zfFAs0R290dOQEx/mEizvFzRo4uUF+2SENRKxQzHp4Gv22Pfvw4Pt7hw62EKX10wQIzd8hSQ4ldl
FJSJYDtUAlxaq0uFvbq3JodTifNwaJq7/VV0vEpxHhWb0Ik90vDt/py5eHc5kcy3p31illLPFXIo
LsHv1jzver/Sis1t6DbtcLaQ/UVrBLhIev5EKeUTlP3PA/9WmIivE+wannj6+6JqWDdoBwcOLdMP
bIXgPMvgmf9Z9U3vKWAPOoXtgvYNcHJKaHIrzQX8+la99a7QZ3fafXJmOEgodCMICotD22T0E1tm
xZMvC316CzXq10LB2m+P7/s+ee5el/3LPNQnjf8f1YgZA0hMBm1JS7sTe5R7ewHnEK3fHtjGGHsJ
0wfxTrVcAVipgns0tpBCoUYBengAnYJIYT1caDoH+NTCjTR+lUR9Qmm5he2DFSmVE3rg+iIHSPgm
KMEuwuHJjgE6YYpA90NQ4CwgAsq3lb8mVw1Q68xTvcdcJb2AopiXNMq4VTrTZ3JAYf7mtipn/r/g
1VGqTa0lPbFBHIxd7FMn5gIQ9W/KX/C8gRziuL3UgKfG+qA+eyy50qxpYv2cT+pjns5jKPHsAR+K
n8yehN0DsuH8z12V5Rsr673r7fpl6RUYiMdJvgZ3Q4OOUQ0C8dg43wOnc93BznQefFHvDyoBDZUY
opai/6Eu5/cj8ZXMlINRY/hq/ja4aKbsc/ENzBwoHpd0X7di01jXmKfLV7fc5rNtiCxNfgoBesv8
BegeTtkSJa4gpGu+g3ydO20RYaaBGpriVkXEmw+eGn4KcArwrfEpZA4sEmAJRylzoPNxmVkqtdPC
/Ug9AUQU3UhojqlhAUU7epNCPfDFGwhNq+DxwAWOhk7hlsNy+HTX611vRID3q7NCxDdAFp2taZH5
ZM0ydNGsZhegnPs90L+zdD/6lxo4cuyACp35NgKKZgfPuEzLlS/V+6ayDkDpDLs1p8C6HeWi4HNl
CZn77JzrnQGKsO9oN+1pQoU7Bse5ofJNJKQaGuj2OhcXmSoB1Pb/fw91rN68MVMr6QA3IuVu1FUe
9vp7q5L9u2jyJezMUw9M3eiZA+Hx+Rn8yeWRtkQcxhVWZnQCXt5B4hQRakW//SpL+gRE9NnXVS8i
Vf1vf36U8mJnY+6NqiorEuy3LWQEMnlE+V4Vr0Ed1isqHYdhNJJnNFHMQKLFzA8Zk9wxZ3YQ+5aT
msvncs2AZOYQyxj6JYvT5fLzNl7zCgfD5Zw+hNP+VRE8rNB2SpT8qfWXs8jHYk0v0ktAFZnU1r1R
CtyvgHy9piJD0mWWSU4rv3WDysCHRmp2b6kb/bv+dZqLebz/ipG3WAJ5u/SFRJoSFPFZQveR1rp5
UwoHO5QBA+PzYSLptn4EfRPd+Vm0oT4eMzcArHY9nHK/QG9LbYLeXkz5ObAMxbl1XEiOSIdJQY5m
3BTNchCNUYFDEFFhVeGICYBwkx0jSjHuLY2WlMiw1UBXcqY1oD43Xj3ZYLsxligvoURx3K50yeRl
2MlRLcA4O4eWkZrAaH1B28gOUW2pt2N0/QnGE91898gFIi59wshEfuRKWZvgaKNzS0m9bLYAENfB
lKSV4B6oWC1iKbpohAM+PHU5H5A/CCu7E6LxJYxnG8gI2z2e5x6UyW3b7NgxfVlS/LylAlcu1ofR
zFQBmmJN0Pk2ZXZxd/T+H0napc6OPvjEJp3aVrfCnuHExC0EvdktqdI4WLyVEshfcokHagQZPRVD
CgntOQzgZLoT7NRctce3qJjgt6/Ot8qQx/a9r8yKcpKtvz97YLOAM2FnesESsNlXDxlNr8rETLf/
zF3mY9Rp/CELFiWL9d4kBMaqmLsfRumQ7WFDFBZ4ZARgHQxbaqq3UQFmzdf5DOvbslRGTx7hbATc
9lEpKomhFYzqJf6JOi3EzdLIiiuqA+/Y7qpujieVMwguefpjmof2JVGgR716zCbhnZzzsGzqgM9/
DZWtW288neqiBNuecNysHSUD47kJqfk11GvW2MfbyfOM+leR5Ko0DaGVT6Gn81t0ex8vD3PrKBe8
/oOrJujGAiYgUbRLBfXrMGnOgMURsFXJGVxuAcUAdN1fq546i9g/auzg2sOJfeYod87zxAVg1W8L
uGKMAsYxynWrkINmyUID3CqYVGt8VJ4qlicXwpeSiNA8sSmIO9vqyfF/IF9jSzChjTlpIaa/l8jz
wZnoS6C00n4Yh2gs3pX/yt1QCeIUt0W19DTpVagsJLGaXTKgVUGq1CoWlp9Jqd9z8B0s5do5HGfC
lDB82mwn946jPwFuXHitvBDg8fOgjzPtaInODf/3pdGcvuu93Js/w2uNW2zOwPtEsz0Zmgx2U7KC
m08h+OTxU4VALMFVNm4KHxtusvZiWovpRriBBHlv+B3Whwq9LRIl4MgxPwQbolq4b17E2kXdx4ZS
p0kV+l3Jcb4E1QDrCE/44pstgVcWcqOdHCI1K+zjvASYlTDSOZ3/qaZbajYRNu+Rh4d6Wnk1PAEu
Gr8td4pmvFbMYMRqPJkf2HxTnDhPHsBaa2h+9bA2HVqkzFo4rbsmqexg4Eho+ZDNZBQFBljx1ase
HVkuqUvRuE5NdlK+vLUjzN4ZW6ukfikdksFh9WiNVpSbDKSKxlwNodA6x/IaQ5Xh5tZudbGz3HDj
vRepwwV74yC+iaagcvihfqmYRCHlZ8DH5xtuQRNQLiiDd9ygrbmDtKxNkGsrNVOfJO//Wl7Q5PJA
LfDeeL70rwNT8RSjcAXANGU6AYu6q5+0FZth/eWvMw6xu2aGqbOCiqO0H5dUw3BhRZctpUnWTFXG
6wtOpvDqal5rn/xShbat2vGa97urXuBrq/AxaAAmwJg3bC9ILxn3mNc7jdkv4pPyu6CrlUmiWwkU
MYU1Oefm1i89MWg8aPTZUamAcMoGub2qHdmHXl1lrZG/m+HpG8iHpda2nuvVxbA1EI5/aT+hH3VD
fLq+qYVPn7YSJ2vk8LiwJSR70S7pMfA9EZTWGSLXZo0/1WZs0bb0SWBU1NDDeHIQB+Nby/BWGGZK
Ad2D26F/uyjk8ONwCy2ebFV8jgNo8N4oTU8PQ3LyOcsO14aTt/7DhpXfxELYV817udsfsW6JlrxZ
rSSIhvPSh4VFPeVWLV5OMdbRawhkL27l1goYLqXI1C0eRtL+31dbClM3I2tn53a9Aw8EBOK/HOE5
0wfZMsZzsK72EDrOs4Vpj/OQ9w4ky7h1QzLqiHmUTXGfkAqU3uRjvsa+vkoENPUVjGcos+PymUQb
ORK18LRWcXB+3qmwrmITmCWddItp23yiRTjvQWr7bk/PEv4HBnmv265wtSa+lfI+jhW+aKG3qOY6
N/906kvey/X2n4+mx6mhHGmnNepsyF311fEHqv3i2i5cQ/eWpkP/qcqqV4hU0WBN4oUmTVU2wUcK
kMkB4C+QZA5SwgtJbZSl01P9vNDKI/uSGz6ncoLiN7XSvm3VbZVRy4lGgkNW5E4hMq2ggg4dz0ke
WaipX+3bidZjLZoI+wpgxKh2DOsTkl9lXAsLcksoiFLoSkYkjBgZvKlvwpS/GYBxg29CczzL7Ukv
t+zn7/sw8To5Rhxw/3VpH6qFNm9KOqMX23chA/Ag801ePMR/rO19WFu9iT6JjFELk5Dp/8BpEKLm
8SeJ1RXsVil31zvaR95iFsv62k6e8jJi3tSNBr3k9nzFdcd67WEjAR9WHJqMFueeY0AKgkbGbML8
7Hwc/iR0G4KyCjDxC0hpedMJXdKrhjS2NfvSmd/tBgm2kQKP5iaEHy4+XGIhRVdsSfP0BP2K6D/V
pFJLqxgGtzeCfu+xeaB6xgJ3Bia5W+wHTYrYlr1GGh0qyArxOzV+kf64dor6hGCCBTfiPbpyUqEM
vVb/dQ+U05dWlp8V/u6h/t4F9Rx9nBOMOGUcB9klbg+Lr/cdvuY+lt6ijhT9GlNcyxeCvl6z6eYO
rk+5gcijhSUuy3nNsbfN6hJdPJ0nIE42fdlrn9ZtojKOBe/W6os+lIcXeKUZPSG63jYT3bsUmDHQ
x2+7doavhp9m1TYBRzw9uKGPNF/7aZPCXHrs2ppIq7WCc90aipVHScpcin92RdMfYbFRuC93+BnP
DQMoP9o7Q0Z75pgH0FZExT97EumQ09bT/HIvzvKr08F5tprNrjzaIrjG+V7Xzh6qL5GsigMzoGKx
Pd8Pcp6ERRcsk2Sd75E7ZDWOMyiYKx4sPJ0CKd4jjL1nkpvFf7Da3ueAbQq0mEYQqok4jGufyG12
C8tggNJfNg7JQvZQ3N52MM2P15J21uo0ct5WSIENdFr6PpWoR97YwbpE8e/dko26Nz+2GIx5eS1e
3kX8Gu6/onq4sd868Eo62pF7q7VdfHNlwoJuE+a5XDXCHTVR1TO21CxwpHjL3qPKAooruS41myqI
OSCNlQNWfV3iGonTTg3ybj1cDTLZRIneS602hGYULonJaYWsYnCCqDkGu98MaqoYQS7Kguo31W8J
e089q67R+Ocgq7O5JtjtvIcM7A//ds6yiz0/rgmFOm7uSiRQ9sDQ9SuIDKhTSWN0wkcDa6NJsjRH
t2Myz1bO0/j6qYOmibtYgk8cp446Fpad1fhpFmxNvkVyhwveCUhXTc1ZHIGiY54BB486ir9u2gSO
wvEonAMe4XeFYT1hrVRHvnjV9Emulws5u5cGsFWSy5QH2v+BgWoXQ1PJv3N3otgOy1q9Ihc+ME0M
vUP+Irh1yOL0mnARUGAPzKlp6nbAUTB0bLzqTUXd5FZShNijp1+HjAiBZ11R72PIwDkhY023ZCOT
T81oTuaHfpIjiJOiv+l4M+dPqkBuRgXuFPT+rvnrp3y60HI18xfuJoperfLmHBeng2qrhkbXZLLo
ewc+c/XEvC7o2IUksEb9tHEleFYgU3XU2P/MH7R7T4a3NS2ZF3Dk9DBKklb2pHUO5L+Wz4Gu2/nP
XzVu3gvEYwSiSQc+HwNKWhgC6R07C6Pk1x+ivjxc18s9jCjMc4AWtwAxOs0/jmSxElUxeEhtsfdL
yQbUGTVVarh1SzaXO3rVHmEEdsGAsstMeKanmBgZlH+LypI0wI5d9FlsaxYZB2z+v/yInwAU+Mp6
ZKpuema9S3s4/DXUgj2jbh+2sNkqKH67stUPSidtcxzU2ro+VR3bGdsLKAg99lYSGubnOgq6KuiV
rGMBxejTwM2a7F9DMtYj5BuyUD5zySvEQnANUFIc4Xcjeqm/QUnjrkj5EftIw0GoG3KVXp23XYvD
n6gSJihrHq8p7QuuqSqcUlMvo1RaJ5JzLgPWOAlxWBPz2lLHDyGOW38a1URYlj7IYTDpcl/q3SA2
HaVkzklTftdPQp7WLf38lLUsSzunGGrh5KfVqSWgQRqAVZ8yD4qQ3qOxtFvtazFaRxeQqpSnU0z9
92mlfMtJttK2yLSFbLLJdNZ/pwNQOWHDqm5uWUh3hQ2raIAugDxHKRCn6S5XsLVa2YnPVCxvsA9T
UzX5mWrxaGgvg0txIOxP2IcNiCkDzDC3pG4u9JlxY8AuBNK4p2+zUM1Jo5MAYHQ6W3eLyWSk4gRr
q1Q+0P7qKGmr3PX6l69bJUr/DkpAxClituRjJcHnwl5MVqGL1fTEflqcbw1cW5ER77+ncFYCb2Ew
AOE/PoxNv8FPJ3SAafWK6OkhXx3fqQOc2yTslszYmOHr7SHueo0s1EtgZYWCFn7RVY0HDILWIE/Q
TeAOW4MUvuUC5+ATdHmGZELQazlk4okD4DLa58Ue9nfShMH8iuLC7b7JIhAaTWluY1zV3KOk391/
zhm398MfkAyPiwYp2h42etovllRhpW39klyz/k1ii8cfycyFtEU7xpnSaSjc+vMtyFeNDXg2oYMz
S1nGmwpjHyLuT89tPxVQk4oRnIUi/WUPV7VO6JnS/XMAoW7hFKtnjdwzQQ5Uzte3ybttCHJMdnx+
Vyuip2nAhIj0mrUTBtKs2LKzt2kv7XxRunGLsP2zaW6OBKqwReZvhzKaGgsrXzOBInVSbKyn8oMr
RF+DU5vmg4QMwbSD4neJrt5duT8B6ThkNT3UiLO/lm9s0iZiSWO5OQtCqrzL3xTszqnsSJ5kwLH8
zHBVcVEFM4qAfRxqnVmAQdTJl+4qf84H445tIkt0BGQ7kfgeqvczYpSA/bY9gFn5kigw6bhJfEe6
o4eJJGEt4+1oQEL0OFjw7jSFNmj1wLEY5TgNYcQ2wt517MGrbxSKSYc6QUCoUnSb1Mya6b9nMBiz
+zhjxU1ORzsk4YMXlVPTDcSX2OCFCZ3I7Zwc9iABr7SubFSyJjM0JcKeETpy+MQAlUE3vkM4FgrV
oSpWG+uF9qAGpYhoa2+wEx0yJx+Wic8vyH+Er86XqZLiOJ6sIJUEvyZJej8/cm1Rwws1PMhAq0en
qwmfJwwsFoFOVtNKgpWQ4nVoXsWw6jI3nkY4hTPR136E3ywyzZ3avJ+lIzkZZ99mMiUPqe32+YHy
fOg0W44AxN2eVu35zI/wyalJzGGFmg5ZmVJ2tXI20DKWYpKVPDCSO38rJG2WupvAUD/6gsZfd2yL
3V6o4rq+4jqiCCQ213n7JbW1BPXW59hZwbZ+ctFlsyhykkUTRM1tSVZrGADpE+uMKQCy3XNYZAYw
oBTi1wBXA3O108mMaCUCyvWAdwScvIxAD5CF3RvWPsLWt8MFSV7ac60rnU03uDq3KPenVTEJ2eEG
6d7k/KA09hq2zvQwtBBcX0lsOA3ZIye00dNrdzw6l1jPJIhctk/CcMcqEdnCryHNl6iQfL+XOKvJ
Ux28jv+qAUNepVtvX0tzO2gq1cCq9Z5TNGidKMsKxep7hoxwdGHtDAiNyUI58fQRZqbkhVVf3gOx
eFDfpN5SO3rq9ntHxztbz1Y5O7AMMo5pxDFLy5pgkcApVMfnKv5S36jIEMrWKA0dNMQ6ixl1iCfv
OuA2PzbiKQyhQXShjtWAECHtxnngxIscVyRYMPowwgf8es8BgtPtTftNWhORJ1z2NtHcG2tMROXB
Jnza0JWn6iQYGbFYkL2W9BDZpJvAIGJFcmspRlrE98JCvInHt5IYujMZYDQ0gw2KMozf3X0g8xIY
SsLUXrHmlwJiKHSlMZm1zdGaGjsQOMhkfUQNC0LTbB0At+X9yDh7pcoLY4WxJ7+64rtDJabOpKDG
aOFgG9u+jOE6oQe5sX9oP9WrkfW0i08EVvZYJyUxrRxGyYVci3adWjvI3tarboZ8apl2OgTeXbHd
J7MQqRrJE/N68P0f7IDmDu9hKe9g8b18cDapSoCE8//HczDfpnLIGkNurekD1oEfrw3ZgX3fE8Wh
v6AR7pNdnTFaXq3lkqkvkHK1dcbB3bwEeAnMjIAiYMCZkeRmE7lCrsaiqIgDJf4D0VSaENzdQR6a
O3ztuJpkyOCgxGWKTocztFFrZZ+w2GdsD8X2zz6K1wYbFvz29jnFLCCxOQ8nTiOlTG/qiB5BiN2l
o9jL+MzzUDwRNP9YM/RD/EVPdIfZdcagUxCkaN2qhaE+Z1XVkll0gLo+qzHPh1Wix+OMy9F+FwB7
7AIVfzq3QCmJUvxQ+AFpo/DnlGpGO0aPFlrFUrWR9l2DHZ50S8bn8EU7ZBXMbLanTCun6gcz68sM
O2tONUY3EveMsXsGbdfbZpMeJ5RrWtoEAQBnmqN4R0Q1+7P0mm0x1qPLXkMHKFl9xJ6vpPJ1YPm8
AM+JEQkDgdil+FNJaVxMpngBZSeIhXctBEfpEPZUvjZyDRu9fMCWYGJ7TAxe7bGTu5AcFUBVfD02
obGzTcrdh1L14an5adWgLMKFsBMqy+DhOMocjTyql1Cv7SLbnBWEl39XFt/Jo3b1G2bAx8e5jVUS
Gtcmiu1fQ53Qv7ThevOX9ZMSbF5baDKk/vT1dCDc2oEffU6weJv1kj/dvcXMAZi1wYKpeCDC029+
VW4qgAE1r9hdS3K+Dy0WcVSaBIzvkkBGp64kuYGagyETMS8X24B1gaFQ9VTBpc2+Dx/OMByzbcsX
uDRJXVbxe+AsWyVqAH1AlYcRHssLhmO1Q3eUynIwOzLaemKA7n+ffzuaHmcSnCb2c0hSMVVo+oAa
QWaytSVnQM34SDb7H9Ie5CScsD6Cm6IkDq6hqlHp5CNRsCKmFHqKUnovHLCMQ8pJq+F+PE6R2tgA
k3AkMvpos3RWRDR0Lp21WFZDh9ihN0AbdetKuwTAw+61/DJHzaPmJ4pD1fTiAQFFUPKR7BpbJSFY
wo6aeSPLBcRup0gJNffKfrS5X5gzBFvm7d4+oVXGKXrNxoxun1yP4CPcl85r78Xu3uEQFSbTU9GT
HQt3qDpADI+OhXdReGW+yT2qmA4AzJCbWox2KFRmBf0JoRdEvFb/fXkZB6hbYFLMFADMhiyFIKin
C7Z3B5qnK0OEO/ceHhXNUk7nJf99Yg1ri9TFG05v8oR3/307mDY4yVrS1ItwIi3yGhKvOisFDI0n
uCkcB7dGSG0vxbaXAajbW0Z/8V/xdJBEW8S/CSW5abXkmUXww450ksPHAljU2GnQ6vUVcAxr8aHl
Nw/QaNvbVdeTyUC8iLqxY0QGygrfV7/aY4og+7pybJ0SqxYSBjRfPvUszKbLE+5uX9SYG1I3yths
0U/NijUNiKdDIxc/o/xa+vr/nxfw1/E=
`protect end_protected
