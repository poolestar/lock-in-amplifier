`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
esfZMsYAfgXl5/1NVMN2HuBLk4mXIq9zMOJXIUmxxCM3ASB4oQAFnvlT0qQ4RqGCLuc6E4dp8YY2
YfiJ3qfTig==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
frxu3a0gIGzWZ457pzmi7vYKpjmibBj5oTp3Nm6xd6yFlKPuVeOksFAqb+1Vxk7jGbsjMJnyx9lO
2VKXV4xFQMpUDAQuLbkh4Vtlfy30FgH+DdYgyNlWu+/ODzAyTBwGnqBBJRWXNc9v+o6I4rmHj7/U
VClAoMEesC6jruAbbGM=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cbNyAAUaXpeCEE3+JUKhca5KQeGFeBJanH6xxovFyeGtuBoc0MuL7wNzVB+LMvIhz4ogjiNfjFOy
erJPWJYNTjakyBQ2KCH+8XKRfXaB/2Qfhk1ktmw/8Nf/WJvgEDtu2+L4gPKqwO93MNdWTVA+E/aE
EBCYg1ZfWdcg/UPLdBw=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
PY+Z0RSXvpKLK3Zrkj++I7214EYh7xr2/e4Nl8Wk/RJ2J3KnTrEGzLus2Svl+SvhU/JJwR8/pRtk
Cxuqgb2MDrHXlSxD+P9HB5/J22qYyCqHMtGZdRsOcTsKGMCCesuCLjP9Hf79ZOFvMD5UMWNYTypd
SD5yDOXbQROe5no4bzSGxG4mwA7f8MsN6m+OxrKBkJB/2o17+ooK4Myvs0AD4AQlgduQYIwshad1
8ZE/VsRTh1mVu30q0wUgNPRWy8fj8p6JpaA8jV8hCsEd1RGRrh3u9yhhQMb28Yu83JzQB0LgB7ZB
gCnOhR+tZ+mwm+CIz89fakBsAJimu/a5OY6MKQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dNcNGxdr//RTutUgFtbRa06+j0GA1Bd7CZ0/Mk8HTgXvP7VVhMJvKvhKuAbTr0+/BlPnahR6UpYE
24CESfI57v75X+wYHFYGhsX6tZbthCLib0Sl/VTasC+DsjOCPasfshwm3hfXJtHrXq+BsUAj2e+j
SqI2/OjpNly7duOdjFzqAXOFIdm4DPfjZ2jQcFNlbTakfh68WpouAv4QpD+GeJUHYkmBgyQKKgtl
kV3c3WXWtWPT6DNWrstlDYiptICqYAAarF9Vc8+xW7gOuASapokdaHPFVyRdYaG55LKcCbBoluiN
J36ka39JittR7uAN20t1F9SkIrGeDt2AOd/6wQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eBLWtB0cBWna58k7uCx8WeEcws/CCSVLQHDhus5dw5ZePa7yqWmtAPvzy3F0qB/J6Es6WuyvqRUL
eQ3fuCXQRyh2WJZ/Kvmg23btMGY42O+kURJL/q4m+kCBbHNX4N/4Tgod+6/h76nVmqHJ2tdXDXQ/
NyPjVMueCsIMEOgWo9XM2Ms0x8mfVwKpoAwo4XM+7wuieBHw+cV9rqJpcpV+YrXad3YbrR8+OPYL
LSjcbjQlXs+TxWG6Dg/fS0HI6HuXkMlNljKnltrG7PX95TytFSyszCrrivTmqPb9TX+lTOyPVegj
yyw5GA01VXWdd1hR2C7kl1PwHuL5GhOEDAzVIg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26688)
`protect data_block
YebvIxkdSh5cYUG/jfEfL+bA4Sf0Nh5YYIsCqPKJ0ezLEt0EDmfnsnOV3X4WwpJq+sE1E4DV+0vU
PT/8gG8B9yQJirNdmlYnxykgnFB2eLhpK2t1y9+me3sfmbquQ3dsw6xD3mk5pH6QNuAsBB69JWgq
vxBhoylAaDoWJ4a9JWO2purHnyXu0GQCyJEdjjEGs40K6j8nJMKpUsq5YZvO3OnVPGT/Gv7fpZXf
anEcpdfNh2uWP8X131L3yVRCHWPY0eex8+gtWPoFyvPgUQZjskUg+zMR6NuMXHvg2oECGWwJzvYw
4wJcwadPJMnsKReQCKjw416fyx37ewN6vbNEoUo4phhCTQRfXMXHkk3g1MEawehPxqyBAI9Xyxho
lBxMIfr1xePWuDqA/9vEArQ5A6ouIFIwfTwFs0kW5N8SlFMNJNGKdcDm9zLoPX13EOgIbD0jwBg3
TzTfNOgbXhkbmPVFcBZotNbCERKY57IhcEkz4+nvkmE+gCAVKXHKR2aT7XimCKU7Fe97E0ZJmzBl
ffh5XPkHuryUeZOAavI9OVcZtQ92lPgyKoVP4gsxU0X3wEYVcKmwcuULt2d37Eq6PMCAow79ObOC
Pv/a1OFckl+vV3mnv0DSNz4UGIM/FkcIJsd4MJO5YH5p7jAqpPfYIySVlRfDqwO2JGODrRuYfsRD
yrge0XCuORLrFMTG9dwLBrwjBnrVdPtSFv2N+1fsfcP8q6to404Zea9aTD/SLs91TzE2dqinVaLq
/SdDYGdRrRLd+EOu8DHm8wVOaJZXT84KV5j0Uv6UTecE5f05bMCEGSEPQe29wOxqClWOUKc9sLwZ
dbgYZBvtctrB8m+xvyaek6eo2lLTuEZa9qK1NTka70zUCjG2d+vff1+LM7wIQYWfTwEtbIL4o15L
xT/WtNBrh9GQjBApBtzgqesLaTi76tM/3Y43UpUJwwbBsY+A9vdakkrL8SwfuHY+sm67QQWKPsC0
UWxH4J9mbE5DeVptuqmCYR9DAMWEs/ritzr+cdeeHKY1ctDTqiY2T7N1e8QWWRWJOhKg9LG7CCrg
uGtVdzN6zqaH/wPlsZoW7eWYsnhkQwXfSUSPGxBYBTuPy0xol5/5/WJvChg3zGbmT5fzNVNWf2aq
eYXqoNGAK6192Nm+mdV9YtVsAW+7mAtvjQj7wmkL9rH/CTdoQgKRTIRyGySxsadKVIS3keMGVDcP
6q3EySW8kzf6zcHHvsus0uv6YyUGcgfv8za9UzinFrGOIfRgInThi/X+85pAwOh/N3yNOgQCnMs4
BGmJjiSRdHtvmBVj85v5SFOtdKICVfl6xptViKDlL75I3vL02f5uF79VOnLzymULj7L+5taPOSZq
f3XJgTC2YD2M0VIr0WhgahrzdRcFO95CR0nPcKy4sXJic4byDipMaz93JHf+UTJBJQSHWrNUzOp7
jDiHOijgS2wPCs4KeAQPC9sAd7H0jRTOCHRQopIl1ESDxertXRWDmVAFIrW0tuiGnW4ewRNL/OAK
IJ8aAFBJEoXiYP9K0QLG2kWem5E08AJkWfb5bETnh8Ao5XSViy48/JUVXGUa7A1WKehThwjc6g+f
tnTSN6KZViOLcG7b9Nrq32eVd6O3NsDXyqaigJpMJbe/ho3ppKmUPveM7MAlnUiD3GNvZlX1/r+j
doA/Rl/Ia2HOyuY28eWs0fvzm2CeVVV5TcLEeqdP49ciqQsN5ic1HmdiZCdHj1qXKfhWj8nRKdny
vWPUHRzR1XEki9dvf4PtEl6q2gNLH/APjqi4Ptm4IYFtOU+a51e5wSgcUEt+0pn7CXfExvo4Q22I
n9av6ld3w6/4n4nQl7YSdjgCxd3vNkrb0XeZ/hfmupCWQPDKaAxVm5fqrgpPaWX5F41Twh3hv1BU
vBv2QAiIH/LqpM8YSPwXzGoBcRt+G1Y7oH1fkdUYqC8kyXikoAK2A5tBX4SnF3x6RodilmhCH+5P
5FMiHayNyzbPJDLDbpHPptrO63uz5btUKKFYjJZ/uGvgdUktRKsMNStWyLJxmcYsMlrQJe7gJdjB
8qsrBuo3zan45MeePD6UVQRFrhYLpZXIw9qC/oSdZUOHqn2EdAthqC22wYWxSUuuKKwPdcQsz5R3
AUB9UAqGZT13HHqhcYIsKm4MwNsJOSyAXs9Oof97EDfQqfICUZlRnJkCo1ZBKmQ7QmlSnq9CIpfb
w5CUwG24jE3LvmcG6UheuCbhckpZ0Fj43r5MnxFb1GEvwpw7B+XH+7ttef3SMCHdz2vJDaWYA5/w
015okTod25tUDJNdQSNaEfc6AsOxHrgpMHxDLl3AGI74unAaqlC167GTyZoZC6EBunXHPQX9pJfF
O7pJjeySuVM1DyKB0YQGbgI6di8k9lmAgxfozJzI2Ru8zqJ1IQ3Yai4dSP/+a1KwcvfudVzJTdZW
5zmtqWK1GRq37cDj+IWA606G7X+qKr2D7qD/zWxqTuRjus1BoMXMflXjeRfoGMyhrjx8IKNKznUy
97g8JVsi+z51PFDmL6LqckkMQzDdqPZUJljhhsMA/kxvazsVn+SeE5qFeCeCHJLBzorbbH+v36zg
CUlr4PkXuRa09H8O+6iMLtPzkda22VruII7PKcx32WcwDhNvoHhUHUQbIPS0Q6IdcORvip59wMB/
rlyqf5cKuYnoG/TdFuuNjttojYNPh07HL44l9a+OXYh3i+IOCB1vyA+jpMIzoBP/XwcBWfeb+ZVW
mraLaDQW81eJP65TDfWU0EorZj02/+HsU+MbkYWEQdbbC4GJZzYjz4WYGHqFSCK6FEm8TXBlnv9k
x0s/zq7kE5c5xt+7YBSsCa3Yl+f719hnFll9JVMc8Q38a9RJyWF0qAqwqON/+oH900BDuFo8a7H1
0Tqil0uo7ha1zER+AZAM37h344fgpXrlXrMAqlwOZUBfRuo45OhQxLlPnoy6xtNRW/VJoIk95rfp
qlK8WV4HzuOw0X6vBMNYLDQPu8nN1ZJ8iBWVpmK1cSoVsoMePEfjjOljmOcxNI6P1hAHrlLTAsHQ
6um38NLaoRbtQlnmLQmZu/yfUzTdmeZ6zD0Uhsh31DoTRappkxm/OOpCrO2bzGzVD84g/QK8HCS+
OWGuyzglZTGCyi1IjpBXI7Z2bl00TUq55vtglRhLHM3aJ/s1GMgML/3d9Y6cI9eXNFuiycEdx1zv
W8hncjLEeZdfOxE6R3XXvGBHLBYsko+MBBFt7Kbg26Kpa5fLEcAx6U7vOjoUDaiHtyne3mb64xOM
p9ubH9GkrH/YDbLOHBp29E7uf5T81o00C6fkT1pq/lSQIKW6YTm0nIeXF6IGQWRw52VuEzzdKfK/
sD8h6JxjGa9yD+htZtKWZF7NqP2MPV8GMs/aDSkfnuSNF6zSTiWrivEhib3L9gc3NEDKCef7hAKz
Ns3AZhY53j/aYcTssgiYLe8A2ZFCB8GDjK73UHad09yY4U+BHPfXDDDLA2Lc8O3/b7luaVFPXTEf
mDCpaKAdA9KM7QO84E7G1F/QLQ/T31VYXRvpHayKVPsNug/TnbP9exuUQ/N/mVfUtomBLiGihzeD
jsTJj0UWIUhzvXlBQTgG24S179UEbp7mTrP4Vq0LipupRvQcDdAJc98l5hlLNrjQXnaViWFcn9l8
jMARa726MftD/+b7URU6iqKknnbP9KQ4Ywh+Ocd5+ivorKnJYWQl2BFaGbXL2MOChtMLSFIxrOTc
4FMvosg/Z1//Iw6LOz4fFMCzGUerZr5l3yzT4rm8p+F8JkqnAcJOzyROccxNoST41NQKvk6Sv4BN
ap1wtoNCm0uml+x1Y3HJplFUYPxX/EuxC+Of8DR/Oxo89jEHpN4lESriybchl21DJdqu1QWwSCFc
ctPOYZz0i3JIWFUzzZmfqJf03gD3qIPH0Z4+OX6xlgDJUXQA+HLkIl+QjlAYpXs690GBu5xmbRdI
xCAyc1Nd3HMnbalUO0x6+LNYdp6giRMZCVKs4Ywuv9zTEpn216wTfPhDmphlQVojQOjqiv7PEsa7
z/34eN3q2sPeS9RLtVFr0NvRQPIeTHdq/IzoINqHCDi+YuE6pQTYEckUhcxLqnqJpM45PKtPF0wt
XBKn5eGuGUwoP/PhKx6RVjgG5nCleo91tru+/9NQnEvW51Ak4yzXZGBrq378kXW2z1AQSMpFH83Q
VjbqSHQbvzFRZHA50eqp4iwgQQd7mHv6ZY7UlPFKQu9QnY3YJws6XUCXkFI+ikCpIateRddzXFLW
74ilL5aJdBlrwWD8tos1RgKEcRpQuoz3jePFDTjahJCD+DFTblCIv/m92EXavWEiv41+pFcrp+/v
vd5jQfI8OBH0Xv/MethtLeUdQOD2Tq29z7ek5oMLzcgVlU4cPQYmYDTjCNpMCs3ZjhRKOHQRATQF
R19a4JeA1iOQv33rc67WGB1LzsGnG3v+KQXvmbBzct0e4cA6el4U7t0VuxKvi+CeFYaAwc6+e5ef
DuApAU4z5VOVK4VrQRgZRCop8f2Hur+e/Gw8pHyfDnLK8SdrlCQaRzccsWQtuFqz5DoOxKUOUX4i
zLwyJTgr3kSv6MM39U6OCfwzkb8EmGWwxZ1OUtE5nvCmW+HumbSFqwTtP0GAVIgdrGSO5rS2UvQv
tNHQaLaAIYgoHyzacUyVFOdCuUCvhB7p2PeHskieql6x+y5+r6do4W1OyY+qAhHSy/bQLAciKem+
o6UO9sprVq8bNF5mtcNI0lnPMLD/vJa2p5bBrC5tsfPrbtVnIK8ZP6CCfzPI7luvQWVTkZGnczqu
ZjgefCPe6l5z7vjxVGGEQPpmN4zq1aauwMvnczi3jlrgxAt+3wQd8CCexYJohkMiDkaBpZKqj8Tk
LhGqIklJaIuN2RqjWN0ZVqkgv43nkQnpw0n/7IMB/Q7d6jIeYnalvx/8N69shWphw5pA8VYKt5Hn
MdvdSZQ2BILa29Hu+mC+doY8rkag+FVLpIdu2Q74cJUpnVFE0BOTBLEZZ9ZexcQ31djIqhdXRFIp
qaafZqzfBz9y9ZJkoVRgBBS8t1/GPl0MlXZsy6W/KpYGO7AJZEsrgIbnqYkXqD5uxTxxEzpCaysl
U4NWb3P3YrFvE7fauSFSfIbYTbRHoKDxDEcSQpQzLO+KVTcdlCCTpSB/n6K3NHDznL5C6L50LtMv
ogukIpXkwQlG03WLzkSVjtT0GC+tcXTQFiAsbx5r6ibessgthK9EKcLU222LJEKg3s55H/8pAhkJ
MWZOHf3aRk54yBnhiixSej/bbBa11YisORawErAzAt40+rAKOct9lSEBUF+Xv0d2DdLMAn26WJIM
I7+KHMyydhOXhOKsEePwjyXZWGDztBGem+zkU6whDvSeAoryj1GDrK1dvKeSgMsU460o+Ix24nLY
q7Vz/bsnvjWDlmm7BNQwHBCTFGsS2AmEmI6dccedbkf5SbG6oKc4IvYPxq8V+NPek8/Bbobr741M
vUqgmGvyFMdiZrZBgd/7I9lZSaq2erKauTl9Et8DImGIzBU25haybswWBpsSPqgWmNFUGGknE19N
qidq8DCp0yZhoxG5InLuahhCozWZJN2X9lg1eRVqhHFHxtbhghntrdkavxmw/Sr4mSTaH/DjlzRj
OHUvxXabY8nrWnHKeK1fzff5cUnlai9Lc/3AYx1h5PaVVRq2NBPTac+pggbD/C36PSFuzLYy9794
we56hDHXKCGyyi4m3Cg0qj5H01m7bvKN+KMGOY4LsIKRJ9Aqzt/3mZ40ijQv0mMwgQdZTrBLEE2u
v1fYz8etY0Dt6/tz4xcgsp5UfTt/VEfvAxILKopWTsyq4kHsDHJmWNlcGR8OxGTXjs/FsEjv89xP
jI47UHmDXjNLi+jYxLx0A4lANo1LHPBo+Se/8GK2xH/55+zqeR5CIdUoblZnFE3Pjvwa+jdHegYZ
D4D6DJt1nJbgVoXde0EtgANLb5+RMGY2KMrfYwgP2btbFRM+CREcsVe3aE/R0IwsyVw4uRkqeGRC
71O36erWD42C8Vy6wc/zjzgbRmrupZTYIuQqmGph3h/j4sul6H3dPfnv0wkgOcmIk5jyoSbd12C1
Ams6Uh3ixiHKxcvov4nEs6WlECaflQwTTm1AMOKrcXV40sI3cPBUY2oc/3lK2k/el0BvKjyn+EpO
gYLGisK5cxl3QwS+LQJJPNvXhvpLtpGLY8n1lh9RqtXgHi8MNraMKsfxcoE2s4zcCh86eUVJ30qZ
IVniPxTpSoc4qe/Ku8cfozoT6T6FS1taBohlaijaEI6FSZnB9Ue6wWCfv/z4kg9Vualh/obsxOBY
wOGD073MXWhdOPRTtxX+sYnp3prz99Ihu1h4M/WeV0ES/oEQ8WFcbdcHMa5LiMyMRfb4JyF579hr
eD86+A9IRLn7GjtU7JZGKnbs8xfds41rErPGHV/1G1NKsD46ywMZpIoSxZEyPp44j02WhNnw99fc
qxN8ENU4RepnGrD1lLWgm/Cls4TE9cf+4YDIWDfYH2osvMZcMcehTxy6JPx+cgIg1fxYWT2nY7oP
XPhkHBT+maJEQcPWN5b5UvVTRM3FmJ1B2bp/8fqgDtbN03vJ9cWGK2oz3F2Gv7VIKvYOnmINq0qm
MbDXLu1VF08PVixBSd/F+B1AC13B8w0iV1UhwCKEuq8mR2Pzah34t6A0EbMe77aswmN2q1xg7ER4
Vvlgq/V5Ko4oNFzuMySPmBB8SHEM+B3CRS1OxEXxaU8YBrP8hPmmwlHjByeN9CFHfk9/L2d/hahy
y4PkrFQrAm2SAUpSmUsAeTuWdYMjpkkfLlCLoFqOVMH4dqqL83YnQ3ncNsneCSz179ZrHr/DKXxA
PzgWhK3BYD4qASb6a8GfWSGzafxn+f2HQYr3lpUKDLZmeWatY5uLLnF6KpyItK6up9BNvxpht8pp
56l6lHMFqf9P0toLd9sUPIJX9S4N7sPrZcPJtQr3tARHJoCYHBnZcSdGTflUywQG9txhaMj5DMow
VmJ6lIbk8Ay3K3jiicjq4jD34+HJAw8L4xGnY/DStCih/o05R3rBfyrymBMUZRxt29Kp4+qwcBkH
Vy+eOO7HX4KAO/lMwrMom7Spta+xPX+ygAHr6lxqFdgRAO1mv1PbWkfd4GmqIn3VpLO9Nnx1BOwN
0L3LzSwGXxK68WtFiJm7fprF5dQJkyfBEQkukI/HpYqbzXYujuNoUnpwo1wCh4TOGdaqhs21if+0
dMeFQl0k7h0rn6F27z1r5oWJylM5U4hc5CoVCW3stf9YuevwzfA6xuG98mzxMwWAxJyyO+QqMYRX
/wF8QwCDAHytYiMKiok7tUKhImKAp+CpWztaJjo/Z6gFQbW6LJIGmLVhIaM9gzeq3xaXILE5SUPK
C4TLv/Co9Weha5dgMq90+JlNQHyrx7IoVn5J9ODukmoF1z2o5/gaN5yvAoy8jueDVh8nNsCAGx5F
qCLnLe5/lzCN/KjVX3sS3hF5NpZRm/Qtc2+kFFQdHQG8gWbBfadKupwO4fF+yG7rZT0rmE1664bl
AtT3KFlh5GjbOW9+dcXT5ejYAVvNoYRo9Oawa86XtUtiWVrVyiKlx+crsjP/PV+IWrip3+CK4dHp
JWC9B/uu4Ri1C8isAJNHbJtKg0zlTW20fESkAuvxZzoyhIiT7bYtBsl2sF1VsstacspJ+pywPaii
eDiR4jio7pARAyXcxlX2TLFHdJMs5aAAmUmr5B1VMabWhHDhs3F2Q1HrlQ5lWRqESfC6oldYXhdo
n/7rWr4nsVLBjqzmcjHX2jgZOUro4nPYkOdhgTpU9pywhm6TU4w6Iype+c95DynD2mP8F9xeJdpr
6ydu2sSiSmXvX2+hG8nUUuEhPqRb4GUpNgBZSbakgO8nWchAmBIK4QvGkQ9dfcg37ohrZmliC3xU
IVgkWOJvkF3AhVWk2ZJTi6gFklH0a7/g1ZFTk5Id+5HCRVtVcxwOyBoXPbQbrIMadSAIL/dBS6IO
nn7mzMSOf1MwIb83QrvQM2L6HwxadjgrZx/2ZoVUPzpki7QfjiKnFV9jcYjudZ2ufOrfMHpwg//n
bMnvoq8/orKBIYrWXFm+BXNw8bPNGrcAnH0BVuVsdYmbylaroh5zCf8VBTrpt7zX4rBKx2GntK3F
5auKM7R2Wnch0+hoNOgYQgnGM9JY5ms9c+xCbS2glfb6gLdObscYC0rpoCNOCM7mo1cxGY/UY02D
Xc3fJETdoCqMX7rZ1W4y0cFXEfeoH9jUCmreyygNQancX+HTjccnzgaAoyIML629J7qyr5pPRYOP
1DfnPDHcytptq7/W+LYKxnPc6U5+1EOqSrLt/MmFdeW6HNwTy7dmds8ES6QD3ggxP1ca5R9m8KN5
5/o6GnjejrLkF4wR/0g4JwZVuxxV+7S/njBtuMzPVwXKW8QqJ33izOfPXjYi9EXfvN5f0ckSx/ov
1doUCV6l3KcVcorQEfTFnxpWUtFpD5byYOqOA2eeg/cnttoPfLW31egZ5dkQm0JJVwtbpZ0tKiy4
+yXOFs4r23zX4/aW7HCbvrMVtjRjgAcO8ycRkiIbKNGRdKh8GrJgohWyl1Kp4RR9D8u4/FpDFHw7
s7IK95Uv1Nmh1FpQi8FkKv8cl+b+2eySdgM4yRXnC/sLJJ3MBrJTPXXvvLekRc+L59q70Bav4C6j
qvw6+ja2s0CBGzrhfrY44vjPPk9aZuPj+LRFsXnQEx1DIVl+3ih+qtizuMmeeIdWyFyM0P/IHEYN
6AgDmvTHayup29Vh41alMFPD8JQR6lXbEKn5cm6gbJuiKSnxuDtD3GHDjsqOor0FeM9P8qCGsVSB
0ZXDIWRU4D0REId1xQXvwQdBwKq/UQK9oybhSUQGxss0lNOd4biiNioHyYX99wIfE3Ds8hYmDxdE
CPNFNTDVKn3w/hCcHW4g2Y65DgOmaQVBhO0LeKTKq4bzN90fhg1aTQy33ldmxVRnho8kiJxMcEju
8+w8g1zcnowthc2ybfdPM9Zgwh4jrmfJqtFuCalzq9WtM5Lw9sp22FaK261wmb4jH94Wq8QQFkQM
hsAxbm4vlcYOmsymJn2Xnnd0fYW+rbGoRobE1FelL3BVx+4mqZdRZACw4+0GKTVWR1Ingefcugy5
2641/2qmiuYvot4aSxRLmN2xD42DU/L6dFag1GgAp1xK+mvhKGF0RWsZhrslBnIxNYHwYWetoNrB
DV/++w7ay5eSs4etNpM5swZ5drzk3tx20z20E3dANRez39r3flLyS3mV+i2tv2dtH6ZdM6GdRQuI
A4rdf7UctYcVpni0Rv4HmgEXHQ0GfuCgiI2GWimpW2IEQYUsvbHtYHProro7sz1e69y8XbQByFS0
eg3Rr24bnstvu7neV8EpqkxF/aH4UNbM3MuCfWn1zB2FU93JDgn9xVAJzNcCTn34c/0DvlJ/k9tq
NWBRhIwMvXzMQ6LDoQRYxfm6tgx/teAKgQewEr4g7XUOqp8uIMVb8c6vThJj3E7qGc9NijvubTUj
CQSv5/KtuxpLU62D91BQERlJpTHDca13Yw4yP1HIyWzOiMfq8er9nNQ2GfxfE0mKnBib+PooOj4j
O5alsxRLyFAIQhHpOdLzyhbjgE6LgTR0ek5+RLZjPUaDKi0LZvsNrh190vCh0iz2YWxaT9Be+cTQ
fM4IqU2elOcxanou2uUV6+e3AGGUExyjq17w2VWHl+nm9uanlpnjp+YABp232lrWALJ767DbRyZP
Qwg6eid5XKawoca4QQtIBLp5QrZNEnKgQkKH5ofp4DstUG8c+KLMh5T3IRBDgKH+59M5jYRqWtJj
QskZETNkWYiyHQ0jIq4H2gLVBOUVQbLKJo2Nd1IOrohRn3FyotYIErEAItNm+n3zvAc0AxsLronb
lz56i7Q1QwkkwJKw1NXbAIcebpERrVGE6Op5tVwgH7AYwed4QLpZjOuB5HF+wdqmZyefHyJJNiS6
g5O/bYfownnu9p9Xtd1aA0YBdax0tWJk/UED7K8gXNzan/7Jt7l0qtrsB5s3UblFtG4P8EyoPo1M
Zzy7gx75+M9bF6FTRCTgyRMR+A8jxCbZSXNy8x6S0XyO75gs3kx5oTGes2OmN9zY+ID5EWsY/cuf
BtdyEiEVHqfydD5tHIsdTp/IHyUNuyRwvxGnEG4e8nWwpyp078kgNblX4coWSgCvqDts48elG3Ll
i0xR6xSuS0WzE42q6tZIbE2V4AQz8+Lka+FvhYESKcBEjafoso5iqOC4ryekLMqMYvQW1n1qfpbF
b6hj8+OVb1jwgkVMu2ox96HcTFqKzL4hbvEmS2OU4DEAX60ZoHXGuWZNTth5OPdHkgiFKrO24yyL
li6cnWwkTpSXUdhAM/RPJS6XbQyWV1kWBWS/JNMuR3pc2v2GkD/q8vMyMcxTZm87EFEaArWvXIYk
RLn9hKwkhx+ifDLMIBBStBd3qf5Rt7ZW/ryy4Y/fvAq/vl7db45+Oh6ISTmiEej4jr5ExwrMhW1E
gpKkYo+i9CMnSdzQU/dWJSLfDtOTfItqcFX6HLWKYYeHDG541zYsAcOOi8ApjM7/0MzSrDTriKEH
/YG9FBbXXBLtwBECr/ZPz4NYNVFC29nUDA1DYXR2ilNui1BL59UiKUO3eMkSl7ewmuavvt2fB60I
Fsr3jj90Rgqn9FdPJMa6TYhFFTfQLE6Qf41Exac+i520359YELhJj6B+nb+45lfaPeKWK3hTkGOy
MYHOazU9UIYM1AepajempbqKvMfGfwcwlNkd/TLVtz+4EmsdeBsaDulZWvKgDSMc/q95T9LbTEz1
vBtQPd28wBs1bst6btrqIWpJHoeFVdCWZ+/DdXQStegFrcXrm6MPiWyIshwaWM4hWG0gdaUVHgr3
KZNRTUpAe2onaZ1e6AgQAWS+jaf9hoeUihyvOstpGhYrG4KnL8f0kw9Fs01KwFxd6DEsDbk86WQf
AY9V0LEhDEN2u3qcva4BEUqSDzvD+7AiRrHQrzRp0ImtCy+ZLrTMk5lIJjXkLWjRA0vQs3Eh4W1d
5kV5POwzVVcOz9yWDBKIlm+kAGt6DSCfZyJlLQcN0F109gLaT2sg606oO9/05G5dXaLopZvRn38g
mrxZDNIF0Fk7IaZF7j6qAPvkEKsddngTYL+f4yseZbWC4OPdANmKecefTjeiFLJGS7FZBi9W7olS
BbM83aCbFkVtFeQ38RgfvXbGQh0nfu9tndEo4b/MnIpmgtWyEoZpvJyZ7kiGYu8eF3ncurjk04tn
HKDpkEr7HcgaaOjEL5XyjSqghF/wiy8DqO8bmHuRaB30y+fZ+VD4jl4h1OkR2xV3ZHw4yoS84rh2
vf3VJGvQ0sxJfHyeYSLykgeYH0TaIKXVbEFbi5ZOiZONb5J3FC88TxTl6Km1ZSNHO5Pk0epBfDa9
HFvVCfD3tbOlcDdjt/riZxjraee42To6zaTclovNYPfjdXqlYwrNMLPuZLFB6xaJcIkCG5A9K3ch
Bk+vBVdvjpiXHM3Yov8zPS/hqoJyo5izHmwX4PSJe0YfN6+3Pp5GWXR37M5I0auCLtMaIA/JPzo0
5XW1362j2RNzYJ2pywhnFor15e7+pXrKZTGqwvfwzfqsX2Ip5SSA1Cod2YsGvjxic8IA+18gjs0I
waoKuPJjH75K8Ph4IXLZgrikH3T00bbWyblWj04jakAjxPqfuDBi1tUrKjE4VdAtpsP9TXv1kTyW
+pOJTm1nkV+SY+nGIOl9NJB45i2aPXRIF1EUw8BVSxlmf0yhc1wtE1mII216rOsQuz4YHDH1iA7q
h3ozBbo6xfsaQ05qieyE3KprZDdCk2eG2wRVD5fV9wJvr0VXDXDpb6kQm3hlGDgCX4yzHzgbNK7j
msqbLOYd7HfONYjiAU8Z/IDeaE0vYuBi7eRtt8ruM5k8sh4YHJ8NfANNszZENkppLIfAfOWU9tYB
5jGDpB3XnJ3hDyDmV7XBscM8tbz3GL1BJUbbqG2aD9K9a/hvRT3S4xtrvEpHWiOn9j5fstmSHGP2
FWT16Uir9terGiVt8W8Zqe5OXsoXRqcepqpqqJauQY2ubDxQvmA8QfiGQR+MPREiRcT27sWOAEmr
/Gfas4bnZfKV1zzNeJJu/l99i5hlYnyhXtl/V8SPBHm1YZkeTkx8uiDnr+fL7njwpPeameRj/i6P
WRqJKUzaGLXQR51W6kKlVv23k9PPIl1gp0crDLByeGd7nuSL9u4BdGIllGjfmf7m3y66XVOzoUR3
p83ILQv0VjydjYWSBZIelsf+OkkLvIw5QiOrhewWIkbNXlMBP4r6JE0XzUxgH9KGYGHu2SC0VL28
4kULb1mLOcztl27GzmnWryIky7VCwcWUd8jIa18Lj69Op/5IVzbJmPPLBEzDuAke0r+wTh6PC0qZ
2/UkCUxtfvbJxonvfAAqo1u8JOBYCLRbBfO0q0bxLYxnr4u4TtVnQhL+NT02GDsm757YHTPKDWAV
K0MogM53CzEqe747xUcF912JEF+tP4Oal0QHu1VoPDB8M/PrRr6rxHXrNSiDM3XGOATNhmxtTwtS
6K9Nnurqi7F+soC4WTruY0Dir+WztDD6NzpYMrou2o7fyEAB44XTfeggPBxqyKVffO4wVKVG74fm
2GK+2IGmrBv1af5Mq5tytLxHXV1imp9WaQYEhxF90DktugXID49Cmnv/UXMcf/jpUDvaDnvY3RWm
6DHTZCFvdoipJ+3vy9gfom8WJEKFGn2Sbthb5RgvlldV5dSHSJwZNB01BOdP/hFSPElJAuqFRH8w
YPcCbrZ68EklwMTb19ny0O8F94/Kpjm1QlUIFiWP/uUs/YVUbnmYjGaiYbQfNVMUIFiPDwtKgUEc
MHPrg2F/mQEnuYVSKM09C9efMQvHvkbqmIBaKn0lyAlISUPrZmosa9ZsC2IuGDUgP3eB7nR98ffH
m7f3IeZFzhu4Wa8GFWCHlmSVgnlyBjedQ/wSopnXV7r4bn/LJLPfyGu5jz01F7y0iEhLidM+PCYu
CwAkkbJXu4FvvOUIirra6tqCcWKyOWb4J7GT/BayaOAWDhf8KZVKN0fuhR/bm1mycXqnot5ccP1f
wjjtHkKAvYWCLmIYrtQ4ToxM4PhFXePE8V2X0iflvfSvHNlvv1GnfaniCM1+2H9Z+Xov+v31AEGX
s17NMi5EixS5HhB6S514V3AbwAxpEJz/j5kQWxOKVSSIACjI067QfQ98dtMAPKqqE0OZ0ykVvMS5
JHkXumY4WOdFRCIOayY4wwdp3KVUc27ZJXPYPt7aVcbW4zZCXG6xKxU/qgqD/JEAMWPxsm6XuhoK
X6KRnXkVYrJ3r5wgqXOOtPumuTnoCj9Ay4bVOIxRHFMiVuICoxJ4kydUdN3CHaxE/aO4VR7oiyRL
VY6HrH16h0jvDC+nVieaUf77tox1VvYztJ5U6/7BIvLjm8d+k0dY5GRuWaajOcgKut/71r4Yady1
yFU94L338Eljl5rgwjdOZJvYQh3BGbLUTkbK7Dq5mCO7Gfqefx34URqNJGIKC/Zt66CZ71CuHXoL
RWDJ+R2IvgEIVdo8HaQOn7An7KPK0Bzrbjv3/phUzJUNgWCvloo+DcdAW4946f6CUiuoozDUX6Z9
Oyy9oSYFNfZP41hKTSZE06YmcOwzOB+pyGQ3YS0qKDHrT06TWWZDW+NIFwWK0+Bgn9td96qQx2nu
eOGFI4hM0SJvmkogva7E49ehnfdqKcT3UnqABWoQg+JyvsuAoT6FmGSV8cxGeU2DTNcwJbHzB7os
suup3xTMf9WdBUG1EuQTFBr0o59r1GzyyGzl08f/SaqDMfd0gZBvxckVySSOCVaLpMKvKNfho4NQ
/kE763urupVfLRPfhZrdciuoq3ojjg1ecGTFpX2DqeFyP8BUPQSiJs4DoPa8EJ23Tu2n4ZYbtwEW
BV9rjVKmwMcMCHa++LBe0V6sbNaoyLVZ/y+ozhGjw7dX/CpF++0uWFo3nM7jZ0khDwL4Ui7ZH7Ov
XePj0E6XnEvce4sAavhTg08+Q5z5NmTsCX+h7ds/2qak4Ir+0ICjc2bYKejR3BJ9n0xA118KwpqA
L67yyyesc3TMMdKgCSV0aUOIt3QdCXeJYYldr/RGeQlUKjVC1q473xfCVu3JQCBKTv4+DVUd/Klt
YrOg7LkK9VqZpbKEB6fVpVsmEsU3CEULdHbAxxjOGOAD4pIHm0tXdTYNEOYUOszmXfrZ8tbFD5Kj
2EqMxPStOL6ccjxtV/AQ5GDGkOGmSJ25+Lf//WP4VKT5Uub0dfqeIDPYCCXFNu1mNfcpa3evcQxa
Q8w1Jya7LfRF7rANdh4/3m3VilE+tPq5VpnDvZ0UFH0RUThO9Nt09jJOADByW6E6O5GLweheToye
/y3mmrDR/tEM2tVQ8zYWX5jZUg+DPZuU86KnklM7mumfpokbEuDGlBFi2Zl6QP87Ks75PGP8vp0U
gZpIDrV7DNCL6xZYjKfqo0bcgM8ii2/cWN+iKKXexuCLL061npVxOZAbc1+kNuINgPYD/nKAvpTD
E6v425A/aH361Gs1NPMvx+zGzpL5VAlL5mlnyIwNOVGCQt/1saibRYMrHy4sWvGA+0ngKYOdwDeO
z96WZvJYNCEwePJ/q2Fb7YAmsw9ypr5EDCOKUzDxDemlonYWd5QjlvnDVC3AvniXqmFFYmmqzV3t
m+mvRdi9v6wcHV+8IuvRQdZ/KPlXv3cVSvL0UtEHY2nQ4tHy/L8PghIztEZmkyuqrm5rlS5LIFyT
ftU41hHG8MPmJKOKKbhrUar25FFx8BxRmDKU938FzJyZTP1MQmEl2/gRMx1RqTohcP6Ox91LeaFV
DycvHPebmB9jt18Le0Iv6Djrac8KJkgi4uxf0qbjWveokwlKo1NKh/Y/CkEyAcnLQybbbT/QOPKZ
L8NCis9K6tKH+At+aZa085gZ81/TVICEzsdKsf3jcuNA1hN0JCg9kBO2inQB3BYfaMDA3EP4ggDn
RoQCygc9D1yJ5kijn1sGtnTL6QqpQI6oNrCr2dW8k5zOMrwBiT8tdAUWPG53B+v5Nv4FMgpbxduu
Sp61WE2hCWd8zrMoNAfeHvJQvq7MqpVafRAI5br0keS6mDLdHV3bFT4Lp6BA3mc4YeF687zm3CTo
dMoZE26+cI0Odv6MDo2Jn1CKflXAZmlA3/Ft2ee8BBQDx3tzxWGm3kH93DjUJeZrcwPH36Ss62BF
/0+zrUuBLG/TbY/PCVeEkar8bTWDOvToD4785tlvv05Jtff7sHrm5k9x59lhaiSrLKL9P9uDCdKF
fOigKmrs38+njG76R6K+9w28n0f3ucxsWNnb/y859ocpJIXZ6rd9uuSrt/RdkYs2MuQU2AUQpuLU
c1ixrJaEPH0sVuP9Z0NxRcuhFexNsqXIyJnoPvW+xKzTpx3gJAMjBIIfHvassJBJC3l6TyfJpm+j
+f3MNTgU3OLOTz9RYtgc55B67maIEqietIY+MV9UU38LUd2uHm68trEwIIst2sQzfPiT+5aP7P5l
XgdKlfDVzLRIMWEB+qhcgXIfsKxbcpQm5BdusZ9oW0ntL/vEPl3qdWYEqdk1/EN7AoP9JkQdhqFS
Mp/8mmjyqIjp5IhJ4eh2o1V3OjVzhb+VnJTqNRJlOww+PqGZKYpbr8uldJ7ink2Tmvv8zEVY2hb8
YLcQhsMFP4R79g2FrZ8hxKgI55qbASNa5At+sSgoGJ2Nt7eXjhDgqY3fPuuGqorGDzzVripLecdQ
s4/VufwQJjDuUBGF+cpr01nNUiSaghmAfbpuN/6DPRd+UcFz34uOLN2KDCSLmvsfCXJvBiYZ0maJ
X8fkBc2xJSy6p86RROOITRimG23cdvxFAkck3SB97zN12FnR40kzaWybQhkX6WTKNhgbtWuL9nHf
J4VVpkVJ1pFdniUxUV0Cver+Vvhs0st4ERyjtRhld1ZFRo87Y83psehq8tftU6y9Fj69sFVMnkyx
Fi9k+yvaAHWZWK51CyBqaojPNNuAvf1GiqG4BCtJwjqvHLb+cYYZH61pWcejzgzV2GoOKDI8JMCu
8MMq+LlC22kjgjD5f49fjevLpwpGF+3ynfYs/8weSkZhXAzuzWOcMyeOzvpwJDOh29d9uwrBbLrz
VhCh+xJNJoDbr43uimV6k0wl2b5bde2nIachhQU5wYHFgzxxb9Z++Xaky3zeOwidf7W2wTuEnUv1
zaZOwSUxXLZAdolUrF2sI5VZwNWCB6CQ1oQFXLaqNTEIM2oHORmxUPadxWDtQagWVMr9agi5t64+
NuDpeIij8svxSm4dSOonVHwrj/iTGEc4npCDpIsEcsQbg8exW4Vso42FFMqDlyHzQQwj/wWoh4CS
ooSO3Yo+98IoWPhpUOk7i/SSIPmVzGV8uU9HphvbKc19WfiWtW7Jx9hsp5WwEdC5juqr5KDg8g+i
SMzflVYahTJ2RSoo1FnzhVNi7Gf7FOVU9E0PrBVy/Yb632ekzEHUGO4UbFFtUDsT5rt3XvIRbWrH
BKHg0OkvJM9+JfTnqZ563jPk3Qyfr7aqloktlLLDA/7VXTm7wa1e0hBfFOMfgFhuIoaLa+T00w22
SYNPPmsXsMPkizthxWndU/1GIwlC1oxTxp1DoFsikz9/s5vJrvXjyYaPXRdEK5X+YSEOKs8sntgt
QEyivNBLk5KroGlhFwD3ALTxWYtitJq+zT0gK5xcoJFC4zQyD3zlX+8KCIWsNy6Jzzc52nvZxYGa
fyXxDPIzsYprHspc4B+9r56gCfErQeyUNPp0YrFF4Lyd4/H/6xFroQvwFvWRNtL0Q1RF9ZyOgJCJ
LVlxlDFhGRyYAXuuLjbtl/Yx2mWIFcBrt1No5nAFloGW/Y+PHl9r5Oh51wyqX3DJ2kjco1/G10JF
09DT+jT2OuuY3v+8cVJJMlesV8P+GkiafeKis12I9+NkVuungoyOh9XQuTynsX7WNMJwG36GDLyl
bjFgzPOyWiC76dYAw7Ju9aPXIKNAEXXLltwDOe4rGikFDNKny5pq4NmY018GwWcOweBOhWgaXYW3
3mCveaueax0tqTXAH1J7a+vCFNCqUS48SmXqZiDOihkjOWLIBICdN7yyN8aei/hSxraZBUGj6hmq
Ahm2CeFKnd0r9tz84Nv/qgd4UC4n+O+ONRcg1HUE+YtHEg0jrb5p9tPJHLjABfp0hfv4u6tSTJ8Q
q14a3jdbisv8nswJ3tWmAyFZf2kweVZJHZfqkin0M44dhEFfvWUIJCDcl5Ys+slkJcU6mr41nj4V
iboMznErjCqqLeoYPNmje9ReefhaciZ4XBTy8MwJ1J1DpEuR3KstNOsiFkAhbirqUpfsSXxzBrVs
a5oCTI207dwaRUZPWOQUXJYM+ZEvNVV4D0+oJy7l1XWn194lS73Z5+vRQ5/w6fZW8D+bY+VzeQDG
pziIxbim3xEXI267WDaTiTGQYvLqwh8/g2tk1E+YWaSar5Xb+GqBvmpz+uBdG5FmmU3kRZgeIosl
wAWoF7lWA+UsaNGbT8GlbdAqhOAgfOebDI9PxCdyjaM9UJPUTiBlCQgv8jtLPgUIthsJop0efXHJ
ilp63cYG73PH+5tYT14E0X1XQex65QFTYgNof0vM/z4DdxDFclSxiVg+ZBK8KaoBCgzCy/uhD1Kk
Kif7rZYzYlgk3NU7SkDOsxKFOxsoTWqTY90Zx9a/pIte+tE+e6J/1W7/2bS+C8h5BzSsgnlRfnlj
S2OkBqzUFo7Y4Xk5JPEfIzipM02TWTFBFGHvWgGxuvcA5vfOk44WAGQ06RAGc88ZM+DOyafu5cNN
k3qTr0XLE5YbPls+GAMfnA0dYpuT5pa+t7nOharunBdIPRJm3HMyDXWerucy5s6QiPdlAPtCHFg6
AhrHfpVH1OutTscfwDbwMnk6p1vAfpc5Tru93Z8cviLWfDRgQ/m771AHWjUv09LMyyDi2qXeHQi3
XRS4dJ3B8gJi/IaTwgbAXdEqeJIOGUXBE5TayWw23O6xQAzDgtPMQO4yjNDUj0JEnSVk/2uqaSzf
DJ58rnFJ0vRDCCXe1NpRSftmkyVVibD9VJfyGm68gsUqN//aqK+XUhLiQZHyrXk3DT156+eFOtiY
Vq24KIKqxaw0Dw0e+n4gLjUKbMg6BPg/qpvYx11Me0nt4+6795gvVo53Cac0oamOradk1k244Jc+
i9jAmIPaIaUdJpcpS5pV7BS4Vz5iKHVZZ07E2yvyJBKSg0HEyHNN/ujHqpAFIo4F4e/C+QGYOZC2
+mc++uco0BlC3BV9sugd2g0CEUp5roVDu5/nPklcDIxok53hPS5TiSisWgIbC0D1tpUiUn2g86UA
FUXTuR+HqEqoN6KkNIhjVoYortEYkaVNjTSGNtTUR2rKuT187DFJ6CzJgjEWEyue5YzSNHV23rEe
UssWZA3wVZALbTi5MKzl/485EO/tV12QveTbbi5l+DHJnJKO3ozYYfSfZI1aGdK+XjRR/QZf3qNp
nKIuuW4YfMXAxX49Vwxky/r3rjPCi5GfhzKe839peGMnkXyc2GDTBkha+4BJf7ZM8IcMMmOgyb2L
v53eiEHstGK/2V1BfIWMWNFlnOk5+0pzCL4xd/IitqyHEz+r5ObTahm+sHbzAwP8p7OMqmUXDDws
vLzgV0PDO6CadMCUColmQCiOKIZfXUZZ4qzuQb+bZ8gVXy/uPAmPlgWJg9wNwvZL1A1iDFANVyyn
cGpX30HYpRdK0awXCq5CkMDt7L7+J7m6DjehUmU+XrIOscYQEmO4z9edEo1DXWtdXjU/TDbnMfPx
zAbqeIFN6Z4VubY3ScywkLSNAyn8tQYAj7flis0vG9STgjNvZG5X4c7MNNt8NW6tmXTPiuvNc2xA
P3hI97uy+b2LtTbYfJD0ZLbE1t9cuYXTaRIuhznP7VFN6KDyE/6AqkbfwlIDeDtM7kzpBhWyknw8
epRrf6eSuah9Pw/4hsnyIYn4Hq/S5tbG+tU40iMQHYHs1Xu/32EzBSS1dRz6ojGYbBIBNoAkMg+Q
WcnkN8PeAb8NwO8Km9j/Vs9AH+fpfMa55smHVioj1uvtrEhtDe/5AEQU4M7nK9V7qtfe5C79N/oX
AqBcLm86HM8zxal13UXkF865egNrs9OIfYGSVsDKbzVdx/vcPMqrfBa+OzGj2dNBCaRThNzm7HYw
HBVs25EQ3FHmBqhwowBc6fgTnfWvDxu1C9lYl9nRzM0uQfodlpO8og64WBwdHdgpeTD+BNqdowj9
tlIrwQs23PX5sosiE52k4TUqJR7VkHTRKupZxDC5BE7+hIGKMzg2EDp7jyKYB1eIFOAXkbbQmw6E
ZrbJ8FCD+WG22ptMK+G1DygwszsZ6DwMtG7+u3LVRdAv/8yxdCu8tgACYA49GdAnjpzrWd8INh4O
GtlgjHJ4F4dVLLwx54Whn6Sh6mAttPzcHZiLCia9KG1cd1nQiCMyvaMqQ5T66U/4nN3yLuoPlqN9
EFp9fbbXw/no7cyIcQqBGYli6jcXODRpsOXYEtWZm9tYWH2Q/oCaBJqRSPA2zUMvaCWVpEHXBXV3
zjwalNHgwDqZX1nZflrEdVRe8ESPsb+VC/hYJPjSHxZMiC4GJFowia6NG8oUFrbljat+uCPP4XPv
odBGa/okvhGMGLax9CP+5vmJQdV5bfSdOT9EnvQpVBY/HYVpKCk8dMMJeULkTkr0OvbG8bklDA3x
voRKLtiRQ2iHB7lpNoDbogDiR7wz8HrBzI1E6pJv7zIm0K2Agm5hHX6aV45I+G3lujAUcgKi1sDv
M/5SaLcpQYZ25X3Wabl6SvbdEGI+jnVq8YHqMYR4thlqRZTP//L+ZwNs0oAWgETja9GqQw3ufV9Q
/Eh9ai5iYtBoNLvndIOo+Jbsnwi6k5MQxe7msbtmqrHY2k4gqcIv8qo/rnRzQCMyarCoJzUHVNPa
xul3g1RK088ubD1b+QHa3LOh3h2m1EzCCr3gZInDqSzReDEt1feh0rTlpwkz31Z1NdtrTL7dWaBC
Mwmq1YBjPSa9cpnsKB6gzKuatD7t2fPKTPAOrqFopRhxLFy0fg3CjRrs2to1GfrNKTdQYtkknG1P
X2XtqCURxsRIVmGFcenVNvPTr7QCuDZ0xEeKlXeKL9Pz/qkbfVoyl70srORRojEIzHsVjlRRa52o
2RAsF/+R2Rrlpxzcrx7UXzVc3HRqCdEEiG/ZqHkEMygDLk1ENhWgiIvRXZfPvgC8FtEodvkPYiQf
5aHljqEK6OIOEsGAfi0vlQ5ZBkAxAxnSLkTHZDuiRqWegXw8vUisRPyROwR5BRA5Y7L/u1CbO+4X
WBils9BYYztiH7mCrR9+KIxC0ukELfYLIGCmGk6h+mjkaie3NFaYb3b3sns47aZWZArQCTwV8rlE
ygI54vXj5Iip65PEqv9mk2CmFU/2kQOvDVlkSEXsWtOPLHQ9vXxoIPcghKXYe3QUfI4bvU9zYEeY
+MRthtyMKc+iQ7qzXfmAlftZrL2VIU17A/xAGidVFfqe/xw0qmkiPC108OSHlgC2ZcSY/GLP60QM
rB/lXTAMRCpnuRhiExAIpqiJxRxmZz4RU9Wugi6hSFt67Gb6B1Aa3lVAK5Sf6w+Rui8es8cWHLDa
+etCUX+swEhl8cHdhqKhB2zFQvr3Pagi61samil1lEV8LReMAOGeYc2FZD7H+ka3J+p+QbIjJ7fn
q01zAmatY+RukhIDklHr4YuMxXTGHbNYQEkxhHElc3x1d4EU/e+DmZrzD1hWxjdzMUCuqNYL3wah
qAMjp9CTtRE5hNMJrqDFTXxKA+N6NPnn6KJySYX2vABTtt/Txe9ctcAXREZGgSgeObxdekVrruok
vK9v6mvp1w/azZswUjw2/IYbMF1cyHO0m2yO5TGCpTEPHmX5vrm0swlIXDItsdLhuP2NGzWsMX14
lLwS4V+S6pr7HyBka+3y5TbpB12U7L/225k938sNnoowwZR/44h6IxUEzU2N9dbn3PH9vsJSkHso
dpe1ZFufiZTjmQRimHpfrUDRK/Qy4e/yOzGXXrYNBbePd/eaYJGhzKMWJUN/eDZusavCk8+k6CmW
DqqyMFFpAyoEsI8OPtofjqapSiHuspHftAhtERiqlfyBp3PhcGVkSgYc2tRUhrDE4Zv1fqrBAzea
4+DtUB9Ore2gzvpvstGWXTRCR1ZsxRHFfBtvL2Euzri4VMp0jj3HuG50aq6oK5bxdNJaaX1HlmPe
/zY90ubtdn9KsU1tRZ26GGCMfUsXo3fPIxqXktGbz+elC/fM+n9D3gctyehekG8iu1mtwxxMnemZ
Oyko/pZ5Tuv9jqv/iH8jdKiD2NaKDNCe98FAQrU2oDPWdvRDZRBDFfxBU5jhCPIMSWI7iUepjqcy
Zn59r+dKs8guGMrNbViUIJXmGt/vncdk2dbAKke+566ML6HoNlUvoV5H1IeVBRy2qFbHcKT5vq7x
cCSQ133CDERVaGhpfIeuVU1kEB/ciF7JGttIqil+CwuFsNn83LOH3sQIUR23qVGTMqphsmWEwdDa
d0gogzDw/dQ7aBPB4uEWP9hVCg24sUNTGq6r+oQyDacRJGnPU+HibYq1ht1baGdg6wgRMUrk1wcV
G5gjYH3RNTmc1G8kJCfInUmJ6/L7zijOI3CTBjx00bvGWI1cLb3hqcfGMXPEtv7wK5lfMkxQvPUu
ON5ZkbJv2pQ4cgURwOdwULU3cyhrcfN1sZ6i64VjxVnbrH1rC/dVerFf2Bl1F4ZY+Z44IONDt+C5
qk5psKP6TAQKSeuejwhNhINwqvSMJdz4hnW9xI725tGT30Xiqooq3jBmvQDgWnza/zAbvdJyQHKT
REMH0/LgrK4Zn9Jc/OL6FsBYeXM8DaUuXRovKpcgzK/ex62sYnVE7OLDm9aTCT1EI6fzw6XE3HLe
Mpim2WJbhJBpsDetY7D3MfbMX5zEpVktHHWr0VwKsv8zHqzeGhWtzUasPqwPIAwCyN38+OVBk/mq
DpcqDCQ8hpPjnQYWyHW+Ee3PT8K4aSCoAYY3bmLcp1RcSuYb0DzStk64zNQgJYS3p5XXZPGFpTfo
RHpLZiohJCZMK/Ctmxx6otedRZSReNoHnIwRmURvvfVjw93XaBEz9Aq32aQDPz65Yt2iOuxsMnpb
L/QgUXZE567Hh1c3wjdXPGw+vDrWntd2/cx/F9Nm4mDycC5Z0bbReWiXvC9BqyudX1ARpT8z9n6t
NtsCJnJHFx/HAY93jeT67k3+cqVwpTCgo3GcFjFjE5fp2OBODiTnwp4o/M4F6dXTgMbPOS+96wVx
vpIBrJMTLoFR+o6IUk03tU0J+CpzkK4+6hdEX25JCmzI/pgJK2Rq191EOAOSTi3Z4dzxUArFWwJb
bXnPQztPxyaPzaGTfYDctrWCQO+K79i8tFWBHPU/5M5WdO93KmlRT5iTUtx1wo5rBsVuyVGoQoCT
T8AXQDsac4oFpv8yDmUxhAz0Ttkom90M9D0bKEFjjvSlr4dKAJkynmSwoWfxcutp+l2HbQ8HAabN
T/o3cmYJlhPgbOnZrUhE5YWsOthe71MKGqh4FHRc1EtZfoPepDjm9hnTfRK6lywcLoXrs0vcfNyS
B+ShOfyESQ3wSLG0DthXkDRoRFTeWx6Qaewck/2kjKIp4QlBdDcb+rkOblkuHRf1sfVdHIEo1zjV
p6nkgapSc/yPHHkVljrXRE3iKLqSSMRG8kQ5wVjlJdS2aDaCLfi0649asWDGrcx6Ps4Mu21ZccmC
o8SxDO/fPWEPV5/70cqVv4qg5TGy/7hGU14bHtyBmEDnh/lM42iEOqj5xqEmEAHZ5xAh/Kdna/eH
0rfJzRpIcsy3lkN8abP3f8SSVbXoLA35qbsjpNOMuCDQUvJdhGp5rHsCmOHAQTQj/yw6NPtamffz
dhqA/1Pk7Nwjjy938ZcE3eNCBuaV2FXneIgyxm9PUwp1fEU4bBwxY4FISv7znd+gEmnrfcy3DPkk
gPftMOPrQye3xwh6GYFTKMkj634nKYwpoFmEvuO3btOuGbpfqMbBRxiy8DFgM7mM3OwC1UwsBF0p
Kp3w78Ncbo1oo6b0PAgv26L7FQUE1q6OJiDmvuUsu4vt7gDYOmI/5UfsTRPDhNuQG27vCNp2bEKP
MTmUf42gTQvgIlCCVgazo+QoRutmq3Bi34pA1XRdYFx2aqx2ZYpdQS4U3JmqjcL2RdxayQ7hLEad
0HWvJb3yzWcr9I/MEupcCIra5Hy4f7NefLh1yrWxWHkBIWsGzclPlZpTupALShKXXSZHEqeTIiwu
QBnBIZOzzgF8QDvDaTDlze7cNPtK07RQ2SFT8Ow2yKicMzMhzsAClp5ZLTXjQ3WCM3lPNb7a5tw2
65RJtVa/F3uXISf7XQUSl8PxmiDKvhVf8qyUZL1cUGOFdujY3bugnTQWLGXr85wvZ/5Jo80Ohou/
vkFaa6h2RPtRIGmeh4TF5MFR2CnACaNibBTNA0FbGJ5bHFKflVXgFK8+onne0tdqAHHSjJ3WDNwn
DXdvLem35duoflOkbJs/MYhNeomU57Ks8CvJtDBxraap8jZoQHlSXUPy84Zqo8I05euwvtX8j3l3
ioI0qWZnjwpukjTbksWP/w/35M8Ir0SQbruIVXjuekSTwXySeEqOql0FvhOnV+/liQQKZ4RtLrpX
7Y9nHqapbbVFDNcRsQMxc816G43PsjXVFnux6yvRZBrx1zxomszqsSlLusca82UPj5Q5d/rL9bVU
Q8fYkMbxyJDCiNjLuOeVuiVhHBTvDu6arXhosefeY1c1WnRW9nXvP6RjHKfGvbf9aIY2qSa2gsQH
Tr+6t5OGswVkly7BN4+FV2e8LWlnqw3bndk5zbaARJkKGjwJ4fjPPIUoiDBRyBxKp+rj3P7JczEG
i7Ch9RPnJ4qdTQ+/TnSh4pnQ8NJLteBAVEz4O77EnUOj6NVtdLQJl0BSI6dHV+OjBL9OHFIr8qeH
cW15kJ2n5IsLWR18PeV+xlOs4gnLhPJierz2b9bfW169iqV4issTD52npcPSrVax4Afh7s1DApgb
F5X/ZdCqc0+8zShCYBTdwc8PMk8xlXExNwOQuFpDMPBqstJ5pyxZHgxOlYCIh5GxVQneXWR0ZODP
2/YPc27ZHRzdH+MubZ+N8d8BtWV6wA3HmaQnRK98dsJLURWaPPttKt7QEL/AgjOP0lKVlksOOlsw
G2Qv9OOafibDglJxvDIyISWZzm1QCod/XbhjO6N8RyUnmzijJsQUjM3xYaXLgp4PuHF/UadZ0WsL
hcXMpJmHL0njIZy4D1zQ+wDLYPoKgAcpBt/o/CJNprl80+ef2dCVks9dQQPebtnECdC84ySByAD4
iN0AmjF4NMrGfcx926ZNiDBYYmbnO3JaXt1m+eYdBUfAiYL8h3oh3YBYsGjrzysF01k/NKSrxhoj
qUBW+gpNAuxsK0NyFgWaUoTF9mCbXhnGiTg3QEiITrsCD33kMunb1x8RJ7I9OjpJEdgrHBDDyut6
f0iZKDtnLdEmBHK46DXWIzXxQ3XsCVI1BVctTS13frY7qGny3BasmiNzpyXTkv0lw3YNOfqmmGoA
2Mhdv/8e0wltDhB4mGAAoj8BHAydkc4IzEVDQRN76p7eYGCZRzaRshXcJ+3YtG5/KOi5AFIvWQKx
QHsCoW0M/SdIJG4OJvetHDhC8qW/W8wd0aluKaSiU4tmv6liYGPgtfPWtdPFaidtOQMSUR4CzIMC
YvDXcvorRp5xL+yQxwSTIsMcX0HYw5fH709R/w5piVtQM4nuqu2sS2axT1DVrnsdAbQrDcBoxjCb
0YBc8X1ZEB3w15seekV4Xu39DRA6SSFx9trypvwS8wqjZR5WGh5V2gwy6WCK52yPRE13cVRR0UMu
t1KNG3X9ukENXqOkths+gYGF4NQlid1j9bTRpIfXYp3jH08QZ7aQdgwsyFSzE9K7FtXuioMoPuD8
2Y8HfeTlQn4YxGcwVJkokqKjSCjPYsK0bwrfFAfkRXfa4AWFuk5Fh6HZYFJhQa1pqhQiodZ0ZbzQ
kV0VlpQU64bKGY6P7450ACsF7CHFc0B1wIc3SO/rgZKOsmWPVMggDnzRw7v3G8CMpFS+dWNV8TTH
R4mKhlJXf6dlBtbM2jlOfQ4x6x4/9DE1uoxjXByCoviuw1Ku4G4/RU/LrOWiXYS7YDkfHECeAe51
hsB2XjYqVhLqTS8gxRUCbMxzw8P2VWBs6W01H/2ED9SN25P+/HHTtbzMWV1mbnbcnrNqmEauyvsy
apQqWfMMCo2mf3rLli2aI7JKPc5z5MgC/VlhfXVFrY66c3z64Ez2Nc2Zp8QOLQCMWJHKz2mUsP0p
VEVrx0yzxCPKf9VaAmfP/8bRVQFcA/Pyky0MZ5x4qWg2VO5iM4ELCESwsX4AFJszrM887d4FfA6V
31iVANvV/0z7o117Js8qNh/eyIs/l/u00jTz+VrpwiHdPSiUC9qdDxdP70VQanZCS1kWaUzq0lNG
ut2xa8G8Gr7F2HQbx2KWjYywtG/WN2bKbRSkjFF7yWv9OuXKWIfGowmGyGgmUOXsLpB7rwasLxQF
PFwwP6Z5IMSFXnYn19bEJ5DeyXavxwJ01ZsIROOTejROYaexnnbQ/z9k5pWkoNFiutW7Fe1fHrNE
mbFj41VOKA3OCYhd2M7l6xMQO6qZyBuG58xopwZSbi9Emh3HR0kOehPtwyAcmSGGO6nH37ba5c5X
BuPfyreiKvOZ40ywS4xvXI+oV0U04eziLRX1wAgiKydEmrhBf0aLSz+RphWVO6lftVBAbUsTE7YT
9cigBbsGOXewGpy1yoUwxEQtNz1LSftRfa6mRCBDuAqYGKA4P25RO44Y9BoIbOzOucmhQ5IPwd0n
q7a7jqjN6wwdVhHXHpMpuunzd4Dif68TNEouwkB7hplbFmgykhHG5a0ysI+Q50JGyP8aZZGWlEER
ZwCEfvqxS5AYtq9WueU46ZlV6BSDV2A9VO504IU1YnlkS+JsqdT3Ijr5ZbJz+mrysD4awwxZ9DS/
o7Vhb4eU94NvYbJZfHue/aG8/SQTf0PU8ZWTfxRUNKpYMLbTDD6mcA9JJRNPRtOGrYIEV0zJnQPw
Q084gNsJhP121BGGiAbpNdPdNDjUV962Uq5DtzrBd+Fa4AU2upa5Z1HN+vTEvBudMdYIJSE1Qg7B
7lWjIaSuPWQFprOaBSIgbRNA9D7tOZL38xmt2ezT6pgaVNnWvCpYJTOgy+u5fKZccSWnOtd7tJAZ
FZij5L36L2vlj5IUXvq0dKjUlsWW11JOJrHrOaefeY15GX80oflL/36uf4KKKJSTWXGoJx2HeaFd
PquN9DIaAiDzXY67eLcWEPMBzA7jY3BmL3K96DWM9AfMxEwKKKTx/QaEALJbJFExuWowvSYFDZpq
fyEh9hcJC34TtM+tOVE2xFW4se31x4S7YH74pECLvQLU14SoBypqvWcBFReiLWUPea0azH/O+aVB
q03VsmFx11L90gXY/m3dClvtWYGYY7/QlDGVukd7HZaqN6UFnbQLXNciYda+NeMihfDSGljbq4HW
evJS2XRDultDr1tTfTXxip8Nu4ntAyJur02lMV+upQU0HzgGPOElDvVCzOx4OrimvGE4LlBPehV2
C289ddRCEphCvMdlIZ5CIF8aLGxFrFnAB+Gk9qKbz/pF63CcnQSEnpX+bjYdTJiAbWcoSlv7SHSO
Fdaxomp4Uf8SE4sHFENhNRl59QWv5WQWAelGCmjpALNjRcmpWZSoKWnceUavYcrdtOoKtE+3nHUg
64ZNFX0MHpEmaY8DnObSgmGog+A1auPhBFERcZHWdB3IPCdDr0LGaLB8k5vCveFcqHKoWGhXHavG
mIuc7rUSf58DmjVCWWWK6w7v3F6Z1KFlr1nRoLK9L6seH4Ukfa5Eiq7HfGLde2SLPLPtWUbH11cH
uRlGHdlNZbgNZoi2DVwlIM0zA8aaqW9EYLCovYnFEdwG6/R8QqQlpc1Hw10Fz6TyGwAPXpXLHG5q
+Ki+zydaX6xnI27h633jD6WCzMKVTDd1PFy19L5ICgyC1Zu+EnXbzAPH05d9hPuqokhJoTHCiUMe
AwDbFTbYLfBNvZsk6jlEZhFndWrD4RzFYjdl8X7ASGlFSlGSZ6f1f8KUTPq0+gvlR3x0z6aUL1zh
CZAGtGlUVA2BK8jhaOhUxLskYYBv8w1Nb8vNg3c0Yeyg9U3JNpslEUS3grukiG1kOzKPsC+avttX
54f2fhuh5uWLQJ0Iki9THxishiur+6pJl1y/4EC0yJOPCjHcd2Xu59kTjdO0Tyvy7qkcfAsDdLyc
kmoRBlW8sZuSZhCrTRu5yn5fMb+v+4km9LF45vc6G+o1Z/ErEP+Yk4boi70Vw2hP5vDJ6efy/J6O
K72YNNt9FgEAZPBbkERIhUB+/4UsmBdbwNWLoQNKEOtFq416kBpBfIi+1jXie66NfJ+TEZ7la9GG
EVbJcXewgfftQkdu5vAVvZkgCOsoat7G9anbsa/ZB+Zm00oIuwQ7plRH3keKZm2PDkURGew5Icgf
j46xJBdsHB9yhlxlqdRhKZPRUuM2b+uvzsqpveAuDeZFzGjIoxiCoIgy3TSpeGRW/fVDCrRCCWEr
8AkzFvMB+MeDOmI9F0uYzkEu3yrAYWy3aSHUPUYX/QnSWh9+UJDexiPLgERsFFa0O9tmCxdL59M8
9bCp5YToGuL5kD9X+tzW77U4fRrf36eC4fV9rG2vXvmNcbdvghwE3yTwZfUw9hqqbJqBUFPfM+OH
Z8Ostg6oY5kQHGbditIZBMtdFS1u6uGSxIcfM6BbbzjeUB0+xXdStg/3qsWbKQiJtL0O7mH4Xy0n
N+oy33lFf4554jvF89crJYYHxfSbuuu1HzLmjAsYB2VTnCUVSdBgfZhVaeIu+mHgWeYTR50C1OpM
3uNq7mRdoxvDYRvx4mSJHUdmSc+jrn4wOsgeztB2NiV77fWgENab36ceeajZgkAEkx6qUs+24WuC
jB8DJM3nDpDXnJuGOzz/p2ILRV7dnzG8xG0OiCj5r3sSghuY5w6MbLfG/2UJw67IPf3cNlwJYbJX
UTl2OmjznIh7HFL0VTNO4zZpb9WhyCcS3OcuriB9aXO/QzyfwTYA3nAzrEZFKb1Phq5z1MuJIeQ6
aSQ095A47EK94+LLGR6uumUyITqK1ryx9YznWNNFLCncyTHugMGx3I1RGB5+RaWHCqqXE4KOUVtC
9ZiLCHsUBoD/1wIKOQ5i4TyeZ0v7ACF/3A+CzxRcOg196HnVaGOTNnDFua0h/G5eVNy836h9L2z9
B6D8Vh6zPkv2txOl3cHaLAHef81jSzW19R0FsaB32gjtO4fdatJolaicjiFc3IEcLwTvN6QxXYoL
REy7N8kF1O2+KcC1tkvAuXx9QRZGtjdzqgGlQDW9wPLuxJtH4AYIQxL9wYvlbf26CfT06tJpjlHN
iITiaEM5gqm6/XOfaxMC3BJ2/05tx1nA1bXuIVVgk71DAOa0fZhSi3iTN/iliJMaanOOc6lqtF1a
RXhJUM/XQCLQ2DDNSwGm4dQ29vew38TR9Y+6bT6fiEriSaPScY1srwptoEdbDPTHhSR7qdlUW9SK
6oDqpaLSM6KTCPUaGWLh+4iCTPixsIBxckzmu5Gt7ENrjrIMsRWQsP9KfT4OLo824YYpQ8+xAlbU
YuQ+g53jAdpCNW4hh04EYYhu9Jblkv66/Cn95M4yvJ3bAwxEDjsTlc0ZV37vOrbdzRcjGBADhrxd
lxMq/MDXPhzU+sKYt5JY+T7SsWWNkfg6V5gHgFDe2sa+dJ02nDIRUeDQnCICXteBUiTDZ+kSTRx7
WVMLY4xzah33i8XfHFD2/XlY+Y0pDzYtiL1cG7L4mw9df3rHn9ln+5ioqUxYWzyxsjQYMOoUBaFl
z735vcQs8fxInnNYB3nOqPEHzLUrECSffxu//ICtGXJVAuW6+6rcACf54cF5R2evcyRm1/78F83c
91BgqYfa23mb+IX4OiHGoyqEZVhj2aSk0tsJ23J6AtGv8f0jMetnc8dziIlllvJZ8LRObmi0/9Ia
Ql5je9cCVJZfBlNUNQLGKA8qEF8v6ZVxYtkMN8Dq+Xuf4GforE1iVuTDCG2qZp3/ichqBxU757nz
HyFGMN7cOuMK2eBvV7WJgp/9JI+MSWYtwckedE2NyGTGmeHU/8BerDFZmQxdaSeB5MPdBZdpN7ID
zpZnMoPV63Ax7BGehX8L0N+tZib6SNYUsjsUmiYcUkR3cyJmkeJfg1xnPzIPOA5k0ocbhNUXofzx
1oVSDtMgXGDIod4KScilL8u3A5r3VyPNGz4WqWKFZjMLUSehMS069w9/5meXEBRKm+0FvHgUrO87
OlWFdF7Lo7QLVCNp9cZd1HQOdh5ulUcqh0juQVfq9XYCK8mzJfSkYb+tvpUcS84PmzSefUSeVY2H
zKUFSilqcUtzNaBNde3qM9qtgzKpSCGC3sfcZm70OlnwxjhJtb0AB7CrqV9QBBIUskylteJhPhtL
e2VWDPU/wJllOFy8FCIJRh39gq1H1k6V1n5aTsKEDy427qrrveaGf5dDJr2cwX0zJLTfcQncNZHB
htFzgZAckSj1vXSdjZSyl6n6++qlxpQIIO8DfTb7MI/DF89u83yyPmNtqG15FcyzRON2oUQnE9Dd
H2S3OUngG9CV6zNA0KAwAOeIVXSJSkcmrOvp8CqpgU7l7lgyeMwrl9pjltvwGW3iA+2ZnxxegrvV
+cpMgJEjmor4gTJNpla+BZyGfLVAncm2SDB5jO5SLtdltSr2LFd6AY5IzK1xkSTbZ7qTMu/NR8In
A7bVYyjNUmLQZ+C7D+zghk8d1tjAsG24H0ZkOjPgqyksHa629N9shNoZAyafMVJdskTk2qrS+9dd
k6JsbnEAeeL8yZCnaPVQiHM+wGekd8mLl13PVegrevJaRpE+no9tRGECxF3W1iwYwJzcJ6x7cQEa
uOOgj/IaMjuxsiyTtSLUEbBAFij8QEI97lNVWnir4jMvf4oKLsJoW7Wxbb6WZ+uLqIxJ1hM+7jdc
02dPELAce8JYaNsv8Uj3SYUU6iw9SDH9FgEmS0530zxrFx8K/SshRgDbLnASXet4s46vKEhbmri2
cM6MMbKYjLP+rBOjVdTTIzdCiviWsnnMjJHd9R/lpxi5nqDGun2d5kypmEr1nOngpYx+/gPIGrQy
tI+w4WGD7nczG/dAQCANX/2JQz1jurLkrwpq9/B1Fo4+fIrXvcVUsKp7623bXfydDC2MCO2NohVd
9wfhURb8H5MWmKmXRaJsVkmWyahBQnyAY7xjIh7gbGzenWa1bUIaA/JohkLe+heSha6KwwL9TvPM
V0TzSvBI1YEPtmwfhojiSmrD2DQxxXATVa3qUb2Fps5sRa3dLpNy6bVCoiNuKYwYw/NdPh7CoRXY
ELV8B5pE5RRkfhFjeTSfoKlSHE6/hipBmW/GOJFXjv3si5i0nBDcJYoiyRjqK8FXITIUDoUZblF/
XPLTCnDKkJ2Lw5DEWdbld4ku0Xt7un6fieTVHb2gAbtgrdXc1UvCMVDW4UobNWJy+viPg8td4ogv
RFLdRU+x0+T3wjWiVlO8WQvKMe0g5hJMGE57ZmOCKNfB8xsrDoN6a/50FoSdVNlJsrX13P/5cSlA
clKc19J7bD7yrkOFdp07+Pl+kSN4pgeAF+cCxAsOm53scwSNTgqsriEhvnPAI1zrybc1FbUL0HNr
i2cMeTq/uTq4tVFBYRxjlnNyVdVw3F/QKRKuFaFZHanQN9ryc90wDBcV0p6enAhV6MqCcdAbN98v
rcc3VVWEMVeO/WLt3+iWviCUVpBnIrfS9aOE0790l2hWWkJYkqQMZtMDW7SuJxPu6azAjt7eUdBk
OgAGd6ya/v1Lp95znOvb5eqviZhwgKiMffgwRU9DhTcrwTjtnzMHDxX/WuEYeylFDL1BmbxKNhVy
oMXTVuLdH8n5i7ar2i17gRL8/MXM9ZrKM43qKoqKzohjoLroHs/ofkemzivED9VpsJsH2NS/h67z
L/IyMEsQL6JS/ZTSd/ylPut1jd0QashWPq+6FeQVf6mL2NdLNhI9NdaQPGF60VIh6wCXTku/vx1u
vKw8EqZ78jT8L7/JU+PI8Fl09Ql1ePr+Su74zMpMRWP5xkpwy5qkhWISlR7XKp4S235lyWz6zcuS
mSQJ3VQ/0u4ENdypDh3rYzDC6hH5yJfYKO/NnNAMrzg0TQM1YQu3gvNxYG/UedtI2hOpLhg81R6l
VFzGTI71OLE1iNHVrkaQ/CxAZv73Urzu1pRshd3C97TadK1W7IfsD7Ru9U3ufNp9JtzEYql9wNOz
26RHBMq+ga3NKJsGMoS0thJVlxeJE6TjHra0pI6hT4dVqXZqL+VutFcWiDd/9KbnChlpzFFSPJ5J
mnUvoPeOXyKPAxwYaU1N8p+Senfelywpj1SS8jxkkBqxfkWkil0vZr1b3wJMx3li/PX6uNL0dCeE
JRfS5E7T/rbXrpP6xlnlh1CXC0ul7QxoTObGrc303A23j/mnAJaFBtZdWaoVirBd2SuNmDtiCWYR
535NSWRlY+EFNmtP+UugDzhntugccB5q5MfE0g04s35FUM/D7b/z+W2wwdjGrHg1n/zBm2etRzL7
DY/zi+jjuqWEjRla9CcFe42hMthrBdEuugqx1cP5h2FnMUExwMIoYFa4i+iHtI8Khf3SB1QLQI6i
seucNvzrm8oMWlSYuE+eJB3vDfTnxIpfV/LT1ge/ailkssVqFRXbQh4eOmmyAXh281NEDoxjiEPp
5HdL21f0D1VlsPIls4HlHD0wtSzI5Ye23m94WTWFm6wrHanxlXFBrhBSyQLUf3XY3yZ3+uv0i782
cd3jvsqiO99XDuOVFawtGkIcjvYzTpLH9oaSapqR/4Ilnrb3S6c+TOZuK/L23XDK6U2qrvBmCZj2
tTVMeF3PE+j3ZuQfJzixJsi73QLgsyNB/eG7ovfu3S6mvcXgP5PU/TmMl2IVqCTy1diDVwkf0FoE
fidL5kmMde9iM9qg/e8eywaOdbjD9Sw/lh1fHGC1EMs7mUZ2cUR6y6rCqhaz83LLursnjiFj0G3U
wo6mY5ggv8+l2sRXp5YQrXkzwG3YWqzs6Y58xIHJXJk4QV14Ps4JZGTZ4TtFl7lavMFcOQT0CX0e
92BnPp0b5wTEn4mvvtYvTrRUBjmzNidKwDeHDjGlMDbbdSf4qkFPnPl3j8tz1e8X0mNbsVhwVyZD
RUE8oRja3vz7DR3R98h/eysY1IMyUp+yspsnLV01KxhMy4lEuezGI/X9EsaPJV6xRVoNrtPTQulG
qLboHGpWTJLofb3XW3Gz/UDNzpw/3/ko0ufg5r5OE+y38W0rOfY2nsZCg615v7CbecvkqCcXFpWi
A2GwyNb5DtOB4QK7GqsOd46IHsNLe1+KfeNxxnzToWHI/yqRnQLePr0/PFntlG7qZPzYXVe5Wuk1
aJGVHS/1NzBaAdSAIBjMcbiUJBXwZPvoAmayl360cWMxqafiQSXSWSZ9B/PaNAgGs1c/n414qo5g
LardTCMXeY2+mkMoHdENxWEo940g+ss8ydWO5IyJPVPJXz+S0nJGHi3N4XVIhtRqKuUSJKDQTeU/
lRGfEBM6R25UnUfh+//JDLfj9hrlv2Mv8ElyqFhnf+yaJx1wkH8vdpBGxs3UK83ccJycxY5+JegG
zJiIBMH0LuDIIn5rLMerlLro7Vib2U4ep/ka+NAW+9Z5X2t+etwxZeDztG/cVJ8x7BQ8ubwgs7x0
DNkPL+3hMiYdhzb+/sHUkspzljDBhuR/xGSriNCkK00mpM0HJXA6GUNG5F9ly0cDKe2Cw57148OV
rsdoq1fUG8FGyMhBl3nDsvGURClg3pfCC7B5jCyIkzz/TbxZyklCStQLIO64F0i6nY6+c4U4d4y6
Wh1ssgKbYtl7JbmKeBP9HxJBetAnXh+rVOlsP3VnnAfKkwft/I47DrHoNiCz2Rl1/dfeZ0ki6UgS
cgFbf/rDkpXUqK/J9HWdh2KS6u64iSkDiDHonMEzkW1M1Z4Uyehco13mdaB8hvE7XX6WRrJB7oyU
5R5CEVDw+4vzT1IhQ/K56yoxhuImP4mZjGCGPHgwzBJOcDhitQc9h3pN5LA0t12ZKh8wvIIHFsHS
OfcG1wP8OAhWGtSuF1XIeVaC0mkvOrFjKJ4c2+E89mOGtS2JRg0idbeCqzek2EpjJWIJigYeW9NI
fM1bCLe/4dz+kGCEFUWeMfMaMtY4z9wdKEcOatIiVrsNbpJDTQiK5N+2xehP8ZXI+x5hjg5K8hnw
a3yFKZm5UduD5SN400LZ1DLNwrivvQ46OYGJsnjbtRjzzxhdCmR9IL4KukrG1R2Fn1cjJCBZVMaF
hecG+DYFf4VAUD6Qa7RjgxiAIA0eFL0BmNeMa0y5ECxoGCYl3VpQs7Rfhbrep1ZGAE8cVvUmRY45
yUVQaQVzlFHaMn+J4qroqZBz8Dh4sxuXvJ/IZHZy0dxZtmfEXae6+26D+wPCMt5cBy6DdGKvRBrJ
q/qpE20UGeGTw0j4sufKNj/U+f0zNTu4zmb2iFOlZ38WmYS1W+V3F3tCTNksjvWejr7nSBvao6d/
dAovgAzBGqov1EF7nJhNgZdHDTcA/AF1gE98ByXy5W88TfndMjc+WjFXFCMjfEZbBAVNn4Vx0GK7
UMJqu9ResYxMg2/L08uK7l3L8wOm7/tKPv1Kle93x4BQUe3S3B1YOJT7LOAFySwbUz9WCE47zBT+
PuoI/aQaR9kePPSlupCdGK4lsUKKJGNwa6RYlS+2TAjsbGt6uqgsYv6OLpBcPLmWeuffjN7Sas8P
VMI59oIWbsdWIjmY+FJy+wFu2EUQdxTXI/qiKCWvFFajFv6yCUKZVv79otsyzb0GdnefgK1f+zOI
aI2W8Ri02fAhp6y/z9hsK6fvLMBVwGnX8RxmqgjmMuiOL/Ty8N73cK/niS0CR7yfYseWGm+pjfbL
coVJPXGhwCPgwPXxM3UiZ4evLJX8vCrl7lM1VDC0C5A7yBbJ/EE10v7OGBphGKBVRqnnNxVS/D0u
GynlCoS4ghL3ermOiGF9LWMy0liKi0td6n8TECtI2xhwqrB/bC4B6XJOU8SgQNattPUb+MzLk50k
1aUtiFB7/lZZ8dFiQNXRJ1vEmzX0IxYWg8S6mGJD2kbnIaRwVRInxBdMf8L9QWaGdFEyf2w679c2
ifQI5Vo2DIDFg867y067dj3T59PgWlY0C6R6dVt4ZbRO5q0xnDoHeYH4G9nYY1yuMrYkpTz8R+b0
FaA7gWfjSYq5aIG5vxZ4OWQ8RxhCz2LYmnRd1OvJ7Nd8KcCO07JJYdxyD7gK+1JDKJgx5kHVnGJg
b0lgqr1+R7uwOh+gmrJmqG4BGUOZ2H/LvZHw/xkfQpBrr7wuHm1mUyECQUH2BAJvYx6Dq1uyb651
Q9LyDmCXc1CQxfAO8pib6PceKXVVj1k+v582dCcwOK9j+ZfrqSfKwOcgAzFPRl9g8cgTYq/1nMd3
nvSeqzw/WNem+iV7e2OI7xRBmg+5gLPwqQMQOZQdMMkwQGw/NrOdL+Aa9190lpR6Sex2zhJ1/Jq8
W42x2D4cUlMUC39fHzXT3Nce5nZw36jrMjWzKgDSyKJFyNWMH7OYr3L50r59m7Q5kjgcdWVbMR1g
7TiKwLMMnyGQSDh8a3ssH88hTwNGLN/mvTZzmsi5v3/jGinhqtCcUr4S9U/vzu6JA0wkMxvtSF15
CIsip6AKy9edH+m7CmdH+pHi549DkvLd7H28MenyV3wqRfhVAJ8ECPZtRQnQBuEsG/Vtstc6EuyV
gTUDjtRPqQBBtA/x+S2h0zSMcM+pCseP4ta25Dnf9NrH9Ovp2QQ6WasrNopjntcFzYO+SeJdvAOX
qqCsXNWZ7dx/UCwAzCFtVpH1JYSp/rymFWvLpM0j6zowBBEjs8NOqyoR6U1uoI/+8EcLAmMX0tZ7
3usMtmimx7qqufmOip7Q/cFq1WZyZzW5rTr7I8HHLHGUQa/9wJ2bnnQEAp1oL5N4kpj/e19bbfci
8NvAJNQabgBunsb3Kf2IFeq+UG/Rfobg1ympaJL2r30j3dUjVhRYFUfRJGyewRmXKncK5WTUt6cU
IyzM6iRpDJRpRIcyT6TtFugP5doyRPeKrZefZuUXE+3fCSbPEw9z27rb/b622WJpr6V3N8+CgABE
CTFkIf0X6IrKfoe6Wh9RapbCIn+xRVZkiIpHyPJmjckYXxhyoq0uIGC+LFw48bOasZBCic/24pNt
UTVtURgTPc10Y5wpF6ES+xrcQ83T6rL3ePmX3/LBJr7wzPKurZjkTNFiklM/iSLGDH7szYcwWX6D
EPOVaxUixEnMEmOGftWx6K1NVW3n35472p0Y5R9vrTw5rZ5FdUP7U51PltiazBFUdE7gnzOqfbRF
7QxxhtarwUHv77nouUwOCq2Ru+Jr2t8/m6eBI8yK4kucNdWQAnSc+TMywx5lAaiGIy8+AmuMN1IY
JM5fXmN3I8AqAcmo2uJudXyYDhdJnsI4caq7Xl5O3lGitqSpY2LJ+GLkhFtK/Vi0ktlvrP7cY90P
56Avw19yCJ7VyIwY
`protect end_protected
