`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
huhkCp1xAa19GTD/MrQ7700+xBmcHqKyTDC43CnERbyBfXNAzAU9CUqfNPDxhJFOirIWv0yQz8fY
cpC2z2ueew==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
K0Vb7HEDNytHh1AcmV0XqdBEo1myp0RAQCKEngK4UJEJ74z/2Wob0uh0z0K/+fxYCvEzodPxdjX4
C20ARTbXqXdEsRyxMb0WazQCOYKyx9sfganvQESYcC3awPPMaSSxGj6hMhx7KiWA2bJ0WVgoFeay
u1HXBKRu1vbxXEMHXbY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
K0ijBIM2uPO9l3rfd7jb7Ich9JFhv7WRcXZiw8JlAsDWRmKO7v7kdQEmDZiNnbQig8n4mYZKS+3D
mliSQA846aZ2THNkvMWn/K1TeT3tNuOkaF+0SmWdEQ9CTT7gnfL9x7C9RuvvERDmCeohU0zC9Ncn
H0QF+lgho/0+cA/sR3rLvuBS9MREgRtLLhXRzh4dvnIpeSMQt/HwiFVzYkwC2dm3RrU3FQn6QhxC
zlVTJSaCNOp0QRA0nWcJmQKzXx57exuuJIV4JiE/qV0tAq14toF2+kyMhh5WZv2wDTC5qhjwZgTI
pzBtgTnpiE22bERTHruJ+/YjIRoz2zgz7SIHgw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
1zCXIUP2czn5r2yOSzCiY5mHzR1PDiAtrLqvoLZf/Ssy+3CH1wUf2tME7aGhZ065dKcui4jteByZ
GCoYfDV/l9VwJr6EyQ1F9Hvi2iLet5Ieo9Pw/vMNkNL8X2w/ikVkmAKdNfAHJA+U4hgo+Y3uQkp3
gx+JZOBuAqk1yLwVppQ=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mTbfMzkG+sfin88PoH2kYiZi0JQ7pPZ/DI5s6isAMevnLfCePc92Fsof6SEGLTfTvVp7A1uXRwHi
vMMF0Ks/aAM+QOdFwl4qm7+sVTrE7UAAMP2BnuV859OYPNRRsWpQ5iDm3YSRBh224I0vN5QnyS/A
pPA+zGiRXMIiYiTezUgSfPtbBzz/zpOcVNsomEvkDQzWwT1I5TL/5QGRRdr1/nK8DHNt0e4IAfJL
wPjnBnMedy0cbzNKNkelckGmLvKKRUJMr+slajjssXXtRtiKqD/2CMGgrzBMEIAGI8mxRn1IqtYB
V3HR+3I9oMeIVzlBQwnJ9tIH/CK20+/MTNUegA==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
PLuU6qjTDiPB6Cs7c0HqWqtCN4uO3BI0ZvmET/bLOpJGPbVwRPb4YiMW6X5dthC2TMnTaeZ7NCyg
vYORdyZmpsmS3pI4XF4IH9gkbZ4dqyhad89nDr2Ubt5do7C9dKeHW9UyZUC/0Js5XQBIKxAU43x/
OTfXGaYe5afmhsL/UATZtaujZ4ORCV8r1aEsSWqmV6ZvK/Z5sE73XevWFLcpADLBRpJwBuWXhr5v
KpobX/Nnr1ntsAiwu0xjB21Gn2mXLuQkKD3YD2vwv30r2IlEVOxN1QiGxMvNP2+YPMI9QZfqLVmR
aPtg5yHTMZ2Jn4G0fPyXFN69e3lvfzwdGhPvqw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18016)
`protect data_block
FdiBo3TnN0Bt9Hkm5Zy9uMT1yetTzd+e+2PTvNoPQOJEJdiBOdIHKwhQ+a9NTO+uIKVoils/eSn2
V6dsUeNK7QfAWUEi6bRgsP78h4XoDJ49owvkGDfj2I29tdkB/Efh3CkqaZybr439R1q8d/a7nwEp
k/zs6EybXtsbQEqRTeATKRBZb/rnIEurzIwjiL+UNB3A88is+D2dJUQR3GRXuz17XqUsSLljqonG
kyGMjd0gAeMPLwd6ZQn2zFFx28zjvSPhQt5oHdov2SsuxFe9X+q3G3azRzXjURXZcUQRYiU2pMxr
L5Kh3Neu2R+NOToMN7F20TZ1BS+2T1OvHQLleN9Rav8EhlNWU2Zo7yhhFRHKqXoZkxaCVDPxkDTI
be/q4gpaDQGiq6AWbd9ifbWXnlyPylH1/h5uSdY1w2ywfQDFrDx5PRtftYVPmDPIWB5IaGFAmpzS
bJ14assQt+ZUfRCjycSY1ZgQtTFQUcV/O9Yq++2B6KqLFw2os00F7tHU4Ee4NasWze1bQ1bhZ/jK
iSD1mf/3pmPjhT8ljB5GyiLagCwfGHOP9VqqEkcpwnsh6+rO9Cp9VSqcBQgt5WJ5kFJjzgVrK1jb
BWxysnJBLqm2G4/9114sEDW6fWrsJhBX7KlgH2CzIxUcEuYQnGErk1rIKaTXbgW/GjLfdnT7KLSU
f9V1Oldua+kgrXR4WFV0/5BOf5kO7J4d/vuTXvzRYbia+Nn51fuckY0vAoJnY0ixurNgKWXNMb0D
LuG/RmmmrL4jsass2VRHItkedqW1WhR1W5t/tPD7buAqiCWXXWI3IFO7k9hymdKLtHFPQMnUFXv+
G5dNLO7QhguGV99WGBqKKkeb2/F841oHwR+/CnjtjPeWT7uEQe5wOaNwIT0L6FSJOHix8JvBn7yD
75W9rbZ4RPO7ggY2OEilQaeGnxN6m0vXs2MWWqqyHQOntZ/zmYytavlSwAC1pdhnu7ePywsTEs+9
CfPVv9YlziC8EJJFdsqvQIQboo8JeGzEfi4OtTz+xdf4kJzw3+b2UT0J6qRSWfJ0eMmm3Vk2did/
ZZP7Gy9uJG/13RQL+HDgQjIw49gfancHDVQmc7Cfaco1mZlnPHKdUtOK9nWue91XkObuJSzpuvHO
+zk3/+j/LoLvbD7u1ZK5ByutdZYzfUyuwtAJq8HIMNUQF5JrmoToUPU9hsz6AREyIeQj6DD1AqAS
3rIiJECCMOFFgujNpgUal7h4QtbhwV5XskW23CVU/sfRK6g/ghlAZGvqNlHfl/ZJBYuL/EMVsccB
vLXLvbWeNGGnzbjB/zVr2R/4gIkZz+snQS7pyWzNfNcuvCQ4TeZIcAbCKEegVrg8hSADTBTNpHre
XWVz7qvS5Z1gP4gPRe+gYDQ86C2baNNnKdGdj2xzXV7KzSrBcFUwbtdn7YwKT4Ga52ZQ2zijBWh+
1xufTSo8KuFP7F9DIlrVk/prMtvET39DKrsbIOcAr0lVUySDtMzYsDTNe8JmwSytjcUMES2KYc7T
uwp9KnMU/i4W9y/MknhtKVK9I0SzIJGKhTIiHEr7r60v+WLIzE7jo06NAXq8cANt2wljcQs4FAzX
2c4c6MlkntMjQGfKnnZsd2+6gyC8kNug30JhnjNit92s6hTL/+Z8sKqayuHx7urSM9lJpmnXH9AV
uKMGjITMsdXx24Yz/in9Yy0MNJYOq+r4gq745KCH0pvIeebQM/hNfG7e9IzWeImUpwvOaMdhF1HB
f1sPd8ZmdBvpOkDt4U5TVoArs/DD8vn3iMnl1OYj15JUnMYKCUBsB0t4y2ZNpmlzAiCDjjgyOeFs
TbZ3PGyP6Fav7Ffn1SxBCsh+GCXcRqTlqWisHn1cHRfn5twGGPYmt1xRq32+uH/8tYTpGynp8Kdl
M4U1QpSrvsPr209ReY/JZk9yudE6aJKYwccwI/fxt7HQeG9suQP6YbXvIlNOjoLXDhoo3v24PIRo
pSaNhPKnHGkyljwsnIVJLnlcm/QjEbDe2yfGHfNH+vffwkdnFy9iz7hbqzMjeHJ5GQ2jcY2UaCZG
BmsZHrW7S5f2Y8G6W1J3gyviJbbkZyPYRDvDEALwL5OScacuePrkow+IciWtPzdygYg1jQeSGbKF
dh9iCBQzNnIZk+5n3Uvi8ewYvvewJqIHSYInkreftPxsaKqsQgDtpBpY+tVmAAm6FrO+DqClOB0N
VYZ81BnHWHOyJOKGube8VWr8crYPbwzN1+kJOHYUV2MD944zaS05h8dFD3Lejp80zw8Bvdsp7gZi
1+OVSD1/kho/Ps0FwlR3wYcliP8w1ac+9zjalgi0cdrOBjbdgjwmaHblFs/s1vIwTcVusv64//aI
df9+1dRXB4Zt7EeHsfjprP5i3BsXQz1m+K3he3ogUf4EKoTtF+f4Q6mFSQUiI4k2m7vyg8utRgQ5
h3J7RvCpJ4S62BLEXr4y99O6rMpeA5ut36AHQEoXHFCZTz1HxLeyzgOqU0kVSdYn2WVwgRvp+glg
GhRHqSswyHZXirhv4lnr1rR2Cyf+8LEIuS9ZZjNaxNOsxogJarSIlW2mwvRdhsbvX3E31cJXLhi4
BWO+oXOF6nuOgBbQLoN9r+Pk6Jgv1s+nXvCxbYWhPCNkcXL989755Wdug53Y3i78QtNbDLj2PjTW
skk2xPkfFCC+JNYAWu5XFo3J7rvu40b/5UFvErWNKeUU6SE8NedKmAy7g4wvR9sI9+6xTWYN2Aon
EpxwPROjCzVhnt05DMvIQAeEcZzbAWF5OR3ob3jZRy06hi8RqWz+Vbr1cV3JqvwlOkglDKFY3C2e
B1+Y3yRDKrOaP9bon2II61Vzk+AhwKZeHlyxk/u5x8Ga3QpEm3LQr3LScyQvHPCEQmZYr4FcM1P2
Mc+zEt/kqWahfWBVxb+XmCcnZ0NNq/Jv5T42JdaEQC0AYhEywZ5zorboXycUBpzlskosMpjRsL07
j5oT7s1etT/UEDmfMK9VZYZ6I/Biq687NKiQ/xA18E+0NOyEbR3TrZbyCKy3EjbG4UMAsHt/LeQX
5Uo3jup0q1sFs1eMUXRuRSTLWboRrIK3xQr6nz7e2T+fgjaVnFwmlAukXaTtEmSwClj1kg6THmKA
MdcxkAkbi4rfA5SJK4KgbOhaIGq2pY8R3IB4TLyEzTnrdlg63JONELRYTnEfboDINb9vIZCY0zB5
5LVQSJQ5ckQ44gbtzGGnZJXhbKlcFZ+GNOQjrl96oa/yXvn/h1MnF8zCgaQipLclg51VcHxSGq9r
fv+kC3u0HHzABqaDfjk75K+kzKJ4bkiv7oWCFTzJHwjt/Qt1AHxCQCwTwi8E3BFhvm2j8Ahn0DDs
BbUJwN9AcdqhZc3jr2snv+gu2i9f4UmxfE/c3CScRs2057kA1whG80fXp2rhmN4FV33Y2Ebtp6HB
utKa4NB4SXbSiGWt6p72AWsHtzfnqcCCEBTxeBNLXkXAO9daeTwRyysZAF8BnKFbQrGN9R1bplcD
CEXxF4HUsYSMN4rx/3qIBWIYol5GIvDVCR1ZRXEojWD6D47ffEwuUAgMjPHgDvP0H+LqQpbxYwzO
3bkUuxyp55WywhfDa9heYVTFEc0QCPDLIpPh5bcayHBZ02JIBeRKwJJZo7csNDjCupaG2mdvn8F4
hX0TnHZfRc2x4Fvf39IUOlzW+tBijRM6M+yfrGC3/XOepVHZl5xnfRwLQvizJIssqWZDPPIIAgRm
QogUWsQRreMWDTbiCoQHwhb4CSJqD6TbCe3jy8zBgEu4A3KivqXvvcODcowZ1JNe19FzFTGGSAu+
FgzgYoQUfpaWoZo/W0VkvBCLyqDa7ONp8MyuVGan6lHM5CI/VX71ZVF3eTofMporn71nkhaT73Ev
kK8oMqX7lh7njA5TPB2tc5BwPpSyJ0cKR8/Tx/YpsnL8m/Z7OfQSh3Y5Lc7nl1Qhi0zfen6LVnYE
krJ+2p0JcxmtPMEMTt50c0ildWXnsxRkrJar4Z4NYfgAgHRGgs/5pWCzLKNj/LFO0Be8zCMcJH59
lNYuJh6ZNF0GqK4zPNvgMued2UgdMFctmDISDjo2gS59IqY5nr2x3AAqoyKoEOG9qiQK/KGw4io+
Rfam14goXhUJ02T6v5Cy0p4BphnPJbVj8B8F26oS4gedWrTw2YSH6C+YvxUwkr2O5GnWU1XKbCrt
/aHkGywA4oHfgjucKH2Bw+dVp8Oiilv4KdsS2AqK2aIH/rZtl3Ug1iSAFueGmSUVybo53PEHdFFq
r0zct5ASh3MHhAjXERcVtiSd78gLr8UWlBWTY5AMzhxejq9vzW72gnJOkck8SM7p8LkNA2SIPkOq
YdB+gd76qmycIZyoBIATq+quIOClynk66qcxbsQQ3PA4py3auCRxAqcYVbdzX2yDQrcL1eks5KET
dNSy35XeckX2luIDrNSwn167s7fyWWwWo1KGLwOYypsuuVwbMNhAsCdYlOsIIninqvI5npA1JmqC
flXtG/9hohpjEDtydwIK0Beh+hkmFsj2ttz08iszEeCA3uipSAGv3JbgfFzcu0VpELHS0SSpBfkO
kpbGlOC2ESgZtlGxbLqgDn07+ig01AIzzWw36DgOeaL4p11fZGH7DEBh3I/BiyfWs8BaAS2HN6Qr
pwArmtNVam1yRGijqscRGdEtJ7ZDdUFk1Ajt2lNDD+sPd3YPOmyjQrFI1PnieeLflWcl9LdmxHwA
SMUHAzAIrB+fnSMTuNi3k6+dK4uPhtCcD7Vl4lNA9mPefFMeVkPSoCXDTJLV545FLGle4Cyj9NIQ
WTvEPDE9OfswF/9dtX4iyWd5XNg4o3FYxt8GiHN/F+Uc8iPvKlzRIEHqyoWoA32f06O3tLZlzqnJ
gWXhbnJRKOxqW78oep4aeSF/t0RZP172O+umJGTrg2tTVRGU6wvg/jmxFVVlzrEKdysGnOsqC3s7
9TTWOwFL90XHvKusc36YZod6m2bZgoOs9izNpMQ/+KAqpIr+AtpIANUAJAc1WZHLly6aihm6nyFX
pUl9zyQ21/9oSag+XB4KGtVwgIsT4OZBx51ZC2w22pMf74DwXxFhQs5ao67sVkv/E5/NYq+JVsrk
k2IAPCQ1cfzIZKIPEO5eJI0t8atWvyzORScr2NTgsJQKWh5AysCZ9WxTFURLDfLzEvWf+UieFQhK
2B+iX9MpIPJ6bVny2XEpsRHubqwdYu6WhHEASyWtVGoRu4IT1U2yshr8faaSmxmYIf6Ft8zX86zY
4eQePG056pDZdEXNuBL8ZqxizG6Ck6yUxjVMea9o15dkaxLljktVxdJ7pMlp46ruvQeBlb8XH3fC
nISmO70TvLQOm+Xwi7WEb4pgHBFb50/EWQwogB63OeFXkLbIQorU4fwa/YmFwgU7XBC8wxHxH4G4
LUmU/QC9egy3HCVUjINfeRDFtRD1/R0uX/r5U1OcWN9Q4HqwSu5mo548Ue552P5LhzvPN6BX7PCN
ZDzLoJnthEFJYQuegBnwqx7Y8cPMUJEE8G36yErCXL1ALhnH24XoM/aERfQzAsFdI75jrbCbCSV5
H/Va/VpQVn6Gr99lLroCFxqBYy4M0nkRejIknMkDc4SUHJltW+2gUzDoyJ9gY8hxteshNAnKTu3L
S1D3bfi4nGh7YfA9x1zmVi4z2DTmp89lOWhykIAh25afumT5KRxM3eH8s/MeIZaqPRAmRBESi+Xz
UmXBJzMwEWvJTsbYCV33EBH5Y6F+Mz4pKrIwUTPtDPzo5XZIK99L6RAkVek+rEJVTmj+gYIU6CXt
IDxZ5/NaCPO4oY2SuqTdXuedw7TNpRxeMVt69iT4In8sNfNjmaQ8XRmXw0xyJ21Cifg8Am0LCQMc
pltSEMypiEGC0jwrwgGl+cuUds8L2OI9XSh4C/0edIjycpY0DvsLGXzFqKY/5OPqZwHDAdLt+JOe
VW8QX8nojHhSVL1nPL0mn5/H/fQhjW+8HfLRPSWNKRBlfSYevzXaVQgE5mIwRe0TTFarN6eDo43q
GF9o72oZ3wv+bDQ7xJm2y1W+IX9mhYHVbVnlMoQaWPw+QJlbTRv2g/GAroMOCqbNw25pKqQUD4H3
KB9L7y/niXl2su73kpsxJ27ewGcNTv56qNh/YPyQifNwCo17YzpmU1yPBO5+ogb2btrXfiojF6eb
WwTtVuzNI2DqVb6LNg22fMgW0I7IOoL6h/xVZJ88VIRWLzRxH6Lpx4w6bzC0OvQqGW68JGxObPar
eJwG8IU67gtrD9kzgAVRVm0OPDx1BQnFMveESac5dzBD4CWCVyvx2SBDnak5T/nAR9Cu9N3p5S4r
3UdMBICWdNi041wL90sGOOfcfOXgHRV/bsDNtNRQh+K1VBUDfCkosz9/jjLINlTcSpMpFP7W/GeP
iJK0htP85WQjhq2Ad2ST6DVgfQaIBOtkF0GAWHkUBwUbaMgp/v+R0GOgkVlnm6OgRfN/8V33FEvp
LLA7pM/4CqIFBQA4nYBYRL+4Gpzo1p5Wk18u9KuV5fLhXYBIodZuWa4bXLT+eNqeLK0/dkzDHXqh
540kbT+sBur2Ax1rQJ+5nECPnDnoguIX1xXfRUJnneDO4hWhXqWekerZZU8jxGkpqNrZzWEU+3wS
OnJZvcDsVmDzmxV/IBI4jitj/TWQr0nKAmBxvOPw8QTT6LPbyYcC3z4F5eG2Rb+E3dNQ5gKzqxoV
4ARU4ntLlmD0EkhvuQ1wZ7HgdNEqpzo+GKUHlSMiJ/DP5tvpefhSteHdlFCnpWktYQ/TGfnkVxdj
S8tzpFtZvJE6rkJddn2m5ETo8XpDfoicEEo7fqqXZM54oTaibkq9+14jlm13PLg1ZdDxRGQB0The
8UXphv5GFomQxBHaIK0mYc5yFRSt+gnv5Dn3OpjWZupq4OcsLUaXUoxwtII1uo//EFmfXIJfkt7Z
3zfDkt0b3HNx7LdysWWIJtsyYolAI99IbclifX1D4hDnPNJPrJ2AbqTmxlLU2FqjC18zzqDOnt1C
KtTKLLdQgGT7gnM3DrrNvZLTrMEpKK6mLeXAdq49INo5jduk31EVjtsDZnpFOtva7N2ixmdpd38e
L1sROqILRICZkCRTqgSFXKlomI7OH1VwQYJHrM+JJIlyjga20WrnwsDpimHK5wlxXnqjQK5AWSQL
2+dXOT1cyXgssw4FwIpWJrYQ0hJKbjAbbSzD9BwS1i06ahjkgMGGLIgDIh3Z9cSorG6LRNCmgMxr
ZIpAXhwxEGFHeO4ZueIdZBFT9gSZon8NT4PQ7nzdtxHWyCzujKcokLMKN1oRqn3FhaBi2tU0sFAm
KxAw/T+pu/gMTMiw8NYHQ7MLluhF7qvXgA35D0spl2t5J5e+Lv/uZAHfxwcv8H9cyntfZgYHm9ke
XN6Z05nzApgmtIW9krEf9YCD0gV1fYY67PK20j3EQm1MSWPYPP1eyWT/yz45yuypY2JgnLbbL5Vz
lg45nWFiEuv3AhklfJQolzC8G5MTzet1bVLGb+OlVBn7edmSAW6eRzXGQQObkkDuEQ7stvA7y0Lq
8Ogm+Pbrwysjs/S2ARVegxJhOEBvmA//EOS253tEl2JhrE10qQ8taC8d9bqPXJzrINw9gOc0rsFP
9fcYPUXPVOqxPJHg0j5iAXILI70G8i2iY3I84P0091Pr6SwGuvfW5BKbN4phE9utA+ligHizNsP4
d6T7dAk9trx10PXGFC11TiGHyia7G4J9RLDDE/N/Kn4G9uvfRAubc+f9IquzwmGakQYYVbH0Bigj
HE0kuIpXw0ik4BuX1k8zVkcME4tUy4A/QnfPOAFz/6WEcq6Fyz79W5PujKPRqIT88hQBhbGm5sJ9
iQaJf4MdvV2q/zl5e4xTokEACDebjdA5YwPdMHrJelPLHTEEEU2C6lS3KFnqPnVQAcEygY28dm7g
60YlPKKnEbZx3biQvGvT52NGdGDjDCIgSCfTR8Q/6jJRoclwW5HtJZ18hdxuETwps0OEpLQ/+vXR
X6GLl4ZvHMoCUnxYpaN4vAHQuDwqapLdxW/+LZePm3YhrF5dHiAHqyC5d9/+vc7Gi8QIV9Fy5Ql/
6TlHEOy0/T8Mtc3djyqcr37lU/Lq3CISDJrYuA1OBPPU+2gwT0FT9H85vlB3DvKhgVz7zgpaO9Fo
uyBVrwZv8dNKsfchuSdyPsh7sw2Pzo85g5kgTe6fFCEqnvslIJ21RgqpIxN56vrze4zJTyNmMO2J
QwmfA+4hOblC/1MgJU+O9PyN1gs8dMepLveOcF+1tBqPqlZlgsnxxRBH09gEXYnR5lDF8isyAxln
uCMsc2K6DqaXX1TQ1D4Yz0De6H1PrwscjZC9g3ckvm1TavYWeNklyt+nYjaxf1Axr+BeQrxaQdmT
CXHFUc1hsjJ2FxjF90eDh+b6urkCHVVzP8g9t1la/B8Of7Fwby12sPDB39SUUrWcBu4e6KuYwRTS
UCgAwILovf7vjytmC/MS8sJwvAIE8xVxLrt7kNyA992o7j2wuNg43qK14MJFVOladcMnyYOeA2/5
ocyXqFHKpy2mFZv2TM3ikMfhPTPSuZSKnXS0P032HU0KP1l22NnwPPgW7vLVGue0JYo+8CZbgxLG
W0FhKQ8MCp2kSkyZERNTcAFTcRAc9BWqdIjMycagPeXQQR4Nm/ErrpTc4PhotXARSi+VZ1KltD7a
yrpXonXJpIq0Wn+9iaXGTnEDPlAICGsnFtTdwF/YxEFDAldC+iqbj8M5bmEEtH13N4cEbnxOAASt
Lwmc5pEX9+eOm8P1AwPZWxFR2FBByJ3K1oOWBCK0oQCt0vBNwhDq5TpKBLmKKoYaB0C9bke37D7z
ANaYp3NVE1kqAGmOfDFiRqkIjuh0mHvWD1JHTqT/PjwKVfeIturRQjPBzB/UQ8oQhXmw/WtmWLBT
HadyCQvwoTKe4noU746UemFmi/KiabPVVnnYcmc5O9YwWd9vmFoyYFmosn9PNlKULZf8grbFpaAe
y21veo8FOC98ByfvRwtpXrc5Y3XRF/baKwWYk8PtOMMECtZdoHGX1XjcKY4U5AKkBIF+IbZ0BCLD
YO8ZnhV9RMkCnwl2rFOxKDE4hQy0sILnqLOBU36DhHEqc5m0KyCutlGLj6ISBhmsItBGGYOV6FN4
kyh8VgklbJWDvKuiP/cIW5dAKIoshinae0L7fLMbOR0fwBUX2NuWI6rNWIReMz5aHGbtynQ2D+Yr
VuKfo3mrVUDviSg05km4C+w/ugMXk4+yHt2o3fGLtiVpmCsaD040WIJlwLNu1U0uaBUFn8nhOcjO
qRfIJJX/WrDw4PvoAqKQtCOhbHwIHVHOIBbz6HWZZi0TO4nHh9HZEz1wzVtzneCtvr2Ys808pbRS
F83MBoVYoDWnBR/zPZdxvHyzMGKPdefAadRF+hlhDZkIzTS4WBPcvGg44mhQmHb2iuZfYsgdWfJk
I0ws6LG6eTbIb2tLEOXgxtw/v3eGfiK+N+cQn7OcFMAObPvJ92XlU5Jzp+1vhW1FuJOgcI6yjKIU
emzxkeceI/AyjhsqRGy+3ys25oWk8yfYgZJCJ63VPgh1s/bhsi0dVzvrlXncjRvg2zc3YClYsuNW
ZACRxmWkFfKHYqMCloa2oAjGskvpgyHIvt4WAU2vGMSKGpj74QTo6sXqwkoSHqyjBOw/hqrbTQlx
UTSIlCX+Jn+T2N9MzGI5LBU6urAschHWILjXiQAZ8/knhJsp1AmbxTWWFp+BvbxDZOxD4V0VJH6d
S0YJ7+yaIWeTpSzYW8/eworEUjBn+Z8c9DV1QpdUvrBTVy51sevndW9DV5iSVn+3cf/WU/sxDmKc
NAfT6gyUUnYQPS8M9Q8vbp4Q2C0i1EttyVC0PxW6HkqQM7g4TSsy9kSMEzH+y10XvKPIdft0f3Xe
9u6qmaMu6rSzPplojZSrThge/gGcddGiwckTcpYHv4VnJ6alNeZocvhm5x8pp3E7kANAkMdN922L
bstE/2FyTdCXf/GBpp/1CvrkGyHGkM4TfLD02yHX+uliIwjtXXhTZsd9/DC9N3F8UF/nHPIMK/zK
EsNpybnSk1zEVaVHCSpwZB8hP3gG8h8x5NR9cqut7G/n2H9tkBW4R8jAHX63LFQ8SDWnA1WOV6RA
ahqZktR+1SdSImmRicQ7IsUWNgGwM3PW/YoQPmmyX68ZryEAGMLPNaFW1hTYVU27yx+1DBm3Tc26
fuve5fPSCKPigbmiYgeep8Pnikjc08MBxemOSit0PrXIRVg3MZufqyQ4d3ufk7mD4yw+RPyA1EfP
505j4mKi38CwWZDHoByhcyOCzyUPQ0RqQsSKhjs1wPalVR4g7NBraWw1MbEpZtVLkzpkzWrSn+WZ
aJVl4/dug1aM+EQtuV9ehQyuNrDBtV7ZjgQzY0g/tVrmZ3nuuCgEDZE5QlHtIvuZDdHGM6V04mFf
viHIsDXNKeG+kra8a1F8u51yr7BETFIdGe1GSGVUuiOjpFp1cfYGpcaDXLVg49GOJBuOeXBeNs77
5c27CVGW3ZQN3kaeWtYC7EjNoAD6X1wTIbVycGPlvMyzpPRzSkFLnVwO5CUTB3qH01XGLlmy60gm
mp7dIzW+M2hGyp6jEWkQOzbclZK/8xjKI/0VlmAluOuvdXaG4sJ3MGW82La3wGR0ZAA2YrWLrg07
4F17hZ1y+J90hIFEEjKUJ1x08N2L1dUgThUOh5UNKxRysTev2EqSMJuWuLLp4xWb4dBShBH1T06C
LxDB0pPMEy52rSd+euKSLwE0aaZTaXUC8sHY4iZC2qM4Y3eoOAjUcbiS/NU0AehXpsdWAsSACL6B
VKges8MaXbyxzWMmTuP8esffRR8aii+k7gx8ZAs7tm32LE9yOy3YWlKP4dJnikzwsWCYNq6Vc+fN
x9HsfXv4o+Rt1OvcPFLBDIjE5tyb8j09T9r/FwZnhWTlQd/w+oiLmn80XnhQawqY6Xg5nHPKg9+W
LGW/UcQOXRZ1H8ETQ0fRU/M1XYkGIoO6rMQaBMvZ7aS05bFu+IJcMEDmwAntAfGZ6+WIxmIQeOsF
LvqLjIFWbsWDt7iiwIA7gSXnZE7aYZupJn232rgmRTsfeTuSLvW1S+bKLbojKFgD97WcoWlGGtef
yDeKlgFFvJvq4RwTWF5UXy9hkhlqdHC3T6qAIysY07G+TOVLj8Ekq5c7xDOJhEtaaGfMSpsOw3sy
umdlj8Q/r81jgPaOPvdARerwYb7SCHv22mn3Aze8nNSIHKoft+OD+BuM1252+266VEUJzjgl7y47
3ws4YhKPh4JciAnsu1scKw6nf/Gic82iCKENA0t8a9vXSUHHYZb0fQF+Z2QKRP8UbVzNF0V+9xeA
95NAxD+A7NsvQrbHqH7gzTtpCpPIVE3eduLNkmSQ95UVzHEWCSew3R5A9JORijJMCdN9b2oqPb9/
Yzl3+93SEN4/MBO8xsw/0DDwf+NB/S+DRmscgQi/b61A5waTF9zM56wGxjDCTKp6wAKWsJWI/la3
9sJaZvQJRWto2obKzDT3BjF7ojiRk+oHTTPGpE5bUTHXxdh7XVGlwsOUTBO5NvrD4DkEsyjEy3tm
QlRK7iaQOo5bSeEHq/D0DPZvazfvo8r49eF2hlBU/S7+5HPw6MzreuIH0rFDnCyaGx0FHWQuHbkS
7S43A+bAje6xSIHF+BneMz9V4Zk3c4WmmtmdFJueeUIbMDWpSKNuWyRmUW6vORVLWFwfI1lsgFbb
zNc7OdZZMXBLItnDnZIEeu40lRwGkQcujErr+XGCokIc6ft5VtEx3sXOYGpZXjFoTHgipLUwuTRq
UJCgdekcpVoivB/q26dO1I64+8va3hPTKeW+yl3jZdDxMW7GMRhy2YqvGuWXaH+t6OXD0kHoVWCF
bhQRWwEGHbPOxe6iWs5PzB0PqCGlyOy1sxEuHtoYN59pEoSnzhEW7RjIRhKX5Yv223VD0h0giD0A
MCABSda+Ja0Kr0ErI87ALmQ0JsRGE6roEsrbsLW6wZimWtiJ/dFq5cz/BjgX1IeKRuI6g07Ngo6N
v0oBXttM8UwAY3efCIthxlTB9IfdCpM7T5KLsxkhnBReC04YpohPLZH3frZB0No/U7XCRe4RKW2f
C+Yk2OUgoNFdVoF/JPs0xq+J79h6InVEMV2NjXwJHcZmIzn+nJB5Xn3hlPYgfhP0XhLQrLNBltYq
cQTL1FsbfOGPIKgS/p8mh0qnOp5MrQpCP8K2KYd6z+9sj0/o+Yvjdyx/eJZEtoFOeSfahYEYXkn6
f/LhMOJ6X6qdup3sl+V+IEDYAw3B5KcfZ/i3IrjywhncARRWwIxXDMAjYxJ5njnsuyYBLi/WP11A
qBtTaTdahf92lOYSjB/+toCrlwUQWZxTYpwi4Q4GTtCDSzTl4TWJN8r2UU3jUL0kOmqp/u/P4VPK
vCVhTkI/SywBDh7v2DXp2mJFOBZw/MhG7HsFPFjwTmhiraa4TGFEOyzeuWI9S1u+kKPeBjLiN9BN
ayC97mjUGV8SlUKe4ZiiYgFwSR18O8QBcU1AUf8m+2eFt3Mt6nNefW84SG4zdKRSJBryITxiUgBa
01rr3SOlg9Z79Dn7sQHsp3vg7OCm3KbqmmzLAb9ODEyOGvlwP1OLCOVksFvG+kPkY4ETS4IJImt2
PR8K4uDlk6YfZNAYrzxgKA/hEAR4TYFmU6QOT+FXE2kKgs6kgDq8xhqHJXjEncxG8yy7lfwCOiji
4z37+C+v1gEBzcrwlyvbxe25/3hrOQfszLt4+ioCpWYKqrwL9DPwzr9xPLIcw3ejeE/wSPmkzrG7
98hXm+8Z6S1BTKEmZPTrFox/uKQgoUVopL7IG4DJL7pqgQclihRKUeKwm14DunKgPfx8qFr1e888
cXIe4ceBesBid9BnF2iHKikMhdvJmirv5gDsAnxch6Dw3dh9TXIPiuf9JUGxEo/qrYWLZeg7cOAk
Y2jA6tvh3qBrs5dJ/jaUhXNgXlYRdHSMgrmuE5clbpciCiP0HqW2tmtosc37MGFmqnqvmLCv5wz7
Ka8O6Ngd5YXZfAaJRjFj2bZ6nk6U9Q5DxWgMNHxcU8OHtbJQo5C/F7MTKp2gwZNfb7I39/c6cJTX
e+dqjk0jJhKgJhe/CPHbTwKYaleYWIoV6ekSWyAgQgQVQoKowRWHy4p0RH41u3jpfSfqiXbFSvXj
95g7QBEogAjMxHGEYGXaEDwwiqIscTySGKem2vykCS+hkmkOmF6uC0w9NuAZPXY1+9mOgIyBS811
dIAUgjPGP3GYJvTxd3JNJ7DQal3ufmIxWSQNJkG5Lc/fDHVZwSTZuKrQ6fjDtKG2UDtrZHe7rjDu
1nInJhevpd8VGyx+tOXUG0kTPDucRw1PQ+HKtAQBESbxJlcqAG3Z5lR8bKvRns4KFqZZPBPKjIZM
ktMhffjS63ZN4+PxonlY4Sc1CEtaV0cKGgy49i2ZnEJhM7agM+WHqodYuB4Fn+hMzoK/NS5gRRER
Q+loBKOQIvDHHHMbNg8Tm6Njn1bfXKKi0BlUSGpo+HCseI9mjqDPSk+LN28xRAS3Cx8lXd6vl+vr
bRP01bZzAWoj51n5t5Y+m0Dw5wlB92lOpdZMRwgEXuMJFlOm0x8bWBfQh8njHDIQqVVVtgzbi9Uz
rb/A6YU9VnJ9QFS6sQOSezqzoruZTTII9t83aksXSTlIc49HZyLzzsWrdlIXqDTAK0DdZ6ApSltP
XKJg6TpnPUvCMIa9XBLsSA6Aabm2p+2fSgwCzpU6GPg5E3AlLPObQES7veDZkepCSJmE0GQxj9JZ
5H1rMs7qySP9N4y0sfH2WclP9mdmer5nyB6BQJ/EJKgofGdF5nlelnfTERIn5vyCoCfzQoibImzS
xEeD5pfdR6De9shSi2xq0kenuFpuGyeA7I/s69+n/jSiG4bw1acHxxfx8ZXcfvv4ojMqgLh73Agt
rKXxwz7If7IXQTuMqKL870dwpn9/J0keKEsxQXZOzUePPqTfoaHVBJXIpyaVB+FpBuGiN0obnS8N
aRp6Kr6dVRPM0tvo1+SGhcs1x7OPbZHYqT1F5YkCDoogMFVvVUlyykRj7TwMcpRPAg1uXgwkoLBr
6Lf5Vw22j8xQhaUUk0vdQuu88CPnfr6Sqeg+tILQRMCFHlbFHXbCiMQh0O4rmdTnGiuZk7bNB+aa
zmcFSTweNuB1M3DTKy54nEwiX+U8H0qedxvurnwfi3MhhQzZTtF1Nku2d7ppbBOkLoAwAbhA+ahT
Mgl5pmC7w+M6DoWxv6DilwGK+HgfngodFdaiAN+wc6gs4NNq3Cng4zun9lRwGfO17yDt7WQREcvC
KsBlx0GAyEmPLI6WV2xfh3RtBCZMP3eq6GduO/g1InACICQAPx4ZqTIB6Nv6pCJmWYb9N72oKxPv
O/jDSuNyMHskZthQL80XeN9tjrRYTx4b07d2pnyDHJ2HsejjkMqlZAADpfyZDIhngKmgR+1t1r/I
SlW7QfNRH8UBWbjX9jILaJOB3P4nfLRaGKciqfjN26KneyhELNwsT4Nh8tmFMzkwlsE7J+UizxU4
g2AOD7IsgSiLJ2Y24c/60A6kkne9S43vrCkE4OkfGRvoBw13Y0CdC4J/7kUqg1YXj9tfbZ/sSZYN
vLRJXTouiWMNPiGS1cZqwA+n8jDhG1x1+P4XYsBiyjtQzPwY+2FwEIQ9DsWx7SZFKgwEnqQ54Kit
1L0zRCMEjE9SqGbnfi85ytI5IR2IEUXsmiQJ64WLFn1JjBN7u2Ewx9n34ILQQ+K2H9CPX9mLm7Of
FkeKsSA0SXXqyCWs94GTSGobNbCTTjUw/nV3WZe8tUYjrbMWWC3khklgMunFporXlJmnDUmdb+Zx
Y8iwLbvMnZCD76JwVTW0ETIYARjGn62dYbyBOc407uY7z+c/Ui5oswM3jHDY+Z1xSWtl4tuqzir6
wLdNMY88rjmM+0ksGNFmVio9nZ3bq22v7xjDGLcWyjvvasWz5n++YJKH95QIPzcTQo9kLt4YUp++
aQGmOlh6T95qYf1CCT3AOAbFvRIcJ1T8EfOQ8WtVM/UMkBIQilER599153lOsSnE59se/KiV6bHJ
584CgmgMZLkbO9xlXbcP4vysecRf+kLv+rkVp+4CyHinSKwwRJS5Q0+8PWeHXoajHZ1TqiExJk1Y
5BcnQ3Lwb1DKvBxnDu+ms35uw0PilOQhD4/IkGf/V77p0mhoU5sJA2kUFk6+DRIV6Y44/MS7+PQH
jB2QC/PlJzNZsf5xLAa868PWBD+w1hPwf+O++vUrmFaMcItfY/J32g9wY7eFklrvFB3ZyDWFdCx8
27htT/eSccXthEMvudnK6xCEVDNyLDPxLUdSPJ7LOrIDfe13NjXHaeSjYiZO1cUcaMeTy13LEtft
QEiHiGL0pmLefwQFcprPyBpweV2XsEAeEjt2JgwqjYNzBgOy3M20HkVeMwA6O5Vl3kvpulG1lQQs
VJbBG/PD67zC3542fLIJrNpXh4Gy4jxigOSyrgNqL/34V7dKhNLOOs3ERTtpqXUGReo6TLfQSqm2
3OkqnA6Y8U1b3QLUBDDnq/iv11YdO/LN0MNgGHBEQ3+hiwbn5lyrbZWEAezRXanFDpNssZBIv3cr
cXrqTP8kl+E3VzfD76BkxPWq8rPxMdE+0nTpN/Qcqi8OYyK8ngHDHb2PTdqbyTrFaQI8t0o0vdrJ
WwmS73AMkSgwPDToTbed4dco+SiBecF9oxdzvWClxBh0NlDipWHFRJYm0pA1QsUBwwOXwwESoCfD
x1Tf+bjO/XMWdNqhq2GTobkO1BoSke2VWawogOLK1dDAKvzJKr+mBmkmjv5J0XxTzv1Ao0eL89XE
UBSsvPBIyyZCVdAL6HejS3SFbb/EhCOSOxX7clXWhKyyAQrU76XPncogXLL5N23AsmMPJIA+WJJ4
OCiAFttXrNDUBJbs1rSPlsIGnjIUU9MD60uKzlI5gUefQvxVX4RBl5THkbNCWpfb0cD2P4E3F3gw
dnszx6CHi3z/aqHGmXNVEtbNnNAT5POhdRwKzPFOizE0n1bI6A1+D19ajCwBgn9mncnyUlTb5Pkr
TAeuW+cwu761aYLIA1Gmij+nVrNg0O7SGfw3iZhdVGiIE6Q/8N6fJp9lPeCEaRJRzvY2KTFTrK0u
YsUjwKy1yNyS8Vb2r+Ct8B/5QkBVNVkA0j3cWSmf71IhQk6UBMe8EkXt+9h+STelYhtrdHTyCYwv
SSfKuukmm2+dL2dwGjoXD4aU993lJ1XrXwlAyquwx1AxbCgxI/DQv1bvsVZh9/XR/tDepy/MGKQm
Oe8mayRakPiUGtStxdckMqznLXte4ipGzzWpdyMaAHRQBiCk1u2KYi2gMwkJ2GwZv0sdr3TTis46
EgdQSzpFLv+am8zQVao14k6tyJ86Ng1tmiN2T2V5xwwCeiIc2u9BYJibAeA/8/nK14K7NrEUpyZL
66gB03iEjLspzcmNeE/hMSqi1qg6OtceUdv/jAFXmrJO6dBR+OQmd7qty3NNK1/I8jKymWn9IKQt
O5rd9GEs6ZQy1WP0+158nH7tmXyyIJjw61oQCDxi7pqBUKhC2PKhFak8+aT/OKq3P7z5dwsfAVnz
1b0JizuvnKWmbu2noS1UyNhAuQM4J/AZz/5rtAtMMDz7J4CnJnKsJXMzh4coRhRlqbGcJgUDXcQt
Hn8O9KNCSEp+JeTCrGJ3BdBtDFnytblqaVQNqP76V/qnKLngLtpSSJJa8esD1i33QyvCe6+GEhi6
H/+p1/YniYP6zlZ72Zt2BrIdI71T7k8w2ayk0YJkCwHLu2yBUMBgkUKjHZiYS9qMbCCwJKZQ2IGF
RpUXGAAVOccyljIv+YTW5GoxrdQSAySr3PURovG+70yJb59cKwLeGgSvHWoSGt2YVJT1JNsbuhec
z+lKMr5g5TqAI9YcKap3/llp/ubiTHff4mUDW7cmFj1PIgqZZq7yOS8KR4T2GAlFsAVOrltQsz5A
GkGaKCjH+8gqntUH8jR/xVZGzdmiqmO2Dw2mfApRaxI/g6wpwY8qrSmzvDzo2ePVUozHadTQmBDn
RvWwFuNFP5+bh+FMuRtj3ffq3TrKnYPbUU4csSLO0dyBUWNA+0B9QuZxCv05iJcba5kRjZgI3go/
LaKgPK7+phD3tCHUoP74kFnyvnvZKsml/Rb01U2lWtwM0APTGgdNdVfDIm09g3zisy7atA+9OUVB
zg9g1PKawUShD2Dresqsqf2IKANOwBU92fp6QKK/dveKj+qldFIbNpPJ63VRY9+srty2j7VdeT0z
do1szYo6nXwKrgKt3jnAQRUa5iMHYkkyAWbBQIRzVxA7/nXfqOfptfNaaQXxRnbPnP5kqw9RQEXv
+WTFixq5oMSdg/OMLEmhpEzklvFN4S4+nYjDNxw1SLTkNPGXhD+iqUugGDLtAb3ewFPaTq5M5xNQ
OxDNeUxCzbQTE10sFFkmPYMmzThIxYsgasIIL67qStOeDdWoEq2t7hxO9X2BmZe+C+UIFIdX3HXr
vhkGBtfNKCJWQXGN4yYxbkx8LH8cH2BEO7x337MlZR4cwbg2PNIDNoUN769+znKjQrvttaEoSKCH
DMcIZx9trH6GkbyvJrTG1U/d1HIiPsShwk0YWsgFOFLML7dRU0ZPH/xcc9fYbZRG8vtUALfPaBbn
2Oq5YPEkhOv+4Nf4Jp+NRLJ+fH9Kp8Pi0YJKeVsRxHJAkQo31ZEwuolhhov9sjpa7OGAq2PlUwAH
GvI7i2kOXX5T+YMdtnI6nmmj5nLI8vvePeHAHaOWR6dWflkAvP/Wc4xOOq5H16TBkGCTin/xYpLA
WdrcFWKzNzDW7I6KCwKvJnfYSB9l4B6Wdtpryj02GPPVtjpPhxHColjVue5VhoY7y0HoELui9yDP
PTEZaNTSPb/jEW981NtvX9U2OWCVeiYKj8VGA46pNEwlnGdyXQU+1ef5QA/xaFuti1DCEUlztMwK
TVd5Kpex7m244KwMsks1l6ju4H3tSrFiNJXBH4aMdY1yZAO3h2m9pJGNIRoFsSNwWFjg4rSJ4CNO
X9c+lpbZz4Efe4ADnnLxi5hIUECIzX6XtY4icZpB9NJkGKdGjqVpe+2EHyIXbbvvaJtxyK/RneTR
l4Zry4XNhfI3msNJi8as+xh9hJzBDgGQq0wX76Pc8DTwV2XZ+ebbWHQdNmucLHvqnvzpkbqTaS3C
5wYlCyjDw7KT4KsOfP321R79nKYLgjZPZD9J5HyZULgdTo0BtAUaeV3N/tPsGrfcTt66YSmt9xxD
7l2dFEoAnI3hdEsIyxZyTG8fLdHPO4fRSXw1wdGKlQv+KMYzPrFzugH386HCvw/nR0vQbiRO9yjs
eJuX3PKEqlX/blghGn60pBjcvbePvcKvou1T4vSudObU8A/U0usTPSYkjFdfTloWMKetHvYQd6EM
w0XKCs1PePmvD1nPgHnut8HVBn0J0HLTQQutzb5OvlYlU/JuPyPwzY1U2BpunOYBp+ATBI/A5mze
k5jyGgrU/q3Bn8Ao7RhKXQ4n8/jZmfxeJoqF+ilfxCO0vc56CTXJTO146+1D0oVm2TDWV4xlznhs
Ufla2QTJijeYaB5a9tVOeh4q7SBcc+/BUjZAxmsPdrY2PX9Z9t1yyszkNhoKUwNmaiKU5mOghXUS
ELwXIjtFksXh9bM7vOpKUIImOQjfTCeE9iyGJXQY7JuWQJwI92qd4+W5kc738tVRfhUj5y2c4aZa
QmdozsjAGDBvvW44lsVnricV9hYGyyueQm2KAfDQmQ2u+k6JAYu5TwnMxiPUsk7LKgIIg146b6Vg
/aYMMdEqrGgAzFT+c7C4BdB7y5OxgnDpKcexVrVldv4QWt3MOyLOIsHd4kzwcauQWIPoDjEpiZmK
oqHA4FlY3ZiWvywE/dcH8Dk37B0erBalme8Hz9C8Bu21oEplPuYdXU2DiqYV0v5PMADXl5L+7yk9
ThV+OvFkA/ApRqAE6V2annx4S3heYTrbuVGU9GLBg50bLmw4XvwUW/B+TXh/N1Yq5f9Fn3TzbcYA
EjrK1Hy27ksqH9VyauZGM0KwxiFS3obnJxJXJLbQHj3Kd3bq6+CxOX/6GoApHw0XGS/hh4X2scVy
Uup39sgDuDeEbSmhxOKw0gKdSxe06RfqhT2DNloC4PxAYIlwse4f+uj7/yWRMdY/nmopSYPkScR3
SyCL291/r3DRVG12ddFaGPgViG9tRiBEtQd+ACSa3+UWifJF1yucyB2+8FU/aKZTWEJAP+xtelCW
4HdJ8T/b8/YuLWP7on4pSqJ763Nrr/9WxSk49fFrJOlTJOYthYjKLWVOUS9wcnyMbK5XysrLDgQ5
39o7HLsNyuDaGY6Soghj3VA3M+WbPTJudxmJs8V882z2Qn5pl7DgxWPamfhxugGg7t4YJhe6Tg8D
IjBfEEE02/7G1W+i2o1AjGeHoqdFV7dZYAzDULBiYN1BDQQRkFSlMYNrF27j4e1k0Iw5iuYJTKft
Zx9QVilrB7c8no4XUoZsuo4Sgss8aaXvvDYNKImiS2BxGZOLqS+YISZ6OOx1CW+L3G3E6Vp8ri1J
l3Sjn1mICeqiMd7v+c2r/jpC7LD+X61yzcgQTjFaesmMyJ+br7nY701B6+8v04QAGwzXeJsZdsdp
V56HCM05SBNhKYyijJFhrsXur+J87lXXsl53k0th1uNTnxdkM+UgSUvYoRJsMesYSc7yKacj5LF+
Ly6dkdTNn7fcTk9rTjK4h0EGdthwGPhEdJy1H3BcA1GdqJDnY9R24bKJO1kDFT4VzaXm16d7LQFD
9JnVg80q4E7VqEQ41kJUZQR1jPH6kMxAx/itVp8Eo0K9Hh66Fk/CAmeYcMU8xVhGqVoovQm0rsR0
ntX9Kv/oBpsrBYYdljcf+pPaq725/fPknpi9a8Bob7kLrcUh++KS7gyuBd51EfEB1YbAlKJPn+lr
YI6fdH4SZ2JErNehIvHsj7BTIJIqESM3L+j873yyjnCn5dLzoF9UyO5H0AUEKvkT4QTq38z7vHK1
hpX3WqwrL6gVk2dba0Uu0n2hkxzQpOZ8bRLd4vUDlyUFxeQPGvA5PKcnT6qx793RzubEAR0sNl3X
EH1lbFesS6Jzuv1+4rzHc4Kd4QSo7ogr4EeC/Tg1HNuGh2Jvy1N3dvwQZx0p7/RZtCTLf5ADhmgU
IjSsJ58Ox34cAhjVd8IVxPsOiB3WCaliBmdx4lY0qAsiBIf2E7o6t2G6ypGeU4YTaJajNDmw60T9
sFDC62ozJpmCaM99gz6QjWzk86GC8opXhJTXG0hxk7DqriKjAkE56KuLv10mg+Ew8HvNBWCo02Ro
jWrKLtdsxNyNcs6JYQYrVxPCru9HhRKx6hIbfnkGU2E5Cyr5k/+bWx0+Snw27gevju+MnRT52lGT
W3Yo4k69itj6PxOzOKystsEVwrHzGoSpewawtt6ZywpiFhH+573jT00wckTnXIAycsmY3dMq4ZVC
kkLLt2bbzAfZrULg+x46O5ZXbCXAeWKSFoFs5XdRHnxK4i+nOuKjeUZ8H3fH0hIFSvnxP7vZNg7T
qXrI19gdOo6qIf9KWSWzKlzVIS97sq3gakvRyU0S4+fZ/VmDNh+IXKLGBPt2moezdb0ZfznoUYwe
JlbW18CGb2z8gE/jiXl59qgRw51QLFQf4XdIoW05yduXATpAWVEl2H2nMwXqTZVBGQ7/iRH4stw+
rDwdnKt1prdfi7dxhTvFMgr12ZMjCrxYDHCmKBzBC/PvC73gvJrRT91wWLfRxKpQ6CJWjLYeCo6P
YYYi60RQ+YKZZwnR2zx56U0HJcoUthZRNtbLHn1uZOxHNH66ZJ8+ULGiTM95SFPENmDMAidl7mvT
mIEtPnr6mDtnjU5Z1rIEavNnpLkG/wN9HN2MTvv2v4XcFBFYdrADhsMaUTGW+00m7eHyeRM8wchS
dy5a0wF1zfEEorG1DzEQUGuzcnIMlPgkan7w9C16qjW97Xm67IfIQpWg+Yn+KRhYK54z4V3LUk3N
JXxX0RSLNkr9ZCtrWqXUBKGxLGngwxYVlh2568fmwQYjg9Bi9QvWVooUXIdXQ6AT4m5z3dsYkXs8
ojmFRhbiNbANgccBaGsxeEq+aJxFB0rpPlPUyFSHKFRvq9Xqg9t2CiVfbc45Paxmh7ChDOQ34WaR
S+F0QCQc3FPHklmbrxBLpmPHC5ZogwBwqRu/OZa9/YTcajwxkOEvrT7HGVZYkW8OqMiAyds1SW+I
GbLDzi3/WfkQA4ljQ613J/YppHnoGHgrBb6ZOZOzdBFnfSxw1grsxxQdfBrFVIzX97y/lhMQ4lYS
CN8nRtMbOtYdo4E2dAws5W1DsvBRXVsn3gbcbWv6jcITeL/5dQ1I13KYOucfd2ZvFTqgG/A1qhSK
wV6jwcF2jddjtuBQpGjdBP9KtiJmUGJG9vFwtXbpzOqnHSFNUtCsmc4eDa/onvGmaX8S+AbjGx2E
NXVLSJVQUjAxpRHJ1JgdoCMVuhlZERYZEUusUk2/EAXkRnvBxOYkdoQdKvqSSGC3D+W3cv99wrX7
FdZ3etxSdbOejHiIvGK6c2A1AXmydRsiCQ9moAphop0SWB5cmqduzC8flDKlT/RDbVhatA8smgMX
OAYOnivB9jupnQSsbYO5ETu/hdeCuw/gw/d5KrPYimjIdBlkQIh+5KM5ooklOieNHN3e21YXfpjS
mQxQWFIMwkOPfn5ozjNybdWGWsOoUTMhehdZw+CLGH7qdq6NTYdD+eZKNEK/BybYhocLZ/xMYorC
Tz4Hb0FrFHgV/RV7yKvQrW3Sd5KT17ilcVLPerl2hagQzKTYRJRDjGyEcSkBZ8ut/M2WzdnKzTtL
YHwPd9h563GIdTAvqQZgKsVsM248cChDAUZqe3RnX8wttHRuXDtfgXzESemmgnOg2/1dhAXaXtnt
28df6bhvFwzPhlSPEwi6axJ96V883shAEmCOnvSK4uHDxEP35i1Fws52QjoaYOtc84u7XZ2UTNn5
kfnTLutWMoJarZhzSfnoWUS0DYDbdCRzLAymkF15gmOXKDfGEaCG/Jx05Ot9oI7ir2KXnl8VynXK
PU4a3nIGU4uTyMoLJdJvMT+3T8mvgN8lZdkBMhTKkrajlCIvF3j9gaDilBm32ZPT9AX5WA0QZ6XV
SmGIN6PXGvYTrYzWyPGdv2+HDWT4pAmrLhklNZeJJKa+fY+aVa544KxU1FqzzLYOEL7m8I1eHfYs
Xz1hr1VpeGtRwUdcjS6Pi+NQpGjyxSvqzWOUF06RayNxcNU//GqqwT233bFSCJySRR8UW6UZ3zGK
YkpXVSaBLxjJj0WjnqqIpLswXUudiyM6pqNXhYtJ7cFG74Mh8Gnijs01rcnvdCB62Q+EwLpDSdfk
A5pgBv2wU0TexTzTJ9quyvdV19fS9zuxFzsfiZmG8WAR5QfqYUfSiNCifUzRWauYRKJMvRUTWHeg
0SosOEhK0ON1BVZgdOUI9u5YTKjET1uUmAb7SE0iA/R9/2t1fWEWvuakCFDw9EvhQheQxLuoblzA
rI7uvrHBxZ1wvtkTwztA40AUR/WCQPsh4E6eZ7dXkxaZnM78TQk0IdvDVIdyen7bVUsTUfXPJMxH
UvSQzjl9JggdBq/2GxwblRSJ5iyeR2ukqydlaNh3g1MuyuOys/nfeRfuy2qXX1fwwSHsc764tHcy
PB5DqEfCTXOuIrTWDjNdmVlFjkW01U+2FKtt6R7EsCW+t47xT/EFmzpLFVbTo7fpk1vM7KVFIm8Q
WaXg96tDrsxXqFEGDCZlzeMpV3pdv8F9XTMYGkVuCeQUn2fgj0Tuv82SoPU6/wVs/Y0nXOyf0ReZ
760KWPsgSURimb5PkVo7GVKJrD+FwRuLA4tgidv6CmDcLlc6rJyo9ajzzYVd/NfZ4UjZZgTfy42Y
+iQRJh3sxqJDARfeAmmEz5mGJw533U+XiCaRpUtqoNQxa3lkQ3QMGL2AKq+hhVUDUxOZiHKWAeS8
FdUpYwvS2hYFRqL9MaXq/pGPcSK7vHuJLpWfxGryE+uatF3Wvz8jXBojotDW/9MpzMtYnCIHiOVU
mDcssG1WSJapseL/wSxNzs2bHEsxfrCFoIemmysk5Omi9Ps0aE+YXNZJPlP0CH/r35llysIfnIPF
oQvr+zkSSixUhNiG/b9JhTgZkEkRnuKYtMpho80WVQ6qJ3Tl/gAX0lp0TgoH2A2es+CY8dXqL/2N
bQ0C0l4OhKxluZhzbVEqtArMFcfjTTmGMYZwmFfYs+8ifVIDEyaJEWfRrqZXIWhz8N7ZHhE99oYZ
Dnsf63zSL5FjPlFx/k04PKQKRMDSzTE8+2e991P4fuLDVg2eGOd0zDRAfWqJYg5fVvh/vFjossJ2
iSrRLiXet+nF2YxlS1vm84PKtKOES4NGaMg4Bu2hQgXd8Jwyd69ki0S22VzGGe2ewDgrfvWVoQeW
wsHseWoHXFl8GWdRsv3UE79ZNgxNsPd/njfXLadEtOxxmRDcJjBTccimReO8+pcbjTO7pwaLovGR
m0cR6NKwPVTagnFmQkHd7gLVszyg69GoRVRwumFqOROUtIH4tbEqslSMK/z2TevGjSTIorZNpfBU
asi8QATxunWTUvts/NO0D9TxkM1NAsRHt5wvw1quvafE6jktJh6WCSpgQlN7EHenXgXfFSFHUngP
6fg9JauTPyBpOl/RIaTBt4/vsIPoUEFVq3kRz+oiuZXYf16aHc/pv3JtSTSA58Dz2Zrjxj0niBHE
Um0x9z4o3MBI5sE30m3BP3dBdalveM9S0hcXbyYHv1gbHrWLFRx0kMR3KKcrqAzPCOdTIuecSZcd
jm2TJsj8x0atjJh8O/BWz0tFMkIZm+w4IBgD/xIaNtnl9VryvKjQOhzXM1vxoaDy9k51YmO7zHYl
SvSV+tWDzrajI3T9bGu9iAoSFmUKanS/CQ2S+CuL5rcbzVQfzqoLNAh/va2jgRNo5OfX1aJH1zfc
cVIRgkTvdw3INxrVl5WenM0s3GZLRKsQhEGUGnsH0Q503V0wsH2pPj7Pl1VQoe4QL29b0sAiyPZj
z9LL5g==
`protect end_protected
