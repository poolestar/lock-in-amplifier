`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
BwdID27ChASGjE/zTvl8Wzi6L2dIUVnECqEjAXJwL7drCiXiZnXJMY7WULr9oad+z9bLJg/0KKX1
1SUKQZn68A==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
czRS0jBmAO95aaC3J7FMqAhYw5oxWCwx8YG59grJ4JJPqAHSwylqjd+z77tfozIo3x4/p9V07lfN
/d8jlDjc1KT+7sM9IH21RTwcPq0lpUSby4ir9WKWsrBOVfBHjzGCGN74hczzTG4+8tQE58S8wUF4
c8gK3PRox8iAFS88+9g=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
wTJ4eXo2+ipUBfFs3DnlTIuSDU0yk90g0e0WXwKyW7+OBsqepNamArtdShLAv9zGvqCig+496OF0
SPaZZifpzQV/82GBxBEqi6o8J10zJVFs5TKyU6FPOovBFEef6vzeJYGRd0PtYmTzDN9K3cQq5siQ
IBaZ2aNvEEo8sxuS4lM=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EIO4vM0JK40s6PZofL0KCfP1lo2LlUQHTPj4VfSL53PSNxn0Cocp9Xpw64qPr0Xibaalne12snbY
zIXCM5PSAzEMM4rNA0n3KUt7ukr1F8niHa4ThjkWTMCcrNXYan6MpU3WrHmShcEZd6enWAUdpnD7
fBkA7WAwIT1+Sxv/iZuUKAOWy7TUkywPDptQo/Qx/BvhJfhNonViXIesqpmk30laV4I+B4nHxYUb
fOp6HT+OuN1saZNXSvkB/s1+1B6cchN8GyCtIytPNFpOeEDjB4/XeAlAX+DTrkj3icz9NGaL6zhw
WL3cLmjCMG1mNiLnlBfZpcidvfOoDlPJkkaxsg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GvDlqLi6q2Hj92rSgRhUIhz+LLui9M0bKlq62era0Cx4OC0kXM4WY9MNvIewhX8BtNNcnptzIW30
KExzfZ7Py+ehKeBXpX1xvHl5H3Jd043CrxqLHYODMV+cC4mzi1lMH1wo0vj2bKpR5zXCI8u7FmQm
SuAe1q1FifRWAAf173O9YeSc7sCGrzk8bcXnnwpG2ao9L3GKjPBR1Dk80/ouQnKTgtQhjWsBU+MO
rZ6qqqdd0NrATg3PMnvRi6l/KQTW3sus4dNBudF+GmrHR1x9AVvlCblfiH6Av0RJ7NMUxNdhctzA
JGCJH5m126Uf4olhtfXxY27VLdqk2hIqqTtEQw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FPonn1ygHGox0+DpfQa9guUUholsofBfytZrz3xlZHFKQVDfIgbypN0x7Pl5vRKh4NBVrQXGXbiJ
CMxlORRpW2eEsqRyBzv3brvgx457k28crfqT/MH2aclvcQ7XkEHW11Rt93iM6/fLRuyoz40EbqZG
1OoQiDTq3/esdeuaZqkjZkf4ul5bTMC8PhodueaDEGBMnUuzq2nbL1GD/dFicHEIWCQdpSavipYj
Y0X+kNYFfln+YG+9cVHPHFMrDHxsl8xolflu+ZyADkoSQUGrTD86FFD9oek2EqgjSLGhVteavoJj
sVXlIYFwVQBjFWNz/miRXbvYX3V7LOeoMGRxnw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 432720)
`protect data_block
HUVp7Eiji4dvdeb1FVibGvFJ8+3tMP0qVE1YHKmhmPK3uaPZwv3X0JG58CmMIe1Kjlp8XkuwUj+5
nYOyU/6kFPOn7wPcX0CokFfEgN1WqqOL5D2xpu8kU2tT7iFzKOKjXYth29c94t4ye11NiY1tohnq
/VPGFrUMomPwjoai39au2aqkNJ/UE+kJyvy4DfxWXStdqRVtO0qa9DgREoTPs0BfcSnYpAbx+KFN
ujwPinB23/betujKJ3RukOTLbfylFzLIFKqxD36UJ/tEp2lna58loajv6M3X7dNa/32/F8ueWf02
wZtCZEcwOHOVECuxInOlvtfbv420bnd0w6yN/BHK/4Dsl6WbSbYecL9hmYNGqpzAXEjBxLqXuzCs
6iCY4x2WIo64ioFf4WrZBg3LlKpFwZ+Ms7qT5RfGJlkF4OMauvacB8TxM5APqA7yZU/JpBAminpe
M6P7YJt4i1+LaswT7rKa2B9Si5IWZKU0GJ8PtYzrXhOPO4B5cKsvOlIqP3Kb6mfECYNa0lDQCpHS
fMl9i6m63V/UmHy2X7rHFC+YoqnaOwoSmejNbvDAY9DpAkJUc5tffBCm+by26Cg1UnncWYw3+Szd
W5TYatQLgAsQekWocYBRP6HBL25/jVksr1sEg0T/uv3d/+f3lZ3iUIEyAmM0AtueDMXLDF7as+7O
AW2miPUY0M/GUJ1dagAsgJZy/r3puyBt/wR0fK5jlRTPL3cnH6Aio+Q+mFC+EVypiiiWXfQo8TIR
4/XIFZpLwLPIc2BYUSpdQ7iP6NxJLSKJQoZjBWBbu6CBXDeudUdnHND+JC3KO5InaWxjnCtZ31fP
Tm6zCMw8wLWo4SdhqBFN0kI8LzwMnFJ72bgfv0HcSjHTVaDUMFQKvexRxNNcCXMqQZx+Do/NcUyK
lbZyHQnJ1AlrUlrfRR7pmIVy2h3NaIL3ni3n+w1JOXxGQiYL004zKZfHBC1anzGpQQ2GOVfQqM7u
3ZyOyXjJ44HR20x6UksDVFk9pPDlm19l3Pzs4a8avSlKNw1nly6K0v9Lq/2SFo1GlSI+JZs6cGzv
8BInKq7VNx0EGzVIUr+vnQdC2sfWTtjbVGkpx/okH3a6fsKeEqVtTQRnqG5x8ZRPgHTURW2hiqtU
+uBSZ0VTFPHBRcXkZfoHc/6WTsByZ0FNp1krjvIU1iJIATCnb/Qu055cW9zeG+i8hQ2w7csVKe4D
TVQfmngAGKSvRbb+ZIrv8kplXrjvLf3lIZCSBvzN6OuJ1SrJXT5KHrqhod2gXJV9XO5rEAv8aizu
ZnWJaztuMnJgYkU6AGKGpdrOcKLpNmN//ajQ3yjXTDVSnKw9dxL8ptOzuh1aPWne27vOH94mDO8c
TD/NL3a4GQGeTUfW/Tmt7yyGe9WJt9n5h4hz8qcG0HEbylmZUTOkaOLdotTXKU4YpgquSSOhCLnD
YT0NMaczpCrMu1X4OOaOpIuTTV5PsOFOdiC8OcvmfxYEfRvLI5tL6i5bZB8xu0bEQUVeneW9Pftu
UZt/59MzqAEYRuSdcPUaWb8D1AbXGW4qq5eeFNphsllYEk2clMQd0nqxNIkI7g3BIn7Fz/LlmAdP
n4tH5iLuLNxk3aBNv8ZvWXFVVasndNu9Kd0j4/6yXL3s2ddVlBqVtmfGO9prgZO43BhXfWhYfzgQ
sHNAm5pgJdkaIPxSB4YXHtlHriDiKgCzkgX2Ky6AUTUruB+2muKrF73FHuUyxYQaLYN8seg82quH
YTIMcN58hNz/N+Q0Re/ufVBM6Lv4tZlYXspJUuJvkWfe5KxrnFCwCTS5u8XV9ugsOBt2WktAwfqO
ytRmMiE9A6ZnyuG0qt577aaL+oegLapx+cuz6HSjdJP7NLFjUgIZKuuIv0HBCnJX2j46PqNISfmf
mq3GNgfAMjNExp4k3yBB5mFDzKxIpKkj3FkKDQUL4mLl0rfieXhHx0vIzwehg6tLx+G5bEcgObzB
I/n4jJ+WZPtZnsT1xkyAvKctvYlV8LF5NrZS9Co8cYYz9fxI+8SxrUdSIhEHqJvy31IlcZGJcpM5
/plrD62ybT88AZ+JxaCxwDYWoUs4ZqK43J/mjPrkKe/mVzY9rZ8ShIsFApSWfq0cvF5b8eyHKvb2
Os9fmcYsuFXTIv1Ky8HgszTS3hC7A3V1Vzo3Cqr/LorcaMyMb+ku7wSFba9ahWps942V0s8CVo2R
QJrD7A424ZRg6/LHcdGFHsIxghzRrn0p2Kckw29FWOxD9KDy+AAZtj3KdoazgQOCnOCwWF/zPMMv
n9vcl85vCbf3Rc/jRHvte/QX5VVDnEBPeTSx/x+mc9QLaX7/ecGrqcbUmg6qQ5P1hAP0rUMRIgN/
HpJJSr+bQpTRNDXcBUTbVgmtXitx6LQkP2JlIEdVybteFB+63JB0L7KXpzZH6lRR/dlMtYgFHtR9
N9tOkeZAvs4kHrtntbyzRdnOhvV0newBeNwotJGRP4nYcDK2W6V6kXkjZ6EG3tRjw0EGTJSvfvWZ
jZ2MNWnQOK1HjCUXEQBTdQT4vaS4fwqshHm4Fb+o7sEZxcKglTDnHmKY9AC6pMlehpZmEtbKOfh1
2WmtI8kzdVB6ll7l1n5u1vFVLMFg3bOE+ZiQinNcD2jsndFa7G+d7W8jPM1vhcqupKp+JiehQEdN
TLg14NTY4G1Z85kyNsES5DZPS2rGJdyTiEYD9reg+4mHAnxoiI1YA0cYLk84wyvDA32A6T2DK+Ui
cms7ZHVCxB7TE+GelOlKAzAS0ws9PrWtLkOveHXfb6D5VLsjAdqPhTmMgUKm2rqApYdON3t5aHGO
T9aXyZ2WBlRolZZd6qnCy3l+2Xzob2uE6qtrmRVJzK1eA5j2Hz8XFSWGTO0vsOJA7yGnCGzJGF85
iv0XjrjXyHkMu8e4RK+ipayjylBUFP6/NMCwlRy9+hoXd4WNIueLYPoWLiMFtAoGO1WIBqxkRSGV
13oDjpmaI05T0i7rFeFc1UJ2uUKxo56yGuIZs0WdY2cmLj9S8R4N4ZFfAyiMSksy7CGbtggwU7Oh
TBVAFgqZEh8drPSQmNF590e8a6iDxn7eWmiyVdRLR0sFxAKGw84+6ZugZDDLrejT94Jl0CPjUCLf
My9srjlko9Jf5xDzoPRGZ7m5QnYPHHFg+oWQM4FIjW/yvFbm6pLFOyFJVvFC3By0AhEj6rjR7yIc
CaLEWssUrc8bGDhf/n6NWQ5OdWUKXLe+jOYAncq4ww9Cb4zfhMu1J5cKm7NReHimYh6VPZQ1X3k3
8lAKdZ7w8dmmmuApK7HxheJHqawiUm9OLXIrwVYy0iSdRd6nNs/2ySZRV9P6NP7GUB07MJixcAkn
n84baKy0XQ0RAsbvDLkXR3eyamJjkIbnVLAAcN6gMq0LYKqmsvxVJnvTElv2grOD8HANZol0gvT9
6JsH27XBtHeNJDUZpDneStZSzFDsjF549JeiWIJAZKh+iAy4g3ySeLr/NZl6lRNIUUivp+ElXiGm
Tse2N6mo2pX4wJKtLBcIH5o9PrvJbVOn3riUjgmL7+4103y9mk5BsVCtjlZzX7jjoTamb8i/TgWh
XNn/r29qju+otXozxekLKLBA+/5zs60CXwNnMifGp+22Tnr4Aou3iBzdEPuoqAdwtFl8/UismWK2
dGDaF6yx0EUbWi2ZNBzey8mKUnARJGtrTCovEzoJqsUoOkVJRqagdQoQ+WC2pCTsd3LkRkyGQlyr
lfArKFyqVa967a3IPBMrlNNeeJCwlPXSu2Ce4KJL+yrm3DTPa5Xpt1/QZuTyEFYqUielASKGgHou
+oP3rnlX9PuBPn5X7SPhML9iV4juqWWRUaCHVFuuE6KWg1Vd9Tnexx9sna2mogm46BuQFbbvrwle
ouTqM7o075be7RjGzityTgZstz66N+vAu8nZkhjUmCOm2hjIGU3C3NCq8UDgE+5lWywKFgTOTfE0
9yTYmJDOVMOUKcgi3L+vtEUEc+8ckrGnJDTH+4R3ZVWileKYTaMsYJiN97wSiwLnLwdFA6lhMvOe
k7pgMCd7kFwcKkLx3d8G+Jnmmrg5ntFk8EF1LW+mLKFyjYwKPIETwsc4TtEyXl7ZFKnVI+3+vcj3
67oojEVhKVBe0NJ4nSuWGKt7AkqCJdywUKs1heg8anfck6xSe34QBCFdiD/NkpR5/nKccz2OO0lX
UGVSqUbJZPIyWVRCUyf61PRIAv8GbWOsZPjj6BKCYWa0GPprRrWaof7c2JV/vicglhEZYuzxVpXs
UXZ7derc3AL2R51cPFma0BfEsR+OtFSFt9sqrNrsgZcRUHm1T9htRn7vY7MZrKT3b3c5Vved3t8m
ViR3V5u/GnJIyBAvMDSxEiKfn0TDf/LHoeVdZGMWR7d7lYLLu+RaUkztd4HAgxWhVKXf3xvwHeWL
VTMD6yN3DKAma0jTsSlw216aPFDKSSt0ZsBeH5N2xTAIx77N1GsKUjIcxBg8mHlAvMkY8VKnqT+q
jQr/K1EBh2sqLhwtoQf2J5tb+OG/Si2xXSoOxcr8qVfJhnxHPG2+MZsl4HW+eb8XALWjFW7M0jta
Sd8StaHkMDH6WNGBGDU6Uvbxjl6fj0Y/bJpOylpm4CSrKvwvaX+5+Z6xFXF6U9t0UsUT/KlAkWI8
X7dK0NKNX8A1VlhdQB3gLyv0nTn/0GyD6c+0jJN8rNKf/Fig3bluV3AbJYe0/XnoiCzG+n0lBOWR
ZHJC3/xy48KWAd6AiDmcH/mtjY7lQZ4KY9Hsa3D2lmj4qxKyu38OXY1+MylHk/R5kzhRHSO6OAjf
AF/LHJjvXzECsSIrvs5xAIuq9wh/EFvfFOGU7jjdciBqkFqgQUzLJYmizLcaQL5Cwpxunc/RaZi8
yqoQOSIaiFMl+e4DT0FfCGE1ZoneaPzS1gMZ5ZYkuUXu4jaCujFIOs7Ln1pLhTPt1tLsQ3xa5rAF
5XfgND+lcxDTNmmFRP8Z+0kyrb7QxLhrspXQjf14dQDX2ow9WGjcwGMbyKuOVBB2Vcc+I+tQlPuV
8XMkbDGMotCF7+Gd3cON0aweWqWceX+g3vm4H1TIKlYj9NiNW0iD4Dj7lZW/1MKIGzNHETVsVLNF
zrhcn8KnsPmgeC/t3b6/kmIHw45hdufx0X1mdWKY0GcDe963H+Fi4/8AxscQfXSmUVO5+bG4yhRb
f5EXSKj7bEQw2BWDuOLAicxG709iikYJRiJ3+qEssKhoW4fSFGL2vyDOC/ZjjXg2tSLQOEP5DBOU
bfl1zm4hYn/5wqs16opJh+J1k1VoVMCD/datgbX78Rj3kNyHs9/tmcRwpKY/4n+kVgyMCzwwDLoJ
Ctaxk6q/Eb/MbasQqFgut5vUOED5qyxBHMdQ/WJvEkjgoZAiTxdnJr102n3i2gUFZe5qckvjhrxa
qXFWsSZHfyCQqzQHvJZN6YpR3IunYBkQh9sZEO1TwT+jnYr8y9ZXVGrNJt5gyPgKkeiO/t1SlDY8
P9AnSw7oj/OvDHuT6e4U9IP2AE13myP8lI/hjMli+W/o0cP8VN1VnT2dgrVgRQhg/xd+rtmTxTGV
g06DnMkoaqvBMv2ZJkiXvfa2MRLGAGR2u9k/5WgeV4BUn9EgoIGHYA8nfHkD0BhVHMZiwMo2UOP0
/oJOnDq8hzWjFV3IQOsefdjOCQSkcYVo4Um4cV6aqr6jmCb0nVfQykbrZsiMeylxdYzEyvjPiedm
yqrfBRhi1eTnIHfRAYel1rZ7nug6tEpFeuUIvgdklw0qJbm2qNcviAWOObUYZq+wHlmVxyWqoXBj
S4WLQPS3Gok+My3lfxsVRG+GB+xN0F5BVz9LEwd+twDnKHURXZ+WOVTO2GaTO1uD4rFUI2nPOyMl
SPg11Xu8Z4Ex+PYt7oJj5KugDivyyxBmfMGoOtpx+hC5/iGb/W1ODJrebAKJE0zV4lyp3v5NYWJw
qyNtB5tpMCayfK6TM8DcfIP77UTXMh6TffYNL0a7AvyKRMSQ1pHuLBJly7fmbhX1QV6+sxhGXCs4
SHNr0jCttaNOZM0P8I9pvYLkjXSe8sCcymKyOGEZppxUvkv4GqQ78L/p1K/uTT5lwUUIkJc3IrNu
HJAryDF1lu5S4TAHzn5aVisD83w1ieA9Z/KL+gueSh/Wv1DV36flMSdF4nYvCpy/ks/X1o7USKj9
Bf6IX6FqXmD2SAq23nj19JcjWoZF+HHh9HSOBOvCLUp+Cm/I6fgCI4YVNcnm8sMqx0Rsnc28ANK3
K87WKPs28pXpAjYPH0lV7jppBMNfXDoU46Bf2DMczh9YmDTPDZsKeW9DLrD9SmTpJLZX43iVHwKl
fbO9MU5Pge4jUXv6gTr7dbjmBIlxHHkgC1KZD9wWBei08in2WLSpeih8xPF0/zTp3QV09txUsBWe
YwPpnWkxXFJzEKfN7jlBBa0yU8L36cV7M8obWyhMQ6FoyE5a6biPUtaWtfG6U1xsJ49PgXuvHy9R
5m8KW1ietx9luak6jH/l0Um0iQe2UmFmyQDJuB2UabOExiBfcH6fNJBzpk+OjLWKoUwCHalD37g0
x/DRKbbHLkJockx5r7TxL3c3ALaWTyik5C9Wv4JlcksVHOXBAXKb23pNdRVJ20/+3nICzb64JY89
5WW8I3z2RoxhS0xgsMhIdGOL5kv4Sz+KwYluAJLoBtZHLqBKLXunLmzbiLfAdoJyQm5AmWTHNv1Q
IktT9GpN/kck3EV8fh2Fd64G5gJNbASkhqmI+WnS4REFX2pwMioULAlCVoehKUT+v2DQ567tFCFn
ITjHGMstEn2yxJIILqEM9MJ0hMdLOQ5W2RS3pynVxSxH/djgU7BPjeI//9nBABLsaQKKSLDT3cPP
wIjrw5lTzh4pY2CDr3eZQrCnRDCD8fZ46E4ENfyuZe/Qr8I7oDzsFRDShLZdUBDpxFVK1C+Qn7oE
EzxqZ9eZCsb7hpEGOq4a6Kajm9OzgyzXNk+pZFQaFl/zfAsYUzWF9hPnN/yspnqUSJ6mT3zNmBDK
/XbS9SMH6fXqNmYXCQC+G/R83RejOxMFwNseHNASDd2EvSZo/gGmtRfyaDqQxUeCBUsSPL2MHMKl
BOaeAduRBmFUCiSDmXWQOf2JWNrDjnJ7hoyHJVfl4aApQXin3GTvCrW9zzpmu5xWp/AQQ+aDf9te
X8OYutDNhfE+wKMQoaMkNClKQCbJyYXEx0BlyZr7fgGv9UEilH5tcHeYGlSRv0qquAzAYcqhmYbG
E/vOc9mZD9mOSo7lRou+T9t1EMPi8zph87bIKGaolVR+cSKpX9sk5zJWVwWMrbT6TiPm+n7lPQui
uQG2t8mJWRB2Bh/vRDGva0HgK4mZT7zjcr9IX2lXzVfuiwZXRnpZgEtGBUdtTmosKYtp9SiQ1prS
riiOnYebQhTIuOC6efdQqyVxHgLZ+DtqXfc4dw54nnPVDSu3qzF0Ep9eP8VHTP0+nUq92lyLEJIo
V9CkaugbSeZ1iB307pcFCgAtSca2sKdX3nfqoGEbnim8TLnpkvdiFpx9Ec0QuJSrzT37a1Zc0p3v
WMKeTqzEPQ7C9Kq1GgfhaBztwr7m9AQVyd/LyII1QXItvkBXNj2gxsZcTB9iDHD+kNtEBwcDhWi7
z8zDpPKgXmEF1wLFv2zYO9rnhDhqkAmb2z/E1QMJOUmIe++TTMw1X9fkFUFPGsUz23HM+eooMsQi
W1caHIEJb7jtJgYMbcOVBwfW9liT/p+irA2IdetjrKvs/9gUxWCVWhusCzM0mQUv2o3iDZTRFJ4f
bh8grksEk5NjwyKSKrbtRWaJUWulMfqWKVXBvyoXDTptKSg8CuIh1E1BBM4dj1kKMGM0Kh6VKnm4
23c1zFvYkRdC2031KV3jtPuo4WgVIZ12lza8e6WragnjHkGxK/pYLxK4LqZe4WbRociZWxSneqPo
JdR9J1funVVQo8k/DFHFKTse8Id0+JMAwHRtjvVwBmUIG7XaFZDmWgKT2qtR0pX1BDrJcJmZscNL
MEm0/zKgH29D2m/ANWV8xouOOxIsekznLNLMgMgZQfI8ouj/oNomQBnw+bZmfT+S/5E5yURmpw4H
k9XXe1KXRO94aSz8fx0/rLEVdUV5LAIrXoVd8ld3URMLxftlB6Bu4X1D81KR8oNUkhBtDieHecgo
5Z9hggaTEUTmIUxGAayUq+0+Xud7CnWu+2jSgmvixPTdXwSXCOmi9PJjeVOR13juhg4LpY3iNS5A
Hbn5r+dBWd6aPoufMZD/tViVxQnJtSsTuqzQy89q5OTmP+sFR5s3G56cU+D9Rc4Uvbzx57V33iQC
4gqgtKfXU/dElMlvy2cQkCEpJ1NRxB3LORqG7Hxhl6XXz7lkkwdsuWDwlmzVKAlmvd1EDUcA5uou
MAdNuet52+6N/ynCSgZzmdGblQTS/Nv56NWuuWVgZ4CKoUud2IcetcBSUXJ+P9H856FZ5Xj1Ii4P
UOaDK/MczLgC8OjVXIpe/Plsp1tKtyW85ha6H+n4RnVLwt3ItcFG66jU/VIPByX04ljvZokJ9tVc
r5Z5HhhJ1TESAZFyim1Ou2zAzaEvgjv+YNpeB80k4/rHk+GenEWjYk/sSn0yq4KAoDTFFLPuXEfB
eRrigLzMcqD1YQwF/V902jBoY7i6/r56aihfdIC8jwYghn3VtLmlMoANZFpN9ivm+3Xgx22VBKeC
2nWPcKCb4y32WxufYAT2ptig1bax6cjJlP1muUC6Gpe1Zk4a51W1b62JfHCOfi704xaVYX0LqooC
VZ/y4tIEhFeAxeBgxHIXepvA1ZdtY7/sC/6juTEBsj4PNHz3diRcmvuXcUVKoM3Q8MRHRo87z4x9
aUawd6QyP4iAzRxtkyE0B1+W1c1JWo4XRNjW7dsq1VSuIntuz52gzAwCnq9Rrm7qB787b6bLhQ8a
jXuaDl7Mvj8LeCGnVB+To1ZzUaEYpdWrDgzI6y15BUr34Juw9bbmnzeGCPeQf9ME57aUNC7IvrCs
UPcRjtpR6BsRG5dQuugbXisfY9D9QdF6mL1cM42+5BfUeSMcKJ/FMZTMbVL07ASEQWHf28Bv6eC+
krT1Pps5N6OCFaF7L11jbkUHXoH4V3Q6lIQS05rNzs3vEwZi73eRuo0R17scN98PPJJ/kM3PKBf5
djhmQK7da34cLY8Y5t1b1PBssXv9eHrLTWHz6n2VLfXE3gL0J3pSVfhlauEGehCjejcmyki0hyvx
pj1c5/y9of0+Hwo3yzniS/AgEF3k3Gh/c+OnT3zfKo9r5QqduV1w4551P/I/LRlu7LW4Frml8a0R
eKZ9hDVV/i8bN2apquz0whGzXzC2f86rvIp6GZfH3tljnyQa/TPs4cDY07y9gtvaH5p045b1m1Zv
jzXGIQ7q3Xq/b5VpzhlCoYVbLGqnmw3P9MW9/5OnoFBR7vQZMPdE8vd0pXtn4xuXx+91bDyKZtKU
cicp7oZqy2e+3CoQ+uRwtbGObRlEhV4ed1bkEB1k1jXtfSjYVmFTOEdiWsCI0oAhVReioXuT7sh/
8GzJ8Mf4P1VMZBQ9xJGxUJFUrYZy3Y04iy4RVSngzNkHOaMprWOQ8w0RsQCEcQ5UNSyvHHwKXDTA
bH0OF8BTT90TOvW9m/Vc2A7cWTXiWX07EjRLDNlrDn/avuc58PTfrHGyecUOYYlnspHs5t8+nkkG
zwuWhOu2WDRAd67JEfhTFCZYSxUc8Oy70rWcAbo6Sy+KZaNyxcmxUBc0oFx+xACi1BtEO+6nz8z2
qx+QrrVUt/AL3RbfDYiXNrV0Jdj6fM14TkpoqrH+ew6eXm3X86UGi5tuBe8/N6SsV1TnsQnusnNz
Ve/NpBvI/6A/mqsWr+0rG+PEcaleLysVlct4InWvccqHNXZmUEbqqpU18eurlq3VTat3uv/n0jmD
EZ6ii8Do5hBUO2GIo8MQyY5EXIbVPwVsmWEiQ4mV7fdJ2/It54G3QkMUrxkN+EsuPNeD053b9EOD
QpsRN2CF611vk+h1PlTCH1weRxopx9sBXXY7iXYJEBCZt2ZPxR/dPL+hNM0R56Xm/NTTZJtZecZB
BACii67lt/hYfHvfD+8A5HIHuSSC88bCSaNFSin/vKMn9F8KDgYuFjtH/JlwH5GNVhApf4MuC+e8
BdfG4PCPCV3BvNAHJwPiAsVmEGtGbLtpBEkfjqNd3qvVPv6STbp93ZtGE86AzYeH2K7lTD41i8p9
FDFYJH5o7vxJTxNf7xQjazrbK6YmHbsclGcDnB+/D63c2+41I3O+M7o5QuLM+XvUvjGFnlkL8DJC
A89QCYOBEFtFtL+G+U5b98xGotAxYLhsNioNse4pr8fgJXfDWtvruw2AMwTnH3pheO957qVXgLzS
0rta313PmjCTvDf9fEE3ddgNys+T4yhunOUfRVzlDHeFCGv4PmtPy+iRoLqb6Loguqb8yfnHqcw9
aUqShQAUXk/XAgPGHTnPyqA95lG5AuubbtMze/lm8jnXrSd/XpLkOZ32CjVLntPBK10mCaJhSS9c
bB7pfQY0VXY0ZZb+ww8aFfVuujmCGnGMG7uxhM3Ob4AS9NCsH3cEide+Src3ZnQyOVdLSLo33w6J
KAljEWn6/HfCyZpfBEoZhcQ0fllpjzm3smb+4qRkry3RWirjmULTCI3aN4JSR71/+Lo2T2K+aWLh
Otk2zDRcHRCSDgCB0XsojHq6YneM5maOI9PnfVSLlfStq6otFPUicZ2fqss1IBQZaF4PjH2lAmXD
NetH4XTFyLURuLGsE8FFfKI2W2FJVqjHektIM5KMkc53IP2YvZ+pl8GkpgsfL9zVb11nmI+zrDbD
3yz6zP4YMU007kFXgt14Wn7kkUQ6CZFZy3QMmozb0EuuMbTfHL56UPaMyHJodCKNDVtMfuoMkEnh
QQjbJN28MaN8Sc3MTB6Xuba5hLF4HbKCRxA+RJ8qqaGyQZZnpFgC8ecUkTnjNksJPY49aM9HR626
uSGpxPN5Ls/hu8/XFuxp0BYoZhW65VhapBjXGe/yosVISmQFniDI7lZ+L0PomHt9whBc0dFDjTRb
8yOvFWFcRH07vVOeAdi8EhziA7IXCn3mLd05b4o9vcccm76VbwpVcgyNVj6jynEMx3qe2fomEvx/
gh6xN1P0ZZAzPnwkEBvaVamRrjmY59jiL7MV8SmWG+aB5pJTpDelWCmQfVnL3wWqvpGkNaz2CGzm
88QNn4wu3RaJmWdf0Ft5aB8lUovZPPzp4z9Eahb67qR/F9wL8hGaQbgDs9flu6U0UVqaKP2hfrjC
71UBAjJgNUb/KW9NjddjaUPU2laQHioEPGMHtrlw1qbJU1/er/Y/QZTjSUPtE+JQRXq/Q88DAK4X
cobD2FIX7/0U8HjO6VxMdfUNd0rnvxSqXFDT+0/Q17tETPD/R8QKC/KnJrzBmKQ4fkrix2KB2EUa
f/ZVyTjh3uzRjZP9mmtjDLZRb51YEC3jq4nP8QgNFq3VsCSqpQr2GEWJAHeBYadnjAb6Q6WeIchb
47EiCe/J/VN1iIP8QmfnDv/9g2X8ngdBfKMfp44qcEWVW/UT3MAG4AGZQdHVC+h9ufWgFSqxx1ZW
bNt/slj3PtjELbEsnO0xEXU+MTS2V4olh9hLyCJzvq7+QsorJOHN04eiqWCZK7fKsQgf5WCr25Nk
QVPMBYTFnJQE/Vm3y6SQtiDzNc/oTQvyuyx4BzHzpwscLxN6VPuZZLY9oS0DpYtdleXAOK+8Bq5C
RZrzyTCSA1iPHd9eMexaXSr0EPxL4uw1Rm6q10cy1N7ZcqheBx1NQpMV0jfg+2dcuGDrK5fnjy6m
3jIM8fa6FaKllLwerV5jmFSzPClxapWphITJ1l7x/tw6b5ihcyVjzJ6URC5C9RqMjvFytUVsZnXh
cBnp4efe1vYtnbfz/XliheVioqiljnrkPvHCW16g/HEeU0d06odZ3FFwlM2uOltg3hMsKvPsUW0i
ULPmi4nzVwlP229Y0HPYKVywZ9kCpYSa0l4SecIKehqvUkqLWeAXJl4eJ1NfYgeceRys+6dd+8Td
IAdOQmwuBNSrBrtkMymGsCyv3KxmgRIbP32LcfSCP98EvTowi8HyGF/4JQ6IAbuMT+XcRDI07Umj
cYZ2ASqwTke3qQp8xTrIoH2kc/62YOTyvmVxu0+XpgsoNdbdMrTW8Hytljv/8TxgowkzmE9EZPoC
zdZ/gjtY048tZHOZucaf/ogZFcAtlOhTtSP8EL0/H0zlzickK5np3h5ktm3djtsJzyb7TMeMJn8G
PPrqejuR1Vn0XQopHOTB5yILQl9tZNdEMTjTo1xAH/45rE+GRNpH6J18r2rimw88BAUxQqziwuhe
FDORFjHIXCCt1gOsL1J0FXoOh2oPNhQE57UTFT3J+fFYTRIa4OU9A13eeDfN226G4r5gc8DkUCvn
9Plgr9FJN1JAJDMRnLTbMkZiIRvKj6auYsKFN3CZW6XwG7D71nHAylek7Ug5/v4xBcW45ZTK5QRx
46IOQi5iZqxxzAtzz/9DhGeUX6WMrEr+oVMgb9maPtmoYpw7Eg1k4sBi1KsTJ4P4NWBdjNpp3o3e
WcONlZpxyDSawaZjPMVPRrR5Ze/N9aMRVaS3CL8RmcY7BKaZjriE6aLnY4ewuKSKrXJcJi65Qszz
Yi11Ee6nEZ6r02ecBhHxniyZ6iqcjeoniaT6FZOC/8onw0E9fy+74wtuUVG6YJxY5wzQcmvPGdGH
4mZIG04shHNp1UzC2aYpNe3dm0hbXBpCqYCVuKTWWm92fL+LqabvQ9AbBwGkTc0xXwXPUgSfjeVd
qRi2oWQ3Jh1ZZWjs10TYsVQl8IKXSUihkRKS5WTZezWbFIw9SFs2l/H1Ux1FO+cfICnzEimv6aiv
irB54e0EmctHzrpV/AgtF9xqOO5xSOw/fA/56rWZq4rWRR3F6OJ60kQ1r2dVd0/FPO4Xks2BDDnh
00rUihEzNMXnchhTYUfdeypPtnwKEqMlqO70dAlXAt+aCVXkVLJCI0gMzvJEjTynMR0x/wdTZCRZ
fr17IoyHmKQj/19WB+vzUNeNjcMTx/h2ALEdf9S63+wTL7PWgCSY004YuFqVHc1+5+KUPDIgVRc6
ZhXNfZblRnghkvnfgtU53LYBjTVouoYlFj5K31xpzSSS3NN8BHbFlKz0f7Z0WittAJhPgJPWXDLA
i6y9dUte1hoJypXJtavLC52tZw0dJHF0Mx6gjNLuez2xNIhY44QK3HaYhI3tcQwkaOt7Etcq57Lf
31rxvW9a/aF5JVW5DkzIzXUK7F/wUW08VQ8EIjb+Q61cbv5fEqZYmCYdJv4cSx29AHkfdEoxdJt4
QanUm4iqxOFK66maji/ukr3a5so2qR++czdKAl3xtM7nKlOWB/klS3haNHRPLzdDXqZ8+F6j4Hr9
7uiAwVrqdzwovCdoR4GQnFGf06OYSEPjY5Z6Mn5sMC9UOfXA1Y0bXzocjBnfvUv5aUC+byvngNLY
y5GU3grziyEdylVnlJx7Bnr2QdObU4BiIqQd0pWj3esGsOtj9GvfCcc+2ENzf8SaPBdalG5dMnrg
OzykCqPm8QNn/d2MCjVtEMmzDehmVtiDRJHm+CF6BpNkUhLoicUv8/PYtrXhuj7dwnLokeBlTPXI
S2x9V/RjfLD+Vt6Su00YeR3JqAZbg7U9rbUTLcCq1crB3/AvqD7fRlRrrBdMn6ySZhh1vjETkjKA
9U5JxWaeHGfVPTF/vQnXE/BPmTtW2q+kXhrkC3sXtdMu2cwJ0bpvdFRVhfsNfCjgOOnKa3zWGOqB
9NYrnl10ILEfQPUDWiPDRz6o1idrFUz9jcH7fnO/GW1p0ylokUsutoYo3ZmO0oUTWdrMgdjnWZCt
04lZlMeLQII311wc7YmzDnle8wVTuMaAw/YzLAMZC2xw56pcLK6fwJTKgq0Nzli6PHKMxdvddW0l
OsIE/VgVIdsmDILgYh2nu4oFkSQZflxwonPw7aYCOnNl1ywZNSMGHSfFlrLn3upNTqZwp4BYMwpF
7shunBqL3/uuslTla2Tyd79gOk63CBlu/x3jRdaxYG1c2tU0f4coGFKwlUfI3fTfaNJBBiaW7fdS
SPG6857EVA1xwaoz0S37rydRGj/0ljFjJGD26G0eJfvux5mPlGOuV4Afs4MpvQNYATHydGBSgrT7
m+A1IwCrzQjvM3bxue8mROziHhKjj6JJN7u9/Q57V0fZyXf4Sz3JkjrFOZg6T4dnK+k0dzW7Gcfo
02qXJriZDVKxdvrZt1aWrfefxJ+oxBCZNqSAbJQzI+Knquvynyt+1BDE7z2cy7tYLx17kny1Z2gV
LC2DoJX7IDAIpxg2cFic6MZ0NJcmICUiK8I11a1ZvkL1+psQ3f9hjcd8IH262e6Q4sJHQrUW6bvj
waGVPIhn1q0H/PkhAPKkOqjXGC7JoD2UcYBRLVJoQcGPvvBp/hLtdoxpeeiNHa1HITaPdcSz6EfR
EQNhwM6x1aCyT0f+h6pOWR4Y9m6wvARzT596MA2701YuYkdyvvdc75Sj4fROD7WsoXx+VH4MRMqf
LCRSJh8Ep54I0NMWDLtHwwN2gzJ1YIRR1mdDqar8q+4p56WoniJwokx4mbdtG7CXMCWGYvpAgGbv
DKef3+pMW9SotILr/xmo59lsWyaqjYCd5MD9IzMz39Fxgt9adt8iY08v+Wjw/qUvBRtTKtiATGpR
3jWqHQWsC/i42xhjcfaqUJLL2UvWeJpSJmLhAdBiNsVVIxh6IqUGH6+ECZv8YD1X5MfJMbW29YBB
tn1Zmdaw+uMRNWrUnWYrzw9ZZDb78N008iAE26whcbOiwa/ObalAAtx2oW1BUU/kqlIt5ilZRl0b
gIxtkVbvwQp0WaeDaZGnajB+QPphOF4j58RV2bZVvY4SzGgV/UstYBcm2H44qOYsSu3gsJfhuhXZ
WiZUc5ZGkJeXc20SQtlxBPFCWNJ0WV9LFQ4eadiRLKQZrD4YRlr13t2mS+1zL7MLpu0/KrgMAJoz
eSTMU9rNNxGdSssKSF+ZYPnMvY/BmTA6Ns9G4zjM/PLrkfjeUVob4BHsZgV16DRM3+K9Nqf85zUU
qWhEvxvO0RCqronTUpgYQ4/MKn8H37O1ZWEYLmvH5UziIjSrcPjI8zGYdeJOTqSbyoFcPuXLVXBC
AOWrAEx2BO8awaFW+XzaNju/hDgIjvqyNEgl+vHiFIupdNle9SHDhjr0nmYH6wcWVCqYxXeWcWW4
8DhLLg+cfrOWGEGtcJv13nmc8+/QzgQYu+O4D1SUXuRsEa6HbgH3tUnrJC48BIsN3BTvog3p3ZBU
6KBtfqvecnZkGxs6L/txUi+mPU5kZOUsQFYmcwbBqie52GZ6Xwq5g+zTDX+bz6pjFt+qzuWvtbi1
fByFEKaYAOk1mzLGC2+bKsOWi0Kaegsn+N2bfbXtjaFLxyCdMgVukmVj1YIhcFylVRO+OPXWX/e1
vFfHdCCV7Ya3y2/Q9Ib7+7zCYHqCa2fm+i9tkSWjHu1et/w+uycef6JCYEDWiu4VwBcQaj2eNbyv
ixc4RU98CqLWKEUGyLUVGxRajXgWj9ow6O8EO7ba8W7C53lI58kcYaDkqwsRqnTi+xG7lLslTauX
8Qfr2yHYxF3cQqS5Iu/4WopB80Y50I5JknnHPd6YVG/ax3kE9IqQyHnt2FtEwI3kLsYT52Ce6rGh
V/wrjL7gO4Afrz2mwrtGMAc/6Rw1tl4sj5wos6rNUGpP6qzMPs8UxtnCENH7WUNx70yl3ElwL/pK
od/cyol+sbnijazUAE/ad/kAAOiQfNHyVxePVt3PvTn9i/pRNYC43XzB4+vp4uxubJFkXFHJ+3w8
1YTBSaakOnK/T83mvjTiRjnpQdX0OHzw08T/kGO2nhtmTiRaboTcFM7jmkJb9zX7PVaMH23IG+XI
aTBzc2pqdEEsyx1dbH1A1oOMM9thr1+QGIRTHbqN3/SQ1U5KC8W+BumWpEw/Kyd3mWct2srhnUtY
KThK4CYh767bpPHFwCV7ekiSiLJOOWbOcwK3b1M9PvsUMcKhG2uNQQHZv+vDF2+lMTZqH7tvmwj4
AqUxnN8VyiH4MFTxIio+MfT1FmLHEOm9q1Nf3R3Bx2SMB6IOZqL4He8hnGdACr+WpUsey8hsdDy0
tDEDwF1loK7WdViciy8SkMzKfY6y3D/pgr75/FVuRTXFindNbSTSzF0NPcLmvywvJT0g+53hcUhb
6pEgJcIRlVqR7FgXD9ZotlQTy8j+3nhNADOW7aIsujN2Z7ZHrMBhZFLYp0TqRw15qFcQVlrfYbd5
UTQhr6oBt/I3zasMviUtWAYaFQG6Bq6UINI2+Ik1K8GQSbBG/cqCuFfyqtrNTLqRLFr2VswsabHj
GqXOiYZs4xLS5v+6hLk/dB0V3nfJEs06cjRCepy/Wyiin2dg7URAuIZ/MwP1+ZPr8OZ6+2nEQ+zW
B0/Au9Qyz+/gWP7J7WDvZKy5KA9UC6s0xg/p3di7n8GTH3Mq2CzLq7EeXq94IA1QRrBOIyHNHCHL
u9/CpekOpTwtgitbMblhSR5FTOKu2cZ8/hzL4fZM7jIK2pzeP/9YcMordvlLVNxmhY9XzMWSon0X
Fw9UGJYCcDm2I+vpwdAljJkQLdsigbyZW0Fm9XgC7Fog9qr+nZI2ct2yBHeqO3iAi4xrRc/W9JBB
NPDNqKCFjQQWSnL9TWb28AgdgHCbGG/+DK/ur+XuhlXbQntB0K+cimvS9Up01hF/XRa2P03Ke8jt
zetIkZpMQ4kQkhxIBxxXNyhl+B/RhZA1OqVlLdFBaOFoHkggtJzMqDuVBwE57mzBNty8ZISYc2eU
z28pv85oOpiV8pBRJe4oI3ydiNs6Ly06vCAzLBLZDR+dZDOaQB/zCRJhxwSU7jm5LRBSVKMbyVf4
sFNDhg0RKX9Nm9PDNK6f2OZJAOzAbnRGKWHHIGTXEUIq008UTdatQTEgXc0sOKjzIRc3ljX5VSU2
HUN9vDl+xmubJZ7CxrpKQYEZtvbW69wGAn57VhF7zfQ6ZYE+MTw4u+rUA5tovieZutXkq5s6Bef6
tlPBeYb5en6wphHUFonjTunBx5a8luNybr1jrauxR/wQDG1Ay5FkMU+3exn5rPI7qsinpU6c4TC7
KQOpTghjzQC1JpDjJVsHCQlks8m4+/TLOO51NcFimU9HVpJgddZoZzNaocJXcP+hthSoQiUfJIE5
h2rmYg7utz/YWNox6eaFGt3nMzm4CkJvAq+N+u1NgcHi8eERJmd3MgdTe3JjPVkvdLZCISKalWYC
L4qfMflNplD89zQUf0VQMDSH5Of7EFyNJ/O0ofMqLX+q07SAND6d99NOEAVCOTRk5hMbHil/aIgU
glVJ8vLcbgjSWF6SFy8wWnvtzcUnHsuIGMk8Gme7LSD3RrFVF7u3l1/KWEgYq1Z24Mue4Hu2Kzox
/Xg3m/aOO3wEK3LM744uhuQV9IiS0vOa/OrYGbV6DDIiG44fqYCNNB15zwYvwcQbmdeCiE+jg4kJ
JAUfkK+LORsAYINocCgtv7outZTKvnQkLdEm5YA3tCI8/6//U4cLlXJQvDWW2xXOG13jWql4O1oi
3BSPbk6Hgw3n6IPuqpDk2HeUUBAv4TS/CbCEYJ62kireythvTdVq+bmyIN2K+DnkV7B6YqZjgZVw
4X0eaCVr2YhpRWHpCbPvofo3ainfNVzLBM7WdAwTRORU0jo90h1Z7gd78k37w1y6PUKHy6nR9bd1
p6OJOAeZEXBmWhips2d8Ux/6LAsTk19lNDK+Hnqjfgr5K6bY4whHnD2zosuBd+M8G7oSxofgiOgZ
gVHAUO+y5mItdJ9C5BzPwMPbdo/5rmLV5CjY6MUz4AaIFQTSOiprlSkVVUhoOLabBJEK8iZpE7JZ
985KRjoLEnW2sKPbaMxOuMz4YrPSLW0IMrUweGNTNwUuF3G+lfNJWPnQ0wv9mCWyn8aQLU5ZrANV
t7+tHe+/PkNFYLS6/eHwXaoz5q6h8oTihkAxMsCGsVHhHAQF/cVMEGN9FQAqao55eYJucFeUTvP6
JFgRQXjF1tXq8k5vbG4A/fZ6/p2GXfJ9yzwwgpzZnvgh/Ha9YUCt4L+vwAtfU8Jd9rJVC7NKGwd2
bCrE7vHBaGCJcWjMB+WvXj8pUscHQ9PGr9GSuPfaGihp/SjffFrYXz4T99UeuwmWyZTtZJkujbRd
3ApVy4o+ubX29+3JhsF5cSq8Q3zexzjvzx+gjVawqLE36IRif51g6/6PrvJQ4b85YaI0Mz/HjM0l
s1BoF9+XI2Gb2ivlvZiVV3bXnZE3MnyX6S4UQnsC+W2ZwBKm6EQp59f6+7FUn+FrNulOsDZ1lzBX
nYRRUW9mSx6C30K1kWKFJprRmVf/764owV59F0wzIzVz+lo1d2jFaJzTrNwgAzh2XnSE/z4NPJhY
2yE6qX4UOOMJ4UVFjRt1NIetC4P6G4ubVm4MbvVjzVPK1ox+j2tn3fIDbSMd0J/RWw2wJk66/K+B
kv4vZEp+hfo8L3ossx58LKtkBno4TAY+8V4/2xTbX4kxTXKmR71vTOO51W1hPHRBfwi00G3J2xG+
65SY0Ljn7iSQu4xlUS88xZiO48GOXib8jPxfFr9qn42qnDryJRequEcQrChi1SbgsPVvnL8J3Q3z
A3ZsZsnhPEoq/n3GFo027yv9HEpF//mSKmooCpCta7wCAYJqP2HLvwbgMT724hJMSi3+p51rE93v
yrTjBcizGDc2sqCtDNM1s0ThcftoMmOZ3wvU1bflp2c/YbNVIcJFH6Ptd97dRUjcesaGFAc9Kayj
mgb80N0PDjZVRBeqOvmsOz2LzPOysyu4aGNyoWvP3QL6yD8Xc8q4MV+Ano0JcTGZFBIWr6IKqZfU
7JQeoL240ek5n1yc8ioLK6SdYJmk+4JmlToRxTOYpDTb6vgXWn2g7TR2ZsJKB0N4rHYCdhPoXHiC
KMKitldPeEL16U0OulqhqF3OxvL5XijMAYnu0+kXIT0VBs5XUKl0HVC7bxji+V47Wkrj2XXGQujO
r1MjSfB7lHpJvQEehVYL9Tb0snHI52vq/UT0jGPVd1hGJDwcFSmpidjfJHY/Z6axy1p/X/xEqkBd
Z2BIBIQ/fd3fhZXOkkeimr+/1pWhPb3cbi1lFYlFFG/v65XS5jVpt9pA52Fb7wfOnmvybzw3G+eb
n1yeG7brO7Zj/zbcFyhVVLJBwpsoLroCsHKcSoPk9aP341wA8g3oIXniYkHZEBVGhpsOoItHOKlP
6hVLCxyPMqawj60ahOcNVY3G0U/dmU88GdKo4GJR5cD5dP3Fes3ARcH+ta/FzWSBV0jxv/6C8zog
tyj3i/5YVQJSkYFetFmqtCMMnsggyMscH034Th8RV0bdsnKN2y2usTtzr4tN3eja9q4pfVg+SKex
uX5T6YKmc2Q4qd2yNM5DjivAqCoHsULPO0qFpZqPGqTzCTiPGhmTvoTQMWSBK61wgWiGAeOqiZuc
nf5uwwKFtdat1KsS/rWSBxFdgmDCaqcvALqs46ERVa0tDqdfyS3IwqObLfkEF/deyWiTZtTAarsM
ty59fh6xhISjvgHysBMCSsE0tM5S1p87fhM68YtGCX6m4XKa3RsZoz1713Gyf8XjIefhLQJb8A5j
DrECn80xJmjNP8hkNuMDdKvbdo8NaetpyYjKeA0iukUaaAbQktsNMyi6zt30GjBbgAzaYnX5msOY
MdsJr5vT/D3tZAfeHidsLsa5KUi6mQKNN8BJsiADxTP61a3KAZzLMdl2F9c0jgeR4kGYliv3kKhc
6zvyxPbF6ivctYWEzL4oCQZSTuWqThAmNUp87LR/ekZiNSxY4h/RpNH5LIk6GIkak9gEwuTYdSY7
6032XCBl2qlRne1RAnRoBcfwR61uTg/Q+DXWfHPcjETi3jZ7J2qwznOuqM/AjUEdMKweFJ1iI0w3
BjlsYeJ+VGmjTBwQf2M/aSEpxZqfhM1etrzlz2tj5G0YEMDsUG93mQqgNc2Ss1WPDjfPjRpuc4Yi
b+mag+A0CmAa589+UtElwjTC/uEBBMQm1yyvTwNlhSnyUuU2tlvCAiLOZuBFkOZpLaBpEPDrOhBW
Q/S6muEMchG4slk4o69/q6ocQLIl2GJNwKR790JSe05g5x90coqI2ngsKFQ4D7MzuE8JoQuUrYGC
wHl+artodXDeFao+fuDl6hBuueAoKp3PtwDWLSiDK4bAHQI3p7vjWCnsbcg1xsXcaDJnlkOQOn04
yz3wFKLyKZQLH6k4GALa1CQswPyj7G4BPz3EYJXUBVGqnB7H/N2Tr/Ez231IHPebbbwvOA0GUnob
29fKJ9p4oYpow0mfQNNYvdB3VfyJifzPn8cD/DwNqkxEzx+tN9e6JVswAF7QRWhBrjmAhgPhqpjk
J80aNe+C3XhI1pWa3b82Rnm8RBbr6/B9pHLm3pIllqgh39lCbRnZkcX0LrMpTcMoD0MgTREuhUXX
CrR9NZuV+kzQhMj7OJMtMbmHqsQFb7kvVZOuBWnsTuZXvF96SDf6kpVGo94R8d65C2FIcwIUs2sn
4yskHijW9YL5jMhx6Sn3hl4j7nLNRPH0j6mIMfqhrMpaGVjksO1IfbBdYZrCHHRUrWsLOnP2k8Un
1J2G2N1xX0UIjBehv4o2deb2I1jAW5j5IjfePPnKdRUzl3f92G/fjkK8fBmQOJV6uxhveZ8j7o1G
SU67VjBex8dTd81yK9ZvEf0Rkx4Dahd0xE9tRe+6OD5YU5wmZgXQWVWDncZWOtBetN+OLN+Gh8L0
c1bTV84pxSxF+aSBrrsCElC4bAFlq+tivVZCHTTkoDBXz5huggCpZJjFZuJS3EIR+NQnpNgbs4OE
Oo1QIwSg2j233jWdJMlTz06AMY2iOySEfjEuscobMjNwAT1PiUwtVMUlASoo0gu1iO3H2cdkkndV
TmyE8yW+Uji+efP2aRMBXtHKGh+pOjVu54mSoFSxJBsa3y87HiPGZgljT9jooqxVdEk4Hs6j85J3
irYtcB1eZjO0eoqDMUclB+CnFMgr24pbKkY7Gd8BM3T6yZmAWmtkykbzWZJ1DCIhQSFtwyHInl4V
3MiQWmnuAQPD7w55F3OwZhFrKBHfptfNn2ZVWxYN9qfiIvox08aEZpVyuvd0iL1PerGWWukUMUSz
3Bx+Eg6280szNoDbYf0HA/CbT/uKKWilAHxzxVX7RiCG3Q26xScpVMAgvVCoWy2qDSShU8r5J5Od
HQjlmUOxqDLyKplH+8NP9Ta5HHEbYscpmmvoIdjIvMu95yrfHd7CZVJYDVif94i+MRppxjKmVoox
ja1XYPS8lrWRWJaHiIPJdGtje+0rT8Bwww2WkxF+dtT9w5Nl/BvRrvj8MLaaTfusU2x9pfRvcHc7
V/EBgQL/mQrKBF9J1ST3bF7Lw8AeHXK9zoXmGdC5ciPdCWeylrM5bWJzhT6fQS6MMAtX5j9u5X+X
Jn+LZxXUoxiRa0l5StvLczQjg/K5tlDrBJ3IzXxJiIH84bWP2h8qPpzE7fgtacJEW/0nSzfF+VhK
9Axvj6whFUrIM86TUXFGCoZRthvnTYVg2TW+5JjSwP0vY7++6oy7Lf8vK6UVaxtrLifxdoheGzR/
swoteCPBu7lvBEFDMeqvTWXhmkOnJsdFn4OuTvAhRE5HXSG1Gl2sLnM0u3pF3ls7deF18vvg+MOB
qsc3gkzgEWN7w6ZbjD0VSBUwOcss8P9I/fdo2WR1gAUJWNLRY/S7sPv73rhTZdIsKFPNLFlH1kNx
XzpminKwd0RxR04iHfZQaZ30r0osjlsH6p/98SzuLWOAd020K8aQHaO30aZOUFOnDTY8W2vsYvsp
lSRJwn0/KXYRzhHU3ns1oxUOFVlH+N1BsqO4xtMyGLZDHZAQV0i/3erzHzqgwnvYLHkAxbBD//tB
y80jksz12GgDayC7m2XT6FiML6qbs+LKRjtxzc1znI4bo3maPS/fCzZ00h9VVqbaSTSBnzD375lx
rr0ZGxb2VZdHhgZNxCJe2AsQJ2J49pkT0k7h50BlHWV7YMkycw/G1xT2n3FA0ZZ5yOVh3Knd7wC7
1o0TQPyShnMgaMsVdhhMQLtoBZO7bSFSaWn3yvj21bFGx+YsV5SpAdGeqM1AY4DIx6OFrpNvpfuJ
gaSXHNDKA1mDhdlA5+y1Ya1OP2RKYI4k5T2hAqlOZWADo6c3ZXpQiVP+S8vW+dMdOOGfgRlMwkGa
SJ8aU6QvdhtN3lSzy+IWsntKOEyTWZBRjrATdzpk6yugLz1ylu+bMOwaI06L5LNLz+LNUQy1yH0K
ngHnM+a82O4LBVTw6DJpqISd3gxXSXkxYVwLLxxskTxVMeDb59mtzOgtBCZVyECoxp0JlejAHzzl
veJOj/tLw8mdrNsHhXxoKCtFWCVhoWjK2/cocfHCumxI2lTtX4oioqfgze0A6OzlHkOxrdN7Nydh
UvJPegLXnagiFDy6f/meKpMe/ZOnq0O69kKT67j775cKeDpMyAl6DggXG3t+scBFHzRYufnowWGh
eQ5uQZuHnFSQrbD4EdJZW+BMgn3Ioe4/aLmZsnZVIwYDcuuP+DDpzMDln7VBhtHZZvQw3BDmTm8a
r20EbEh7ST6X+EW1N6Xr+iJouW1tf6sL2tt4y2clbIL3rQGAWbyqCUYV8UumR7I0gqMsN4/dSTGY
G0J7mQdtcAhhA6F8uXvG2RnF7hDIYUVtK/AHqiMQHn8scTcBBm5ZekunreyRcTkdIC2iBv7g++1q
i6Im47z/vzXtZMvmqaUpoAkh9k4zCNcQJugrGWfSUkMcNOJqkmXQ1ZSHCtSgFhgwIncPRXDH2uZK
J05uZZWG0mxFqH8vzD1OHbDnWAl/Uhk3T7pN2qk+5kqMsIW+Sjahlg2BLF4mT5kTqBlhnlpYVB3z
LYDNMCIA5pK/+n7cLDsEmPJ1ZGXdifBR6qXPkCTH4SCst9b7I38j7WSu5ZcYTUs4GC3Lru5ceyce
qu8AvwkJejeYL6lj9dnWn73SPvTtYFG5pb3ZyP1WtV3t5q6WHpLHe8uxI6eB5I/kFwWGvDfq+qjZ
zI6ptpyrHwgg5q0aFi+uD0J712QurGN5erRbi5y6r5fx4jqvRms+JflArDAVx9NHMpUjtaResPxb
q2K7lsS8sQBYwvXJKNNwsIWNHRsr2vEnnGo9t3EUYw1SS3n3xIE6lwH/ZsEUlmmUw3Pm7LR2y/OX
wovxsy2IDjnk1Qepp4zgHE0c5ZwFb1Er+oTDIoYn87OdLmyYK5KurJ+WenIPUv4gPju5VTWNmJRl
DkbTp2Xa//nuj26kTFAyc0s77etf2PMGawDBBsBSlABb5hnYXEf0neqCtax4AwJLQDDcZB4y73Rm
fdKt1cY5Wuph7GrxoIGOfHfyjmVEUQ6esr8T/1odu/WPWbSOiQEZl4D5zD5CgWs9Iujic+R36Z/J
BbIQI4gW26QdnOWrDpbK2mYUtlf1GVL05c5kwRj9sXMof6jgTfJx2Y2z1KcGlO2XD2xoU1kza//Y
/e4jeK1wcfGro99cWqC9L8V57bdgR3+tihh7nRb2vX0XPYv+LuxHTON5sgueLscWp5ue53wq7dlt
VJGxPI5UZlt+Bwn7iTJjnxDjetU5AGMedKUmfSsZnZksDsxjKDd+l7q0DFmvEwIlylUGkOW2nTEL
urXebob0Yw0ss7pJfi31Ad+hTXXjqg30ZaMHOXkaVg/Zb7iGsQc3R1XT/SDOveRJ7e/GQeHP3wU3
08m+8yaUqlZyOXKzVGw39ugURrjKE3xuF/30YyK3UkvkJxEmKJtToQ7HWQc1fqKkoiLa6VI7RviN
4tLpJb+lnjSHGHDZhy1yQQ6DkXkNzFWs1mReULM9CulrpnmudqDmU6stl0h1aEvP7bcS3H44ycHA
SYk61C/1/NxZBXmB64iXq7Y9Mhz+05YqYtgPxYrrhM3HPdLinmkX3bdYLxprbs/bG0YeIMFiy303
pOIWCdUMoQU/1MQ5EVhuSB/j32n4flEzrySlCOPYaynV3EihuHJ+4VkKc0v6grmYWjjwpsqiUT1c
0Xrsm+Q/lXzeNIARN0NY2CWBUKIP4571rum3ZCNaySmZrp5Z0/j6ML5IKMOZuNKoia5X42qyivM9
bb8f5JLVjTcWlHzC95wJHbO7Inw2tMrq97/4VZ0qFfIx3GBe+m2OswMQPBnMWi4GXVMlALfic0mx
Iw/C1nMqsBhc1e1welrPWwQetISLoOFdPlPyvzpP4La/0p7IBGolq0rYPcaI0C+HfIvEdJE0oEkZ
LX0JNx6Hy0OG5MGmJvj7zTxqgs1/Ry4ANxfjpJwlI8a4Edv79M/BOB6AoBmYKXqtUnyKX5kpuowt
zW0ZjFVvAhxC8pOY3MLylrg+zbHmnOJypsMorxSsoHSTneOoo/QpEZs7oZdBT1x8TPt23oW+quct
kQJqmSieNkyMTWn74Gi5Rf2BuDAyIVH9Dyhj5UQL12saw166Ea02n1DI0m0bfTbqP/O9VhlBYrMu
jZz3h4styRPVhR5hq6m+OYRq5Qj0cDBgxhjgC8MSCGL75qDEaPBB35WL8CutPpBazUTkp5GFzwNK
BUEKIzwk9ZFEGuspgKDk71Z4riLYr8yEfZncs3VcX+NqzlP7ys39GM4qJ/mQzKW8zzyzeO7KGNYR
4IYFA1DSgL2uMy2woIZxy7Mv+vKQrvyvcCgdfPSVzLlfKKujMwm0jc1uNHBKbuZhXrG/XjB346aY
PNeNKN02TK4tUErtBiHYN5mLNZ49GDHql99QNF4GXA9i727/S30tGzwHPF4QBpTrHsGwwNr3QCiT
8EanHOcFeNBfv7F9QOUBHm1+GguNsQK72UeLSODII9xFy2gL9imL509CC8TKGOXTNNIEEnOhlVS+
O181/8NoaXqgx1BnzFJsikwTEmh50KeRwJr0Zj6J5rgtU5Li8O8/wZDZNvqWOShAOZ84/8fHOwpd
bh6TBogLes8tEhWAmOnPNZPbDZsk/0tGp5lm41a18VH42PgmNfECGkfhsmcZz/xmS9Pec1IQDXrQ
UX9D8Cf31QPoJHD4E3wkMYP4Xpwm20LBSxzQv9pscckTzWshwefCWSqBY+O632YgWfO6aUMZErFH
QyyuRhPyNXVYekxX89xMN5q/a68QjCCrf+mwozri6OcY5qzP0Pe1GcUYF5VcxTwsKCp2z/culf/f
HCJ66J266qOji0OrQiASMtR0bvZvUPOd6H0ju59oKk7NdTsT93yeC5Lp1yTHysckBVUGaAMto6B+
4MI2ILQwMtATHjvEy2SLxX8AC7emijeTGSV28yEGICnh5x40WLkBfIha+RbvzYmy0EvXk1X7HpT8
/7fONoYERZc4QdyeWMT4GPVeDxYveewtfTCy4fiJ250v1zSku2ZVoR8WCljBqtKjBE/WrjZj+TWu
r28Ydrk171QWYd8XYcPTOXUuIgP5qqGLOkItmebY+kjSr3Bac/wDwTHt7kwPWoT1NXbqyv71Sfau
5oYFIX5q4YY8vgLwqt4rPJsbvzAGC4QmFoLqBthFhFlGBFN4nfgzvfrU+0pAANtgJ16pkr/e4O2V
c5ly8c50h4/+U3FSbtweBzI7b4j86TJqUPW772B7ZTkS/C2Iw9O/qTCa9DmVIoP0gTGYjm2AZc9g
CBc9nzY3ib2zduQ1U5NlVcyoVbiSfMk+GIDsKZ3ebzHOI9OD+Soc3WSHz7czK/1figO8GaALWzOl
MshJwuSa0OZHJG8g4sD/1sbsx5Lb04CrY1emIl50eXDNcahQFO4G1FiWrwR6BkA24h93OzjUaLWR
za4zD6moXhvkVzDZslxC967JQcYd80jEbhr5TXZDmkydBNJ6qfA9tjQMe6mrcrW9In1OS3NfbfWm
HZ8UdTpEaPabIzqYvkExDL9sZqBLmOBi1hf4am1nu4qak8usv5GbUvXa3ObMyn2O4WPwDS4uLg6Z
xIZsljIfQb+AZszQbk74hVS04pPYqoMvvMAiFXr4ixGblpJhq8+2y3t5cVcDcirsfxtFoeJuETq1
1b8FJs+24b/LtvyxYe+dNAMPLjUQk3Ju+UHhqLL6dxXzK37wlVSztidgpjLIPbzOdmAUixx0MMQT
e2ict9rwSDc4lId/QSuuZu96bXkSHKmav7liPj8Q7XJwXYF7H6WGV8FV18ZZcA4z/VDUf124NESv
vevOu/e0/wfXIDN53mlD36dNzJ2cmpc4mP4Y8x+vnrrQc2fOYuVUotSYvaRUwCpftYFLLC2We7EJ
ryRxja4XcrgVi/O5RM57+HW+f+RNqjCtxrEdzMIUiCFFQxwu9sfrDYoCJB+riKCN1nHmCamdPgAU
MkaH12zgjNcwShait0DzgvIsCTciuf4f88uDo1DZb+uMU+DhxKxbvRuhyMQ2Hf1sI38lW25w5n1b
xHGo/w+ztzcUIha8WfwNYxA/wEwPNae48ZySIsPCQ+sZ+6WEOu+mWu9HycZHNerbMlyxJ8LQuJj0
MD5BgSybO1DKTPX7+XmrDBfn8MjvY+2Pi+8Xb8B9XuwCHdQbsh9CjGMFG9ZhPzLhh1qDqDwjJXOt
vAbaEXedmBGHZKZGs6o2IZ6M6Nv4+YG5cAeMFB8JUvNGerrcE1L4+lgvSax8MJlr4g8L7WNYAKXB
bvWq8T7y11E4zUI4C21wbjnvPwNoe2Cve5yh6cCQdzUQdY0IvbGKaRVfoTODxvEvUUyRUHifMaJ0
1LqZOZ75tYHkLlOiy1w62Z4VW6t91BrkMYReu+JxphXmTqGjsWRq3zcwpXyeEfuY/dhJc8f8invd
3U2e2v0Er/uwq17BbDOhW57BdDfI/9Yqans8U0YZNspNVvCXZ2dSAt0aFDLFU5sJETg+UZDe0loF
93rPtNYY5DRnefi4fnyz+0d2wuvQGwIOHMgyx2NriOQt5ElmvVjq80qKvV977w7oCqPRdY/ZovLr
OtC5orb+dlDbnzxMyrO3hp5QFRSe+VG4x748sYi+qYMy3CK6JULgZdRF7TA0sIKvLcNkBsVWfEoK
uxFOwfRMrklR6Bo29LpmwE6+2oy+SItK3Pu8ufV2ebBskojcTC6HyYVxnKWscgv6K0iSpLxDJ2Wj
iveTS+wj1yhQY+6fJA0qLJ934DEjs/Lj1OXnDDmaXdAGnwzrRMKgla6hbhi9hr+OzniFQ8kEv5fj
L72qRceZZH33vkSjGvMcV2Y7Pf4AN0QN13QcY4evHGgreQv/pvsV99lGZp7HlTIlCdBjMjCxFIRb
oiIN/T6kYWR5N5oyw+r2CBlq+W3i5g0/Fm/Sd6GUhBUlKr4CuBgkWl+r5ThTQCu8Ks3rkSDDXHjW
rjB9sZrVYM2GsfOP923eIDnlhTs3uR4v2fB6CVPdmAe677rybrjsEWdfgJ+ZK7W0xRuzH9K8Y48A
vJF8FLE26VS49l88OpvnEBT0QxAVMAW0W3Ur2hWFJou9Ryoi0bnSpKMXPM7UemoUiBkTjhL+/p7+
N628QvtG4Qw1GU5u21LOHjIbkG+tQ1AyFUZqVdO8TkHyOc3zgsa8I35Oc5F9Ix3SLYpk05Hojwu0
F0e/ZDr3kUfOyIkI8a530uP2tfYguoMRxr6GCofx1Raj0hkbLIp+P77j669ud3EZC0gRh05A8gD8
6OYhdIjY26cMAYPQq9E+hjJvxZZJfOHGmYeWbG5c40p062GxOlzO2+aQsDKkhxK2O/tDLywPYuxa
9aHgcQ3aSOufvoXqlsxW8RAwcHiPvhTWw4pvtNBw1SRcz64Fl0u73IRLWHpYU6FcbnV3eZkK7cNw
AOEhCgjgP9Nh4DUUvRsz8fCsFCbHcGRWTNVp4vRu0WPoKCqhEkifpoHGZ9bpiTz27MO5uJj7JJDm
mu2gkJcFVpkgXjHvjGLbqKuUvS/CjsAqTGMNFY63vB8IgHPfKpKj8Qxnru/U56PZnmtLkZJ0I+FY
vXAy1ue6CasylqDQX9HjtEJ34W7BphvkQ1vuXhr4aDgHuU/2CoqFsCn+tFXVPD6CbN9WmAIaBc20
/hIhymkbsIGQnwR4+unQteFz0yt3dvo54UBCE9uQGZ08uFwdr3LQp8YCd+LT6d4UMTDxZVkZVWmU
JCHgGnyINqlcM3OHsSAeChOeEuKkVIlunlmlMKzZkAxGRflx3/G/7+qoPQKXUk0wmopLCMspYIPm
KKhTSBPfIcb6rdum1D/ojCN1gFSfsjtLgaCOLGQ3uzfcst9LlN7toxWauQfI3JRFjVEyTUxNuA+Y
958I9pue4XeGipMAL5kQn4SZ6uczTXWlsm+0OBaWFkvBM+TcmuLL4ZfP57A9wvJGHsUcRtp7JLgd
OQtM0/CRAWcHFkW7lDenpI2P14o9CL4m2Q7kClcp9rqYY2vXDxIwh1gd7tdz8IwdNyEdWT45xls6
f+OPd+/QDkZke1wzf9RLLcQx/c8AIN+zDyO78J5dc9edGIT6URNQ/dD83xJiiYxNyIRQBpcGJnLw
Gy+WvLgIHfZf+qFJrlYQkGcXVk8XImZjAon9tKrnR8Zm8y9e/GVM8gcx9ZY2edfmR5s9p39wUB7G
VaG2DYlTtZWCS9hZYV+XQBdjjsDknn/57yMq97Zfc5qodrp/8diBglDDnv9Zelg5e1aht4Sszw9/
CeZQ0HoZW5kTmEr/GfwE1AtT2Ip0vHRGGrTmBTVzniomMBgFwwK7L3707WzkNr0sFRAbHSyqqekI
ErhNsiXmm7S3lIGuJHAN7QsLRw6wkiBhcR53hGfwiToa2EJKtT3JwhqNzdth0dAA7/NjRXVhTSMz
WE639pw5dcAmLnH14fiBscnQnV9KM/n+mQsgq9OFPc3DIy45qVXgB/ArRFA/I4TgFPLAb3rVzGMq
Jj11Qqzj51vBDubeSQ6mC0EBBQI2HOeHaq7zzLV/BanScRSduz456N/X+pOVkFKnusCER0xTKG05
4DnVJDEc5J7GYHrE0X5L2gEcTwY635fYXa0OB3f1W6YG4+A4I4WTlEf09sJwvmjRPOHu9kY9A3eA
/W2ZHyC6Cag+ZaXFZDAzexyPyM9qqEid5u1z7kc1X5cq5Hf032SWr/oX4j6OPnxza6wy7UClq6JS
XpCiLiVXVeBWsC97viKBfPk69tAevdy5DzV78ZwweKsXeEfDsUGokfgH6w/0kR0DA5VjJkSGbY74
dIGxsCriSrXsbDiYejkBYApr8C5gh5uHNv5Yq1prCimb9aVtRlfZ7x5TjU5kDOCE8jk8nTAZE6u4
g9EIwQSwojm7cS7FL8yIyFANKGniRSyFH4nAo2vZvlw3MyRF+yURI4ZgkSak0VZDTsy9P5sFuBUR
g/pn7n76BzmYID2Yg7vCkr9PcCDyJqhrLFVRJhzOf0LH5HMs+BCIOOatE1i6Rz2OwFqLySKBBdRl
DCQr99zxuc8rJKM9z6Y9Yw3hPG/NiJereBBtxtmrxhx3tcg/MfALO6Qms6mPOuHQHgOnnWCoAKqn
9DQPrXFoViF8sHG32+2uxRGSTnLBUNjKADulFUDMDegdFGkzMscM7zOyCetDQbvHPm3WDdoE0wMl
awaDd96ZAQzCwp0pqhZrD+dR+fks2IyZ21GCR8tuD0HW5EqkRObNlE9vBibvJwmNdR1VLUi9jC+5
BAJgOxR8diaBJLU4qsK1zPks7ub+EoeD8vkAPphngw3opCi7vW37b2MF+tyej9+Jh3IpuC/2U1SO
6W6TCEDTR4DbXPLmj9X0G/jTjebAQhvsM4MrHVP8u+esdZ8HzG9qxhfb82gGFQFUh9G29pvCqgxo
EZHu1EaDYA0D9oqAvyd2pYc4h04SI+TPCafJhhfeVNbTRaTRuKzJVzkJ4SWc/HMC3dd1xgZLDkXm
+G/FVk552DIC6HBwbKnMgndv+YomMCzKyFKXrR5aaUWQN8GYdTwGWTDK3Ri3z4tKLxUM0fo0BZB9
cR52wVq6RG5xcDtw8klAKmS/R2q/Vcd/l2XwAaDHkJjR6YsS0IpaZi0XuZipg/E6O/K32pZjJdo3
lzv693hJwncfUs6wcGNlxR/V+xLfp5t/xbT+7V4Q/kZdC5/jxQ7vZkQQos+vUSSGzEhOyXRrRuA1
qAdueb8VzHW9Fn2rKUxrmb6aqQCPFBvvGA4g5HdzuEJQ5KsbbDxtSIFmlc9cfCRrLWIMh8zt08mP
J4/ZTvIhXXApxP4bBpG2S7v2APc+USVc6IzcOAFpM27LZDb2UCZtuGEpS5CbquNrIPd2MeaSv4xs
s6uFrmLUwm6QzLlSGNJJCB7PqYnD/zYWbpzvr+kI9EKjnpfcGOI7mE8s2+khw1eao7bfao3w7U6w
R/9D4k3q0vZ9meU9tpchvPesdsamDCBpG8KTrwDGwVmJe2xQnavWqEafNdYW4SmdRN78MSS5xtKc
gVHTR2SkhLUNLvgAT/nCdZ83wjEsYAiEFTJ4SDSrWsFefLKLpiUVpcXbCPZ3/3EkO3eMHCGN42Q0
JBTpErX9NR7m6aRYoPRjxEbasYhWXD0OIw3wqrXoG61M+jgSa5irBr5HQBIQlGP736F6UFgvR05S
h8VRTG4C8ml/+uGe2nYAD/umtO2ZS9nqLLb/lVTJxDtfW/BA2QfIHFUMYY2hGijWWLZyWlWWVzzw
/1nj9Y343Z8gotVsbc53WILhzO7MlnlOgEKYej1IIuzyDgKRvbFQZ8vcuA0Eq1Z1OpWBktI7xVgk
GZ5u16ApqNaBYDTpwee6/7o/FB4pYzSuhiX7/lhSwViJs3q8ihhMEZZl8MsnHnCcsY+3ove4qgwg
9G3hBr49WA65Kz/mF8zBzMO6iOScVcQD/bkPsYwaZd+6AJMSFfOAebhlFIjy/hvgl7XZqtTCEl/Q
9BcKFZ+IbOAIoiYn8J3FrUy3K7s713u/wTh8NV8e+jtRMz9xKTL0vl6zIoYWJI5Mcu1YdFtUh5wx
HoSzDvjve5R6cNiz4LYhkfa26z8DV0Dlc0OALvcHb4fFYDzTdtaU72zpo/hNketBaFQngu0crgUt
gKnBXzbQtxJqG/tCjaLDieZtElafQQdDR8DKOvF6dbxIuY4hIz5bhHhOTUAgEJ4b/WBJSq2rav8I
j7e4YZWXYMjiCU039eyayHrMGZWbgLQOW61qWDutkUY5btqqo29hX7w82D1CVrFATMSSFyF46Nzo
lnnYVEoQvgaM6PWnjxiSVo3FvoYr4xQG5YyCAlm+AV8QYseXGW4I1t5QwfN+nSk07ICmDr3UcJ8Z
XOBom4PpwawQBiAm4oiOURqFBCzb/pZHrQItvHm//KhxEtRz26nWBDuhElcGL8+IMJrp95L2rv+y
w2D206pkRGwDoV/q/TK0JpsZ9OPK4cAQTFtnOguHr0AGoN+8tJDqWGS/21Ni4VEUgB5P/U42TKoe
i69LB4ba50npZ9OGSXX3zRJBLRsElMIssNOZ5QjNNYZKcs4Q+SDMSCj0SMs6gtAQLublkDvzwCqN
G+v5VkZywRgyfmWRdnSHBZsctKaflAKbGAh2c44MXgoLreINYWYckcjvYW5TOkj+04mqlH73NwVP
UyyH0ihkvXbfapX2DGFUnIY84vArnVn7nlKcPzx0ksyAhVG0YUClOlOZb/SiZ49kzRWO890nfusb
L6bt/5/jYvyahKlX7Z3F9Jl6qqsInjIEgewPTc+SNIVDZa6CzKtNuQjNcvfeCwm3DJlGRGmSqCPi
VfCq8kRR1+ui2SFdqTIjRQwPARrURwqw2JDaziZOoRLOREYjmkh6ofmhlQRsU+oEvpEWyxo+LKIL
0xzXhZ1qBiswJ1PAT8c+eh5NFdW5SUvmyruGupDWKCEvnQ00mBNUdU9wSZFO4P9sTBQv4B0j4csn
Me9K2BTSffr3wehWxgyF7ukCyPh37rAKOSxnljMcRIjxv6x2M60CQyYLHgePIGRYYkI8xWXFgHsn
MO38aX5bZiZR2iE5qWrFUI7A2Uh2NHuQkNV/uzKRwYhE1ItITTkP0s6Um6cF+N8so6m7ivoygRI8
kF9MkRi60gZUUmIUKNT4gdkfNybcuGv99nUodE6Z1+ZfrqOIvDqsK/o1mRlE9fzsTBE/ze/Nk9nG
+Ww0g7DLzUN6Jj1xRuFSs6VWlSUyruHG8toZvYcIXlPZRnGHNVY2iixsu6bYRizs/GlZyhNMgrFE
lB4W8riOkOrIR4X9UKGCKDE8utuMC8cE2q4mTqJhk8NPmTm/2102YtLEVLGJ3SujJaqT13gwng+7
VwhsEnyWPwt6HC/6dJTdehEcpXB1I4XGgDkNFhbEnYy99X0ul3yL9w2paIgpbvaoQGFCcQqDr7t/
9MpiSw4L3v7tKwnfsn2RjoLDZ2VLx9G18JNB3W7ywrF/BrNookgTlZTYl4euYmgOWxYnHwGmj8mX
k3oa0HTngnZ3pTUSXc9SOlEhxQWn7o65NR3eoWwYD+L4OlUPNoHYkSnH1KfK77fR3etJRe9Xhsza
5/0JqXYr1FLNwkM8rgbPKNqwJDzQP4lvYW8vsVVx7nSHm5ViCR9O+VrH6ZtoP+dQEELgGuyuGLds
y6D5axNitHr38ADdugOX76ZVx51ezC34BiHzd8fa0YCmX1GfBpHpBgYW+9kOagIeUoSsl8+o5MYj
UYXwj57iPbuLEoX2Tclxwcp9XDO0vGC4yj3ckV8dpvu/al54KP9AzZqMwo3t9nqjqB9vN5855fcM
3Sfoug0ZnRqfJYUkLGICH9sclWI3r21aNxlOyV6OUFcWo4n/vLYspPHzofg5G11spZhnEUncWMOa
C250nRNM5RNpYkwrExVp3C17+1VufQ2xGHErrcUJgk3I9s3q3bNPb8PksA7C33jdE0m5Lgm4KBMA
A3EAWO0lczXY6F2hBsEKwnG0nhmVFRw/uqnlzMwqAIgRn0vY9pITr7JGsBPHC3J1Rkvu5PhJsOWV
/vkdTmi/USG4bExqbqcxTx/iy0AbZrjLNbkIXHa5+H+7f8Zl7z4f4qeyQjjl5vMBs7vWIIEKVW9k
MLa0QhEvGtWPZJXSC89GgB/5BNE+fTP7/bXdCbrRWPwj98EGo5/opVM5IwzABm5jZQa3sUwEQC2A
OmgjE2poOx/CXhoXZfN31bVygfVmNZZcjDC4XNEve0I6jg0/wPqTapvHpQL6Ku4QUDgQ+xurFF2e
yctQA+JXnc4RDA+fwEBl2E5icZJYoTrzEwuozC4LNdJyLPImMvVC2/veMG+LSiKkolXojAy/hpSm
JB66ktBYmajByt9AL/StCLvSaGPhYBgjCiuc/BvdwY6piYTQlL5v2uJ5XYvdAKgmtN9YxaoluPmg
W70lzgnFRsiQJT348KVMdmREvrKYGiGv3DCx9X9qQ8FUR3DXhpitf4S9o7tYFA6GWnSGNHbgdJsJ
iVpJw8oYyQRsf866ooIfIZDXcE2FPKNi8ljeO3Zw4LLTyQuDhVBEnWFVVH9AC4g7qgWh7k9pFC2G
ubWkbJBXAD/ySolbUta9mX1/jPmanBy9eZY3xpjGWGXwclrv7tVUjR9n4YVGJDy8OdwaJfevwEmf
cj0SQaVmMYeCDKS6wXFYzy536Z88kYC4g0aqNUrwnzBVMa8X4XaYES8gPwquwk/WY5brywYEOLJJ
D/RFVj4tO0uV2LbjDRJpdvwuumjvy0O8UYSHtRn8HFoPz4sehAFdFno/4z3p/wGMv2MloXKQWyV9
rX8Ol8gy5FYxVLUwlap4Otqkf/p99UMKS2o7CInMkauXmCxktRz21AISRpBQxsOMPhVH82R+dyCr
d2TPEv/iKH4nAMqoKarfdmXygGCdfhiLdKMOLwtycJu7W22Z6IsT+KmtEnKbWF/JqkpkhBQFAJqc
SARbJrkIbENAHrcyc2NYkAJhi4CIWgcVQI7YU5Y6+ACnaoTUcbFicAmMGYBrBm+k6LhhzUZiCspt
z0C53lvcS2WRu3rfyVeyeVQ/PRPHfQGzsjhbEGZ+txK8chllEK4AHHJxK4SviYa5RO6PZkHuxFYQ
g5G62LSVpWHo4MonTW08hY6gzkl8ONf4+pTjqQ6y0WbSqYQUNsnKsgUs6JWOhipgXzUWBMzW7ZZp
e2K/m9D/0VidDcidDJT6zeoU1rWQSWQI3b82hNUqPnvYKL5Qm3ISy658zJzGD+OEX3Ezd6TEZB6N
NQmiUD4E7GSvQQTYkT2kZvyV1B4+Hbou2SvlipL/crN5SwsKjU9acpp2CWWOCNoCD+zLd1PM8D8B
aHmWUQd+gdIKwzziKeCEfvCz9VGQyXOYM2JKA/ennTcQ5i0aPpaFMRCTVa277L6ozaAk3sdBqqkY
IjocS7Yigc34crtx+URg0cBzLhmnTPbqLtfiSTHTZ/dNQndfvd2hDEFRfwlBNEgyUdO22qR5DPCy
jQnMRGwPhnmWVkEyqYuhBrGm1dSRSrz3ltcP7bUoImPxzhpcHk/aX7lROvISwHQ3T2GzXvsE55eG
xawFVk0YKE+C7sutetSKZ3bKVepJYKQZLJyy9Mn+PTMNNwSpGYVU/9XGXUlwtjW7MVckTrJC8fxC
E+79WTtsWo9aPN9rPD47xvp8sdhpxpsWjRJKpQx/f/n3tVgvhXFfxRxWCs2diTR3MWQUhfUVBmW3
hn0Hp0syRvzjwwnnC1wZmevh35scQ6w0M5GY4X/QzfPEKE36V20JhSVACO0UaB9l1Zh1JTr3G8lF
s3+tX489iQK6RfTuoL60esTK6On1cvRpWrA9yqrN/4VcbLA8q8bze+80LnnEaMc29OvUV4kxeVkQ
DN6uuuZmRg5CvoXOKpycYk5B/kDfckkcmhLfIONRHywh0CMctsK3ascbERnH/Wlz4mgxWx+qNO+A
tSApORsAjCR4LGp4AmyGoNMotI3xgAEGcxTaO2vltRLbWdYc0+6BQbloC3VdSd2clljtiY1jppX5
PoIMot44rlsqNfvedTHbsQGevOBOricAFWB+82/BsMb0VnuOYHMZegpC72jsthTvZbx+RBGAXkNI
EWFSOsbUORfrlEkU2JT8qMuyBWHblZ1KqA8hqY7QOT0nWHCv/WYjVT2eRRZhHgleus2TH1od9n60
DdzqsvHJ9sqwLPQbT+4zg4lG7jRgJyUKQ72EcVmaJ3Aurloi+IUBM0+edZnUOOvVm4qW4MuCgMuE
yYlBtsCOuK+kcTyT1es03unRw5o7XDhl4gcxJN3bhgn9MkMnKXtEgukU1vTsO3iKo6iEe07xORKt
djp7+Y5LgcB08R/B1QUYZo0W01uEeuVw559cL0clhk3e/35Tmu3sJMZC67BkTVWgzPJxRIFE4WNu
+Agi9Oz1ejm14aZS8QnQVrqzmeUQPm1NEMtHyKrGh4W0Hmm0JTyhUk1GveTjzHekAE2hb4qhEJTc
9almIcwmOXUVkmCBAwj0+02DsiQhyfcJYaGsYRFlOfD8mMjQU+MSNI85o8/L/d2GKDRUe+F5BuJn
IG/X9zbgvboPUYgtV8AvtAgR097ovCiyotnuvls91OPL6OLn7deGR9Kb0JChyqYVSSd/G+5DcB7s
W5DpRZTMpyuR9cGDWVoyXxt6iiOMepSgqKx4grHthShBrQjyt269pmbpV7pUpn39gsZRk11h4N+B
yKljV9E5pm8R3LRTbP9yuQ6wPY3QPDcMZMDPfvz5xp5FQnOuD3R8kczt7agRpc6M6v39s79vlQjn
TZKNhYAu91g6dEF76NKMbovE5W1L94k0YpDzkxKslNZM2BA7ZrZiVP9Wm/0JJcYoWRvQfJ9ZzZX6
/qdteI9rHyqGvzub5emdOeRayhU1hoy4MRRwCeYMkAKsjfnR2QyhzEphfYgf1gMmQ2P8IQC5unNo
Zp0drTGCRYFrx0Myun8X9ne4BeuTk+s4Z29AlOUF4TzHZgUm2DZVVVtkYjkQI1262Gl9idSO+MY9
Z/Dm51gG9bPbO8ArK3w06CP8scNKMXR2mHU/KloVJn0t1nUqdyEqSZR2kAbq14I2lVM1a/OneIHh
JYPtrvgzIiHgCQQvkfjao2PUeAVGQJQTPRcTTEHKyXX4puEdplJgUm3mFtajHMjVTGw3LSSfvwF9
6hayPG5re86O0uJpRDURxnj65kS9jTZxBjvS4b6nLw4meYOlYzcIEi2qP0VcB3bY9i9SHe4CGjAz
4LLWCPivp19hNuhxY1iplZbt0sUPYtvXZzFt3ouG+SrRIhO+sYSOcz7y8j+NLE6z1zrMbomGcMfw
DXZIJ8jRojCih+HZsvVtmGFEHRBhHVngeBR0Nw1u5e9guNAZr7TvAmbTvgTlNfr29YSe5AwVNDHS
v3UPF/CVoRGCzld+ovxI1dlPD0DuggXvBi6eQbeMWHcP2NAnEIwuLNJpx53QCGE5gWUSsIyzSM9J
rIaJp2jWrkap4G6C0o2lO7tVuqtyywCSKEDahQFL7paG3LWpzZaOZ9/0mEnSbjy/Pg06XA3EJqyD
aPcwP9k+xHqJsAlvh2KTQizSR5OEKieTR0ntXfRlen666Xf5N0ooJj8K/Fmmk4eNyNrTRjX5TDlU
kR+r5/RkmHXYO8prd7fApKdzaNZgcdyxvhBW6PW3bTRWV+nV3Xo992S8ixyzKTVBrpNnWup6NWUf
EqGmUWQXEPr1Zox3kTpeRDSBRqRdR96lce+erTYZs+tUgMN+Z6ZvLMdQRTe0nBpqrRoravqb3FL5
TjmKjRQFdcJJNFQiSh+vbmzXYL1DQSLXZUKj68seOY8UQDgDuwH1UzrQJEXm41AOQKk5vGSpwCBk
AOuhbovurw30LfdlrsP/Owm/xstGMUmXUH/zDMt0PHPeBKazsVmturdzpFke57ExApNglSFWftKY
Bpt2s0cpuo4gMtO2TO1uR5ffFrnIRyf6Ese9V1aJjIp2ZIPbSvKOaJpmx+r5g8QtNk00E9LHBW1w
TnZOKLeGwM7uF8C/lNnKYUWfn3eofdMHJzHhVE5hzcPAXooLYAe2wt+5IOUCpvvppgilJzTuzrDI
7K7Z95CvnJ8sfbkkyLiRy2qrP9xhyoKipv1M9K80Mjxb6qyifhzfM1DXKBG4tTlzAE8+vKWt5HPS
VN+06iKYNS7EIVNk2L5RTDNOFjgTy+MC0mFlL2QKWENqgCopNLiHVb0PFVFLSZ6EskvJSsFLnBmP
WnyOwxIZgMQumr/hBLb+RpeR4YbGoHOeG9PoDzZG8JpCeVmrF/gXqSw+drUbeT9JP26N4vKF4KCZ
Gfhrzmr8UUpqJPQVX3Y5IprYvVSCjOucHxOaBloBygnYgA7O4Qx+tI1a6Sp4H8QDrqrfdj6aqI6O
F1MpqRfUFbXlUmDdT3ZatkAjJBrwL0Yw+Gisk3GVSpQZ3e66WcWEdbygVqejzRRECefQ3vJE/SX8
SFqQFduihI2mkBJrDryyJUoJRV1SbAhhT8CNAY5Gzc5C29JKjv5usKKsfEbSqEIyoVimvMX9az7j
8S/xvPLVaGB3nuKlVtCJJUdidHlZwNd4XNBU/PVJ9w9PyQ5stkBaS35JoaVVfNsD5yO9ys9GxKMW
DLVdkm9wZ3kNYK1QkdZUHXWYzIDWxEFfQpdtgBkzLthwfvvkl7Il3hzt55tZzAKq0vynC9PDdsRD
GrFr3l2EyRwDs/jxEd8IQDuolwYtMY/b+OrJ+IKUU3AGqwNBGZ58jdTF1m9twakYgxP3EJpXkEIw
tRUbDTGWjeiUwcDHTEVDY582RtBW5mGgF8Ydb48oxewHZtWYl/5WFMR5XlNjj7u5uL0c4PdpfRzX
L4CSN6ydQ+0eJiYZFN8bl2bmR9pHoGVIfS8E7Rgi3AdMfPUobc2nzdWWbLrWxI3pdzpzi68Opcdk
+P/LUv1FRRF0Kur7py4Q2ZzWJiV9VPD3QKVZq/GCxszbZXpZixO1kBq7XLz9MkyXHxcHaiTMPMtY
ICIlJtjOFzejvOw/TZplIEoVXw+u5bn0Mc7koHNm1KHlR8sklBiI5S4pImup/Ujy1FJSkRrAeNr0
cAZzjA8S+eXnShFgp25tQ+x8Bp4UctKKzQFpXdLhdyzIf4l/47djMPvoR5CZfzToq3zQQ7r7i/0B
S1kX5b5uTuWr/9v4pdVtpmqBXN5PHpYMrummMc/FDshACV+u2K6mAvoMCsaFAVDuqc4k8cm1a5UO
j1Ml5ZhyQm+Dp6BTuW/VpwB+v+4H+ZaTsXMlHjh9ffWsJjkuAVfugqZmHdPiLCp6w2tNQLn1uGnJ
zDl9FZNM+umKe6dp7Owm4gCUwOPDCrHj9GcKuJAbscDbwKzxZDM3KN+3CKv7E19jxeFpPC7P/Gin
tHaH6q12s8YwmWqgx2Poze0pxjCLor+kXiSraQtK9sURfA4YfP58AyBpeUaW7yCiUR3s5a7CzQlJ
ExXGrjInnNEwELNSehZ8+0SfEAJJGa8lhQBJ6hWHn8Zw2Y/k+c43GRc3d4urmSiZ36NVl+yUuwOg
LDLF4IqUlpudealDI8jwWHfAi/yBkX5wY6Uloe4nPO/of20C7UnkVCofLP7v409rJYMAS89g/XYb
PsY542z2igcrd6nnKBbdmn09DNuEZN0PeSfrxu2t95YUg0Dawjdtm5GIWL2XldMDvqYmT3m0ZPVr
EDR96JkGv0MyUq7XcfGLmqPwfWES1CIHN4bpzJZXaOCYSeQ7iQbhohl8mxBM931m96ZhvK2HoFph
Ll8CgSIYRzpQ71+iBRWoh6f/8LLY+YrnTPFenqEqbEGn+eRDA1jeGaX/B+u+6XybCsHJbUHG5jrY
/diCo88WEr1kmJBFapNqVlc/9uDZAQwrMMCFeFK27MbC2tFCMZkzA/ZzNQmJ60MFOFXpzCnOZpvW
kLwDUAI6CvSBKYb/m+W9mYuyJlh3qas6MLvPpFd48ofxSKyvNSmYqLf+CbkMAq3dgUObIUsMeSll
DrL7zXdXzik3wlMZfuWUpwITj63iyd3u7OBpiFU7JIuU190gRlPZnDeigpy6KHCXS1Uy9s6hPjd1
/wV1vylhaCoGame7c70Tyh4qm1XFfGBt+6zeR5i+UwZJsjOy1JdSNKVH8ZO42ZOE0Kozv5w3VJgR
z1eCQU4LMxJB1DtBE6DAI9OUOTC+nPMwYGLp6Truk6OHfK43xpCOVh6hHN3hhFiBlnFTFnf7QrOz
0WVlATIBWqnsQb2/R0enXOiRzByIbKD85OZwRGFtbUcmPpIFnPW+d8Jt5S0Yi+do4Cb/MhV2PK0J
Zx63GHkeJda7LYoeJo02oGulgfExmSTHv7SQ3oVpJ2PdTBLb5BX3HGSEN4w4NkT2AD6GRfabRN71
8aflkooy+MHnpgUITJ8WQKfGHAhhf0HY1bqgw9Vin3RGIsFwq7V7Xsrj9b6pem2QQcfiFrUFWFTK
gkQJMTdV4MZBy5+omLOBUHUOdNFChMCsRsi70Fy9Dwh4Zl2DEqHLDkeQDdcuBb58j91sAGbFFHNC
q3Y3HOHB6w4LO+tGTP8RhtL+5jv5uM29d3+fS9IMSnFd7/rYvqYf8XSgwyt1XDgSLT1g/eStnCt5
qltP3IHDvA+7Ysf7cLtnFr0MeuegtwtrxM1wL7H9Th6+mueavK30MJThu0MmFPW+NJPgYRaPLlJ8
CsAS+JrJdG+L5xlXxxteYB2PS9hlU4U19QVJ51jqKXCEkA/e4mnq5h0tqx1X0Haj4nkFV+Vf+rAD
yiDNqkaiW8zxFCplads2SquY5HE/9NymWpW2GKOabNh9/EVzdAdl8u2Q0gLE3nmxRJVYRRji02or
gEgW+1dvzHUicHfgSdO4vDQs7xPO5qSYZdY0MIk8nfFa5LWqaYESzfnFstiAMBvx1z8RjX0DBjrT
2ZiaYzIFg1nVAyKAvMV1HJitiDfs6x5VKw8gZ6CO/NU5NAvzbywa3rvZNwtKCYgiQnS0Vxo26DcH
PL9myX0VcTzebPxmMIueQNGQxohzaVbAsSO2pNhxmq/ckn51jmc9oNqBEHKdYWghPuZKpmdYd02q
Md0vRvKTz966KNzTBiVydkFI88fVW7UVLQuMy9H7p4zv3R4lXizwkg1Y2A9bjMPHbipMDsusfHBP
taVcoVXPmpemvSs5kygBFBaZz7H+6z+d+9NI9vHWrABzyjepj1W2R7/8y/B3yAoMhd3378ws0CSE
GHopw7BDbbFyHscZd/Nmo8ji4TW3yi71IMFe4yPuyc4Z5Z7Alek+tBDcl/EKPZ0Tc7J+xoc+tMXo
uVzCO2R9iUvG66rDdFEzFRDO3j1dZOpBwWhn6qslHZReRd6XQdULH0E3WxopRDA84d81FQn05ZKM
wSrfcPh0kRc2532HMVP4iYUmzoYbMfdqLS+0+0PPrnczFfA7iFmqM/4LbaEVMqJrauBnG9rV+Cui
atL2B33NTsqj0m0IR/l9OjHxmDTamsOUwwHjZchZcg+Igq6vG6D6DjY/abDRYdESwwdV177VcQrm
cn+hfCi9sVWzxBuL7kNStXGiaJufKsA+mlwI54b2k1MYgD/zXRKrhQrqpxAgDoz0SXC0gVGhNeyy
hWdELzaraUfm4fTVvtv8o0fM2XloclDPDgL7q68SKnmyOpVQqa3m44NxPXAlOokkDDqJhmZFYoHD
UWVCTgOV4jHdoef8I5FApiubn7ISMxRr7oxty6AOfMzi3TMtoJdnChVnG11Sjn07zFkRWxD+tIAN
rI1fTzwgFPwFfnOwFwbNG4+eAFPVp+T0b8h33bgJecNBbZAqiT+q9/Y6hpVAlFLqEJVFBH16fqs+
bNOoVASVCl8tMnks8mNKJHQCScTniU20K0mg0i4p/4gbQPpJVhli2u4E9sYiBMWXczunUAu3DeDh
f4NIWrkBC1GCWY7QuxnjsgTm2GQyFbdwjd8h/Wpad1taPR9hH0pA7fRArBcfpjLLN4HazFaLzu/v
DuNw0TCPjmiR7DPXGvIrJ7k8dgk7Ov7Ees2fWgqjMApNeNbUiQsbz0KM0+UavZ9BHY0ISM4lCkox
x7mPq1Yh2X9SbvsgiW1dYEm2oSyJgOXxPSrl1EAIbUIhb9yknDm3XUAQMpu8FqtjAgkrrVVHHpPL
OALcQmKq5kdtO6xK7jF4dHIyLo4asLBatdK8FWElQrh8uFpudOBBYuriU6XWfsUvqclxBoZLR6tW
ub0TXKCpjlvJpwe0CecGeA6wLLXFP/KB9pNCDT+T1UF6eRIEdRJVVCwM0h3sNf6h0bFGe29HXtt/
Cj6/ZaGoerJF4UYEH/MEFE2lIZYRIOmTSFBKcBg/l/cLC76QsX+tGEoNtA5h0y9QVl36JbxMOxDj
ms181bOivOn+jhnd93PQK5q5U9OAjhNgFdBdZdDzWtGbfkn/wVwdOvMLqcdvKGwEz5EvhWo2cW+k
5l1IcZL6Ny0b+vvrhIWrul/FmyooHsYQWdpkue1lbSabKjINkG6GyP6MCRR9WUZ75Pj8VoVdKQ0k
zLIjIccK0bkQqxvPHw2lb6GbxewcpmsALg7pPbshEVa7/u94udHyoMmjqRJMwMX6koGQ2Oag/nyi
fZjUNHfWQGu0riszxzNDbfJ/uiylVwsWQb4SJYg6fUO6J/L5HdCqRnx/rAMkffcU1EYIqlPNn3C0
Tefq5Gdd7u6YvLIOBuN05Yy1UQARn5pZ04QU7RjfBPg6YOuVPVhgnYQMSY7fzjDi3GFyTfT2RMV0
eubaZaXRNY0huOyz/jrfD8WLFiR8eYBCRixV+YHgP4Z1yfd6tqJeBxHMUEHAtLyxs3egNu8ADiSX
qXdD4TzkGlt4R2LcemoaPvht/LouHi9NxQbtjXSiazYqTNn7P22fwjeRglskklQ4i85EplYXUV8T
2qasLZdSET6QLXoI+PwU7lV+dNObcJJILx1WHmJBx3kg8zFxPDAfY8VN5HNCCcmASBxATkJmL0Kg
DKGB0A7u4E2fIsZv5KO71U/36G5kd77/oU9fEftwXkLvjHAQ/XtL91L7z7vwq016A52CMdh6lrAU
M+KAi1pCwud66bcl3yv0uMrHbRFmrX6x/hP6imfUMittvFam1adAIx/Ql5neEMhu2kUCK8Et3SuZ
weDnPm333ETu+VIT+WDTb9qWAiQjBYyLkpqWCw0MDsXgbwwM4wWG8XOd/m4c2Dqp/KxL/Kd3Qcg3
Lr+IdlzMq+9FXQBEZUa/u/q3BhMm2FvolMGfA9Js6jmDwxdb7RbfAaGWcQVcAfIJvBbJvY5+D9hu
MwOu7hY+qxkox0TbdMVHsIz8heA3fiWW3MfOE85KsvXPyq/O2HNRn62g5lUbO59pyWkhKSnzzp5k
dvd5R0HJZ18pqL9TrLeuIU468B8Ma7RvFt5Se8ql9DfUqFTynSt+ipxH54H9mWXFbGqtWcvka81m
Q6/YLmOnQrj4KGtYSbudcUfQPNgwoWljvimB8iEV1mcZSxAYdlTITUH2BWWdk4v9JI5YF1VJaTWH
W7O35Q0IU+LXSUhsdwEn+SjiN35mcyGI7ZdNBdG3GgOIxs3HxPXQ2L7kshNkXCmRENQKKc8cTK7o
sWv8MpXg7ftLku1JwIaslxhXKHxhqiyTQi/WbnAmID2KlQblKJcEZV2exYOOTZt1egzMPbEXO9QG
R/yzsR7qkz+B3okjPEBn8yAqzIlXNBw8MmgR3TwjjnSmh5N6UVlQd1HIaCP3RIGjxlMcKbpxsQBL
yq3yY9uUAoUmmhjj6SF1I/xNFqAI4fy/8PJv9If/odA3PAQFhMbVKeTT5/ugCshKOR6p3BVyHY1Z
rB0wik5L9v00dgum3jMRumlygWAIaCUwN7O0+go0OFr266seW/+f9N0y7mg7ATUYJqsPXn8XRFHJ
JxLKUgLCxkW/KLDBijbDrlcwHGw8ZKQdaQab29pC9SbTfvU5D0fWSJ2+IEyWfHMt//26OrM9UTYt
OMh1LXhX2N7HLtwsbeGp5paUb8gWlHwXfU708MEwHGQOiySN7fxqPHEb8iOmAuOdaMS2nGKmtiua
cVQqSzv48V6rmijgkboL0YwvRbZ4HLtS5aET+Dkap07ykOBTJ8fkcOBUeA8QvEQ7J7mQx2L+8RqC
iJExUY1fR05ymxarNKyjEkik2hQo2vth53Hk3sv74NCOEr4dRdTqE6GBmlD3eiqGpOW4jaEZ4X+C
eSfDFJhVk8Luew+qQD29SAzfRKvtj9FTJQsALLBV5hhN4OPlYO8DWHuf3Sa/havJREkrUzRm6XJe
64bYwo4Y1RDAtpS3BbOI5DVA24YZm58spdGL0v4mSoozStQ6Onozir2B37x7AmhmThUFlxeXtevH
Ih5CogYwb8TTjI0d6bqMYHBVEYa4bHFdH2l6d2EGfP0AwyR6JIMWWvDKzTy8A7JV76h3KREJX/CL
4eLKLzIRPYVwukS01XhmbxyPVGVDphGXo3/07BO9vuUV1d4t7taCScFgULmJpohNObr4dsF2izss
5SBUNTVW7qarcxZUyC+qKq0yJT3ECo+aRhKVI1jDxyERvRBa10FBCdWwCiB17lfx9Jq3tSDGARPi
PwErIrqEJIG950Fie/c5+XpO0K0k6JBlE4I+cELQjfoPXtmwdNxTsINOSennDh3QZ6phffm6WFG6
XMaWipliHHG9Jer6MtipP5sFnhFfXyuaZW3dTaSTYnAfClMquomeix6bH8BoLBxiufpfduj0zL6R
c4CtgGm6PYCcqcqruSkdKh730/LNWuGBrz3aKfPj9/IisCRYI8800LUWpQ7qKn2yazs/P3YKbTYH
dgu2NN17AZ7D3tZYWEStnzRnJn4Z5Jhnt+GM+Y6d/5e59+fjGF8C0NsERKRwMsXzuRD2frQRPqPv
fDft6ofzpSe6PQPtEyF+vEoL6fPQH/BfRcHOKMDsda59HohJSN5u55jY+GqOWlx+szw2hOLKwSxS
TV8WSQquHVfapWQf+dqiImrpfSQ9fPIK6Oc+7Xl1I2EFRCw0mDwgph+Fb410RO70Kv2fYnodPcLw
mXzGU+I6zyRXIx08GhffJya9E0cGM0e09mjSF0P4IvpN8/WeeWV+wYLKqZkNztfgguW8talzRwLJ
hVT5DjAR8i8O09X3k8RTETfZoxa/vN1gbp1sjHEQTkocTpdjHuEVFczNwr8f4nN8hA/zgIPhMo41
dw3guSG5H05QBxE+/bBYlPyhL3qmNa1uaSlmJ6/OTgPME7eGPcxQl+JLtpRl+SibAf+Do94mVMpN
B0uNgY//mdLDNc+38v3x6zQ/qFfL6Qv7U+UbiB0n9A4iRmmyRoEutQAXFNF4z/91xwkeHi4XvYV7
rKFWIQ+YXU4L73s76fSBMKILddAtDOc3uNaUIf5pyatBdNV99+xWQrMYmHgM31afV1rDu1tCwRjq
IiJJ7jE3pG9nvNIGZBl4NbUhUO33CTGoDTkBZEAGZPhijGMMgYljP0+ccCM1SCCoLDtQGDkaEL0K
tv8TKQhyMFVuCwvDNUxECOgviKM3ABxO3z7bIah992Oc1Gi8aNi1UZKPxswpbQ+XpLEINWHjqIy7
/+1MWj631FViACPASYClcfLaG8rOJPUYfzQzkOfECU1leiZxSRwX3nA+vaZ+PRngKiP9ZEayfLzl
omsiJ0bYtFEenTXCvgd9jpzBdKlRzJdi4IvB/tBafR0LiX7dhcKH+6bo/GU3t+b+AK11RpZocYE/
WW1mDCvHQad+ZpDORgu+y324xWY19FoOiQfT98GLHGS2n7s1bXM/kwjgIYz+i9nfogTaR/nLDy9l
DofCxtm+y4bje6VDECuq8cs35eVKi0s4ZtHL5T/0XofO0vsalMEYOCM48zyfNA9WNarDQb02xA3t
1ESbrDbIgGvMavg1/nZuG8hmL6UsqDyLtjC8glYzdC+5zbKDnEMwjA22/FY+6tRV/rKT7unzjwns
D+qlz90lVvhSD1zku652QhKvwx8RvLm7NmI33RDTBciGKG8zLuFcH0yuE/08Lt5NcFbBHdAna/re
klkZyJck8hFISl2f1sIxoR08qAITWA21FcWbi/S0OMr26L2fR3TKOSkLPhjLtxWhpn8F3sBOdNvK
F3+hbSwMRRMGBg0/M69OLzRhBEqi2BGsiuFGJCfv3IGbuCQDjgYlAOLPzPwI7CKyQAHA8t48DIzJ
DHI0O8gw0Pb2b95+9dWEL3dzic8H0FyQKqGicut+exkdtvVNyKBMy5pmj2Huiw7ScQW/PUBi5WTm
S3c3fOAyhEqrluhZbbeOouWqNqw1SObOeKtjNxNYKKMDpgYfBZWdtsSMZCkhHRQBS43hQREkwuOV
J9RCBcLN4S9LVszQy6Hf0EWq9CtKW8i21j/tK67BF+VihIXgQ6VK/XZVOqkfVpjLjsbe+p4Bp5Q6
vkjkHHHai7Oe07aYoUgVUPFn5curQxfe6PHFsATEzuncb4fDMQgQIecZY1ZWH1NOboH3I7H6YUwh
UE23Hdru2NivyAw33dKwubp84S5K8h9+E2fNn5qbFLmYT92JlRWVHf8q2v86KVqSNGjmnA5lCle4
ziCbcBFbQYXS72pa0WgMJwD2chGC2UwVQOhwFf2ogN3JqVPL+ld6ZMWzS1xetu0BKtiPD1KGnS8B
07zMW7/QzXIe/G+bwf3s+ZG8WX1jaAIJsdtH3zYMN88hXQJEJW3exNTQOelAw6hElLt/JO5mAqlY
6C3+B+Dg3iIBsCURBExsuLT80cK6UPDIIVk6ovovkYaANc0KTl1NAq3oVDuA+pxjuAylLdksOwHl
S/IphD+U3QYn9iYGUWbxkgtFbkdTaWbt2wJXF+6kxaq4nZzGfPi0PJ5GKR16JAjW5w2Yfs205HzR
ClpNNu64AwSotrUQmfL8ER87cStT7I4sK1jR6ntGLnDrWPnD5P6XlHKzPRxErvE0KpnOhOe9oRQG
100YuKn/qdx9uG1N2BpHQqI5i0PA+jU5/LHy7PKKyzWbYko1ETcW8asTVJ+kxLR98SuGp2U5V6Zj
v9g2lUVAGKej2MrYzPgurwDN3m0PcZCvKBn2OFtP5+hoWUGUyKTTVlO59lBcgGCIVNnp1A7oQwGF
uKU6AgMCE5kr/VaqoKj8mM6hGpV//RISiD9GP1PGnmZD766cY2dzp9u5VRwx15LztSDYAHcJUwll
+h4RBDSdqCNCbnbINrTfWiwgPHGrk7NsR+6DQ9pForMiJzG4LWYfjS3K2Ngd86NQkXvwMPEquiuU
QQKCd4pDuNQVPKPEky4tVih8iSt8mLnUmmlmrb4kQJVeWIkV/2Y06NZkaBx7wh1Zb5iIpp68PcCS
kpNTRLvV66YCEfnaWyQQYH7UArwcO+m2h/Hyz4HZexMJymwEXtVYMThNvKjhcvKbVQ0q+GCx0bUA
plltpRJH9xUbi3Zkq8Mk5SKHEdW0GOwNZEXPfbNGySTMp3blX88KCSuC2MnmtJAgNLuZ83iwS6Bs
UZZH41gW15q0pJxCSHX6CCXu5UDLl+kmub6nGH/mtmc2IRU61nOj+7V3NG14osiKJpZGFR2zLFar
J1pK7wiMoE1R7ATbxXgM6ypNrE57emMhleC2dmiCZ4kBWLN/Zonz6gZFMiU+Y4eGZzcr6m4RlNvB
WHeZVMN7q7Il/Z+NHnZaihu99A01J4Pibp1W/htC/D7MViqBEDFjMIZ91L2y38G0ihLjYomuwr9f
PveLA5p5FORnPzQe0dcEx2pvFih3xbBYjT+vBvhpuP5VcTskjFtViiLlL0fZLHZbnh0mH879rr/8
F2MqVf30z0QW4FRqoMlgimVuaAyMTCQ4QZLwST5icEs9bbPKRWlTCVeEeUkr+qGh8j7WlpeT/8he
nIVKCbTHRRMnd5VhSadRHIqxWnIWTsi3DfyIby/xgzffkLvTvnbsUTkdJu54GTHpw/HY9T0RbPTL
eqjeiT+uyIzKWE7JQ+YAVNesP02CPrB936hplGB5Fn5zzop7rxjP3fK4vxQ2V8vIJ4e6jZdN0DiM
JJFoAP6ppII+tp8euxqPW21h0FPwXyswPRG8LMFQLtv9pG9cfhzeFQbkNpbAdTPy5DFp+zRY+/1X
Ob1+BBmE4wD1qCVnlVjrgOQOjDr6U2cqDcDF0Kbqh20aCAlzPQuUVbuSGnXjyarXhBLSbFPjP+tB
ieOjqzM1UsO5DlPwJDIUP9SIyR3ktIiKq+qDiUX7lNwHurWalDjDG281GtqYjPZei1jejVfdb1zF
IfGxeNu7y/xar0mMKwfh7mQJYhOy4/4bYrbrjRqSZtS4hNpor0+ko3hOSirYcwZeT6JtT2HI+s0D
Nxv4QzYFW45Yn2k7zvHIdmFnOqbpQENZ6xMmnkb0Brr1Ukw63P3Ifddww4JuGhTIJDJOwV/3myAZ
shqDAlRztnfjPz3M9PD8o82RzHt/eBThS6eM//0FjShgwOuQAgrP+rjsiIQrBVrl+jlWeFv17Sfq
hDQrv0+jQW7IRO1WlooozchHW6O2AexLS4PpYiV+fMSWTYWzqRvDRhxZ4aoPpErEVinhxyezmITQ
CRAr8+fbEOWHHcaH9exH25qy0WUnXHLqJUXq0dUTlvJbUnGIy+5T19oVk88CLTCga/UZ35vpltCf
hJ1AM3ztblMPZGvZU74/oigAumqB4/CfXmSlu06i838q+SZ09t/qx6+6N1PnTSCXqPZdtTBBkNNY
PsaalQ1PoY1ERusQ/dKze3qgKXgiCP3qSDTpBn8rHUUiQX1+6RNLSUAUr53UVZ7suTKL0OMBq9Tx
j+/U/1mrNHhbSZDLcBHvVzs0XZNvC+NzeupvCYMMWBHrY5zwUmYpyHURzjDIUl5BhnBG2ULcdRqU
Yzu+yOBLli7BZF5G2c/AVyaOzPE+1ysODQ9O/r8M8OFfM8QmYXs6XgPi81VQ/ZBaXHv5qm+QJd89
rAtKOV0PkKYUsNOChTIqWnd+pgtR9y3KyylznbCfOOFJ80Cr4qxEkjZzjaIiXX25/4J3huPwlBJM
TfeHldcDL8zoLTuGX9o37TXDSQRncRuyCtc+kejAGaU1OdUXM72hl7FyaDt8jOmAZZPfbN054AHi
VpuI8o/mZlcnP0nkKtonXJxjEhQ85LvNTxMnUIJ1SckFqARj1eWQWz3gSaghVkpimfkahvxYgqNq
MO3Bp7RC6wiI7rljzb8IK8t53+Spr7CxzK0Vbkk3xe02GcPTegKeSPdHmuY3dTcFnG/Ab54c+2bl
X2E85lmcftTwbEUoIhzDyhz25PMv6wECQ3LXkiD/cgYAUWwu1lf9w+ILhAZOOJtonGm0r65RMI1l
Mtdwm703dT8O+lyTvDmg+xkGjBESYvOFh0xIoDJ4O/EIIcrFQAL6ygzGnjdt7ZsUMkjCafsfR2FB
s5DnmLqtLceRB/ARqN82GFfUilCBPjJUYlI+te7BqlnxOFVa6GcMO9IU/wjrqksyjZUGsakyN5PD
1hQ2Jtwj0BH2G82GYk8snxjy01RIVnql1wzl5VfsxXlE5ZscQBrxSxpy5MwaBl1QBsEtJvOT4ZvW
q2m/7BHlGjXMzXY0jlqtumI2Fh8zI97MmB1qqCmST6TCcBld05dlBcOyWbH0teYZI32UMZvPUndM
+qZDPsaheK7rlEtNg1L3FhEfuqvFMqo449eY04v5adDlwIyqbMLSGS+clU3yMoKV9wcF2g1CUIxT
kaJrd8AY9U0lldGqkzcoD5eo9yyhLtjHSZrNsWSdx94dPjfchmzBdtwXUWG6QoMnlPgTbC+Gep8N
kliCfCSaYwd6TCiQGbOCDAxOldL26LnOia+E+q5bSHPkPaTjZ4JyMHwRgQZmU4+u/zryKD9qkiyQ
tyhNRKFcl3MIStwmYcW+Kh3oa2qRAoKkL7qFIrtmmgXjLLMXFrK1+wIup5J5uUcF5PfgXMnzxaSC
rEPFZr2uddQsLkMJ7z9tkEh8NTCgqh6az97/H1YIotNuKR61TY8xOt56gaBW5iiGv0fMmB4E65in
3o+iGiWklSMR14l0Kb7AmYBGeOJ1W6RBkJDfzdwVI1PWeIv6P3oLyHmyJwWbzqXTOXy2/sPMLmsC
gWjr8+IwHIWejOaIm7puxGYLZ6qQXMBdl/bWTJLUIp7StCyEZuYrBdzG6KTcBdXYOX8Ja6MvSoaN
Gqez6KqxjOdeeRgkecPfDAgCMjUejLnz72ZPQDQA8YXoS1VCR2VdZn7YwbO2jOrpfaBB3mhkGKMM
QcTT4VD++HfeUg8RPRCLPr5R57ObUM0KZDtzGtkWPH8D6sMXk3E7tuODJc+r2BpA/QEmxm5RemcG
NbrfQQtmipRmNB1997fk1iy7M2K8VVRzLiGeDhMdVbft80whAXF2YKK735ZRI4W9wKjUC22/JvA1
p6stvWpLCPkcRQABFZ7cV2NGr7g/gIgQCPhv8YXgIkxeW3vLfoxqetY/JfOnlYcKuxKt3MJbJAsx
/saHISS06e1Q5XpVkpHkFenwF3MN5mlhfTiFkMDOuUaF80TGF2okTMLk6dTQ7pmlchnMG7+0DkXV
D2LXYzkazbtpGgD3QnUxC1T3JhpDa+eNRen85XXF8eywa1eGp4MToTFoU68EogmMEJsejUIuWln+
TD9gHw9dN7LW/9Xr6olHZeIXbz+aQMg12EtKX5ZtvpjRybUyF4IAbT9crDxlLd9iVy7eQWazmz2o
JoXSUrYdlHJ2fl+due11XrxXnGlAYk6T/1qLUaUUNaA1z1+E0YOAj+0kUKrQ0/EeEPzWATzAidFw
1JZfLgM9OsVtjjeRaYscBoH86oMFMwnJDdxFZQx+Di6GirkIDS8gkEwO6fix0vgTpWSI/Igfj/Xv
tHoA9S3Zu9hyDhaGXWMWkaEMeWMPBxr3QIZU9WKi4iaEo9R7EcGENcmPufA6F+UkR+Fj0OgJFHSg
Pp+AhYNaanqk6KGx69yejxISC31+L8Fy4zUhQMcs1EfcFfxEJj6kp8Ywk9gnP6J1XaQqmm1uIVZn
Jw1pBw+fg3ncfCwciJiwm9iuj4YwT2t761zJ6E44wfTpB3uVtkcn4gPXOoJjBXj5L/DD3QAHWwhc
rnFsbbyPbGkB0Mf9nF3cochboQmV1gigU1/JhB/QcSV1PGR6vJpFTQrwE/KEiYIxXIIRg02ehhOD
jeXxGYpbZp+wOyZrmh2LgaFPa5BZbEyVzoBJItwk3dLfPYa2F4Y8NpUr60zlApqA7Ixb4ijd81KD
6nN7OuvCEytrhe/Xqc/rNY1zFV94S9KWfSrqfFKV+0Ge8kiFAk64aiaTqEaDnkDLfVBBCgKEMkFl
djEI5d7jgYA0VgAHNScWQguWxmwG/7r7L1zKH5Vgr5mo9WIWM8EDA3ldXm9Q+89+BNzSkNnQQs4Z
k+FD/qbPj6yX3eQn8bCCs6lEfpQZZfl6gg6I/pesrEWmnzX4ru9nhrcZasNK6akOPbtnC+9iJici
DOgL8odui7OyDCvGBs1Ij5S2XdGAoT9CZSJBbmajcyqln9nbaOVa+sMP7ks0JZRQu76/WtOtPutJ
RFUGbVjnaxhdZwX8XS0tl4A4p9ZFwyWZLIQystmiwo9nokFUs8swr7WKdY4hX/P2B7Vf+XwiL72e
XgVBjMd9XRAyREbBE7FGX8DUyzsz+e6IpEiqzY33rXMOZsEFoAo+4urLjflKospat3Z+xnNQScXN
7afKkYHdeHcbQ2ggUtdmlapCWdHRjbpf+lfloByEVeUrghRerhU10Orr77eNhajz7hduX/4qAQHr
uwnKcdCnrCHLDXfw5WC4OexgplkwLwtJT7qt//YaPQ8GM26ZiB5FOLGD3TTppZysXWqvB0lQr4fC
NJlU/0KwC7+GLM4bQpPhjkT5quSRpFZyiqSVgg32PHYYvrdvfAqHyZ+Xa/9BdHhsxZbDa8zul/gJ
YfLMwAmaMDexPe08qiD8r6hwdCzHHFe2aQzE6ulcuKeOOshM7tICBV/fIzpHSZK3cPao1/wL/xRR
nURIPg74mfrHctoHzRaLkNj6i9QmswZtVWfIh4gMdRmmtH8eM2KpTJU4glyqIXwoFl6RII1olIPR
Mf3oChzJb3X+CO48tHXAWWaIvHsDy6ET9drKot/+WSNvSgN/gAwpgp3sDJKock7KtVOWhcuXPTYO
BQmIiXMh8KTe+RzRD6I/TM5i8iNhz2cdp+1K/wU2l4X0jkVizlappvlI/d8xXPGQDDtHv+JvK4eR
Vl0nOIhupqKtmnrGGPHUIkmGxfdT1C2pBvRAV8xOlXXu/HZKDM6cGg1pEaewLCaX+5joZuUZBUUV
X799xqcJohOrKttvEyQSlFE4SU0NlBp6+lIhkZstzjVGRvBqRjAuIt6u2mPSrBS4lPHwdVRTX6B1
KEdAlEB97w4BkIHQX6+CK8s4UyU+i4qrdWWny2BR86Uql7GlTl0VCsD+zgK7CV9dsh6AYvbuacmK
TDGaOm5YQsCx3RjZ10TuDYLygtfDNQX0pCKh6wdhHcPc/cKpmlt3Mq56wbOKDR/9AHu/v3WGqCMM
udnAWleA92bE8/U6eb5qKmRLrnTeRgO8HaDBkTIKCde1WW7OIr+Vu0jPAstS7KZSW/q6+ZJgXNWh
g2nezwuLdm359i8NjLZI+/p6jcU8uzD32FSgUKhYVwjD/C9tjZ4BWK5sRIoUzxpvNTSiunclRty8
JPurB7NcDSP7HOLVMoQlnov6ZJ1rOErEMYfLP9j9pE0dLmBKvm7IfdBgRfeS7P+sCuN1azH5be6p
UfOUhf5/NZbHMediwKwpO8VA2xqKWZtcmY3t0O/MrnI2KeL51OCv+i3P/fYiwDiq86fY2jN1bb43
yt44Q4ZF0hpVAUzoUFLoXFYNkwFmoibjJDzQZKh0Y8Yun4nl2ayWVTF8+vecJ6tgWcNaUY9Q1/eh
nQrxZyIQmsD06eKgFEZVd/GubkvPKf9T5fTk1wWHOlJyHho3LC/cX+39TBpKePk1UavI5WHDJ2B7
Y/vVNZr012Bjp+jv5IbluNhsUt2CjMcTpicPWzg57EVFfeV/q+mZLFXxd40RLd6lCPL8yTu16MIn
niNtCbAB6k6s0hVNY0ZDqPYOwFwZuMSJupLcON+rTUK0/wa8VBSF+RnCKHoZQZWxXzG68isqng9k
mmB1p7Oi+vVEJ8VUAIEnm/NrONl2X7hp4QXqQOf4cFGVFGyd4ox2dXYQvltW9lBkxXD0yC9ELwJ2
RsY02cuJUSax9wQf4e8EL3i38sxqb/KS+/ih/MOcbzF1d0OultfgQsWtBfMmS3/hOX/mlnPS+CCA
uhuoi749Gd4eSxKuc9htzhcB1e4U4YW7g1fyTMziQlpd1jkHYHXrIj+YTFNv+wLCju9d80g1VbEn
kwZCUYIdyvHBit2Vdx2RlYu1dBP5tIuIrQAor2DYuM64whP/fiVNL1xkjEibTobYlVAXq+giogRi
KR0x4+erpo94GlnAGW3rSNKEVIExAnfBM277cYI3ze8FhY3ZUzuSxlinE+LVzYQCxZKAeit+poGM
ox+nqAKKg+PQdrl/oxPDXrCcCZjiQ1+H/sOytOQjE2mw96Yz3fIQcTu/HysBvmkx0oPgf6L6tbXC
Vypu3jmoJEiU1Vpa5Alvo7j6HyhsqFnDS+M3mRy5ZX5X3BBUpj3gLhMj8WNAbLNZXQZPbFtZOvqN
8yspbclk+AhzGDLqUTpkft6xFLfxadKe+CySNGYWTtQqYmQCQlscKQQpiEYpl85kthOFZk1VLpHd
iHosRm0L2qmEo+DPzUfVqxsDonDNj3J3s3INeRF3hT/nk9tHFbk+dJu6Pb812xb7nkeve89Cg/Z7
CoqoMgZISzlmoX3VO4Hulufbu1ppSWDxZWZMEfUtjVkg+Z0O9i/0v8xKhv8hysKxiotjBSeJE/9v
Io/T7cXbIo1v0XQwiS/FI3UnhGQtbZjqP/QH5GMi9Lor+eSv1nK3lROXBJpV2veTtH9dyW+2zNDq
bzqMypakkJaaF51/WpeabPElIZ/dfJ2Ocz+Q1Z1sb42JdCPcKZzJovlFTAxk+Lewo27bmifPGwtd
s+J/K+T1OtE3c8Mle7xPlnZFCDQk1SQvvmlNHECk8OKDBv4WKPTrk1mt1gdy9Lg9pnRpjJ3z3kBj
pfJiG9EU/VoKxm7Lm5leSkZALiQugnFOyutBxk/1iVqqFdRQVLX4itVgtbvtP/fEKdBcDubq3reo
nXJU2p2TmssLCWNdz73Or5U1aAF+JAdeXBwZPw91CV7SEErII7EHoVaaLmsfebJY6dNS0dyD+LD+
fQgh6J2jvxRD/OCNfxClhCtfeDnJvdYqs16hrhsl5T2yc88Asghqz8ortirG5u9Q8jvVsN36qq+E
8kvjQxQRkvjVJ3957IROP6rCSVNBueWMKDEw0+5Zj1ryIocesk9+BwuV+oGVf/wDoORRCQyt5b4k
sh/62Jhr2LNVy2jxJ812dqgmQIfaVB4YIeMIDNN1bM7ltuT4L8TCJZ1s5HPNzB414Orz/9An/8QK
c/1rkGP4+u4Q8pIyu3B69Vz9HYA58EIvaAd4BXMjgOHIpIUQzYjxzLiFTbNuEokZk36sI9DhsALK
44mnQR0i/eJqoqUzbhaUAChMAac5FEQI1jqDR1Re/hYs15CgGO+wVPf1bIqMoNqen3hm4OF+pdd2
CVhADX5WKAehKy077G8ULkQTOHdeh36kiv59hPp231RSAn3djx/KDCPQexyGxPLr7Yuss1knrPoQ
+frfBgT6jAWDAa//mzMJ53rPD5e2kIpMVUZ/knuIlAbSRz/LddHC8npRK3dRbZ4Ri1mPeWbEmjrw
2RkpVW3E+luMHX7rk/bX1A+d5V/sc8D0auNBOWJfJwFYNSbl9nUlU7FeLH0jT/qAn3mRN5vc25YB
1tzWQ5IZGSJc27OyiEbZ+yT+Fb+qrmG5knvodJa7Kg3QzbwzB2y3GHppuh8ZLq8N+w4Q9A3kDJ+b
2xok/C/NWKeS04ICtSrgrowFUqNaJXTELITjRi94UU1VQbVSHbdr+38FsvMP3xFjAlFw+2JiSriM
6zOT0I9kODv96qcpYVkfISfPYm6EN/PV15ir6bdGU/4K/IugcksVRu0Qi6bWmYbq2R2zSVo9yn+H
LgdvwhyZDzayfjo9+ELdtxrEvQxevCUW8oMszug4J0N4WRWenpbwNwqjYUtv77+046KLRAxj8vnH
mxX6u/dXXBS3eOh8/hZjRs65OOm5suwDVtsUMrzLpRgls8hYX6dBbrICg+keOUQ9+Ni835cxGezo
ZxcTbDQRVy89jMwNBVBH55lyAVH3LW94EZ5ywrlpajmSAVGJQX2fBQmoD4cJIZC0bfPS4LeoDvrk
V18f3Ee0x+AadEzVAPSUp3l30Ws/VZxJGMaGmN1RCopz35/KO8k/sg3C8EHnsNSNWnIrusZy73xk
DtXuQwmsG0Cby40h80HCIJgvlcbs3pwv7Oky+W2As6vm2f7KKfWVi1nfrnUIGz96xKEUVaI53sPU
3LDVepOvl5vz+vXT1wZ3/7Tu7N1T8aguXN4hjtl+/BIvYacsnk3y/MALETdd+Fs0PlVuwkKF4VaG
O+eUsJKcVNq9sev6ZhRPq/i1tp5HYZrThZ+t+I/0Vu7M4ne0hDZIX3Ia9RW806FxnfD5ELqDIULk
RVtzjO1aTGp9nzZD2kZSSGcnmHuYeQ1e8JikvYqvJwSm1zLxFJVy8fohRhzrBAK2u3wyCidDo6dJ
agLdpd/LACgbaK1o8vWFE3JF1LqTGQRhfgzUOINLQDguX8CDEXVpqaw6SOf8B3jKRAqGIlViX6aq
bCozx6Y9bP8fS2g/OW2uzG3UJ078UmYGxJMxlid39QQF9LGKNGKpXo+vi3T8u2s18GI285jONBEf
aKpZRtO1zU/QSqpJrpWl+VjYIUxSCGq5iGlA425kzIWnPV4gjaH2NCGJclCg3xKDtVlSJPW47scB
LecazDam81rvtKi2962XF/75ZvxuNSCm1ry9ojnwns/f1208yTElRwaIj8yiJy4dFIvE7GYAKkVZ
ZGzMraHYZnyMUkostuiRauYlsRyj8nrWUwVslz6kZCZTVaKU5ukPEzl4GVezDlITeU6rjFHtt3ES
Rw3Nvb2F7eMopDKJCyx48wwryE0v+NwDevYzxCYJbh0vO9X4W90nLIehjHxfOr2JeHjXT/bTKJTy
i60hNPWPvW8dek90SbykxXlhsKLMUlNdY54E+md+EKXBweBGFfW3gciN7MosepXWRRPjrgr1mOHk
Cfp04BYthOp48/bx1MLmi/O+e3fqWP5EA5FyQ1uM3NaKXrD1Q5jQYhOpGQTujDXqXuS+nl37nQf6
pKBB6LHTgorw3FWCYCb8pYagtztEgAwqFpeuN4ee187X0UR9HLZ6qQVaQH1S+Gre0QtOHFiDVyxJ
ZllesAbmMmrHmLmEX3vVLy2odLlWngxfdGhqTnW+OTZACelOcYYb3tluAplIbC4oSLCvaswAO/rJ
/qiGemPmlMWrTpQAiHlUVbJI7OV8emdV2xz2V6tJdAvKny/yVU5UPai5maFt95QBa+5gfk/fs0JC
yo25XjxVtqRaCMB5zr84lWfhwahTlPPJnvl7YAmeUtPQqQMPOVoVILup53jKswYpVKyloLpWyGrm
Qyqp62urFodwVQ5GmgtNVpaHXhNFdrNnoel2/DT/MVbRMqWZl6KesYrI6JAUtavaVUiZJVORjFNg
klc+T4GyO3cqvTFQulTvbibUuSparr94W4Mmp8rcMajPIQNlT3sJKrwH9ihO7XYvtwUmZoeRrWmE
HfRfCstYkkDMW3FQUadl8IZCKlxha38yZMsHHFlkvA/8yMyTlwgnxPe8dVn8c3oME0RLEy+bB+mU
/AGUHdQHoG47cCvGKixR3XZnP3BnKRWrcTsxHWAZFagJVtngMJqt50I/jsmxTBtOt4ay8z8AqxqB
VzgZooHnZnbU/l1G4qi9kFshX993ZQIi4d+HfR33/7ejXVnnpqozOtXhfKsik7X4vio0nhSNejjo
C0ndyQOFtgZmpx9aTIn/TUsCvtiQEW5XtTTJ2B+tVlWBKyvt1HP72oL6/necOW9pHeyPoXYR8lS4
aFbEcZAfhZxOJnk8qcpC8BoNfFQxPwF8v2phVM+vgku4PToJLw/iLIriq1Rs+/nbRe/Y62SIH+Vs
necDtPcIgW/t52E82Ko9y3ZYbRmK67JhfzC3pW1Wj5qnmPrgI0qZQsMv0IocE6XXUtXqNOQehbia
OIb4YgWzulHycEVUfPtSyjdYzYPhicO2HV6HcI2xN7+KzhSVqD7Je7hm4faTEhrHavbk7IoISYbl
K4JGV2I/YFkR4woIb0fPdLuqxpii1sbkQGcyWUNiC1jT3wbidqxIa3Ynj8fPRVe56PPVZeBqQ0Y2
OXAVHSbW5n+SSMXRIxQa6NEahvkga984MBesiQTIX+mmysgZV+lrhoA8e5Vp2av0dQoIoI0ocFol
Y7jNKy3j0DA0F79QhIeyDxWQ5JVS07Qo63SxcPayZmomOn2zTYJHf3NLx+3PwvXijTTsGHbWjBax
suogRjxVlmf9rar6+K7MqxZQhOuwo3dooorLZ94lsZ1OmUS/Bj2rkeoaH8Fz4oj5jxfBDTuf7h0L
TZHkuwD2AHYHilN/GRFagoY1sB43DMpvVNTqBDR2Uj373AQKtCkcduyg0TFyj1NL9QI8D6hyBJ5C
G3FOWkA2qcELrlpmhtxim3ysBz+fQjKaNPWikRMyzYHOMxrUCP3nWfwad/CVubyO+oouhZ5y0fjA
25TzF7YF2vrSUfYa55o5doofxWgD4KO14ZjGNO7442ENDEEZKKkBuz4TUS4Q7Ojlho88Pq3qhG4c
pC+1qm/5/Gaa2PuGkxGpIYTmqiURT71/d89rWssoK5EDOpKt5UWH7c8Kf4csIlkoTwEMsifhfBtG
awZcbP8NhSWVF6wx1nUkxQjJ4dwYUOPPqoXJJehcbNTCh6BcixMnP/G98ofna9wMMdlmEEaJ8DDt
IkOeewJokrH6AYsPgDgJ4pmXDZlbTHcdgI/TAp22PBj2R/hSl60OkeGNAe1VzWhf6fghgKnYByXE
IMKv5eYDcW4vLjwK+xvqR8a4z6uAI9QJ2NsDIRRkUXYzWMQOWFcOwoTaYa12ySoJFiP+wqSS1Tsn
txXtwqicYPMcUgq/CjGUS1b1XuUfpHYJG7LJTVVTCi4fkCYKTWdu66zbqZCPcJhTsIEZ7docb+gE
SHfPK9ZdWXt8hEC7KvSPyhj12hmZ2L1tkF9VqzFmqRBtUFFRtcyfngiBeD1FEDf3bsYPJuFJmgbL
LCwBjnDa2qbI5Tm8tQCt1XVZzM6u3qmKp6avdrAN6P+dRD28gqVqOtg5wbokPzDuZ2xD11kHuI58
yRiYsKDwxozfewO0W+kTIHta6N59MZb09J3k37xTIee9J0ITr9k8Ur/QCJh7V/7xa1VAr5iywcqy
2/ZZHyfVAmbj6u054Tf9zh+l9jGSFlOTbgdO62cFDa9pHrkJYG5fDSz/wtu/MxPom0DKl6Pr/X4g
HbedGy1eb990yXTBz/c0H4MtluH8f7s0pHmcd7R5KrtF/nEONPbtskmsN7fakIsacz4hWCZS7V1Y
Lc/71SCF4tEnQIvqrTclyiwygrfWyVJZb2OshQ5OKtEwzFRQx1qvQCt0UNV8MZaFnNkn+8nN1tUt
+Z00op/Woe02/QBY7lskrIvjGa0bayOZh/WKSsUSdsEZvI792O/6EbA5WqqHzz5OW+0uPEghofzE
Hb6L7NALE2q1i/y9acY8W6+HgGCkEhkIbXvZb1iv47wCvttXIEtmVDWehfEogrjgNySMgbaRXjbM
dwmN8A37QowMfbwE6Bz5qlCOxuuYAHh/Sa5ZbTRs90+Yo8+hZmStEzIXamNzLFA0f/7A3i7Xu1Si
CUtfzNM3Oed/F9FOISxXGaNNReyUE/Nxq8mLmAzL08JhDtwd2TkD90cL73qE5RVaf0xybJPJ0Vhc
rUt/f4682M/RvQ4iK8KD0jbMtnfnsgy3fgBhD1ZK2g1o5ImdpM1LRG+ftTnqegd/gr7UBLXNYdvE
EwLil7A6uhTOoFbZPZrq75WFEcHmlemmJgQCKfI3iZPv9rsRYkD/48aSVMpsjCgSK9iJ6cDF11YS
+P6/mHLCPwCjJnEIOJkSO0x4ilFl0c993s7P5zzyDApCo6aJLVTdxYzZUdTmkfFzP2I+HPArC9Ee
hAEWxrAa4M74bIxTGGvLwR6QB4NEJCXmz3uvYXKF//tOZKFLwOXXT1a5BNe+bJESUAu0ME979/Y7
D7i2D6yqDsI49PbKEvoO5SKZvLmkfltRtkdc2KTcFCkmmYN9FSQboa9FC4p1rDLep5aQxao3+gZa
YbWGsD1cSGH3MAGxQtGWYpbp3AP6jY7ZvPZO927VHkjNR/RdzeBqoBdLwSUyY6z/QKjFz32ztGQi
lE7YYTp7HnlB76Xcrsc7vCm8ls9e8S+rEk8ebCW0/N+h5yaFztYyCMwRTecw6D/SCk1v0/GCgtvC
Daq31mnIhCNqiGXZn8+nyHK2fJIKVv/ggIH9IeAXoitmX0eNtQZRYkgOixm1W9wHM71tas5i1aIP
3d3o3P5d0PgmaA8KhDsqsvk5MIsp5IXo7a+twz7U706URfcxPLZPhQkswjDy2PGs0YZ8tUPXP/jM
j88EKt8jbi9SWL3IpPAGqLMaLe1qiU5+2DyctOEMMeXr9qccfMcbIgqppqJX+3wFKAurmofOAEZH
ffuEdqoS2UM+23yA9mCQ6FON21k0emzYJSGH+houT0tlb81pVYK81cu/I1niFKqmXpLzcjzk5DkO
hOc1xQc7kHQw3uRfEyZOEusINrn4flnJQH2UtfF6KePU83Q8orntES/bOTKCjLCnFMNLIwr1GNvp
czh+A1hQfBkgRlMHJ9yGEeehimBcovYI8artV0MiFQq01uK99Appm6K4z5l0FlxOiL54VF91htfL
mCu7NYmOfVpECfpFaZJuAWbJPTTD9/sitgKDUncioD2/+0/q2wq5Mm3UY0pdoFIiXkzyEMFgT3xJ
45Apoe24EHiae+EjdZKdsW6PLfxe/v88MGI48M98cBaPQFVOs3q/0wMhztR8r6U62N/KISrj78mA
7Ny4ysUo2l1GPOW6bVHWB5TjGKTj3xXOJwXaHQsEmmxBZ5oocg/YB5oR0F8S3X0lMJDCy/+AZpHu
mDlnE0ZR04BbMZ79cUx1ynUBO3558NWHtg64uz3XPZowVsWl69XDRaFtdg3CVONjheqVfkDULr0S
h6qSI1Fn8gK/gq7CMzRMyLiMyABqexSW1dQ08/v+BD++eSWV0Osqggvtpedu3GkzvROqkG1qQ/dP
GG3lbDW2ImqgSXWtjZS3sDpB0DfnbkZcSpexEnJ18uf850KNR6uwpJbkyfYFd93jscceP+BQmrkg
W1Yt87U9gFhPCA4peKebj0e6NQPQR2DuhahPmrAD6JnGAkKFtbDW8+hG6rG4IHlCnFifbYQT5d31
ojg+qzX4tLic/oi5tW9qebs0iFe4dxdyD5j0fyWJ4eiCHb/ojFIv1jVdQIsOkFdUCzFP7JNoAFtD
DwkCBa5AFDx5rQKT6xLrfv4FoSI5ribLRL/8CmTbFG2UYNyuprFOuWi9x//xLy3DqGS7d2302A0C
lJC5lB8oRyChvuKWQG40bMkoGXDvwz8ZTGscnGrxwnRvbKMzaukMic/ly/ypc0yixJ3I6jvR7G15
uc3923pkKICtuBtnaRyuyz6Zkax4g5f7K0PRYip6dzNPJFsec+ovMzn0nno2eKv4wNdQ/gRUhbbd
fXvbKc2jDDwrLhXIRFIg3mkasWCTBOXg+1TvoaTJUvbvlUJ1PONGrzlWIkKmxk4aQLRIZ4t+vRf1
Ykz7pX39VWr2cE6w4dZxtWEiQgxaxOrQL1UT/It3NLFlcpbKoeQduJuyakRMX4TKMidW1/Bu4KBk
P4k+SbMNW5AsZ3pFqax1CLBG9nIANRbyU+oiGs6BJ2Almw5Hh2eSPVqk38IfF9tiRwvLcX1shRBP
spVP+WdYQDFZGJaGh8bf/Hd8VDp9MHv7kHsu1sqstTdXq/4YzyrhE4VNPvY2gIMCgVt/i9MQFR3W
muMWgHyDn3CJ4/zX5JWv4UzLvsSyoMXGQWXxjZ8q7QceCWp/kLBxZrOabLEufvLjcCRkuKSaTa5C
aFo8C0J2hyQOpJMEClpxbwIm3M0EXBzUFMrzpD5Wag6doa53mJwICicZbUrnKvLd2ullrAzIr+Uo
W+ocVOSaWVreFeJDRp3m4a721ioqeXV3O7L5s/dnKT3ADR6Pew7TsJC8jr6VS8+Xo5HMTHHoIYhB
av1Mm1v3p1siWupaAcqNTpMCNaS4UmQjY4hxR4ysuqubCArY1Q7EZ001ebGs3ex1GgK9jUC2jS4C
xhlIqyfawvwp+vmU1M0G7J+ZHpjpqnVKOxSBO16wzrrVgPORRnKy+hWigbwglhhwJrt4N5/K+EM0
8yG3xB7k0N/PiIplrR7ST4Ljl0MTO0n/rZQ9QuvJQmeFrmVPAhtmpfUZBXe0WLgnPUl7F1JaYeVm
WK6GCHH5gCdUlhpD/TE2Qi2y4ZxZ7H6S/hlTj5RiRzUS2xAB4FAqydyViJXWVa4R5V59dBTViN+X
ZL1daHFbZjgBYsW2mCOnE7QpZbgxZX5IHmnXmANtWWJWyOMR970zDH1SI4CfoRSZTJ3f6+YVvsQ+
F3MDiKzTLPh6ns7BuaDavPB5/DHu4diF8+n7pv+xGo/H49Gx5UDekmibfILpYVObBglHSAGtyUTc
KrDFldmnEtEDBWkglIY4Nvhmy75IIYJ/sq9Ofn0vyFN5sztiGfUy8LBLv20UY78wu5bbktJbBhLT
9fp5rLMq5C83re3Yh+s7c/HDb74IGjC/19kwnqRqzv5ZIm6O/xOan1PNowMGR9fm9itbwm0B+lN5
7s3MSR6FXAulHokEYOin/xiV728H8OCuxSfDCof5tboOaqZzw528SH4ixHDqjohCFf5aUJdNqfnw
xPjX3+b4KR5ORRQUmaRJMA8qSVv8I+B1ONn4iZ2Y36KqlUV+U9WJLS7EBXy6RdBBgpaiM7/IlGHV
LWD2QYd3Y/H+MPUfZ7OPVOLXxWUh2FbF/ffStLboXbK8/tfxRvXKg8ZuWC+wtnOzpViNJUFC5oPZ
cKnu5nxIHsTlMmcOPA85ur+6BTVCWID9lYohYU504PReiMe0KArFgiTxKyFWcjLkb0PPe7EOWzhB
bm9518AVk0krPBgtZT+5OvOZV9Kpnh3uSFfC5+2Pc2MMN8JCdBGJcuSDPUng8vM28jbjxM+vP98/
jFIBOUK1PQ4kh5TyLF/dMW0dxHoOsdIHJIF/GdYqfL3euwq+5lelyHdDFlI3ducZZQrEKc4L3aUE
bGLO4+vKHAaG0g73Cm85J69NR+PxuWx9ys48ProdBz6s673Wvq72syQCm4rtvWSU8hGjnqs7Esb0
nf9063l1MyPE9skq36YjXKYiLf5gxDnHYzL8Rf4qy5Qhvy+1crlq2augE6ojXa2BsA7oc84Dlumq
aitVjYdOTG8UYTCRwLvyGqeg5wBD8HlWfxIdH4bnqWQHjyIpvXpSoAqCSX7usSFcUP94V65Sg4Xn
ak0knVKg3MqKKAM3DakAmauzsMhEtcjUwtFpo0u/QxeT5D22meQscZUBZ/unrW/ft9L7OpU4AT94
TpZknQGZmMLbUsuVa7x9c2z+FAHlQzvFJtI1el3OxnbAxRUdXZZxtkm0jIsvKHU2aykGGyKPt/S/
wh/vwwoX+/6Z9hEEUV6B75EdBebSXqDXtG1IjWWCQWnp+Pg5EH+eCf2NVueQzmJ3DJXCe/00qdYQ
CvB3a0om5b+ZZX0aWIVmM4iw3+42s5gZ1wjPzfWXukussYeNdyzhnMmeBu6kDHTpjk9T042OtIx8
XCI+X1PxhJxfYnxxBTQQT2OU2I8SZ+BZr5RZmJEN445Kr2lHch4+XhcLeSuG41JBQ41CiwGIFSCE
l9rimGS0x9QVKyVmTTON0V1adY2F4MIXAwkii/2hLbADnuoIC6akPAnPQoaQmzOcrsq7hU1DNmpT
T79YIeCgT7PljvIquvUdpgZMED3Qsws4E5GQeusplY8cEHjc3F1oOaYHq+hZ9sU23tViyLVl14ba
GCuEh1M79Wp/lpbVat52jAajhBihS7AFajFz66MAkEnD/UbKoB0fRY4kAEyazq4rfuXtR2pFSBRt
+Y5eELikfmXNEX34BygeVdYMCSswc+e5e8I/gGrfOwHe/wUdejTph2GnF/8U13H/wJREkGXaGIxH
KaiPHMiHPpkfLpn6v5K+C+xIobWmIdh3zSpms4n6ylZdsMIQwKwFsQB6k5i+qzzwbY5PKvMfU2i9
c5eUVqP+9e8HrWjdHfo2mus9rwZQpuQeSzKr1U5iDBNMLgxy3A9wyqBS+RFdhMVPTka2NZBELld4
IooQmtwg7iZFcgKJM3SY60yEd7diQOCifJHnFHli8BFW2JfY2rqeRFf/t4KLELdQOadEOFFgqruu
w408eTnRNy4D5J3ggeh6WPU6PuG5fTt+gWs/gXaKdMRCfmXwO0X+YJoLghWKQ1Xja/Ct6PwyI+lV
7vKOWTDOkGK/AQrmfCfKmHVyPooqm5xtvMgFCy3gkYLpXx+uYJaXI1kXaa8QSTG47bxquV/w88iN
7dDOvM2naBn8jM02GyaS89hQ/B6J2tggcY70ML0gb2lUo16RxBbtxzKVdKOZp3THrU54hPsC4QHt
kvDsT+Rb9TKtojf5vw33zYaAoS3mZt7sGIsjCespTa3grQZZzLgAhRQGcchgtIJDPo5qGNeJInCs
Z3fKkwYPzOGktGZndRphZBURrtUNcieFWUnhMHNG6nfFFugbhLDz9ppIilJXk/85zNWQuoY8FYkj
UcFz8xheocMfxWu+s/rUO6wVLO7K0C1kab3HMSYScwm/JoaOgEmQJDpOA6IlWxU2kt062/awHggi
pbKy6HplZrJ/sRSfbFuEaKjCMoFwcCsNxHyACtaxmD57AYoUlj61NPoyVMNUoXmuqvd2yUwjbdMB
0J5GCf0nA8e4GKt6jLI5qnl5XXFyQHD9Xn/S2rhyKWXFV70guHYcBzEdr6POZQMHNqwpbojjzIWX
UzSZewb8qfihTcqiCI6CEYon37dEWGVYNQj6x4tq3uZTla/7WsfJzSkLS1pGROJ0TMibUeitnt3F
+uKAOcu33kPfwX3jXyXChBV24OooSc5uMrPcFwkjqDCcaV09Hxgh8ZUFsr2iiSPcVbA+x+oobcVh
MbxGsrFPFklJqd0zkecTNcoZnmYotlgsgjmnSWTfOPlN12LktwWvK0ZU8EYV9C8cmYUyo/jZwVfz
9D16T1YhHpdpdRaFsiLZcIGsaGIIV3TYwjZqDdKc1HouC/3DYUw1dNMV2378sxgmkWoUn+Gz7+bX
BsLwQ/VYxFlNP4Xxt3MuhiC0Us7GtcGclil9q3pdOjmu49WGAC6VHJFxMhqTP1Akf004IJdrUBkI
1BRQpqLjhKDm7yz0fiVsEyR4oXJukU4CoAa27nCZkFgCajPUzeMHLttVtKAM6e9aWsNdEMi8ERyD
cVfmnFyfA4thLUQMkVwr0qS3HOG2B8NJv8MtIyDkGOJX45ZBshCSr3VRVOJkWuuWIBr5zeOiHxxK
5Nfq2JenYE3CfU55z2yWo97PmSFWIwmro/2ok5HO/FNGG9ZKQs+fs01tAbDtA5IYe6h2/SXy+VgD
x3EV3ypgyhJamE68vmOrd9M4gmX+qZZ/R7xZ4/Met00yqqPaIBYrVt0sIlpJ1FTGK+mmwqPaAf9+
2efwxcgoSbWH8B6OS2ts+Jzb872JpLZaV5qF9b5phh0LW7ERV+m3237fTosrqijtIMLWd0V0c2Tl
vxvcX2+gvVUYCNVNcaNyeEtEyxGq/NK0491DO/Hi1TMb8odqExnyQja97g+tMV4Xd+xct4dg1tuR
xpDiIZw4RmTEEYD10m1yNtimeejgVMIbB0qaEM04M5C48KEEGuSkipJObaYoOfek6mYxTxrPc6OV
sHLjsO9Mhe0vbs/yELBajpt39iuviG+VZF5jFPRLQZ3IPunVIOZ4VSstQkv1Fuqadjy+T8xY5zSf
3rVOtyPt0Ce+pnbywelM+h9TDpCFYY+FcF54tudbvz7NpNAXoXe0kVdeyXISdlmF6a8d6PMmubZT
W1Yhgr858dDGYHlTvzlRN+GEIeFvPEqsKLChIcs+mZc37BW1HosuzhWOOGbfKU5ENchBI6Ch8C/V
f58XwtfDR8jozIjHrcUaoTxZYtuWfYvjJ7LzdP59A5CFambXhXuwZ1Wu/vgG2BS2NSIugJkzpRn7
MfR47nVbkZKJRxG1umfO/orjaFp+svhZxssu5rmoXJkdmV4Nx026l7vD3ZHz8Re/vniIjqRDR3y4
sC0ROshh4bldX9XgoV8wB5Sp5poWVoHEAgIREoS+CFyZ35peCkjOsEvPpNP+DmXfqQmvbM+B6tHe
zJxf98okd+Ki7N8DSGaXB6oOXdrUzQsWuLHrH+zHMa3ciQ7yzvj8mHbyJCIcKymYnG7BjUlN8xFq
BCMoDr+i0hbWf6O0InYjXMjggYGDtrZ5PsPFFoONfQC9tE6kE2JNuNQYdm5+MKvYFze4AYC9SwAQ
ylr0Yz1ZmRofXeJnCh9P20SEKcbwnXUGnpUiHsa46uaKQaH35mVrkviu99cSqE1SY3VgsdTTlT3F
ZWnk8xL9SSVe0TnqxnXRL1ftOS/sbK52Zb+bJxWf6JacyBKXSKg7fJoChxv7XijY0imBKOcP+3hV
sbyWxMiftJ1t68ZdpJCZA0qcsCXODy92aKMnVfYBN4VrB9PDurYHQcEv2qpNXJb1O4LyBKSFCtm7
eIS1IGnrcBdyRKvm+ufbMKxvI+fBA2sgE5QdG2PugufSrynCzA+Z8gdpUboRujO350HwdGt2iPLE
5eAOk87grZ5AQVhXmaBvDmJps95y5R0SMIIWdVP7PGAyp3Lw94L2uCAl58Q7GNWJZATjYb10EdiP
hCUvJ2842DEhuE8GipoluCFRL139OjDm2cj2iaq+G29/JKLhoddCf7uu5R+tLd8babvGomZpfE9X
fLEZMp214HJ9XWzUFBeUmFYG/l47bVqqa74XGaGobWT9uOisoxqHC1UnVl2JtmVARTJmBA59H64P
oLpVQsbrSzVAOs0ME+9eMF4DOx2AgJ/wz8PAkFRmGdzW8nvKFUpLxqVOw+6Zrvyx2ZINlZ3yjZfk
QZV7F+3puoDK91s4yWST2VEBZ0zWFURtNUO32lUo5AbEwG+96MuSe0dOXcDetqXFhfJX34yiN551
BicCB7A046cg3j+KoTdK5e/ROeieuAt1OswJEMnd0UPBW5KbiAukQW4VCK6KxRAAHtkWGPTM3bA6
qrnVs+1X+QLPaNO+FBHDq8AJrnWgeQdkXghJbXaQ+MbIgDi92kSpq00H8XIx1onymZgswWZJ0cut
IHm7O3toGbl+FSM2m0ARRcCXrpg/JdwThEg32S+IpYo40Apsq04GpR29dmW0PBY4u0ZlbtmVXiCS
NqCIfYDzAqUhRzK60JCtBkSGlOyK88kasT8y/aWYlXF7A/WOznHZ6XLCfLajEARENqSSDpSekPQS
5jSxKJAwEdYeRGYTN+C/Z5CcNdd3kcNZgVGGqDweESiyTQInGRXZjGmIV7AH+nJgCiMVyXN+zYiD
M1zbTMJJSGJ6GpkUb8l8i03CC7K+fjMi8VJIatgplNX5JG6mVSBVTW0vGb7+nGWPag1btKGreRHM
oNu7KmsTi5n6ONTvKQsU6uYKxM4JFSZfE61qPjh59VokeoJRQRTtC+rVltXaScZhg9lQTs2jf3Up
li8LxXFjf86o9c4gOxpSBTEXC7ed6PJUeMZo4C6VN6nU7RdVo0SlVPeL0Hvs+pdq7oil+lpj9sow
D6S6OnHo09kwqcBOqPH1GGezj0Bc855m5y7RJhLaADUmGWX+zipb8rEyb7DGlGnsix98I4tHy8O9
A/YzA71grg9lHUUmrCT2QYIx8z3EtszUcNXfffj3oCbtcS9fcwZMEcdpiftNIN1kU7c01fkn/isW
Xm/fJwpZCFw5GCi7KU/tVlHcNqhyB5NlKVqQJZUbCj59+Q7aJRwhFaQeK07kZxpkTBrbXw+K/Gyq
cUBv4GeKozz4Vp/zkRL49cDik/dyGd5O75JDrBklN8ePMQYQyOsrexZ69YAgBPxv1hj18H1+rgW0
l7PMV51gn7RVWg4qV4Mrmakf44fJsw4AuFG+ZQtB2lfdzDXIivNJytgV9SBWAfgQtxD3U6XwHrJS
quW/Y2srM9PFVb5UlFYs95Jnspr7Yq/nGXFrvwF4f3aKJxTxNmbs9S8fWJtqFw6jhxav97SQAJyK
HOByoNC4aissaf3H2nADaf8d9wuoVNpyc4GEdDykuCqxhtXYw2o1TACCfqzgJrkSPWbRDLnll+0j
5bY8RcvQUc7WpOkiODkHtRb+/1a2bnyMje+QdD+5S+pWGRYv6PdHI5N61X4mbJzl5nIItUsshgGV
6cSHH68DjtimafwGJjm/bfxOHk4zkgvj5dasELD1lbaAqRMhFPs1mfy6ESc8QQ4YA6eMhc+rgykI
RMzWjYxQbxXvlqrGJq2xT/m5CNQawe3PpGREXCe87CukH488EmDB8UEcBZ0oyZppAVIc3Md86UjK
aTO1ZB4vi8fFwtsZ6djW26EBmwZf59GFbbTBt9LU7B2C5q5do1dAPq4TfQ1LV2lRoX/s1J+YOcKZ
dUnRQnd3gsTl2t0QMczXBjp6WtTZT2fiNgXY63Y8EuSDS7bXTBj0L04UX/nl9bdy1w4LJolqHENM
vGmgRC0Fq3I4M6eRqT6TgOgfNqxABxjnju6sWFOL09QxoNoPklyImnO0L+bvnW6c4DszzRm3T9hF
CgwvpJ7bUVhxEY6F7DxCSClFjWImRuU82kpjeWs4bqhvfeuYnD6l25LMM9w4c5+Xf+RmCicjx0rS
ivw9gV4ieNvqKu56a8pdPx4HA8RKnXcH7mdqpBId52EZKZwaAin+WuzgM+CFWvpjWptdzCj9qpZL
EflDyHa/uRdrMkRdHIOrcMKDv5tkCcXbCGfy8SeCm/WiBu9Hjr4Ey5QwqMYNChYbfTStpPV558IC
qvR3I0Mw1V8pwoePJc49QE4aUuvqM69Uv73r1EfI4zRRrE+Xn8sX4//9jQT4X5s3WeUNrjqlzIQE
qK1nQlR3UFTgcDLGqN43pkzSJgFiQQnkoU9bFEvfYN3fHjTh0EKIIG/s3cU5TtNQEXFql2C7GvuF
rZadoQYNDjs4Gua4AitybS6SA4sz0c9RhEu3QrLdBr3yoPcgdXh+MZB3L7kLfFJ+jdo6W+TbixpA
KnRDyev+niVPfYCBjo+M6KUAFUUJi9f8651IgMEc35XtaCqUdU/87TA2R/riDppHaplF1S4bSLli
pVjet5CsjIJbIzPBfvJAJ0yo/KoetExBp0K85iDTc7WnU/rDj1Ltq2+bxycyGjiHt6v0niZXixv7
cbwvD/EN2Qf/RXIDBuvS5nbIAv6KFoMLI99xlpNzrtSEE90oPlV/Y6oPOtpyIcXlsD7HWsXJr9Gl
AqX82d1QvkmlsF6vw/2mJeqP9G139F3C00wOOQEP+wTB2uxHbwkdZv9+fmibwIdygT5xJ7SVRK5E
xDdndpbUIw8CmidZ2YaTe0TBc2Ppe5PnH4U8swCZaSe3buxqw3y/AUsLXd7pOjwZGz7XrfTw8K6H
9YIgSthGOFHQsukeY8FMkZt7tHEazl1Ho4dtAldCIAmvUrqogZ5rl/qP7S+DDvm157sCyqQ9twJ7
E0bZ90tc2URhcXY2fcwXNy0se5SqlskNwyK1W6mlhg1tmNhp+jSzx8mW8C3lVu0h+QNewyZJy7E/
GbPCNmj1uDFBc+H9FtvPxxlvmaMcXWzXZEKXK7VRU1w5DF7suxNVftY/Y/ra2FYFhSBHS0SoigWm
azVhmO5VENAh4cno7ROeh/gBHKtcb31nnMNSTiW7NO9ojMO4IXowUcl9KFNrgyyR+on5ARt4kwmS
7PQoPaWdy5RepFfJ0Cx8zkSxpo6pLAdjWYT4pg3Z8e6D7kvuvowrJ14wSAgVotQM8M53+QDhph+l
Hw7lvlFgRPkph9J7R3QSBfz4cQodkICX66elUnR3GqssIhIDfq5kSvkFFk8YrPtUaHTqB3+TgttK
qDoapFS0sEZI04wr34K1ebrHE28wqrkKVjIIjLBnsNXWLFeQb85Ye9FXr3f4vFp+h0muOwOTIky6
9RYmVF6UdGwpLRKdpAarPlUOAQaU/3sjEgXX69pk548KLvNxgXyyVPZdql9fTYUAv3u2l/9s0f0Q
7Mf6f5Kk8MgGO4adK34TxnMMl+g22O8zQc/AJ51JvHV4UJpxplyj+Gd30zas6KCcUHfEvBblVWch
333nelFC8oJu883Pj+9ADhfCbqGS1IzJIiQJahKjnTG7IWlatfl1tMxDbfEmg8uNL4TBsgEXdcAp
FL9Lcbq6Gs735PRy0u+b3osw0UjvU9r6kcjxRVPQB0uYjnBqPAf+sS7LmLQhSYFZnftXUQ85ZX3b
L274+k7rVUbet4syFUU/qe7k9bwGrKdZ4q3lUS5y0dM1oR1VPQz0oX6u9/RV9I6W1PISogs7Lj0O
ASJzxZAi6MGLC1s6NC+si+MBlqhRN/QtPamkC8BxSAwV1EmaDNcPyHRMGzEGoSKlAs/4lz8+6OzL
nnpB9ZXsiyjwovbaEzHMAE0eVUbYpU8byvQ4N3KDcopYyeMCn3DLz3fiIu4C+AqafzMUSPLCEuME
gDkMxfjUj9jiona+NVr//hLjsA+MT/zhWHf2u6SzTCBIrYyRi+mvPQuOILFTWtlkl1QBhp5zt0nh
5o0MEHdEJdJ5j9k/YJllYLzt1rqGuNIGRIXG+QgZIla3O6aqhQRbKT4QHDBiQgXdXaQlkmlxOnjE
gI4XDdQebP0TkvTkiB66njWrYDmr5QAzCPuJ7e6u4Rc8Qgp+1QtZuJ56ZCQxd5lhhiGBo8BP5IYX
+kxD3fdhOwG39M3kiZfKpOm+I6EVQRLUaLkgsRrYOCTsdyw1QAvSe02VEtX3a1tRy/fQf0bKs8/C
El11BvJjYcgasxVQ6Xy9JEbul3v7ltfMaYP2HaHpOTrGb5H17rZ7wWXSo17tx1N09PgCYXgCHy7D
UKfqmqfLKA81YT0XRdfIYASnivP8ZVl5mYg/fyJUCt+YkWhJJAYnhW21f5QlFvlIzEUUu/z/zy9o
sL3uBSlVBl3uRfd4GPQfPYwXvCxJAukw6hxlirweYm5+UflBPuKN5zws9HAwBKtU7ObxKQA+pSHj
MAr8+X6AjmzPqj62PChnnX99eUEqeRgoER+waKoKduSdjsUuAwX5NNQAOAe8H93hn7gB+VNuxNWu
jVWJC3TBzrV/fFyVlRnb5E8K2Iu9pu7pgl0FIetEwwExGVpIYOoduR/Tf91gMtiq/RiO8M8wcvYH
0wChoKU0KethFOANwBzmnzEQ2CDQXUA5NAicf+JQ6vN4iiWEGNF02vIeb6dnzK/dl7xeEGltDew9
lYULZgEJGSA6e/sdlBVy4qjRdPT89M3vvFVa8vZDJUunmGjg+TzLfN/kUaNXypYfMClU+b62o9Jc
0QEV7y5ke/LwDjsA+Yez0wTqdpA0s7CTXsL6Bd+Q92q7UQGWNMtNndVNfas2OFCg6wlZAV7jLYOe
QMYeoknoEwJIJXfsQr/WC2cS7Ru9bClDrE1IPTCOnn+fGxLGoPGLxGji7N4Q3NG/HaXgmtWdagGY
kK5L+G/WVcEe7GSWDq/LBo9lYkBvCPlPpirdUDtfAP1ZUoQK+a1B/Zqp6bUXYvVWd1hJEkgEynIP
gkbPyyrQvodb8WuGWkTZ3YDyvbqi/jurW7A/vri9ucTV2ssIUp0NxQjyAsXhgQ7t77Q1kW4bUefd
DjB/FRmc3a/mDMjuECwLUbJQy5FgUZAq94F6t9zrwhCXnwkMYeCwXwP5kWIO1Kcw96yDqEqmNJ0z
0J70vmOBFRVqiIN+C6mkCjLw8Kjbe4V1VY6EA8AnU6gPKPXPv1+ObXk5z/19Qeu6vkW+m4rT8v6c
UqH6ArHkdnuSsSF5DUCSuleBUkH1VjwAmXdWUVv8ovmCQ1INQZWLlNkhpuouK23+3uOXNaiIVAvZ
65huaBBjGvLcr0sQpZ1dChZYODt6g5YR5zDEctFE9BUSNEMKM2x7uVpjIJnqlzHnT4Apt7fIen39
+yAzAUARLS0B/6SgaqDedQ9B8Ea2XVMS2FGyi1Esg1gk/dgOBZ70/TFa7J1b3jFpLFfejk1+cwWV
BCxLbjXa7EU21alqeRUuW54tyA9zUI+y5UBoV+ac+tQmDgbi8u7OzD6E7vlEW+OcH8Hx+LeelgfF
ylgH3OJF59fTo8PntbCUlWb7RX+yqEsq2EqTxP4RknRN7EphPLsl6KymvbY4pnzFfg/vaqpjyNks
U3mmvsSFE8POHK4bCWl+XfhKP/zxxWMcCgou51TBDe3AGASH7MRkAbnDhCHUqeWWwT7cQHmshFX4
ccs/JPkeRrST1PvcwtrTtWxJqPzYgXz6Hx/1TQr0OourKB7Q+ja71+4dYIuo2Nv20MeCzvrYS1TQ
3Da095S39sfJqArNEMRehDxbG54IoQ/ItjwGdXpzPdNvbM2RxLSfcf65znuSsGkg58fof5/RrrSe
HAureGmTHvsevLtXN/JAL4UF1S7xZexrtg21HqC0TwGsHUtTTGVrJa9P9GoRJDDySLcR2LUmPe9k
zIHb9M+Zdndd0PjxHY5qd5dVsiQZ4uTlh2M+MjpyGxqEzYwr5sYw16jonCJw98XwOdGPW519JiOq
z2BA4QDszMbQ4OYtxxTPhjClx6P6OEKeHD4tVfXjjrFHFp6437LJfE3zbPYFYUrCqZyafeJ0aDen
uPH2J4w3EjqkCrwOeaS0tCoJcZaa3OJb2Gv1Cq/FTkk10BALgza3MFdvz/J+XdykTxvE/V1116Vi
JfN0sGh3p3WIpmIh2P8Xn2WIR5D5hcEosSirrHvo5YZm8HXp1MKE0C9Tk/vJUhRBrzYkY/s7EY7j
JUvQO3IcJmFX3fpM8PiUQEGTdnu/SY+pABn5TTxSJBVOjYaRxNYyih13qSIv16tiVPAqiyA1AsXy
5Dpu2O111z+NhEM6mHS++dTaxkYd1jDhlsssy4+zkpOVx7JbBqYEbtXyJ+E4LmMp0F4ghfJ0skT0
+yDz5x0PqSsGapO9LrufLN3mtYU++sSup/ngS+NKFvssYLzfiPwz6idNFE9AdZP16c1xlnhM+Zu1
CAb/Jx3yX3xa3g7a8RMuV/WbLvrbxg6lYJ+KCAn/Eh9ysIDeMnMaW47iUPSc+SYxZ8hsG1s/5uQV
tvxtymIUjqfG28QuXOB4YB/raUyLfbOwuFt6zoYWLBnHO/CDgvF697VNPa36eBdlAm9t4QlYf3c9
uGG892AROIC5OiBRJeocyRI3v9BXO4SBvtnw0F2sX5JK40k7vrfvQBwoTcqvaG74IvAK2GfBBXoS
LvCE5mdFzc3gqAT44cBdlODdoF+KRtgr5LirElHO+6+akgr80xaGTbvGh6VS2MAicAjDZuE+lkIo
tS3YwiCDRkScEAyDc39TIIjreASPhkaqfrD48cOzyLORGBKHKMiXuWen/sG5Pbu0Q16lKJ7mzBRe
+W82ALq+/bIe2sNVUtEWh2qezaPECe03t18ULFYGroB+tzlp8lHeYPLpOGys6ujTsuX4x8jBNoMh
f+FnurjrxUGzNLzramnMIhoFoqV8D6cHRHiQAPrS4qSCQ8ZeKubH6+XswVqm4KXEcUUB1Lu+1UFU
NMyVyGJrm/0fnyBAhqGPswYrL6VNFhsUNxd/d63Kefezz8hD/eYndkQi8980jm+QfUL5Q8oRXLlS
tenzNtF/VDIy7O+CRwojiPgByCQP6IQQedE8QAwq29UhG59E+t+xnTEGovDhMAgeRRIjBMMbRLlI
8rXYcJZfCJd4zV+dVNkAT8Qyq3H4W5K04G/2ZWOpXJH2cD3csC7TGmjCihdM0h6veJLqMZgZBkZ+
ldSSkv/CUGFknQhv/nYYDK3qK/VZSGk7omjXYhAHVLt2XE0JFfnyLv+AYEX2KOCBOW6CNId4hlUm
eew17BY/CjM2kRsfWrhOu25bv6KephYFSbjgMGHswJYcxHxUsUJRuU4MAJvBq9gfMsox7jrUKTyi
gtKgyAvilSUQ+E3LOiFDbZjN42i32bx6KfP/+KAwYAagtpnP6PV4wJDjw0vK1ZUGtbF6xcoCIe/5
KclZGsqgktCEgqKFyb1YCaKgYydquW4juJ3aFiwuP29g8SKPewz4ISurLeUzLLyfdBe6ImLccvv3
9Sy5Y130hPh5MF5+HryOenCBfnVcc9JNmASwJe6mQgBb0CDbZNTe6/ELcBEsMW2b/Uf6bwOcrI84
wMwXHymCaDuyNI64o9pmUUsFN3+RLK56F2Ao4C5EHZhhPtBWbenmf74FphC0VR8RzrNGqAN9lZXt
lV4PDSe0aelrURPHPHIsWfCn++xv/Jlxw6gDe1qwyd5urOLKiEcIazb6nRke5zPJCiTFlV8+qqq1
jh+232VA5v6qIjNVw+c9SvEQovD6SX+B5623/K5xF9EVoQ9uaBdQHRKh+YR5sNgMLRQBrSNxj6iG
jBxofBZjcNxUyr/NLX6BWewUhV43IrYBih6spDpP0tLBxqxns/Um/xNZ3UwZziqj7rZs7FckYTex
elNfCAaLxUvwRwqbpJ+5A4GrQl3v24GJn2o2fm7fdT8ilJqyqzvxJBX6wPBATWzwBjTJNqrqLgl9
xSTK47/e9g5hKTTuu1CdxG+M1/wz4/f4F/6GpbMOSCvZsjaaqyXVxqTsvsWk0FUwPLvNOAkzjw6G
khQyBPNO1snqVDC/YX5uBBA7lI6yEDI44M4OnGFl95aJZjCKf5Z5QbJGZyRkyNbo0iAzMYE2q/gv
+/teYNiErbIpaxPnpSVetF20+LTinxKf92JyA/McZ/nWtX9DoRGodmongI1tEa8hMJgL1vcE92sE
q06XUB7HjoCYQsuqfSnKjkiUADqRvF3GGoJ6i6sHJlhtKa3VRNI7E7p/ccu7p2gOUF5X+cnqHUCb
2FMusPb0/at9VcO8IYHTdIgZVkaBglybYiyQea5A7n/oClSd6zvNyk/XxwB7bv6YYpC3OV5u0+qA
C4soyX304cw2FGBAjG9cCw0reBg6+Oky6FYU7w3e/n1iRpgCzpbkymSiYXXjCMq6INoZz7OoV7wl
/vYtG4ObRxOhTETaKvSjPccJqDK7WURCbbg5SaKfaBzpkPjI0VGsD8x2JcaIbMbBt7xnCmpV5GHy
nBoUhI+NpPrdqYUui0ACqVgPnJ77mWNV10rDii50cVMuV6Ldjz2pRd7brKvQk+RdYivsOx4PVAqI
UN0K34ptvl7cWx9AGFyWXeObyEQoH9xEuduGvcGjLivrFHxNKDRfUI6NeEBFdbRQ82bNrIu0XDy3
RlQ2eSpVHLjAVOdKJdU7FqCOmRxHYbxdNqe/u8czM/XcfpoDos9bOLbinV4KZRAYfV9qDT4mj1G8
NIoUB651wmlJ7SZ0mHHwoIDyTUwlcEtPv2mtquNRs34NvXuflpFQ5wfyLbY9kEPeK3kqn7xM0mhN
dhBAsOP9zHq6AtOvB5IHwM4W/5q8ywkkMsekD4k/4tOP4ZABGFiQgr85QrzDJ6decxLdTN15VuS8
U7rQG+LokoB4IbMYXSAUsIxTth3PekRN8DpGGTCCTC4qej22JJ/uQZOZzjQOPmThZGEm+J9yo4hg
Dogo2bIr12BTmRB2xxb2BAtPlny1w5FWflAiuHvkuvr4+AIdJ/e1oF2jWE16QjSCgzpsxiwjvVrl
cBdmRy8NGxO69PmYFZed/LXxU0YqQ/zM57SmG5nNzar5PiNUGikIyf5Uyn5U5eIq7DaEfVnAMg4n
HalqxkwTNPJRCxNZtcdVOuIAVQFDI3bRjwY95wK9ohn/SjFuCB7BkjH5QHVQkAebEFFj3VymLeZX
7Vyy7M5NgoWYTXuiN6fixGyHS/kOHbIgkzDnihCIiS18+QC02+Jmg5ni54aReTEXuke1AH+neQS8
aSFreSs/CJgkvH9f5p559TqHFKAaw9zXz35ZVdCV/t0f7JSDE5+51sF9p6oodvOdj+EadOHIqb1u
TIvgO/LH/yWnLqRyyJc1+NffBnAHOXtjhmoSI2UWtfIMcCdzoAaJ7q2JSnVxL7XQ9i13WwQT112G
CTKeTfbIQdiKntkWlTSnRnDreirRRzpEppzBBVdff9x5lHb1ApA+rJXGH5d1LeZixWHhz3aE0lQB
ctWyfKgmFWdQnmIYiWji1LxvXgr6OOTK0lv5nMWPYLU32XjpVfxoHegoYfqsQI52wEGt9Ahybbae
GS5ThfDARGVjWqggRarNiBaEYMzax2ooOVW3xvNn7A4l+6yB77JGoCCJn8qWi7tEpvIBnm8MSCe9
CuOG4PIlDcwN7SlHn74X3c+aUYHdAjimfgSJHcKc4jK13h7SAwDM/wbQ04dxLYzoF4e2muYWvm1Y
Btw+YCtIxsMthiU55HMbh5eZyQYLXsn0DoS6iGfeQ7Hs6flsM9YnACMPZh6pbvVfqunYY0bDZFWk
E4BSZDgd92iYV29+Wtxybaeyn8iCCOHXxBuKYmgzDn/qwWinP8LysxVfBlxcELV7fxIWRBbGw0ks
xPawXjZ0BYXJXxSfX+LP4KVRuSRAvvRox6UUarx5jmzKp6Zv1EiBq+6brl/MEyusHprbpr96BJ29
A1r62TQxaZgbQ+kMD3b+LtChLmGS+EFKX1GCVpPOtSF1LL9G6BVy7quLjAadTCKkGxFvp5GK7Xqd
9AjH+tgPOJSbneUe6/XlS53Mv2d3hgprVkBOP2MJstiS8IMRbF4PY0mP5bx7GcXNm1yW3J+43oEU
jJDP7Ij0ZKlDLWNZLbJsDr46slrAQ/FHk4V4E4Q+kOrIngw7XBg01FlqWejsoGvnI9YHmJBkSNVF
kHuxW+t/Z8+n/AlWFVqCt3bY0VEjLvf8OZ3khyvFohUOH0auHIfjYU6D44BAmjcA81AkIKiDe7m9
AgPob2idenia+wmytRn6qNtGCXFk6YTGMWLXsXj1/v+GBfN22cJJcQBxGrUu0Uv/FC9IW2st3W8A
BVrPXyF63kt95T0H5JjPsoE6UqEUU+olM04KITrtvRxB9Ok90I/SNBX0bZtNOVmlJ7rE2ORbZQy+
Qrnfbc2PfQkCX4+lbzcSscfN6KEjykD2a44do5xAyaNExT91u0+W4c1w4L41Gw9ohUNnDr/vc3Wv
ODY3mZtnPx6DUCjQxuVrKoLZ3WhenhkI7itQkiCG8mmLEH790X3VYcoKwZCDE58riSbieFOx4OYA
XYnS2+uPTuTM/EJ0393qKhIWYi4VQ8gT7eqltPwjObNqVWN6kA8Yjdi1/zi7e1zqJDEKb6Xc6Lxz
SBaqn5JDhZXUEObZOo46mVrBf4XSfvPvWdSUO8W6/Rqogc1w1DfR1WzzINP9y4794UMsbbuTWyEo
IPPhuTJTuQhIDfiFM6e2POUz47Dfhd0kCnqDl/yhsaDhhamlrIxt4Ah7aiGjb4hwdcJ3AQBPjeCl
8AOx4L94BIxiuJkXy3nUcSuxKa0+ToW+t2bjb0Ls2sTTPqZcr2xaIi24rMEIqeMRp1H5iPoZ8LsB
P+vHqp2Wwrkz7LnBDT2UGVu+SFljWELShkaYWa5BHxDKmZeOITxgiAakwwbTwaGzUubqJ9q+CuQ1
94JwgLLIjfTEyDqT16E70REeDucQFzYVsjdpyr4wREZkVzcJy4ME/kojZ+68GhYY4ktYW2C8VX2w
yITcNUlwHcq/8G9701hAh8vKe67n21nxrRRL39XjymkmQf/Guo+98ByR/2NnbZwv8ROO/fW+8Vx9
tRT4CB0fQl5Zrj2k6PtJBdg2SuVgOqOm1cNnioMQV0oct3rel6tSMyJchxfU9KB2hgC33ubifN6O
/xQOK2Qb/tcA0ihaxKzUBKjnTQwZhoGN9W/d98CJiWZd98NTAcQ2YnPIPl3TLK0YO21VW0jZ5sJQ
n/TM2LwlMFP0fccs9lIl/yXimLmMarjskmWuDk37qogmayryJoyRAGW6gniufkUgIl30aS5QP0Er
mEKOWNkwtec+4Fyhfj+MSx7y8wWEmr1lUWFkZ1OreUfPeTm2GX1tduPwghwBuTCvremjvNLNH5xT
+j7uxWBjj7QUkJiAPKaH6BuGjD384bdC0bAcVDDvJavYgY/d581B/usLgraANJ+Cm1hSJifwOh6m
hMGU9jeiMCSknU67ZGPf8JGuJAexy20ayNTcF369ShPwfJ7svGmXnWEfoZ+r/cFN1h54TxNbvU/f
qIlA6wF3iMp1A/1JN83Xne2vsOgrNfUPmrwZSA0Frq9peRAO/c+/bHWPXZgQN2xL1eYfzauAW3mi
EHIsfwuVnQOeLdHZotbqqcfbiAfzuY8GdkB1/Aep+Wvby2ZdFImrSaAIkNBbOjA01rwnoVRC6pcn
MSlwu4I+x/jJvqcY0f5y0FX7gHc7h0BCFq49srEkyGXr1JYAoJlwFeoLbo1uC59010vTetOV2nHJ
0LySmq2LDdlRddjQiroM0KCapdzgs15G3T12r9+lOQOLoeuWF5hsAPcs7KCHi2Wph+mnVDuhO/as
OpDu4tlk6nCpJBvAmViI/hCzd5qzX9EL7StIcL7mGpYkDdOSy3nRRMdbrr7NUZg2vOVkr0Ah+qEX
qaZh0jhXD75YLcdL1bdZbozkL1HdnGS07BZze2sEzcE5HBxmoTT97faD3ccvRU+xfh76Wh4I/a2x
g4c6Wcsc6Bzd7MlfD/PlByi4MgPlAkTkqh9mKKc40o+QWpmBrRfKkkVa8favcVuOVgeKFqfmn/Ar
QFSd2+N9GhVtMDRYIDNSBUxr3oBaFKqPxZgLTs0hyutK0BraL/Ol+7Z+MejnGT9A7qSsOR+S1oeP
T4aFozDZlTqMMNp3LvS0H7l+bK0QJDzugo1U6/AsSKKIueJE8G6TA59Yly74uqnWh2dsPA09G0ed
iTVk8ES+J9lXUzZwk/880tEF2ajxAMs1IebB43fxt0rwKZ702OKjM3W/CVajWv1Tip3sI9mYfvoe
J2Ur5KgAZjQoKAkMsMDE4HEoSIecg6OS8iK4iKUGJTve3q0KXpojY48vXOdd3p4D9zdohDA9c0/g
X/LdUVgSuZefsPXY4EJWcwQ6ZuyK/jgM6/YXZfuwWsvax3505hdkg01/xTQ7KahHJ8alFwwvuZ28
NmOBdaA3w6tuN/HdWLMFIyjLwoGYdv5VsrKKwaL/JEJT5QH87+CcnQmYGY0g3IxdIxrDcDFCu6Ra
o90WHsSF0DpDyNUcse0SiyO2wau8/YQNqZYBATSh+TtPUNaizqRZSgP5XF9vQciHYvYk5GjPJOjR
IOCr7MSniDM5xhs6aCkn8RhDuBehm+aSIW28V2c+YPFLpa65Ls8bORdG+EoZomoLpmwedhUvVH19
gkV42EtT5+yjYdJaB3VcKXrxPzlbgkOiKfY8qekehjjVnjYXBetBhHNOeVcdNdP0Mlt01LRREx1l
oS8BvCEs9JQfvntuqKsRGgNjY/Clw3h4E1Uqz9fSWtFnjrRcBTZjIR6Y4RBAcGqhdLt9QeXsXuno
+8pjm+cy3Hop6am5jO6ZgdS5Bsk+lG3i7b8q2f3CUk9EcDoeFfu43yvpTD8G0BImt8LYmGhkCDdR
ig+N90c/kBCwcVFE30weQeDknITfTP1VrMJeKg+VnVj4Fli/QD+QZFMAZNS05doiKoKOmsFSOJgk
H2/KQyryXOB/JpnmEhNXSdkl4EQZP0eKLnsCUGiV8Zxqy8orGm/c/WmfBXtVXey1HzobSi+jSmrG
Q7PSVkE5QsNiPWS9HVaw/a/dVr+Jzfh9xONa3U4wm0u9qgy3vgsLdeRxJdpGbmntsjSilSt/nSWH
04HeOvuImn+kPFZCa0+RkIV2EX+O2qmK1hoVg4vKsNHfTacVe1bF1Ad+E1VHRCRTn19vozlhnwI7
DFn8/5QI9RJJT/3NomtSbG2Lmlx9Yv5MP8TjCO/mBuAt+Hz+7I+HaettsxjmCfTblKU5oQSJ6xu/
MTncEVxpEuGf96TWrfnXXL5Yh3KGwVOEsc/LkrL87z4uEXdIbsEAPD6swa2b52+x+Qy5UZdU9Mks
i2g63Rz8R+S8Q3lc6CbqzQ1RWpZ/T45wKzHJOcnftFnrhYMNVMuoBzkk04AABJyC1DXdswXJkNgg
+IMi/nKoNG2AdJNkaRNKTum/wCmnej4tzwc5L7v3r+YTo5tTkRVF/1M7crjLhBGdsGdZM8Yx203q
pOZ0w5JIWVzvAegVqgc8OEOkZNB2LAKwn8Hh2NgGqwvs5642ggV+UcpwagqIQY4Tmw5J8GTRewyu
J53BcAbq89zlIFpESxak9atV2RRLk5xIgNy0bII8KIjLpf1zRmbGJzgULuylxjGtdmLXhzlWrudj
ELi8sBL1I2sNBlSkYAF/Tky+9QNyRsNGeFErnCu4x6QhL0lCJ6MbPYIIGlBDtEg+F3Zz8zPzOhni
IH/e6m7o2hI4yCMk+Z/Fd3W8aClq3pRNRj5KVr8dqcAub5ZXkUzkS/K+0M605CUfgMcWp0ZGdJNH
zVPA4P1NPZflu5r0ubx5ou+mR73PWflMR9cmddcgk/PDI76a+ZnhAgdtETo4Yzyx7Q1BXxOvJDDQ
1LTkRnMhzFClJdSeV2k70th7JJ38YPy2mwjDM8YnYQyq5QSYb7En4fP2EJYgBPlyoibFMiNM2SK2
wxkOKansxxbE7H6P+37ozp/lgXv6nYPc3fbWaJYPjmrfbp4vU2GYX/OyAeEU/0BzLR6PTpfYh8IL
Kh4RIeZps2k/yLIVHOfavs12GZKjFaDX8wJqTqc8cdS4MqRi93RVuZwv0OHmM2AsBguAXqAEGPii
rE4n3ereVMSTFjxMOce925HhSN8Mm0KRFcWi8CFQEvq+qFvj35fYgtS2xk4zvmmdasP5D6VXM5CT
eiB+/C+6JPC9oDnlu6n1zRhzkjoyLTXu1NMhqIGyAj2Nao/R2eRgNKIIpxo7y3DUdaXSgiRJCqf3
f12f2bK2XN+8OLTmwRbbIFI92GA+H2gUsCWMCq6rmkl1ipgFos1ADvbX2NboXb+VBtY/Ido/aooH
goQ37Hv2KrjS2LAcU0p6yGcsBWvckLlpRxdex921fNC7pcMKDfovB0IT01yVOeh7eR3dyEVX/IEj
ZZoywjmrunIZ7xsYChbz4YHN2LetzeB9i/xsVPc6HavJLCF6T8DCqGqc1MsuDIouKTU7MjYx1HHh
qqO5SUPHNk11K+XRSMkCdZD+uGWk+Rh/0mfthTHzZkvtt90MGOaazFQYSN6CGN/+fT14rsP+whhp
8d6aCgZuURXhNWe0uGXfRgpq4WT8y8092gqfBInSIzq3tttjZIo+5x/ab/qK1Czr5al290zZmIcM
luGAGcYriNPItpei+UgxS1bFBToJmB6/94o3bsyZHv0pV93Yc+FmG+PwOgf/nclxM8SM9np5xxix
7rUzPMC8XiLm0auU2xRbLA33LPiM3E0xLbpDbFH7/VzjMQn6DRUTriLqfPUDJqS3x/jRwkiCvfwJ
JlLRm0vH7Ge/SVHbUonaRnuopGzwLYRF4L/QL+i7Bwj5lyXPGP7yisZyIweuhQgTVk/JoDWwKgFL
i3AW+G4+ZOON+S1Hvix+yoHA04b1akuWvUsVwlNuQERbVmrX0m5HIkrsS/UkaiFWwbWUlCkFyOXk
AopqdNzKHMnVMbI4rWOvjE0Ef3ZOdLuDo0M+hBlqmLquKp/xhJjtwVrj6hHDtOoNV+9Dp8HJzXo+
YULFSGuPguf7rfURu/et4MUcsfEVZoqNzyMQf+xplXS+7LqKdOb7sBwcA0k6tCwzURT1hua7+NeM
tPLgZBI60tylyQNovn2RVjxrN9Uv3zwRya0Szh414MPmVzIFmGG7b2Nrqep1sh8Sa+0fWPG/dPmW
SeLE5Lp7tRg2S+5RSxTRrqzFdyNsx+A4GlGGE7dVA96g96pza48qIOVi7YzSkfFVQoI5DDgtEsft
6R8vZjODSAp29NqJsVeDZA0heyKoq6p6K6stwDqOs+bshN6/r8IEQKs2dYst4da2+Oxaihkil0j6
1nJzrc4kOftATumKGO8meCJJnzsHkJGLM8KPPPbZYBdpCV42FIUBkhtbXFPX+nlFmrmhMnZOLFch
LfL3Kq/H9hldHz6eXd0XLsupscawgl2HSBiOe1v2eEoJUk0VTk8SOBZOz6LirWBWphX34PM5Ez+w
iWY+ihm8664dLXzEA5myHTm+3jDG6m5sJxdNV0YPW4netDi8HVPgbX51j6R2xOpcb0HOhcwdac2T
//L62tMC3e6l30Ug4cqIW+qRlmQJyVVQXeMm8KB1hIGlnkEXQBNvl9O85Vx1CfBZ6L01cMArJaFt
oML3DmKZ5GNt92VoBiDEFRYwXv3EtYNEA5JeBK9WPzqaBvSnFyLCs9WMQbYVWZBPFvmh5FITiPyV
XYZbWHNrHiDFHytxr2FfWcuCD2fkYufVRo76kMsgYlycZ47FL1h/fuCmGMEVnyRtFBkgHMyXynqh
41d3t0owEcyDAU1p2cdeB4YJIe4eFo+Mlq5+o+qv98Arhl+xXuxVxryCe0EP/3dwyZgOi2Hn7vbl
LNMAbyKQoU7wh5SeDNKOzvxcM+KSUiZ6x8DLOww75BQa0VDegAe2xUC8MhhF/KasMqdALczYPt2/
wyK6IYxuHOrRhHsY+H0WjuR/sRzp/NYIhM68hKxwWlYC+COqTLmmkqRYtyrbbIHCHiwEPli+vAZx
E8KK34/lWuS+ERq+jCc0tcch6OMcTBX0tSLJBAOJuMjLTMWkE/gmFoytxGbfbnBGYfvRnO6uAEMf
Pd6VYs30QcOgzbZgtHdi4/fROsH2svkNE3xksXFTqLY/dkSm9/H7Xv8ErOYuoHUmVoex48mMGIrT
knR5C0vC30lxGpYQNZx04+Zi/ufoTWG7tPz8hsLX8P2NrxCE78B6GCK2NqxofPPrd7opte2BaDQK
m6MjRI6Zhax8eVqaxQ9YaTKqo5B/Ng46OFYJQ+J7xaMYWtQp1eF+ZHGrq19015nvX6D2HfWcLWSP
MWPD1w6jPetkxZMxp4hnk612Y+Ewl5hpri3Lg2/fDd2XiZR7UlpUhOYuvLDrdCCXmpInWV8B77Bg
EzGaO+/hKUIg5hVUpB9Zwm7W251rzkTE87sJ8w8x5fpERyiKf4VUjSRHfvh3OIHhZRVQIcAFMhoz
o9OKJewn+JLE6/DxyFA70booszrQdgQa1za2a63iUEbrYZ37qk7UkMtIHcEkkG6uyxF9/h4syicG
uQls1slrSgH+D44A7HlMmk2oV1a8K7koKKl4lzrfNO2tAJ21lzX/6hevDP5yXKvEiggaTGGj8S4b
5QdH3K9PN+ocXTVQvLiK5KLW5yXY/0AE3c1RTwUjjd5wXSZ+i8qtTbMSWu8+8QRwKzPAaD7LN53s
s6Id4ZZ/ejCUa78nTbnDhYmxSl/1v4AWCRIdJK7MyKrNuBrPh7EeaWZMSZD7gxWxqrD/t71WEk48
QFkDhSqEWf2g35YympHPPqWoRoFv3bnLmQdBRSJzb9AqctouL8jJhMHNVxcKDbzKwAQ5bN9mrD/S
WkFloj3B5epzJfNe5ZOQ4sXJJWqCR36jwuVf7jwFMKh4FwQJD2AVdfewwb3UQq4ERu+6iQS6470Q
fWm9THJdQQohnqOAYdzSugQW4LaF8lmbqB/+WfT2K6eB+neQ5nsijsMjjxb7GlKMazcKseSep0tU
oNx4mJuudCNZ+TTdKTlg4VNimpnlzM2LMrfoaYyjIjK0sMlX+tacRYYFJyLrXT/wOtxGfETITzxi
QT87NxO5kpdfYA/ikSZ5iDyyfnPjiSOP1fIEvosDkts9FJpjUMcNh0sKDY5R4O1Bn3xGe3E5+J9w
hSZjwSoCklNwI3p49aXmO7aOmGWPUhb0lXFwKdTZ6OAT79PrDt5tTdwMpZRNvpkWiQRUA8Osl+cF
KphAMJk0S4yIPwaArsqJ55ruVUGqNlpjkl7GX0AkKsFSQMyCkXfJhSKWzNMDUQ7IWC+N8YpguVwi
q6YqKG0QvxxwgP97e6LzIKPqDAaVA/nDwARU8oiuUU7sRjc7hyAXSvZ9dDA1oZByPpk8XNoVnOW8
dhAmzfq+OgJeJ8y9wfTiqHG1UN3UivxocZCfspGRLajAuk9urmBzeV6id1lalHAlfGBDY0OuBc7O
nOSSfaWRzsCg5Un9GaB9bK08jfbI/Pn7RdoExcAXpSRgp09Rx2P98oiI0U8BZLxySMvME7R944RK
Irbs4QtRylcrcbcb/uaG/eopd6TpAi8QgnLa09RZ6yqek9ZnEHefoL2cRjKfBY/Ck5ZZPbT5bb7R
3uCUP/skMEvn2GCJBW0jHvWOWl7fowsFWVqtWakkB8zImwHG9VBch94hHskxpXviv+tbaGyQ++ao
ZwstyZ7o1Bi1fkySMj2JYDzWhD7Z/GTnOGvFVhjSN6TmXLla9xD2PadXLIvpXSApXMbG29RwM0ae
FB7vvQbNB0ncdEyEwpYKfSOG/r+pOHvDCK1nP+26Gb6SC8vONN2jHoSMRhvn1s0XgVKNVunmlkaZ
GhwsUqh5Y6kvkZHlkdxtApID124C1Duvas2diwH9XnE6Ow/DYzqZ/QUpZkJvhb18hjgh3xDX88yc
rFqFXkF55Dhjt5dZpQ/w2GKPxleVXz19YCe25LzVnnp1wI2pY6BREJZBQgSo1LPMMIgV+QpOcoW5
xyhk/YOvq5I6PXDnOTTybUh7o58ojlBcY8+qhxp5CfJ1cy2CGQ0NyzHwvyOxJryJnkULGjw0XzWK
XAKKKzMlX1mr434Vo9O9ORiSmZxe5t6cJFsUulaLKWbv9sKsu9yHeh7HSbelWSrI3E0+kRmWo53r
B0Ar/P5fL9+SSxcMnBTQVyubRBMNmmE9rg07rOeHJU0Q181oXlhYXL8oOeEDU48CWVUeQIIBMnDN
N2UUELsCeipgvs1+IRBhNc4XMMjGHuCZTUc77HPfu420GcYmM9DVjf5nGsLH/NQGvparFU3YMmJY
r2Fkut8+mG7WvwKlS5AUpJR1i4dqJHO7EeeGJ5PVcOBqVaHANRd1adKumWPZfkDmOypsmiyd3GeD
9xb7NtCsqKWJAZ1pFg99oIaqysXHu68b/cGf4IIqT0eR4PzQAWt7TXSC1s1NOi8lS64iAs/oZwaC
4qxD2baHUxGod+TBVd35r87TDnY3dNCdoFqunHw3IDhvLFlaevRgHbtW5vm342aDEq2j6BvWPpuq
6JIHCkgbzXrfVAnMevbfxDTBGtPIZPEjqrnzHiQ2DnVh/Zks2ouO5WYnrVLfLr/s3W+Un3SCztLT
33uLM+iyx+VYgvo0MFKugj22w1r5eWgc7SwOWkVFTGCO5Dxk8r3f4iYu/gOhLF2ynLpHBLK6H3CP
coDH4vIlvb48VUxVQYv/rHbBPtqgLCzu7B2avXDGx7FhhxK5VFcyBShlATu4cPVph6vYQ+rL7O/S
Z9Ub/Ld93SODvuvD+q3ydSiqfveqcLRmuPys/skixrZFzngQHtoEIbgC0UJEluzD8eKaEs7au7A1
/ccelKiQHBQk80ALRnz51Dq/NfXaHw3m8iS91N3/mv9xPw7iZ0AsRkHWJbxvPARKrIadMnyJUtyY
ho6OMQ2I88VDHx8ud+RLtjfhUOJJ8B51czZ00xhUQn7aY9x+/zRul5xcfMVYxDZD2vC7VFPE+xar
vMVtiQQcdbH3KeT1Xp2O/m9ShCEvDcLnt1yLKW+UBJ7r3Vd0Namz8EBA5hjUfQfk56MU9XH9Engt
0ir3jPeDLJiu/jKBQ8nbITtUl06DKRrHCDIFlEOzf1yFWTmf8X1TTrsXtfl+l8IHG/W1dwQ8H1u1
L2eduZ2kvJ62yZGWM/YAAqgK1S6ucywVerHkI7lL4pNktGPmBWppucpq7bp5ES3bZj5RZjqgVYKx
IhWw1KvHSwWBeIouixNiNiOTq5PLxNZpiG6ZOuS0usFKJ/0ABTBurOWZf/kW24ZQ9SkTCsTElz+O
M29wrnZdDAQzxd7AwEXIxH/VBXfpyIoXlcL6JYqlai/sswThsCAj4ll6b9+/JRFqQjCHQiEDiEM8
CYfWCQ8utntztCrfqVAtrhxf/3JnWaCPFEkcY6tSGvvMsyX+BVBln3/eXQvANC7v1HSg94XW8vL7
XeOcA+lZP0+8Jt535Scwcflggce2DCysSSM9XR7KsXhqE/inpLxNmCknpTJpTiWj17bkfkBugPW9
BnL5b4nKpTusU1uXr6eLN9wyGQX0zC17kq3SdlzdES6KL9wV6xwEA4thLKPd63PWRp1QDXj/mgpQ
689hTn0ttzHR8M/haDWkscv/1BuGRfx1Gl2xVVvnJ6d5hVL4DO0amwilsbmKOq48ht5HSiHJ3gJZ
fqutve3bm1ENqaDNgvAXaUF7xbsERa3Xu8h6f4VGxvNyK7laVvuJ8d4nEk1cJ1VW5u5ui+k7dqwE
aMwSjpdA305xZq5RpnROqVNIDFnVpfIzatQ7+X0QBK1XY8r2abl4coAF3BcU2bvvgduDQirgQNJW
ixDC2498qWxtS//ODybimaHe1ja3iSK6SXqLl5J4PZCeadapLETW72M/+Eu5OnpX04JSRspSczdS
P/h5g0FFjjPiXULfRO5hfoTVuN/6kuf3L65zpxRix4HMRpKuVD4dlRD0U+Y63yAPD9kwB4/NMxYd
FeFSnUx1Swt9tMX/xZEIYigNPd+ZlGQPNrt6WKsF4b57aORwf6HmaPNPXrftB9vUw70/gv5q8ziA
qcmdV8atYG7F1S0dZBsOXWvcPnhxdhasO3IIhthIGJOHsZ2yt6U7VW7osddKzrbezLBrq4gpi6hd
xz1NafN+zeCJh1JlIYuOp4rAxxnlJlBH3inbtXDBz3yyxrm1WBIvugGPpAmhGtCkKUpA+t/eJT61
1tSZDL0i0UhoWv3lPa5SNG8OR8gAvbHAxC6DwGP8+Dy2+x0X9NUBDMsE0F7FidPyc/PZMzmPM4yD
DqSZB9r8lrj7zcFWUJuB6PqS+xfSeGFkR+Vlnxg35whSD3C6vvv9tnbQD6wC4ZhosuxpDc5t4jQ8
vs/2bVGKo3xayPowKxw1huEsYHBcp6CPzU6PkiI8lf6ee75//M4cnwfHg8gV+8ywbtffI6qdh35h
6WIwrYGmjtQQ/YgyeAKPGQeyEdKdqm9rirGAKNGsF8D1BLeoWQu9HmLqm5ZmxdnAT2cc8MvLi0Dy
MdQVzprfN5lD3JGQgPaHvMJ+F2DEUjx2MfBtmnpNT409RPFRC9QX8X5vQm2JVArHw6oKr6Fk8RSS
BzwBrdB44PWWqF4fv83tWpUBDzpt9IkbqGD9QJcI0ijg2E94BVew3fnNhTDrnHiStnRnqLkyIhJc
Lwht0tTBxhe8hbdwjBVQz2ly3uoJfCzbvVtHakF+8U111OKRNQH69XTaKY0xJQEZOFaUUWcwTwJh
jJWsMNQHgf01k+YD5c6vWRRON8BETNtDYu/JJP0Ca7IV20CEuC0P8dPfQNfXWQCYHRMmefwjFWM9
kvBHegw06qBD35xFRIQ+nV1UHoXyeP/JmIN6T8WsITYvLxWzLXUUdE8MJjGK8OJUmdODi73ch2Px
ihvxW9CiJmgN959i0EYsp9t0Z8Mtn8KjulrUhL9Til3hyMgYZyZcVrNx2sWVbauoCvxyX+C/5eFR
zspt5qdswjj22Mi78FRWAoNhCexCoJkSz0sx3pZdx7j+P7OMIBGyoMkxwLHOt45rIA+tBc5A82N5
GOMPW7QgUWQMlVaffKmCN/oQABxbOxog0qEYmde5FAFD+qPUTFWglXwSZZRuDg9/rISZg1CaPMKi
3+3orrzVgyT3NoeJynLcNF/oM38b9osQoFuZJLiW5ZCTpVkHk28ZwkM138iTYl0mynNk3DNQygn6
ezZS56mWIuxRMX/JOr2AUUUae0+jvyu9ON1M0yIfJKFnNj0+sRhgwo4PJsoVT8H/p2/J1cNxN4j8
YUiP0LIT6ZqvASEoM6y2ac18eaEhWmgW+zToUhW/L59hxcdv5YyCoXijbtjtJ/YwFeeOz6cRVRV1
ZsIyeLl3CncByS6d0G17Ym9F6ZwIrfYtJ0cLCOywYpcZfdcOa4SVRPme+fLt2YAwz22JmQiRSVCq
8Bpc9pd25lE2mex7aKWfreD9WNTo64woy0g7hDprZkNpiaEjKybhDSnRAjlkYlKjlGa0gvnB4sA4
Ui+a6pL9z/rhxjcfhNJyeLPk6esiTOtzlkoRA7FdgQmxuD4oS5m0lLHVdpBS3HxZR8GHZVqF8USP
qY9P7a6VMgDdcPBdtWiO1gsCw56Cbu5f4HY7qE/E6Mq85qhCAMT/3zAcZRKln1pF/NQ+jedwKUHz
JTC7dKlWvyLjfR4FgT9oDGamiwxWU4VSoiT548jTbt+w7lsiaLHgap/QqTm6v5UHxCeczKBpgRjp
8Kz1Ga7YrEtIYKeGJeweFFJVxD95eoEjOF7zxB0OZLMJOQiLsDJd2quNTEJv4NpHZjF724oZb8wo
fPTXJXckBvJLj7BpEkoztCd/Gh92nO7YjyEiNZrUmC0poyHIZEsoQUCNwlHDqTl//2SMuDbtvO8C
7FRmNo4QCOPqpj4B62Ly7fCGOrZVx7BjZOwVmpllXCJ3YQ7Cps0uS54G6/5O5F6esVdkNF3PB5tf
DQfRk5wqic8yauvf7P0sdfbdr/4PU1vkxSK9Q371U30fLbrLdxz7Lk8t3fLETvedkmMR6deDdJGj
pjUhZwzCPl0vJg4Qr6cVc0iGCbDBLgp3cbL3ZRVJ7LaB8SvCWAn244bnpVoHhFrWdp9EAUS0uQuL
dPDcpxYVNnPyYSHN/8pN1kL5MIPps+jMt2aVd+szQvDWBxzMM+/TRAQrEcIaAKzt2T6O47djqGB2
iEUshAHPWltkidTlPKUwBoWHpZBBk5HAVeGd+AB1ckjPdvhROg0zYCIhsixHECXfTIF59KefQRT/
SlIakz0z5PRJ9YRVDC6jA4VX3qmWVHFP3+FlbS4QWq8epxHDh+IbDalgaYu7bVqHYno6mAo50sJR
VQCqBzV8ScJKQePkBlZgsnbdHnhwvlyTw/SGOyhTfITqO9JEGY2JQEGpaSUJh0Li7F15M9KGjFf6
X5fzcMyTlcyJxZj7skgDjzVU7iRFNqFUyy5Bno0uEdbxorXFuAXMR9feXwA/9aHzGo0kuo8+zc3L
lqXLYOdyKEgSlni5NoIPOAkKnDGDASwt9QJWPOrMPxUGVkRsz6vQ0s/z9LNEHe625Tqf65vOKfvr
pAQ4+E67z+E/MPoqtVe82At65tyalmIJNK8lh1d30hdB+9ZO8QfWjklc4fJbiDU8RrFy4kfJeriD
W4/+fgQVVaq/PZUum6tx6JUN+1BvvsYo01QrQ92kevJgJ+yVezmTMDWHj6Bj3pwB2a0s9/An5Zev
j353ruCTYN1VjQv6HzS3f3Fg/TsN/TkVNF/zk5M/P2Xo5TN4ib1wj37saPhA5hNKEAGejWJ43Dt8
HliBdBZOHsaZDVl60S2H3z/uLjfp6+087LlhU3mSs8rc6MzEQdLBhpzqVUow/gZsCGr516tmAZfV
JmCq2xT0F+7fXDO4y7VA2dJ0hJYNW/mErlzYZW7dFti0/MAW0K6p1Vi3g0m7/e5HR6fRL6wCaoeX
u7pzKhLry9Jv+CBW1HKJ3rY4sva/bR17fIb2kcQf7naSMB/UXRmTtfz6CdrCb0aiWvIGWQYmJUvW
6Ppa0HHF2oc3GGR/fvDijEj/bgGSrFNhXOnGsjnEY5lAvJoGls4g+k9rBpWkuF+Fvp6U38Bj18XP
u+oQmz6u6cPI+uMABgEZUcyLH8NDLkhCMrKbNMJcK2r0DuKfTpi645HtgkXhAzopUl4Y6wOlSiBg
6ftLLNxHkpsDE53h58crX3lw3G+5qPwS9FVoYbnPNf6TeEC2HVBsoSWXWewDKzR0ygZWNeGzqupq
UHN0eWQjwocLcu+vvFMEvLpjRxPMRz5g9g913wo/LRWZ/TjrANe9Z1hCzvZQUDekw7kv3f2cpUS1
PZyxCa7amZ4b/66zSWjogdwHHcM45S2ouD4nFqwpLOvL0hEpqESud9qRkIFJjvlRi+e2YGVCFDSl
WbFWJcwFHYSOTT1JaYIl01TGgk4kREXt/hMvYb4YcBd3/zzkl9Up6FuxpXAEdWp6tSx3bcfbE/U+
X2jhAwzAxf5r8LlIgiaPpke5ZbFbAHUAc6O2fEnQCZ/3e/+FE2VSWpFSuoMBEdjCuSrpBwrCykzw
mz3xyd4t8VRvbEc4CLhwiw0H9WYXey7iuuhUNFXKU26AUlubFGMd5g+A1s57POHYKhxGK9E9fVgC
PRM72aDpZsTELSYbJfqDPMhIZ/h4icZOyZEBz9eAoVB4sgR2b2aPY3Uh4GPoEXDdhFUTeoT4aOFO
pD8TFR9A3Y/tDM/SCtdnfO+8Dsv4YahiEXNTpguKyaNAwM76cb2i3yLtSRqDCnFJghVIMyVM72UI
6mXbEw5Ng2fNKv892nt4lQQDhfDPTGdXPBzAa1nygX7n6qQtknyBKrQ+48dXCm6j0BRFykH8GmIo
PkFcivhmntjcDX96nZjwLd5wrrZyEVHNW6OYhmuM7oEgIPh57uasyeFxb7G9qzcZaL4A8QxtfH/x
XNiEFTHOdDWwVJn3NglESooVOb33PVruC9jf6bSVjmX/8s2eYw+M+ahzUFEnIFMVJstauGgcokMy
yxqURhOi3Ov8f/7XtYyzIjni2moaqTGra35Ds1+oLX1Z3V5Xt895EZAoRdwPfgSCBjdJ28u/W0+N
CjUW3GBZJflJOA2TPWuhVYoXDxhnCmshNrzbKhz3z0oSmrRaYOqV0yQVC3CIGIDOiAv06UkU9utf
aXS3CBrOD4p/x3fLKsZ6TqxKOfLxdnWlzcPltITb7jr9ls+YqhW4Xj4W0bRdY1qp0aUghqOXG8JB
WkD83T0j6/ZPo360EUiE6fbCAZJZsMV5/IcqaygwnIK5MDDM9T5A4ADaN/G30fxhXXTr8HHwqQ90
xRr4we9XsaajhRRh/Ia2wx5TfmkWdRJW6YV2+lFKnYxkHtn0UmFbI3FYrT7XlDVF12YWgoXEOTsr
qpfnfVUD/wpB1irhg0W4tfmTgxeFLTwSCywKn0CKGpLoViLOAmXwCncwd79rb01x1SMSVFgZab2O
sEClj42geXGaoJySiJ/ef8YlQuvQni6Wl7liOszuuCWU3ig0flZhHUN9A3bk9Zh6TS8ARWQPz/fi
ULhaO/ZlexMQrO0PUpHnfu47p8yn9scRlqbqLDUyxjdvlWnaO94DnmL+jKqRqEnL17j+sM+r5SEG
L/UtO9tS8Dd3OwSTG9usBwSU4RDRzOqTlbfnG6NYeM0mqPo7jWVX5xIwDAXTCPUl5yKdja8WTY4J
G2dAKhd8OSy5zDPKV8rCAPNw27uGFqB+lNIH/QVJHTDXGOMjCVUYz76LuiHjbb4+yT+pLTX+Y/aK
1EanAPvPitA3UZjZF0y7W+ZnqtcvmtcP89ljqQNerCgfmfODW+jzog+e2JJ7tu7Hebi2XXI76XgJ
/X7/ECPfnkAOrW1zoBaOT3bhs5KF2UmbHAsbw9QfdwDmyVPgahjOUHVLKzYb4IbcXB2VI3boGhls
nPQKy17s8dOPtEmdlUw7aA0Y7bGv20h1jQ2SQncBJ7QmpZevVya5O+2+9nM2G16HDuRyqzIrEEFi
IVgQQZz6/ApbVGoGHyn0tPYhRM/8DXQ/wa0eQCvHZh/GPDB/hTDhgPxtLsa3z1sF7WBWAT9z9Zj/
vTiBTLNP0w3xqTda0GBt+4mxvDC/JSnuylMlVs85RbxaExn+1KYBSDKl+v/uP+vMi/iC4oaJJZRb
XuglUIr75HPoaPLPoTTn/FUi0OSxwZecEICGLKz04n9hBMv5hcg/20//6i0Sptx0JhVt9OqJlOki
gzdv757NhNox1KWHAcmu1Lwm/fuHHXjJ6ziEExa7CCiDBz4MKgLyI+F0w4zZqzBReJAI/sllBqc7
05lQ6C33bSR8BjMgIS1yRsWYM6CXlFEKJxVCEl3NNubDGsooOp5fu/ThD2dBPBzEkqD7W9sKa00g
GRrL0leYk0wTrx5rwFSwsytR0VMi6MXj0kL6ngD1ar4Br2dkDn2EvGlcKSlFGR6TMptzakc4D97q
MV6HjVsuMnUu0FqhQBM9JLo1KdeYEGd/J85JMSA8ZJPSsU2WHkSlRbtCbEoEvhixUyBEJ1RHPXBc
SOpifClPl0Q1Ci9kO5HVoo0hHxfYf8qF/FJqgV/CLQFUCKpzwRZg2Ku9Ngf8Zf6RlZE7wJfbr+z2
ncWuZ/5RhLrl7Ls829Nf2Ukgw/QuQAkOvyMfYjSjfGF+UwZL1A0/zRsqNu/HsHmoEMfkkkk+4OOw
2Qqurwj26z7YzTivDn9PnvLrM4L48QMA1l4BRZkcSrhXQSZvFYF5VCtier7nuTiYffP76ta3GGAx
3EWBm48k4ZBCXm2q9VS4QLtVVAUq5Fik+D1b8IdZ5w/bZ6YTqkFaZZyOrb+Id3bIvysCPKucm81R
cN+OY6jHEJXNMaivcF0S1Sq9HrR9IQ8mO2qMhpaEFmWqj0IXAVRwlPmm1c70NgfpFZzuGvj9svZz
PC4aQd2VsaH6J7uevHXuZby5wS5Uj7wTETv0rwNyH2Ok8MgSS8HjAr2xJT4Y3e7xqkeF3ROp8f8T
PGiMngyMMwmmW5wDIweFM12FseZPeuIg2m3P6brGZRU1Jn2eP6zWiguRzhZeAbYG0PuIqgQLEneC
QP88X/PZYP+Y8nAjZnpfIH41rxmI2pTiTMZinpDXbFzBU4Gf/WCPdMVuc/ZBYo7DVEN+2Jzu1kBZ
YtIfRrqal6WP6eSJlUT3M86o4CmoeNa9TAGIc8p1uugH/ZEJibOzfD+z0iKebfs1ASBwZLz6445Q
S4OVcFTqfyuOx3wfoB4WoUgZb030+85fCUIbWofz3XHnFAsC53xmKdZqYK2o2/SYBdqY+HVkDLbz
uViIN36soasPnqsiDChmETX/QdTB7Pq5LoTgWvg+Uf4UvJkIR2YhdDeijYhV55vemNtrMjJZd+jT
aHAGZXqAdHiMZrmfcB7xBgCrDeSYe86EHmn5JpOqtD35Uh9cO19s5Pu+0IziUuJ9TWnxt3CbWywj
Y3ud7wUXMYX3MoKMS+CWzILJ2oshc6mh2ipiqhRjtbbEKjx5940hgqFvzdp0pfjwVCQBEivRSO4L
cgUWgm/nfzsyA8HjWPLS4J0Mx6kbEoEKXD1gq9sWNaf/cZ8IxbZQT/5ytw6GQjJKnEyOL5vd3B+5
Zl32Di/J7Olm6OsnOTOBno5+mYVUd44a7pTQXTrvkjMw2TLRF0b2IQRmuQKT5MzXsd5OFfT2lPq4
e+4AjKRzFezTnT5+AQmE0b9qWFZxkB1esXVfVW1qzlp7m8nGS7PcLls+CXLWOwlFniDLpKDndQi1
OgC7lfWqOMSm7mck5+bEGG/RFfYIubsR8rFtH6NcyFhM5G74mfUuL/Ble5mkag5nU3WT4w7MX80M
TwfREW2/+tVW5ZNlmZh4TIrK5RnIwGxZUZ62iBPTDjqDNKXSmJb/a1WTBxFdZCa0MBchUGjBKHuU
tTVYIubKyLO5xeGjc6oQ07ufVe3Eg69QS6mqYa1Hmg7/YbzwnuSaItHcQaovLGlrW9Ga+dSNxi3o
LxRbo7s6PYD5Ccm40QZlHQcuJVrUggQpnqK6bkK9LN7xTriQUVYuRa54JUFn5tgTQH0EHsbMtW2d
/GpyuL8JmOR2Cy+EWsyOMAUc+KcNRkNAqnIg/vW8BTykHXtO2zssk4KfuM9httOO2tdmaBhrEfpw
uia7ZKQ5I+4LgKbvW7WnMB0s7jPwRcVh8h5OsmpYbrCoeka1rLwH2SE595heyaF8v7fj8agn4+N6
FBuTjgH/eAUK6qZ0Fz53k5w1ysHIp3Xp36pMKDRVhwMKuPZmWvS9Yz7EjkHJHeavlBiZMB20TYDB
b4J7Dqr4u7EcD3hahdmQYpBpSi0wx9q8Nn9yjbU0bMWwp0F+MdV7TK/NTJNcUXlHKFhUYEdeTRtW
s1BXFzmKquIYNsG/50rZUI22SUKLRAL3DKpyrvS5svPEWU0hUIQ1vukQPqcxLzkVU5lZxmwzsZXo
wdlaM4SXzOa5ThFpGmoi8icSrF2NrQOyuOtZHcbmpt9C7iiEginHgqIxhieILQovPDPpOfe0huNs
1s0nJXIfg6RTNQHvB9ryFigY8gqaOcpLpctFJt8MyjWbA0en1+4oybSVOKCFacIc8IUrHBTfCBfR
enMzXvQs5DtrrywTqLUcPJM/5kOmYRvSym9qX+lJSg9817nixPxPWEaHBeiVwqATqXZfeK23GUC9
CbqHtCYW9oqXXidTCPWTbfQOJ112f7lxCbSTvRk0JuozwSxdfP+kLzss75JhZYuLLiy0t02wD9qf
c11chjuIijzCAwBbfx6YhDTAhq3u4VQXBdtZTUtpGarKxbX6voGNOb7OMNe77Q98j5gy+NpodGpF
z2aJjNQqaSXDCWGk4jurAWUjsQOgjn9N0aDTnZTdBmUEH7lNCJ5eb4dWiomFPRJjIrwupqwgt9Sj
2SI+2GD4065Tf4EvzPuxQAVJ/QqGH9hiE1oe4ul1M76mquOP/QKt+CHYxwP/J+WkvvblLvapuDbA
scgzaGM8wnXWSqywDd+va/K+QCOo12Cjjp3RxFV4TYLKGL8UiAJd2hmz7nxTqQWC0snNlA5dHTLz
X1bmb3mzE1/t/FV+tJu9BF0Xp9lxPeGKXSvpLCttChNSEp08rg0/QLSO6XEKHHbNbI1czJFz1TRC
CVcRuQrmnEppkifZj/KlOcfJTAQFPAHG9cRmtoZYdUbN2lXsQKzY3FUyUpgFiPI4OpSPxVYreQRW
czhhGWzE3G9ZHTOdJEhZiHOiwvNSiYPvLgF1EeIfjX2s7CVfr6//O5YGSVwA531pYlm4cqsTLEs/
HR55nwYLG56w70yEFl+w/FgZoM9TTVybmDLF5xSCsqEzrQGG4Gv3/LKygNn691VPLFZ9oMwxt+H2
hnPuvttQdYIl/MwkRfBKQB0KdgButokQhZ5C4gLq/D3OOxfY1YKXHWlAIeCELJyk2lUDETc81UNB
62MEJmjhLgG6jSOpTQi39Pw/RIRGNU3yYSCoJHn5myfIk/qFa8uWc9GaNAucOO0b9oq2++B8VhFz
PilSd0spxb5eTetdmNK8MC00MI7SYVc/FLwSx/Qk92zevDs8tNPe0IiBkZQtpJiPhb+uS0ngiXKv
UhGP/0P6KbFSPJ1a7sH2X9q0E3hcxZVQIAc+zQxDF4GqySu3VUkxuHV25Znb11cuJH4IdHlazebX
kHHjhn1TT8lV6NrWCwtNBcjTf6AOobwCmJSIR4GalxW3hrt99uBELh7x8GNTzVJ/Qc6GRq3c7mUN
BZhYoh2tiU1V1rNXMG/M7SfHcf13cnM4ud+jcTJcrTaE2D+nVsAGEPjUS4UQgS3eiqaJkMYChUIA
TZgArjhM/w6MghIO8a7nGVLYii7oe4FeqgkOskAS72eCb1+HcHaRRY9zeDnQ94P+wc6MkOcpYIfL
+WrYPeJ3Jrqim2ABs2Oj5/kpEmOAX5an6wuyJFNBbguOwFMJXidWJ7QSKjS6JNwv1jYqtIQeiV15
9ZIHo2SMXD0WFRL8MMOX8UGRCIaEH8pORXIF336v5SF+BAHYohathiGswEwJOjWdCmqDAPRaovTx
mzC2t0fm+o2PFSg8h/scKmMkNjAlpakkeX0lVd1K5t8WqPLhQYKDkOiVw5vr2Fdeh4fRG2BHRm65
FE8URsk9mrdRmMvxXpm2+ieru/6DOex1h1SRBW5qb1UozRQGop8Wn9xceilPcA8neVR3KygeZIZ3
nEHcxZqwvMGVRc9UQAMmvTBlZ+hJGmqz7PvqUZreLH77cXdQcq/qjTUqxFmM9SUKVe0lxlmwXer6
L33/OEvvybvqF1G68j+RZKfqGHpNKnrnQ0jw4k3euPWwpMAPp70ZsU+OA/mGujVca543XMS1rx8f
EVYmDsRwErc1FIAXAPJtFx/guvyr9Y8YKirUfoQ4xbL7KWfToi3ufkyhKMV8CvQO7BFMed2COWLs
1iVrEwObKXIDDtXQIQajvQB2+zLegWGKpSDDI2WjmNhlADRLQ8N7XXGnHe+KMsWnrdc4MQqQuWwY
lizg5jVcJwyl2LiCkFqifdZ1Y6yRPg/Sk7d2kimAPmyTo6mrx3xSxPecIbPxVed2RRALDjkgj7c3
px2J1WnTiyV+sGARgqalfpmO6piJVbVHdvkpsX6Y2e1/FuGDtTYGmJ25M+djnizjY47McER3saQ1
wpvm2/hXOXCV1/J3keJz9P+BJYEBj47Bm5RfDICNfTiApgZxhXWtJDKqPUrBM+mAgsBZ26taFSZs
hDclVubi9Od5GnJXOELswPWCifMzR/MRi2wcgQYtGMHX9Hv7nMttmMYWaF8y0Zv9tVHCoF3vSlUL
veIFIGNrMyWLu1CaPpxIu9qZOi5pdlc9BpTK4At5Pas16pOA7Pn6KAlzhFG/tl1mHt1ugQVuGawf
YxG/K20ST+muMj3cLgJKqhimGmQCCDENy5onR5mMv3GOF9QZgjpUPn1PHjtV1GUqUaba6BgXRme8
LFyTajP1n1XLllqzW8iSQvQY1TUCMJOjjk/GONX9D6XwWg+6KLL7cE74uVqWvyKU/lQcjNgGeQbt
I24iEHYLMg1A//AKmIwyljqIPjr3M15URuQgJJGBscd5uKLsOmqi+s/J8cY5sjIAJD4lDYhSROBF
CO1ZCaYxy+6wxqIuSfJbJnGJnMJw+b7cg0WCCyd/iK/SGjtmnlwvVpt9E7NKTTn/E78N2jpHL7j9
1oN8b1QUCIblGSpZ1se2z2KrbBj6WBJflxuiWB1ZKBxO01s6XzU7QL3uAfUR5U25wKDfEx2RQBrE
W63N28zmaGPOgn/lfRyKrgQ8JGWXzE1tgaYobuLRw5bdxksMeQ2pVP7r4aXfZoVutVNsSCKUyc6v
L1Di0eeyhs9rs2oppjEVJ+CNPnH1L3+RCrzfORZPBhS2w+qjhQlvyMy6gIFAJZDVlTIHuSpUmevy
etx5u/l+14/6WtoBoXaGGX8MDRMuq9oDFDMq7JuGDzBo6zPadhECFBEZU/Hq+gmhQqlEE/3A4c5Z
JVXmcCzgqIoCW6Wa5hi6f9XBareD6STOLIwAweC9YeWW4jQfVZuMae/Mvb2Fbww5sUnz76qXGijW
6StF27NBG7KoYm/VEzbK2N6ZajRQWpxgTFdI9qRv5lWmgKDQmmU3w4RNXPKLmOMc/br7z0snJcvl
pLfMhzYuZ3c529sMvnsXIlWMcp2Qdv0Q5X0N1VKU2ZnaR8zvIUq3zFzzHNFRwYlYamx3gKWWgvVG
DlQCMeloU6WCC8uUAN/yVxkwZh4X5+pwBRONcHkMnChJ7ahtGpZ9k0wNbbxJqIhn/1RQQed5BNKV
wTaPzCQthtJuQYmLOi0OjGAkLNvd6R4V8RTFJa6quUo0xxt3JdEprMdPeQ+i8JuvpIUr4S3zRpSj
AaFHeCi+eGmH5KiRtUXBQYIllQjUOYou+3AzEbRfn+KRX6FkMo7nSFgPxk92VER2k51BhftMJzuO
tgfr9BSuvHWip5qBz04lDK/ECX7lNO1eR+dDhiDELf6xn24cWIwBEyFFFHI1TAHCIIRzQe7JeiN/
ugTzWrk9LHjwMonLJpPhKV3i+P+2YcxFKlXWz6n0jyMrFoRC8m48MYp76birMP0jUmIUffy8U+Q2
kNFK0uAPA0GAF9nRgCi+Oj8lUVsjFXvahZKybLYDbr0JS3UfVlrHs6hSp1RMKBSNoQWqt601R/MO
LlYlfUctTWugsXXfJcQwn2et1KVnrgbuyV99OFugBpCcmeJkV2MAEPWthgsEpMFAJm4WYM2sg4E8
2IByVtkJ+zJxar3+EdMbUkdRU14UFm4vaYgvaBXibqnxql8ewPye84mDGNeOCsG1VzYLGl8q+JIh
1xN3Zpd/iZZLwmaZ4ogWe4ap3RoomZQglbZDDXbVN1Hh/2i3iRI/29tX5azQMWZ7BegQJn4LumSw
+/8Gt+cRB6tLyE5L2POWiNxkQPYKYqf9d95bakktkauRMyDx2V/5hQWnIS4XGTEA5+rYA9QTzB4l
OlNXGSnivFDaoij3Ug4X4Fk1wPGILZhlPweFmBYcDR1Fhi+d5BDkOeyAQ/tFXIis7N/87mcka0u/
X02kLf30WqB8tjWpsEjt2KSR+EbBzMEbbysV/GpK8J7bfL4b6/mGM+6HIFuuig0T2uaI8u7d2O0+
vRvOOxTVQqrosIwh3Mfz+eU0j5g8QusTFKbeaR3HidVZcaZA2kyPiUWImwycO+/1fVIIHPKCHb5Z
VHXldpSE+VCwfutjg72cQ1sH+SyuhF1eJssvgA23NADDaIsVcYaZFHcC7a11SAY0L4NMHASYyRQo
7x79nPuPFfFTYEB2M/4J5D3whtRmADnIUvjUQ64x1bIsvBYM2CanZGLQaCL9wA+39Z+UW4I60zWH
dunaJmj8t/0xNv4IfU54hdigkSJ8cL1Q2iozaZNWx42b/wMWiU2sRN1MicGwFMiBUBT2sNR6aXJs
QIXkn8zIQy2HOCDU5Nu6kS9pt7SB3HKXb3NLLl6i7TsRqvx3UWnxiuC8fNX2lTGQDd+4d8YlcMOD
PXGDauB5B4QostctpOcTjPEj7Psee/R28jajLFiLht2lPW4ZHx0SEXEcX31qgNK8s4blS3vfm8Zv
YSm1o+uPN/x14ubVu3lrEvnPl1mjNUL0z8ryZ2Dt+76yCPSTlMgQm3s7BxJsQhJBJm4YIZmnUI1N
s8/jSdeR4JhmZNVksWuWWJgaiCwb3qcKfBuNP1rZEbl5vIM7RVJbj0tbfdCU+mcRD3eUKZhs3fw1
QcbuUaSz/dcP75/WTfX2hIah+U4OyVqH3+ssFTOMv8XoBI0FlCX2ZfwTxYnvovAa933KzC1fDJDz
HLVxwSkBmTnuvDqCbyO6441LNVfzZHSBGcTxzcYU4GgI/67VUu1HEZ5AXSarPPwBwXLdaiYldGpX
XzNzV30eO2+YBfuO0JzaDbac6e4K88WXq0v0j9naezOshPookTexcYIYYwOJDwyIgvPdJBf8PyOa
89vhEB7OuBjPzshBxk4l/j0mpgl6YOygSrlvktVpO7ny19dpKoX53ip21ghEnpXxYOBMbX2foYp3
LCSj2Vfke1ail/XJVyZbDv7MxEs6NnSHlzpe/XsBzEePDXuz7WG7TSnXOwxX//0mvl/SefkHLdRt
58WJ96jem35gNL51HX2LwBfNloRgD9U7d7RMqgvsyo3qIEWqDIWOdyGuwdq5LNOpIBUhZSTSCv89
MERaBZoCxTBulXL94XcxFrokbBPW7Ou4pbBKIus2cJElbHjABDDX3EIuY+f+lKgTglVunvPzi/oZ
BA55tr5i7ssyARL18KWPT4tfSNHhYLQN4cuzs5rYO0y+MO4jowcOoLn37yZ35Y+R7RT4OqIqX3sA
Ess4vtkDzB1fwyuKyouH9jCYvlKColNOSKHqvmp4nCpWxA8NJ5gFeRFDsCNqk7wJL+r0b+YhOewC
fqTaDLoY7th3xD3H/tBoBRJnKsgejGw8eIx6XJl88j9Rud8psAx4eNTYT0XDTRflcBzUZ5zWtxd8
IlnooGx1wd6l+HAe40XJOSu2oNrySNA3UM+pvY7n8LO3g1aWVu4psG3WN5nFNVR0L9WNsn5+N6JY
r3X4z/xr/iWHkNHBzCW3fNgEnjVuoUM8dTONWkAKeCObKPbXcsiEIPpLRnufN4BM8BERufBNVH6V
SpxStIQIkfyPJurTuRhtzU9/I3StLd0+idcICYLg/PhyqlMfSuFGg5QNy+jKdzpbtn+buGfcU2BV
Ri2MRN25g05c/dYgimlFTxzrBlqihOaMS64M8HNdyaUv/IcTtsooocJm04RY8+B45wYgTG0apPBG
QT8h532hIciyUVccXdd9pNUuTrnhOIC5rvSTxltv6bnB/LPN/RQkhFMemq5WQKaSQsW03fQJb5nd
/eAVa3WU63LYpcVpSdOqUWiPAZA6uyM2L6rNAZADmNTTmuJViwi+qwxEpzZXuGTANG5ppYsaVJga
mj0j0G534zwSc7ogFOqkYzhqQ0iAPbZuQjZ233r/50MRI9KhV9b3UKxOFKVQcZQf2vP7tXdSTKKR
JHgT0a+vb5tY9NkE8NcKmbklwcurmW6bSf48OnJDqU45wLme643x+RWrF29IfTCAHsTGgFF2cLBx
4fN5vE0RNrA+Ahbn30YgN4KqeXcibACo4EAQgHI5cGYj68kj+cariv9W/v8i1dFvk7QSzfmdsp9p
M8CWNzkBXdK8FCUsmagcpQgD+ZwYkHWW42YNe744NOqP9Hh0byk4PdEGoYYp97eGmVaQ2kuai0JT
+bo8vtKw4xFi42rW/a1ibZZSxB9GIFEQhPgo/8SjgltKtj9v0+cZrcfuiiYJSl117zneLZo2b2R8
UBQF3ksl8sG4qq2ZCmGTuo7AI4aelBMzOJ/EaXPukcFjEc6J5ad3QsWoiQMRX6IZPtdYBgmk3dbx
jzuyv6+bjeehCIcbHlFi8ew6kbIjOgbLiy9LDTFayT6aYRgkPQK/2yJoYERNpO62wB5KyRVZRBvf
LZOi1pdvIR8RZji+HGVDkb/ycv9S/DnpCQLu7Dd6nL5twkK+U0g1o2sh88mqDGnEf8WwO0VCQG8+
gb6kTmILGTMztpdXGo9d1v+wkc7S5J8fiRnIWlvVQvr3uK+25yWpW4fBdUZlTjIwYO4XG/moYBF2
iNERVg0OwOVAZ4oVTGglJp5a4j8QX1fwM+z6NNK/YoYMHqzaOxPK+2GagNq12PGzBGrt/2S+qVw8
c9FrfP5uBuFh/uQRYgfy7zxZXupzvsCF1o4Z92mNcSoarzBq9MWTaIfQCleBNms0d16RNjQ5HGsz
GNE3SoSSg6QHQNxpEQO8IMH4I39pteSw7xZD2/d1Up5O7UgKgwyiiQH+3VpV+ao6+NALcEfjAF70
v1bi2ThzzI/u8GNybwSRSLNznucL1rQ0qsp3pxuAGil3EP7EW5Be4otX3uvfb2ADi87KyApw0HxM
XXF6E3r2/m+LT95yGqPN7p1K85730HinbX4NPqH8Vt5Hhv5heaENpNmlEVYrJXKeG5oD73ZWmdMu
AV7XQcsP4CXBk5MdORimm4zrHerPoCcre23INt5DrmNwsnn6j/t3tpUeEJT2io89MCiKyWa0dvNL
lkw5BpSysbAzCH+/pijq/1tTRcNyn8RZMdZP3i4IWsqdIlshKCnrlAHSNJ1gwrKzY2sKXZbwMBt+
so9Bmfmbr2yqz68UiYh0jRdCNC8ZrNg7IoBpCkM5pSf7CSspN8J8+RTmoIcbDno3LKwH3xWjo9T4
iL5Qx++VdfuayIPpCJ/2/lSXrpMTMRvrbFRHkCeQOYTC96tqpeWlLEOJimn7m5l9Uy4x7IYtjPql
BCmO/FZkLhEkeaK5GqxK2b+AGTIbw7w9Z1JYHZwETfroR54F5euMcwVMEJDUNEmW/TUdL3daOoNU
qXvG/JnEiZwG8adFy+foJF5CteWeLFhgs0H3HZC4ajMqnaoLAMt3ri0dmwqgVQ8Dcouwld9+aPSW
/ogfigG/B8NdzXIQkq7zb1dIVveFwfMMhKSoUyuc4jxNvylECKCadmFOvAdlUuIyjFUc8wuRFXQo
r/+fi/4aflZD8T4NRgpqlzwluO7BiTyGd0bAm1kuJjO3tZ/+Hwsr2cLRsjfaezkICkf9mw/BSKLi
4cP/PSuid22RsAJIFzDlprB87o55F9+SACNcCb3RVjPxzJG9wXmn33EVdm+0UhT+MuRlG7DX1ule
6PWkNLVl+cznkFBxQwQCSF+6ZjMXcjAnXc94c/ZeqC7V+qyrl6hiLHn0bEV1PvQVhTb1/C2csKMZ
vGu7XMOTPvX3jHJlXFsAfJCFTvgDPs9a1wc8bzdKREt1uVUxMYNXeKAhLIBDT6gJ+S23IbCeK/g3
urb81ubqntsgPhTsIAeTti50Ff7f+XRonabYdrB4MY30TZc1TK0qrhlOsuG/0Uhxy9xVRR5u5YeN
kUKqE8OJShmyWOxJ1HeWnenXh1r3xnx1XMtta/y+BmYrMY6jMlSq1n7EiuB8Fafgv5w1+SqVlVVv
2F+b5cr+/ttr7HpVn5bVZ3yyKlxinqzm7EJ0pfWCJ1BCeQJSReTS8Zuh9uE2Hi+eMKf/UUAtNAaL
HVMQTgX9RavlEdcwigMJDn+z8Qx1rYINmnl6+Jxl7PcA8WzgpNtdHN1+9d7GGH2LTq97Q7CdFWXC
KTHlsAaPaV14xnAneT16sNRGGi88tphoqtC2EQkTWtBkHie4oEf9evTmMnlUwWk6Rd4BntrAS3xe
SUjGQHj+Ec0iAafNGD64R4rRVHw+YsLUcOVj5FKzBugkEWtzeZVXsevYZIgnMc0GgRU5g8iIN6Uo
ygukf4X6RTZnNDboYNtQ0z2/wvaKpzfLQYyCIpRUf3Q8gSl6a98Nm/RGM5pPHq2fKIA6AoD9F5Eq
GrZeb4xi9guKsoTo3qRXyOuSfj47G7E21RAFnS1NGy2wktfH7A3PDnDQO7E7HBfVpanJcxXqHOzD
sAn1tpVGMQgQ3iOH/hVWnF8C7JSyXub4YkOYbp9EjPxj8bwP5sPZpFp+prBHyKxAm6Yq5c1Vtzus
uqOKX0bhoYtvN309rePA0zWphUAkZBtOteVLVg+d5xB+OoJeiE1TtO6HBQMGtaoD3kdFGFAP2Abb
PQJxyKaplm2t2nsaYWI/8bQotIYsNdW6zJcupHRgyOXkbJlNNxww8NXuOYJOsyUUwUqdmwDTFLNW
GZnXtg0xhalpa+qRdbQvXc1rnhq4VL6dB/4nzCpDUlrqGr0WXgFRwInpgh8kUuYUZc2OeN+/mNge
aVGlLCngrxDnyxEeYkNUtyfW7Xvlwu1XHzWyC7Ufpjgjz/ZG+emXOvyTeBrTfY9rBgZ0VfSPB4A5
j3mbZ2j0R/ROulU4klwq8BxMO8OeukghoXQgY8VctrH7cQ5YGuO4KXCS5f0DpqxgvEeZ74dCevVe
Kn/SCJC+lPDdttYNW1fj6lT/VYhhQKUqHd7movu6CIoFlhy36kE8jhcL4TxspAGKVql43L8i7yXc
k/Qe75qb0BobQpCGQsimH7qdLMGf4YDlOF3cHBIVZK4zNysG/lKVZOXvTIUpwSjI9gmQr0jIudTR
+D9OknfbIYBEOxcjvpGkF/RBCaDUhB+BKHPL2juGN/mLOGpOuIKndyJ0YE6Qk3xZk7qDmsl1SU+I
AG90kyoff1Fz70f2vY+T3i/uUoJ3R6uapg1c0HqXN950uf/FmmcjVLNZ9EYHETADY2B8d9b5sFJW
yL7RYI+J/2SLkso5k5xZ2djA1BQsCxi60wMqoQhUTqkBzHj3/L9L2HsUeZPO6qdmSiTkGufJHaFk
5VLN0wDnWTx9N/kE8ITHvQhcOzLRofveRAQBVNnxHsdhgAQ+SvYln6it+S4aSTADrICDRELDgSmJ
otXFb+ggMxeGzzMUc+UnzRJY52N25dC7WGMOJiLqrrbytLYPCxs5GV3l2Uw5jZpV7NHXTOUC1T2O
pC7M9gSQWDXhyDznzrmIZUUk4vtsT11UzWc6/9eIQwyfJlSqilL21ZZJaDoTNiGoFWL2eNc/qfpL
SMtRqZF4W8lW8912eVg0GwYUwqKnGrZMnZyWwvLV2guBJvWUFDVn4ImP7oVSrtmfOZrGyBWZOYkw
07aA+KAZ8+38vABuKblT0I27pWzF2YMaIWJhnW2cdT6TlyykRfHHyVx9RL4IM7ZnE197qiFvSk6B
JxFLaasKR97RVFT2ZppMURX7JjorRh51ncs/6JiBppn5niIjjoqCjM6ZLsLoH2bcy+aqD3G5in75
JaRKs3+b4j8shqB0UdCeEm/g/y9l+6LvcMBqw7cXPAzP1gHY1nfJt1qEKe3bQDJn7bisBc3BXJwm
y+qdgk0YcGQByF5fJ6dIcg9R9b0funAA+slfYwJNWGoLgUvTZ8/CKFMp8NtERUjUBR+ltMov9vjw
mnYQfR0XD6hVg8gYEHxHskZVwarA4mcGhCdWaUDCl4kX0+qufBGBZvM68kp5W2T1AVkjTB1+mmBH
c8jd9Km87gEqWTAtQVN9I5X7tLmgCumf1u05qv4X2TQwg8snz4VHNeA4B7dvi4S2cg88qtup/ka1
3VSTWwfgqQn8alRwg4lS4BGEyRRlCzArKRG3SkHztb2zonVXDXpVAZ3z8GtGLjo4olQ7RS4TL0YN
+YzzayfQMWUA1vZ1D8Qb4ngAdTFRhcBFduidRRRCpNSnjWAo67dGbooa/Tg8EwrJv8nZ7KS6Sm3D
rZ1/UuUhf7pfWa12xXxS+68rM18olPkuEylaL0+bbMoNtwPywEeOEHP5BnNSt7iODVUBxn1wTn+s
rvYYscDt3ZF2j4ThX/NK8QgOcEYkSGTiURzb6ctrS//50Xaj5ivdZXM7qbQk/e7FjU0T9ejvFr8x
RLpLswbK/lFp2tvtBlR13ZK49J+SiobKHfuZTHZGJmsCYDkx/nSigz6O85wZART/12jgd+rQBYKV
1rvm9fS+Fsj38UtU4xraUUbs16URtdp1VyhQ0l2Y80nVo+bGBfmPLF6sNVgASic/jAhDXtxOofmy
6UulB9orW9d5GEgQLVWXea/HTmLQj6GYfFfl1hQKl1SsJfzBz0exNBAU+gAVHF4odH3QFhckuJ3s
fh7O12vh9VAeSWJiVWnExZT0IkHZywfWKZzfJRHypxTrds9aY4FwmQfgASqp1HngpGhIEmnGWJ9Y
eqtDhRRnAr79tF0dJnQ4gPbbdPsNawKqVhHUL0Wmvm+i9aaVwzG70jdEew+SG62Z8OGrpyB8SF8q
uQ4la6DBKXgYrPY1fLl38mlf3x/1xSoNFq607bT5o9R4lNFQRfrpKOuprTtwfAsPLeHCQMTXMTLq
AzQAlvqcqzsOOQ/ycTTXCazDF6LO9PklrkdeD6gjUARzHUNGqxvkg64JI12MsgBte5vY3aRXbWzV
tcs+9wgAU2ifKHWA2HlOr/fSEkgFaMVgGAIW0gBYuS3N/KOplXLyJhsU9mJ0tt6UmH/sRfpIzW4D
+RcbRroEId5bGqdIKpt2UgsR4g59pd/JdoBIBUWg8FCHEw9pZc/NhRVP9Ew848tZcatdLQiw1RH0
a0FIu09Lkv/m5vRt3U8YcIiD6k80ac0Wqw8Nnp9nbA2O3miDzukWNkVlt4qsxHwf91/JcbD/6htQ
8E77Pm6Q5rdw5zjQQIpUsZEo1Qs5iuotf/UX08N/aIzekMfkLrBkOCs21rfQozbMvuB7VQZIwEL9
SFiSTWu84ujB9GK5QwkwqO30nccOjJ0mpRbXwXpgUv5SwTGGkpqOqwAH6nE520FpHQsG3PF+3z/V
i9nOb2e9BkYZLInBScK+wuGphqciGTKrDr8Pfy/jGYE2Y/T1INh48GZiQTBSHZIUvFi5oagcAsrD
UT2jA88v4mfw2if7grlRnb53pmOuPf5HZ2hG/vgmBTwqlRZd/oUDNgzDs1RQ6h+8xFc52iozfkcC
29hQ9xns5DVCKMhDTZOZL4tAv7auAb7v+x3AW/jxVQSW8vJZpdBPvDOTSqmo5LNJB5cCcUY8zi/1
kz2Z0Cod1bpL9XC7P3x1Tc5Qfprp/BRDOn0B9AOXCKyHIYKbOmA4QCkL+OPhoWcX+kcr2h59BmkM
3Mo0oBGDjRmyW52MiOoIDB99ehkZR+rm463CIVqd0BZeV1nY9v6brn28mZJJL3GHRYZy+p6WAppH
x22c7IGcpTbMJj3G6oyLOXCenvfSyFRqE2o7JTFWykmgHv0s22t66qZIjKs90NVvYztva6QP+cdG
UpVoaPMe6ElfV+ru56iIZlW0khH7ctVXGQywe+Y6fQszF7NrrplVHVTakwB4tJeNoPSGoY6wjOmt
SzKv0sEPe3d2GUvnfnYNmmQRpA024scDTQSLlJHXNUGoA1dAyvywk4QV39pNvQ92RQ5R2y7p8QLL
1f8eh9YNAjP6mkkMwgf1mwLOuo8Vj+jmw6s+bBC63zl9mRM1XR3ilgBo02g1rgjuxx8iGmUPRxFi
LKWYO3MCv7C6RkEwtY2ROPLKzDneQXhuMhzHAfdDhtcs8KIUc92gZv2lvpRY7pKQ9rvqLlWdz4YT
r4Q4dalHhF8d8Q6b6w+kwHy6xc8JKzUNXM9C1PuKUiTneLjIpKtopYQ20XdsSZMa4erYNyGng2o2
IgvZmuLvCJBsOUj5hHbYCWxwfjtNzbaRPUpuQknMO22fyXrnZ/Bq3I90ZIFwPm7jpGRbvOB8TvF9
GQrZ4vDpJpv36Ioz52CmWhjCL7l00bFlLEfgxcO3eTiSBzo2PDN4AtLML+NVUR5SHMkLL9Q/fJaY
ya6tnMEIuMOj91wd1b7L8QJQ59l/ufxQx1eCoL0d2fT0fDbPHktJmECk12dSIU/kATknr9saKJEu
a3yp6qsKgZuIeMp3ECS/hxXdmocNC9jCGiZzW5KT5WUruOeGiHLFJ12o44L/mRlA2gvTsj9p7eWH
iMwac7d7ig1LBMU2bsVJ9etR3py7Cw32M0YWTw5Ba/hmR4CjLifXrCVmcn4ezucOpxte9k82CN96
NmVBETdMEKYVd3cPUB6OUWh7L6Skvmr96JEExJq74ntOGYZbObavK1DeFY7GJ6RC/kNXGvYcpwuO
wr81CXB6Wxl2pRTMmXy8M/h5SD3JrBeTx4WO2OEZKHDjpmaQznxXOTL+5T5W0oNoaxUxp5BI+cjq
z6VXQO5bAsTUbyKV6vLydZb6UEL4YA7Z2ypQtJFy+Dp+TsOYegkFlPTZDu25rM0W0CEIXNjA6/ZP
tNmlZU1LdzFppJ4aAkFflXJEcZEn8faCZoUyAtafz64BwvPiiwsyV2yYvQnpZCIgExR5P5z0k0mP
+2DwPiVPXVtatAxoBRImNeJj9ZF9wVDqg8h8j3b6W9a+cOONPcu57FDz2RbsPY9oCV/u0PtGYukz
gpxb3G0owmTY2kOC0a0b4oWrhYmMN/kksA34tdhgs9PURUkFYa48mdquBSB46kAa44kMbJe+vsi+
AIjngqNkAPx5FqLmo2Kd29C9v90IdEsf/lJL7zmkp4Gb4bWjpYnMxbyrfyxOD8gTwn2m4PHO/9Xh
ET2QzO1ddx2CtleoXfH0F64ORwUW3x1G+C7eugOh/dJ7jgLg6XJ5UgZzibwfU4AlUHe5h73SJxko
sYvZZPasOWgkrY9bnAM0Eva/qZtzXTw6CnQk39z6iHRZTrnGaiFUphBJNqoCdcV0+GAaBDWKlmX5
wLe2Ds7vJaSghw2faYiQ6lUT/zVe+STSH2urZ+Na5hHCItJ6aCU3vu889gUxjkOB1F7WSN+x8q2F
Gude76xMkgFkUEW0z4XIetxOnDm7aiEKaHSYK2XHV4m3MkcL/iIgt9TF9vp9KPhQhk99914b4bSj
1SNGNhJXAPtY/rIJI2HsyA3/TJRoN+VJC4YgkEGiyN+v+59+YNB4eL25DL9Ze+9/qKmYaEoaxfwW
qsqDehG0qr0FnjIJNPYuqg5691e1dBHvRbOBUZUoP72fmz5UydhObptsO57UnlJwCsKmPH52/4LU
hbNzyRVxwo3bmMNIrKnoi7V/4HUBX0Z0X7yZTdAPq93PTuAXMM6Pm4iBWbdsJ5sSEqU4NNHRMpgq
E3QAzS5ucTLUCMBYXbAUfYAE6tVIX17HYIPRJmgtQ8/CDH+TLwr967rrNI11An9HfcCK0VD4bjiw
9a2oU8VNIGKIkBiiDs4lNTwcIlkOqM5/mMgck6WDs2EUZK4T70eENxYWTeJfhzrPvNczL33p4QIE
7D1h2SoMWHnkA+Zw5Pb7n17QarQQh6VV1ki9sd6BRnd1KaX7yoZrK7m2sCGRk5ZtS2b6BPh49NGA
RO5pg6Yz/jhwYYnkpt+ne1IMH4hwcH+e0fSIHkW7fG1lQ0abLXobBGZBLFKxI4pwBfydH6eex6Ze
mVWB/jC4IVhIKqZElKb4CDxDi78ocKfEwAnNQhk3wFAnc9+80F6akBDcCNnG0VMuGFVWT0wvK1va
96h4fIDxOAYmOZ5o0DK+sVMXlyMFDQLZQ8TA7wctkFhzkhpT1xEDJWPi8JJGHgZ7UNyxwqIICmSm
0oeHAOxLXF0QxPgcOJ07hseQ9ADsQNfxfbngpl4YecZ1LIAwh3NPCj+G/Yw5/l4w5GlKPLdZuhQN
ev8YidAji9HyZEaIo5MMXsN7w1pZD32KW4pB4WP8srwxtlLytEiOdvCQ5iSsaYaegk7513Adn8JL
iADUzl1PkwiX8HpJ7yeHA+leL8Y4GFL7iObEHaHJmm7v6pio8ju/RP7QYXO4yA1ub1Lx39+hqEMK
ui/bnWFyNBwtLpL/jxn6c+P9aG65F8ZYiKPZk11qJ4YJeOXe5ZPfvLrEpIXxvUNkmmQo1g0rcH0V
VnzuleJaqUYbDXzPwlN7qUqNwgqz6+IoU/FjbMBwlcqx2g4+/g7CmMbgFXDDuLGYbdamy4SZ9chM
+fLzsCpPvEQkJOoHIJcGT95rzJTBHawPiLtYNtzOdtdPVKjaqLac+R8epm7zRLIR/7MT3LjKb7yr
2zCKY759ymFsMchXKCxa7S+ueseTnUe7NWNYa1ax/0yBw/vZ7YUppoRxdUSAUVRATUsfkYISSb3G
y9HEiISJa5XJJ38lZgCD7LYroyzDf+3d7CaYhoi3kYUdqe9pb54WwmOXc1xquqq0R0GupT+Jev0H
c124olEHfUIlB20QQGcMvDNqmgFMJKftY4jrtgplW5X8P5q9N6XMxOt3+EEPT2CA8NHBFxWnCevK
z5gBnCNDqFJXVsQ61b+t9nTPxMa12hfFC/gYphteMHK/zD5OBoN1vICtWoCIO8RpdkErW4qgNk5O
o8ZmOZBeA9Z+Ut8Rtwq1G0X4rkAl2ycoVJVwyFXJlrY+6oZnFRT1zYrxVDXrG/S8cqFGcTJKEIgK
9uKT/qEt80uAVs481nZgeixHZIthwRveViauII5Qou0mXndVB1nuifok2oTxByLZXau871UioTvL
q0pXr3lkkcR1TiQYLL+lGHwQ07GiO5DzI8xoMyFo6J9r+yvWjdmv5gJfJIokGCwAralSPI8aWECy
2e0M3sw5Ws4YMQHTcbZkkfWKPt4Wgv4nGVGQAWt+oAq7dGe4LwWfW1WFWvHMgE8drpBF1yseu6bp
svGo+JKHM86c8XApWGyDERIxJQL8hS3m8I5HMS8j6tmKC0SUSf2PRx6frP7Ut8og5ef0hc8mPSx1
AQGSCbPIenKGw7k/Y1GvDY6AS0pGgst0jpo0SJXnR+3S7PKl65gOsiX6OCMHYLvm/PNVgkV1juWt
GsbaWx5cHOqSgVwd17wQ9numtUYPgiqYeBvIadaBm9B2tKTz3lSxhbxu8Z5vAyh8QQ4vU4v4IkGi
5362WgF9hqKS0AAeRtDGBIOkGFuyjoSNwDs1kZKYmp/C8XmbVammkgLf+WeWHG/zJ3Aok/ecOo5V
sO5Sm1p2mz3n7HHs2e2PDv1dH+zB64PzQcrtwtJTgIjJK1ioxi1xQiOMBx9V0kZ4x7axXgcDSEIO
nqW1zTGDCqwIwcQR6RzdFSvF97Kb0dQiIL5hMmR2t/t9ketvcutgj1zttHMtHzH7rA1zlfNsqnD+
1HiJGRMQxKwZ33sLeMl5YcU7jobofP+3AiGzkb7GtETMDmXikrKnbonkNQvdgUeXuZESW6KjoWFX
G9YJI1atVwJuhsykp46k5XL7KgG+dghcRsmzNpSLz8PHq7RM/DjFzjUAsINFqAUR/9xyV9etRhHd
xU2cytxh/guu85LZhnHDg12aQ8FgQ4GI47I2kWlzvQ/2r/ZnnRJkH3NFPE5GsBQU5ZTDV9AstFwF
XUyJRwS858ObQ+j4IXkYSSn7gho6HRzJcCJdzEq2mBuhtgw2JR5SE8HgQIBYh33r1e45J9yhR6/l
n7x4rdZ//9Skxwsawq+Fv36Q7n78TgK9uwd5z3fTFxerslrARXyj85L+wjD8BJ1XUdpXGI/iIr0c
t5Lltg9eGetqSjNUbCpUd+AV3ZHMztS+YE5JPg25OmYBGA4bGHghV8XHhcpDfvWMHrnmlL9KRgmF
2Bptpb0g20wRKaPeEHrTMslgnc3ERDRuZpBEJ+jrcynt/5vfgB5ggtakYteKOI7WjQcL/KGA6huW
InsUalxfAMOBlBZ5STLZ8il9XcJpffqY11iX5hyFn2BcixVNZg9dFLNlWASlt5upNyGfUdN1zG3r
THF6UGByJTo5hakMk30A1BITnLl5AfC1NlNrLl8nRA50rGANFB5B3lKmyUgA4a8bu+wwFOi1Nbi6
H4peCV5EKiLsFeJbn5I3mkGAlw0QiEkZ6kXjSkF4GSUsxmOH9R0kzOQlh/df1mh7ACovlIMwPyFM
UW+VWZSsB/JNOANP76+wJf61+LbbQI7wBWDRSH3+n2NwKxuNprV9geOJh8L+8lZOzSWiejUOOtZi
PRa99jzN7nK2zt7ShuU6yO4eCH6AvudhfIlftTqgl3htStkO/AbZJT4chBve1Nl6Del/Kke0Ab9o
idTrketNKrL2tNQgVOdebM9ZnkKi4+HTyABaX50eAOCNoocRzQB3DmeVurvUV2cBIp/QlkDIm7yb
4UvoQABehl5dGxBoRFIaOBSZpv9UXj9b2cRmAnrpxCqUpqL/VUmbxG3BnwMShwZ4b6G0lO3MbJfi
6TddIHnmoCDim0Plo6S1URh9rXuhIOvS/dFYglbNN8+0sVoXYCs29ps1n39HYtW2zrgZ6iOrvI/v
3leoLbwCcjNQCJB4ah6UpXtMmTFiwyzdX8CGNyD6qfala7tEMZLbncJ4bjHKeBC42JY5vwHEA9ZU
3e8FXEKdGBzbp9oNcxOVB/vEzTAjRCFVO4XY1AkcaxyU1j23Nd098As/ZBDHq8NdhLapNY3O4mWh
7izebfIwENWBBeMFW4H3S4BAlx0MbrGUjV14cjdlqZjyDgLcd6u0AqbPzox9HDebcCIxpzlFhDTA
IsYRz7DVOPwPC1Gx1sZQEnyWmEg06IeakF53/BSR9t2Nc4Ei717Dv/CeBEv4+1pKMdNnZjcCRt5N
V611VHvnTa3EK8lYUlgP2WT5LLGJ6nD2K+X1EFWZ86hxbzlyYcsJxQ/pwN0KLjxpmDP6FTH/Hz16
JEgn6k6FWckXJ3Q7GysXIiXvq3gjA+DijO3A8ydKDTSdapl6Mb09tPY4sC5dQ4Ry5/Dhr389UUfH
C4L22GhbezHDFMcUm22InKtNmtkRaHd9kYP67Itf26E5kAX/ycZ+bgQGk/VdIrqo1UrJkpxpWcFB
iSjndDDx4LYq3WAOkBt9TGBp+zFFIY2AwFKwIji8l0VBMM1ELnmKwsuY14Ii/9DJer/kVp+NFKXl
RkBqOPari0J2O+14aTlUb6y+VZQcrmyuwtDIn+mr30MelhVciDUzJzQ+oaM5fbbucTO2F0fsns+V
LMd+nDXLmJn/7ZS0TArpx74k0Ahot9jKNpxZ/4eiv0axtE2U/Kg6jjRNze8jSny9N7FBTTzD6wns
mBf1KwFUHzl8ex8rnO+zo4CpgAnOoYgvWCEM/OZHhSzG6RUmckDEOAtFqBbY3RAuGwUyzWLOpuvp
bo3hh96+P2nsnkW3Romg3KG1uFjH3XlOAaO3zUDMAssSvvcpD43lkhsmeFOxKr0MpEd4QI82HD8W
GofAODZVmfDtGTVETUUL3GmMrPnatTIQRXAhaUKjDYQTWHgm0h/DywviEdZ4kZQMq0q6UEePzNzg
qGxrIIGI95EHYEzmDpCHF1PbdUpQYzR6S1WjVAs+z+UGUTKiJ05Zp3oeFoMdj76Cla2ekrXpc8JN
9EtWe5rAdr1QcC7e71vjx63OErJF3irwaX0EUPHrewsmHtgjFYwKC37nmW696G0EVUmQFYMcfJye
yHABDnKHCTA1GC/wtzKvMx7JOaFV5BoZh7ULuaMNfJdOG6Dt5ktVHpVCzTMxNkTLtyeHRSI2tff0
qfxgA1j4tDf4PkPl/gTrIsW6g1s4AFev11+mzlQ/DB3IVpJVG2qd/nPpe9w0vpyxKYpj19lJwwj2
4Uf5EBc7AmgsDOcQnTBpUaQXjapkBlnbGniYozWKEAR3yN652gksRoeSplNSmGpMwV44Mqd/RYcM
StdRBGowZbZi/R+MU0/1i7vOVqdQQRZSbt9jS43UZQ+z8q2Z/i3dWckSpLARRZu9LP+RJf4go431
2RzDuQia2dwFbmLffFgyXzdQ69Eio0sjAc49xCIzlWQOmPiDw5gTa90j3Waom8ejMmlDE3ZHZ0i5
rUumbGHAjVkViUPK8djc0/HusCanu1VptiJMga5wdQ5zFUqUxkQcoQvqBz1mirXLesQE7x4DOkUd
R24VUUZ1GBadM/1q1zH0QwTciAAxg8H7tTlyY9eoGtmojVbyso8BehVu/cZUezrJc61svLlqloEZ
mG5UMB49xf9RMv15jHH2BRwI+E4e93Y3WCoIiw8PhbvACFGHaiWcbZjDP1BXYpmtpBoe7yOpD1mt
KXehqpqDXH9oER7B/P0L/aDEXFyMw339VBduEnDwrdjQPPkIOIUkKyZFf0LOo2VNP+OhBxKaCi29
7EqtL2gdQKNfL5odEfWHrUe+i1x3/2Nsuc9eQjtP97xlMJC2Ha4H+4THiwz+qJR3OXfVOpY3Ii7o
LhWth4TEsicbCiJE0HoaSxdxWSyKi3+qg3LOlGA5VpAgRxGkXmKFtp8orVgAzBmUMdcd3feIjw6H
M2yeDbDJCqHmEeqJNJPW75qNCJW/qLSeiJQ2BaGC0eHPH6M8IwuaAHYHd8eT+/n/C9nf6KfFskpR
cqBxj0RIZH8nmI00opjZCKVrsOk03oVhelRA6A7erdunYXoyCduu1N/WPC4ape7ZSQmBo20fP51q
6xSMEOYj3gv+h2GQmfIn0Sx4epyZGQHQ0K8XLmJy294fjMaR5ea5LsBbnkT4Bz55gN8ndne1GnIs
SoMVg+PluE6b2JPMv62f3gm19q9AsvTFit35uj/WIYQ19SRRMV4EF6qLi2GXLXvd97hMA3U2pmus
w0SoSpXdRWCDZ5zm3DXgVfF9o2MOlG2d4Fcq0TELuvutef9pN1j7Bj1DVqc7OxJNJrRuWMdxhFEg
NeheW5nzGUCU9dG7bUcypFZGlR/BByjh+YtaEhzfmatSdlmr9FlGLaWpCsrJkWTha2N9PJUIG0wq
/w6gVJwC73abzlHiqvNMvetQVFnYUJtnOnbXVhC/9cmBJW63vr2/TSdFVhxmPwKkCx/35obTRWsI
gOstuxmJSUwci2A6YCMb/2bG3RN5LS2OBdZyCS8XVFEBNePZq45uC6wSSmQhN1kbvQOgUpcQXPgm
WD7XVgn216SuyFQCdgQ7r0m4GgdnpAWt1esnCpxtL7a0QRvskbn5bYrhrndox2tax/pR8DHeVQWb
X3hhky5ScXu6JY/quhKb6wyMZuzpIp43O7D1THbqoV911R5UEeZxxTnpnSaHDVo3Vgdz/2IZg/hP
lVlW8F0UfOFBsPB8Y8wNU5mCgKX79mDhYrJ2we+EAM8TJHRdnwR+WWSboSa1mlgeCk3XgXezBuNj
P9z0SXuSsIc8WAelC96H2XgeN3RQMfQ4iTkz3XPTeLbws/30TEzvHkTQwW6DzSaD2RxfMvKmM+SO
Oks9ntBiQoV83DXDv41oPLvtMtQaHox+f/i537iquo9Xh8IHJ4N8TrUtTitXro/sPO28WYCbh33T
7PuZQG6Y7YkRfn6PYSYxbISQj+5zGxs6vttN4mRQecdzO7Js5HDoWdU1wpJ9v+MlvE+CIkOcySF+
xlFG2KMmeFCyp9HTbB+nQzUzt+rN8DBRAh5wma8rZlNYpjNLaIT5E/sR/UZW/QB4rN3FT4HfAlg7
/KOZPDncf1DV7lvimOAoZdBKOJeNNDkmp9p2jGVCUt5YNp6PAdF0ul/RLtNvVLVOaaukBNFKzrJr
iVtTBSU99dsBJeObhf7DYTOqfu4DbaFrYJOrpIWVV2ax55MAy2lhQt8RKUfU/x5DTL5vDn5TiTIJ
1VrbBVu7BxVQAXZkwIf2e3DQlY1U8TF99WuPIBNv13H3dAejOP4Q3S0Y9Do4BJFoLX58bUJ1e2Z8
TzLubdXedRbfRDMQcnM3g2yZTxTNI/aqYVxibOo8Pp7cEFbT4iHXdKb8Mm1+/bsEGsTsIxIlKOM7
pQPFiC7ox51yjlclC9xXoC6wc91SZ+Jd1CHVCToOJkc3SkozYSCD10KX5+AdXNx9sLxXDV8pRUyD
Gelj3KpdxJiMFUo9quxG8vuZwRWd9XE2k7hPiLoZ+hJvfVSqaJeoyKtQvAOIv/2LA5KASnht17Pv
DYqrZa5os49lEnZr0fp5cfHBzGsj5leIDiEoDGNNRd1XksCfNjXkw+hHduxXRvxdT5MuoCw3sNpA
Tr7Ee6ZSU/ryv6pg7huk9VzbP0jE6UdDzjh9keH69vgGnds2j+MOIrqu0lrVO8rsdpr6SAc47T+z
16iRzBmpUk5t7WyqM2Yz4F3XGwJabOMmWhSY/U+LBeJ2HxjYm1A+D2/ygs5MSkil+dJLhR1NPwY+
kj96yVvZxYYvXteUGD8cDc56n7n8JJzcCnSdfAFS6sMxOLYFzllujk5GCRfoiRpOz3h8Duq6g2HK
/LbdwkzM4ten++mhow1RmvP9ZoXFV0PVM+h/Nze2dJnxMibO7EMjkcwKMuAb2PvVKi1yki9nkEv9
XxkvJ3ycjLEHczjhclq6UO9x9T5cd7EC5kUIGBS2M494UEjCyHrp1Vt2C/l+bedQQe98it6AolWw
+V3tkmsmQ0+3Gyu/nSbqyKgUSmYJXwGXKYZZCA3CBn4JrViiOhafUXD79KF8oZMGuxICWrRy5oOg
GaSfcunEpgcNz5UPLB7rDEJBQRjj3h6EoCnwGq6Gcm0L8mUNk8SUBd0Bv3DRr/b6o/j3bP/WK0ja
6bgoi6Gjv+jAW3hET9aJkzw+QCRQBXtv7NabvrmQsmop77GvMSZVD5LCs1QRnQMhw78eKvnKcDlz
mIrcjsdBJAQrq83Hcc1Lm8xJ8ELYgGuuLzOch8P9WEgu9FbmSTX+NPZjSAnjaUvioH0jKh3zlje3
HuKuFWchfLZIAoXAgZj4WmG5L9fYr2d7bkl8jAgHjDhfvixlBv/CsaWHr5LMELAyPrA3LeAV4MBK
aITj445ojYJXtf+IkawZErJaAcS/TgdQJcE790r//Jb7LCBQBPKtFSU55wQDAXXqDS1mww+Y0Vd0
sydtFAFqHLgoz4H8f5BR0nWZr0AiMD9AmVHxLe2SnQ/2BFI1vo6Atvgj/c6/k4NMMw3NmJC34c5V
dAHsvQame1fCRICLmm5tna3ndO5H+IYS0CcyPHhIFcTaqEWwlR2BdoCm/LagsNUdVhGb6WxWUVFw
fa6fkhBxtLNDMo746QQV0WDCDSL/aCVKIy7JWcsg/28g5SlSbN+rGs1UhQnZMykQ9Gm1TFEuHIo8
MGHW4bOI6mvbDxZTqCz4sPJgYBL5dk5BrSpXw21Dak5PMBIInE0IkUjTgBiFloDlWpDFcHVZZqLG
6p8CKL+qWPJxwJeDPyu+w49p16FBY/Oru5z23ynIU5Kkdd9PBIa4tyhqAT61xPYz4LwEBT8xR5jL
hdwvIQWPtcxfjHlJT1TnL2Gy/UgazaqnmLyv/LKRPP0Ey8uyafX3Uf/HsR/62fO1K9laGmmpVPij
nfZ6R+2ggmc55iOUShunWcZo191FQQq33f7TuGWkFA+/0K8+FeWQYMi2BvbZBF2E5iJcvESL1r7r
PthrjCfj++S9r6R9TvD9Rd7Mtq+oRYCglD3OvfgFHMM3T2+BNwAnUAgcDwSOy/YwOuyjkLednF4V
D9PP1FHNJC6FySwAHm18L1Of56G4HqBG5e5BEdBH5yP0iwCxniQmTcxLwchjUOAiNAYnVQqVxPk9
m2ojVcYSDxtK11MjvGJKRpBqUa+sEWOn6aThQJVeqqRpb43piIOV+Rax141a027NkNAzRuozawdT
kzw6PafdOP3DR0m9gcQJjk2+ib25QGk7XtE8vzJRcsc9ABKtMguSkLn4wgaCCHEE5LXjYhDPp7Qd
dC7FpOhuubiy+9XGBZqf3nSmUub4wP2WwJvH7+FufXa5iMn53NMoqEEaTlLlGJP/lz+OFb93BLhM
WmJ1AKO80/ByqrCt5741siAYtoM2HmmLXJMgAdRh27OstGi+/hmj6DG9XvCSnfIZ3dlBZ4R398ib
kdbI8nptbF4VBdMNDjty9vw9Zj7FTUPjHioiqmIDxipAyVJMKk0MQf7nyRBfLPtywhKua6mZrnP4
W99+HKRY1MMv0GEmJorK2wujc6tQqVvbn+Z2tB5ZUF64pF38LTpj60zIyybl+b9l4YlePnpbHSk0
4hDzhBxn+8oVU5BtaCcdDcwsRGYE+vXYIv0u97NFVsgfWP5KcCYZQycZQmOhOZvQJmgUKmMc5vd/
GQ4eUNCBEj9id8xm99bvrvQiiwU7BHMwQzZXzabxdIGpo9QYP77S/9MH1LpOgR/M3RAWwDAUo6N8
dWtNwIeHJLs5E7fEglWakPcAwKwR+Z8/8s7yYYw8YUGNbElWbX2v3yH9X5ms1KqFVcbW34VXcUTv
b8e9O6pEcEINmNzJcbyHpJ6Ja7jXsyu2NHqUANEkAbLPlnLUNx2vqD9OCix0jLf8CQW/aUVyX34f
slz2arOE6V0umLQkYyS07Jl1WlHv+ZJmvwMuNkQTjRuDAX15pzR0fK6ai5dz2i99JvvsZRneKkHe
JwguvPnFh+4KB/vgBkCiVqp3nkmnWfc/CDO08fqLX88c2PojPpfKYK9fqXR7cSlsdy9imPX4MYms
25xjnSvrf4v5E07lQlszU0U4meBBw4Xm01IA9NblzPcYEsMStxe8TgyHSK0swKt8WD6STToSeYEU
MtQ+uAU2QyKLPPEk2+iIxMfbk4isUbTSneSJrt5/Q+CUFGFxt8UNh+S8E1VKoIW/ZZdW5rDXSaYz
HKRMuoxoCv+hmvfTWvRDonpMB2/lW/eFzqQGNzkClqRqdsBEK2+t1SyYOgiJPEfpD7NGhraweWNy
DZL8FqN66iJFa9G9YIAoS6FOfKz3zq4PgfvgsczRvhYuJxj6wVrLPOXOXMaSaxsue7YAJFpBebCb
MVFKBYmbqsPpNU+rZURABopAi3iZQ9hooRBjW/Ps1y3tmQQcGIP0TZ9eFYLWEKznpFufyPMC2X7d
NyRwrLAcb4n7my+3h1XquT6CBIloEKNKhOZ2qv/6N/CPtIvvVCQMhNlVMG0tT0qgcWG3TbMvmD0p
ouqJ/g7LvfsHUqWech8wJsZ4o9dfaDnJPcr+CwFSWcNleAzML1PDHphCNxp6PNctJvMr4MruK6ds
FOjH5h84XdnbDJaQ6xo6YWVHLYR4CDQjvEAmgZ/CMohGwHjtFLMpOkyPM8Gae4le5rGZid1VjB7k
ikkILPILk3ycdWHzzb5Nuxt8yh1ttEJtkGs04N5TiR0oaUMN+qz5j6hjXWXMFxOZvrFLm8K4r3M7
OMP8Uquxa6HbkBC6mLztHIS9ob76VNECRb96GZnQNGobNj/mhMzIznMiomVG4rJRGm8GMfyX40hO
oCVWJMky66/0jA9vmv4P54+zzUoAk9e8myanm95AJ2bJW7W4GySYcGtEWDtepqQh4GBG+MfS33jV
3h4nYaR4HGQ0Yub+oDTjcaswpnfqcjDYKBBav3FmPWKNlox119rD5r9ag5uBckeS5/y1690vzWA3
CLP9GSgidsKDHdryqZiSvwXY444ErhpTTlGjTblJyrDJH8xolN8mJ6TgQ7uI2ymcwgRbcioRRmj+
FKjvwRJP9290jKs57hGTLE5lnorDI93f49R3XROD7iahEJrnwxEpEEYsEezK20hq2vxeWBQuwP/+
/i94AHRQrY/xXHODKd6IsHq/Oy+H+nxbQgWWnvAz8P8gQTgW6TCRQwyyJ80MZPRMO1Vl7ufhD2rP
duSWnzxZpQBJLfN82Hy1B12FI1JrIm5L5NsX3ReIsV49bVX/yED2nsNXvUJNGXnlBQpxlme5CH1B
c7GAxxynTT0HHZC7wjtz88Z1jsT107FEDkKN8OGmozTBgzAVBbEjKD+0Wsk4I7Zy/E2lUVnSjEvy
zA3SImeT9ruTTdgnHeVDHMLdRIoiCLwj5kgr3EC6f532u+J0AqAVQAEilryVnouMAgL94EJTwQmt
SV/Iovie16e8HT8084htztCZ3/vv4h55vdstwHkpVmBvSn47FKTSZnuqt7OdymP/TBD4laXnCpWF
fzkCmmpQ1ojVSEjEFpR8Jj27z7rSqe4pXW5XxCtmmyG6GwXwFSvrGWDg9u6h3Ncyp1vURB+bBc9j
0TxrwgV9JBA1WZyidmktYW49ebqD3X1a6G1KqpQ/ZQmrFJXazz1orQ286nbjRFM5MVD4M44Cj1TV
8XEsAAEdkTD9xq1Lz0S1rM3LDuAw58lSA+2z/AbiM0RZEsYm1J13lSawgXXN0yVIWeAchTdfS+8O
LT9fXqO8cuFprxZ8iQtCUMqAe+UNaZoL3n/EYh41koHu48ALwcjA5hJDdjvdkCXkN8XOcdxwGlqs
DBwzKk4KChqMfosCyUvlwWIjRlAS9gf6jrHLLawiMSmdY5NuzEkYuCXSUO0KMdj12afw0pifiSnR
Jc5wU8ITlsK/xsxBF+hdOSJRAWcVcggr89V88XV7nFDt3eeXrVnrU9TJhXvStgQbOYofr7FAaoOp
3ryRVLGyt3Urw/lcawBTl20nj/1SsV8r0fERR6Sm/gkUWmbtTxVYcBamPCRCj8fWeS2kxrvpDbGK
dstEB+0Efw6sov+NF0HyFBbQ5W4dXVYhFOxtsolSiqFGDTeQ0QSehrv7+2/bce/of0r7mfFHSVes
hnsR1wgzfZpDe82Hqh+aCnW0Vrmm2UoDymC31UdHvhVtsJxOIVTx5d6W5BdHwYbnzWRa1RZzWQPJ
vxaP4Ya/wkjw15LBvD+LtiOUv85j3CayJsDbM5hp4BNcAnIY1DTo607PoYoS4ssf4p5V2KyMlKA0
fEL/VHVf1Ecx9ZlUUsZrh0546kO0ht5GyQZaHBhwJzIyKjDj44mFQVoGhVaLBGGqOB9JE2IAV9y5
N+WKCuAQiwFKddUoFMFE76UapHClWfJLbjf5YDIIM9xICqrBdHMP59z1E6gR9E3YXoxLcS4caKrc
jnwBpjSzqem4AzflTqF/GC1KmG35pDRrTbRoTuEjGzD4WMDr82IC254Dpb9vj16IvBlvozJHXJ01
spA+IKXjLZEFxFb/yq1kWHgt1xpZlwRQaQeHb828E7q6StkKl/N6QabacmvM0w0ayqHh1qJw7e1Q
eiMB2/vOM30CxdJD163bdweuLx69cvK10UdBu8ZEduhylg7hiUQZNOlNOJ2XOogBbRk0VAvaLH11
OfNvddC5EteD0m2PVufAGiy9bWzrFVn2Drg4bOh/hiNc9n/PdpUxIrFw+z4d1WHg3sAl8wP9mzBo
2yvTnyfppXBexMZghXTIvD1IVA/ILkfgtf1CuRWkzzXXWx7NZ5QtODi+Dc3dl0igLhkv6N0fLB9u
x7XStPkBUSRaHulQUV0YQNBILqGLk4YquAOczPvJoBGlKdzhcI0OqlDqQ/pfb8pscLVSzW/tk6X1
Vfe0fbR0taiBZ80GDyOY07LVIVNp7dPuGpImp9TNpjm2Qr2oORabhI2L7ZIHLmkzt/RLGBci7hwA
h46RQSVrMe0HGp4MnIHGbERAGHyPICkI9ST6pgUrWkgDJ2XqJxVcJb7zIKTXOhArfjzEbrQ7FNJG
XIRJVJi20rs6xEeaTou0ibsOJVP/ZUc5FGBE4SeSCJuXfU1NrhyXQT4MnAmcafpGSYw9KCjO4PbC
Qm7pNTv29UZaZTY0Kb+Y0twDOq09FkJ8IYoFAMe0Lpp6/8DEqRF/EbCLrX9dTnuNbJSu9STc4rg+
HCoaFG/PLjbwp4EjqdttAQOcBqslrZLhZyfC1EDdBG3oKkCD/5vAWFZ0JpMOJSrLNFz102m2JiKp
umZB592cuZ1gO9sgimpd3YYuVXnDDIz6NKfsgsFhVMb4oY6sUMkaj61gueR98UJS0pvTII0XAUNY
PwkLcDO5dxuIYOfyIh8LNnnwX/2H39rN5zY37iGAcqGJ5uQfHH8XI1bFmL8DxSwFW7j583pWsrap
Eb0scHbtWZep43NuGKTTSkwlAdOj2B1LSNJohY7s5L4IhVoKNlg7pgtRaampDHgnd6JVlJSMuUWp
DxzYYgx6auun6QSRNd+zpHFuNZ05fWO6ASQ4wMDaObURIaJ62s4m7Vx/iunb/zDea9qDUxGAHyNU
m1uYKJOHcxe9UgDaNg5IM08Ak9prcNGtP7Gli4VYHA/lmD83GlkAklak5crt65BCFbhfZd3Pu4Fj
wgSK70ZbE62qWWTWYYSl5e2gI//e8Z6pZsaX9z2o4FPCYifW6gW4IXeBDdvx0Rcag14I9c3ntHJb
ToRdL2mLeWnw0B20QWSVDTFEP/cgTrHeMmIeTcMXqRttF8MWTy4VMrYGVVBoHzm1u5Zr9MWyWO1I
7zUfvwyov0mGtEioxsyjmaI4qKH0OULGzDNVCjjniXBCpb6tKBlIUW7OBkMkus1pZWlfWa/aTDxL
ss+G7qdboHXbIqeJ0ozf/CNVtN6P43Aev26vt3FoKWj4eoRREBIEAYM/DRwgqddo1TDZQLQnOYhn
cm6yunPLk9VUZUmiF9UuD61wf8Pv0bmRPnXmUHcLIAnKV/bdyOs821OtS33y6wqjzWTBFFPQpWHi
hIPPWWnXhYgGY3d1obQpNHRpidhKC/W47M273+sQFJeNPs2LojhLJxDawT0m2Gja1T6IGOFpaOxc
2K47fpu0Uec1J00se7MMs2lg2fQuJT8ABL/PGOqAGC8i0BIYgV3C5RdamGYqiGOPfZInMV3r6dzd
ynjH5Fr6AniqMvGosRl+Z4hVFr8gqK4/eE+hFIvYffx5AEGLk3eHcRdI800xPFdC5+IUFgt8S/jn
OZd0G0R5dk9CJ5Yx3US5RjPk2VaYwddHMCKjDUChYCCIbFlnAtw3I7rWIQeuCrOvJ563QB+SfNhZ
EIRfdR9ZxI2aWqr3f5qJl+nzTG6OQ0ioQY6gwvI7xGfqSncmSu8UIQK8/IBAid3lO1y67jghqJvQ
xBsOqdULDNv+mXxALOY7KK5OcYgHM6pAClax4GCGrNB5Ea1TCj4vcL9qKEATKgBvLvki1sCoyYbg
0INXW8aRCQbLIF0717C4b6i4g3Bnjwmu1KTjor4Wn5W/9SLjP+ORJOcTBheF8uU8wvW0wnv9xhVw
xoZkaopwHpwqLmtxu/qLCEzLqDJlWhgNiaA2aQIgyMD19LYtLit9fZaRN+yWjut6H5eHRfx9/KLI
DSeViQFpYDiwHjFLEHab/lh3Z7QJwURh9VqJjxq04niK64vi38eL4S/IgbSr/2UmlRg1EEhXe5MP
98oOyy3jLMdVMYfbKbO30jlfdJ4XlDTxJaqCmTEiStaDZz9P3852AIZQ8ZIGJv0Akh8Ock8LaerW
9tOm/FjrbIIAhfw4gGAO/uDainkDFR8PrcZ2ll9enPLyaUikzs22XMMtfAHCH9aAO8BBtBZdf24E
7GVd8+sb2Ppyg+Wl9MKOWgCIzh0cqpCL/vuF4Um4KwW301bTqjAvyWEURMoWuw0JvrVOYSjTZ2+x
X3t6q0XDzsjv8ebfxpV/20tsoskPEUVhqelLnsoQI/qD72u2nb+qlvPfyAoQDZLiE8Lj524TjKsR
JWREYkRJV/yXJk8ACLhLbBgwUX0sfXosVB5wwsC9zNl0UMVdnoh+mIIphBDjYDMDEKMhVH5dV75Y
fMmdmmB7w8o/mu3U4mCSr4O5Ft5aXt1CAIJ9oScaJy+BYzay2visqfsD8lBqfJEdMfVGFqS4mR+V
MZkf/3VzO5L8zoEnejeAK3uE7yozshg8JsKd7rXUDHRjrcGh+zp59GYrT7A/ZjWoFDHQnl8iPSSm
5n4eGkTRxmHj3jE/F+tjEzm2sKCdc8cm8BXIVqcbhJlvO+JWF9s9nHD3DBuwgYjJGfitC8X3Qz34
ZErLazMRxjgFHsHx74i4D3h1er84P0gCqSOUxkfeZXOoHNHN8kSn1xUpFVRtROMRdJ3NrFyuj3Gu
TdAn0WEhmpSXuySNpLySVb4V+zthKgv92lNQmJF+CXCaw6oxwueTtjnFdNpQph5dXfY8e6Q6YG+X
XfGmcPgkME1CXsfu/k2SDEWxoYNKtjp61nxtXGQiMQNIHykYPto58Yw7bKX+w0W/ciBlj8STXs1c
9JnfgvKOzFUX6BZaQ9+HUMc9QKxXdKC7B7+TNJpO26d+nPIr6CA39kcKrFbw5AM2j2w8V5np93CC
duA/P34CTh2FEjeAlKnVkBPimbYCYsN0XnWVDEP2ivul//bjAdTEcMDYi31j14bOxgZkfm2C8BOi
Bh6SuwRGml7uqRL4TWF6tsMpPZnjX1H/czO7j1iIKASy1P5MQ1MkQTCqDDoL17brvmWCnuUIAws1
ktnz+mmS/LSwqTn91oZqbabMc3H007OvZCUAtrxS13yCNAOF3gnEIXrum8HOjYq/H104uHFz4sxb
1ZlQLqTI9mKaK1yteDL1SXJcfJym0MujHDXM8TV1wgIKLdKPK4H+WSi++PsLV8Hq3EBafAskqOS+
NA7gumyoVqitOcCefTM4L3Vs8KYpsveYm/XaMb8YravzfZIiX7ImnWUwXT5XrGNT3O5aOI2cEpSH
pLx4Y7OJuf+K1yDtby7G5PtKz7uuYNn10dMuIlfsWTGwHkOwwe4HyO89O7K+wul91Myk9SR41oV5
KfHAzNq+mFU4CshewdKDEb43dl32TTdasv9wjOHyqdMrIbj5+pRBz4HJMnTCSMkN6ni1Ek2oj3vz
3ypbIymJ+HKYt7/ziOpmlqX+etKBKs3rYL3okVbheVSmJWiZGbFk2KRZtH48vtK3URelpYofsywF
5sHhTKwJchAO4FhaUW4EFHp0FycsFsCMGAx7mKyLREcuFgPZAkepIMDRyJQPpEZ4AFYnV3i1gnMd
CIruy82YTwjHFrk27Zo3KubJ+2AfRrbEO5MFbG5OeUSOA6c56MUs/qCqo/QaIlTNxSRrCJBRd4fh
1B+yalikGlmUsgibycMsZumBjOO2VkVZtUdoNgQPOSkmlOvaN6RQY6ou9Ftdc4Wst71QO+5RoVaJ
t+98VrTMkiFfj1Lakbak9PImwUzv8BUqwM/M2EvpOWtYHTXvAg9BMbWYjLjciGSfagcAZ9R4qcPi
N08v5eugofORnYSbGwb5d/5aq1SimxbohCKl06Yd11QL2StgU3lMHWH5gEo8+3+jatOHevlkmy9L
EF/1vZN0XLzx3WaUEIK/cNkI70i1RMMd9BRM3goG2a3Hlwli8DryzuXwJsYk/CijqNyEkJAUDd9/
G5gWC+R9J41pwhhxJrNiVRQXIbAvf+PdLpHwBVM0+yo/TEHcoZAbPijuNSGIZV0+sdo7xVrfLSUj
8r0jbV5E4NYzcSjTaFzJQjdbsdKujowvttcFl512WekQXjHcDSnC/j2ilVn1E+2eWOhlVc6gvuyB
jbdWhNmxGK7aMQpbUz0yxdsTx6rseXL4DwTdacNiEf2F4rW4qv6zYDEVl+0NSZHvSsno3ZwTTZpU
X1SQgslgFEfhL0sl5qp0TFH+6xvaAfObWb+PSI/ACSp1tSUlJhZuxrhdiUMl4kapzDhMKVCaBH4h
wCCNh+KWdD9FzlOL34tk7mesNGT6XlKU0cb2YM++ia0pq3H7Fo3SADyfjDRwK8bOTvnQS5k8+HHS
q05qebjSW/ayanE+OhSC/FuPum+cflsFe9CQAhDQ38CP29Ls+L6J+twEYm8/zEI53uR/eckxxYWv
z6qsIcbig7Db4duY5bJl/Ew+N+xcYhgrdQom2MOtSQll/hcyuwAwOEILP8WB3vS+B2qncQWn7GQL
D0eDzBtyBDvGUVNh0ZKjyNFcMV3PrlW3XubqgH7UcgqhE1BY7pHnKd6hniDFdW0kT1cNDSUbU+nL
ZDCv924sf0VM54IcYKgD65gX42u8ikOIboBjM8g8nPKU5u7sIANL80r+xzO14lRuqnBVs0saHZk1
z+Raj2p9PAPE8EteDty6EKgW8gJKfDry4W3UX2FfBffV9XwxnqJrFt5eJ2LOGKGgeb302qj/rHAi
nf+yEv0CBtsPMfcCV8gwvHVI1ogC5mhRC2tLXkwrTJs+zlAktV+GTZKNtZuzkI/S31KmGgY/g+Oe
UeQMXhEzEPBnYhA8DlQmrsgzov1Vi6B/fFp9SvQH9Z1t8lOF4opMxK/T9YGiaOg+5JHI5azEqEkM
1ZWrYpsY6aoQcEFUbjIGWFfyXinTETKzpU45E1HpCeaXYZAJKvGT6NQDsc5EVCXfk0WIHQkBcX1X
nM+dp1Qm5AuOGLI/8uhDnUww1D6Gb5Amf7XQc0w5viwG8px582nWQZI1t/e41MYMIjrrF6NR/fvl
5g+Wi64P3ykAGK03d+iJvc7w7hquhWJeR9SVHWX2riMDrFIhO/Cawc5g7g/INP/j8Ck3xiQ6xxGT
qX3q/4X34sMKiu2DkhOp8QiBBBf0+E8KRnwggEGpDinaduGjoKij4q4S1kLHDY0KdjhNM9rR4qRq
ac2mwkD0fxfqk+aPwumiX9Vrn434IbMyAuaev1fqfKoaqZw10tY7TsEQ0Ncp1Q0U5ZuYjFqqtwwk
jgNtpORnWX2HIM8UP4Sx5VI1/LJvl80BAj/ukTA0tKNH9d+JKFx75agKl2lKTIaibCCzejy6pPK+
gR33kl/i1t/VDTOTiFBGnkl3+fIV7U4jeJ3fXBnA891qGUvI0KL6UdR0/u6c8xKRVGsl14zhXqJn
ijVI+0tOWf7glqVwVPj9sUWralMrbNbjo8TpESTllhLcZvAEYgid8qy7BNv5fHAezZdWnRgLVQuX
uvRvucNfBs8Vpsqv84ZYBiDYA/nsqaXZBcUO82VqiQk4B9ZMi2J6fkgniIUBcVNwrYp0zYuZrttB
SO7zZu/H2LpHfV5KRT6xlJHECCF5q/YKDF2ecTrZ1i3483Upw55onq8TSeaW5UEin2ysymH1IWR2
sQ5KCVdGxtvvNqlkk0eOYCd6A96aLIkTn23rufA6+08nTFJoJ2K2YimMda3MXooSB21Z/6KwlMCs
OjqH2A0l73928rBaCzRTqkniL2uD3pc6Zs/4DetOnO6mo0OMhAQiwSS6FF4DdNMkbmtH2IWRzG/z
ZUsK37qkdtDNzPClNpwfGxtbFFc+Epckd9CngiO3+8505SdQNsy4Lr700WVb0tVmIF3tm49ixKmH
qCCf0FKk3rSs6FttIc9E29J4KKvHa3pi+4p3eJySbvgMBW0+rDh0uaO+UvRADuw3lme+K68b/kp4
NBQiCeRM26K8tZY9TalGio1Kn8mW/NA6hWOYW2mjSv6pzPGrfJgOGaYz+bsqJmpnB+bI4jf5Ydqv
u+9g7grBtO0YWPXhq6z3OaXJiImkRAHIg5LAfz76PJz83emdQBWOkgEsCnBwmOdNr/6unkyvJTEA
Q9BFmpumL9qOU7wsIa7ktieHOachkFQ6OhNcnj42DZ1JF0QzTG7i3/0HFaK328Ut61ACjqR0xFQA
28WJtIEFRHbvjGodH+B4PLrtB6DDiBu2wVlKa94ExfiA2DOudvdLPBaVQ4wDPFPVzL/2spy1r6xz
EaDYEbkuLh0byMJVrTez9H57HuSis4b7yhgLEBcBRQ4ymG7SKIGax+BkcK7A4ximAglLqP5B5L/+
c4jB7wUtwVN+x+gwPAJ9B6lMwZwl55QtkTc+lE0mxgb4867zC3mIAlRKIctFOKhWDRXg9/BVJOVr
CFo8lCQYtpzFAYDXGGAL79LKNNTEnJ1Lb45DmHk+1wuWJYUsDLw3yVh6R1lsP5QuwIppOpgSbgDI
vc+7mjOPgxidcLu5gzGcSQfRqSs447cJMUobtZ7R5bMWKnvHUUMICZYQgvLockGxhWPxhJK18ODe
eZ+fetHLDiynd9uItcxN4wxtwpidq0aUWkCfC7j21aqNNsgChJKzPm2sIhmVD9z6WuZWYIhOf/vz
aNARAMJLOYo2S+BdxS7UYIZEj1H76M60dd8gU5+df8f4eUhZtCSX83q7VE0Jh3rxhedKPH3TsBDP
0rj8XX1Xn07S9cn+BVk7LvD2Bo+3Y56MXZebAq2w1V9W9+Tx+p5NOvt9ml/ASYYfvThEtSu7er4w
/SlqV/fDqu3G+LTIWxOj9vJWtCAHKSKtYcLj/mu6NrH2h1hSeKkFevKv9Nbu/fwL+GFTMP5+2vUD
NVXHIiYftqfvqMqU5tP45rjdZU0gG9erN6WRcK9+Lxy8umnFm37uSGlysoetKW6Z5Og8MuJTO9AL
ig+QTWmHMvaKvosr/1Q2iIN1qmCYor/5QhL6AbDUhHjqUSZEhJY3BXUYdt1l+gOt+EaK5Z67siYs
1LKtjEIFazevNieJsIle8gmdenyWKg4jhBYnR8zrxyO0fc2NC6Jj2qhnXVF11A/1Jmohea5Vc/3L
ANMt+F4XcTVEKEa9U2uhE5V/UKpSbGo7KSmVgB4dWU2bA1y3faEVYrIC957H6ixKWdy+LNSwfCM8
dq5ThpBqKJixVF9q9V9nkJzRwb+WMZYlSHLdq6qmsfCgrRg9uBDBWZhYOFh89i2L7/632SUk4j8f
wEvG4I5M9knP0G7rXToPJVjUglCpZBlgDZYfwViI81DUeGDytWulvSdT6N+UrrjA799Lmx64tMsS
sAQHcZvEPRyCZjtfBQcPZg3f3yN4Ii5N0e1LLtm5wk6ld5Cx31RgajuwA3E9qgPBpycPhJ1+iNIw
JFBQ3s9KhKamLN1NhWKV083zaJvElxsvLudBeOoQOsvfDiuS9LggLipRSEOEDyaPOAiBCvBi/8+Y
c8XaJ2ZCtlQLaE+SacL/UOR3t/YQuj3dkzni4FVtfhfJOkM2UruOl4F06sEonHx5euT29CQKaHsJ
SNezcF3aTBWl+cIFFASfw4Uge0pAE702Iz3qOwK3duamKMdKoSSTJqBzyC3nunoAXETv8i/aW/Ed
bzzvVNXJvL3KNu3GFAfTroN77RiBycxoMUreRBN05zwaBNWkoTjsm5/LQKirXF8GsSmVwE7lR1Gv
I+cjBSE30kvR74yu1NoBKis0fhYzbA2MM6/4JZvQFTcISgB5qI2i3rt2GePQaIr/16bRhPeuBi6x
O0PQkiVxe1eJcYzUVbXoIVhk++wsiCdgcriL1JXJ8aBsEtoLJjr3mPDVFN811Vh5/XuuSUv7yfT5
dQ6Z/ysREc4RnhMYFLxxJA1j8zwvdMnLfJua//ETPpuuWCqG45gD+jB5AKK6iVZWbgbNBZ+VHK0l
z/kkjxQJm/Z1jasnd3Bt9h7LsgbK6/7W7Xbl4rOjhvIhTDsTBcPxuek8s5mG06jQ7r6WAA34zosA
4r90A1sZ6aLTwRR8UDYoQgJ1qrSBMXcEgftJAOhAL2qGjuQM83qluHZjOtldzmkcJeiFo1TwHoUW
UQ9HqLPpyghF+WtVinmm9WJzatOVrcVe8tRhsEFSQtkFw15isjWpQLDumQMzx56ubF8H6JOXC88l
auqb5xZNIK6XTQLxvPvOvBs1f1I2x18zILh8MD1bB5QAeQeKfGfes4aWKGHmmBIQzOH0LVB/2u0T
IViO0FXss+vZCoZsT/rKW1/Xe53aQy8fCGVf5LaWqaqJ1wzvXfkgejWNcjLrNBNUe/fOgu4PnXQ6
dYmOaYkdTOdfW0BxpFbKVpXNXh1s62b8DkPqnq5XEVUTAv1lYfUjXjgU/TTnDNdlHJIW+pY18vXN
1GlSlUizbg3wiIOacRf8f7nTNlXbZXXxFIWFMaBrktmA2BcUdQtzAeSS5Q6t0FJIF2Wm0ghc8VC4
tOoN21LWgUGd+7SSOA4FYmOICI4fMkLRguadzg4bCw6goAhnUEIMMUiBNT3KEfAmlxgREo/GgkQ6
xz6oSwzIhrRFZ3pDR9pm5I+S4pObGYD6YwZmT/Bh5T2qKamEZwh9TE/GIuTee1SHO7zOZPCd7kAp
Rm6ucHO1EdmF1AMT5cJQnKa40ixfwa6Myvi8mClUojeCQDLJWyWWlPTzHG8GMkFhNrVF3ARCZeWQ
sYpE9totlyyhepeXpiZJVEcpHYLX8oIKwygw3oRQjqwizTeR20NeODvCzWZKhMzTOBlODRP4koW8
+kTlmLJUHX3RHNj2CxxqAqAJpjhB+VSynO4ZX+IUCGZeNLzzWxbtNht4QuDfSHcnxFM8FPAcX+Qg
gFKAIPuzUetfyPvVnvE2mfZESh0cI8Q8yBwNeTllKUUCuEEk9U4b1ZwxdRJT4KQriCrGYDHeDU3m
t+Cc1IwpSML9CB53wf9ke59x1B3K7ubxNzY/yD5DxBjiaGlrw0c6b/iNZPZIHnY3APEFk3A6pTDv
DBjQ4J71xuUghcmG0RgDN2YZxYsDAxa9it+x6zJASIzUiIROFtYYzF/EtmBQfbMNCUfDi41498bn
HURtCeTVhMXwmxQKSjVcKPSSzgDWgzw1uxMGompxb6kvGYa5Erp6NP4vzzb2yWi2DcbP36TbhfGJ
FreIKUxdX4rmUnCfmidNrwcH5oF1/Xrdveyo/gyzdAMAGJDc8CbL7C7s+rRtgIukvEfKxdh4Exlc
VKGodqd0PAvfVdWN+NYS3KrEj7ZSsBwqM6l3OToyOGToD7ojG7xwIkPphBuXwU2pAILcN/N3rtNj
eZ30fGwq8nIWSnWAfvNAy6WYAm0yPVIFWpbI5iNZf0uUOp+s/p4G4UYLBGwgIHYaoowhnK2J2z7c
Z0vwCN28NcHCr1ucF9FQVRBqRStMCYvrCZQUguNEZ193K2QW0NUG0ZlwpMXrulVVvDhsSuZIVnev
71PTXjF16tAkdiWzDNjD3IvO+8WoPtBxghTT+dZvBYQ+JRwR1xi6AitGm/Ql/+lA7GKiVQG7V6LU
dRJcoGOXBcAWtPqAAK2hkhnTGeVSFTqM2c99HPhRClA4cEZV9wyjxHhqnNLZ3psjrL2be7EzE1Dv
HjT5ijvLF9vAyQshwvdisekoBtl1HoueEOkpZNyLePfweAAIBQw53Wp+fkJDBpQ4i+tbZ6RTKC/o
6553VuWfS0Tf65RO9h8sLiiPg+av1vUQC8Xc6PaJ2ZEplNavGFoQ+5t2xPhyfqs/dmz8dZzjsh61
9FQnxSfi3W86tjTrldGNeDXaUTmBUsi29HbWenGarJsHMH1gmd4MIgeqE7rnJstGfR2Ll/jiD/em
hmJA0UB5Eb3NfHUjZaxXac7fkjI1oqPsc1GfugrD3zfHPJrILs7dPjOi9LdcHq6Gb6KJfGv2bA74
YMDlhhEPWtWFq8qDFrm2fI289fr4nIPzTdsVBvl+fORnUfjLL6CWX9c6YziE1quVQxyjxsIAKNgI
FfW8D6DQz4rVXQMSxPhZwoqb7JwRTMgHN3iY1G1TWLpXjgVvVtLN6OjW6WqVxfBaPijZACE7gKOh
RVrZu4d405krfAdmkZHxa69NMsFtck4qXJd1oJZR1udos97AokX3DL3okCfJvIKhBSIqox4T4hTQ
84fJWIE9n0TJiDJzXiOJW+gSLBlkyrBf8F7n0EstQNQAw9CJABFiptykK2PwaKxvlewJ6vR/IcFC
cxyEzEyQ5tesUQt9ewNxwCg3DnIkbDocmPtRSsGA9uGzb7TbXXOmEnihRGLDXt1o4KBqHqjt7qT0
zl/l6u0XgBlqRpbkz/54m3gpBvo8dVc7oSaf0A40BfkQiXnlkMGQbbJQAMbrLK0A4uEuDCS5I9Q+
1eQbLTGS+IvD0lXmQLy5ZedMWXj3Uwml7j9YUgVw4S7sSGxJS+1OaB61YoLrl5XUfTmcUQGqIulj
Lz7UuAf0VhfAvk1OuS91BrmJ2yRFj3FOQzT/1dPBNAYD5/Itnd/9k4hHDalSFfmMHYHW6rVKmzGQ
ZBkQh1Ju+ORYaQCX8nlfNBOd5oSn3bL44mSa8e2JPzhGNHQJWS3zA1Qh4K1Oe5TKQYQzpBpe3kqw
4461cViUeWAfWsFaoIMM5hIBGWGcdkXDfgbyMIu+3FNlwWnthFClgvLlDI1YID7Qr1NWrfiD4XmQ
2566I4OvdVdC8XIlE00Fp0nCrv2sdKReqaGSqirC/pW53vWHAGz+t1xN2LKyEkr/uY60yszGRbF7
bkcsvQk5O74iXytNUXQHpL8ewu1Az7ehwo6+AHsw32LYh0pGmLLuN3uZUwO5z/NgYxPY2s9fGxGB
0fnH5bSz+KLadJtQzabk6aThrjOT6IhRVBPKMTw+N9tB9oS2lxCNg5XAQ08QV/Jxr/9q6R/9D634
wG8j9+V3O28+MzX4MxWXbWxKIUJGnnYf8nrvEd9dbz4W1zqhioxj1V4Zyqyla0TccJGJnKlNuDs+
WRCneYNUF0EcFrKkkUFjGh/aH2IJFhofkIaM5vEV26YbJG+VdTq87GF5xrRChh60i8dzYb0cdezD
8h+hbHo/ye8GwAcrZC5lzYgutczqm7TY7UA2EbE78wE/0Jq37HTxn0knIRNA/lWgrXvsf+v25fg+
0+TE+AkWZJL6/9puygDOR7KLdaaGIvn8hn0jxs6QIwHqqN9lc5mKGINlOsb1jJqKKEhyeyv5AE1X
yg+1b+5d+Afki7vQ5zPYc6BeeqD1J745xx7A+BtaaOaanx8bNLDSnF0535AtyJu+IMJ0wwHRYPh6
Ck9f9TyQR9j+nO0M7oq8h5JDyo2Z5xe4xBhPSjq9PLhXV+V8I9OQ0Sp3d6s+1+JcUeZgxDkZtHvX
GGi1eWUy2PN/PFpKAGIRSosASYDTpcTMZLJJMj9EfcV6qrR0ChdJPHWPmGEiDYp6elB5WQs/QDjF
rzUqfYtUJNHgefrML0yfPL02FkIZ7capulLiXeCxXT3+LCA5mm88ZVpTbNFNs7m/P1UNVuEIqiOg
7ao6OMPU7M4xwWCkDx3rfh81xOnXxMXA4vpE2nKmk5TChW+8XUM0zP6bZn5lAFTTFLGyDN4EgNgd
IBczE2QrhuUMIUXWDhEqxxYaEp3JJkGk6uwe5vdxOKv46dJITzEyb7TX9nLxl4l1FcTwdTJMtpBs
qKRkZwyUnpNaxcMx9iA5VfvaAkxvVEp6Vst/okL1Q2MQ3rqIHHugu9vwUtJ5tCXl/c9dvRpuxiNX
PWY+FeeAXortD+5CF+ufnJs1xI71euiKZdW6ds91drTdiONjpSeYc6qL3DoZwAOP5nErmiDDmrk1
MuMt/9WT+lbIajrpZnXdNfVmWFOeTWTWtyYgJNczh0IMjLlGlxSvjMbSnUUVoa44xAvREgMTwFgZ
pEkqgaBdOs54v/9OVPQ6zKq7FsVLsWYthtufSXcNgxml3D/kxaOsTBsPA5NTnDvay0usX5Dzy9Tx
bIuN0cxPZfi4QfQ9yn9s+BQdxX70f8vNyxpxY2KbheHO6MBbjb6zHusmzyLmMjxvSlS0BcOek/Vp
Eba9cFEXTtqdJ0E8/dZtjebmdbunNDEN3k2SqKZ8iN+pSJpYoV/PSVa0LMNwD7ph3LbPEx73yoox
zwjUaj01wMimVxNY9nAASMv9yOUvtqhZWfIwJkIDiPIAqB7jq/TkfsyH2SdeotJ48d/Pw9k1Hylm
6eJ2U18idqbZcgM//mDtcquNG2kC0+VLMX9yWkksWEdt2YYFwQIvv/eivSL39i/6sSh8ZPQj7aSW
vuK1Pbtjjd59FOS13iG/XhFdEoftlpIemHxI1DbjgxawAVZgPfE9UZVzuK0YCDgiaeAb3sffs7fe
p51pbAIXysZsO4N7te3QjtdUC/IOZXpmKSV0Gt4CO06MaB1PEFWnJQ416ObbioE5a1kozyAVYLbp
JTfe/TriKdtd7z2RWcAvls89QzhbrR1zLXpTLWFR7tvYbJpFhFEZ8h95BQPsfBs8drhZcQtFRmqQ
gqBT0n2ZD8+jd2CugTjsxBiirlI/mg3jn3ri1DItnTLD0QsW/P5VWmWbuLczVIgAZNpB6FhyXDt4
jo0oevaPt0gv8NOPUPOeaKO63F2BELhzVFOmWBskWVSDC8YqUQb1YXVGdeEtJFkhaXX1XKF7GiGc
7JEAwsdJItQUoDBBD5+wsq6BNU0czGuUAFd8CJ06XP3i/2rCVuJoriM0PWgtkNl8vvHYYlMoWg9d
PfbNJCeKVq6Brnh1rR3XxVH6uDGa47DFV0matc99cwsQwmfNFPp8Ab7cwwhhlf2dJpO575Z+DB2t
La15KmNN9FMNv1E01jn95vkq67/2IU7NztdGCguTCpTDMmrhMspDq1cOH/y8sIadAFSH/O/XmNsO
/lZQ3k9dK6QCAzO0zc9lGewlJX4OISztWf8nNx5HEL4zhL8JbCHRpuxhsGzG+/AIq5bL4O5hGQ83
yKj8Dk2V7q4PSswixFCY3b7PCDkAy11LUkz+5z3eJHsdMtCAhXkg7RZGRSxYPZFhv6UGUjYvkM5Q
/dIyI1MxAHeOTjvK13SrK7CHRi/mr/+FAWm1IJJ7M1CJzfBf/qX2b4iEbF+4VD9SKiIXpbOxi8Dv
gbduN9lYP9dr9BH7kfD3m6+MLAS8WU16pwC6gnOdnK10Nn1gVsTTdeiQqkKDCO5eNgYmJfxR0Gg/
hRUHPtSamU1Pgcoz79Cs76vS8IrpiqNtcBTU85ncmTYhDPRvyW1Fc1PSNOdolpABJ5Rn9ePPsits
6EhxtkFbjAwMQXMv5PCkBpeaztDqfWbVx1fnyMfLKpRyOUexYpORx+niCF9lt27F6w11D23pC+hv
TbE8D2dgaySkTkHItUs+zR2Pgi9L0Rv1AiU4IwtRGO25X0tQNSLIzksCmzCEG+Ay3MbrsStFX5TD
jK+A1Rm0Hpzh9DJSs8sl0+bUOXfZ0uNxXgcoDJu0UJlqqsLLNEWaY5adtBRlRejIvRcx1PNhOPfa
0pCptAI4NR2hx5zHXt5ruxzQjx7/LaVGTrKZtdDzttqoU+C22gFW4e0Bo4s6Ru6xQQxJKFsZCjI/
sMvSnWA/EXOgCw8jLLl8lEYkbOJyGZTs9/9SLu4ilCsvZN0RmnUjzyMWF5TylS26QaF32Al0soNF
msSoo079d/EEqoOARWkitTmCBt/bcrYVr39ax/IQtYBQVPQF9BN0iVU9sLuc4OBUY0XVAudugNyU
/+e5d5fBSaeusibhVY7eR20F4rhgGrDVYJx4ok3hfgfJ7SUgZlXTZN73Kj0rrSm4FtaaQ1MWLMyW
SBLSKBpyGa/dC0Pc2A0evG7j1B5SzF6hT6OhUpfEMbVlasf9Dq8LMgH3n10rKgc1AJapybMenH8D
pGByl7U4ywv5Hc6VOah+6XkWu0oVThPkWFscxtHnvNoR2LQErq0pOQ5KnME3B3O3wNOruNUxZK89
4TpNA65T9gNNeIZZu88C83VmDkI3H2S33kih8C5NC0vLfdrD8L/XgUgsQ2gVDceq9wgjyEU0j9qM
cyGTHsERuu5kNci7W3KZxEQZXobfdyV1d7Tn/SZJaj2c6RVkt6hpCb5RX7k3LX/V18I3KES8Qvlc
kefV7fGYtZcDLP84Pu+c8/+PjX7V12x0mKwbM7CMaZVMdKXRe829L68g3fixADP19HXU9UovNgUC
NliLFY91QXKQhso5gq7fqYyIYyYHSRWHLUAXnG8xsjP2pM1kkV5U+R1T3EXHauZ9OGQ+R4EjUIqz
vEnsFK/95xYYLRjCTC7Tuz6Q3oi/3ARMGfMtO9zGBKPAYhdBV4ourfn5v8pDxQMhgMvHIgOd4hFO
Nw/oNr2Rz8O/zg36Gm7pKJ1aXleV+A6i+f9Tk+mmXUqK7Cl0xRO0DyaJr4sn9WqDvLYj1uZr3fpu
7Okw+aVp3cWcOFwrk+v03nL6Dx9pFdMTpzIg7zLTFdiCpFTesVDThzNlM2srElU9EybWG7xSpt5e
EnpBi58t9VePpK/ZZa4aNeFN/txX81Tvu9Ed6NTeyM9vGbWtTp6So2hwqGlFlZMKecYK4fS/4JXX
yLsAlB2Pk7OYvsO3WMilQwdOW7MdSOPrKl5b4Oc/5cmY3KeWbLm14b3t8yz0f3X0fX6QRU05PqNO
iNTi1usd1dEu9JZy9qB/DUCEZGSLkngr4ms3SgGWDHtI94A/U7FKhj8Svt8BEx+CSjjBS4nfSfb1
xXQp1vbFV0O05XCuRcMeh7l6um33VmDoTgLux0vnScsA0vKVR1hDFxCgO/HpWBiA2kjXL7Zex68T
lJSD71rBF45rHIUVAtOHqSjrcF5lYlHTw74Myz9WgdTnBKAhTaaMqWTwSnu7h2Rac7WhwWcLstJu
GVYaxN/zsO4GlTTGWAaX22U0h9BLW8JSkQT19x+9E0BA5oM4zK7XcOJAnLtJmN+FCnk86jrr74Gu
nR1lzKpgxIlBK/9aUlZeRsWS+YYpFRRLYiTpqIX4B7z9x9Sie4HqEZR+DwjvASsmeFkCYuR3Nyo8
dSrsC/7zXmEY8ev6YbwHojO6D1eP5fCq4t3DbHIUgmO8lcK7SqUtocU2KMBwYuIf5ktqx29qP67C
1POwNPp/izMdbx4gFR+SbYx+splUQWYc6roH3Z7RzEj1YkKRR2aB1nkBneEHg7OgcN4+vmBO0Iwf
QXFE0skws8s/h3xqkN1BGyRtTt7SwwYQ3pCKVV4w+Xo5dnhODmw0rWgVwbQ5oYVemAvUNz/VIX8y
yD0neYkW/nAU5CY1Qxn5UKHe36maxRSERV0R/Bg75dvIOBLYr44g+PpO6MNOmNk+UYF4urp/e46N
bjHZfGN6lTUT4r369CaQSWP0ITc7t14oUAVieoAMTx98CgX3fwmNLfBiWPXMXr5rQrMNnODUjb1q
a+ATQ4CkwZbvy11AUcfl1f9JBPqAAa727aEiA4nSJg0wqu9hkFBDyi/zbUzczsQjD7flr5Iha1jz
T/TMtoDjXPxLzs8bKbiqdPo3IQF9ZgxBlminbBpiXNKd6/7ZXnOXouy0Mn+Dce8n8wBqi+aiUSlI
ToX7MqG8lF4uyGkce7g2GBoJlJna/y7UFGumoOB+DgoekOxwoLAAOlo09Y1SjPuz/gSrHbJBIm3D
O+WI5hIBMPflYfaW9AnIyApWHZMjIXOain3fEglWnefS4pN0eiFMdcRs+SnWUmzdh74WnKOXY4i6
3lUrB1LLtbqSvnVedCwc4InpqTfFCgv7sGkWA+DEspKuhv39V7JjsBoHm5BHTW9po9B0fycziugs
blPIkTXQkKRi+N8LRdnPt9OLpmcWUANhv8hpPHNG/GcMTLO57s8Xo+SOSp3b714Xm7zuXfEZTJlZ
0i9sCjxK/Uc+gAV967MLXVL70EF7+K/puCo9y2Yn8d0T3Wsux6xHIRF8D5JKYKiQ9k4ewO7TsLRp
4/eHFm3NRQOqPHqulocMjhq373o8DHPeNzzTXWrQ5R6RJcBSlGAgR08de5PYxAsD10a96EdIHLQi
oy/GdS05o7J23KX3DAjthz5ulFlTD4nAlNN/gcEX0lkOxqLV4AqEI+fB/ctqn5fn5yNTO6vD9JMc
6RaIYM3jA3nWPx73VWeBnhGpTCYvwS/op2tWkBDsaClZ+lRzNJbkfS2MQsr7du0J4Gg5XNc5oT7E
0MqlVDeAeXH410w7vtz6NhKMpbSIhQdKnJnMjy9VhwVege3nJgH56aBccvuqQoo9cTKW4CDgUgMK
TkXQ/sVvxqg5x9wesxUZf6Pjd37OBFM/G1oNCOLaNrWcuj5WvkP9glR+bI6YApsKXh75hAFdUmx8
PpKBGzPnfte0E6mQ5Up00qPu8BgAvgXbKCzFnUjo8th2kKyu8gjUOFXScDNHaa1sDpSVI/N5uiFD
/aOlo5yIWwkCqO5Q973VEOcd3teC3X3RjH/8nbkiL9hrnm5iPbw8KkBRjwkzS3b7UeQAG+e82DU8
Wi1sUTRHToQFi2TaaAPt3N5oX/eXJhOoZBBTm0DisRx1tT+Vhhn6ii7zkslH0IZmK3An/XfCE1xT
Ms9bePo+N/960wWCDSwPiK/t+Hx0+ZYc8gxFoYAKFuS3sgee9Cjs3lHzunFo5qaznr/fTMt6/dvN
Zhx5UoN/0F9UA17wNJUsE9ufJpuXnDy15AyG6SvcMx75HnfpWDRlxAQj67KoqNcJlJ6eoKYjpy+Q
GcQJkfF7/iYqspMFDr3yFDQ+BH2zcvyIQOlI3VSc3bD0u03UvcxNo8LVJ62Pa3l3BKafX+Bg1fNL
fRau7cJXmBRE/vWO6UKlP2RNOXqwjSpzzV5fn2LVkiSpqyvu6tNK6wZf2jTLNQVV2BmKcfs4xxcg
pG2GFO0Eien6w6fwFa2+199Xa7Aro1dPLqvRSliA3N3+1eilbwLopweuhJT7SPcLSAsnbTUj9mCq
H4tXOEOQbJe0sJoRU0yd+efY5Ewx/n5XEDVDhnVHkNxhdfBmT1jf7Fdb/HjiULItRtbI8QU+2QPN
ZzE4E2rQA6Dq+uKMdbb0E6V061gD40FPc82jXJytBqcfbF9jZVNH3b5eFOkDgtieucQGqHj7ePyR
H4UKFUUcrMIuS0ATqGA0/gHaICvGhBSABv5iy90cWD+KU3pAgwRXOYn8HIjjl5QIago2yl11GkYL
ewjcU+ZWUFZidV8eiais9/LhxdkhAznmuddTpV64VfHW4NVOPp7cnqoVcdD0A4UDE5HwDrZgCPMm
YJVJ/5fLjRooVUBKwLgfsnwKCejGfjbtjsA2hCh+2369HKp4g+45VpoNtnm9i3F/ri2DxyfhC4Op
NDvRW0gKShcS10MxOQLCiSSlKdL77lt/0NsUs17AOfEJ/1/rtZqZRTdkmUDiKjFOzyCOh6lyHbBy
8K7j12HaMgxcDM3csbumonCK35cO3zm8zD7ezwNeSpnffovHCivN53mstqVob2/HwWeO9mwHhrJe
ZRLKNVAoEXNfLfGhDvZcmTT797k+kRh/DM1k1tzg0erBLIYWn/OniOyHU+3Z/MH6r7xKqTk3OfFO
jMnOldaR5Iz08SYpuN4haloJ7Z3yivrcc+vNIAAgsOGKhhrzVFqcxJrqGMN8eIVbgtHcwi8ukBWq
OI/0kQ8NqRBrrIOIMQ6ZJu+634k0oOzg/gWVLqClkSDhC4QCkWzVovxOcLdRE/Sx8K5vkipYR4dh
/vRdU1buL3mlvrbkwlZYIAcsrzsv0gdfl8Ix04zX/PsO2sdOFeyKdymUYQM1K1vgfQncF+od3p6h
eKaJhcjjPCdw5qc6XRNqM3CErdaqizBYTFWKCW5KjDfRP/6kFvzjO3dDZQRhzJ/Iy7Ixj2pbnY4P
qfWBh+3ljjhjGrMcmnASSiIHsFuVX02b13DFkE8P33FMZe7G3/2FmeXlzIZSBNVDBtC63cSlm+uF
aurnEJEcOjWHee6nWymJJJTM9T9+hGDqWx4N1y2Ih8+PgI6QxTEatDxaEVeon19qodvN1byhwjPs
44xJpkpw/dycoYgt5tz9GNXeZOaVpj1WVqXhbmtREbz14ZW53X56kcMUkfvqFfpQz58Gcj6Lw7Tb
Qeast7jGvbz0qG2Tlb0N5aQadx4Wwdc5pKKtOyi9PHGEea3y0YXSllkl3fWzjIBWbWbJbGbvXj4r
uMaMouEtIWfl/gJeYqe55D9qXzh3L0vSkHPSzpBS8D7iRSRzQn82+jaXol4IMu0KbWJegEiKvBjz
xUGuF4gD7X4K7dN2QeHmOofFVsd5plHSugdiq+wIw3Q5kZt/7sX+3KXgjG9jU6tRJzT4v1DEa/Z6
81px7/n4iwd6KEyfkMMNMLOT6AF9VwwySAH+P4UCWOQvpt24/kdxmjH9Em0sMbvZXX7V1TnnWDqP
cmkK00F2Uj/dE+9b40qunX0jsuiV7YaU8N1U1IvSqMYqMltT6Bl2jO+nfBbgJMVSY9lEv/53uOrW
vDFbWtIUwpynKsxZXmvKb0aYw1Cks07ppc8buG4YLamnZkj3G3i5RPuYSxXS2JcXFWcjmBsnHvb8
CrOh0Zb+hQC6RNE458BeEYEdfKuqLhKcwQXtUtMPYgDFAnGzJObqFIqgs6o4cHTR28qXxidgl0sN
/YyxxGP1Y8yFxf53CIXjkLKwxUZrOnVE7LfsY/iImOS9Rhlm1h5TbDneGkC58ASE0TgCl8gBHUZM
WhvhB+kNPAMtdaceKrPA8R/Ik3HzwOSpUaJQ8KCmHrwS2rjLI8cH7DqNpPsI9XUpB8VNVPCnc3N/
wEUrklBx0WzmySbrBlNrnmpfyHBC9uLFxF+LblpzLOhgCfsvILfTGKd1SCl8sAytJAcmoDu7xVUs
iAMdRS3BCpKci3mI9LAeQSh3sZ8Jykk434FpNWyELKTbilzRaKYqFSmyGiE3+n2h8xQjU1m+5kwX
f28FS2UHhDta3iPUahCHtNLOLleB6BYe2NGu9Ia3n63F1Vigt29p3/NvlD3/jPLxX13JQtzz4IZM
phy1OK5AoxHgRy8Qi9gVbFoljDlMhwOSEmATIRl0Wy0q8ZYrpVpL1velNjbBbzsx4d8Xsijk94uv
ekBSeGMABcs4pKqdIyQVJIIuqaY6+92fg9nofzh4A9mJ11BzKGkWVAV42FRUqRsyTlv6iqoPWxqf
aYvJ09kc/ptwU+RJYdtkn1pRlqU4pcFB8lopg9Z6TRuNzWBFteaIQm2oUCgDz610MuZznump3qju
GERXElZdECe26ho6BhxcUUimuOpJ6zwzXLc2FFJkYsxgYn9McHxpcVOW6NhSl4irr5+a08AfsfYT
ul5VhfRXLadbSKaYq3otIFpuSWmnHQvLCHhxg9Q3L9YQnLNh/NBB2R9gRPDJjZActUswtZYJAVmL
G4WpOqDYtR816y1Jtoq440o2S/C1X8ZFMt/zrK1L6HTCkDqwF+rt9ok/HGERINnDYcyh4M1ghmH3
YJpNm4mr5nqhxxh83HUDNWShh6grlfhMRQZ+uVuSk+DvZqmYBZujnUcKG4yDQ1YIEbiG6y6SOjjY
r1ems25B120c6TjngRZQfzs6aPTY34S5yzYtpkmLMdtQdD9GF88aiCZu2GmI6olUWaXqAPpPwCmi
8+5gAYSBlXdMLgIqOxYeMicDSBkGj0BBmKjKkScDO7ddkoXywnXuMc2LBLJ4N2GijeKRp1SNs7ex
qipybNFIVLv1V6jTWn+bqbVPSwrkC2O4mHLUvr2bMK6Q4qRpZS6ODELxHzm90TlMWTjmOxpZvflj
qtpCJ5KrTTEzKK2yTzClSSKfJzB5Ol9mFVLTK44a9e0kqGvMsLFddQLE9+A+AKKuXcOMEVExOFg8
Kg5MRnuymIycomnIek0FlIMrMdK3AwniT8IzwelmE5mQtX98QjAvCxdoVjkRDqW2E2isAshUKwgp
6wM1B+gRdRJvpqEZJqPlBeIDCTTOYk46yl2sP61+28xpOB3Bsy6akbKJ45g6xhPTrvsn3tWex3po
+bzLoM9cB1f3zYoPoEl7OSYHdSdXq0eli2evAE6q2C5ikASRYk8SaqkQBNgxtJ5+YK43niaW2I26
UGUJARMT8bjv+3rvYYqrvWCFNWsNA/9EW7ue/QfMKz0rgPy6P3BKIq4wvE0SnLVGZWd295m0W4nc
KSRz2xk4R0j3k3nLSgweauwt9acCKm55mZMn3meXs73MJUktE2WaP1kGGXMcArRbxULymJW7l4m1
O4Eib/08Rh1GUw+8kWxWF2qn8guUOImqNHczYcDiQc0H2SpQj8WanoyocQA9TWOdL8ocp5lmfaKT
XxbWAmeHj/0xk6qx2+tNeKSMrwTc8D5F8Kr3XWjJ43p2KynfJITPDzzffe+s9om8gsvllASX+HKm
deVYkvvqZsjFtBZZ72mgEPqCqWrXeaJ6fhO38I1v8YB56+pSGgZap468wxBlKD3DrflUL/QA+5Rs
oWhjHrMuRRSoTdlsVjWBfCo1JidRyKh5kWj03CcKho/PQufcCCq5WJ7tiIX2+zeFHGNb24qjDxpx
rixy+Czwwea8IZ06vGq/xUorKKtomdD0nqgQuvYrrBqTy0q0B53rJnH4Bz3JW+UtVcFYkji9k+oJ
5dTWgH00so7mD42SJId3HDafs+Y7LwSlEWn7uneWAGD/WP390qbAQqfVvXdxPjE2cgxDjWf3mYi2
qP0gVICS9QIbEJK8Wv+wZiH8+NFySzrORTdiZd2hmcQsVOHgb7t+6DEJ6oSafXRAzjr3tzI96rVd
JeH7+VWG//NLlLxpvva0YahOxYrUnnq/0b0ZA5K30eNxjLiyqL0FqlLLRlZIa25OA0VaSPwm1EdG
BEyRG6d1WVz/Ob3qEzp3G5LZdttx2KIj3TAxF7fmljbQ1lr4ONyT0ujPfiiwBQWFu3FikmvodLOV
tU9FqBdPXOYx51hBCL6sC9jiWlH8++epPI6NRXvNxM3uo8N+ybXi+Mf3OQ9DHuSrWg7KcoLIyRDA
3s5PX8zBELammopsh7Ei5BbdcBN2E78/sQGm02i+4DUY/njp+NLgvF/s44/dSUM7qLjv/ublqqDY
tmpyo8rdc0z2QvsrxfjDnJDz9W+OPro7Tg5STdyKCGowhKgS8Zgz2zDIOeowvWR4mELziaXST+pJ
PQb0PO1hvenRLCi3r4XzYrDIweb06ozr4XuPgXfV5i8/XsAFWKlxn+YEgpYE8yrc5HA+d/YHnJKN
ilV0fI8xmYXfpXKyCwLrV4ofNfde0H6qvubUMfL3FIxooTJfrVYND5gHWaYotLFZY+uqShO7njy5
RZ8Aruu/UOYVriK7QUREuoTJk7aK4iHeoFpd4XDvZ5jqtp1u+Jbbnpw9F+6Sz1fepGL426mbGnMd
t2Vf+9MdiyCh/mPw5CiGo3hEJFDg52i75JaRhRMtZXYdXh5PVSXVzbhh4WzBSq0QGtu/jPRLC27U
MCcPCJIyWfe0r6lOBI4bBV2soxNhIWQtJ6uXaTJ4xiHjvbB0t9ewp8u8R6LBLXuDsmuAOWUiyEHR
bsmEMAt+Vl3gYKmCpzHCCM7M1kekzBUXeK5Eah+14YDfiuPgN+mFLt4WKAL1aw2bJ+6MkIQkA9bB
0A0dj5q3+zly+zBiM7fBwXEU1TRO4KWismlYWmYuiEg0kV8eTWl2HtA1d516os3vyPZU23HyFSL2
IKsvHsgE2g84FwxjjsKEs5el2uBhtzmluV9wrwgyC5HRGQqavG5k4LkvYOP6U+KJAdu+XXSW9FAJ
0GkC0daUvNm1bJ3Cafpb1+UKHfG/WMbeIQhe8U2WbOqTBh5HIz/XGOf062PkMjoMlc2t66vauEPC
sUXr9wvn1J4u31IAkgKmUsAUuGVimcIHCE9IZdsMxbiWOdgAhCIZAJxKkpaTKuTnoxAhNdfnMm4i
8LIeMaihR7cmn3Sn0E3iKWn1fV/fxh3SomyLjfA3AevQZhA0rqCKPPs+SEWs7Ml7sdr/gRaX4EEN
baNGpSreJ7418qobstWmV+h8SX3CiYsGPxptGZxJVrg0peyxcoHcgy99Vf5qylrIt1NM/XV0VtgY
JrMZbwEIoaDKUWQae8OmxN4NWhiFbgCEbD7izpZRRGnTx5aJKaCWoMm4AVNhpY076Yv1DKj6v3XN
jDVQR30md8p4vfUch6kIofkvLMi10QxaC+Zv9UkA1IUDC+QXMma9xIjKbNaWtq9KP8vzmBmtyy0X
G5UG7cFRmajwmQ3ow+u5eKF9iTwCY4ALjtn/wlTVGUqcJgwVNQqFKSs+tQcQbjH5gm2UN6JJbnq7
qKDI1h9Co/UcMvKIDAgU4+WAyysa6B+DwnKGlUMkSqRBlUchy/YNYCra19xEDIi/MqoenFn9NrL3
PApthKiRiBtFgAw5OskufaSJtKzwC1v3PFrnjesuaTfaiHCMY9knYObfIIDx84V2/5wRMILiqI7J
UHCJsbLLygv9EtzLIHtX6bjE1Fgv39LVgIvMNLc1qy/5s59wqEEqNHjZhgtG4EScmTmO6/rkcoig
Jrfg9RVBEwUda9fcrOundyQoPFWUOFpcV5EOcRxB+gko7IWf9NGVGRSu1ZweZs84W+dz85uKgxoM
OK1kXEsSdCJPhjeYCWt7Jyh7CDiZj8lHx6qjJrO+rvSWN8U+b4nB0rk04SmWCcqESK6081td1Ao0
aW8jBmf9FevOHuobtwZ3N0+0TV5baYAvecNeBfi5V7tM0RRw/GRzXcO9DMow+651+FxTOeblF8fZ
lIHewsYXvHpnnQySRkVZtoT5C7n6hqt9AbTZrEOw1U0GNYzS+oadxMt02XhSrtfHt5Jp54zMjLDQ
+HrAHftEkVTQ6mh6z2gFM+vpfGD/bTfXY9N9XFlNdX872WXAn4T/F21X6Z4XidBR2t3wPaNDi18O
0ep/ObFe5ry7KRT4CCuQOtBjW8XBIte+cNjo0WLs9CM+/lwLZcmswu8BXiIEJPt+yBmIw45JdjnR
XpfAHSI6FKcKNsOhxPV73KLAz0ZPW2ODbAGwzWHs1Gd050hMJecIgA6f49OyYl3/PKxIA9SCUVq6
PZp9R2UubdI+fhJR9b1u0Za2xh+U8QLY1ryXkgX8q1jeZz1xURfEPn9159KPFWi0inKVWbQgp2O/
j/xFaq3OUKLlu2WIMpEg6wZZH0akIVA5f5E+RfKKWXtohtS/px6z0wK9ds/p7wHWbniCRyAPTZAg
l1mNKSKIMHtTg417FuztcSUJjShs2Nnh+vNqMTkwB1Dmt7GtBLl9XIx+liTWY+SM3LdscdJo0dc1
oByIYDGeMWjdDWfYkS5jBk56PczyMpsLYOziRO1UJC09QdJz1S9W+zejUyrjHJf74DQL4Sjk+jfM
UsHeVJNLXFTdTU3aHq/TrJB6dJBzn9wn187LFbTMHNUq+vOrVwYiRqPJfSft61yD7rtDKTlQrF5a
UrvpDz9uUXIlEhzqWzPuE7CazCnNv5ItDKmf1tLwkgQCwKd1H/pmA1JfUREjvYcBbFAWooo/tVzd
qoThqhXuGazDnVTrsic2GWSkglX/GY1VqRAoIDOP3MMZK+L16+o9ujy95YCdKocnWPM6Pd6/iKj/
98+RN6Ce3dYKxGVAhvRdrgAWUyNmMUeZfSbVw2lGEX5LhIXwrEa1qN3eENvI4cvw/mabCmrC6GqN
c/xr1oHnmhLGujABOY27MrQAtgWtcs3y0Ny6nF6rucC9QpIdc4Q7+OWXZ8DuB+HPL3P2AqMXf77W
vFnmG32Sj0kgDezHRoAhSDPbmTAjAbFCJdciIMg6xavTJ2dMWW+lgO/dBF8e0xnGm+goQV9k7lgq
XgEZ9J7e/qFov2Ex6pCDzWaD1pH9H68zF5AZGM7Pnp47hHWrtcyptTMG9mOwGezdewxn4ctnylxl
/uBhI1duIHyK/2Z8RojO4Y3e+LtULrIaJGc5rWH1ChMStd7MF/41zjUqwKWkjnhpQ8ySa4J3iwn+
+p27CS7Y6lygiZC+/sRtjnAdyW9EIg86gabjPvISXYz9hxh6Mbg9AHE3qMbUiGDmNMQeo/I90ZUv
MU/AaQ16mY3LTjU4eZhM0S6H/Rcb/z8OhIQtNYVvUhvQsKe4+Q8iG0PBFKzAMQUIPO+Pq9qvxHj0
ySt2IxqhJ48joroAdKwiQUeIyK790yIxYg8jZID7Qun1q+ksaYVDYadTAx9xkTKicSn6Kyzx2Rlk
/hNNU9rJFJj9QzAHoEWBMdygLBI2m+CaQFjEnrsH3U7At2p8SGie08+j4cewguLkeytB89DQLlPZ
V2w+ZnnsXnLe4eYRE1jAJPOFGGp7sN2I6GlRAUENhWwWwaA+oFi7Xiopvmy2wKBovj/8rcx0bh+i
zvG+Qg26XDhis7baJVwhhyAJykRlIscHCz+yd+/kAi0w5cLhhlNrQ86Iv8Nd7YFL4RnvzRhW3Buy
vozL+9x78gY8V/XA3p7+3mfCt1doxQHxsmLK6BBrfBUqx58gQJ0qQd1l9TPI6u3p1zsk1O7kSgok
qmDuogVaJ1KjamVic3DRhXTu4MioNPNp8JZ1Mo/NVOibJ6wK+dZCiG94gjJrBTcZ2rb6ts5Lmw3E
5Z4hthJFkGiao4dhzHCk/QzH6lcMThx74xU7Lx6G40lzip4Z0zd3WIlhsrTeZtrsFcH2dwnAMPNs
nw5VqYkENvYW0weqicUEmcDY01cfgqVeevtTYXEqzcA62diLFtFLMabUsSEmdGHwgIfSwzRTN3n3
u42KSazWozt+wJSQfum8aY1fTBjWdBOv3V219X8fEg++D6NG3NachqjhIPeD2yuo6l/LQcG9AG//
GovOrkcVofK56V40SgB//6nD5T5Su0WmgVKG2f5lhSU3CFLuIwuxd2EsgGx+EU4d0aVgs/eixaD/
MMoJ0oDzR/+WRK/JnoC5qYctcG2rMk0tCs0L40TEtXNFsOp57FPDECH4PcpvyfZmQpqU4Ffs5Q8k
lMo9EtpCksJ9dKoMLGHjyWh2ZhX8X37Dcsg9U2sD+FCg5hLDFKiRTzIkmRD018IIkX2xBu1wLpub
LlOd/tmn2jrTNwd86WUXZULaidZM8pVsx2vAVprp6dxcVlqU+2WfwtFz1LBTg1eQHHbj6v2Kr2+5
7VyFvTB9c3VIQg3LRvTH4YH97BRxsqxJAzLaaWwh/BYIqBQVRNWKfo8smvqEKL59DEW1GBaxQCe4
TsRPG+xhltIqoYKxxv532Qnf6VotqILEqmKsZlW07gpEqwVpyAWz2dxxNcSTPg827lYtSs2f6vZR
G4tmUcoHx5zgjG71u3LvVDj2gChxYt2twMM2sJuf10S8Y60MD8kiNoPP5Ko69umEThg6YSpUsHpt
n2XFmbJskifPrfn2sB+fdcQs6a7bsOqzOjKWTsVMq8jB/4Uu/MDrWPAnHPxdqcyQKnqVAaVT2UTX
8UOmsT3PgKdoLi2Lj4fCmRgZDiBNB7mPb7clcMCj1SXkAceUiwHIIFKoc5nBCLektM+7Yu6e4Fb7
bIsWtpUjmIwc/8WN/BRdfAPRjyEglZl+i6rGqkQQBZaIRRM6PmI+5Its2lTnLCfZYFbFbYUqyQ+O
GYyAwLpFNy0aShXH7S2PCs0CsM3eAI0a8osQz9USlLvGjcZljDCvH6Nxrr9q9BJWeQNinzvy4LuO
ACU6kwQPHzhl7HBOL9slJmaBl5plDC7DVzq/D/Csykwjllrrk8JsdjXXBSuwIMQytu5HU6Rt1FxQ
t+2yNT+gWcdMEP/8h2jQ9QPM7qVte+363f7qj4Z64cBX7MzLkLkGcq4eXmMjFJybjeTKpCB0kFQ8
Q7TjmrJt2agzTvhIJMW210cLEW7OSNyKKqtrsHXEg68LJcIUeOZt5yOBjbCMcdGhumM4DQsOj6r+
Wg1O2Fh4l2B1tSVKKD6RWVoB8kU44WvdyNHS1VMjylARHaOZnnbz8dwpF/3KOkHpkpNg4dsy37qM
4co0rs4c/hl5OX1r05Z7CbbgpOgPKy3qklnX8c0ZSx6WKo94jgsX0Lk0XWchS3rRB1AAphL+i0Km
pQgy4RP509OtDpb+9p85wC3gU3dvv+3J7mq35q+zntynEtNkp3ESfwLu/5VPEAS8Qq1N5vTOixcn
mnngpgbOjRu5cxXg5caUpxC4gSqZLUihee80TyQ+jjK56sV7jDLvxbeRrMjuinpV5iTgqC0wO/dR
G+l8X19TyXxFWbeUIgygVdEQmDvfzrI4blll07E28qfzAVtW6Jm8VNlx5hwgN0+eYWIKR7RAKbAZ
Fbu0+I0jXPFm4QQC6q5tIGykZfEnHt3k6yhodUWjDZ4zvUSJBcXeZYONzsrC1EXh3+YgkVrJtqK0
Nhr7baUdcDLK+vb2L9S+y6v8I/ebAx4w/+R1hewlC5U842fydkRBFgoPCC85Y1CkIgSWdaGoTTJQ
zL8kUDJhpn98rFYtfh/O2IKPuy5DUSJlIk7XNbqtVr0g0b7qF349mO1fNqhnqxO5q1pVSSmCGYmS
PIWrJMOS1ANA/N1DkU7zpncdQF0/pjsY3w/7YylP4LOF0CFSM8NMJ7yTQz19PgH3RLRhOgKA+d2W
eDFRztwbLYslg0HDEDRy0wmqsNjhaGBYHV3N914CEq0OaT12S3+UPONPKRgWayAThwGhJ4prl2hn
uAcdt0e5ko925sw+TZfdf9Kqhs/EVlf6ZyDpk0/nDIc5dJkwMdYFfBwYBfIz+KnTTB6MOQTk0qJD
UpJ2yz1TyIl5VoCOFDnRnyRGgNkMaPQ8Dqo4Lnfqw9d4eLSuMkJkvWMW6zk/G95QvzMq8rB4pwS8
jLggA8Q+yxH8V5fRvKENMe0ulTzOA3qto/9cKpfIGR0M8lpHfsBqY8Kh6gVYaOZClayG9f3CBt1M
KNSLE9bQKy8kQsNTzXnZqSMLMoRwdLo1kDh0uH0DSwDoWSkpqvba/PXtlhL1Mq/j1kb3SiK105QL
l5b0eQH+0sOowJv06AHsaCRaw0jDV5wR8aOvQwWwbvhadb49yjLKVJCYgdOAyiyglPwT7A9KhtKe
kUpThHaH7lsRv8VDBAGdmu2JJRjKyawtMHuQrFe1PDI1s19rGcaq1mrVCVN93BHShy3iVzByqcV4
9vvO/U0TfqvNizP+25c8f/CxdAzlW/I5UyR9wDAI1uqGIRdonSJvovHgA3V0ekbBfJVBn1TcKB5J
7HyXI8plokdqwkDy09QZ98IyPPJTidA84QbY77TLmHxhU8EtJBqjLdVeD9W/TYTwK7m4EoXzncRN
luza9IliFs9Y1JHfrp6d6xWY1zLzhWu/+ntzCfxqrAA0hQmUD6ci3u1W6aRtlFE7NSTZo+0MaGuG
fulCS8VQWk4vF48cYH2oFQs0UTQTsI+DEJA6Ns+sslEN9RZmDOS8D8IT1WRK53WUfZVoYaofaxRy
pikCblGiNaKte8ZFWQnV/2GrKVLaa3DmqZF9iDHAOTuPHP4CRM7lKSU2nDwVn9vHqnA42HjD5Bnx
kodDhM50d6PT3L/knGUCgWy02Qfy9W3OQdXZpdNVuXr5saE79U7oEmvZNDoJg6a9BPHiB2kqtvD6
Im6de4g1m+5b6BvJaPLRk/wNgMgiLasis26QeX9DeNlqpKyo4iXxbBJvtSFJOaQB2wrtpyRwIETJ
Oz/0vcEa4zuukmeP2OMrHIpMHAlSmJdm3Ec0Omy8Uk/IsUXtH3Ppu1cPcK4EMATvqfsjuj7KDBnU
NsPOomZesLm6wgKc3ZtZZVhNfoHeSCor6N/mpkocItbrd9GnaHtb4ol1/2DwGRmjT2o+R/Pjrkc6
u9O+whuo2ICel2pXJUfP/NkTMTUcTJtraikEyHAPab9WK+jFmXBghMa5CkIOSJteGldmxq7905Ra
YeGJJo1VCVyWglzBRRa21IxY+OTsRBZ0FtkvHnWo5xvsKtB9gqeXxDvB6eNDqwuckeTAVcNb0Nou
Ro8ISB0ZUqa1CURt507ybywLPXZI+BL05IL0IwH5A1cP2suY7pkky7xu6tHYucxwYfu00TskqJUB
SQm5rxW8RAHp7lZqJBsy6KPq3AIAAHAQ7WamouAtJ3igihXLQ5Ss3d3YTAqjWo/Q3pQmtaH8byXL
wjKCRlBuZ/ogGhKh9YbzPMagWQDPRgf0KvA4T9L2DYkcLLDinph2Ns4/IE8wfo492M0pTjZwNaZc
h+2lide2/IHwHaaaYuux1GcSvui8O3orffzcIcG0wW2jIyNjjkwGvSQDf+f7LV6NIUkmAPOoxLoJ
o6s7d2dPmipVCggNruvmG70ebNgiBChxsWBDjevg2I29R/SWZ3xZBIPDdI1oZw0CmJ99VNP/gPI7
hfF0ieJ5+S0T+/MS7e31xbnr2Kt4MNhaI3KhszrM8W+lgcthqw0lHY4QqT84i0yGki6N1+M3EwBj
ks7flKkJEKPlRDbU35nfTtAERWqEwAKZoair/V/RLcYIFHiDZgjnLCU/GfcNEMqcCJN59ZIAhntA
UJEdodJEfQyjQUvaVIVUKK7vU+crYgpK2JzDABdZlErBJEw8B+xReqXkHEfLvyF6PxmQDo13q+pM
XipcH6OfvvvwMF0n3nxVooU7dfbE8aE5WLhYDBS62QmKqXfbOkQelfpnqE5XJSudP5Xr3Ksy15Ki
DkgRdyPfwe+tVqB/DUKPSanuEsHNBK5tO7XkOEapUvnyl+MGfQSTyYoyw5wm0YvTlFxjeyqMtO2l
Ujmen/gtcxp8Je9y+21C6PFeJQGJ5AhdH4H2T+vt08VtxODGT4jN3qQjHE69dCMWHKbfLqze7ck/
6l3M1O4ifz+EpiJ+RzvHxiCmB21bBdBKSJO/3d9BgWApfDfWXvLkjcChayagtFvq+MxP3IXvC69T
Jj4n7SXHxEkbxOrte8Xulnq5up6Pdh6V6/B8wsz26DYoNXiJRlymrs1ArZdz2s6lff7gI80AVMoa
b3RiLyPaIQJ/qw+FHS/R2J8GitOxaa/DzePfuL5SaRrdjRCAFRT+9TvRXwtOaxxl4oF4Jn7d5cAv
VOf8R9u5GsYs5MG/UU9QN6G7je5T2su9eia/fooeO5xprVdVoEva/vpbTl/bj6ZYbOTqJOaFmHOM
F9yyUHVewzR8Tfz0/+G7Piaq7rVWDolyzxWzPH/QmbjM/ZRK3z9w6E1CQRLO2r00EtxvtrG2GuVd
4/JgMhbJqxx3ciCc6SASfG0EcKVqSwZE27HIYLnvnRyDpWL0odpRmYhl6hBu+OAiBfiCgwubjuij
/3hMY8EUP/iWdpvr9G0V7GJILl3uWa/jxwW2Od6j6K40r8LYfxarB0/PLefWRMlDAm0sWZTJSAwh
HzfzsrPTukFBUwF9xzcIQhLu2N8P7TRztK4avxLXk4ccIhuLxCkbMFJvNd21cvRB82XEYtgdNJUL
9/7HkVaUj7Uhab/NGLkM+F5pMiIQr3HhFmMEE+ApETNLCFEON8KU5M8QjImqTnI8zo/sqNwednsp
UAvKRepZIILBhrhozHoTLEVkP8BjjzYOJ3jhgPGDoxi3he7vW7JlEXQJQ8mhrbRRUWqPT1PLSHgS
c6En5+JZRzpWIOHl7OA7milbFVNlFJscf0fkLHKYlJRhdlvIknCapaFZ3w9h7l1esSjG24ttYdGe
Sh/+Id/hHPTwK6+O0Wvr9B3HscIjeMxWBq9c0W4HL9dewVnUjnldekA/ziz22Ui74DwqIC46Fkmj
EvWXje5QDa+Xa3XyQnoe271+L35N19GgBT9k3k2Ucl6/8MgJzmQB1WOg2vo4imG5bYx2SE7Tdfoa
04k5No05NDU0dfTLP+fZMbn7XkNntF41algkV4Y9u1zgrQukn6qJUq7yWtlUCENSLqgYvo0oOILP
3wBkxIkcrDJ87oTKIUjPrQQCYx9vrRaXCdIGLslSbGrLXtXpnyQobvVExcY2ZZNdsU4gp6GMypMZ
ablFVIv7UoN7oIDLpKViK9QOvpBZnI7f1Axcmxjh+f6s2eghqMPNu6FZIf4LJlXUPtDdUjfFADmH
txtwFRniPv3nIplALsu9rKMA6vGtANDZlKpVBqVXLmdxIQhixKWFSa6pmGeOaozUEee3OM6aHz04
dkKtrsPVrNbo+dG9URmgLf2XIjWC1IxigX3OTvZ++OpFqqMWatyrIrKB+MhMz8eb1RElHIzZlJvr
UX49UWUU+orlfwrWyBObGWWKTJToSNy79IHLmZ5MYY3dzDl2E7svz4OoqzkcJhgwZNNH/zwGBf0s
E2ugJWxDmXXB81kaVLDy/x6GKbkc2XogZ/6EqdG65Mlzep3kk4sF2bgp1AkT2UlL4UymUM/Tl5Mk
rBtByJ2SAgsED0qtiWoaDm5uD4+tVcOZpweqXgg/408VvGZDnxBMXoyo7K5f3Z/2oeJaHr0yC7SI
f74LvtjDjY0u6ckBLGkm/Igx4/Tz61xrGOCoAUxSkPW+rxU0//7gzgtznqtMblBcqhWC5CTRwqlr
6+roA30QPhTplND7GchYZ/WJ+/kALXBBNvnMTtGvhQiufFU7ghtr28q+cVEtqr/NWHkkJRbV8T06
bMhvLAZMSG/1x2xAKFl/ZdpbzZOHje38rl4mXFdoHWTurIjdsfjcoGTRVRBYdC9ewzcTQ0n84o+9
gKGFGfirnm/RQFr1gEqBhiH6NE5zaVhHLHyXDBHdA9S6GLwtp+1r2r11KtSYSnCLuf4ldOZA70kT
hIxMs4/h/f5QZFJXfra1UAB/ZfHQ4kzyCWEaaryh2k0dtDSZYe93ICnqYKJGhoix6+GImPaFL4uF
HR1rOmJQGi8kTVgN8RjKfD/BulYGC2F0iFFyEdtKJvfzeosrqmEONW2NcTJXOgst3Uxk+VRxSKvV
Ippu0M3/GEMfYuE37r8pHoXBeB2Gcl3/s7RR1BAu0sdQep4Gx/4FfmkhO0UHdKH2EhuW0s2xwQdK
+3S0k1g4mhSFQqtUK6c8Q4lZoxheaDGkLaVjkBy2ipqTGnR2top6+r9MgRwgzd/uOAPqjTGN4nhn
WvswoCX16cJolshKD3rksmVcrqRyMxM1azW3Oq9AJQiTQMRQvunpurSNHc0CcTm5sWSnqJlPyBXD
+CHwZocnjN3D8E9wsMQPfJXAk+hPakpU/6LnZL/+KI4XyFqrbhDiqyQ0vSaAu8BaVcQD+ft9W8+v
j+vzArLfKK2QhkAoI70JtYTGc5hYyTx+ZKG2mqhd5FTETOG4i2j2v/vHukAmCfvE5I8VIYP+o8yv
A2eIaB/JJVR/vFOT9gT/eYfZnoJCT4Xg5ODhiUgOJkfyOxtdG6PC9kG+9/w7qIUKe3pmqfizUzpR
qi4OLsXTfdymPXEZaMrjgNJakJ8ejE68EjI7ila1hKbUDRBsYp8r/WPGBJtmu7VTu5r59zCkyt2X
XDyzKqh8ZqhKbVQGX7wt8iapN1G8zg5NS1GOoooSu6/y5fKHKW+dBqEwMc3K+MyKVrO+6y0qeqsb
CEen88T1Ku0IyTHHxOZbt0xlzrkV+3I7Dgv+Sju9AMlYtnewA16wv/2L1nGt1bT7mZLxsey5+onC
ZxcSZCCbHJYZQKrUkgHNa+3AuY3gkJ8e3dx8vk+ivC1JClhNjr5jTs+sfrv7lqhrBJInp5cu6/7E
IvcL0JLB/ovcKGq8GGbyhJX2GJ3HPeEeER3O2E+9g0tkz6yVcRiwOjkuxCCQQ+ldB015+9JS8sz4
bFGfoUXgdpF1o+U8UO58AEwHw6CnzZS8IEQGfTrf4XxML+//4kdmMDzMzYa0OruZxgueEICYACx5
PFS2tJqNYo2PIJkl289PmKBvwBYwsgoYSV035A4K52derE1HuJyNUbMuQvgUWdom+wqkjbgUUzVZ
bahBXcjlVmNjXSy1SNY/QYR+TP86MdXFZEro9q22FQRVNQuJA3FoH9YzUvDKu9eDQmKMoWgrXOKn
/1YiaL2092enzm5emX8KLZtQcq6r+1MjY9NkXIucepqx+sA+ZuOAbNDqZtT2BwXoeXcrsQKCwvYv
IlA8dlJ1yVQ7FH6ug3h4joBLd7Mv+hfR/+BLn9HFAdKk4zDrvXmyDAdChcDpBRFi18bkx3DBD69c
cNQacIZzokzI7k16jvl9JpVn2Ytx3Th0fTKDRU2RGiHAOSNyv+VKUOI2ZOXg9dWWOrlnkap2S5Td
V2RiSOYyGrwXJLEILpaJmZzNM0z1RKvnwuSUURd4d421g/Hn6PeHVWrRK4k/sUyOKNvG6umxU9vw
e4qz9oTBJ9kAbAZ2DHyPCAYK+K48XJsXUobUmPpm+QP2rNXyMgDEIJbdQU3a9HYAy44en+k9uyWV
Ii8rpT7e1zI9RWowUroMbnPVfnq7//XqzrUKRVEl9UrLT3kZTLFVxd89UDNrhXGbACF3HaLE1Q6J
GKpCv0h2pwVPmsxe6RZGlJvuaIFBTw84mZSYU8bfjgEMvU8ajK8kUg7H/JoWjvzsmnZPGI7MyCgJ
3zGNt5lJzJMuuW9rgcFWQEiAyO5a/Tdp7keAhtrxB99H5a6u7BuoVE5R2tHj0sPQZgVyJO5dsXbI
grTHorASsY9FEuRblAYa9SxbkobX9iqpBxzPaZURxEts67OAjF3yjply2vtnCislIFm/LfuQRnhg
gq/N6/GN/LbZ9a9YB6nNdaDdr+M1lBMUr13hFzCEdiEuc9oKGywC08+FQxbnqc7K+O1MRZIdW9L7
9aa0eZFt+PWtIBjw2nRuu746jrsM2gJhq9QwczER5cgx1mtNBVRqGkAI0Sts393NU5pA3g17FY/x
3w+mbAW321cRWtsqI57n4uthSPkHMTPzhItFSE9+a9nb+e4hAqBfrR4q2mCizAkZQzIVDVIwUXmh
jm320G3QqzNzVIvoStW+SrCE1BAEw8T8MqOWh7b78ADg4/mwWzEwp31eeGygj7yryjN/0ms10tJL
7zYlBZ19Hp/3HZpBxXKhDb0DJmr181dSjwwA+q6R4INRKc/R/wiVc887thgqj3fdmZmXwRktnm+z
0nRm/pUtLfn5tmg10Hgj0u+swDtlu5qR7S1yR1nMyWzpovczBxni/6Q894pS/zv/gi9FbtuZ8WJ1
g6fjKApCRGouS4FQyv4vFxNgr9eaNIdSMiXGKvGBJAmK8xpd8jnf95ap/PIpP9U4N8Yc9sRxvD7H
duBTvHwbYVLobb01uiq7gFRlio6dWOGK/dytk/54P7zEg5WmyKTIS3uxxYiP93MB6BiRzjCDio6T
bmdYZ8xBL7+r2o3h1q7vTaUgYgaTSFuiTPqIZ98MK0IP6wi30fKPsHV1kIy0kDNmdaHi08DOWG7k
PQ05OJZ1V+59cQJIAp+4lmfk/NyURVBF4V7dNq8hgsyT62FNIvbQQaHfNgfPEiJlIqj2aLTd2rwT
xqRoNeaZXamvIWyppFunOxPy20pAinEB2B3nB/Wq0c/5gp3g19Qcg76DB18sT0LYbos8H7Y8JMF1
USM6v4uPyjUAgpJXChS7ncTWf/ALF4T34Dz1+YWPgS3jB/nhaA8LsyclvZYdLEBXHpqEil37orEZ
EJHFviwY1uwDhYvO40PfXnI/8r1O8fdtf6uSWENyEN851RgrVpLfWmnfTgDn+O7MGFBCoF+jYs6/
RISflEkdWMAM+KeZQGFzwQ2jEm651AowV1P+OsVcmuK6H2uZwJZHLc4mw885CEUVn9fUHrNoJ8L8
mMzSEKEmLZ3XcKll2WT+/jDgwUjQMEM1ZbF9AEVMlRU5OAuAO3kJ8Q8xEaz7k1VGkf3ReY3t3cUO
8GhQt9Yd/F0DX5H2O6MdQWh8NO53yLDQqa9JUqtRZBH6EZkctlR0jj9nKiUR4u9RQjTHuEftQF+u
5jlH0Y/b1YBfjKVDjMxDqZP0NBeR98/WIwJkY3yorz0Cv/RFV1BiAar7Rh78VHIaw0S+NOLAcieN
ZJFyNrHMALBAI3BVValLQMb8HbFzeQUQLo5hjIs0BrlrRnubbxi57klrWs7WIuqihHhL5EKG0ERm
gNP5hxUtC5foNmZPCdmNUsaRVzdWaQMvhpZqeUTQwefjRh38kNS9wX+CiqyO/dhdupGXuPj6lD5Y
QyhiKFUJtzK5wKFrLmumaogv1VgyoH3+KEqE6Fz0xzKxtYgcF+7rcKB5jRrkuAk4xJXy5wMVDa7m
jPkDJuXmNUJQOEyD/c6xcURu7yNzcUFB6nCJn+Kr00EJMbDt4fTqA0M2/HMCzHHQkEu5nBg1FbYo
pvwp+km/l6gp1Ytv2FSNz697etCKqbIVHNAYOnpXG+HmD7aIRr0nly7q6U+koaMaICeQYNObZa8O
75G6R7o+tfdVxp6k72CpRKTjgIlm2sRWFCUPCS3MHAiWEa4raZZWMb6e4iPjkgIK6/DKLzhDe+xK
xmUi4fjmd1VtnY5759lovZsPMf+2uebiKOrKd6je/cVOzX25tkgU9rxoAV6NwYRB17k74ikMPhJ4
5WaooGyjPy3WuYzme47Ww4QbTewCVLqHGDagm5tKa5CWeqjd/QbEwG5SXr0QaZNPOdkrZDmwdAOy
uoT4pFfI4BOaCP3R5wkxW0mOfIDsZYTUpgqt4a8shmAjmQvf50gNOQcVoMCYyKzHDES+DiyEacAQ
Cjn4Eia0bAMi6qVs5k6O5ZNp8SjQMk6wFo8Wqu91jjgKo8rVmDiCxwiXg3cPzb3TuN1EUG+mniEp
nOmtTxDcq4o5jw+xb01hCXsX5FpDElXCEcabwWkfVZDMqd31O0jZSvveRhPL9lgF8X4Or9KknE3Z
dpRvY6tl6YQ0yyw8VHdMF1+xoPxekHYkPBgz6hu166R6l6h51/WoNL+0sm1byr3YLfBUnJ1f7Q7R
ign9uvH54FaUsx6tTawMMrdvk9TIgSN0Bk9nYsS1gjfk++FtEqsO6MIyxRBFxg6qLLUCaUIuUXZj
kyaAwbYsSMZEBZtW9auroAEtDrEoECTwi7R1a3JAKsV7AoWHH7QdkkHK3tPV9EvmUjGxd/6oLRkF
NoKPBaYB3svrAh+OalXZuuNK5f++RkJHWI8KzzC5Zp+7q2nsq1UNGhUe+nJzLuSqeVBAab/YRXn4
p9DAPaHSXrRLA43PnwH13rUpfE32qsrQqXtqhwMRwbwfyNKTbbpk8XE7jzWloFgYeyJJVLLiaQ3Y
BTHT1zAIwqCHYD/VPQADr/7kvPnGq5oti8vpxLT6MCp+PhNRqgexxxgBpgEfXIig6Jlqc7DAh1DM
LrgODk9Hb9fvmHDvRYC5GA38ZV9X8OZKWSKEQMxcpJjJiYxtkt/BhbF35eik95JfuYUx1SRvxZac
H6+aaJFm54n/uf1u5M+ha1F+BsgizluNUwSfvFsBxlIuQxFRuDa6WQZEuovYW5y/mqp2zzpQij1W
Z55i99EFF1m/aUUDIBwwphfJkEv1AvbnqfLFq4cEtWl6YSXv+KdIcjb1IBsUWSXT03/lJx33fhz0
dXGLjLycUptYG3Qg74wxFtJRfIrDCHqhMHqZA9AiRlDDvfWGX5Ic+fwH1ElP00c0AGegVCuW/VDK
fYGWoz3jeBOBV32rMZWmlTiN5KTISa4m0GLrZsiwvxG0EdvAAfU7CPGFqwJoOcVsu/VlTAYaOUph
LyERXleBx1vh+pYSzI0FeU0ei2JseTs4KPTmPy7ikGdAKQJCku4K7J1jwIk6DG/RKZW/QzQVGagb
EJOLEiglLwMz48LBtDrJHRTV8lCgszDNtQkiRc0IdYYHwmLSTAniHr4o4zrr0603C3sac63wAPkj
sGrm8ysXWN3YZ6B4FAR7sOFMDNoXJqoBpyj5LjpmL5N+Rgsg0K8/jMLHMX9c23Psm3uaTi41Mg0U
jXui5SSVRmQErDOREgpyfUOlTdN4kgcKJPErQDFyb5xkd9FtDsDXbCuL1B7cy714vecgbyA+CLi7
BP0Hsj1e5K4hOUrg+AEaZVNLom3I10YpBetaZ9+IiBGwOTuQ728xAcHqQLbsfWkzEHByGnFs81Vi
8oCoP3tNCVxQJNNyNg6+fLDFqOiA2JCmLW8VfPoMOMfog1E+KfIHC9CMF/1Bw8mcNbLhbuOXnbqe
buasUlnDUNuv14mktltGs+opqJdfrNHpnLpllZbuDw+zOo9h/20nB6iI4vOKuwfbPVvNxXwzN4UE
gSfBC0T3rlQz5jrPhrpvbd5tqU+CAWYT/HZ58LnWluaRP6dT4gwToJhm7u3ms53Cur7F7bLEGOyS
i+g3gbMBCmn/zyv7QD2nUEGyAIyeeppEYfTom4DKNcGXVFlnYYi3kYPpJI2uQgrouX0ksHHXBaw1
0AnonisEVKSXhgFNpacZ/gLRxfebgHIedsQMMGeMcXJ9f6XIPkmO/aM4mAv++U4s38STluSXmW5T
pgRrFpSTJZypXwHN9XlhW3Q0HbuWBomoVTuoR9OeD+cETbPiO1Zpoh2N1BswaixQDM7lOAeJj9c5
ZKnG+5g/USpcAL8Mt6g0mdZO94Usakx/AmDsI2idPFjGjoJhO5mG7KzfeULS/+c3xgM4RXV3z5OD
sDcfgXHX96Wu4jhyQDWGO5GNS8hP08r4C2QsDHg6LIYZjxG2lKPkxkrIIyVlx4xK26grTDy3l6AC
f8GKfgrr6iGolak7+7y1V8QK5VMofq5+hQ0i2RhQzGht0YcxDFguOeWPyU+zEs5oRISalF7pXBMt
hcYndq1zmo2Tk8VdGIZsSyKAV2nMetvK9W3QowYz5aZKKOZSNMKS1t/CfFqtfCm/qZI66UGgTvmR
lL0PO6NtVjLDmA6sJ420DtKnItwrFnSqKYFCBzA06lvRqLF4XHrUM7FllqiTBWF5Bznb2/JheRpz
1sfFHE/c69eeicHoJTats8JS7GnBV6g5wx8LoKm11S1lrnkpDlRbSm5EKJUFfngN2hiI5z22tJvU
e9OXw3btfHLWxcPbJjtxoDNOK73rnKnFT3Oo5SqOW7PZ49dDiRnHIVeeWyoKXx6u1yp43nPt0CP9
53pPVjal2WRfdhsliVknDykASDoqTV368uId765hsrwUlIYpFuLkwSKcJR+tMDGR6FdPTKAbFOz8
qHxXaSNU6V9kmGAKSQ0f2ArgPhcmW8ktQco9HrqHafEu6j6U6M2TJM4VpJoJtI/veJekW9KGRIES
/0dguJvPsH0z3t+d1D9BhVAAbhO6SaOJVTa80TfS1/EridE+QeSlrLby155r9KRT6rucMMBJzdUc
hvu5Ab5SBH5qXG3RwH+oU7v1e/bnooGWoZCVZEaUWbkqpbQW4vkvh2GxHN4AbMb9YK9j7lAWdHj4
cNcmyR53a5jmHL5JTElMjJTZmQiZRyG2VsexSPCx4Sj70T6iRtv7NG8fYIzEYJ6S/E7C+FLlULEy
9eadUisDrABDJXz863XuuxICUcWDUosC0p6/vPNuJSL8Z8OSCHjon5tm7r0LIkeBe02fcxfSm/WL
lLpXhvaItxTGOVdnxJ7mEx0guB11PUdXLRWkHlerP26WcIT7ATR1K8x3cAkVSibdvVH/SBvwQpeB
DSxbuRkoi2ftmdQLEqvr/N95NfISROnAj46OrviWYtm+DY2z0h7KpxJRgP0/o/TSH4hI3ZxpjYfe
8MzkI13JUvOdrrAWTeyWvsV1GTi2WpTrAhK5/wSJBcgabBeGd5i94ilaK/UYr6YLHHqTHMnPQFVk
ifU9+QSJBqBd960hrZycJIPooUYrik5v2IxHM0mTTHpHnbNZeit/gaw4pcuIUUNkakrJClMNYNL1
uFYOYBzOsSwE6YbEeX8r52aI1srh60E/hZHXyOBzuD9rUGwGnTfycdwO+U/Vhs+SIbqRilYt+qsG
II+qYhJL8voR/reaZ1/IT699CLGqtdgjqiZaGjezyzBPuUUX01PsSufj8fT8Aftl1YW6qzalj8od
Zt3ZhYqlGh5Y4b6Fiio1Odp27/dnjXutkYbNK417K2qnxdftta8ZmhmqwPCOeZf1elabnMhcQaPT
9vYJAIDSdHaf+/c+pgGXSZ2paPPBBB9m9Vb9/4bJvFYhDVdpo2vjM+uhHTaNqgNvX2KReopbQrTK
Q+FcP5ncs/Jybj5hLcRvjROLmdxUdkJVV/HO1rCsMJrpWJpni5wtoJ8C0XXTUdCxnbzXuXuximY0
j3zL6Q1ytRFISeA9AvWY20FXrUBR718V4RDjG8zn/x0UXqRPA5vIpgHsWvcHSvVdutvdw9GluyQs
ZdGY2c0lBMk1PqNZJ2HAyjArHFhDQX/9tKhqzxoJ6Lkyk/qWbUE64S8YkSEL83fKWqHjV0Sy9ifX
OPI5p0N66qYZy7/2u8euyPVr4/rJDZL2/k9f+M+TTAE2d6FRoZhRWvZFh4aJ1a1XzEB1EJZgDlmr
FLf81rPuGTLFrXOm8xoD/M9dr8j8Yfb7XxCNTgqSki2LsmC+gDFSyUjULc4upQfo5TWGwE0Vn0T8
uD1oAdLmcnpjCnpESFcExmnkNwVKfGQg3nkW9TfXWMnf0413h24tvq4RI0j6+7Gu8Sm2rGSt4pN8
RGZbEQoUT/8sXvgK1BxoaBIOPlO1MMWU0KpEo1N62/mtethr8U9Llgp11C+wEN4orHFlG04D0eVI
d+w4tgl8C7JltwNZQFaj0SMVcZ+OwMl769Rr95dBmcxWYf3lksA+SNyKYK08wJG3SyVH7+T+8Hb4
0RGAaw2JtI36tQlvE+hLSGnTa8fDN0Q1JULY/BF8Ir+rSjsLzFdVMHNpnc6WZExyrBNDZ8gIEQBv
Nw08gc3Nmk6goGXniUu/Szfu+COyJ+HRYlQ8qH8YW+f0Ym5zbGLa9KR4xwDMgx+Wyftk1IeKeDfW
9R2F35xZs0CRCDx2lw9cdIyWUUDLx6Y0ibKeRfsTaAjld07yJaVp2P+/yjEvA3W+4+/Us8ELMvdY
b/DrtZGn3QomfsAFt7oMfhd0OrStWKhoWRG8zs9l1Q3u/sGBaPcwy73rvWiC6Bk79BZu15dMrvvM
j62hfsqSU8LcRkA82/vIIK6xw7ZaP9DGYsR0XQa8iaXZtHDaVMBIl//Qj7Sa6HUE8Zi3fRki+h6H
jPBhBNPPdjYGKBsDTM1kpotD/2qTUvtBabfCdq4WHsZ0Gvm46SWMHuiRa/UokP2rq83mJm57Ie6B
b122Zc9owouWwVMPHVxE/52QE6TUrtS8fpo56jQFaxfPhEfK+Jo/CcM4aj73Waij7OIpPWnBc8x6
NTcyDZo5DByH6l+A4g9/viOqm9COH2oqOB5KmzmgSfs8avP1L/AdRVGa8cEXbzvhTXI9zk/0AhCl
Xv6l2do24MsfUG7luFsLL4xiZue0W5wW4SvBozVDPPlM6ijTyPyMv1c6G6BsOZ30M2a320Pjkx6B
I2Yy+Ec8Qj1Lkco6FtrXHMfrtd/Co7vBqwKusLJiz/d3BcDwf2o+8Go35Fao7LFVQBUN7AbXy/1x
yXDfZFA/U9VSvYK0Ngg8rVBXaBUQhmBPj94FZiM0Wu5nCkKYMeL+wSleud5jQXrEsyvwOUdSHauo
eHkmJjKeZGFpU7qJKmvHg5eshmtY4C+YlKO9LOSY1bfOGPlJPTFhbBk/yjdaE2O/g5fuD5N7fcPh
mH9apMb7x8LfYc6g3vCY7unnOuH3SjVdJpjExaObh02YGvVet9CtEQ45y3ONDxQ+aISepRDsUnvL
68smiwBWMiQy2kmdJi3Z1Z0RjUV3hJBndKkBv7xF4+kN+I0/DERyRcPWNh/E2Llr1G8qQVSOjEor
pGdht7Qj0fzUwT+tHaWYDCFJqVpwIBFDMJpFM2Avqkw9FYDoEgZ/l8zt8gAzW4Im+4I+N1FrJKFj
EFHXJ31435//AoAI2SNADzlMe3GJImkEunCTqtNG7cz6idUjJ9YMmHy808dIxgx2UmBEgo0MWYKn
bARz3I+DkfsjV4Un9NRNlStir5HJ6cZ6fbHH8gmNRFHNedj5z/FPzKSXkwyemqJ60XL2FeUeaUN1
nPz0yo1PRfrxe4GMa7useff+rt8FL5Dkm1qilaRK6PzpQYCD0UtyXLeaiAYT/lQqWogTs2N2FofO
RvWGCHxFJFNMseg4FdJsTUJuYKIsZ4XLlt8acFtnPFcI1Y9KLXskRAOUbl0F9KJnnoCOjJ/FLbZX
eoJraAxz/LTDHvktbtmaYhdNinMujxeXGha0MIWJbQhdKwHLwSMh0aZH0ANhUL7/YgqQV+NMEEk7
BMkEOHPX8qrGp7x+XqpilqJtJAmHTUiCHEqsyijh36PFHN8SfZ8EWd/1mclld5DYdxeBA4D51Vjx
buSVl8i0RU1OH0X4dsptYjqkbtssV7Gknq/Op/1FNVAvkl8v1wUjqZ1YwDMFXbtLryS8XR5nTB4y
TukIXP0r777s1eIyMB6xCN0CQUUCVP/VEaL+Bm0+XHDmPMqdln8PAVlIKdMgfzlCTdZwlsOShw1x
qlP1xjv1i6ovnaWzbiyrYz/23n5MOWJEO1yDSgc06BSIEOgEYuPd8KibdSikwCPU4zUU/5gjIKKa
weDgPTyrxFfGEgydonBWb4PNlQI3hPRzsqjAGZobPRNeqEpZAxXyyWmFbZe0mwcFo+FuqaCVnzIc
N+GlTvNGXo1wfVIdXe/VuwW2pnZqdTZibNTG/qdDoLnlnmo15A8Yir0n/6+BhWglmGV4pYaEw1DZ
kP6LZE+H4RGckhYEQQt/jppeGUAvRvviLT56LtONUFEVEmVN2JA2UteIhFk8LMk1oZEKn89xz3H2
A7Dhw+1JfNL+uolpafhs91IxHcBZ8I7u9pVLKPIq3eiyYh0kI+xuRbIpglL8V8N56S2ikdCSVVfJ
QtHh7xh4Pk1RpOOdHs5UWsZMXwxUqK2PPROAfD/UdFFYBCeUJizU8rJ3WgwU2xKXGYziFdyJV9rA
pnLFlbITzFK3h7Ibods46Vv+Bi0ss1HWPo9QMGv3k26o2By0hXR4CkvGKY7e27w6JxiZgKJ5oWky
QcuFs5y1Fm6UxyvYXGWnKefQW15JtlPIEUcHzBWp8oMGRgzquWaDmnVi1k8+Hoo66n31OJpL6+IJ
uwemQNBGAeu/cVfCLAtX2h6jO7yVxcxCadPXuA0zpGUtd+3RmcXg8WiRHIed3lOkK78I0cIsjLCN
XICkXw8zmxtkfmqJPx2/ZP+VrxIpQ5Oe8sG3nwDEqlChSAdrY3FU9Nawlz4WmJ0UPrGO8aR4PgPm
Ks9BFPjCDoIN29/v/B9LGvpfGsxBhV3G1Ar4OzWH92mQlnATS1INr9NfhFbaKeIcOWcAMMR4fXR0
/TciKOua6+iEx11AOK4QVUwV+9McGzfP6xRRdeMf6NCdBNvS8Axme0dDwlNVmELHJ5+FDuqvO/K/
QQ11m1ZE94HYyC99A5JXc/2xpwd74N6/iiBYEFUFOh3kxj6aZdNFU9g4McNHGXMdbhQWBTYw4x9q
+piAP/6+H8BE/HSIs6QgVWKNW1JKDgxA6r706ZrWlAfIsF3/KmxXvFR94G4E0aKehz1dgv2lzLSw
xpaQQTq7hdggAS79HeYJN3YMy31bDDlswLbbeOVU/JyV/90Gt1EgP+tLw3EdDQcEHnNxb05LvU6W
p/Y++0udwvjMcgQ0Q5UqOqIFmijTsfFZfFIaRWgaeJ6lNa62tBXwNVaXXUe44NPw30O5TOP4+2bx
Gr9YKAn8kwAgofl3DKb+MWtAH2WczNyPtF8p/4O1bztWckBgDtNklp0tAxhqXuLIihS9jDzhGtMB
vsWFB19obNFHSh8TpFyV4urxtolhZxxKodkCa85VgVLVuIoVYg6eUFjqOtwxWHFWkFlv833ccyyj
izA+CJ//55cSmEWE1RJhkl5pwRFYv4M8ybWqTYJSL/ohOiFvjSuXhdj6+sbUcoiq9wbQGe9m6WB0
zUoyXDisHvW5PNmcP9LJgACacbGf7eN7950WX0LBepZHEgOjM3z3otKJVt+6v3bkTGRJpa8QyA3l
+r5REyLI+ZgDek5CiKUdLNynVtGZshl5/vvCDTjaGcCQudJ4JpLQq/L7VTMfiBOnEPvOr9uCgtNP
4KN9VGMkDuLUiFSJnf+2wlroLeuewXLPQhTtclpf0anmHxnu1sK/HQPgsfAomrUuNaOjmFc2qYVA
U4kwFfgeMs7YY6Ba1sQfW+Xfrl7nPBJ/a6B2Z9RsUR2X+l9gCK+nI2rLbC5r0CsZfvf2rnYC1QGK
2z308J6YoUDrHti25YM4jNSH+Evo789F4jWc1a0Kgx/LE2mEAYrvkpAkyWPelHh6PPT0kTverj2h
2SYjGCf1wut2Ii+rHxW7GWwqWGndzNVJaG6gbKtOK/BwAfWtSE+j8cE97Fc1HhijGklFvcQt8DAv
1j7w150L9oVGSlNQPwfIjKGm0FJRtX3CadpTmNV20i25jCOGeLkBMKtTmM6QL+AIsyLV1KaIo/rA
V0NHc6gbCxwwuQXmP7Uc+CQdq3YPierzjF8l0FxcgQ9e5KDpHjOkHWHhf9wzJb6Gyv5O1qwo/2LK
+/gZbp2AVn7Lx+yWX/SYhQz+FUtY3hQvsgbPtdd8zKbRUvtNlHg/K5F3ptqSimZSuZzGPUBmiUFf
bSPivWvW5JzKZ472WAa1/UhAou+jjPKMPeSPkvP9l9v3I9xE4N3dtqeOmWzmvfNPpxfIindj+dzn
/QBzeFKuS5Ls1RmP/X3PO0T/4c92qFuUTUSFWzCeNLBYS0dNqv6hruOhqOtpCyH05la38BQj8hxF
JIe03YAJ6nAVLHYKqPhjCJzQ99vCdcEe3yUpmk1Pv7PyboT57QgIjSlag/SyqBzNusjZt4xUfHah
IHZHGidSxUawf5CI71nn5LhQB5JxbPNz3MtNN17g/PicHI9IRYJ0PAnlm0OwwMAcfz0AOP6Irjz/
tiDMftiZD0j3mLFuxtYRIX0I3y8VHeU/Ub/5wWjH5kfSyTvptLsBuw/rYU+xcximEG+G8+XExEhy
tbXaieRAcygB9D5WYJLyMRwBkWw2jbzYMG64Ti1+rkYmgt8BVtx1faXdwAzZIJ2U3kAAwEFodE+E
ySvrJBjIImEm3tWJM7xoR5PM7/CqPcsgI/+0vsVmatTCPB2ikJf6oAkHkFtZ8DQDnbNJc82BJaPS
C4q29GtY2aOFu4ZKwzSe4nBQKaFSpYABk5vbNRPJdpfPBhFelUmVelCZ5tuDKZg7z6GFQJTb71WZ
HuhwS1jWIemyyCtOhwbN+YRRwyScIx4zoFM4T4ZNXmIJl7RZW0za20kSMyYlDJ2ABVaLgKt9ix2P
kVN13S8TcHX5w6dThH3yyJoE3lrgz0joF7Z6MXei0Gd7erBmcy/RVhzbGlmp6Y5Q55vaiVkUaONx
cFIkWLdmRdcOSw/YZbQyL3uMJr45vT4enIP6Vu2eEbNZiS8CE/d7bfW3yDEZJdiiDFfUA+tpyypj
BiIJvMiahR2+7yMpEX3G79HnYz09TbQ7kTJ5ARjs8opXw4X2Of0H8vZqVQ/LQRiA1wdQpwpmR5VR
VKcUctUXpwYlzDbWVKv+tp946c+HYiQZ84MO0+cOo8g5loJxwFCRkbUgEwiyXXhekJBKbrC3rtiy
WJYWPM1Ch1iVnt+CWM+gKI5uXfS5nJtJGeInlC/ptymWyf4p1NQCvK9ac5s/bgRtOV/myU5L2znd
fowyblc0qMUQafwocBnrPLwgVKjyY7YUIcE26+M31s/qJK5XTjzf4lxxlJLh5BIDSfpqytsunyiW
rMa2EotrUtLba8WB58HA6JpmdU0vSQVQ5b5jN7tWN72yCD15PDnUerq902oyLcb6Oebr7SE5OKCe
DRgdLkK8USvSdENT53tmrh/BLBM9gMmi+Qt7Z/vsUUeUNMBqb0uOUTi6buV2MZjbnysuSrIWgKLG
iDXPaLgPJZ6MQbDxhjjcSvWlNpuM0uFF01acLEKQN/VyxSSiFpVhpgejlL2sDJ+pMk3PbupfSy/h
/WpkKTtTquE8hFSGO1aCnG65Gx7CDoid7jv7vn8PZF7YD0IGrxEmk8TUdFbKmvUk5vmcGb/M7jLM
1YKNW6xNieMU3NvZRtfFBSQhV3WVGJKav3WX4Z/Gqb/+w2b6QvRQmTwicfc1xZsnEDPS48iIMhzd
SF8Uq/wWbE3eAx2Ab3XNk4AHWyYeG31N/Kvw/x5Yf7O5qnJ0xFKHO2pkcLz4kvFURMOrF6J2+l7z
34dYZdP4V2Aix/3Hb6GOcaBQOwSdnslOYzFAdeJJ4XIvVcG3V5+9xjqWoxu0KCHjcY8OpPwAKvac
0tqRoqwzpr7uFIOegtewfNGm1vABh9dIcNqRoGFpOtWX1kAKZQ1yduZumCf/NjyqNTujaHD5DBey
xAeIGQPjN+llJtYbNtAyn+ETzzjniQi5877L7C9z627IksdlEbqHvJ4562slUcADlwleB4sS3mtR
07XFpsxUg/OTS+/JPED2M4faJoEa94GFrBa5ncNNIg7VPyRyOfEkmrX+/N/QB/JiEALDK9R2F/S6
fwRHk9sNhG47oYQAhGPtrzbEgZRObLLdTczh4wj/RJ/rYi3W0YxqCshUS8q7+IELhE0lE1hHHgrd
TkEcSgnOAp9PdQ+vf0BzBMitUf6gUt2UI4f7hl6zB6LQpq7EIVODTAmHS1mAm7Jni90XndXvBgHv
ia09H+GI7eLsOa5uXVRCFbx81kBzjY5oHh4PNz9w4vDxiNXrDexnanV/1zeE3NSK/VQRhfYWFaPh
VSZ0TYIXA2dVnJVgt3j6d6BkIp0ZC8BdbaHn5OYJjF8SpMCd93j1uWSHiGFrSHLG6TUAFL+b3J7J
qIauAhFnHl0lsXlLnkuN4NGk5jaIDj1fnsYjMBkcJrWA4AiCcZ0sjcbfBTMB70yY9WD3mk1R7fAm
wCos9uT6N8J422VtMCNXqcA+5TaM2IA/uEn7MBDHsHbugqW/QFFwkgzPiM7IcvX3pp1rzbEPzH44
Rwhc3lc7d4wupFQU+sTduDTSDFOlZfw+8IjedVtNZzhs8giJW9xO91XYd1yR3m4mCoebULveFXrG
0nsXJxmjW8LvCRBlJcn9oc5F6IsO9ElaHnd1Bsq2UqcbUMAYMdsosmQrp4Calm6hVbhJyBhHLk0P
wsOOr/xrBgvAnFzNq5BVcidAvIfsU493jPkijdMPiGz80cB1zpuvY9bUX+RBHqau/0+juxq2JSd6
cZJITsOX2Y5McRKiqEw9hixII5L0hLXYKOoZniLAQiBXchu54hovsA2zViHehqBAOXSlbxAuFyw9
4V0OPshwO9Vt4ku7xiyHHFT8Wi8ckKiGeD9MDtJ7B+ObsuJ20lMjdVlL5PM5HiijGoKdwh1weqio
hMfu0w4vTT2P586O9XkOT9xJjYvNjiDx9QkDyvHCRtyt11ZRGuLl7+aaDaDvFnc7oZuieCzjuzTV
LnTp7QIIvYZ62PqL8hc70+EvFtuhJrbhHs3iQk6J1mI1ApwhFY30BUGgSm2zkthaGv1p6mlGf8em
g+dgDWsodx5HZKLEgo/7rii37ztJQo25ACqF1tti5CJsGYMLQXy48EQqUD7fmD8/k49PsxKb0JEU
szRIHYE4N2UucGjfbMF2Hl3IpXHIxl5mdiQHPgyBRUgneqPtkrG0zWbBgS6ogw/MiVzYs0Pe2BXx
8a07AS5L3zhP6iEok/jRcImloYAjYuaEDLizsqi7ZNhgZHnrg3oMRcTW+baI/OifaXdGtMJ8CTNG
XqkraTQuYfjvfcxhE1Ccx4HSIsXuL/yYom3MHxknGa73JMcqrcxQfJhml2yXsh3TFL2Vlt0/1duP
PU1jx1dkUjXbMNwALtZYYX/WyeqJ085NLOG2MeFWwlrsgbvczLSU3kJx2g2JdQpIBPTHV81M1pYe
XVlzeQGMZtRBjpIFG++gU6Pp6K8TwMjPJg/lThkhq1kXbLKfe4AH86YBViHJOE4c4UWDRZ0tActL
eVcJkoxqyOVqC4/pATSpsGqJP6ezRuoQZCjSmOYuhPhPIICHMDQChH5jnVFzJY74khg2hzEIK3Kj
usON6XhO1UVanlM2/mXyLdUXAOTf7A0z9rl6Xn7e6bLtH+fPfWOIwX+oKXQ6XmBuoCEexWFGDcEG
oiGBooLF5fuS9Lq9Fe6nP7bRnkCA/0Z2yHEZ4S6EC7noXiuvu8qxHhYw74MSXy50grHdTjx8ehTx
kJTA7MuzQBB0znZcJvqUc6H1zEgKwhqXngKQ47/v3cncDiTmzPoLZaJR/ZaQoUpCv3BXC3gieoj7
ic3hZzSrXD+y/l8Cjwm+b9cK1psb9x6FcqO+y3zI60HUiadIUPgy9/PoXFpHRu8R2Kum7jUTX4Co
vfkjatjc8YAN5ZOmmf1WaS9tb02ydvnrSaLI9UWGXbSnJOrju00WTfzKpZ71ZHgV3i8IbB71OqpT
pOeaLvGt7oFEF7MRqZtSko/U14Tm23ut3E0xk2/NwL9K+RZDYpY9SPucK2wALFOnw464Sy0z7hsq
FCIdn8ZKBynYr8z1tjLINGBuGd2iqLFUZxT31t136vnMaSBsaCBN4NxuTItnF4GQY3165xidyLhd
jm1FaIgsdI31sdkyNGyjR6bSUQ/pOHyhuBxRFwOZmocTnrYg6f1mu8rUn6HjTn/UgIi7mEx4bnEC
Du32FZuXByg38qutv/yYgNOoHQpCoYXaGEUvPBlu9LTYueoNc7PV9FyzP0+H8MCQnBvdzjERVhlz
h2AC/V9b21e7ZtWIjG0ShK/GOpxUCGrePEr1E38HCGcJmqpioVFSSSkxsmk79STsBagWsE+M7bgg
96PF1sckpEOWMPuFxiK8AIaQYTpcGvSXGS0sJxowEFHVhWow1PedpfrKA6Wwl50XhJYk2VCht274
R1Z5Ms12cGntIiIRV/sulVBXs+QJPcjL/I7aZGNYaVSdYlSf3i7WxXbRqbBQp6nhKtr8aoG5gnt7
4DYrLq5EhQ48hnlYg2rzYlIkyJB1/JiE/yaTTh/D9NsHirXEgw8fsTlWsupE1KjrwopfuyM1yFGE
sEwBn7GbxGvjG+l4OxL8xnoKQPjhd26XTPoPJvHQSmQhPvAoivSsMwTjAB3i/QIvA8L9Ujk+zKhN
KgNBDT/vG35Y2M7004PeTRvNvKZpbSc50H1joR1Y30sThatOui0RR+W5DCbHlcfg2/zhC2218FXk
KADQUEeTl9/0D6HPAyisI5VjuUecNKDSbXf/Mv8qZkOzDgR/C2NDyNGuAsoKAmFdUT9eJtzzPpy6
BZLWEOjx87EjIyQ2Zx0qyvzLE3SESF1feqqbhexGbEDMRneeePDIWSmPNzRZe01wghq6UurbUqgC
bObR/Hix5XJc1EXgYtDBHkRWYsOHnRLFUQ7juOpF0pyYko/N87o6sVYyQG3LcvGYpLO3ClLJ0nIA
NUqX+KMgBKu+f4NmkYvLUp1qzQtvWWPf1Pk7uqmwjEdt7KTGRYXw8jeGbZNtp8CEBB6lC10EU9Za
epJLThy10hWX0ADHt/CEiBk/JI3zY0dfxbcWb10deMKgsRqkdtuoRsRz/EjTzFTsxYRGA5P7EjCa
Mh8te2nPMP1D9kOnsh8rIeZgFUeUmF6ntiajZ+sTsPjSmLv+qqswqN4R7Wmkko2QHwfuJvkYXKVm
XAmqBhgoIQAAeXfyYEoqSCxQcwHjYZJAuYWswqRrvVbW8eGzAcl4iBhLl1ny1o5QfVAW1mny6jrM
AhAdolh+WBssbS7JiSa0xq/kopUWmsqhVBtR5DotqEWUOfmlcXkfA3NOTbeoHHgrW1X+TYXyWhqc
FUvLsFH1UTs7RwRrzFOJ3nvCWay3ZtnW4EhXSPxd9cwj27PSsN6e+L11tCPfLHUS6vSzs1QFB7CQ
lxt8UCNtTA/hfytWQQgh2va7uZQpAP8rG9u/wuAZGObxmKJooDRVPjs0gXKDl27dL00GhiorUTH+
01hr76sMH+tS9fjJk3cuKQgamj0u6jDi9ZACS8VpXyBQ05OLsDtMKil791bY1an+nACKGSnvLv8P
T/3k+5x7hSa7i1YTm78h7+cTSmul4IB2IM/UF/4CF5RSOqg51x6zsR4hyfuesF5daQltVl9iemLv
UxP8LjqQa86HmgzrPwoxxGoyV00RY+VQ8REA/Z7TM0LgJlFb22khC9fNJJqvZQovmD0O9rh3mqBd
zGilbhIfD/KfeTcWVI+JJo3eT28UaT37ts06hrdPv+toj+AfOsfcQBCdFJInriS0f/R6K3W9P+31
fuheLBghoyP/Z3HdzyYRoWaPX/LlUv9P40jiwbuT+0oHrorZ7R4sVYmkuBPxUzdLXkT8AD5acaOE
XyNXyYyoCuaCSifPyCYeLVkZgqtdre+F8op5u+wWH0VZfc+J8OAwW31EYupi1qjIUU42TTncIqtC
ReO7tEgpnlJj7Bybke06NGkaQZ/9wSmBFnfaKBaSxPWdwptlzQUeXaiYCyWFHJnlkf++hpl60d9A
PD62XgDQRBtdo24NTM5l+BRTSLH4llxz1cQ3GF4gCwI/bFqFcaP5MaTkuVzXzJxzj1NosT1KDaUF
oObGso2ke54JumVyEPRkjfeV0uebiw2JjU8OVbB4rBDWRxuAGtQjhluxiL80xnjvucPY5P9cvs5j
vfLhXWOnBhnPQFqykE3yvoSmmXCn+IXYZzvtavFuTpEo/2rPml+eN5M+oEAh8ySrLcXvBrlDoHvd
PtExEQVBYmLRBcMdIIha/uZoEvZoSpfimKdMd6LD0TCkYdEzbSHVoIaxPo+c3Ey+i/liNnHdO0Ur
iLs30jDDaeuOkf6txlPoOlpNCE0yBcMCiyi+M6KbX8LXc0UzEDkpRkDp84qrENORSmgK0S+/nR0Q
8s26k8OrI0sBH2CTdEvDPVKv8HphSkgdBF87A7Jzj0QsyzwdF750mQkT5vdGWBnt9F7cScKyCxCG
WKHGnlKgO+4+ta/fqrevfgfyAS6UnM3ONrFCF4hPfcDspswZfwBm3HHpX/BkJFFiKK4pckidVMxw
0HzDMZnv2Y9eRBgWH9wnu5vmucc6yMo14aA5gZlyzULzGfZseI04kXm4fi/c/8QT2ZsQQ2Gzd09X
lIp0CcVQXl0VBSZJ3DHSD+6ScDpEoYuYUwsjM4lgLDtnwltydI4fLtLl5v9ASd36N/GZ0glbDIi3
jE28O0/l1m8qu3eFfpJ/44DsVjFZ2ahbx0qUV/705hrK51l7bVoHahOhinwUn+XKkaZ8z0Xl/Va/
sNt5Xi5IULZrh4H8YmyafRrcUa+IFn8Ei0v+qkYpzOr+UfqeTKdICfc13+rrC3VhcdIRs+K1jIDY
jHEHTkM1i0btB6r/y2SyqQ0MTpRA2siH+7Da0xLtpTTtzURC0OsWiknfsfjtjb/+ihJu4skDu8bQ
F9qXoxqjepBm9PswPGRVEuhGSc4+C5IWkWThKd8u3IekaMKdXemttyuNuy5kGOxr1OX2bOWhHshf
JnsBhGZo4pVzX880hilHPcMHpKskBxBqHJYNfU8TG6tMCyJ6LgU9yVvFDJD1dVHUqvgAde6QzIbB
T8ReAsnyqQnJ1gmtoVB3DxCu8maKMiftKHeOrh8KJjOzHQJE6+nimP40cGa7Y0FiCFhD5D13yQYT
BgrRRNmsDleVsYTe9Gjy+ApjVl2cdaZC6fZyjxFATq5b/fzRXrggTFT1/bYZNxPCcBIB3yGhzPjI
v6Bd1jCID8s7HADhjqxlftS2PCRXfA9YuJL6tpc4R0DFbMTWOyeV4d6+JwBOUDpywJv3eDfOynAe
LteG5vXGYpxy8MiEu9C7OMp3duFC00GtTupNoZgBQTsDmicRujQSJ4JGv0GLdOSnksfqwwwF+/Qk
UxrGc3hRaWkRV65LZbkVPoQIV9gaK5jg9pitnkpF5QJfyz6YGCcnCKYvNzc1EGfn19aQf8hrnCfh
XEbZ+J3zWtvMNKh0T+HwmHQXw0SXArfFyfDPjnBtNg9vnxiTz4koZ7qSsbAaxPLFM/F450nAVXbj
OpyVFj21y49T2go+J/9fb6IKgAdTmNxyoKkdwkDJ6Wlolr/KkKGxCwowDXUSkzeLpdwmRUITRCJO
0jXGU4s/bFj8DPKCQMcI1cw/aJeE0gugfIFEvMSicf9a0YE7OVZsI5ByjyDekSvl7nFxDdSkOzzM
0IV0050YYKzfoMACJY3l/7v4iUnVXhcdn/Y0pdY2pBxwYa8hrrEqRWxrE9snSbTVR7H04UhV/WzR
aVIr+vVteA2kSCAyoaCDc3mbYd9aTVcIFpBndBeRUox0ekJ4ybepP4FehVpdTMBI8Jc2nbs/OlZs
VPGC6n1RQCO/lN8Dg8hRCeHVl3MSXLIEuNTO7+yfKuFlQGOCOv5YPFpYfwIDWEcXdx7k34clqP/n
Q7fEkGeBdLTwXkyOg1eOr7pbFyMTFd/cQ9uIjGU+STI15Vy8ZeBpGTspFiaNjGKbxuvqWcvwTQ2E
oYSegkcna4rJI5qsMUAnYxd/UAj4N9pNaog+ko2khla7H0sAGsLvyQ0ygJkFDDBPRfj8UI/6373A
a1Sz574CeVRevlgyub99VzH0ObgFXYxc5+y936wIgYZ1/GdEU2tlCss+WuHUAq70wizfz2euPUXP
pInpVy8rifRvWkRSSEOvEwX1VV1xU3dXGEL2vVG7bTTszosrW8XdieGDlWbR5jg1hCXOJMcVcGMs
cGJmuaF9lyNfugyyGrodGjHasUUiO5lcBnhvgZNvlYnyZaNxPWGGKWyqeWb0BBbbYnbNQh0GOZsa
6Q0G7y+YpMKsH7ynGYnsG1Q8Y5Feeu6cdp+cMaCTZl1gQlMpaA8RnMpscTIkQMhKPsWRwe1vDtcS
fs/jS7GA9g5nZ2vNO6xSkp/qNsON9vw78w5PAWRYX0pLP77lolODj773pY8hiXdNgAd6CYYmh2ZR
kJ51Z4IgRd7gh3HL0wMEHptw5M0RVuISLqfRuHubDm5Uo9bhsxD0KCm3mgxqLmdCnW6MhqYBdn5s
irDwu2qPDgq3lnt8kjNxZahis7yeoPa5rmR67EbPKaiLXfWqEneNKtLnWxVlDdLPkSxX76roWlob
JSMPDkt+S2TgWgt/E/FkoCBVYuT6u7O4o4zem3fmvGbv3hffToLmBRiWjGeR1u/zaZDls3UqYh0E
NbpVjz9gAkLoFfQDq3KU3j6JhFtGWAe5iLuYtREJlXQs0iC50CMXpvZq9Lj8MKHRl0c5lhkeyClx
6fP4AOUmQMroUWKSAWo5D55SRBYl3b4SfJyL2ZfPdlM3HrY4pMNrCRgB3i/rdX0/fGJizbE02Nah
Y08SfXBGCf/TsqpKCc8TzYVB35I3Zg2IszIWAmDTosSxJHAtqQ7t7DgRL4H3ksGZR/VGbPrIuSOG
H+52xRUEqFZkXyh9YEQbfRNAcbmlRPr0/sBgHv9PG2EgBS8q7TJtkfzbWRFPDYHMeSFhF8rjLsIm
SjDkc9PWLIdl/QgYUc7TCGirChrlJnHgbRavmLl5b9+EFFyH81ljCoZf+5z+p1qyunyWwPY9oqfT
qvXiCF8OdWo903PSZahTQ444753pTJsn+++xxYB8bHYGK0vx+N3kgmAc/+QKKV9OyZj1UDk3pmjw
ZRtLqM9sx7KykRxzxaz7hlDohr1VcWw/31JYnUzzlzl75HOp8ORkQqSLQpXDz70uyAr7A0lD51o5
t00nxwLQwdxMwh7PteUC4UtEq3IaJL0gPOMCL1q90Fac1IvGHf2vdNyh/WaRWOf9fppF9fUn1ya1
A4/DF0kFvFyMw6SZ0myW2gFDF0hLtWuqjm3tTCZJqwYPDjgREyPMf5pcmayKvj86/PsVMmvyVxfL
NQIvNslWG0lThQ8H+hmvEDurLiZtzGIwlCILY7z6F5TJILU120PAy6WmxGPooRKQpD3QnQQFjOtR
Fc1wEvHtHtyIoSHjOBoN56lo6x5uR+42P9h47rBwsqKxCozx4QcTOc5NJJA3Cs5Lmp6bfgFVRbcN
jyci+FjFBHvRAawzDIr6DsGqepbTccnr+WTEs+4R/OfO1iYV0aFL/L9/LzyHpEWfJKH0339tjbVR
T7kq3FNd/hJ+fYYFVQca2A/2mab0ZUbsf1yGMwGwB+BKxfPLDRcwTPqFHuX1FGkODrrb9c/lN2vJ
1H+cA1Sfxnv1CUQocP2mYXK0q26FI0JhD29ZedLwlr4RskCgjTOCJy0QL8C6WRWePY+15UlM7yFi
5vZ6tWb5e5EQpWQ5bAxDUluSphqh0lXnNfueWwtJXTKykJrzYFNL27ieE0r4le1c8HOb7/CW2/oN
koqaGyZ5xr82LboDBjjfXZAQ7ed0tSlUOFPfucCQ9wUbR7V2kQSmTp0ve8AjweQS8srsRxGkjo1U
crF+FW0Pfh90IBg+5K4Z+6WTwsy2+SDzdNc9J2MqBgvQKvorO9sWfNs/aREk83WsUJ1FmBWZMFar
Y0gvXpb7DR9cBXaSRNXecULNGoSWm/f71RaWCTz6Is3GcWc/sCrChcpDcpmq1x1X0GeqZRlgDZXl
37aHfRbe3ns/02Y1WIFxWoBQF5aGrYJoc6qq0dXLsV1sMC1yd44Y/kPv7TBLtgkKIRkBeteE7O3Q
G/XMFZgr6kJkww9ufTX4LnUtiDxdwNbpy+HdcqOUy60ufZgG50nRyxB2au4B2qI2yUt+2bu5FZY8
dhydjElxTEmt3yOwtA6n0wCkCiXbXHzIRioTeTU2nZGvJvAI/Dx9gChC5ZCUeDMEBWX4a5R7Se0U
PDNnrP6E4cq6wsoWxPPkWBP/rf6xrHU3lgVKQHGVabDmap7pAXDOfMU3RQr4C3BIyOrHrbB+JH/o
pfgV01XQL7LKDgcEI5IgTjAghZb3h276qxSKZDOCStcuLbHVtKcnlrxjkJfaTCsOrKEYl3d9r1dv
dosqO2UjjdaLGX6jlqjFvKvKN7PJG744usg2ISaV/+wgoCKB16rNrbuAfE2CZNx2+AWXVQHdO3Fa
KFBg7UMN6HG9lWnK6s0S3lx/j3YsSpjCVuHDYxipEhukjujV84gzufvO2XUKQwFO4CwOlbxonNqW
nvYDXG2c8N+MBOIpxtbXmBX6+nYPQ/gItN6HosEsKd52k+uUOgD4PxNN688fNU0Zvw/IxgdotcUW
b6O4c/yjLa6fBBlOdV8yiW83IYrrW1UToEIoReE/H2mk5MttSaQwn/hPVoPl1JItumKsmqD6svxc
pm2FmnQ+hydw0PAT1khHZlPTiMire510e0NfYf63335fY9yjigUPiadTUQxNhekrWhEi+IJfn1Ar
R/GpA5ZDT9jRusy0hD86/fmlchwcNFKLWZjSYgAf+8A385SQS0VD1EAavqA6Y3YgNTZhrypSZ9GB
b5q00p5VWXpA/LSwO4SdsDauXYraUruncQbQ63GDSSJ8r41eXnxXT9H0p9nMYO/7c0D6P8A2i6ed
OQ0CaYD1n/C15T+z0YqY8V+7BMjiFMPtP02bWC5CQxdV6s0tKBPgahKaBT6oFi8vOIzWYqfJlV/3
JnmHo2gEd1H27Xa6lRk9fFYb9nMa5NcEZuLIk1z6JnG7k49y+N30y7dwh1x3ZSflbxGsGiVjBdpo
9IxSrsy6e5DXh4DFfiA+8hO9zyg2FFLV+gGNpPDQvX/0nzf7YVlZR3EdqfyHPZvYFOe1mPVHkehK
P0pvYJycgS6M412aFdiiKy1sKFfvcmnlS5vGk9SneIjwOCqLZJGYlY70r0/DFngOMVHEV1d+KdHZ
ebq094ggXith3RjFsPkQ2sIuw1brodpS+KvT6OS1/fbTdRhFCx0fQuaEsUGUUsYUnnyumblFKzM5
bVJle5Izu8ff0CYmLLqnlf4G7Xnw09O69ece2JguQjavLplV5bssALKXBQNmeyUXI0cNBKWZT7Py
dLiYqhshB7YWA55C4q9nKuo6J375QWxW6Z2BQgA9OrzgoRzrF/A12R1eiLv1/V1DceLbIW/+ihmw
xF6hdTW4Qe4OSs29G2OPJbwhZiR8R0Sk9sHJpH5LF1qfNm8y5P3LxrpyPYBkZodzEAVlJz40hVAf
sF0E4sJKbtCDUtvL0mjQxj+l+CXRfgn6DDskcoqUzXzUOgU00HxsMWjnJpoOGnlEScDbWkLwmSu2
iVMb4zSVpzZIJcw71ybn2Dn/4sVRmRmtz0y2FytXILfGvfEuMo9Lwxiul6g2EMxMbZhXkUJQKmhW
ascJ0fB+s0KoujKOmRx/AHAaLoyMl1B/0XejfLJgSLwkgzD4zDRaUmR/P3IKb4/wtgKpG4aEse+J
D3CvWmlhjiffJxX2Vm88LzNPgVPzPNR9Q+Jxdk8cU5LKolMCob9f85LU+Va1lAJbN9Qt7juoZLJ/
sW0WCMg7BaTF1XcvHshIIWG7t6Ic8N+ME0yRPzzP8mGjnWexcg4OsoNH/HXu3xuLeBm/EEv/kDZT
JIzaP0f/PdHJcGRtLwnF4CEgjB4g6G3qNgVoV8a8iR8u52n4Bm5miYYJam8LuayA0cKhi0Y896Dl
BGRX/W3WqSY8xwVggD8VOo7lBZm0t2iEZ5zMkcQ3kk/4PwP7PQOskzs5siOdXozcIlzx2HrGm9z9
wCFsMYg7ofabz91f8wQjerrVudce3Z+YDCaJF21rgGL0XV4wQ2mWj2fTerzgqHmW0f3nNw+zmJkQ
0YhjQxBLgTX5+qzCaYQlaSPZVBx47NxTn4N8jTpYRDM/GbY6I2Jsj+YadeKFWydFRLe13Qn+9JsK
XI/ObnSGobR9+L+uyWBl8bb6+AVewuzvvBbIWgn7nzpiNa4mqYNWgwgosM4uWvqkmf4UdF1VP8gq
cOVC2jR9AbKX737a6bPb9pJQH6yYzlntuDJFjjZShaGxA7PimAAqJbosN+JYWS/XMCoAltFNg8Z8
ljbDWBB8aA2iPd71fijMjl3gDtvFzRX3qoJz+xrYzlwOEhRHLju4/WCW77CULtBNkKG3iBnsTsyJ
5AoF2lnI87hKkt6BszyWDBvrQ9tQqZ7JecrfozBqhNtM6Hvg92dUWWMnA8MqbZhVDSsh5WfZAVq7
9W9tY/LOJ+5eafWhpAyKJvN5rjN9EiKLXM3PQMM9ZUCqfCAmnaA3cI2NdNtqEq75j0kNdIVdqixK
k+xPDGp/Kept5PSdTpCI/9z8LqBPsYIPC2+uSueBjGqXqvAj7XtujCkg+mIWj27YH6/m1WJ45iGt
RSGzIwiqs34e6zJJpLmZAfyi5I5MYQFieZ/9qqKYXNmiOgWE+GHUU1dp4BQrGrrhOSCTXi2ljQoG
KeWiDwGxPC6kBWm2JjE4khqMdCOt6SCwH2++DIrRsTKB/GPuG4RRxOzwXPmwMqmQX6e4OJK/WDpd
CqnnSPYDy+syhgyCuiG/TM7LnDkFN7lX5FECktnoVK56DFRI3ohSS6U6DluejxUx2UUeyYe9VPUZ
5j+XsW9rQFM5wGhWsTqiV98Fs5w3PAStGShEKoHN4351Sd8n6FvWtuZCPNmUAeP1r1KKeEMlwiwG
DcPkqgSI5BbPWFGWCAvayKImhcwYGSlunKu8mjylHg1ecP+flnUd8mqLbaFIODYmHwGv7rRxDmde
N7V0zkG7quVq0aGRmzlHqgZE+DZPBCocYtkb682DjjgXEuJaG5jGfe3RX5V+m/SPwD1eoqOzpEeu
2Kp0rnV1EvPSh8uvubOcEefWVYsfHImDHGtOolJ+PKtAxb5DF21LacmAfM4NWX4vDbllbGs/fNCR
wD7WCEAyW0gh1NjJj8HPXmSXwyWnzAhk6OAsP9OwH/3iZw+ua/ZN4X/83GOfqBg/SQxOX8nC4P8z
4ZSwesIDaBH74vdQPwhjKHJuk/OKQ9Lujd45p8WVjMS/sVzpXCzglMsJ8ttNMJGeexobIW3qoi9Z
T1PrX417tinCctzHzFSN4eBTgDko36aN3eHNejMEZ5WiME1/zvxfon3gcdggf/yFJror6jqgu2Wy
2Q/ejYIxsaDQfuFWYs6+taTAfQMuzF34DWcLFrVkScsbLLJ+prCpH+l2SVy/aVYapV2Plym4QTYT
yzhOc3jr21gLnttRdgh2zvDGFWKRuXMugC9ULIs0FQwadEjuXMfEAFuCNSmkWfYPLznukA6Jd2m1
rm7iRrrqvnD3PZPs2tJChJurlErdhpN6FORFVZwV80dJZyTCFUlabhRVjZ42eLTr2+l+J4TgdGN/
6J0kIF8O3WGujIF4QWdlryxqQMaix7FatYt264Q+CbECNvNGFxkUcFi4zhMtyFASXRFwtWfOyVjE
KlmXiBTlsnEhu0QjauBYwRYANWY7FBGq3NVx4VbNcSm4wQZhLEX4orPFuWZPIuYiruDgVTCxrYL0
3Zicc6CIGONe1m/PsV1miQxHOwatxismBs0fsEXUV4X+6ktqYsChNcxNQBPB0nfirtzTXDjxtaVd
s+JGxVebKb25aXFTcfqCpgP8P6xNMMcC+S9MX9pyZvaJZPj8SahGKiqnKd/Ab6yQ/dUc8ycR60/s
hulbmuvvRqHhCyNibt5/zWueMNg8iCbRQOjEpYNQCGiuZ+qYL6cM21cMORFD/5KSRVsZIfT8I+wi
3VwxlPvY4gxkWEC1+1fQcPz2DFUXBAUknk3ddVYaLBE7vbg0lR1Cr2PefOQskfcv43F0XFsNsKVT
8xh/dqJwWiac+cbPc6HkXpvGXTGxx8UQUazP67ztfq3E7GmN2rS8fJ2cW6C2mSYWI4pi9Ql2+QBP
PqkuKM42xx/8J1NW3w5JND8K4uDQlUF7TQVx5VAuRhmGmU6sN+BrWW/1YPb4IrPoK3PD2Hxi2Xup
e2Vmw3ZLEhaN8gkMEHJAZImhD5X+R1ApVE4/VLAXBQkgM0WyXUcoJ1+lFZSoREnqYAE17e+OzsCp
XMh4u62l00Vwc2TaxyS9Zj+yMR7JhlEkpQiRF/2knuyhMc6G2hGV33PsoWTgsjYENt/NEoiUEN9B
AIHABYitCkcTMWAD71OGi+YOS+2WWirLCn5nqW/9eQunK/bT7H3PnfUrvIvnnU4+Edo/32Dye3Js
hJ5IyxQxDo4ckJf+5cRtXaoJODYEUnQMs+R6RzeewTMU+jOgGjkJ/TyPUFptSmERl8gjILAUWAO1
KrwdRwQaoIKdB+V66WbewvWAHV6MOyJrRf7VjkZF3ZVF8z+1OGsYbGVmSBYifVGcMEDW6zy/AjO2
aQwfBUOC3pM4czq+OEZrkUqJfgQffO6qYLKR/LLv8ZGPD62ZosvNmsxJ/5ugAeeDzlQmnCTm3izi
vtg80E/hNokK7F8h/+9qvhNunuOTahzWpDL5i9ZwyT2c77S3rx5CJkNB1ug0Ermg6p3NBd8auoNK
F7GGqT6XZUd3hOyZIjO66PUE+mhXUbXFjuPKFtwDFx/JSrZCYyOmijg5eiCvyI5R5AVRSjr7sYik
oCHkDUBOTcvMZi75k8idWgSuKZXEc9qEJ4nAfB6rqjV3PeHYCHIae/bpkhtEKGvZELz32r+ziuZn
AEkUJdJjxhuNoc2ctoFg+ZMrixOJwmCv6oSDZZqHdDthFyXX8WEv9YOKo/2J4Bc3WW9l9xv3P4cf
mQDgIn4Y/klBbHo1C0cVEDZ7hG3V02+Pfb/uAkeJF54DDveGa+1i03KM00RlH2nbcz3N/Zq+WwgF
EYFuaqUiUmF0+tEAA00TEYtETijje7E/VscJR4N6MHIP9H6WIO62ZrfXTZby56yXNTZPjB1C4is5
husnNWNqo/w4G5XeoVVZ9yqStfoB7NEpb1NvTVCltEc8azDDgXqD7BHgIG5jiNES6rPyBHzPMCz8
7Y8OtQbSMV+h3evy6gv72lMwG1HQbMy1JyJn4Sb1px2QK8bV8pIyRKNDoTUZrEl0Otvx+khomYXL
klzgFLfQsg8+tM7qonXcb2msx/f68UEVH1L1FKI/yoOEE2TM/9+vbfHHZyPmQZtCkh0NcB3rUkJk
RKrGpd8ITiC+N/J+mSXysN+I3QakiXJBXbs2KPC7kxrRDuN1LBG3kHPPdOChg7nkMYTi/T5scvkj
Qgu9uvoQOCWCezNAgYD3Pv/PWJBtf0OUyyMJOqwMAdIKnfZEP2rOyuSI+yamGmq9LZZIUUiq4utt
i1iAUumOPY0co/GzLVoVRYy3zbDjgQICx+BNc7+uS2O+xCAObEemd19cjSFb2HUO4AabYlijoKi2
KTMnA61fPPIqXL4Oi/7H1XwH3uPIvJtmzGUOTwtIyEOWq0t0F2q4/yiPb3uY/QJxfnwA3tuk5UHO
jTpS8glvx60IH7vpgX00njoGLAQKnDvLz59eaLWKM5ahJ+i6sfAZIZNo6Ulgm2Rmufn8Uo9wCV0k
x3QT4/xwEWnNP5BtNkqBt3g3JLql47uD/tDJb+uHohrKy17Qc2TNNg4E3I8JwVdHSO1wV628CtNn
ea7jbXX5A89VHKyJL71/O1gpaveqntidjL1olRtoXiIum/qcroTkGY9779w1W5jC9JFbgE5YCi6y
06otsIW6Xfdk4mGBSNN8qCd4b7usZw6OtYX7Lch+ow4iQtV28SmwiuLZZKuJ7G/B1AX+tLz/B6pR
22iW0aUOxOj/UodZ7ZghNDkMxX/JgWrygsBjhJPW3xdfmdSKM+b8tTsGZCOlP819X2brKd7Pk3cb
Pzi3MlrE6mftw9Yez4AmjdBAIXlwj8Chh3I7XFduxLrTVtusDEpj9uAWSmc2Yq7vuy17BkIecMjH
0GdrpzWUsM+gS/F9HQwOkcGMtYKKmohiFQaaz37Dn8/BGY1ZIRH11x4jHaPPp8DtIQRODhy8ukdP
nX9dYx0aXaFo8H4MEyBiGFxtE14OVoWXQof2mPDahUVKJt1YgNIguhjico1JaIrijBKg7V3mWP+V
MXera9MppGlQOAvdIzNlMPasWzFcV9dmMOj6CNau10yXOlVPjM3gSY6EZyK6/1Dm0BPYis2aq97k
I9jvQjKMwLLGhPSdl4Lbaroxi/5xDzQi0yAoARBAVeW8SX4EQ5AaR7su7sDZB972iawQE3lFVXWj
eE7xr59MbYw4AGun6CHcAw4a+u4XcrZCBl8HLAEmptx3R9ShQcLxn8oFvXqqRCMsaCSoZWHZ4OId
HE/XlsSHQOatFzECKtsCYP0E5UM07GRySr7r+rq0RiZxnIjT6onNd6G/MRCet6zxiJWS8Dji6SeG
D2S44rFWnfi63xw5k1jcTtD+M/5GFbNLrFzyirqSlbWkVw8lCRfxeoIW7Oh5unZa+vL3UQ5m9fEQ
lpUHzXm9AvSuwhcyZD7/5Uxu5qTsi5LtCP5SYIkkxyEAAtOAlbbRKjDbixbQmoVbZVMRdwwrtZ2l
bPh5zbyrd907ZHVpCorEQ8UOqIWfC9Z9oz0rgl04klHDtuk0x+NvbU3UkfosiIFkSgH0z9HUzFsW
yhSSXUXBJpicQHNQAmTRMMg1UbHmcQsIV5iVClGYugGWGcmiA6n2Ufby3p55z7Qj3NS/BFnYGFvp
qwVCViBm6ta7vZFJZsLawjIMepZkogyfPG3P9yl2hDsuFCv8M8ni5tNFs7j2xiRIeYHX5ighJwDc
2pvDnEGphPqKtOis5oFFUD5H+H6JEk4IR94inl4Myj09N8j3GN07RFuZ/LplHkn9AmJyKQCt11v9
i5LuTHnuYZx9pu80X/eMJGOQc+RrRxA5T9OBqIhBZ7bp329SezpCLLTbpPjWutAp5N+g0wS9DBkw
L8MUsuDRoDLrxARdoXO3kWqC9++RjSeI6Yho+goRtwTAgIM0vHEcJVeP6Pd3f/66Oi1NuFn5J1oK
EHk8yHjhAm2pv7cyZwNu9S3y15wazLMLqh8U8uxmPPF1VUUIHOzXr2I+u9bAiOahrKVVL2Tc/Ues
BuZRTU+3F8R2hEOkl6RFHiGPGPwrv/lmkMUYct3mLF+Y/xGknfgfgJFMhU5XTSan7p2tMfsTcsiw
0USf4C5ajdHa+HaINMT3mG/ITtJbl9dRJtyZnrMYomWA3KoykP8z07EHQSUFzhpD/vY6RQ0xmzNI
llOaxm3jj6auVGAkE9XdHUiI/Y+ya9VMqG/1BaUiI7YyiziWLm5yBfY81FrRRGqds5tUw47nac2L
c5XvmFIngTW2H2IU/i5+HflhLdCpHqfbWYfPLsPXNG8iO9GkFLuukx/iUxAVrEdWGKM68aL/hYWT
dXfsxwV1MrxvqOKWBLUmvVCFYTnJcgAriKiqQ7HWH2W2Xqk6lzIZ1w46z0xDtut4hDXL1QDmKAh0
3VM+Nt890bGUKeNIigyxiI5pOx8GqOyXPKOObkzsj+vBXy7eoUR77fSkVJ2JcpUY66f7WTXMdfHC
k8BnCnnBH6w/uDh3MtWgWScwmU+ntkkUWlLmn4+UBOo1Mpj4yHkUrxqlzvw8CkAgdQqtxas4mjYY
2yOETixkhjI2qeqToQfe6MdK+JQe847E0YAlnJEQktE5PH5g5hvNC7Dd2rf5j6d50CGL5BQW6nF9
zjENiOLvffI6Urtj7hA4P0MMNAawoxc19CNBrqQ0ORfECYMWQNpxARJsZIumsdzk1b4exUdpbMfx
laelYX06IG0TzeOnTjlWTs7F1LvIY8vjy6eYoGK6Zn9gEArPmMH9jARq/22r4RVrIE9odP4dlenD
1o7yImsRaErAftFYSB1EL00n6PW1PYL1PC152SHFjiN96LWPlF69WPucp11vXd8/sTE6rx8uN05K
oVsJ8wtc+aDRgm2XNTnfXrDVNWW8jr43B2CuisJF0UUO19M+esHW8VyB4WKCDanwl/oLxFST2KIi
MvYms5k6WPOvheWxbk09Hbz8wH/AJKXqafcDZOUJNTPPtViYM00///h/jvlckN3Mo3egjCBUdZyd
zgwzIM+q8srydBz8ZF+v3MhDpU3zPfwzX1vj/kSrUdhLqSyam8DiP4mVIVl8IaqhNFItZtCeVXvw
PX3aS+djccjG+kZqgSBvqS7NGjLdGN9xZct++lULWGVbIP8N+WlF2yZXBlo7MWt6PSd5WqPz57I7
q7QtMKjhvq8/OLVqj9vO1FUDOYOh/VRv1ncF8KI3pOKnOiETVxaiS6v+A3/5U6Ihjd2M6arf4RWs
S6d82bFOtqTbBJVL5eAWPzO9ovYYBn+pGvbFaU1z/lKtUAznLPtaXl72dDMGb0AaE5zOQ0Hp8CoI
6/VoqNXclvz1lPHHp1yNTdKDg+47U8NvIruzMCWJlEKmwN8OhMHZotFUgybxGCObYObi/061Xb9x
DPRaBrORUR6QrjY729Gq1sv0Sqgmc1hhtrkvQR+kiGRQiwawN/1HQfwq2Q3J2vWnUxyqGo6xgA+f
1CzFUbFL8qfsho3KE2ByLZPEo+rbNpYp7ZN1nEWdHfNgH3/LUveOBTGdYAyX3XvQmfkERsWA29Re
IfQiu6D3EeGmDpOeki61QGqMMdkZmdAXKKbcrYK6N0Hzw17iUmTLjIshx/O6RfA7D2keYv97VCVY
LmAnMyyEIHEQQOTOTkpBI3aNtr6nv0xZllIzcJBNSAaET/udlcnQP4A3OfITZJIDTr0mPH7USF7w
eWsB1D2Wne6mxzfsrF247LqaH8XZ3lUNoh7ybl31C4mgx45CWYJufvo87ZUe6qgKqapFZTAg0m17
6hug+92GtPPr8iiRPBeHhbkdsENtsBDS3eRlKtGau31ERYmoS5YFkAobba02PJmjbEXC4kt66Rqw
PVg0jOKjl25tVus9mkU434iKECUI4U/zEKuqcQbAHoRCPuZnvTKzywlaaT6FTjo0FsYzKEZ25Klr
439AONh3xpeeWB+vEKZFyR0ZEniHMHfg3h1x9URllO0uwiQqeMxTWamTo9JfPWKRHmNWGBU5WmGs
K+XxAQK57ejxZN7B+H3wD/Di9XlTUum4F09a3qrcttwPEdjBRwz09exn+vXORW+RQTbQrwvQzWeD
WiK9V8//4zomhIuFz9IHkt66Y+GfyCde0PBzQ2PiVYEyNvbo3VSjv9S+VFhAlp5tIKFsjE3ZyY7a
EPhj3CjDPoqZvnV4qRqcyfNNWIRbtafML/W+dLP1NZ406XKzA2eCmHrYhYmPyjGRjgnso6noaR97
6qocbtfb68MOHfKpEIEgBPUBJdYf83D8I1Gk7zE/mVxm4H+VK7UUC1UNgnez2UKtFs99Uxv0k1dn
BtLpV5gVy6ry7e5S4SJ9e5P0WRq8e1CPv59X8rb9oGq7qrV9KWzPgLWTVnQnlmqzEfVhvecLkdZZ
XX0amYVqNOuAgQlkbJCe7qvKzArqPzd0YS8svnoa1/rVRbQSUumKgGKvSao48k5x8LYcW/skYCxX
B9ntXzuhryeSYzUQ/XS5hICETmkND4mBTmKG0Yzb/sZ81KQYn01rBjvor/eG4Td1fUaN06lzMmZ4
oVf3BYCAQsRJFTEe/MG/SJHkQhSMRGUP0NcmUTlG+ReMvmJdRvleUWVL0itb4bgm+4AdE+IK3u9Y
kmOKeFnh3HHDWqhYLvG+PnXdwTXCpeTZdAlq4jehCzjr9vMPYL62sLyaTuy73JMwZFfU+BfOECUW
JncakxItRe4OQh+hR3hS6LiiBzUFWu2tB9sHevu/6lRu6TmTVfoK0qGUQcAZLna2c5IKYHxvDLJ6
whw2IPBQscraViXzx06F3yUiBajbeclEYAtwci2mRKDs/Si3Ru8eEleLX7RWOvKD3eLtOMgBu7AW
E1KSkqjgjUYiNj0KCntsU0IGXgBJzED9+bg9DP208jcmG49WI03pj5wJvq2OeK/iW/tVsXlj/v4f
vRoqsvBCogtSlbcKze3QyLQ0uF0P3hyDBEuJYZxNlpWpFQ3wktJNHs73b2nqd7gBCZ3chQ3tRGK/
ONqF8cF+qWlbmkxyFa7az89qA7gQtMGPX9WoQCOLTJq4ZkemU8rE28B7D++Xtu8L9Jox3tDymSjF
vAGpSu4we4BjLYL2d0WO6xoK0YrIowZWqkmqUhFedAPKsE2OqZphqdXdEx6Ms8qQg4W2vzDvfw01
mh2gEeoGCmIQMzQWq8Bzo8poJ+GvQ51J8Flh6YA1bIWeqNgEP4XNo9RnikByg0FNjG9v+ksjxdVO
x8vG6UWJiBw9idpzZ4J0kEEpJlgp/sey5x77VU1NU5HGw5LWFCsnxDllUIty4Y3EKTvsVLvC+Gw5
cTVM/wFivNFbMXvY1N3x6KgqI4REikSViOrr/tjv7F6Q7ylMYIN3t4o3tZW+2EumWyeLyMd3iL2y
zghq1aEgOMGxUHmc0aKcNQcpAsWfzSEk5KKjyqpERlBdEO+DPdpsGG1AWuqPCf4ov8V6kwJ/MEXH
0m2/wQ39sxtvcyqcqO+XftLirN92fMinKo22YBK0LelmIhmDPzeQZ9266O4qMoaB3AsqqaFlX78i
hhkyooY57HehNsnnifCv1KsbTNRMWPqLaYQdG7HABqZ3XFAvFEGBboZxl1jDtr9fM4oHzT5daPEC
1JDQMllDH/pQWjuBFKx16f0tz2Gn+tflGc0V645hF3Esb3m+hFM/0PNb4rjo5og6vCHreNcQeLNS
gNmnQf7N7JB46sIvFUO0/xPpfV8Nds6JMX+2edpeu5CzuGRCtwrEVussQOEnQcRmVDEyhvYiza+z
oF9IRPXgVJdBQ6vIEALywEXM93afkWnSRcsbi4+nbARt//wHaOek3COgUnvND99Rx9eTslhPMzGX
xqdNXv/S01ILjAo3DhcuYJxEPiH4uLJ6oSX9Z54+lHx6Q89yQf725E4XTkGrUspOA4ui4Xon4DWh
xcLL7jqzOqTjQPWi8+8MsYcLG+fygLgmYZiwosIrfhcMbWJXShQlH35zrFPjK7cwgeDMLAulOxoL
Ksylu7qe3s7HAeSc+CE6bm+pRuHll3FBrjVnjixuQzhDvzGdRXZvzxGHxRffK7rgidsA8/7GCnAs
1IqngsL7N9iKgy4Q4hPmg+ivRprxk0c7CiWImuTw357zWU/MMFkCe2F81whs2IsnQtvyGT4eiXOZ
RIPSDJvLzzzjJKqxin95bkc2KgT97YAfrxbnJSXsgaUOa4Zq0IwgzNbcquaNS+8ceBm8vFMkC75v
LR9UcZnHMF+zBsIi5V1cLhBPl8AB8tIE8ZRkELNZXUswOWlVVOOr+cTILEIzUYeOJlFod3FUNGs+
iq/lGcc2YY5ZVmejq6AZHVI9BS5gSHkmPCv6B1xUV1ijeUx9zJ+pygWGT+D/YqzTs/qjKrNDiIrZ
6Ss026XrCr1WWjm0ijsbhtVvjWXk2zl2+BjHE+p7TBm/sh4JInNuIsvLQjxIm91u2WY70qX82QVv
Xr+GXNNdJuPBlq1T/becgFUF8gBHkjSiajXQenDI2PlYQQUBl2p3HzpMksFZAHYpl1lWvsKgvBSQ
eLtm3X9JOZohnxgyPzUmw/Oh/zkFvJ8ChtMrZWl+sVovKfErtaGeFXqbqGMjgwmzAhrKSwelcn3q
3ueuyDWDX4rWu1MFEFc6zLAeVAaXXnchSKY4LuBAGztNG2mmKH7A5FNCEE25OgwgXE/jrDLLUi/B
TEGwuRSPN6BIsSSgfDH7xaVJxoaRiwpKtpFzz24fCDLep6je8RcesmAgMZnGe5QmOg5e/nozJ0qG
FemDvcFHuQIs6erCsb2Nlg2ZnITDr3TTJsyM+pkXUhknralvFUk4K+UFa4+3qxA0zgC54tjlx6CN
sN+u+3je9ZfHKHDImwaMVi7hlHcfC/bP9n08apQ6CmQaYPYnmQByOTTG08pOtE8h4bmebWCefHve
sicpeT6PZ7rJW1AcdhTJKM0Szi1rJ7o7yUD8oRWfVhCJnrbpfATFaqp7EGcQ1kaM7h0dLLIKCYfG
i1A3NFx+4zQtRu3bgLPon9SauNkOfrmXGpcZtvSkJEYXBc7ZCwsFc1ZcMY42sZ4VedVSS+BLvnjd
GEcsviySlyVuch3ibdPRMD2X1n8R5RFTZBorUDX31IZaBa38jTCmBiTIWJLwOghQd/aYZCFlf37t
a55VAl/fdIXJ1bVUwumgvJtIcSwQvqumyOPUs72DCCAMGtozxxjVQzHZklsyZRqSg6v8rH0jD1qX
05PkoZ6OJjkxUwrW8t7U6Y+DK/O0bSruJjWhL0WuPnF9Yw+Ko2tOJOAkX/CnTpRpcITIvoYFSkjM
gg+QsQOcyhrKFUAs8E5dGFEAk1sIO5OcyYxIjmdXRrKXp3+EwxZriWjrPco/4MWRnn03lq/JLRPo
UuqW6uR+71PB2cC2iibQ+Xv6UUBiJPVldn7BbHv9p49gN+GvFhE1KS0GKmDeCk5bpERw2Z1rXwMo
7JwC6Rmm7MwsEd4vfprOa7aY+15Y4OXavltMv/RGp7Fdo3LqQVkhRI0hzmg13EKHSaUaN+78Bnjk
bQ7vp50EYULRi+4ypsfQb3UaJKbfp1dkOcEbxyFJAD+GNtuGekuKqyXlhk1TY2CxogyH4OnRUv3h
mo8VIcBXZw0SfPvBfZHClmjXpatRN6t3G+HSBglY/B1zkIPfC8XwHEn2SojEpTqFBobb6gpeN9YL
9iVFrtah/PUOj7KvE1toKzHXQz2eoU6ZEFplG2lsJnZzRyPbiaZDqSdZZMRJIUscrA7AcPhLnUPt
PudNq4DduxqZJuD96heCAFLD+3iDcm07mQorw6tjwzuiY8NDbORsChoMUXsz0AG9vlflTfbgGWrU
ThP7LFQ8nqlnlPBma4ArYFU48bd8OxYqImokxQMM6QconhBKX6m8bYCB7uWkavBNyi0f6j9McZ4z
gbWF8nQsddfuFgM6OYAygynm+kcipGENVDbo2kLeuhz/5Juik2LLDa2TkOk7e2Vz7SPdSlL0pYhV
//c/9v7RvE5zTPlQtqVwS0wCX7Yv9ej5Vy9J91s9f8LPUQY4WHBMRZusfjZULb9aT0PSxYCodiTO
MOfA4O3ldjuSwe2jXbrMO4u/foguVy9LyMvRdHk6RvbPfyM8Xqw4J7V6WX8qUjq1fRUpRSvyEBR2
ZyLbgPLjQr/7MTMsLtSTpPDeHuhw7W4GU9BllsimkgWpiYc8hSyCTAOh7urT0Zia1CGJ28aZkq9h
DlbVrPbEYXOzqF6za0B/+yNs+uaUo0XfoiHKRtX9BjP0dVp/5feVALn0sJ9fFLVTP2aKE9/z2aF7
9oRuSzIKTwE09VOY3+rrGBoFycMZfW1VdsAIRqUinBQesieJusnA5z/Tec6ECojBj0WG+iR0l1jn
oc3r81lz+A+Si2dd0ZwI7mN4UT8zRicWMa4KOq54rmQ4a9KKpLoMz8FeEXC6zS9amoN3rrKQbrgu
KuhISN4xdOlXu16ObUMxs5eZimTYxDd9E45ae7mO1ayTz93jByLIkV11d9u5fJpEs3Ou2ApjPUXk
KDTNbYWWFvktKfIrVTbbLcHbsQqNdUpWwsz6PLRp0Tehy5iiFkmpsBT6IIHQAnJkJ0ONngl9oB7U
iKMqpob1tWEv+7XWo3xc2QO+euQJkw94lowkASNT1bWsPpADhZ6GpwilZpdJuPAvUIBUHyB+zawe
Dffd8fpHQ2sVNXXbn95qGBlq1kgVy5S4hBFWq8WfinItn2SmxqbV+dbGjS50umhy2mq4kTAoTEm1
qHHScIGPerbjvTtFyJaeyZ2K24Pd2kCm6gEtanWjqWpuiRogdvfBDy0rSFMmrGkbiGq0HrHCqPYP
DmkBsk8XYpXNTYVKXDmowYBQriwPODvaooDKbb+PjhMqObxrLZSYPZhhZPvNYyhG6v+NrXGUN7LY
0zp4/cHftw0NkCY4b/Giprqh8/VYmYtnCYR8ajbxSQnPm/fM+ALRP5LsNhZPO1l3Qmvnl1AeJxxG
wP+qcg0FucubCy9so4loVkx9osdu0p/Z3BGC6ymtY/2TPmvu6bl9NrUH1SlibgFndNBOd7fbkCjK
aIVaHuqfAEHGtoETQNTxblWru6hzHI/rqslp/Ouli6iaPWKl62rtNZ7R1tMjKkbz2jgtZu5jnUUa
UhhLIA9fb0L3izVq4yJv3ARYdN4WPlzxgdQ/1xoLd6zh5sSY9VwnB7IDAGeT1Jmhl+sG6J9jNpmR
NZRiztV8Es1LCbhkd5ijS7BrRDhY2hsjgFR3kDldfYRBgM5n+eRIwDOpYlraWOntyEsNkvdgVO0B
PmkqYnyYAEpyqb4MQaoITMS9o/Dx5Z8DTt3hIZaU/J22MIBX6ewc78sbYc1p0KWSFBWxML6vGGJ0
VUyvzdxBart/dKpGcU+c0WnAy5FIBxT3l+3laOKEVeapsMvpQfwXXxc71k0qTbCrsHTK9jFAVnCO
EeKoEr/GL32HQy/ayDI7FxAjqrykEPhXxDR9jCMOOcKoYYCq1QygxbKBNIlyzN6q4z/Lj4xBxef1
5U8x/6RlobesEfRkYp8RQs6AZn1j5V7gZpiBeJLn8zhT5x4jKdxZtSd6PuD5fRInJ7wq75QDQQYF
NV1QhnkUlwy2bbAsk7iVXdPoYoPn7pyE6txqBuKWcM3GM7RLzy3v97hJHHrSBbKrF7ZcNEqu7880
zVe4vpDOeMGnxFUYwpIz9Rz0hLLKvz+eEnazle+ZxqVvCiX7uUYQz28SpYBrjyVFbiFEJ9jdDd40
Jq6FvZcFlMIkH7blAgRxyXkT0m7Z+HVL7JKyS6lfqNYbCkg/VVPB+GCacKjn1b7SGKKIzdbPdLdY
EMMW/cqX/AQ7jx5ILJagC6Gvs03EIpeoggLrmoMxwb9pUjRxkaoKAjvex+rcvkhMHPuW0z4feALu
hHPElf5BNVKSrwONCDMNnbVUeJve/KJgmMHC8tnOs74AYLYYgHpBXm9r5nkS3M8fPrXrZv0qd8fE
I6ALQ5prtbPL7gccwVuj42mdm1nxgMzyN9JWKh9aqfAJz40U7WLAB9iaL+WngWz1A/s/UxvZA4A+
CpdO2F9SQwIbDGP389NmhnbKw1EI4GEeFfJqTPDvMhpePthtQaOxjuaZTrc/zk6PWC++O/F+Q7BC
VKMrlmYcWpkqji08KbcmPYDDGuw+qJvuybZ3A21PXwNqG7OBFTOsdqW5xNZeEVFH4D5pZa7i4SOf
+gDB+ImdQCJiQrkKMsV97/1ZMwE+YZWoNm6g3zs0xlt4RYVS1nGsP9f66tmsM8pfdWNAanm22ZX2
hoBBeuQtd6wma2Bz55m2w4/yfdCsCEbXqeK4JFchBFGv2vWDwr1I5H1Qi6jY2eY92OaL2rhcJOrQ
MyrqAe/7XIbkZZ3PUwUNVYSf/ayIMuiZyB6PCIOafi/KRrbYyckmRYTVSgyPh4sQZb2YuLD4GAGP
3s0Cz1tP+ndEJdKKdzGnFt8R24FkxU+uKxRTlFG3Q6Ow6OAycNt+ou8u43+d2PPTWO7GU6s6YZ/1
sGJSC5Ej9y06pFPJuipliCSMRreXVL91Ecxq9MehT3UDCRG7sqPsWafZQyLeZCDv0NvaFXdyTzNF
7kVS8RiPcSunAjADCNUdwZGzKKUY/D6hW4ut9j+KuyiLRECjCOMJ23NPitPXaumr+Pc7AYKznMFW
1WJfNoufw6qITBFx7ptv3TSdujopPMc3GnlE1U9Ch+bHszdYkwJHrz4vrsTETJqRgoHUwvcw6ua5
JSsGv9pFzCkASTMJiGWZWsvaclbarAtVq0qVK1DKxT/tiHHQ2ZImW77alzQ4HH6bVZU2fNcjX7Dh
ZST3lRLDElcp4EKJcEcxb8fJDt8g7FhXQ5t83otDGdvyYi4/hv1jh0TBFJj93H7GZbnOmCuI43Wc
ZC4JCDwx49EgB/szVWdbK823EkQy+Ad1FEmhUgzf/0xDkecAF5isUAC7smH9pDtciwZYLutpIFr2
cCaBigVxZJwNowZ20JvU42otzVR/fjSiyBSEvk9XUKGWoiz9CNKt7i/S5sunhut+yU+pUGM1A2Lu
j6yoVmfPj0C5p/JkyquFyF6Lb/5ePRmBeU95WmKoiVwzIiYwz3IJBtPrPLuJTlwGmMBsn11eOLki
Z+nQL/+wxn+N+I3t21hq+yfCrqdxh42YeXtomPKNCQVVpZvNGMwIVBeBgkvCnE0jKZ7TBBuCR/oP
lhsAiqfpSC4D/UuYhuUb1JATZfcI+4xCEijbKdrHQVN3X4SvhKXtNGwpf5LTXdcF7gfuNjzHwMBm
nVPjDN4auTH/tfshZqGM2gYmKbZRwVQiJxeRvemgNHgyxYF8Sfu5/LidDHIZLVbz8MJi7H8NTeGA
1VHB95AYsE8Eu8PoT+c/kjBYNt+5xrSPr6cHDUdsw1Qg6laSb1ujJosI3gP1NuU9ijmaWxwLTr+l
nJhHYeZmbQiUrE1u6w3yJakLoZCmTT6PrdEgiH7CCoDv01gWpb8ANifk7dJeDWFl6q/TgqsGjVpV
oE23YtdJXuAvI/HHWL4j4xVtdt8Vq/N0aDguHrb3JjiD4serR3HL6GVnHYW3pNuC7ugLCinOxOZH
YO/WAkhwenBQ6aZ0cMLkfPTsBti2Oz86hKeb56DKEESTM9hTZ7YL1XKAsK479ZjH2qnCeMslDYan
lQ5+gWM6O7+A1/vM9zBRpPqvj/dfsiSHuUhIu5DslEU0JXN2VnMo05egHIsDqPJqoYk1l497ZHyh
nUXiul+7TR3NO5CysnQ1HKmSAFAL7I5Bxkkzn0QccQ1V5sqvYHf25J9gVLoADVn4E9AgTdXqxzz8
ttR8mfEr50DYdD6DcSJmousckpP8LCP+fdNxIESnogD8i1riogeJ5jvnVjmnD5bEUcuuuOWYh2nU
i6ALPxUoFfeZCbL+fGYaGIA1I0UmZ6oSDCOR/nPDs193r2OhNy7eVE3lUwvBLutUJouNKbbJ+rHA
T8y+Jb7SBOECVSanBQfT9JVuLt+9NmnRwMa4JMvdim2Xg6UQXjHIXM2WIrJtIXEzHLh1CqeKZlGA
JfnT642qQo7BN34lTgqmWloV6MGO3N7lbwLIaQcwkTYy8RWxl5sRvT38+/1OgUFCsUifAMg3cFY8
OQL/M8Rnau2SyGTxObEWav9fSIAZPrdWVYWEAmBol65Ae4khhs+i2z4U2mxzp3wTPIasxwgbaEsk
g18SXd/RknRLoP8sYCzo9AMKzQbZg4rtqHbxqvZs77/jiQfNhXQFSykDmlaj/WmKoawk0prrjTs/
/xS11vvAtMDXTpj9+rtA/yT0C7vSxJAqit1dt7xIobQ1An1B+EngPgxegHx0DPEHee3FrWQI/mSe
5PHB39uYdKZwdf7DfQFWJkP9KkNCFD9owC50S7bKHI/KQ4/5ZMuFqxuLlj/strUxujSLI+Ugv62I
qCHYCUpOG5KxajuJ33k+Zjp1YKqEO0zD7RaAbN9yfbjJQpJWCo0GR/YMdzxtOytdtgLqUdf5B1IO
tMjBuutDVwu7pKE+y6Zcb3hJdUUkBCViRy6hSZrqM1Wn/Fz4POrPCgyQlz9yPmH13sO56zvGpndA
LOATTNuNtXwyd+4qQWORTeyIWjFLJbshxGNiCUbzOQ5v/1Mm7epeLHYuuxwGX3//fplU/8x45jcl
q9QgA47M6uaKUr55zKnUrrROk0nS9Lb3SIutC5mGkUCaBIAIbnaFrnwMHQ+8JS3fdR3F1aKkP1jH
E+PahYlV2Q4sm4R5j10QBf9HaWei6HTQIi/5O93mnnBN4JFP2fT+j+PmudQTjm8thdCCykSC6Inz
TWbs735SCIqkv2pWepVFUoow/HL7ttp2XoE9PeOu90IPFXc8jGW4eLLCX4FyXq6dbv9FPu0FzhR4
qgtnwbPoXL1V3HAjK1laqvqEPts+3a7yQwL+BvqIaZjETBWApfEW0ndUpHXbnOFjxk6s/+ZWzEYT
kJKedr4952dqZIIV4esodhZW2SXqt9JaceT9UXQe0XuBuPR0d0m2S1WPC1IzOQq6IQelzSj1bXzN
mmz1LD8ZQGhaHO54Z5wR5EaZ6+dVNbgqtEDFhn10aE8d5yPSf6V7VgBABdF3zwkCzcXMpmSNBLV5
Zu3p7Dkwcf7bigDNMFgxyKd66szh8EDtocqw+pRD3ONCkRc3SjBHY406s0Fcn72VqrKzFwGnvG4v
CmB1GrO2VSTxgMAdK2bEntd6PQxUPX8dd2tjvV5cFdU3NSEbXymUxtUHiNhk+C8U2XbvfYy+ftIu
f9yMB9AWMuDJJc6qGto4Mkyy3V4Rz1HEMFormkdqY0dXW2lWqJIShv+2jlBeTbQys/OSX2KYZG1l
KObwagzCqfQFQVAYV6H+EkS97gk9kLEkQc+L5mPlt/4mcWrnLWqqN7zCZstNR/pzBIfjXie0yIOR
i0kBHkK2AKgv58N8OdP+VxqtXWkMTAK7Uds+fNFCX2N2ZgtHv29DaEpapnnRg7XeihtdRuMB9DLc
zmqdFvMTw8RfIIywzNM3nGqbheFjBRixSUO4Em1MQWjViG+E73XQ7ZHyIEcYF5ze/YR+6aCZypbN
Ypt4Hg+PQSyNl91Is2A3IkW5wgLQs63XC6WlQaX7fakmgxIBw/Z4C9Brfhrjz+DjV/krSe7Jkq7J
PpXwiRF/KAqrdGRatQ6SEcPzJpJof8jv0dlJMOIrjAUvfxMsJZO1Hv3m6vhvmPu07XkvzGPEZWAE
i3IkjSJQdaJbM/e9MlRBKc4hDbIT+77r7KV0rUM3qVCJv4XAPVaFmP+MfCTw4wkikSB88fjWv+Hi
VdW0NoWpBcnc8mqHkbZ8Dap4+H98WSDmeKOj0lNNBPuhJvqfyBdhkgJCRgKccssPHiAbEplOJmm/
4gozQaKoRFXA4xpfcjazGFGKr6H2ZtkOtZbX8kGFk+9eTCKIPrtHLDgKceM5okcI1ubBCef3EZB2
6lozbq++pyhRdMUqOjpd8N1qBR34FF7Jhr3rHDomsCHiLwIoMMfmKTYcbkXyREYQWshnC+Qsm5fO
xmHhAHrXldiAAiZtr1iTxYufkIaX00pZeEp5s70PmD3uiae/y+Ru6yYzr1eSfB9rMFREn8zIsUQi
vQeHOfNClOW4gyihO7wS9E6KU5KzaRJRvXpNnTfWlRhXQErHJi8PCQnjHRMBk7eZHwpgUqUCj1oF
rToN4QqWq9pM/Q+6MEMOsb90r3iSWp4P/cX9cafvaR1ViPefUnZ/eEtqyssUptOcpyJw9gxpz+hm
izWMorTHN6MmFNj7FaLSJW9Bcn89GbK/zB9vs5qePNZwG8B7/XQJ3xH2lwOp7dXYjhYNOESEbwMz
pPXJZJYw2Gq66QBuvVPX7hyNxUCuf2FI9QI+9I92EGoAFTsmeohuLOiQmybeeX2HS/U/hBNJJ7kk
gnrtSRhev+8vjyXRcAADklg5+ToCvBIjAL0cjatHmYKajVhaP3QWZRuByKbmWKd2Q3oHmohZZqBA
Fe8tTraQJrKYvB+i2lkXYYZN97Rj0iMGYUyETPryRTwS8tH8scNkK67ip5kuLPsp+qND9cAoB/Ll
IIKyR2FkEJ6cn6/8sYEeZCoMqhUjayxwjWuJqyYaHnOP/mYvdS4ucVnvgID8DuQuRqt74HiCcxvz
NEqKJ7p57y1MZYhpxmiaKu4rPDC4yD8V2NlkAr7gL1wBR19713oPY1odul8Z1y7jEbQ+4IEdJzU0
+ojqz9zadgcgXrkbVOPWTizRYCJCy+W0DepJ6vYGmTAFMmZ+gb7ul6ekn+cAGVWWqdqKiZOW4V2X
zN2HDntqjvo33aWhsz0EGprfWzuUYnogmHgrp4yr5DQG/e4dGbbSXbWgZXAcVSb4L3fJqu6y3VAA
qTAcdDzhjVBCc/bqwOXKYc4Vbk8JJQr14mcGdhI/OrIFGWEItH/4V6p4DZKAFoVldeCvlDc/383W
T6onmETollS9XDjCkc5RYK34/LGGHESq7clBwo4vSxPY4xIBMcd531JIPAq0ew+dQIbt7s/9hkrx
SxoyEzfWUpGA3RaGjf3SmGHiBJlv+FNwKxcE9qjIUP0MiFrqhiQX9W3tmn8PtGRQ+2iozYxESlzO
22t3WV4TVpBHKefk1Dz+tvBiek3iDU7GJMWjZSJ9iZzxJAeEF1YTaH9evyTNRpO6yCiY9IMbXLoL
g5L5X4wb4TOl5w4yGvO++DfSX3IHch4Tr0oysFqWU/BQrEf9wxi6JRWoWUAPwhQWTFMA1g+wCBIn
sRHxVsm1NnCHr60doFOKa6qxIFopQthSWqKUYAnURdqxOMTLrbCYPp1/pPLk9IM6F8+/4Os1ZD+L
FnJzC80DAAH/8ypmshfSZ+Ph/17tGIV4nt6YOLlwP4xoE88hrGZOCPLjaDjMa0u7imbLkOstX8ne
PfpaVnmaz3UJ6Gxcd4YBucMdBiSVuK4NUI4ugHaU8QBG3kajq2Xk/jVk4h//RDz1QrprwR0lpQT1
GTbbS1ItScdEkX7j+oi8uUi0abyKk+8iZeNjNxtgYJOS0JEuD6jMO1dcqzhHFDOj5v2fYXc/AuDj
SE0agKRl6YZtZTFblEWKi+m/H0naesP+XVzt7Q+inGBm5ZjzNIklTJf4IAQK8Ene5RXm2COS5Oo2
02QQq/PODA1AekmF2EOVTX4DdIvD+1er8QxUj6L4RI8uXynto7NRfWwV5GIjb9a5YY1F9qhH3IcG
p3ygAZj/Cjm6qJsFNfO8lvDZBuD0ADhJcgMnvNW1/x8+I1RzmnJitzwpZ2uu96sR32zCuXQhq+g+
ndrRyqmDhnaMB5TN2ePDT8k2ET5RbrG7IPG5WkONACh3wW3TyTeUDrWLn1OALcUQHcSrPOeCT9jE
GUoZZXo/Q86+PqYLZQBLL13U3VCCfdusYwW9oLFn343ZwN52wfRG6ETVSM/1XM4IwkIL2eZE6v3u
Jsu/NkPWjO0rSxs+j11xN7mn3SB22CpSKJi9p+jx7w60VNvYqcluWA6O2iCOD0HYoFX0QQRODDCj
jh7XDLH8q5mkXYxEJM+hWyaIeiYi5PZwRSquvP2gWg0aTOZlptMNdGUpa6WUiWdPfLp5bFcvf9CM
n8wH8p6bB05UOobwLRw5/oBrtaillGC5cAbXXn/bhMOej76YS6Nu7ujp4xSszam9Wdf1CgQpwd82
7hcZ3m+oFW5EnmyXl4jYGcvNXj48Gf+0luUYI7vp0AwQPjV3RicNVN6IYm3//ETQl95Cr67W7yt+
ux5jPxEjHJUN/RSEdN4BNpgaeqpBHLZzUwcWJB9tyL7sOUQSLyQmNhBa3kDOdZodYWOhaAJ/C+kj
DUKgdWCLSgl7Aud9cstQdvULipRm4RTIcLcb6d3lrnDtLSn+O0YvkFE3NGxJiPL55NsAWse9ukKA
o5Ruhn13YpLqmkYn4q+0BjFAeBSimH+COrZLCIwdWDj2bRyq30h3BNePtYvS+0YLk6Kd6Qf0tLFd
VKmQY/szY/r30ZGDKIlS1sqh8aHQ/f/dUkJEVP4R5Z2wkjcy/Q350lSK9frz0BXBuiR3K6OYsaFY
gW7q2Y5xcerT2DMfcCHHqGWvVjBQy8TbmewUHEGsZ9S+2aMKHVQWGXFMqx7u1nqOwL69YSoZDCdg
tfH3IJn1B9o9EPcxV+jVb0HsO2JSwDgqgHi4Aw7mx6ExZpr3ISzl7WqmUO6UcxA1kAp/SG4za6GO
v1u+CK4e7xsn25MeqKxfhL4G0pYPCuNd+myI8Qb83HolqMSU7xsXHzy38QYmM3k0QWmg5gBJfGGT
S/+2nEqowMy44GjNidaptFLAuvzjHcoMKEKB0gIvgVPpzEDpUatTRI5lYvPztv9YgGNBMJHCS54T
e1yYuuFXQ49MESwn9DtkiiD5c4KzTEACLVOkjX2TDIDU3FUgE7kTdtzbGwt2WoGQGHcbZdyZDshn
CFeFlka3JB45LcLtgY0IYDkIkpyyQn9ZoZWVRDlKz6v2s13ZsptYMTGrd6+m6nVYMxMAPjhuNN6a
BNPyBC9tgsKaopYQnpPF6UeX2Kx9uNS+l1eumtfazxYec9KiLJRvy37TU8QbZgD1jL9TfhSnBGQ/
Ibw7G99EgxdsDiym029prQRNJ6LE//aFrNmY3mDQuh+iEnncMdPpeQZi0o1jyp5O7/xjMI5+qVwP
J/W6JbOzIYu+DrFxgRQH7Rrhmo6FQXCuFtX3RtmMAI6LRneoSsqF9srfD0oiT1nD1QYfwXr+gVD8
Lt3qUsQi814n9fHfk5OwGi4/dQBhy9I24MsbGOE8AjJEJrjOAupeVb+kLCFMrTbE1SGaMj/IeHnn
BNcuW/GITO4K2A9EsppoHBa7VtyR8TxjRHM+JIhz6UxZVL+ScXx2dVcnqjjZWm1CsuPMTIFEm1+X
ve+5XQrPJZdY1M5xj9pzo9gkjnCYfjdW7+qsbSJPOIrhIETCh3lyOwmnH8C+yUwVRmULDxHsby6x
7TzR2yPuthuRUlmEwKaIzGGDngB36NrldwrKCnPmdbEen6lauPZbJKt+H4zIWJql7WXtwsHLvFC0
00sYPb/2PhEiIKIuFMRhzvZ2fciVZHd1lrkpAv2i8KAjwwE1sKwdjtj0NukcvFgbBNve5McbXAwA
Iro77m9k6HJhqkbkvLw+o0yiqVMmmSNbRXhqxnSsGI4tM21Lcs5Rzatatm8pQzk1PMxVIyvzuwj0
N1AJ7xVPeMcUb73rVV/6pNhPSsXmBdZxRTprejYGCkwGgcmMU6bo5RH+FUth4eujXvyf1OzgcKPX
WCmI2luaR8S5Qzq8rJ731EDv+MZJ0W+4Js6m2tAlc5QQcYtKahX5YMIUF5tC+4u+hDMIhkXBWvNv
1GSbFsIEgrIXKq/GtDb4uxanU9CUUOj8ChXQa3/wkVyjjczonTnL90BMM8F2q5KwkBbe8kvopptg
I0KRCBUEGurLufDVb8zgNXVtNrjJZP7qRc+ZjCo+ZRcxTz27ITwA2vxNuBMUPAyPkWGso9c9Gf0e
X6/F/zvEfP1YAL/Z3WWhm6bT5OxHZu479bpUHX5WFhZJNNFhdtqY5wQHslaHNK7/8P6lg+DdKuLO
LLAq+WNZAUdXkONeLcJ8CHvkVXn60Sh1I9qymNpXHU5JtVRE6cnGjOH6tcqe5JUDlLFCzxRdivvL
2td/ViZ7i2vqiwsFu0d6M8F4iyBzHh0lIjYSQi21s59c4TCfx4xYw4BVxYfqxY6Vy44U2flRAWz6
K22O7hgV7crZ4K+rC1Brsiv9ZRqzMLdNipeJS5i8GCQtvfR/ntCRvJQlE4cIeL6LqILwghBS0Ppu
/7UG47iOgNU2jxnby6HO1eRKUH+2XT9utzXh2pe6ajoKWRPuW2BJkXs3mjWNbXMAlbHbL3aPgwbU
K3PGHeBjSWvLiP0jf3gUntk5x3kqeoq3gYoyQGy+8hcBZDEmw0BNPyKybYTIRbublKr//nQaBz9y
fgyjqt4uM19orDPKqWSxiksYCH9pa3V+Pw3TJjLfGcZRO8LldriHHhsv8v/h9P7ljG3j8kbF9hQM
EkkZNmMdHxnOi1RsPr5S5EH7i2rAXOIM0QD3GyDyrC86JRY/xnGSA7v5//rXLLO8XbgZEDDBZrVd
3fDSqVVHfeUIAzon6WpQ6v8InykXNvhX0GWXT8mESwhzsHlDXTC5jQVb/puuxiHqNLTixckBjLJC
0aMAQAJt75SXY9oxKqhFae/7gF4SK2pQKojGupMsGpqpRFPvFONgpW5wjl5F8mENdKCvTM94FXqc
BVnreucIhtNIa3q+WVq0DAlLGj8/1+vWXNX0GsWQyTIHtIJyixU20tPPzdX1jrIdheIRx7qa4W1L
WIEfZO88+ch3o0ahqZQDg7fV1LG+CeFgh8IKi6cCM3Ql8QK7mrFthIZPxPvstyXJN6paVGQB7qgx
3HJxbzvkR4iK+gF8KOYCsSgffBRwUxI0oPnOfG2Q4BavIS9trAG/5sRPH6KNoHAytooGLTaieItq
UzTM+BjEtKUvN+9y1stY0XruMsROmZcPCl0OGt62GtC6M0pK6aGAQz5i1MIPi2TgXJtZo9CiAagD
ZQk2vFVUBjIv50UszUvOELVSncvRVF/1RTzZBSeOdMGwLDjbSToCiKx6siQTxi5jrBk+v90Wm2jK
N+dd+RmDIhGiHFE7DT3GNC37NjvCjQ7dpL4UFQSAkfB28YO144nFZrIXkRqCLDAowr3ANS7aXH6R
TyS48zzOMU5hnuJYZEN1H3txa0rUsn3M73gkl50Yl9dhKo7nsO9Q66eR+MkgXWMKYO9pLqf62FlE
pMptWZ0YD5LA3C9uhUY47IXuNyjotsqdF31i35FPh065SdgEH/En1e8RERx124TVNcRadhet10ag
k+1o9QkwM5VByj4NTFKVJyvVrZb/C75RudM46WP1YUXaAZtajqfTfoG97TBO9KRmPXj9csftvHA+
FnsBgl9NRXk76RlswE0mcAz2oRLFRwa6oHbtdBBEPsRWhslADr6HP2F4WXJR+HTf7AWbwqYnaPQ+
vdWNEbFwHf7EvUt+0qAcpnRW2fylHXzu2RC82mGS/GFNcD7PoLAkAp5SxaJ4H9iBVfNgiR0c9YsM
X5YZIc8EZpBwWLMjKBQ7nRs4v9KyGj6qt5uq68OzgQkWJ/LOVFYar9pMTI+xmrIlU3lG5GEEKv2u
LN3dHvVN6QBhgV5T/W4UNqFi7x4YX/pohiiUI4ffiqULWw6wQzXFCNKKr7s1kiq21FcqLKXL+ATt
milMWBnQkYVy7rHDGTlRCTU5WT4VYiUezxj7CIhJUImY1eVivgIelVN+Tuk0ogA7hpSFAga3Bc8t
MV29VljymUlqLB9UCrRyTQRX9MRvgCOcQqZbT4s8fQfJ4meZ7592ayPc07jMwz8B0CaiEnc+YWHD
AxKbTHaYJVj64WDfaaexlR4JHhaGwHo7NgO1PMDCnY+BRlVA5RKj6EXModJpJYuW5sOYx5z9a+E6
BrCmH3MQKsllUVtMmi1FBfgCuKdMs7Pl/hpP91XOFtZcVZzbHFKP7VOEybjyWgoKylcVnASzdK8X
pEvVetcXeLj4AKqiqie0Q4/LwIlhqlRr6JKwytvYN3yERUDPZXmcINTrkDv/25BP0+FF0QqAvODu
HQwpxaRFe/3dRhcPh2jpA3QGv7/pCDOMsM/e13ewKT+XImWCyYb1RVydPjjp5TvXA1nyjjcIlBDa
dua+Or/odzm7hvuh6YnHHXIQeNjefhTH6b4qErEfBv+jw6DQJyXamLt89YPhm9Lw+6FHcfB0dwhv
LAr2AJeofjTLjHBfIGGHy5j5YNiXhMXFPLuK6Gec0sJclcMf1YPCMibICjZ9CWebLefOIyv94uA6
iNFzkuUgs45PU3Ew4vRpaFbemOVkBBmhqZ3HS9UFPgEQtIGmCXqoKWISpQuKA5UcU6l4UyxglUFe
rrzCd3JIBOs6mSsM86p1bkfjiB41eYtdK5diY56Z8N1aVLmoG+C4QgzC8pXuovwmXh+TVKC5UJe2
KLQDKLjlfqEU8bMjlTJO/W8kWvZMeLkU6/GlUvpJ58n8Cw53duGusdFHRlgYJ8slDmILdGZypqQK
H+2RMOEqMIEwNAva7QxMZKj23l198XRUrYWT3MyaHjVCCY7INcciDxT3MBarwMeFIyl0BuDkan8f
fUyZms2VsfhlXQ7W9VoYKbaFir1Sy3+qni6jwEoULTcX+/uZP08uFk00RWcI5K9WvMGrtYoCK1m0
XmfvNxHZ4RmaVakZ56FKxWWjsqfh+6laCU2mLS/MrI6xBytgaNony/WmXsySSw3sKLanVgpebgND
qXAvT7v4wKFVr4sPFKswHGc19QEZZQsKYGojbU9h7DxriM5RMkZFzijAiFMTRLCRk67D3yzy+FrL
NU8b1uXvIStj5hmavUHTuckSTh26W9GKP+ivWyDhtAqpwLs4kOlkY/Xk2I11lihwX1JROqd9zggU
p7YOILWBcIPZtwHeivljfqGhle4IRh4iVUtrHl8H4/UPQiiEe1L0u5DhvsWogq32GOKpbuN7CKA7
EhtWagSb5tJb7kEIFY7iLfwSTaXlgdu/5pkikyQdAF6mAICXbKZvbU4J+8tpZ5Gi7VGDIH0+yzKw
Xv14bHeDPO0sg0jlvJivQyAcZzphR3yvzI0vOZQS6ekNxStYUesMYVo9TKETO+ERSpnCEVdUPBU7
S9sk1viEGoAOlSepb0RbGRRU8FMhdO7SxjXvytrg6JSFkEkX+u/Iyz3L8wVCVSqrm36CqwtW/MFg
u3XJl6nzJ2+rsyqXEqAmub2BMqWW+X9/WpTSCt1mNq4+1YklJ03A5w0zPTmoM2PyCuRPc4AaxwWo
iby+KwM30Nyuft5iPIBXf3iXwoH6qk4XaWJcBXr23VCFKENJkG/cV3Iiu0eiYij7XPwNgaPP4Mas
t4u8BFvmtllnj4Jlhm00gwmAu/PUcvUgvJX4kkN+5XL2DT7IsOE9auTfzfZHV1hjBOpDJatndnAO
XFzopfadWKl/Pbswc6XfzN0OeDpn0Cma+F1kQKN2xjY5By9+zgvVxzTE6/Gya9W4U492V5T7QfxU
eYv5vVEl8y8Vra55zRzVe+oNRBDQw++0LYhQ6oFukv8QjgxSZj9PNflncg1Ho3YmE/+k3A2gEr6p
Kypr3ecpkhAYhX+q6Ul17HhzssH2IgznfO7SePdRqRqXpWrlcfuymxk0KYX9Juk7EyedaCn73bBJ
xO0iHkutzzDvVrL+8GwE/v3VmihPEmwMa1LTDa5Ml3wrPSF0nsbE30EOLurwMGehhGpq0yjtid/H
7nZzCSiVsNWJHUuNy0iiKk/k7/JCJS3XdcEGdg4p1uC2QuEntoUnrvTwA449kRf6BDdU2q1vDLe3
saBLVXdlXF/EQBHgvxdOQEPKBO3BkibYTgM5/2WAzzyVmBHl+GXa3w66POzh63NcHgfeQVvuHghC
7mba8F88+AQIU7C3d0g3OX3vLb71XfKXYBeq1tgtAvu0nKtE+5Pf6pMDd9BFOrs6HW0Y+2036Ivt
AIzI8Kcz5JqJWFho1WCYe90PaHz+dJhAtprOwR7W9irpaIR0fUmnvJX/G6ePwahqLQKL+MKIvErT
/LVDyORgWwqW7SEe6bN3F9q0RgXnhFOGxE20SCfD0sbYWbt/N8iwn8f+qgjgcvFz3GAaMl4Iw/AF
iOA1hFunue+Va9Zhss1Bw2MoSQ9oaWU0FHFHLST2aS0pLrFVMmaOW5JaZXsKd5Fbxpj8408g3l27
kOC0uxFTgBoqE01siMC4Bd8dygJgqZkaQoFZIWWDyS37VxOGDcvlHtue16PyoHP/Cd4IJQh0X77B
Run8CW2Q9nmrTiNmW6m/A+GEKBTUqydmmKYcVfOnk5bBsOgeS0Sqy8dyRe5OJdrJpRvQCc9epnJb
LEY68ZGNTB4VU14gpN2WFUeTaam3Sx7sV+IHKS+aDac12tf8PpvPdatbQG9UN4Q255luhJIEKM5D
C5eZyECbBUMjKguOiDXmMgEmAGwb7Akz+6z67FXsX3g4Jot0qvqFhqKTnT2zI/i3/3ycDC6jYaCD
jgc/CVY7eMyo7E5wsGptmafS54/5x7UfW0q3OL2wfTlY/nYGgnDe804fLuZjzvwfN0/BDR0IolRk
i0FxiSt6BRZj7Iz96/Eq2bm7yqE/iPCQIxBCDshaktaOqoMIJUT/60Nz3eHDUvi1+p97AgKBxsdR
4BlbaL51eh9Jg7J5XvVsboC/g3FPYAKU9rSqedi0Mn7g1QE18okD3+MN08kkBZrpUU6YZFRyX7/f
LDQOFNobCxXZIarF+nBGhgX1f3ulOi8tvW5qdCDfM3NDnl/YUEfyk2klCYEl3lV22Qskjk3DVbg8
unRM2t9OB44J+mO4Kl7xqBCk0OzrBXBDtIKZtpKWD0TdhUKU6B1uqdMB4sZvcpm+TM+TOUeultdX
UK/SFOSzs5xEDSbpsolQvw8f+7thTo+5Oi4NV+x0ynVJaHsKVW8YM3sB9Cpv8hUjBZRgqMD47YD/
23S21BP4OcwLNkXwj07j8jJeMGTkQMtyriigTbSIYOplpnFqQacQhy98zMEweglU6FeLAOorFuvh
uI3bapI3r25pk/3HpT1Py+uqOctC7S1sAUCAt/BU55o63bHoR66QoJl5a1SKCeu575Wfhr6kWTYl
Mr4qBHOXBeGY+5/UTNTK0Ap+MUsTna3HRR3jM5lGg92eRpb15e+3NawNf74jG7g0ADj4fxrewgMj
ed7Yla77vM1XxiveOXnaIJ46SqRH1pfqh8c6c7nSFEfyh/bVujhrUSfhB9LEs4VOQtmTgkFlstFo
+CBJcMbhw/LwSCT/XSvSoiYigaYR47c4mHQwII30fDidMTF9x9cgwG02Gn1oJDShGqcXMvJeuaWs
jYoC4hgSI/SSI9+zOhnHOvec2QljaGn6zyV+XTTPLT6teRu6scinHgLacPpRDGKJ/KyoEBwCYgXC
6PuRHx274ZQdeSsEuWs3AW+gpC1a5PdxtnCOiWpIohF3x6BatzCxCgw0xntNQ18eP6UN/iB82/IM
eVHwCdgqyOt2EkZUk66u0UmLEi5WWZbNkw8/+B75ar5dAf+9k6vKycdsblUkmQIpwh2tapfZX18p
1blvoVT4hybNBj0NTRrgyGpYPW68EhPG5sf0nYIUOfkf5QzcBNolnt5Wj/jdbnE5s6gSZri8vj+g
bPNMohhjWWJFuIM3ZqrTumZeRiTKTVjg1DSMcXyAKoX7lbKGJc8bPafZ9tRVhqM3XKnkVyrnZMLt
YO+45gPTgmwiFKSZVPMqyk/FXDNQEb1qcb85T/I+M7k9R7hRzJyu+/bQGXhGxXIIsga7E5BkUpWw
RYvX8mivmbL8zxzYb9ZIbBLiDn+8PuDe8qu0THSNRcgAUhtoie2I00VHSsUmH9d+mAXDVRSSkEyy
UCus4HWs3WWrHTXQUzitQPceJlxlCMyqUoBKjvBOGNfarMFyewaaAsxZlvR7m3s5hrIjZFkkjv0l
8vhPXMZueMOwDRuLFlrSVuAMDQTj9swLZBOCnavmuFpJoCvZ3jS7gsd1m6v0eq6Hsk9jU+WlJaBU
OTgg2psDB4h6XZ5yjQlGRXvRWYHZIkQ/IrpsB089zZZUjPA0a//RC10KvJjp4o78w4acXeA8Xr+y
gOnlVZsUe2+gSavo82NeXr2eqZfJbp7k6pU8peSnfYV2cegRyj7t5vK+s7CiobLoH2Zj159HiFpo
NfUfzHvJ4uhoyqPa1rZgBSkmp483e4gV/+fipwjP8f3uZWmHCBEpvj6jm4qRNw6ZFHOuht5sXFH9
DeamganooZ0ZykaQGhLECUs+eRfWrYCPijK16s4e276B8HB39mMM52AAtlyrU5fq5ps0aH/aUsox
E7OxWfGzEIpP7S4zUT4zVhHOXybcs+soKzBNgVHjuFBPM5J+5NAOha2cSE/7MaouQC3WfyOc70os
TQm18diYm6IVSAqwprciFhOU59ILnT/r6z0zU2vA5E0JPFrbeUmyp7bjHhfw9azuNcrDZxyv3OEj
UIahSzPpGSXQOxolVlPqWR/gNcqBExrsaFaj7oWWVA3tr3HdZZCSOF21IzOVHBaKW5T+Z6LogDTL
CrKVLLZb9PzZdvdqirBlsoJ73FXH/Oaw/CbGXW418RL0qh1lRyrBRQlkiYbAUysEJ2y125UooUcW
UQo5Gqqo7Sqeg+5EAd7vsPaZ9eM8P9nncnEKjb9LaFEpTBeDYn5F2Furl+tobeLH13EYlaUgPu2O
1KflWpsYLsHrobqc3yfgzfzbvdZZmnXpynboR19R0XEDBoi+ZpAz0e8vjQGcUi6IaJLZ1co0Jgx5
/jTQfqpkZl7Fv9mwe2tjiEUe7UV5ZvEQnnFE7e/kfavkPwWN9Bg9vHmMknJB7A+zGv+t8K/zcKe4
CJDspBp3W54ESSGMyoLttPbJvIHfc68I5I2RM1gjIxqyHraWe0zP60poK0rqs94LuD8d3iMAnmfD
jXD8oJkTJ44Kanxz/ADiUcVs7Ic2qZw4u57bg8eDKVS0Pos5svOgMv0SLwfA7qyW52lSnxCZRVmj
VAmun5VI04J2Hxqx4xiVNOMcxtXbfe3sMF+8B7lyhXsnzpKh9Bl1NhhLSPhD3xa1dvnK9PFQSSRY
uMQ50+MJrqGKGVpyKEpPAm23LZA4gAyrNnHGQg8/iw6hUXVlgM9Aa29R9ORvzht29BfbVMG26p69
cgKQor21+1JtRm+7aOg7iy2uXsxUVHQbpMjUcrF+BCRfImSDA2J15DvrBuGX3op0PP/oyM9ycnRr
gUFLB6m9uUqtrXMX9KBfkGg0HFRCzxskOkWX4KZTe/WooaCGfb3E9Ignhyn3DLLtYtrHeGzdjJg0
zTxExfdJwYuQQj1VnrZzMNuaHIW980rHi6G7eYtRNr4PK8GgN7OasWHlXGUpeoSj6xEOIdlzQm+n
lPHjJvb8bgiGmHp8dEf+ARqzilabqeqKqRAEYDawdTmObn+rWpirXNl7LUcLnZNpJbSav5fICMVQ
fkqhCyU9jBo31ZUbHAJh9JsY9wtKU+uqa4SGJt91GAfaxT/N1HoeAAbsIVrBQa999vlDBhrW09mS
BWHTuvfRyPDIhRF8+ZS7elicd2+z7yGKuz7GvK+t/Mv9zWuN23zwJTTL9dyFSjQFOCsgjdAZjpxo
ruMASUT7LuuLOhWfS8cfSkKWfVRmNCfc6rUuLcjIW7EXds5ofajwEb4FcRSlQJTCF/Q9qA3cdrNz
XtrMBKugn3XOQ9QBh9HzxbU/OEJ1tAumnm19H6R9Cw3MWPs/MGuvtACtYF6aa1JlSDZDHg5IHRYA
QN3Iiu1OkKyAoHe/vs18sonor/GRg3hJemAsDqZcVTJCbed9RqmMJ3PLExFgKhKAw5B+0Z0+BaD6
nMKQRNo6Nofbj7bB4/T4bO6pYUFYABbI3RlaEHjTFwq43DRCu/Ybc9byf9k8xjTpb2FTKke7JzRt
DxTmRrwgK4ij0bFpQAbr+Jq/b/PPm1LBSmMgFqx10laxKnjUiMJIfcZ7bc7IQSmkieJ5nm7M3pzo
YqAFqKVktdwmU0e5HuNqC3gfiMRtvKal/H7nLQKzayBgI4P/WnuoiH2jR4w5anXTgFWw0eoejXxa
+N3MVKINdqwk04vkoS/m8uOi1ZuRIBO0ha5OdZ0VblmGMd0zmDdjA/rbQ6Cw2rJRa5BmH3qN3hJ2
kiwGUdXngPCEj2Jz0fd688c13YSmQhhTSGLwNLIo0dPqV3imt+lgTVynUrO76ACYdrjpi8WHxSKm
YWD5L5IfZMoUk5586F0fUv2CnP9LazSDCdZp/LFV+a6veHIqR1vFSGoHGo+RpcPkROvLS2HXtoGs
RwVtTv73d8f5lZz3j3ERMf5YEfj/QXMTFJ6lMxa/qdZzNQvOOppKm+JMTEdAzd3I5eoIkulJ+6it
4JtqJYWuWo6/SuStqUsBs1dFEdbi65kvg8O54JK3BQyalKiSwEwBEZ94xV4jEi4uB2a3fNHHvMvn
4OGkvfGybWpzYTlaYZt8YZCPjfU2BbuWouBOiJY5uaCWYScZEodhzvZf/QTz1GRpx+rqb64t9q28
QfsnA5QX5fIVp5TTafFlcrG5nf5CIceXJWL6w3jWBrMXBKltIOuPyldI4/1iQOEadfNGhmr8DZ92
TRvWb5WOOB1OeCzNFuQRKV51bGCbd+SAIkPkYpumzse5cCZ8Q0THjR9gNTrXvTBYclEw4wkn/xqL
wzAtcHLvvFzheArYp8CgEI+r+ceROKFf+7TqfuFA8027vf8scSa8ZCQOiI2cEJl+nAsVF5cPktpR
ybaI/JMZik9ad/ufSA6LV11gGyk2mL2Ksz2aRQIrlfllkKjheDCb3BlGSR1yQKBH8/tSKlOqrrIH
8TIa6ssHx3RyvNSr8slguzvyIfakbrvHIxRXL7nCn+lzZ2Vk3sa908hCejUhSerer9gvYVbLgljK
1URojQYxyiU1TMK94A+tOYNOzTbosxhKZF8GVa7ZymVFmA+B6HXERU2LjwgStyXHepmxXoInCjKm
2QOoDPpoeL6jXX1kLn6RYK1Gs1kIR/xiSl4UzEMId1+xYgRdUqwz4Wf6l4CVis3J0+ToPfEADFNm
OeaInCaJiDbPbBiihv5IBAWQwYP+EhlCsXaojOKLboM9CknqlKRKXuVbWunQFJeesBYCf5jyJaYH
PfY+qcYdyIKkdGksjut0ZVlwRQmAs+cMW8NEKwLwNJgtWUxpWM871wHDZYu5MhVE72MVpKLbDydO
5rup1kcfT4iWUO/+PnnxMjmItMPBKN7wf21e+kpWGIXOlRseSXiA0wfNb50CNcdkDP1sX/HUgGsd
aJkNc6T88LSACegC8O0VuBWtYggEV5n7JkxQqYwbfI1TQQjsSEcu+Hll1KG9ngR4CrD1VYFhL2HL
TiUth3S1p0FBWqroCm7C6KhJmyEOaxISLsKFRxmO+nger/IFDW3yNZbu1xlDB9N9CCxITY61eDgc
1tMtKwVvh7LYBSGqjtFpQZDE5Q+AvzINpx2IV4x26lv8obD67WkuDK4aaL09d4k5bvNt1iNynILO
PMOBoIHnIQcbqnB8ePcdUuN/c2rsWEkGG4mRHgY/z4Uybc4DVlcWHaJQ4Zl4bDJiCxHExkPkfPRU
B8GO2V/hC62iTcBcdDE8jmJBB16LdhN2tCAOIkxkb2HEy8ChKGTS4PmaWvMoWs6BtOucf783gPOp
mjtfqS+ICccpxIg3B2Fgm/c77OogWZVCP4UWYChKtnMvQCR3o9SbvvQ6P+vHCAdrfuSGQG7rWIV3
l3U4Vu4z5dLEUsSPFYgd1tQB/oTJAjI1oRTmN04wcJnwa469c5PuIEorWiWHKw8s9gac6kJBkEUD
tmSnFEbahNUrb2WhdbYQc7KVbl/CvZ0ViNHso+TYGQBx1tYK8kGY/SI2ndw6E7LEs6DPWnMQvFhq
eh22jVEZYbPPEV40Oj0887CIDmeuhZDX9Lfaoztr592NGeZDbIgytjBdV0N5irtSubFruLRj4vwV
abxm9j0wso5wSQUGGS39PIipoDOIQLjsq38GiB7yZZB3Rad75UOI1gAAuz+7ndZ+NhVSLff41Ofe
DaokAR2vyvutMUs+YsbxCx2xUgd6FXtlo0nN08VxPwHB8iBgKr57dfVnTrptfhnfN5YZaCkUH8sO
lLyP6S8lCbw2VPHx/DiDoyRkgwmemgcz7e4MDSr6q1AYLFTp37PrHmjXR+WloJY8q7MHcl1FP/Ap
eFPVVGsRfyrIjnqOBkMNwhEL9/COc0Qjey46zIiYqTBS+Umh3Lz91C5B2bZvswJKd+7G+XBpfRn4
UogQ+To9ZF/3uhfsHsSR8W3JDp/+hGrrNFgIPa13A16ys0Nr92k8dGDBHQPaYoWndxJ/oU55kjx+
dsscx1SGpjP+1Lc2ns0EPnP27IZYPhLZ8zEWaalymdtLafqr2cTvutnB+X+lKFIGy3DSBE5Ex6a9
R73A620q7UWPx8r8DDQfFp68FvkHX0ZTAsGnwO6j65Ph2Pny8DI10uRtkOxkR6eoHjSgP2ISFWnw
XmPhROJvhVytlnLyP1abDwn/Fjp8gLgOqfR7sXFi7CuS76nkhEbm7AI+knhptZ4fxLZPUc9RVvus
aN0XoRjdprjtfPoku/SaThe18c1vacgr3dhc/SgZ/x18KHZRRrqfE5sqI6EBFdj6LpXU6HzdfdHZ
eUqFuJ/ydQ4fcPEB4UL3hpNOSk3fnt/Jh6ThWkIEvcIroDAtldBhlRGuqgmifBDoGZiQHKEd0qMD
mrIQNZTwVJB5VsbsSeRl61jo/BGeL+hKUhKA83j0tbudNZruEITOcAUBfSKH5B5h2/xsQWRX6Pnc
CmrmjVvLWpuvScOfyE1QQmWKNb/K0tKZoM57sxU1IClLp3ueHeuZOIilXI4s/3vN0GguEjEmpRPd
deguTR+4Lt680AibJh5q4Gx6s/37absU1VPhtjEyyw/yWDCS8uWvg2g3+cOkmO1Rm/KIOUBxxmi+
edMSy5qXmDBEmdtMVkclcH1QA36hQzWlUFnbR9+9w0zqMQfRfkfU7bPcD43aFz7V7Pb1oSIOMA8Y
goafNeOqlQbskLcneaAyhLlTk1bR763bTgTQ/XuPrhvgFvLtAGegha6b/QxIYVndKK/OKxcsERAA
WSckK2D82JDrFdoDvv+k5JPPU2VCRx5uvVJPfWiUnF4YGlHCZ2wVxgu0sT0H8KSqGpDpvchvfJRX
vfMnSvVuKbL05SduWeXgCRSEC+7MeJnlOY9101NqOYvA25y2IknSg6sZSHqWaGaqT+mjN/Skthzs
LV1QlEXduEZT52ZT8DHTPAMXbP2Z4DpBU7Vfb2bRbBjW/zgSR0QvYJpmZ4mJnL28dP4FoO/39vYT
uA//WxFQz2iUVZowEgsfb3azZYk+2INXDwnA1b7OFzMpZu41gK+VU/rMyB6ltxI0n5lVRr50BWTZ
oRiyHz3WnRuByxiz0XXS7AlDKGDRav2VQaKV49XyKlTPMUNHfkQIXaj6kYpFmkc6qoxRV2PAxrmQ
EPrNDE/7fFBmJAK12w9d11YxFvNPtO6JqVpySJS2v8t810YazYuar3Vk+U65fwpd3Dl0FWC/Hx/l
8evO+GHfjftBQ9wHWj1RvYFuCiE/N9r61+vuh0VYd1tBa1Rg9IKVYhkE9RBpL1st8q6fJwxMOm+H
JWLciHlrHgVum8HrcORqA+tooDysRLRUqCjuCsf1ojlSVp0Xjdk6O49mEVAnnUI7pemG3Pt5/6d1
ddJuJWJXuJM8h1jhUiS5RKJ2PydkTefhykHdNKq3F1n+RhucD9KwqFet6tCdgkQ6/+2E6tVTWHy9
Oru/2U2Fq3tyj08JX3C4dbCSjz6Pdsz63krEj3cQaI1yqwwRTnsBHisrJ1ciJ7iYnCxYKkO1RzvT
HoAtRErfFLMjZJ53lnbZrsB6v9pY0Y2i/6TtRJadmuuIvpcB2F3I7nCrFyvHXnAhhkeMuKAFulr0
L2toJwgtLxvufEyfiAVzpC1TKPqU22epc/NU1cfG4x4iAYaBi7iIXYFpsYg+jWVzPDfqN0mwwu2Z
dVZtc1m5KnstaKpzOrUTJGOKjoqJ771Xh2MQXR3fDAuv5i9vB3YlU6qvv1134zKCJTsT2WD8HMMn
Vm02D4my8bckxj9SMaf05SW2SKMW8QHck7XVNVR2ZWMp19QfGjhN2yooatmCdqfyqeH1GSUG+DrU
1wTiA+zp4D6rfuqFD1V3i/UJw6yVFkBSMGvkBGFigufMV9awLV3JtbgRZZtJKQb0SK5tL5CqJOx6
PN5N63TjBLxWoASL1ML68MbOg8nkX4i+i8Xl9me3d4w1NuP2uveEXMnc74bWVb5jHY1f45ZpNVDv
HyGfk6cIm51nRXbP38hsWZZEwjXYFtm/VpisUnZqYcm7JyBrceNt1iPSCEue6dOO+AtRiawilyri
jTP5An4cuZTmZhOeh2ncNLn4EntTClJIgssWd0SSKTznWihKkMr4TTSKIajkfufhTWXq1GshjROi
A5ZXWrTpesU6Pr8J+MYnE/+uRG/Hv4BxsBDUu7rYE5/JQew5V7QzUB1uPs0IcFaCcsELeyvW8m8y
DZqjAZDfKBaA0WzZhiMOUa+CZMMn8zjlVnFyQu8hbrFFNTqu9yJXAf5TBaQCQo+Wb4JFKBHuKBMb
zMlLDryucrMUByGWwX876Bre3eB1kKmi1cgmUWUV7c+0t2dg/OxKw9oBGmWjcDBOSUi/OSJW/PYC
8SaZgu9AUfyxi/Lm1nIgG45N1MZh5PvjJgdJPR0vk3V6nogGmj9bBEB+mPekvaQnCp7n8grER5Bg
+gdjlj5UMz02W82iqRZWQGv0eiMsLisg3mcCw/YMfv3mJYOdtQ4GPkZOfuOFB8Rhn1LwO2Om4cDu
CupurjjGaxnaj3IzYuv1VMMUH2JSJ1gm2SnRTOx+zpwKx4NFLtcRlOt+JeDrrAaunKMM42NvINYr
9IejFkv8EC50PjK4E8cZtt/zmsMz9IRMpMnpb2NUnAXLx3+pnTi7MHDtlePRrahW0jn2BQGQnksq
ZvnP5iCLSI4tD2UiaD5GRy7P+aykBdH5pEE1gCqFz9WV2sKaaksZYLbxN2M77jff4IJIvyR21LEK
JnQhTeKG9oDCUQwTX+DO9CPFQ619lyCuK9oTxDETOMgJkAvfCj6ERDjVik0Jaw8DiEluyAFQGnxz
6AIlWXpyhFzg04Q9i/Yiz8kw5Zz9pQhTgZDkNzbebZoQ3LyoMgQvV1sd7C5ZC6jbkKe6qk0gekLZ
1GASYGfq+dPz+ruamA7qskCNGuoH/vab/peusJw0fsoqEftSUtRMqgHrDuTXujsxDdza6oae6qfd
J+zIvu1XkEHcM+g9Sp1dgI7xafGrbwW98pk0JvMmSDGq9bkUqFY5A4nwa5xFu6sSyuSILJuZc+iv
OgyJFNHUOgbFn3sJw+RoQ+elnrAJt3DjDFDRIsrlC9JMMPmHKv942XlAWVOgkA/tGoY0C1Kxc+7B
1uy/dhJL1M+Fd9GwNE9EUeUD1W30dkErsyarMZMNUjkw0wDcR3ekdngV6U7XMk36kcybzRPLnbkj
TIpM6KG68kLaJpS9oKqErXdP2sHMok+/oCPJi+yElmjgI/S6eaoNetNCvjHplgZEnOW2di/gyVw7
C9D8ZUjBXCw3UB+A/tdr3wzcLst08mRQ1pTde5q18D96z2oTJgQaJtpjcLBO0SWMWH9syPZT8jUO
QVULSL+TahNp68kvChFE2QNtVY6Ik6UoZaOLxzq5g/F3NKdSTZR6x56qRYEXZ81X7u0ffKDutBt0
Tt2UoCMwHPbNjlUR44WtehB7x1xoR7/8hecz3pjEw478ErgS4OAN1+0ctcdKWCoCJAfcHWiv56os
JXB0z42hzozUS6WqBfwo8c2SPfYG8zRDt9RIZOFJrmt3LP6OYgeHFPxC6L9bfivjDP2D+J5m4Qru
4cyf9Cjoe5iFHHKBDqXcnLOdEgQK6lI8/SQYFBcBjLqzN8CkDcx8GNdTOee29Ko82F7WBQiPWiUR
MNKiv5nCCF2EeKQmmhfKkRggj7Bq4wpepkNkh+h4/aRfrFn+ad028fc3SXSejsGeCQS7cUk4xcTJ
asR2buYTbwD2B8Y+/Qqm2eY9lnfIfQKeVnCdws5Cqks8nym+jYDmhNajOXgBZ5YpVxSBnEuAnRPU
dO3rDBWDC6+qh/xHOOCN8YisVZ8v48hecuh9afS/dHYZmAWnSCBuSbbdfAih7Dd0V8iecoFSRrVF
wRKSnIKwqnFxD9IjoYTOWhFx9TdL4ZqP06/ZcLFG05jTwgBdZxSZBPugvbey3PdDBaLqjYyPhLue
e4kBRlqmGbQcOQANKlfAYbIjg0ZmRrNBP9cQqZ61CAcPwDMf+XHNI2D6AiIVxYOc4Q5YPT7j2CCS
LCLJq1fC7nlq7wJqD4Rs5/+DnRmf+CLMXx7OMBnRIyd+wq5a75ShilTvVP8XTnn0Y1AkQsYZKmG8
qhQFu0UM80zQww5Y7ZgKaL1Tg+O+zpvxxCteTY4wgrV5gbdSYHwATnjxKq7HGeHRnkMB5uIfXtMi
cvAXTRMU6j/39a5LHBRnXEffs5pU2v9WtQDzlz5ewtZhvMLWlAqVQ9JHvwcMudLnL9x//1aXhKUW
3SbUKEtcqyfjy8y/2NPcE80R7BhyCtg5zyHiN7ZHl6jj8Q9eMlATK1tWGGHgGkKwcs8X7f5BPCBC
0Xh75gfTJEivD3f6rHaVgXPqJZ63CpPJ7vOjRIb/893p/wUSfHc5O4kv2wOqH+qG/90aBQC7IXFw
o7k6m7vmS76uRP/ASyPRe/zmEw5UPTuiNOdG7mAv86EIGGaUvZf+FxMtX3L6IfW+MpCjdxOEO9Mz
ezrh2h3yei5gkZY0YWATai4tJ4c+XgVuLbrdysL43J8viWzNDqDtE2xEiHF5sBxFD0Kn0pmyvPf9
NJ7g/QwPQl8Pe+yt/sQiDBj//RdEiPF5NX19Bv7p2B+avQ/BHYuXK2ECrNl9+H7DNtBIZAH//bed
L7OK0+GcPD4Csv7F5uNFHJmI0tiyBgy2pMUtXhTlMCTpqz/776Zn4j+knQ1LfTQV76E/Xt6X7U6Z
/INduaDQXv3myA1Y/iJxmbB4SNDJJDdpzQMtQTaVzm+BRMGC/9VmAiZfOrUoLOLAZoJRgBEB4eyO
9T7qYwYy1WqadBT7qOo1UIT3BhNqguXotpGsymsTqOAq0kdnUtW5309JqPnGls3fkNjX9RbLiysm
sGXEr5i9qSBQSruSYuSfS5Y5LlmC8TO+FkaSRs6jAPWpDS8tcv+R8h03ENNdZLUvmw3n8gSsz7dQ
Qd9DYwOSYT1D+VhWcIEoS+kByMIRFauzium6xcrePoGqiN5AjQiyZ52k1cU1givDr74VEyXJSzoR
XwahOfKIRuPyt2rM81wKmGGuBVF1wsJVH9hhrpIIKJ/ALh4GP+mMP86u1SHkLSImVZTPsn6ae9ac
b3+xl7Kl4Bs9R0qnXm5NpP9ou99k2qEu0ckenXsxc3ITf8GoHCpF0LSNdhBpsAlmF/UYUaUoyMi3
VPX1u/guxumPaaAqcsH3pxWoioy689I3QX5i2U9U/UPq6kz15JLzD/aZWyn+APxEfQB7PKBggEpD
afFlM50Yn8pWImEt60qrq0dxCNcqYCDR5snAh+BL3SKP6Ql9QCk7lv3mNmpk1KTpYqNkS16PargL
odVxKcP+cVb2r/44Nd+TiJ9epfNJt7pdwZ3y+gDRvS3kQ5XPC83E1H/tPTOezmOlBvnm5lkXJ4S0
BXSHQXIkbomWd9MzllHcdnWDd3+YRsoUOitr5M33h975LZKBUdNCQZf+FwwUNWLiobBnXIgnEXmB
udTWDMMX7G+BOPQYTMDfqmHOCL4B4yabA5NVaM/yMPhEqJ3L+gY8Wj4/U9baTATYMakNLpdFBJSV
WN6JlStq/WyCZUzPmi5gub/OuvKIWWn8rDrOwF0HEDohaKbYJSyzkIVk6jyPngUmA1+g6T/WBdVl
qxVTawiSqZivNmRoTssQth2RsL9u3hMM/l/C660IULX36DCqCyu/4mhsaNFmHuwqDJVtWuJXYwvA
8eznnlIyGAK00pugVW/ahcoY/L9C7yVyr3v+PqN2DcwTzbb2P2z7FhNKt5zpqoMUM8y1NlqFduvZ
QdLsAy1q7g+Gp8Hxf1R+PDyuwZIEX7fuUs8HuCRMOuics2Zz+9xpUNyxTthQQoHIsRpdnyXx7IiJ
fGnewMHewODTB4c+ziNXrAK3MdvvTikHZ+Grv0CF+UWUNPrv3jSh2RAFYe+cpejR3NrcyX8Jy1Cq
xpEURI7we/B1c9XcocVT2ppSyXnFZriKT1Qc6gn252OeHHUuiAp5L2z/Ob/UvKR4mFJzEHvfTmKe
8MX6/1N51e5ICYYKn52C2fXN1/iL55puC56khbYPFg9VsrV00ZZUTBvp7rtLB1yJzA4klSDlodPu
Qv4wqx8U0fIUSiXXVviMB2UT2MY3bHAv722vMiEjNnnCxRbREoDo6gPgC74R7k9F3FrDtDdhs0a/
L9fR1sVqSdyVVRG7OCY0kJYf4SW1IP7HEAYHO1KJkBxiaT9xdAueXBRMo0QvpKW9lBOsTgNNU9aJ
cz6lj51fodMm64+2skvUfzOOYnfXzcVTDHYKFWNY38aWQ73EecRGt1uGmMoXk/q6O8xQuuYLCyWE
H9wuueOJjquLSpEX6uhdyuGdx3wKd80W2kFSvkLdPXRqmotBw37pnZN4Bubf4uu+eDFYDVFW1Nt6
vryXZvjLd/GUwYJIl+seivtYl1cW5g6IBySaTaBALnzjLRKXs/DsbNqSBNS8VuJDALTYsEww8k5O
/dbZKqU5RfTdYpDAvmyMv5Caj+tsF/erVx/qGaLF8jqXYLlcz4+pox4ALythiFmWjIFFPjnaWgQ3
OnV/mFkoXkGwSEdq1LsjzeNdLy1UP5Y0CWRd+lKuQ+blfU3sKZ60v+OYAkLRQkYHMQYXpRs9shnV
XpjYAt9lpWfIx9QcksT6JD3PRoLk6O6OfCSyMrzpUQ+Dc/HJL0RvV0vfN5yDEa/IOwjzGlpNkp8m
rxHcgH493o+GIGh5bYdQBRpSwsAxqIVhgckSBB3d5OLPa4NN2A5qS1VvgCdMCuDWYZcABeFYUuIL
Pya+sQm4WNR0MnmsRKNki8eNF0iGhNWvznYuBxFWMf3cvEdxVN1VSy4QHtZIZ2vVTkZVcdDSZleJ
/OEQiNL2RySpd/2RrJ4dWSxEqoz6osb9DaPninbQguvTMoi/dRBYUwBI4P2ASYdAaJEsZmHgXqmh
5X0vrw1bKUfzGbl/dhRNC0Qft6ttqeT+IBaESdoiboeZ/QiXlrQBB0anc04b4EUjiZC1gFA6+tAq
SXoqi8DqTyZbLgrTWfjm/qCWZ2nBjtsdehLEOeRzKym2oawtLRp99i5G2+FvSnY56DqNNVM5Thb/
1QrnwsNygP45eQwB59MgwPoIHsFCPJUWA7b8QLJbjwRddACwdhYgsUQHQxs3xg5uUcVwh05Q82CO
HGbaHEQQSgzluVwAReGyzehYS7gsStEKnNmPKs6FzAfukq6XPqqZXT3uiEYWUbY0lxhL10RSdlQu
KBXO1N/EJ6+qwSXblVPPyLYH7VuzebTh4tqn+e34Ro2Cc0DAM/SiuBgMIGDvPYmkknn0S0r1Jnsb
BQJdujHDliqKAuA+A39M7Pli8C1Wg4voW48V3mwADRoTcOkmRsO16h6aGBf1AqwARFwWo20VtoTd
mrjmJ7lWVmYW2q1wXeM8YTNtfTS2vXTWQZF2PBzug4Ij8Ri9Xsmx35KcMWlAvgowHRZdfiUDBTtH
X/Rr/HAmiE8IfIyXyg1h0WO9pqTglt1NK9OkGkRPuoNedp34mTk/WqJkhZMM1cZVmJ0cUCNo7363
EBwYq26KUHREwER8+7S5RDGOIkSej+g/Qeco1QkQwTijsMeaNoNSXK66FK5ZYl4qNY4FT6faaUXs
ShIlX5GNfwWdiFyNvEMO6QEFjH+14/D0shfp2ORJ07oPQhTOm2v19YGPpCnIIohXKc73Bq0rdVeu
2Eo91gnRKtl5XOiLeyBY0Lssw6KlS9Zv8E1dzg/zeoNrQflVqQvqHmYCqkeHU90ja5ucDaH/rZlE
FGzw6o+kvB8mpZNomTjdJJkTI5lKGYV2ro7oPaoEu1T9QPjvS+SVHTk8CTkPPQ6nD7aE77uSe74B
Gn8BQ380G5yQEgnlzrBW/eOwwqwl4JFlMfGEIlexpGsM/uO0evvZdZohMCLL82B1qao7wghlEunr
PlDVyCQ2HVpfVs1cnicK0Y9tPpotdEcgpH7ofEPx+6NNdLAKJacDGGw4DWI/vgpD5vee5RgsD2iY
xnd+r7bRq9wHtT+Hd3GM230gb6yBRlUYuo6cTnLOZWW6biMxxeXMHcaQOzxpkpxQa6gtOZdVzQZV
2uxiKJzKa3Gy7KdupgjMS3HJGeIsZDTdKHZKEqhKJPIfi/zTiQkau5YMkqeElInI170RgekcQe0H
dg2ywP/R8EacF5tMHBed3/ICDPkw3Su8Q1RnEYDgA6SlU7ENtS+hMSOmgsVa7mXozsBgvRLz2uOk
T0W//fMKlCPJA4icVpEtIL9UGGIUGvcy/Wa3LJOhf/7OqCH+GE8q4cZTpGLI0XhrTfu+RcXYZ+p6
sxjCwrSQbmJwrhFj1jjQ1nfkMS+2qlFo72VyhUtVAS+VxGyKcJnlw2DTx5TAyC7AnOKAozxPAumr
GNr4kNiuOnU758Wj2tAyy04mlt6dIa2fTR2JwXVF0G66yiYy8ya8jdezBEi4XOK0Zq0h3Uyg3TJe
Yp/Z67uzBRy3G6UtkFlA4LvredeCG4TtmIT1ERh8bj7lvx++9uxRnFeyMF24CyRt+m69p1WnNXPv
c2RCZxmBTmvrD2iM3UW6q/yqmvDzJJWmgEqaguo7rN8/7TlBm/ZfdB9typxKrtuonfmh6Qa47U1H
ywhO3NL0H388bQPvOxV+6C0Gmnbhpv08GF8CK1FyUmUTCLvDAPwWO5S2bvgEcKJNEHVTQbThu3E1
Tqw+cF+zIsjgLPD5+q+ykguydR24Age3vx3tnEBM9PtNdC9DqotWubIYG6sPK0+OyFT89lX3n5zw
xM8u+DUW5FdXs4kNrSybSBg7fNXRhI7WEpCqiL/CEJRZd3cWCrdb/XjpKDgQa7ePtDCUHdXVf+We
PJCN78rTdOKYDyNY3gfEq4Z/bZkWDV4vK7H9Ef+pD0kv0KoeahWxrEuTcpNiuxIlp2s8IN5nk3Rn
HfGjicCCe92xToHxRdfWklVA1OZHDEQb7i1QT6nkLdD4owHRXeufb6Ot/nwcorzu9OqvdfQH0Bke
phci1rLRWm3ljEhbuloJyi1g5Oqwy3V5iMZgKWH7AFWVcVhIDDQ1SYLKr0uORRVU6wMW2F2oITMa
HVWmWiaFF+3rJTl57KxqotcKbTX2xyV8nanaw/v+oWvZZ0yMArL/0k8gorbVYku+HsOfQWMTOTGg
FfgUudPMfrMU+1a111a5FcyQbOHLJwpIRabigiqYEypY95fO/SlGeJXfUlNNFNdfNB+bJ2p84uQI
tY4E2lcmP7Wd/FM+iI4OpBLn9+PV7L4PCehp9YBp2866/JdEArZwMIGl7NXWRH1aufqaZleUQrlc
+yYLDMOCGSPBGpmzpv/wPn05aM0jZqX9R79dn1/tcLk4fv/nGITfk2ojizpCcdT0qqz1IAJ80nI3
TDhwnnM5lw5SdqC+QY5Koqfw3LgJqBU0IKbkkgpx7Xwtazjdy4sHwfbz8HBd7focT5oGJjunGqmq
oL1zM3eHuRHZQl/6//s1xTJ4WpQ2Cds/GWP+q/mhhr4r+ld4Ri0lWnkFmeen/3/oy+V8bzz2xPRo
/qwcfG7pwxvwiT2t/Ot9mFjU/mipuhfZrxwUtda3Fdj3C/8tXc5tA9zHxPvxZkWE6vwpJLjDuHkO
gO4l4yPyhD/66cUiD4L7kpmPmPeoRcqOIFBktl7602P5x/j6LQOjPc+kByQvLGZVAFczNFcuNkmm
HajW9puWmKF0IwMymJA6kUoY8GW7ex7fZu8owKDDDj0trnCYKhF0ibPJKpkNUJaMw1p2GQdFTeNW
9YYPf1uWqc0ys2MXyj5iVqfd7c4yOqq7YAFZbSZ4F9bwfzx8g7ERrRVQPx0TUvOTL2TKCmPCMh5J
oAZ9BBuWddrXysI6JR4Sj5wk0GCbUsXdflCbHKCKD+2aZAHzCzyO6fsfjm/QveAPtkltc3SUVsHM
7k+hmLCKoExn8oIlsRz2fRHgOgOpvtEK9iG1jGtOT4u8oguACnNPxnejNPWaQ+D0NebtbID4jt7D
eiCoZflX9N1bU0sNWOFtSZV12DULj/+mJYmbuMYJZ8cHsfpC5GiKZttJhK8CII9pnqVLIddbYC3w
hNVWz/Ji/IXt6UpmQdUO8vbNazUvzsQ2Y+SxrU6ENV7L60tel/Sz8pe11kGTusHMKHP9jpOj7Nxk
IXzH6Rh3i4ciqTZOV9miLNDN9mmooh6jFrRrM+y/sbl5FtGu7SJzyK7abbJmlEGt6NYdGRyEnayX
Ultx4uNB8kgnDyjUZRZvl8rjLfv0jdK181Q67rlw00GgsrTSrAqMJ0OO1lYHj6cpN7njrBIPvKgJ
ycAcOvlAlmZa8LdFLfwU45U4csChr5pwEtQtyrKsIpCjv4AseqsVE4oTlfRtVby39oNquaEBOvoo
tG8szUE62/u78mniyTIXNiZalMRr/LTZI+z/1uHTRJjVgNPyBaMKoGPwAsdukqu25DYtME7BcP2G
EmTBwZHUzxWsPO+Qw713DbXUiNOmOTIEKmyLw3ulU0uT+3xmkc+m4SCDqupCy1Nyu0rAn8m8zqEx
JjsgSqGEp+J0rWM8bRQfP1MtI4SiwriqIa6RFWJ3sfMv87Sx/y6AR2rlLyN9jwhXkfOmCfwu5teh
rmlujiKxhGz2eXdMM34bc9Hu2xgtlx4Z/vImP0RtpCXxT3TrYuBxRSYsPPIy7ldDkT7S6kzH34fb
memkRHzGogO2m8tTW2nac9SEKOzNNLhYM1xSlgm9WpHUSFs1bBJ4BNBj/9ZbuC/pVGYQjiaR3ONu
CTpYycLdofohZH70dzXQWEw6J8N6gUiOOiu51ATxN40FLcBTxv5ZGF/16HydL9R+6Dln3W8an4oC
ThyEf2MTjfZ8J9REFXdKOB+IwJSrmbt/St0p0KV8ZWBqYPV13YH29Oqo7ejLzKkjvLzXOlC74CMS
W21FmwzmJ8YI4c3rR89f0O60gfWhVPhvrU1mS5KLfcDqtNGeyibgZWIRqSDopTIrRJ/SRD9Q6Cl3
81fWBtH27mZ3oamzXbjSIqdr51lAEbCTM8DVqyvOliNoO8Tre5uSLUIyNKMbpctVNZTXvpx/MBx6
jEfp2dFX36PR4XsIChJMyMZqPKpyI3VmQ7CdgHxMJ6hlbRgn2zT808y4MJcChYJpawN5+/eLlPjN
tDDiGfX4uuTAznc8HhN4QLRJP+EVSkbYx/Hl7zmzuP2EzHJYo7dtAVmWSU2G+fRwuxBKvAVbmUeM
YbGrComSrTo90LgGkDBZWmM61q9d5YAFymKvrQrtItmQehh+7Lg9miVN/yGPSMmGQxh8HXyoEgEK
o5LtKUaIz/YNfONd90DuU/bOLFwZY6OdsCm/8jCn8JpDK8jAV6y8icuw3YDrm/rE6pvZD05r7rab
zzgH1ZU5kLta2N+qcWLcVXljE5S21miFpl7xwC8IwTvPi3OvByIYIz6wM/VOn0QA42ULAftbnkKH
bDqkAL+DD+WoQN3MEyKZMt0cFfyAMvWYNsur5j4GYYFwcHd/O/6tcxVqx5ePaCRu5YJt5k1OV+lY
8rm1qF7aZwY4det/47apbgOEQMbEO2KQijqfBzu2TFnazBhNAsLB4lmZNzxlUOkwV5BoO1hwdHvl
h2heXX6LVqglRgCtBImd3dTqvvFYQZsawhIb36zqJIQtmm/BFmMaqm+S2/9m+m7jH0/03rtWmldH
dN7n8nuU3oKnoipRmCXPV/Zr+bC3obIEGn1iaa02doRAVe9wiPTe0PfgGV6Na34QB0xfMkrRn/fT
JpnX8YeMi5VZ58mC4TKbwueDyMo6c8POynDDX/V1xbe3IFqHjEchzyH6n0FKL6SXc0hPMFvNDawq
v6QWCjto+iwZ2rB33CZWibrsDdQTJRkw9BzXRDcQ3poFOt6aoACGNYOrMGLBjs8A5v8FS6+7xEQq
Jfm0HKmzqqKTPCLwvM0FE+xB5tCR7afh+KIVx/98llza8qKh68tZYnJ/tXEKpYo/nLU7Qov84Jyu
7CeeKPY5v3qTv7/7FyasUc2fO7a8RI9fYESuBvKJiTFI/5YsTcj3lqncoTNUMjjPsZ5M41918ZbI
ki7EYRaCljowTdc2k4twU3DthaM4KxRk//H5AZFUHxKqHICosNSXPV5VBgIaidxF4kWxID2Ni0ew
oZLGpVq8HBMMt4lMBKyuVsG0eKiyiP+CZI5wUjokfzpqHIxK9Jb/kOCHWCNEKgUAOZFC/2aEnSNC
L47h2apnTaXWJ1jejs31dMjjZKVI5ue5hEaq0lHo5oZlH40vAuSAlCF7jWOm0UwBp9j/aFYl6IWf
2pDFqqXDAqNkJclC/L8xa3c7gfR41kJUHytf4yw9BQW0lIX0ZzZn759rq4kc5XmSkE+V0hT5mm4J
2eLeay7tUluySeOOKsmlJhrpOmq1ETXsYCduyVdZ/sebqlJ0tjw2P1QPOEid+CvM1Bf7/PLkh6B8
DbH6ryozH5Y6pMT06HzjzFPjcjtquuZ98k2SFNQQQBRn1VlVdnNkvte8Ml5RYrMWy1TxA7PgWnvv
iJ/Y4fdTYrWdjiex68iY1Qr/Pt57UgPWBeWDTkySL33Hn3pEHIFXXiv/5D1hHi6NYr3wuL5VLspk
AXJ0m1DxE292+UiXCPIBQlKMzScGnEdx421BOf2Pb1DOM91NOacHypgiCDkpGMFj8eyo+7Y6f2gM
8Mx6es2Ok5ERcLGt/wSC+Kn/pX5BJKgmpHiXH9mWyhJZHpSbe5V6gjlHEl2cTNLiZYfeWp/ARBCa
jGuSpnVnNhz+P+LXxp9SaSfZ7ynO21bO4S64GFieyNJ9g/iHjxzIDHlnYm5nTHgt1o2GWKqjOSxg
BUoDzzQJhfYIbV2DkqtmPQkN3KrVsEUavX/en/MVyXwuaATVKvllYQNZ2X4eS64rkhXtmu+A3DZy
7m4UwaJ2KgS2fNbkWfPNtoh4TMU/Q+lqKTTcBSEwfnKmg4EbC0e5J6UrtKirevh4jA36eZbF+WVH
hJVVtpxFnqzJmMn3zw3pIeIqvPEk0yBWmSA4ySXXBA/dl0O3GiABoKPbgBH9cdWGWI/WtLjaqkmx
qxnsRoijopo62JtU4F/WnKhwM35ox2TQwPgMfpLpoWhBzjoL79GCJGJVU/8DlY7nK5M87OJGY+Ot
ADYTLqXgr2Z05toQ5vCPW5G+bKnxvAniApObLrOIAZ1E7v8/3s8c8h6sEkRN905VJsnUaUE1Poos
MZuU8FRh616VhUDoESymoMMKjqL2cYY9odOI9HmPwVYMNk+5f2ZTOYfGtssfMU8d/X7yEO5HITU1
GUyK0qlnam/O3HSMSzdJkQFIqEn4GQvDz489FZ9FuVnxdVp4PEpIRmnWjeK9fmJHnB8e1e0PMbI5
NLgcRwU7o7qTrCVBDNvZWss7ch7/xKhayb3mJVOknXSe2+dshBbeMjhS6TXv3Z1Ws5hWgkBHBP0u
u2HcoPqq6qUhwNbbpA7WMhLg2yZnO5aISfBLWZ+iM66mdS5z3jf4439BNXqYwFtAmHuZuFlRPYep
rRu5ZbEU87lIvmicnHKZyNSWv6kAuVQECmLQ1k79jQqV0/sI0I14cT4854DTrTOjIxDgWaUNQfPv
si84IOuJiNZ32GdFjTqFMXga0PqH1SfmJjk1rQSzvpXz0cl3dqsz3gpdaCHPYR73nygDcpOZW1/t
Zh5mxIy1kwGwxpjxJ8zNLIccXRzXS41BfjeUOnJdDwWM6zOAqrFrlNolnsLETaWBGWVj7eGVPnGc
ILryKYHzj+INj6QtjFcR+1SLIMOgxaLuXCE3DWbgfwOA5Q5djVU3pYCh+R6jSmOTucUucxNCMS/S
VDneuoEyjFHFNRogN9AEnj8ds9m/3+kZEeu40TyYyLJmn9Jjc65ZgY9rk9fUE1m+p1q2O6ubT1UF
We5To4xoo0iMRELAD6ZPdIH8gcsRqeJw92an9dv8Krn0inuglhOwcusninGNEzASjIJ9etgnyJUX
eSyxPf6w+LbsjKYeWDc3MRD7omNgsKlm2WHJXQk95aFRMxOfhfAL5wn9lfQ5D+7kRe07PhYMVqA9
NAmcxXFL5zVFOTo8E+pfqcZwn7aJKzYN3lH6Lu/q7+FY7EOpNYm5k2AgV+t3Qs1+Gt6+euJ+rZKJ
uC2qkJ0W4bZn1ki0Gxn5I5XyGqcRlfiS+J6jX5lgiMyR4r1vI0OuhrcaM831tuDvibBzY16pDKgn
f3moBGaTbm/MMIqVI062mw0DqO5t3JTxTewA7pvXqMSrFdgO/S6BopkES27mrKAVmbzbobCHxzet
10ZZmO7nrO2+fqohQqEszWmyleUHVrFv7JRFeBfCOePZBNbBAyNM5oMA78JEoEaYTMLNUmCyJt+D
751yv1tYptQfh1o8zJl2pp6NALU/3/3A51IyOgE5Ki1Wk+Tp2AxgLFu/ZmmUVRKfWUlxdBLs7kvt
dKzvtqHha+QuLXC4eb8rA5c/RCCUjdJ6DlIX+i0IIg+ZExMYhrTxpq866BCVfZfg/cD18c8j1xY6
Rys3dwCLPtlcKBz55/zdeBardLBb5YW9YwdmZqkl93wQOEBS1M/tdBmpqM8dW8we1vu7bvTFEILF
xfzYcOEOesHofPrxyQbDmQ15sml3VDEwtj3ZwTL3UrjxOM/RXVogtEffz/DLGCEzaH0YBfOue+9f
Lipu8iNJkSJyuXe3LslNOakZyvwKz1kUCTzP7vt+ddvwcWA3GF3coYTece/BL1HwOYlyNx7JwdI3
y5/Qvd0ZXujUH8LwGP5IAYHOnTQffkGmSIJUj94mO+GCrBm99Pv6h6cFEDIy4+aFEYXL0s+/2Y/8
AsMY8Scz5IOJy/ZN7Wc3QP6lB39CcMV0HdEDCd2equu0gNVz9cj+3l5rNxw/bOc+soNRY264auqV
ScW4y0O7vIyhj+gXHwk9N+xPVNAO5Sbvn5vXX+Nnd5uM6p0o92KuhdSkrzsuS2C2jkZzPIM2QxZH
eJBYHm2yOO4T2ABebzxTX7RU/HcJ1kfsxxU2c4mnhVWbilfEDy0M6nNxAhVDw9kWoQQdJNv9e9AZ
O3IEw84amJ0w6vPQUWmUVMiIszvQPV1k3TTRbMZQfvANslpTUCkJxFm/CA44VHfz2PgEBCmf2JQb
3TwYYhXrXgdfCTMyeLI+WtFhqujYsAvcYK3fKgQxMMbGIdBcXUZwdeFbVHFN9izjIzzQ3gz/XpxS
uEq8wIZUt/xgeJWCNU8jQBGeS+e+oE0xDR9xg2Nn5iQeJPGSmHsvU1LO4wQs3F3kvu5bZHXjqj9j
L1HezrrRxHgFUPpvPB2F5oHo2PD43sUvhhSbi4aKSs3eZ5Y9893rT43VvwV8UbccO+5JEIUVT/bb
5CuDF2DHiEg/XXVePNNJ1s3VLZh+YIx5GYjBBlJmaYLrJOgqkbicfb87Uxf9KkZh8EP0P+dI/9O+
d/A8o7zQz7KDzlSAZ5T1lN/bOuTGU7AuG7w/Lsm3zUpMq6qkYwol7gRJKq5oF8VW70mAcViCw1FW
g8ZnlY8zrxYdGbcj1as4R79cRuM7dW1xERMs9mXCP5AcwXn2rHZZ4ZtUb7KY0y7quyJOblKlZJ1Q
LwqMNtljR6VGsSkUiFDqeszWbk+QeU5okwoArs5xRdPvKY7r9REIRgZHk9CAVya5Zk0r7P+TykN0
5fCWkBS7zO1x9IjiLELRtPFfN/j+P7NSRxe3dlNNrY17y8/bkIBWGGX6qHBlXx9tbdLVcvLvB2zt
ZEMzamtjNuUKU3kKp26SOk9JCq3LcWLpiigjGgTmehBnYhbfsppcyxCAg9uzR6X982d9qt2odhpO
tGDAHsaA9vM8CuvsC8SeCKuI2aFxwKIthnWopqR6IrxXpBwS1E/dXoeiS0JjOFUV3kZHM9NMa0ld
udwFso42v2xZl1KcGzT0dk7Vi4FQbWJWDc6gemsNAF/sdBk9jGuN/V0z6PXpxrgHlRPgjCUMRT7i
0S9PLWKuzSaXBsHFX6GT/1dWq6qeOg2dx0518bxL9bFrGGy1IK+GAtF3fzWY0bnFmqa4pY3yBP1X
8uzWUk2/60NEcAC3aLSbrzxSvnykenucD4Ck6dLr9yBZ0jTSG0Zz5azga9Cqpt/VGySqYNMmcjfT
TUamNB8NBzdsYpZd0xMQ7c8VE5IP226Altdtvv/ipD7POkDdRE721QKB++qBwkMIkHSYOSXReqUW
49pE/4qVAxWU5U1X5vpq/viUQOzTRsRwP4rnYJMdrDla3HD8I3DpHhrrI7nK0Eeev/6AT3FQsGyc
gsiHXWuK92KFClAgoARWbkXlvZWhPqDH5TpYeMvp/NFuyTW1Ili7zeRw1xppK/4D1Bg28g/ImxU8
AhjggwdDwuj+5/0m/dqnVUyg8KFgJv2d4CpwU+bcYTmA2TDKmLHS1rx+LUfeVy2Au6H7EBZcC/Ui
GivONb9mGc5PQeaD8tykSbYRQj+T6/jSO3Hg5WtCDfe3ikyzodWxbBMu9mMb/mQ3pp6zBQq+NZiT
DYgoiDRGa8VeZwIpZn6JqhUyD8G0g+q5UIhOuNCJqfq1uT08v7CsHDYOsQVNSgSjS7Yaos/jtD87
1Xmqe1bYloVpM+v5XFqAK98JFqMAliGCJwes5kS39nuJcgbVmp9ZwLkykcAI8njCE7OFceRLxH3O
RzZStZFrdoPEYo9qz07f7K3H3JcA8auBpw8I0Nelx9wD6aISDUY1lqGtWPX9Ah9nmlCLZXngOhll
eaaCPHq+oVD6Sgi6rwav2ZBvwiGX5GQXprIsUrBEv5xVGKHvMew2sqwHw7aCDt4kpFzB+/j6rbY0
PzSrKwoAkmVGVvUHi83pDuFQGCJkZkYwVa3WyTqleyZdk/paEwMGsmQk3hPlTT+5OQ2KvcqgvubI
MEoSaWCSqVKHldi8NX8W5fQFB3lf9uwHzExRkq3ra9ifGu9bFMk/KI/tIZtENq8vt0KWemL9MlQa
eA7tT/DSV41vLS68bo9BkEAF2SwoGBOSNymY5PrNEKprJBKqGldpcBoR/qeJ8BMU5Izf0mg4FqQH
k/TBdn2pOnixN4S7d1i01ee1EZS921chs+R+eDGaLQMUk4u1Tr3ppBTaUAVqfeEaGuQRy7htO8RX
PsrU0PEaQOZTgwOyeudc6qMEe15fotQNCjkJAcMq+uYj0+fAp6MptjPZzD7WhfxO+WFNJN8j9Epg
S24F63NNbZt36cfY1xrUnUN+9vsbExcMv6GzZHPl+Yjnf6JcrREwPhm5PUZb8aXm15btZfpPdrQc
6pKyDLim0D48UcLIYQX4SVKMi+WvU3MnO4ba8dTTLn4DcjU7Y4yw5FmluRX6Hzalw50+i3X9DrI/
pGThzmu39/STKPT+s9RPXEm5lq1uu9fdhi86x5ljsZ4tkCXsgW6+S/B27W6AYtfW9nshCTULAYE6
R7Q1Ug9dGQ7KfRPHKq91ocE2XS8raRPikhfKegDwMMn6uZECPwdIvo+NwzCMlxcYNvOcLE+U/mUb
MG9XslmFrP0ebCyjGma7dPx4m2l9cNBPhAjR+gdw8cOZFxnrV14mwj8SnINqTiw1/i0vqjVDgYdS
GkQCJV1+NKlX2favX88KBXSMP/70qLaG9iIlmCukBs1H+B9V/hBxxNsSXe/GcOw9uWvoVhlJ1x3j
z4JX3lhsU1Org5Yp8AgJa/yTvsTwd+hx70rDto7brWmS45Cl3jlxLIGB+q8icYArPNLxQmyQDh3Q
n00eBmDGF7+GYwz+JTF9XhdqCYExhTl+LgTtWyxNR5P6P6hAVmNgFZ6PgPXzFQnAXFX0w2hdnA+d
Tc74INp5bjG4UndKXvLuSFcgNWpB1zhSsr+YXef//UYsMMetD9haHxLp0i1aDsTvl9kF0MZxis0p
P5del7976meNKIFyOQ36KSpOwI9sXFIemg7jVMsQCcWcrKiKxw6dqHOi93ZGaFgxEq+JD3SqjbiQ
dV3eEBh4Ynih+wz8MZF1GGzgqV4PK8/LdPEJwoNSXbB3MisIX2+LMfFNkqLoxr5Cd0xz7m59SNCE
ddcSU9IPppEV75/E9IGm6HpkBYekQOTx5+jCu57PgG8SnducDw6q3xwI9JgCqZ+uFuAM1fPV0png
c8o+CD2pho6iny0iWLrYAH6dlLlJi/cUeJM7hWPPyc3qhLSdWvj92tqo5aCJ+pZ1hjfeYxrf0jMI
0XsLHS9sbMgaNYvUsg5SVtFR98EJk6BBQWIOWGgiRl2HGmL7txIEL9NwtEcqdiLv2PEd/abTumxD
c8MLIepZ7puhrz+hk+cLfPYkKCNh6yBGhxoUphzTSukIoMivUzFP/IWIy1xhSsgSuW9jRrkU3pxo
7HZYwM6W5aN2MZhLfTJvDNDUORLm5ZFU+AGULblkPIdzAaWda/3wQ85fRnw7h6zX9DrNawad9zm4
1GDnC3AmoONXxgEP8vN4TrLatUX9emQSuQSRquq4v6Xq35+pMaj0V+F91swh4TiZDcBR/7oZZUq6
cFn1+zRITFBNzco52o1IJdkrWoUK2RL2y1LIo+s3KJq5owlucaboeuTAfjVXc5vMpzFxSAcOH2J5
tbVBcO46Z0hhXuAeBUFlfyE7eFPOi0F0zqNuJ80t/mgjKMgAj3jCIWVxDPWtL7QPfArsesZpEplq
0jYA6XrsQBmG1Sr0xgPC9J67pjms+7/Jb5b5pEQvZWgewxrJy8bgEFHwgp9vYKI9NUojUy3wfMj9
MqQgFlnRIyurmaeSc3qqnuGP3UCAAwjjgczdxlfGrvIhttBKXJeyci/NBg6aT89kP1DL4Yuw2Vs7
uTbTM1PQIFXc7RuwVLamjGQDIs5TXrPM7mnGD+p21g0Cub4U0SZ9BYY23AEVjkWky70PN/RrWF6s
MDWUCWSwc22t4s5MXbZ6D7vwsLFG5vYmmUXJZA/5UQbdcfD+ja6yqgeXBRK+yjJ3wMKno2QXZNRJ
PJ34JYz4YO+c5SQl9IdAfJau8EoDfODuk/R4i2L1YOTkq+nU20Xc/x+GUnHIArepLQwmrUuSsSST
LgYmc0aOx/+4h3R+PM7v+ONbkbaaxke04ogiltm8oTt9/31yNNGZMRz6VotnEf8PM6qtPo4WG6BD
nNpHzzRLSlYAwVdBCIqCUv6wdz4n7vXSBYd1O7RN6TG67K9cogcKAVsIWV/WkduSadX6Zr8nOdTZ
BWSUr42iibZGph33ZamskPte0V3JFEhihwI9G81MH8xL9vlVxe+0jwLBnnXbS0qPFX8ocVFSDpmf
5JA4ZxJKhRal72ulni1SHPMWPedwx0a1Uf7bhTn6iSV16vf6a7Obmy1cUMhC/ngcGo/L70LpB9y8
H4ijWSBo8kzRHk9HIntgulejaG6HGlS+zQfUoih5jH9VFBiqxanp6ADRZ4mKjBUTqjd1hV5w7TXY
Hnsu+Ydx6jEC3lAvedhuWYr3C55y/u/ouNfkrwsqtRxajC+dbVRIsnTXNmViJDgVL5pxVwWdQZyH
GeUcCVgWnVyppuGMUurtHPm60ew3TKkS7xsImP0CqNSSLINvGPKCXuQgZK+ehOeBTTeDmCdmBz/a
TCcRCGcITZkGWllTE8/6yw9Un0+dD0B6r++amtaGxqtNWaotGdKGQA1SbRIMnjqOFEGIjXAKDVb1
oyBJ5JfYaNz4ey+OjvlE5DUrupS4GTfqlX60vs0kylFSvjlJCAOd6+Dxv980rJaI21V7jUo3Iv3r
w9zjPvS9WgVCiNhKW0/ZmU52/GxtSapKExI3Lcpr0/CvhY+Dua90kq1wN6nu8RV4qHbqndKnDbcN
Qiv51rg2Dh5pprH/Pa0/jV+C/fOEOWb60ly69LoPqmseOfZY0mlFKumae6SnA2cVaO1/HrYvKNAW
o1RYJOYkuyrSL2wzESHwWS518He4QoD4gASdBVoRLD7BhptGRqZplZPdPH53ksaBamcCJ0QIufJz
c7O232lOYNGI0oJM/sGt3mSLidRiZzvxBk5I4datVH7ml9tLrUeug7TxeyV8GWu6ctCGzE8aFlYQ
6uixa9fo6w9LtduKpse0hZ2Vausb7r9rQAWdxJePy+mdCsX5Npu3JS1bD2RJvuHcPb/m5T6uR5nB
MbJhapgMuYWyQaRXWXrR5c6HSBJv9tyBg7+xQNPWiNLyAbNVlaYHMVgy90zzzefJddwi5Fp/L+iA
NJUcd1thX7qIV0QUzgcCH6MoeLL7JIlFyT/LT8gQIByQmuDrbmgQs3okDspdR1DtPvgFa3Vr9iNQ
PVai26oBWiD3W4rQJSL0I4Rhlh4IYi2zTxT7odqJAVFHczKLB0xhksc5lFeIIKIHgtwtc5vXQj8T
fp4Axs2GUb9UHUEc9npa9nxuAhXTTLgSxq8IYZRhDJIlYX3VnLJ6w7qQdBtp0cvgh03FevhS33Rj
L0hftDLDPKOEn9azAHEWSkqZxdj1ataHCK6P4sWPVqfC36s7Mn6fGRgOrjtcrkq6SBQprTeFT0Zx
rdV3UCnfNhSHFvVdCvyLunSTF/TyPUuNM6ee9LRN3atfyvD9hNAmNplIK0m/DPISitoXx5CIp+rv
lYvtV5YZKiZJuM4U3q7LFtU83huYYMuH1x/AOLOVcSY3EEUr3L7SdkxaBn+ccHX2HVc9TFGZwa3N
QMku3p4x1Hg/F9qFPFwcEzu28Is4dIFXnrQfz/t4/cnVpuUAc0eade8AwImZgrVfpqobbhMA7H1p
H+YpwT6Kt+FNSGIBffSqajPyd1TlpOsIU4leL0fD3tq4RVm6g3EMpzU0JzFzNFS+5A+yTAVVVDOv
YLuqkciKokzq2PQBEbmCOOv9VTqgsLwHIyihv7IQEhqOcwKWZfaEiygK3i6opmVnZlgxU/nKdZkg
32YWqNJ0BSTOcKq5HVlQC3tTvZkLydJSHWvhFeb47+RFyjmqZQTsc6WeK8MdEQazFnI3EmZngGw8
WQF6JvLNhWsXtv6+uoiQ/p25Qw1W+5VBge/rqxZT/m55zktlOf0H79ONzHoF5dX09fxvxaW68qA6
HTCoS3t1lO3mywPKgOj+4oUa0PI94G2Id30m0RNgs+dMl1RTLKY34QjRrDv0i1Um61P9zgoeP7Sx
lfzpFB9rbqKsh+up91y6YZPW9KEe4wcTmG9gUm3Ctu7yB5Refo8phK674jKI4ZAmnuXKLl5FCO7r
8NpIWCSgMLtpXAuBynjdBGn+Yi2EIfdrolwAKtSa3RdaAkLTI7oKIgEJgSp2/UnxSdAxaEOJKuu9
wSey6wxyTWEcMxNJukelseLkAX2JJp7IchyJN6J8wQGabsOV0DXBIes0McqH6B4kEY6TwOGBK9AQ
jPMv2cnliIgMtasxKsYKANsdaFTOfFnUlKVfNyulxYwRjVAsGJLHfJgdQtddvcWvxOg9tc0Y8mNN
SqoPAgZcQz7dixzzYoS8B+aXAz+Kgs6wRzJ1oxon/w1j1tspY+3jb5S33gees3maqox2PDZ1H/ww
wZ/4fOvrg4O4yEQOJFEyUnZPXqw5NxSKfMQLSI6J8YMAeDkN32HsVUOmzCSXr9LnUrcx5rJ73/0z
MHervTW1KgjB8p4qdp8xR++6SvzhgEL+2yVg1sL+99adE7RuU7RVEm/A8z61Zccc8ZK2Wl4sZwmd
sm4HVCM5t6xr48zed+QLLYRZQtnHIQGjiNtnFctXH9vcMUP4NWVJw6lyvVELJeShrnF+vaqxJVyV
MFZJCOljwH9qztiWyDGgmtSo+DyabP05rEEbCaVCbriKMWezB5dsGG3AkSdcTDp99hxF9CGbZWOf
OYDNJM67JwREzFURsc9q8YWnJHQKt04mjwr93+WuQbnVI99ER2TR0v9iky5dMYwcOQmiqcwT5XfN
YoDu5rhL9BRK3SeGfcOwNX+vncPaCosQAgm/FmWGMwAxwPDMk7inspkKBp1BExFotupgHs4XH5Gq
aQHdt5F2LjT9Yie6TbZpLbWyKm22/BlRf0+PozXb4X3m3nuxhnN8zPjDUwwHX873ipgGQSplGyIP
TU2Ry5vQnqLSSliQU7Mg6t8Pc7+GYTNIVG/o8J1rq4qt6tOTml3DQVNFJW61J0qwokx9yU96pUwL
YdPlWy5eNe9Nm9flPGLQhrhDmtDb5KPD8t3wc+1q6nSxfX1i9vZBJtPyqU/iKxkgPxlgau4KfuTp
chS6rX/n2n7ThY3oGBWlhwB4gg9J132BAB6Oog8PKUsHaxhPS8E7izuAAztyMv9kEeGTgoHpgDxk
Cw34f2owGDH2kmJbnmTIQxXWkH/jlMbShkm2Xk5vvJpTwaMdqb8y5wd2vgpkmdh7DKeVxCH1QPtJ
iYIurm0TZYm+ALkv1I7tENCkdjODzPBOlr6ecREKsz490epWJnXUk5VWn3X+8t8DoLcIb3a20M5O
JjZok6GSA5Xj3HZnaDlzOWpWudJMg6h3q7OfmSkE7hNJfLIyjzGNOJEwHMMVbXpxMp0qCutwwgIz
i2pz37qrTV7zTapw1rlGmcj7llPOYlQhkuTlmxDJOg8YKar6BujnDbrXjQBoZCx/IqSysKXhqht6
DBsjyk49p6UJw/rGGh550rxcudD+3fiSM45TIgQSUydGkphIaG7i/mhSiv82/UperVhoqva5USyv
5+2M+GwnS6xHMjkSDpY90gCQhrPVaE0He26X7a+FZDSBrHbZkZqeN2OyKMkuW5abfq3ZdV8tDWAV
wCZ5iC8hwYJfP3u7bjJK7M94Xnkz5ajMc/NBkr2MXbpCPa/Q9eJ3Lof34NpR0DrlewWduJSAUs7E
hW/D2HqFxID7SYufyVd8K8h9UB57dTJuKweUc0W+HZqZ42/A54qAh6TjqcYQpQ+eFuBf96JpUM4J
LYkLi0P96E8XTKSOaa56us0F7zawYnytADjHzhf/8mprFmGzF/sIxnyYaDavgNuXZmDGSpmS2R+G
VcWvRAqovrN+FWVc5a3uPNENVf+Gd7z/MmpJwXVRlXKtAj/EmmrnUjZc7zF2753dMoiszexDCMI0
CEo1Ceqj459fS4TfzDI4vawlwMiB+dJTfv16c9YxTtN5JX/QxL1QNB/W8ArDRn3bw4CpFzRaNCPY
egUpBl2v8xFNi1fkDxTqbAHNKv4q1UJy6GldhCxc+eSluLYtWGmr9gDxSu1001x2G1aczf5BwWRd
t57231k+b24H3Haf/zQdlIbz3yeZjr5AvDr0OAcb7WGcicDNKymWhWLVbu+AtM8gubl/EOTQ9Ek/
EaQUk+qrK4JO5g/FQoma7H3eNLXO7WKNOngLCNBwPlFov4G4DpvK6huCf7paGe93ER7QEzprj207
3Ab0GmNrZkPNfCZBz+1V0e/BEECRojmSdKoT5Xr/kRtyQ7Fl1xqDKVSKQmjg9hoUVVq6j2p1NUPG
KMoNcDn/oejX3Okel52hypwt1udiMEilGAO8SdALYatLNT9gxzDZGQ9YZzRaUilZcMSE1Yb71ncz
HlP1imFDYhgrgl0xxkfZcpcO1yyUyigV/PRT5jiLFvMbecPhEPgaPF3HmMf9YzPwZiTkPs1zkdt3
gmPc0g2j6rAcp0+/2oz2H+a5JB9ctT7A8MCGOdsO9l9sl9xXaOTzFtqXsVmrt6JPON70EDBVRmLf
kYBlbvV6y9Zth34Tlq8Qg8exXAkZq0V9z8UzOgHPL7br1OhB1IztnD4mwHOi0yE7TYWkKIpbvn1A
fqb/ChDKx7VUIqjd0DN32B25OfT+FWbjxuw94TV0SWKCmQd3CfV7kXqno86RYnGgpx6+AbneQmQ1
b244Bz9XPtmzKpYMPDwsUTkqkAgBFBbC+JGrYh3EjfavszrCxqRmYBdXloztlw9T6QpqbCmFJM36
Tn8guhT2W7bNIc1eZHFaueC+7RBCNU+vXHGWUU9Dh64eVuvJU0d2OtcMs8UUZYSvCdrPKcv3n1O+
lAhhCe9znaOT4axVnE8NtuK1r/kAOpk5whAYAygLGXk0wW2e5I+49RM0JKVwgYMZ3wc0UTfqkgES
6kCxVQwst41KfG/eZut12Klr0FNNugdRAkLFXxN8s1dNzce9i7ntDJz+k/NMfqpKd6qncuIlBRS+
xVYCboPf5heDVozdQJ/IdrI1/F+eHX6cwmlMzOXuHTLnV8LZDnGlVwYSasP9ZmiWAHTuWtGBAErk
sGJNb5jKoz4c8/hCy6PxTENWmao6s0Tw3CmZoF12z92ttb2SqUN0M/k8Fu0Z4UY2m/WawuAucUsA
E17caYPxP0zZs1r3tKRN+o2UjYCOmxIi5heh3FkKSHKAzJuD7wP8gkS8eBmnog4ylDGN3rJ6nXLf
D3a7XEFKyizl6RVAiUCZobxpe8y1aHEvG8ciNfTKlJO/0ufzejmR6kaXNdqI1fK40hT0cAtN3pS8
Xv9OsCmbLud2y6jso5D7LCyYQbaVvOlVJF3YiqcOPighPbLBJOdrLnkqEjK9+QEPeYRhVmRPEDQy
gsk82QzMazYbvOREfCmjjmTiLv3i4lvQ/ssVDOkAefJ8R1iAXcQ/WaHyol20yZy3dAS91Qe9K54N
H+bOjhtJ/EelgLF4+ZoX8cXOtBAttgcfaIJjWAnUaq0WdvpZYZbAzwHt3M7jq0JpgdamDyTq3K1E
UWfgbTNfLGPQI9brIb8xR2GiV7a+39MEtsWrCNT/NcvrnXC7dXDXx1non1pUnyMOPCCoDA136ZS5
uVMBra0YCv6H6QOnPIHEnmN50TkS5ZN/hFRTqXgeBsDV0vgxsc2Xl2cLogDNbO8l3mzY8n2ru3j6
Uo6Frdo/sAh4V8QWoa3zhk+wqV6B5Ws/WRt/IsNNe2qCPLaoK9pLFqU0Pinrfdr6Hi6iNDds+20W
v43EyEzmK8jCF+fX0xOTUgair8ONOwjnk2awxCvxTYDhJK/jQ1oXkbOGB1pXdshnZ1xm5UerWPuJ
bN3AKDfipp6tUGwTnXZR1TDeAiksKVQWesG6Nacp5Q7/cGzCkgwzRxfNSGR6GwkK0zquyCOMYRCf
BnBxVXJ3pnQIl6NJaGKBGJUlfrRUrWfYgOvoPMjlYRhOfDWtXTC2NLQzq9nz9ixHgjsT7OYpRER4
mam4W5se9mqLJJNdsCfcHLo2S/9C5DWhpLjkHoQHqMbnSU8zyBCVBuiUQtdz+obc5kvj6AmUh6pu
76ldy6RNsgdxsKbA6UM90kEUgW8cPjn67Z6sQYz/xeedRe1xmMoN9VGf9dvK980Xe+FojMeYkWzZ
zVzeT6u+Ol7Ln9Np76JzN79evTaYiMZJ2R6m47DXRqBy/Qp9wcW6AIjB8YZF9Vlns2nC10xhToKT
W6Fj8eXnKVaIeK1JOWB2jLVFbXpej/EzsEpCXSjxSW1ftFqbuBCqz7ajJmRaJgEnkog+oImGxsrI
QjER9C2oel24jfqx2LZfAEEYxBeRWVX/RaXal6EdJXk+egwhTVWqCTR2ERvwwPriGP6+mjrLuRZ0
01goeRpNBLFOoNKOhSVe+zY1IPVAgTuW/mi49x+kiXZtlKAn6P2lO+auyBWngEFYW9rLASn2/iiD
DvaUKAjuM6LRaOTHaYJjHoEua/3f2pr9v8vG6JI1jUxDLeHYZ1bj9OGtzn1o+FZAys87+ms6+Pa9
yV8Oeq8y4PfIyE90Mi/0dPcz2DdHcU/Z3E9A7aSXLNxQ3KwGLpWc6ERvs/47oMhbhg5CuGraXnj5
d2Vq/r5WHEY3fJtXx0Iw0yM4WmU2Qj5KOj/2K6AWkMsbNrho7TxwrVG5wTMJp4M4NEZ8qhj1MTvr
9WWNt4ZjFOaFJeJ83AnFVoa95ROtvI/hl+Oc434IBr4/VnNDOrdTqAhb+SNfzRz/kiG+MydS99wA
7sdQppXOFrkrUxNJlk14rIWNtA5MXEARR9gQ9B1MPcc6lUIQkpogdeWkZPqiz8sQcsWs08jSPqba
Ty9U+jQYCB3PyTFvA3FCb9VI+Is/IhACThWpkipztjQnll3fG8jw/syGmtVPNzzaEfVDRy5AlhzZ
XRMexM1b59J9+emwB6bs1vMNjbStt/mB2/3bLuFRKJP+5u/j3WMN7/Ld7EJIOtoeB6Fs6B/G9lCu
NLfifqit5CvoR9pn0Of3i9u2GXpgUceCBTwh2IT223t5fwZEQFJjjwLPluiA0XX5VeP0jVIUFTyU
iOjeAGG/IKK2zFZVecHhy30WI9LDIsL6V/8DMZrpBtNxeXSHe4R+90xgNUREC3riW7LzKDN87sZU
Z9wl44Zm4T2WCp7UYR6e/6PmHKKbc9gvUsYYmv12shtY8Wog0IFuXAqMfnVBKePQhklH3fr/525M
2f3v+YOJphQEqIUwG749jhXfcItsofvwkexjtD/TP9Ijhj8iflosWVIZlj7XZvVqwlUl+MmulBZt
3/BBFtORDwoPPzNex5Uy5qrvE6GiJBLNHpvk7IS+lybQV4D687az0ZaW4ZeBC5EjZB5E3cM1aMXg
P+su0wsPo2iJkK7VmuF89Hn+AFqnJVK7d/mmVtya9IRTmrQ/xJswkXhwxOSrg5OS6pnlrqimx2KH
DGgnw15MiMB6feJce/dbisCeXZDjN7F1Ex/MzwPF5d2CvxTVZtuyoSGlpzv8LBOiWvadwrq+aKzf
e1xwGnE1lmiTgyd6ODIw4a5D2mdZivPwr4h02DPH8VGMWhZwVhiZmQdYSEBgyUkHJ1fiKS6G0WMY
pS/VYHRC1hI+ShPcEnJ+Q5ZZ6PByAtyrRv9KgS2m2t2mvAwbvJNP88AJD5gYh2aFUpRMC6MQXrt9
wO/kKLXNG1k8vjWa1jZD5FZy2kQfHxY48FsMg/p0fYvpH8pbzbSpq8JJooEeNU9R4hWdDrJ246qV
av/yeoJsWRthpphSDW9xqwRofVATvMBegWJ1fyxhqZfozDcVV10YzVWNCnXBiwVaBbl0MstK8/W4
TQx1R2vFoAGioVWy5hTLmW/VgxLEKI6zGlSmNkAY/m3Da4yPA784e5qGzPh/+Ug2VvqGHFLVxpau
7vlU5lFHnhDR08yEEzpnA3MW+ioBJz3GEAWFQA0XQk8fNnitAudbt8wilQJ24rOi9Zrh8+J+A9Ju
09YJiNsTFnqqMGsHN9Ov2ferGL6D7s9NasC2b28dqrFe2HkJnWW8C1I1H2qI6jSAxU+bhAftDGYX
lv01tu4Q30Yi3JyZj4jsHYBsIMg/6BIZ1nbVySi6wv4N/tW89KL67xIfDJfui1vgM8fXc1wphVM4
/f4ljrlM6NwsEk1lYyH1JspUMENVG5z+8csHrTp+S6bj6vzinM2BGQs1myCR3cnGoEoug9k7uDIq
tZs9Gt65WVaJYY/Nevumvpo58XV4E1XATOrgA4VulikDkb+TrNNRoMfh10vI2rOiceKA0U7oxUkZ
iiZI3x5ALBuJW3bwYb8SEwZPIDsU/fiELAKde0dED0MAcPdPH/UfJmcoRMcpjNR130MZram6vniM
wG28PbB1e1wcDSLd3Oz1sWJDXZdn5M8MGd1jNeIPXcocEd16p4BkLtoa7oJgfj/4YmUCB8hHHP6h
1xD6WdATifQGysTsIBmoxS5Be1QqkFc04EwKP8Ki3lFhXkOjX0Uiufc4iUN1M58NIhmkiLxj0naF
mubVDbVepKECgdQzDiBXuHg2SdMDnsP71b5ZTTY31PoOUCnOFl7kf8iMZ6eR/LFTlnBSOEUimDVs
TdEHhiBhYZwRP0DeDs+q7KQNN6Q8F2fvvP5bIHj7A9lXSYdn7hOIfptjcDzvinZJbo+2K36jqfnT
+Q+z0UuuI2An/eoA1cjXJVi/2t2YpX/O0yRYivLYGQsN8byauaxA6LxdhqAxZqNIwKBUV9NBss3t
xleoxMdNc/OD8S2VC3vekWbZLR6kSIoZ9EFKX5U2tlvQXiF9DTWw+yyucNgBJpkiVesarnVT3KPG
fFFCUtnHhH1J89vMhjIX5gNLs7xDPiPRkiwrX8K4CqIdmxcDxTmYLZxt8MBAf2W7TycnuvfkiLNd
lRsvzIkYJQW3xXCgg10REpU0PPXYQcB3BDx7LJKKRpTDdJX/vKN1Xh+i/MkwxKyKXTZmW3PPOROj
0ArXLfQYOqYSrRZbWMnyu7cjcN7YTAjP/090BFvjMrG9o8PCNUlbLoX30EJJvKgPVOAHIhfGcFUC
un8R0hEI5ovXRhX9va7lWJKoQnJNX/Ujl+ey8FRMcaskDk8ivoBG/rdDp6jJOGQ/DC8amliiFKaB
SQ6KAqP+2JIHfsf69oiW7pQt+GgCsuEiVaNa9cozr/tPRSCgfsgOy54M7ghxXtv1x2QxqP3E/5o0
UjpELjiCKPnk7GJQrkQ14B+9IjiK5gdR5WFSuNvRbHd6Mu8KQx17GlLtZ7xjmi9Lrl1BqfGy57QE
JXEN8p4+RS2ZwUbRP+3voWCQcrCGcL3jZE/L29UHEVhYmu50q9qNTtIs+X0rrnWxAo1hRiQeN7qx
dDCYWsLsnqFUia1NODRWlxB+6RquwLghqB1bsMgrchmPm3lakGkiTQD2Rocuo0B3hLhPOIeR/8Db
he7fHaVNupOd1oNtYWZJRs4V+Ta9fGltb8lv6Wnt321iXV6Ndy15yrG3m0XilkkK5z6+x+t0hrv2
OeYKSNCaSvFmp/Pcrfus3bmHE+RoDcMZq5s/181EeMdj9AYBaJxbWeOyEuoIwYmz4FlmLgpLbvAS
yzrtwJvyb+VepE1CFdaU+oojqlTRky9OgURBIb7E6CjAqthMattbuv+rX6WnCsdcxbMC2nSDDi83
IaE2xwk7TwWORdH7KQvwV2OvY3kXdUzHTKdETMdOslP9Ro6jAjJ5bT5eJmSaikNdY3Dw1PdTaBlP
olRtK8+oCurVavPP9Tv5lz/KE+5YFxapEYFEmZOU10bfiG4qzw+cujTwpIuTo1ZEQYtgruojgLlU
lGNB1x0+sotIUVPFghlsTk4o0cHpiECLVu0upDdbdGiTrhAaAgscluXljE0rLyvjPbVfCdQG3W28
QiFeul3dPOOi/e6YiUu9bldhlRIxsT3rRYDOS8NuGjREwZ7xWo3qpNP0SwSStVlKjxs4m9Ap/TdW
7cBRza9n4+ZDahwDoMgoIeHFQtyiJsnq61NhKcoLEnEz64RftVlDLlKT2zwfFiM+UeJioEEHyThk
P7rT4TXjQKswepiS4txomya2011xKhGDv4Wwwp95csheiKPzpnpD0PK4V6b+y6L2IWD8HrbtKthx
n+vbALvu3I2LUtpY8eTk/K7E1g2Zy9PsPYg14VLNTLisvdahqdbGu+dEhn4e8Qt+jFeAvjyTneNc
bXxB/D8vgvAkFWRmidC4f5e2Blsr9yC/9nwr5n9Hi7/DRypsFoHnk6qYip2z9hkTls0W4JznApyl
XI0ulIdmKg3uBer1HaJWD1ogF2yR0pHAUG+yn5Gr4uioz5XBliZfTCclIb9Tn1Tb0Ecc7qE48pOh
F4dRfwCZmbIHZw5XcGyQVFMGg1R+EyUsEvlb/L9ti1pTyRffoJNn9HN5MSgfT7efkf6zaEBdCYFI
tQw2Ks1fGIlcBTd9SLTx+bJlBW7FdvIqpneaFEJiFHr91PlfDgvqgiFG2/3drIR2rDwAZKJ1d0Dh
F1saUD4E/DRb6sfa58fIdReOIuYsf37rcZa3h5iXj56TE5azYIGkA+U7NalvmlcDn/+jYi1g9zw0
h8iX5JUufR3I15wKxIuSsregRL9IPo2NrR4DUgQFWB+yYxSSQGxd0dDXwNcHlebqPLNMmJVWePD5
aPZkzyyaVjBwv/mvUr8wByo4v6uayCgwRpKRIkfl/U18tTdeSc3A52Ti5gWtcPlaZGDx/FocqZMu
SHiPhqKRN8aPu8ljePRwLm3RHXMZ3tW3nZkbAG63sIMLwBa6CUYkxrjf6w0Z7gdFJ7PwSwAE4k7u
JrMMDdW2rNuxBS4biyVFASK7Y3yJJpSoWpGRIQlRuIztPBKma8iBW9yRiBHkYrYULGceHgQZ8lxQ
S6IUlCqeki28zA+YEzYUzbFjaHE7rHKqGu3+aO7eMYChxjkbxAip6k/gBEUVCmCjViATvTk9KdYO
+Bj6OZv+L/WxAwBfFFUEsG2XlxVtc956/a8PZbwqukUArf0v4xrw0nMVYyNwKVrwjrdczoRca43Q
XWFB7k2htIeBE/Naqhv6/ejB9sjTbq6FciwR086oN270hLUryxIpeuOgEcOmNRM8V6e77GbklA/K
RjS87mCCe6Xetx57TRC0aZS2WNDpYu29gm/cBV5upLSocKrf7x8K8LdT1IGvut1AO4GK2sMmI4vS
hRAV4NiibWFUkVHyb8Kr7bv7e6oFoi0vhDR6krRg/ZPEJMUoaKLuILY86K/xj9/RNPuT4OlkqDzu
if3J/ujM51D7kkXqK3z4KaIS8VvnMbZ8lyaDqlfP/o82KqZUWEP4iiSSyd9A/u9MViQkCJRsC/Ff
hqb6kAoAWsZIhGhFG+ODSQQ3lVYrGApKlvxY9Qxp2q4wAX2YFJPAByISMqqL9Vb1LEWhf/lnLyBb
TPhCw1/KZVj/B2RWcOXZ+C9U8LFKBNZKu6xGmRjn0mPZVAWKszK7duj64H5E2wfmPyeYIHWhnxba
HWxc11En2ljmLG9kpyDseoaMG0cy3m/ZncDzYa6OFkKeyFk1GTtf4g5y7hg1qi1R4kEEhT74XPCh
ZTOcSInrjWE+X8w9xjKJAz64birwKiFr91bLJloJ3/0uii6dLbMBts/fLic11A508l1cPsomM8Gl
WJE+gi80ZeHMAY86MTqmWX4bVTclIIX+J8dXF3+9bMJJSFP3Q3w5K3Pgp+WGplpyvsx4GmpjBH/g
4cX4LKYUaikDGgjOh8hBLvx9VdugJUyK+tRW9wnv9qX5cIS/VYpd4kEUcqbgYd9rBx7aROO3T1fL
TQVCgv48tdRKEgjnUWI6yzX5lNlDKDFsnR9a04z1e7I4JBIHWGeKD5V74U+4MvCAD8UxrfbtfdlO
bsMpndTkflNMYgGSTNoZLAhNqymC1ZmSuFZnqhw0cWQ9OCSO/T0L8nT9Pkjva+zkY73tr/nI6A9s
XVM4ZwG/S3gKp9z+DrNrp9eKY5BsHt5dStE/Ly7m9QfMCdR/7grHhHL/UXoVgtxdMOksWaTIGVpv
i4ESVp9iyBl2Mg3CLjeYhKq6W/fJki0aC4DBG2pT1Jy5stvHZ0IhGca5p2X7b5grcqJffEGZtAGL
VdLHWgqznLY5wRy1WPLnNysG62QASZTlMvi3BWvR9pQQGBqsnKFgHPFba2XCQbSFC+LvjAUAruOB
W5qlwMzCk6JUrGDOx4NG6ehXz/dgQBc/Um5iDGPCsBHGCf51PY9gn0dvE0oAJsiqkoi9i3DOfhmD
bqCUVBT0IFTScWyQToOhaGXA4QCtYBucoZTJ7+NsBsDDLY+Qpji1nOP8V2XwIT3EDYUb/jxP24at
nv3jqNut2ZZQaMF1lEOXvadRpmX3lfd4H59xVe+4KO9LpkuzBrA0IGd+g0CtAeCVY+GUnVpZ0IJ8
QnKvFPHCLwMfd7ODnyg0SdKBuOS3WtjapnQGLKpCVh1oQGz6AP9451qH5xzn6W843/axxjDoEdal
Eq2NWSzCVp4FaEuqMQAVwEf60/0ufZxvJCyorESiYySrFygMddCUjmYWfIF9Ak4do2NecFZX5f5c
rstZzRcgmpqSDrG1khMUv1QYhYqWT5YU99B/MpMl7XrxuCI0YZr0x6biweS8LzMJBmlPRyTiyOdf
ronwGdDD9V1PgGJ527z98re+fOQA3DJRQO7zqemujYMCmcepyx7Ji7Wky6qU2W1mMS1qPt4YtcGF
IkcnyxJDdpeuE0+10wPB3ur04iy2oFcfyyJKnbmymw1/rU3N5czrzI8wWcZNElxMN5rsPbqY9SZs
SndkVqDWsFrjOTWP5N17zen5jmKdEijfMAJX/RiYd4/ExyTIb7NHSM9lujHYzrqeFs9mwYKzIpfH
sUiRZb96kNxjxB7aBO7RiaktqknyespFiKBqbUG91VtJCGY63LaviY7GFli/iGC8nbu9yje7VrQ3
fXpPvzDX1OMfqsbwW5F3YMevw12P9v4f6BqBW93iDxXNlUPBoCn5G7rii4Vi9ZjCcfKx9Tucnk6N
+faJNzChpqsZRVaTYF/1FBQMJNTay1Co+pDF30870qJJoMjVVIbBgV3fBV65pgi37yjQGKy2nLB1
S8gsNy1fptlamBm9t0wOiTX5MHbLzzzCFf8mddR0zA/eaM+6t8cR2HkYdCpP4IxMBUzxHwpOXOW6
Bnm3USdbXPTA+AsbVk5UwQu7zLUZNpILrC4rnHqUeiuwkTYt5g7Ev8S4T2Ty4skyi4swtmW/Pk2V
vNkFTUiiO/ALDEC1IcqycDBXfNtu/KQtM4MLGlE002nULlghXbxLuuoqpW+XXwdBN87ggjkM55B7
lV70jdtFiD1Jth7DtL9JZCJXJVOmm8oFudOHtWdr0AtyYJQACgm/mHVcpsVFpcDvPm94psynW7iU
Rlce+2D9NmQPKkpIcsEas8cTx1cO3VCK2AHC/WUFoFAGF+Vna3xr8Ty1fh8dERL8mYlKU6+havPO
Mt/GTOyZ/R6Lxnz/DEZuyQG+/gQi6rxZWFl1RphwppFxJadPVl5MSENCen/TOk77hujZ4Q5xH9Px
5Cwz03s4H9GWhRopdm6zr4Xp9MmSOe2uro9k8X5+7PBhxFYGXtLa8wYAmMF6Dg/r4hT3iDkJ3V0B
9TYZwXi3LZT4nZcMwkfC9rCPdtjGH+7sQImf9h409+Zd4zY9j+UTWiTiS3oedv0i523G/FOs/6dV
aY7tO01z9kr395wV3fPopT06opP2iSo7Ejg//4wb7MDXWcAeSvPf9ivF1lNLD5V6OMTfp95IWuXn
xdssLzVYkAmr+d4nyegx2KtwTLiZhlxWgFgUGt5Toa5oiObjxDBzu+0oUN3DGDAkBjMW8gDfCoLd
WV7IiMyPNaVonPeRmdFepo+/nIc/tWa12vTKJ/976ulAnlKt1GBOkUTSSCYBOj4NcoADOqw3FCqW
it18Ow/PcnVvpmemYkPHkc5lOdK6eylX3u0nfHLXXgzyRJqH7AjeOjhPSv4N0XkySU3GvbGuPcm8
ZQiqdSfNG0cVVAmWCRM5MQGLP+ggNsBP0yWT8idGUVdsFw+V4sd2ZIOClj7Yll25OtmBvuOFbOUR
duHwHjuK5NPU6JDm1lRC9VrdFSSfZBpAC/ACu2WWzUebZfF1zV7lob8hDAM3UdaMF5KjN0EKf74o
6tWtkVzkpeaUiiBUWuz9wX0Z6PRuNnqONordwMT195xuiwV0PNBqSYdcNZLeFXLFDA1YDy2sdJ6H
M/qd/VHQEqQrAIe1axGF2ok017tM29YNine/6tltEc9mIzeo8OoR+qnt5jTdky+YFs7UVDvJyNU8
Feo+Yaf9Hst/65OfvUVIub4hpygP1OMgiaA1Xufrh4QKfToabuDcrJLCcBqyEMlJIu/ze0UNcWXi
e8PsJjjKx1bGB5cmKGI5pKIQuHFSrd/L0Cm8pCyyRY6L67JYcVcoio7PLQXst5JPjggEx5NTyi1b
a8fzJqduJkNj3UWJvi0gcktMnEijX67VOOJ69k6zjZbNYLoph/2laUSDKaHGDRjmBpu5GoI/2mBF
u4Xp8LT4WVJbH2CD1Vu3wj53KH4dkHLHux/W/GUDhykuS+v/TIPHsT0yO81m+DlnSrSguMAmh7VA
rKGpTIJSmwI/uCqS4ZO4LRWPpuAmg4UvjfvEpPCebts/lndGDH95Rfgf0zRPL/hGQk3ai/IiuwpD
vKHYUrQMnEyNv6e6EolE3MdQFnxbzrrLEAmORCJDcGt8JIFpLkaa42LMAOdeCoK13xEEHAtdpdkZ
xkbyemHWjbbQ4+1jmYrMHmc0NwLD8bBnA0uDivR7cfXB6lG7nukMVrYu9QSLRJPZlx9g0EBaENMQ
zwKFCFrWFvE67hjEPO1tHIt2sGbt1v2fdu7R2l9q/a6LQWlYQB2lUOp+lj1FhGpY7L0XRq4RL4hZ
qAxXp9ZEmP47tVxFY60QbUyKvyyzoA7A5aNFj8/kfD9qTnv7DcVwu/t0qXBZNZ9YnO/Ft5nOGhWD
RcTfZEnoYh3gYgHXqBEfwDc8kdW0ErUuU3Li97todP+OmKy/d+ycvDyHEbx996+xb6eJ3RZKBf/m
94IHsjraRiXK6nTKwudSVBSB6PEELnMYSzYzKeT04IEVQoRxAKZMbEVdM7xOZatTBDmJ7S2d4764
79pkchausBp9QbP1+SuOYy8rmVNrEc3Dv61Txq4nOj1jbtt3BUpGPB4kj7G50jjQoFWo5pZH8RNM
AK14h0THFFjUAfTFAqsyzDGLqfc9rJYoqYLhXOHFuz4GVu7qdEo53XEXxM/DMYIZMk9g5dtB0ix0
yGnOmxcxENS2/Vm0g4WBFlLnMzDAWsBxGwA/d2jx7llk4NpOqUhAsEpD3ETjrNbwSkUxUPziWpEI
0Ie4ae8zGIgoJBtOfltfm4JFwxb0CFVDGz7lnsQPylBdXicseGvYcye6/VJdQhESt8sHOXeRnK+V
6TgvhNI3+KaUM3m3vtur/Rj20MWluZG5mDRxW/4vDWD7d9CvD1d4jCyx3zBYkRnhaU9taEYfdn37
KAR1xMUgiLGRS+dPEo7TiVqgj244fDhpNNaNZJMKapno30cB0XoW59aGz33BbniMfihhpP0Xa6Rm
MzJVV93hhL6rDbuxcpU7kJ6+1E24n83NfjQXdwwKBoZaA5csSs9zs+f8WE5oKAwHvqHb6Bnvw067
q2GQNdZKrYkhkJjnkH72ItNTCTozcffcVJqUW56K6P6bRPU9GwFZNnY99sagNMnuK7EeVbCE/nZp
DavNUo7IL2mfJ7qTIMFWC1f9yA1RE3Us2pvcGM6SDLCoOYIXYpQ44MgYgYB7dp6CGgeql7dPVnhh
pJNZllUpBEuScxKxorGsBkqGa+clULjAuzh3QfmZYg2WbpGG56K0IVtubO6uodYzs03B+54/2ZnV
bBo1yu/xwtSZw5wmqb3exCaIWeT2ECoppZTSMnUPXnb6MVoaQCZAbGJKnb+oPFikmpPhHAjO+vFn
ng7G5Sq0QQ3uKR0UT+HGu9wR8WASEWlm4TEL8yTHXx/4tKtRwDeDazFkq7p1vL8iF44tddn3oEzn
Ev8SV5YO8jZQl2IffQzErjKbABOpgieMx0rCsvI4VG8AlXZ4uJtVnXxpSaUtJT6UkNi7Y7vwmHLp
HqsjCrF1RHZ3UM2X4sT39fsn5hKGB9FK+kcT1R45TqCkKH6/Xw74pZw/uOsXWTIm4PO3gnvurleX
MaYOqrjkXp9BZ4OMUVQDD2BpBI8eUNEJMDAE/bOSG1y/hhqN0qFvQY6k0f+UWOf494s7hB22d4cM
hMiFj+/zAYM/oehk54y0DziKxl6PcOl8ZTUTgI7PLq7vlOoaHRUjy5K3eR9c3erWISJmF+hYK+bh
edrFGQggthex1Vv9XN6Q/ELbkKlxdPv+IClYXOzLjrAWtsSF+yrQp+UupH7RNHoqt/sQw8lx2S6F
520rDkVAvZ2dJZZo5RVVxSS25hTrdZPrwhhBLBIbXZppKTGaQAREyvNb+SvI35P/Zd/4TypHADOk
ddO++8bAb1Iu7kmp6AIH0o62nxIH/9X8aHzvm0zzcWVyP77VIfVKojQSzOQhGD6A86B3aOxjrH65
J99Tv/gPDlb2hPFkPICptIpZ3ayrI039qDXau0M96/OSYIXH/D3o8lA2K+JJnhLLpn0ZuvD9fdVn
U6s4sTCPttFnDMYQZKUzvTYN3ep4AOgPSFroMgvBfhmUguapdDicQ0LNPuE6hVqvS2vZ3aaBDXMH
wyPiwWhPA+j2Hibw6jbL/IHhv3ZzpnRkQt935EKriyUXJI9uLBJW8PkeYjj4D8nj9qmjMaIuDyNB
Vj3ErtdP/Slj7Ff0Ms9v1LgSuyYoMtVV64EyLJZQI0OL6IW8CK3b5HtKydVgBDppLZqEoPjN3PS4
Ivi7/Kg8Zboq98kNveUOmw11CR8uBWY6aTF549XllZPXrI9a2bgMCSzK81r8iwZPVzzMEq9QvQ7s
6KnK8wynb4zghoKLH4q+PJehWldkPz2Ta4dFb5t8mHcmshA53CBk9JQoOZAQgo5r/9m6QAtY1spT
HCVa1CD668Kxz8fGIvMa1QttqyPrS0wAFJmWGrFii5DreoCQu6xv0Evqi9ULvs7q0MEArpXVPLP7
Wm0RM4zHWypb90D4onA3D40S+gqK1nFs0GrWbnBU5c3ulLiIrxPjGFoz6i/D1OKoQf8/4gG5XViA
AuE2bH2tq8e4ySwuyo1A08R18Lb6QtbHx1Abaepj3Y7mvZEtDPCHCUZp/I01o32/omSjvN37dNpP
Gvwhx5nMULMxu4wdpmIChvOfNYMHNunkxk78qa+VHPib1rO4a0Nt1IAA+dL8kDKiQwzyLNK4BloC
I+P4UhNY+G9bJ/EjDE8BLSUegWb+5mINui+G4j6e7BtipHRgsiSGtiZVgd6RIDmg6d0b28Y1xsj5
8DNmMgZ87hkV4h2jb2NaOfYF11WwDQcxx4QzO5xeFz7pjeaJFfJGObF+Dbt4Z8IT2FQyDWPf0Ipy
d3wcuHwzKwGG7YDpkRROfrOlRxT8MXR0iCrwyfi6mrcDEsyJVGNR/zcmjHOOqBirhqySqwG5nhNw
QwDa0455ayaPJb1pFwME+/a4iOXQ34scWt1dExSk+VWQP2JUdcFoq3bKw4wMfMJXtA5kAFyh6MyI
BAJaBdbGGvUMgKICjIG6znxVom3IkKuYVHCmHYapWLvmRSSfQKYF3NisaOkxP3/rZgBoHR1ALKWZ
9Ff0dMZodQD8cu7xXm8GeLOUuacdazflJsF72a2xWHI3bYreipSNSi6xXAykU+w6soOHw6NqRJt9
SdYiARxrJdgFtfYjFok9eZDrMJOzPA5n+yvh6vNVFvIJAQZXfX6/AtJ3ajHbxVPvNvfRWvoUmGno
VlFPFUBCbHhrYUV2g/RM76nXLcpy7inJmHXmL+Gz5CURjL8yXKJ2yxFLNSdsoqlCk0yNxXQof1IQ
HooquFV9DyuPukUkEpdymOoQIyrAxW4OJZM6ZEMZbsSuYfxo3thhBaieTi+mtiMImq70BvYrsQSU
zKnhaCVbFrfYlO2VOpHXIZV0POqULj6oSsotig71TLhixKG/rY+jzBZmO1U6bNIYovBGWtkWc6XP
YTyhQ7OkND3jBwcBQr6i8d2aRXOrFckYe67y6aSCI8+l204xlawODIPYJLCwSMQVgjART8m02K4r
vHWpP+0wKRLmZ+ypnXrFRJ6OTQsU/ovTsrLMZawMrbUfPsWUWcbxBP24D2v8Tj/fdzaRhh8wGqk3
qPyIlxFjXHCtKPeNg0u9vGXd+ZSMqMOEtKF5IR2Ju2jtfjb+HLuzDfEQhbEoNc7z8DdfmD7pyLaU
1itHlT0yDxp8NqOeIw5QgHj9iRp7s/4aIhpTXjMtS1wviH0/+PFON2+nG81/lQjERQCoj40q7N4K
igCWDL5fF4lXbdPSnhpSqrn38dJVIqMxZO0wOe22jardxR/huB+2PTY5poJsx2P2NP5J5O48RGex
akBuLSsqJt2BExQ98L3TvGkdJkgqeaTzFp9WdAsCb31DYab9MJjyvxPBukmVcsWSysbhJyO70Yz1
q8JjQ7jI6MZ9OLlgc0aFWIGN5Da24EUXWWawTtRY3bH+Yux/FMDn/WSl7vzBXqI4zE1lnk3Z6apy
wJUmKDyBPbvCs8dK8hB7E+iOczZZRRycuxgt5LrmAksh15gp1ibwxR5bbnKGp4ftJJJK43/zKLj9
pUh9Je9ZmbA1xnlVOqhtzlqcKG2n38J/SVSzPyFyDpkKFBGqRUjOFHUGczeyvEhVCk1z5FAEgkne
MTjyJDCYKBYwb7PR/+isWSUb+zFT1PVQ/G3uJD5SmY0VsUyKJ18Iftg+i/fxpMbOC1aEp4oYZ2R6
gx84cqYoe7vagyWZh8mduU1QPgpo3f+fKpASTHsmnRmoKSeTjQgv8kLdo1RCvaCcmhrrzdertHeD
+JfyA0zyBFkqpQhlTu1Vl+QeP4+nN1UtzaZV+6sdC1cYgljLgP6ueppW312DN2LlxxaB9Zdy2wek
PQd4Zzqn80ere/kDu43gCQZpspnavYbrl03qSyBUiWPFonD4STi+ZukeL1gkrQDHbACSdAQK6CBv
Um/SxWYNI2Eq/R2AwvOm1zqCuTzwLgFqaFwh3Nxr64ySPLgfG1GvZloFk7CqlfWbiPNDtoLWaMkg
pCM7NkDPH6SjNo6Uw6SjGH++5OwZyhAEnP/LP8grqeP6Zol3hBwUxHvDaS1ZaGbPk0S9ei5Xd+7G
IiYUqAP1DOtZLbtSONFtpKC9kLbzhvV6o8/HGZuz8avA99hcvasFXkS08i3aN+J7tWtjh3eh1G15
BQ1WlOPqlvf/1r05pczBaQXrU3MY6Z0q8NC3BjSGRp7BCbo7UEso0lTz+tCpKz9oPijPMDzeprGI
qTGeDrvGC/bJLFg8xYwPAPnqbn9blY/ASxf3ci0zhqxV++MZLjBfos6Pf0EGPvSWqOdeVjVE/ZW0
7gNWXbP2oewtP7cZQ9fehbkyusxfzuzxs46z1gnmXNZyMt56o3z90po6VYtJOvgsBq0qz1ExhVg4
QY58b4hTCRLHAt9ClkMgJUztRdoY74aHKpixE+xAJKGWbHlW9IjHx/rRdQAlI+wa3dRJgxhIp120
GzB98cXd20vJJL+sEAdEz3gqrIaLlDBIEuEqVhxbXE/LN1nKPprDCaWMXW7U5h7ZBNXmdNhQBsJs
zBeT0k6IXRsa1GElaB0Ck/5UuSvSOltoEZQlWcEQJ6Ini4ID04Y6PSlxVGVumT7FM9UuIUAFq/k3
NkdTBlmQ+pAncgGGFFYEY0qTzdoZ4LUtIAwP3EfLMYESEcUtMBDzVWKuKgb4rFmQVYksL9jIyoP3
0kUXLmnlh99AbbfCow95t7vwKcakjpOf5wgoAwFTkILBTjn5BMO+ftpsSq7iNMQ73UWOC084ddjt
/FoqTXuo2rnyc7zb2PU/2RGee+Z1u3DmyhZjBQakHBmKYqodoXjtqktTvYSSGwfDWazFVpeX+Nlk
1kFLpxgJqOYwdcS6dTnQbhK0oCcUm2Q6e0S4zE0vrwKxtnhb4XkuoEWVuC1m65QExWEcFjKUgUot
SLDwSr8cFofiRQp6sZ5A8Dg1yztceDcCN21Ff/VM2RdNEorSoxVnxENjrVKfeILaUYd+zU2AYH/a
Wj5L+a/45i13i9W4ppclByA1ONWKuyopQQwsPmdmOzX21T7ErDpRG/qS6HiI+/tYKa4bfYq8YWt6
XuhUJgK7iA46wxT/XXIlAN7Ek2E1kfen9oP5Ih+ta+Q/pTdQuRyjARp0lqYaV4jlYz113XGtkrym
x1GENOeqIq9uvGQA4IcpjHPhERinVDXm9KgjY4cLnUgpn4V7/TGXyZUtl7+v968K4u7/dQoDy1c+
zcKWZmz61s8hG6Lv6zzUDxK6RjhINByaA4OQAvxBXot23yUNfPkC29xj89jImHmsuLM9iyNnLmNi
ClecNTgTM5k6CFUPWdngTcp/EF6AOlAbo3SixsTaPDHakK5v3DHGTQrMJkMRm5CBcK/slWdKOnTh
/m1PquV5nB8HdjF4+wF91Smb5qQwvF3Ajc4a+0zItbboqgGBr8ftj+ii68RFkGkeVNBGj7Y637+/
LeF1YlT1iy4eTlBVD/Gdju3q3vx2pW1cvADAflRHbJRFcD33H6l2YFjpvHKqYUAZhg3SgdLxl+nm
RBxjF7b1BY7QJs+iaDh1Ko65rjPRLZAb3taQRkIa0ffs9eAprd+PRjSmqim74s4LIYGwun7YcJma
YKbWPgP1Xlzm5kozAXG0zXSYBvWuGT+wwHdxSHcfxKZFq7MuCcQlzK0TZRabMbzt1Sb+lxgZVg75
6a9FEVq/mXO4fkimJHAZKxLbxpd1rA5dNGxToPL5HPeLEz9irLIKUZsay0C6ANmh9dPBoUtAkguJ
lKzdMxEC37dzDe8gk32BUZz4RC9rs80jrkxIyXHgl80uuKokZOmNTDHNtL/c/KinEAF7KmwpJGbd
3ruDIXS1YNnNvwQZ3KD0Kv/w/2zCC7dI4APGODZRV/LphcHnixowiL6X90gSTgKEM+Y7ksgH9YEY
/na3p/pkvVgulVvfTCWw5v+41BFT6bxKU2bhVg+AhcCAYbXlilfri52whQUYTIzMvVaR8rfeFE4f
491J5p1918538f2lMEca5gcpEr+qeTT+M/8r6N4gGLNxsJR8k9/bbZevsmOhiX/2YgLHsRtMJ4Y7
6pA//TvZZfUUYeenFyixtPz0T6wWYqPrALYNtdAUKnP317DnIPoToPb68sum8+809LFW/S8MerNZ
ryBusc07u3LpTpmPxM4VCHya3t8xAwi8wE/CVswaO7IZHbIVkkfEyCu34SiHTeU0iaRKpFdK4OJR
5zNwiGbKupxhMGTwaC1lPU+tpihym3fNKcGwsSGfWaQbdjoKluzIARfkfhkIOsJDB3+WoO/oLMin
bWB0KcR3jh50hwJRCPZX5sAQLmPHJc5LQ8q+CSdU2uNaiMpabwZgg6WOG8aGeHPGB3vzhp3KGAky
9OCraEzQfU91HoWmm2I7UfxmfQ55rKVgkt5dY6WYoKFl55lDL3Grq9aZz8vdLq2PLnxNbkvLACQ2
V6Ot0B0crV3MstXNX7dIdq930pgs3R5WGE2HuvFzUDIYfZu3TT6LBRfGYVx6VmAS86Tw/6103ZdW
ypTVt/5ei5W/hIg++s1Fd87wBGEEBqbnBGOHukGq4ZN3xajglIMBTeqDd17E0qUWMLcbsriPVSi9
y/rqfsXbjAyTYTi+9khAuQAvauMujoFc3WbenzTrslaD3dT/eYojdjzz1fR7CgFdfQYhRWtwgAQY
MrB01JOfptW+FrmiDzseJAX7/kO7GcaKQRyUA4QMQ/VXSbxvO5U+vpXvUw1cUKvVl8vTIyA+TRxj
r9Ad1zWq8j9GDrf3sqM/X1zR2BF92LFQQ/pUR8An2FccYlXtqugZorrWve99LcXyDKxRcS603CCs
P4HH/6RA6JO3D6JiLHF+6tZUcoA+IaTRqBs2n2qt256wDbHK+ceL3IlKDYBK2Rdt22Cbd4fYZWOP
hyjwr77i9ZsF8bMnB5BcROkvtibmgn1m+q/9x/v3y8uMPcxDibCX+jx/XSYmyPEn839/LmiHvB8N
lSDtzqJe5yD3O8DSQE81YLLagD2Hup2gm7wSCAtVBlruqMfBsB6/8vvd/jl5/U6ZPep+XKobZEC9
QQu+JlEQgyLlfUQrhZVTJvTHOXM2+jKmK6sqWz8ZCSs5p3TBsAsSEiLnavAroGllx94dtUiU1+UI
L9Ldzj56UpMInxQw+3RN819A08546VSZiwnKQ3S+lwEdVRxKL/fK1vVouKRGG/968wZpSNvRNFM5
g5VKS5rOEOeEiBbuSm4+4E39JsXJq9BOiwCPQfMjb5uYlNUz9YgaaECLF9KFN+gp/Zanmufqx2TN
6ynXQJQemWInDPg4WI3biMXdNFHpZ0u6CZszzLrYROb/1YcBcC0ELORE1YabR5777S1orpvDeCQQ
eInFdjoCqphsF+c/AfPVy01aHzyslqfN7nB4UPR0wIz0xoTl7EL8MKNY/DDB23kbRbnjUSBndXAK
PfXThV+jTqf7my1GCSRC6vTElkr/0n7vNNfXJxNJlsYrHD8dQDhD/ECcJ+BnuqVvdkzky9iWJckD
NxBdnvz+8J9oOvFzlXNpiDaBvkvJ2tP0BCXsNvbpute5FDrVBeGtLof6+g9qo5s9Rki0o4EJIKWI
4AoLRwjlbF5I9pm2nR2/StBaQnx+5qsed5SFvK9vYzlYDA8T/qGZII6tGawnbpxQBkNfuG60gwMi
GEphM5dbT8ZPpR5MDwhVBQ1yj87JCIer/uAquZJkZ3v6QojR+WI+6VaoNdobfXmDD6SIwoC9yuoJ
CFClgb04fKEB4KoJRAnfMWMwhDWSLjPd5yDyrwBRhAThtA1g05tbae/p0TaGI16VuvN4IQlMpSnI
h0yCfq/sQEaijVCREszMKkP5qvJL1zGOzubHQ0nxk+rWYssV4vTSmPisDRDtdXgQZe0zpqsw3pN8
5qn7pq/09vt4CM8gTDhkBugNAVJpYDPpt0cagVEE0cPpq75fab+OontWA4ZIwTm+vLvgJIioK/b+
jBUnvbOrxCNRzAZzq6vojXXF9QsRWL0qkI/OeYwDXCXB9IjTjbnAANyeIZBLrismuKzaGGsIAKOa
sUmpoSSkaWpw8smHWl0yNsNzZltvcCZ3Q0rej4t0rh+h1/ohIhAUQTs4ijUjpxboWacW/h4xJ+nr
azr6CYLc/T6jtnLDVSlWvW4SqPNs/yqTFP3vYWwpHk2iVMvkdrGk4uuNUQf2br1y2K2e2FolJtD9
/W5orWXxquaaC0QpZKU7/yRFkMQ9IksDTWLv8j0LSetx78rvE5KupXJx9Eaw33Ji3aPYUOzwB8Gp
DnHygyEa2v6Mg+m0Bo0ujfik9cgAkqgBdsN9oZ2vMOL6agaITmvyccoa6VWWt+jctBPmlHJEFoxf
ekMVysnB7ANVZRpekKnIcILDy5nILZsnBL/9C5M++L7OExCvSrCoIY3YIG1/omN4NOMnGOFIDtq7
1hgjqNB7hMsOrvWdsZE1NVVngd6j55iBulVf8TJ1bEbMq/66eS0Nn5UD2EtHTK0H28WbmOM5rJX3
Yd1ULkCpkW9NCvNzNCooca5K2CD4IcmThYp4OfIX41Q4Ntn0qvGrSY5ika9+K8u7H5k29gBDosiM
QYyDWmQ7LlPyxa6RQg8iN9DQqrYvLfvd0aBEzec2VJIntx3lH6GKzk/6v+PbkiaqrZwGgIvZwrEZ
078U6czf19hJeGiLhSuSx69ISjWYCO1gtfr1emzVv18aWtpMXTcEVFD1KKzB6b85C543G8a3Ltt0
9//JwP+crwsJru1mKRoG8RqSC869/2vMw7r0Sl/9md6rHyrRbPaAaZibbaoInEDfV/2Aqvo38iml
fqypNv01o/Dh89yFpSuOj0TBcCUKqGALx170c+TqPRgjnc7npW3RcC7u3N/ojUbP4Mxf0pOQxEM8
qE1Y2P+7Be5hC6Qd3CgrfS2pqVLZOfzsR0oG7NHzEtmM9woFsC7PJQjiRsCB2geKL8M5Krz81k7o
HqdRW/AuJt8zroKe9Wx0XzRAVzqPZ2J8WFBmRSWvZxRCkI+VAnQuMBxwbKe96VoRnP/khcP0jzJr
iyN3BdZIajWauCPeMp9/8DtPUFFdKu7v0UVPdl3xB80mzyduAoYl9I+ElQdQOLIdQ+daiVMbUnmf
zAbm8DgWl63pV1kZe8l3++NiL9R9/aWtcfqsnbReBoln7tua9Ymmhi7dBF9GSvBJfI7Xn3kUZHHY
/I7kyCuU+r1HidiMrY1jHqizYm/kXRRsf6KdUic8/O5ikjxkhc7vM8wKnBfFjUcYadMTYil3hD86
uVO0lTyK8ezq9O9DuOCw/WDt1du788/BB+EgJaZJPgW0+DHDEXsRh58d7Wr34t26a1CWYUVxOFHG
a5hwg+qZnBoQ30wUmTztlweEXPCOJTnLq0zJNDzbY3lOwhsBmLEmTep+GRwa6NyABAlCcGKngAzs
51CvmO94AJh28VSdpHU22gg0URcAKB9N4CDbPx4hTjKvuNtRNvXgIOd58ssJCj4c6dX7GaCPv/7F
b9l3c2p7aDYBWatSpxFMPl0RjwJQi21NHOMONPLuMXLcH9EhDMLL6lj+VOffmtk4mz9obl9DCb3C
/WPi4copXHYCIE/pCRdoiA3v+tu1WXmYIxBjgriUoHhB8LYdkwcdPE7dG+AlLVCxxp6nb2ja/KwU
h2cjCKqSE9/Zv5Z39Rqrh8TBr5bcDrq7z3d9RDq2I/O2wNguWOgP77NDEUTPzD9Mexpz4A7x32w5
fEVokl3NrAPm1Qq6UAC1vf14TqRaXSOvwaSM0QLCykHkJtORLs+rpqe6/7AHoSBpw4Oc0Un/nZeT
pQNr9V0vohyc/IwTbkwWXcsKoEckLvmkfhKGCHx1UN70t90jzgzpwGmRm7eUmdACoyvDiCmvf8YB
2jgdyJ6geH9KMdLVcdyee1UaB1id5V4mOTLCnVeN3+16vROY1OSf61kxkD1Fdtvv183rK7otz3iS
LoIP8a9WlII8v5ms8UCF4VX1fHtQJySQeeG0NQPR3nBYBOeMC4wnEIPMkdJDzaDsbOC0DjLAakTX
ux1zpCf7sloJGxsV++SoOHdMITeOGJ5hCtyGowMJFRJVHOwAw4Egdt8ROdarkdJaYFsRsTxw59Od
RI9eUCNh+U5f3hlaO9H7PgGRAWN9+jlxAuBfDNo0hzKdYo+IjkqIP2YOHJRxdO5dmsNDG6GwuC9R
GVZ0+L2SDEdLRNr9ghdyuSKofzN0ZwI51AINiB2omJdSlhlJv1DB7yKtwN8DsRaxPwGwiJrILtD8
WUNvlzD9FEiS3uqm5xvmqnaGvuRQCl2hbiFmxkOHeXJerXuNecpPg1JNS/cNfJ3JuTHyeAA/+w2Z
ieH0ppDu9f3BhvEou1Xn7Q9WvyknleI1aghhG1LiIpgRUW2k2J7LfvTGe2+NmSjlUn08kdcRktH1
wAnZKvLj+/s4GNQQl4DPcOSfZhtRg1EKbPBwG2f2+rPMorRtgHG+PKgWuc+soXGmDpUJQp91wVG3
1YNKuKcLAk0v6MCkNDzGLgM3jUjR/oojCiYUGUPOcNqqE1b+ZGL0YY2Zjunl9/yywbRAK4gSH4va
Nl+iyArfmTvXA3Ct0s+Ewih2gkpGw87LmdBmv5tKBsy1wYMezEKtIGRLqVKlkvuSnGg+Ex5Dcp6n
3SpVl+jQu73YEFXw+e4sKrvVmS/b1eMOuEQc1v67boTCdsrRtohZbnTk8FXhIjnlfvWmPA4Ik2zm
H+dCMQ+r1Py3Fi393rEEbxiyPSsD5pw/atfZXs4/A5c45/6fuP9UjmVs/+dJLn5h++2hiZPQTqS6
mkM/ed9f22KWsjtFQbDHrikcuHGLoUiazuSKzA6gAOl+3JBiKi811a+/kdZ5l2Ton8zVkDW1JpKB
hFV76/jUuDDByqupzZGOjhJuVZEPW4Foviwo0cwm6UM634fPZ042JNq9swfPXR5wVxO/ELKIc6m9
Q25bekkNX43Kfm6h2Yi9B6q2fJxdsU2u+lmTLAJRmFHprBcHkNeDL2d/xyBxLAYqtCmG3vZ25oXM
T2ZsFgv0pAMiEGwCcxiPBK9Ue7sKOd/aB1FqcX29Qt82e65bb3wZGAxzLK9mHT0kQFDCMivzYTw4
rwUPcvYlNlgwC2o/0R/kYGx9zIfJOq+m4TyM+a8ssOLFmCdu3AiXlEkRxuwNaj5hRTpw/jdX4E5q
qZDiBhOzo6c+s4EfKNjz1X7J6F1Vnk0DRis3bQJ9jWl1oic5YOXWb4CFvsBRsB3yfrH33ZnN5tSV
IVOAVZlcVqZ2eBS5dW75IVQTXNjRy7xpRpyr0NMf7eJnWHNF1DPZYFsiD0D/rzmp9YJeYxDRF83Z
yT3Nc1nom8LJ8CsLXpQ4E99Vn2jy8wsRISzDIoEbFhlm07NpO+t8n6YFnLdqMr/RUktBtLIxiqKj
R6ia7l8wxZYDtfL4MQsywAOg9gtS8vL1t8570SUtYkoSH6nwiJ2hKVwzR+ipTgSJfwil/URf1TZj
8xSMZsqDxxlmmT8IN821MYmlWi0Riu3PcRMLt8RS1X2EKShmNdpe+brMP6boKs1q3Hk+WxJFj5dJ
I4reUQNcLmZP3AcuAYnGnJVj8Le9iRbE+PR3B/qG8tnJxDmUcCKHBVzuk14B88PMRP0wcBwEFxM8
FeZqPTO8BYqu2P1Rvln2hPZNMc7cG5hdpRvVt7eldwhhzr2QCnnRzedBiuxYpHpHOQZhsCVA7tLO
XmJ7vQxw+pnjqYtgk98BJYq13VehWcIkYOZwpYTqPW1F486E2Kko1rAXrrZ/Mn4dIjf7LZWHeppO
gvyFB9GfbTX250UhVFq0dSubSn9MO/oYG5XGX0EmlbJj2PJQaQC9mWcGGqBMMIzESBS+8etIRadb
YqH8QvpMXjiUO5v0LydVmVNujFdG0qjnW2MILdh/L33oFQOI/eEzPd5KZdNmBk0p6KdV9AhiLkZa
zoJmEeirKN3dVJNsaL1glX5gpsOeaTpqHfIqd5NMHolZNEtJxwWmO/xs0GvuZmrbiY7ETerypSt/
ninLmktzzxQVqms0095P6Qj/5yqyT+cWgE5Pk3wbuVjwueCc3wIt+wP0Uf012Hm+4QHmgziyhT4t
d3vRLq6kwTdVHdnTIHXONRpBDWVYb89YuyylJ76qww8Slh5uI3eCCklPDnz0cX4g1T2l0cXkq1uF
13X+nvCW25R5OCakqockz82o3wG6efOio7ZBbkZxoaapWQ/awrLo5UHuj1QCtN3vzsT4IVDBVbua
pEU87wfJfgRLW2dZUrYDTcwOcugRj33eBX7hpzFDdb+BYgzKTM5nQ0eR3KnE356GQeAmOobFlfcm
wWZr6XGFVcWKI6U4JOs7Nhoe8HylwNWruhU9gsVGeIuQyI+kTjoZ5uWiNMVChEBeIUNJQwnuVfOt
I91G3DGr8c0JGFNNvZNpibGAyo8KaPEbONPGt7YQPqevPkXH9wSWN4GStbfcmRrTAx5M6qgBBYhp
RyY5hcmMrEP2t8E9SY/yfFoLCOQd5cE8f7ZoJTEv7WVXHPe/T6eGZBuHmFRS98nNDiM2B5THQSvI
xU69tomrmIDMpx5dbNi01+C+AtQMC0JBiDHG54kRM2xksurXSuEDoIS8F6uFtTRiM2Ahq3Ofmg4L
k/nMGZ+99GeWwg7FhIV0uIBJvHNEbsqGNxhcg3drn1Teh5KkO0PQWR3YPh8PbFhwuKDz2XxsuVXA
830gnMW/fsx5linqOB12gI71T2VTb7bOU1mNw1vw3WyOXWhAvv7bugTWuxe+AQ3c5eshgKMrLhpK
6SkkUJGOj4Tpc+rh0KQGj8Omrg19OmgGmNChMFgGA9dQYn48L6IlqpKxHcWsTSz/7BgzwSmpDioQ
Ydzqf9/W0Ib7URFHxtLlcaspQPx25bMyL1/sAgm57Wne3tipFRfadON/bOBLOTH+Kq6KJlMld9/y
j3zLugkfLycdhTnwnP/Bd3YSQtIKv8jSIO++ON9sCOXFIUukZEz2/BFRnOYvGqC0/aQ1hNJ/rQHh
cb6DgiUsiVg4GzX4mMGWV5ZoYReqOZkDyqA56EX0yjTLAxiZ9VxtlSdfh/YO6C+uYKUdFJ09MhWs
1sH8Q3v1zTWZXbezwOM2FKFM7EfDZ4fcPLVWEEiqJI6SyV94i8IF3j09yhjShxejnxOyiC45qm+/
Bant7z4WR49NURD2pg/AETac96cFJvuAP3+bx2mQ8oi5VyozMoOrX8fBiRdneOI/uYPtm1aKXzkZ
xqMTi7F1jb/68NhlFsDnQkgsTfmo2kR6vLS8Ak5s7kzQvHRsuN/e9ZspyNznpbO2cwhUAXMh43zC
+wkPEDTfGoTQ2wUuOjMKb9O2Jc5BtgR99eopJZaett8kdhflEnbyPb7IBJADy10EFoKj1ccw158W
AXwJioC8RWIAd238aJHrwwqaT4Z2N3zxLLkGIupiRN8A6NbFbO5ukcV79Cy9CUW7d3dMIhGK8nQj
OxRoGVs2eUS2NJy23p3hJtguXlhq7k6qB7e3kmNLD57zK6kl5r5V0HlTJTg1r1NYuesmcg5IfRDV
i16thr1Ge1PdtAjHS82Vj77LYyLDaVeZ61o6WJ3kDO6iDjezCjLwdG5ql3DsngCP1csy6tRxcj8N
L+skSqZ5AyAM+watqYdMkzYVuoeBc4vFoPKiHc0k5B0EluH2ftXEXsZi7wJrxwx2aafdMHRDwME4
ImOsXfBLqa2QQfW8WSdeOdiqdgPFevJXAqk7hzXHWjNktVxm+xNOipW6luRp/TSVXV1ZdmMl/y82
qIhzkQnIr4KNyBeTfWeLcNtp3POHUCYCMHlWSlaI3AZZnx+eSB/4aD0iYkRUtqxjxTAis6sSMPJ8
jhE7DaZF0L8Z/bx0FkgO4PT0uI1Rb4kZPWR7N4EpB343SJGerISGFU8BLHM+spiGvKfUSqO7JKnV
KQ24U0VdbfTVw7p4YfLSg7B1SgBOoFpSq3pPIet9mOikeliT6Y3Zegfhf/CU2QYpVb96rF0wFgjO
FttG9nGlWcR9uVkBzhRu3Z95nT5r7psi0M21lMFn3ihq9Vk2hM5BdTe70EXPuKbCLOw/MbN8pQvp
LgDtlTNz/82D/6zMYBsnROXkSePc6lLTVlo3QYR77ZEUp5JE7a3EFR2z+ChFIVcDDM/GgoGIBtcb
ggtGNMn9Sd7Q/D4EZ1FP9NbFprYv/tpkCfC2Nv0nW95xn2USfTFEGMLzGneZH6BaCeGM88dGvfL8
FF7SiCG+cRzzwVW8zCXDdeHx2BgWLr1XCRn1dR2fadd7oCN80JBckiQNnhRXbHk6A7WKdbDrqeTO
4yv7Tf7oy2H9wwYYU1kM31bKSMFoT4zt8k7hc0EkCKxETa9KsydJzY8XTsR3qqGr8QLcHb0dhnFJ
Kep3kc7570S+oM5G4hFcjO7kInozfadKq+eiTS6G/0AGYl7/65OJn3DRqFX5XfclCFOwNk4DcNlh
1qYzBGiIhdkIMmSevl7Hh14IaB7jdXfylG2z/w5zxUaJ7QUfN5o/CaL8O0r25vvQOvrOC30NmQbw
fnYrf0tMBkc7bxPz65m6z0hD5xUuPz/SzVEKR1nKfWvFS9pLjWYfsRzOv18Wl8hJW45MfEBECc9Q
WMiLKBMNg4g1HKwT9WpYmClO+mZ7677RBHy8cEV7ca4Dor4QJi26SC7coCkHk8GOgac6FkDPsyVN
dIWU5y0KgkFRELnXREUOs6Bi8oD9TsYfgP7Zy6tGZpJCkMzG0aMX39xoFuN8TTQNt4WLwO+rWemT
aiAaqIi7pqbI02Mbk4qmd+wftAp0sRX84Bd/Usq5LSPKh1Dy4UdHPwbSHmHrxwu5yRNrWVWX5o5P
8mfR5YyKI83jjbD6jfKG4OFHREkyW8qbLEc47ZfiCZf9Nj6siabdoqyWicMn+zDZDzoNjVgqbXN2
AjR75ZNYjzYku0B4STkXpC+awNZ7wCXGT9hia1WZuV05daLyADZ2AtmsqrNRXpn8Pg0jy9bqCU0x
gZP4i7Xvk5EGd17cQR7drtStr2G/2anwK1SXvOjn6j5TQDklORYQ0O6+eaBD/qZyrD9EGHaZw/4R
h6eYHyHZNvYAjhxFolycbvjgEmBVpDB/slRVNptZtMesbWiKwFF+9kYJs8HqrDEl71Ooq/UiEoiO
0B1kH7rbVoZheNlNBqP00rSkT9CHzOFUTq+ID8VdEACE1CJF9UxucrWaRq37tgwQpaJx7Z5FuG82
yYHNlZBXBnISnY73QCVwQkoggEckJHYWEwsALIZ9HT9m4SoLIo3K0utM8UWsumLPb8PY9nroK0HM
i69jmRui/j6l63XVeRGeGYkjCFvrRP/BTjGCoEnErg4SmM/oMwIyY78uZa25frhsRRvUF93+3Z4A
j2WfskendfdOnfYfFeR+mcF4ugTGzWrWkowdDj8PiUXwQXDgh5HjWJ56Kgz3J+Fe+zW/M92FwszH
c34NYee1zDbiMH5BA+b754qzuw8JAjum2hX65hO7+66Rp1O2ehUcGIkJARo47gKq2O1MdNbbRP2R
tHbkr5xWFdxe5hghaYswIK3rnKGTMoYHruRpY83HYUmBrdeVY19v54SefnR5cW6cMbMZ/Q1tt5J5
gXD0e0OPZWRlICpKFIUCNrSqJHQYWNgZRCg7f01DCZXtCe8ax78CYR1Kog8fVrKIt0CYgjTXktri
B240uNrWMwnXFZ2Zq/UpSA8OzsQ9WSTj3AvF5qFJhPJQtXDfR3z2ms03WnEFTSHoqnw5gMQnuTHQ
0lrPuNvJ3+aex5iVYfbA41sBd7DSI1yTpZz5N8ruM8UJkVud1MDR/TVfwqQEcwm9Qtn1mKf8c5md
CmfGHuv8udZvDAZ40r+ZoHOIrRDAjn0Exxg9stqjKib+ZbOibYTSdvY6AY0YcqIjacqvJacqwUmk
6zL6fIQ8F8yUyVfQu5zmpmIhNeZKFQ0I/3+wC1mx0v7hoLqJ8xSdyNKKOqpbzd7dBL+nQvjZXlmS
d+vChKg9gpIvvCr+sZQSQXa5V+kxOgMvL6DVn0/uHhMpu3FrjyCqwC7sSViwtpnBpOyYwlOWONl9
R5kfiUX2LWzrIjV65X+1Y1QKkEm+k8ihXYfQ1BNEnbJi8wJ6dglGv1J9x5wYZ13XXQJN0iZQHsc7
EPwdcwFjGedKI4d/jRT7mNeB+CXD7ot2guND9Vo41lz3iwIAsfJCgEg3UpywEW3Ll7Hesv6LEj/3
+R9dD/7nHwibtfY6zcH/2KJMTzsimcM/ha4VKmpVY6bPYUTy35vGNRyJ5IWCA8qbFcNFd8Gpy8Ii
JF6vPrMS0rbi1Nu4wybaQjYd/qP7sq+fRmy29MT7dhBCLalgeIDNUYt12QFkVMUYlauGa7+IAvEA
lUV9ypPuyGNgo72erxfCm2hFLvjKKo2Gb7tHWJkvgpFH022hp+jJG2ncIcmFbVhOHOWApQeub0N+
/eQHV5lodapRk2DVSiGEXYj+SjZQHYhBhtBoO3o97PVF22auOjbDgqshb0IuBmVu8mSsGhcxa4W4
d1Nl9NZmUQ/MWX51a1mC4XWyhmDOUf/c44QUHYlwzvvfgYC4tGN8jeFP/1qzzDC6oD+5aPMNCnWm
IfewvNtG2GEjzcWwDD9eTZnaDdKZNNYSRbIOGMZBPGQginriZSu9yJfezuyRhoc4tZxpJ+OU/taA
igscLB2Ylcx1p/arG8cHz2CJYp2IrT0+yHgHCNKLdvU1O4N8Itcb+sM6aFawhvRiWCCKabR72J6L
/AzP+3dahGRe1lVgfIwS5ODaGae9qNxUe7muqnminz1+q6G+WRqPadzGk30etJB60ySu52RJZDeZ
x3rA6Sc1s+t2Ss0BrHRtAhRMWqufnTs7+VfHfNoB8XmwQ6BZcx/xvOjR8VjFv2Z5FWezOoFwImO8
rUq5lw9SlFvBaHYP8NMgaXBC1r4WyQIyrQM1erCW/6OTtboy9EXM3hjFUyhpSHElfpZOOVp1xYi7
wUvoi5NlEH/f1B/fbArau1lLKsTBx5zTARxWtfBtH6PrJFYV+DcpZPvxcsUwx59J/p9AcYVn0ABj
8p7i4O0gNtT7GBWxXiuc42I+T/akvQwj5pMNhY0VXqjJTWAXvvGtnSovRuoRurk0t+xTBgh4gCTw
PRC5+xvZi5gyvciCj6MLjf8CTuQpSDou2DUiphCUBcNoOHCLIpHYB76zwvBfZjjAeT4503aUJvFs
jPlQPsyeEnN1W7lgVlPkvbi9ebcluaDOJV33TECICh5yFV+2DWUrEr+G9NEjQt9jxJNz306DO/Zr
fIB6/FvnqlP13agmKA2Kkpx3EwK6eZrAjpdFDHEYtGrHk1gp+JHTZQxVtsUP9xhpUPMp+P3EP558
x6HwOHPoIMoOygVsqTL7pbN+tvZ5cSqUOGVHbM246CdyJmiPHE4LefrFpDQ/n0lX1xLm3cwwaLBX
WU3YHmQwLaiCkEckZ9096psPyKYiRUInTTKF+roklYgLpR8+D4DmeBMBXKStNWn+/TUNN0USoGXH
plkY1/MPfHJw7dXTAFPPXuL7odY4TnZv0TweqLcVUsC2S1RwH96OAAJF3XvQVN8CjgMM1/Isq8XI
afnA0fkT0puloK8DxgngfrZLpHTlvVW5qqwLm3uY0MtQU3ANrRyvIeAws4ky7Dkux8FqmUyO8Fo7
dg8QtNaSoUMCxQeWduK2M7Zhm2pRl/DJHo9KQhTbB4eF8zH+1IJs6ufFsVYwztf/2VP4UllY5JYd
t5K2rNHfMfd/YLmUUyZFzvYAZN+vjhw1ENAwMZ8Wr4IaDc0IiVNxn29mTgko3wFWvKi/iJq8SD3a
DyKpKKV9026P4+iNafLe1Sp56BIt+7NiKQf51RwcmQ6FwzPlNaO4KAV2kCXbarw6NvIPZ2lUZJ/B
Ii2LGOP6hE2ao3a00ZlR/LSXs19agVJUP2t1PyBhVN/0CekqPIj2tdlBcK3P2RKhFx1IOibXMxno
+8JtJfMcZ1EH7vUny7L8leFFaM8h80/4Uzf6QF3Fsiu1Bme4tiROWJWeuJ6pt3HEZNsitdK8jNfo
OQX5MccXeNl257vBtp2LpuW9iihnH0x2xs9oFL1GTKmGurSFnOj3wjpzM2ZRMHHNJ/r/eZvMW46L
7AZCTmmo90vioJpDI57kkp2jLVs7wCiAK8ioxLMdbVLLKSOyq8XnU9JX8oUyJptPv0q9upQrVmIF
kFG9NyIG4f+LLbNwRMQy/ZO1lklxGAv7uhGhYaBvhJGVc5kX2HN4tQ6ddhn95DlJuLjD90CxEewT
hd83W8lZC5Ot3BAzUvaK9vuT1x84KHoErbQGkkI2LyuE1cvi66M25I4DF3x9JoblLc8CMzzWYfwV
4RAoRG7lLUqVR280OXSerFm18G8wRT0RMvY9MOfUFZUOqiy0qn0saJWj8MUjG8UC6O7v+a+eR8sN
ITeOB/00OMiIUFcBeB6f54MtewnUDztZfyTOwMj1zso+BLaPWkqr8rxJZMuEC/FvbfChCBrBJGK0
bmZV+gjK86SaeMqhfvCo/KbWh91vN0/n4gq7sTcUeHTHR9PXWAIPBOvwWfqbxUIYl9sT0W0DxR+7
jNKFIymtOg6frRpBdI7DGhsNIxfRmqVLtiCqRR9EEAAi0pD4WCt5GJdYuzvqWVWyIovJ4TrXaXSg
7oLfvFPXxmYl541pzDo/1By0KEfWSyKJk79UeUfGTYliCW2uN6Glj2as3uF/ErAkprrCl4r+9tQ7
tm9sudSkzK8RaLd/aU1BheKgQ/e6AfI/TMDr51l6XUR+D3NNJJYegYU0D4ZjU8fmXo5DzlUNNIO8
xMKIaDMONMqVQTHlChjr3BcSghjguXokt3K7d5/Q1Lug5ymZj01VWhkw2Vl9sL37fM6vRFF4/rEA
QJfLnrH8MFJWCj4BL/xfW4MkZ0PcIORv5nfdZq158yOUvCgCahb+yhjjPE3ZRI42pa6TsQg1LnQQ
F+GBdcQkSADvokVYeYNmHlpsn7TSkXlJ+kAqvK2gltBScDasNpyT+SajP+H88pot0hwtqetdsOhR
ELY8t5H2qIQRwMh0kAzSjFnI14Fy365Hzc4E1XJTNJRWR2uo6sqMMilPU6H2wjnzW8E+A2jyrRUa
fT0+kYWXoFvi7tsh83c6y6AKZuF//mBgF9+jR4OEP6USXRhlZTrhHMDbe9rGcNgZSMqydeyLLfH/
MUpROIhq2FLWGpcBB7Wti5YfS9h2s0mTHXrIy64QtobCdw7Z5D53rniyKrTB5lx8mnxP/R0i1xWl
jt0YshanK7WxyMHkvX8cBKKz5Ew297MeEzkerCTVi/qpIl4NXLbV/9vd3oyavPAIPeyvyH1BpFem
eSxY0uRBObQn9vsoFdPfDWviUFyBQlCMiy7EsaW2EAN0v0DIY6mCtabyAIDmNuZnDBdoxfucUOcJ
cpypLBrDa/c0W6Bi9d/p2lO0MNHWvznOZqGRO72V+mmQLrIwVoxbc5dZq4g0kaMkEz67CB8obJkf
M1eHVdeD9Blnv0u0pe/EgCJQwEaIvdA/nC+io5hs0bWJK8YIUYgye0Z/OC85ik95bh/DYF1+2uLS
ozqXDWa30w7CMKa/GExtAmvsIcLnG8gHmFAfRmJT0dmh3k/tWYT+n6qnUHPjhUA6docmo8SlBHTt
NOPNXhkY4exxOlDpDSnhAmylx1oMgmDLEieeAWtPt3mJwp/f50ZCLVMLWtCsyAu2078sSRJPsoMM
M8Lb1yvD1yQWzXK2LtcgEVPJsqJU+ZNgxwYfGFVJmC8xzWyC+PfO2PsvrKxkfZHq5CO2cvAwdj6D
k83N8fqtUNWmR0KebnzIpgSOECuKc0u5bA9hoctAgGSH2UDdvIBZaJYhC8aYchrKolm7xeoOY0Dn
4yhcZf5nOi/2dTqV9pbeygqIVtkB0gk3sVRSwx1da9GjoeVQZ7y4qDTI1o1FfsytJC6C6nIC5M33
q2rvHG/0rYJp5r7Lz4AbKILRyffq2gW/g2b+BR/FqeiPXgOCIlY1Q0FbTBvfW3w2L2nV41BrZIvk
EzYjJZJzerQE+0i35kR+NpHHkrs/rXl1q3DChVNtERF3tFdBxB1p9h1wZPVX3P1+OFvd1TvyjL/4
rP2dYhUlSxYZhFSQ/T7uC82pPWynpG7RlDZk/8TpVKY/BNznmkUqDXF0YEn+tefDyZRQKg2bsu4o
IWg+UN+GFyWwgtBAiD2ghIvix+aTKvH44arNmNVp7XFgE30N+k/Sbm3kO9KVwsRpFEToMRqGqdJZ
mkoHuZDbxjXW1gtJzdqTcCpbp0Ug+Waap6HZpYBkmIrvHIOAHzdnn6C7ErQh1fQ85MA4G4IZasCM
vUs+b6UnsqUPKjsly4l9rSOKKW9evqiAik3aku6jLepyF16JOqADWyes/Lk881vOSJOQGqC8+jMg
otJSngkf//ixTMw78M+aLKxch/1A8aO4PaaPrdR9zH0n8y2W4y443bt1goERXUzOVHgtuhWP95Uh
k+k2qVC5wxPegHyf495t7RE08zEsHyTamQHJrEJqubbeSSfVqIRrwxY10lWL/1pHvrRy2nqBF4x2
/fTIXoeEIvSp8QJhX4bDeh+Mp8ssqLPFmbPKfFQyQnLldAsqzLods1hVM62oGd8xzUHc6ou9Vywk
uAGwd+wBIuzpYRpc87mV3T6DvzNMvDSi1QXtq/ZOZitDjt9dYgdxbjT+F2ISNjkqctMmypl91V6s
+M0am+8UR0ebn9FsZXDQr9JaSd2edq6fDuZrrt/+zHFJA+ssdcS15TjL5pAmy7mtW5gW+rWKCtn0
yJnJE+SiB+cMSBZTkftkw+23XihIr3/8tbUXkgG25YAbCBKdiXU3hoRdThXcPX8jKIQsH2bnR3Hy
47o+t0jr746OwzoZ2uWMIWCty40GwoauOxIXZ20F3WC63j4AA0wTV9FGm2WK/jKnNTMUUY3U596V
t6WPR0rRSuTlUpcyii1g+OYs4AEn7yrWiIyBhNVZJoVLENWlKkzCx+Ozfw6QAKy9hQl+u/DhwAHR
myvh7Pwe1Uml+DOQ9gLKA0OqVsUWsFU7LBWktahwHP1MOis0Dy7EOVB0z+2kl8rmN2/fvYlGdleY
3yjwDkZQG+9H5q4NoVOw/DEINrDEau3C5nZ0G2B8fJ99bHKWDO+0Pl8X7g8MuvPeN+M4uWxmPSXQ
O1mh3rTFIfDl6gOfRO8cbIjCNNPupR+R7xlRiYlU/Hl4/F0moSVsD+SeLUxQB900l1hmxHPq9hZI
cM4OOQQNYJhskkz683w4oAMWXmJNHi0mGj4Z4dKBCnUGlRRvGrzf9+/IvQJ2ptiVXyNv3sSg5ovD
oYwRrd8cqDzP1gT04KAzdtAVobPPnNCvkAfeYyvuQ4lVKMpRaI0k640ErC45N7efs7csY6BHZ5Sr
oQU4QxYDGu4B1/v9JfBkuaCdPsQ0dh8acbNMgVLu6rSe07alls7uaLt2KowKX0rtocvVlcVH/UF3
Dqmw0XNlLS5tMIlkE7OLCovX9d/ndGEibTrO26FXPt84E6g7E7vTW+X+mRrYEqFCsNX0YQVnnS++
t1XinZWtgVgUwdsMxScKoA2UrWIdpLRdWaN3id4zkdJiVvJ2e7RaCPG0O6GKa6HH/58R76jTa0Qt
wtLT5SqUZzsO6JsN7vEAlC+ctRK7yeOJh53PxbUrllkmKN7C+ioaz1e2Nh54BWasVIPckMbyfjMJ
kuMNLhTYIpl15BJiKMlOAWZsd/xT5IIS/qnNyWFBEPK6He2aZVPjl4kUalM57tq7nMfEVGVVSLV7
3tSLOXYWN8HRMV7AydIJEXlBxvlBEaRvDvOxdvHF9D0s41YMqDRhs5z7GXxfvg3XmYHvbMDtFA/P
BfNaVzmcfA4MJL0X4BSERzLfKbkZbHRBEcPflQ3tTcNiJm43AFYzMWdKEKGxZkdfKYn1NuM/aW2u
bXefJBffeuKnlREQzYlz43Hjsvw1OWSblvWx/LL+ea7ZB1L0nfIqTnEQpLpHHPAWQ1x5+qnl+eKY
0hjIAZRpvb7hLT6cscffxIk/pM2YjLI1YnUstGfAUnB6DogXuKJj2ueuG29l1afz+6f3yAhumLx4
YiQ4sPJnk1Mz5AbEKapknG6q2X7IG+SFQGzA7EHlRSLvpuHHPExpirrUyTI4GTjOt5lZBSNoGh8N
N5jctiSc76wj5NcL3bQNda0cGnLNgfw/3Tlo6Fd/xKaY4IoTLYdGarlkMHbQdguGkY3Xfo8mhbZu
DeNN1KzZI/mKGuEljQCJMgA4xnyrXyduybIWHHIhlv5zp0tKi7x2sGDIuDTgF9wl4jWKeod4Oxgi
kStFjabNgnQhKNOQJMqhToiO0HeTgb7DS4myxMCOs2BOocKac4aTZm1MPsUVVrDeH70836es1GVP
LkZ45EK3plACfnh08gfZdCvr2J+Vm+Wm4XpZ58+uyshCzJLPUmMJ1X0f00DRgi9V3Y9ilwcLt3Dy
wuDD/Lw35lYMuuUxq1PXKvrFnxDEgM089S/YPi+5ixiidJVgSpSAMA2c++sPfsMn9U5HBb7Em48V
FD7b7sNkRG0DFDG/K1IupELHSupFwcu/BPdcInUEKFZX/d7hA7rP2oL2/2TngwdnfZ/Qy/TCD0xl
LD08YZJvh0IFQ86ST9SMDBR2dnXsIVVQS6l7FLGOqOOcBUVqPPAiSkWk71YYNXOo7c53gvkVt0Tb
Yn3iVs/BJvcA4mR2nu+n2Ejft4/A9YUwkHMVtmD6HiGdWDV2xBfjKAirpdmVQ7OfC7yiSeatdLd8
mHFH0Wml0BawDkMyg/EIjuDH6/3cof5VpVFzGJaf7KzwavBY3iaaHrsMlhIQdlPVnVDkFpGLsImT
9N7hBamBgnyIG6rYiXObSKEf4oMYm18k6wiC5GjBTS6jP3Hyb9RRrgl8vf7HYSUsI9KxAQFHkiUA
k551II2BIPe8Ow5mYwGPTLrLo7QNRwequfJScMAHkssCo+uV2iOfmocjqjKDmk8LS2Bi5YTYvyTZ
HPP3fmj7zLcH1XiMBquVOfeyojUimECYZvgRO9rOpuHZl59eJ5up42qQEux0kEX/bmZUS810R3uC
DlepkXN4EJEx2RTSkgCb5ohN46/uXgtOOj7oPvaNJMV294Tceza8QHUSCoseiQPF3ha6akLgjmQv
x7NUtk6J4ozUhhDh2MlYroDLqLXEs6CdLjvJ9Js3RiLF3goeRuldsgwyaEasLM3HXOgwjqERHE2x
3Oa9BYaTRFSenqph70WlY6K5vVEGsi46FZpaUF0sLjaTurOK4jXSOrcZWUM3FBmaP11iNb53rfMy
sxr8HEPPhIJT927d8ZH99YuTWqaLDOG4dcje5jUW02XVNGbvN2ktB3lWmfuJiRk3SClU6QT/6dA2
UDslEN3xxSaY14wB0r69pU8LK6B5/kD8/fnPyTCpsscBy6xvkK0XbfK9scEYMzS6d8IjkBdM2XXP
wjc9lWn7OkKeG1MT8Anv2rjyV7T7i1d8HRnj7ELD9QjFEcIl1WQ4q8eo7CtQzsVKDaGE0MUv+Nm6
8doq0oQKliRDRB85H+V/E16+cAKWqQPiFeqD4C5w6hQSYl6DBU38EzLfV0cLyhlSq3m8dZniAEqk
HWX7tdYwWegd/ABdFSq3UeCKT5PuhwrEkk9T8nSXY63RQiEvA3tbY9/LebyWDNlBjjPh3guIslIL
GveI6gKFLhPhT7x9T7b722QKNikW4szI5id2baywEtRSYpUZSLfNNX/V2kZzMo0SqsxImZC4aDFc
CPDTjW9d+Rqk2n8q5Ob2N/oNl7XqUjfhk6ZfZEhFW3886NZeEE4r9C92ZYgJpF9kxaTfiGMyqhNN
pljVDfey5xtCBTIFMTY22rUvUO5+CPG6+A5ygaVirna8GC/B2q9M679eIH4s9AneM6csNOQcksJQ
biE8TvbhE6u0TnAPbChRHMOeBIXjYox8+AEsUGaoHIpu4MMs5o+hnxNGN/1uLw/8lVpnBpa9x1DP
Pib4LCF/zkXJwOPzs/yP21QrFAOa0Fz+e1hCn6Zetlg4wyZICezuVJq+vAUAG8mA8AXQ5Id3yNlO
j0XEGVRY8K1KJmduiphsOo1ToT3USjNI1vV3CnyW3RRMyXlnGpM5jQpaZNjhBLfrUpaO6tuciGQ0
aUjZwf1ZtOqcEQW6uXHkO6yRpFU/sEjxfCbDyfTZeo8kFr07LTi8Jr5A4SXZ1+vYUnj23EB0PuQO
qzY5+bx7qMx+WLE/iC5ou1aC6LBPf7Xi9SBZ3E1pCnRYcgAQ0QzEbqXxyLPEekBC2zaTzfXuLg/5
9HExvL+DhmOEnocKD5iBbLcuaci/7SN2XXtgf9gyoEUB1dXFoNWhkt+BWjGicj5XtHxRNb7N2gKx
F4sn8QwoKay6getKgQkXI19clkQjUtFZy5SbvVUA1GAiR9czws+twEEZUehizB+HArqGP8+Gbms9
4ZeAtgazTrc8eRh9FqO+ots2kxwItrEQ90o7AKElmTpyXit+hOCR8c923PSXm9PmoVgq7QNCotEr
9+hSdZMjjGXHpfn4ZHXTA8VllmYNlAVNB6m4IHxHEYDGVi8UBO3urzavTq4xltsSgVjbGhQHjlbL
yFBmnPLtD8pgK0RTo5E14fiAQzaJO5iRTfE6YHLjLXOPXeBNkgso7IhOMqrikZBBc03yYsthKtJw
8G8v4M75RzWnrX1dv0netqU9uHsi7k6Zevvj4cDONs8bukrX/K/TMArlz5hS3l8pqs5d0g/VZBEc
6dUE4LIXHknqadcOqQQc3fAUNPK2/7hpgcbPV2cXBsdOcjTK5XAq1pQjE3L6/xkcGISut2JTMR7L
j9+a8Vl524ZsU/b3WwQAVg52MkXj1omCu9JdDK98Zg+Po6iq1IpL8VXiOlEa+jL8/1Vwokkso3R1
TSN+ailvNcIs2zfNjiSF3qEzVJFaZxlP1Uwp2aD0yjFAnbw2F7vs1xcyvGqNU3vATvV9lmcjk0ZA
nmFY8bxGqUlmCrRD2EWNbtsDGTTl1HnV7xQQyqxPV6NSMbC5GtRFAsGw7R5u4U/nTdEgMH7T81ad
V2lJxuIpp/4Pfr7h0Uk30tp7SHK+8p5ffzJLQPoVDpSYrDPNeAwbfAs0VWZekvRByiI2on7y+j1i
awqBesddJ89fgwLenJCjMqvI6jOUUTMGc+/J9c0XtsLZ6bXXYYLSMsPTdiUGKzfQZBBjMKbj1xnF
ywATlGeCawCKQ0Kn0k4kSseveJrg876+pFlvtf2NwuKXYz3QQKcrwffV4IUhmsEhDOCM5OHji2UC
jAbjieKLvzO4ymfNK4qhjlsjuQ8kiL8OF8tCk/gArfUPp6BbS8BLrzCW1zsjdu3xC4/ulFONBl7c
jZndtK84sUBYJkU0Ks3gIJzKNFg3BCS437v5ZkLc5y6Ia1RWeqOL6bP2FqOwSOAGjPyFfGRW3xbz
X77vFYRsb9LeXe3DKMuB6gEDJddmCUqYeHbLi3nDApmQA1WCVV8OoozGQ6uS5soQiYQYIy+b9f8T
CdD1o7FAPJew/CFRnDBrCFiumqR6hyfMNEMfixAXQJch7482akg8LBunBE2a8jaT8WhkksxTvi+w
qU91XAzHyG79fh43bZobPonQpHmeNHRch8yjwOIKunsfmEKW6RMfeNavRvvLgQUNgU+3npsRExVH
fG5Wob+xMr75kdeu2lor+D/Eu/gKU/QGMexPU43yx2Pzn2OakUFO0cQrYfgm/YygBzIlZrRdBbo9
AfIDLikAQpvNQhlxWkSaCMUX8cD11x9CcM5JRn+NGYRlwJxqvCyqfOa8rFVEWKbpji1yaW+Q0FgX
BOsKl/FkJvSzMxAgFucpAykb6iPNApif/bk+rEcWF+mlMz3FTNz1kTSmFc+9V4xR4h+pyBhlooCg
8AludQzmNxCGJi6TbR1HECPQmt+k5a9l3V9neMphpPWqtllqMmGFe+zhCtPxN5ihfNtJ747hUp8z
4PEx66P0ib32fWTVQwb3+YO1Goj4EV8lgNNsYimJAxuc8oZ6USBMPx7P8j2W9tFRA5nJ0qvqZ8Dp
VEvEv9t2mFAgs/Ym4mECYlL8YP+zPyNw2VKEdsVDSLsctFsviZxMzKxE+av/+blpRVGVy9oIpAai
MTjizXLGFtgSBgDiG3zei0LWx1lU2oBI06CUeIpIy9VDW6XNTnNRZAsVFa4FQpK+MdXIQdcPC0dr
XJj8+uUHHA3zx5PIyEI3cqdJ5sHI+UfOwvNpgVXHVbD3s21105Eqe0ahZusFedw5YGBCpRUoPd4r
sXpFBCn0Q0BMvqYAKEMxFe4csYHrJQzvphimHlMw8m5vMmCFGpPTDtf7CPuAqGLF1Aj46eRgHeAs
3rxsz9KTyVjXhoyOvb1V9KyRL2aFyFqjiFw2kQFGknIk1/4GVy5uKdTQK9ZsTu3t1Fo3FDkWBjPx
MRI0aM3cZ2iCpx45qf0WqUHD/7SosspXXvT8eJfHlmaHVrYqwFUNW4Tz3+1kN6w7Qp3BLVf4YO1c
O9O1EB89JVMHI3lFlYSkVsDuLTZvk2GXqLuBxfWCSR8VMnlw4kAln+DOiw8AEQglVqU+VB06PUj1
ZTEoGzqsXAu83I0uVe3KS85Q3IVx6urv6SKZs2ux5Zcm/XQP1SoKkdQ7EB42CXw6mRFlgE/RI3lH
ry8TI7Us93jdSQwstjdqBdbrGmr2i1kVIKUfN6Z+HZVD1gHDCUu3OkClncXVrtgPYutQJC2+Dqh+
KVK06wJF4hk4CLD75Rrb8UoI8tRiMs3xXoOg9QBKE8xVxd+VbERpldY146dB5WVqJcFtljaJn2cP
WbwZ6xKFm77QYKtpeo2KApFn0okp1QrkmREu/wM1SHuD6taaCyz3hj9HAZeSYtZC2TUhDCyeKbf7
ZuOqtyf2l7q3kC58bepEf6MmJ464qGN3JXMcEeg6QM/M2I/+86FCy3UPcd5UuI4dHbP1JOOldhj1
SgO9gVgzMhDeVubEPA6iP8MQ6BbWFUJtKAHokRdw80ijf8LGkZw2wMitrlkew3607hitrRVvgV0Z
ZCzdA4bRGfVziOEWZ3SBz/v79LDAdgN0ToZQZJq++QVy5gcfIDvcmebFwHeZz1j4r7f71IcyTf66
hthHm/znWaaAfVvPoiQWVK+DDHybNIpYnn67ssPEMikjZw67mv3ShJTbZ44VyEz6UtBHN4xFL8VI
bUGW94rk9x/DCVo2Wrc1TweZS/k8Zi1fbANpx3Yre8FXPgK2JL8/MFl/xNmCz3fUzstalsd4sbxR
OrlIy56s3htdzJlmBVX+4Vb9VgbkiP562BmQYWN1cAxJpihp85y33GuiGMISVifzznwW9dXAf6LU
hfvLjIIU8idFTvOGWDBUMIKdVtiANUdrMUowEe7OGxh33akdt4pe1HcbHRYrAPBIwCSYAHkgAdTT
Ggj1WARJy73h68oDh/34Oo98Qxr9j4zod4ODsqCWiIS9bRwyHNwEG5x6UqBz3yxZ8jghBwNY824g
wa4X4U2/pVOxK6uY5PXRSJ4F/3XrBZenH26VSVDl5A0ZIzd2DHePELQuHBIlpW0TifKj2WKTjxG9
SWk+tpiRXkENgTvMgJnNQomo4T0qq13sPcFjFftUcINDek7qCbxpHO/r7oNo4tKSl/mqTvK1o6Mx
NYGO1EnANm26MkMOpw84GcjdYN4T24dYgfI9KcJqGRnf7nlY42cSgK9vz6ippzOk3oZK8CMX9o8i
9Z3scWEW3nMrQasbFkhDEDsv5nSupncrgSziQnR/oOO4Q3SfSqngqYvX48eoNEHzRQhdJjmNK7Gs
2jnoEtU5+gnbrFxMVyvKNPvwS0TtyMnbXSP2MRWXZMR8pYRufy6WFeV0bYZs1Q3MZWotkoYhERfY
Stm92zUolsfDx16hv9HiRe134nghqp8NIha6ajJcSweaKl3OzzGn4+InjQzojp4CcG1KXye2F5Vl
8TZWqAykVX0oKkn2yLnXy6VvU3MZ4VaUajmScjxUsYA/TCbIhWSiG3VUnxc9gMsAgCBG6pijvwWW
oaxM3rm3SttMXikirtIFbxKJWFojzES0cniTXtcijE0bbFOa9TWTNYnaWrMzTr7Glus54s9mdfF6
qbIwx5WSeIk1I0vVcbyWdZllSiQgv/AMAE1I3uxy/4gzpdt39pslE6LWfTvMj39URv92STlKDypZ
Gh8GaZ2/T4mrYg5F0vLpPgHxWDTLBgGnFPykjVc2KR1vE2qP35zi+AHoBA+SP++slFcQblW5K1Gc
jLzRyRwN1KC9VJh+Bwkj1O9xU6uGJpGzLU/N6eFty2YO3X3hg2RD+CKBZzH0XyFzL/oQ7PGV9Ok8
B2U2UXfnbVMkb/Wl8SqEqEzkkABErAH4WN3NnUUcm7OAx0XI2ZKSbLVcq3PVPwOWvnXQW6t0pMrz
hqQ1CzXYm16BRiJ0hjZO+a/U/Ev2p6H8m9cLVSP/xH9CAV2XScIXUT2h8xiKldlLa01VfM+aTSuv
uRVVM4SxLuUmduqxU/5bZnviBPV8ExdIp4kqquIlFYUatp4NbiFbSd2mUzPm4iIz3qHI7RmE+R3S
uyW3pzfJvw3rfgrl6uQOUvlSh/e4nrYrO7v1WxGq5M7zGiGgYWACzUw1d7xlFvBNq8Gc7YrIIKZy
yNmtncO2YZ4SlfuiHl6mTtdT5ANXHiFLc10L+zhxHxA2bqtGkZZmAW586KSm5Pvtvrwlg9DvLFMg
vwcJzmu0G6K5Ez9Wfr47YyhydBe7R4tFxixhn2xky+I1zWXR6rBlROcEWHHU2QTgmHc4KSNBjBiM
mbHihU1FOuwdh/Sa0aCOQpaP4xoadlD8/nFEATbYRDhaGrzaol7NtguwDka49tCyh28q/gp0qETb
o5qXsWRSQ2YWw0Z4hf5lex41H0YBxNi4W2tPlsWdcOnvJzHxvdFGBr0v2aGbfy3ucQcTORJpD8kx
jSY+2yAST1u5WowxHbjDe3bYmsVBU0idzgZ7uq/Mu0D8BU4l0TUsmV6jcSyOrmvwAEg8A86Du3+i
PanUrHXz/jfNpKnLEa1LXxobpMNYYNLxhtGMHDbp9O1UyaYolRoFCIfIHPdy8XtoQjwMo5f16UAf
SOJlwqdb1Gfmeah1VuQ2vLMF8uVkpEB2wNWXbUPTcut+du1gY2fBp7shwzIJb0AK1v8BH4KCWNrF
Sm5BOq08jbhIIpvZtMiMX1XkL95Q1qG7O2RJA4Yyl/ySMGjN2+9o71BKlnEEnONoTGhEqdxPIjSE
YfbMJcSo2L/93nD0EJRL88vVBoq+bI2uHge/guZ/rFiF+sEMeJpPQW7anLnSWjGvKydeOZV2bPpz
WNN56JOOUOmzFzxKMoDBuHl6c0kDpFb/3VbL4dhrva/mLfCzPxe2EOmD9Q4L2aogvUgnaJYJwVZg
9uJJ+j7TtuyGKrVUkkzaj04goWuhkp9jncbWaPlMzfcfhZTC/CPo6SJdBdTe7TdjcamS4j8qEqzf
9AO8UUNUp4kFeUYE+JAzcGDHL0od/jkYWGdMA6yc4Njmgc/H5kPciIn5ipcOwdJizo78RJzR2VXI
PiqgUZS3ERFyqBv172R21WOOSAEJsiXSDvEM6O2aQ0L6Z+aSWppSJxkz2H7y5Nk/U8YtiogZn8++
dfUNrYFECMQZGmcXJEKz28vCcmmtEKrAZpguInCg+z4TaC8oqMbV53kLSn4e1eOONwf/G1eB/SK7
q4oiL87hZz/rfdEUGJ43CyLjjLS1UpY5I/JDILJCVJTU2JlLxRsfZvbLp+SVob+EYqYOHlBqOnjs
GeYZqH+xXmmrRBqqW6Hpb1g+E4sEkfSIdIjZTgZ+/SHO+/oB0uc8xKAXEZoij9dwswlqDme/ayzA
zDJ2/NpKfe8QgL6YMcRLshl0hxJiHmZxHwBJ2Cv8l8V213q5mxoNLcy4FHACg8D6Uctmm1eI+a3K
3mCZVzjkof5CwFO6qKu85oL6mu524EOFEfKrQdfOwNrpKT/uoc0m5m/Y8crr0SiUK4vcLIms5ZzJ
IyAPRGztfOfn5hcGHR53qTNgmhDyxT65XPwXrprifxJcHiK36DVIVFh5dtaUSi1vfunwgESyhynF
oBEeK2YNv9NKnVCjwPvAf9tiZ+9Mk86vg0YwUQSGomNy9r6k89NiJSoIQPMJB+8oJAbKbBopeAGm
nsbXVN6R9YDIcSn7haDtZtywC3Ac1qau2F3pNn2skspv79ANHJYKhPMhbnoJOLNJNR8qdgWD3AMP
yOEQy2Isb1JiLJi/lKIbZTvDXVxm3+0OxXaLT5UwPFJBSdr/AE7v7H7MMGa+Nnz51TI2HEH/G85S
uAAIEM1ydEowLf48shmMCkHs53papRUsV7ZGfJMC3GZmZANJluVYNdqp+TlTm5jBFG5dg9OD5N6o
qLjY3xLQggwwiFSyM85IXWwI9cy+9V9bCbpVCkss5yAUvFz914QbiWa6ZotaP0DKhK/Ua9jwLwrI
pc0nA1jFoHp5lgc5lf9nTCU7Wz73Du1D3lsTcBsAPTdL1yDf7IcNtbpv17JBndrcp87pgE/aJy6x
wWTaafAVhN3uRAR9WAQSoj0AgFB5tjv1YloVg1LF8um/7gHwn19Zs/5jk1qTGT3mpxm4qJ0Ne+eN
Bc9oPN8a/CXzo5bxWMP51gLMr+S8oV/NwSIUgL3Wu0D15CaTD6aL2NgfYIayjp0vPSFuQDtwCfX3
bhYHJ45xaV/cMH+QVUhnYKpK17SppfAwHf2jStb8NHl6hpxm7XxGwz+mYjppUHDOlBdBa+YZ68CZ
Bm2wcbHbhKwRoBa7BiBDGJsSK8+X5hkXYcjbVAVqN3Ioqvu7dR1EJOHsum9WokA86KAK4ueMaR0q
7Ws8y7t+ieUZ91mFl8rwpCGupTi4b9f9MbreO9O7V5HmWNyPRtzZlXqmH5NyD1hUL40H3kJPbIWp
4ONqdMdqHtIRUt/1/lGB5zk0Jj6f7zqXFxGJOjBsD31LzvFVpH2icY6KkMM1GQ2/q1ZVAn17I6tK
mtw2HxJ9XvulRpYoul5WuwhYDKCfl9OHTa3P1AHIxyNPAoW/kmi8bdsvZr9Z4zv62Wu1jVM++xfO
+dj2AlcbRtwffkICYBopCC26b4eCV0wx4sRBtGvr/cKxbxPFfw1XtAfB0Gd/STy3rbjDpM8o/vvd
GFHDPnmTSoQJl7y/1cz+a3A5Aku6ei9PyBSgcUxxU2KNl7fvxobwLjG99WaBHaugt0iLZFZNcSRM
Y+THdzPFnceu2hQSTz1ZcSf+9SArRkQOpkv8IitLqzLGdpGS57cQdxrHOTZAOTbG+9T3WgCOtLum
x1J64iit7hHBg/0toQogwuuBlgNjtTFH5N79HDuGJcNjO1a6PJpyUkrfgmLrH60LNI4aKIu+dCZX
bTalAuAt0ykBKne36FyTLuhq48aCwLODVqtvXl5UpdRvjEPo4jjvFZj2bVItHhstSlsjZNfCD4/k
dANZT6zCyXFg+o8PdU3sz0IOA6F706RV24fyYST51pUGqbJs0abWo//N8lX+rMCDL2QOG51Q9f7j
z0TU/E5P7L2z1a95INEK3iQLjheenxStlymGdZKip+0jbCljEwqhSUb84wO/Fcp21tZLYmyWcvDJ
mjt06qfYHNnz2DTar7BTw3+yNslsk0w0UK+MTKLI2XYjh2l9s0OO1ywvl2oGIfwaZeMWkbV27WeC
SavG3RgbIQnailtrlU0JaleMJWv/FPzBrXMoXougisgwVS0vjATFSDCqpII8k4nJhZIhbtXTbwXY
RNlrftQdcIH7Iaa8lEjaPf+1myXGhBchAoLRo1ZWUCtgZ0KVUbMQxicN0gunBY9wAS+6n2l84pEK
OfmrcdoBhs7xoE4hxeQWAzcfm7tO+CabHk9wiF/Da0cHuJ6Mvd+F4ngITNy0n5QclwJHjLysVjaF
z7d8gl2xViaw/uwwM9vRwgu2GZr0+KqfQgGScKjon3rTIMU0eS4VwmQhJRtN33fa9iQE/fP6q3Qr
Bpj63uVPzj2clbrGRwUYoSPGAPzl3UZjti56piIUjkuImzcY5JKNIpacFVcvDb7Sx1ivclXQpGcY
eDqG52LankELQSaz/4fdwvOENhAMrBR4q6WO5ZM0NpoH8F4BzPGPc66ZBSskVUJwLugEOy8vmXyO
R6oh5KgBCc9qQTRRfDWSEJ2GZsBoGiRb+EDsfywNTj3ruHMHo5b7ZExBdjkXx7ePQC4WhRMoLJJC
zGeMwMWN1Pzll7Lj1isR5FG++zeKVHjKb49QaikBSe68CCxghVBGf87JbCtHYlccdQoO4KDLUHyr
20qvIZTZzRZFmD4JyFq9CNCZKTmManGFadvMMSY888zQcNAl/uQ/M/BxE9Ki+tdNbzX/FM6DpZke
9OIZEC6I/oY8Vhd08a0CFGcM6IhPWX5ewoVhYTk0XjGSVZ5bHrKxejmyaHgmc7UayNxVwezEh3tC
IK42bwTRYUnlzZX0DeR5GrFvPZOs22JkRPcTeVetNoWbwsflJF7d2qHgy05Ni7NqIKhqmHF2caxX
2YEfM4kFdOqLYd60DS9GpSaopvfQEIzjUb4ekn0aIXRT1ZLHjbGIWiWjCuXL62oXJkHxImV9BllF
ZIBHw4y9agYP/dTmoFV6yfVuFPlxDfbBPK0SBHX48olH8fddbE+07Eri3T/+zdo0GmLvWrnnCigR
8kLPOYyQ4+ozcyqwiWMIrDDNJsf9d1x+DTI9hGAYYeC+IK79esyS8ondLWcygqBnhMV1gzEu6III
UGNb6ljSZuaEw3wuwjnWI2cCF3Sg+a9uKFrg8zczWeMWoK/43TS/Cci8nwgRvtP6u1SpU8imjw96
Wyary2W7IdFmNHD2F4H4Rg5Y/HjqgFSbv9sdi28L49Yu1LTtUR5p+pawj3bOrhOoXVHK2bO4F8+z
8VNCmtsTJKsg/9t0uBfxV/+lhSHebuxg0UR9rSlCJtf14vHtRVRePb9rydzN64F9MaAh/RbgFnZI
jdRn4DqmrNloMMkmuOQUDgOCIKN/jMifcIjKLopmzoZZWyH4kYHdKLJFQw/K6eHUGnbbUjXsyRGR
KPlF+7nWPp6CY+9QUp4ASr8k/riguQIXuEY+pI6csv0cv6I/b9kXgWNWugLkq0NMxb8b08PZGtz+
gKfKhBbywaSl6czk13JazMImaNi8xZYH9QblKR8mHTtB/keUtC22AE+hrsSk0J1GcbRLojahDc8D
VzbIRtJ+545Wxn4uk7/x3VI2eIdaad593PZKxA15ToylnE68g3KrJ7/NiFRwZ2vFhqef22M514hy
TBc0lS/Kcy3DbErqkMgakcQEW16nJSyjnmeK+h6YezXXGBksIYSizO62qg/1aL6vl3nEKBngqUgl
/vUOp1boYxcmCHDsR4lgvBY1Z2donAccFndHvIJUqyCkmSdVtUOX0ZvMsVSbGb9/3jG3dWjus3GS
7CrZrqHQ2Yl0cNVDyyEUfdKttV6NsjPaRQa2/lEOeoAPe2LZkX7wnxLHE9iEfqxT3roMc+x+8TDp
5qxfi5ZJA+1H0ZwRa/TePnCKU7T2/lSwPNBU2+khTNXC+eEbqVWd6RyShmujLO7xNpdJrw1tzKgk
yY93oo18RH1AsJgXJQNd9fv11NJltqJEiEHPgCyiHobREor7aSJg1n4y6uFN8orhCcJyY8KhPXL9
qzVygGzxS1JfARTGjTt9BhP3fOWE+kNplvTnf/jWldelpmW8K9wa4Tlpy7rxTTr7dqsD3NHRRiDX
wFBDj7Mj/67nmlu6GKF1k9yzLsuXCyeKYzVZh5SI+FNfhdzwPLTgRf14eZ1TFab8rcTbp1KMg5Jq
jzWShF3ntIAAXC6HlwxxK/swjLySoRmrjp72+O6cPhwqvu86h59GRUAzohWNnBk793MjA+1r03sJ
Ui0eBXrYjkKKWA5s69T/aTTrPxKeSx4VQbCNJEjDg16wQemi8jzIkynMLAFtr9o4aEw7cVhromxg
C2Ge+uDOpIeK1FSAL2fTzRuuA/IT1S7XAcRBVchI9tC56atG1vFiowNwctcf7p9fS8he8/ivnpOU
k3kmU0OdtFR40QAK3cJHA/wzbkHYAu8ivq2sISZZvX65DZlvu60xXLu3YQg75LY1Dw+J1rk/zCIQ
2S6a60u6vyXAD9/8ah1qdrunvw+zc7mD/KpDQk2xsBJ4lfDRzKafS5HYJ/4gxnAP5IMf/FkULarc
g1yexPTmYzJ/E4D2ZD2MwwI2rqNCJ7FYsKBHEiHvbCDdXNLWmjDpI/8Vn20vmNvE++PndWEJ/QKk
eis3GcMnNeu5ABbkoi/jQmH5oig1zWWeBjAo00ZlULBoBz/aQ2Iq6DT+3UoT0rMbV6aBXae7QADZ
bFxAyTSdiTw+ysobohuuqRZv+8+MG6wF3x62CiWKi5ZA48D0ktLXpPFESui1gilBVJOr6pJoF0PZ
3ws0dfaFoDoeJEKMM+NzHe1RJYHisxVwm/CmajNd+fhSyTAN+6gJdEbnLpNehzKKsaCsuBSeDlS9
Zu0xgA23fchgxujbldPbOvPtowDTrzVXP9iJBdeoFObSajF76Vxst8l/WOIcfi7GDD0dMzSkGIhr
P1HXLep1t+E8A1IwXzxGHaPmY5RH2+nvVo6mLxgRlhjnMYUKNp0Syj9YbHcoHRkxFw8NBI2wTlgq
IpG4Mnnzts+sV8hzFjsK+BrYYeNjCDs0g90OQnQpuaJ4kaaZDdwGQpzzK51Vb8pd0GtB7rk3PKsn
B32zedQ6tO9gyylM+g3tFVEuXRBKyschdYbSLASAYgck5xqsOl5wjueGs006rlB9gbzgg/wWFeNQ
jhdE96fbO8uTUgQLSI4Lm0ukOGQShp1Nu1CDXB7YEA++y4G1LSPUxlzii32JZAnqgbioE6qttH5j
da65B9yEOs1FtRRB0uMtjIBCA3Ji1aKq33vvaj7PNHpl0nJkf1DWh9B1a+Em8xLtlXJY4fhcpr42
u/+syY0Tl+HhB4QdLv6w+Qg5RGTB6sNH9O/O/zg1sPxjXLQxY1FrE87caCCS/TiDhTcdQYBVOiTQ
lNd2hX2agoyj1124GkQJ7lqV72vDxwiiu7vjHOUiT5YOsKg7Fx616pV4a2akKBlcp9jg2RZqCK/1
T9ilvTHwxFMcuikRM0/wj/CegXQt8a0h9DAoOM3tGRhRxXUdIBXDtBeBAgHU9a8G4Dlnq7Jc1PMG
m/EWIarpxUg/HjDdsQHBmNkuKXmmoO4m9E091jhkYLNi/89lqdJKJG3VVPErxQBqPH74EiNgFFWi
ZxqPiMHMs5bHvQQii3qbkjFxGuOXLJWQBKdbAP4PJ+MjS+fhQ5gJCoLDYc+DXc7ROJxN+0Rjr9j1
k8djNuPVuUFGOAIdiyZqWsFHl4RCk0/X2MR+C9mHgM6VEaRqZ+TwvRXFjz3I3/fmc4IVyQJzXR3Y
Dj1vVW9Qmn+hqQN0nurL95suguu4Ry3I4jX+nXcvTRAw4uaYC7Aw7nf11sCT74vY56nbx5h+w6tK
skvnIsQ6BPq58zo1CiUL9zAB6Lk8lQPo1iR69y1TTKMP6p3/Yd4LbvWiCWHfZE2pGI/z6WvRsaFO
x/MuKiUmf8QY0yVyZP+z/qRXmeIoA26PhMgT6tN9zn0TexpkVcTB+JZHa4f0c4i6POvM8R3l6Zcy
IhERLP+eG5IqGITtYvWUXcs5TXGkySSUkIxVtkh2uLb20GdiuCPnOjh95ZiHOBXToEiz3DxGPs3n
I7EsaPHustiU/hd497O94lvYOxuWgO5C0rewQJ01JcyBnFhh81179zB3p+nuyVRPcBMB5TRI5SgA
aUwc+ZsK0kYiMdvbnxfv2uDd7GgBOnGteN975onLnVCB1//4ujGODkWR7/JjsIFqqNADQRJXecpJ
VKuEZaESy0BFyCktwOKcZfA4QInu/Cs+EbRkK7WuU1HVz2wn20OhQTTVKPHKNKmDt2mkPL1fkv6h
pr9fb8aDqU9HaBq93RBHfWz9/9Pio7po7OaPInMJcptwmriauCsLN83+E04+W08QNYcMOgQGRBtl
0pxbklM0vDgdxhusaja9WvRlO2arXbypVBATW3jUzruLpUQjZtMUpP/GX80zpkfZHSBqujJhsTCt
ecnYWeIRrtp9ngA+2GDD2cMbGAVazRp/p2Gp3qLC56mMKS04n/kCLUU8lQQsc/LjyTHc93tBzk9o
POFgHUPlwT8a2eYQcCkYPROqJbi5vEjARTi15dxEwiP1EXgJz8+pygUVBR8FWwD1NC1YC4Aw4unD
lTSlrYGTj6Bff/dD1A7p/GA0KdaV9LKCEtC9F3QEekyohXzESuN9MceGvJH+IHwtC57nuGh/fN8t
wtxI/+B5OSDI5Z+njAhp3QQ2FHzkKjR6h8Kh29cx0EijgzgVgjEQZVfBDuqZeATCkKF+x/6gxD1X
xU6tYWngRGCCBkiiSUnIVvgK1NioW19JNZWPde5ULMU2BTVwWoEbDPoI4J2CPwlUn4D5MHaqI8JD
22TK6tNwZp7ZA9x5JzAuwZfueUzq6iX29UXWG2aSpYCQ6AKlHqfK7ARAT2uB58FkqUm81Dq7ICS+
LVwM+Fw9aBDAspPFDuPCVowYgdRAWQcRXhZVjoZ7lovydb11Ihj8pgFWYf+JQYaalrZyqnocXJGm
AwPcCFGzGW8rSFw5T3qUXYJmLgZ3+R0Q/zcA9G79KGxR8H2va6l8c5KadpXG+lovasNj4r7WQXvE
juW168A/rK52Uq1Jj9t0TtnNLojj1KcJM4GaHIA8XewgrlIzaTB+PXkCx0AB2/sbKa1cn36yobIa
kqnVnf9lbH60T/em/1R5Zv8QdHlme2USClT9UEGdtXTkD5/UhDdA0g9XP5AJmjLxkxclKzyN6O8z
izF5HaWnq6ed0AEyL7TI6xLfpFH95ry+6KCBVESXrSwggsLI3Zg3gr4/Nv34AS35Sxgw0wmX+O7C
UBS29gY1cgi5a7ylK75U41eblmIFvckxtxaKkkF+WU6vtpM4nqerAQnzFfGS6TNtHGFZKnNCh8sC
GWElEc38O/CtrfZl19i2AQkpU8K057pPnETy+DpQjrVLfpv/VPAVhf66Yz5WhlMs8wwYdlbgQZar
Ye8HkdLHlg6/6KwwgrcQ2Z/kRE3J64Zl5qU2LEqbhbRxN1+CWDJ8iA5CszfoELKDjW4+I7czzUDb
Gd/j8Tgy7Cm3hLNlpmeXq6ajiKdjqtOeTfuGdG+2kCyZgmDo994diEnL44nnw6WKQiRw6sTvIna8
XEkV5cg72Ci9AhLRefWY++MZds/IW+jddcuop4nhCNLVggGfQiZHkChvwht76wYfOC3/76tzXWmj
quoWGkYsD2PQAkCi33Dn7jcpPgp6uodnNo1h/pJs2Ofy2up34e3RlXNpd2NuGyNsAwXQMrajYqb5
nzm4fVV4mCqMjQkvnJRJw4gnAs885HnDRSXFeVLNFwbi0fCC/rCKLs3B/E2k40RsK04tykVgd3TC
vNG3e9FhJWEVx9ToCMZRNUdMPuZQXt5/ppOuTdbvCbID6EgPHQp/PVWjAtMaWSD8xiQSGqwKRDLS
WwK4aGMVYqE3iXt/zWoQe+YV11wSyIKOFIohGy35g2YR20gMS1m6SiA5t0+wsKuyeW9l7PMg9tzC
C61Lpo8Zp22yH2b2OVDp2EfToy5Bog60TnhpvuhWfZ4OwkJJRHpI1lKlggFv1mtfZt+QFiYndw+y
T5NII8PwpN87v1qEJEdXHuLsIVbLPKOoUrYTvRtRa4LGM76h3Aoz9qmojYGZFb/+S6CuMCBQW1se
/5Wfuc5UtcXX5z3+5k6mmfEK0XQm+F0usDzF4BTLYnAuSA0gGgLIVKkpUXXCrjEN7Z4IHQqDsjmN
nB1nvIC6DWmKMQ5x4p4TB+e8PZj6M5ctTX51ff/qxdSCROh2UMZRXvrvGeX7dyto/0wfIEtrelnZ
XGm/soeiLPCpWG05z0+3S3bAwpUzyI8zNu3D5HAiZza0WN+L/LzFG7KEIIM4gvO8c/ToLrgdWOHZ
Xva5FjEwafXL9nLfLW3MoYhuiD2YjftQd5rxRNqmGYs1f7WpvWfSqVfQQViijjY8K9V16td5Wzzu
jUYmla6PuzL6oON0/vOUkkfCAAbsd7YLC9lk6kW8ZFtBEKl5pctWbu1EHzpYCmmQ431gfSmEovxo
FXWJ1kP4hp2DPz8nH18d5HWyGse6RcCOUQavF6SzQgld1nwLVvRj4p2mtPI2hjDsyMdUAO7M3iU6
MNaDlmEFj7kV82Vb1IBPoseMQiSftkbR2gzUvGZeI0F3DcQOj+wGnDtVnYC5wO74WNp2/34YIVfM
N91fkZtXYVIcVWCFe6PZA40ewarwur1411sExTqYejHE8JqFQm5JKJ6Hc2Ms38kRCYpTSuknX3RC
axd+3J2etwMbEIzv5oT9qT815pKacjJ90vNCopXJyf8ks9U91QCuZ3Vqf1BABQ09/V26ffppQHbK
tHYCE9hcOOGiyJx0Z/3i0YzDohnlHH4vRrKvgMG5e4Ugwig5TgrKSHfOl3Chv+Gk8ao5WNczmCW8
OH7DJDIjHcCbKSZfrGuNP65YqJ65K2Z1/5AgM4dvr87twUvPWyXoYYzrE8PtxPfFEQee4Rd8xRMk
DuUutodjjog6rlfV1vDeIE0Gci8MYnaFfStoPyH0VW6l5bt0iPXvk5TS9qlCFa9jYG4ZXrCz3zJ0
QlFqUEMVPGYZi4rREX8oowdMp70JhL3jLW8PcVDO+45TV1lEVA94ee908M3IVvb4fGqO+32d7rUE
Gr9h3R5tvD15B2sX3maruGDNO5V5BYup+474Sb5FNygH16fL2Ylb/HhuOHmHC0YXdP9ApRqx955E
SbSRBykc8Ut3kL33pXkJjjpLEt+K1Rn9l8KZxGcu/wtuVOIbHtz3pST2iwzxYey1XXmEL+DcKW/0
04njLKGu291CrNY9m1KWhofcSbX4v5u4qXkvvDxTAaIDvoqA5ZXua9TIMuX7t/Ie04whvXAHLEQf
uigBmyO3jag3UYFCjicvrqteV+fftn6WRbBGQaw2KlTSY+vQf8THAPNUAVsdkU/Zc3Ko5NMLv3/M
9xG7hJJlXyjlQdnLgLwenAYVgeZVmCWrNqqRBVx9SMbe8Brk4g4KC0nEp2zdCCLEu7gtZAbCdTTr
wNJYhU7xMKT18MZzshR8siblUb5TYCREfliCfyMa5ewYQGASIPsJsy5vn0ow6p1l4T2o3hro2v+n
xeRw56miCgEQFEvCoO72INJEntqDrC1dLiGo2z+SgSvhXJrTCnT9b5E1T7U9iE+l29vraziz6Bl2
+btfF4+thB5i4+tGzO1ZLO+DqpIJkHXQMVRGeLq8XYy+co+dA3pEep6R0t8DqpVU3iYMy2PPMjNM
25xu3kW5rHfW16SOS3Fkr9FG5ziSu76v6M5S9VRAulvmD14/1H+b2WlqewRZWG4RIss86nBUJS2Q
ZpGCoCm7BjGJpBmxBWvfCboLJG0OhEwwGp3xLnXl+fpavMU/V8vW4tqH5ejG6M0VbQ6l8hWSK+Ev
FRKmZbqTvmFbec4wLx4q07FNUVL7DmtyL+sqlQvO6qKb2ftl/J9O9Bo/77zJvKRYPb4BDyqlZWkZ
4/+L5FVHHNGd0QgDflb4S+H031H10DMUarTlkbtvVnZbZqukZvIAgSBoU5QWqgiaWM1cWySfVRdo
OFwpvQb9F+a28R/E0Wmgj5uSLa4ISke1fpylPbN1wtBMfJpCpyULWrXClF5NEmMj5ySohv6Xdhpm
Ep1m5cQGEd2afu37F+vv4JXyRw9PXq9ZV/K/C3FS9krWqNbN9vGwgpzYRwt5Vh0dAPc3WXhNkt75
TAYWxZU/MQ1jVti0Vr4MVraly6b1JHesUxWZ+KHxv7kMsK/tLQgEv5yHg3ViJEobA40NDvE6faGq
WzMTerbXxTBAr1C7AI5lhaCA7ZDBzXnrnS4m3/536sQDYfaWOUXZ5lxz8lt5UMbpSpAWNpuT5+IG
cc2P4MynyiVxOkDptGaLxm3HaWNxhAq7u6NUlIqsQxiqtS5kOzNJkyxjX7wEIYhLnsiuSA2uUD1P
vD93RCzTsH7AjxRLS2f8cYrLniaUGSW8ZToc1BD1j0DSfbOKOC3wDQw9HYgYH7VZbgKXanMd/FqF
5q7uCIqyzG0uO0o//gWdl6BHOeS7tvf+WRSBf3xJdvJ8SzPdEr7bA8LzqxZfxVulsmsoOkJ/KNRc
C249rxoG0PWJSTdh3li/e4gbmdtk33uRot1wJg/XUaCjEQOltMJUa4H5IjLkKX9KRg53aqP2KZfj
ZKVolbvHr2UXeg+r5YyAgf39a5HlpCXuT7pa4KHHqypEnP1XEk1RLdC3za6NQDmoxV/Vh+yUJli9
TY/kuVsuZuyTieJZyj99NGELpABYKN+DMhox+bir/WOlP/1AQjrPaUT6s52aPvD7Qx10oqGpPz6t
f1IjEQ7vW6z8y5mHbsPfpmtkb5WAxGgMKdc4XfGnXyj/XfVjZi53Los8uG+bBS4H1vzQ/IoZ0PAO
f8W6iQJPGySvwLmKg7HBkOzXg2X+pU1rxgK3ccW2IK6nSGVW6jgJ0tge3is1MPlwcQIGImQG98+j
yrMxg2AykRy1e2kk8Z1UiMX9iQdsSMRCgpKucWDm8UUX8j2WeViq9u8/Q2N9dVCX1wCIDt1Ks5sq
3VvFnGSKnKgv2VRW6ASdWWrbLrzUvsNYblk4zWMmsyxjxHiJgeqi2uvuU3wRUAN1Hn8aB5MIdcqa
QDLtpSHeaqklOuXsYP+0o4J+sojE44AZ2tEYbWVf5PPP7K92rv24KzSqgglpPPXTnDk/JCW56yO2
Fx6cx5UA0VJ4YdHyv1l5ejC9+8/SBTA7xqUl9LpFdw3Ofi7nXya6g+euFV4NVqehOvt5xNL4DStr
qITPlCWprJQ5EPEsvsbuN4g3noVMdHsaL95bM0+i3p7Y/RNL/jGJpp12uhwaU4DzeTDKhmwxwg4X
F9Ipl6e/DDmEnDgcPHNMBYYWmrS1zzNna/m+8TWBcIyBeer9hkHIbnBxN55Tvqr+pHS5e4rzHjb7
Q50oujG5kzDkGWn7XcLSekLglAE134So63YBjHYSKTFJtvftm8GXWKXzmWXqZ3gkMsDnSfwtBGVE
c8iSZodFrf7mvJ56GKzY5sAyWWPwH6UodM0wR08zSAauLhJdIKnfynSB2OzNxyfmnLgCgZXO9FA7
nDDLx7b4hfeLRtFifwR5RvloMwb2cTIxArTp5tP3qElJjOpb3hxbfTSOa9vQKAREuiWQsRyA9qv5
CCXDakwAyFff43eao5Pd3yN3blh/5WkR0CrAZyCl9DnXpzwcVY+EtNLoG8t9E6fB6W/Q5JB0EPJl
oXYuLnsMIuGBAqnx/HPXHNmeo0gNZapHVo5Bm4+k21SWSGX3tb0o1C/+rov52lcf6TPmsHwJUR/y
F1FqyOGs5LIwAMLT9m7eJi1BYn6XJ8nKH9cH/+u21EPepzMWnfSzHLXrZp1gfKhtDNDXhPxct1IE
iulFkCorGhc8QKa35GTTySiIQ7F9hCW5+aLPaly2dZNSl581qduv3KxCeYsh2m1+bzIi0tg5Mmwd
4yz9h5Fu9xz0uTh098qwI4qnfgi/0WGNZOxYtnWBpiB/Ac2KjfTbnxlGtv60fqDa1bbwFGDafvqJ
IxkiQK0HBkRaWt9nFTH40spBZW1tsqAhgHpYZZDwqMobokkvuTJlbIFfZ4BOXYZvo14baqZoZOks
LkQYsXszFAvcWPtieVqFF/PYmJvTNdgPF9Q7Zz95erPFq2j6jvQzW12EQLDFmEqG/GgC3/u37dTY
c1vSdAvg0yBYRb9IJjNr4IPyJRUVkhPwIC6qODUIlQBB64zGvIlV+h/FSr/dE0m0WJdo2wghuq6j
+cOV6jYJ49nXUuRB+VzEAesIFe6JMQGPzgjkPVfvSoRVcixl7Ezd5Yql6hgFGqOvYG+YmyviEysL
tBfuCqCVJBFLDPkXQgetD7G4Urzqy+YE0jf8dyFxfB147jPbbiniV3rKHrXZ02Kfp+cCGhdj2QlZ
mLwK7JALFGxl03e7C0eHA/Qmob+O5ZMRuEJDMr4Su4H390gQVqG0JEXcMaWjMYfKIv5cdb4/k7/j
nI99mj3Kn+MNjPTS63JKOldr/Bdpc5saq0TY4k8E/5WtTOxcKvCZhABnIYMX9A9SSajhLPwM2Zwe
PpieYHysdbyZl9jmuXrkjcQDxFcZjSx/yKwOp1Bf512jQ+haAAw4X61RcGpGBpE/9Fe9X7BorhN2
I5DklhuAMrX6E8DW2IY9NSdDaRzKrfRjGBGe2Ss16dnQx4P/l946t/yoaz/iTXupxbhPGMnWETyl
HdARr4VLvuOACB+O4wqKC5NafeynwKYv50gMQ6AjeR8tFUT+IDqyZD9Saag2mc9Jg213GXhuooTL
JyjI+f8C/awFdSQsqqr1hoaX5VlRx1bytdvbzhk7p6eUusG3SnVWTBkU2Jj/DJaI6JcMzvF3vur3
T/m10DzAx2UMfyRbaCz58VJhy5pkdf5qzTpXIYLdeTzmYkgdijDA+K8pbCuOO/NOdTg9QhGQTQS7
62cJ+gLj0626nY9vsdoc4JnUVCRIoeWYs5WdTPvSwd0beOw4b90Kw8zKPjz/Ju3ga6qw+8MfF12P
/VrGWudXNWof3Bwra2s8E6IjLlO7nTeeKmAE9Qo7qwm3WyZs+/KLwkgmHe9JispuJBznWgrv9XKf
dDwfvsSRTWz35Tg4d+zDbCq+IBOa3SkcvlZvr4yy+rsm9LOU3VRLeELn2ppSdIgyOu0l1r0QkSu4
AdafbVOl5x4DOvZU/kzpgg3SSKXhPsb96JosyfwaCyz4RzMiEBRpDNn3rxJPflqxYsTDLk28o5gF
nIGnesV2y/BRkI6Ai8OsWc2+8Uv6lNufJa6ZmXHsNHev8MCCPY8hcjHLpkqpigpqNMsF1Mh2t3u9
yS4Zy4inDzvam8+v1bPh2VhYrk5Xmr2NYCzKpMKMv60TtQi67ILE8g0MjAxd/GPIS9NMRfPJnOdX
Np1QPLlGARXhLrjIdkasK2zS2B5LuMw9pv1j3zwy3/3fKy5k8ebAuN7sdsmt2cGERMTgeWCl3pjI
B1BWU5qsoplUn5O2YGOoIiRGDyhQk5483ylTi5JNuAPunV06+MB0HC5CfRTDkkUp5dnl3J5szME6
HCvtNZ7nOQ47JYXzW9VYxp/OCoJM33+ZXzwm0C11xZba8U2SWm/s1FNesmJPAlEWgn9vVwoOKR8l
Hlqz3wJhSzOpxon5KJV2+fyObd5tLTMGDMfEdzHmG4w3BlVbjMoWuerIT4Mf5YZhsZSv/o8GyiHA
8bN2kVWWQWIJUL/c9LtxZdhIFYYJu8wH/RxFVhjg3c+bxAIoubCcVapbzUFCECiaF/KP4MvxNbmn
VbDXkP0F6lRU43yjAv5ph+BL4ePmKlWVYqGGFaksq3LWcCghOsntFfKAEc0Uzu7ZgmrtimiOPSHy
24y6Z78uGaw0zFDuSlPYE1pQwbiZhmQR+TmN0+dbVgISBssQyfHCZ9U46jsO/vhBI4zqaKP/DiSC
BsDqX86e4CD9CK8QtiqxUP2Lcr3KJpTKRPFZJAdbpJ0z3hJ5qyP35pzOkg1Xzv8J43WC0quYD/9o
SNtCUw9v9RyAOPcgloi6FEVdE6zknepk6kmpKxlcP+OC/4Po4ci2ssl1YuczRtmPqsTSZ85eef/V
VE+UDg4o5E8+qQBJgW427Ltto9SMJjZM4fgphnEW26k6ufESJ0tS9MXTC6k+EtHhiIADRPEHClR+
W0tLA09J5xXiyaeoyAybadFSs/f1HYFrrFfjHga8rB0Cq7rm8iAT9yC44ggK6tRPwafXuS4BNix6
55qBZFsPFJdNqzqIG9M5h5gDhOX2kbycsbAnd7GV6FL/sB1o6TdY+H1U7Bu2fBkf+d/LIuNMVst2
NCjXWH6M/6QaAQDJUF7rYpxOc0kKrbqK476Zaqzb8onfYtEEiapd7Rgn81kD6yacLxDOYMxDK2o6
HOC4xpUy8kwwcnFB0QB1Ewuk9jvl8YKsBThNY7bo7Df2wznDl1Hi+wiwmo9dunNJPTf6X7OnNa8P
sfxx+2CFOeM8hK4uoPUQsRHtGg7UIa0AWSeqqE5/jcA8jkjBrpDzMJyaIIhjKfFZt+Rtj81y5WIy
ZrLMJvIZuxGw693R2g8OXQjUl1e3EY4IFxQiXnvnngRODYT0Yx3cBut+jJrqLiBjjFWqmBJxvoGv
WqTNBhaeT+L9DWwdORmAFqzMcSys8kDZbSyjLsAn/u1x5K5ajzIaKQWLzGaBqHAfq5QZEd0+TvSy
NF0pF+chOiwhQN0KUoOm592xuzdST3OnmPj+I2djdp5bCa/D3sd80nv4Uw9ML+UwuRPlwe22Tz+x
/pBrBSj8gBxvbT5A4D3HYvYdEK1ewthpJ3xTEsV1CZ5b7coQ6Jk5G1xgvyc2YPBwIDFqLmkrr0FU
1xSFoawGr0CVABNppv5H7Ntzx3L7NGa5qCr/bpMEbDmiQSdC7OSdkQIPAwHfjpenhzqdALBXaHhV
/MWKNdxds1uqaCZwbapJL33gJDXOYJtsMhfeS4LsP4Mvv9hgfh8qXjFMzWLrhhvM2uJVKFnAyGxs
DjEKFmkBzd7sm6ybLrY1mCOjIUiXf+m+ke5j8n/T/NErjnxxJRLmQgqXU0UXYbo7iGXNfixgtB+i
gqtoO5FToCNzPRZl3Qet7TM4nzfULsbeCSAJBROywMbAEhdaxQwPQElP2wjZQQomuni0JM4LpgcR
bjwfsMDjKELUxFLBQwj+5HQ5MZKmXpAif4Q3FMXQcMxlOdMWHaGdPlQj3mdaa3QCHe7YWNiI8bX3
9F+kq+YuStUxZOQOobAIVgZs/VYoF2f1Og1lSZsSt4Zi7PzibY48Gu6of2DKZFZ1zdGyJIHfw3p3
5hPMSi1xkSlDRgjWlX5yOlBrQlblGk7DvizJ/f8CrbLTk9WAZ+mD9xU3tZX8naJA5Q/SUyMRujBS
p4kF/l8HoKNckDMOfQctEZ2Zq5qsm16BEgdGjOZF0+fLWBQBCc+MxSDDaenncDbAjHiEoJPD4u+B
gfxEpISZk2o0Oqb0p92okhILpwVj4SE1NjFFQoNqkko8IBJbuDOxNMl8w4cuxnfeFapXTU8vrNfQ
Oof2cy25InDjyuNXM58j+1EQEEoDft3OQx8fYuFVjwkwSFT6M/dPqKL10oT6hltCeL8ZGAFJRRmw
7w7AkkLZuqs86gYqS503BFtFDRR6dirFRPMTbi8Bk0NSC1o5FSfZ5TNa1+h/rNMSMqgrNPuVft81
5VXvERk7z+uv5yP6SFUSDwCgdc1CZGDWDANtH4XSuPRB9xwzzrBBdfVfUuidiz7INYr/0YRjVhhE
K0m9NB5aJUFJICGadU/8BCEWh2UILeVPX19a31aKuHbby8yESGYkYh4TJiKnyXobh0YDUNiK76mJ
N6micK/n1sfNbYPDphPV71G6emiJ0L5C8Xdm+Y0EbLGhSE3bAMfJ1LjAyZ4BEE6mgMguLz0jrrfQ
+Z0xyrRJtgJdk8TN+ovYZdcv1v4f2JmxHAE0yfSHoGCxzIJiucilj/e4g+E0Jz38bGmoiKHAsVCJ
xOtkp7BRsCt2pDSgayJKGVBFu9p/a56bbwAj23xLDnEns4zYU/hoM217UOfbcrtKFUHWW2wDNIMw
CUvc1YiPtytMO9EgdPkhPa4d9RsfULnAoZU487291+bdeTe6CA20XsVDUPxWlUgDUW81/HFrM1Kv
PehBdDBxufcLcjfv+8jPY2kV4POlvuAL+bzKnrdRKbRcCohllNaNAj+yHmINzPLyEjC3FXcsBRy9
Puh3Dyto7ekttAauwoyt2PEMh6bm74z9Cbb9abbA4A4iOCRp//PcUCgvFk4xJPNwPmO3cNYPJ3yX
V22O3nLjCPL4Ft4fiSBlsUW0IK7jTW2SsxZpOtVkOlltXA7+3ufp5yDaf5Onwy65oWC8aNjZ78/i
ezotkh6BRn/QNNawnwHR9FZwsZHHsxtUouRavHB/B4S98btFXHlzWdGNtYgiXQ9sF0a1AN/7azGY
lahSMwBKPOzws0Efvy8Kv5BwkgsODWwuKOiyHKbPA5AzQIRVr6TyaluHu491eB3OzSgvI3yWeUvk
cMY65pBcUxHhtWARV0XRJmRE/rDjolaVvCsLbDUQUV01AkFs+XOcLMZC5JY6AagRFP8yTTb1vZU+
s6WNTDn8UZtjTTtjnM4NiGLgXpKlU3UfQkNnqmwBZDcYc0R/PYpugPXBHtbSeazL6IcBIr+gV7Eu
RMNPUtV+oWDaYTLWS51A8dY9MjU8G3iDcev3vHzsP93lLZFs9ariWkH0NTL9UKJzkl91emrfOXyg
F7M+5xCYzeD1xThd6jdOf7ANx6L6VR4rtdPuETuQguiiSrmBcinZbj6gP8ncc3HIaQZ500SvS0Zg
mCTM76VDUwNxRNIohtIU/AmqbGf6nynKyBnFSNS71pqTk1/94X/C5sJbULJAsgmMaIt2/iA1UJXI
ndt86WsuW68II62+TtXQZT3uQtWx5TgAyIK6VrwprRf1rYEdv4o1SoBZk6uNyy2MtFKFJ9MV8fQ3
bq7gKyxs8VeyUAIw0hbSL616TMdmMYnMZ1yMCvGUgifaVykQahg3kp6z/CMcQOFuhUUde3SRyUZ3
PyY6YIWJ+ZIY/ACzngXrUTAK8QXAHnI7kt20pG1q7KkIoz4KUqBEUBZRB3t531WdKV73gg+sRwh1
r+sMnuVFA0MCNA3990Vb63CJ+PnliBCfhPe+wj2+FyuIa7Iz/VpUS54YcRjHjGcAS0OOJ3JN5Cyn
RyIL52hs+egydoL/nM28Celkok+sx0NJiRC9wUED+JEiU9Xp/TSAefI17mDVWxsGsq2fGJuQntNx
0uOXhmrvrfSGW64zhovnJAsnlF/Jbg8g3vhOc1heGQQNHIjCI8SHGmOTENw0QhstlGLwn75QPuwH
6YVnSby6lw2QM/kXr0Y6n9K2v5ttK/cpRgr2rvCHzQNGpN9ZBuX22G1ztTyKRIqDIqUJKE00VbV0
bOftJ4O0N1Cm449kD0C10SN3y1sJAl4EaFim/23n35RcFpry1oPk+dMZkUvZhodDJnvoDfHmq61N
/4FjTNyy5hnCWofeaXmBzKF0YMJPMYOH7LTymMZwnk+jzfHpFMp/dCB6Bu/62lmJ0JPsBs/7ZGOv
1PK8tuR3dEDGAZnFNzV0w/La7Dah4ZWtU07UtrG7L3I3oRpAraM7INccVw2NfFzrsuFd+WiYu6TL
cWNBKB0W+/f8noOV2AuKWT/P6EJIVupkN1oz6zscRBX+buz9ImYJ5RrPYuHTf6hm51KuE4luyYe0
FbipeJTD1NNpEdJWr9O//48VjZQ5asqte+rAczeKSndh25l2nOvqm/379aCOAKbs7OdgWfE38Khm
ZkUZYNk8gAJHGBe1EMclZPWpUdHvZqPgu3PxKsYb/fnGH0XbuRHl0PUMnThkUeaYMhjK5sz6sFPd
KrGRSjw3knXcGKY3Lu2veWANsicU5bm/HDvvV0vC9j5K64QejnknLZrrA9owGJCoBLM55NJxslfd
swAuPiK+bphPmQ1Pua8uAFGuA6lZwbIFyt8CrawY5nb7NJJlT1CXYINcA4jJPXXmKtCGgFEzNRrj
5Qf0RWp8Wz0+s9Zs8Ps2ARFEhBCl5hJIZfuevvGuGBu076ulD7LcWgQiPW+9/OhvvM6O25gA4s1o
OGanh+lxLxkeHjUhCqnM4kH+I5e1HKiJi2DR2yce7JUEtdAx65o38aHL6y52VW+fKRepmFmKr+t9
cPDmhOLfW/ztcfdRITBSx6WiXNOMe0q33Fmc4K/JVbgYuzJQVXVmAM8sBP3r/B9/wrOafeAVAzOH
OXwv49/C3ITBtwzUw4RnW1go9R0gMt1HlbVIJEekSJ2VglzaIcSABzQ41wPuSl9E0k1/2SG4taUe
BMqjDoLMk6aXGIZDIqLV0kI+NakOyDcRHG8wDysbiL/p1KrDW/4j8pdfVAF81KLHFFxx4yg65VLS
UyUuZ5MI5c0Zk8C4pcEEfWCiqC1em259PsdDPoPUe5tbUD/XQZDkeNU/G8Ved0zeX5CiDXMt0H5a
OeSjWJQr0e/G5MO+pukB4wo0BLxwWL5y2ZBWNw1fK1wXFhpGU0RAA4i3KRLaZbO3mVs5dT2OGb5N
8n0OPiqyImu2nD658NhawoaFamHYqYO4DYh+LSDwRTUxKndU3Uovv027c4JqHLCcIufal1rC9irh
CT4w0xy6h81aQTAm4SVc9MPJII2S0H72O8PpXhtTJucafvckwbMnftKcgQh+ywaBdZqGgKllGEud
JB7xlM04oTb3buKOZiC6XhHrpDcCjL/bO1URwGu54GOuorQoktgYNvKEKTbs+KsNRIH/J4Qd5/l+
ApZRKo5tfit3T5fRychYDaPe30SBxrYxZDFpZXhxMuIX76wnKQ448He4as0lyLbKrcJxCDVWlur1
KLmawKxcmnhxwmFcJSeNMd5qOEipeui7xvFZGMDDULNMVLxsIwzvmvw3NvbR2N1dBHTScRKnAtfi
DXQIzRdpS7omWnACuC0cAxvKvoBIn1HNMAEFkJ0x10BcDcKPT//8PN9VBQHLZGnvAV7f4goRLBR5
DjxCm4W3for4UNmVK7cPpgGNm9pNtMHXG/xRiBR7bZbqpC7ca0JaRLju2dzS2l0nqVt1WB0s0Di6
Xzuexk2rbuXiIMoxjGGc0VEIpJsF01Dr0QanRyMIBEhS9VuNTOO7wxSzfwD7VUsV05Uuiks3rlCW
Q9CF07E/yT5exTbdAUl50TkM4p3J+lRmO+H1yc3A2bfkPHK/CpO7/JVD2hHe8rSWog7E42c4PWov
lKc/DfQ4LlGotmAC8b4luJmqAQ9my4hgpfV9mP1xEcXsTKubk+kptFnsueZO3icvQNtmi8dNcBxu
mbmMvt5PBSMQ+fVoxMSOS95lLxXQ4LoOa0IqM7hS2GxPeiFXULu/IZMf5hYqq1dPvvndjjjWaUdn
/MrBKj79AOwN/f7lLDSlbONme6AyL/UonI3OfX6SxPcvI8Qg8NIn5J0vqQK5FZk/FYiEW4xmvzgv
yI8/XTuDk0KeSL5KXw8uX36ZKlPfUabv/RyyUK0tJ6m8fPuETE/a7qrxCTXOk4eJgDZuJsqK4/vu
OYiPSD/91qnyGnvlUkmgiLaP8CYii3oOVCUVuCAZxaiMm6ZnoJxrAgYUpO/6f9W2M6TlnnMmZbx9
Amc93aWf8P3lLgQt3f+HvNdYfgA2aRMNFBhXwGdp5nxHJ+N68OMsQrFTulF5PUkgtG4GBGtLfe/H
MWWB5znNPUd/RDaetLW4lVhfOZ1S9Otmn8ilbjRrV4iF+IyuY0i8hWgLLwNMx4X7rf0Vr8KKaHmU
ojX4s5SZD/j2pRUBRl3L3hXlxopgNB3L8B4PXrwEcXUSxjIltmVoS1b1AoMoKuH/wILLJV/4Wp0+
JNXu3cSOxVkKQcJh/JJLVEvQkNKxm9UX6eO1GI7B0/XYMPWR4jor718NvyiC0bKw5ojRdKQVUs18
qY+xyn6+VTEUBQ6A9wgP+e+9oSV8VkKo2VfQRd1wwNR4UN5Z5qKjCwn/Gfykz5m1tefVFucO7Sjm
2OP810uoHiGMoKdp8rO7CZRfq0TcRc0Mnq+VXsK3CHVz/l9/PGuF3oAXrEMdSWUljBdhswONAUxp
tfTOnEb2nPdCww4fVxLZmGQPJKiHrLvSBj/kJdsGK6s+7StSQ7sJwaMkGJQRyw8Bm52wZb9nQymq
5ROZOFaiRV9mRaWrw+GAO/0Xh/keZBwZQcH4EMpGhsbRUvC6f5/LT1Fz5bhCKpp+0/dMr300HlUK
zTiSUAiglWmAPj4AST3QKqwvynx2b6aRHycPmphf+fXmlzC+zHtfMobGxxMuUyuO8I4qVyRGGDQO
YUVct2omZQ6vBa4bppmZ12eUtt5szHP0DuO0Z37bxqqqzKoy502W1YG7+JpYZt5XYDbcbELA5V0H
NMI3B8hj+wXQZXA4/ZDwL4dfJg2Jmlya8jjDvXqgNe5ciU+9uYBQ2V9beHpP/aVLkDHO4XYEGnhT
UUA5YFDEIY70Kh1FDXm4Q9FYDo9HYMuhc+r2LiuyxuGbwCXFQoVfBu1cfAuUyKOsZgHyZd+QE+Ab
pvQXe6fY2AROJblESjhscdXXn26qWn/E9iO61DY18rpm718orNs1/r6tIk6KOgbFJqnKt6BlDNNX
VF3c4T6KTqAUzzAdmBmuVxM3TQ/YKPiFZAd2acxSDCNiFgnTyHTvyDMX0vXYZgS2sTZuuoXR3/dk
edYJOfqZXvuGGszBn3MgA8VO3yHRwDnkEV0qWFXvTviLP802DxCF+mm6g7waTEhI+8zpT+cYAfoZ
epCR8+L508cQIVfiH+dYlmkUmOr1gZMfcM+iwyPNECZ33I2S6orgmARnj2jhFuTOPaAyvJ5dP6V/
v04tvMzkDzwXAPg26j4zUU5D6AHvnnePq1SqOV7c3aCTkSz+QFnTIvwoWalZTUqsZo51y+cSkuTq
Wr9R08cR+tHD74jRUxsCVY3d7g0Dr/4WdVGgNdS3PH0d8Xf81/76p0mfF/gcTmZpOocY7rcdFr4N
5VMAJIHia/Co4P7Kmir3USp6zhF4MRENzeoMZWe5ab7DwmTLp9RSFTIUUfR9RcKT9USNdZyszRNw
4/Re5c9PMo9w6T7InKDaE9rZulJyoFLnortox9ceKV/2wgkLSuNj6y2BHDGabLqlqqIp6GwdgB3n
U6II8qra3+bkTvncrVY+Qv3dMMoihl+brpVXYJdeKanvXNJ6CnKyIOq39U3g/j3MBjWbSo1u0CK2
90hdPz7pRoqYy7iFcvPxII8uc9wGrAMMk7TydlN56RssTHH5UqsP2o+JUF+RKg1MCR9t/7Jnu/Zx
PCBM3GpwaMB+65EAgKVNJpt40D0oK67flrgdj0/DX37MZ/nkzR2fwNHn0EPwHL/kG4UlgIL6vazO
C8+WlLGSVTV9txlw1mzsibpgVu8FXQBDOBZE5e4afIG9QYr0mJQjjRSKybgw/E2HjMXhRcA7ErdS
kjr0JDYe/krftlQCU8ORJ0ZDwjkU7c8tcqEicCFyctjjPoGzc6AJDmpRRWFCvLw8tkz3yivQoUWy
I/e9UqBlGcT0qTRAQt+Q9VWME/xY5eNNPcIZOUYXn0cufkhuOOaA9h9gbKckGWBF+75BAIp3EaSv
UeA/9/wEV4LvGJo/3Rzq8yBg+aF8WXbaGeJwFpMlhZHiLGHNDLmZUs6n/+LTNEzqY56fOZ+RjTUI
XR/zZ1NJ4JCLJyXswAL+jtUgOsDcefMAX8DFgb6Jr1pwRrqRp5RJlYTyZJ8lrYqCxr408sWMxq2u
IsCbd/3DBsIRyA2wXjGSNQ4M0O/nmOzyVzlEmEci0DbzRGzTaHFWr15D0mlwWwq6jadRviFAjUta
WNkX/INtLl+oeIi1KH7qNjwVK7rUmZbPrZRh4LlH/d7xny0IhpF9oJNHsOYAAA2YPyI5iW6T93n+
iKAyqaVw3IV82GoQkPZi2Rm+t6aPgRkzFMpFFPpMnnxQX/x19CUTehHpjcdvV8x2bqxEAbDfkxTt
rXlvWuY+7M432V/UIoLitifvUxpE27MUBgIa3ZZdgKr0K+PXLTJZ3hPLJWoIVAKtjJ9go9DkPA8Z
Dr0aRmnIcpkY2pFWjIa/bSOYyhmZLOEGmndkZVPt+1zHm6OCPTW6VELbuZjgt5OtgWzfI2C1LFvG
6w5R+PsutxTbWfbz5O1yzDKm1WF0Rn2LWbfI/4bp1IFXpOTJAk0WLfLB5nJxXH5L0LSzKDEfuCpC
WcTT9n8LakiVl4bw772bDqpnmZ6cwS+hdt8DKV+Z7cZ4yhm0mOmVS+p+IVr9ZcN3u6dEIXeX6hC8
zeYTK6HXuYP4ZqsNTg5bmb44BJ5OvAHfCwFJiqq8iOIwSYEmYpLl6dqGvZlg2/dPfgMT0Ii357JA
/pZdLgCUDs5LP0v95V4NzEyi2AJ29kERrkEx1KuLkOyenH9IODqlRDWxg4zN0CkKVdlxRM3r6Jhq
2+l0RaT+ut8wCxC4YhV7J9nQJ87ZZcV0gFpdDC7ZmKFay9J9giU/EynnRzhfuK8P6OLdvMtjhLyL
8XxQf4MMONvnrOcf6vY8xgssFGZPB6/o6BWWFdRaGyUVsX9GDq5g3uo0F9f39IC5v3NwzNPAB3U/
bysgjXEctvlzySo81Y/kSaEgcqE3dyO8YZmf/9/QwTLwaQe36rlxMWBwos0AfFsnFr3lT3tiBrWt
c0miALVOJY/izKzwN3WAXu4s8OFzTcgCuwJ4Z9+Jxo5omjcrx6zInNx8v1v5gC/8zWm8U/z0S0wo
kUm+PqKBxUZdEcnkuUg/pRNxZTDDgKxzsnOfNcm5NnSJrnIBWMBfEhgKiX2YG+CX+2QcAuw2JjE9
w1ASp7nuzjoMR0qMBclF7v6MEs2MtzaAgzJW4QCrhJOsjWntQ/fSBDScEx8qPh7irZ3oBbKP/X2F
JEaHm9Z+2xBnt09mq3wuBuk4AefrwsNwiKSXkH7hisc93cpOiyFd660PH3VApsMRzW7rZ+YCh8K3
ItZ41Lopcwq3t22xJmalI1L5RA2eneP/l3nLGWeT0uzbTlXKuK3L2ar0+9zQMUX3YR1dbm4UohAs
pVyrYVyMqQ9Gm0to+S5jbhh80mzjgdMhn0gn8FBDWWI4i2Cmw1LgZqillcdZodYkS5IpHWrT9Uge
vnownVd1DitSm87t0s8t9v1t96lilBHRivFfYo/pI2BqOxWDRDCDNTED7OcflUDMZLXGBuLBH+aE
3/ViMzIh6yQKNpdyXZxx49e0EOvzFGa348En/JQIAaMVozsLoZa46sTLZOS4GjYEez4Bw53RAwDN
zH3KhBQPzxPpme92vc5m+GvVKXeZPm6rCJ670lzHCDamEoJ6I5tzB+Xoxt0fiX7cg2Y7h+tyrFeW
AUHnEGSQy2AsSsfM/xOJmsf7fYJQ7zahHS9/fBu3m6w4Bknue2OP0nWxsnQtlALEAkb+XIu2QhvH
sKJz98ucV6IrPKDB3MN/mJJRsbl4iqvk+L+LAZi206BEicVngHefEh21tFOJ3J5BQzEYkvoGyhuK
KvNwH2mKTTrR0pF2EtwoYTDxK6hpA1SGUdtlyb0iVS/OnNAvHtflBtfFWGwY45JPRgrAWBSh/dcI
s2cdzm4bXhUOmxwupDMDcI3RHfGas5KUWEtXgHQyrXbXEHPRgqA1vo0m2IB5PTeYri6iiWpS6KWx
TEAYmUMDdFJZ5Sb6vVhAwL5u2YGlUvHcVIdszla3cJi0zF6CdX+RuvanZa+sKvLafov8H1MzDOuR
eFTHpGLcXHE2sDIuOVqdJjWwrIiH/6W9cVRoE8yiuyaKCxybb+s9hg8HQ7fe5aMEZPCIJdLcXkDP
KnRoFAsX35Fhw1oJv24imRR5BtFlW63Z9MyyicplpVjCNOAUR2XsDhZMs6zQzEqIV3wXM7vcj8//
RbLZqaql+SKewP3xAJTaj3HgiN5W+nfJc1hDob/AIP2ttSTYk7ZwfqDHVVxAyUjKIo+ANqiWV9cb
a//8UNSd0dRI37aHo9540xaID8gCPYwO2kU434KGajnnpFwmQLLrnvGvxKgdAcDdw7k2hVQQ6MKn
aO6rXSLKQWb5ZWNTH65+YuwW1uhOgUQon7gFzDO3y5tDYPxq+iENtKGS0PpuOorTxQ25LJLZURps
dhvHqioApGWo/Jsl52xkiec0onkO+z6PUdHTXbiri2efFwucyEgl7jAmbdJ1Apa5M2cyAZ9NSA0S
bT+TfCchm4Qxb0KCTK0f7l0GwNlQAN26l/QD3Mdc8hM23GOu09wKHgWjlpYVEJH79yWZ8psdSFiL
n0krmIrFz+JeomeXVCy2dhBPHlk+Q5W6rfnxKMH6VHoDT6CdqpMvu6xFUJ0GpbjwrgbVbcHg8ouB
3OVoB8z9UNhQn3tG9qNyy37AiSMYPrXYaL1K5m5pdHMKWxP9SD36XfegsF3XbProZeZ6h+MvtTg3
HWoAVnpUVZKnynkCMKsq+7k17PBHbQHFDuJOneZZ1PV1ZBV6avCDrWj+5qKLEVzygPpLUbyd95Jp
bXgMYXJ6m+/GBGBsVJ1gBBGSUM5ZyO0ibPqHIMX6K32QA1j9T9aHQIG0a2jxTHJIjXDiQUN4v4UQ
rkrbc0d/0KKHn1mhF43pWmphbaD83N30btroPucTfhiRty5wqON3lQiTPFFm98Eq8U9DRLbu1nLF
pH3gv/UmvXji7oADuMPykh63v386PdAR+EURqnsUHXes/mHMlOamv3iUqfNZvKklIhK5EEe7tCsE
iTGn7pvU+n3g8/QE4P0K3f1aRDIhv9BGsUdQSR+Uji9JMt97AeahpkP0gFtCwNQ7aplFW7Revt+N
C8Qroq97nvU7OF20WcaYbTDqo/q771Y7T9ecFlZAX2Eq9m828YlS46D4h5UbQSdi+Cu0gfzUUN4I
OjZogMDAk9+YZdUP+/dUv1BUPC62OJFP3fMV+ZqSNIZieHAtwnxPthDwfbY/ZxtjmxmrU/1e96ha
2gkFp9Y/+75lerYvnSEHcJlQJpBmyCXw1xBXtevq12PK2qSV7y7VY8j4TIDpnkNuTTkxXa9RfawP
LxayD/FHf4ch1Xz+Mpwj7nEzEO/ELT+zwdiE6hgI2wFgOkZgC2XWRbGHQwcIGjR/7icJ1sRtEG1m
3i+ZLTjSoJRJP6hZCTPEdTnM0v5B4SPJ/tGaWJ23IjDEr1k92cJOMQiVEiLFIEDh/BW+jbV9V6qY
FC6LvOi6kf4fi3Fl580N+8RHpt0XqRajdmELJnZ6LyRGTF0zk7SiOgi4aIPElx6KIVKUlxMsur7l
7TjfMGecJDUUsil9kWQw9mg2jFFn65B2AnNRon3SMCaGrUu1mra/gO+2hI5eyq+Jflet1GZsZRv7
zVpGbpCobn1kA0hqgxtWgNH6GthmE99vFjv6dOa9JX2tBCwlIssiMgc3FdNmQySnap1xppuHk+d1
T3Q+3pTA1QC4ZZV88LyZ6kb8Q4OR86XTfFebYBG09oCwPLn0aKwzYSV//mBwLb2u9Yef0dXGpPqq
PHqUm5eSbt1HSaX6eHvXbMVtC85AuIPvqgB/AHBaUgzQsJmeJ79aryoXd3S0dWOEro15GVdpRoGA
n5kaSf51L2DIonEBx89Qn5B4zHHRKMPIFRiL8oXIG14CLG9FPKJPy1VkzN9Xani2FaKajYZgcJ5e
L2eVjfPa0YMK/QbywacqykaCFFwqP/ZjtXIqJIbupWiROBYfBY+qKUWpzF9pawf/Z85G28jGnwUp
qj/6XYOm0nquDfr1YxUkRLJP86hK8iR1WDzr4z7frcW74wVhEa6MPFFb6UCeLg6ROJxtXuniq1Nl
gkSR5dOxVKeRZEKL6O+6OzlxD4dJqeD7SJKu9+Q1F8SE/0AqHmZYIyMnaxXkbI/R7H9P4mDv601d
ZcuxuWgzGVOMNl6vSu2thZv0zgT99m+6Q+Z+p3oIm5iW5R9/HX3WcxPhseu7ERl7/KwvajjIhpFp
n+Zu4J3zWmoeOiwc25q+HRDQmQjvVvuRHDGefCope/gU5gAaBVVAKPM8f+cC8zn2+lyoBSDY+/cC
xkAQXnuxOf4LDHhr2b/NNY/kYCZh2ceWZnuONlKLk4Sov3ZGG7Z+L42HSPMCy8FKb3qcZw7i+fsW
FpLJ+z/FfNc3zWVLPu5vLqNOnyoS7bSuwrLB2NlnM8GdnCZKF7zB2WJeYf5Gip5aXu/8UhbvJi78
9ygzxbgHh5Bf8OQkYweGxwN6fLd9PSQemqZW/Knuj0zH5koRgR1z97Y+wPVHxBsltADWwiiIG7mY
4dx4LebpKA6bWtaMbUvkW4zZ8ZcgPM1709GvhECOinKUZNvihSVtaJ3lEMBrKU9jrkcXt+pSKz2G
b1VpSSpOVSA8QE/zThGYypFo4pJR/kBeCoa3krozQoipWwA6id4F8pjNkyA6YYeokc0+L4rqtJO9
znqhWfK3QruIiljetXF0Has5C8huTd0czxeuci9TEtxK6Lmrmu1eTIiFKcJva5gJ4RT8QrIEVwQC
3CTWNPAQQblNSQ9RSWf5AnGL8ObFkcRRETUN02JJ5Z9ViNXyH4bAGWS9bRkMU++YobOr80gneUVo
a6G1h8MNk60dcttipjZXIljRdIyi10yIRUNQO3K6GGHqgI2fb72/RcAcuJWlrybCtKKXQD6ESae8
VvrSo5FMJDB1vZ8VUh66U+9elkWMjzwLGgX5RwNjgNJ1M0aSVKFoKa9eMx6zYRSbxstCftreY2c1
ctTg+qZC0MoY67Pryiisb888yHUg5Q2dWVA9yHgpTedUGJxzwudqOc9AONQJcDNT2HHW23DpmSig
I+qw649z16ZXOmj13dkSg/Gz72Chqbh5AuBeO0DX1aJMMhYbJOnS3yhQQ+4RQ7DOZfJ8+CWgUst5
UjT1mChhYfvSW6SQwptBPJRFLYdcwdYq5l6DwE0rns28CiEvWlp7iguUrlbciOkuyAP2vEHchfdP
iVQYKiWmvPsXkisjPFL+pt1zUov4yrKCeWWrqoYQxrUhdwiPB/niXiKCfWOzqls6lnp3LAQw0jUH
w8GDi2kzTiDjEEqDFvqcwtZ6MJXwQUQJgE4QXZZCbjMyfJrcOrDaQX8RRP0Pg/EcEFoBOFfOK8uG
pr9sxLWl3RUE0fVbuOhtfv0UrTyLK1kXWt4OYX4tQw+dEFQJZrI7HxlxlF/C6JkhfDAMb14OHZH1
zE+pry1uU6Dk84i7xAszBKooRwPvvFE+YSrl3FuvSQjU+c8923ggypVZt5QxFAhNk5NtXnK+QE6E
z/SYsI+v1wBD+qVGQoKzkJfVHBfhWJD2IYnB8OMM9Lc6uuwUxKTJpY4JOh/wZ0+kBJThf437eaxr
Wt7M1kEkYpMgn6kOJe+dfxO/6mzuPjleHqgNbCdBtUqtAs1xWyLHJ8GGKRKgZjAHtUooJC16Bg5j
RJ648lmRvG7Qa1yf3T166+PCvw0VHEjIMMKD9frd+za8FB7YjCWUIDvxorZfGeCW6iQ9Y6fuzvbe
7xcGFDzioYWd4NuxWh7epeiuaU5BkDstjudYSZA9mzoRrSNalYmFMzjGpYT37zn+gdpGlMqmDM+x
1d7hr3q6jBtmos3sIVO5rYbqAaDyC5jlZjPbdJqBkW/m7o3ob0PBZ8vkIpEz37/XWmGwq9K1KvLh
kaacSFR0InFiIsloLaTL8K4jLBjR273cdJX2ycv9T5O0fCd6K7nnFphWxh7ehp4CZ8iqRCaSTt6d
TdwQ2mmzldN6geWCgSpQl+/6C8FCGhxv8r8wcX2AvLUpKa4GrpRqNBzmxkTCQZBV9Lp95XS/ERfO
J5EGtlly71vPkbdy4krooxGuvSfPbN61nEVzFDo5y/qvx8ikn8XyOwZLq29LivHWNFuNYa3bJk2t
2WpOz3ejpu2bIGTrEX/3WE8RQwD1CjWZ0m+FWp5BLLKhHlTmBZVBzjzIFsQF448hwGB4ykvEi347
+n87sUDRla5SDoCWKvsA37laUqMTaloHTE9ACzxfJ4wRQyceU+LQG3Mryi6J+uPhdm2PVCqefp4R
WFoHpAUZqUCVM25EJ0yKuEBTNTe6LYA/Ci4F1WsZEedGXywRH4x+OnKh97VzyzecXamiSYZvonsr
2+4tC4+Cz9t5xfgkQ8SA5oyoVh/Mduz3kuXgktlRZ5Ei3G4kmrK4jxcQVnE7Wv6P6iEhZHy5c9lh
SZ0QZbV3NEf7AifBe7XX4yazunNl1tmiWXtBlRqJRHgVE2E6/nE9ZxRO+PBYBOat750jzdXnz4EM
2aHUyC/O8vVR0ILNf0248xcWSS2Y8OxKjGi2M5exkZ/V7PC+S4d222b4tCV22qa+BOLklPuHjY0x
vZDPtvsnrKbzL2tLYbJf3xHbrSQaBw8637SjFydgc5i6RpgoTF2AV3NrUdNVrR7eqaj099P9sQgv
1iAifIcuPFuV09AbyWnosa1Rtvrhslh6AnoEH3YcWD8a9Kf7ncGUWDDhvLhgx7p9yEy8Uo4DSPjM
XhAJgwwlKXvGLWPflvR+vRWKXe+MrflYXBRXzrUQTk1ZclOBLPBrhFdNHaeRDX+Qz8PduRTQUk6M
m5SsKjoFEREYbW4XiEy5rAjc0DcAfsc15Go6vDwy9cuuC3JjxaAVm6cNCovQFw54VZNup5rObhsg
Qsb1fC0kENet9fqgwf3+gHaGFfmiNZbzba8YvE13CC6WGamjYqZy6dXHUj9WnDc8CCgSaj8/tGsk
hHYOwio5KFYCRnIqmqlMd9Rjuqst0YU59if5munrprqfzTd25C5s91mJq8gYPS4JkhTqiWUAk3fN
5N2h7YenWN3y0RJsIMDd6IX+uylu8Fhx+Cgt0sWAE27aFtwp4Jj7oVd331880IJzhPMaXpSfuq4P
4kx4+xS02WAICs41ErHRavMbIBD/hHbXv3UdsKAJZyw794obNru1D1d8Lp70rC53yKYtyngaarWB
b0xSAL6EvuzNsnWzNcoh2/HKxWZRjOLNZZWgBNyzS63Ako9Ahp+6DwF9ALoc2tbWkQ7+fhf8lQeo
Oc2Nb0BM1bDBsDPGR3cKazFrGcWeKW6u8K47MkLmCWeh9aQDn3jMqX2XVAXjqb9KFccuiOXLGLOR
9M9pF9TgF8P2FZF9gTF+Y0LmfMi4ISfedt+agb6MoyaChXRv6VxK0qCMrkJ6oAfrj8PpOheCyHn7
WgFkOk70HXtr6pz73Ngaclbkqsh1XhtDfVXp/6eYdIZveZo1dEgJe5/lt6EQi18zHDnvMcRKqiwg
/XcDXIZi7Xli9meT6K9v1ZO5lsD6om3Zaomcsg9eFtpvyehdCDUu+Z1ORnHG4y9AIk1SiBzhc9uL
NeiZAHV9abUZ+W7SOlI3qVKoQeGW0AoI8YB/ki9jfEJJvkuRGILtQRtrbPFawNrivePl2h7UNnX1
fWWiWn/0SbMJM9PhBdzbbMuynodXsIQXxylnlyb6upPtuN1XRcVep1+htjL0+pqph1nXfe53mQ+V
x/7Xl6ISJzrSkQEtpCg4AHdFNhizDW8hYTqZeWnoFTOg23bFxmR77Y9CjtIYaIlr9MYrMQL6+4lq
dW+6GaOcv/Tm1rY5zYWrPRTr1iXDKXfumia2zOSgv9ju5mjmkdEgWdOXs6m6s9LxnDjs61NXmJez
8XoZIovyU+vzem/dklJqNGJFzofENLjEwDsIgWUcDpGGmiYxJAn6XXAl13ddNhERP3wfYppS9usE
aArvrYpgqHfm3VK18hSaJ4InTKczG+I0XRoq0mix9GdRLRk0Ecs7bqDRYOVLIed+QGABUghMR6A/
1TSCJwcwsp44vqSSl0yErnnEaeS3vBpVZQRfKyGpt4AU+0OH5xbQx0nXghgIsepBKu3uvL7LoywY
Jf4o3Q6Kb2EmYiHaU7joYmn7IsiZnorYtVV+BSmE3y1T1CIqQEEh284/bafq8WdHz/FT7pvDqlQc
A9Gm7E5z/FWYe9LIHbuYECbu8VFdl6l99XpUvr1w/TEWP3lG1zDjsjmtoYl0n38gT4F/uWAAYAfu
Av4J2xO5FIfeC90wGCXLltIVcSzNlSfzQjxHdGNccrmxddTOpjroekUOq4ADYmblB7CRDlXq8aPg
Mhz4ph1+Kk8GvP1vFwpMb2vb5Lvj+wy4QIH7BpgTK65a1zT3nQrDTDcLJ9j9a3vPGT3ATSa21Thi
ulOO7O44L92FJPAjemscAwBVCNkuPkhHmM5WFg7RDQ9tC+anbGxEeUED2dHvsH+zKcz1kqszRQTR
Lgv2c8Nw8iVyxCL0G77q2Oxt7BUlUCvXxesXuj2IIZK4tFfTD5GFuNVrtwqGVQTrTPQ4xgLvOBRt
WAYSx0vAxQV9XIWgUybGmRhoR5ZhJiW7KDO80/y4xKViYm7ecEAa71aW0dRf6KbmeS8oOm1+SulR
tbD1dQ5TFkjXGOzcMpb1vXBfP6mTSv0ghcWUSvmUwdSplEH4f2jRzFvwaLbYiLDmPrRrCyn0ReZk
tRfs3eXH1qYr++bODw6Xm8r4mXOitsVkyLgh/8uk/dD74Rl5wu/t/KlEJg4PzIuAz3lp1A4PHSIp
1+Xsse6XNN7vZTPdWiWOcPToBVzb2CueJIjEZWZB25VlvRGxygPzd0KWDv6dq+6IdTNr6qsyQrDh
6eXk5NzaHn3Sm94noHJlpzz7NqFPG/2vuCm56bBMOGPYbBryYlqyqBQ6vlF1QH4L4xon2UUHVBQD
3L9YEMszhjYJQVbBuQ7BXN1ykJAEEC5cw8oSjFxmRG843utCnf4lEmwPpvo7nypoSagrej1I15+H
eGnd+KI37aGGcA1G6OqIzo6LuVysboU/VJZJ5LXY2aKi07SOW9XsDoLa80BGqz57rzZ9Fc2FI01b
FHhnY4cnG+gYDor3bpCn2XIfeLbLx8nTqWLkjLjZ02nxTp2N/qiSr8kOx6pZeOMD8DpZcRAL0cjl
bR0wCaKW5X96qbdYeqNL/U/7HNsBZKehFsAN7W2wIYP/VNHaLbXvn+LliXOGQxaK90qSbxiQzzG/
cYnY/TE/W5M76/5/8BY/CWifPMXznVMU6L/CaHRe2/P6mnP76R8kjZ9HT3qcnaZW1vV/qirtfXUn
VBfDz8C3tG0P1gevcGz4ORjro5kYhRRQNbBxI0wKUht1c0rSzqQGLw3f88Fde6MkU8D4l/yNBgj/
DYuuN3FMAa0rssx8PuHySgPOnZhwe1G/JDRjACosdMSPdhh881bNbysljfwor91ZI6MncoISBbCQ
WGHzj0onINnApnOt3zEO/uCicYm33HBc+XR5n2k46c+FDJSmbb1NbuqAey3AB+uCZ7MdS+cjsGgR
BdGPBWZ4DnVIwKXGHeKga/uqSC64Y17VsMxLMnUq7mLnpVRuTllRt+fmuYbhQ4ng3vJ0v0JiR+zB
CY24ldbSpYEl2PjRpuCmqqdv2ZC6I01aEadWHcP/w4lPBCygebP/nIiQurZaw28ILNhkcTSThHfJ
Xp0y0yWFmCM8Q/3197D4B+HtvBRHawGNQ9HpFOvSnkryc1eoxvJq0ozMrnATvL89nw8jX4iz0K2o
Ok6ABTDMvwQxvpLn18RF3rxg2XulFFzN6i9HGMPhCfTBCEd4p8hhDd7GmldizJJgdgo+5Od9WYQA
z70UclPaIyBNtdvwUxNTv3kfaa5m0HcyJTWzp61XWS4J+387k4OxnCkCmGVFyiwVYH5qkTjoSUgd
DrUjwNA+qkMr87KdBQPUIHIzEJ2Fddx5Jnw0auD9RDwDBqfmAvHyzcxMpBdNaK/slCnSlmr3aCmE
MNkFKxa9ZslQi/eFGiHdOHfoWk4OiandKWoN/61i4SYlQHWgcOXhTkxF1DN6EWQRHCZ4wpEB1AtO
hZLqMO6B+FHGKIDtEuvGHfF46kmPaRP+oU+wM8lKZI45zJTXh3qgx2onsCKEp7eC1jBNHinuZOg6
hFyC4u8a/yyalscad65TVmkJcXaH6JvKpzql/OVqtjfE7csZEHM9ADvXG+p9ji6UeNbJLSrCHYDl
F+iTZMvgN3Tzewtpb8+57KWlWp+Ytntvrbj6cTMUVnkw57FJaxtPsagpwGSybvqgHh9bpirTOZvZ
RR9XBl86BtwHlgPq7vxyW0bxlCPka6DS2LOpoTRFU1MnlWtj5mPT6CYW0nSPbXbgM/bzPNcHU0i8
0fZFiaK7u13FGWwuDDaifwbi/KsIX+fS/36+fnInkxdFmemlobMeV+j7FiGoN6gitcGsAtrwQCnp
X42WItByBDPWLrz9tC5WNw24SQKc9i4eXgz6uUoeAQTxlBmYWE33I4mwIpNVhbY0N6WT1rHguyFv
2Z3SIO2JwQlGYAwvRaR/pAw0QUFKGmkFubbcIX0dVFcOdOXS50rb3yXnUv62HO/CkhuWsOl71XUg
nvLZKZAzDKxM5cTnRTw9oIYMqPYypALXZJVu0OKE1fm0wFtWzcXiHxFjw3yInI1t/I2NR+xMX8px
EiqAZ/PpsDZXtXpTep4OkTuEhudM6Mk5fxE86q+BNoyGyFtagH5oPv+rtVs4FRzRIeSgar7DIocK
vHR3yucjN49/bKTkHL0KRB0F02/zuDOqkF6MArIrnP65xfmU5aUKmHQ2JIdL/Qi/gms96uqCDmlI
eoYpgotxZq7sgR7G2VuU7eGt/7H9TJgHeT+ShfVIWxwl/Zys7VRHLAya0fMKH9k540dyjFkYz2hX
s5U0w9LsO09blQqBfHYs7yMkwNZ55UGDZ6BX7G6ae8cEnzMPcaVU6PAn/Q4oHgWCnEQGGyHIYhbT
zvE9N5j+YDwQKcGO/u1rqCCYLYsk4MGwP6Aen3ioW4ygOtmLM6FaRZOE/ZbFz6sMA1ZJohfg5dEF
8zbO4yBPihMDsD+/aQJ4Dovw6eZN6TltLdw5LXunsWxBwgcDMNU2ywNSOnlPmwbxgR3vJ/sujcdx
Qek5rH7mp4bvz/EfoWFF+3zM0k9z12uMdzRigXTxxxUbfAZHGAg0lz1iINHvP8+cvzQxSWF34IZG
LyGLwtiGFYzZjroHi3+wXHsCspTr0gbTWg4kgi4o/2JZ9ihc3pP83+Tshf5G+9p03slo1o6SHscQ
FDdqkiA3DcBhEsa6YWfWsIuGGPwHDsuWnMXX4AQM3RFEyASB2lUZNNu6pM2Zwuvd0MSai8/wC2eX
IS2iDKp7wWKpxrIK5Vg+ZWTSX9kK8Ol0iDxxmvURYMU/bRvJn/V8Lq5S4UycsurUwcE8dlVvuUW6
ieldBB9BAoi5ozkEDz3xZWHA98dcDGfs70K0QKNN+VnXjfwyNEpNgIZ+cTtWwu/FMon0Usus/JkQ
DCF6fVTDRHm1YHXCKix7Bs9b1YWCvquox4NaMwuVc8bv4eA+MrU6XTRzXxSAe1xNwE8zJRx4CWmh
rZgTfP3tkysSdbXgp+8mAWE3+99F/bVYDAyAyonoCjdMwtjz3ptxjrpWFaBUYqN34ihcJiguou5V
vkKSwYsfoQy+hrPreuH3i+IjOmuJvkZfFEssyGkijKuP8EPk2w70C1uCX/nRbNXaIv5fCeMxcksB
OjgOfSq01QZNI9W5b8/Dr9nq6TpEDYE+lOdWBqv7Geh2VunkB1ZDSou003JuwVEAumMXrkqA2MV/
elk6e9oyT5SJRZMUcmLLh6nX1BL4QIxsCQgcFAkd++BVddxM/8AzedmOCRL4jbkkCtM0Ohi5veUm
cUHfHc2/ptxWWjVySMTpTRiWkZep9jyzuPPkMeDHLdJYV0Sxip+r+13WscwztTdQLwewd0CXZ+8V
EXbFEpzwZl8UwQ24EzE6Y6eUsX5seUcmQvrn9GfbNiPFoJawrIv1Y56vJ8XiT/66pUSWkXA1FAad
SZS2EBIpFVYP0n36I1Gl6vT6lie6IB5MncAgCazNNycs8TwWgS709r/Gg73TY3rq+GYifFrQwoLj
Fp6l9QT5na7XIsf0ZSPSHQo3odWHKlwD4J/tQa6icPZzsM/DB+dQKb8/yG0WsF9/pQx6YuQsUeg3
3lkRMJFC1UCkkR5Chw4477hRGpM7R2W/s8+YLIUPDjQS2R0hJxCkA0fUeZBAN+0YPUcuP6JyFcOn
2fallhObcBDxSAxBJprKIeVaHsHN0ESlkrtKghSAVUKi12q/9GmYt/JsAp551T9fCX8AfVIwIi6D
RASW2ByTw4YAAhv2FGNYp5LQi7dxZoQv1Ovmd35s9nSVnzO2PLNOs+iGY65aEhieVNLYtE9bnTJK
EypNpX+u1g3XEM1rZfxc7dmm6kr5lHY/dypeoiYv6sGiluu8GitZVXdhu9JwMMFTrLaKVA8U4j8b
1HVD2LiMnadvZ2eoEDVxacMrckbAqPVD8Tpjox8yLoj9iGRinj45pNyhjdDSRVpszZQY9UCT/aYV
Gr5TGMc8YD+oQjKwO9frk6wSbYEFKYM1zKioxJlti5tOMTpYTEJCe9dqDFXEHTObaYntuMLnfi+U
TqeDfY9FjLgOSNPHTXowWz5j/m+mNAUKnhsfQGcIf9TsZoV+i1SFLd7xVQIEESsTQLQgrxRQg4mW
ZpdPAjIm2IkeoyxUKVpF7Fz85QXmt0Rb/uh8UOcZbvh+WKzW6FmFWBXJYFPrUND00A57xoR2EmHD
Uz1Rl+EFWyJFmN8XH2SdtYwiB/8c6TI4x2Zg/+dLEZ7Q5j3qB8/WKehgLSqttMTVKtykNsq/hFU+
eGkBxQnbU7yS4pxsKBaiu9/nMFRjgoDbKsZVR55RKvUmAITg4GhUagf8ta6opYZDCvGudn9c0BnX
SkH4eUgygEgCqrRZ9xAPBj0Rp+GSItJQnl3ERe/Ky24k6CRaxCoL2F+boiJl5HSuWpHBRE2G4rcZ
SJVe8rHuddeMQjk6eQZgYP6csm0ciDf2B7+023GtxUV1lsBnkgMlcAEQzsxqiunJpglwvXGD42RT
caY3D7Tx+V1FaZTKXUJUGZ3VAEuULvIjNcy1DpPTBQWutlYTJPipJUGYlPA61nIPZR/1JqZ2uElX
hu6ecOOWyrB6k42Gko7NqUFOGeob5JhhMNct+HhEvhEAbrOfcr9DS2R4qAItMq2KDa1pRi60yiPo
dAszoDtIVvIcQYkHGEZ8crQKzM221VqYl1KeoMSHRD0U3OkCjKdWzUMuNuqOqijRaqzvjWTzkvvC
tOLZN2UpW+g7GuEMZpnEsfm8mqwX9p/S+Un8pg9TqGj7HjgVlZH+Xl6gT4Qd2qBHhe2LNM4FY3IS
7x1fQchajSZSPYE99s2MxN1Vke52qwNPwZoPKaTHBs11BmVIwC27LBUdwUbuBZbQIdoIHrj2ibq5
xuRs/1oZI5btphRf2uVXdUh4bavQXuMohUw3+B/OpR5NN2C4kDiszf3e4rvW0mtIguO4e6fSJlyg
KMHQ3xoXLCWMWYQOD9kRETLK1cXA2JhX10QwzC8AGY9C9JgWvc5nQ7FVdPf+XXqGURODwcyuZ6Mx
8/Nc4YZFHCbZvCUCKhEd5Lh8CgjSoUnh1LjE/WpgnY9kimewUx/JUnl8a59D6/XYKucu1y88Vnzt
3v2kcRwhk4ApIbVgwwNH68UFoT3vP05vUNon2ky0pPfAlZI1rURPWdoq46z7VwovhGkswJkwEwl3
dgEZ+Z+AZEHB2TKiT/1YobH4GCb4QNvmaOCsBnNQJHCZfcm4UJxq7iQwjTjkm2XnfMrv3H6M6X2P
04urkU8s7LprEHMDlu98AN9sqOx3CE6kQfxolQWbdvugsqgI10MKFssyAr+E01XuzWskSMU29jXU
FxZe0XTDsUki3fm9e4lzf9TUP4lC69ZLCQmE9Hd0lDcWQNMwzpjDyuUBdYTGzFbLSEM5cquWfuWj
c05+h+7N5tavx1jFu4i4IWVhDs2w4Uir88Uk9AvZVAZIXEcx7wuQB4IUrjmAO0jKMMEvZZeHCbHa
zWbG6kN6ZPPPcHuWMpd09VYLTWh+rAkk2KJAbP8ndEv8VhW0HyzNP1E8CCk/uCGmSLS2VGUQBglh
OpDF7kTrd01papFQTlk0mNK1wp0Tr5wlFrX35LCwxwP2dC37KJqZPDxrHeEkBL311KZPMRBUB4UV
r6ZuN0dkS4SaoJaGdgLJZSoXtWir5YzfM6fN/Sw20XU6FKBM/JPEQseUrptMeDDoZwgS4DrvH1yh
EBE4KsUJPusDcW3U+GDOikdY75vBxn4kZCn//00Hc0ImM1RLmr5AUpjvKT/OhQjyIFhokBoHdeui
f+aXDYlTw7fSkNvNDYGvlKZ0Ke/ZSksZMhm7b2Ceoqzr/VpNyjhIBgdU1zktoEaASiqrQ6suno5I
w/6AtKZHDl2MhBNymQFmfJQtCrTyutk7rR3Cg8LjC8D2P9GLmjWpTLxJY2VxxsBel3PH4UD9QWeF
VaEpagUYMpbZt60chPwhv/ezTEqUoEkLB+5K5x2TQcZFbMMdGSs95DoQA6FoG0YXPcIHxGbs6/9s
MOcsIe9qcgJfF6FB8WObEHaYHKGoAUoq/ob8JbRK/6zj6tCtwXKV2ADWgCXn8ssYvY8olOpYmdV/
UoB+WY+04I5+nGzy8Oq8lufW9fV0oXTVaBEoHyWO9IHohcOgsDOWMLNL1lodRbcixJDL4AvyUU0P
1nUs+mLb3no8XXrKToAzp8QMfF8h9MlG1GL32bBak+nntRHAOLgPENbr//lPI74ocNvNL2eaQT/H
JO+VyvMCyUWuSCFZOxUItcKF8GB2waXqOXht3m9L8RK5lrBo+jkoe9Ql/NaSq1H5fgD79rdR3Cai
xcRb3AmfLwqvUVfeY1VGDwWMVHGnJD86KYSASvQsB1nnZ06eueSkgr6jop3Ql0R1nnSyvwduRAuQ
blZVQZvXLPREGeMGwtDsiNK0KolljJL8ivuusnNbIf74wtuSXsGFGr7kooe4DigTKtvoB2qQL0NN
Hv0S3SLtgjVhoLxbmP7X9VfizScjRBNjDFZ9Q88xSlmSefEKWmACwh9OpMNjhqIDgcufafPXujX2
t7VhFwB3MdC5Ekj/VY7F4mv3qWrI+InZ/gnYZoPwzGvyiZrqNkNgs0XjIM5Ez5Jou3624LYRI9zU
D5VZw3+cPIcdS9y2imiLWKL74H9R+bwWo0owdkoBelxT2atO4UkJtr33qQt6KNxHoD9zJj1nZhhO
BHuDFlOQ/B752bD4pLgOi5z8SbLY6nCuNOf4PpeTQWxvdRd6FhmM61GFdsbizd0zavdhB0eS3xpB
2EgE/4ELs4bxrjKrhyVm408pm0zVQvh01i9SL/gvgkohcxr0zHnw7o3O2TEX4F89BGp8F/s3q1t2
HVS/Dqpq9qXZoPhO6UoQxF2rQuwTnG31/rLD+sXmku4UpioBHJp03wVcMn2s9RC2QIXi49YoAdnQ
g75v6omhU81jg3PMVaJ7unU+ORUhcr7YeLiZ5JOuv/FSfww85T4lGvB1GxrOeVvM/04hOVultRWB
OFX5810M0cdsu8PviRJlfr6LX9YbwWrgTwm5Rw/4zH70oTVMC1eXokzM0I7fsl4sOMdRPgAf8MRu
p1ZbxOo/WZc03+N4NSnNtOCoIkCmMSml/QhD90tsj4zE8MPft4BER55PCvjza6LqIRFxT/isu/vW
tcY7R2fXLpnU9w/CrpRP4+Bqj4jBR27Io12UlBdzhCRGNylMj8LMWZSS6WILVQrInekwgtG/DwIh
/Jn8I7Xrdmuf7NqZz8G0nGNSauCLuibYkd4Sd+jjMgq/zr5LuPeYw95Avajq3Zwxuw43wKYds1i+
qxrE2QU/CuIkNykrKecALUjYFkrJwC1QgyEQ7OkYb66dlCvIcj6XUThElGOVPJorMRaFSo522iRe
r7BSsQLITV+uiRq9MObS8aOcPgu4pe3N9j29BN/gcrwNravbzTwBCB4f7WHayWZtihcxxuskgVrK
IS9xdsXvoKQ3mMDDc8PvA+ddwo/voOZeZtRYmYbGSBuFqLAIwzECDsmUkAxg/aLZ7OTMPj9mkac6
NaQIZLVz7sw2ag5xkUGjxis/yiVbMXlqtWsg0bZ2UefeSVR5oiYHXfAEzHkLnuAWwe4LDaY3wgoy
tQ0e4913FZmYsIGWE3XK+uS/mEZvtSWpibEM3QwNfmT4LkZSsAakPdb7o8B0gl4FhYmMX3//CmCk
bojjBGwUH3MS5NaeG19S7PaTx4APGIPJbvBGvT6eqBMdfC1NWyYnAfc0DO3g26awxa6HF/5S3WxE
h4vVAmK/WDVn00cBRXiIo9Uoe/fgaBWqe6KgNflCMxeA4/rEySyTtZMia+6BIgzaGR4jMEj7XBk+
DzK/54WMoiZQJelduxBbhnzxx8bvTvuZinmA9Axsm5oSmXN/Mj4zb+qON13wYsoxUkpDt2hCTCF2
Oq+2FQ5oGIZiZa7CDxo6cGQ8kmgGZM6yz9lMzkag62tLhcV9aHEtYAp5R36skrYoAYJ8nbi3ReSx
AN+JMMQ0dGZAOfkefsLrZcG/94o1/WjndjL/mHDp2e7rRVtxUaVlBpO1kWLX+HBoaKxOd4baUw63
bKY7wW1rH5piP3yr8QXkee+iuRUgOiSSj6O2VTvM/XpsoI2Iv46WB8gcdLypGiF4QLfRxDQD0Q/W
hCZjw9uPdWXuKe7c1dO/uMBqokcr/aAMtpjLrEWiasFB7saKwnO/1+jphogXrkN2pJtYuAHmq8qI
v54b4KvMK3SdsG+cD7EhE1SCNW54S9vWxZglmawdMBCj5zrhwIXhWMBOrrPm+Cky86o5Lt+jXnsY
9M7QTamQI0aYmSIZ+O3MJl3CN4e6MfGXu/kpqtQIzOwx9W7FQbonPTp+YpdsYYofiTLzd5nhW/G2
90CgjQR9Ht+n7kmx4+gTg/mybFpxuCU3dFlN/8UaLDp60BjC4BC6Z/I30wWCgRuBe5BCOmUXFn/s
JSPxPx+hvQzPF3LLeuT7/xNpWZOwrdzOlXQu/SPgmJgHC3Y813ZOUR1aP2d3kL3HwEI12q3CFiuM
0RAm1CAby9AfxHY2qHlbVOtsFgRk/G+GQuWp2l3OnjHr9WpSnlZraEzJjJaxWzjxvj8olUmrwmXj
djBxCUM90Rdgggr3xP+SRYKGx/vJcsdS978S5Epq0MAct506ATNiqEiRsnCQod38NBvam1hnKF4C
ILw6U+NXqi6je0nuaKvqmFOE+kJu0pCmLkaRoK7iiLazT0OWqkDWpijkEs7vI28bV1aLyeimJWRN
+mEHMYrDe3bjH8wHsdEPXIeeI8Ywqh+gMDhKAwiqkaEz+TWH9Kkq0I/Z+9EVR3BSGy03+gmyFxHz
jFtz1l6BZmq4Xe9Ek5AChz+lQINh61CANI2XGPNdfIBmjbUeadphJicD3gki105EqdTTqE0jrbVP
NPAlmLK+oZOv/sp9kbJdMDb0I0lNDSIhbImVvuchWgBsTJIOFeyhglebLz9E211hRJ+JQ/WN6UMy
+j4BbtE4FyzzAi7N8p5gPqaOXFAoJLJnAXB1Evhkmd1IWQjjTGAC1DHc0rUtutR8XasfQPDznhKl
TgCPHAXO+LMzQldTeoAH64VM40rXNPVD9n+kdK0p3N4C29AZLv/60nwVjmleo/MggArKDEi7qnY4
ZEyQogcSteczqFapIzGR9BOMlL1TVybEWZn238m9t1c50+awtNRArJ+3S96YH2CPm2CjmyKemCZ/
52JyOopudXst0rwJ9Gpxs4pPMiWdR7hBJ9flmCP4ESc0/dkMal1vZZVAy5g0j564EtKsgJ77zN6g
GuMxpvQ40Xmm2YnZFvX9U3mOJGwfELzZws6Ajm5OKqSUauV5mPFV4HJTPDFIBFD3FhZxfyUygbc+
ljHgmrDSrhgkBczna/fjqDsKhOEwDK2rG6gQXMS/otrnLY8gAxcJ/NnsJ81NY4LfvOAm7AEHfQ2a
zTeR62Tee2zmFHzt92goZgFOemws4cy6Ky3vGF5XR1D3LmLiA8C75eoMy/zoamXtvyfTmW4pNbOe
/X7bOsJ+D9edndeb8Zb+Xai8RG8T9mNo1RXP4oR09jQvDRPhFVpjCKmXrMyF4KzbJ9iePUmMGR2K
sJgozrX9RdY/8X1+j7u4G15Cz/yogrOML+z17ACGai0MU9861F0IT7VEZQDdS0Vg5cAlvf7ACMI3
HU2nIrVPjYAulxE+OLBH0il0YhXWNr0r35NRAsiZ7db7T9r9v9xGKHyRXj3xeTfYRqRlGvs2We39
3+t9dPjlZ3B+3Gpn5UNUz/AoxAhFB7UJ3llk1slQlVDMoM0uLvWHTDsZ7E7qmuItfjaDaUgLnYab
zH92BbyjqvJE5r+3T1/n1vUKdjkhXMVTs8t47A/aMRcLGT2KLWFbTl/jDgBpr/SqYQcQo3QXq0Jy
E01Z7EmMmp/e7TYS2ewDB6zsxFI2uLOEoN6ovkN9H5YleME+WsmXN+K7xRfPuIUbF4UUNxm4DPDK
pXIx8ws4ju9B5L4jK7mpqHQU9woV5xlttQfy22wuUNcqYKknxFTik29U1vGjISgoik/Rv0vgFH+W
FLmSzc/fFwSBesuydP5w8PjRyqdFo1hlZ56EKtsQzqNoS0lCSmJ7xxXIoScc7KF1+rxUqR6gkl68
m84i+Sa16lCfDJvLa3wV35XFCdpURtZenEUQlCpP+2CETJ2qBa/iicnn1gRCn2zvChpIrDOB1fLr
ymy0ELPRK49AoPxZVptc8HBagWQZaQGPHDAHH6s8XB1pTYzXf/Xtr/k44f2dbUjaeRlpEFJC0+/B
Cq2XvR9icnCjUUWe7bQXhzaOf54RpkjhI268ZWxoWeatnwIwus7BMThLDwNPGCsStPjRbttKbpTL
yb7HiLq7SPtoC2xKEFR+9KWbWHgX/q8naAgIv1i0MHGGHRNikujDkUxxm0CD0ebDIDwhpy1qycAl
VWiaBlESXvh1UVQKXg/8ctPtz0azFwxCrt45sMwob+55cm3WnnYd/Xtv7Ok/2rCGr02Z1/ZyzZzK
KLRxIB8Oy2IJyScb9EKbe/AoX4coOhqqNPFBB6/z4U+/lXcViYvLe4Dkn0WkUhKyvWTQ+DBF0RGz
qxadqNTO9n2Id51ZMJfXqX/PW7u24v/V9MGJrCR1uQuHqV3BwzTTvJBBHLK7I26uuO2TuyWP5SXo
XcOuiKgaetquhRHLtdg4KccuFA8T7HtZP4kC9+YV2RZVkMqcSCDlAYS+J4NWNUZKPT96MiAfCbaY
qfhC7ouhvf/9gsLMnFnVgypQTrwe4uORIGLlH6KfFidRchnaKFW0U6052s/6VIroU3pJLufp1pyJ
59/BT3zacL3C7WsswpQNzGNHsYiRh/uTPH0dhMiH1YM5OmEmUNUlDuh4MAZslfSZ/BS5qD2K8GIt
LiHKW4tu8OIxBon2OdDBTC9DoJbFwWN/HmV442Bos0FewuDcOlwH5uId4zcb8endRPLPDZCa/eAD
LGGLan6zcBSqT3j+LN6TdVruNY9FDzgRPRP+B08EnW9M9LPPp08lwZbD7Tja2kv/eSv9T7IVMjvy
CgaZCIXdkBS8cn88JQaEm0PvhcKZ75cmaFSf1TRCd56cBUCBPlARddc25aUiN5UImCQohZKQgvl3
fsC2JrRqNRHA7SPB3ldysFmAcKfnefL8sWMTnfPqvqgmGLvQxFKZhsvT8eC0enEpFwoCXu9OfaYw
SgfmJUw3a73ASINrIoxHdb6Zay0KYIIRu0gB+EObEdNbrbYNeQz3wMoejd0jf8Yb8SJqo19hfHbJ
GmUR68JJKHzctLm4fFT502LqmL7YLdZys5RAe+8T+5A7OrWHIjGv5aAbk1/R6g+tmOLT+IsNbidk
UH2T6R8fA8CjtGK4c8JpQm8g9KekfbjJM7hsCjTDrfx1Me1uRDnmyRIClQ0oTBGVjNxOoUqa8GMP
H7edlHcfCNzLB9pssPM3lv49I3r/3cuXBOd9878lgKdQ/uhn4FPe0fHwRD45u9F/7OYKpUJ8Mk5D
bng1ifMECT6MzzwSP9Z9ggnFefNvR3gG8I4BVqSfErgsQebj0xdkbp+8Kqbfsz+OsjMKywE+yGsW
+wRItL8y5S129uzwZsH1LP0/Eeyci/MzIgwqP7NnYl9MowR04Yxs9WuZDIrag41h6Q/P3LH35rfJ
jCHLaajoenVVL/vfuDLO414VYfy9cKEjbExR9MFZwXYKtpwCOKGhzy+MCSwaR18rbiRRWlabvNlS
h4GDOS27ZpO/Amj4OpoFS9MWYJXCUOsMOcP5XJOvsjkiM43+qBsp7+2nlmBu/t6YjV54RYZOug3c
J36chafpuKWQLqRKS8XdbXa8vQz4tGpDU8srAHmhqsG9GyYR+jAoMF9EkmBhcUXxGzn7H2I2gIf8
Rl0U8QhOcSAODE6/HlOmFsq1VOIaIqZf+YXdwiTrGTnZjnBhbM0uQAAevu5PCqJOXGm/kdmlmlWX
m3LXYLTX3UDvM+NmXH6mBpCx3jm/XR+rGtkBvYirb4j2oNpFwKsTOE0TYuvX5pimvtj/RFEwhrzT
QTvWqT0447KDw/lj6aoCmTS6LkaVFjvOZfJ+BwdHW0OZS7NzHzwqdIATN+Cznu72yb4l91lmvZTy
IOZRIT9aKz1PPvPu1+HpTiXX8Bvn9N5XuySnd0gypekyhtSDxjunAA/JySslsolqPsNLz1lilDcl
Gdr9xRfhT0InGtnBuFnSjOwqZ18RlkKOlOKpqMeZ61VokDgDIT7o4gaACPFGZaSKKZbrH4RKFYyK
ApxpzSmB/Bh60VzxxO5vSnnKILezcP5WuPw2XSJQhWE6k0FL3zAx5Z7a5Z9tDRgs0p2gWI0V2p6x
cf9Vsh2tBeRyvv0ioOvS96aiVWL76zhR+Sf5ORkwGFzfzPEHhQNhokWs513trBp7emLHj4N7p/nh
5aDt34YoD69SVUnDpqd5EB/FsABUy3AHubuWWSgWPxvueEOWx+oo6TvQBdlo0F3FZe1421wQ2I6z
/zt28L0MdoODBtVD00pY5S+F9Leu2XdsH0gEftHYtq6AoAzBoX1L/Sm7d4Q0vqwQGHB8m2emUlOw
lqbrJuaCuLfuYUg5XUNwTblEuQ36qx9G3/WLs2XF7y2ECXRFJIzR22PDkBbVKP6gv8vOTIwInXoS
zvUU6qzgox4bgSW7SoR3G7Ye5QM0teMYHNYGjbc1/rTeiyeidjRYLtHRPHUSQPX+rcN6IMPyRkoG
m00rRLRY/qx1qi2Y5yjeqskqQmBtk3WNM3NKnWPWSzy+3OAcH8Y+lNO71olblU1DmKa24Rqf7KJ3
vObfBiOtv8UZCWuSLu6+3K+uDCdp/+Y9HqQfgz0ttZIMKPwr5TnVe7K9/7cy7oyWMo97/E5Myk7s
UtC72BVwz+cXTg3+Y97m3UX66gqRN5qW4v+gdqe6qYhhOaN9IxNur2qlly23XoVpiuJuMuX9R7bc
LfjxsDKjFj0jI4qQicShgJzcxDtgldOnaKjxhooR18jOAJj6+R5hmv7at8yh0rlaKqRGu9DCgPzR
eDkpcvjdFsgRZ11iQ156dYwqzfUNH3VajLJkGESokt1ISmW+WjRdasvi2FDEW2oD/3h9qGjnLTfR
ge46m4uySk3Dv2EP4yWPMvLFKHIe7XnC+2RFxMuwEB5MzE9HLD1l7q9rAv4xPAQtXwFivgDJBEw1
vIBNtv+A9hKi9hh6nnAJbnRxvs0BEbLBbp3VHLOR7mSUemfeRU79vS/hmQXdbnZmP9+OSOhCa5Js
j1K9TaTenOcUign+KgiDNYJnkXQskfvSMQG0NBgFJ/zg8Tv77hSnSpna2qXmgO4v6lLAVZ6iT3Fr
xEYA8nmYFxRM3MGf5bz/mYQc9r5X3xiHXnlz7O6npNcPYv2s/FbVYgeqgHKlgG5mrMZlWqJJTR1H
+GMrfbMIEWLjqwFA8ntfdxzY9rnIH62JnbjqxPjgjI1CyzobGGsMMKGIJaKiYuC9Ez2z+UX2g89B
ZzbH+MrErHr8o48WHRqqjH1CcnL8JJ4gY6F3aqzQkBg2cJ0cz+IIRJjmuc+ujaA00mgCQcyj4KiP
GtQqY3M5RI4omkdGCmqAuri+7hUZXpOS9hj1fIF0w4Epo64HvxIu56YMlVDwskLF2Y6MOFnlJVaz
GMi8Qh8WXmL8BnTPvc1Eeu1QsPFLJnVM4tM4Gvx0s62t63hQfzUexrAFroweI/oL5TtnetvodQ1R
5ZES3WTuRBOTXudrO2uq3X4YOeYfOqY94MacAVkvaZBuLaXnPjM8BqpfjcSnZtk4wC/Cnj+EbWaf
0T43THhfFc1IX6SKVLF491Qse8iHzqZHsyIH68We7GEWNcedGXt2+kTHtV0Kmas96T5BFrnp6EX4
qYemjI39000fKPHDcZE1ZoOM0TJt8UYAIMNzfUAdQRlennif0ukamagWUWq/XEasHPQtmo1zPcXt
RapWCgFx/eg9i23ayfqdtQl2L85stUwG+uVJvIBWLa5BqYpVZd39BxgA/BooCjl5ZseMQS4zfSop
LQcsFR4obKwDE46tnYIo7gq0u+4H5DP0IrJa2tKegBtPmiM1KW5dZMoHtZzxBKbhy2S8V/ir/AUe
hT9C8SCYBNCrx8F84SlShCoBbVdwZGFIKp6Ydtcp9+QPg4jWd66A8kLrJ1lEtB3CYGp95Y4c5ciD
iKbmsd1igJrL3nRX6PFcnl89bIR7iw7gmEz41d9ue6yVMU0fEBvHFyvN6xYaLSgaXZoeZK3vsDBH
xy+NzHIfV8GLYWKRmmhF0+K/PlQMHE3eHY8THltZFyi0Ag5gaMSPwURAhJwXvwH2Vzh5nv/XOfZl
CnKnhlcYYzB5e6kVUMkxDjOcTWWncQZlj8juH+EiIvnyKtzMl0Ss7nGW/d1yCdLxigsZy8uQBvQI
nNpXqRSizr6X08L881WyG9dKYsmhp7QHhFL9gGQc9xapA75geBLhCUODU4DGiXQxbrqMmG3huD3r
bGJYQilwa83+7YEtgZuS2RV0dpCNXO8AjHr9W1MzoBAVE/eW7PUmKkLHiJfytV3iNizlkpXjbefn
h1kg3nZuVBtijtgionPy/UEF2AvSgxhPbS7bWNCcl/jMSdil6ioIr2kAR1f30PY31IoK5XITof2m
fPODQ/T60QM4ZCvs1FUGbUovLC5OiVn4UDJ9zSz6OKUaLbE0ZSNoFqiKAkrf67peDQg/rjHVwxo7
XIuJproFxVatgfpZN+ngmpmeVbl+P99YYuGIvCoRpqPd/5HwwNNg20b5ASv7N2k/tszl+k7pGMKE
yuWgDzPSLdKk0W7Qdd1beP01UXhRPaVHra5UtmXdcfElta3OsrEHTDbCVPoppgwOvxbh8a5H4X3L
HpVn3lu+h8ga9lTqKN73gjwADERRqh7Ik8YGNAWNwlzpMsxhcr/ND5RVkheU8IlVmyf6B+0G3dS0
8lSw1Q0zHSk49NwUQjz9LY5GLTok2TEEHlL2VPSLeGAsatWerroUEQS7162RbltLD3ZFY/P42/EU
s/0Bg1eyxaGe+I31HpxyubN+lTdcWcF8DUnSaDQzcvLyMBj4CPPfTWzlkuGWf/WftSaa1LK3GQB+
dqMyT2fsGsJGB17YxHT/5AJW95P+vAVBQTHqi3qVVuYwrGXZYvUY9WDYWH3tzvSo8/7YAD7FTuZ5
ERxis/8Tfso13ZRpo51+lo4V/V++OJPi8HpXnG59oqY54u4s8Jecs/2+qLZFxZU/ya+7mU2huWfs
Uc4Z+tvs7jZHYq0YZJuUen5IKDPBFU9+P1PF42rHVHq0PzZP2NYnrdEhKPMNCahsRJ1YGI54IE6b
ZM5PRk+w0T2IA89iC3BG/OjX7hfTL1RvuJm14vWO32efSfBUBc3j5HBQwmyOra07031qzAQ1sARt
TA4gc8TI65fFxLioPghJfWhr7L8SLoVBriU+Xzb2K+RHT9whjvTMBN6gzks3hvD7nPUXzYlKkqAz
cw69FNLV0r37jBw5gfC44TadAvrpBbWptRQ3ZAjQWDtF6LRAcd77t4orvRu9nm5ziEaYk3JQOhZ9
ZffCpPdvfGLr2oVCjvYmEVj7zhwz2ALE7tQ1QNNTNzJe6v5ZJdOhY34go3+lP7u0BExAqlqKuFAU
dKg5pBUuLwSXW2UWzYDCr9cvxYpc4fYvUo/4CCGD8A88TpPsy/ZNDqqJXe2I9Ewnu/bL5bqLv0Jq
AsYhJuVtiTcxmX9+/VFPLlQ+kLqPLnckEb7u8qtvNC4svo6vMspPbEiU2cbfH69mOhLR8b+D0tEd
L9CQFZYZ1P6EEEu6Okc+xcKYzWE9H5vfSQB7Vtz0UU3H+YK5DPKWnBFLzoEhM43wX3RG/6FkZdTg
qcW17cNX5ygm976q61HAMhN7mEoQ/8m8UUUx0C9P08SO5RKhr2/PnKbbXZmdIBziLC45b/4iqtaJ
lbd/sOUMtsGnvVLM0qmSgr3m1S/nE02FUQEUd5n6m+/ZMvl8+Al7I6qAVFrNCChzb8fCfRSe67mO
OfDsSt5iLMBVK4vW6+fooT6VqjzUkvCjS9nj4vmhtivTuF7WOPunfzgk1ilfZtP8Z3+rYSwyoSGm
RGkVUdLc1v+0KhhYDdGxKFTBwWKymjX//+Jys2TrVzjxKeyroyLELTDOSWaXUcE+ILOlbUH1LrKi
TcRb6eM+Vvz8iihMJXxR5r591BSB5efFLZls/D5biBnRVYxUsSvSAkPQA4fmBEbb5PRZ2iz5c2o3
5n1ycHbhFaQTq0a8se888nQ3wazU3Hvs7qrao6pU49Aln5RnZMLzKGbAEW7f9X4DerRcmU9beZel
9Y/7IKUtnIUibXULZ9OjDSgU2lpyvenmefDjv0f3Xddfz+1K+6LYnxJ86igbno9D0z1turSoraqK
LPCQX3j43m1+HqRPZ5VmMnpWNan5+jAbXrJLC3gJF+PJo6QAx/7PWNPolqg6pWMOGlPyPX2ue7ZA
1QDwJbfAg6ugA814RVD3jZguYtCNHsd//9pWHtKwpp8mxTk8s1xc+NybeFQ0JZMwu7QwIYvTizE8
/febL/+nHvsHyIvu+FR+qJPbNOL2HnF/wToSYbyDNKAjhzkndLAmwPyR3xgGnJANAUzvVScalFcB
cLWg/lns7ywZzB7P7q2aDsYvPsEbGe6c0FbWlABvpEdH2vaghVtFKO1zB+FvimV0sZbgQa2JFVJc
tnQ2KGHEM6c14HFDERrCo4UDGxVvkGH/pCkXHYns8xAbEn3OskhZGaWvyXZKrMTbe7ioZciHrMmy
7RbrvNB4Nlgtk2O9nB+TsyHgaXObITSGKQ2QjgC4BNczC4qrvZb4t2wlkUjfgCcc/lornsV4CnJH
Xj22SPlTMAFkGalFDokuYqkearz6LHOcVvq2c19DZMDKL5ZD5ozPMikyrZwHyK9nOl9oOaMmXEl0
JbiSX6Y1644eKANkKi3kVVFfo3jFRLcqUo20TFf4cfWaAHZpWYU02iKoIvC44U0RahkGqtz5wnIj
5Y3rdPGByeo97i6YPBNTOwDxoMtPhcgU0mvgts0i+/EQuPWIxAYvn4wnkRmfGjTFzwsmd5E10Uv0
RO9Mjz4Xo4gQNJLniYWayigQifyiORhP1gu5hRNmAw/M/GgOc4pNdoGavJ8E7PQiNhQ3qit1Xlib
gpY0/4RVHn1lpuV068FnOehdBjMR8rASyduTrRnydoKerMLXfe3ktFJvH+ts2duVbhRU7EzOegw4
NgcbguPWKkMIKllvZzOzpnV01I+MvuZlcdO9GsASkhTLcPvToIDg4Oit5Zy7TBUbmMXfcgxg9Er8
T94uMKrcFCfel3obD1u2D33yKOVvQL2wh5MMuVuI5yXfrT++3MC2ckWgCO52ZzLMsMzmSDctUEOA
NGqYKnE7rdYx4/ZP7SL1gBFld5nfLYgCnr3ji3c7iun4CTz/1jaM/Ngilg7Si/+ctB5V6G+m2jAX
O/Zflnq/yoSwVevu6m/2GoHSdbrNgI4O7lMJ/ISddgxSni5SQ4qe9H9JYhRA8oHWUJdRd0huZrC6
ccyK3LJ4CRuYUumJCEb1OXABfRIZVtHd2s5dDf3jn/wghGkGGFOl+NXIYO1P3DWbj7k6LBhwQW5w
f20wZrFZfXz6kDgd9M1IXU90va/hN6PRZj/5xHi0HgeaEN6rGoWncDcQqGuYAtXDJm7jdxZgCsUk
paSrnOdl5WH9bdVRNu7oSNBpRIF842NgjWQnPS1U1IalonEgHzy8Ntl37vQU9rY9Ef8SfwkHs4fp
0XMlbsWi6H9qw1c6MwAV+1UAdIcpYYjekW9htJl2ScUfZ2kJ9SrMq5ABL0ADBjpENN4724uEhMHW
dAPoGflchxHViEWsZi2qUyEkH76lXsajz46bZt7Wyi9YWUMg46PpWeLXSKZ2j5EpFdBpfhecSB3Z
gJ1tdmFAXiJAiiKiOuGBsIzHqg0JxvyrnN6kEa7ublkY5E/rw03LBWeZQdUna1n3iHnVjCuEyqqJ
Lg6G++htIz50shjWA49APpVdIxHrtjr93+Lthdei299JCoXXyButIdK2KYpQwrYadC3RzJuFBTk+
sE4Lb0jcn5j5ju6jVfUi4SY7r4LnkgkPXCbrP+/V3/jlFP3NsGbDwclG5Pz5bQbNgxUfC+vVfJPF
s7pixdasW4ThvleqaYJtCpiiLlve+LPjMFfQw26ORhdBrEl3q8Vr/rrWFIRpvnRHRZYx4Io5jalh
1qWAf/GiDa+JWO5J+SAR2JykLFnI5PAwjJFTKT/PRe1v1MaKm4yU7ozKIZHhayoCmZFLxUanohXF
3cMGj7+F1AbD6V21HiYIG2dm6gpW9U1puE23ls2C2nhwVh9paLECLgfGGmYaMQarxjzogoOHlXpN
gMG2Q73EWrP2/5/6FLIZ+B41FQ2FRvEkOB0X83n/ItBlzKndJn3PASgYavf2DSUtz/Bc25nUH3i5
c65xaKvd8PaMaH4G7PqCyZ0Luc6bk9i5CxK1/OyTnB0nAIlcKKadA6gUXqWvxZT6zAN3oVHXZpO/
9bPhOiEUyLk9si1M0dApUSiZLrZkSGTkiGU286Aq46uHtD+QUCvBukQUoeHegIHv96faEqxIoG5N
8Nnb/3OdFgIaJMMdjaVDX9+9p2Fav9/zgINoSG0r8r8WT64Z7GIqrCD4L7eKVZBaL8xn9AqDZnwH
KCZ3WEenyhaPUCOeSj4V8e73wBjMt8/PpZ5EB0jQ4E2s1UNe4Yxc9BZsRO0vIxGf84JEcbG9dUNO
H9pzqOQib66eeSJdlO8sbnR8dZDvBumK17IGnr0DYa8Js4l6WWlxwtMGd3aoFWWLJJ4cc1t9zaSF
/a91JF9ErG3NwOllCSfxIEhzrMEKOKvp4n7ZpBJ2o99IDp9/xeNpzh1Ps9hY0tDBGiNBmqdCDEp5
9E9n+AKqx8laSZi9vzVzQ99MpFHiVg4Ub+5OA2xwSSg8SPhNevBaYjeZT87SFBIvU+Z5wMW+vlHv
QUpS8wv2IB5PHn0DfzWsXbX/+qwl4czsvYP37BgAOgoatcm9XzhXKBgiRz3xvD4rsYyFJfKHyk85
fM1vT5UF0qqX2WME4KfW+1FvMHpxr8QmPQkRGsPLWC84mTvkS9rLxwd2p/RR/hAB2vUm+RncsFcZ
o1QeB7YTJd0/MOk3YiOCwP276MfCzoC5vPcq6t4KWCmasTKZ0EcdjQBvofktKMBgNzF5gYvVhkgt
//M7DskJltZrYxMeE+RUzFIBh8+Sl73jJSJIlsGXUcAX8UCZVBvoH0LpB/0e6YncqkNjTlX7q0dO
JNwgSCZkl80CZw7YJf/mixWB6oIPKuDAT4tF21z/waAPIUmp23ToNjxGP/dgsH8IvtR6HaTERonu
Ijfms5inqjgoYtkXC5UtYWCcZ4q1LNL4kkyvEU1X9z+jvIJNe23YQsCuA3UXNvLOASbD2euuS1tX
9Gtrh8rl58iCPv3gysriPgVN3Ve64NpFSTzxu8XpvmjqDeByD5lOOdQB/fvhoO2HW0gMmXAaef7m
jHiGFisrT7DImGggaYtnDVmeIKx+PwfADXMVxS6QdfAi5vyAvFqkntjaSUcxKQQxiwehQTUimMhi
g/UG2F7Mk62tROtWvkuznuMiMI9lLo9/DMjJhlCtHegQwLwoagcbIgdtMUMG6Vfwrb7XBs0yr5xS
gVgoWQHeW7K6NC8+Qk1G5aHG6d2vYbAZJKKV8wgmzJeJXgtn1cxzCpyHhSFoufPDtkD9gRwK1/rz
dGK+tFlLahOFBZwtuccR4v0fICJ+zqGREE6G2tI3xOCqk7CS/WveB5/debuY31OBRSg5JdpgXHxM
HA8QHSbs1tSjjMdbw4hN+tg31iYVszKAjKkoyZc0ctN8WZIsepU5AvMJI7TsO09RhnkV9DHqQxLh
O2hdp7CDHJaK5JIVbbW0WMFVg+FUAQ544B+Hsz+N0mYFuS5BRLsjRIY2/Nde3mXetTm+EJuqTWCP
J3muEqBWrCWrNE+2LMZkmn2oWnHMY3EpyIKaQy10PACKOkC5pfb3NwdKqB666BbOu7ly3nQFZwvB
3G6Khi5l1zPsnGW/hYUuAONE3wIHm0eEc5bd9qc6HaQXRBwoLGktAO6C2SK9qfNR6Rd6GBRfH/Dh
n6g5Y9YNbcEt7BVvSqTQtAqzU8jTtdKN7o5K/k9REPx/iGsqUbN4yJIKLpIXi7FJFhLJ8h708lOb
WIrwLRyPgAUcDFGj8Z0OjTV4dyBBdVb0YpVnOh7BQ15WqOkNsiW3rBMTjaqZOPlOQ/YetVRGU6Q+
/YIN9W1CbKs1WGNJImnC5wy4P5xRP717+4zCZPl9D5qrkahknDV7HDSBlwGOXHMzbRP2ecOVlTiP
bBbZQCwtDWAMIY5bHlJNyVs4DKDnmS066xabzyNEpiC8OgMK1OuL2zT+U8zVS/y+ujhDDQsyBRCL
YV2jgVIfdn/bErOWIW5WJofu/V+zYzzy4u5FzqM8KY6P7VvD1j2LjsSxYguYtMmkvffO9KFkBcP9
hIYJz9cyCJt6a+KPwGXfkvzzyrgfcslBg2HdQvWClJFhp4v6p2J2WmG3FKxe0KE6+O+1wsPtc0DQ
Zo0dk7z+O4vERMZiX7uIxWRSzgJiaHCX+DTr9xRuEF/UvZgki7thDPEqYfYtcIyc17GYB1/Ql2Cx
AVvMdYraHVWOmZtWsQK8rW2SSdP7oA/G9yGX8LxOv4A2z11vJOTTnklQqyiP6ANp7lXSHWdwNRUy
yMR3S1cu4QaLiyJLJbIgsxIGyJCX8o09hbuJdO93SmUstQUB/v3avfQMaky+MWD6whZ93mpaBjYD
6/EM4pQDljsdcsv9CrYHKn9PpWkcsZm0gLtHKIjj2a8UsSPLd6xuBaxgHOy6F4mjTP3PkK0j8VVr
y4+gaX/GsjyI7UT6VvicujXbZkAZZqP1r2yA+ekhnFs4JtjpyTxOJvHeHk1eZc5iH6Pa+CYgYk1s
qeH2IfGPaMM6alV+TpRW1h0iB8sqmqEadMqH0qxxdOwfbDB6q+CG36uPS8F4xVQflBU1/IBl1t1N
sgTa392uNrrSzMiwxm7uYbAVev/Nuw2udCIED3XIUtvg46BGJi6hlWUR7RE47EgJbSiGW/sRJjQ9
b+DA/+oPy6/L45Vtxxk+OGdaV7QZUmgNusr/umzEs0+uFslHgo1STweF/0sLPqf9/scHVabi6tKQ
K5KpsTnAVAaG/wmpU6YlQ4j88bO4muEUWXF5sqFMLEu9qW9x+flifvv5LVZxjLNZzYWWpRZmpjqw
gEulLXIWAgaV+zBxrYiCT1jqHIxq1Qkk0RiYrYaDCVt4TmlzHtqN+GoK81CxDns9DhDqE4JWDZEj
0dGl+iPtxakt3bG+vI3+zINYvSLaQvynlwBxwkbx5mxUWf+SK6+HcqPyiHPZEQte/nN2A3cvaWD6
d2jYibDO49HPIJCtTD2tRS6Je5Mm6OKoPBa8qDpSGY0D/G6uAJy34oMxY2a8sQRT6lJvUJrPZhB7
7hUZS/oS7EMdRS2bdATvzePO2je3qwdrmDjzWmDU0EWfklSGiwig8c993IddKa0eR1tEwlFdDeVQ
mMi+ZNPSMKwvFHYfFYgLy3vv+LRFT20d2dyomng4xLEbAoVBc5D32Y1OlgTaIsSPM0rNcZ8wDBSJ
0E4KhguS7v+1w0bsSrQMSJwnZCXRUvxo+Tp4Mh0HX8ER8iILKP+grHGYMQhWG/MqybxPJWka1tHE
VLmh0lBHUwsGYPMqx+JRCAyzJBdAcqmZcAnUMITQYfpIUgNTm0qDSp0xJxes64cLkGYsZc8YubS6
MC3+sjidhkWtqZcf9uEcWsFCGc9ZbxO2XhGr1eFwic9G4Quj3Ll0SBZWERt6GmO1/PKVeY1hTg7Q
jFl8FSfN7GFlhkFVSkmI/KvzjYNtCH4axKMuiSRs7AaFbQw5YJu1vFcd9MVJ85ilntPKorD8GYT7
Yow8j1IxV+YqwFqiW2t85NOpJwaZL17ttH669sdi5dcCX7M1uEXPcpjAob+YU0baIt1/VdgWolnH
Xr6zKA49pviYSIUHcFByy1EvaHfTCp9FYKnJy2d5FP1xs1rc3eUp8osIj3MBG2LP+rzx+8fXXbKy
/bAJpK6cO9bYYqvWMz19pI5V5+xloU7pxG9nNQ+AoCq+p/jOfRbzQRhm2CekG8xozsmbw6e75YJ7
WcY9YGttFYXGvRP8KUpypfqnMuRuqeFU6sGYep98zw/MMld7iB5OW+dJoadQcSTw7B8XF14d+cgy
iw+MGtgH6DsZosB5PzMR/OhrodlU0qtGbzJ30eUuw7NP0bSBCV0U5/ee7U/uXEptVpkY8ls0wa32
2aZZB/tvUKas37IvhCaM7rNO+7ASOoTr8c7To8Haomw/mZmQPz+s8cj4VKZRI/8l1Oh/7AE08QDQ
7Vf+NO9p9XYInSglnMQjGfVXwaGk+JtXFIpbexSnVAQqGquHsKzYndzbXB8rvZZZ2NW+kjk5k1IG
O+gBpdvgFkXOmXVU0eFYOO/HBVEpyT5NcdgYoRCsxQSbpEJIAXwLXN9GuAWg2b9t3PncMIMFhhLp
NQDIiZ7pmKxa8k1eQRZUkBAljQz2j4CLg6J45qMqsgllyp+qwVTeCh8KSsKbIYLEVStGV5fK0Eqc
7Ignz05xzpZdVhZ1j+IyRHIDxd5+PJ8SGJhuiYaV7mnNNkeg6ptpjT38Yhwtt1PR0ZdAp4J70tvO
uNUKV9FOKzuJaR2lq64rx6BfzGeLxo4Jvk06oc9F8+Ss0Z+vNWSvQ1C/scE2uddt12rBS+s+MKmN
cE53/cc954pmRowOlmbGcUjTMdSft37hk3kA7TFMl2ltWcqDtj2c3jIeyPF2VE/UhKAyC1tM8Px+
Gdlwa0OOLl8j9IAYUHbzDjGS2H02/FR70okTfR2oH54iEzcBt2wjxBK1YVn9Uz92SAE/W6RJUU0e
/xlZm9JUd1qaPJvY6JmkNjntbhhv+YTyWDsFE2my+qKqMbNZCg0mq+o84zYIg6iVhZ1fVZE6Ssdb
cNUk08wIaYPk7shJD0XBzGwwI2OfEGWUI5Nq6DWhp8Qn/s04wHz/Y8Ii8om+Iz9hx8F5TtSudfRN
1f54JBgNWOD3IbXEyEYKP+5/1V51MmN2yo/ySNGznHHEaE9cMfr0COl3VyR9bbX3zwfWPWCotgZ7
pwkEEEMpZLU8KG7hPHXXThg6CSdEwP9JnJaxvz6dPsMNv8YvZ9ubsdcntls/yavYwe9wRjtNrNcP
M9X3mNsCjKBWG4ixj3NOhflXOtEg1VEMEBaP1JjKLM+NzpEFVUH/x0XAjAfYp+23npz6FZJzNTCo
VtU7C5TmG+vTiVfrmsezbDxW74VKy4FnywV9tTUqYMG8TrjD5ITpsSqlHQHtoGMoVe38lM43rflw
phxZFoUPwvt/OPyPRdI92wNbTE0W5i67E6hWVKNPA+9u3JR0m9tyNHXNGFFw8aQukiF8vz5KeTLa
gK5Ap7vsDjvJ/gFOw2031inJ6PRXvYAKrd1vbuglN2B/WR8RGP5GAYhpuHxEPZmtJ7UWRwM3sgV9
1hRrjHPxCBhmZYELhACWVfwJk3A5yVBHRikieW4A+6t5GQDT+2GjUqV3fE9H8rTGmsiMsPE7o+GS
eIafRTjwaAGVqYFxMZoF7XzZCXuNavqFe9lywd+S7VSiP6MIibFRen+vz1z9yTX93oHh4gF4+B5H
f29fmClhrwV2g6h4fSxGpTf4/CyuUN3UtgcLoSqPS30zqgZXKhb10FQtkpnezC8FR7JzTNjDIUdl
bc0fpaPq+txuTHzLTLaLhK5O52hwvBMkNblv/2+c47h8PrCUiD1JalNplfSjtWWEGWQUVgnAB0Xi
Dw7PSknP9067RwHMoIzLg8B99rzItMPxTUsE0XB8KnlY8d6KQmuyYOsgmGun4c8IJ+EL9Pq/em5C
J3NuGZF/gnRqYOeSOlQfmUPu/gxgmWLSA2XLQfA3vA8jY4fLIXYjkOaBj6NcrOJugSaz8CGR5td+
YhaoRFijRmEJ4EJ8IZPjfeTypfSgs4Op8X8O4FubuV6/eagme1705XqOGgkI8GafzcFR2ZKSVmCJ
Jl/7vNfWuZzNhumITwh0H9NGfw+nCqSjrNSccttOrl0L65U86tZcqZWLHpmmfQ+WZ6RlLR6YDebB
GySXRImmLvrctoBEKSg+V5gm2wwazsr4nMfBZbEDRcNTV8f+5gn1McHtxGdKnN/PuKw9+4j+Mx0n
qgR4STM4LHqMvnmIFJnlvxGWhgrdt44c/RvE8lqWUIyQEzHbyTNsqGyIGZSXZsAo1Wmn09FFdQrA
itt6V7vWxz0mX9HQBDBjJpi8NfA3H3Cfzg7WqYYGBABFy5D+vRC60tWYGSITaZB40IOtfQKks7xm
IW2XX0xPj37ouDteKPsJuXBhXjFOXlsQTBS41vtNKYETeeGZC+V/bm0v7s+mxWXkHSWSl4xQ0p/S
TN8M/tGBLOuF9jTe0pDqWJP0aHC3JvUZHH6t/SyY1eAJsO9OiBGW2mnBMlUYt/u/x3qMsUmjgKWV
mOlYyN8RabiUYadnllOw9U//IBMQYKibcMntfqpTFnO9xY0+GYVOkRaxIvymLLIb7ah0pun9swfa
v6CFOLn6tp/Ao0tmbmael47x/v7VmLQ5+L0MqXaKXkuWAPH+3/2VxPvMLaR1MKnIK5/brW/ybFgi
6l9Koz6tAYfCp5VqSIDSVU1G9lv3KR3qzlZ0+m+n2RHvcbml6+BM5XS+xeZlxvaeuXjH9KT8zgCU
gAIP+7QxJmbO/+Oj3DvKFzq51xVkohEchTIra3+PHgJbP/QQQHbfYEBeizBDucEs9HZ2d8BwlVlA
K0XOTf64ie60JMcvCGvlLWhEfwq2J12Kcu02SJXs2ItIvBxHlD5pycGRnzwbbnMe45cnWggQwvFm
mEqWFBQlXi1RpWeUO0WBUlNZyF/uEHcv5Wn8hFJAPDIWGc5rDFWDZKn+o7kzvnrhW5XpHh/5yk8h
34BAerFs5qN4iFvgb9fFUAi4S1EhzAV+VhC1dT042i449MSpuLImERdlK8kj7T1/hMqTs+pFaQnk
yyfrV4VVG/zT2Wn+oW/QZbCFX+HGJNrlbjAxGwHFEdfd4iWQwHFnJvk9i9vCOXWE40IOKMneDTpM
KygTAeLQsWoZJS0jQmFQpeiZpigpe4h/fmfSCAiXSRpT5BOUkCTKLGU3OMKaBvFGULq8BOMGmuW0
jgkEx05vI+chVB0tweU48AbsWhzl7If1/p7DoBvw2lyUHhCMczQD6RJSse/QC3ZJk97megCJ7WcN
yJ4oPqww7Ctl9tTbvesejpoIv5XrZMJktDCL2CcF8vxecNwuEmS2oxY6t6LdgdVoOWfUH+4Q7plO
wRcmvoq9OXei78gzqgH9OczfycZ8Nd+Yx8IDeN0XDJ8XrRp45YVL/cAnW/L1z7M22V8V4wn0MXl8
uhIj4DjcZF8vk40xzpKOj7FOdd/ApnJIkfqNs3xAHKDFZjzrWej7yMSVNv+opX0znZ0Eo5G0bZIz
cFNYlDBJiLeK/nyk6VK2yvKYa9gZJZAOhvqlN3QBDAVdn0GdhOREV5mGBH7h1HE3SoIhQP5TH2d2
objAdNR/sivtqRK/MOM5XRgDVN2HdCkq2XU3qtWQDf4nV1xOiWIXVdluy4pKdgNwx1fGpLQTmG9W
yX++BnWuaLH4rhuUm4/82GfrB5AXbdhouRVT6L2g4CduZ/btcvELsCZ0wn3LJ25aM3QEtZDMcKDh
mDWTB5GByWdZ6xyCKfw+tiqhJrYHFD0n6jXEd3q93MRffG5rIieyUAVWBv799465GSeqG78HngAp
/PUHYHWRF5/xv9jTsgoeg6CeBJ+0GzPYOmxf4LJhX0YBJvWkSE1XIvkBxNiVQyMeMIYlfSduq7gt
rA9vAnrfpPTlQzyrBQhVEEURjT081WII/dGYPy5IvQadmI89bLkCs0fPcxWe+J/y32NYpdF2g5m+
PohcHD8gA3sQFH0bxWP/u7YfVMX1DD7xGzo/fvqZIJvnWVkyXSKLvOfA6zv9gUP5Lrwox/GBL2+h
G7uWBcNtqrx4Upy+NjzHPRE1Bl6KEoQvfIGOnKJg9PiTySNV08N3osKuxrMzFGOX848MG4dx2dlk
swOi/NIJxDLMmguDI9ouEd0AqRMOWnyf+XkW3QwIm+/L8qfKzJAFmMbzVGC/fxEylQmtHdn8DkZN
Ug7sDBK0MODiaIvH358LhrXo05OPQkL2O93aelqwD9xavouWKRj5PFupDZC6ECXz0kgtkR+3CubI
gviQ+3gYgpFJfs/luTpGdoaa3GTiSe53eCVygyEy/hrm+/fxbk3Xz1xiie4cMka2dcAoPQHPI73q
FwfKsJ9ssTLloqwpKNxscuLppJaz5WL0ObBVlK0OHTtofqZJPLZx6Eof6bf3pDNWg0KEh2QG2DLd
wbZfDkmPL0BfnXdqpcV/UkWanHQvevWeqBkqOFfCdphYKPVBMBP6wRZgZ+AKyB/Qr/DGc0kP9O4c
X++UdJGxNdEGdt9sUYxevk5+/oLXNK2WX/s7jLrFEhHlEycVPs/gKoHtDKiZ3UgcdXaSyFw9fSUJ
x/bSRSp7Vk3yqUQgJhAfC6KPA0z0LKy1WuzcCsn++fKgDsxO3+KghKmUpNViSvc+XxFESt9+duA4
pmQzBAHi3V6HjHtXlygVEpf1V0/u4P81FrcT81JgbnlSIFdFFkpNz5u3E1rbEsfweK39ZrPIIqEr
F3GWYVlopXS95JB6MoVdwKshrC4yYQLQlLwMWVJ3eCXgrDnBOBEw//S0isVs+Fu7ZFbYR2hI55+M
J1q+l2iTCw8YQ+ZOp4xLKsvE2o9vD2Ez2BDqsGwIoFT+SSgzGhQg2P1Svji+GQ7/Kt96bFrOHNOc
tQXEdv9W1uLPQvOkxa/0uYDXjUyW6FioLjwCZcrJ47+tDz82yjS1mQvZQ73ED6+DEbMxs6zTzpFP
pQBBIt4Ij/UzcnXmrZRw/91Uy43C/vjo7TmHt3YkirOYOLVObM2QwuPbdONjf8fyQJ52UYUFlp5q
H68aPcPtN2LBkFDDc4zi09yqPr94qGJTdzzrVvUGbp5NqM2opfbG1M1Lp+nMHKu4veG7elQkpIiS
TTBcuylZFt0KlEhEi+MUqGfex+X6+X+/xscdMN3c1NOYvMRrujbf3mak31jWiPB+vOf07wZJHFm8
1kfeVncTVpTVQNdA2QMOu5+wig4k7aoZapULGiI7dO7N2cYs4KwAacberfMABk8fII42p92KH5fX
h0aioKsx9FvuFB/LRryRVahsxmlLB8g194STaSkYJY3i00xw3RHfIKZhMhlWBj0LIi8uTNfpy1A1
Rh0rv+zO52xxR66oKpd0k9FMREVfbFv2yclLzb/UME+hyfsqu8dWDZPfkEA485xAtu1uszngwDYv
ud4gg0XUvpz1eLr7qIeTVitdyYRTtXtdxhOmdZcZSUmFPkxHKCPuFZx3l9yV85OV2WGCHyjaqf9v
8k+zqXGbV/z5boMXuI6jAlGk9p5cMhcDYHhkND+VYvH3pq2XrkHANeQIJCKdlOLlQyUTc7HHkGUH
7LSi3AxdnwqtxAYD0QRkePDyoeFY9d9z7C7vyBMLHoGQUivyolhl0dPwN+20P4y0uqTMt9rwgFmm
zoCF9m+eUQkaJc1S8jcuj1wR10JvJ3HdrrIFP/RItTqAvA5ZeCaXO/HJsUx5jlxnAa/soHprQ50r
RhAadZ3JFzqzHt/7M+6An1GK/qKCp3eqRpbIDTxUqTKbr6QLHSCPmrHQzIdoOhz+saPX+9wB09dg
OK18uDeRTq7x+KnAxn7aScLK/hPqlMcBuJfHDpT6wsao9gMGEJSvDxypiYfbAr880grLsozv/cw0
JgjJ+zTt9FAPAWMLDJk8CseER5bds5CQl31z2ol+/ngGwTif92hTqQ7AoOdSSBwfNnFTsih5K0L+
ARKrAf2pueAu3XA9+S9vYF602u125CaVpJgPNK9SXjqTo+/Jrn37Y/LvAKISp5/f0c385ucyp2jJ
I9eJChJfyM95Vvi4z38xw8+1yBBW9IuOSyK0Awl00n1I7nlREciHmhq+iSDGVzlWlyrlSV1C80ED
bIA294RqZrynsndhmTcUecWNysuxf4sYfk4jT52veHW1hYTRV9k5ttQ3iwDqcbs3jJoCaNF72wrb
5UES6RXDb2DRuGS9LxkcDDiGPwmMUkKHfOC4jM5vTrbVEfBPWskoUHC1INiil151/N2ajthCsBbK
g9BvKNRGYDnjUiwPeBjzIUCMPHy2knxveRrCPXUIEZlymhyo3VeuZZ7DKbU5e13meRISL8YW4hTP
zsSCPMPxPfGB6lEMQjjOBeVJrUO06zxParaByzOiu1jUXpkE6yKGQ2REgpIZp2+VjCUf9xS5pUAh
7EWRLycWDAfK8sPoUztmqWSVGIgx+VKwwYz0nUHSDp1dJ9vs+wzvr0qsaVwiasnDJ0SAADi5AbTP
n1AgIKM3RS2uIaFmAFUdxkupOsTeqwfXFgov7jzzOj6WiFh3ugAxXyJx1sgOtnXoef8cur5q0vCs
FlHhc6QfcM2Ag/OTzl0JlJtE3F0CkBHzspNVx2bIIUpFObqQgqkZtNXZR3/wn9pjEjHQa7R12YJw
ugasVNs3sXywrLdPgryi9P4BttSkf0t+X9jkZi9od24czbxdykav5ZvwT72c5DuniJ01uWMLPKyn
cGAJQ0oQB6P3284RxHCxYLv35oi8saHtqMw2S9lfiYO2/3AafkeYD+5YiZqU5N9w7JeEIDEPRkTP
dzlBG1dT/gSn8q8dcSKP8UgjKTvItnMvpbdGGFoj73ba5u9C3Hds6QkyyUoyJPRBo9p1uXXrzmwM
hIMgjuBpiMxHfExPuemkbcE/e2akRYWxdhOcX0USlmnGtYV0afeVwrWG63paQNdNZQp/9baSTV/+
DRiasz1yI60TOZMQHZA+5pud0kFh6b07yuXeCIab2QuLt9ZCDdd6evgReazC5kI5l2pvT32vcLDQ
Ex70tJWmUDAu4d1cchdBSXKnwJWMnFeCoAlfyMM+Fv7v21x5RhN2NqWDfSe/Q31n1HnP7i8O2RUP
bkgcpfCmGHgqouovCIBMzJyp5NJv14OEXsBCf51CHOECiRkhcBb6tfWY8DrkidwzFyKkDThNY2UI
gWV1IfBKOZJ+vs1KpMjCOdKIlczOspWa89P6gumxCYTr6rG0GZ5/epZ6RmcdukahTFuwyIXJqUdp
mYUo1aH69YlwoylP21uBVIiZ6CnHwnqe6HgcaWf0KwW5eEFojwJrjLu/b3AT02j+jUS7T2AmtBvg
Z/ZXomJJY+YRXPAiCCSS34WhbQhfnuXMApvRoaxaXHVhJeRWhMvVRfS35ZhtU9GsGze+C+9YMN2C
vmKWE06HtfYvAv/hY7tflct+aaftB6j54are6dhXys467eVtkexUZALtDBbGT840qgM3Mv/t1SiX
IE7fsJej7BSzfQ3cJq57hHZWKnf0C4gN6At46DfDQk94iRWxZM6uzlfVh6998AGyU0ieACOudUuq
Ey+lTJAkwDZXCO7kKSfgROTmGGKZUkBqslx52FTUP1SJUa3eQKLXzh7My2/9qO/S5PfkYiQKGlLy
6SIiGLQwL4uJNQp7BX3SVDZhR3YGnZ3eOQ7UKQv4Mn9yn6auBxxzVAuy0JxcDbRKYpl65nbVIlID
CFTjLF0V/l5b3Ra8Ph/uSPHEPZAVzuqZnc9LDFD3MxB6KsDqArH1pXVTuvg1S+arWjDrNyLPeyQP
YWeiuB6QpfSrjFp2FXAZg5VELfhIGYRysYYYmYtXrZVRZTr/hl2vApDVGFTr3MLRwHTb9B0/Zm1K
avS5M63VCacpuOeWRpG8Dyj3iPGyaima/bktRvmhDMzoAS8Vu5uJtSdjYgKolovCxaTyRXXO1He1
N8CwF16Ajdtr3ZAV40AfZQq+GxKyvf0LwTu9SWtld8mAcvyS8IxoLF9qSg4/y1MK8seaQ3kEUBuk
ntXuhCQtPilGY/dPQfSGuMAdLrcN4kLygvQle1MC9em4/eQ+XbTX81gS+rhC5mCjfjjnwu2DChwO
xdyWmuPd9U7kNQnlKK4qWEg7Y+8IMduMJgpbAvCvPx+nWdy91P9ULjduT4McpHr/s9TJHqex5fz4
Ew5eMsHslDoppFCUdwGB7j8cUPCOFE2LzPOMDP6Jo50sOcJeW6oAFdBx9ofeozOME1xlQmmalhQD
M54Po3ujx8OKSS7M1rdU0y4AurTz/SHf7eJInSK7+SVtYcTDwH6TBQ5g/WMe3f9fDfAL27lu9UGP
iEVPNDujaO1E9WUYpcEIGKIvK4OMISMS2IG4kv6qdsH/DW+WkfH2/N0qM683fyM4iEo7l9SrLj6n
enYUniUdFMLNny2vjQka4CAm6hnY3UomidSaJ2paCOhTzyxAxHyirYuoYmrum8D0E/kgZiRoboIP
MEajyC10T1dnT7pz0dqIMfkrFSLDI+xy5+KARumxVv9MvEEu5EneFt3NfEFY2D/OSe8IPpZ/QTdf
8gdV8SGtjYBip4CTjKW9oUnAvZlsK+9o+OSAPs4/IaSu2oZD9Op8riFb+ljGAcgtJdqNroWLuxov
PbeNhZu+fTztdtFROVVFCWqHAtSKZ2uidNWHmqPoD78edfK9tRDE15zrTVr9Vyh2cl5Btf7idKvR
lkbxxXjnVxYPJ50ibYxYrrLO514gWVwbOTjTFH6aT3zOJhesMxTV3Sl78ITphjiOf2Lazn/TlJKo
JmqveHwrmSJlDwdbeQQZRLEQXObDcZEoUuocsJAKSEx3Yb+GuZWI6i71Dam6u6VKvZqup5Y/vqSR
VtC3Lx76XVpr4m+s0mTkl2Xu3EyXlv9HvbysfgFu4WGvtWZ3FWZFYSrgpiMLBVyLMI7MlIdVKvRl
/sCfl5SZRIBrO6iUoYGg+x6UvTYhfDjhEFZ4MNIznB6huYWDYZZwAM4vYwyv/H/H7QKDYTJDMvWN
EHPrZqUFnRhKfVg3ssm9+6bAUZJTIrnYsofB7FaaNYrYcD7GnHqiXz2sqaGaXsQfyxIoa4rLEQGZ
2r0mM+mI4Am1GExB+3fGESWAkIfgnpLHhaM1nocIB7xLgQMCHEtcyVtlSkwp60Fs0tYG5FH9NWaU
lrvYzJZdHFvMg2ANXsNX7MYDumOMuB7oEiiICPL+cTbKtOwJfbBksnR463G4g1ybWP5BrEEvtsKH
bTaGjIgjV3KIoYtgMM9Y0vb7flg+MXY6nXmk6lTzLOCY8ygbtdPDJdDd8ssq8XtzgMomU5tnGK4r
osjPdocUek3xB4589zEmUtFiKdNejxo/+M/tuPyJ8O1Go/B76Dh8ihQ3yf5v/mGwXBwNCqWp5Znk
2Z8aMJ+1//CfXflDEjXN0mXiQusVieRKSQrVxvs8xUohS1b57rlNbgvKuZmawgDBkuieO2BP3ovr
TsiS9T57+k9b/85/oFKpjYYiRmUm/veQOkDkg1zX+vJJc0qi3XL80y2A9kfEb1jq1ZDEA9FMfJq3
D9da8ENsyn0Cvf6FC0genlz1Zbc9C7AuaS8K01ixl0zytF2RBLi3hBG7TuKxNctWvol4TCsmP/v8
PXubPI3UyEHhTGvKLdkTj+pIE//RhnTkMdtb3iMB7WpBDquxJJpi7I6JbbBeHQenUJrgXhk2WlFw
PNthCMZLQMr3EjJHkigMC27hl4RFFvGnYf3FVn0fbupYosE2rG6gBJVYAEx++q3S65aCJ5KA+y1r
eH35d+UyubCxIW7Z8DbvF6mu7zzflBtTZbzuQi123C9c/1G6VlAXImZyoQN25jUnsBznHKxqRUBX
orc8zw1cUXu+TenI4rattX1Cfvm+U3ew0bvql7qfNHhWmuKvp4X0lR5dKTzkY9s1j+ZGzir43IRu
NwD7sHilHzH+5jtf5/w12jpzQD+Av/GkREE10ep9FTIaIw4plcdUZ/+TnWXtaUIgZkjCSUbE4F3u
I/aSc7+99sVHSSxB1qc3lYMv2R6eA6X6+RRLvYq5AOcjwjXvtkMDUEivjD8eenvfmOMy4mjQTioO
Q8Iuml3HUz6wA5gzTIvJIf/Qmxyk5XBqNnseYoVLg9AJz8JyLgaAgkmNDEBX3VTBe0SbD94akotz
JLqShattxWsUETDRuBCLs9lBuPNMQgqWAHAXz5BORBhymzJrmbQ8sruRNZaQPqXi8gqblggmRcZ9
VTJQFSaHgQQQFX2uUZ8zxyFO4mhQlxjLkK5742IZru6S1JYGfUzeQIZdwvLLpAtGhwpb61GP9aQI
VEP5RqE3ywxwyQMac75ypDYpfw4Q+sNFsizZ7wlkMsryCeN2XjWff9S6VnAPCrFSWaF1C+Cp3fwb
2lxB2HPAhPMcRwvDBDrXsgcMqnjZ9yVOM33Lk8X3we3bumpK89bKouDIoiwk2FWVMJuyIY8LXggC
KVF9XxwmXOVvbibYCnaShgDXDiJO06WAbI7hhBkj2mtjqEYWgyyuq6O6f4n7aacK23USJNI2B9tc
hunIFGBUfAKfsOvUXrALmg8izJhrZDKt3jsNLOw0I9MjAJRYvnlbE8HZI7XpvWd/aTZwobgwyqjU
fXWtX3Xh80O5uy0jGpWPOmRUXFqfY2jKtoGlk5E9TCwxJzKMF6upEvKytwf2pvvijhdgriuJ1NFW
oHeIb52iPKL1WbW/5iKIDwRdljQpKHQT0GNUbMp7MMRXL8oNur3IQVmWpMgb7aNfxci4upTYQXns
ceOU8yzXpYtXa5WdT9bcVgjWN2ifN0le/UtNbxu6B+mpp3E3oMEJiX5BASp/o521MYKy566ngaeC
GJXNeuf3ray+IdgRwvYV8Mx/y5Dijytwnkw8cGMOPijGVzg1jBlWjZ1BJHsKVGvQUPXFO+PSm6+K
8Eu7eWYnL9ddi46GL/06ryRDteUcBXg+Nz8VfCvwZLw7CuLLswcE+PuJDd7D+NU6rdun2XQO9osB
Wp6KYtUGmPVmrG7p2SPE1HwOHOuc+vF8/gZO6bGqXTs4jq9JXQnwoXY2pDfB7tqf3gNiUicpbegW
48OLAKt/RCYS2ETgK3VPOun41WbhY3lnMXtLKPahpV3gNN6Z8OYY+ArUOpRBvwvPbkrp6q5WV003
WeKQJZLC7cUEoSUtHBgRR81jkJofzpc/K+8hypfxRowOhzJKijOGhu+RIOr045OUKN8/jrcwqN/8
wHB9goTtkL8gzxZ7oa1JkqxGKpQlYqGnt2Zl+sxpXGg9lovUYDqPNtLlfw8KAKy6xkKe3xt9vbHw
G2cDpd66fxA8CDhqd74wHNDGa7/R5Gk1Gz3JDyT3EYJ1uzIpbD61fi50sbpJs7V4/DcvRyJhrEYG
YdGfAF3oCVGiWnMOgojjfI/I4XBxf2hjfIxrH5r0BPwDX8reKNB/e8gFt/LqaEywZ4FYhfhx+H/t
OT/RSzUBDKQQoyIgTp5Al+SNlAVdNKTQs2EIPGBAk/BAb6h0SBJDD3d8Oz4S40Rb96HSQkJS7Ea4
fII2P03YUTmWknX2JdWFTmyjIQX+KVj5ohv08HkFyPpFr1YQkjSgOivtMTRK8Xn/ULyfFuW/QL49
hHNFnAjt9oc4NsL70MJIL6GZrWg2i3GXGa8nXZtpvNNj7h2m0xJeU9fyuBwucU5TM5ZiFmduNv87
RI79XpeNmRGyxe5Nm5Go7eZAEMaJh5jTFh9OrS3NGC7uS2lyr2vYxzQv8Qt8ZXLrxti7Gp2+e2vV
z78M6LGTXaRjKDkeKMO9IRATaw9VWTYidskca+htZIKeqmd8uSIyPI/r9uh0j5fy4kvGiGRweilf
Io5qOEw23eDlr6OiGSVdpF1F0Qb1JKld3KJBf2OGAmHwaBL2HJSqPtsNyQPdlBHH00VIg7bnbVJF
a4brpfFZJ3gBffCmG850whSHhxRK7qeA5FxIboxeHhftsloxqH9RnwVO82/mMXO/1cSUY0yXp4/D
pcofMcEMRDYYNb2P422i+hOEBHehX76AfqjRUg/U7t13g5FXK+D9NL9kcRA3ajNQ2TgK6ag/6//H
SogmJ3MzceB73rBiUk4OMYbsfw4rl9TrwlXUrcG//bB7p7pnxe8fkPTRj0CuAbctcSi/XO577DHB
IpvnYN4c/HUDWL8WJxRiKxg2vY7iFUat//+3KvKKVMXwqt4MnK/6+Jl5zq7QSZ9y47alRq4f7Ioa
PdgbNoUrEmmiakM3cqCHjp6yqlzVBUX8oaS4IQewDtKyjluurYI+sN464V/34H01TK5DBRjL7+/k
QIghCJK/oFd1QdA1L8wF8+EPlnVPHb7pxBeG8mzryiEWp5lBL95/7zsyliiZp7TT6AinMbvMnOXP
jgXhx5WWPaIHy4UJtodHzFiyouA8XqIMGt+/AoS5gu6L9m/6H6IiALP+c02Ia3+LEgg3g8v/yIRa
uZQA3vg3uEuvZDvVh7RLxU2VU2MiNRUB0BL3p7m8/qwIHxkorT1lxbZ/gZ0LErfGYMYHH0QMHdcA
V8WdiBXwkOlJLVgoDLIh4BN77IGGFdA7fihOF4oWm/szgH4jsjDo/Xw7QSeHcCfeZhdJn7k3pGaD
PTZrZeMgs1M9NAIJYgwBC9GNBrR1mnyzWOi51HzeO6x8ZMvh4XuaDElLQAVXeh+o1qnxRc2OC86E
wgNWTMmH5yMFkzE1vg4EuUd3qS3HlY/cOGYRM4sBJi/5HNWqV/KnbxlWRNhB6Ye57bEuRR+WDzhZ
T0dJHAmrzfnxRFl7/BcRjj48duXOvPWO2bCpr8FxW44rzgmDJupqp18JWbyuBMm9N74tNlRpPJiP
Unv85Tg8+WO6A3wx5z4p/x3bi9oMzz3/Zv67VMhRRdIzD0JHIJp5mipQxtGx6AYKolWTNgHxrG4V
RjZFyfxcFC7wTgU6XAlY/bUJa0QekPR5WcCuP0pR9W4qgCjI4rJ5D4iNov9B9azcudTx+0zwzxsG
sT1mHyWUTRjlFHtKJr5n1N5fv0S/vFd8HXVRLf9NT2oIqmTpYkWjaXPQZhN4r7LqEFqsIcu74iiu
D/dAB7ZqSOK31BraX9Y5zVDI7JiN562CEkWXmIdB3SKRYVetxtG2FGgemd7SsHUvBGRVHO1BpU0+
bvUB+E/3IFz109zrEouTLxZgsxEMuRGGPVP4kEisRJA147XYmUUAB2sIUmK7u7JNSsDiY2zHuSGU
vqTslNE6RcW40C1Xlg2NDMdynnY7XvAiL+039jku6IPw+0/+r3McPHPG4RKf4+VeUg5ch4QWdOxv
d0qIe0KI8s9pqTFIIjM8fYzXkeVaWHPzrFIavOuSMbIFgfe8nrVp6bVpqR1E66POt8h94U4xOXSJ
/X7Ouh4t/teW+hhWHNfvMaKCWCb0ieWe1ieb8LOCAZkF6Z+SyCMZgE/nOhfE7Rp5lJeQJ3Sxojzo
nYlegZ1cJ72/nEiwhkWBqujZsLzLzLG42e5Gc0fjsNAPTyz6LTle7AEZfFy8pgH/qVHbxFf5i7h/
S6V0wUQL+KJ4OBex6Vku2jj2hQY/EwpSqYSpz4LmKcWxvXtCj+95zmVVR5jdH8R23Dddad38RWf8
DBheXroZFyr7q6twDqhTE9qGIBCvRFmHD87S2th4Q5CwVJF1lXAcd/db8quoNacNQ5dfHWBu/9lH
1qHrMeNkkIPEfkfDwbivEfaoW/UH6ABB1MNX5TCu57QxWTC+NHbUUlhMYhdNTta6SoWOoTjvqR8L
5I1PpiHsE2C/ZAhdsQsqPpNt0lbh8OpJ/t1tD9eB35fZhuvpga5vuHYt4YWAucI/exFcwJAl98VM
HfkbQB1WyWeggtFSCzSPeqg6Q3fjElUtTWHdNkXV0ljwnZwdTg+RDUCfant2f5FoqTwf9luEubHs
yvT78VtCT7/aAMo5QAd/Q4XhpTNIc1kARKXwXb7PmGvfCj6o3hc6fXAuNOIuXTgEoJk1+svAcG2E
OL24puLbae1UnQAORHHGs0KE8UHQfjDE6dwOu5q0MBSsI+vhZT8loeAbxJO7KyAu/6XDiaQazhlv
F2kkyw+/e2+ztogZkXf+KF91bS+Bgh7QDv2JXl2cPnzV32mBWOZHRTWsXiZyp65I1IHIGaU6WV2o
hSIrB1u8mKY/cwLRHQ/dEZpLz1mHLC+NSiWyBVP/QHdlM8ZN1aikooMtUQxw5SV1ebSHjQXJJV+I
7IkZUInL+KuI+h6i8y2XdnfjFlOGsFerPP7PcWAo8FwcnjDsq1tkQn4LbiSnZQQYbZ1yn04tCA22
V5gyPH4BiUWAu7WVbnid7qWRMefaPlwLeViqG6oX+GWm2yPmmZP4AY5wSihX55I9N16KFDql8Ztk
A4ZHT3p9LyBqKMHxgt01zeDSxfqBLtRErfq8JMMDeNmnx/iOM54hi2b2xcW+R8LvFsjrSCJ667sK
tlfr25x6T0IHwD8/ef+ilfm/521Wkg6wUGiLM04o88P5jw5GUd+BkIxZi0AHnDV57II+GLpQtZnB
J7mqCg0ByzhzQ2eaLoIrWj70Yr2mho5K+XOVy/4s8n+R/aG95MM0YWKy+6uyA/zgwFFo9o82Y89P
+G8BaOboy+HSvVPaRe0nXl2rK+JD5eNC9KGp/RIys1K4v+QW0KNX1Sz6RH4lXxTjd02Y5FKS0NI9
2lbc19veAVjOCWO/leS8Fpb4NoDYbnCjjZ0R7zvDpFSPL91tA2EuEjGOSXm6qzczM58ixOAodZdG
Ay0lmPu50MnoHmg0wmBhJPIkOV+K0cnfvJrnDr4qQEPB6oAvEMfPXNQ5061Y2RTzRekVzg8uVFDl
dJSR1tj8+/KtaU/6td4RgyyNs3DLl+vVZHi+8QS/bFdg01no5H1Hfz45w/quPY3BG0kDrqdzo/LA
3+56J+ow+mxnFKl02LHis8xuDMnOL8lrxWiAepEf1D2BssUXk6rV+vgO7mfxVBL/Zt6h6rGQnXf8
VVyNk43CB404PL7arli2TTLB8dBKs6dFOUcftT3QhySNkw1KF0DE2J2ca79laQKyorQOzUa7scCi
wx4lbeb4PK61C5CyTFXTLS8lid/bgjfA2/zLLgz0DXPrTTLkxZxjmvCp33/O9/p6UuQHwjRai+od
xPVFINnhpQ2AinFKX83XVda6bFoW9k3Hzmf1SiA/HVX5G5V3lz0u34BKNfnH+3wiaEW/BSL/3WKs
r+FfzvCbyb9N20YIIs6KTFgEOjuM1EhubYLCbNvUmW2OpjvqHUxf0KnoxKainZQjh0+igZuWT0Mb
2hkHzmR7F3flnr+9qDVq617BJUc7+cKgI9Kox912+TK7c1GE6M4u3umPwslosF/aycDUgOKLuFOU
jyOzXHuP4sHAc+AAlLPOrOAig7Sh7ixxbg8xWunF8rdXl3pEb+Sgiio6NuW3PioXXldMsCgLF3Wj
DC7yEEeRf39zAADH8td6bCOzqBpNVzQxrU+yB/iFRgoOdVBeI9bpYfCQJ+4/u1sZrgaHBGfZWAPr
RwUACouEzTt8+oUYQ8I/w44I4buuOJKvQrGHifiwjGpcNff0h2Qzx2hS+nZc3X7+zt/s/EEmzpAl
h+ReMHm40sV6l/tVdrtt7lsm7RYKsGynCELl7IZPPzoWjQDyf6kJXjLC3sqeQIoP+3PuYkybahHY
sC5zzNCdFJPxtdbT4t/azj9mjcime9Hu/bPe8HxVgSoH1HwOz6TuCUdzbVfw8xWzzjEE8Cq8O7jD
GmhHxy9YnS8yeU8bpzAl8guEYul7rjeUAywvpQT2ShTpG/pFBP4BwMKrhi2vAI5hbZS4ilvz9gFb
QJZEWQC2pZ6owSSwsDfgxu9apLTeH2hdKgpmkIdDwM7R/znyzMVLh+C6lVEM1EaRLrO8CBb3IFLj
kHFsR9+7UtoREAlRsRxI/Fo0q5RYylBGMYY+1KXmfgv+hJG43pywvepA/crf9H1LNkmjdXYdUYbn
lI7fhE8aXcwHwwACJQscW5QrmgTW7qhx35BmK+9BmjgimKmDyZmVQ2xP5DGBZPpzhRNayk+tQ3xH
bLNftfZtRxglPDHNV5pgeNj2x+pKJKlE9P1Uy9bVTWWlEpjnYbGc9e88yacc9nni5KUXd1PdDB+3
FG5g9jNtn9/p5pNWOUl8EZUtpRj9lTdGLpzDAzyYuSJRMiqwwFRThlj/3K6MTTvuXC1rhPurwdH9
7HtSLZQwzIz0+KJlSbyT6TlOqD3eOw458hMeLlihXQnix6oIPSSm4ZUetCJtmdkwCa045WhQWEaX
HBLUD0m0/MUm8NHOJ09MrwJ9nwejk1EGBfHbZ4GC9iNl54DRgc/YJTFjhkmgkB3aXhXVxTOxs8Pi
qg1uAUlnl27YfocU75hZl8OeyJ+vAixqLIslHOTNVcv1isEPpfcs3pgi10uymLCnAkxX0+269phX
3gQxjh6yS/Ebr2ez58mohfr6NKaO0EqvSvKFFAumFngiZBjlK3Bmw+8k3Z/8kojwO6SKwHUCdPpj
J/0eQUmmYPxChlHtnsVHltm5GeSOPXlGuG9vM6Z9eOCD0RkOuTQV8g0GG3ojlGkJIPkrywwsouXX
+iH+Mt+Tt3G3SQz8AnaaRrjA4kF0hfRWzLGhOp6Hsa22f8+6MWOdeCMsxgsEzbvlSxhH51xRN/ko
iAiB9cCUzMrlq7VWQWUmm7wtAWPd5hnEqs5OjRAl2BDMUVMh9sOvsoWlwN835QHittjuwszne1B3
zPxYmItx2sVlT3XJ4jEpr6zls27FiMajNAG9MBiFZc/zxcHjli1CCmS7OgnCN6yDvnTU9/IyYv/n
mS9czWItUVeQHg0q9aSwQF0GQR9c2vU0GTXjugRGP2qCk53i2gzkFFzwt4t9oKQIzK9ru/Jx5WrS
chNSLwXdbY516S+lx8L+U2ce/nhNhu3bSbvVarNx8gB5k5zBQ42sNuOQL9zXvae0IZDIpxUxooSz
TjLqnUKPb/pT78fn0nGhmOzrrudjpZz5ThY6CIQouUtyBtf3JH9IDdQQTRJez+GcesM14pARetjv
NdM5p8cjXRcUSoJ8EhXy6T/KFAumu8hUJxr0xQ4pok0u1JwqG9dZbpwr8TeNvR+03jiq2sf4Ee+A
8Wu2W3juAkBP9vbfUO31gMtaAQHkZjgIcUqhQyTpQk9/rLNqeQjZvFcWdvESrsJ42PemZdlaeVYK
I+Ao9hA3ODQW2JGG1Vqw++aceR8HQz4YuMtvRhesztRBHvXeAeCkCdD0HmiB1pXVlGCONNHo6iea
6/g34moZ3gfhNNj34EaWeA0dEcEA5S7YfVjCIFF+Jfn2823Upo9eWUB59adhw29GMBNuPWcb6HS+
xd8gS2nQKw5Ub0RW8gUil7LDhSpQ0BzpdSJytwWMIytexhW/ma8lo6FXrgW82DS1Oo5mAnRaz69Y
XbfOjKoMyzRoIAmCnuApIGzQWwgMigExuv89i9nxni0zjowtH/mN/jwUJh/dh4nPPFr70fPJe/ra
JNfkmb42rAdYgSswtdUUKGGKyQwO4DjKT9Azq96sCnWeBEtCT0U3QFmgVsMJ2P7UrKw9/gQHlSh8
OnG4DHkKc8AUTaJxpw7ejRxyb/CVVIzZS6cXt3liOqIk1rYWypYkiy67YEB/qrarJGjf6/I15chR
FhUNfHYtWL0hPkt7D5C7fs2uDdterhcz90m0TVKCCTXu4+4q9Tey+khVghb3L6mseeG4zKQFokmM
nvD3UXObTZl+UcYiDj8WwoGdnJOwCzK5tVFNS8sdN/VO3rPs4UotDoSym9HeylxDzAwEbXJW1Be7
VVjq7QD7QOK3d22JXOpqFcXdY4IW7v7ngeGLkcSK2moZo0NDmWFK4VoOEBW1Mgr4Q4FzPTuyXK2E
J24XtLbxjfxVCwzf4gBKM3vhMlIJZ2XAJkEQnl3FEymOEvRBWJtOOjuoJv+Ccjt0tHfXnx/bstYS
TaM4V4d6uS4f0T7vJSwBFA11L6Y5uxVdj0X093wAwkOlcCCS6P/4ONFwfY54d4k/YwGtzWZKjrI/
PFEkmLF8eNks+f0EwBYnVglDMYJLjFxV1NmOypDMvfXldMkDWsqSDfsCOrGUP9omEUb/g4Hs5eCJ
s/k/D5Ux6KYGruTLIinpWfiCgyEOnjTXL9qtfQTVjYdaHNdYmaDUZkTkY+HJaHBPXzfk2Zt6eaxI
J4NKSl5jNIsgLAvvygdbwB+JZRss4nsNTO6ZW2iddB96WqRNPsuHtcfL7G2HD3xoWM/LEcKDCHVH
JwLiylBRbS/Cnw6sWzgNGaSYHJmoINV/rmrrcGTeuICKPPru024f/723uMEnv/kWHeC3LP3YgL2D
BZaomp1PhctFEU2FVezHUD++1/lkrWl6/rEqEukvatIryeIujh8Q0Snu+KFU2u3/JT88ZGVgStPF
QeDBiPNU9+akej6CVssjRzspdJLGOxdRy7GuoO73GUyPG6tMH5Lq/vPXcjY05Frs6JPtjlw2hfpO
poK25h2WZTmijlg4QXduvBSdgOv00VDcSobclLrw3l0tN94En3+JQ751f1rdIL46TNphukwBOQjw
zMoiXb25OwEk9BppwIiO/9r36ytfJAt474i4OPK0WcLegOVhKAmA+LCY99Gz/B/mRNtBOo+/OMFz
PNNVajF8kuMeRU/V6NB/dESMfdRt65QaV7xdPUpGn4AaaGLi3XtoX52fV74Lx/VbdlAEcboTCaK9
YKNMdjGffFyb5f6Da+/v2N48QrkKVCEWsFIZHPJx3KhIf8kKYjIRRh4mgHlkKBFUnPA+4VvScfFw
02EsBOx1U0uOBWSdRVLz1q4iRbNJIkCMuBV4paxdkSHu4c4yUk6xfngLeGX9gR8BBO4bL9TImx6b
DCRlRVyPwW4b1Br/M1PAnZ/K2ohweeIJe48OneT45/0FeUGGlPU5BK9fgWJMyebxhOcbrMH++zRx
Eay6YK6Xr+SxgwUwHvTVp/lE/fAuFzqyh8k5F1eWW+849B4KUP9pt5bYNROIu7KOO6PvwwGObQVt
QWUU+HhVFSxC7MydZ+bhQzdpsk2+bmhmfpdF0ICm62fUShLgBICW2AYFey7ug1EoViSicfNk6MpW
ftYdhO6oqfMvbO527lmCW2jr+jskCX5QUqc9B/JCJ8hXh7d0TA7sK4ZXuQQFHQ8AbDxhH7J72BlY
yGgHh74DyMVPYXZoYxtjIRre0BLoWSQHyDivqcA9zi2w25CK1jA3BksWC0CA0AMc6L3YU/1nDpOF
aMWQIfe0Vhn6sdVck/h3LAa/53RUdyV3lTTXIWhU+Am8iJ55flpjnFcc8sVcP/WPfyX5vyRe7Fcq
lNUJr0nERGe0JOqR1HjbLcs/BQH7SFzl72bNtorA07N5NALUd8s8yB/6bktEnVXWGcc3LRKC1jcR
F7u5d6Kh4NP06nOFMwQG0txsswJG73RNELEV2yNklDbEMP91MdZeaCy3rAgIhAPuARUdnONZhzIn
rpLMpkzAdkcIOQW6dldTuZOUGN4UiieLZBNTPA073aLmJFpekXeuG4dvQSHWr1FB/jplrabxChjC
iCRr7vNdrCbPsB5FTzNqz95WvSffBVfh8gllGIz05A9J28MJnTuVATcqwEnxj8j+/QS/U2nFOpVR
/rA8hce3+8srH8wX09MNZHo1CkJl4rxK3K6+83w5pxxERSqjG45uQdAIx5Tj1rswMXLonhHuQbAL
Wk6FjJF/TemNWEW7psYl5Wlk5vbce06qYUsmJMQ1dDN2R1DYMwb3ojV0IwUVY37noZtmH4LoMG2x
adX8SsnO/11Bd0ho2/aqR+kF376M8fDQchCjk0ezGidU6ZOMPX9+YEH87HU+8fltYsDQz2Ba3DVw
AIzcBVXGRdqFzibZZU8/nnC9n3Z3WsQFetClEqvRJH3EPBH3Pj4//MGjL5wAvJRf4149xeASFVBx
LFXjgZPptHhxUoZ3QNuUDEI57bF7E1Wt+WAVQsFAJEECK8+vHsFpMTFE+g8lHUIkN4YkrGW45Pqr
BREQByR14jV45jvKzMC1yorSisPpYogkXCPnKoZO/NdYsHP2c2mzGJ8/yhrqZnnyzpqc0UNUqRVm
UtFc8+ylqg1Ldqj/n5DoWkZRpIQS3FZKhQl77Z2WW8aa5UvIdGDxsQ0ZBRxjf+EJwqujzsRdXBeL
IZ2M0sjtwpw/clN//MRF33Aq/BgX/cncgleLZWaw+06VqU/hxKRtYTwx8R7g6RsdvVnwBXQO8NC0
Z9BuZvfipAYel+g7b4OUIyJrZ5ok0K9CaGNXjXDhX1aJLjVjfAcU/gun8DXgH5fNUwbVkHV/+Djn
EVhQWmyAZXYuwzrQ97EDer3VddbMGCCtDTvEX/oPEAM/WA8eWX7oWVP10Rmr4vV0nRlxvigzmEg6
5fa5XCpzFMrpjP1bVP+LxQw6jvpdWqgIMTZPYstHAD9mja+RBB+4XXEQNVK2SyhdLvLg8DXl5zYR
uwlCfyDlaPg6Kd1aIKzAv2tSdFZ3k48pKTcbUsnWBIuq4FRZZLiJqKtrwZLScP4d1zjPKP9vS16z
4TATEUJoKftyxC1avkIJKDgM/PlYyimzDOjzulYwroujLO4es4jFYU/qJoMF/B4HHE4Orlaeovv9
/W9tX9sDeXW/BazlmpY60e1/uKVNdK+s0EBlYG9lJE0CWSvBBagbFhcKB+Iw22h5Og2CurEOksPr
rkMAfknkvrpKRS5DxQ8OO8A6bcHjOAHsVTxMVXlMg9gB4qyyl6AVqJxouOhc605L6MCCdJ8QvuZs
ob/6ME5r/H+9M+Z+1wjiWzXonnfQXogV/LEW1qejD8Z9K2fhuQbh1v4l8SiIN7gQX1i6Nmxj3hOp
oOEvMWKgIPW82dj537j33/Du6iIQarxv3IhZpeJ01aE44HoeWes6xGFtV32YQjpSQ/AWIMZ6VwzX
XNm4TbjKOpQsQK9puXOEFC4oHra9mR7pUPs+yjDs+TPK4B0+94AOQpzTvkF/eJw0UNrOX7GuuczF
0i26yZdxhkp/uLJHAgcZ7lFgJd2tWNUO0xDw8++Ee2Mf7rBYWqNOtwZrM/bGGFtPwXuTqc+EEmZ9
CesVR10WQAaNerGIDiFj8R6+Wrs3rx/Vnn/jbBE1jmQZqaSJ5UxhrKH2aCaXOjIYWPrFU9nGur1p
Q6GA8wepQxzXU4bY8ihW8eoeGv6/w8BQetinv7IW/3xJXYUrT/gtZX6WbQsJsmfhF4L6DHnatIry
PxWFQVSNja1vM595CmLdYOqtwNLlNz7d+9Gvx34UROAh86AP81If3beEmjbMqka7EpKsBfbjl9lD
Xv8u52XmmtW/jgRaflH3CuyLWeJcMRqzGEWPyy57VkHLLyFIcRgqLSS+DcLAiftanKj4HTJarWC3
QMazYw99od+LEdtpkaBMq5C5eepl1zFck5Dway9rHN8cS/sy2WPkXDP+m54ce3Srl+uJd2B6yPek
EGSUmTAsQ908cOEqXBDXLVSZ2F2qWQNm9/Rdv9/NL+ds1xfUsVu3Q/q2UE/vye6dlbaE6shecY5K
2OyTVb2srq0l4K6V/sIgWMiQ7KvYKANaP5vEog3Kb/kpjhq1h5HXn1LRhWsuhhbjEzf+nDv1J/er
jr8ACddRnmdFvcCO4zHquqSoogdahoRBcBFE41fRo1eENML9leMzEAazkmfqEuB9NQCBJuKFvuBI
TThszT/Ev8/UKUo0bbh3OydLCsmgcxqOUzY3w5hN04kxewWhttb2NEamtSLOQpwWywW38imNDdsO
PPdGHM6PZhHMCMe8rEdprq7lQKcmAKI5Bl5tv00Al9GL2jO7y8AdIXbGeSYkPzBeMmwDclTH/p+h
NLgkw+sr0r+efJNzb/KUAYuReuW6vvAJoc68FNdMbzvLTt1GN1zLF/Qezdczk6J0hFTKynfmKJo5
j3l4W5P02W9yRtbX30jiHLOm10zChM0mvpwCEP/gS2YqyT4ZhhrOeYSrm12uhY7NMPX2+oi45WUH
O9ddd40l4weNZPPQA/yEpEQ0ZoxivXI6XC3U3onsgcf2bi3bUOuMskm+CgnFHU91ZbhxCKTP2gV3
u0aApaxp/r6Qn0YF2pHLEQHpRUhmjgmTi+fAqGDq/+bMQFZuiL8uldCvXn3yAVO3FUucqt52O3Tx
7jfI+THcxMNYswrqQv1H6sDFQTJd9G4kAB+o0alq0chAnGZoYM/kXnwpYwho0YbEDAK0zzsYjetP
uK7510WZgnLTP1ZLFAJPJAivy1BwWNUnZhOsT7F3uvI95EdX/UO/mUV33BBNnmw64yAZ1HDViqds
trePyPLR5t0KibbUg1zaTjXiOQJG1Dz/p+OnT5+/J/OWZ5d+BhQ5oCTAL5RDSGt0bB5e3x3PDtq0
3UrJtp+AfIw7gUU7E2VHrCC/y9E02qrTPQzY/jqBDG7D8iOGY1m54f8MO2ujhYCK+M69cbebiock
1umyWpIe0eAFqD0hj8kOuiagy8V3kQwNrAoBcfrGNCsZJ43NTBXeI8d43QJQVVnMYX7e+gN63ni0
d9tEhQ+e3z+92cNrFf79oJu1nMbH7nsiUy1+Rxsh4l6/dC+mc7dwF+IE/tcokVDqMrOvgAZ7ZmNw
FmWDtE/lvJqWvlF3lhgaGz/EzUAHmlet5kWiekIyf1rTU0INtSVgnhH2351Olif2RM+o5Qv5Cu3u
/HyDlxSgl2rVdt3/UkJMiEfOFsQ9rswtmy2H9bfiTAmyM5bkdSjBgVXxk+MT3qHi1sRO5MvMLRgH
PEUOz1KqdkqjATZDp7l5G8AM+dOKneUbMlCEYv+xsYqAQCLjGoYGhQ6loLr7OU5u/gR0ECnPr/80
aTrM3/Nt+Zbd3IQGktDPP+LQfremo5Fzm+ljG4NmUT6ztf56uyKnSggrM8ay+0zVQOE1EiveWR0v
xiRdkX3gGBe9YaHSZ6cUOmRejtEPTRZX8Khc5k2LCAm10DNrhQmtA3IxfMRfq7CTFCsG3fp4XFAb
g0Ft414mH/EnCypfA012howrFltWdBli93OnDjBB7ABINlwePjJO/v65F6oUDsbmdwZdffb7NgiF
D5d3QjPUooOoC/6C4pOZyJj1NE1H0tLtBO+SDI80irUGuws/TFEhxZMGDJjhcK26UUxxG3oQk09r
V8SdSMybzypsZ5wraD3Gx9p6dXGNIflFyxo0WJa4ho/3kHUubhi8ZvKhBmttXIUpGTqYD2IM1xc9
6VVIdEsr+D6JVLy1etgq/7TBQI7rcB9kNXjKc14wDJRGvVxMgce2CbO7bbcP6XTeS3TZguh15575
Q+8jewKHbn3aLfsKQYewcWY1Sbk4sMiBXU1T7/ReJZWBSJRD5pCGbJplBMRkwoO77r6sOEO80GSN
B8lrA8z0aRXY0STy3norhxKFhQZ1V6+suuibpsEToM9zKYAhY2/uBlChZlqf/D4QKEceroIvXkan
RIdQtgDxc/EqBtGOihGT5csvAlxoCSXspKSZ9/PI8ht/KGOnMqGZWmadQ52wVFE6+YIuh17QQAZy
O6s3zIPG/51Au4HNIVPEsliqJYpUbhfZcEyBRSfZdO01WgHtzEgBKxQO/a7xh3Et3Vz19VR6oqKy
r4ZP+CnFub2UgrwvygHw+ltu9+4812OuA03fNkauHnpeF+ypPo+rvIVmYAMHsbgpdRZFG022lxZn
n/nAKzDqNL5V2ioJnhYYElED5BOy/NhqVAP58YWdaEV7JnNyTqWhI5Rbb722/yDzoe2KdWwmgywy
MQFljEOOtDgqHv2j5xGo6g8nJ5uhPL6u5dCqTB6JVI7xeuym39LToRvvgWxSVDjfs11iCoViCYnm
MvM/JRNtzumImqhWfNxLd6tBN9ErVIeVQRVQRuVnsnOPVcWUe7bqRuX018zEVPttlm2iCp7t7khT
Gug6F//2pVYv8etEIBfOlepiY4kxYbQEwiMUaProCinGqJkGNrqQ0jzwO9X4/j4usgrC5KhJoNdX
mtxPT7TrhcRxJ3PqA1i0icuGL6DQUpVyLsAw6zUocbut20pqzdjcDitP8Sf2DbxMn9PVfgWema4A
09ZGCcYcY/rS6Wlh0ZwhNDCpAnAZFhYl6GD7n/+7bSHBC8KxJeRl2SC5BHceG3iR/8M9Sg8gTkf4
FWIVYgPHNyPRnas1M9D12G4+W74tCmMScn+HkBHUjia0St0UX+HJ9NOup0aR8uN+YlpjXyiKL+7p
/E9yzHf4h7MG3kkeoMx+mfMPI3OIOWZMsbk1FHEJMbDOr8+ot3tc0FHMpCZVwqBjSVVAvURzgPXZ
eff5fLsHIdGXgSnsicxs8ozfCFh/yizX7wx7DKHHUsQKKCfHZF41YAwNCRWrcWILQgHfwwtok8xb
FwM+uWWt7+hry6XmgOS1u4RCYB16/pCbNZysd4QZkXqDODlzrkxPOzQem8U446xjJBFQF/n1FpMG
PFHbN3d378FVFye4WRBAFi3eEAIZjk/YKHW+ijV/4vArFhxnTUR/G32meZla4f2aidgVhVrlW8BX
XlX4Iy4mkBEIe1pipzh+UKPbtuzIwWJ1/0AZc5nCV8iTMlEHuXQo1i2uQbHeaIot/c5P4/41cVSS
7ehwdSnO5DvXxTctiDyW4Xo+tdAxhfo2Aa4CCLuh766bklpEtuyrWJHe08BFQlcs8dA7Nzllcc8l
P3sBakSxib+46F711QG1vv1KSkGS1FXlC6y+9AGmxHrTO1gla9ckahX6wvaB11tPgo7/uH3mrY5L
FruF0DUn/xB21Wu6W0dTYOatUgneYoYYRd+44KubrbyJP5Qq8XD8GCtMTlv/zOPcJ4Jzg7YyG4Mq
9GAzGxM5wR6p5sCFyLfbRo93DADnzE20QLQeK7H7kJT/JGmaMF+TlXXbUxIi19IhvvcQvDstivC2
v1KJiL32hwdsHmdoDroizOYJ7PIBIO8ZouU3FuCtL6zpem25tQdNbeLQOuM9XOBPo++eqDBepWJD
HjOCrYbDb8aLtNV2Pg2fOlvzm9U3tuykLsqwH7HwEM/7wjTxXvqxmiH98fM2MiMX6A0TdWorXfj3
YYW2s7SZaaFr4Zmj4KBcm9HTi2vO/oqrq7H1bFc2zIaKgT4h6MshAuI2KyL2i8KUjPaT79fgHnRw
SlQiCYFX7LiJ7wIVgWLXzFboOme2KiSXkW4GYfE29lOgrwlxPl8Q00KrfVZwAXztKc0LTMLtfqwp
Ux6Bnqo0PyKAWpOjpd5R+c1MNCvlD+aEBwJk+HddJFcFp76dG/hwvxKCCLvK1z/LXhs4K6XrAoWz
bykj0XvPE8LhUxxchxjJpdg/0w1mHawXHDXmrDddk1MCedCwr2UKfQJlf3gBr72Q7wXu5IJGsd1x
cqsfPonYqjGg3NvLY39Fvso36jHF2JthhnsLjAr8WDBm29LkHfGUsA/ZIxTsdvNCOM1CNB+mADPW
USD7WU+bv0YfSlgD2D5rTXxH/W5n3aS+C+OD+LU61+z4LWFafRUo/e50MumSE5lWtKQRBX5Q7IE2
oPE0Qugi99YNEgTK9pcnaE0X1FWcoCM4v8Xo13HXPgeXSIsh0Kw30KOd0N6xQ5ScCbmR9w1oAiPJ
pfpxizN8R5Cq5DgcT73E7gLtbA1FUJaTSFenOEZBzgmqsMA9GM1DL55oVS135/lc+L7CdaVrZsja
OKpVuFQcCi3PF7p2nfD+iRkKcS6XbfJe4bKEQmIaa9ENBsTuazHb9/X2VmRwskuJWqrceS4Gh83P
6fHIcTtbviNlcCtNOOLCPhxzS9gNAVCMgBwD22uuZcPNT4pon0ziVqXN9kNexrABT9hCJ5dfsr8i
fzPUPSNaI0FLT7zBtXUbmYna7xf6Qsisu12WEFkrQVyPV9zJFiKD1hYXOmosDyexAs3OWy9QGMTj
qy6fgtL/kSN/bNgG6aiJNMONW0TLfTofysBWwcxbYhwtA+BdJwa+FfXCc7yj1DNgrcyH49kZTIuN
A+iDETv/raxGr51QkInPVHsa/JUtzV57bou+uIkxgBkOR6+oesP04YQgaC4s1EI82nfWodbonOmG
EbgK4uzFlAip6QuGVzaWkTWImNPYH0PLe+mkcBf0KfbcgTiolvRfdOSKEwvxJlONuZYRKiP3QRdB
HTRTBZdZxEA5ALJCRX096KP3TyF3uu+gtRzXk4Q7NeO184gk/bFVMq/BVpDysQKFSNE8ycSJWRoX
w1JypShhuVfu22SoWDuwV9l440qJsl+id4tOo7ggNIsVJwidHquUmj94OKuPRZeufOtDm9bGlnOH
SGFf2i1Xn18EyutdRKUHEUsjrzPZLCXV4vNy51M2+buWgI6CqbbvxlwK6ScN2LBh3BFuIxfYlFPQ
7ROwsu8H8+1mixSQQI1E1AJvaBI0EnncCBL0ueYwZiVnNTjuRysEaw9Dx6kHpgYD7rab4BEu+85e
MU3xduJw2ifP5KBfC+X1ghnyYTUn7BOaIiG9nhclymY8hL/MLaH0uIz6hfQhYWsf4dBl8aVlNp98
+NHgN7javyNOsS7xkfaqoIPUSjqoYqQ7hVb3THpDRgj7zNAQGIUAZPGUXpfTDUXK6bTlzZtJjWKs
ewUWkQ2+lG4+uQ/5CdDKDdAfO6AZZ2clZkkcUQRrpndNlHXKJddyd67W3ASJ0K/LIHTdvOstxWMf
WxcRZl2seBK08Cr6+YDco2D+JpnQ7m4SkxbxTBH+pAlrpFtvrZg2U6bVXuXbOxJU6I3OyY6TvoSq
wi/azu/TXePphuu5BaFI2JNrO9wLeHTJWS6eyZga8d4ChA14pvZxXtTHKHIKctchkJ93MVvOuSXX
IH0ztNovk8vQuYpb87bGDMCUB9KlgIK27+8lNZVtFsJQRr+wlcce5bPWLiA9d32Q8+NkEzA2Qb9Z
nIKgYklueHJETX6HfHYRojbIYnLvqLHOzwmZHO+p9328zONCoyCTz1zXXvSWTRWbogH8nFLpC6rq
m/voMUe9/IbAkZftJRDs6gNV8hHvJwlFl716JUhXHsXEJficj3KqYSCcQvAesnPK6ZiK5FsDzcRX
C4hU1/ya3m9rVIUQ2BWCb8QYlnTPZA3UrKl2W4EN0fd+0Q7/HS3UIgQG2Zl0PTneSYmev3epA/mS
0f17bjANk4LHjLVBUrssVTkZuP0kL9rEF1q+tR2/ssSH7emBb4FfOFTmXLAu71QVXXcF0qzMm1h7
L19pNSZxrtzAxjvWe8YxroNL3QzddggI8CXdt44/3xb/9PFvvZo7PXHuRAPVabaUPzuhtB7tKCOQ
8KOILBFgtG1vwFC5wD9XWWiXil/YHfeRi2g9uQQv7U/aGr/EjiVUbLngzqAt4C1HnOzQvakswQmV
6tF3XbyuTtYetJF4zaMoBmYELQkUm4cmAYE69/JsEZCJ6/6R5sl81+znwEpxLWTDfRG+PBZxb/jp
NrvommTdTzboZ7D8iowuuaulmP4ipZ4Fb2FLSUweNotyTzF1oEck6LASb6i7vMHG24QqYkkMllEQ
tYL6Bl4ifeRqZSxgRl40XYh9TQBMCHoRrMK7dh9asOiqlfDFXMb68EseogQGNqn8+9Oxio9CQnvl
rIPZYfvZ4xDegHenlc/1iSCKDGh8UrvChidlU8cYHHLNXM5xx1VWIb9ECdQmtErPpjlsDrw8L5xv
kaxtXT//RfaK7vy/mjIyTB7HRPkW1Y5SHlViJ+8F3p4y93rxb3CKOQAtfI0tuLpNfkE0Flah1GaA
i/Aml5OAoOldE8Phq3ohq0wrAH4soglT0lLWE+k7EijqvKqSkveAK3jQfohxYjEnHsNWus9RckKt
hLG9ohIeMZhT4Fc2NTbQNdhfaLmfVguY/1XWkOyZqpJgAspGMoAEpHjYHY82I9Bgk/O1Dct1KHro
3X/xf8U6pk29Y995il7QMHx08zl4Gp6aGZ2/fH05CKxI/D8dwe44DDx3UyM0IqO8fNDRo19KoOJI
zQqukt6rdh+mak/8CDcaio26NcJdSlODa7f27Lj3vrB7ni9sxUFuSwLUG1Pk7alYSj8fPVGwuy8y
Nq0+1lEdG2ViUcEsIwJqW6aw/lpB9W4Iy01ocJ8b05ltnuhUmgj1G0juwa2vm20hLfacyuDTK7s3
OQlSs6ldAkouHc2G/P6BZKWx8R+E6EfS62ms/JD/sPtBUyrOjt5jjkgsWIGTQ0NJgXByiIrV7cPs
K6IT5cm+L1zzpcneS7XRjecUXvh/Of1TCuVuC+nKI0XijTytpee8G8JhgussF2EtmNcOtgMSk0Z4
IUE6eTczDu0XDPlYhqHJMVDolMt15BkSu4xdKf7WlDgifg65ZyjYHs7rRdGmoSheWy6gHn5Zy8nx
y2mrB434UmmD0PBhrQ1/IIDwnOML84Z1xOhgGeEzZuC5qdfBQqmnC1Zf6d0/C0mfdTNdw0T6u+2p
89sAxpZvVvnv9vH8dZuqeViwkv7icQrqeYbI5ZvECJS9pzUwTd2n+Eb5ZRmQp7et4N4wz/jUQNws
/POKFSMFaL+Pt5o5K6aWmCbQ2oQcabCpi5mHAnjBCeL3vnr9SzxncaCP4fWPhhEsdQ1+Z8TqwMUR
n98kQY2BZpaif9xfAeqZE8ZyhpP/Zwm4dZ2qtdCz/r+An60o7yYWScO2shVMEDATFKrXjvZz2R95
P7247mljnR7+rjrGzm50CM1Zy4YIZHUNQOsns1alzNsRwDHo9DC3Qz6HzipicqVWIXQs38PZFBJo
WalJE1+SSxsZxVSax1polfPZ4yZsHvMBWa0pTJ+3jCDeZT9BgX9KcyMJXDdxW4hIw1Uc6TGPCpUW
NnHP5yDcfP81ouUUyV/Fie4wUARSOwe9VnhFMtXSAO0sYCBbEhidAX2blyTJpJh9s3XSPd6SPQhn
L1uj9uc+GP/hjInvXzlCz9o5tG+GW6N4q58tiQmWnWXXSl4RGWQnkgx55+8ISO43CN8/RTwJP3+t
0HUosDKkIwIB0d2ihhrDnJygYlvNHM+02i+zkLWDI3JmHuQcD6bSAcVVp93u1lrCGgJ6BSjmd8mD
D2oCFAAIFYQ8JvcgQFxOMgv20TzYwkF+36MdmOxzuMhlij7IO8X8F0kRmhkU+7LjU59lx89pVs/p
kjKsJy12qOM+exy+PpI5Ik2CNg6I+w80qf3s1aayzQ/BIzxa58L+qVR5YkokbsCtN2AWhK1RS58U
EG8U0m8UjPoRRTOc02AxKcFJkszk28LqHF+E2zAHyv+bnb47FN1Pv2+BIjG18a/zbWl851MqUW+X
DVEILgTHkMeVYpTFUeOg63OamLQvqR83aGEjl5tyilceINRoEylDFdNqZUgsuyFE1WHGGMSKCWH+
jXOcqSO5Ogyei+VINT/atpDMXxe0CB8p27BXqujvWtDZJnUPfWfSrVMj/RJ59eTuhpzMebkSjRfv
I6JN2r2Jfhva4VQw2qWL6FtSBAQCNJS+7t5PL9jwDHirIcyeAqgk119kpe+ayvqP/uZhPmO8d3ga
Htzg8Vf54ugxDSUslSgJWfrG2Qs1tqWVvHuyxjYG3ETKW+XJnkC6K1d92hGdTIEqnb6HmZfp3GeV
XExMn2J/oxlrTxzIPzezZWheSYimiKcLl4OQe5VERQexV/p7xWp/LhUiLk1XOTmBw7oRYNC61Ahf
jVIwe/AdiZxIcMJEj8GLubyI3/eas6XxA3xkJvjKcN8mwmUVRDoWgzVlqRFtnp8jiKaPv3nOQrFE
8ecgB6Z7ColN+P4rtbcWqsZ0l0I9xRUnsFlpHEPaaaQ9C2VPKgJ+xtY2hnZ9s/WyIVK3G7n+Pxtg
BaTUvr2Yst0ss7EggosweyRCfenO6fSt9Y6cAiBS0Ae2Q0yX25mNUQpOIhUY6XTfSjv+nD3ClCw6
L9aV2omw/k826jora8OlGtd3tajSIBogrdEL6DiHcExOl4QgWuCwYw1x7ptUJtisCsDMnrVYirLl
WybDxXOXcpTx4Wjg6pqLwH4BduFUPbwFKvLsjNqqGAJse1+PhkhVbePOtc+e9Vs9E9DblpSRzTci
Q7PhwJVTHGQe7DPf30mfnBtleGDHHB3qBxRW3oNvam9l6JdG8or0WLQjMy+VxU868CjTXtKt3+ra
/Abt+2gtxdoXft1+3/0ZViZ9fUsaZ0E3RvNV3fvE6m8gquH3a2KtEhhOKGHqVpk4+yxKJFdU1Hj2
sXkh7SWbJ+ow+ZwjKsP8IHC1VQIKMQdgP/A3+JYxVsF6QYEx8E8qDvORpBH0BHpPf7ZQC720oBg9
g4oNaedwMDVGvMuMlOg1kBrobmsOzuitLOHpuiDXsR3XsPBxrtm0ugslAl7MJHn3RbCL20jSb59o
qmoEhXMR4UGJor/o4WsjhOdPjIFybKmP2ap/UrfnW9jtTKvsHRVWr8lSPSskVOk2lJZGEoS2/v8A
5bmTrufDfwFFO/khJhCAm30ZodHdpMRSo+C+UjOUTbNg3sj4LwIuYM2ou/dK/5JXtXJQubZKhaPI
2WgRX8zI4VvGrAYztK5DCd72nufUg2LyUrnqTA5cvdkMXYuvKa4zLj1bvaHc9+otrFG0H1OKpRXL
mzAsZlq/tElN0R55ZPgVyqWHX1VdGV9DYYraqmIagrmzSW+Elr0/F9ltO/Ju6nflTqwb0GYG3dD+
cOxS1vTwon50W9f2u2Q/KY3KdwVL7pPvKPAVPKBeny6drUyKiElDhd+et4YHQLF0bzD88Is5NDma
oNMR70J/89zezw/rsYyfr8HC1G+6nuTZIxYAjIoI51lphuHvVq3Aicft/9T2uHtDC1cMTqD7Yry2
f7ThezXQeGatBO2COEqLHqcVDeOFvrmMiKIBftQmMWcQPrYV2W3japfRXM05x5HUb1PeX8pzXnxT
AyVteFIMz+pJbxf0Tf3Ec6x4npMYYpF6kEG/JHzd2lxYE3lS5uNK8Ici/8Rw93zZoq1kolJAnTPu
vBYJg0SNXeXfNd2zpGWHVC3KBCfMfMpAHXkRo2OXADBNJosTxcnVrQ9nunDNNO9SbMZo990XtMYL
XBJL5he0yCUUv6tnxB4GBttWOi6FjDkJZZAagE5jUQKpCw+Lr1ZBKmSC9Y031H2x75u4ueefk38n
5ObQj5yGY00et8wZ0wt5xjOPm6gErXwCKQx3SppmHnRGRWMxG/AHctFcWps9R3brVuvIeaSchtt9
mMQBqQpK5PwXxbd+IIZ6+Ag4ctSWLNR3Ioi04vo4hdCOZMKONYGtq74/9X/wC9ULr0cHEKMgdV2B
M90qsf1lmWPptnwbRWhQ83i4HRdbXjmj47tlnbJ+s911ptYPzFVPmDDpl5licWlK2TgRPnxlB4TH
BN9Qaccd3MDxRXxo1l+UGbVS+d2MozkQJ+xxOcNDCA+pgq5KgUiMuXH+EYvONvFXg4P/5nP6poMg
IQ87LVMdDEdV3si0j6Spd02zRhiwCEoz/V+jmXqFTrOWXq4VUUQ5gi04h1bxqwA+lbtGqYG5Y+pO
WaHTNiEsOX4bYe6WMGPf6tqtRXAjm+Jie8Gm4IZQVmOb8IO6VTWm7rpbTEdlv6g+rMERumjC7bZ7
aEo3DRqR/UXmCsQ67eou9iqMsQjnd3zTqYIPE/zWvZCdIfYBDhsxWQ2lwUL6j1a+zeaf1StYaA05
1dfy7gWM/VZ+inmFRSZlF+65lV5A5hvrqx0Qm48UGvFRom9OR1KJC8rHQ3WGEdGkRxq6ARes4rzP
UeFmZtxVLqgcEEd9Gqm5Lw+DOelOgM/alRAebdP6XrTAb3i5sUOH6puT3nGRgBeBedX6KikaMi/q
WSh2o93FYTJBg3yI7yJHwinqhp9tgunTXp/TstXVus+X/disZ1KUucU0ZbB1NGePDyJACw8hEzyt
jZdlgG4HJtGpy2aR2yLY+DCL0oKTkDiH+PMEXcYAiFcv2I77ggXP+HGHHRKJntljCH3jOwuUZi09
rEbQMp3u/2X42mRVjbMv6dxBbK9fJTyYoj3pti85Q6DDDaA+JlYw7n+4YsFq3eCmwaxaolL/uEIo
3eqP8tfRLok90Kk219lkdh4Iff833/wY8L1+3KLdtnVM3XhZ0VgQX4vhwW7OHRuEc2a+4oMBcXUo
9WnaUE+i3B7V1roCX3nXrZNsjZ657Lwk+QkmxbUgV4f/VpYGC05NHJzxIvofDugkJqCYPC482z7p
5/3yCrKajWY0i9co4WskXwDUnPUBL2m3feTtA3S79SWE/S3Z26IePkgsVKawF+gNpflTi/GSQsDJ
Owe062WqeUMhSYB3BVJItLWS9a3YEC/z63HcEJXW/ZmMQRQSRDnkgT7GzIBrjlHG2xxSrvfneeld
HblvYFOfnw45rfxHv7TEmWL8kwBii3v/eZnn9FFH+TnjATVK2Dd5IkLdtXUfofn/vZkpN7PCFWoX
sX8pVTkAeSYSlDr0apIBlWyjlKs6b5As3C9YtsMw7708AuJ7mc0oFPPqMSu0tfTFJxuxdURGe1P6
sh3qcv0GxjyBH+AMPAhZuHhT2iayQ1LN7ls7hTLxfcqTr8gfHIgTiilJ/ASXd3vn0lJY5VEh314w
s6ygi41nBM2V4Ao80fIjT2Ui+yV3FA1v4HX5rIm4hbtp+0Hsb5i2AKIjM5UF+0kkmIyzyZl+b4em
yWKk4JiJDjVdkr8zQVZ9N8Y25cwtyuSukBv4T/P80/5NNYikRclTvaiduk34klOAzPDM8GoUQdbY
q8wpDKe4CxZyquQW1Ar9I+/nT5E2FbNg+MgOEQktO4L3r31sAiy44OYUu+1hdCXuimlrz7gTKN25
brHETGcDlDnTEp6dzTNkSKdBXIW9JvPRiAOphPbRfgxqikHZI9nanmFm1dvq2zrsHhaqVBfZDXQp
s/lYJPUERFyHAFe/75/EC139mWOdhpM2H+m1xM9flLOyV0FBVRSP3BJwQkRGX9v1b8QW8UxYtJGK
ciREMm9ISCB4g6CLqojdCzKk9WSWdKT+7Eax60+UoYWh0VLSGIwITZmD6GCUc1fqluo9UqtPWqrg
l0lq8/jCZNckNOzj5OaeZqS8gH/iJM1J1gr7re9TvUIiq65Rt8QStyuxJWvqtFowmHzVq9kZPKSR
7oqvTN/NHsu8gUMsI4SEbZHdFYnchSEi10WedIHq7kKm6pfrONZij6ia4no4IVWrRuEbUatsQ0o4
+u1Te7Ktc4ULShPyik01r87KGJ4TV2ZOSjyXoFh+V0+2QIxSrTvqQmQmXAA/5oqJctnc/5kuzUAd
/JVm8MD52PZRu5fMkjeTVfxhSiYtb8qCO9jliu9lvrpcUBwplWNsQt/Jt9Sr/PxKMrzy8a5ZNuwT
WsACtXKZHqaPicszXYpSTAvPKD0r2fvcUthCML/znBI4HKAkYNLY5ErCiOXhBWr8D0So0bnEJJHP
mdAz0n89rrbPZWRdLj+mnLPZZumrGo4wvp7Qt3X6C1iHkZGchv2WHHxymH7melSvvrI+Kz7JKqq0
I+8ZUF/Tj9l0YG8DI8L4V+QALf/gKW/eZSyvmpiXDwzxfDlbOFnQOFmXwRKKW46xurFOpiAIDVOU
jXSX3Hn89b0clbCke1DhjUy6uS+fETpHkJfheYtmHAWt+K27dqJShoCDjy7L8QF2lTjeZK1bQVmu
ctdYVoRHSYa6CzFcoEipvcPjQP1Mi7GE6FwD6Z5WxHUXuUYaPnsF3UCCex/9ql2imEe4SiJu+a4h
A0qVF/Qm4YtZjhmPP/DptJNHQlLLbtF62Sn5J3BTreOD0smmUx82titm/ZLPkRoC8uxR6sfCIDqi
Ip97ubNz5vNJg54VKo4uvwYVHt8v+z9Xl57SyWW+CsU+JHMwWmw0WPG6xG9gLlsOxwVN4gKsA4/F
K2BbtseOH7VTUT8h+SCg5/gOa97z8GUoU9uw/anTm4/MGkEOL4q4Fj8avejq8GgNC/vYEH0RvEjK
5IfyQgUz5c9FfBXufhdltDj3zvkoZJ+B2zTRdf21h9sd1Pe8BQXOsO6oorw3p0hrq6gXFsvhJDIo
l3zhJC3XAMeOcn8rwaBc9qGmixB3M++uHuTQFsLrb3Q8NmjqzSuf5lwQSzcOp3h7QHdbbKfYaGQA
Kt9Xp7V3ft1QaTxoCy8wsvs+dEriuHLBmE63CzWq+5ce2AnhIDIbCbW/O4zprlCMQpLZa6DX7JTl
FlUcLcYrRN7Cmp5IBKYseRGAOq9+r5i4GcHZkl26bI9q7wAgv/Yqa3P+0dlxcfp7VEhYNRxuN9G9
FpCVnL/IaGtjVgnZrgLJ6DbVEYaXnzddhRSCYqUFw+u7tI3u6NByTxhzL5tRyFv9VRjN/BnojDGi
R5ub/B/axD2jpcrmhcTMwX7y/B17xCGZslutU3KNuXH8WNv8gE+ThUg1ubw7nBZCfHWslGWQ2+Lm
itVkL+dThJ54CHj4Az+syUfCKOgZzgB9iQ8pTFOMU4S7FUxKkeiHI6ZCrTz1x6lisJ883vHL0fkc
4s9gxwxSa+NrK+K+evKKE/ofrsWIBvGxWaKP4PdRj4Omk7Bp9L+VxnRDCmj17HW5yJngJesogTex
+0wrQwMSI5OcJ5WfA9BYP0npY1gx1Kdj9X/xSGJAfrcrY+KCuAsnmAhENigbcrRAoryM0G7ezBZy
FQHsyVt/AQtxkykDpWtapBL/2gVcuzAG8b1vXyIngdB8gq41oeb9bKxvAc81F6Dkz0/ecUyX7wF5
f0Ud0C5ScDUR1YQrW9c9yDznCtqqIDUkrPptUeiYaighcJWLwlWfJyZIGfqlsWHQ3xlPI02+z9Jt
VPAFdK3+Y6rfBc4pUViUDcF62+xMl/P9ENE0qELlIDsHCGYLmrsmadzw5LDTrpGqeE7QJ77nArbW
Vk5jft7ou9AslZaCFyoNIcXl4hreKo5LHI6EgS8PBKdbEK8Uv1A2JqtpXaWh8qzlJZ7N+OrOUgmj
UK98J/pzJsvTKbuVCG0fI4wPOuehWo1goHIjRe4v3qzLgjgaz0WjqHF52Et4TsCGvb12RjA/XcEq
aVxBEnVBW7KkoU0ZqAwwzsepZ8tu3kqHgMzC5nx1o8EJciAqqkjdSDBhjrIXWRIm4yCN1+zCrNuq
6oEJViLx97r2cUJjsrwUr0w1jykTrep0//N+Y4rEE80lG0t8v6FYT6QbBP2Jeb3tGe3y9xM6EUir
7hqr4U4YmAIa+8kUjg6un4EPn1wNxTM60ANVgdvL3jFFfGIB2z/I/2JBVcriTOwpmORyOotKvwRM
6RnTMy97VZhboyWY0IzBMhUoABgNRypKrV/3sZHp3Lx1IyNqOJP4zbZ7xJ+KUhxUxngKWx55aH55
zsJg+KXiQJ29sTQwgJEiUkcorKwxCf85sEUQRXGYNloNnQGTRtyh79UIaMK0ZENyJKHZjkkR1puf
0ixq+vRShDA+8+xhzZpOjPF+LhULvWqirH8QMzZOrW7E7ynGA0zHukPzollPwIwBNBCKKajmt61T
WH3a3oc+2G8cqKL1/iRdcdHA97SCBa5CcAKMAD4W2m73XMhgQJw1czHxYWasJbq2KgCz86MldtDP
g8+iqETSn9qU3sTnE0cNq2bwiOjbg8xbKu+WSrrqnjbYawNPM4fWt/4vCs9uLMlAYRhk9fxem2z0
j4FrqK8ZBXNcQEknXPYgJlAEl0cKAI7gmNOT9ntXryTGsy2U2W5Cn1kmpAKqD7bklRKNj/GjsjGf
6w+H0hw/cmA+AD3tUsWrSKqmTjP/ZicrVi3OaOdRHy+uGvP0oD+7bcut8m1Iz3DTzN+DBbyqrlEU
t/ZafCOY6Iocj8SBsS0RXOic6mL1DCNyJk8lU1F0eYOHndn9NjaLyj6q6bUnHnRKBVLXa7WZTFlC
V6jePdKaCJmSTvW0W3FzUIVrj7tUiuleTOu4COF/RSnRZhMDQVLvllBMb45zmhmVZHoLLWnum7dg
5X69RlyjkTDIzwubUg/xxeJIJ413gPo1dQTM1RlqPoo8TELniOJQ4PYtbBGspdPphOyPnI6JQOB9
dvQzCsimemzems2UsJ1wfTNDpPo5sBV8ZaVBSP2Kl/iIvlpKOWY314Y9bd63qGHX1LG/gGVcvbui
2/niyr2LmN1cIuNan/rpH32LEGvNOG88JlFSld/Wrw49NXI6genkMPejlXDl9caPtV6x3K2atw3+
VEI9oHwkM9SWZpSExzGzC5ZkfcF9GlMIGZLrp5AhcNsd/oK82bXd43kWhPtERG/aFc/cYCsE+xnX
83n2MB3U/nu7OfrZPAgHHN0GrYUuZ/gYLSKs752fTQAQiu/blkvjLby+tKeAZrop8py8VHhOpJfx
Y85TVrrG0fqD+SQHSo3Grwk2eW/5imhpXB+EqxaBD04jodNWTLAJqgyPZlOLJc+14g4zLcY2CbUS
8N2S2EhevHcMYYmPenmypBbjshUz4l4aGwVruDDeAyUzGUKatUv9cZAbX4yu9/B2Mwczrna4bz9r
xw404/Bgk+1vxLQbX5FuH2XXSwTb+1fm53YnZb/8PY/wjVxrGLq8WbtILW8HoWq45YI/xqo7Gs+3
it6yZ6J8hY7lxxvGs5xmtp+IvTdtu862JhU4W/3ocRz7ArsANUSJc91xbIbM2ocIyGWT0FvO1dwb
X8D89/EHtjsOq+Ci8FQfgN6MATjzqo+V7LFlSWWgMoj83TSp8+yTYL3/wsS94aSGsYdHNzzUzXHw
V3bPIpqLmuhHGzdfe0qVImFI2A1yhwirxVWOdSeAOuETF42aQotsTcuc1IwSNM5wevcpS76xTuf0
Mw7bXFjYgmzMn2wcXw70XV3jvoHp7SUpbSzQV6wlV696I8sYu+V/CbfsKAfhr3rITP0y195tSUB8
dIAHSGo6bgWllkvGhesjNpkyBQoUhYUN0BJYE7WTCqBR51h4Z8NJ1JbBdveJjeSb1CtJRQ6Rz/HO
Sfn+SXbCx7pEdwV9XqfFnHl1SjhxNEbxWCuscX+xR3rg6OJVtYmbGSd8Yzj4fm0wyca+hYVXmHlp
47lrDj89xoAZEXez2gQwA9p4aFqpXb6ahhMPpqNjxVHtkqTIFa8VH7oJ6zZZIFuBtX17DenSKXY0
gl7uuF2bNrLOtX+NN7sMD95rB7uWTKgW7dUQWsmfES3bDCXziDCtflEa4jTtOZu2Fi4JRNtesmwd
XqNrkv48w7AVSTXCiz/3UZt3StaWvo4oovuQoYBam+b39FJpK/knab68cYKTQSGJCTPJw0/LssdJ
Kd3iJlS9D5tXWz8tASvHGiO0BEC682FwWNinV9twl5aq2Z+tAeCnYiz6zgsWJeDIOP9FKLWsBJsM
6bcNsOe4udj3lNkJ6C12wn9IVUEbwDq/aFOgWTiTM+Xg1/FuCTVI/DJWx2QmPHZTI9ZRLwO6LHUN
+1aNpScSgxV3fP7zRfvv0qo4JdY1atiAYG/iwpSSG+3/gshjyLo9GhDJ2612iW38qr5Mu5eaj1Sx
TC6zCRtDtpdtrXBJYewz2bB4/mABjnW3pWhaPKdPxTa9Dd9TXjTfJnl/2ovdriZkQe05IBcjk7zy
7Kcv1QYnQihpjf5ZibjTg+r6CINon3p1k5PdsLHJgwaeotChDKLpj9VAoNpz441cAaJFv1fK1yrE
XYqmFjB4qyc9BP1dFgWI8IpvfBxwx0Y+A9142Vg7hbL5vEC7z4gxlVlt31P4bb5IGjJoXWhe3gkp
bhMwxddTJryVlkCtDCXKx8ykiAkm7jTI8rG9EeGzn+/0J4ouhU9ln06IQ1fyK2Cka5W24MI7Tfuk
02beB/JbWxk9UZej4P8alEiSJSftUPaY5ohQ94ucghVbrsWtQRdzz8ZOonwByzSQKjCFTqTZJn+z
ZnzuzqLEUr+jvP+mPadbmdQk5Nh5HRFKw+PU8vYgPqJHLPeEHdliCAhrm7lsCEWYNT4IwcTZH5sW
SZp4jJnUg5wywzqLG0IhNcJ/NSpyALnoqpTIXCfnVVLOmFByx82xJcEysqQYyRP+eWZCkG9mlXCM
VPgEJA3P6unkEYlxGsVMeQ9hLlUijYpcVsyV2ahn9ge2RYE57EIMW9wf0RnocaPUJyoH51sgHP2O
Bro+lcZqYJQHE3f3srj36o2jzIJbSb1uqpB9YtBwx4ra2G3AAK+EQqc6d63gymVdYSXlpG4yr1mf
FEiIo1fOq3TLaUQtsVnDPrVY3iu0YZdyXCqM09jm3rytjDUPMjVH88ryCWgLo/sCWkp7qFShd1BB
zRKiblHC+X8tumPqm+4dLe7FHy6Lx/nb6GOWk9jbc6WDMemxNbCzyqX6OSVDwH9VLrQnAonBg5G1
6i7IdMwZypM4olYdq+IRKgWLDQMTucnVUUC+8VMVgp3sqMlfMPfRk39ZDrU9URz151IS21c2kPUZ
SsuFr+jPnoqZCrSQ8Kj2XgB9Bxx4nnST328vpqF5U3N4kZV47pJJBoHYTEroLLB7Q4mexv6WBh6/
0W5wE3BKltrmNvn4ANzSau5/k9u57PhuB003K5y2za99wD6lXw3JaAN/WJjsGN8VEV/lWwAydAUa
agDLV9kapBWFE31K1pd5NQ6swHJMs/SlHlFmADf8JhFC0QK5jfxFJ5mUQhGI6s7gM6ozLZIEqCp8
i03ASkYIayJjDRh3472aftKaJ9u6snRSg0fEhpRCmBk7tlU3N8gCKmamM2BUTiYCr7F7BKg7L2o7
7p4/2OH1oQEZr4L6oJnn5kPZsTbSQEpfBkisnLgjTKhNC5tY7toriNEZ1dyd3SzxpeYZjpnJbIg0
JSkPith1zN8NO+G6vZ9+7o1HkkqJvrMZGFKZLbVlWVpvd9BCPgq72/qxbPYdTyOTQpJJbcGvqINI
1ZhDHIdqoESTPY1Zavi/hbAGqLTTU3fyMSwxGWS69HcTeDVzYtxaYloXQWd4nQUqVUHYNuYY0Uzn
aCycNMkkJtGj2lhpHA3yr4v4xytvCYesnmRLz22pESwmtgcS8VTi9IAtZuOAvZwsC7B3qMDyHbxS
Z5uAaDPx08cKSlHhmTitY05gXW3cFCKd1oFMd2GwpvmxxDCbAS/WeEAILcrCF6iKrKrjoLTchwP9
JDs9POX/3Crc8RvMUuVtpBGdufwSLAcjdtqsxJNpw1UF9bkVJoflTl7msVY3shgGMs/lBfZeFN0k
nvffZzsvKVYaZkqP1F6CYitDZoHGvgOPhhDR+LzCx3s24Yj6ESFM7Z8qXOxi7L0YFYyBE8ccS+Ru
l3qYhYB4Y2Q2xJ+PcRGthyLRqgiHyhpCesPPGY5Tbbn5fcJODDoHDX5w8xpZQeo1yc4dVBAJLY6q
Dv+0Ed1wACsyqhvUypHOR9DbXjxPm59t/m+Q/sZrcrGf3x8f+7kSaYvyDkanCao3dSYNfyFqJ+8a
ohXn2O/AH3R5srIr3a9g5Wzthpez50vfNFULRdjiwr8kqcoUAKUTg1G54EFW9LXiyFbjY+Q+ut2v
QKIQvW1/L/ByUSqO+A2KibwucYq3deGNbJZ2PNxYngLF8keM3oupAADGiRA9F6FtlDq3voSlkgFi
+TJREXkLfD47sgIS9NfCrkm5uWOoEEHZ7vV7i824t7Ena3/2JP32CM+zv7sUc+xXzSvvvAf1zQKz
UsW1ZutyE/V8v1jk1lR6G1qK1d6+Tr8sLWUxWRgbE3QLmOOS2MCgQYbqPC2Sj+ZErrYVA5NZIJ6D
h3joQ5FMMelCxYOqUuj8VFsDwND2w5Vo+1lEqnz+pRQVyCc36zj6CajNcgz8GQT/Kr/yXam5gu2G
Zv0AdkpQjLdkNTo9E6IN6MYeUtzwincy/kPaJj6Wgtwf0XsRJgFX+lGEyotXW0vLPhNkmNboOO2n
KrxImxdxtRHRlwt9Lk3sK1nHm3QTr52R9+fY2qN56zuHkZg0KN+C3BYHLghhgcs311HggCpnpxlf
F31EuRqFtQ3dqekoACS4ZXHdJmHp2v35IWAbYk31FCdEZYPQ6jXvxxLN+MwylJlPfTPtCyPyhpfi
W5/LyGuyy+Bm7xE91qoXJJe2ijby1x3bElMunRGCfzGkPY03A6sCL3pgSSyc5lhGp8Wd0+XgaBMv
BLEjI14ci/qUedqjoDRJnZNKx8jKIouvRbMa8ni5IUHnuOASFOEMBKyUVPKhX33IFAIw3oK1zjQ9
D1O1PGS9G2Xf6iHJMI1becbJSBM11WEXhSbk/lWDCdgUyqDDuMTMYmVILrCSm8cz6Eoa6kdPOsZd
oyMy6W9qtgPEpbtSaAwEA+GBJEMhfmCXWha8MBJKh0/dC/1e6I/C+xV6Ya5wfUXCCOgJaJKHZRJk
7GgRWBVcR9+IUwNdZz0cKmzD6Wj2oxP/bGDCaX6Y+BZmSozbq0zvbQy4RvYitKEE4/Oyu3KMgt2a
Jr/pPM+LkbmR/wMaoRRNrMnxUVZhSH7paVwUQ9+zhmh0X0LiCXq2kj+0PnnPCMGm0qGf28f2TMmR
lec851sOgJkSeq+Pi8JmT7bTml9Y8STDYPUza981XpTH2Uj7p5zAAdgVoo19WkpULOuycLgkST0E
KyvgL4TumhDWkOGTWHS/X3nK6qtCmosv4YlJrFSiLrn44LmN9yRWeAEGxRaRW+gkdftE+E2596AV
0scQB8mUCzCN4yFIUHSl4taY+3q0IgYog+8IpjXi9aZIsOl+1QKrvhiMhyJd+ZQtVHWrsnic7Rch
N5XdJw1KDO0Epmi7si5R4vAJIBZgGba2ueNGCA4Z7m4eKnuVj0je78nkw4tPOMWI3HIcnUV8hBZO
sDAaKEJMObP0stf33LiIbwZWWzVHMzK1QwRAs585oshZrx7itXdOb0lyTmKg9ebdJNsBLQK+w8rY
PJ94Yecki/+7kdUgqIkW4AHTDQ87ZRlfZJLF7Lnz7WRm7VdTv5WVb3fxQZ3h4Re8PqYi1xr0CJeb
WiQtbhubvT5Is4DArqV1cvpH1rAGbQUM+yzUxfOpMOeoMUFJ5euz9P7T5+3iyVmR8C02y+abVHqS
pxRaos4NmXeWC0bcX/vnYqFm+/4EmbxPsMg5xXzLtH82Fjn45qhVG0VRgsRvaU74aqlo0itez1Fe
7Qsf2kz7lXLzILSU/V7V2ckIL7nILl63eDcOqZbg3+KQstR/a+A3RuJqE8zARweNBPVtW6JSJwx/
EXB0Iru/F0w/mP5OgQpNQ+fcLSyQOZaa4DX1VBCGc4Ncj0xdftAfQgiUMlwl+VUaYwnCt69giBiU
wwcY0hObuYqNHSDEm1Oh4Z2XapUnFIDkvCTCsUoqc1BEH0Bd3iIBZnYmi7Sc6o68swAcaX1hQNGx
F08YNdwmyQ5xO15ZTGT3iERmpMo3S2yqr6+C0zkSZmjwtivcz22fISuwZFvIkOp75tdhpTA0j4qi
usVuo75Zh3+k7yUC5EQ032vd9Kz8BP1g79B8fBosYHwK+0cs55PVInPcUlvvzh8ZUiRGxyJ1tK4b
GPy5KEhevO6I70bH3dwaXT0UwgzgzrwjfBfLEdrmvQhkWptCv9ufd0g1er0MVaLjFc0xwScTJ1XT
JJx58MLYG2vaiKx2A+mLGKP931Kv4x3Xw+l8uOA+HAjQ1uUk6GqRkei6hpIVCcNWT+Iw2rkskGxt
H5xiZl4OIctFtMPSkA3/7zt8yreZpR780FgRQH5RgR8d3Dw0iJz6Gc4cgiTcf6qeryKG8k6AqC2R
zZXIAE/iHJp6A3ptztVemi7X5Fp5ssIrMkKkw/UePkt2C6xcxDfWPbSRwvpjjA9RWUEjNU87yME5
t+AxtmzCGCE3le05e7b6fUgL6h7grwuQUt5Gw4qRLcXTwhWlzbDMjZCkkRLaAvSlHvQM7c18ZyJR
m+p7qmQBWBkbOZWcIovR835ewX+x/ctxD1AoUp+HdZJ+UNubVxf7YuYgIPS1oLtaKztrTMSIN6/7
84u7sIQ/rWvStvhk0isnFoMgqY0kJHFfrsLdVAGzqvpokQdgQNy06T6JYbG59KdyOPVVp4kzPw/g
zTtHEl3AfVkzWMXl6sIbZmtp1pWn6OiNJXP7b0uXqe7tyHT/v4iMf+yHsWjkw6bRAi2O5hTfSUK9
NjjxPx6jMTNsBF+XocqR3D/SOQq2Gycvo6VrSZSUMYAgdLJgbBvHDqDxoByKS4uTwmyGQSxh52j7
vX3zR3Vj+jOPpiMkNDGSnyXyonGh4XXpVnyOHIhRlg+mU8i9mdFocjY4ReB6MBmyNhB4TLf/Els3
psYvcISwvfGPfw7ktys1BpSSBhISgKqnWgWucpW4r/KAecmdc01t1VRCAYmBamt/MxKMQ2ldV1UY
iOVsk8WlBGi1RSYrgJgD/DM2jv2QA41otssWcpSUdovSM/6pX9rFCG5oKQFbHcYANLaXh7nbAMyc
ia2RDv1eKWkawApivGrw1YFDEsJq/85iU/fA9glhl96GsdB5Hiz1i3u/YHviZcOunpjnOnsGU6Zb
URFDG1m/n1HS1U1qyqJPdQTpge1Mt+Z3+HuQ4JZXxkYSG9wrZbpQrTllIiQ4SZ2hDRLBL/AzNhU0
R9VAj2WZZpom+KVQHSv6UfIa8MziIvTLrRa2Dpp/qSJ9Z+uu5X/RsTcyQMlWxb+tDlxsEH3k8JVQ
+d0QMUQIxnbhP6vXM8na0Dm7/9yuHhCkLCokO7h/JxgROL/LMsbfHuwVZFJ1sB+HnUh/WacZD3uB
0v1SpYD2MFqCJIpwLc0XYJ6gIg5MDZphywgz8MGfXHz6h7yFyHpOloOWjmA4n10fl55c/L8LckJn
2POU5PJ9Yo+CsDUtSRlyvU4FtPXnk0w5WsFqaWacZx7g8+X4qOhSmVhMkNqx++2v0QBh9HGltEOF
Bxy77CV3q2VNCJIBOQYZbQqtWfUoILzDNHtspa8KVPVGLvNwMzETJaVFxG0hsEd/e4uWDaa1oA9I
iUR/sZOf/j4OoBHnFDAeob1uBMenq66s3Phc6V3bix0XzlBVCWngru1MFDFH6C/jy3Z1zvs/P8MW
O3nQUjmh1mtPyAKOAg8r1ZeZFncI2uFPqhJv24aJOH/vMEFhVt+VOkayyL6vqLFmAfTsq37ZnTT1
CR1dMqdD/j1WTpEEF13OlEmjhiZokMKDSSlPSPvaxkbZ6QTPBMXJlPkIq/V3NPrkorc7Xf231agK
RyyxX/p0bbqG58G7cx1iqodcrUO2Nuxhz3TI/CvVAbx36hEuEIkawiN+yBs6ci6tIeWYj05kAJb5
nRI//duL7XAcsrIBhZgviLtzYj1I+GUzZ5bbqssaeJ2NWXN1ZDM7DiHZQj4vDh9bp/F2IYdZhN7i
3QKSe/7IJq4dyoetXDNHegY9n808h9z5ywP/Uo7nWgBG88hJAS7nMyeNcah5Jo/QsJOpZq3KE+yZ
1jm+Sx79AaViNDNd5msCcPqqnYDKyBM1GeQyx7IseB53zoNscXGQ5FSel5M6LAWA8x4PwLbe4pKW
6WxQkyZjd8kgzRZLb8iGDkpHKDtLV1ZOlxp8tQ4c6mKWZUiracfcO9WPVUYWJAkqowrVhCubsmz4
abHk6cfUtGAEJrZMztBR3OM5tvXnC7kN63iLdVXBzssso4VQSeW5VWWXtnJVZuS9cb/62YiE5Xwj
83ci+93c8Lcc3vipjtMVw/VlL9sVAbJZar8EzXrs23eXXK1RXq+og8DG2qQwtedECekjTQSkctHq
4+4QMaWC+kSM03RslcqHbKI6I7sZfLQfAEuf0cgBb8jwc0iB8gwXkDsoYUZLCxluLdb1Ks0a1G4q
RQhAgl/y0aFAPdDcF3+q2Gd9QIQNdQ//7UvpM1iP3KPgH3hy4KknKwAKkVoQNPCOLeLwN0IH9PLE
re7ObrK9Ep2dyU7wsxYbgw8kFqqDnt4apgW8BlpFfOaTMyrzdZ/ncVS7hcHQziRGl6E117rnBe4g
q5z/gzuJ1QXP1XgpAedoDFaLXtF1GGyhfgEPL4952/tXpoT4ZtWrPCHzp4+DDojEXCLgLp6tAADX
tJe9F4Vt9GRehj3i4wvkUiquUlBLXXzFG5I4c/fP2KvH6UCDzkC4vVqDROodh6yhpVUVxK/zbZqm
QRFdT5kDnASeB+EF8gJz11LiXtXBAzl0MR3LCah8tqnpJI5a2XS+WGuyov62WCLQLxYz7v3qhf1E
hNo6hOTg3paEzZZDItJZd+tLFBZ69q8HGtGea6wdcBesWonc3gd5fsfZI93AB4U9fGLlbxvxvZqn
GTiMFnvhy4bDCyOcMpirjZ8ZcvSshbTHyFQ/0WO5Np5+7HbgcHt/zRM7dsiqesDbxIYDcMoqWepy
d5TjkqnI2szD/lngUF5zA4rkVAC9UwSuc8XaAANK7F5GfqbuPu/FxvX60YkuhmIibX8qOiFiSjPF
hADkWRr5KhYdrg8pyFXLOv64kwtcPCWGulGmg762wfZn9u9bZJ9UO9j0Ta90irnuo6/WpKEVdb60
3dQynLtD5jSWERx0CFVjgAJijbJp68OSjQpFiShzQN/DhltVbDQDaARWjVEWFdiHECd6yeo1aSw8
rzBia4IMLCchKFZCVmAnL6ZRWGwZThZOXVGc8jg20f02gSra2jr5wIN9Fgr1FeBKnw9fNVYO0Ahi
WP0cE0x80EviWbsKTnoZiUXFGHNiKgILqWEJCaWbXOEPlhafJjjvcVIwEr9QUszyUI1RiJqQ4fBr
cVF8GOmIcVnmxyP6zGSlsHPdch+cXsxi4mzEdbtV25N0lMXZCez8+g+WKzFFBpTUsipIkgeCFPtn
QitzKJVNCBIQ4ZUwHdh428Sgr5ggdNZgi9nI1yxFVtbQIBtJVy/kzTPrY77Rm7vW3B9fQn7HTQUm
enf5xveeHNRZDAzloVEpZK1n5G0D6zW8x0iwiwt08ro8LaM0q0uCBfWn1qkoExKSWNdsRaMzZpt3
/p0fTlmrNptS9g4xKPjdFt7QNFOzlbGcPM+LbtdK1n3GIWyzcYDLw0ysdGQp22UNXSfE/RmkKjBa
zi8RwpQFWFncKKKu6ZlgpWAeySpAxTrg5RRdslcUzz/S0bkl0+mA74velh833ct8EhItstMm6hm0
7BvHGeSW9cbDFUbkmRsBpNximu7fyfianGpWKPPdKLQVs5Y260J7Z66g5n4hxS7WQVXA2M4PaXeG
VYd6RcehcH7cYMsh9k1OPR2nvtCi644bApA/3TbR2Lt2Q8J85agFO823rkYGhaWQOJq1vsTJOeJm
w7CdxpQzqyF6vFjOR4e99f3o/7oxsm7eHOZYWtoRh+xIKuOoHEGUNG80XGBVTtiZy6HACXVDJnto
9IniN3v1sGoDoPtjbJk/csiM88JFhDYihsx9vrvIjovZ1qdlGzXaTRjaK6jMFOH4+Q7DrERLG2v5
jnZw0txwsxSzVN3+JwRWsbI6i5sLVW07kVN4tY2OMHxFz7DO4I15l6MYC6K+HQ9T3kdxvJq38mRU
+Pqr7nkxhuNbEL0XLQDmR/j2klK7bM21s0VAslMHLiu9+Uf1STvuJ6/dlokbT+pfyzGBgZrX4ZEd
OFedAZl7YTlMKVeZ1ZGnWANEc5C3M7TBXf3s4ZshnZGc3f6SK432QPtWEoKV4Oo7njglxe+41ERn
oU+IVJg0WWisv3/z1DfXLOFDgd1swbmDjYktgQ3NYHjH8K3NPWt22gFuhD5zLUR/uaiSh58ppcEM
nTLWSfv8GX7poEGovlF8SgLd4sBjxTWnzz5/hBWMdXEnsNS22T6YPzo1H7ajgRD+WDlCC9lFGZ/r
z4bqe1OH+c12QU409zj/td082lkLhl38XaeoTrD5zgnPrkE6SGiiKzSQntn4trjeSgW7I5lADKTA
aNlNjVOl2JeZSnON43zm0uD5rPsl59L5ynBpqbRuMufY1he3gg1FtMRYFcZcY/DPvk3BhMDxy4D/
3JIDEIzVZphHmlLIc+o0B8Fwx7Z2HH2qQHgZlElZtj0D0UChGvmnbgyccXhWVaSjhzy7zebqqrvA
RJTnuGb3hLBzZv6Mg+TshT50C/fYgzh8nuFQpxoExSuOHGEdh6MjwrxE5tvEWpiarX059WZ93+Gm
x5SraVy+c+dv4KgipqCC2IdMvMrMbAxJhCPrCZbJYdePlAQXO+F9mT1X2kmBjOd4PuHbBDRo17eY
CGQ81ostUq2Rg3l74jCMTGOXY+lsAY3D2C2J0Z5w9Yx9P/Z9UKdOAY2x2NoBP9MnwTLO+fEQ49ni
L/PTCI33tGZjL8HjT58H6iR47pS+i2K6P9tPNHox/rKzA5KChz+ZHaNcorKJ68yxktTsJiUDsUya
718IFGgWS0WOrEFaV9YKw2PTVZUyis/WedWN370DAwXpn2nTBjH1p9ardm+WGuGToe72+yAlenl/
xOXsA3Nbmp0M66P1+D35OeEEka2XoRxyeNdUCzRIH6vFKilFJy/r/3yuQMIBhJca+1eAinXlI4yJ
b3Sn0AvqikiIhYgNkQJMYYyMA8aG/9WtBTnx7H3t2nCeWSGtnXncuJRf3JVdM0kdViJ7vpeq+6k7
Y173AbLsKPp0+w4eh7LTDVFkeAc7V+y5usbDJNs0If7NZMvFzswYC5teSwleIF9cOw8keY1tsA4D
xvwqp2Ekjm8DSk/GO6gss1Vcu7ECyH1qUeUc/RU675QbAu9P5MXgQ4U5X0G7NKoTfoZ+X/2fqS0M
HFtdbq3GP6Ayarsfqd0X+LYEjraC2GdQasCyJJjaUGLAeiNHlWBk5099sIHRiYeAup//4SV+uNXG
OFoNcmiusg5KGQ/zl1T+JrILm20Zi5r8YFTjkIVR5fWxZBelKyJGW8mzy714nqkftU4BsWFnA0Vq
W5Ed4VfBqnuEjMkuwb6Ot1KOD4i4z53rJNtIMzQdfBxALeOxRqqyItzMvaNIDl4m5nlcZY8Nygmp
X5zczfmQ3X6zCoUIdT+1MfaBqaINW98umWdjZhx6s8TvTsZwu/DR3srIIQKR2xwmN8v8cP0xi/N1
9q8EKwdNyOn9e0w/2xKVh0pc7+5627bfK/dUhHGk96CWeDFd1CnSMMSYnsqLMcm19EkLa2s9N0mE
A+df1Z6Y2iFzQ+nzZwi5wdYfGBmak9Yr+d3x0bK/UiRQfWR4rxKBkjk5bA4GlrL4v5anHK1iO4YX
cvitR5S4j5kiBNz4cYgJRrujhtOLWR7Pf+V6cnZ2En7HLMUgvEqJ8zGDjYM3rX2msSZ+q/KvoxZK
hrhrSxx9F+UhuIO6uDYgBdrU52iVEF7gkOmvbm32Msa5lSwEGEI2FWz+9TQAP1x4JCzvxHgt7a61
p/evY/VXVPg/bTpWyz8mk5nplgsgEUBAgs9yg4bG77MMKW+n9if9JAz98rA3A9TpzFdxIx80EXVJ
ZBefLiWMwOjLdz+wSb4SmJuK6a2V6g/izX6ErQjJQDAq8weloJ/diYbZZ0/n12nUO9AzVBDkNWPl
I7a+yxR84aCn8DeQnSG4hUY6akDWWfUbwwa1AcTLvMAUCL+TAavSdinngDK4a92cNm8GkAzHoVoh
lW66sMIysrbtaTaPd2IQPIbvgJMLogqYM1qyuYZzZhetpTvLWvM24rAruAZfR11d4ka2HX3/2LPy
aN2wyBWooLpNRsOcchYOqkD3+XB8X2HxDHBk1q1/M7v1/Ws948yD0ffqefjPS/4q7Q2rh2oSqhYi
yDsU7m3iGkj/04Qia68sspBx6WTPvTU2smBttLI6JtNJdf79Ckx7P9fXZ2GKn1WggAd5YiFrLIS4
oXDD6yztxLv+fBqJZsUs/DWOwy69Jlh7vir04zEvbft5CLEk5+LVEUq30EvRFSbfB4m7/utvMi73
lw+oBqmd9UHfms70W6sJN1/ucScj6Jgxc1ejms4nDVLxVyjrmU/StVU58pyXpQ4oOr8bOpnNVrT2
VJlM46AfEpoJ22tBseDycPI+F8/Jxoakrdkm3nuU0ZhGbBQB1yzq46F/BaD69FxmLvnwnhQ0PDXv
Vi2f3KzP0VRPqDOu2yAtwqLqJ7XqeUWckhO/0/iupaAvoIOEP0uB3dznjqb7HNnXzuN9N1aRpVpO
BtH98ZDBJzJpAu4uU7oFw71eIhqr6VbZ/4clpEG4dVN+8reov+Drs0lnZkfFk/p70aA4ohXenrMJ
fTdV+i9Upplu1pUW6wpduc/KSTyfL/J7SWwAa27v4OxN3D3K0RazL8CxxgK0xFYYX2U+dypBF2Vv
9PmNLX8RPg4kCC1i2FYAutvURj6zlBjGN0qEUf6Jbib2aBAIRNTzD8guOPFl4s5zbpokLJ1AuHP6
XDXLyKGYNFku9tZM2DIB0KrFt0JnRAkt3Ppbs4XHuDpkUoPcU/O7kmf6Gj0U1Rqu1ZzjrymwNZVc
AMvGmqiLnKhDgW0RoGdyzi5vLuLH/81TZhJxz08t3ReUo/Oy4gkqRxu3Eu0Kaom4TtywjLg48kYC
uEdWeTAJzTQfnC+Cl8QBy6AIVR/2N3i5eNEZOQF4uQJ4o6xa2GAXLE8O6TOWEXmL11n/UHhhq4p9
IOZO+KZDoF9fFZFLsqL3AerCx3qc6aK3U+MmPvWZLm8iuHqFANyaItxAqPKKITkA0klmdyaj7Wrz
SAo4zdFnGW03P19+0fvDq9KDlGYZ8aI4VQj2Gqa8dbuSyvz3Ja8MD6Y67gg/RTs3ZRGanVHqJkIZ
tGy8EYfVLWhdcXsxTdLDbZGOZJd9jFhjeecMs+4YZK3AvXWBOMkGa2tpt6YMboSHkrfmK00g8PAQ
09GC1talR+TLGFRntSDw7Sd3uTqHWLwGp9Ul0DgdPFAxX/SYy0DTDTVQIigxpaQt3MYLLGZNRJMF
QzGe0nktG6rHuKCsOgSSmB9yMTqXJemuTtcyBQgepSW3ePj3mv5llC8RTY4WgLpbFyZb4UNHxS8P
wj4nhD7FHAhqUQiBnsJDJ8uQubPExpJvj07NCXBiqSGCl7gpXuuE+OfsKBkHqYuwXCyfupHuWDzh
WzvQ+1+s+0yv9slMLf8MTTaM0x7l7aR6ufHxiZ89p5TzsVsdkp49/Ehe5IJskRYYU7n09UnUmdC6
8wc4z2xoBZerzKNJDKfXiiRADZP7KoL6j+M/UCrgudogiVZjk9kFLbRd9zQcst5XMWRHqSOIEhz2
22bROgZds9XuloNUj/7O89REA5f2GAtbamAv1V1G00XjMOJVmKHX34ArLUq/DL0yfHSDxJxXgtdA
Lgufum9Th5n+UZkgH2WFFFZoePseAonwSXs/hXg64dHLAkjcLV3I1dWKCCGf/9kcQ78hI+4LbAp7
oAXkz/DG5hs5YOkAsPW4AMW6uCgRZZr9SH6HhK7ov8do/Bh3wKeJK/6moSd/kPKt+bRbkETQvX/1
LW1tAZj3cLkYAFzcoWuWxUqTrWO/WI1TXMn67M4Xk1QMywiwZEXGKkNeqfWo3eMQZxgEk5WBigCU
rgaXnqDiCxoV/F/4UOL927qGE0xxqOSd4WRuNVQRuHMVo7HU7p1qIKtDc0URa33/1za43Yc7asDm
77FOkTJ1+L4BYNUtPPWzx92VyyS0LcDmr2h4YR1i0H6QCDHLX4tEi18WUFJ736VJ3fJRSpu6amrs
o0nETjG4mal2gDbbZ7pkiXfyZddS97uA63r0pJxFXu75RmrfgKvEq5oERtoBWEtz24v9ok1O1V5j
YqQHaUBKCqohGt7GwKFuGHqBE7bNGP8zYG1ecHv+cmzXp7ej9QAXxiu0+8VCj3z3Y2nTe49md7dX
fdfjL0P3ZRuYE2nLaXHrzexywZwKv45MLLXS6ZZan7LW27N1+bDGMfzQVGSW0g8o9gkEilMZRnbq
QIJ0KdNSosAa0gWzKmTD/j+1ehc1fDIFlYQakhFexi218Od3z+brqlhl3MWRkqGIJu/Qwq7qcRre
TaEwBGhGwF1YbKdAzatH7UTRXxqPZUSxo05aT2lhO+rjy6ZrVC0Qhg4xKsZTg7gLLoMPq+uEoeXd
J+uqcoA+j8Mqr4AplO8vEU2Eb722LvZvHNqMUN7HJbcUCSnaP35eIgz+Ehne9VilYiccQy9l5Rk+
5xnw+hYNmsa3KDjnP3F2jw167KEgGKBsSgxeCFfQWDybP5zHzl40Onx7JA2wLJG+n/YqJ0ldAVjg
xusMMGJ5WnC3qbeqw7l3xI4ake4WcQRjfSws6igGvnZ0VQ5rdrcFAkh1UBXjCoRGCKk25EwtU9R6
w/On3FE4gqIHr1FAYKRImzb5VhnF2iMGBhoy8x+UdPhfTnJ6sG+XxwVe3WNNLkU6z+gbQkI92GYb
xiMaZAfs1ofw7+NT4TmXGGpAdc1VK+EmuindisGl0fGsU2rl8Oxq0U5bwHd3iicrGCPR6Y2uNDLq
7PcjfHsgYoTmj40L+Unwipq7ztpXYUrJ3zaqOf6tB8L5McUZLKJFDs/MictYR3OmaE/QTftI+5fA
T0TmJOsGGoIkyRDLZcLxklTbxFReyNzwHTi1tsMx+Emr/Z6kNfc931EZABwhhCtAXGUMIUDyyRYb
Jcb1SwicHn5Ub+72q1Mkofq2NcghdeAgYrh//de8QdP0mPmsyWzq4UHOymRsu4Mr76ApZb2FVsEO
ZT41cFmA6LLNiKa5yLRoHp6A1VB5VrE8Z30ADfPrZLA257g+G3lFu275BsWm4nVoMEx01r+aoRKH
g53GvbJUxiSF0J4v8ifpPlK5WhHlaEumyRvSg5zcjzvyOSmhA8dEUz0jkUtd9nnjGr2WdyrkhQ8b
+cuUSapBIvOg5IXJhO71bk9bxhpnj8gbUhqkZF2zrxqLMXfM91xLNHnAm/4Vj133MNIp1JK3tITD
giwVZ2fPDxeT1f+k6EiJzNWpKpeuD0pUwPJbhVEj6YtYBjkUc+LcV7euoK3LxvFOB9cl7PPlFnCp
FFGPMDY7HLhtoxlF1THLDiKDMaHJtpCjgSs4Fg007GaMQwexnsIQhWoxQstSqMGAwzZE6Lqu0XQ7
qH2pnVS/QSBbDLRjtQRBRTriWe5QCJJQTzw/DgveNne43CMzFAWvuR07PhSiG4qinTDhAa28J/qQ
B9Q4TMwVlu+p+p2ELR9KFZgVbJghujc1uDPX+MsptpNOs0IQrNtHm/zBFZKwz0bEm9EhH+x+u/jA
LjpwSLYcDSYEhAUoVNSg3h9PXb7Tm1w4Y5cqy2wVStdyNWT6v9ucEO4J6VrcdowY7E0Shxf6kIoe
ktcC6yak+/oRzxhuo9rjXgtPruvmO3PZy8HYxnyQ8zFbgmmN9QeiZ8Tw0PxTcHb6G3P9MFX4Wn29
iJyu60kYDnnyjRZ9WK+RaWg8CI2KVXsLcbzkuSGtWipQZc9aARjcsuv6gVIO3FZXkIpwqfAxwVFX
gLJHn2cvXYRamMk+bNmvspbS2tYI3l5FGknSF4elwIjcoThLt1jGcS6oBNRhrFrRQnyQeLK/NIJZ
1ox29ku0RvgiPUsXrUK3/uUeYsI2WwaVjuf1gDov7COuMEhaqWhb40WFmHPOyyaZdcgVTcHK9uWa
oP91HYC8+Lsqb3XUoKwJg0fXXyATWMUt+T3L2lNzI5QPwQqd97gvNUzWpXLnvSMbpzXLmFxyNUhd
Nv2QJSsP8mnbZxwhVKwW2yYIHmJS2P9sAvNR+H8YV43jS2QEbpOE7OChxxTVuJDbg8RLBPIbvnLa
IESW0JkvOOlrxq9Yk2SHvx13RHj9zllv79hvaB9eGXsA4oWL02yiLRXywVIZ/NO5tChryBk6Gkx4
CxN9koPU9Ofcu/CpjBaDhu0GlUFGtMCDDr879ra62ie2hdhwUOpciSBle0bRDv05h4BtnarOlJKo
1/jrLseoYJjxdqWR7VXpLNw2e4NttqwTxpw9LVKKFYsN3abgt6zg6WGUailoQWLKgcuLuB+ZxThN
9tlsRs7gjfPuBHbnQEpCPMQdihZzR7giU7E3Qh6kQi6iPP9DplLCZLK0pe+fe+AdpialsW/opiPW
9eTxelPZTUkByOJ499lE7xZ3ls44i/82q7KrImx6zR6HpZFTTx9oj2P5PIOTczDqlDwQk5HOckw8
Ip3u0poaFKTcfJLq7+/P37PkbxrN3AG9oEDYBtFf9MxpNb9Y1XRww0LisTCIjMhULcaCTs4VEa6J
XMTBuzyXfsV3PrwZQtxa/JHLHsX9XW0p0kdyHozqIFEV1eZj4yd03+0ZxTvLnbNvgW04kKQgMmBj
hjZG+XP7UglTqtKglafeW8RmthNSFUMErCwxVO8zg5KQpkya6v8CdDMS5suwglPBZFTJ049cVjBc
4HNTDJtrUVyOwFHNeQGjrx5RADIv/K5GIeoNszkp8O076Vp5J9I5WEDd8V5hX4j10XP8hzjG8fjC
VroRkZS74KkvazQnJReXrExN9RolgIRv2oEdmIX6/RxSKMLZsW3RHoRm9EOIM87N1/DmI0b/XhcY
XS4kSppRwo7mJT8MIP74uVkQ+PEEhouDP3oIIaBxiCapRA/QOphqk0dhvIIuwjJg7kwLW2MUgglR
3wgse0nqGowgBxPTodTcteO2hlUSEMBDV/0niVdoPPrDUiq/OkGvhiiWDrV9zTzcYhJCffypquc5
EnYSbguieILZOentV/lEznsdr2T5qIQdjUt+bmnP9MeHG28UHvw+QpIRShun6qswOfFKkZOCtjao
zUUyequDpsqEnHYxkTv9/IZVLvonSBCNnb21vBZxWlDshvn/08imq805V+AyPqEGnXrpfKtkYLyl
1UuYbeVFN4qqeggQfavtdVIZxgcoMksckD2ZyJSSOG5YUf0Sv4N2YXaT1CoDPjkF/0J0/z65d7Zc
QT1s5xS9IsaeFbo+RHUEv2jrVzpkVV0tevV+h3TVSpbMeUqW/0hUca4rbR9cJrqAWq5+2Q76Nv4D
02p02WN6aKzYqQpPODPBQUKqm8bVJ2cJtB8rcQr8kl9l9kQtbq9iksvLEOlg4kTDWPpd4ep9HKG0
ZDiqcFb18toJQqbPFqDD0UVqAn23E9Q4Zv5vRVw/uonJ8LZo/YHO/hVzpNQXtFm8ORqWjG8JfSYg
cS63tU4hNjJNXg8cTBFqro0X3bNYSWcovVRiRMGqQn09UW6YDvUMTjz+7VwMr0onSuDn0xzesP6+
HMhpzgUzTrMrBJByKuQge57BCrKl76bgHaOqRdQ4CzhLtu+ifQxbO0sZiajTz0fHPeP2XRaRCNgy
x5u7VmZcdAczRSRJtYCki9ugzeJWvpwciu12ilyfMq+QBs3gXTkaCJFKWEVf/oXQ82QcOKS+XEdp
UY/F11bPLye9Hou4/knhpErqEKzjOTu1EzVw66adhaP6jZHR4PvZvkfEws+dMGgpRLRN6AKLSRI3
vMpvZ7gA6NpFqrZZtcSX+cM9iFcJKdMZPkXRn6KMS2zAS4OcHzpmU6ZhCREYQekR53UDfrB3k554
+zF6hGmkOSv307n6PKFFLPEuJMfwiQn46NhUIaLN3lby7If41I5TnxhhW7FRBLhmi+fP0iDxPeZc
Ms3rva75VX6ftV+Jy5TqlabKb1Ts7Xu2V6MgB7mdVpKLKFl/faxywfXUAgoq8po7JVFm2xCChzCB
Th0AVzwEQ/b8BtfQ8k/EXccj/AmnxOANNuFQEUrgFQkIzuDJ0uG8Z+z4UPnFduc+VibAk9M7Zwl3
qyI0Srg1SoQ76e5oPh6vzeDGagW9nZhMFw84tzE/akHEy5CAAyNrm1xUkMzZnducT6Ce3OPF3sEw
ObqeC3ShP1T2KxLJa2wnNiFjXahuNIUeGl0FQDBIgmuJFmllg3rBPVQ+NElDfb+48a/ZE6xZweUv
4vWttHes5eYSs7Aq5QwcE5+JP0W/wu49mITxfxAxuxlwavP/f1wE7deXxufNOOztBgI8OB+CPXq1
eFzdd3yLlFjshdx/Rf8lCQ5X6gi6AE4hIIqyauSIh4h9nzIK0ZNyzY6B96xzFxYldZ0ZR7kuJweK
T4jMi+jcYKG8y1jU0mKwv9XGKidKHy+sK/0Dw0c1pF5JGdWhY1sJ6tHQhQf2liQsoYxmQfK3Dnwc
+X+1VR/OAPdXjCPQ42tcVMJcxywIFSIsuqLohk7FNMtIzEOb2K0c/Pt5g7GYUGAjymIk653a9R/7
iDBJo9Y9Hgsz9P71kWHd6uCKXcYh7DRK4IJt2Z2vM+X9S4wPblpgK5165OiL0GqLW4E1IBhndTLU
MsszoSXaGoy6l4Fa2l+yfylsFWhVnbiR4JsRW9Zi2N1dG519W9ZDvP3RXkCufO5tbYy5iDFka7EP
/m0Vx7zkoCj3ENzp3VzqTqzPGNzADOniEp7LIzcD3PnydvT3fjFkK9ISypqVogPHbrTwljJ8dzwO
3fRu93rn1deptDn53sjdvKDhRtJq4loe3Z3eWqbOhcUk6CLqDIK3Fadk2ZvDVsCfEUjUgZgDlOUC
lLjYHPLv8r6sLcbbFT569OzfDq3uFHE2AR+AZu0FYGa5BEqvnXU4WeC5XUrOFN8ylMW7ILseR7fL
xRI11Oy1disgPNvaZdS4xb4h1VCYqN1AIKfE5FhKrGw/m4JnQR1xNxRly4xgOa31MImFx+UxGgbG
ykq6vyfGIJhDHgfsFKn72pW0PCbibT4pL96XijXCQWu9P+xJcSpmQu/Uvq5by/30UE6BRETmG9ed
eLGqp1YwuQilUEDHqOc1EGJ1ZHmcC5xxZBnAbLeVawvSA0jDivJmHVnbXMZaYiApJEphmDOkScUa
CEMxzf+pY3Z511td3U8k8licoWze2vE/6KutXPWg2XqqvtG3Hfh5znfiQfyqgofU8yt83OYYNcW7
OfRbbzxwmO1AzAcV2WcSxmzwaV//5slpJtrmEobpwfyqs6PnRqNTGrOxnGA3GYJi0JEADoahKWRw
5/UlrMiK1+u5M+K32FA8BgCfeqwX1KJ6GgtC888+1GHogrlqm3mCJ06/1zqZxuMil7HmAUaaIptD
hXfrNQSsony8Db78+s10gxIdXyEjyQdF+K30lvY7z4Pl6PLtcbWv0DlqIDO+DJYTeJsCOjZXgQGC
/kP7fOf7VZzBYoe0degQGykxILnCBKC5Uc+T1V9oL4ccdXG8NxnIwMGrO80naiwINdubyTDUIp9w
/8+vyLEtXsVPRmadzviH0UfKMhWWAPaAjPZkja2iJZakW0L3+n2FCdQy0NfDy176tg5mHX+6vpzo
H6dUzRP6yFlp3l6qnYIrhpOQKbrNWrDD4c/5kK6igaFjwQ9hMtUw8XHDM9Ys28rBrsb+o2dD13Fk
u3Rjhvr1+P8jxltOtXYvs1B2AZwFMbsEyfhNf8k7P1GJhbzXrYklMmNBA9qjAGeCoSGpqtnFKFi/
Qzo1XY/vBupdZFNJLAcwi7Tl3ovX7yzYo1YJtUR/JuTg2M1wwYfBptoA3gW1LFDSK2+2xsl2yoH5
x7wAL8kLpBzuffG7FsHBtj9whgiXZH19m4Eb8yytcYTZ+n+Pj2m76l7PgpVXdo60gr3GXF4/JN1T
fUD0lK7lG0kzkUC6mX+9vKkKJgTIX/bEydW+JEnujKV/L1T+LUXRN/393Zsp+FzymNGhTD2X8StZ
3yXGLKAmCWXBx2l73rDj81uy0hfNsHZg6uv9L7ZAwMuQ17oWT7AMVDody5yEcQFZNafejxEhRro1
shAh/SGG3xFyW5QlQ1BOiQxCDp9Kxlws8E+bJMIn/hdlcZK1hSFt6l73TTzd8cJ2h3cpgf75eeO1
GHfFoJDyPqm7nAaB/OSd6DEVGFcTCfVoktozeNjGQM6xx5Sedszoov3tATJMgTkvb5/pkIgHwLQE
xJXSgyTiYtE2QnozFTY6gDVnlyC9u47wnbJtfwV+rscaS/JZijHjBrDhmutNHUx6cWHHesGxjtBQ
BEaVqjNeKFwgMWCgLubQadcWu17MsHTodZvdyh7WE8saKXrOCuaL6nAykHuY04ARSBNUDsPSCwFn
5vigjJh/JVZqV/JBVJUPCBvcl0H3cG8/W+biKGElPEM28yxWpxTmI5yRczgPUbEzXE8SEQur/6a3
Lv2bmLqQ/y3hoRzDW1xQkF16339lTwsujIwDVuAfTSkfuM+QY8MIkLNtOP7u1ei3fs4L43hx+//+
D8Rjg2M3Tsak/2pr67u2Uh85J4zr/g/zPtHYunhYlkfpOEySEebBqe4yrclNvVHujvJzq9F2gYXM
Fduq2f2IXRl4irK8iGOjt+jZENFz1q/61zSihp2r6scCqR3/e5ZU3yLLeL/OJoLpjMP/ugW9sa8y
HrPcVpyYwOMZxb0MsmHzLu1h3sxIcE2R6SRJ+pUqBnoUqe5cqjo8wBQ02HOJyBk6hE582yrAKvoB
AjBM9BOs72ro1gej5pga3LHRRrFLxv6KpD9G5kZa9QISX2rnNW5lqCJDweJMUe937VjzBCkgn/Wq
gR6K8yUYLlJS0V3TbH0UkwlxgrMOHMkhqeovi3X6Wc8GJyMC5UlZd4eMJ2dIBMsS+6skfhuRlKF1
dmuUr9kjs0X1LRKt0CI7PKtkzKXDSpX6vH5a2c3D2KsWGgIcelNqQYbH91wzpCgyRKMliRI6gF3X
bYGrCJgqatn4xn4JupLhclQUsDTYTPMM2/pH0dEGMcz7Pa1+lKdYvb3QCPvnxoEtWXR04Oy0IP7/
YmYXcGQx6tEA7yFsA4z/HjbCS2N85n7buO95V8f5VTlZAkHZ+pRweELUkBPX6GfKin7uTl25+Qvl
chZ/t/F2cRSkH67/Le8Jn0tZheNiDV+Knn6Fx2gfT/AHyhi+G/+RaPcjBDK1agqPX/QMf8otM9NF
u4VgrARNfgbalNZW+HmI7ic5KtY7EZE4nfqjSBTG7Ms8qrwK/JP4+QyPnVJki9Y3vMGyIam+IiUC
ffv/w1JCBZFKdblT9Ehv9+3Fw8qEbkFFqL5HIf2yYvuDjCW60rUYw9Z+JoxAvcJvEPfaW4LEwYuj
FbPzupmPk0auhMU9bdu6nSJimlHj1HguifLIhX6xs0t+5PJIKYwSWStB8yWv2zjbPsZhJxNDbfJT
82+Gl0bJNszrvC3V52glXDsa8YLya1Tm0f+TEGpiYOD2zX6PyryFopd5LwTf12IGRWM1lylLRD42
rvkApy9Z6rY5Dspy0x5zT+chegbTk8geCWBCot+s2Fxra1no2fTrGuxgAGymmfaz37ITiIBa/91A
yhjXu1gKX1tTJ12PbCXhTVamti7gWXK/6r7p0D0dvHuqwrJZoTG8FjObH0z/ODuN2wq/E8AHPO4g
NSxyBF8UZUlqO5Gmpkf0WEtrhCJxIw0K28gu+a9SHY6jKiqcMiF9yNA7dRlznDri1bJt6YzRRxyO
vvH4a4V9UZlZgqvH+4z3UFDV+InCtuku1Ype2+3LuPi2UrRL0VDTvA94PrNYqoPG9aWWa5/ySAAc
vN4t/hMBVh21sPDmgIa03vVK0J8DUjYm6SCEfUmHJ4E33cAxQXNyowU6CUpdNRII5kF38Rk4sVr1
XGEfCKWJW/Sqa7XkGGf485ZYOqN0LCanhI9ilIrdEEmXAoUCfjWF0CWpr3LnsmydAgIWMmV5/q6x
YfdE+sji1GDktsmE5jHsy8qp0gDY9Vhi88K02iCepT+7gjpO8ewdTH8hoi9I4PflDp7oBTltLBGd
gRk3ZfFGVCnMMJMQg4+lO3JnYPGmDnFH+kJf1b4fOIFq/GlYRpDxXdCR5sEHn6V3+pTCHqWGcaPc
Tj4QHkYe8jvFT4U2HURtzfStym4g9bAHKMabjHLqb1fyBo2EXZUVpQYvbbsq7sgMHeMPwzVuMy5S
07iWF3JC9NkS8igb+AWOTobMPWQXUdVPqCXUhI86R6d3RlRFuzSxWoFM2wc8ukjMDSePgTuWQMms
ENcGuSLbQHn02+05juNEAivI/WorFCs0/XS43NSONKZyxd0FGrxROMx/kAPpumYZor5nNc8pkEx8
AGIHW/FL2IyYjMKUnnT9pZNtv6VcjJspH7Aa4uUPi4HaLFCuO5Zr6NemByJ/KcDauHzLVQCwDMB7
Z0cHRCSG7Lh6gOcDweWAGCVPB9lEEugZMz2dyJOWAUeLG2cGM2dgyiBFvDogZs+Tceabuy8VfIaI
SJzcHJzIK0YW8Ng0nTmwY17ZE7qoiPB/x15wOl9BCxFissNWUXFdz+Z5tzx8ll2ILkPJXFgFevWq
tPtK+ZYZ8TozhrhkaXNFt50PFpKqiZGwo0382Gte1kD6cYKRioHztapgdrvqkg7mb4U2C9ff+K4B
lnnmTDCKh0knosAhCptzJX/5Kh7BKZ4SSt2Sknhsr1tJls/W8qp+aDHzPhZQxBtiZ2g/NpuvosId
N57ZktGqhek2EkkzwKaDfrr29uCywZ1boivZFay5f5ReP9OeATaAsOpaZcVdUdd5htksWtBWV6EH
Er52c6AeTtA54es7pTvL0+xNNKEphQMViw0MzsxYDBN3vh5OzryfaiA9KrYIHDBX1uB4Qm8WH88S
o1tzV9t/50yK26q1F9o2F/Tsa23GzBVNuM0z17hnIprs0td4c/laKJnU1lSjKT6Bgfvs40PZ76ov
j06AxlMB36DLSYpt4Xw1G2tTIim/pe86sp/CLiMQtxe6xx83K+sL/kkDunSh7D//u7IDRbTgI+mk
LrPfVQBoJKqu+WLt8lBbs4vG16GwKlbMBSQVXlQyEVUUVdMN+EwVk5wKWA7nkp9+g0SGUg0GrTk3
RcVp0oqGQi4r+ir8aAydfj77v685IoIrlWXlHHFQNDr3NqGVHuT8eEzLvVpMuXshoK58kBV5fCby
1dS7CssCHKEv/X/Q0vrKk1a+xhzpozEPh/q68Hi+exXCwICONG0nJO1XulYbTy08BWhyUmf3I+aC
UkTQmjm/YV+swQTD/kZ1ljnty5dwMp5xDRqWTJApFiCXq9A1vU41p7zSOwMA5VZEu5wAJTox68Fi
p1on3en0lGCjPT/9g8fRi1Z4am3mROetY9tGTAwQFuY1c6WLjhz/Z5ew/iRce6wMibwPD7evYIoi
M+HwB92L+Xym4Ymn2Lve5w5aY8NdYgUrEDpLpjQ68IkEHV9/JLIx0nGVdNlnNSuR/EHUV1pWdSSL
RZsM+EtU6Ai2KiRMANtKnyyuqZ3KG4ek5l8wSEqWti0j2Ihj0E6b0V4Vm4LrTe8WHLXsXxrH+apy
NnHPQHQCs3YTrMgzVjebT9uCpkyksnY27Exk7vZvSEj5tz7mlE/sZLPLCBB04r8jRVvMxJF1viP0
8MAPpNsdDfTdHnV6eKWBjA4u+cLv+09FnBapfSCsZAdxdI9OLjRm8ImDFYmVbBXd83LYJjFdxTwq
FayxhmKMoJqv5F4N4hS6Lmsz44mftizQcAvx6jI3E6ZedxERwbfH20mDhouiOpRhbttKiXdvn292
LthO8JPM8LWYFysSCpFCNiJFxWq++6kkbDF3ExRfXb00BAboPDUcA37KOroqGc7C6W2XGZImPkbQ
sfzrjzmlKTor4aLQ4yKG1suXKjbQPu7daZXLfEoVQPN0RqM5Yg2hcwtG1SFUiNz1YILiDvbEngJZ
Xvd8FjvnrHqskvGGndhI98bc9CZvdNnKXV8b4rYRtANEjTSh3j0SWE8vvJMGlb3FvzMTCOqA4sZt
ui7i1jihlPXR1jLH9v7SdB1lWWvzl95a6E8fAJa5uo2bYXzEm57F5sJhiJE6HHuGIRdMOGTLJwZk
wzOPUurKQx6TPI6+Y+1rhd8IM5zgmFt3y1TJlhUqZwyvm4jLFq41g0QFkCTbd/M2206JhqDu1JgO
vApQiEF0dhW2ymeOvS12T7ITCBa8jCRsumDZdDmWhgLPJBWgMYgWfK91EkWEqHTumtrOgGxMd1iI
q0F2INHagEX+FUQt6MnmKCBb1dXk0cJZb6BFJCzXLNrtoszTteawirO5oJuVsnwr5uDboYuug6ez
rSVsxyVFKaZooLQAYaXx6xcZ7TzcHDgSG4CO/hImfF0/BAZFMPtr970/PpeArSRUeZngT8TaOaOY
mXDCnjGR6r6vdEl5t36ITABb5rz4S5r0s83PHS9l9AkR1lRYkgwAhCoyYaW9PiCi5USxbKCgwdoc
P1QXTAOzW5LQQNQ5ssLox1hs9tAkID/HdUF/6KflsrKExYqijBVJEZscm1Uld56GIhTvq7IzZsSY
9N4TfrW7Gow8TAUqQfS6kKybnWHmwSLPNM6eRbyk7b0mRql2TTYNglNPfkNKF1Py5eWdQ6dkdiUV
vd+ydwI8bjguD/wyiVv9DULCAMLnUUHWqALaIObideuFsYvi0Oxq0cFuDkRPw5DTjVfpLc02D3/4
FOvPRDD5Nu7NLpuW1C1bkDXemtxsYxmnRMt67KHxfsotK/mpfHsYDHR9Qm49rvLURArQuKs584bp
kxgUQFelDaWlNPh34VO24d3LLbMKiTitkWHWgZrLfbb+t5RR+4ZIcznsHaqNaaRw5JTa5gZPYyAV
Ue9Rym8Dt1SmaTwSD0Nhii/0wk/p1zBj2oHcbpYOhnV7a7CncShHn55OzJiTpiFyXaWbUQjjhK7J
i/mq+59FYekuJX7Jwu+z0nBauCjqmu4e8iAKyXGk4nHUjnGtVPX0uorDikqWXDhjC3iiSQR63KfQ
+2sLa6l3xulKtt2W3MaUbycJTNlkwaqOY58fmppIM3GE9GSSCTrutz0C4X8ivoguY64tw6isxnKR
5i6p3IjjDAHKtZIVUNkRrrp9weR5wgneUEjk4q3EbX9LTgSjOWsd71HpW4wp9XGzFfwuDJAo956E
pgpsUgcLTM3keobf1udBDc9cYHspQC/BZZGqB85S1wov62Ae+4O6VFLJUi25HCdQXqj7CWZq6DBk
2Sk/33dZbItczNQ6NL52Nt9gv+TnnOTzAEZI3+qOzrSHNdD/VGhI7NkAQf0BQP6ZBTvjSWWASAaz
9uXXr2MbFz2GeRrwZACxTR5zxbiF8zyoVkkrfBoLQ1YvQFV+VkT8Ztc0PQc8HqPudOGlYnxB/xpy
4z7hJdYRf1DexUuljCxRRNh1MnpO0zrkMkU3ajIhbCIFfEX4aQbHQ/kyhsDtKP4GtvDUSO0z8w6I
+dUPW/sX2XTaPZHGizZAfIBFZlNdd+2VbUlHHlACMyl8bwa6KM/WRxiXSa8jabGg2ukN/Rin8rmD
FNzYHamEWzIDCglPVC8kqv9YxGuGM/Ii0+t39uCn4lTxi8YPt8KBkCW01CFPBQ0xo1cR2nwMzyYQ
rRGzCjcrg0BH9KvsoB/Br1tUsoBnKf3g+F3B0Hyappype9rDZGdrQSA37IBuHiiO/S6rpeZCi+WE
yGMwCVZZHRWKXI33MQpGO7gVKsKSm9JStbCJI0I16VKcIppb3620qbPp/cno10z6fSORAfD8TNcf
NOutaDQbOxAjaUmsaYImdlBY7rCjvX6n/LVo0W0XqLH1ol5gte3ucoh0avI4v+IxpbD5Gl1kGJbe
N3WoUuObYlvU7rcb89RwrBxSE8T7yH/rd1GDL8DOC7O8zoW/IugAM89mp1fJKnS7+9iJQDZedTHa
nO3f/neI6YNDU0LWm4+3lyTV3DpmmqajSnfWASdaPTnROAo3IyDpIPU05pfSkhDFkrqKJDCGasAz
FHiZf/7mB3LyFSWWMxNhGPwQJJIOYuLnU+RpJzNjQWW8kbozSEEIoth+jKR63+NCNZTcEo1K6lb9
rGoqlBJSHMV1fYekmlsv1Pj9C01wqL4RNSW25KjzOK+H7Q1XC/0yZx+q42XHiFcdluA7ie6e7oPw
ObHbLU64RYMPOc042LwavnkrBf7MfOJI/7Q+lWRRvdsrC38O7qef3FbHT200E8TlVj89zBxiguAS
043fPvdQEQG2Cntbb/bMFDOHeRCUXFbfoQhcRgcMn1a74PaMzOUDTKzrAKgbUMvEaVy5IrNxk2DO
Z+eLGbYDZGK9h+pp8+AwuVp9lFEKIttn/zIX5PRRwIGSfTM83eOTWNMYLIhRYyNxTrnFcvrC+qK8
R66RQ2SjQeZhwCBQWdAIAhrexjke5XByr4/exZA0A+JMQVBiBk4TGKuU3mXkoByEX3dX30c2X+SO
jRTx1ylFdXD1p7BhiYfhWQSeyGbd0VUTCR0zjLtUBUOEK3lQNE9ECaw8ZTLZ9pqyxOozDMgx7O9q
+rhCrpLzEfD0XcpgBfMqHCAvAqvCKSWC51Cwy79hVM1YdhGllSJWNqDHy+TWvUmqOr5L3ZQRKScQ
uHjpt3z97B7pw8vJiTOa2B7KW1G+IsCBdz+QKxm3IMp/6xqlNabWjk53bpsxCBg45YCBK1msXE2b
AaZW2cXa7zm6HDzij+7I88ELTYKLc9H7U4RDPMwpsH1wY6aCLtlA6yBIm7RtjcXbZtdk79eblzmd
6suIRsHfK8WZ5SayOFlK6MVsJBqWMaloOCRFafnoQedWvz1ypXonqNvg7xY1rx7fTTLzzcyXKIwG
CTummaT0uJd304LGAFbACnnbb6QATGZpc0mdrX+H4A+SWAYyGeL5/pF1QUGEyf9yKLbq36QiUh1V
eg7CQQJQPHowfPps9OcuZLIcT3BqAIn6vK1Bb2HfULevq3oEUwBMLH6vrODNmaxVtco6LCZ2GmWM
Wd3U+mHuKkGtpgMRGBnu+eHPm7jrugIoZYRUcaNA8BwiCmoeVhuVVlxomMkxdZSvBEgnyLZsRCe9
0lrRT/DwqRk9eM62cW6ID7x5RqmLkrScbArAztKxemEraZc4A2yTlpcnwpEGkQhiClLotBsuZt1O
d/2hAbcZsYC8Mc0EY+Y4jB113FZz8qKr3pys1ECLUNie45T1giWXNLcZx9RYSaXcacWuMDi5N2RA
nNr47olb0mO3VzwfDBZ2aj3wULs85SyABQVZ+qAdETh7/PbjpKGe+tNqaLRQqOM2X7PPg593C09P
9/7LZIMiiYkaMlQBy4Kn0TPOQeXIBw5dl4KGFHHDoDSJxvlKyudc7AR/H4YV3TKnJ1mCpbX71ONA
GkPXemijZuvWqy9s0CwKhJe8sszDB9hdEumyrP9ZUo1YZRaSRXqtllkBZ82Eo9HDp8VQRsljxBAU
Zg1NjTyI85x74Iz+Lju7W4D4nIxsKP9UQItQem2SYgvh8orJ0Vpdu/9O43amMSrfISMdAoFAKOe9
GQnCU11qMK6RKRJCIS19Kfj+EUXgGiu0q3m+/DbUTa0NhYGBSmtij6F9sOzMMMBkP6XX/gl+NJam
wJ0Xt178LoLm5A5vTFD5fGIYfXu74nCVe0OuG7nU1UhFQFxZ4TysIiA+fStriZgVv4jArhdU1eok
5eQPYBwICvCHbBkMq4u6r6PFVoBs7QVAeXGMRf61VQU+Umr4PvhgrhmOBXI1x7POCpnYRqYQd+yJ
f+6i857Pk8TxPpbtB7hi30tCiTuokWb4PYeIitlVWb1ze1+gjEIToOqeYaRhP7UT0C5ICKq5TmX0
xv9nWOyQ3Sgvy7S5rJ4aFZ6WRLp61dEmt/zkeAVqptduSMNvKgp21wJQL2fiv9rah/d8cGcAlCdT
swvxSdosAX8emRszZT4sIsj4dTfxRY++GF7+5sV1Df5so2LO0oGbO6G5l0dyLt4rVdrf3Z2GrImH
FZlT9OVRYCAF1HjF2ZrL5hPBnytRIEP3j0rNcl9eWGRwGm81DJSVNGOK8WaHv3NPNKZw8AiIJObt
kK0Ix1DFuZsRHrgZFCB45T6TkwUUQqn5B3PiRmQcYHWqPkk5iZ/iH/I0ya20KFuD67vIIYf4Xzif
ph2jetJJfQKrQXBwzgWvzJIai4ObZmNXX09lewXdzYM5cu3zNoVvYj1UT+gPhj1L5GmWi3SyxqVU
ZlFg9N7qM5wgPYg72pSDUSxhAHdt/ZEOvpMkPrrOFpyCQ7MSP4swTytUMBsW2C53pVZ9XKBBQRPW
+3KVZ+yNTKHYDki6k7isQ17xRxE8Y6OUb8vg3RYFrMZeHsXiskz/E0O3lktfYNoBU0fZlPUNYnCg
MCZzGHD52ak05etSQBCvoVGhf4T4VQt2n0JBY6Y62Nk1Mx+cyPYX1AaUIofh6kP8mh66qB7pXe4U
ur2gmB9KDF1jlUGcXrzCqlwkKcBpn+0o06NpywO/0Ay7OWa+8Mqrj43n/96GdcAsSwdktBinPneX
VPhq3nc3YKh1GI2y3Q8SXQezwTsbyjY1eYLUpxI/chwGsCurS0otwDqKVa4RMJrOhDRTbn+1ssic
hHkZ2uPnrhg7ksnimgcDDIdHmzBxeMAytux1pKO+Do0KrdeQYTY42ncl9V4pkL1oA4ZpQSTjRpW2
tFOXia5xO4v2+iqvmMy7ktxgHCAYIeApozDFGKCRva7CHhC6sTlV3ADxX1J34i+AohfAEtuAE3Ps
m82ERPeA9tYCV/jo5rOS7O15YAwz+50ag+4Rk3LyelqFMLgYMDy18JkdzPSfeZYLALGt2q+Aaz6o
nZzWo9SM5DHNwMurhAkI03f6n7Fmy0KviRsS9/OAcICMCCNBkZMArtSUBJTbPpZo7q9bwwuoIhDC
ykoW+gsOxQgr52SNVBoQK7O/2zJ3QyqwKRntJQlkhjV/QFVVof9JQILGfRNnWtwfcjFTFQ3rk560
ywkw0wb67j3v9938i2INMyw6+gZdUXhHMTCDKeR9vJ96COs9ILPBdDgWxZ4zswv7lpxuLJYRpqOT
/JeqGgtcc/TawPNgx6ohjUplMjZNWDP7AIwFH9Gj8FCK397khN5bU7xB9UmTFl+34AR/rhsqHzWX
HF+suAJSwtr2eHuSYY6HtTFk1UlxLg+QZ163cq1bLyZnKtw05IKQ/VZ73WtJ5pN78S+xHv0XmrUr
G7QDnISckn8VvTO+yLAhMhJZ7gJMDvTuh2hQLOhwKWzjJTmqluhUfm0DsTmn1wvGxIIBM5EdJksD
PZ4EQE605aSG8ySi2vLxv/sA53v5ZkCUkaxh1u1zySgpea/rHVmo2U9F5rufS6SWB4PkKuX5SDuF
WaIC8W8HFFVaXkRLvhX0ng8YPUwVA/dZMfLSX5xtCeG8LfDaAMBzGnPUr5srIie1eVDUpjR1S5ns
2LjNR/bBtXlKopb87c9mrmWbPwMIXiohsET9dlxd83Aeth4rwCTxGcsD95ZLbChWimfU80r0YWIj
xKf+P/4k/VdVZQOOUnIdIsq1SzHukeJXW9zpb6xMNbvzGHrafStPWrMDqvdRncEK0+/hqVyNMOuD
bLJF1zojik5X4sHGJenj9PAppPxwRbTONMeTZ6n3owZ6Z3hPFhnvWzGa5Ywv2AKmYsrl0gqQGsrs
kwCBtpbXLcrxFfobdDCNLATjQj2TmzXO2eNDKCx5W/j7mXC5yAdhhV7NM63382Zc3L4gCUA5994N
9epHTTDj15tunyFo601zqDjMkiT2J1ICWQjmqAaKzCe2hYy9TwV9I3F6Wqeo2s49wTpAyS3x2eU1
OFCE/R5UCCuXJPyOVhMEACe5PKGklPUcZFcEi+U01xh6FcgBni97vlTSw2wwBR01uJWntqQjU2At
55U+Gtg29oi1l7C1XEdR6E/0qN0eL7z6wvzRjV2DFRvwFo2JxDLjkBqEW/FzVYHzIF5syaYzKBWT
AO+qYKvsngi2SpiRa5QqnSuPA532Y7qe2Ukllro3kjQaLUli+LTaAVrwnh9SK8+7ix1lJrQIooph
FcevIZKYA5Kw3s+R4OfkjKLGciK4wkyMBjn3q/xbSaznxb6ypryJVVBM2AOOOBmHh9Tgp23bwoug
B8DG6CzBfnHi1/9rRMdLJeICfOJYRGmlpx+Qh0c9e+2i2ieQ3NwAjWuxd5RNO3iry+ip4fVZy1nc
6Ua74mJ7elWybkiMHBKhcE1Tke12vIcB5MgewdaF6ZDYJQfNJxKWdtQZXUjnL2lkdG8ktif8sbkz
e/fBEfJ5OYvDmf1maCAOD6wH8KIgl/f7vZWS28dMCocC1MCJCxcMeDUC0eykugAHaVwke9yZTo1p
YyM7XrAer67BVgJ35GWi6CV55g95WVfq0FSEcnuN5PelGw7p9JvIInmMKdG3JPxU4h4qYGHs0N9y
O9nV1lVjE2+C4prI2NezsqCYkH+B1srCI2KjaLq+kspmj3CK16b6ey1RI9BpGbVzor/9R87l+fE2
+at1MmIS3vgUhX2bVyRPMYabSvBEKPtXUcTlxk+3rt/8CNMMLhPEfVsv57szsb2V7idzcEorp8Pa
fd+HBGs6a80NVbYs33W1SAgicwsx7Xc/lMMa6IUmidC2svzBwgNrIC8XZgQGvNcCBn0/IApSIj7F
cJ2JlXMVQ87VJ0uInhzoYNZ0nZIBNyggiVtQ/OJai4HbPjzwygtcEouExXGI/R7OrTZQ0QXmYb+c
2l/bg003JdGDpZedJ+H1tQDl6TUsipJ6+JX5lGIx3eRfqjEyZVo7CSgcnmEb8mxAnBTrOeKNNBvm
9WHmthZDUdALR8hyhbRgnJXKUTkyh5u6BqhVDt84u7AmnLHW6bXVGzbH2Sc0p8FTegIjOwQdmEbE
I5Rjo0PeXl2zvRsjNgsaqFZcg3Vk4tZYf0CGLMmIHWyque7yBEb8hN52Z9QgwymBIuuJ33Xbqg5j
1oK9hzx6W/X0NBGlljiJ1oZB8+PaTtMkF0CHeZ5YNU+uYwMDn7JASq+ZJFj4/8knbDzqp/bEmMZh
6zWpHWna16pob2MAcKMTDuLB9/T/Amjf9QxDC7S23foxFDRFFVZoMQ3h2BUu0R21fxkQDk3XJlAQ
xirzmYfl07683yqR4E3GXZSwSqI1VdWmvijp3QRva3znwxDtXhUA90cL5X56WeRhPzPqfr5oPLlC
3nE1uteAH5U4nl2XsF5PTDvNDc/tqF2VqA4UdJZrhrEQRtXmb27lZZIjC5s3N42T7JDBQTKUW8G6
PcqDUUUAuTzuVYS7h0Nj9X7z8LwAZuVPj4R6mdEZrxC+QL8ZS/NShQ53xI2oc876FT39JjKYw8mX
H6Vts0EUVMEyTtOry2eL4c30SSDZ3MGDQ0tMu6BDOZbWYxgMwmuUXi8TXAA2s0xaV+SiVRQH/UR3
VCTgWWYyErHntAuSbumWSAMV8L1AJwDf5DQl5myqNW7lyL72FWIbAXg59Be3uCB0e78Nj0HQrbx7
42ud7yzMkqByLpmHHWhCK2B03BYO7hFW1DxhSB877Y9WICg0YSHgM3ykI6LNyY9MpDqf2O5Ottpy
0y/EAKW+kW1GWTHqeW7bnHK2L8wS9Or4zK78nF46ZKX3wbuc7jFm1TxYo7IfSUigtDgMrb8xxPQC
Cs+GimvE7a1Z/JaNIeo6Dr9LhfcRABKIu3BelQZa0zNpMYQUEF960EoTF8rZlnXg7VFJ9YYBjIoV
Xu2Y/76uI9rdvqUkuh9EdKszAoOCDyQOr9FSqz1H9HMMlpsLOjEBTlqT7d1XH+3fPFDvEWni0gv6
iv6D3iP/1nRLcheNN1sDAglfthf64hskR8f+O40tolUZFEH9vIuPfGeFbaGeS6tcrhfBh1AJFYvJ
CRTVcgYCCt6mCcsXB2U8ZVas3BNpLzHOslz9hEfdi10sJpOfv4vEKvvMvMoN8hxMPm/KcpzvVo0m
I0w7TGSsvkYSCJzaLhE/2J5glItvpvU+fEG7bGcu/+m5vH/Mfdag3ga9wDF+E8+8r39mmgTrnwMH
cKskq+p+Tnz8JS4klrSIajOo6V3akzgACFOsbojHIH/ciyWft+yht2ssDOgGIEKFWugsJ3g4gpom
xxGPOVGYWWUMZU+Z4GF3HWrM+9e69Epr2GarcCKHoZ8/a5HXn8UdwhG4OAvezkd12+qeQbttoZvC
E9+XW0h0KsKYJ0gvXVaa+wmpnAtasj94G8Js2RgU4TBoRl2JNHTVxVFcnnBiYfQUaWIP57fSGR0r
Qr4NLeilb6M3WKTs+F80YlQ9asZMnCkElUAex/HH0vJcYjSSSJZhwBGBSufnpKCIyxfhnDAEhgHH
/XRLskP1V5crLgSwpV909mUabUyTCTzr4s0tzO5FpNUTzn1vXCueAL+oIXvCfFa1ITz3f78Uqduw
AXQ7XDOeLAux53t5quLBk4h3D2B4DBCwNOpdyBL2xZP8GddvD+Sa7QfTQkM14ku762RC14EkZGxH
Q9DSbSwTVGtU20nW/ZA2/kBuJCokcI8tGjuUIaGHN7yHSUOjqyoSGRwZ3bpn4Wx3O822qgdLP7oR
lmLjQcvYlvkbYjEZoxXA8mxn/BN3Z/q41luEAWGfIbpCSL1ydoczqjfehYIOT2Dw1/qN9Ya/43HC
h8xR6FbmIU2jEgEcCzRXLiGIvLnNea07eGUk3ASawz4bE/iRChiZWhib+KQ6vlxKW63JvBXeA9AQ
xRG5eJqU2Drm6hjHVIeL0ZWxUDm9se7NjAFES4HtY6atyUs9bhi5Ohs+Xzu06vJe4fDz/mtz6sbN
YF9D89ijxVNIr/NhXvh1/h9fB/rFsD1Q0RS2Kg2GGc13muzxwcGkc80K4cMeaHAAqpqCD+7KVLmV
TblMip2u8kX3EMr241cZiPoFdyLYAii3emFIoWHdm/Viy6qrAYfTOhCUigB9I7msxPvM0IrTol7W
dovV6mMTGrs32ZqijjvOnY57atJgNOTUWEnPqrKAVCpuhW7/0sfWi1Um2sodxsXP3o9Rhsfglk2K
4Kuli/V8QMc3ZF5cv4kEb5diSYEuDJvobL/WxmasvuuckaA4lpt94JItUvsjB1FSmnd8LHAwaOwt
hmu6orsR74j4Ki4V0eLfkHExb6MF2a/cNLGDyTsy1AiYbVjdh1awigqV0ceEM5Ie6F0/17HP5KHo
OlKaGk325JwfSd5zLwRCdnWsBp8rKABSGKHzmaaZv2OhXwafHa9Ve6TyKiBKgPwCc7tmRvffbKTU
iFKQ80kmMaooOPQS64vaVPKW5WAE01P9IV3tj2R4T1pEVwRjtGKgksW7qt8Qtp7W8K6ZsvI+6Ulb
dE60cNf7gGuKr431K2L+nAAp6/UUsEcJhVyvkkuzEw+v84lvYiG6MsMC+bIpbI3GhG9aNylUHKjW
TIVyuUXqimC7FQXCtNI1HIk3X8/997mbjZZmrAc+owXwzSiTrXzOx9TQs11HgwbqMEyiu4KTGyc0
1g4Z+NGfQavUeUlEdaxp5tEJmiEP14hRch9hshAu9n+HdGb2JK+8CRoCEycT0BeqZ6kEJ6T8tB2W
au0bOMaPA6jCSWr9LGKZ/AEEcm99g9GZyRNNFVNQMnA8pYC91Nn5DG1z41+znnARljwmFwRm01TU
Gl6DbuzfTG9h32GP3EtxPneotdOAUy5xQj8FthHkKeaxoP63oZIQL8XVDsR0eK/WEb2HlFWC33DR
toIYIoJj9/ldiOCRDu8tGNrBQmda0fc1FQkP8HG0dOIL7VE5rK4F9N7/sqFHDX130r6XVe1lNpZr
9BIN5IID7nT1CjHwfSWFidVdyVp6RHSZ4DdxLWwZmm4VnBpPXtt5wyQrO9Nku2Z71N//BkScxOsn
X8wTvjtBTEZlp1tf/xmGQmYC6BYdFzaZOGQrv83j10cxCAwVVJDLciErdDgU6GBYKngdrNC6g9Kh
iT7Z+wXf+lJY7Ol8o1NZ7xQWFQvu8QdsnYBicP0dfz8fUXYYD+XzwcbBbWvablIoEBwZbffJgoTu
z1c1E94lOe0dPrGoM9Zt81qrTPRwShgJmhKeXRQ4kb163tna+JVzf+v0S4IiGiPMk419yZ/6w8qS
XAyLmuSfcu1DxAgR/P/60T0gBKB8GCVPLz/yy0e1yDTVploS54ahJX4JfVW5GqSo0Yc2Pg4tfyoS
0Y24mK1fVOG71dkgM7KQhi55deincU9WGTXEDPERqXG13UEdwjD2ZzhV6qSANj5b77BkSaIgSZQY
Zyk1oOeANZhvbI74lPbPbKNKjiYxK78D6OrYMmBx3u4LwplzYYKlG9X69kbFOvRewkREUXfL8O9K
gCxRc0+RSFT5Smpds18OqPvQp0hA92VJlpr6/mge+Myymnmy/BRRHGg3V2Yo2faHP8uqJSLZGZoB
5E54d3k3nViq+TrTUJt98dByLOtWJFpJIk94qPoDLv+LIhCal74EJi4YzK7oPpdvaviJ9xgYqy5r
gcaLo2BzLEdtWLPTpj3ambAX4i+ytgCI7uuY7qpZacC3dUUgkd1U/9iZLdv/W9JpqjO9ggxGc7cs
QtCvlUSsEr78q5B5j4PEuzeNQn+5TwQkd3zrlZFoNiOOGTfENicj7QfLnuYHV3lmskIylJb0y4Xg
4YVN9UiNnw8JFH7aHSvf/byiDWjyKerB9gEU/zTvaIFftz1wBqhqX7LjCKH/inHJTUzI8aWQuC7Y
40iXhzvXnO6MfhyspRiFybB2wfFVrlDwaDqo8wT004qo8GFJtG1HUBh2xEt26TfWUo5B7Wx01AOa
yrEVlKcxTJp0LZYN57Kg9FrYgoilJwtKWBIimsymjkQPDsNtiKDOVlH+h6RzxIKqZ1CYxq8+Wbpq
fMTCKcNbq98acQuVA39nIsm9hAda8tL5fh96V1oA4K6TCl0qikbMJdQXWir44U4YaiVQNNjdp2eW
jXihwKgzcD7UUGcZr5g4clF33ns9d/SbPDfRtGBu93mVXahbfk+EPyHP0EyacVeXO2c95cHbDKov
Ew6shUYpSyxvdhlfRCHSErqd6AAhaZVMCSTdNRqPhbD3plEN3hmjiBHE0ALPr4M/B2z/QzL46bjL
JP5hCzwedBuIyUVcEQCWbgjCwZfUty6DIAhEeGm0mka9Sx0yTrLBnLTL/MvBklrSQlyttecRdtxF
GbLiX/XVUPFtRy1BWtjqK3iLmlsniWpknVxDlEWeNR1pmFndPbWnAi2cwLTc7jKD/N7U0hqj7Cpk
zH3JQkhuBKYY5m1+pF5jOJiTVzXiTf11Vl9PMZzPz5qCMAutzG1/732RjKzvMH2mOssaHcIfABHe
3gBU1lVnEk0LUxKDVSPUcTJhvfdXW6heregV6ClugVEmtgTIbtjRO+OgULIcjsAlasq/ahtgbL9o
P/1l+IXco0RUVjIqieDMl6N4nt+0m+bm6ri0nNLhAva6ckO39cjHPFeVpnXJtN+0fZz7u8Pt2Qdy
KDfSqVlaFqkSA/9+hbvOMaWLJ4GTm0K19+iNMIRUztsCYvR0vaCQPvMVZZIW3KCE/v8VRVj6WEoh
jC2CD8XQuRfb8JW+rqkGbwFO+ZMTM4JY0yaBbHdxIF6RId1Welm7RnIvmjRg+viGUNGsUSNn32ZI
nxBBSXU32vd+WEZx4L/OKLChYX+SjK4jSOTljGs9SJtMx0B6gjy3XRqfZpIwV7HzOvMWCmkwZc+L
OsWnqCMgNxFtDixUTJ7HITsVL9zA2Nd2o10NEdRo/DHeOMBvRAu5ujHnTU73ZB++NpOIHN9p0+BU
BaON/6cn60bOe3YEP3rLTQHcw6zUCM1joL5+gc0PPzaVxAUklWF0PcsQJA2DJgOmJ6fjrfxoaifj
vyOxqoJI8/XDsIOIZV96EdJSrxa6+SKxJ8kIe9kBGUq6SWeXXexKKgYtV+hq5vNgQxD4s0MO8AdE
fyIWICwIsHwW2ykaUF7R3kamwSmnFrSrRxGobkSIBpn7drJJgedyX8TyU8yZkkrdbtiAYRYR2aou
WWVSg9IEPOIDIm9lf548Yo1OjAzN7Hx4B8+qwpXtZL6emtlh+synlksdFNXbDGSEGB4veHlDyWjW
iDDVEuabRV7/ObuJqAvrHddRM8bRjeXoWcBZqxWpVwXY7VXY5XiUuELR5PkKJZdqnHN2nHOe6kwB
Gcnh9V217UF3hRk5pBI+l3EkN6Cu7+Wo25aNyJSH3fdi5QwBFw2+hbuSQKe5ct3wAsD1Xsc55xwS
KCGZqPfUjY6z+Ob2oJ9XU9H87NwFgQgBSAQr0MMaYm06USu+m9t7U4svOi7lKzGU84auE7iUkpAZ
83UuLvLsBfPOj7Qfav0lsm1BlqcDPMpFTuQZkONXAV9v4XQ9CSDMoORtc7FSS1nfr7fMovHz4gBJ
+leLFpfFx2iTlE4QYMi4A2d9FG78+CBsYVPGHciUX7/SIH68I7qEkht/RfbRchFz3BHGv7RTburC
MeBk6/9QjQ8HPAtTdLoRtWq3PE1+48cskFF/c2Bsg6Jfqp/PVt4xMw3oug180oAYRUAJtyGKofLu
qIwpN5XRlhT3ytcDxqywcbKHT0WAekgnTpJIEoxj5xxgdAYkh5xJszJHHb8Rtfo8f7sEnb0ksTHu
LXi6zyY6uvGGX3jNXKbxPX1PKAJ2HLlX4m7q4wtT7N6hO7KTkCe/LWtjYSs1O8HdzTiwVMjwynAI
vaW9CL2OUiUD8U8h+JyNdTMdmaaTsMbqhMuuOE2pTL4oXioYdf9oN3nUtkRptn/tvqi/g7HMSzbW
UlKNx6zfTUS8cJAuB/l0GHOAApAsiyjZOrcr3bBOsV9F9nQxbwODWOyFjFU2fqj3mYjDycDcmZ6J
hl//gY9U5Koi1S6EtQUU/C3/UEm1vVSZ43UBiYXhKSv0s9tPoGJRnLmsXdKTbbyMz/DeLfI0EGtJ
T/u47gSUSnlfXnwF1h0JLsT8odzDCLDqb44rIprDapnGWyAcm/tFJfMQbCRt8KuyXdZNeLfUyncN
+LMyJ4WLILdoapKHMXTxBAMbOcl3DbB+K5JPZiMR8nfQxDhjMlN+AxFrTgDNSOd7FLKQUxSiFUZy
tR+xtnmV9JQSLg8dvDYlCJGtnrNS9jwFf26Gv9QbzMWd+8FzgYqCwsXnLL3xDoy1czR6p8wbjv8A
mSwfzEyM97cNGQdIxyzkUNZ21AabM/U9Lif4mlsbjw/Kz7FlJuln7XehdzT3zl2yyw3095x+M286
WdxNjkLOX3eETW96yzKIvHkp4nhO+0QyvHPyaTAS2OOcGuPnTbcOwJpztyAykC5Jhhm2/bVQ7yYh
7H+xAw0lBUBjFW4PXGqvJ8kLZNSDKB3pHLSYJO3h6Ct5MOmcSjgpxfqcY/a3SkmX0cU+Ywk9yvmG
FT63BYA5MVm5JfsEw+/9XVjJFolY2ubm45uzCcu6/t80u6i9vipR4bjMwP7SOB/UNLByXo85tm7W
9f8Y5ZM3Qp/RfA0fyQgjjMZP0Q2TTfKwjkxvCoAKp/mnTq7XOIunPxv2QxZ5A+qA2+MJypE07uuy
g3vyEeHRzr5uFcYKXMLtceuoZfNQ/wyaoABLhj7WgQaCyeetEFtg15nP7e4SVlFV9ZVgXALoZ5ap
L7lq22Fpu+ojKWK9GaaevHW32nx5tr+r6xlAK6k42j6upX5SlwF5ThVuL19p8/OeUQJ0zXuS3sQ9
bY18VKBaoZOH8PZ+0HSQgpt7wTP3XWjdUtfys6y1r+8EUkEZjKJjzSiT2ljTBRr+KjrUH25QHygW
ikD++qL09puKCM0/LbZPkUhkPvZEniZ1QHi+zILUM58pjhD91kv2fBEaToEBLEGIKZxu2GYneQct
5pHBMrQ5TEfEuLkyD9Lh3cCIcVsFGsRwjiO1NQ8UF+uvSWvjDqMDN2+dm5oQOVvXyFJPHouSfYtP
Ptq/c2WA/llH9NpQvy04y9/7hXZsvpCQnmmcdmqfLRk4LTygqY7oJoOcMumaXwMkgXxuH2Iur9wW
ZMlM115f+LJeBk1bGV2akXQnP8la9Fmh2XmySmzSQXcxLme2oLag2MCEWRzzt1lGnA3pZK7jCemV
n27w8Cg/r+pb+wo7zAhab23S8oZLESeDUl4qfw4r+GPYertVFnG/JIuD30ELTyLKID1X0BAL5CFL
trfQNdHt7mHRDFVL+2kbx5CoLXZ6KeV8hMPDPnafYmLPE8juSDziBybsbYWVYA9iLY3/ah7NVEv4
GFh7uWRkDrotfuuZA6mMK5aGTG8EvNRkhf4OhUHNRq6zA86igkttry70c5Dibq0fAspqskVTo3TF
3w0PIsDRfDoCIpy2zObMFYZi4005FBx0jBdxS4Dl3P0tHl8Mri4aETeXFYZkeo5L/uu8WF77Lqg/
X0Ab0LD7BJwOaDG0yhxXf0aNvA7Ej5txaD6UxvKjUW7EX5n25ZPq8Wwb9mvNeryCREqm0/68gF7t
UZcQMJn7MDNLWmezGYIWtoPnwruycwePg1NY/kyOVNZbSaAtSdKW/7bFgbpWF/QcwJPxTgsZEHTj
EgTtoS8zOsJxYdAIaXaCLo70aJGT10tVs9iPoI6KJ/KVJTg6ejmKDkuylUl3jh2V5ce4yaCP+ZAP
TmOiXAF033dGBfiaGzgZAbdhsYLQafE4p8PO9CTuOlT4pct+eeNrp2fZDstjpW1meyuVpqCAziic
Xnn9hrYA1HuNk1lCRNMKkCZc5+Hj0SYm5l4zZ8/AMISQAxHFx92tm9AegLyB5+IAqN8Ld05ZjvGO
nQloSNXTADysu3d7FoxVq8wHVoGZC3xIobVeXE1AatkAdEGU3z6zCvUerKOjUyd9nQ+rB9F+0w+V
wFPHEt8HRH+b+hJnDMwo64eZE1FuXmW+xKGVz3YgeNi9u8lciOeTjMI2wa2voH1AyTxElVU6rwmV
sn7NoDg5xQPY/vGNd7baJ/jzKrKlTgRJgz0UgmLddykU+5No8LU5XuFfKVQInD1/THvX5GgpFSyC
Z9oFCt/zDfnz1CA2S62rejXrv95HWitaw3+lA/UTapgU5clsLbsEo2mh6AgUOhFlw9o8VG0CjJOe
ImFmyoFq5YnX6T3GP7h2e0ZL1nEom3MXaeXn0a22sPYkndxHcYWW56DfryLQ5bc/HT0TJ+Z5OYgf
Zs+zABCnLjklcO39Elb6CAsycnW5oQlf4lNnQgSMR9MjivhHiiklWTrvWrwUJy3vt+63hyj7CSaZ
rbz5BC6l2Mgp8WysEJ9C9pJg5Q6ly79hl3FvC0e1VawXULYMimXuLMnqa8j3fsEp+CeOi3XsVnWF
Oy0VGBNJYG94ZAMy7kj11RML6SdQ9otTpYS75VwxkNcUHitFi/njuFSExqpblQWm+76x/qIRC1i/
6DrVYYNT0HuyY0wF5vbeaBHV94bAabCfD3dPvyoPqBbFlAhUcngB/Tz/vbIfVAbxp2BnDE/Jak2E
VrfFV+fHBvsqozjE6jaBfiYmfTlMuB0EsHFdPZEbixtG0KwRthVWRKZXBswr1SGaHwTzktZ/h/e/
kcZORXZ9Vr9kVWc/roe7n79sc1XTnz3vPP9spK1NDUBStKwd2/cZ8+Atzcqe1H5Yq65vve/703l/
HrZBikY/pCc2QkhcVlihyEkETVeLg+Wn7s6BaRZqw9nrplWxoujBqB64fKGRqRTGNr5Kwa/QrJ4L
fPzNZp0ovKjSflBw3V/DaxeaTI2Axg4jmjl4oth4oV+rVTb79//2tdRj9wrh/JiT2iizcqKG16vK
QqXDPWW3BTPvRVUUgnAgImsv3hQQMP+d0+DtAPKMTq0hQKpfUZOWTbeB5a4Lg4eWvoq0Fl3KOy5/
RF0satBI+ggWV5LCdnOmIaEomrv8B4vODOK0qk1OrB2g/NYdxsOrLFLRBoqVUII5xgmnrPan7bOs
OHYgsxq0sm3pF2Nb884PUPnyPHrRiJ0YlTqESPgDjjCd55mrDMhaFkBhGro0BWTtBlm2CRohd7uT
BVuTunUkb+/2FxgVsdaCc+f6wDZT1RoI3FmO848ZlnLQoOeEOlXS1gdutQrvIEmcnv8IUkSEtfI7
kT1ZMII5+ewhsYIf3Tn+EMubbAg6ciONkWGxmeWSem5/YsLwmB4W+Ek6vUsZ8CL+6TGeF+EKY/Jz
xUxnnIvoFi9sxB4VeFWt+TwFw4SKCyYk/W8uvtCRFvsAWvFTC8zzoFHkdjc0Dkpf5JHfgTL64wtl
nixKTytG9/JIZhtrxhomJv8YAc5xa5aEvTfjIwTKMHyZc4/RM8X1MOpfsw5VIBVDd9Wf+/rMa9fe
bXUAnIbYTeX2QB4+1N/LiB9R0Q91sW3jy5ib8EOvH9etET8HNHZJTO0ii0Bdlu2oQyP8XCJ58QkP
JNGVvqqMuRYFcQlEWOnIJjNMvS6W6mbvoYBkugX++dQHqfxyhtiXmvCcUhoz1eG/AhQYy/ByCWlY
APzaxj8eOvoZWEL+WWDEWujya2qkBZi1S0a8hjtexoNEOSRyqg5iX3hrDfGbT0JrGS4P57qTgn4t
krhleACXwOHOT354YFRodhuJwNwlIUFP1+ZX4Kw7mz7L2taFfHod8GWGhiiavTEnCNXCCYNCKg75
IXSJHaSNIHfIaBBggoNJNCRL3QrQP6r0l2agELKsUBPN/4pN5E/MeC4ab1GBwNddYVYFZj8b7/z2
IwBhgg3toplkd+Ufgen1cHGt/JTHJqpvcMzVIISWAg5lBQ5mRrZ5g9HBS1rLutOMsdXryXP457Ru
2Zwqtp9ZctlEF5Tr+uJrazuN8BBKrg3yVxFF2Fk2uHUUqUwQAj1uZeCSWfFY57nq7bngogUH5ysU
qBa64VH4Wz3rNGdf/zXRkrXreua1cI+nVoj+OkGhuKfQhB8gM6hV/RU6RJQM1xKce4MJbx9wDWz+
Uch4LV3x3w0aWvz1BSp1yBKLho18T48h3RTY1fOl8kf9aJSWbo5bPHYzmKeQ6TCGE1cguRJpIYg4
2eAW+DbC3t9TsoI4zf9IiWsb+HMG0RSE4W6CrLy8z6WtM5vUqE2rAbxaUdGPcomzs7uyub5TxqNs
nDVoUoDiqaV0HAK6pUwFgEYHrcRhlLIb26noEHOGgO4k6TOmo0AvnhMw21paFoRMgjybK5YTxzQn
+dLO0gqIF1XkxRju63/+UXAOl/v9OunkvKO78bElyj77twSYipYCxUMZ+CXlQBTzII6RnUs2TI0+
Hh9XlfbotwWG1t1lS2Y5wXzRAXO65SKjq23U5ATYIQH4/MmuTZ+RGYUBLNwCjCL/6YAM6uUsEF7l
IpPnGwJ+0q/uOrWk3Q86yOgYjXuq25ASL6SleonyC5Ia6SolHiZhRYpbpoI5T8Jl0mE7BWhINbZU
WMlx85Hy7g2Ej6PRuiKwldSlNFSx1EMGwaLYbqzF4mABjpsALK6AWkc9jE0iKchFcYUYTYnX1Tw1
+HM2K1pXNxe+cQD4SSCPsOjQ/bHPyLRAyUoCJBxnH6lUhX9SWZhu6OCrk+0ePPnyxj4pcPyTOucG
QzStgG0van9AP9nx0ZaFtJxs7wX8MEa8C/xMokPJMYLkqPxEjKChMORb+5fXRoXi0utqrgnmeDMj
X0XkUxV4Jky0ZsloW8VMEKLfsAR7D4JPScwnOOxbeNZdpW1sb1is6iRY7wwN3sTY4ajRWu5PnUEK
AvfP8nUz9xpCnG5fqJVdOFywCXAHnF48pteF1qgFDecjKa8mAMduicmcqorYak+V8ILm28c6GwG7
JMh3WB0WkAu8zUvXDRnxgfsdgLJTrsFyE85OwCjFYeWG1RCDDFwPuABb4XTZjXVJUBuXRs3pnTSg
VyyuNn3HEgYRJR4dVgOQNWGSK+alVUNA/e3xE4pjra0l5YidG3GUdj1LRbWPUHW1oBpRkblKlGDn
luvfFEKu3PCsQtD9b/+qEWcUfSlm4q4PjJtOdiTD84IoVybMkzYpxMt64WxU57XElPLdrWuernH7
jnvHPG2RDSnw704e09IkWxNvLBv267pt4TTpi+sCD0knuhDTmKeRAObAk5oYS7kPBxe7FVsdZmzx
zD4C6BTrP5jv0AdCyiZrx+Kalm6CU/I8c0Uu4J2cYUD+3V0HgOSr2E5Qb0fkiQ9R0IY/gJCI9uMy
VNrCcptvG7u/Gv+OAt25nARI44UWEDLMQt2KEfQWCLwzNe/x4wG0mQdx6T3dUT0jsm2BWde4C8Cj
SS61H1DffvTiJr4vJsWFoxd/sjTZAHTwYfZdv9uTLkbfcxcTQkBuyqmn/5T/fME2F45IHXNC394v
8E8r8aHx5wZwtF6YPR3LZz5DCp3q2kzbnSF0S5M4lvetmhX2SkUI7zh3dEICWdMqVG2bM3SlwSv5
YgnTq4vaaRGLl/nLChkVOmasjXsQagdccP+h8gSx4U1yX8FyeAWyfj/g7BSqt2onVQRwa0qXv1zo
fpTL2PKTPCzmepQL5ikfp6ewKOW+etFQe6EgcfflRX66qI/dmnHe/G7px7+h18EvP3laeeKTNFt/
fgH4OzYusKZ4L2Ipsz18mT88ENQKmuLdYrx+gwWrDsOBpNRQelVtgY4SiywUHf/uJnwIifbJh8rH
xhHldl4K9rFWliyz0k1VeROZLU+5wSNGEJGTXSZk6JjAmfOgdLJsRGWRhtX/eLaVva3Bdk3wX7KA
++43hFkKX0KluIw9w9XrOhJ7kLagfdpSYzMSkHk6CLQ1ugt91TFcxF0gIlUUxGMJNDV89EvXGhYI
23TU7LH4Sv6SLchVx8JtSosBS/vVaJeY1o9tEfN8v4t8i1Bjom3WpJergsgmoBk1wyw2TiUb3RPm
PQGwL4dyepclxJiVrnHXTmGdiTyHWmdNgzqDqbmkKCvxswlyGupDIzg9iQllEkMP03nqQVBWTQ4J
qxbAmMT4LPRMzcpovqmkP+p4v55Ky2lsDTCmdPfjz7L3/v8qNNE1Ht9TLvHuLMkY0rMx9q1iXa4Q
pO6YHzwiOoHVbcmuR38K634Iv2TCHrb5sAGhkfMWG2ik4rzV7rrRDUET2IKpuKiRM6d4Rfq2vp6t
zTQY8Irmvzy1lT1nLzJ8KK4H8TLl8x4ewcrZHfRMCAp8RvTpual5ZjUV3csUyCRxemEARzk2gmQj
CSyxiPHNcexaPQpMUlE/B51dvXar8toni0ejzffUzJCMpdRm2Skll/QNl61GfynlGyS3W/msQim3
HpckMUzhUygQSF5rdmBqOzQgAWvrA0BzgQgCSW1KmhsrHKduzJymniiLxHV/vVtdCOW2Hx9Wfbnz
eq8k4Syid7SZX8FK4GfOKaLreqAh8Ga8cPaQKthyaM21ydsv6/GmkmFZUGp/SxPMn4VhQzuyemlq
vlA7njCAlpVjf8Qhqv2eutNN3+NMgAChzUWoKZzB96A5DROnMjLF4mpzsyrc6S2FDYWtJ0rBWRxj
Rvfhlcc7mW9Lgi5SjS0kfXHinEUWScwV9itaw2UuOUS2Bs4E87clZpmOob/qrKDxNX+R4xSHHk0N
GnQg7/NHLB79ZmW70NhEhr33HtuahfrAbXPuhd1V/quzk/5+Zw+2QXNh+wMVLF3/j1HqCOaDEazy
E6ygLVvVgH8Bad9aY8bSemXt7aL+dd0dE4C6xqVzrEW9BAD6XqRWETBVwqVOiXFAzaEWlpKQD+kz
5Yzj5IL0xthIkKAPA4T3OciIi5jxJH7GAINIT8XHZ5cq3YKQ01uiEePq+3R2m6YJ7WjSF7OkmN0a
GA08KrpL1osjBBDiJokXTnOZ+yrV1OySoCoj6J29q1fBlAoomb0sX1+Lv93cpNcr7elgac/uUC28
a0XHwriBzkMrIYfmgUYZT7y1wwyqa2xARKh3CZKg2JSaQA/n/ViV1TEmyXdb5yxYTPeD/gFd0J/b
fY/UCFO8gLIL/8a3I4OKfYiVQi6RweIZsSJfcOWLUER6HHJHx9yjUZ6ZpbyNTtOYeBTBGmyK9T5I
dlwWOl4olm5fHtaVDSS/6sEpCqtIfTIw+3fDsRvl+Wi0YV124KTGPU6i1lZIkGCMFi/6hE7UDHeN
TwFu/9+JXhaVENSI4TXBVt7ktQPRujKBXy1OwQavGnQ2pmJos/cKx7ye2+L+3cdahoOw/ThMrW43
Q3yKZNe0G6zI8WphwO2/LhdcO+u+TuW7op+ccKkkw+/koUBtT50aImqm7DcAOInnV/ELa2c0AV3c
EktNrpKtWx8vnbX4WjZ8se1GE4szrQIphLW6X1hAxyvPYlNWsMvPYyZpsaxITVJUZyrXPcuJgEpV
9/jR5i8nIpQXgT49h6/MsvivBuEABRYGmN1MQWo5xiMQjJG6o0j1nl8sPjf0mF3Lg4rFXeSywYD0
FwdnyQFH5l9KMsNjoGnMZfy7QVvCBrV/0zWuM6GGxgnUgJeq3Z3fM6ZkdqRb9SZ8ttnu7rWy6VHC
1SbkfU083Ji0R5yif4MZIhTf4b+yvpSBtWcQZXHDvrfCdfE5H96DHx/0/t3C90JmGVFhvs02cKka
JqPjvijiLd/+4gq8rmJHB/ZN9sIC1xRQG5wpZXzUgps/881MkQwHRJC/X+YInMMFxDzSpk2PwGg0
mIL492lBS0DajcmLLbYNiCC35FYEYVPHFr3NcWszPX6OZ5XZkEdB5uH8U8Z/tOm3ypFISYiJxhdm
WQDMyWM223iDfZnRIV6V9OjcY2sRk71mAKcYcsm2JfvYn5ImrSUnWPyHngJmTd/pEOxAi5R4Qkrj
WwFf18Zt0OmThwCWafLOBnniwgh8uKm70RpVxIe+XB55F8KmGYZQ6s/dFY08Hq2BdTV07GOvUiTE
Uv2B1d+wsPCbIw+DOevkpWVeFx48Ll6lRBFvDOik51jHesWhqXg0bUuZseGAqCZQLeDj/ID3XvQC
qQisqRhLIabcoZkUICLz3ms9sMBwtrNCy12NYwiwfqBLmeiZvxlJbHJD9H/Uko5jBB+pxt5P4nJo
8RAPEJLk4K5mB33wddysKH5S2FE4TWAwHS3hv/DfIsBP+WIcmZf0bPlPkojqhErRHUC/Vti/NGUG
xiiHt6VZQC69hWSrAzVb1w0rr53BkF+7mLBBmoHxCsCYiisLIRUeLUvR3+yGnuXfD9YAwu8IKnQP
p3xZ7ElVHPhJMpT6YdqCM1K1uXlNdnXOtdpvduWo4ODGsNPuwVZr3H4VfbnmI4xsc1F5xcFKzx/Q
zOlfbHV8q2SUh3CdC77tH4Yz/RCff/BLueHtFMBCQc54I2bcn4aznu40PWBp8XflcR2lAqx+G5j/
4bjjCwZOkA1huYsHTn0JZ5BeE7Cy7Hyy5xN89f83JiF86jNfi2sZ5OSDA5o1DBJvVIN4f2aVG38i
LxHt7wDFn5n8X8J0a0FtjJqzKJgMdwBrZ3ly/dVxIzkETjkJfAHmao2jXWLaXIg9YwU4Xp78lbsg
CEqQjqEEf8xVAkMdnzitibW0Je4WnABw0iHj6YF5bLs+Q2M8dIn+P/17/Za1fXPSffxtQMDJTXKp
edB12DzWA6lZ/rDlrZgeG1RgTAteEj73ku5FS63QcRkR+ctDIt2h0Ytnyclx9vEjaTBVbb3cy1KG
pMRJcNZSXvYVY0T6kAS8Q/HiaFR5nIzuMt4qgvagxdCkGCuiH8nHmh9oiF9AFKLdfnyDTzW5V4in
21aTr4K0cJbz2nXdoTx2mMrpM0VnT4Cl17yHkXa2jfdjwCaH6vescdK7sDzOh+x4w7gkH3jmrrHM
8ZR5J0Yg/3m/UCYXpop5tla0JvUGZzJRfZvpCn7BLnitsseG2IgKFugjLI2YcC+UMLJNij84SGVz
90peEh3/Q4jZfXXT2xgwImbXLuwcxvliOlY5Ii0pkR8SyxcSp5vILrO07BoifsNH1kglZ/bjMlhp
g0NSLeaZrcgvDwrICq5bma2N4YmlC3UYiAr8qa/SJ5i22nG+cW96xM4F2FhZTXrgvH/7EfeFLfI0
uZR9mn7ZE7dQbijZlTDJAhU48kuAv+3++7fCNvtkPVNMZHri8pvv/M106KQLDLyQtNjRBXyaNLY+
I90I7WjG9eJta6VXChfxqZMGxyGfKDM1WIMTJI/rHujUcgiG22h+8ViBMqNYGqAT/kr39ZQCuagA
5sC9A7aKBSoES5CY2ijFkAltCv7uqFgrWIdcW9bWdsjXZFVUfL3vbsPt2pS/yray9ANgofFFWoII
gjvqITItgCav1Kh4SYds+XzddjWUkYWDeWCFNnI8VZIEAFof71VNocc73ZxLp9+HUbH0/ALx/2ty
d0za743NSQ8+6y85vu+T3mGrhhNfey36xu44eLQQDHMoh1rSar2kq0Mp3BPwGgThya9RfLtQi1H2
HvXYcWj9AmlSfXDdj/t/r6BI1RfawI1YpoKUSLne27SQTtTZn1tQDD0gFVfA2zhobOc+9Th3xRZB
4F33ISt7rRpRUjZDoJooxO/9sXV7w7RCr2GpoEGsCXF3LMiTxkcDW6kYTwOglwF4islUg+4xHUAI
13duuNaDuxKC1wB8ltJvNVCCmj5cl4obI9BeZ+8bICIkbgmayO70QgLajAdTN/1gS67eYLa6xAyF
GI5xL/ex//YfNgLbzKBM420JhQSZ7dgbLw8egK99wDvEeDykj6Hjz5KZhMEVa3QdDIh7G9/uh6Bl
L1Ollor4W4trZrFSOm8/OnyC0utBjha2u42NPrsoVjW5dJnEjCL1ocZEAwtFfl7wssHVAVUFcjnp
6PJIKrKWz6oRcAv9AXgxXRTpNbNHLQrOLhUUOVozHsL8KRR+NsprRdgirmSzVCp+J8rsTsYY1kPj
TUJdmRuoOua1mCyPZAWjStkd24Bm2sPotD+5wekFoyRXYQIVagL4WPzXL6cDn5KVO9c/rZtPbzZe
qefHHQpmacG1Mlz34CiAZHB4HbVkoWhtJbIJBj00E7LQw1hn8TU+KjDi2grp6QhKS9IMiaXEl7+q
x/N+dIqsmNZxGllV42Bc39hPsCv6oiQRNjsHsENt0BgFtNfAQ1NtOnM3mF5q/C/bmalmzWIqfhVb
Ph+T3Ttdj1R0ex/HRYdFTIZL2F/y+rbHzaJAcWpItOwe/bVqZPIWUwjssKirDdKDMb6Ar+ZCNkNQ
TGmMg3+E6PXCbOQWp5aeWbQaeH9bQscOLc3m0BwndEn/b9pmbqJ1dtE3Daiq4DN8brh93UANcVma
3u8MgxRG5Fgh7FqzWC/5e05F5KzxKQXPegF+hOunV2JTFUrZFtQOpDq1LivKILfvP9trv8RTP4W7
enL6HjPaPr4RLfyztEF4LpmtD1ex5XlcPOyho97WeEwvw/6/nmkBEsoBf/dJ8qiWjFjmgdj6lxJk
Z51P0SIkjDlIfCprk99DQdl1Ier73q15r0u3/FlXdKIgKl0GVCBHyk5YmzTNxCPYlooW0sGXalZY
8/mK3HERCoB4auUfq6+NgdlHGiTaT4rUS+HVqh3gKBadurYFDAjAmrqOFqPHB0nIVivbZgcV4R6Q
BA+l3Fizh92CGRQUIpBKdc/HEOZZ3MFuW1IxVguB9lgyqWnTUipIK21GrwOUuZYr7tPi3xS5+r+P
q3Ez8M4NeXTT+vwJz6oJ+mOoQoqQ4klnomnvMBYxfnd9CEYnxGRnKiRYW+fGHGcjpPtTUEpWLori
rkHlUj7YH/DbpS4I43G4dvFZ9n9UjUC/MbUSEnskCwQ3vu42F2LcabdpdwnEFN9dBdme9nF9Pu9t
dt1xBLDCIrya3OViTa50vpVNCKb6xhV521mEZ2awWfeEfgOJiJAMe3U/DsclnvvyXhTKv9bsY0n2
LBRxdFS8RKw+Rhlv2LEh9ttK2Jj7gdY4KED/R5Vv6Tfiv+VujdRtZZVC+I3JposHFDrQNysqjFmE
TdTHXZMrFOm5HHW8m6ROO5urtzwpKFtu77llNjZUfwjX2NUjWMvaptlEpaPB9k0QsswV3T2bZat9
rGGUGdRGIWskiXhQdItUXr+uW/Ijs5jepO0mLtxi1pw8adKQvCu5nXT1+uTUAPVwRN7ngWldAg25
AwoE14bHVjYNaMh4VBW4om3jB2LxaMkyE2QwXec5mFWyfPdWQ0zifYcFQKMG1TaTY11TGm+dEfu9
soOgadNJr4qjfhdBsPsnPuCAqwsPHIyjdLywwsF+2bf6pY6AdIpUnnf0nhGbirWhqO5jRFx1Xdzc
w1a3wxuPQ4DiReYTX+sEVo7NM0vXjnYRTBukegIEcSht/a7U6g2s3LmzjDAlPfqbKhBjGbLqQ8mj
qgJTtVpDscqHJXaXODFeBrqi/CQMBSNi4I4fe+yLZOu0WXK6q35kdf3mJ6hLpZr3P2eTEZDxHEDw
XBL7T4XL1sOp/J9c5PMGUNS0ZTuWANgb+zbJpOdlu7TUl/9qxRYpppbHseJvSN4QXwZgYje8rqvo
oclfVf+35gvv78fbufog+xqwcWA66NjYLwtkbiRk2PSAvkltgnWYskdB/PytGuiS/aCN9WWlZ4tg
h1D3qf1TGOo8Rou5FKl6qXz0Kj9fxxj1p0K3h4aYP1rMwG551LIV/lHHizshzjNllCxPm6QA5io5
O13JgWwUDBCGbk+si608eTtA/yODYuUyE53/yHZBEDTvPfkojN/7tLYFdWB62A2D65TIaJOFCl0r
s1cmoS164AhUMNUz3d6n9AemM7cDA5rSLS8mKpKseP/8YQx1fc0BteBCxZyPP3HkH+flY8G+2aLS
3bS57lYjjXROV1/95KkLqBcDg1fFLwwz+O/6bmDl6ruYFF0wsxzeuKu4eghTZbrkc9tomMByl01Z
Zev8UBfgZU35AUrmPpL+ejWAQtxr9Qmn/KZ2C4azGWnZgR0nebqAZmjWii6najodJrKeOCFSEgdA
AgeFjcYF0/FB3DRtjDXvv+l2PvJnfMmg8F6AhfUfN20/OMoMsheHcW+oh4MC/9peIcYQ9o78GTcu
L9i9cM0aaMkBE2Oh98IzkqtC+YTZlkN2hCNtbMwhZjrs45AQXhH6VIEHaEa3OUH1WA+TkuCSio7E
ZijhoGrBbb4L0tt+mIKy2PO5WCOyQwnRsNjWk/QlLeb6FLS9j6aY+sWQxs672eXpvzDLm0SHbYUk
mXVkr95M7GjKA6kMjcUaEUznT2fLopzc6sVa2mKrFAC3A4msheDWP05MpPNO6gDJ/2lmAlakzWv7
9SJkYgYf/OftboIy1vnImz4wRfT5cs9VNbm18r4th3QwLxdnEPO6P1MP52xcs4AOGW1akk8rR+3z
ZA2Yt5S+Qws/8/NHNlD8nU+AS9J0oYOXgh0Cve9f3y0xVl/HM/kuEVHNBa9htNpAKpYdWYvABLRH
AIVPYHMjmm38HjO85eItP4E2lu7UUjPrg/f6bG+E9ZXVj1qFZqsKMBXZ2NT6iGQPfhBOrOzdKLaB
PUQ+9vy+Tu9sNE6NxEtcOVoCkDNG9w7nuh07idDnoe7XVeMGzbhdxHQ38OQwQDrUU0zw944yMfP5
8PPncBiNn37Ge4KCCSXF7/8+ZWhBTNShP/KN9TzTzZo40ka/yxngsZzNWRhfCGsLZ5lCz7eBjNTe
x2vjoM/mxfjPVUVZNjPz+kmJmxgCbTtFcBz0JzPU+QkUVnhnUmKE4TpxEidQDyWgS2JvEPOmBePm
D2gHO2T+aeeA4oWE/7G77n3yj6NtitE9dEp2UlvEz3Bx38xjxHn0l1YpB3qT5d1b4014BHZbqwQQ
L3N55RstIff7U84BiOldxZejsKUOY7Vi4yLt4CseI6BLVafNsri/5Xt8d85CEgTFee6T9L4cCNtB
CxkfhG6+8vtgiqNH1aF/nDHV2Qu1LHIpD3iKwQvuxEjJ/D0mHH2wmrhSdWPNeMR2U4XuPAx6ccRF
qJQP0Z49h95Q0twBr3I6+kf1D8LrLHxSbvzDmioNvujHw3Tx9+d3VcjCNAdZom+y6teFXOn9HiUg
55/uExZ0cMk9zsPKSYHhAJxEAI21d7Is6inRt+0iEKYpBfT22wv4Bn3WlIDWCgPwZGCHMXJ+ohiC
9alCM7su0TIecjAK2XJRrgFEzJJB+ctk8DdKmPH6nZuzSdgx9msSJg8ekYb0Uv4cMILfka+BnJY5
FPyDOG7DClhbBng0yiMv/3ckQMATjevYeCglfj5DmX8/j9cMXUWUcRxI9dxR5iqs3ZAcVOiaaDAw
HkwNleeIlzchJZmU4MFxKlXHVqY5NpBaNneCyiAlQGWYQlVFDX5teljcQOSguXU03IQvAGndgyl/
vuN7OdjTNDGUtzf564cfYNiyG+EYCyAWPaXUaCJg/1vEMbIz1ghB4HoH9os6pt3oAEX+6oYTVH6u
d2tvw1a8WS92AT38FukycbF/1awy049AG+jjBzqwAy3JKaZ54I4EzZ1WJLyKSwYBp5XgWCYpvcHt
htIBMaEZ/ELpoCcyF2iDVE+yZL35EOWTC+GkMO7JuTnX2t9Kd9Fmah1G1KbXJC+cCf2iPcgDdGJD
maSvtkmgbxIzP0ruQmeZHMCH8kQhBQDV7WEl6mzIHAUJ8BFI/ZJSCC+azwxVTT1jJRVbmeQcmSHn
A4HeBu41xCerV74m5lSi1ieImcpvPfZ0CZ/Z0a/bt2u9ycxXD1UvVJrap7k+4QJwLxnRnW/rh8IY
G1VycTDRy7BtSQoqOdhxj4kI22egN4XzSdK3u62wFNk/DiTB4A81+XCqFQ5I7J1+K63QJyw/hvYc
nIfC0vCx/3nYCIlGoPIUJcmweSb5bvPeEw4A6xS4Aiw9DAX3183/D3D3T1rjZBe9N6/CAeOnewjp
fqbJRE4zdxFY7VcsZnMvFTjVJ7iCQipiLn2bScAFSNvzPcVDU8dEkpb9thd69D7VSamSySE7W4WD
CTnR4YgLcK+mXoBjUkJ889gd1Hm34aKUSG3rEcTYqMhG7+puqhWYMdnc7uJp1AEv5J82ErLPHLyh
12ExvQ1cC/T9O0s2ywNfa+j5NQTSjPi0FyHCaRiXTnt4687xxvsaOlJlfQSlbgEauzSJoXl7G6s/
XBQXs1FZg5eHGWa15jdrObetdxHJHAbslJuf2PlKbDgZlDqfkDRtxoE4xiLE8H/cKt4untzzlcvu
FUPpfqhto/xH2JBxnD0udIewJPiRbe1hXUHz9qRs+bSU6n4kWn55uVxdl+OdMokHl/fLPGRAqAVd
Uay3YPg7AbwdYCXtyF7YHtVJ2ZRGDZa4LzO4WgwAZzULjW7z2IjdWqHn1Nfzd8P8OpQcJDL4Yxq1
5D5dyvl+uxvgrYwgfVNNkrXOua9o7NzRsRccECJl3n0wRiS4+vNDyG6GAaAj30XUSeeHQsWwoKzs
61AJDIer+HKBbLNSCzSoFTj9o0BahmaWujHuOlvyw6H9OV/r8GunJZ5A5MjElVg25veMI12gv152
kmvCNR9oHY8qsyeBt3LW8NDdh7Ifh6tR94rkAJZ1KWBKZUQxF3N4yMKivbufwIIiCr7Ipso/x3Kb
ezBZfOA6/55+gdqz6SyxPJxX5g5NaW60vmYjJlvzZh8LEHjY4wY3dq6H6c9E5YmBAiGM7eHPc/lr
vOLoHEzci3laQGA05BUFzAgLU2wmJZhdwQGnTfsWB/xyuJClaFb/Med65qcyW83pLuCBlf7Y6scY
xLEWgnFxCcy28NRne8TTz0NqgboILd85+HDiM7l6QldTrcY4rq5B35iYgPjMPDbKBmSKWVCkOHJ4
RxYvCx8UHifu4MMof2eg32LrhyvK9/i6es6Om6vjFLZ80DXZUHoh5IcRj3bHdsJ1kOOTB3Y9r1R0
5vMEmbfSHx6mCCTAXBFT4omNOf2P0zMpcGnG7HqmISJMxwY+Lj69V/wJivkdfLS3ATfa0LZBiShP
McjWunLPMtjVsq1Fe1ddApvD1XvO+5jU8Sswaba2w7vfddjT3V914gQzjKs0C7NMHto+00NgWmy6
Y7mKUYadkRUZ+oNI0JaEt2Q9+4xnb2S3gtbxlZMdzFhXSr7LyP76nlXoq4hZi4c1lOFP+IKS6Zu5
yw/Lerxu+w/CWu6DRf9Wb2e6tKARwnzJGneM4dZOX8n94TtI9wM/dlwcsP9LjWtOFTmQ5pmQJMgV
jRglS417HyRXX5+cTVPvnIDkBUi5Opfv3owwI9MKe6IA5t1uwZIeiMeWol41ct6RV5pCgZGIckXG
7e+KTLgYuspliPfVDlv+WysR84EcB/M43hBmZXspq+BXrmoR1LJipMd467j67DqulyZyo04hdR0I
SSerBKzZ4R5qlxFgzNY2q11BeiTu+WEm0M1u9QJ6CEYcNlBwPqWuieLXHWZWahTz2vGPKybu7GHE
2yjEbuYYhxx8j1x1MB/S6+oM+pW+IcZxGvzUTU7MctOqc6MUtEYKIZowdzjHw6kVC3fM/Zqe92i2
6YN6kvC933ytSFjqYiFsnGldoyjFq/Tv6iSmaiIFtbFfuNgWCuyGzbqiHHRpxitN0jDfAEaeCLg9
6la7m8GiiV3mDRIcd7LHg+22EAF+TzwVologP/lwVDBLMWKVGTW+rukecZfeDzFiMi76SyVx9zdQ
dMW5/7QcVedWhNbw8kHVKFPv5z4cfKXOeaqK8Sl03qfQBCGBa5kLEWljc9dchUO0R7qvirQpOQgt
Ohe3ZLkO3z3EFe6wCF+nprYTUXegyrU1dT4u2KuKaZOH23OodszC00sKZDJlD2MwF5dJkdkHj+Fo
vKj51memKJrr9N8fuHoXkcWAQ0PquD/IYlWP3OqERW0OxmQhK1tKtFSHm3YqWwXmsf0EXg8QBEar
jXk7YuixCqXazkeM3KMvZhGHp0RAmhOfU2lojqxjeichcS9xvZuNWO+ajjzXi1YZvO0CvSYrMZ59
bEqTyO+6kkMR2nmfsKp0HMtE/TLD817JvcY7pqPS3NJHUtFer7cSOiff3S0dad67wqDPkDtiz48I
lToea2+YMuU4qZk0kk+Yf+P3xp21KnqlIolAyCDh6rpgwLLoxxKsdA+WBuWjnGejp6zeDNn7+XW3
nnq+BbgnYRgxwbcea+TUwda7mhdBF6Bhovp7cQjzheK1MoEOId4GGnTjRz/maxLQrsBUn8wVcQrk
F91095A8Nzjr5v6SnDrK5xOYpaQI3htWkqR82yKs+yepQKBBrpbfkYFHbIi/lGG+y21ZUc1EKwJH
+jwBJ71KxYmEWjzMGkWTph+mawD3FfhIwhjmAh7GX39esDPMCG18Ry8CxJYmhh9Zbcb9ZPO1uxjO
8WbCKJ5uZRmy0qPGilsU4fTvaIIYDbAwfOx6XNWo96xSY/MQSeuFurDwmVLt04vPgiXnK/Ku81mf
2SDWBDkrQ9Vrd1nLVzj2p8Xtk3skxGy2rtv+reFYYobtwjdWWtTM4iBWrqv2yUSP6fmzYNfyJwud
m+IVwdP70L9hq3ZMlhKwUC0oWZ7tUOuqgkb3dAZcUiWi/U/ocuYuRLXfkmxH0kUfL9iRpSAQIdji
bigob1PP2BW7gA1nca5TUiUeNclPfdLcqgsd4f1Ana+g2AGQasPL2Hz90k8jQ7rb9rTtR/XFxnKo
TE37wUx07u5KEddauyEfgfTtaadKFY86QAv6bG4YZbgcBedrD+mLxtA1OKHWTuAfqtQjudgtB0R7
FdjwKnNtw7hqBKBQRsIsIbzkF7s15RjtpKcur4IvJg/PA8qP0QjffQtPeh0DrRsab7npf6bX/+f0
J24lBg28AWhPu11d0Qk9hLoFhpfSwKTTc2mrezeCKR9d3cfGN/8yALH5F4yRlHihMAP7hHSE2DFD
uYr0XXIqwHZGJH66m91GyzxObpiQEW4NA+wlnh/auqGrWsZVXG3RCawF9pTl7wHmkx4xls/21B5T
l3u01BRqFixHlXb7+uBdTofW+icOMpPT5lI+uy4hso7V3FISsv9X/s+JZDiBj7v7+7UdjZBXA0ah
DamRx90jpiY1Lfc+hbNtvmXxX5i9m31/gkZeJRX6Nl2SJIdJDWzqLvd5zkWbjqoCVfgj57A2Iqtq
R3U+4ucHdLUOAc01ZJSLDs7F0ZjCLasbVJjR5sn5gwCnRGQLfObdE88ibCT53ZPXYmAbY59f+EPt
RnZ4LDjkpfVsmufCmDp69yUcpkw5X7+I/xZvxuItUJIRx3oe87dZPl7l3gtWFObuoJC3hohNeb3/
nL7uPhj7Ew36d1Y9GVpz6ZRs5xXQbOVt7IG/E6ptevemCx4TsUpb+5YqHhCZVY4nE9PRPBXlDDfo
WG7gSBS0fLOv61PcpJksEyKLsI/6URCuKzLEwKTIurDnCKbXrAFbIk9dtLBX1nS42J1BeNK3KZ9E
jnjlc29WxAjsWiztBEeSV1ux1+e4JXsiyowRZS1kkJim13LfL1Qlm06wcLSg6i0STUtuXtpvq3eE
ieNVWNQVHQiEcBdDCTvySAINOl/c1zVwfmanVeR1MtFA7A7umYR8COKXhs2bfek//ABepOHrm2Rb
dOrqEKNazH9A3x+GKPGzHkWk1PVBIMh+D7B06XNm0/pLnpG2xRe83GHkydhjkUCg8gsgt0nStncH
WQ4C4DU3Ny/ZTqX8OVsxCNpCPU8Jyn2h7MDVhOANm5ofqUxRwdlqR2wtlKEIxPkNx5mDv0QfrNyi
5VNQ1WgVCOhA7U4FgVxeZHahRL6dCQ20CJyw+cv5/kQwtohqibkXF4VUdosPIUa08iKZ054e7pnn
Z5Fy4HfFT0yWZgVWZIg6b3K8Asl5hJkClDPpCs+kb87iLSNhMfUkSXU8y7nfue8GWcmAfpdyyjwA
myeCQ/m8/5XpKzRt6SZG7CfgqjP1eYwxXjpbJjFXqyl5SdFW8INa2MGuh9IRwtBDqgBjO+VhU4hY
LxMMVgP5S5+LAf21rx9ehQnDvIRbaenluHZnjm6FfIH35A1YZfvSTqUbiEeS4hiXQTeMhKumaLZs
oYYEearZLWyfgddq5OXDVMT5N9bxH7Smo2P7Ho9RT8ceMDEv10oC4i9b8Si+Hm90FRMwTPOmSgZI
vFTtT0GqAU2t9pE7kYfUEM+jXjmW3ErBYdIzALESZ8UwEWgpm+Nn921XHduC0opf7+7qamEYshW+
NWRIi9UD99Qx442VR9oL6kEEjo+zkwc6Urq+pq7i3VmGHC2eR6OZEYdR2HDibhIJQixkPxSemdM1
3hLXa7S2mktzM2REp4Hxo/RwLeVj6KW4FEFuBLYK7ZlHQqge/k4vRU6MCpkIZ1RRDZZKy/HtuwfD
Kg67xPBjfXXscHVDa7NoB1JF0lZPM4pNVI/sR65r67NdG3fLP8LnV2m5kRo1Q/ustlMB5G5Pqpxu
PVILOY4O1ep9hCtqLkmRQv2e5I9E6JfmW/HoyKtY08geA7pEiNETiGNf6T5jxgnk1AZ+PWnZqRsy
jZpLggKTAybM5+oAQlR1vjMd9LtCkL/xfRSbNMn13DbFb3QhlarFKk1MQnrFnCr1bsm6TDu24LO5
ceyX0Kp40hht09aUOc+QYH7rV/bqMCEnrJVq7R9N/KbSJHHV79C71EsaSqaewSV90O5At0Uzxpe0
Xva/46SRJpM0EJiZdAo/7uYP3XXPL+aEMtyzxqJdZ8G30kL3bgVhupwioIvwrfarsij8sL7tgg2Z
VwCnQ4IiqAPJNrcwANl4M5ra7ye+ZyiB51voZz1KdLKxYrP7NnW1oPdzpMJPebdFNqGLaCfTldn9
Iu9sgzy/jzawLtEKa/dr0A05X7jGVdqvAUwg5/miSpw8d/KRBCOhMnRzbxMRw33E0SPhFZu9sC5P
ozCT58+h1rjxJJ+7mpDFGgL4KT3h172xPaPypYDGcquss63m+7gF4qPKk+8J9qc2iUu0Dm9N23xt
nfAdxXOEKI1N4cWPqVR01NLJc/8dnpA7b8gep8NGEo5mMFyUrX+QReW7uct90tL956zxCb9bnCje
qvKkpg7TgojxER/Ftu9HH/oOsoCBhS+tnehjgsXUVLU9YGRrl87PFrMwbO1qEVIpwPzg836ZSJmc
/CNPMCADJoilXsh1oBD6LX74La9jozSKCqYHY1Qobo6oirPr9jaHjHD26Y/4hT0PcivQshDj6Xyy
lWHZB5x8HbkKS6AUR08j5BHJ1VId665GQBwlRX3QpJ2/Fm5Lig26hQQVl+eNTyHrl25aZ2ZFCLNy
aeOERUeBl1URaqzaCHzO4awPtg+z+a7ojQ3ZaAA7OUxq9hVE7GSQZXGmN0mi2bHoXx5UHdD5pqSp
cU1ZwavJ83rHRJUt7Wf+JTJbAJ3ybe1oZ1PLaNlU36r5y2KlRkNlPYECYeOvaukohqvOVQi4E07J
3eAmro/4GSRtH1mqg4vjvmR93upzMI/Pke8Zk1/9xIdmm9CBFln/mqFBVn+v2EbZzbMQusK5GRVu
ivwdoiLjeqxZNZFFbpow5k93xaL5IaM7JfcJxaByZ6QiCXlUjUFpKWcMk4zKJGlx7Q74ik4R1boy
DbwYAKnOGMoKE65+K85r0n5PPRihadXe09UWyHZ4TEIyNg5RG0P9PC76op+6Pgunj4uPcV82TemJ
0D6FcpzoI6pR1XsGDTQNrl8L9gJlOWvzzQSVPZyflIFfmhN9PhspUDxUPtfvjNpTYnalGs9vIvXy
UtqgPpj2F3lUEGwv7hG0F0elPOJqVUcTZy0UWvKtZ3+DLfHXJXHGao8ErUpVDIWsfMyiL0SLEdoC
lsEnuJZE1N75w3/dXh/Ym/2hrVS90PhFh9ME/UVd/mpAoVGAfDgEgSDZht63mWirt9B4p2O561tI
xLGfkJ2B4d7z7Tz13zXK5qKvcIwDLl+h7jURMbv56u4O2L5Gmw8qPf5rT/zCmIIy9yfE3IKlkEle
bMg9em+cKNxt5sgV9wpCq7r6Z9diswxwugZfhuc1ueZ4fX92aIRIMcGq3MEN7MatQqidH8yFShNj
HnmI7auft4SsmWxNGCC5D9QUWS2OOhoSClCiNn3AeJZDoPNwMRWEgFSQidbZ4rt+JES1qEAHvDJu
IwrGRtOqZK20A723TD2TMqS4O7Y8+TCpHJWS6bPIaGbyOf+Ou7JHeIfJatH8d5pdrl17RUW8lY3o
xp9vsSIf8yWgtdGS26Wx0X9/CV2suwFGmEDwj8aDa1EEu35ptDj4ZdcJP1BEGu8C5ijBcs4ZISeP
QhGuLn42ktp4POE/MqFc4IdHpfKU2uJlzRuyaISquNbmhNJi3QNeUd8ajNi0kWtZ1ciG/wb8Q6nj
H2J2UTCx3pjLGcrXY4HaGm31gdCEEqZtb/eyeEBwKv/MUxVbDuBzwqLtLfYBaUdi5KG709coK5GW
ZTdb1PcCQL6tz/hE7UVeBuXowKikFj5LbTcNfi84giKcb1rZUC8LP/YXhPY4Wl49AjAO6yDmJao6
M9+lT3Zzul13Nqc7w5wg2376BEIYNY9IO5d5/79N5x9R4MMprG+TV0I2zxqPMG2ADoXhGb3fw/cO
FhkX0w0K0edsQmlUkVuQd3QozPqP/lKngOC4qRAIWPoB4ALXKduJHqqLarPN6DkcCY8IDHjuQ8nB
CsZkqZGNk/vHf6faJWnuEvrROMdNOwmKlq0l/BUwJ84owWD3NeaG6ekimoq4li5X+RTKGXqeONVe
0M9iFFJtcYBgHAovK8U7g5GY+WjSXH5mKaV2ibkOH5ZWS2/v36f+KFzakjuLONgYb80RJlKr5ZpJ
ia/HnEetQNtqsI5uDzOzTBbgDNN91qr83g7BQkAiD5uo/fcanhV9YC4oe+cPMTgdz6hg9eY9S2Dh
Dp36qyxWiMycQ7pQ6Ukpqbt6jfpH6Mn4QwUos4J5i+r2eXDrHXdWW56iNdbr1ji5+yfnTD31t8uq
ahD9ABElZoiU8qkrxyMCrFQNxVjZlwonQV6Dw4iH0LbltqYEWbVhRa7eSBeZ+2JiehO6tvQPhJ6d
EzTDsZf99pOVq9Gj61wPPg/bbK9dDCzicCV1YPEvwejbwX0eo1xoRZk2/0OvltXAEkyH1mq0F6G1
LaJIqMxXl1MHnzXxjLQ7GJdDH2xpmL5VLP1NaI6JmwoWFMZzHGMUjj6CkII8ecC7mOziy67FHkcF
E3GA2klCv19+rc9JxFSHqBIQ5L/S0n4j9rraTFxSZei5+swEHQrLDHlPDf0sPwiQNeNCgMd0tFM3
inYpVljrEFAsX6WBHjsSnXm5QIgQyv/YYH+NaGyGT9+4/bl0j7gxi2nuYIrBRuNcXTFXodTwpGSU
msZToGOb6yFI7oGCpeHjZm8rMwu/gdQEeKdkNkQWUrF+D04guamWD6gWXXhlhF1dmJMX5ph0HNB7
W8LBtVJt6MQeSZKGzhzrcbskPydR8xE+BtvbfcONAcSz+awqXdTUzzgTYCfkzDr1dOvIiNWG5pOl
kLwVMfYcwk/CHnRbuFBwB265YCzzBNSqIrTi2F3XRoZAzInj8fSvtaSACwjyNhxkTP5+8AZp+qJm
mJ7Pps6KIjTxCBZKyBEI0FGlsPFKeoNRlCfqVw5CZmVZmsi4xIfb2mwhBrW45hiLUI83HpCdaOJJ
2cMwkqCLox5Fx2L/CgR/0uYq8LJ1wwAliQ7X8dguSLp55hhBoH5UqxamiMfAFKv8cKPsZfI392zD
HB7LABj79EnUAgQZ7EDlBO0MmugKLiRbAmSlLG7vVkC7Vtx6e/rFErWyEELsIm31LU+nu3pvlufu
FOHZld2++fpEwLJzNi2535VP8MbI73pqFDvUTOKHfvDgzdPHB6eXCWzWvQMroF8LznN1bpmjDRGy
dlWwaSUBUeN6bc9PNUVjenBat9jILatm9uf8IIwbE/SKEbW1w4gVk/iOXCjNpSRKrHvBLFDCX30d
5XJdjoLNKDiBA9IKyxHPN51pvrxXjp8UGeBE1QzSVgjgeLgrjIPsiP0sPk41fVF6sQBmrf5Pts9V
4rExKR3Rnj0QZAorkVaaNYMrA55QwRVRvTRdTtZfGFTu7K2um6ymxqLzxgf+Ws8LifK0PWgwldEM
NPzexaKNPg51QnXo5H8YYAEeJkgfRS2tDb0ZgL/z1ATDp5HMOKwtCKNYsUyV+zcrfs+AQMaM3qx3
PAgugJp/DCcyQMV9KDw0EH8IHI7upRnKKBPwLsfai09shTJ7w69vdQwVO4JpZ4Bibw1guNxKj0Wx
1gLZYoGC25wKmYLv61S4QjUPA2VN117uDw8sn4ppPkt1m5u0v4A5FrJXvnjhBtU305Q582KT87ax
+yEp38evLHTWz9BtNGhNoJuxmXbQztxRskWa6a2sM5Qxrqn/xxhVKqLW7uMqaXgwNYy+SaDDd4sU
+WiWCKx2PcTU80q6dbQn9TBaqDz2UcnW4R706T3vmS84M4aAlYNvqIzq1ZypsrdC9m8SjZiKLB83
0P2+ai1s85TkETOm2Oxm/w1ufD8hpZw1FIVghiTNK+ScKRjNCCXsIK/PeOtotdmg75yllS8o4oHe
VQrElNWh84k1BrN2tOvTlpFaVCIngnHbCF5Y7f4FAAO7atAbMoO9JfS2xl5ylZM4PHZbaDqFxvdN
cWTjT8lnfEP8X8gwk0C0lSNjSpfsNITUv9TFwIYfEzb4yjBx45rKYX82IUhAH0JiizPdkKF+qJaU
OKfmveKK9jOTZf/G6pAxjoKGKWtQvo0cJSQ8Dsmg+KEJF8eI8uX4Syl8z2+SfC04eujP1P5Mbq6o
XRC5DOrs1TqDPM3c22g/ot8DjItFtibheN6Dc5fYcNFoz0YHhEMlEtWePaUrmsVcZu3MKA6W4FZd
X0+8Bvd8HgiRqi9KnpFgJS8rTPB9H+LkXv6Kn42LvPIhVb90R4AWA3bKcyV2AEasZZEX0R52VaZB
Wjao6b5kJoHJ5Kam/CcEwiPUq4xgkWrjibedWhceAkdkLyAok1rjqNx9ZhQBLWQ6PBmiSytPBWLo
lm3BOX3I5DbmU+S6phNq0Ww4L3inVEpTZg3vu1uuIeIl5ux3aaDqXM/cS31qZW3KY34S9L02qeZ9
hAntiuQmvNGSCqWfRuxTKtbf1/78FmS00ln8vWs7X+QtJo7rpbmjG/3vbUPqcLF+b4cvxUlaXUPE
RuFV600gxvxsm0ByAPrr0ohAFOeOQQdyF4YoM553WTJnLhDji+H2/+LhSaGA9HeE6ZnC/u/ptV7/
PVeY5ny5tbM9NgYSGP7iv6ZGzEhzvveaFfKPY9yV7W9mhmfdndyLRDEi3ojGyQxT2bTYPE7n+N9d
UPNJgaGb53vfySGp9YN5oJYeBoenHn3UwaXnJhd41uByg33xqsC23FlESdzzNKVDbHm3rCQuKO/W
Q/IKx3URri/AsTwo+Vm2MN628H9hr08mqWPjIS/gRD3+HukRSJWAwAnitmkkQkgTtgTiqvXH0xes
aWKS3V68MmhRAqc7IJ+DxK/XPoAV7GFxs2rkDa/M4FagP+kz45uVpic3u5vjqw3lCJ2ON0mT1qLN
YYDLAsjFbXexk28X4LULamW2QZgNHBkLpzwGROylGW9G41bxehTi5zfwCQBzGfUolyra9Lc9nM6e
dWk3F9EjL6pjU7tt/ZBh91zK/xLUE1Kprq9D22j5u2zKTcj2HhjwcY6tzPtqN/9jomGjfmegNbKj
c0oCtbZwleBdd1h4QycP7OT0hpNtXkSrHXQlxebjTMpmat7khlLzCr/KY6yZqEVJ2WO4FZjCx2Tb
36EsEuC8G7Jb3Tduj9CY8zkh4Hwg4YBJOnkMtgLLh8aOtnqUBCq7gRkrdKnZrkP2mjikGoVlH1cN
MZwYarUFEN3lbaozgFc6O8PAShrt2k/UULn2gN6isLIWQcOW3ZrbsnOy+k6fvXftZnZf3rrKq+WB
5J0rZchvOxRdYXIfyUJoRVqEjcBGhJdh7m2ZpgEI/oSB29Q/TYS23xwaY5sVfo+wI4YqCUiooRHe
qikmkVPyIy5t9mFMcTkRCh14T91ntGj3aLidbVDFxW72kHg16N8FwsQJQ/YmQHhKYYzt4ovQak1/
fnHObqdYwok7QN6TZZKm+loSzIWFRa/QP+Qtfk7eEqBaM0e5EeGpzmyTQ9KFAJYTsIuoIp7lNmFR
OpYtukLdbzXvkerv7KQIp9Ew4hxDKA/bgqINy2JV+kaC6uFvvDFQ1zF6uLtj6MXAI3tzyal/cyC6
XmzAygNg1oEvPXLNrTCjyTsEDC5w+bzmmBL21ApBBP7m8bm0TSzwX9AnM2d2bVzw91XNUZvLXGOH
35rgUTiuSz3MtJB1MBPpIk+p9ORF1IGkYLt4bZo8EOcEQKGXXxT9+PvivZ8EjoRBUfsIKGzS9zRP
7OM8v3jigGMKBhWSLfJrLZJHTXRv5Un5lpBv3avez6fa0exGmtWri+9AAofg9Dx5CGXnsvLEDDLT
t5BNjOexSDO6DGztO+QHFlnwsdcUdqlGhwHCb5SWsr1aznce9CvfnaJLXkpiPlRs1oE/9X5AiU3N
RghLmSaau6Uadw5TNzSz9CJBgnxAjh7tpEzyMyZjKxlt7TRX2byRnbDE28HGkSkldlxi3PuwGAOJ
T5xCXI1ABIlmE5gsbIdtEx7qELc3nNpHy+uuXcGBsMDNnt8IoH4Tyf1V6TogfUfACUYWnmaD00ig
z7enRW/MbxsDDQNGvzyrG8O4zIx2SR2IYRVkEZfHl/ZSKloisZpm/q3SayUUyFNohZwiTuRzb9ov
k+zRIqCXnlF8Wx1Kcuk5oN3p+7BwygMwQTx+3LhCvNzm+krRpzkCKwDO748TYTnboBWmAtGuh3bm
/m5bR3/drm2CVq6YQCHVE1QnNT59njw8bujHJF8uQNUnxyj0P7zXFkEvHZ0ZZi5xUnlSrYz4hQii
MKgmYAnp568QxfZ2wm8O86kTNTJEN4mLdXKTL/9WqQwPC/UgAA5a5l7gfqaYSKH/uJBW4+4TeL7j
6tJvFIN13YulMMW8gZ70012hK3RzKGlaisL7M1NoyhdJKQhNJHhIAvBHF08I7U7t6OifZIwh5saG
L51bByv/6Kir8Fle9/RT1A+ODxF8BGE0GLfMUOfOWYyVmAZzTr2UypqL8oJHOPaaLbwgI8kEYZ6S
fjXGlGoMOpXXM+fzpPSY4iJUmXM/YSjI+/bPuS6lb9AiP2VGkNc84Dwe/0RX2IhKZBWNry+G6/sb
K1oirhVVOKoeDBmNu2NGjKPGwfumY1myK9miDv6VFHZzrqjPb3SdIucgKRtdt3zJBLujUQzsZo55
iEITTcKbfmaYnogz3OXJQmZj4n4/RV3EnVHgO0ttu93vy4sQl7e8sBVVqbcpV7zh/J6CN7YNUn0k
N2wGfABB3325gRb9N5hwVhrXlGtetQhhjOjtyyB0UhabuJG+Nqv1jo+vOIw/xxYtvTt4Ij1RZL5x
tX77g1P25yTlI7LPu2yA+2gQX1jgGQsIvS4GWrc4/Sk4EYKM3fpDBh19dfIiNZPw8r2v51AHFbPY
WZ3DCrdbCi7uZTz1C1jaEJt6BI2Fj6giErvClO4ru7PhLARKOqGLZE4rujTP9KNXIiKYRIJvyn06
yXUOwMuNYT3ZoIqcgfdp14X492nAbAiDjAlnKNkwUjR5uVtEwnUQ/LRRap6LGwsqHHO1LM2mul4o
7JeZTouWENHOIhll1X74VCotEj8TJZuSSv/WtbAihOEE/WMQyO4XbbeI57xppxaVUIsGoHLdy9YD
57sRnj2gC9G9+ebNIQ71NP7OMq0c2qXCgUsYlRC4qkm3Shgnprmeueu6X04C8lNpqTJPKOQEPTDA
ZnBMV7z7YtCjAIeKV6TitCUDo+rivPgZAiomV6BHXjx+tRBpqc+2dtO3gC/GDN+IBKSHNhT3Niqv
CmaMOc3VdftaSF3NoM7HZr5zaoaIHew2P0H/OQt+QYKWSM4EwLydq0f9ZHgeQEN9FdwRKzIIsw+K
s395vjn9S7rMRnp/WlbKWfazT8aRgIBJjsaO2caxwrPB/q/3DMKMGoroozYMTc9f0CktEjhr6usN
Y5NTe83ryDH8bwvRl7XbnYmx1MzEVxpiNfVsk4uF7BptHc/eBKBwRC4+1/oMV3jdzcthcrHYxbdu
O+SgBanuN5VXGRZ5XOeF991bkqF8HYGFIFGThJgApFFYbGwxtkOxjbLVLFnOxb2gGD+uQajMP4hi
9vFD/f7ZFBNPE/sTMlTMuTiSUO0CkZ+GqwhmP1cRfDbRFn2M1E417gUTCMC4KN4zu0gIgvbHNleg
E9Hy9Nrg/HUDk3+oeQhBnRhc8umRQILG2bzV3Aqo+ZiLl5JlQ2p2qPuqVSgloKqH0yfFdej2jvxA
U9ZUnCBcHwxDLaesKAv4sCcff00Ut+K3Fl/3uHeU+U/dgp356eBAzM058vhlCb6WUBXWlhxnPgNr
hkL4tDozKrhncBPxyNBAHVWgspvrLu6O1KsnvrU8XyOlBshNkZ4RElPBly0fqzRtpGIOfA0p7saY
5/hYwWQFDu/GeOWMjDhAxBrwYkK9E+mfmqQgOYkOGCMPbIrVbjZJF5zHNcpJsbjrGYoyriDKhw/p
mvzp3jKxIUohr4tD2QXO9VPZ2jXVVP/w1caLGWo2UrFydPx7OZuE4Q/YnanHAuXE7/ZqNuR35gfU
nUERZRPLgUO8z7rDmQPIDdgp/4wNEqia/aiMZRh4x4snlLWJiNgy+j2XOPWRHXK8HUJ4od+mIcf0
QD+irwQk/ZrSzMFGsXAacp470xqYyARxuY2H6rwdDFO/zcK4wn/2HqKnhtgRbzIEhjg7EhI/rkK0
cvw3gkmmEdRyz8Ee1XAhKYwrykwYY+MI6t6++N6v0vrRVyqxsJnRVkZrMHM/+ycX3utOFsfjDSy7
Z3QGfSgSLmXo2uhlDS3uq4IlGiaxOFPbR9eF3zqMeaWSiOwY9Kr7aIf9xduLHDvrntoKfi+QTcUm
EvXNZRxfMzDur+08Bza33GRkmQd9LN7+o5l+mZ+HtIgnKKWn6SENVAFFgNcGRznufPEgvqyS8oMZ
+N2CMQyPPQ7cGhVdHGgGotS7ul3TuKlgiXlTRYld+f9uCWo2EkgvHv3tnSQA5hG7IRVyXut1VyKw
KepBRZQxeuD+QSaVf1UXjVI8lWvS1NvRzd+wATSeiMPivbdRpjsHNY61Gqkw6oiPSVTGFDzzHRJy
3zW2WM5dLfdDote39hXcR8MvRWpsHeaWLtC58I/50whQAv7x+VOjI1uFEQxWGX7akDtOJVqcyqdj
aa3bSXjNkbNaxALliIIkZmfzl0Y1D4ZM4UirvfH/k7ovgaa7z93FnSmNrm7tepkXHR3RzDHjf6Pm
k/bDrkx9OAJnMsUADcsuR6xLlEZn6F8wQt7cROkfXa7pOsyC+8l0q0gh7Cub2yR3ofTlMa7oM494
XzXFndcF+Vk6/r26gTMb8M1MCOyCqwEk9OFbVoWs+uck2LLyWq3otxYc4g8EPz2KSUWt4/kxBWfB
hHIRPbqJ/bfBkGB25e7+cmJjMt9RnHIvsGqK5cnwpNA9GAZ+63LWr7vDZdYXfup2koOuxAtQH1MG
MQ+74t8gFL2SWNPwgXrX6n7Nk9OOom9o2Oq9aHUDQIJwzSjmLS2X6zouotV2Ju+mIAj6fxLQj3eY
BdBLnWLA0aOmgznIYZM0HnGMKtsdJl81nDZDvrqWo84/6D/Wudn16Vzh2N693hZt/xjCziHib8N7
mjuEs2jn2sScg+0lfh/rh/iKp5ChhAqBEaUeyLc42CNJUdE+d78LxwOhHdfJn10xAtr1199ydwGE
YJyKR1ONjIbxefd/azEgDWpKH8NwGZxSEbPSItmXitu3uCssPMNpsQDOjTndhY9R6e37chDLmS/9
y/faRCTBabZNrmtzY95blDcS1VspeKnG3iFDYNfOqM4jUjkPTxZnkQH33nJxZnnjqyYVQJVnL5Pr
oYng4BTQ0PmCZ9b2VzUvzSg0mGim0VvTHwFU/Rp9FYOhnnlLH2wp+q8iKcnHfjZG5hcQfx31jbM/
Exa6Lb6s6hySJ3t/jyYa+CwRLffiHMRZhcTC4tIsWVpXMK0bne3UP0g38UywdXsCkFTevj5L9EQY
ASNTYJmo+Cb9KsbJ26xtW3SVGngmhhHdINGxdMfAr4duGjTZFH3YDaE5uWlHiSET7sKU2gS8vAq4
crrK/w0WXpHsylmC+YR61f/1C/MkAjuDNZZesqqb9mrozXiJSkUPQ72wH9R0+s0F8DTdtnopNz7e
qVd3yT00QDpCTzKIhRXHlviiJlteQ9k+cT3VMWEMbc9cX7tyP0oLOWrltpBS3dNYGsRW09JvnyTx
WXBxK1Yls7eCHxNLzSCYQLjCp62dac3OJHc2KpG/FevypgLP6m3v+y2Vxu4ZCgiRqa9jaEyyD3Ff
t6WP5Ol1sdLe3DT2K1yihadtj5DDIca8qLtTR6nM6IPCrIBmPStVDK3+jFI78SrIKYYM5BZH1sSO
hIgK5Imse0szRzHXOV6yZnSa2WD/kog42QIjQ9V8OkC36MmKtSpjUNtzOxdCEqFIqkHUf4Mr0FMP
YbbM8yN+5xCU7DKtDmXwEqjxMFHHENXkDA2Myj8zTu9O6Ez9KVNw30eLPIULnHXtky8VFYHIXUSe
auACYLM2LWtdKWy/VOlBBNKM6hRRM7peuY7zjzxsOJtHXBIEkoqHX/Bgx+wx5pKB27yBOUmv2d5K
iKSdWcA66VnkrzVKhgl8DOqHJNVtFYILy9/oHZ55sQSvtjUfa5f8eSIBlFTcwXAdT5BbiNdD0myy
hV/7G0nGuOTV2mMS3GDJ3bBNZ/yIOl9NxZ5ePytYMTP6CE7AkSXVkrDoIezCvFSb1pXIjm3+M/DM
MGClVS/aYI/1c7bvEVuBXvdhruFqLAZ60yokedrqD/5LzIU7nf4wpb1gig8BAD0YD39u8Ccd7+Nj
56/dNDKHSAGSGyPAwZxYmymsIpIJnum7+hfosJqUZMGhtyFKto9MKuAiRa8uMQPfhH7aleYjvQsZ
c/GEMNcyoGHiaETbt28Uh6+gVxnW6QsTnDGscGqS3p3/U+wqIKLt7H4RjEVXzyI6BPEV50naH9sq
ZvufudbkOUzOLNwhsjX2r3DVVmiwQw6SM9CqD6b/5wLkvZnS49zlK44QwGyKrR6wHYkyhZk1kDaz
70a6PtMgi0SWkTc9Xn++UOaiAqBCdRHjWIfNZ7U96+6ze6A1A48kJPWdJGqAk+2VfoyuA9KRqsZJ
eGIQ9g1frz33KN+JEzP97rxylRTMT/q84Z46dJRkTrfgj9J0FjhH+jkCijD+OSZytyIgtOwOfsYd
G7WptNooFHwrCY2OF6WPF9MInKLDXBGdZlrfmgLcGO9yfsyhMWKk2gJomMCV+QiLAX5wM7Yw1jX0
z7/VkKcQMcU3JJ2qnBA4rmxpCC73902H867nadLUqlgoAJML19lHvHJsCTTdvWtNoqyr8D5vAOAI
v0c7OhE28cmo46M/MA6mdTIBzfndrVXnlftE8EANekWkaARUF45d4W52Yf81OGZd6Loy2befUfHy
a2mC0zo4Up8d8bEWyrL626t0D3tMqha2tQTnnm9xouMl2/ldjkQYPiD5K0UwNTm9U/mRdp2tsZt4
YEdgEvfzsURxM0TdCVEnm7tL8f2Pug2JnoUzek+nfFCZmMaCVc2F4uR7QBc5Ohj0iQoTPI3UFgiW
IbFkpdPdPnmw+0GYGu628EmnXfaHuf8a5y0dLXOtj4m8Q1ChqCI0fOGYYTZG5/HbKl54qwmx6bhW
eUxSGkSx870/9J600SADAHQ8z7xfWvoSUBiAd4t1slzTqlFMB/PuA2UW2TPNbVXd4SzD/+1YVyFk
Yusk7r6S2V6I7PPZCx8jMRXXOuWgYOGXWTEjBWMHVSSoXGyOsF75atUjAky9khebU8pnmehDYgni
2K15q+yzFCBPJqXbrGsjnCgMCbDPzr6f91cNdsb5W5emvn0temtuYg1ew7TIbcuhjm67J3KuxoOa
tcvtMPw54CH2tdddh5a/POVGAJ+TmdTC+iDmD1sO/OmGnCDawjl69hccLismaUhpeQH8qbOO/r8w
pEJnaOZK9pc+q32z0pCbLK+/C+cpcPvP8CqfYMvuWKeFJUoJ9Tn7Qm0s5WNjc7yWdoM1Jk6SBo53
PVjugCoWWhFkeBEB3J4pQKEN0NS9bl+3W+1a4jGXPfMSvXa4QgVV/H58ORGl8nk+FY9ML7bUdy2P
J4vIaTLK3LF7SKpiYAq50ubld82GVJKbyWhGNbzxPVn9zZIDNZ3x7P72GAjmhqkVBqiNtNVdUXiZ
oO2Fu3kHyevedoK6kG/W5LaB4tKJCR6UnG4fOHiDdb3sWY6VMUUurKD6QFpk5nKu4Y8GHWKWom2d
WT0zYtzGIj1/gZfAsFq9hhaSGL74OqpGZZRyIPcQNw78sMWEPLKxoHwCNUQJv8lOTjmN8i+21ytD
Yoq9Xyg0dVd8+Wq55Xgy6GuALb8s4CGa/BmlDN2afW9EnWOUfI5P8HQpJAbQFgVVBDSkMEPk9k9L
6UAem/OerKXXI1Z9GBM3yB+ppbB43JGHiistL9pT6fhLnGyR9MLkLOGGi/RbQw4gxAzSJgwJwUxH
+JLMDCG5maZE58BASX1vpN9lOp68DgJeu1NHuelaHNr6o8nhJVf467UdN06hM1BODnOq8SSQfrd7
u8Vr1ChVUJkHNPGqAYzbnj04VMN7HCn/G2HnLd7zDGpjprdRBfHoqhRFSd91C+yXGnH3g5N7z/uF
zAKeUA/5AZxktdyNi0C/Qzeve9uNj3WaGo8nofUatOv+vzn2h/ndWc93EWGstOM2JOdNCA0Jgw4O
7FD0R8iuKdr/BGQeAhm4jK00AHK75BC3SvO5MQ7cxFjhruEgkdUpP8ggTmGPkaSc7QC6TcRaVtVa
m3cTJ6A3iEyZZWsN22OuZ0/W62lspmq97z3CbeTtJ65qdj2DxHrYKz6B5JBzyfhTbnU6YJKr+nGm
WkL0jSGcwTSaJu8W7HjLI+2KLoHl2BmlDNQGnNyrP0X1/dr3/8GJ22F4GKiYQBEEJdCqeYmy0MlY
bvVhKAaDD/teXJzacY1C+sRVu6HQtp/1nZdnkpgYP22ouj6gRI88V9AwdfW0P4x9JDXeXZlKhufd
pjEOQF2AJyrCSaHwsQCxp68bHlvbijoBebSa+1HUln1v8w+8eE9vRTsBaH0ebsbe2x1pTkKojyKP
Y3ERdCnTvCsiQ3pzlQbnJzQ/3O9QA6wn5iT16RHKp71f93Sygzn+Jk+I5s6kf45WgE55KDnYWZVD
7n6ZBpkC+FO27UjcfvG783zc+4jzwF47NfW1pXlh0uHpSGQ/5tDddZrDuNijHvfTxKDi/+3Evv8E
zObV1YYM44eCiJFTOwOTxXvXkbiKNXk3VrzLBOYg0kMT03beqBw/HktfVu0tR/Jv7WqSEuJifp8Z
anejgXTke3LVz7MPPBARyvRp0s2kEWXWTII/ZYRHja/keLpCVP28SO4bh0ZW7N+WFS6o9xjVZiKB
0zUIuZmvkO1yHF0uWnUHKHyMQKmh1G90zVnlVTjxAfPU2/wHRzGplwdXwOsZHzrxtsUeaMgcWu7X
29cmjbR3J7ZAx2Yq9Jb1EDmPxdjuJoiPxJSucPMyuhm0bB9YmbcP1i2xAx9iHvYjuqG37gIGC7Vy
Y9vKMcB5AR2fT9nATCvNyeC5LCd8UERoVUDUAnj3uH8Qb8yZDQ7R5w3IQDoXkvGvXTvCD6q4ASrA
BkaVlj/6Yhx+92cxj1xwNksSkYX6TzgGmWI++OHT6ASDWNg422sIfG+kTtmvjurfBywUFfh6FOf8
bbkNGLPULKsnBP2gueXBQ0/XW40lwnDkCQYy4RpH/O9tRdCGe+WAJpDxD6w2qglYZLLXGvw1jZ7t
rellsezgxNJ6Y3msCn3oOtClHhjlERdpa152TDPEFSrEFFxwHtA0jRoXrjKOr8vrlhIs9+fwL07Y
m4H4h14JF2SU19hk/8vLXYEZjdj5MxtzyD5a3Rb9A564rvQludDUpu2Y0vllo9VZBGSGPpvLtqRg
Iu3WDyfuybnmAlo+l1ekrJemC1+SygZpWwpGKd7gguEkzoZrCoQIxLSWyJgsbbL0Vac3xXxTNkGD
SpHhpFoMx7N8IkjJqo/B7uXEKE+D+UkJ7Dbw6JWY4wosfZdc2dO0wRFDisEXBaFhIXQuqCXbe3o0
UmNgpZo/IUgTDM22D4T8AU13i+py32G20ymxt1496ogE3+/ruQCNgJowoLT/6w6jeuda3SdStFyi
7EzhfR4AT9xusJ7/+ws88KnALIp1syLcGQakn9rvruHWEu8TpLsFEmU6+p2uGzw7OEm0LAzGoBhN
pHMYR4Undv1zgfgSoleZYyFNWU2iIqvMU95/JbR+P01Zvegex/a8SpUJSNulAmUSMSb2e4/TcGO5
3PFnb9C6m72n0EU8y1OKqbypO/XRyycF2qshAwFptl4Li/PmNNHgNy2u8hRta3G83HZ1nK76INa1
sRkmwvVm+n8m69xG3wEF63tcOVDo8M3ldKKDdmOB8Z5qLkjQ864PmcgAh/DMZ7oaCDrhOCdWYVi5
XKP/IPDB3RhPil2HPQ/hqZ8J6MZMsqrMlGdhDdEdtfaTvSG1m+wtRpBP9+5zFCyDhqXFLoExoewc
ldV9qDPkzGFHO/DIqSg8sTrYD1VF4E4wcdvutjp1zMr6275BrrCIYYVZ/PmUlGUJPy2SlDr6wO2g
4JJa8JFkdGmQRvUWmgCGaC1dmwg1oWwNPUkSm4tUApAanAZCRhRg1C7E3mape1DHqf+6gnRLd9Wu
jghkbf8ItotnCUiB3ApavYgsYOnHRobM7WIDmNASZp/XlkRm4XdMZfzYoB3tOkp1NsLHRkDNfo5e
4T2rRl0hNYtz0BBhh4BxFPYd1+MSY4B/PeQj39sG4f7a3olZLWP/bWejNPRp3TriHf06+QUPbeIY
kQW5xavWlau0mtgTBC/aKXMN/IJIARlPtRrZuOYEJZ6QLvLF8VxiYBs1GhVBujxfzqT2aoI6LK1r
9r3JyKd7BVdpdQwbUuXVHD9y3Zh6wIalq9mOm5q5XS6ptOG4qUeVxUELh/G2ChmZjhZtOls61Dnh
2fiGpx+uIk02RKGSdAO3wnM+VdXPzyM2rW14p1zC/24+8vc0AfgJTGsgNOHj5BVu0QDbf+AO/wjv
e9Pm0fEIx3SPjU4yOIklj13d1X/Jhr9Inf9mxqsokrOJpME+WW2Zz3cB0W6DGtLWP+s+1KSZMtQy
mT5pAbGMJkTNIEGd1sSgyzAzagu3jSefZ8CQFxa1stIvhZMXHTVI5F8gKchu9aDcbi7IRS63DSAr
rb7xVjQrYBZp80DigkjY4WY9/hKyI7nVtc0H7BOjYLzqEOALncmZimy8vcsB0plIaaZ8X33Jt5zm
iR6U9kIIkSAGv4tNro1WoCEQFRmDjudrFyWwees+dg+bEwomC10s/8CQI9+3FqtnN/HcQhAeCLGP
Ca2N8YaQy80ExEfTaXuaP/wGtdGTHYu9SteCCuwojFPjiUdNuwu0CTyRLF61JxQQWOYfh7xY/uBi
iVoE6uMbXTIQ7pbZMnSM/3kGGD8dvAOQSccj/oOLfcCdWLYRfAcc9ZTUZQ9R7tudSsTGPjuw5IRf
y6sTIjKzTRJa3Xn8qZr8C3iwg7zCIDc+T5Tc6+dq8JejsJXQ0iVw8dJhBrex+n7VeDnxs/Hw86b1
dB5W3QOQuufBHIjQ7LJ9NUemcaX833C4pdPx8H9sLbgAvxWPocrPiVmTuMUQjf6Sncf2VDwSr6wO
JJcV2hLeIHEciWnqoal3O/tVucTQ4DADu/HWKVRW+2B20iTj2pUe1GM+FxcP8tIX4N9MB76jzIfS
cFqZdnZSLMYYJxc4xKCGGQOL7myXh3VDwKbaOcoPsJcTsxeeZXQ1P5TiTE1mUtxDmiPH/+hhS0gN
8a166Is5eQfpUCo0Fz1QeDm2EO1kae/f0ILp84fBWe1Dou8SL4w+rdVX2O5PAlRyjHkyxTuGrtPg
CcGHgGBcu4fS2t/N1ixpx5xKzf0ejSqIKdz4mr1u+2OqUgGY8GdMrW+3Ak91ZO6UqNsZgsYif/k8
Y6E9CFrAVT6sOuLmqrNgbWyNQhdAovurtJuW5Lpl1szkeCE6tx552G48zTPdq+CLpTtPF9m1DvSC
Zw6pIt+F4Y+twj1kxqzlyTX4rsU42LK8LX7AkJ01VyIruHBul8Hh2rKhdeFSdflRbpeaXeRfB3Vo
ycEQQg1F+SiRD+GJN/vMIH+rJvpV4G1crVkzr9Lo7FEsDkCDgeaMt8nT6MC2J9d/2niYY3hYY4wV
QqKKN7mmvNTKC1t1iAZ27aXaABZ++ZAO4F6+bTqHxMbiWCMTYRlqufKHCzrNGuPbFrJ3XRhrbTDg
b6x02Fqn2Vp3TDTi+Euhn8dExVs1yBoOA1GXsZi+gUoIdVX1ok6qYAvFIuFQrOG/Lufnfhh/7TLn
T7F2wbA6OGY9mlbQUDf/VsadbOYNyge0q8SDykJhc+VSIpvsgpTG3TvxnEU5lRAIDGsrGuYeHenq
VC3SyJgNFtgAepZghoC3e1Xwbh8hdpByVfUlWAQJEjRaUv5RfoaAqI7tv37Rdx4SosKZzlu8UC6K
qT17laUOXnrxoFTs24ZLmTxtlGSpAXfLhHhHoN+YtTZylQbBUU9NdtJQRIaqYlzTNRRdr+Qlg94v
ITnU7WGUvvqWqeHAdNWvBwVVFgzdctyM0iGXee9eLsor8+OFTe1AW/modGb19eXihOkm3uZzqr91
uLxl7aKJALZNUwTRSMrM282GHlyxjxsCQDqrN9nyZDuxnxEkwlKg19/Ni0Ud1deApC8/7DoTkXb/
mtlD71/1Ry6tVsQ48UoPbzLhDnYh6wU9zK4t6cpa+q19m4FN/2pd2bpv9IZDnRjS0D8JwTL9Co92
Oh/EKiNfNF8D25ZN37Mv1G210/wOPSG4yYkwAsTdi27tLRhbdOKBvvVeeUGpVSel8O1Ed98LaQj6
tALBZih1ixdVmyPq0IN0wHXBRW+m78msZCfYx0xzUkbxEItguroVkMFdxiEV37EQzsJ7/TJTn1gB
tI5PQkAQJ5BiIvWd338k0Y5dcaP7UEonQ8ulO2SB6hkD21nP2yxsTn8EKqZ/EsDL2kI2pDWMnt0a
ZD4K2MIFl1s5KeFJbgHVhHPHzt0xCGVAnSmsHtlFY49tzvlzXZdK3wP0pHQtreUixI99XgKFLEw0
jS0J8D36V27uQ1gaR2GzeNNEyhzkEHajhEK5OY/aFA7I6KiDlbtBEWDzhf6wbxRajuPelOtViTal
NcItW6KPtYX1fbqT9UbvMdSzGtxhcH/L3Jq+Ldon9NoPNMTx+NqNprJ5ICMs6z4VYINExo1soCyp
qJu08+VS94CXkDibessyrpO87UZmj2NPlBjVdNe6fjqAESPb2d1gMiVPu6MFBK1avBpTPSi+Pd/w
lsb+rKbPYkqLfYz+7wc5+BJx9rfvSurg2c7n8TT8QE3wKqMG/xiQg16++JuLXfbXsH13aoYSpYa8
TH1v2GQrhJNnOxjO0VKKZePA3cniisfZtMvkrrOSBsXjUTf4+a6o12BtLHoRIKSWoDw3wDdFicJQ
WV9mouFvjWP3GZEA19VztCeGgf+eRjNVbwXTGuL14fmkTeJS0playETYgSiZx+tPicAOWRlIlCry
xOIOfTQxz5mUOF4yWPWGS0Z9ELNqbBc9m0edT/+gQ44gfCjMQm9x6JtaUDslWMaIQWbwLX6K43zz
9ahFAfm4eV5Q8p9Txmsep1Gw3RCe+xOLTaFAzlNycV8Y54G4CnjC791BadKV+yIvYI9vWYatEJH5
KpN6i9K86NEbFUjzvfPL4BFUjh1q1x+hp+Az0AaXtiixjcT6qk8n+dUJ5z9XF8DbbxByRx9Jn1PA
6qvYUNBTe3rzD0iQVgRRlUOBvJU/Ns/3ZoGHkA3mzj/au3FZQ34eH8giY8fgOegwpAuoSmVHindX
8/veYLzNa0pFpUZXz7hh9SaAKsD9BQwJ0l047iaQqKdVKU2ChGN2PZ5tbsRIfnd4y4rwzxxLdOgo
uwWb1oElvEsptJsTOc+gLTqDBElqKsFnrfxhp/hVE7l6ipd58sJsXQ/38WcA0FIw40XEgr1XI36h
UWQrTeEFSsTDbXKdQcLU5S0+LcZmHOP2W07yySyzCI+kKR6cim92hYt8He3EByiHwDSiQ01iKcwM
cCfpXuuC6x1CTkYbt5dp1AomZ5vPEAICpCQIcUTZMKY80pKKM1RhCJKRp1THlLzxTFXwueDepH0f
vsKTd/L5qz+8eIh4vaO4IQY8jO6VUsi26ihWSmNwsKE9zxWSyckdA7HmhjG5YWWUhT3YoEhUlFjo
lo2MhLijWrThAUw6pXZfv4gDfu1whRPHUm12Ei3WtbKpWm/cxSinyx80I5YsrHE9W++IeUI8qQgR
I4Go74XkuOux2x4qSsdhzeY3v+PfNPEsCxtNy45r82zXEMf8IiEI7mW+f/TVa4OuxWmCZi5ZmSQX
bfAf7EFiIReyFcYf71gYuTl/c0u5RSM7K2L5MAVnubDg9P+n7jCCmYIY+eXeMbfxUtfow0ZLSh2z
VwWakeMxrkXhsokAgWKxoXMDMuUxZh0yUIirn3hEWMXcvhARcA5HNdcW0wwdtvCqxcvY7PciuoPm
72/RLirXjSIVjUL8aF88QWqM7sRwjpT+51vjmG5/5Ar1jp06xu1fkurgU1qxEqpcIxPmiVC8zrAp
3ei116CBtRjJ281E/C3zrvU/Wksz/JP9u90UgZFpSb8pW+pwGxs6a/ktQDsF8Ygj+CIiqm3XyA3+
2JPUQL47P+3D03iENGQEwUACOsxmGcXtGlF/NeZSYOi5Bh5tBaK+gJlYB8RUgsWVZJbhnrzPIqBm
ajtUtcC1jxHZoWxuZ3XAuc8QCn3ycgAFvWy2M/wnFzFYNrLH+yiuW9kdKb9QJvZ/BcRXlaMtSy2W
bwV6IuhZHscsxOIgAJkUW2H0PWKX+33vQd1y0i0GDvB+jeyvShm0dqML4MzwlIfC+JnFM92waB+k
C8ve1DnDvgIHmpaRoAxUwo0LqAE4/zU5vemXsLlWEGapDtMl7x3pHBRASHWoDeta241u9Ra9jRhG
vYFzkTsLq/zkyzW/afCcAECMvDAiQmCJ8uzZrvw4+8vDumRHaxiNZm/zVAc8baZ/jFJlxruoEc62
Gzb5+EZkjgmk9x4Ke15EuZAKLXlYQj2ntHgJMsvhNVa9cr9UsiV30QkHiBwRFxqNbBAUyo8kjzQn
cRQ4n/cwaeX7uTWWS+gU075Kkr0hjTbBKlGBdssPwGQYFgMCO3gHYGr16EHuZ0ENZVDsk2bU7ych
imELLNBpdgs5cNVEq/1t3tlkqc7Ljh6l+bw0mxPGm1VnaW4bcwXZ43gMPyqXySZmdRfkj/sim006
IIsvGnkw/jIu1O6mWXzMrea5f3o6zmW84XfJfOJcn4r/kr551nkEjhVeuwyGV2Kn/idhk1g67MKO
+Jqp3Z6GAq0Tf/wn1s6EOo2r5LU0OzxfpEI+EGqFnxkTmBck4dZZ+4Sei99AXqaNW9xbXwMKdojr
SrGuWiOIYRfmGy+6CrciPoOdlV4guq60NjMtsT8+TyY1opYGYjv4Fc5ThC8QfPVsXeqZEpxG1Nbb
WzgUoBPlxh2bP/yc5LcYwAL+8H1BgODW4x/KCoJ0p526oaShmVhcCRQnaIV4OJ3ZDLgBWAMQK1z8
srJQLfO9rLsKBZZFsm+FXgAoz3c55fAd6SDABtuUWVMIPp5h1K34HNWTLdhjyTaFwFSAO8au9tID
RRlOku9CmdRPqPj7m/W6KJKRnHT7Ue3I9vmOaIgiOe7FwahOpUgtbWwcW1YT9SP+R+6IJAm0TyfG
gOfwTXjFBAsJ59eWk62ElPtjX+DG+7qpPsc5EKVjKF50wxYHuQezaQ10vQ7QMlzZ9QJL++jn2i3m
aJJ5i5tmHiGycq93Yw8A+yXLZ3uR7z9oZhS8+YPizFD0sXI4OhgdH5ckLeC5z9wEstIrtDi90EzC
vSdBlFJnG5ZFx0H1cXQwT1zYWjOGz7gtAtSO4Gh3iPil9Y0RUI6eqcsapHZ3G9nXxqLoUehxMyU6
P64cmY5AffpsLt008+ViGKFqpxgUrH+u2w5FfEOKxupCKi6tCYn3tLmywIzFmGpFkmitOvov+OXt
NtAeo8x1nfjfA8iv1WKPt/LcU4F//p+QvW6Aq0p5quyFH7BHO96vfmjiKpwKbQdCP4PMN7yw+1Fg
YiBZ+rlzBodwXB146rquBWD9Os5P6m9mQm/N24BKq0MvFpndLJdDyr8x3sjMTmECGIaYlZl3LVJL
eCrjjs0CcVhsLg4lzSvnpM9cYegT1X2UMEZ9Du2K4+R/KDC9cjjUiS85ZxzCvEgg2le5+YniDwIU
lGVpy2UZjiVXv1OwdLvaqSJpKRJ5SkwCJ4i00YVe3gnpxuq53qVWuoYGca6oU0exdNtYen6/qRXX
idXeY4jZua2eFM2KcZ4gCxfDvq0/+Idur8ZALhZRTQKz9cxcz4I4/VHPENzHBoBCttcsuu7LP8IV
OXeU2uqgI/mCBy9T+buortCbXGFpaV6IQ4lWGtXWcn7X9dh+mN0osTa/DUMWqURjT7AGnq9X+tf0
0M6Uc4W3lJ7XGTg51jZKFwxhVkrg/0DuJoacRiv20D66mEvJI0JnchXVaraImfr4PcalQRZyE7oN
YCrucXs9j5I3dZrXfxY2Cg0EKQiq7DV6mF0MrT1scthL0YcUyT7Ui2/mnoEEgoMY70DOj6gNbHPv
YfyBck+qe0a5+KC1WP/6MRzR7oaLx9+hHYNwad/8g+wgYKKbcCZjWYfo3dpxz7KTMS/r/G4/czTj
ndR9BtvuA5uc2xGeKSjKPdAJZ1pmCZ9TLFem6wElFUVSIujp/dnRX8uSbAwQdc3yOx1ZxUmtxmMX
hnQp0K2vjt7Q0cMjLYaEkF8jx7f4556P/a94lo6OOBD7sNdtH6DtnOow6OCrzurLhhswsnGl/ufQ
sByc0XDDm8vZj77zJot1eikzExjn5SCTi+vMIrEseKgdQFglzOhy3tTuhVXnWYyQso9v9l4WfC8h
a+lHINBHdyD0CFrbKg1Xuz/qqvjpJCi5xpeuIfqM4mzY0iSRTXw6kfWFWG4uktWGQce0W5bh/RHR
IkB7UhbWBeeR1/g2cXXFoc0T/bVBvZS8suLIWe50kBJDQJhBfd8gikl1XSIFc4Le0E6lTc6crVt9
v/ble0qCdG8/jTnoQ8/f28NdVEPC7XWYZb9kGSrIyUxDqZSyxdVybXPuk/DMOdCrb69Cq5wT58ZN
xZmcHMNp9iFgYIZeKZV/hz+9j3vV3YHQvR76ksqL9tgzyDCYhc4GFQO8ZuWzWe52QhmzBoWnfhTE
AZyiWnm8ITkifHWHhEuaLzego2jv9Zq8WEodo+iuMv3MSHrM6RN/DN98AN2bR7+9vKg4E5ufp/9B
6u8ti8KUE+5G25JHh/1m4+i+i92heR1wA9d0xIQuz4e95chrYTYW7vX566NiR786r7npmd60MfDO
LjfwmH1KG8qN0V1mu6srDiP8kOoYQnm4pu+azZrF9mmjamtDzwdN3oGBJZQjDTTmPdKog92Mmf+E
5x7zZzF/lWNxLEPM3eTmFsHodY17riLCf+Bfi5Cq+D42N9jk9W+PoS3k1PJ/1kA2KP52joAcBqYG
CdlFSbQARZfkX69QW1bAk1IgdD3ozmM/oDKoaq6DP0ZyMaaZckj8Q9Z2IujnHKGTQf+tLMpgYCUM
kg/Xte87/QqOBk4mRjQn4y/+bIzobjcaMrTusF1aQPxyoDnpJ5AhrkYShoRa36FTHsAsJlnH1eLg
/mErTiypx2C9Cnn8ikflyENI25NpdwuD11kdwHchNImFJOqUOzYJY12lUIzyhmfAziAv+x9gQ4ia
XeEDDwGLGWk9WgxWltGw+kLXXhxpNtV4xZiP/96GEolIk6wyHg3PQT5c2kCo01I6Yt7p/z+mjLyk
7VZr80REOqmokuFXLcJJ3CP4I4QT1onLUtSQKPo/fUGeZuKMHpGRK9o0uzobkfUwp8fxF/RJ2KvX
C8ICmnwXccGFCiRdAXDKXbCEiQ0ynAG0RKxlwy2zB58Z/Wx6IASs2zQ8F6TBSF9r7y+O/24Ud8Hg
HimKgUJPVnUg3/VRYrEj/cw5KwyY1Uof/mQAuxFdpOqUZcD8/aMH8FAw4OYH8kOGyt+3zhTl8uHS
N4bcuvBsKpL3FLbdXCV9YfWbI6K9FtvjLC5/JkzIpNl8tI5tBdeVV36wU6nMfc8M1UVa+r/ugPHi
pOe1/PDKevZ3ndermnHudWc/Tq3x9xzj6k6k5aM5TuVNgB/ShCRt53nKTKXa6wa/OFpenyVBErkr
sgrnRKaLyFtB/YR2T3hTfxJJnhwusi79hiA30LdmbyuqOyWmDLaWW8mkC03mNU9AB8Yk608EeYCl
zGfpwu/sMi8jSejxzt34Lkd8QYYt/rRSpsEcb/ZVEr7qFq544c9lIiAHsP5/fxece54jB7QOUvBU
SuZwH1pfKAjonzjoDum/FUOEouKzt2rp8j0Gp6WTAr/ogTkVOXGuH9hTl0ebVJwcZ7esnQpmNKHe
fB3h864G1cR2i5rxWYSF1rp9PEgElL9La2VHxLrvw8MNBXJXZBqAZ+H1i6AnyLyjZWoHKvfDB0fu
4jze7chVzMA93vPy5JF2SwCoiNYd+aVsf6Y683QuNk8s2qWfXOsBdTz3TiSa7s71c3EH/58Zlyxb
kbIAYNVsDJz/LSQkOP+aVY3/hK6dYug3u4eCUPV+JNUW0bgmn0GbdwriNkoeZvBBQ71VLDNThbRv
iEVaJiwYRdcSGgLJgLX1lyFP+7qVKTni8JBoCjUj+GexJGrAlzYUi6sJkzmJIFwPEtlc6+nGPjry
H5kGVIpJx2HilBc/7KYKdAAGLN1/cH7kxIAdwkBUuA1J1ujizGiTyfD5nTiBbXG9AkekaNOJuyjJ
kOCCdMbt7kYo5OkDP3Z0Y6bt1R7ToyAEVgLx//vzBxvI2tT3YrsxX5WF1spKI4aep/cnpXQo23e0
orAAiMOkr+maklubIluALDqvfr9ywBp9J0dcUYXz3Ka/OHxpiZJ0+/XJk4d++S5nmgef7uGYIgmA
CDSKgoo1O3U4URzK/yXngOAUZvoMqKBg9I3Rwz24pMZQkZt2N992D9AAVcuBVJMA5rajB93eXcK+
lN21f+EU1iufYUKBwD74BwTXSIVrQpyQ8y9Vmo7NwizoPyXNGHlJZSXW8benZ44KB5ToZeOTiWYL
RXMXXkb/5bmSk+PRjma9FRVzXRyKYCmqxw5b/k4ncNsJzK5uKjSyUzw4p5LaWrm90Axr6EGMxA/9
1Py1VDqOkRtMdrxCvoCkbMWDNRDobr/mumpdozuCzqspdII/jycDArHqHitFi77Tiu6vkmrnLb7O
75zUvP//+8Pad8oRR2547K1eHLkidLYYMV8+hauixf6fyFnYzlq36CB1sgRwFaEdLbqP/2S2pPxI
k2YieJR0wuh2uO3kyWflKQKoQhP6rhxBq0HPSgh1K+R8AMe8MowyDKmpWh/FV+zQEIUb+MQlkE4v
npu65CNEDTTzFcbQH7K/DIV2P2NnfaQ0vb7abvo4FL50ezaZEmi3XJs0xYjE4lRK7S98tI+5Liar
qsUfF7IX23mo/9CTBxV5CxZi+NrkEaxMIjDJHEoiC1r8BQTdHHI37O3jp1wMealzpfRW7w53Aj7V
SfBGZUnfytcHSvBg60P8yub/syZ1fCF8YzpU4V7gS5fDpb2g9UHy8kz964+h5EYVXH2Ev3k6FYVQ
rIongjP4y9Dy6QD8kcMDXWteI5WE0dH408+TRly1IgXsn/ujWM7nqcSCa5btZ6x7jxuwbEaO0LHF
jZRjHijgiiBoPxLwfOwlfVK47Rjdo8UYbSMEPD7DXeGDkU0JzJarXwx5bSYSVncdKNCnduwp63Xd
fZEGLKVP4k1uJ3JDMkWZJ5bbiSnpXes3DfSdap+dcgesMdGB2Xym/FwsUSCHBYRGfxTUE4Gp4o/N
QPBkXuldS1HFnGmsAidPUACTnpoXvTgd1QFjYKq4HQShXj7U4F9ngPvI6u59SSJfuo9i75w3XT7l
fyYUwIhtrIOOyfPqzUFNXrItb9mnqLEAZKzNvbYRUSc6LIyMupXBc6gBC4OtFWyMmnyQ/p6kqHa9
yWPoU8UlQ+w3vcKAWcYZ9p/IlUL8TnRI53uaavC5rc9Zbe/KoXN+2/SGrDtcW4XjpmadUBSm8TKV
LNnqA0Bk/paAe3CKoH4vLlIFK3KjkLdUoXBl150o4GsJ5ACnX9A+hM3sos7G/i6MYsCujPrZh0wd
oHtdDmLqWCAaxaZX6YZqBhHqMtVJVrZn9tgaQ8UxeHrKmL4k8K9EH/7poJ1vnkPMXvEBbKbMNJB2
pOvVhe9ZETAuP8LjnjETqgiy9FMTKU3I4rcE+cHi/YA0GGJhOY1KL6/0MKNl8zXXN0oX/KDXYj9s
K1DmPBi8URHFSqGdj7RU9+XeW5lebjVk00Ta3mqHd7E78eiCSuP8gA2/s/jSrZpVrHCGImCDZKVk
uEUIwV6s6ZJ4YLdmMoFfAlcNRggtGZWKf5HUfcYKMp0yYZ+g3Vn+C7pS7P/3JELGMAWbXjKEiy60
0MBg7PXSGwswQBS3ZU5+YzJ3bJ/DtS+WJBC/jXdF0ftDedP5tiAT0SjA8wHKx4DjW+l1pd0WbxY/
gwAaib+QDLmjwi+sQC8dJiL+BNUyGpDiAmrLncMBVcfLCJVRMdZEH3do59Vo321DzMYYRtVuxulu
sOKh25RHcKgYlFz/ksiD2/ahSvvtSDJvSto1u++GV5Mn0B/d/ap3KPkiX4Q3sZwoe10pIsMO+Z38
fGXcW7+HkzVp1W4+RB5htQ14Pasu5+PF06h4xabSs6DvCQhwad4rOWAG/yb8FJYdoqNPO5WlnEE6
7U3GWpKTeZB1m863i7OXkW9HIkc9GCI5wIUrJHzpxDK2mEXiGSbAHh05yYMa+bC4VDnYIDIByxWQ
ra3xwosDu3u/NvFejQ2XGLy/8er+UjtGiQH36XFDCOYY6+kKnOKRlJsTGPPDHUarHZCSY/QEmGma
mEqf5fgnvOt/Oe9qczpb0QVJtBjHcdKdpcLIOJ+DJJkJDwVXRExzLwNXuG46nSd7O8sOTo+SJ+cp
uyshEnC1WHBabPplZN01ZVhTtr1x8+4bg8+gmic0qiE35ljjbZ5bT6jn7f7OzEJ+ZZNw6d1z8vo2
32Ni6+e5rkIE6eWyAhS6ABgNkoePhK07KYD0e7WLsFu6bH1eOIUsWotO6bhuppHMJPsWPwkNGjEt
5bTFu97FWoykNTVwpwEjQrW9wkb3xG6SSQtq5sm6IqM3LzSCyHSgLvSVoxPADJnwZCXSbqSnyQib
MXHXKrjL0LjFf8eKzj0/pqSye/qI7DnMre2zcAlNS63kYTE5QooglFW+4HURePcNFru2LkzrTBqE
N583MhaXqXQYCFFwOP0i0ljzG/Gmetd2x2Vpl3r5c3KUl1dpy5lJbBVvn6RLiadQLek9qa/NTSy9
RbtteG39fIMrLzsoRZ7aY87pDy09/F8A01OTDWFlNxyc/M+4EPPsqMR/01+jtkEChxWpeKjl+CBT
IluLSCVnm62wcrre38TumGkYtZ06/lYjIOhnkOxWJW6CPLAjGDo1hFja+zZgwmO1VpNXhfQ8WhHK
NrV4EBV1vapw+G10e5W3AvwGGRgAUQn2ll856Xp/PU2QseILuMptKajxGdnKicaPtvTvOti1zOHx
EVZ/XBXMkVKtxqXWNfTDLlZAVlbG2yKEuJm+v0p6DzFPdmwlllp7xVZ91fz3XZYePDLFsKfp1tmZ
DtNZeXB74YGjdNzw3mr1PNenmWcoRdQFEFqwYefhO/aJGLNBJVOUxnggmrvxycfsPp1DWrHCV/Fq
h7wQ4vUcOeWnA7IJcVG1Tbo6WgerHoXeiYlkr0A94AtRK525oaxhmdFpusng9Yj+6+LKblXKnUGN
mxK+8hB5jV2I2PcDgdjQMYPVA8dC4DIuwqu2lCypgY5IOFQBXFanu9/cnJDAVKrnFBhtdNJowHiw
tKlx+CMQPcEwXjIWKzpo5cm6BzBy6J0GaRDD5AkwViGZlhYTy+mbrnL68pxLZQqNnzRtMB4jrZPk
X3km1R8jx5CdgSfXrhoxPZgoDmABb1tSFLKeT/lHusx4h1JB8+ALbT7z0gnL+VoG3xSGbIaUEMtT
i5P2gzp9fc5SXn7T4ItZhntXzdSzSWAxrOJhgGKCMGB7VWaJ2cHzyaqm4LbU4xt6Qg1kuSLiXBbb
vmwLwWb3lQR2t2WGJo50q7pKyVYLprm8d6sEvpOc9iteXqdJl9+Epb8UTCVnmqfBT6eY17hYzrOa
6ZrytoyGsAByhctLEXEdqP8vb785GrXYfwGMC18e7YtCL/x1wv+1KSe/qPfANkS3o3uzxesCVYNm
Hv0gWFcqcHoDjktmmNaOnCc5a+yn1s/xyNRORFk08j4KXHq/ixXHTGcVN8125mD/6WBNH/4cha2C
Z+gTVhj4BtBaEQTO11kfBd5DcQNa7Laa6hlSW2/SLJ++RvhsUhqN6c8VXYadmV1g3nffNG9Yl3FW
kcSUQguu8NkaeN0ITbgiW71Q+1aw4UO+FEHfU30mk09je85Y4nY3Q0ZJok3m7V6x9aGowe4MhVAg
R/4LMtyMiSYl0m1APBIyVZEqhmt5SlNiF0CwU0YEHaON/BnDntG4kbiwXu2yL/noFUg80rqZnGVq
Z2RPxpxtetrpYxF2CZ+C7AnspiId7b4inqcvL2XDvZlBIc/K8+8eXW7NMPEVhce9zvyfhjZWmiD0
lKwanx08ftM649ySFZmzxVANdqTC4MFrJPH/+nrlqIVeLlgMu16yfxcYC4XMrkMjYqOYP5x0CP2z
bTAS8cKQd+Nycb9Y+MOfBqZIISryWFE/Cki8RTIT76aVlJLM+HgbmQvnSE5W5/Uu+h4fhTJIZv4Q
fg1ShgA2QT3Gga3ZmZjDTnWNAj3Y+Suime6H+/LnyhfC83x+xp9xaCTSAsN5l+NPr6ScA/Ttc/LR
q9elrOybhSY+w3YxwTWLEIyNnomdg2gxuusINacjqaDOBMR4g7bQsT2pEvXHLXEXzdKeJVmoySrM
Wv4SvbVzIahBooAq/HZm7Pu7s7Gu2SUADAuxBa6E00E8fDgHfllhLBfwVMYmCloxId7JSY29yHQ7
qpBpCHALfuwAzmF/hWZT8tGq8ov7uu9b7q+4NgkW2gPmX4g4fIX/6PtjTUGO1SbARYhXZ6P31Ns+
XepJegLBArmiDy4VYdPFSt8AwkWj+NhCwT/yzwVcj+BT8NY1d4SFcR2vl0ZXxZWOmimcrRu+3IML
PGQAr1Dr5KrA5AQ/fMkvHzuiZBzJGWH1O6FqJJ9x7yJZ5PwVrxKzMmLHkQ+cva9XPzo0RaBjr5HH
ZEdMgfBaupED5m6EgwoRQrPsdIbUwgdtvRQZJB+HKNKMeyZ05aVJy0QlUl9EX5Z+bnBYq+zrg0lU
xSSMsrfUNvTrHatenXnqhs0RT3Q1qgDWXd9bYK/cED/qNQo6eNM8j5oyGHMszcu0ATELvLgj136c
5ZWvI2YE/sBGya5EB5Qih0WJw73iOmuky2zKeXlNuG+VVAVbLMMQlSelPWyaGM673JbuEUdlj76i
gkPeJe41ZLL7xAW0Loc/NKzipjsvz+eQg2VNeNmwT2U8PTO7g/2P7L9T+RA1EK0LV1oAAN5+VSMC
em0qilFnyYazCKFgEKsDyZ5aT+9FRKeF45FjTDHtZBb4cHN1PazM3y98IER3eSOQhL5WGB2Bz/et
zVnrnDZUvoX9jcyn57WwWEmS1Pf3FU2lFHgnLtgZ0gt53aU4Ug8uz72gsgCMev9hXN4QqS7dgoxU
Zqh3nDGkBz5xbrFE70wX6ICQVLJWLfTkB61zy5Dh4BSiK1o7JBu3MMDn79dgmJiuztDJvir7GBt8
pnABWm4bGYiqkGnKefJTbF6elYcGJ98jpCKNOYHp7Cip8i9hNxjvFrcqqCN7oM/Z01zQ6EquazHA
bLWY9xfCYERfnLG68uDAc5MjmpzRxprlttgDH3TGYiS3MiRfz2h+5ADtc0eC4Bpxpro3JJM31gsD
T6sFGvOwqnDOkZG31/7I98l+0w8GbOMgCPr34PF/VBrqQoQ7G5CNbVF2Dpg9Xq6FoV/PMH4wYyCK
tmZIy53T1ISAwh61mDAq8mm/z3vndPe1t3TKLlNtr7xaspb7N3rW//hbFyUZaP4DxIj0PwU6YO97
LRLlFYjk9/ulKtVispL+jbzGgk60ennVP7TMa9KPZNXUrOsra8lq576MSRY8e6NyeYPR07PdL0jo
JxajLYDZufY2giM4+NqGAz1AAmn9hKNva7l77q/GSEhiyCOrPpr+G0krJepsnVWtH2wvdhj9oy7u
qXbWUWA8o2uWmytGNmKQxq27NvcZF8aJymmNG22v4aW2eIOXY9G75JvuTFWh7ngkIpTq754H2tH7
PmSTCEMCqKMLaZsSab9/u4mQqxzVu3eULoO+5eBERzVuMLCDXOWodL4t+gYOyzToZV3SVa3jXt05
9n3VBOCQ9VksB2h2ALhSeWmZ0SD+G5v5O90hazqVCkvPCoouZf/D9fK20k8R4UcUlq7tk+5R8+QI
Ub63/38aO16fAZUQ4ct6hVOm3x2YMT4gObNZtFhj9eVh93bogwGhI5Tswvv7hls6W+PPNd7oWONv
uXRzACfLWJU7jxfs77PXa+2zrh2Lw3SszqbYXPO9MxM/jtAFJqVSWydbM9+mpOT7hQSlLUQ6IZyb
wIWR2YQZbMoOf1Y+0Id90b6upCtwCUMBY6Fm7nAx7lc7G7jsHP+jWcHKl7cAxtqHZme4w/sB7aUd
9mxOmvRjQZwwCs72dSkl23lTdwUbHYEw5zPeckwzSwsyPimLk8PrKn9bGM4e3BBKRRiJPfu4Tn3X
wyKmdm1v86dABrivtFnxNp/+Ygzl/nFwRMxHbcT7BLrlgClZpjwzpaDY3EN04sUg/85dBvgAp+iT
q35EiCO49ZK/SK1wWr/ovBDiugqeuWjdquDTrc+vj+E9wu9bsxV99dzgK4n8m6xEHO5u/FU2A/6U
IOawsyTs45GKsDMm8zU8S23bV3WM3/2y6D2RPPMk3+SDTBi7PRA/tD1NoxMYBMcYN9cerkiN+OL/
u8Rkwv2jFjNqgk3fYfGmZhGV97ixgno4yeR2bWGU+jvlBUYDFE4xf9PQmIVIvf3rxklCqcRvQ8LM
CcVCSzp5DzHA35k8pPgv50tzn7h9rzquVfQot5TQX4troOGE/co4oZ2S+CIAaDH4a/7ZVbsvhIWo
/ytX4ASRg+UBBQOGhD+ZroQnKUgMMXJywq8uhoGwzU2ZWcmxuzRgZmjDuzYVxse5A5i/QjF9dD5P
jz+ktz/CtKe2CO2takpvQWhHB/+hz7e2rXgCOvmZK6LPXN5LxL6lMqe2FEMFCrPNXnXP03/ziDwN
UblM1eVdkSqIN+1+lJAHDu/F+5KKc15N/KFnrsLKTFJ8A1lkFOnIfQwLkXe9Q56k0kQXpOmKubpx
nuSVvkUVUP9+AMiN8nhB77s2FW7rdr7RO56EbJWlSXxdtnqyppri4iZ1kUTb1OlQ/FqSg/spRXMJ
WAavv7QenxCicE5uh8SKXhcnOsuqe2HubQ/oP5ajxrdOkCxBUomGeePvyz8RJuXxc3X17OUyte71
fIN+tLONojED/r5o/1g2kbVp49DnSxNeknKe6KcNI/3aSgDS6tpRFxDyi9wjtDEhy03Yf/3UH495
2V2vYSd4ITuyzpcP+fvP84R3vQKtchSyCifsIdmqyujlC40LFuVXa5QZ0wLKXM2MjHvivMD/QW3W
ToyVleSnyU9jh6O6fAFHiqCM9E14POgvB9+QtxMQSGSClBOOQ4ZN2MlxjpiUzu+xbLj7jpS9TxSD
VFcUublMeINNJuxFYSmz/ESFC4stX1qnV2Pwoh1/VcWMaZrlYXiMQtZEWprQyRJqIHm6GjSoXcFT
UCvYg7dJZ60aqNHC/PKen209TyxjHODHlpgOsSp1PJF8qHODIY5mAQEZl0MPZj8EpnCusOFT7ztu
uxVedNJZf2LXufsplC+QN5QzYRITkofC6Yc8k87PPJkBgNvb2rGGpZBMrEgco5aIo7D8TThXEk0f
H0iseGgHblZ3nwH8jh3CKuJLpOzTDvltnmg/Gd8to7OSydsnmmnzxLi39kmqT9A2iCdQ4JWL7ZWf
oqSAjmDnDwmA8CLifMPdvmmw0Imi+wJGWGEY8gqPqBqDBA3tZW/++plO8luUfbDURVf5Fuqut7E2
MoIbnH2+LIEhaAnJEdzT1/8QinsAoMXOoDLKOnDK33FBW5msuv3l/NwemdwRlCt9bC3aGVtx6dYj
H2nADfiPCELdM+OA4UUPtcuX4MpOWIIFX232vk8jQCHjtpTRT8Xwke/QQwPzG5xl38/qujbeCNZf
VW5wvUb6dRMfiPMHMRw9EphI3Ak99c/fU7wpjls0hV/0stNt5LQo4lik7TZahhWE0HUa1kLa6w9X
V2bjPnE1KUTsxbcDwNZPrR0RxI/LP7DU+5uc+T1ed5vf3usAulqeMwYRF8VJ10iSbi7f3AyIX1Vz
FzTmGgFDPUbsjT+pU5/Il5mRBeb1iCUAkSlop1BO9bWLPjRLMYhf0JJ12g/2RhrTyW95Vx8O4m4f
keS+Ydux3aKD7Aa3VQD42jg74uvRpAZLtXFbBhh4IHEjN+Ax617yJWN/nx20dKtDzd8ozTdoBuew
q3gdOcpv69dTnfhK/F7u+5BzUz9skcOWarvgygK4U510+3DLxyNHWJtRb2EL8BwffpMesH7wL69/
1JSpCBVhRPPV6y+QlXsl65tlUTWrybibW1FVzIIuEloAT2Yim3u3amoorXPY/QcsY8r8JnBmUJzB
erHvUb3h5gE1ul0WAD6XxZhV9DTrhhonyEN7aYc/L6RhBVtBLRyBwOX/DjKulC6SrJDvugZlDjlq
wTPw+nmDQaPnRbuy+rl3lBTL7FQRdcdnuJQfcqTEXCtXsRxHSPungrPlzWePWeAz8bDFY6j9Jaxi
C68DwWLshhBN+YvMWnBMaE2GSMeGSeh5Psl2rI0i1Xs9gf6r3W9FKGhLaz9mZhdoQ79cfyy49Jwf
5l9RN3pvqcvi1f5NTkgKnp38pJ+B/oqQI2LeOSuetZkRLK1dwcKhGZwlFAiy0ZKweQwx4LtSp4Tp
FxSq6G94QLLP2IMxq7WV26lhVL29XsuL+HkWHxzwhJaEFeLCUKi4WEiarTQRApu9SFsF7XDXmumX
56vdEsycfCNrFtSow++saaV7xUOukP/YP6btlo+mgD7YpNB0dMIDS4/D8HFrxscwhRrU8NLMFOWl
sxVUq/9HO56jL9/iEO8fK3NmpHrfm39jHDg49gryn/bVS0wwzXi6tECUlhnDB/8BBv/u9jXL8iLN
su3k7dnJxYN2mfLSFcJvLGT6yByuFO0d/U6eXYJ5c5pWsmTLAucPgewbfK1f1RVfV6GOlmGZAGlW
qXXo+gN6jl0AesJoQYDCBXYfW2BU9tul2cj4hzAJ6JkkmMN/hEO5YrmqPqxFZxiaUfrBg0CTAwNl
5jKloWkDZAWoQ66oJ1CDq72ilAygNgMDbtcFd6bBSYmWUWmKez4ZX88clUgXlv8qMKi4o2Yv0OM8
5Zm06BsVO2u+ORkO3wSrKTelFR1UD58pwHKey1uWLSmrpZbrSYwCMSHSyJmmmBMTSZ+fYAFubp8G
x+xAlDD1DI7iobhAuNylizuRi06sqoq5PLSTNPB+XTs/L6Jz17KVz9CwlocK5wsqabZxzisE5oxA
2jHdvyjiPajNFEtNEyPqFvHqJI1sdDQENNdHjHg4/dAE/5Qf4RilDaBy+qxMi7EwBCsCruYJkAN+
ndgCvXuEx2/8KqNb9Q4VXG4pg5iFoL43enjjJ/xc9nrzRsirOC2pXg4PRsoLLJL1HHMj6ZD2Xb1Q
JaP+onMw2WqsVd17AYg2M33zl+HNg3WWd+iPDb1wT2A+FWJ3XaGqyOIaJIDuQNpaCiLET5XCSLnP
Yi/63YRnUzyqhzfyF8DSfzAQXGgwatZRuNM6ZUvPaJwPcmL5m0jtbl98mWVa4TNMBh47W+99KDI3
NwAdQ8CrKo3c7b798y7T9KlifY2iZZe7876pEo8rPtHOpl58n4H8FpSbNJjkPPcGyh4gxHeQAUrB
5jVE1Mb9XysXSLQZtBYsxluCH5OJcVd5rM3MqwvxbP7ucSO1ZvvvaN0htTFVdbBBIgeZohYDQNp1
+kZQ1jELElr4DH2WZqWCncdz4IZpdFkVlxWyXq9rvGE/ZbjqVGjK8maSmz3hZ+DK1E2v7izstGNt
oqjsfa5yxa50fT/jzVcx8EUmcDzs1eqXdHdlBsiIwe4fev1AwpxWzRBVye6kTggd9rH1XDamMip4
kHwEK8b5ySqTPPUU77KB/QkEqUyF0fJBGpdySYibRaF/6YCtfudTIzxAURZBJo/UXgq+jMTei1In
ZBt7LpYdpH21w22n+7ysx9yzWfQWUoCj7AXelTTVsFA6VrboowlZAHqCT/r2S5L0SZ7APkeidJdf
DAdmsK+5wCLSiLRN0ZZf3xIYRJFTyjERb1JrS2yWQbUhlOSqeFtEMGQyOYRbYac3sDHoLdH+BLH0
1WzbLqmG1pKo23sAabXDSlwIv5dZSxbArJULuLEvzRJg4GKRqBmkpOCEs8Lc7gPMAgIUo50kvzYL
aTeMevYN8mXiqQg3aAIfz6fd2kFt/lZglJ+CDvH/F7Qqn8ik4Vm3SfcqM0Y8IrZaGz4l57spIN/j
EjEKMpT2ksXhSAL+altkoOQ5WV/52pvRKW2S1ZBk/A4cyqSjy6TYWwUFOkYJVuhbaO3DMDLFWMqw
iy2CSEWvQ58G64t0LXm+1e6zbPF5UvLsh9zNFUmi9AC5YVFhWEwb1SLIUkTvR9iNfOCVfblgJA5U
bVt0/1ef8VC7Z3A3pBHRHhk+j61Hj4j7cQH6dC/cAheejdQ82WGZSbiwte2EPbiSp3dgRGpJkFGa
JxFc40q9IfIk7V6+6jiKt8SHtw/50jO0u5gXeP32z5W+9kgOfVye/veB7UeFkMGu8wl1IugJDPA6
s1x8D82Ds9Gr3qOTb3LdcG3E8pBXNstxKt+2d1HU40OhWZW+aVpKiF6H7yxgQrkZkrPq7R6UjlGb
sMvNPdeyqFWp8TuBVH6lCdFx/bhcbl39izGQ4SWes5eEfEP3AQnVpYtLIfdxATQXEdKNOCdyQXGU
HfcNRzOUn9n14oKWAH+tjRR8dpZqjLdNyEA+roFLQAzUlfK2T+7VWUEeBMycZ3b+jRK9/qYtZfMI
NZkELOuPuyrL1FI7fwLhVclfo22A2JFXBzVXDZ18477bCpmW1ket+VynfvdJms/uIFdNI/o4QPZZ
q4iLlPkR8lD0TLSsb+fznOtqZ8MFHGmETimOjUaoE9uUjYmZSj/LxJwdZdfKEsbo2OlCMLAEwtdF
HbK2CR1+EgDAy/dEdkfVjEhaikKnn05aPw9DlyI/m+zgSgjnKs2MPEoL7eBX1lts0NVkn7sOuqVR
y2jN8M9qPMZeZJWZC05XyOlLvuDkG8Z4gS74JQJ4Qgh1l1GM5erz/f68gTb8Lwv0Sirty+kBj4Rw
wvmKwlSRnpfPsCvDgFi0Q5Q2XEuFE+ZVJ45gcTGVwe/PzYE0HxSSSPs8XkfHTChHTt9fZ18a6FEC
lAFCTiWZ0RYfjJ7fcnMonRu3OUsJAztxLGy80IeJ4QlRRVry2u08Errphse9ot1eELgfL/3QYuKA
9n8ugb2e7FEtOT1vsLBgxSSHBj41vF8xLUWKvZLeOBG16qdd3TxHxRxrBdikLBEz6TFFn4Eou7dE
Ost334EjP8FLOuMKhnUCP/6l6JHLlCiojrmGGrMAypSPlKreAY6v5ZAtqs3urF5zqnPfrUo00aiz
qDLVRMVx4lOhgw8bWtd6k9QciBL9GBXWl64x3iN7ArCfQKOSdQOCSMb8cKsgH8JMaDcc1HWZnVkq
npdjo9bjMJGWihk6rsl+51cV8Dm1qcTK8WdHETp66dO4ds7ZMY+FcIcpzG6SdZpxjqrnQk/+n/Hf
w0HtRnCxnO8tZ2quymSQNr4Iyl+SzEPUs1MeTk47X9Ui6uVDrpjNQa/cHrzps/cuDSsLigXA2hlL
pBDqrjHsyZcZPfio9nr60BNojha7tFK5Gx6tEsSrVw4TiepkDofhZ2QaHYPF6PtExwY4FcCFmW7A
oD8TFylAoi+mkDKnZKliWxrvSsKriE/ohL6+oVgbOnfRJI/d8vY33FRrXZ2oehvKEKXrj3J7dgO9
3lTChoKND51d/mJtlyDC0E6PBd/nVxC2xVfEM9x6pEwSX5+TbgijQ4wetFLlRzKqwvr0UUXCbIdS
Hm/hn9CmYNTlgrXUPN300h5C44PMNnDhhpiOFIwkJngXHDWktGDImROBWwjKaRuFlndBihX8Sq1m
zye0/ECi7wTb5yc6A7YpbZwAWMQqm2zAX4+EpLg5nFXNIImljswpGbXBLnfEIK1XWC3cvZgLVezo
LbF/jXiaAfOoaEbWEOdcgVYSSoc1809YWUfFaKnrvFSm+AXDPCGz+5LCtdik3sU9nE7MvDHPnTgE
6tzVH0S5swPh2IUWR0GMMU746Dz9TrXyp589GH1redobjubllZwBAhKhxR9j5IXR/82xumNos+UY
KyrOaWCWlaxjXhH2/ePcNzK05t+0U+EgBXJSGhfwxH5bmrG9a+dv34GpWxMQZ2sleZn6jdTJvNVR
PE1VG1tUQsN1XSUdUGNPKPEGvldcVxk4lL9yYomyHKYn2f4LW57KP/uFGNhNzbLc29PVB7ejRzPb
jc1i82dH3BK+4XGRdfQJg1LYDbz391bM/fljQR1PEdKLu5RLYGyYdLXGmQOsrtO659VOD/Osx4kr
IrqN9I4pd8qoBbCEQ/NW7tbYqn0gOaMsofViJ5xPqxF0TD828BTQ6xUAh/hXT3CdEa4js8J3rSOU
u6EuhZvWiZuFegWiE8ApA+J9F7k0a9rzT7fzyxSEKP/h/kW+KIGhukfTPvnUvwuBceZpXjKTv1+F
RNKETXeMR3LBZZz+SJqtLiIJdHXQon9ug7m7uvxgFnL60k1cK93gjvZWQxXS6zw+9iAL/7DoJIF9
Vrg2BnKacFlWXI2DQWL35lbCXkkPsPWdbscorrh6R9Kd+UB6/1RhwSwSmGMQt6anM7W91AE58tcP
Rc2itJmSt1C3MTzVRP1uHsRJ07/hSSInEgSNbdVdBSlLTfLaXr4nWcTVdwAiJNvn5emWFPFtKW8Z
fG4g2mndIb2AGgAHPUqWtQv+BNr/kMpoGfDYrozOY6itucWZSnMyPXPEwLrmFq0m3+iezL85VWRr
Qhbr4wbRawiY4KthxpdCY/ai7XQ6s7k2nzL2CHfuTTvAoKJ9TAt4VCObe4C806kxdvPlryofxxYq
Cr9eemnlWzy55OQ3UT+QvhiX2O+NgALlGNK/xOUYmELEQREVido3AKJbCeEtd9o1sMrM/XPcPqh8
D7NICvxiZxuLmnlV0NuoXkLfaPWXNIUN+R1G6aJlsA4znG1hszogQa4+y2tHk29arGpGHzdoF+pB
h8Gx3fdevVT+q/xDzKUy8fC+Js5bSmZIwWEpzyn1CsBziOv6Apyc4HTaI6Mi75hapB1u2TsHXxh8
MtjrsN7KybF/+2T/3tguY9uZ1vgkAWcngtswdL6vyhkm5dRKWEhUBW2Bjp5o7BZwkX3aqWjH9Rz/
F+rXxw2oMThNF+hji2jR1plRHBSNmIaV19VEopCjjtZDY0qzR0mlpPrf1kInFT6enxeg8tPtlmil
DQpFvrqLbcj7ntxQkKEqOkMKailOQpd+kYQX/4woQGCzwcTU8oT/sNGDOI92jmO9Layf8pJVXfvh
HhG0lvAK8KvrcqP2g5GeLaND1FfXNLORaSZsNMVw2WGkt74nfk1d8hnnPZhygvTdvjOF3EAEFhB3
vY2jCHCnHX4ftkUWA6CNh75+vacmoI3wtfrd2ulPG+EV7ACuzw0KZR03fl3zJ4kBv1IJ1cwcjw+h
M7Z66Gi20fsHDghEM4OG2l1tDVgt7Jx48rA1rX79XLygiLnK3PBn2xNzw/+Bk4ksEonGYOoWDLQ+
h3IRIeqwJ3pnqD2P6d0okviuBvEdTBstyCEGXO4+SLJvp42O6N2SzvLu2ndpewSlc9A6eflwQat5
8aeqY2QQHuqja+M7/IFQslhVjPjInaoQe8Dh5wqQ7pMj55j/Pgc7Ija2u1mzEozLIgsphAN0LqKr
SuVSD3xqCie1c4XakUYOIrsfb/sJmTQCX0RXw8RHCkcWBDNDwaAlu/iKpuJE2HNqJSC8b5M4k7I1
x91rqtzW0bDKyANBUHdBWshm/Ir5cjS8fjsSxwYHQdkZ4en9tKc1yNRo9z0dXUlRQKO7qsEoc42k
nlql47TWLMXUQS/6vhE99hEeCOKpwY+f3uLCl18w8g61NHipfgXzdBFUAfauVPgbABT1pE/jaX9c
jY33d316SSTnaj8jZ00FDz8RuWlFAE6ny3g8JQUpfUy2CsChudsqDQgAJ5tknnDaFRwHvYakFuVB
SPGlUfJvirHy9DxXnSiHGasRhVVQBEl5b3gbLpDmvGV0JTioa5HdrdOiOkYLFnxQoVElPeoqcpGh
D2yYhxET1fryuAKjm/JKnPXsxqXdggHvdu2deNfFg8Hd5HQBNGqMDxS1gLQk1si+x/MsSUS/pBBZ
292hHyYcSvpH+VB6DIYrirwOE+W5igcx+3EvzArvW3XOA4TIb8JEUIxWXq9WgaJuCRg8CvERfpTx
M26QBdlKHlFDBZoZEBxNmR9UqRpvHZSUC1L7wFU39pfl+3UGiLiP3/M6iBD8JCBxJOU+jIaSByob
cDk2WQRaN4z2iEHqgUWHKAe3ptoYe102nhEsku7yza1THM9r0vZ/d3l6PK5AcAIN+8ZZpbyyEr2Q
BhxuttDZeuDe1l0tKf1Pb2J0YcCAlYGFaYdUcq6mh2sxFzP1DjtbnYT/GANGL1NVV0e+d27ZtHTW
3EpeMu8T8HockTscAwe13fww7BuOpWgFoAWW9BPN0A5HW916F0c6CvpTWwhHOBo0rIyTDjBdeJMM
gFSS49KVVbOf8MJucC3d6TL0g5f5BkAt9E47nG4c5GmjxmmjX5zP0xejBGl6q8Ey9GFGwI0qygLp
hsHcQ7ako05r43oO4O4aq1JCChJAIY2Ahs7Sk/AiUJBU8/cmpInYKtpKa9CWQYFUuUq8zCjmf/71
YGMnbwrYlpX4heh2iz5FIt7smRtAtFsk6IiaBmXqdBMcSnR8bfRy3UqN5rp3k8N0SVZz4Gl7mfX7
HmxOADmHT84dJ4LbSTirpcpcl8o/DzbCOOjAoLeY9JUqE16Ond3W0zotMe2OXIk1xi2qn3uw6q3R
1fQ25YGLaidi0lrCIygOzoxA+3CCpp5sVGuyTyjBHXIW8GP9/YAYKuRVdlIbrNaHPsklpU+ZKIHr
cobz8DoxtJVAMreFFX46CC9Vs/i8kkPAI7xwZZzTuYRmKMENNWihf+JF2ShohsVfTFvLKfwlMOS3
HvXsjGCIeaGpzxbUeGDXxAWsmxTBUte+x7d2LLeCdJj6nPIJiEu84s486fKvIO0Kpoe5qGXXDZB+
Roj6xjtzy7oS3X8thftywbxNDHzNvrnWxjlT4OYQ6t5xYhTa5k5tomlj4/eCj8Ic7RrB3WzDsLwU
HBafYB8ZCFxxwxchqO5NW4IRkiZ/rUoSrSsRs2b9s9ivXGrSp98xPXl9wyHTEwJRafycWAOXQkmc
vX82K4Eb+8Zab65h40ZuqWAp4LIo/n6Wcbmg8umkXyyvrtBDKVLcJzOs0fbrMIaDH08KZxiqu2GR
TgCyVW+wnA/KxamKbFY/4Qhi1M+tsnYhA6okAaE2/z8GM/rIdps/lLh7jV6h9Ngvwwc/5hTuFhSv
4UWr8mdI5pbRuzTgjhmon1A48Y90DC6qxOP+yJVtnjirqdTnFviUT4yU9syKn2k/faxChYS+iJnb
Aud2djmPbGiJPOqZ331olfo71qzRizwP9R2Qc3PMZ5Hhlq/TFaofFbc6+FCqFv3iD6+7SrG4ykM0
CSCTkZVihp+Hmf71Csy+nzUGufXunT8+p62iuISQaNTEo/VgQvIrMEytM4pwJ0UjyNOq29wceegb
Q83nrp156YOrRSIm4NKg7owAcjcnjIhXBEHc+QfOsQUpu+w3UXJLFErDbVVoRojN9Xr7dBQ1RQCN
+F8OleIUH4vYmFUplb+H3pkIKaGw9ROVV9Hic4gSU+ch+Rb75VC9b9K0wpl5Xri3lovCi7bJ85LZ
4SPQcKBD2XekF9/hhMaHQ9crXYufrQvDdYqvF7iLc2FpUovl5YYJiWXr+YBj7cpLLjbu9PPirtm0
jEinU9aagJh7bwcnFXOzhg6V0O9Z3xELJsCBMlRIPXRtgiHrXv5zknSiZ4DHirdbDZDLzpvo0Jf0
fNfSSgha+gxxznrArTmlfnwzQEzyeBdYdCBUyVB/9jqEhQPwiq457tXVlHJZ4Mz4ZBIthtLMMmrz
q3nhE8XsciOeHRXoLYreN+HL8LLTsUv8HFPyS30F3EN+hlNnhrLkiHH8qL7IyZD689sB6LFsvo6/
n0jzdGsOQpz46nKTmH8pff6GpayamhOO3QfpvI06l/ucalrb7Q9BCuGyHMSJe4mMJo8GIwecc402
FDtfDkP7ie6wYmsPj6PnldqoQxKv0CopTdp0/KrcE8uj+xqRwkO1uClCim8TWP2eNtF8QvubIaDm
GrU/Ic7yAtUWE3oVV7ZGoqVivJkWcRvnA/SZMT1GxaMS2OsYBy/M3cNzqKKekk1U8aDyBwNTnhY8
nT7406ld7y+M0wASsPymVDr5ZAIdxLNS0j6gITzhWvgDq+HPzDFRvNiUv1m4umgBafd2eNTfXij7
1b5aFo+cSJHE7sUe57XY9ADrjsMtbVvLN5mVQvT1IGS7UdqvmrMb00rNUc1CXQUMyetXiSJ98ybW
pX57RbFM0Lf0oScKZOIMH+kcQILUb7SCO81gOivvCXG4qn+U9Mu0Jw4kg/agFUY/NbufA0mfFP3A
6OnnuQmDtdUishebDsIou5wYnR0t9C2C234hUSXjmmFsnuQ3gjv7s/FPVi9vyBsxtL6xp6OzMwRL
4IyHoOmRYGugxjn7uOfqTrzx983DLHNdShgzo71BqoihhpZrH/+sm0lMkWb5+W/92gfSVd9Uv7bU
VTJ5zp1P/cKVYFjvz/j6WSOQI806lZn/zU/9Q8Wsc90PQzuc9b83FCGRlJm4g1FBIr+8wLwGCepm
ZOndhG6ULNDCeyetxnc+XMFnSntXWhuwBGWgimzmJJy3pcNIj/ti4Z5pyiER7Axb/BqoHuaAr0Z9
XqmJxNuL7ga3lGCKiOdppsCl9I2zvHjK6dMmZ5V2/VLUMpih6I1qTAdwuQdiVwPxOjIgNUmhv05N
IIDGgV3DFz5fJNO+eQNEytiZlJF2O/Lpz9iKt3751smZugfim0nLbFC94bOXe+bDUdLC80bYd3DV
vry7DwrlDp3BOQ6L5Jz+BUVdrIk7kQM7z9pGiwTFklbMs/86rJem+uZiNqj13udVpE6ngM6JYsxZ
tCRMUQt73qKZlZ3Gl0+36FPl5pkbS2BmYWUMh5mtzKhlDpraxYtOoTklQGHV0wWx0WhMtFqzpv1Z
aIY5ynPfHgXMwirCnrsEwzkJs+2W36I/SQiy6IE+Ri2xuY1AijpPR7eHl6t+Qol8IoP7gsRjUp1v
LbqDr2bDdAD0owVHqiQF8FiV+6OykX3fhtgYiMvJdR7mpSeDrnu1+SMNS/Amf47GuYB0m2SUIzLa
ZPOw3o83JQGwJ67NhTdlM/KvNUrGW4YSP/bE+vx9gkkMiMMzCiHEaO1xb3uSCmb4LvQWTar6nSmE
N3CywP7PUqgA0cm8jt9zWFFuYfn+eLdYETjl8+J1i74fQ35jrzPgJbYKC2XwKwI32fHbmBxriVR6
y+x/q0cfBW8E4yf02VhCpJQ/jBR73bQ0SHwH8lXov7j2X36c/3gV+h3vd8Vy0eOeK7EwH7wTSdlt
etGqi1im2dBjgZysRVnoWoDMeNJNlBo0O5wDLcXC39Lbl9DRIkxhVOPLnXHQddEkN9jvTpdAfEVv
q3MB+Osg76EyvFgimWJQMmoJRjZiNf8/g4L3EC6BBYUxU1HyBUgOqHXUjFPlnnguRn1ihWS7+DmU
/2F006udJctD4eKlO87TNo9SY5WV4YdjYP1XcJC5YqFRu/2f0bFGAD0BFi07XCdWycnSRbXCzXjx
7O7dhG9AuNiiMLqG5kmpg4ZQ0KqUHN3EiaIes8dPz+mmw3lTcCv38JAL7VhmGvoZyvQIZr2bUUAt
i/TqWfPxpsVmv2zDQvAvW+5yol91LtBL4I3/Gp/dmWw0cbBALeXHy6W3V5x5VXCqoGlV12+x5+Yz
djH56Tc1US8y11KFMUc8snqAin5OPuGnk1Vdz+wjTROucVTFmaXkUxSi7zqNdmneKBsjpcGDKXQN
2y0/0jFX8Z0bigSf79Sup/G4J9eRJadJQjriXhzn75LKZOqGxflDD9kWMh0bBcYrhWCyfWSHQXYX
IALi2c8ULNZUK+J0gsSFfjdxGdUt2Be0O2PmnhOTdi26iEOBy/ElyA+v8lXEGKdkA/zLpDN6p3+5
PozkJBwca8ahQD3ftMrjB9i/wpXf4i/b63aXC+9ASmW+WGwvjYnezrbLg2pnGsnjd7tKU1dZ/gmr
h58QpJhRkdlsnb74Q55+oNbAi2mDcc+Wk6nxhPqUTxWDQ5zu5e1qjUuQmAGhsHtC9NIonicHpyHP
nK2h9JwFkeiLhPOnFMTUNI48T0eZVUWfEAe/o4m8xZEVFtNt3WCV6v7/XaprQQaEcou8mXhbYSUC
g2UnGqbeV3dcg9ruUO+miNWYqEpqn1nqbVnQcRbJcW0sY48strruy0w43oo6i6k9GsV6blTQMjy9
pF3QAJEFLHPj1paMYcHY5i0kcBNC0UgJh8LH7zuDiiQx3HmorIs0oU83IxfKJ8UJLRN3bkMozCDH
iJXuSypx8sk12hs42htKxrCaAwx4TPuuWmEzfwFXRPTzRv07jteVkWVITj/pKjFj8jCfS2AUUzBe
ZM2PgyWe7h1EpIPToh7MIAweLLRcCawgveRp02V3CkBChOPG0DQfc81v3NdibgpFDZD8VaH3O3r2
iY6I/nCixrAo599V0pORwaj3EY2XxFzs1MwJQnV7oKqbdHFYYGj3q7ZpMtgb8okKw6+JHdY7mjJ7
uy7QyjzWMuX2IfWfvZQnuvhmLBd1RwlZ7B9gaQdY3+NCsVQYa9Y3qoNvHvqt2cXvGR0aW+i1GJ1F
Nr/mKYf6PqTC/039VSaX8sPeZ9P8Ke3+zOrwS65SGzDgVJwHNfAu3Og9umc2amLpZZ349Cn+SgYq
AP2dxQQ6aHBgJtF6bZiA7z8vsMMSFQuApl89IpVu70iKAfJOhW9gUuHrqAiuboVuejVkFq68LV8f
332RV5JTF2JdfFyUkQLX1lqIn6lPPRFjB5JiWrQwFV5yAWelBnVTJsiCJBKa5f54vseeZe5uV7e2
VAMVDJjajhwaOji8KsZrS/hp30NASS9/Zhfn465X/s2cU3xce2UKYrEZn8wjv9cwwxEXYgZIVpbT
QLr6AMN1eDtSYGk+bZF3F5cNlq8whP6qdWnQ5D2+UCrTgeIi5j1P/mBXslflibVTY/Gj3/Cl1Alr
Rk14qyDjQGPVZCBZoEuRDXmfcZ2O3gOQIEdpJ49kfK6zyoEePmWr9UIUc8Am09zOtciWj/z+Ony/
eCms3gBizK9MksSNDvQ1PJnx0IaOFbta0oyogIHy0rRjGdhjqKbNR8jn+gXgOe1mxQl+V9tPRbiq
nOEao0agE/4peNA8dEpgplAMJiQBUM/sNR9/t159VzXL+0pH0G5QtBjjyUzGs8Iy0BsqA00JLE0h
9acSHwL3gWsMKyDmTCHlbCHzL1AnWTbDmNz7VSIw4pMtEUCPjQYYBAb2UvEWv/3pV9dwi0I0ZIdO
etbxuC8857JKFxdiZSIaeZfuEDnNayh8RqQpLWvYiQYPt5XJroR+JyLlP6O20WT2hQ712ye1z/Qf
H9l+l1Fzlm3MjC/V1agIUtlrHkkB48lN1Dh97gtmr5OrfPLMp+fa9Me/XvNw/zgSavlFSI3sAkqv
TTL8IA8iKnXvmKvrBAgL8F+AnmAcianYjTWDB2PhM8ROW9ATLLSNADOkFd/6n06crx2yadFgEfH/
ijb8pkh7zcLTYQtJoxQ8qtBtzdZ7KXI36vs3hhp3Td2np0JKyz31cwN+U6qp447a4Z0yLPg5z3am
iKV725Yydxi0gLlmzhiyF2Hhum6PmkW+dE3FrVwyLDNA5levLqR39i5lNbjANq6avuG9ZXSJIjul
l6R0U7oRVdQ26MWtttsLdoqvLiPrkPML9yspuRAYaStc/Ypf2AAxbrS3OUR2PK16WwnY45H1JXba
WQ31hLtMLPjlTaIds7Igo3agG+57O1HvuThRvHQyUZQiKgdq53YodaflxM6P6bwkKhNVzW7IowiE
xlhWYPqL6+oKSqsEQm2C/9NOHV/oR/jy9YPNI+fBw5GWfc94TBS4s0n5EitJkb+KNi0jVZq5qjR6
fewGMH9W7sEZ6JWwFCqwP+A6CZE3kwrajN5ddFXhn7J2Yig7eVY25Bn8llFPhhBRM9szGAG78cc3
hNy6l74/f4b8o+mcxODSElH+Qhk5k9WvRTHjKwlKhe3wduxkrMpqaEZpAMkBj0YCnnORYPhGdADv
qqnuwHK3Xhab7kDoiZE0xsCSGvuKcV+c6WX61Yng2ENLsmH8ciNN9B0JhcGBBCPa0MKJ5rD8lbqf
yASu1Evzsw0MfbrC5fxKYqbSKjP81jl6WRQh+cALRUKcfzgjKh1ynzLKaxcP8qvOH/e0Tm3FtMWh
j4Rn1FFredFPW64qU+H/kBSd9OstMuhZ734+af598YP9IdJWArhVtUXtlSWvHOrnjuDhErKkbLtj
uIdNDTcanarcCKh4XXOx+agg/y7GpkcmZbgGlrMzaaemXtTgKMt64FT1J1c2JbBjjUNgFQDQoNQI
BWF7wanjv9KVfWbaf/LwBA3gjuVUs587VlzkiSEdgLzEDnHIjWC/wkRlwvtU3Eh/C7rjdFuygpC0
B40FyD3XgVScx4E6NSpD621tNs2tp0k4yqszpTNLCMphEmB/Ps6ExKhSCST7bW6QUqRrTmfxejXV
aFOeGgI2xdN0v+XgYXEguBDqFvXEpzjAT7IIG53X5PLZIJTsAGSu7gkpX3QDUeKwMfBJFRitXzjB
bb/uohi+z2b07nSLAn/JvVzx1WCyKS9r7+R/pupTlbwd9oYHNCH+C+HYE8hZ25dwrs/L4BuVbISm
4QYH/4Ae06V+eqsfKXHRDb2ec+ocTzjYuUswzt5hgaczAiVdZ6V453Cw4q2+b1g6k5cA+ysRwZQv
+EFY9kmuA3Iu/HMCRtvE/eclZD9lejo1Df8oJPicxLF8QI1v0Wl8tpEQY9xNJIs14HTNXHVpThq4
j57qg5+n7GDXiai8777M/ceA6sufqAQe1rQOAmZi3M10zEW1/nAmwinFfsKlgiJb4ihXr6jPG9Gp
MCW2X5v1LGs53A7GxDKAZnvugGgkKlDIotF2xFuhpr7T7zdwRlvR/LSI+l+gRRjyskorMh8zwaFo
jnEjBhnFbgh3T0Q/m+mqJ6HLVfNIJyq42GEiyDu+QZFpu0QlOhckNTJEodBeUOBaqzYGmKZzCc1W
hfNdEfRGXjIKhe9tpgqQibxcvXPzK+d5EiSQlQP3AJr3KjG1Iewdtn/o7/cpj6Sz9xRmFeQYLf2A
0jeQZb4nFPRQb4CVncvtAjltiENs/rrvlMVMFWoIdc6AHBkwB5kDoGlB7NQr2PeDRy1tUJtby4eB
Iy0uH6LyXXN+YpyL7s5W2hehYirrla9WYcVd0Lqq4RFqar3zJrnUJLfniG6hAt4xECMxa3XydnIB
pjCHHBUkUw2ntreAFNUUpEEkyFaZTY25guqn7CRGDZG+hdFzefmx+9sLlUSbB9Vl7AiG7k2QJay9
kRh0FtYiaQmW9EwTdWP0Uaw+CAFe1+YM4162m6Ux77N2GXuI+CrCjQWDvavtudkDEhVt5zp0D3yL
pGhvCoTOIihhnwPdjlP9byPXM8OK1Y9muzw+dyXKyui5k59pYTfps6FaWAIhW3CR7PA70aNZqR7o
UnDW3q7YSLYtmDW5vKiZI5lCOrv7bMLHcdRMyMD0hdI1Gw10YzK1K7+N5bMxim0br4Ky5y+p9kIz
0ts4/8VuEeBJS+uh6EDAicV4IHFX6CbNPAjnRpEb+UPIVM2bHvST2pv9aROhrZzsYlR4ZCMsGinR
2+uv/CvI1JaEvRTvtanR/FhXG/+aqQz8rXsafdnkSe4PvJi0ABbkT7dqFdtI6utkZmkSm0xYc8Iw
B/VvmrasHRVg33NjswUq30HABWGGxsZ9j8v7kJDNscH/sgbV9MDA+mTJvTLLOXpycTYMbNwp8D7K
46Rj4J1pTrPRx4MDGXui5tlj3yqsNj3+zH+oGTMhdcLlKDD5ueX30hMS1pn0aWnnVUZL73PKd4UA
e1VEeZ5fyRJYuWlJ51PHnzkcKPfX0yCqhsrExumsei1SN5ktakUL188NkYpPNLZLuu0gbZ3kGR2b
7Sb957vLqhRngGZ5JCcdramOE0gcouVMiYRiAxNTncAvaUTT0898hRwaI6ZG7lnUnbQ0hwOCdVMf
p5ThVotOJvW99hboox+tyG0tD6KwupKXX/H+uxb9QvoJ/RE8F8vfG/JlGD/gRTLOiGF+XyXpZtpy
CYvieUpLe/u6oQgAKH6Zqc56T3O8McvtxbdFjcfSHkWi3PcsnuKoB48aVVfND8es4NmFpLwxDPX1
eSVS68Va9eToZNXSAXO24t8QW849wODGeB0dT8zKgu5hd15dupzeLJXyWqnM06Hfj5E+jQehKiQI
TzNbqQnpTIJZFhx9OXl8QAoS3sk6Bf3RxQPvlWB9p1zuz4rltRciGnyhCOdUm/1S86UYZI1qGlqL
WPIRR3DooWMtxPAbb57OogiJUjhoKO5PWBgzOgXyTgT6Bn6IpcI5/wv2wg51fFrGSD0txuZT1usF
OyAiqNwKPGV0jwuXsANbv4Sy5Yew31x4dE/wLRJcOAfF971ljSj05V+j0c4SDGdshUtztnTDcnm9
tAbp1hIK19p7tkUxdUpFyuq7rxdwNEAOrrg059MpvjFLLt6zKvCNRkJdyMDUYHirw0afQm+V5eOi
LusMadtfz+MepO97T+u0VyMFClPa4HJ6de8wHQg3uZYSgxDy8+VutBiEw0UslyxKRCgJbvg68ggp
5izy2GQeyjnojsY/vG786W9+V3AD6uUAufhtPuYZj04AFJ2YNIo5uCq5mcg6XVzdQcQ+8Berdvbz
NTIh4gZ7UIPUr9iam/C//lFJZ3qhlRoaAUOZNg7hd33kPoCLjl2VWKVZdlkXm1FFiClqHaMPNWbf
v0jpV2iEuwtfdN26nZWG+eyEG06bkfNEgiznFSZBX8BrCsTFmZknHiW5hV/vC3nemKcwWxRZuLkl
8JLX5JZ0qRKkaqGwKZf7O+/KRUQv3P4j7+e2iuiq/pOoSf1fXRPmQ9NqBfOSkTxR3ncdb3VY9xBU
1wXDdseTZCX5Du8JeC0NjL8NnPmEquPrAjtZvQ8zbk/KTvJAx/uYJUiUwCqNI2ZUw916BBsADzQk
+69mmfhVL0eQPSa+qTpImxqrupKEsSqIakaLIj3/nwsEtdbK0TOsXOjpDltWHG9T7yNmqzM1ryVL
e4LfPX092G/rO0IknPzhXOguD/cgdpWIYimqKghD8kP6U86eiWSswGfRYm8pr02G/qBLOJdt7sN7
KKy4lCPiy0y9oKRv+dYoz/Denb77dcW6JbljJ1o8A+jFGweNqv1un6RScG2uB3cXZQXdYlnzMCTe
mAVqWZVlTcSxyrDj7H+mnU2S4drZkNng66DdjLiLku2KkosFHGbXNQ4JuZZPjMAecKlTj7xp14VU
kXCI1i1S9bqTTOK5E4Oo7MlhRm90Ab1P+QWWFzd2+bGi+7vXgBfhdsVRFXRmRYF9Sn9/iu6Zv6Bc
MgQOte2jXZfu7HkZOM5rsmqCVXLj3GHWjtJJvD0fkPviT/B8WMjNfc1uAyM2mjJ70h6rA5+IW3vQ
e8vu1Ph7t1SWVVCvruzxp98dx2601xvLaVSRFF4X6zJMVKR8CORRNz8a/ZD0+npGcN+mtJ1ePbTV
XXazMauJy9sQW0imqPpnL5teAMzv2DXkG/Mx0txEtjMLU60hURBxl1cHF16X6NHQsZ2UkygHT4QN
6nPGuyaZO15vSatLcY6l1Ev1J7AlFs51Zu9M6XggqoAoqhEzvKhRDWkjxmwpNfxMB+aZmNssybQb
hpxEXljjfWctJiyC2LwVhvvqRuxZCnOEXMuMWyqlm+pIKrK0g+/+ZJJDmduq6UwEiT2muFi7YsRO
FvgYRCh4Kef3ZIAl3cR8O3q5ey+4Np1mw3OQkYegvV2cGKJ4Q/diUhHL9COlRbvT9qHvE9e31luE
yS0AWSdnKp2JzQ/l7/7hAO42AqqNlftsED+pI4mpLWUz50bzi4YsBPSRi20Ydj5KlOby9pxNvgKu
Wl6EVtcCP7Vq9cP+Z9BGYReSn0Prec+EJlBUx5CkEFe4kiRZrXR8spYqssTUy/UguXUvnBJ072gE
UxeAl0oe1wxZ4RXuaMUORT9YsI7j4dW1G6hFDelsTcf7uj7yseNtGB/pjfh2WblbZT5p4rdeEA2Q
8ombL/Avx37quE7J0Ll2flaAAcLIMcsZ6qe7kjPDtYDXSj/V7/3Y7upFaQQef6zsX+/zDYHjhJIC
tFByLxH3BnrbP+ZNgbeNtIFE5SGHokYgNreHJHcDEdfQZRqFpzmQ5/iE3/1O3pBf1bcsd1gu+VVR
RUBAL8T4c71S2CrPLWngyH70Zp5OSBtt9lG45R/aeRYfst6WrP0u6XYDqCjKJs65BkFokNv81gqK
hM/iK0W7YmsN38QZYdaCUtsoBxeNOJTrxEd44l9HU35jUiIcw+O7gJa31+WoBmJpw4pr4geM9skO
smLLr16KstjuE3rk+hDGDzxgHX07rYpRLcDjwaZJ5jXKgLXt5UwBmzqYEqWSPzAp338RK2h6l8il
DsYnzzi2ECpAGmLRyEKBH1pZjXqy/7gJbIgpoc2AeY7eFLf31/mpaOFZ3Ctz2749tuqFjnHhUES+
KxspFCTvZ/mQ5ZZwvS9d5Fefe3664DwnFkwtfi2tIss+QKIQOHH176ZOXc8Rlz25fcgFeMG973bV
+HDromHDg/nA4T0Osiwq5DxQZENPtmloTpTCrObTTaenlfXMvd7AQjeCYqYvV5+m+8Ru/DYly9py
F9ATAuzafEFnQ4vxVAsqLh80G0EiiHsX0ytYnOyNMZw9mjrTZ9mN1A3r0G/SW3t8fbuTAgY9GOeb
PnfNqI9wi06aoI0JwX48IiQz48LKCwEWgPZ548toVJak5gKgR5mCcR3V2lOfGqTHLi9tyNoYbgyv
Xg01xWclkZ+s87LZdMVqXFNMtgvJjkJ1PGcXpi0F8hgqcLYm6MmrNFmphX6wh5Qsrpwt9fWADhYu
xF9llTuHdRbLdMB1eZk++Fz7JrX7T22hPFZKGJeDQ2c9twIHgk25fEy6GrBa3SgNhQ0aTAfEH6b5
zapnMhPvG1DcH42E9hY0ithFWShVmwc2EhS/VspV0X4qDkVxaMYhIj4cx+UsIajXaMYMZrSZSfL+
CdxLTwKptJr4f7XPFLJK1hOghZHXMW8kqsWIrxr5NzgLTa/KR7ez5I1l2sUEkP0Q/gdThQC1sxPh
pXovhT2eNHq/Q+ToH3pR6CRP1XaBOhMSRNgXpkY0x4MmXRUkE1GdZFtleutR3FsF0lsXWA6xhbpo
aIpdU3PsUBdktjBfdmhFVhimt6y9tYny+ZTDsodOaWs/kM7Jhf6xbaa/OPavJqxL3oTDZUiHkb22
CBdmPPHYgX9UYPFDObnES48+VMprldqVgBURNXFJTrkZc46hyp3He0nxrjI5XWpHRq0sCWad85as
kQlHZhSF+PNDuaBxO6+5uuePs4iEWwdNaw2G5fm+iRBX4ByB8f+VuATJ0MaViBtcy/syKbLCvEcJ
cD+Qr8px0nA8j9NDH43tqgF/g6l4xdGG8nFKHbwf3fZWZLAOVIAQUZcYDoBV10GgyRjdGttrc312
2vgOESRxgOcCWlYW0hoPga4BZVYJaqxsawL9TE0wqdoJ96MVy4Hrh//c9J4uSUapJXH4Tn0sWC6r
luJ3bq7XeY4FRpYnri4EG2qCO3fF3GAMAX5/DHZ+tFkkkNORdjsCy1IuOogiKGR4ZwCUyt03USRl
6Z5KpwHQFBHWiQL90/q62cq+ojHnXo1bVASt2GF5Pc3AHy5YaJ6M1N2XFnDqJ0CW0Z3bQato5wl0
4nMWt1GF1nP0L0XtrDGEj66TDCJYNLGleAFz9t6r/CpilAJuM9rGq0PobbZeBPIf2SCyVs56e9yO
YtcWwAoEsT4Pwn8EWydPC9q5rrwMTFOz4J60XLocpD7+NKNoo/4s4Xj9gGLteCNedmPnuAvbACuj
d11pTwhpxr0aiHY29Q9EFVmok26UYmi9weBbMYOXYk1GY6scOPknYjnB0KmUklVTRbPg8EPCmwNF
yHVgSmF82PSjwkIwRjz4lstq0id6Q5mKqLnbC2A8AD32Np5k7m3Bg7yMXajABkGjcMTTJUaj4iWz
uN59htTUh4NZQaPaimJSw8GMCTTDKo/tjSaB47Pe0/qsvaSVYE5xgfDANYJlWy1LpUhuuuCk/qr1
r0PZPQ8viSdaY1oOJ2aUarpmQykPo6eJEKzL962PAGAXsQSOUkxPZHOh/4hxmYTnKRC8vhh6NQQQ
r7j+sNRfXa8bLZ8HYjgWvlz9RMvNyn95WwguP2JvQbZ4FIi7RxXTVpR/K07RIaskz3IHIXKlBlGv
jvTUqNNCHuIRKnAUU83ESQdgPaFd/S3sL52Bi8ovVCZwyil9OjYJ6nNyrlV60i/zwHOQTdYgD0kJ
O6aLZ5arubd4DCuCE7BwTpOVul7otPj4rIcaWeudUF8yW370j0voQiYlQ/F3BsGbUyX6YZe8qItY
ft+xFaoNtVkh1H3xqeBrK0kBrVaKYe/ycuaThJs3AapKS39y3XoLn4XzZYhivXHKwiUYLoIagSyf
IvZpQzgQmcmqvYlE/V745+IVbiwb3eSSZLYVG3zHcVd34VDxH01KFXXjM3j83IfHLEfRJiQsfkOA
ZoVW+JE0pcp/cMNMJ1VhVMgtdqUOl58EPWkIkW6SxlVqvAln5k956Ony1GbnON+s13F5Ef/2zSIY
hu77G9X+Ue70tGFJwechrX9yAIumyR0rIrlAgWPJ6unAY2gArNfXCWoHaQy3d0kFhCzTnTwGFWqe
6Sps9uXBBxSj6PxkjRNm+1muYl920ygucHoC38DpH2Gv3whLxGEGKnifCLDJwkZgordCm0dsVkbW
iNlDY3tsiChWqGTK+XVQpq6Yacudojfcs5UwUBfAeBzm8aqAaX0wleCJgw4hFaGQjvFv0Y1MkFhr
7jV3njXAC3/1JxsZShgbKheIsEjUfLtgTMqM4b9En4JXM4Zn6+PEBqCPKJGSvWf1tSWVN5pVAFxO
Wke4AnYYzrYeEPnO0ibGy6OcsI9MgMSMebCKHDuJG3tdIH966Zpm2ncSOacffPvPAFGNUC4vC2pk
1BbV+UdG9IVg9dSUXFwQK7liMmO1OUpY7nsmNYjURhYksFqwmZ3/SID4tnnIyChxpWLRK3zistSF
GDukh+NEaz/ud2o7stcvk0eKD6PycLTQYXSr/mvOmw8AGvTVvCclr5tkx5H7OQyK9gymFHsMElWA
IskjJoeKQrtSdCMxuzlRJyB+A/4NpqHy2P65oHkvgqFljOnIPftNS+xea2qD/aL2HLX361mGbYgW
3v+6WUChb1qtgALYplsulRtwZSKKCBO5nZtD6uFcNEjY2ArGLQWRMmluu19uRLbx8Sv+5G7nX9Qa
bvAzYUBklu7XvfUujzr9FgFabTV4zy67oxGzJ9/miG4l96n5ToSb/vzC/nuS8cOMWiASHtE6lx9i
XFDRCQa9wjNX37YlIvADn2A0N1Hg26AeXyxBx8tvT25AXw529rlcq8MisbDd5rWQWNo7FDTObiHB
CGQg47Uvd1r2Pjjui29Y1UhuIE82DzvUkgxUzwtvXPcH4iuzrxnRsIXPArPJHS7fsFodyF0+Q6BI
4e220SZ/WAEGUoDxuiZiJiiat2N5Si9VO99XSZu/5SmZDPfJhnnFFq9d5xdJZMzEQv7+uj+QKqTd
dNv3hg97iYFyeimuYeDXtpXzV/cLyrcct3bHfVGfcQ8tFD235SVOj3pDXlYXXAfi4KRrGyBdOn/2
etXeX+tmCGIK3AfwbVNjfy/RgYd5d9nzroyZIe0BOTiXgz2IOIN9HsfZWIzmjU+2X6icrhlMIff7
e+sDbNPPIYINwVIDGuIVV7tcsUWB+n+DKk31sT1ZPfw0fTS5TaXAIM3PEqLR9Zq8KxAcR2+GoYcO
H/XC48hO9EKgV22tpgwl6yOtU1DhxQDO43iQlouzXjJLZ0U76gc1LhQY7cwRQw2Ub0Uja/r9tfU5
Q1qNJRF8luTvZrakVxIstkjelXvBOeupqrX/T2GSKSlc6s9RCmzz01G374qp5/oRY/7hYJkvkBJf
J+ZrFrlPbwD2g+RK7xHMBZJ6LWzbSlZXwo5NUY/JYeIkVZtGnGaI0XazVTnFx6nupc9iB/FuxdMJ
DM/syELvfH/e9mm+dE+kzmTrezbLlZOWjqejT/5SFnBxh9RRh6NK3VVCrd4tCxJwILhw5z+nzJga
lgHLjIV2hmv5+aUmUDnLuHpckG1H/0Lu33ZXHYBJyCtG/VSyNHEI8SZavdBgPdUsO4hRUyxGY7nX
pUV+9mFw4xmC6kbRxnks5iLwny84C3vzjq3+KPs0tD0zKAzrn9BYA3QlkcDf9JNSc8qVfHbc13+6
NMpzQ/6Hab4unJEqtUQV4UuDCTLZw78DtFOwRH9vkvCNPNbfbPUkADCLhE+kGGhL1BJFbhjywpCx
ovNkPoi4QKD5oE5c9NQWJ4lNqKNxQLLD9xVVTfbbegiYsYDeskOQXIeXTOjLhMAUTejquxZ6my26
nJYxBun4+hxV/b8DFwKXcCPi6XPi8BnZoNM2TCcxbt4SsDg40QbQUEuftgvDVoINUQ6jtPlj8mJu
+4wIFiPctqplEGWjLcDPBiRd0oGMrifzVhWyA2jbuGne2FvVesLuRuuVFNYqAvvL/l3xpvpvloK4
y+a7xgJ1E7Y8nV8163i+E/tOELy9eQLnQdKVOddMDzNLXotwDhivBvzucLskLA++qRpW6QY6kJz/
K1TtB6SKbiUvT4grxzf2dw5gkMUzxC181EhxqZWbdxkmyxYQGWdv9f0F+YDGC2Dnv7h1uvnqqgCP
YD0wxisLRRXLaUSkqhH4ep5zpaiMHX08yF+ep9VXCEOcR9pTSCCsmV9L2e5OpCskakon2UOBCeoj
S9dRhlmVlNzL96n41IKny8El81ZK3H39s3QVdOM0WoPmYu7gNSgA49pDq51Pm/q3ahSrVqq5T8ed
VDWtYnXedHeXHuTb0jqdmd/7csaLfhwHm5jIpYg9LUjmKvL5M9EZNfhKt/L2hD0pOKVywudA4TVR
ML65mty7uTKtao4gIzObzbI4KfzeL+lMQju6ZAKXAIliQHs+4dngZxUOC7TZFsFnO3harWBkZY/6
efarx0DwYoudNWJGN20OL4L8vytPzVIZW6vSzzXUAlyS4XY5IMGJgl4vazYqBfhRJ977NkVUYNey
xmlZtLUGLyrUlsxv/hg6Q15h9yI3/v19D/8eYHT7EExi+Vf6GkguVR5hgT1WS11hVO1GLJ4jUsuS
tkbLg3UYXicWXp6MjtPaFrY6JzTuzIRWHc4fujeNZfCuTk2YbJJiQLAHFPb8xtrAv5Rv05WWUQL2
2F4sKBrhTNGFEuJllV+SLfKvfwWYsNpPP94xGKTxCFvrTqR+1kqquCt5wIT6lER48wyNIXt3v01B
3nyQzmW/jLXtcLT7wkKbe9VI9FddZ4ZnfPI0zwwTe9O8JT4Sp3JSSZA3H3d4BadwqW4YGSDLbTJd
Uh0omCHsJzMZELS4D/sRdx8pcT5soUJXBW08YZlAbYGqwNUyezK3AMXQ0JnsG2pi9kwBvp2lFkW5
ovsGU3+BdG0zL1BQtnWsgO6fWNVpXcBiIrohLbk43xo+uL/KDrEfnJ9Xp/4Ta0tIl3KFpdvF9P6p
urTybR9rNyCn60Af7ulWRU5sTWNR/+LDJqru1vaX0eS/Q3J12xL6PRaDizRn2pJxWj0dkKcV9tzy
XmwrQx7VTCE/Uf7iaJYPkblpdTJoFcyYaNAJEnqXcG0eIblAgmONTNNVhFo4TFMK0xJwlaJ+TJhN
K7YrfRlcr9IDm7YiVp2fP9IBnkLbEgPfLp1CuN3OEaCkHYEXoikcdW1dxhjc3BbcY7m5lumoYQyY
PBLGMYVcXnugDPwLB/SziHfsASYjbgGNlARerTmsPz8PmQ/2brRDOmYfQmTVtLN1i1fahZIzAmTh
u757Yox+6ZZmrjjj+G6kubdvg0HZlQMxkr/cYx96iiCyZpD0HQBgbGjda73GBOcTawhLEYCNmF3C
dPAKHhRw1NfANyImLNSqjqPof974Ftfs+DZzdvVGIdwev6GXTnpTk/JoydnHtD3naVpFykSvWkDN
eXrr7K54GAynTePW2MgQXZ4vQzPEoj3Ia+2NGEq2Ls+N2FTDuRgWbsV3Rgw2yCGkxyNTiwqejg+Y
vgDcnxBLJF/5orQ9xjRZqzHCeLPmh5lVCnhipDSsiFmctPNBmGDOc9uNiVoBen8/gbhQF5AAF7o0
RkX7dR9kJYH4ve97Zwzz7baVuPcq/PyVxhXZm9yuipyNB+4kMXVsODGKUIoMBVPLGBfbKxmQpz6v
BTAIN1pFp+wUSeXijrrUPt21tJ8D+wdTtX2UaMKAp/PsOx0JvH4/zyGR8b6q9MYOY5i9klFzL+B2
e8FPH2+Qh6OrWxP5Z0RnTZ2+QBWWLg73mGb05n/3mmTqJgJ5n9PYjGYegkUIwLJ15q7viLQ5+hOj
NuxA2lAggiCV091UphEHw+UWFitfLS0RBsxL2v+61LIc/uhohlEtr8kw+hPRJ7n3pusdENvXvK9R
L7RgxpPS/mvue7QqAaYfDmb84ctdShzw4WyMkGxuFwgnFc4hSB0/2m6zPcXiSVI+nNH0F4Vi1DFi
tK8bPpmoqv9mT3GHpEcGnAcLW3k/pNgrfa4MQGxlcqeHQQ25oJqYJ+ClbwOj8nfPG1StcFVyXKBx
ot8ijEjVd2Pmgq9FJmlfU2oVmHie/7t9ujreRQIquS7Ks+iMjYF/0My8mcW5Y8ymXhN4nL+QVYo5
4ug4wrC9dfreTjqESBNrRJnvP3WZgh8gwmDKYFgoUMRtrt4rPX2PD8wPiZbSAGHQe4QyvJai3jAY
KH1oWZRmTs4ZXR3OPwIR/XP1u92ZDe8PVgk6KE5cJE85vHC+D2++uzl0Qt73yAyA9WGeL5+V7HH+
Uvt6lacjionj262WQX8e/gYqxIp9Fvo8MpCwIf5Uxn02f/93Q3BGqhucpfO5mnFYDH6Si0vxewPC
AJvBa4CxQOlYq9q8Sue3OWShkhzp++wOahHhYPxQaS6jebcSyq/EtS7VHPmgyJYw2jLm3bVQ85du
CdK/neKMkeAyTZm4kZ0ewsMOnnklpXibZMz4QHSZsdtL8pJck2Paauf+0d7YcGmkPbjBNIwWSDAF
v3t9eKfxRNbgz7nislYayqImgDt91id0nVGfbCpn7PE3vnnUl1jYgarSnH6gszTXAH9yTcDkHxR1
TgExwEyTeIHcwOLegh2acv10bGplJI2TXILDEJVAn1FJgUMoqxRH4QmPAN1qrGCfr5EAwLoU2lhJ
Sk7oVqgXGuW6r2Tx7w9N8j5SbZ4aqzJA/xhTkRHJWA5Ht7zPxPUN4UrLigHZGmi2KzBj1CMzJ6sJ
jCj5EpL0aeu3iow6aUiwBVlDnM3z2V/H9tuSdYGhPWfh7mJO0AStN3IyrHTpW13E4+ZfGHXJo4p3
4IrwtAnqgheNXdd8lGUsNK8sXeaTfHeY6VkXK02iDa+vP9N6c+j5U4SV8Nuj30GeBy2+xJ0rB9Nz
+X72tE//XyUFQPuy8KBqkOep6DQb5wanGMFU6x/eEH2hr8RK4QwzlrMJA1MVPkguvxb6kbynvHJR
mcojcO9WdVuhorkLNbd+FC4UloJ6briJwzR7bAcLEuDRMuyoDbaakdiqLQ+8mBWR4koxBMue8uV5
XB4Te2cESe9OpTlIE0ZnldfvKIE6sCAxuNQhLuOMNgmhMtGDwJxb4PuVeq0cadi9HPZ3Qx7GqOmV
lXy+usY1bl3xHqW9B/73s6S3RwILrZnd+uKxc4s/hb5QDkRPhAC0R9S7q5bHGmv2vhgkG73jHCdD
TgOrH6OX4Ed2d3/sNlejNz8d3H32ryK00aZc5UQgGYNPhVMBeXyuXld+bXbM701eUcGpnkvz9LYk
O52QMH+wZ5AwsAO6sUgfgNcymbTlNVJlw/XCfU/mYkhRiVRRFFucFXiFaR9wf+c5FhPzoL4ZXqKm
refFQ4RalmitB5ETLAN75lXiRPxQh1dtUGo29SmCzT9oLKEziZjii7ovdwe1jJcKjgMkK1DqAK6k
y5IpnRtQOGxChypGflM1RsqywzCOmGCS0PXNXQ9vWJZM8HHaFzLgqtrA0HSEhQdwKQdl2f/b2Lp6
W8FEcGZMsd1mZOYMYijYm2QUPEhEuyDMEpu+F0aPZcN5+lJxjlF19fUWc2tnOEv9pAu/DRQp9EBt
AhD19Zuo/NsZ6krdS1DkvBmJWWwktP4hSuDJc2V6SEDyXx2t9Bpt7KHYY7cS96T4neL3k7tucocW
z1JkFxV7cXMB4zBVV4Od1Ozt59DdExmYXskRMvA+3CCQQV1Ku9e3PaffRkKHlyQamevnPk8HV2tf
ibHzEdYbjASLj1lv2S7UHMnQZf+2d+ylGTsdxvaL5r8ZPgcMTDIBno0YSmQ5MkV1T2gOan/mrkBE
0sRl9m2x9+UATSBxZXYmW8+i/yJBi2ZBY8NGAT/dpVM5x/uBVGw36Qitlx4VYHGAdEcPNzK2QRHT
p+6SR7B5XWXe12ZtTvmF2iqZ/m0uuDNx0LVJXCHFE9mvfo1C4LxVVxrRTi70wm/gmsv7rvvKwaoY
S0JX2fkmg5VYtVozKvpC9joJklaHqjJ/AXodZWkHr+97FJPeGI1bRfbkH5rAsHs2gM2n73CHZHDS
cBAk0E38gFgsH1IXz9mfKLG8CuMh8NsxvZFh1ewQyDt+o2R0/snIgEueQTXgNHkB+iVjYYrlvaws
irXe1u1SBufWAJgAfdUwjyGpwSSXc2pHSJ3dS838Cz+6lTJixZbtaqYsshTqhWOynOk+0fi1AiT5
sQHg7YEMwGaVf2bfs4LitYv51pNgPmwE5X39H4TXBeoiEhn03Nyf1tEUv3xjd2wUJEKrx6++Fkc8
e+lxNRy/bu2ua78gn6g70+1i+UI+oqprTxEDyblIxv+SedlE/c2jgM3sFsNHVX6lQY6G6H7upBet
lMVb8+xb5FLMBxN3+np3b2ACcVgFXbCCH0IRlsPkBTfeNy68wmOZzQUOYbrZOLbd2ifajpa6MULD
nGcFk8Rk4o/VAckIPkSpoG/A0iBdXCkPaDDuvjsDFvtzDOvrIEKtkvyo7RhzLFtiINCL1oY4367X
QYuaQ6zZ4cuHZF6INXbqfbqMdTKzn0dGrA3LhauATGiz02kLqt5bu7CWFoxPLKd3anMIUkqNbMjP
UoqS4ynZskTNb7OTwjuZp9Xwmvgw3gU2TAcW0UPODaUBfsz+6zY3srJEVWou6RsJXITmetOvcuoT
BuucNop2VjVy4yug1nS0+GFDF04ZyNMlGK10//pKGzry7wQ4ZZFYI/HMxiFYAAo5x3YNnFYbvZzI
v4NcQjZxf9cAOhCLuAMFyKAcsTNEPAo1zY7BeUEXnk+sIcCzTq84AKu0rLByHT60dj5mVSHGYy9f
J/x1ylbcmo4cQxwBFgHF8PXz2gO8BjQXEosdFgU/EakILyKNF3JxTGVdPEFvCOeULG3bj4418l6H
YAtPiYnBPFTLGQHqrg2ir5UhJ3c/Hccz0DZpymZmmLxgHn7Nkn/HzmnYo0W1NAkXAfs22E16LoUo
EDN56nY8t6rS7bu61eZSqKoRDqFwzltlHwQNr17ZflNRO1gweIiBgCJo/nju4XxPxoKz0+O8/57M
tJe78jesi30ibbJBbU5p8nfP6bRRBqWmQFQUOI39GER3Hcc6Q7WmRzYHAFuCc4fm0HihRvCv0s/k
eAUNJtnyash5HdJpU9JMLpcLTvIn4pNSIbAsgB0Yogd6gKW1cQDtyfBbfjKibxbjAglOzE68JwqG
Zcsv1N3Nhtoeux8lA6+jeSWM4AKBBO6YcATXIZdke+8ZZzC+Flc6ISyvWuytV+G5OZ0RmOIFH+IB
qXlXGOGk51wx0OkDqg2pfa3YPbO+UCMtomh8UExYo5M8brzTxk6EzqOqLQX1kMJ5sdqZd3uAXVCf
RQZ8tLy3qhcNRuMWy6xj9Qf/SFoiASdH35xeKuvhmrlFmMNqK5P94mfeDO1Xw7LPmp0fMyS3rEOr
omQHihOHZQDujSpiHZ/LQj9b//z/KnqaFYeCK3cd0nhR90Wl++IySPUIyzB8jRyRhBR1vhi19ZH5
XGMt3Lu17mzGIynmYcwVcmjgKqJF0JMZN6x1usNM8WlHVoFcDeKLSrpohirzyVvb6nB+KgFFC6r9
mgDM8MxoqGXJZHGq2hRHyLo5g9FV11eoMTaMzK7aREBqEr+tnYyskpkIE1fXpWiT8lzKMQTfU9/t
S5r/30AXfO6Bp5mSgIn/czqfWzM403eM/msmnsSJ/NJ1Y9u90GWK+H5skUE8KFts8uOY3B4GTAMz
yx8iUeY5YTso8yFDEijXLoH5DBseYq9RESm9bApO8AvLvcnaBhIldjIqCu6NeiIpbMoC28bIUegW
pDGiIWg/gk0wP+oqPvcQHcktcQAZdzWGxhsAMkvDTV80TQq0P8VvXchcXd9F+KW3toC8EoxowaAt
+gVP5HUoNop0e/qp6lPFJiWDMjbD20qdyFCc947uVLxhwrKxqftHMo/zS4ar8tV5s6LuQ+SzvSit
xe1jzlxROR619dNxkeiuREVv+V+WAMLQIgtTLdqgPYGCWy+gr6yiKO8Ige7Ri3vl2iwRAdReejh8
pDAlVhFdXHKpR+jnq1qNJzRwp2ZwnekH5NqRUYPjAfuLXl/1tHV+wNAEkCcm4DRlDwESMvWYEiN1
O1wbrXwxCpJNcyC5lXKk0Kq3tT2o3LFhwWLhzq3urh7B2zF4FJSJnlu83tZe6cziitNCoz6FmEUo
jAE7eT0kkhu3VS5zVm2ZxE3bfKsttczSxqr3ywNSlqVDDwCp4uDoCtRLkePKqyMmDpCPOLvG80Fm
k3KAg2MtHvCAWLGksSDeQMYej1F31qYz6quXa/WvuUOxyDBj6wjXNk8z6rUoiv25tIvvtanz8KUk
PHZKPD2OzaOeIR8Xfh9BzpsAEpknlK7FlQ1TYgmPHxkXkn6x2O9/sjpG8w13oDCYILQqF8VbfzWW
z02iL9DjnjvquCOFAUHIAY8mWr+uX6R1yC2+iudlzSm+/ow4CZrKJ3o7Yr++hL0RFgDlTLOE2ykF
q46uPWHFKvvb6/Nw45fNNe6He+ZfY1nOYUSIrKJ2AW8NsTee2l+guPFgTR00AH1KXHI2JFRoqsYr
SD4pHGaQiSaDe5n2MJ/eMeBjDTln76DY3anwPurObBi1mHn7Ba0Qa26y4u0trdPyJpf23fdGBDDm
NzxvhcNtn4QAo4nbVEYaoG5lrWE16C3R9k4lbpYcSbFDKFYkbEHyDa3au75LI13hTNjm4uvPAbLd
tXkov6fkrqLvgrbsxuuZomgbF0+VlJHSS95jdvP7QfqmJbFpRy2X9PfsI7Hvi1cIRvnN0O8sgRUE
cdb+85HUfgg0NZG0fTL9wNJFkP2vLCqEfVjzdBy/+Jymj0LNlVbOY5EAlWEjuFwMfN+Ccdx8fB1Q
J2cgjB6HuhLu0TRStP4pv9JeKRtNJdhQYyHetjZtUxlbMn5gGN72Wyxvp3EGJAqKWVD67QReN09v
dOcLED7v1PdC4BplXcwsqbx9n0Li3dJihrNTUYrbLsYoQzV0M5LYvD2nThiKAmWOIhhCm8NDi/+D
1YI28i34aL7IGmQjbxFE5FhIXB9j0fQ3AD8vQfltb9osdGvKUNQu4Ghx7ZLA8xXyObfRXRYyspoi
dLPsczFwkTM88sC0a9U/YevN70ubk13ix/lj7LXiwNUxeRX+REbfBlenV9YgJvq697j9/LIiTBdz
85IX17gjbmG8O3ww0t5GnZEvg9lNZddlxPNCuEBSRtqfdU3AvhMfbUP7pfDQyTwDw74o4c37BCfB
T+SHczWVhuDAbD6nDzpLqBrsEdj3bEnbpcrKVJJxMYJIDQnTMIFmNpVbaCfOYyH/aJFmPV6zENJQ
df5ojqhHDCdcwnRBEESUN/N5pvcZmnCigYASmqU/njyo+s/Fodz0becaRz0546dqEMt6SkpLxpIi
/oOpLKTkDK4xUDk1Vu4zrHs7vkyMHlMWTdMplSl7WdZI5vlEHADY1Aw43src382oo4NCMwKMUGXT
xFC/7mgEqvc/hYBHz3bNhme9gCrK2DWYVwLFgkTG49mWrbEJa5kAR/WUPeeUhDpVVMGsPXOLJmIx
I4J8nz90z0SZWVL/A7qz6WLlx1NxFYFR6cVCK+B6tH2WZxCEL68MX498K4sljlXvCj0smDjjrcTH
xbFQUfLbXyuUJ4giyNlJSRy2x2JJIrd4wgGZLbdMCmhEBzRLSqQNUx+XLu125v3S1IkE6Es9P0oU
xaieWmDxSV+Zrw/aEmNqKaFZRX1xYe6/TAGfRLislCk2dp9//ptsroxMZPDezitmlWVgQzPEk1SS
InUIfeGLnCeI50xT4tpX7uIESGpRSY36+KP09gy9kD0Icw/GCx8i5N4k7qPVvT4Cih2KdcjxPcEJ
241tc6T9aMCOriO0nSanyhvWc2CX1gxRbhxCQfvpl4fJCSpczX2GWay227ivMrNmh9DGK+xtWRdv
kN4hFYNzZLMepVT8pqzV3OF1GMo6pqh+eMJTY4TxX84SITeO4vR+qQ4PronV2dx97fj4IHMJ13xp
tzmh9okWM3wmsBWjT+RSOiT+rZ/XsUIbuylEcQRGpuopfeeIAzsfHgWOUZYtuqNYS+PYxPfo/C8Z
4MgmcKLFq9GWqgsLR3GQyMFViesXtmVFVicV/HzzhJRJRrbPNf8EvO7eh/UIn0yg6h9myvZx9vBA
5TBm3kiTZ5tT/3lBVaelFe7oBo9qotcUwoa93QZnBKuZJWVzG8uTxlrEQPgj4WZD6PNOGknxTMLu
jCr9BHZJa0+5dW75dz+PXMsFEOKmURjfLiuv4L3a+breg96Bg39fe0cOhrp5dL2+yo3HNX6i3dFA
2wvfWQ4lpOIIxkD8UzgN0QZtXsutpzRfY3SMM9tyS9E5mETr7KrsJH74tLZykZQ7q5ArrclVU9KG
p43kBWizqStyQ+gmclweduwqpuJ8M0oXduJ6RJdJhUDvuAz8nyX81Mn60CLzXDx4JPuJuws9lprk
d2SF42oImkRp8ZI2Sn3gpiZA+lXAz1uuawpHUfOVXK6+ipUft1YWejmhzn1y5xij+A1Vg6irJOM2
/Ukbi/mlSNcB31cp/UyNpYzQL3Xt9OSX6RpRCNJC037eJ6OSuHeHuV1eV432DISjvjQ2Pi6oFmqu
wFHjWX7wsBhgiE+AAW3A+mpusWE5jtHPvXWB3p1yo3ThHrV2qOiA70IdDpC1TjKoTAk1nBkX22gV
bFx8a/9ekoMnAhOvyqYr6zS/KHM6reRIpHBwTeSWReTE+fsd3nmKwaawHazZmfGv+/hNYSBFQEVH
y1/+fR9ZusjT3kBIK8j9NO16uf8OyNTUKyhvZJQ6UBX58KOcvQPhEnvHiGC0w8Wg1r9qxcOA9b/t
TgKdum8noGxwpZW1VfFda4ZYosnVeSiKVuVdGEooMunV0h7fIarqACvRY0zSs3iWoSjtPne4eHOT
8WfdN0TEzjgYFjeUD+cMlF3txi0kVfitKW7JY4mZDSH9UOVRpz++CIN6nbX0dFxkfJKUjQwQNSvG
iY2aOii/EzV+mTMfFAEypeqwTRer+S+zcqgC14TJwgJoO6/HKnNcuy6fNo1oy2Lls2OTRGwIQsoa
QHsPerJEbnqfxI+6rdi5u40RmjY6HAqB7zhyJW2zyOIUgY23Ao7KoW3+tblEBqMCP2cP54yf+Cti
Skr1mPGvDaWjxE2iCMJyeNFvsV3qPOCuuJNh1TmBXiwfPP5SyJYaXRe41hEVtKpr+ebjyN+SB3Lh
Jb95B1vodp/OAhGUyJ1zR8acjK2pwItB6oOmw5lyfh9ylqAmCveFfHaxmLE0F2iDzxV/8aA18lIQ
RgK6RJ6M0egh39VsVRosTKivFB6FUHigTVF/WiK/ncORQhKjrP8reqi9qhS3b62B2ke8McacIoLT
d2NyLJPM8tn+zRa5+Cm63h2CZz2xGuryphB2TdVxClfot77wgo/gHnl/IDPtcssIlWUwgI1R+Tz7
+LiGvUwb0746k/zRIv6KtHsbx54FqIWu2KbjHd3MNaHj0LBTL9mJas243cYXkvzexeTCuKRVzZIi
+svCtVgE3IfTpCFoNjnRYQrQPwvQkc+IxNS8Xc48SmSVl5gsCmNIbHO2UwifP1YIAU3oko8xtS5V
QIsSkesL36UBeSGvE2jl1RVEX3YaqP5rRRNfSGN6oD2qxx+4y8o5IQSjJjzpP5ybdufWCc0qkS6h
DdUid2XVi6JlPsTP0RkZ/8ZxwMscnJD972rVATbiD5z4rVa2rb8oD4xXyet1f3pZShUPih3H4j1h
Lbfue0dd9kJVXs7Ydsc8Sm2TBmpNoCkMPKfyRMmesgA5bIUAT4aBqnvvqsoO8fbUEg/TpIntrOIq
noj5TVTGgI2YPZPY/a+7hv7G6OfbGdQkEEJD8pLN3N2XExXsTmtK9UBqlwT2Wi6irqb7koM0lX6w
9+Rqq802upoW/EQY9JanYTNJQy6LjiHWlEqVyrDP1bvTXLwqmszP7dbVhZDnH+R4irZrSZWtR1V2
G6vNtizDncOTh0woJ6geKhXkzAtrF5z7ykOXXR+EnjqtKLyNRt+ufzOuDIE3kOkSHN7pG8lRcDNw
Av1aaXBsf8EUoLzzf7itfBV1FTrKwx+hp91S8og1BjeK6FpxVHB0WyznRh6r7obFcUDnuc9mwVH4
KbbpfWkT7D4a+NewJkzsajD3WR3HBfC4TsZ9TsUaE1W2ORkPtNV8nifCKotT93id/g6sx5c3uj0E
31UUDV+uGhjECX8oZjBJPWzyeJYpavAWHlWpyOYUbcFUTq6VGPX9SNk8BHny4MmPL41/toUMre1+
qAyJ7ugtwoig9fZ7nkoVbQlwVpBKHPQTbAuxK0bvKJ1yCgGraWN6z8bSAMo9sa5l+blkf/FhqlDS
XQEFkbvvs7tDj3J4uU3idIjKWmzFjhPYOpmH1qpCsGFn+NGdBBuvrI0kCCVPKpEJPWMlGQNxmAi4
jqAY5GNv96pWe1XGYv7qtfSkf1ymHvRiW2hr0Wn+ElyX6iDnOJpINv+krR4iI0Jankgxv4jAZaNj
c1scYf9xvHFE9S/G+uvcPZ3OKI6UqOK+edOinJdA0tJB5XocxZ9YkeyxruDvbYCbCv3bDlONILOl
hsp8mFITT7YihpbA4tU8B4b/N70AswGjT1cZ6T0DdcbUVf8Tcajy1cXKRXFRQycTL0YmzoTUETTd
MuJ0muQWTFU9XMBR+erGY64ryHheJFl82458EcZlTOmP7swTpNKtBWS0ER32xAvrHTv/9EQ052se
2OLwEFgQtbsH8/KQt8MipUyHDqO9U6ScTALh1v91xZLgm0GqqAzE5CX6fcVKrnuyo5ptmzFqD5tI
bQlshAxTnKHB1rLVXVyO14wYA4bw7yu4s6TYlOznCVbbLa2BhqBtI1CLsBba76KP/OOf1zaGu+kd
HnOcj4mnUJsO8O5VeM52AUB1+6pis3nOcG4ruCHAiuqsZoc+LU7bZC49UEVu1KxO9QQuZvlZv6Ki
kYGSsWj/DDV8a+lfe6713h30/GEvZcG2N9PDYkQtC2hxsRm5mSZZ9aGlbZQx4j4KUFwZpMU3Sivm
v5uA/buvwIo9DDm2//hksqJn2007fls5stZC8AXdtLjBXtMdZWE0sV/OkfG0fJMwBH+tUxwyH8Sa
i1Z0HDqtbGJBkg6G4tEJgpDABg5ldkOFSqctbdcTU3z3OIQpHw5h/LWSwoYf43viy9rT/hUkt62a
veRgoi7JDPSYQNlrna1vu042ecr4PqLamRKkOzD3FfXr7KVXXpPxpNEgKz9mAQWQtI+WBaOLukMI
GylmOdGzpOkwx8F4B5kQ+FVixoCNUuiCL3j//ItbvKORghYKqRwykylQQlhBOvsuJB6H9eUlB4ya
Ru+m2B4s+zolqEHww4cc7VWjCSUDRNULAQya4ly1R0I9OAiXvlC8ib3LpA3pckEH7AbVW+DwxMiQ
ZCCzwCfkTJNrldm1kEJVCIdhI2SMad7/oFNGpnj2HS3wAmy6gRqJeprz/5ekcXuiCMlbVVf2inzK
f03ZGHiynaSrzLAthAJ12AsXsEg7lgd4bUT/FOI0pHGXrJhkDfg7RwIEXt8mIhvwSh3psvabsXdH
BkJvpB5/G4jTY6E+7dqOPDqO6zP0b7HliDGhKXeVoaYTpxTgGH7o5i76j7jM7Cp6GOBi6y3kXz57
wVSfMAd1G8fggrxg8ESvYxw2MPgdw7KL9jk7JEhHdb/igyx8So6zVbBElkYS7PUWEGWBgBfOu4MC
qqYA26E34p1hYDRDpfKOrtlAco8xBDubbBq407p0vaJ06iPHsbLLvS7lmkdqU2Xpu0gx3VdcBVGP
ShhL9F2DWxhm75HLeCgoSEmj0mjQ2CTvfurvd4G8pe3Atx2UeH02bPOlruSqSLBv48kVsRx0sfLK
nbtp5ei76NvT/Ebz0FvpJweK1CDk3FpMX/xQcH6GpHlAjqbvZ1UEDF55q1SaP6FBFiDA7ioOG/BF
CupmPiakzq33f/MRFefxvacvuiDFxSUEjPW2CCMUKNWtmXPzhcdagffbTJg2yMDqDOUYNPUOklUf
lSa4ze8NSqqasae/8l1Mx3VKT6sPaZEePGmcJ4orpA+wne3B6iE27T3gM1EPpno/v2O07D2ABDLy
u4dY0/rXpE3cAqrUy/RYdV/cCjYo2KrFuK7qpfaKaXTAwKNvBAOb6u5bCFZjYbivvTDeo/+Vbja1
Rrr4D27wjQwiXTTG4mJHlDqCXfkCki+E3niQ7gezkws4o4DRWh1LiugUOlG+9vYPZdgEMzKBjDFt
a6rDjxhLdsfvN2unW+FF14z/HUhGnZIUHRo0Lym+4pWhDI/LfORj4vFJKEa2eY21GcEfOxpxOJtA
fPLlBNNeztNINecJumRi7hzoNp+eGe4MiQe45qhSSlysZriQ9BglOnJLEPEHLpyxLs+B/9E75zRu
7N8T2aheGfD9kLv5/wuT3PatuQo8qkEyuu+BGe1H3nBLaiAAciS1HV4Ti3112XTmcssx8B+T0MJP
hMuCjoaH5gWINVN1u+FOObcTnzpGMSfbghC9ZMPzZssHsq5UWLzEKa176zbncj3h8EeNUTDflxAI
lnI8DP9qt3nHUB0kEeFK09V/Ixk+A7/P1s2SPc2yY8e8dLrx5J/QKyJu+1tNpuxP4/UZpYRmMMOx
j1QLEU4N8JtrcsJTlAL2bbRtUSd9EzdtHBX0SuWyKSSbwZxEpxdYLhOw937eZ9VaHcygbshhMYd/
vr41dT3W/C+H+/Fd49m6rObpENE+z0R9h2+kTRmZ7eXM6jwxoteIyFUaDXNkhWMWDjoo5J/cS8yE
v4q3hAAjzA57YiTgf+R1yIsAyJAd3+n2U6z476T4w2kWYIsm5oREdJWRsa3nZi7HUQzf6Wod1DWn
D4ru6g1hyWJYAWsQRC1CvEFdLJGQ6Hti4gUSuVTwspzCbZVOT9Tm3BcJCyg+/uIfgL3ImVHlangr
3U8orV7ySuRo8bP210Ye5ojhqTDYgxiW/w5M5XWvNyOruudqL7kPtjj6sbn1/Nel440RixX4AVH0
q/jGByARjpygNK3nXrPuNM4W659t8QOZBVBHEg782bTWrbnfIHC0WDq8VjOU0LXd+I9PWhEA1XIC
+dPQhiGu5MwY/V93qA4Ipup4WWuxvCjWScotoSuL9JS8qYOh/mV3WQafXfUWL1JkL4Pz3VmlkueJ
9Lw392sMTvp9KgkpsFNdNp95CUeMoVWqyWVJHOXdxa/koT6USyLMdrWf2JA0m9WHJW9Go5dNhiJz
YAUqH3qsCS5bMlaGgE5tNMJ9AE4Ck5wPyzTwdJ4EcowZzk/jSFrAnFDmd9sHUvW7ZWiFKNSDNapa
rWPBW9LLFh/6EJ0BaS9cqtONGVvKTuxuiHm+S4GBhcoFnlkWH7TlkhaUntc4DQUG2/UCNwwwuLOY
HGsHTOwnl8+jJw92tBcpReDI5KmCeehqmMRj3h7XuxoTQTfCv5y+ix8BGlnq5bgA4gDRWvgLkxQ+
iH99eD7Qdrd6c7UsX4GLa3176dXkxwMhdtYsxkV+zaDtw22yyiTwiSqb2ew+2agxOyf3ylAx4aiA
wOe51MTaQAF6ntgRMfgTlIGvFMnlZkeuYGFyo6VsOPmjYWGqm1X00cuVz9m7peRWUSgLI8zYf6tx
BLP1VhOQl6koR1xfv5sbu/q3fnjKTXScgsEACYmvwFe0p6KK2ACcxKoHiQLEeUc0jnUB1r2MT5zP
0PVax3IKg2uAvbWI0Riuzvtx4QfbbgzyCDrbc4nXMKf5lQyUsckp6MWDJo5ke9BwB/HDtoHFzXlH
xlMfoEPwiItZNwdB3n0w6bQiuCxGwUMpOvRpTH7yyEmsUjBClL4QuGDEYlMQifoyP+W2MSX4dwVP
Ngf+vDf0/4vmXl6jOrj6DH7+qAwLfGLM8rKFJuB7xYNzCx0Y2CUz+ODQjzPgL8EQ6H1cMKLrUQ/b
blXnOFma0uOSgjiIff3jv/z4WKw19mnV78RaZrN3C1883/uhDcAqhLRL9gteX7GkGXx2ZWDLFhUM
J7LIy7CjS/Qv3HMRkqrsKMbUklw+FUfpNudnP4tSmyzersHQT8v6bkRwrfiDlmLGaZ8OBsFpZmn6
SegkU3D7o5/PIepHXZkdFaXW5ceyZ/XK10Ea2/OxtnGU43/G80K/UNIpYOcbRVdAqwFTqXiCWdG6
OXAdr+dTmKi6dLvYya0oNR06GhiHelX7nem2+3VDIWgD15XuBlIFNqy9u3FWu4gzbrVlHOTIfwIZ
HJ8m7APLd8GHC1NmlgLutMTf4RFq1of8uy4IL772WXAWIG8ulg4zRKSo2i25prg8hl5ZT0ifQXUj
KJjOT+WP1ATA6ZTRxg10ykkV5A2Bnn7nxcS9C3xARgUbwNmnmsz313fFhYtPGYKk1GCDa1WCxHS6
osfAMom+h+LT3JFsX6MdkzeYveSwdD8kIHfISWz5AzfV7H1mmSg629EooC92o4DVyjRtNxQZwhTM
kGmPyDh2xbOIM/Qee7xSkBgPR7lAaWe2RXD30Rn1LuG9/TTCSzk+fFhEz5ifOAXIcORKuiOAghW7
LJtZiMBJaxn3ramxEzDoI3MDoa9y6BhqdmyDXeiLiPyJaWrr2qqgS/o3lTlIM5qIBCAPwEjnt2jU
GypZLgCOJMNq8LPJuQdqkayadm9zzBrU/lqvKW2drYEYhXoyaKgjYImbQbuOYWeHuMgV9KCaXdB8
liZEaZMNglTnSFjL/CDt3BKvH5ZmcPCmihIvFC4JDoPnnnV8jdtJkxrpmQp7BstTkxEg9S/kINHe
QegIxtPkOpzK/M6gA2hNK6N8P+AMwiF/eIsYwUr95H5bu5UIsSLxQfCIzQMCepxXsLbpslabvEd6
e9JBaBX4etHBgwYd+YZQzpea1W1+kfDnozjhAi3L0MHTR+acAua/tqmE91JEtMCKatYKPA/xHuyW
gAEjd2d8KG7UpdrEcYZIFwtFfSmGQjG1aqUW/Z1Klje075hmdQ6PA0kgr1Ju8Bl/moK4KhIvWHeJ
tzliR/wHY2Qvglv53fJVJdfYPIkHfQOqou+E416SuobSI7jUSvYfk14HfXXlQMkRXcOI1zwN1FWS
w5x3G8gyCAOw9PoD0Oxy4IVgCBVGMK34OyhJpJ3jjFB0ugTG95+5f+1OWlBRDRIHya3GsYoRNqdh
DQe8hhrhj9nOAB6CHdDMlFFDesLyMOoAxhUWW/j1V/ZUkd42vOgZTdZ78UF6/qxchmCYPhjYNSUn
AIJUPqQhRPgHU2XML2xdbxFEjHraYXcX49IWKd1IhvOE/L2AjpgfDfRyAcSDPxDZcZ9L5LIH/uTs
C48ilgUoahQXTL8XApoQNIrPZfYcHAqkhJvS/G2LnuuXdQXGFdTZMl/tcykFGgQVXI6cYBIh0sH4
MG71vgq+fepSpvbUPjuG8TS8rY57qSEedlvnBT+gSUsEhFq9BJRdxbCErRuYawGoqy8UhVCZRXQV
jLuiS1J9fPnZC5rNA862tJi+WJbRla8H0hB7vQUNgh6uEs4YjMByGSIQ55XlBjfN+7ZMsXmk+CfZ
fd7FtcttIyK3Sf34eFRJ6jGVtOs9+HoXtkw4RV6TfK2lUAyiIwz0ZsctKftYgyNe0y9j3rv6Tx9c
LBMLl6M3EFExPLmgF6kELlWRZVYx19fA7nLxmC4jHA6XGMthihE+AVH8J2Fi0uy7F1wMA94VcGAo
WkpjHa60XM9hT27OBDkshi0ridJSxofDZyV9haCFtBOnfGOY58/BcjhiXFJiXal7fojsKntjeOE3
Ot4RNDpORyRTOw8fBKq+BboLl4NIfiR80QvezCE8oPr3EHiU/ZVwyD/lbDycwvBm+Bwy4HdpocWw
cJPrF/1yJfnNybPsBRws+ZEMdP/gErkECucgghp9+K4Lna6sKiKXe6HgHCjAQabYImq24D8Cch5S
jXt7kya3NHTspYmSIcMuPxCnLo1VkIUANmqGMJrRRX6biu5XmMAaKmOQphiAYtU4TJrCf48+Wowc
jeBY2xQrOjSiwaf9eK/8RucOj+MbaXkiP49JcoWCByAx6XCGRed1Fh7wTe5ZP2aM612VdS4b1irw
ow19S5mYCLkSUokFx3qdc2CYxle9NKoGxG6HbUSATAvqAi9hsH4x3MZFbWM8xXQqlsaZ67m8cgR7
I0UjdCAfrkWyBGLSABLNAbcd9YFwbHh+graryJuxSoHgRlRpY7x6N98WG+eP7H/7LHeTBgxHe+jY
smH9elJTZuP69/a+cpuLJEjEmVS/ys9ZqzJQO5ExRu09LPaYqeHro89op9KAFh1zFZe8Twmt36PM
wA1C/uJ2m9XVtLghwnca1PaOlMSD1b1wNfrSx+dc4Z4Lv858xyAnTa+zsmpJ65UeqM7/sEYYugDC
uyO4yvhtxbP8bbYwKXRrzF4xqxAsX+E/yCokiDYVWGDA2RUaXxLyFxXiYWdqCwjleDC4wI/Y+2Rz
/Mn0cKXai/6iIa7YU4IrvfIUKPkseBmAM+5qEAE/WBbVvGTJwG2qVaQ7NxQZI9ZbokLHezKsYhPL
Z4yi/ArNjMiwOnnQ7ecvz+qr4L4q5nrCaVYy6Vq6RgYaPYRXpnfGB/ymmck2V9SPnFnry5RFE57w
SuOwrxgkbIRJoqPlj+lETW+GHzj2qtX90GbtE9sYwm6cdMaU45B2mQNnATMo7uu/WJyY72bDaM8o
0e4YeWwSZgq+UMXqE5mKlcTyuW13389fR2qDQzG82Y5+uc92ddP99fYbyCFrx8tDUysgeWhNlqA4
MyEIOI//n3WurwU3+omOSaLG8tPWpYzIHyrKYa05htsTOVO1JLQdbucDrSiwyRqvWbKkwSD9w32Y
F9UIm0KuOpfg4fC7oA2OlXxdWtjd1awFWIVV1BgUnYCefEo2Mlx2VI8y06YH/OQkX8IuSD5kyJ6r
ORXmWHIRVmsj1NSK7lAVykpjWpW8CNXpVlXIt0Gv5Dokin5inEckuZOIl5VfJ68XctmyIgRMGHXf
JyvBnKtoFemG5rhQWtWxhfEjV8fWGbFJfJ9CswErEbp2MUhteUvVlFTXChR+M3p24J67i+fqt3O8
LMinZG8Qi5sCaF6dMd8F7sthoXNPGgfhnhJszCCZWJmvV2KjcnMPT8kccygBrfa3bX/WHLUVslmi
+KI4Wi1Nmf9LNFCYVPf6rk+dYQ3xcgtkCVxskhrIyCazToTXT1TOqtEHSuIeHd527Wlz2iBxQ8p1
KfZyyqsGYOfL5LnWRaNdT1Jx2Ui1IOKSa7ArVKNdc1yaO9/+mA4hpin8yjd5KV+boNodHB1UPTJ/
ErmlCK539mxCSbdQPUvjE4QbuWZL9hT76jkmW7/mD1520y0g5VJ3AcLIHAICE7HjcjumSQaLjWmz
vEW5/Hn6qTH038Vfch/tervD+tA6YGd4W8ADNiXSnlU3wHrBlE/X01+6RIF7Gj6QOA7lAl+naNgm
xuJ/Oq9mywH52a5pfD0pFiYYBGrPsNVx8Fd5N6JgKjbgkvnFn6ICkELERNR0MQ5i1XimdgkySeGI
9hgRBv59YTdD+OL13eIubZca6nnixYkO71sB2sPtGaKe3vCBGU9NBg8vPEu+KD8eps053XXQynUj
+wv5mXCL6xw5RvV0SYqvLbYqbSJtZHGCl5/KUxETdQUjA1Q/a2oxla5wpNmJ0rFqxyXpU6R/65O3
y+N4ByffCHUFRIr9c5EwtSRArizLUHNXJEs+kd0B9nu8dZQVSJ/iso97wuUrR3EJjkoBWBkjHMt9
OqfoZSwkwZDsPQgzHBeKqdSL5IAkm9gAgxy+ELjdeEPoC03lTorcQ0lWkNKsogq5mqrrUHZ8moBM
3j9QE6CrZMs54AwLT1mH7h0B8vR5fpVmjuDT8uZ94U02E/kmQJikiEHmNzoJGObKimUDtUA1wiuy
YdMPDa56sXoqlHWtrZ0e89Auig4MeEJ/aMmQ3O7oMQ/kyccf7j3pEGfsZeIxmYeayDQ3RTKRj/9C
ZvbUmDPBQIUx+nSb9ulUAbktfI270mAM56SrLP770k015Pa06YWCEv1PBD5T799wOKnFenH691jL
Bksk/t21utjSmU1WgmPO33DQDBN5CKD7nlQ+FMNYW0g0hGRVXL8PPyqMy5fkWRb7Skl0L5b7LlSI
LMoQRPhHhcSvUw/uqCa9IWp0/6kC3FVgPkXZJsQl39Mg4UKHOAlW8ms43+w//aaLZ1ZFZ+yNOx2t
vZLrMUpvFvwrhU7VtZwJDHfM/uP+/qukv6QQvFGTa7mcBcSVsewENd9nT/ArB+Vo3UANWvlj3fIl
lgn27oO3p6xR37LCKdB18mZuOaojX+PQ04+WkQDAX5HJXcj5ZL8yYxOn/XRO3qgYWRe6aewjAs43
8amuxvtT7qiFcud9sO3hB1p+w73tVhysEg/lkJWrAy4LrwDdvTE0jDBdM+VHC4faGEduwWagwXsu
y42VFfu/JAQOWbkVzjNfaksuS9sfNqOU6MX6lcbeGA1xUr1HXylkH/+Jy217X2SVslaBbiL0qcKt
BwCe9AF+EQU53OEdjzR97oBtDVplmucXSa7BudtNh7IZnG7mPMVEk9lEUfCcdpQKxgZA+JzfY3lR
1OF/Lu26OL9PKumAABAuEYIwYPm5oJd0yqa95iYGp+F7I4lTPJl+mtm3ps62VlRw88zXhLh0l0LO
Pu2ErUsZAgq2GMMBJT2txgrM1tQwJWrBW41iaoRFtxzFBHnst91EZw8vJabDhSqzDmf8yQtQtv58
H8Y51fu80ibkIEiVqEJCLe8t+6Lsc/HcFn7WGHjZmaOSPxjnYcb4vwa7i8esjtUiELalyZh5uZpM
q3L+WNERH+sSuc4AUlUJNy23B49aCsbxp2TZ3moYNqtBLiPmg1CLBNm1d0ac5BzfuO2O+lcugzmQ
kpIKne7Wn6wOUGmLrgZHIDXug/BUcq38uj2HXVfHm1cDZVAleYV/g7DDXiZAvd9vQmb/fPiabdhc
+Hb1o+J5W9kX4KyJeOsvjEv06KoGTLqOIvRJOLJoj17VjHwWsCWEHH0WAYqAdj8DjFbbfi6AMp1P
1AfqPmWUgyCXROuCCrzY4iRFbeYS7JNGKP7D9jV3OSlAn8p0LVV69q7/IuTUOkTSZ7LPucei2Rel
OIK2/M4Dxz8M051cLmfvUu19hdg66yndJNxChVxvafuw/WqOowHfoifaK1vufSILj6CKko589QH3
N+8bzMvuh20VjsoCD1bwEFXamNww967KEpoOy6TgTXDs5I5ZMliw/OlWCk0N2aRh+x07PGlXUyNo
9ob8Eh0/n3bRrggYXX1jzXf2IoSmhchAjrbONUaRJcHwaAC8pIpu/1gzdr72Gg5QCoygZOVjMsD/
hsdllUAyLTqlx0t5dz1dPp9d/m33nq2UQTBEmmC9p97sqc1Ebqb15RNZNP18e9E8flcydxH6M/WY
nYxms6OjMWr+BPkQYSBtcy2YrHDse1EV4EmrUyLqdc0akTZ7hYZu+tv2U283cP/gZWavQ8tc8Ks3
T/V+1/diYFhHnaoA0PZSTQ4RTw1gOZ8PssDQMl63dHYZFCMoP3iSjXnNVBjbeuErmIIj48xMs5H/
MtR4YhNBWCspCcG2CnWOTgRNtaC9fLc0aZkcLc/P1K08QYS7Ua5bxnKR7FPZ19eoWINHNJFVpTsT
7r3zIQn5z7lI553TWsKyElq6JYzsjK/7oOmGWRDIEzH6brd8RVykdyvwwTWBmhvq9/TarPJrfEb9
3stSHK4eTtk3ggUQouo/KTqKmT0VNPZYctKa6n2C+qOEwa/CgUZcXNWzO29IrvCeLbhbiIkYkDYA
rBYgcSy+kxqbOxVm1LWUxTGXdlGKe1gKXcRSRufPibLULoPIGpREA1t1kpYOC4VbkXQ8gioydGkP
sKdvd+9gkJvEK4ZGQQYoNZ/kACBQ7vgRMgMr6B2471WdZlzwt7h21g1/HtNWN7V9sj/iiQhlbUYk
Se8b1ezE+JJyRd38wHjsUudr7UsNf8u5XTPhp42xufHrrSXkdNFWa9ipzc5hEnhKzjqkf4oQ0SXn
xZmeAfthSR6KgvLdDoruhsEeiOOxAEYHXrUqFkKagUoZzg8/xm4q7yv/V8Y1vu0InTDm8CJZbuEO
Z3sqpjcGaSWzr1hgZZ0xfv+LcTz9vhOx0wLYF8jWzRK2sqR6SzOrVYIpjqGrHUARcqSndQac6yyU
0zzQ+eGfq1/Q377yVoeuNbVWS96w71BGlmVk7APQulASndme3Q9Om+8myXj+PyScNZ7iXo8MEZvY
xbSoLDve0/DWPIop1leldN4NIq70Hy2en6SRg2dMczGV7GJl6jD6A7dTMlEtDTBhuSsok8ZIAJG7
lheEqksKZ/7YagdhlOKVU3qHJm1m3hA4y+Ju+NMziASV6W7qtJr9AZQ7FFk+OahVEhEYhky6THtE
szMM8s4ATbpocn4OMSAUrarUmMFSV+XDJXAvJ5pMKHGiTHAv7vKKle0yw/XH1S6yPthp863S6ZSL
3esNvsnsgX0aKJSlREN9TpyHwKRcq7j/65NURSh4MNbP28mn/a4EEgKWtmt6GVFsDFZuSDHo12dX
FNf8p39KLPeH9MZ0IX7//ljKmxll2+VePl8Bw4DwY0tkMMre94WRNSCgKF5/46+ozqOUOMG8+WTI
4iJi82J2wiypCX2AAiiWeMn1s6P9dn7v4RUJ76ToEJIIFTo7BbzSjhy5I+H1cscgD6WOTvAUafpY
ouxaUfQ7nL2Ii7qOMv2LVLcE0AWwblFPc0gZsCB9hTmnGbbepcFFmEBPpGxNyTdHimX/ICrKmoru
OJE7NvvCJgmm7kik1rhQlM92peBGIukuIxAAkdwVSBerHBr3D2npxXlu0/PX0dunDEZOZsDO+8IN
jk2TmqpWjWWwABiHigOndcuiSbbmh/4AKOauf7rPpRVsRV40Az8tWBsjFR7ZSQrd+ruU33YQoTyz
atblNwa/asG3UzK5ocRwqEZkGPkl9QhWvCg310Q4Ibyb4vYpL3muqWjSWncnDM8qcrcnG00ZHCAf
xIoYM497QHXWbE6ZFcUPhjD+WmRC1NvxD3fZuv8Wgc69fsZHTJiR89LaGJzP1/0gPTOXdoXmhaBo
zG3O4fQjdnmYmwfToz2yAKg3PZFl1ToLMlCk1sW2afNOWI+M4KpJqrTMofOe+ROCm/G4m5nkhW2k
zbR3Uo0n2ByiDsufly6p/UdOsdemsDrHkrIh60ijZK8PdK/xKUT5cdoLeS0W0UvedLWov0/WGrwV
Pn+reITTmpDCRS17uAHrmz8zA2z3qVZMVDLa9W190OUjNP9ue6IYDuO8wz+H1PtIJrVfuiKNE2x2
3LAbOzsbhVOtZTQV5J10ZWhF3jdBuaOOAyCOtke2pSFm/XhkaM0d52J7DAPIrmAQ/NKtU8VGIc4P
ePQ3jejnPmsti4/lRNwQB1UYHGu9FldT9zmwAAoScCtNH4DOUh7a7Mo4ga4aN8WnS6pdwNNGtOo/
LPRvXdgn7XJd2+1K0VZuUE/+5n3zg/+FpPdDIaKJ2xlOZJf2dbJ6LEM9sZLiQlQgSYn1sN1Yl8+s
q2EFG5mRkyYJ5MpKCFqgfRodk7+9c0AscwA3QpJ/S1uJbLYSXq6hMb6BL6vtsArHTfLQnDINYUFA
9i+Kt2KUobudthZl6nh2huApp8lptNsZqE42Tty3toyiDwRoGTPaI9ACQi0Rs9KBatlAtCZIfVZ/
5Bmj6c73kNogJP2cI4PMHUav2DuYH0UtXQ9fDKIT6hqY6fHlrDZ9qdnjDILdjf8NIPXDwb86VcjY
uIcqs/dQBgkXRzlzRjK7ckmgZFJ3Qcola0tQiq0mvMxnE+yh//rzuAU0yYLZw9u0uuXGv1jyZmyt
ZDV6B+SBXq4WYje6CmzL2PUKhQF+uDBek8IOPLTEfgl8S5jnJjmBHn1jOaWxsZZ7dDALM/gEZI1J
svc4MNMRTtRWh9bhgN79POsX/iUaRhjoQieKwvtUPRCVGcu0c9yEg3SmGspRKtRLssbAUjaXt1ki
LbVZGBFyF18V2bOSvm9r43AgQAFlNCT51RT/jPfrui6FUXdAlyQImX3JgAwl9tcAetSXGcLyaOqI
R4oFCbcZ7QyEnhjJTXXTK0hsVcDDx6xbSiHsMxVkkEPAhfnyS87FjiVZH2kLTGKtdVxiE7/CCOnp
AxOaiKl8/tID/PVWiAWAIVY8CUqObsu4auyZbd56xfem5RTWf5PCDZPA0zNVydFWWIM84Eg/aF39
Vy7D5oQlsI2rSspC6XUAEw4JP+c3zn2iSctap0cuLCcEVW1/w0eu22zRuOl92ImUrHtXuBlc6BX0
p56CHA3LYGmnBpkCpT8ZRl/K55kFK5EfREdFjvTgeAnSduDx6+Q1xzby9bXZyPzIm6Z29axXEpdS
RFj64BtIIf1ZiHAaJ6j6R8JmO5m5a4evgECJHAH33ncQuIKEw6gxCcWr6XPafTSaXLKi3sHa7b2y
+5UiFfqpjdvjuq6vgmQpFx4a7mJXrVf9ymTMXz3EIwp5LK1ToH/nb4Z0cMVvzCrYJAcUB8TPymTy
H0WNAHYVg6TBOC2+3m0QNXeSuYnt/A44nG1EJRmQuD4NT61KsUbEXqkRJbAsvDvSuGJxFOg+kXK8
/mZ+LNRUgiXfbEx8fCrCsBwz2PvUJbK+6YFOr7vfFJRuD3KMQSD1Sj+FxoaIjSKYYHr9BnhXRS7Y
totRw5+2rOzbXhfLQkDi7JxbXUEycuuEB6dPAxKy8iEx+ESYHxx3Uj7wh85Wldl2aPUQeB/PKTBg
azYlxkekWZaesdG8WR74/tqczyFxGD4dVprhFJXv8b7nuNNvGaGswYLnz4sYkFFnUfIBUDZ5OgsT
xaA9lyLkhAgukrMgxRPUhhFuDtsrjvvvxBoZo/T7/0ReitnAKwK/qyic8G0auuiLAcc+5NzM6PBp
anva21/K4mK3UHsJMZbdsBYdDuMBFet6DN/3lQQYlY8DBlv9mwcO+xNHxrPejISEwIbhZ9YYf1oZ
4KI5bSArfatmARvR761+TYPrtA6EhgQR/8ClHRlO9VmIdnv7wFxWCBB6syNqJyP6Sw0/Ywgz027K
85A6j6V8F9rTw3xZ78AB5H6fU/Bx+kTv5dfy1wbt8QUU9DNYlp7qFMj3oFaNs9sfMraismWmDyKe
RfQyHC9OY1PoSfLR0RXvCn8/VuElfPI0fjbah2fulTYfj8wswV4cd0Cd/EtwUR2nXuVqeejl7/Os
7/tJ3+iF+NEQJQEm51JirS3pe0Hskhlcwf17h3TAUtcpn+GMkD56rn8KeFTonSc8t1rTb8CvhTZB
cSZyPX08J7zpG1G0T8R64nkobaxa+urCW/XTThoFt7DqZqF6p7YtdlGvtYdNi8+1fK3KTBMV5eI/
I9BbfCmSMNH5kwpg7EM3jnRzx6UvTqhe48m93vJUzn9WUmU0+63Bla4+A+mMiUfrjqPbKwyx0gUL
b3LX99F29YY8FJs80QFOey71uTFkyIG+wGTq8q91JaRC6vNldmDrfVwkmAqwqxja6Xt/NbcE+RHO
cEDf6Omtjpcfeb94bja0iyLCzrRoXPXOOApCWdghFyq1XwaOkHMMtmuniSPMtioVcEco6ffNPhPd
a6F+pLtziX3nqU9l8mQc20Pb1YtRUSXSE4S5UkEN8FFqstuc66tYF4+kb4G+VavXTm5eMYOfMf4y
AYfrTUIck32byXQLcp57quFOZtL3a/c9NlT/yXZaThztzz4Zx5S9Gmr2NagxY3xdCrrUVoRmEvbv
8s8XIVvcZsR8CIIT6nhaJreE1uhFLSZeN4bXwUkY9S72sE5pskIqmOf+n4T6pdJ7u/ii4g08Dwzr
24g4zPrjSjLS/A1VU0uJeS8tLIdSEVLsltJoTbfd/ksVrO7ADDZCbQvzY19pjteIGIPkGhMYgjdj
c5mytYNIRSAp5R47nV4K79LeWKBT9AS7IgZK66mNx4+lmc5QFElWJZcdYuB+TMV/0RLIXgB5bY4W
vK/GDQJNtaMmXHgArNlMJ3ya0Zd+FRp7RKVxAIHnl68wr4P4gXIhsHgh26SNlM1iPcsTSwj4gipf
tvh08oLt50wxnXtorTKfPgRbLVuOAig2+JLi5Pi9N+T3cIuHy8JixfresOmdcv9IAizOdSyjUyaw
D8EOJlzOSlIfIkBg9GPaKhV6FKG9FpfjpkWSTY143buW3nSbIMdberAl7uAGStWQ2nPd7tTt0LL+
dTJjoK5IiqkVR2i/Yl2v/YWUy7ceKH9Weuc2bMKH6Urz4bR9KveMr8eU4O11cY9dbOn2TVzDtmjo
WIl/9q4d7TQXpaObW4i8hgW5UOnGZFKUta+bIOOmD+JHfvFL0g9ihMj92cBtpDgvWDkJTzRNjN2a
LPKSc+lrQ7eP0YHaM9L9RhE4v1urf0qSi9aAQRQO9qAj/Z5ccJwKzOb+26959nRyxRADrFVexLhL
T6lXLcRZ3KZoeHagWn0xBdX2c7tuDccLemK2Pc/zYeTvoZ4nWdlmXEQSITIdtFrTD2EQ/I8LbAuE
kbq/hEjf+bPnmr5SGRD8LSkUl303SBIHwRkuZRuStQgEm8/oZRUZprM4vrIOHHu/uab7T5DwxEdo
MX2g0IUZq5AIwg0nYzhLIbo5Q4BdeW8e8k3z02QlBqre/GYslhP7EN6IUOvYQn7hrv31uHMDfoW5
yf2iIt0UkQNCzP1F+s7xBqxOi/vQRMqqAlevcyzao9JCRVws5V32Nu4rB2z9m1YgmTMz6VK0hBBH
qyL8mVFVNrg+TfhYjv4Dce4x0IJgb9b1YGuQryfZMatUm7DVGoUGqimHlwYRjcSohS7I4bMUwqWu
1hnMeWUV+Jv27FXzQEWRMhs9prwRGNXGuRo5qtIluEdfFxmkywc/8+oLXgryUjdU9poc6izxlNp6
zgl0mx0s7QUTGeWcm0dITufuTR5G/LeRSYfbCSZq5JxeFoxFF4CNhl4dQA0dCI3cNNlQZnjVprWF
glj1LzWrPhkQli7kmmabEn9msMgQSHNNG/F4Jp4j+w5EFwKqF7Ky0gdlnE1r6Oa8pTqsp6mgDiZa
UWRs10ia7mEE7dC4mzuqrDxIpPy2VJySqSCd3TZ9y2BxGvOFpeKsv4qm8QnkVV4ysnkhMxMEMWd3
f1v72X6qwjQmr2o0mX11/jsmouk5YgCENkn+iFW/nM1nuXp7h4JKk3WQgjgNV/VTX3ysEEJCOkL/
jSfuY74seWiwbPpXbBatsNAKpFPrhz9nQHnn2UMMMn/hv+HnZYke2vTg1fkPmb9ro4Lc+AiZ3nEq
jxaIOpOt3W5f/dvqst+EqlvnY56hKooRcSPDVIBScUg1dyfCMit80novdomYVw6IpCXnjewobcxN
6C+yruK3BR7CiBhkAJV1m9IkfPlg8ZAQO1hxw4JsvXtM7tQ+PnmDGkssIeUvmJF4EDERPdWj00hJ
45tuT74fcls9vTAhZh9ZnAKCy2L4NspO0oB21VFyFOKRQiHBGGnCaRKkT/o43FJoFZ9MV4+R2KwB
5VG+Qiw/igL3WctJFVfrn47jvtTGCkKvvWRFZORbOkmTPUebh7tl8PJxZRG6od3LIDiWswdmkpgY
Lu1u+GeavqffvcUqN+dgMO0Qcr1r6SHyIgi2IJw9gC3G8wlGBI4nNXSHDixiZa59Ps3mNQsKD8iv
SFPvq1ZTAbHoTRsGeSQNis+pRh40IUAsgSUFKohzSkgME1BUvEXiPZBHS5nOdux5jZP0aPjr1JZt
hPsSapKkWgbAnJMvb1Km65IJlCJ4h+aDyNKL7FLluwj2Rix6ghCGiK0MzE7/t2ZrCDYDLC8lCbZ1
qk5QwF9Xzkdsfu8u2nKVJGxUk2kXwim7DV/8Rb/gthja4bCwMx2Zxh30iUF+yZX9t4dff7cGmV5C
6o5KU3pdioOh1o+Kws0/f8RWrn/2XlF903edpoK8VdK9ASJgiKpjeaq54nfsnN9FwIjrVz11309w
VVwS0xRl7Wl+zmEn+0ZsCrhpdnZLuD/J9Sbz2PJpPtT+zKpbAF3/dGIe0e9ZxsgNBkfzba+y9NqF
zFVyKGIQW7BjA0SeHeYQHbqH0cobo0qUFGYdCesY/ecpVK6rXczQV9Y7jDJ9kdSSMo03ieus4NyH
+PNSHw4Vd6ntAPe4NNZv4Zg5G8nlgpJvlfqhl0ToKrBFqxqC2SDlcWu9rRFXrK6Yl9fKUpKTwjv1
1HNqqH102yxc8bhQci86+gxufDW00fdsTzwShbrVg1j9sqS8ArNi+0X0+psU3DPNj1dLdbmHwuSm
MWdO2cEpADlZ+A0eDVBBsaYhlFel0zyNsVaGkv+PRgH3rlKRLQWXe8k7R/EqSvtdCVuJJmjhZXHE
mWAkQ80bHwpEgiFm1tFXYD1tSXC0gsbyE8ogm8stpGTi1U0isvx4ZNU8MoiIpt2J69dq+Trp1p4R
qfe2b7pRchm3j80h+FOAmM6MQlwLNbMIw1Nld6xFTo+mKFhxhhauLo6qAfAYlMV0lKflXaAFdbS6
y9U8992813tXLyO3P3p6YsM+0A0ryUoh2f+7y8JKkvCRpoksbyAXTTzUs8gjZbp61BmYftJZqFCX
arOiJta2u7XAGoZdgq2RWz80mNvAhKhu27fSgwz/IAYY0mLZ3f8EqsDyRDcXP928AJF1+jj2qJcN
kV2t9+OlesZaj46yhSNGbTo+x5CfO7GDM/CX5UTbDzvJg+RloUveSo9O8axVE9sq32EDlb+p1HzA
q5agaZ2BpTfrZJzoqL9thrGwW5YybJlSEHyONwU8zpKrC9c9QmfbhVpL04U+npzaWMs7C+yx9Lhq
odqe6YircAIGWjgKQyBvJBHwoMl5zsacpwZgiBlenBLD978X+kNJZcx76J6KtLGhDDmDYq8bD8Lm
KevS45JTVzkk3dFW7KiJpOg7BYulNaZJgRBGQj40UY9RFcQx0ufgYmGtt9k5dQPXDi94VlXK8OKG
VSXQZID8IwaS4qDLbud7Sm0O32KeVnVjd9qBp4RBuxzGbn5bQ6KPY7o6V5Y8qrwlyWZGvIItgSUH
1E4NN27MUCAqPAqmdpfxMslfIiGeW9GTfNqghPMkRpSxzuisGQPR+XIXbqVa0gkk4h4ANtUzpyE8
2ILubf4qVjNZgLBrQEhGLhExCXQcSVkxseRDVY6mMmj43ufqYgHGFAxDDwXtA2jmIVCkhrUYUpdU
7lo34XxQObLq2lqL1LSYekNyJG5RT0kBVTFogCK8jj19CiTQ/kBtZpREsmsyKKFRrF48Da0d+lA7
asBoqN9ObsMaDaeUGqAU+ploiK/9oakwPsIIh9o/5WwvPrggt2qqGcCD171UdHdKSyLaVM6rlMlE
0alXsbN/3blDZITHYPx0FOFtIn4ccX3uGgarSasgyYMtfCZr3wk8bjGFo027VRShteRvS9rd/3iJ
wBbUEFPRMO6XFFMyYXIpKDvYCZ8eGfHRgD36RhTGtP5ql3tpDnStSCYOtmWTh4oP2Wc3T0dEr2W8
gVCI/DeOiPDiVq4lW0BWxd+4o7RXdO8APHFBTElGCROIk1MXHJ7nupWM/rEPeVtZln5PKHH8aKQm
1B9PLl3E6vf2rd/RKyQEVVJCdwmwkVSsICroIwLqmSVRTK7OrlthMN7hcS6lEQwl/OZngHaBmltC
78kJX/sZ2QKh8RRpoyUmFtwDe7QU6ITrlZOi9ekFkFwegJZEnyK2YxAngl9s1iE+wPep+27BLEqT
JME7RCI1IffEbv9ND+CXX2Y68m1BuK6clgFc17sUDfdzHKbd89/d5IA99fzHDs+jWdYurwXCxmhB
T/faJy1gQnyksWumJycCHBzx3Tz+1aDsLD3BcMnj8ZU7bSQ4cFOSzifOAiVqqGacSTXgoKCIYwl5
6Ksl6BUrTK5EYK23ruSOU47lxlRdXdX4ls+pEfXz32COAhCiZPetG7+6kj9oNlfaiRKQysfGYu7b
3vFPGy/iO+LaaD4o4AH8ZwxEZpltXnh6BInqqqIjwSh2uxKWU6JwapX7nOirc3lNyqAVTS3tsNwd
BwrgjZL4690/Awzxw4MRtT+f5/vhf15W9liGSbV9ByRZKC9U59LnZ+htr4x/YFpxZ2U98iyz9SWE
xQFGT7KrCjFuRwWOQnRS3JnIE2qyJ+J63LcJQHabyfeuy/i7et0pTxXqJyoREe1DqXocCH8gmtce
z3QdSJ+LBHRrvlrp0qMfKZn2z6A3tGaHR1FXVIB77R3/HxydAH9kmki8yOV6hCp3s8DtNEZrgQxB
EoW9iFFlO2Yv7tcybSIBCDc7Wq0SMPWbHdRS7WfEjwhUSSAJgPEKgb1cxgxHONxXwzowealOo/oE
/LwKSYzlqlSdjnv1DlbAk4I5nS+9MgpwGfJualItj9UGyzNDQajo3SpDXi0aVS0NpaiIZkw2Wbah
/wEEoXLMzTctP4IuHfyEWeMH6kOSQob645JVx1hsv6xgl/aRo7Qn0zTdgkfwgX9Aw3QVSfZGDNuV
f2JX0wGfToRUzPkAaoswYyIkIcKkQOFewz6wFyNhT39IdzvfX5D8Ohw2HYoljUNP8w4FwsIw6AO6
JaAnJN7QpBtglbT2FT8+k+IaT+HTijaMIQRzORHVfZnffCC5ZAAlEUJdM/MLhyuGamTt0VFtEF9k
EM4UQKewfQAhJJiUONgiNua7tnvj2XIYuJpAgJFWI+JaGiZD09hx9gh0Hrms/sYxGXaSGiZOUsg+
o853FXQfbC64TaxZJIxNcQe38IYK7u8VuedN0MGp3wm6O/wEqebOyvkM42rlQa99xmhFxJqMnxWg
eNo/NzeNVYVXbJc5uye4tkwEyVK6lzZOMVJ/8faoiQmFRatLPdw3rC+7DdjZpj/ADFvXbpEHeRrU
R10vRlvZQsemTDQtnrM/rOh0ok9cAPcfQd2LFspuWgNc1AienRAFPb06Ex2D5RO9X6fR3GC0EkGW
wnvzImfLLiJAZyVxw+PKdFjsRv4uNHwkUUDo3wS7g795qUOPGRVCJqphy+QsHC2VoNjJ8sc+AnEu
4Eg0Rm5IZDcBDt50CTcAEBRjX9486KMnI6IUIKMNW5JeZqPLs7g927xmJ2qOO+eXsoGD7UbO8fga
8BSbMlhXNGTSCJl18otW5Xvg1KCF3kkJZVn9Yy6wL2P0XrKwtHwGQxk6/inJEvYppWTJeLUozw3r
qPqDxaIoq3PAeqFS8m6pkILWzYuI97g8CbeWhG2Mgtd7W34CS6PNIN5dhVJfFT6QKzT47XtBLQs/
dM5tGrq1JdSGkyqzH/mdY+oUyn0XW/KOn+jND2I5FTgSmG4AXvoms3tgjNMM0AW09H38g2jazM/4
oNSt8WtB/zRutEvVppm0UP6gLxFII8CahfK32W7I4/wLVT87zXuw346X2euqTulDFSOCmptaiJ9V
SMkhsRX0kXREnfMras6zCujy+X5vQFmIRi2rXgd2vtZlHgIyOEVBaIq0QqhIpUM584KblAtP4kL5
V50Rg+2CeqFrPDrXeJaHDllwIExp6e8Olz5KuRPpr2Vhe0jEQINoxeTMkcbgD0UD8ilHtmzl5Wwn
bqr4WAQ4GYN7LhBwVvVbCZ0hELNbmnS+4fqmVqu67Eh0MLRVhV5jH1SJZ6WyALgEFDOa5rgL41SX
4K94mBWAvapWsW5dI6lg3n0qEcWBJHp6syxLPZTpxBodw2XytCrei0X9fhokpCZvvBwZvBo/oNFL
fqJRJPwuyanZQHTA3XBPCIKHfoEHx0nkVby/B+IpK3efXy2UlZZnF4LYflE2nYDVKAEaL4r7a/Pj
bvEJPW7bvWcmm1hd5LjwIwtDAvQGtiroBmg0xIgBq2qY1G6qQ0GCjeBurRrAAqkepx9t5ZK4RJH5
hseb19rVCBCCvGwSp4xv7tIm9t5RAQ+7uC2eIj1vgz3cOWYEbl4usDUcW3CmK40XbVbBL4vluGv6
Nw95U0Ea83a8aicfLUwQnV+YqSg+C75oqQ/rPjt/xlEgwnFItYpz3HDpcJmF2xDCZFV+RrjjBlRL
mNu9HiBMqUYkQLvii1ljLtWQey0wS0dMIzNTx+MlV0qr+E3OkUdbFw5vgNEsZb7XvSkikoIqxlcv
exs9959+W3a/CVi90JxTjvLPvItpwV5v6dDMeE8NoSclRDdZ1bAGWNSo9czqpGAFarNbzDTPDXl4
QGO9k6fAXXRXw2fKnX339ARdZXjIl/qyYad4tk2B9k8P4cdALcRJCSrxfrdPrJSUeI7EpBN3SWaB
SAr6ltPe8iArDz12A9nR37ILxdwnUxjspetYmBa7FDgvkzEoDaDWi1NvXKBOokW+UuIlx5R2lTHr
oYjOW3PCcRpDn59lh7tF6JDBWgJOSnzUfk/MvHsm7s+BKYTY+1lklo2InNIjrJRI7ODcWf55ByXs
a6AQOQ7ZwEh5DOKm7qcdWRbKkiaRoez22bZqaCjvJB1p2ZUv3oWnHguDPoZfY8VbNuVYGfeYMFgx
a76XhPTz5nWalSKdasmhhT4a5d8/KWeDPRUSHYVLpAlopmutsW9OZ3luXKpVmK83BXpXIhzdci6M
0AHQTMi5b/MOqACPcJ6jX8/X+YdXnfCOwwxgQszOt5h0GeWtHkxds89f62+vq3AEmSNJ8zuCYSes
zemx6OYiQ8f0AEwMwlHL4+7ZItDbOp9tJqZbHPc1R4jDvK+mHcjWRE+ZRNokmafOk7U9VOKQyGZc
yOAD77CvIYwlOHMUw/SJM+CQHhsj7VOuUb3unQ+bYAPnWXx0hg9HWYne6mWvqQFcgwKYSuF3SRrh
LeBnQyvsX/MbK97NZkUsbllWPhbO/tSayZhFq9eIp0hS1hcpdTlLJd6ZDktUaqv632/M8umDtb8L
fG4FivPY3JNu3elSz3I7rzZhrUYmG47Hl6/dezfE7SEtVs3jYWIBQPCF9hlXvKokbqRyjXlLqj6U
+AWEh/QujFAvCNcVvY34x83X/GG3Mfv3xjXmB46KfDvww3KH/HIbU4M1fiAuXM2VkHcMY9g4L+oi
driZrcPKKtWsyibB0heaxqjF84Dx5UWiSNqiGsHtAjDFA7f2dS6c4Srm1fIgL/saqi+Ld6scLuii
kicOGG8jd6LwmWLG9cbxd4DjUvgutenVq7yEL9ppWKhfemHNh3MVTdcbp+f0Vn7h/4wOCC+BN8NP
PKkpqoSA/pZHkRGN/nP7Mk8KAjA9wHWVMxaTmnBoghZd5+of8g9JWDODT7mBct9jphiH/5cM3/oE
UmZ6uvUhy2HlP7nHugo7noGH4pWlYC1v+LYBMboTeTxvbcZmiYdW5v9hBwd7bY0YNdTtSZWzVgJ7
gTWhgmuIUYvP8tfBZFvQn14dc4LHEptDK7XoPNHBb2FVtFsnNLddkgYUrzxJoVDlSKigMzpOjXFv
T4cKxPm3Mnp869rqR1vwdQTAmnM2o/LR2az00LNvuAC7RVH7850IOEF6AkrykdpT+yjdhF3rmnc2
jEITt0p0DPYtiMKyQ2r23lKYWl41vY9w8uvdRsHmennopBYaKnFnBjmqinlJBL9igTjO1innqKHs
7hHSoaG4ahulyuDBo7TPD9p1TfDhOqJRkCNbMlieZAUS02TEOZIME9gfC4w9KrBFiL3FxRhT0K+Y
DpFLqLdhKe2jJD9NWlTI2CUNIKMuXyLntvdk7IBXy8LwcH9s+9JdHWpLhKv209+n78ZBAhu3E68B
WCrGvK8SgEkKvk9mnCItx9UHb1A5J8D2RQpQl5IzBcWdr3Sm89jabOJ9qBAszmEfaLsdaYhGGrIo
8pgoRD+GTE/h/KY6GHws8w+jaF++jYA1uQvQSQuI7EFddErjmzzUg49m85kPdusBY8Ss2HJTD6H8
j4hli6kgzBSM5gfBMsav4EIyDnJKzV1pK+xW8JuJzk/gSHdx0Duyu8kEHB4XmkHjD8sU1X4vu7qO
4cJeF7X0lK1cIRsvTF/lzupH42+VpfGfWw14igHoDCV3YDlFRAlAjZoXny0MuYcWfBgv/ziI8Rr5
3bxRJvpAcvgE5c8KUV9PRug0miDOHmelmEN2xd243EvlYVfZ6ejVpbZiWMcEv2lPK1XVYJ/pUpYz
Gk3K8Uz/AjHPXb03mkCL9doJdBvG5ROT8lva7AhC4Xt2RCvtQ8G5krMlkF+pNHbjpIfTm38uaQrV
dGd3H00wn6TAlxDYeREeRPsQVwZtOy1jwEK00JvTO4M8L9L3UXqpZNIk5i4cw+PqOEAhnRsigsxI
3/n5qoPfbChNl9XXj3fvrU5eRfl4Q7tt+BqYwUdaicFkXuw78mthaRMns/D6r2yTKw3b8NX3SQgE
Zt6Z5IC2ZmzvqmzWdwc93u1lBbiZy93hEuw1patM1iKk2zh19r7/03GAHknE2cxEpF8z5BKuOOki
bXuomFCsew/fy91Vm6MUGq/ycyieKkssP+/WHehxmA3oVE/BWGX46kPA7cZxnGEuNCzo+Zfu5Xpk
KuGEnfFUwqr6f+FtxvgbXCVxB+S8LzXhYsJha+0Mjgf2b86Dj2LunkIhsWImTTyGQPcgNGcHwW8O
tlBkx6km/whKV1LMRu71iTOBNUYI4+aOJQOak7y0cV1BTto5DXOqA60Km73UotwLI2jJIy4TzKom
KdSoJh/neU544PrUFiesvylAlOZJ57JbEOjDKlQw7eO64w7YgcCiAru7EBFvhRscABcO136TZpsw
nSkXt0iEZJh9szQlI+t5gqUmRO9aSUV7CXxYfoMCJI1zMDYqwnNpSaDghCCKIWBg1wc13zYKDUhY
ORxmMFhex9XHQqxnS+i3HkiTn+nac9fGinGwDRox+r1lX17Kw+UVN4nA1WZtGDZFlzjEwd6icJIk
ietRWPMf/7QZg6DtI3weUdFWZKr+qltyLJuWIByb+1VREAta/p7AXd1mO9AEs8sav1dzijC76ZvF
r2gJebgeuSXmG3OxO0gTd1VHN6nQ4dRBj0HAj5lBY8WU3ZuhUfa6GYvsmdN3rt7yqJ9gPtVUZknw
dy+Pw5KkpWt0bqK8DA1OdmBVInwfrI1sosCdg9qVuI/C5KEcu9Qu2Fr1K5nstkfAMrhzgk+7TVE6
sOWEb07p2RxJnIF5KTz0DOxRMdbjK1Vxaw16GdrBh3ahCT19+B3vkzVHwNeU5nJVtkOGRzAbGcbp
KPvppqNpG+nqRe42DWZBzv8zWZ2Z+EdAyzD3FX29T0bOKItKSc7cFAuoluvlE9KYeR6dawJwyxAS
BpsBMi73vvIbxzL5T9AFCM7Xpbjv1WG/3wtxGDg+LyRemoXmOmEvd5XlPGGHtv7RNZDkCucF1gWK
1ue2qTJLMPpObOwP/o57pEGodT4pObT63N/q6LBgZ5GuxV3lZqwuGIbpU9nz2YimlKIgAHKs7w55
DzEeJSRYOeo49c3O/V4WeeEvYXkzB1HTwHrPVAk6xgDacrtWhF3b00zzW+tFIPEom/ShSBBxyBZK
Pb1GPFDpI2OR8XxyftzAuKK6NalvtvelzD2kpVGHh1YAJTTOdrD4yNIl15CWrlas2Qwju9/ZHhtc
DNovoPX4gsWgu2c2tv7U0zTilyb6XvVdD3u+9p9GvyWyPdleMuReP61c3LjFIEBEic85bd7YE7Kc
GOxs+nHj8XFHi79WtZEMvhhautX75J54MfZJXrIwijUrnvCxUblJ2i/7ukxI2Q5qVk6qpZaAvvYy
w+/XepBzr05R4v/LVJTVpdGIa0LNS2CdveYZdt7HTE4IKvlYn2yJN5LXHLgtyP4PuB1Rigx/1Z6M
INiojaCxiecgk8PXQo8bRR/wgI3Ap6fBAp+bH+bU4cCnP92vuvgpv/xAWYf0iPRdGv3cSiJwR2hH
7pcf7MhQ17oFK3NsN4QDEvbUCMbuyD/SR1bUcTMuO+XAs3BRDaWO14X2fU31sAqqBmWtsRA+ze8k
6XpbyQDfA5JB0Cm2pPkPBGUwHRokxZSijYITFq1TrXzuwsBlZQMX9vc8VEhE23lzf8FaGYSg0ZWV
N5kFkbbG5QLSIOWBDosbO1bF+PNpeXRZCNaXuDz99N1zetUf04n6qCqgNcEXHMwihScH+LmOJ/Yc
HXcMYc+mxhwPq97jjKPtJHlF0h05KWBAUN5KQKCB8bO2ImWT8sqbE7R0rvmzSxk3bcq51+gvdUPg
Pjs7VsHNNBc5BZrDH0xb5JHQul2VUQ67ISSH14aCn2dE4GBOpfKQRp4KeSqgOHPQEWKhsomHb+Fw
0Ufa3Km6Y8Q0QM9VHLm25c88yJwMVRaiYE2G99X39V+pyKHka/hlgAYJRA7zl0r2lZKSRwnGnHit
WFoKEvUDUaAWeRrjSSRUD4zQV+a5ppHOlu5oohLqS6Iyt4vrE58nkeSKBkKhDnyxVHKLTiFi1Z7y
HhgtRNHUsX9Z5ytoHdGpgrWjWEw5gxSZC88iUZfi0VO2x/WZBQQyhlqBrYSYmT9yArWvyr5agzeI
0j4KTX32BH0hdWJa5ijE2uv8XegNrVHWuc2DQbjfH/nbwIcEhQB+NZtowuvsnnr9Aj1CS9SDiFBc
rid3GPrZtERzhd/IesyDXdLK3n5ogLH6uHmE3bymqhOOsW/eqV3OkFrMDwSbjZMhxbGpCs1LOCNo
Oo27MelLkpdVEY4Vg+QTOTYuzX/Vk1Idr/Rh/97TzFWS24bearUArn/VJpGH8PRfIIkGxZRdQ4/E
PEx0uIGgzF7B49c+kxTr6gBwmyUGsXoabEPGCUuwlRGzJIzRM89vBAy6NCiLk1lyvVrCbilR+7fr
p5ZJzUyX5gOlu+KtItqY51iOth2E70FnYdEEteR0h8Ep1p7guEgIs1KzB8ZJfaPkTLTCJy1E6HKz
lkT2G/sXAjZoKQuxmIMtyO97294CFIlifRH9A0X+rgKEPPSKwVa1++eCpQLllnmllg/w7EmsphyE
FY/d9wzMgPzuAhK7ysy0CHBfVNGxFrFWFMRUzb8wFrALKHImvDjhO3aEuMP6pHZrpkNRVYM4Kpu0
Ow9apnbvRkjoHYUJ3uIyrpvmAIJmXbMXIH4Lm5985aNuIHpaLz+Ka+wOQvfWhuCkqH8jjpCXtemg
ON5oLvQL+cUdG7UxRhdzEsp6nIcyTnznCBhKOoD8i32VLlQ0pPnlv2+XNt5SdfXB9jWQyqwL2G6P
MR/gpX3iqKc72llY+1fGdz9T8qG7MuY5CAjH/wn8/V9MBHqiObnCipaaskG/M1o9bGXQQl3tFMhv
zqZFJ0yFanfTkuOMFwMqwbdcXxhjyWaLGYjPEm1avFDbi++AojpLJhyugZgRpVbnmJYRS5CvEmJp
2etQgimLYP6f8C/OdfBpZG+qwYjyZXdZTIt0JOWCTLGVT2IQBpuYjUPjW2Qs7RfQJnC2iFb3EIBn
PiBH0dWnT/XqtziVEroziIRN0GREtyglGL8JUhfz6pZCZjU3E65k8kf7zob6GW0mJWV4ZmUIT/5A
Jqz5SgFcjcLCTNang8a8lkYzK/0v1jp4m3hkZ+zBGwoYbeXD/NdmhPEtiCQA8Lw4TBj37gM43A0y
WZvpDw17py6xxz6x7Ghd9/hvZE+XIcCe/1a2Orbi2S/8UfFoNTigZQoWQxP9mT3j6CVIM1BKl5S4
1/bY6B3SBF/ovSUW0+dc0OKUrkbLArFRnZHQ240DjeuaIJBPtX6jvLU4ioAZl7Mq1Vqt1JefFAek
3sCOfSAeN3pMthsqeBt1Wt0Wf6eax/F3J19aB4nBMG4Xppvx0ZIdh7bZalI3hauDplzh6Zn7OwZA
nIlqv0zxEMlutupe6AiqmNJywrPhRzzIYEZ9Lb+bqsLno5euA3M2MYwWAsFr+Yahi6JtMHQei6q5
JjTgPsmHnKVW+5EDci0fI4upAhzUaJYqNyVZ8v9QmXN9SmjFK9XOB5viyQYEnmdzV5O4iayOgVlA
c/vdKcYFhBfE3bmmAC5++kWMPKxrFu3OS6iCRIoVkajkIMJY1l0l0SQNlsgEiQJO6atlTRZBx/2p
PSQcDHIlZQaM7oEC5KD960IiPzmw2EV5x+8qzg9qzAYVUrgD8RtWapIyHMVoz9atsgfkSqJohlYc
Kys2BYneLt5YFd9ZCa5AJr27Uti6ocU/oDza9fnvEqLJNNNlsLZD+hf53tNwINFZzuho3WSS0A9S
uTxesRfOH9BPRnxREilFp7WXrPV9BfOAPrVAJI5UoJdDyeiRaUnQbYOlxXF93t4GnI+MvCWotzrV
ichR0+FKHmO0rcbi5paCAx/nQRNX2uxf37ihBX0ADjKogAadpZFTJ/5nRm85jVHvo57m0oIR5HWe
2Iur2S0787+DVBrnhPLD2ROS3IDXBCTLzoaVwiRCdrJUMeYP1gn9eItV32QjWlskKpbPnJsksAGD
f40uKwqWQuNfVTbDhKmI/eVVovS2EQ6brCjzXrfHQciPqdluI4Z+GIWVBSStcsxui19yiYJtMLSf
VkntNZDdH3tIgzknvqS1gn948rND4zQ60HlVTVKvuVD3Wn5HOAEaQrdJsXTO86t9FU/p4jsX5rz+
vV4ydwICj6hDgensqlKkmYzC/hsiNYLThsmZ59IbKO9JLfGSThSvegvlAnEIfufniwR/TnNpjm0k
Bb7MN13mkHQKNPeZDMkrjnswoy7TfeAJVy+EDlTT6pxMhLNTwbRxKVaMhRkOr/La4Y9RB71/ZmD1
UJ+4SkaQ+FsJfXEW2jRFm4B6izXAN8yaxvu2IC+9hu2C9q5rc1vgio13S6dnQA75t27LJVrHGa6B
FlG+vZAdp1CoaqMBBI3pgV4QqEX2QVu44WjrV5pbpG6m9P79fGYfu/oqypIGQlUH5EWgARqZSIQe
sqYVhCsGLzqAKBJtnZWi9GIK+5IuYrPaTZTaS+9ApFS4rqcPDuc4dLIpREcBDrNCtPlTHA0j4m/B
I3RgJGhibDxdViEJwx6RJ6JnK7BXpfKcMMsSh5FRJK0sbJZncXPac5TasJtyOtfs9+lcyltSJlnw
MhZ4QY3NHYrN/CpAf2suP9Ho2LS7IhehWtFlxlRphspearwznw6/A6cgGowPtqi6R9XerdGUuo9S
7ewCKrhUlA7luHz07SIVD/AROv4z2dU+Ob6q3p7JZGD6288EipjJBKZOZMqVS88oRg82YAnb/zI6
CUeokEXqiKa/esDyg+4hYav24t0sXfpKi3jIaPCzeR2R//U5yLnVa/t+MBCnEW9OQ0xk2Np0+bEf
Y4UPPb41lk2MhhsRIatAFyar+d7zC8aqT3rJLpOqL79fzeAcO3wEd+OU0ngiroug1GCV8Rtgzxdz
2sh5dwxZBf+g+BEijMfvVSZXf7g15ZosfBTA+M97DtoSKS/CxSUWdZwRpkIJvKOWV5HJbUqAkCe7
giRolGkqwoF8+3GAcdKTvZ6qDs5f70OyuVhjwbiB7tKQn7waEvayYGuQm/szstlEqltnw4rdhJN4
XhCk53VfGhCRblX+ECbjq0BrW+aIMSFTfr/0UCH9t+IRbcyslCszKtphijriTKxRT/s5rtV1QLYu
lmUOBNMaVpaIvUz9zpWfWhefAl+OZQHjVU+1boTfUmJfxZhoIrJTBrBkrm42O+5zxH846Tdu5Uob
d+YDDpWbgY2KJhCn3/5TpnizKg9UxoAO/PdHscmm57A2pde5heGSz5P7s0iAXG5Rys0qgqlrCVpR
1S6kTS/TpHc3FtBPJQ05HIswYlpgG3EvjQp9t3sWxSbaF4kY+//aJt2McwvtoOKCyJW2cToRDiP6
NNaOeh0ZxdYVJWBf9hjT6S74szF6a91aE0m+9AAnaPwsjhdlSj/iZGX7qR599e6xs3i132MharB+
4AVXZL4JqPWCVF76TO+N8uB3k8cVSGzV4oHfd7cPTinuxgpat5qFb9HbzyAZQ9ydhpmaCY+a3zm6
Chx5VyIQNUHq1ssNZk6nOMz2mRQg7840uf5hGzeetYkjnT7dH0UDd7oQhOJD9WnWOJGDQ7fZk+HS
g3M0JlIHK+ndl7jgUmmRFVbvgk5OdQwmSs63SbstJeBnfO5aSvI/DgdgO6L2C3vaU7QEaTC/xSqj
4hhtENMRVDSGyemYvq7kpT5/k2AkxCd/AhKZoOGhtNxWdrvBPB/Rpk5rLfR1tugimbBGmvv0K/KB
Q0GcDm1mx+CKx2ieRCKqJevgYqVdTKLP2YqEwF5V6pKzMLo4H5I0hbVW5ob6xvBgZcH+Eg6jgVeX
7YtQyCMbsIbkQCkEvOCJjuyWYEK3F975NZHfupPZcFnWXMK0I7xgc5IOstPzJw2wJ2doN8HcE9wI
FEdm/l2xbSbMXBbWvRGCBTITe+4VwpNsc6V0q0/3S5cockx/qIx8NxqiZIios/slxnSwx6jHBOok
rkPm0Ui2lq6ElVn47L86bEWGdnGbpiqxC9gEigc1BoRtFrlYFsTxOuF+lAZkPFW7iH8k1/ovhqDH
vyuhFApzQw6fY5/cYuIhxYJPYxycaAqnqtHyr9Qj3eS7MWubG/4qH+1jVXNUeLyE0MwV91zd+qmW
0y+6IF4dT7az0F7m032RMLRbfvodEbpoIDZ7h2RYdw4qztshnue1d8tdEW0JD/DINXGolx27cwnn
z9ie/d9vu2YQGwxxky5mHfi9MTJcMMFBuM8Y3Kkq7fDn3LEMbAf8RmD3ruAy0Nxb626f66hfxZ0C
LD+k1dAhXe3+OBxHaO8R+7KlK/1Js/hX25Mo1hgtv3qUnY+Cew6KVY8/aVb2hxnYo7UcL9TZDNNA
VQl0LBY7KMdTybvFKg7dCNV9NFVNX8YV8hMAhyMPprg/NtGQDQrKVhZpe9slWbHTALQ6R4RoaDND
ZEpTC3dfZ7RAKqRc9OFWJLpn0xEB5O3wXT8aJpnxdJpaXf6MHGjmsnxgkhSt9qgexxufCY45WbEY
82F2PdfQlp/KRgPpiWKI0DlKl3oVlF+4vNKl0zJIsWWxgWydEQD0WP7vPEvrsbhMTrhsw7xpmC7v
1z25qaWZBCrkTniUpe1Z4eYtJyFUWRhET59xw+Tsl15VWLGiN5qwtNwV1S02n3y7aWD6LL7x4Vdx
UsyEuuoyieiQ8170/ppGkS9TFb9uVwBXJ/BI0wPfrLCJ4KxOE9qyK1581JPHebWbLVJnDt4+4nk/
/1l0yuV9rHtIVUYNJ4kgT+3vVtm/D50lh1q6wKr0z+0HfygvNCsgWLFNATFkMVTUc82b0zpsErcH
kr3aaamFc/D0vJgj2rGMhFgD+WOx3KPOyS2WUHn2KqFntHA0xdhvr8F8hNrAFqo6093qnN03Gs4C
8XMx2MOFGKj8knNUvNhSeJj+DMdRKizl7isDKVJnKCgFm6UVpZS3liMNohjKhkAVCJSJeU7CvWZk
VEyCm6V4Fc29+6oWFxXmQS+3dNxCfTnpJyto4nfZfVzo5lrqntWgop3BprK1Zgb5Z/g2N3zNlAoC
MwJdLElk77VJrEA5rrpODPOKey7EDUZVYSS5U8nwzyXII1tLRlSEbS4veI8iJo51r523WA74ANeU
ddjAHn1KmNyL/RjjL1W3nOJ0JFf8bsISkc2xKmVusWcj07RB5HWfmXa/XJcNIhwiduJf26nwLckn
aw4AJGIIQwO4v1wGI6uw2kp8qTWvjItQhR8JddLWGxcM/Dj7CzEobGVEURSF+eFwt2TUjTrbW7hP
PoC4x78X0yb+3qRCDAucqLZgphW5x3hPsC24PC487QLR6q3hTlGmwWakbejytlzvWahjDG8JXu+b
1ibJ6iL5IbnTjPRjPVe4DhucMppNqbgskYMpu5w0n3DpIPZFQK4XtQtg9QtRD11O5sJNudQNYn00
56eE6ue9yNiz4LNg0N5tmzKEOJwHAAxPOjbdrCf0bvd3J1Rb/QUcA9J6H+bM/o8CLp9KR7KD6xKr
b5BA7cdQFFaVL8r0ZAhgy3thhmfpN+VXYum/XA+UwIdqdtlThjmxlESmqikwENZygW3LX2N8CpCr
Vv+S9xR94BuILYn8sPExoFxV7/F9/KffIzZtlAiy+TFW1v72Pon9218udWKb/vGwyK0P2quKBhI+
WOzx60zhNrkk49G5ztBuepCDXK8JyHEFoJWLJy0rncuE9vv2r8fZYWR+AiH1WJKf7jo/ei6PN0MS
nE0rS2KH/fkGTVjavoxuatRBKlH5dKxOmuMkysLuuvOWZEAM06/ETOEB6y6XG0TROZLWU9XCnFcx
fVfZA39PtYFh4stQ2KbPYU10qHCaH0xeRtU8UblEWqN6sjHgJkuhUu7Nt5AdZSzFQ/votSYrbvkA
I0wTjVmSb8Q2kbR+CxoIWtmnXQF5ECQ+GuwK19dVQg2piv9QdK75r1+m0nsc9vMI02zja3nx3f6J
f1n/Hh1DAIHgaSf4fdExTtoH+oNFkf4f1lGaiPQzjaMYYMC4J6cqDVNexnrBO3PNwlzoGSGHTOWm
54IVGAtQQVHYdjc4xCle9Dwaz4B7mHVXhCSSQXzEF8wkyHuMgNz7TSqP6uXGIsry3cVb+La4SJHI
GZiE3n5r0lmSGV0yrIVRwGc79dulIAQ/7Btf3sXy9L1FFRpuFu7ob8EEf620m1UBFTt1ZVD7W+zy
P0Ctq+jWzsWQAGRucMh9OpVpR4o92O+aLpqw3VvOsHpD4JGKJgp817yfiZcZZFl2ngKA9ltnQK62
cboBwops/QydiYRE/pv7l+Id1bOc+sMukHQza6AgU5AjP+NGNvcasO73cug1GGAX+v3pZ0O3MwlO
PDlaaiD2a/lc59bfPwKRNqyDC+RkEOR7PdLdFmGQGQjm9QEAbIEH1d8s9vp1S7ZxgynFroOp40gb
Wd+b1rmmFWDYIf0K2aV8WoLC5Q/xbrgIiwSjTweMX/DgWnK0FWxgPJpw6afOAdu+BDSE/4FJNklH
jRIe8sFk573QqC13CN+f/iTZBgbJq2iE2nkri45PeJvJmLF+RJaCuIYRFUSMPgCFVmFx+0Uiq7i8
p1dvh2Ky70oy7pWpKmO62ogkexTVZHTofluTnm4DeKXCBo156DrYBU6ip/Q0a3vS6Z38p/zLJQJL
ITfhcnEQ4ZCoK5RlcaduAEz7IG2dEFEPSKd+HYzH/ypSypGOfGHI08ZWI4NA9PIuY6gZWq2iNGu2
/GZVKoLgseXUBMoX6HPLMjNQbpYroFZrX1i3433KWv5PNLpJWxZ4q/jt7IBfjNcTLNaTHIm1Io/Q
V2A/8EgMS1pLWQJSqDlam5tR/mefMqBk2U/8dPr4sipihOw34YT1btQ2iPklvrA1zfLJB9eE9pF6
RCfPNa0z7QHHvM08Gw9w7cuVa2HD7LWYpvau88rhXUUXDLVpWg7kUzSgIzjnx4J7/EgwZSpngheL
LzUIWOb6DunL54JpsV6wcJ8uK1KynUUUXCtO2qAYXHirPJ+ainmXT1nu38PNtQbxtats8AnXiSzp
YhqIx1OTadQVgUcrMwSZlcJrWWpwynXoRFo3U9+2YGH6VxyD+NXQRo9lbkcvcgeQyRfaT7eUZ8Sq
9H+KXPRUgql+eIPF4hLn5xdxiYi6vlCc9Pm1iBJBfL6mM/rd26dMQn7/DbIfff7YXH0G9v4Ban1X
hPlMrU8rECjALg9HOkACrn3m6uLy64/GChJfa6ewLPhYw/6u8H38oB/wx7qhVPtepP+e/7m6Ne2A
dMoDG+uCUKFe53cxTdPtFrqLPLlvOuSlygHAs3TSk5P2NAEF9QrrR7pARJEJ1JQMSen6YP19TmiX
lh+M57h/OTaE+CftrE04Ifb+B3x8MX0T/gj1cP3BN60VEasg7/QtEbXFO6SlO0AuUk2nOSX2TWnx
0EGFdIKK3DfYojWlix0+LhRrXKlfM8JpuQbyZx2+TEExWbYzAEIdWz2NFJb5/bBPkDCYe5Y3b6it
3bP74wnHSBpBx3X2tfC4sbk+GSgpzSSvKLaGDtvMQ24PX4jRFJ7n/z7Pe7vUmwM6HuYyjFmpcjPV
HK+GM4bF2mOVlUeVpwS9eIvrs2a1Mru42gFVhtguszyUIzXZBvqzMBAuTL8djL4bVNU7yWtK+cKU
Zx4MNO6aRd+0rh2tWER97+/goMgZriiQbTP/pIxpUgCfKKL8t6i8xyFRYeq7ba7ctDiXbegw4JqL
uv5UUCwACYEYE+6rRYc4DS9qArxYKm1RXUCU4UZQwckND9ml1eQS0WFNBXg5O6Bh93CPe4qxrL4h
ThyMnpP4cqivjz8YQrqhb5ZSOz+j2eaEPyuEOndYSIizDxkZFNDGDgO8QYs5VLbqAaKyaJPhvj8P
CZTjkHsWgGCIt9jPQ+Q3D7nbbpc+/mNhJrF9QtVzDA0LshRrRkOfDqQ4Hz8Eom6xKt/BogUZG7Pa
jP+hjvjfpjm3Hlr+M69HAktxXQvFLlEeuGDdiHu3HOj3CybLXZ/w8y/rtOMBJuFKWiBwOgLX/C87
OWf3WzzeWZCSsYoW4W+w1/PvLU9ErZxlQvYwkFeGot39kKmJf3JWJ5fa/+y9SCoj3A1zvEQe35Yk
CQ69X8qxlj+Xx61esauWbGMi0nWn3pwmD3GhisSftml6PkiFT0lDdkIwxXy8E0W6fL5WrjEnUggG
nSwhXRbn83dW7zc41V2giB33iUbuWQ/z3GqWA1VZCh0q2FcAkA61LcBQWGPTkgjKuRUfu/6egis5
SBlWyqETgONP8G2AUvwZt1/RtGGafKhGq6/qwjHZWuZo5Xvbh800VD7fFIaeyxin3YD0oBdGFI7G
p5QhpuRPhtObISOf6R1kazzIcjbPl8x8z1NoHOMTHFhyI+vVNPCBWyD5bMEJG6QThm2kfawMkJZP
zw/CMpewWDlN2Z6hHPVC7if7ONuBvyKLzrCQxtC3svhzYFZ3yFcFStn6frJu0Rt6THq416WXcptk
Ni/R9Cvb1xzvAdfd2fJNuM3Pu6pOvmrrc7vM7qOEA9eERY3UhKY7cUEqsYQ5zVCaIqo89AADmko5
DkAzADvF/e44KOcDKUUdMtTu+AgFKQF2SOKEMHHoR5h7Trlh+q5wXK6DqnCg3a0kM4vS3k7YMZOb
W0u6ZlgCd8Akh/bW+wlpWc1TUqdF97ZOYHTFUJ2tuZGs9U1KyffxrKQqVdO3U08rzx8KaTpbtFXa
ElWtXftrY4WobZKQvEyO8xlwtrjAHwXClrnQFFwOlZCbq3QVtybjjgcnc+xl3KZwtbHoNTGXJC6N
26vHJJH1sjCogBw/O7/3Cd+jphQlN0D5hutkY3Sn0PNkeolp9sv5dbUYgwGFKRgS+D9UOFcAffHy
ERntIe57/gZBgUFMwL8ZsJZL/uAjcOFYzH0qIC4AdWIcfa9ptlXuEjqrPUo8pxIBRZdc5zwlq+1T
/HMVZXGY4h2aCYMTj9116H2w28O74Dq8BM8zRoxk7Lfdg0JRhD+6aMl/Q3nmFyx7pUypsLrF30G9
fxFSjZcB6FwFLObwwywF00QD4H/Yy2vy0bICvrbKCkjqtmJ6bZRmXbPNv2nRmkakMxt28GlkhXZS
L1XE5QUIdqL4XpH3OKghmXDUpv6CJC90CD2zDXygkS5lP5agngnMWAJ5jJGeJl+5fZzn/jAuK+M6
wVMAMzG+nKHI5Hgb/a8AnSvIj8l7wrz0w/DvFdr51nK1aiICxerw8tRWHqL/ve5PycjYogmQjCXd
OWOU0DUcunZVT0iuYamzjfbjMqI/SU6slw/6a8OolbKtibmA1ollJqLO1QT1JD/9aFd9zjP8E8CY
9oPkf5siDOn7QkaygOj/DLpllQKYPosO3KrUrk7f8NEfcepqUR0h8j+oci5y47O1smq51XNEjbSV
u7/4jQHZSrKFgmDRdjlAy44Xpc4K4so0PXyWb6nbvTzUBvUzwIH+ruWFlvqDGrltWdtCw65O2Tza
surzZQzgKvEena70t9kuoxAXBtaRG+Y6wsU+HXJ9wWvQDIWr00iKb+F54kNJTI0kfm/Cd1AhZP3B
Puxc/b0SsrOtSSlWPiRVdgMbPeBiyaoDHitJ+4dWUeW+HCSzVLgMzfpXJzoBzFvIe8xQSipSOznb
iD+WruBkCnoRW3ED6WpzA2IJRcu5fMf2jWNYkIAYJPDQV6WPgdfWBY5uzrEI+06SkDBgNGAP9/IG
HN1Z+YlBn7n32BjdeT+jAz8V+0OgLReUpJhM6tmArO3CllotruH/IKXhZL+kWFWD1q50TPjDK/5s
CC0CWEyHQ0epLUejtJJDBGgkuIV7JqKt6Hhn4EzoevLVOJXXyhi9TGbV49UXETxKpV1XLTIdJNAs
xmR1PIANM9UllM+TFsMGFQjsTQNrZRJTLq59hhuOCigIUksvpE2/K4b1JWCOmjT5zvugmglWArKp
J4pGwuwGmdK1mx76Ph/jX81PBV+OGs5FwNxgAzxcChu2kLdPGBH1UqUf2NX+aUeRR1Xu4i+mSbxo
dsnGiQcXjKU3y9ZDCznZzUT3ZYVvSw1B+fv4+S6rAPbOHck6i6qJkoIRbPJBW/Ah2917VpaYoIk+
YL8bsB6045dF+4GjFWxvxOATNL+WR76i4b7as+Ezg1KxvDx2A3KT+6f3gd14eK0JM16B664XhQiZ
k7Ad+9GnYsy7+hklO1JTlXQOUWjIehlvHQpCuzYTOZV1efXHak+lmN50HBxyxlFGk0xM1LrUEX0a
kuak0bp2F1LlF53HVHvRJiu17t6R/wC2iepZVmJs6x6U7Nw6I90z+ZCK+UHvxf6LYASPXb/XL7hh
9LinhqVgB02JFSOFjAli66fIlbbKdsjcILcFUo617FeEfQGrb6nAUSFPnwwOrc3Gjr68Sn7aBKEa
xSxkFD1MV2V7wiLRAFqQiFjxeQtjdRZ7POgYCGJGyMAZ6NGWBEW60UEdpZ4PpgZWEDbEaDkkcyeq
RIgE8sCQZhM2xGNnhA7juMO2DwA3YG8k71gWHck7MZiXo2TG5AU78ahj9Nwsaq4/Y3sQnyC/W7c7
TZBMIT65ieQU/DBfGmYo04uBLfHOuVjAvHium3yIL+8BM/ZbUdi9OsZuEwmpgPmGYKBjlTMKK6Go
fLVcstmN1x8E+pCQKwldoAkvgBBytPmrQi27hwiJ1OvmmDX6BKlo/ccHqSgtq1CxAqyfvDDx7OO8
CYMRIT2XrnPN9alHyMkOv28+scBplHqI9cviyL1AaDaYcXGe8z3kF0aBD9ztMD8AOyFPzR0UaaNh
bU5xtfSVJvvy6gpGTXSo97gxRSYrQNG989Kx6Ut3MImCb4z/9cULp36hzkrch5/iBcKyY3Tvji+D
Vk7cfAxYDEbZo8Y82SCJpWV2mxXLgseGy5DtlhwZHNkuYa1ijD+RsArsTVZEDt28rlXTt89rh5P7
DzgmAlHQEI08JMyDeynvVIq6ZnCQd+8Md2A1cpV+Fgjamt4d6YeQq7R8dz9GIlVkKxW3br5WTZPq
sYY5aDtiGkeRzYrhmT2kajvvViFCKPdktzAiUzVSrYeoeiQTBE5sGEVdRcawMVJxWJ5wBXo1k9wd
Ir+2oVP0lkQEH5c+eA1AkyXvKgdpyCvmoYLaPujGb/oj0Dyfm+JpbfJDpIN6KOp/YR516I0jOiF1
qggmWZcAK13Xo9hC+Lx/s/rI8BnngYLhHZjvPvir2iFY0WBeVlw1c1X7CjA4WxYGxfSggJ4oVn+z
VQMLi1xgId+DsWdXhq2cD2ThEt2VdMxyzEr4Ffse/Itq1EtZupPOJ56skxk4MVpQ2B4yaaRAPh7y
fq73DdaZ3etOaXHS7HDL/OE9Jn5VVD/UF+HdmY7JAWaRn8dQhGBFFMUd3SSgUi2/dWuNTm1t1WM2
iRODWOlNWoTapCuEjV9teu7MC0TkOA4TP4yQnkhxRapZoE3VEdT/gJxmKv1DMTiWw6tAK3h/8+Ly
z0Wcnr2mASesPv4q6pigqoP8Fb5m7bCVlwfqt5uiCKwEQJ94mzUyj3UdJcq+kmprLc2JabLnjsNQ
TXAOpUgGAGpv9/xYg/ifePIoEoaac1mPb2j+UTfGT6+tc/04UBUG+s//y65IlF9/MZHGdNYgTFjf
vkF6TEuZSVA+cmQPq/qOSEcmF4naT+x5F2TYZMhwVrjJmglm3eS48EgLqwAl8VHmWZxt+FZzzlfH
YOD+G0d4DPWiWZeyEqHCRdOGRQ5A7S3OwfS2q0IYYOOaEDcCQRpj7KkWkadYKxV9QH7n/or0YEep
mKfd4Yh8w/Aq7AOL6m5c/6k70xHEENDDkaCFUklnxIkvs19mI+eclmYxImr5HGHrSDKbAYiDjMzz
IlmRC+4cthtFFa4NMDQH8kABP7wHIn7+eOV2HtqjZLUKjUKlTJJ2R5UdANBibk0kQ6+/Qzan0Roh
cAuaPmsalGNPB0zmj6CNYK6pVr9iy6OoZPshWciQrk5IdllinEHJ9TiUWmlMrnHApvMuhzDjvz5S
rf59mQlC28QqMrd42zBUr2BSwyIvREN1I6WQIz1KzAUEx4IBMRSUrB7qZBzQMKSrZtubMFH5OIVx
rF0TOPZy6uJiePtBZK9pahuUNIwLBo0sMmzs6Tceqa+5dXdA4/0cE0TrrdWCr312AsUQTRavbzOp
8zdAok2ImRmPn2QP8EeUGmaTEv4sNdBksAyYJaxcWoNjCt4QnBF3dS0R/P8Lo7LpPaFHPnM8HDi6
V0GQq11eENcfTCx9nO32rBFdjB844C1+f6HELjoEtEMWwwnlifGMq37kC22XPU3+FGpPh6y59bhj
w7aWZGPctrCJl6ImQ+MdKC7oyhgxpZ1mkugypAVFBrp2naVNzxckCbCJu6+MGRwKDLvXGjsGZBO+
NMiSlAVOfrSeajc6puOEKpABkbFT/Fg4rxPqenYQ6dvywn9KFMel5JWQ3rqt5Aj9eX6ewyNX4DC+
89dhrJghfNRrsbcz9omVUDxe2+71mw0EjagUZXDoMtJZO7In0XMwTiTnPjSxEaJGO3CgO/ckHtz2
OnHLkuNqCKoQ7M7laSgXed8hySZkR8sAnCv83GB3JS7JFq+3bcK+FREaxx269wj/zz3/j4ZC3AkU
jM5abP+q5adbqbuMC+iXNarbGv+xZw8VmnbBUBz3wiH9nrB6vCOoJyHPvN61OfytBpivACs0DUqH
JCneYlalYvJr9e3avE9X4cB+Z78xZmSa+3tJszR6AWsLfqFslIq/b+geN+wU1F8C7QJdwBpaaTIz
QY3t8CnBMjy16mVFvqpzM9ZcuBDYsocB8M8rfd4LE43BK+qpWUTMsIizTgLN7/q1R79th4O/Luja
NnB7xF6sZbSilbLCdA3GS7lrkhLqEx29ojTULe7+27IwNyOpwG1sWQ2a3CxfYdkBswOeBMCqe3rx
/yyHxHMJZ2la/P0Q6KORyjLIxH/KkpAomjtKbM0uGEONhpRqQ3BwQ0VNK5FNBG+GwUQCBar/2r6u
O827k3+9FiuR2otrNnnfKbVORfl4RFzYQ8ungBlDtGLdEWCNanlNJUYFDkw5bWDVHwr4FjfkNsgP
sIxIRgr8RXuHTbhWrDnFc/NApUKvHBDaTIt7tAuXIXBKtjVQLWCUepkq/92AX0eGFEIjMtfi5E0n
LebiB0oyxHDAA6xoZ18sq5J2ijsuQAsjttjulafQT4EADvGlloM/oKLPD5y+S9jP03TPoWPX8zaP
fdXxSwxeUgatlonvLfKDme6lSZ43UvwDKXbraNY2V6HrLjlDWyea5FSUns+rdoxt87j4hoaxa6nb
6wHQrmw9ky1L1sQxe/8YF4B2zxQvTGg4gwd/yFUR0SmfTclvM2woUICnwtnuXlOegs0StIj2SxFA
MnRE8LnPon43CcO3EUxiZkwB2k5+DTz+nqqYQc6H+XN165sBw8DJzbBx7TgqHkuJl05RqgbQgf1A
4dvPUGdbrXXmyabxfBhPPDZzknKa5GMga8k+QlDes5KO2H9N9xxcQdeTZ9SHHZQRpN+ldbuX1Mt6
cX1xH0xIj7MAxK+p8i8XnSkvjVoMlO0xPiPNipP1ZaHAOR3X6aw2xY1GaIJsePFwJt1WjhKnVnzV
q4V3aCn7gdTKI1XzLzlNH37RR7PO7tbA1eu6FNXkqdt7IXtMeIVFiA7EetkZeBRPuQLPfEjSQXS/
ep+qsCHLFkX+j41r8ZioPTFictggYdMs64kGGX5N+t/nl9ZQgQVeTgpxqW4SutzQvcBaGrVKvWBC
Bf50DOnH0RduToKTzYniZsWDX24ySkLzkxBxdlFWorvxFGfC8o2qItvM50aSY0AtAL9/Nssi/qK0
ktKs1xgMMuwhMn+DGFMrogBled5H066gj4puFlwKxn3LpoBSJNG70oNkl0Y7N58kfbUT3+jMltMO
QXAwEvh0qIKX7Jnmqm53VrjQ8+B7tsDJyXkyubcv/9X4Xo9lxK9VhU8r2lixBAmg8ZajjuUsKF64
lk/1kWJ6nZod2zz5NF6pRpfcQrdWaIhYBoNwm26LZcz7574F4PRoB6zxbi0Qw/XZKg3WNMKitSuX
eb3gI8VBJBSaDI0i1c5V7zZVKG9M6uInWdC/ikkbsUNvAMSAzRJYyUT/q9tx/ounNXUnxRVvMITx
kqDdGWWwaJ1CNPNNBhbBgJtugLaS9Owfy7flsZJgY1zo9wPkpnKqlu4+q1Yc2yDnf/kNCAsLj2yt
jE4KiGejhiZwR6c0Sd4Xo/SAQm55+tTa7x1yH0qZNMmHeftN8lRwr1tFwBFQoPMLWBGmRv4E+5Ys
NAKHhEPJwDkJI1xP5E8Y9zcyfQgTWA/SzfXYazUH0aSQZg2kj3IqgEzL36vTW6P6L4tFNMidrRIn
PCCJKnoidDwVX78SVby4efdzY5aYbW6EdMgXRZjMc+TP4i0fqoanjcBiY6QnI7n2QKDL5Rr3NFub
x+nHvq3jQXLaCE8pCKmodTpsOoXK7SFx4OhGnf2jY9JOlz5koFfF1dJboIB2ODANQ9NZPnsw27vZ
enk2zKXOry+5tYltPFjxx7xj+GW5HA/ApyAuAGBb8dgLaWMXx1ZMoI/4NpPvbipBIWbC99gKp+7O
qpTRAXzj4E6TF+Wa00aqjUOVkXmB2Iougq12ctVHfLHUXVn9vsFT6QPcVVWtDsVfPMKbKmBXart/
LZLGqXHmDlkpqry/6Wb+5BM+vGIizP78Q7BP1xNoLD8xbsWyx/JwqUwOU0JCSQODrrEHfX2Z7ftd
o+GVaZqdJO7Lmcr9QOkh0MOFohowaLon8etCHkK5pCxXjNhBzMZaEsfxyxC9qsCEApRsi3ByYcoW
KBQp8L5yKKn7tKRl5b2jFdNu63/GBLDuEJ1It87faZNErRpzs/PPq2P0GbQXoMdmqfKoLfwygqxY
2XM74tn+Aq2hka3FYMmd1jUC0uHOG2hELOrmz//zxKAhI+hcy5CUJuuCan7/Bip3N/Gq5np6gb+v
Qm7nv7/RJUXCz/uVp4sb/TyHdirZwFBNesBDl7hBn1JWeh+JHu+9RZ8EmxSYzJ3EjOULUYFvQR4y
CXzS1nc6LKN8yvGHkiN4TEi7rmG88LFpA61Mq08p9n9+17eiLq7gXtgKMP3KLSZfufYH4nkDTc88
+PdQECAaoT8m7ErDmZ3+B+g/GHE8itMNrpoKyn8QNcvkNdwxslaYVEVsvnYna+YL8VYxJf/whWxi
m1/NSJDzI1oHQXK18bcW5TYiBgJPpyqAjE8ArjWpyeF8xqQ6Zyqgu/iGKCWF4ui0X+OLHQGY/zK+
8toGWpr6LzcU0cTxuXr9ntO2EPjR8TvepoRelchQPD2itvbr9u7LD5ha9qZc9CgIzl2zM910fqJ1
KfY4z9VgEFVX/T3kD/GUp2SWN0CIvVXdv/9/kyusEcOf+B+8grXzc3FoRXZpdbKiHchkQYKyxZ8I
FTxHq39JoL33LG5w27JTPBPQM73zeZWDD45+uFFUR6AjdZMa7f2KiaWPO+fI8c9fuA1zQvQx6v/4
Vrt3lqxgCg0TjOwkEg528TRcsNcbGb663uoSeChULhQIv5bTItR7O5UC1uab+Rvx5w7cZ5X1j1Jr
JLEB0qPMNqIBJqILYwxqMppUXK0eRwGLBrac/6bumHhKta4zERNon+8knTs1O1G2LsC8OvOFR25j
rbWncv5u54icV2LGFTknizdpEuSx76ahDKqA40zpNjP3JHQ9SbA7QFrk7+E6AWbtpciq5OJqWb+q
9UiwQKu5qkaasYUV6RfTVfv73lrqUWBTd2veqEWouX6Z8c52TTbDvzpFjGGIeY4M1rJL5ZfH4KGC
iyo5woB7xwqiJ7RUmJFa7Z2KVITARoa1ouElbZzl8mdIe0Q3J31UeSA5T1FWpevcjvrgXtwalIka
9/304isTMoaFHtNrc/3B4wcPgshHQ/uanzuJQXsToC8m50LBlv4GYoCLRG7EZRHvwXTpmOX7s5BK
mPpxVRy3pzvkjSxJDb6DdgPHKqdLrTiDzyIYWCuwkfaGTbFUFtOI8j2pdNazyu08KnCb8s0z9LAd
PkNLp2XTZxDn/uOOkFDInptrDIwxHU3V+g9CYR4NoRIRYwb7ULo+VBRXMhkEsz9lhJDXjXGp4iyo
sGjXSOiVmMdYGJuq628Cj+gGH5G9J4azi0QePfcJLaHPbNuP2puooaCEpqkJxifF5xF1MxUygXeN
+TmaXjcG4uUwblXOQw8h3cX6DnhK2S1bXQfoJXLpzPaS8BbRC35JbrqgSxWO3fW8J9x1M+h2a6Qa
KQg2/xverzOmgSG8AxZjJzXR5Q70PouyFPfaGEsoUJh7QWrRwwR1ficP6LEUI75ciJEq9tjgWQp2
4+7M6NQNxvwVUQ9hyV0hqLKuucCX7EY9QGoG26LdaEX3jsMqhimghQOH3dSHDfMWa+uMm4ouVXyF
yQ7GCPso9V/FNxYb8oP1dUNM/x8JTnsYtaJcNZxba5POAI69Edz97Bd5JmBkOWg3Am/xbfJVfSK1
ixR7KIHdkgIH02jnzIF6yh7jZYaD5GEIiAG2YNMsX0rrZ+8hmJlNTzmetX11P1QOhjMEaQGs7Ity
RaHDwSC7G0PNvprJgoRpLRxe6noPUWai+zThP/gxNzSw6aE+m10aYtnmL7cmwBzBtLsGTtxuU0/9
isN+BGTK4UvbJK0qOKF00icitWvkLUp5JaXJkCZ2VWBOqYJXbJR/7uThWX27PUOYwDOnauiC9Jx/
6ZPrAUJayt9C3yW4AlhUtsaCMjIqzT8lSEWtmWfhiKrXTICWbnmNt7xJc97g04xtyKk8D00MZ9vn
tJBx9a5wLdGKzmZ4oqVsVa6PT0kW199uA93daUQiQrVit9mbWksrre3QKo6WKtU12zBtW9Tt78Yo
BtHsD2SSgmDIJ4aXMVhCYGFE8i70kufBSLRCiiBlGQm3pOYeFs/AtJZjBKIjV9W/j/MJD1d9+vwW
TFXF/yizAb0Uu/LP1aPlP3uJrBoEA/80rdD7HkVhfGa1xT1L4lpDGY99r4lkLgtD1dUSgNZRyjnt
yctJ0jLLtkDWmTzelc7iX8KyIZd9axD4PHqyCeXBsWYKUu84odiRXURIKdDI1bAFslM8h+/kuCKa
La98L5h+TNlsV+kyrKBdT3NmdxvtlGww8ZzI+O2gqfBWe7qgdKYvOsWMkgb2kwMPjHmf0O9sPmRX
SwkhdqaPKU3U/8fQN+XNXcq5P5TeCybBWannhkmEoX6H6/RUndnTrPV1lGJ+C8w3f9/UXGqSnO7r
c6zpEvg+Z+Szg7p8nvepOtQNMUgNvosUrgAjdhnWDNILQoHGpn/yqGLV8FwT0L9weKFGZx/Ces9r
DNbhlb/BuJqPwiSqCDWq3h0JdcLtx+lI4IGPm6QJ1EZ870vQKyOeoiWJEXxLrGtovXiW0S3zPgyZ
gqn3br/JaoUPuIwhigHe/1SAiMjDlB0eUGCHq7ME3y5oOvblzLEkCxq1qeTdXNYKya6KFQy8Fipy
LnM3QNN2acc8aOoYKSFtfnCE1xX5CbeD+kHY2U655OlETCwg9BL+Ew4LXlPl+j668anr+taPuhtU
dY/1WtTBPgSUQK2RaB++c6abyENbgptNtcRRpxHdKEp1xEBgcL1xSmbtePbTNDwJVgZO9S+ANsn0
hhcIlV9nm0I6ooCD7XGXaqWtvuonacEqw8UJfVw5PEBdD2CXrXpv3U/JAWd68Orc6wsvkhkPDh/K
UZU1eJbFSweemGi2TZ9B5jvQJdtmV20FyeZjsIxratbbiCnGmTIFGTBF52SKP8fm7GgMGQJkZfAS
pmu4F4s8IbIPeRDfaMuykNKEbKal9nvrtpe4/ycEi5HB5aM26094BddM9XH6sJRJC1PayAvhCRaN
f5l2luY6OG48kC/uSnqf4bWGCj5M9Bg3B0WkU8NPY49wXBx9QLM6V/2+bL11AorOgynmPq74FiBK
lzP3L3ch4QCGiRirZNhcLu8fTLXQwBM9F8fEFa5PYqpjjdBv5zguBZ4ILHhzOyCbq3+P7MAm0/Eg
Xho/rl5Tt+APMDSQ+gqijKP5+QWN7l8eLA6f1y5ctdN/7Xirc0/98Dc8rkNxPBILGEz7MJN2eurJ
gGYXBIB+b2HhlN8xbqD3ktk6jOpCacrwRXqJ316OvC9qKx0KFXDXuwAYHNqEZhSvNwLiOwitQtX2
YuVEenIJ4FfvAxK/wrVsCNOMEVi/Mgzp/WgUmXqSzza7kl14Gpkv+ZQkkMUMit4U2ofJxi4kSt9E
UBWj1whzMY0B2I5/OPu0RSrFH5FJyvboLH+CxYlo0q1U/sfJGX9Wff1d2qfNgdXyhs3ptavbxyHy
fsCzmBo1ZyiKRxB9tR04h/2e+XVOMyyn6hvy0op4+pFOew7nE9V6Ijs6fzSLbQY/sUhhYufvxn9n
OJ+xQF46ne80RZoqaxtLqGIxqos4lfGw6kPphBtHa1ceXGbJxbvIp/31wDX0airEPBtHo89F5Ysq
jVw1cC3SCTF526eMNhm4d+UxnqzCd0lVwZSfyHzvDbcFT5MLTvSjJ/MZZr6aZKB0YA4ezFZpxDbE
MIE7UWhrNZ7aTII4jHChEYON5V+9coXgOIwa+15y7Kn3cdp3dPD2o1XUECuONsC9EDXxvmOYFikN
cizra7goDuwLqWZyHv2h+XVACuVwi76zvW7fmJSF6/SxaovcOlXhEZvJNVt2aOEErR15MZPGCFb1
7/UTDjCG56AfQLEtKGFQYBGHmaYQ2F4gBjbVb3CgnHcSbFur2GVTBFBj+aqjJKPUKfldYyItraCe
5od4cvgwdy8yPpI1esyIkls6Ku9/yNz3BMjppQMziZdVhi0FC9k6staDifJ2STdbth0+tiVzBtew
NyZZlnRSzQyDKxkVUSnUa1CeNdMwT4OKku8RwbXmPQ3jjGshwHBH35QozKcDu+p5OVdx03TK0b5N
lv4/x9vz6CLaCO4f9PETKHEyQW+nqTQ2f0FsathaAZO+v7L7a7GgaH2Rt6Qqr4GvuzkQWVi1xAM4
IO4ywCbZgWgQLfAI0OJCKE+uvoBtYgkOUozpWkhV8Pwbyl+4pr7jzAsznYdqxXKISkKYLMh/FuDJ
JxxeoAu1ZoVROXEGkj4zOtfDBoUmdQPfEdk1i6klRlu+WzzauMKGc119cmQCyKFDBdg0pkHqWyeT
CU9jHSVRfTDrnO9lbpiz9cDVQWmIhCESlFgpO107Qe/iFp2ZslIE18ESVVB104WjG1RF7ShwAltx
wIe/n5iS7f6hXnP5iwIG/W1D8QGVhS5Pu6pxpNy40xqjWw/m9Lk61rvo5R/iPHVQrJGMYP6Q10nT
j3W8wpNr1rweAQvvC0V3JW5JmoKq6vecUKdUsoEm6XR0Ty375DjAplQPIYEiQjex0JQLlAOOBCFn
Jw46r8UqQSBd4cWy2fgcdU0wSYGxyeOehYlWs4nulnXtJ+Y3+mFzAbKf711REj7KuBlZyTY8XBAe
XieP5EHl+lsIgukqpgc8Xn7ouK/f572PIKmIzwy14vt4yqqBcqFZss2K29QkQiGUhxy0QPk88elS
jhM/MRA7vVubvcNsNRQwG2QlDY6h5zlZvrFMOm+pHbBxd91mzfKeGLDfOLy0AlWd4GQV8BihpKJB
duzhk1rYT6zr6K7M/kpi/2UmwgFKB6wM44F/mtdrnbtZJZuxyOP0RDI2HEgIHIZABErsozJl/YWA
838NHRCblOfDKZg7tu3yTMH6eMNo0asoQ9IqjX+Q7+YnuW+Tyi+JXcZjXqUFkWflmzThkhss+Rco
hteHBzF1KNjdeavhO2DRtbtOzjj2gBwwcR4rWmxmW4K+qP/4rl3TYDVzal8OV3Ll+dUzbVs6M3+b
ueA2F8+BPpO58iw0vN02c/VGEZuOAfsxMFGqNDGdDHUcOjwVEhChBqXFwlJIZm+HycziOstLrfva
nFgE8PwtA8ML0HhXdDejfbRrc8zUCZM/dk+ZgabQS3fUGQFg7sKmR8vByi28ozRkdf6uUWZiyGEQ
KE+Jls8Iz7VuIds5Y7B4Lq/kaOmSVt2rfL/EZRPX5cDroin8ITjY4BjVhhtdPz24XMnZeFqq297u
viROiaoOWqat6F31Q5clJzx1jeRAqtPt7c4rkEOzyPapzHlfWRp5PfZtwdXV3Kdyzzpw8fMk9YYW
zKEt+WC7/a3NgqeQq8dSUOttFEAPE+KBB78REz7dcwlmr6fI0VJKxmxo5czVN8uAeSDlHw63td0P
ki7//aVP6qwEMED4YaO3bRVSN+3XvxSEl8imWvIxM0gBHn9zy9xbMQtEmYbrsyOOV4Rd4Uh4hmgz
82ygF3PkCTYOQ9IC94UHSgvSGCxcoTRNbKRgEnCyE3LTxtFej5kojzcdVa7dlqq8xoJ7wcLWox1A
zvBpQg8VwGuR7jF5elk6NyPk8xl0cZ6gn3ERFN8VEDGYXfVhPdhaNpqmXvVcodjJlIcZhAxUMFt2
h6Uqe3Gr0Cu+R++1WYzlM5uGImcrXo+zx5p7Ks3ca6jd8SeSnghOE/OBO7bUJRoIpH6bt1KLvxeL
5EeNaUbFH9rVqeCcLx9jrOMIKoBVVaFeYiv1QSCSpO8ZVaosEDwgf9PjvNoIpJfH+3FtuRhjPLMb
/ZOaIihfhqpSs9z2PbHgE6z0OJdZMoPZSpPWbSVMef7l/2n5biQzULqdSXBtjhH8HtrldzOFZSP/
5DCuTPKIVYz5j5wEwLc3JOR1yrGe5PCqwLwa+7++R/x9IJUudVrjZmOY6uMy1UrGqfrQDi22gHJz
bBr4g1uUzYqK9QtO0/3j5bWqp9moASD/8cpj1A+1YbZaJN2EAxrThniMFY2lwftdbrOJvQgGDBga
Bhgl8DfqWAzw+EiJat6ySaPwlCgaCfwB3Na8u1047KunEHDi3l1Xp135ZqOxSLmggKlNSwgOphMJ
yumAQ2sVbU/gJsc4YfLEhW021rSACYCM+AqMiHXdcJ+fAIzbeLLe4ltUcD8k0iU2PYUg+rsSaTkf
PaKki5MSaQvILK0oIwD612RUVGpL3TP2SaaUegEOxYx7OpWFbkzafmkjOOzUf9TYK5AslAUT2zOJ
0Di1LaehIdS4qGBWoAmex2dOPyEJRc/P/+XwIqsIHktyBFc4js4pURXlXaFnPyzYzqRCcwOMsm6e
UDMXgI87or1B45i5vIOOqfxvvnZg8PD5MVobxQSMwhb9Ld3+WSZ056Nk28E6Ez3PFziSUAhSVVoo
NJAc8Tyuer/NaahZa09LkqYYyjFMZ4ZGzJBtGD2KNR8yzT4d3fbOOyJGms1OI7XXiB2Ih1bZNK/E
lXkLujSD8g5d79Eq84S8JE+4BeD2vbqZVrp68cPNUlZQwvBiU5tETSEZ/EOzvJvyqFDzCeAOgy7x
L6CmwJWdbKyHvrdLxXgDLyZH/3d0WXo6/bsIwl0U3PtwNK273yxPF8TnYas/tuIeDVxKEtRmgid8
U1aqEOUXeFm32rQqzbgXuNmhU83Sdtqtv42/XLXIb9E0CSW9RuQQ1uNLr4laZhM2Gds8u059d5pL
sdaTjH0G09MkbyWSHwMcYqhgE0FMX8k5rxJdO13UNgaDUVw4tpACa2xFdHykuLpp+9C7AcZPP2pn
zKk1cQ8U0XHL1bLUGWZoy+cLoCdF3UmYt4IFrNEyHGczWPANbEXQGbXItErMw5j7CJJU33thl8Nj
f5aA6DCfddO0TB0lPoO0r0qWSQc8gVi7LVSX6s/NckZI7HG7jGnoxkZigukQbJllV0vfijWh0oSu
AeEwEbgRAkbEcWDv+9uUJL+OOQUrQJMOdH2zLMpUObWITMlj06gqgJJRUlC1CyaOmKBFpUia/arR
ZxL1QEia66t5K4Ikf3+ZSJWOz6Sjly4gcJSzbNCONEafhn313lvCm1AKvtL+mSeG14Xg63COiMA5
Kv5XGVDJwcPRPgJFdCONmeNRM0j1qpOJKVuruSlJUrSPHwf/rK6u69ONKFhsezLXhI4JmcKvMUaW
qGz9hbW5LI25I0/fBeG6jXSaU4qEvcWcANSrkIHFKajJ018IIqGk7eyJEkSZH+/dMcjt3LE68USc
Mn/9kDJZs5h1MMPVJM2xK71RG28/7//2mzAbYMxHfQegBA8NO2BjaFvoRVqlwISCXNyrkwav/vLs
dLBSwO2cpX7zEMFMQdYjGfwjclE6xUMLOoxjw+w2OGblEa8iX9y16Zy0odZv0CIsiBm9a79W3yk7
IzAiUADF0UnMOgydrDA4Tmk049h2ZkeyHLlHg3M97ekg5w48ozVvYDW/dnpRH+/VlllFsprAI22Q
90wODlIDLdiszV2NaAUC5oYTwXR3RCD954BbG9T1SlJjtoznS6p1WPN96vG2kG+TeKGMFk6sBH0a
YtIBvCz03fTOOIOPhmKXo0ZpoiupMcDXV0MEjojEYJtu60u3RrTXHJAbryJcj32wWrNhWx86ZQPn
fIyo9EFQtmBZA28Dx7CkQ+uJzPr/QBMWv6/t4e1B+bZCPL7+S8SzbMwqfyC4bvY1UDv/VUUXXOH7
0L963xSJ6yNjExthRj6rmZu5hzWWuW7v8YpPGiFIAv4hRDbEyTpiq+oVe/+GPOiCsbiON1rsLpKa
rPNAuieJ47yL1HgYX3k21r05bWZhvPGSvxZ1NOSdAinn23hjDPz3hxcs2olZ4mflbC05/GOUfspr
pHbXiYmgZVrv9uIQUA2a8ZMrboBUXldUXoWJVPX/GtmIz5RS0pBVaK4d+l5hx2QofNMuAFh1Fitn
1Fc2pR/oj7f0yg8JQRiRZiC9Dn/czWgB7uPxXlYHT12o/lE3ydHPHmAij6KV6cxaNkbBweNUMTFV
SynqIhX75fNB/+paO8J2TPcBx+RcSGRotVhLvFkrGqKfnG8OQLi7zOblKBBdDmgm7BNn+0sVNbPa
3EkkCefLSY+wNBcfb1Hryg2+H3+KPifSFv/KEm8jI33x0McoSaNWrQuCApsOz2Hfljhr2csjwx8k
FGjAWAY23OXP9nA2umgKienY5dfMERbmN+1pKg/S2sT7HClMIn8W6bEd0+kEnhcN5lJm2GG7lBrb
IUgGW/w4xinStBbG5FXjDJMw5uTirLrEiMQzcMlvYc/8FeryOe+xU8+DgZTTTkkYhiQiV7wwUh48
WTMV8QStN/qHCuqP9cIl4E9Nms9sQSYswtRR7Ih/eeRCS421+1R+71ezEHwbhYHZ4Ro4COhaxPlI
WmkpqPHZkZ2o4Jkf0PbJasIZQKQ+q7lezyci4Vn58p9EJiLQkyygvMvBpNuTWbQ907AGA5dm7+qR
cw0k3g7Z0MHXzsCTj1fCBdM1laFOkh8z/QrYPnG98gjBxM9JusJM/Zj9AhaeffF12wDcTAt9HbEr
YFyfqjCpst6mhUWq1AaN1s14Q8LVtomW9pFd628/ACTcIHajfHWNpzAdcsZOvGcTTAAXQegvQmlV
svcXQYjtd6vGVt0Q5XixeJu1VaWEdFuvHhcQHM9Mb6O3w8O9H1dTKJAck1iQR4t/B0Q0KE5DwtM2
s8gK3nKyaDMgtdZfTJJHnh9MpyKa4clfN+K1L0Pk6keabY9dVmMmfTzfu/Bzu4AMPfVaJgzEaCJZ
NAjwqRyGw26qBvuEqoD76Q9WEO9J7vocskvUvPzTu6o22qxfASlfn/tq7VKYUqU3SEB3yQkUkBby
tXOjXoTunxncEbAsrvhgM+k4uxFxMDUOTW3JqnotXwg1wX+dgyiNFY38V9t7ykjCn0n+6oNg22aa
Wcv3yyGlsWdJeUdwlIs2T8SqEoRQQkeEAiE6KJck6JhJnv2XbOCaShgGC31UdRBaWCdhKiauaQ/z
y7r4YY+e/VlZc83vb1PsawrVD5LW789oailkkYVrFrhF5JkDQRSlVs+cqYxXZH+cF2MOCJgYHt5o
pAL3sLjsmUDr9MeKc8VOZ06/OGtq05rR3Vxbn+ZozgeBifosIbNqptQ3S6fGm+a1QhJNSPP1gR47
q7NESU6/U9nxyHFCABVJwnf9yJ/irtFAewmf7uLQuhzGOMa8rKpPuWIZeMVjuyE1T6Q2qYLQ07WO
s/XN1SGYT/5iBP7WStgYmlwSKpuh1dMazbIMn/WLR0h7Q69Wg/DJvEjqCialsew0XQXkcov91EUY
d6hA7v83qi4PDwcrg8S7pIX5qO+tNdnHVDfxMZ94DwI++3fd833qrjCUpP1s/oiZ/RfbCCAEzXXz
MHk46hDk4ndpy4bnq6YxRTREGZcXY1QvNtj56lbYAnwuN/R9BblaRTbVUOFHiBoJiBuAPArNt62t
mmHRAquZur54mmrsT+b5vPog4Qqg0si47K3ojBZj1VxteoUNzqTV4RYQYpkXICmHQFjVsPsIbeLp
nclvDE5/EuOwIiBv8jKvIiTZ2AbaGij6HS+MRmaAZZTwdxrzsrI6wZCqvsAzrBOyzer/H4zCl5l0
144p8+gEyAFLn++UBoIirrWVrS51cuQYtDxJUMhdH/qrU0jEvTL72w/RAdX1KDNAWu63uzQZrYPd
e5ud59cb4JKwl5RDM4qmILdaBtO/XWZxttvr7H5ZanuXjwZJOzDorghvdN7FhWHXaneoQPEEN1P9
Z14VjB881n1/kSIbub0eA5MN+t8ui0F5InrgnaVL9td3qL8xW0lPGCAGTWtHobBJRSG9yG9Eq/JF
q2wNW+rzzGDUoPZduItEiQay1/eC6LPfK/JfPY04Ench/zlDIHVM59GJHM51VOuaHHp33l/pqu3f
lkRbsaYPhCTHqR8ZdiEJ9l9RaqKU/5jvvcxeGnEqk7g2y7Pba98cGL7qL2WBIafQhS2hNLerLJ3n
KssG78N5Bz1xAN28W00j54452OCC1TJwU3k/59thPzbHS85nrzCUd6VKU9TRzR2tbdEVUshZryn3
WeRjbHTueHZTIUCXqz6sbpIu11f5Ig483KlGfF95SoOGsFVbvZBLjWtjouWjSUslprlMJXIMO/fk
yBftRsssoJjoBNCSELjqwlI8l4SNUoy/I+LbMYRP403daNKTAE0x4Vc/qlPci+mofkgj7QRPmqth
n8uAyooAYHQvj57yub+2d02HGUdkKjy6817EIt21otOm1g/CqBu5oJho7VfxXL6pIO0bsam0kdFy
lqknVjmNf6IvGMtQlErIkkZtuzzGePGwYOIgtnI72b6o38aolZ/RDFAdCGt6Yct0uKSdQzNPwLeY
ArnOp4GaznKa5/wRG/4+e67w9KL5NYltyhs4cx8idOFOZ/uNna31DLMIu6K1eQJh6ujjMDqx9coN
yWhsxU4kRgAzFLBcKdwEqFmna1FuDs1wTny7EeSLT2zo3TzLjtxCDpEXNxY4bnAFg2CaoeryvDCM
3MUCdBx/yp64Nmrq3qlunBkgbhyY6GaYun5ZlL7tJKxr+yiqpnAwnGF9iUgm55j6nfbKT7GfqURQ
m7pqFq18r2C7pMP6gh6ww04D6d/yOIH13Fx+OFAv2uNSBWTLRKsy6G5rFvHA/h1mjhvvoQ7SEsT6
9Y85B/mLxAhrJ3g9vqnwd30e7shHdKn+4oIHVTsw2TSM8W/7bFOLA+3WZXkjVbllbAOvnzXL1reL
ugPIubM/Jj1Y2mwkHjjeRoEfWPx3BmTI9MLIuJ6bk8p0kDle5QAQZpftUKF54syYzDhOiS/obtxN
+8KHcwU3FRbioCtGUJdRw/4yyitpIVZd1YJ+m2P38qUmodp4kMIxjKuS1wNqKd8FF2A6+RNMHso4
FI8SEzjP3Razvif0g8ivxyOHVoapuWw0fgDYaNkN3OI744ez2XfRBjfBnT97s8akUhrcbpZU+Gm/
xPIacUsOsemZtRgOhzWMMa3Z3S5rsqDBfhUcUOvagnkMSKca/asT+tEaz/u46jlliv5qswLQbDdI
HA3vONxKd2xI8NgiuFpbQ0GDmx2t7tu9a1XOKS8DGD9zQWoxTGaknpPqTf5dhuFVJCLUr3TegF7t
yVX9RZTD6YlUX2SchylOHgccomUfwE1pfYa3sxu2ots5Yi6UNV3ROjl2KalH7b/srmfOxjM/TWpF
Nn1Hs8Pc4cckCAu99JZY0ThN3Ppm/X854/HNDO4j77npu6sfxGNBOOYhDcuM3NZCDv5gg5Jpqh3n
J6X597UXKOvbkHyGoYpzUsXO0cbVE+ynRca4tljLWMFt+92WErwnYl6hDL922UcSS5f9DwWO9TNh
Ir4tplNzpLP9on3FimV7+2EHUSNUvXD6ZkhH0b8ka0M4NSGH2W5ApLnwvgKrud/VmcqEGAp0GcSX
4oSMH6ROBVzRHIXo2GBryL/eqGe51yAjKbntJXuiWA08jL1CYSj1CgYuWMAe9wQ7Qpx/dX0qwyp1
jjrcEWOkNvATyd9PfaYh6v00V59ZIQ++7p62u0bTA1Nwvihy9aq4t/uJ1ZU+4YRV2WzhhazabhJL
KrVZZ2Tf2UyRZkspbUJzAkbqLNbUru9LzObrVpKacJi8lsiuRIJfYCclk3R5kvZXZXuIVnVDlz7I
IK0toW4kec9MOyjUrD2eCIqAFVL7UR2ppWh2EJYaJUyy8lDHaj+bhV8uGOqqT0KAqXPMzh6XiaCy
kwOYVgfMokdW3dPO2hKqsofzhFjBGs51j2Eo54yS9LkBHV0kPpXIgMpcBUS7a4KkMbcK6x0Xk7Xu
Cj24BP3Jpc2Vf++z4FdF6qfHTsGxc/ds9G6jz38A2Bfg4zAlJYAHNXG6F5X0IWDd8eh4R5zCvUST
DXt0EeSVgC9ZMA0ZiVqEcf758XqsfcC8cSLNr69wjkN/6neLI9sGi3IvnSTUm+n7VYEdqBMF7whN
RELRi8cMQCK3ZymSarxp77UYSmDekmZMz8psgWkt6nFjRt77eKc18bPE7F7eKglM7KlRKSfPbF0/
3nACTkTiSRDMrS9ZtNn+Om7EEuXaWCXr/Zn/QYwWIS013dt/NpKNFsEJ3BZD06c6XSMCM9r0XGrE
td0BidNybyhD3PI/2U5xc4PcRCm7lE2lHEgCYI0Sh9dVzc6aIGjLzWfbfVPZfR1Ksqu1JckbjbOI
plUz/8ZoKnmqNByoEo4TL/DUl9dwa+GzsdJCtzylPjgLWSbR8H7XNV3nvPQPnjheqeKfXZaLIHzN
C9n9rPuZsGQANQL1qfgM/NHfU5m4hIwz82rLflo/vbDfqOkPxA7o1j9zJ3GjPn56iddl+djiXI4T
ePP6WXJotXSKdNR6BFMz2B5KsG95MYKEiQt4fsP2c/U38sMU5veRO9PgeCqfvUTtToMsGWvGYH+u
sR1103x+ny8yTq+0267VLr/2v/NZF/uI5UR8l9PQp5+I/1xE40YXDevZlVbGWJQjRT58s+kMOGAr
IjKV6Jyap3erUVckFqKkSqYVFO394EIGC4hkuWx5m6qto5UdLUN/OeUU+MNNr0isAXaVZvnb3aRD
0lpCW8AqAF+S7fbuPFxoFseqQOmvFzxot4bgQxVPZ+9bH3isoBMHasI96+4PZfSNbYB9dHfuLi7h
jpElhQkSNjpvPEIL64rMqEr2oF9YOibzNxa9+3n/i49PKUUHq5MLcma6rhw5iy/n3XxJStxcnUNl
/geS4QIeVF91ZzLRQvRfMOCBdtuPVxrHkn8U6xVSA0GNhRIJWGbpC8VT/eEB5Ygg5urhclLtJvzK
biPHlMxRETBOdidCdqynPy344MXe6EnUxKBS5lFSLLGoAiBE988J3eSF3G2OnSmGKpSIiAJ009oW
TqO+O5xIxxYqy66vLNRD5c11n0DI65HROBJrxWO8+Fqo4NZpxlT3xzUnQUCIDUkU2su1XXfLSs8m
ZHiow2tuOxc9ky9yh/Um9FXejmeCycNQzE/Zb0VUQxFdLiqLS6nYXelPm4bXfQr9546MhPXMJ56d
O+6tSE8zrZxdB/gL837Jh+q1Y9/KMSBS3d9oMNDTwVG5ryCo0uqypCJKYCpoLXFaDdpEA7kAu4J9
8O8I3gruw35KPXGgc+B/y1o+lBN5bRUH8jdztX3lCYAvNVArh+yeP2wggAA76Npf7svJ6C2jOnsF
zb3BSnUiVengHGpT1uAlI4BNoZO4ppf3/mOIqcl1gODtaS6wZoSb/+cZQ71RarnaPPOXok1218Wv
xshBKHwPe63/rtbuU9NOIORn6NKTdyr4aBbDJdS0bb04Xzzqy84WODCks6Eavp3qjK7f6yLmuXcw
Vg90KpOvrAJpdG3rlQuO5lB5x0EiXIh5Ivm7sRoNQ3bRXoeag8Uva9eF4XssVZEtonFKXHDDBU2u
VgUKW4j4TZmiSaGUpE80Ryuyz9wZXHO96CXh5QDiLvF5L0EU7cNJ7uMCJCebeQC6vjvQAqLcgOae
fMjPlpmU07fvDwujsKGbJ8bQF+hmfXHlBpVfW4+DwYvB1Z1xI2v08kYAqa5lAegfUjnkUB55IUZJ
CSjCLjdb5R7uK5aDUbHJXoQGPHLCIxpMVbcJXuoSzNHHjLbgrCkTsm19ayXWjaoTL6MBJIH1tkdo
8lg1maPszpy9kS4O7U+v14EpCHFBSrLOA6/ZV/IhxhH5W7hMZxPw25KT4tGxNKbS/AoFWWO2Z8Kg
NDPv+2JZt+Vb99iduN8Ny+FxFvb0d52PE4mxaC3xu91RAqe4QpvjVuvxexqoVYyIf+MJatOWw6H7
lachnOD2S0C68DeGV4qaaTW7l7MHTIjXenHnvL0RUdDMJHXm9otjG2EHGEgdzvetF9B1RQB8Xf6V
X8S7BHHerb7EbrqKHDaYcwpGU7/uuQ5CpXo70sCQlprNBgNR1r8QkrJG9rPyn+qkCBM0K6wPPNKE
Y0H0tn6kzL4NQLEYN6AKQ1RmyeVY9aH13wMa5ZaBC5pWVNMq45xvQlUr1pFNi2Cqw9dafwUpd6Qu
l78ls4h027rRbdkAJwvX3tmEa/S3ehlbu7zzc/nqzKFSJp7A4BLfgyqLqhove5NAXZXfa6JEQpSR
bhhreHjf6Lt1kdEWFzDZ11EqX/IzLMOZ4oU2X6rCha7Z+h/tw86xUJ6acAarWZ+cJGzRt8ZMFcyE
lXQdmDSD5JjPeDqjhHpDmyQWTXdLabrq3QKac4Ul/m5wsLuGdJIlwV5Zq7l3MvzG9sszLFlBbgMO
C7EkBziCnRiDPdOtFOBnfXcwnL5UWWb+so2DGObP3sGPvvyaoQkKvqipmni/PUb3HBvzbfGk97Cf
NyY36TJRIbDoRzQuTj5TIGKTZoIl1dX3erylYx2NRCf3XIxNmuHG15BGBaX71f0eB8WMXRXHMhcq
V3uSXAkk5Sgguxt4RY5GvklLNjmNAi9fsL8j3ErBC8EWAaGN2h734b1zBpN/qlpXMDzBhNjBBgY3
XBWuPdYomF2tDl+xIvEWAOSm5h6QiyjPbUvmb/FZYo5Ts851h0DhKVMUeo2UcqcexnaF62buTAVD
4C7bY2bHDscq3z5zDEQe4985PlqHqC827pYd0Qq9jRPGZUR4cTLTkiBv+J/wzPvQ8GinH+P/JVq+
BjssVNpb7sYW3txBiKThvW/Aqm8Roafn+5JEFGvZb0W9RZniNBeeSWxIAYSmXLFeb1oTidnbfs3J
ockjJye0AwfBWpH78Y+q38WWq+GUpCbTpHvauygHQIqDnRPiTy8Gy+6MrMn1PpjVtmEMc2YkxhQX
foPmzDFo2DWc5lZ61GF07fpf4NwquVvSwbmfCRKy3Auo8SxFGpdF+y+QOSdGkQrF2M6rreHs4uD4
nx2x4RqhqMzgMYgl7LzGmcizwiU5wXl8V32TVg7Qfdqbp3KuwF/QTo9J9usfFxjETLLBFxDrSl4f
FxfJdqrX61oPWL2F2TodaiCkvSEBk+cCXqfEnMK/lu5FvzY+tF1mFyKXbcRDqhCdz6raLFGjfcp2
JVvjA57nqporVN9zeeq8b1q/l7GbdkOfEgr5Tp1eiraEY9gNcMd4kROazxgKNUIGh8QTYn4aB1I5
9jeHNB0gFd7HcPbmgICNR0lhufZGu2AiqQGGiS1sLdr9ZlnqXRx5dt0j54Uf23WSkzK5kQp72Fb7
VuSwv+jZNnAMNz3Mzd282Qj9SBYuGR2xDnNExJQYlBoE1gEXvDNKnczE2UqstB3fzAZeV+blrFSK
2pmJON99gRzMjKHuD1Ud03jOk3BvToDQ2ymUo6vHHU1mU57PCvhVjxaJHtj+F8CO2LwrQCAgmxw7
7xR4YjEhkYYEO8WdS8WsauGbclUJ6hFAAnVty4OzHyBbyEmSESuje/Ll4fDW4a5HUcbswIMiUWja
rfhxY1bBkKhrvyuUbxWqLAv3qgUOOGfuea2p//I1LLEZKkfaLpaFvigZVD8uYliOnaRzymLVeuN2
y08qp/s1TI0VdHlyvsvPHb4xJ1TMKZMGUYS6Msafz4xPVKvNxf58zF1a3uli1h4J/qWe42LebVdp
otuoB5ciQMT937XEVEg9XQIFdn249adhgUvVL4mg1b41R3UxcwzdhUvfRxfFACXZPa6rN+CmYSbd
+iSKBuEGJbDh5h1doGVBU+Rj8gpGJk0PC5Wcai69Ukl7grOU3vfUMvg2azh7kHfXdRRMX60NTxAf
U3aZVH++LY0y9xb6glTegnVfYlA5/b1/mSPh26ZnbDGH/E0EurDRLWz6VVB+evJgc0kW0ezh2IMD
MR+lifTfXkIOQGdlXCyw9TWsafOwXof7yX6IfDn4zPeOtMPEyYfTY4p4nE1RkH6bc8C0/D1IUMfY
w0ljFr+ub27uXJMbFeQK01CsfdMBJECBu481KacJMLFMlKyGbM2EDCVh1+JKpXS77H852uQt7n8a
kBdSj4bhg5PVwkNPz8ucCw7ARpHPWuwrOFLd7RT2jEoz74fuDEfkmfCHY//e6EXMIH/EiX5GALwS
Py9E//CCoqEeuUuIuJI7uLqg+x6lvNLAh7i4MKgfaLY+HFaWshQN7pTgp0J2Xn+IKsLj27Xe0Zdi
J+pituldOSjdxhJ+jbisSQytzrz8emIGQuuvgrLR9ocd792cGXGN4wCjiT/nrqU6LYgLTOiLWWE7
16A2ia3CNiO+Ll6Kwr8EztIZtjbY9I6Zrjc0RSoGdZG7emiFNf++WrtBVh2giY5bQnzYIaaWna0C
cjAAtTeNduoUNoe7KqlsLjQoJGEyTRWMHAX8hhrAWLvDLGBg5NJHXfqOGVE+/HgJ6FtycDhqwQ5n
4jWdisV5oizToorbJucnzWguN31JxFte0wRG6saD/XKCGagCgwzjEmW+uaKe17/27aQkC2ss8mBB
6pu/cPwoVRxnTnvu7+8QuuvR/lDH1aB4kA7DO5Fa/+yrkep4FTRmKxDOdpjrTxAZWijx78oHyJj4
2KfhChATF10nsStkI0VVKyZoIUPUqWqNZVXhS95cI9UJ+yZzx9yReF9Fg+uErZ/SsG5DTtWwPQOt
WzNLzxrkvatck/jG+3v5AoOyRVzz6Aloo/e0b8P1qhMl8p/fn+ShdbVFVLy0YuOjlc3JgCgMk3A1
tTVZqrMm1a8ABjfPNCMCHmWSC6hzqRgc/F8uyWPLUNyqw7MGD8qtv1aijbWNMCLTQTaKdjd0LeAF
W2Qyfw5879MzQqxkWjDhNdDMurIPaV6JFj0PAJpe8uEBJ/wD80QFSfyq6kWL99BMTIvWWbRYYM9x
xqJTw2WR6eRE53B0k/6heRynNywytl8xdcQ2hCLVyCkn1nJM2sKT/YNmyIKJVAnIRhbpOY4msdRc
olp9YD+BwukV6OwtL7f1ci+IMUjaNxDslZ753oZYgI6qKrylXdSE5NYngE1qZv1vqdVD9oYr38Vl
qiUxtTXBv7SEUzLSMNngQbnb0UxV/xfWKykrRe8+s+u/3H0VAN1fOstcjroyGy5eaqHGkC1w9YDB
iCe76eYLDONXC4j4FV2YnS+mOnRRZBxw7EJi9fYevoKNiED9JBk41AD0EowisZWLIzNnjE+kVAE/
KikaWTvvNl93fTVQkDoNxJoO44uHhnIRH4+9poglMdYoz2+vaU22WDui4iO1LK+RzB3hjcjzl9CR
vrwALmg2Iak2sAiTuwHjOWxpJwiVwjC83gUL8t0N4FJSLNAMA65ixWUpK+TjThV5Pqi1+g0KHZ9U
DlfWOtc0lWpxKmDkX9kIvKfLkzOMEwWz8b5tMmqZpZk0vRko+kZd7zC2gxX3WzU8/OMKnKLKf1lF
qK6jJnCXARUJfTSKITiExaY9o1GqBKkZ2XLIUXGD0C1Js4swpS1b7HZZMhbNldCLOyvc6cv/po1I
3rjHbGwETuCF4/CcgWzRE4FjMxUlpjbj+A3OTY48eSdoIWOriBrx2g8mQgLosuvkRcsIQ0xeE9SW
r5Afe+AP3ffTQhfKKH6vedfovfPY0IoSVOHiQCNDFO+0ufvWun+rsCS2H7zP8YK6yUmFk8SNIhVz
u1gxva/jRBwFWVek2QlIN0I2FodO+PCsSEvL0jSKK9ygADXLJ9koRr1fd3lDYjR97xgFzSGMCmJM
miE/tKnwvBW8kYbueockNb2h+r39u6PLEI+vly2+pWtlg7uFVP01F9Jt9kC40/6csasxwQHEMoeU
4z9cwHDc9mB2Uxc/+0eqRhhYOrmtFQBaeuRHOxEarV7Du/fCrE3+2P1ycIyx+H4NqQJY2wdd6pck
aVM6ANBN2DZvzc6IIUVTNKEF0wuF8BXnZvxe3Ko6IiUnuLw4mIwT57TIRueFU04E6AI7i5LfLWfU
nhMBFZ7vQu7bie1bncmVgoe2A5YRuXzxgKltg0JYlN7bhHZx7rNr+vhU/4/LP9WzXp+/GiBple3Y
KFubLKYPpVcszs9fL8eV149CvRAxv48MHD3vbepQxaca9Jy7e5Un2II7IKxPmVR4f3LZYXneU3X5
Rsw/2LST+JUrafwlGGfGoFlOkejgHZ3E6PKsgZQ+0N6iSj7niQ9jONLZfRShIcOtgiHtsqdJEZzy
OYtXJiYjR8RKWH3zovz0R4jJ19P4TLkFtiNPT/iAFYKMusXno52hAk4mI9HlhMANPqM7qiU/cqip
DAZirjMV9RMO/wYhhOTKQf1AnmsUDBjCy8BeqwircUYt03cyh18WcJoN6j1x8R3ALsXSfsRGZHcH
bMoL7fh3ZvkP2cu+iV4+SRhNhoRQH/W+YtJ3O5uCHvw9ZVMEpgUwSU29yDQGf9xiIBme/yjnE4tx
0T/jpEtSpLZ82Bd9le0B4p36p1Il2MgD+FqNiLjQVSQq19K6ua24vNc6r8yVDoPTKJEWlU/wLnFv
aFyvzfPuQFwqKsCveSlrq1iz3pX++Y36scbYkwXgqRSk1r5acc+z3qZVfD8/R9N7nzTEb9oHhqOe
Xjv+d9D1BnHzZHrk0cIEz16/kJE/DkWjIjz9nmF2Tl+coUVro6PPzbA82jNWj5XkuGuWtIB7XQWZ
z9LrfuLOWjqLuRm/huVQIdyboYv5xtTQ5d24fcZokKgMVcKVgrE7omWGuScxel+FGVJyIy6ezJKe
45bo1UYutInqH82KNYOGFtei3EIiTXpmI9VVfcZKlBpNhIpTeTm1d067+9yqXFJPy6aOOVVGufsB
QYdUyGId46140yHTpmt9hVwJqIVJABqs1q64rtrDGZdD6vXSmEvbCdFzgVE6G6cEQgXDJRUvvi/r
PS2OQVejaMQ80QRG+ft+h5pL7qRSuZvZ/lK4UuLwwlcQnrwymAmTipjPWPuJoTeNDl3fVwYHEaDd
IW3SA7BAhvyu5ox0li0V3jATP1ljCX3Bbdk0idKZL/1yyYhG4r77446Uh88kt00dc3zFgKdcmCZt
903ihlFghkPBdYQvOVckHKnm/Hhi8JviKLPhfzTijfBav4DyDID4nZQ3SujVffydCGkrf5RBAjdw
xqHxyNG0868no+uzDAkjw8ljbgX0U4Nd533cjcjSbh9Sv6iJSe55zhfVDVLn+oqhbGitDZ/ayOMg
95BcPbxSQX6ZkwvhguSHv27O3xD0oU+2CcuPYFD+mR/icGUM0HyYBHDQjXbIQl1U7dXybYm+HEg5
TygNIFILzg6q3JkLPmqNhmX+XpotK9qWxQ+kUaHciTIda6B+dcYBsXiKygTNh0NIcU1WItcs1r7P
RbU8T9txPT6o+jXoT7W4wO79Pf99MPTNwjZoQ4nfdUksGaYDJ/vixGZTHmh7VI5X0MBuSwuH7+wW
i2Ufv+c/Kf4uqXEVlte8AW4mR/f0fy7mieeiTqc1gfcq/MzzLan4SaDd8Z6rHwDNBr+lF+ERRrld
R0vL+IKvZsikszdhREGQcUKECrCjVbOUg+YkAFQCiXrdyBiwX/U4N3IO9x+pYsdwCbgMEsZ+qIBV
GNc2aBq/rF1X8B6eUJjvBLIe4xDYPcZsaC8euHa2JfU+mv1OLaovJdIhLlG2bTIziQ7L9lBgZGU0
Brl8SGEZ9SwvPoxv/jYnI4rejua6lznVOEKG/Zn6qNcxINbf9XSpB4ZrRXha/t2I+SOQfq1DAMT9
Pdu0aknWOG9onEjSv9ShGejHwFvKRevyTfVRaaXrM2xB2pFjbJ+9VQoJJX82KRHQxiHzAk7gnZzk
8jML2qyOShUWFEdyzQ6UEKThuRD5Jnu63KidoHtcDzmzqft9cLnMUAV2W7d92iMUP6DaPF1cgLLz
kPF9FAdon+dRovVODWYmfpnYs7alcZ7s1DVZcYAaNZaKs6FXVCcVNLuzT+Vt6yGf0tZ7PFMzofzl
6xzZ1ldzsicZsW9bQBgw6+uf08vbbYcMIMhbEaNnmInVvPpzl9Uglsi/w52TLX8xw96RR+X6Odsc
7u5KR6M93A1g/MA5o9OnL3nY0Lf6MZTHCf9IbQrOAUJ1BltQUQOhi3HmhNVi8uCj0NT0hrzQoInt
A0nGENEWin4VnMFmuKFTMBBBPsw+uDyFZL/jsNy/ct6zG7LDTkGBSxG+2G4qXVd9wWoihdOZKwky
yI656SawNQ0FbcPCq9sjfpekQs9m5HDAdMoeV3sP0l2lXDsxhMuvDsNGPwhrKXQ4OT3xT4fT1aQP
r1dKVZ0MPPgIxLo5Al+lsL903W7VqjkzsnZ4dHH968C+CGvFm63Uyc8JjXNUzjo9Y3nPG4OuaaCQ
bdGNNbRF8NCt0ptoK3wTnk7iupZV8MijyBWEG+7Sd6suRZ/hhj6BnxlJqjNo4yeGmfawKL4JWSQ0
zTM0tyNW0jEcczaKcm2TgjdlW4zqUCNSbhnA+F70csYo+tUoRO0ydj/6TvW54M6QgZUPuGSOFOa4
XqDPJNghTEANYeo9jPf8+W8vJlXnPfeDFj0+kE3EyF/Gxo/+X+SkFE1b4iZdG/7Szf/TBeT61CGy
yRRolyyQEJ+6QDJiGaNs9gyf5IN9iSt0dnsgyIx0TEZ9LnIXGP8m/w0DaqsVezOBvEDrTl3szhrh
2tnkJ/ZpENNiAwll8J3hqJ361+CTciBnA5gZLDntQCwYfaMyOW/fPDpMhaaEf5sXwloWqHhHNlt4
7RqEEQ0bm5DHTcQQPJZDyJa2b1Lm7SFIVUfAy7t+NX5PgZYu9rMOejBB5CetRfjd4A9S+2BjDuaJ
tqq8A+lz8KrnysqXEqNly8NNfwMF4LwrkrXk785bjjaiycEDlyqgRCj/xJ2k/efKlS+/C70M+Rhv
7wopzDpCm5heyygJoVMv+fyC509c8Gz29RpW1xqBjZcin6Jdw39QWv9l1bJL9diAEv3tB9Ln2aV4
53Zrxq6h7JUXQA86X+hFBmI/u+RvWwUpH5qG2ZUjdvEeRFao1va4trB+9MM0rRaLzIO2hHssLYDg
rVk+v1XC2J37C4CQHTlC8S5pxdlHITH61m6TV+VTlNH92uWaJ7nLuzJReP3SCYHEoPvU+zYpKWMN
ANl22c84qjR68Fj6IpjWWQcfdYOuau6i3pmZzXw6PHCML3TpSaSH8s7vUVrN+4oLBzdKXyoY2qYZ
NE+0vV/ASZYw5qXw7D7xS5eviBOZtEacJY52lotALsf0rS0pqGC0xA/538qVXyzEHG6xd8Bw0UdH
oqEUKyBVg3JBTg5tGDL+RtVY4bq/k4w8YmEroFHJKjhar2P/qr7NiMog2gp9TUt35sz33pY666Nc
hJQLg8QXKND3ZcurQq68y3tkc5I6DYC1zgu5kHNm7scw/QKtTGXbndwDb8tfO3DkPLKQXz7XrB4L
aNDDmbuICUIRmuztY7qH5mp0seb3+seHcSt7GY8ilchzeLut5qvz7iYp/YrAO7Fhs7BRIYLCuKQO
F3izaGzQ6YlV+zb9J2NPhJDB4kFC7op5n0IOkux0GZdhmbWEX26s4UUvwcKxSMFqSBAbotr2l+g6
VMYcb+OuxVZFKE3N97IFJ/ApEsDWh+9Q/hioxS47HZl3kCc2Pn4fIDKwYwaou9sX8Ey3xeMucvsT
j/Y1JS5aQqI0mkQ3A4evqWlN5Wv7a1Y+uiN+Eih/WMtzmrOcHp0ksMeIzlJylf/j9FgRuNNGDAiq
q/SSa1Joio3dLtVif4UapqeDrBJFb7pJgB5lOQmKys2r3oyHrxGmkaQde5fVaIf37ckhi3ou/GPo
flLrakpz0lX4VyXSZUFd/F1DAlrbl2OAZPuVbmv/fbONHsV1t9rTfarH5njgM7XwY/Ytss2QBD/N
F40JRdqeMKBlUIL8Pxip72p/BI++HA2uWP319yubiqv7zraUbksDqK6ckLBSbMqP758+iB6aTWsd
ynCrAFEgOUd5B6Q77IAN9BYt40wlPvkvIUVnVFHMTq03qQeXIx3vl6B7t96OkpbXBdG2p7fCoZvc
eOZ7iDjzXzFtN9areneeRZxrOXgz3idXMzOrssssF8oY0vKp191xaWy8CSia9dGPc+KEYzUiaC/Z
XiyhJpJAit0JL5tKnnfw8iFud833WNyfJLy9VRVVzeKi7GjqRZ9GOnkPNqz/Hjrun4YuVNT5reS/
ozyADXTqoqSoBzy36AhI5IDrjVeFlAu+poRE1PRk3OWOTRWT8indyxZf3TP5qhbiUkw1kzaMN9XG
77SNMgroTAFAyEsh7PheUO9G8hUJSbT6wmXM8aPIlS1mhfB2Zyhl5irkAHIOCUqrI/V12gcc7cbU
CzxIYgHYMM6g4dlTSKxEwwLDZUXs8pUaUUT+mo/UxMNijewaTd/qpZC8csnU9CDIcrAEdwlHJjAu
6Vbl2tliX2X5XpMsHvuv3fQUNLyCgyo6S5403vA8SdlW+hVJid2LCkNfFxcPwFdzozxW6xJCxg1j
XF73nZkMR4vTj07Mb4Fkt9+OtNIEm2nPyUyMqlwH4fss7sLn8pr3Rp0alVjFnsb0ZXYR0R3pGDev
dgqLfmLiY87ihj297shGyrtt+njXjTwhaFkVyOSgytlhic9szWWEGsUAeesXcqUlH9n/ZCvbldId
Ag4Ht6udhfVd/Kl546NmFUom7PcLFMB2ISNuwz9/ixA9OqKkcnrqdKQ+XnRm+Z4Ae/hNT46bMWuG
TG9NGAlAPnYtLRGtlv7uEilZMX/Ta+CGxqpr1FN+1csuzVAPG1o3kfrNV5BMcraN9PUhKubOCgMs
gtRjWf0bf12Qy+xbTWE3VdBTAuQR4KVVaFyxOeuiF7S32NpmjKNt03pGkZTq+d7wITmB4PW7r2dq
Qq72jNECElR9vBoiN3lvfnpomGr9ZsSFKiIHVg3OjkA5RSVc97HwrGETWgKUTV1JD/MsPXlIy6vR
Yb7LvrKTCf65EAhdgTGszG0eteVj8QSmPh4moSLExUulfMX55SE1r5k/6gjWD6ZB4A0drQU6pdas
UAzzZOfSh2QGXHGUr3zMxWP1zhvHFGkTERMEXpLJZEXtxtvFw19dIWoY7hzZczWRkXWd7H6UF42n
ZU3vTjYtrpuhQ9/CX6ETEM5UVPjDJ0WftbaPeiMKXPtLGgKFsg9PLzZYew/yE6kzXCthkxM92Nvr
RNKmQxwvozf0zH7Ak3gs2mgcpKm/mWAUNRXqPfupYKqRqzoT4YQyJJW15jIP0tB97MCxyqK7QvCB
zTJW2fc7R0zSG6wbpBQsPFmomr9LCP0b5u1NUnZoG63seha/6qBoPurF1ofHti+u1S/8sc/mKE3j
bASEwxVt/QODemO93gROMGTyxFyZEnYtTyYTHIRDORfcm78g+hfP9yFVBV/i9fC7stKcAo0vk5/B
abrqeCGc/nEPbbFGMp6nZHOfpgW2TbZZM/A+UaT7+EXSDk4p1Qzx+UKGDw6e8++bincSKaURBl+/
Y1DcSbF+RFVK/G3hPBgUExkDiTkoXNL9PgRUh/tiHrkYOrrMF6OdJN6uB3Q/UJmJYDQGThfuuSFR
KST47NXb4ru2vMjuC1Oa2P2EobGRTTx5hjoE3dmOICbV4MhbbAyYuh/HhyZRvgJ6dE+v/lmL//H+
P7ini7yjVaAKyfpHU32AwrcPJlJIUMDM2q2Lmy2OEn30WkVk1L3IOLtMewNWrkf+nIwUV9yLh/Ej
U9nsVsbIr9QfScO//ufk0fCdUnnNLBbcEdQNK90hRAgfcJWBSS/x4KLN1//mYyHL+O3drtmMi+tL
ts2TWgYcl+cIArC1BWj3T1qgAwmyR0p9R/9a1omVW79j21Y3s7/8Yg01coG2Q2IXUkLWecg3d/aW
LDWSVVo2uaFjZXiIHHbwv53clNEUSx51HLx40sg7QRoRr4JhsDqn165DAqMFauM7KgUN7uY4R9ok
HdhleSZoAZSMLL2JYUg7rfLLS6eoQvOByy+L2DE9SuJMGK+iVIzSRUFJsNcCTrOJNTNwm3WeEqUg
GPbfGv/6O51CXqq9crL8vIhQFrKQ8lmOV7ZSVabh8E65ybu49rl5MEOFhcQBwdwCoWA95Uln02Vb
2ch/6ymyE4s0rQJDIvgxjVjX390i7GT1yN/K+40DKq4BRSESfXmAepPCZIIRPcXWNyJsGbfgKcwJ
Y0PSadJbjd3eR4Wc6Epzyi6MZAlKpSAJDvHLrEQ1lVkUf+VPVX+b13NuIqC6tdeoo0a2RkMcpL0l
UmKoDxK12NPmejHI/4nvWnyPzwQULWxIB2gXJwDzNYMHfhedE/UVbnSHwrj09OQklidEo8+MtiDW
nUO7GXAXr2FSIxlTRS2wUKFFv0xRHWZhCYY6iSOWMdwLz1JJ9v+7g7P1v4VebCAiqk5xOItxHkXr
fLUS9UTkswRpw9DhV69UJn1wthWYtT4RAcm65D049s62248qeuT1cqhvKYyuhEe5easF7sO8rYsN
OsJsVgJK5GCX4NUhjqStvbqT3PRBI/CWinLbfLe2+/lCuIzMbXsmKRAaeiLDD7xTHBNezkYo15Kj
C9L4hlmTYz86lSfARpCdTBW+lfS615WLMMSGalKVbSipYJERVG0vmFtIiK1QuMV9boMt2bmH+vhB
bpz/icwAs+aeRaZOO3waZ5LizsOmy0t2sJqi5yvTGTQqF++yA9yV8Tm0ELChWvmUrlysBaZUHAD3
kme4hcV0jGPgyDxjCXWXLWGlig9Od9dko9Whvh9U1khby2LiXZEKPEQgOdbk+FItPHQ+6W9f73Oi
O00vJSWxPGICgeQGaxZnYGdA4Rp7QqLa4u8cmCACk+gVBK5tcKBtyc+7fN7TRtB8Ch557SlavlkV
kzmS8SWLElNgiA2DdbZc73z2lOIqQ9FmYai9fWoFWOXtBXJGhjYB2eoC6LxtBD+ZivmJ0HFYeXZx
bYejEmu+N0uJ3w3WxXlkJ4BoQd1iJpFqrdOIDYBDnxv7r8TMsX210c5eZVcXdaWYTpTwidJKdN4I
d0a+7KHRxNtyCvvdj9RazxuRMxUHqABQ4YExUWbr4PQ1hRhgYfJ7pAb8Yu5jr6MVqXakN7Omg8Z6
DOd61xrnVjAatvtXrBZlFosc1140IjfP4l0Fx82n5k0e09i8OBYZzWum6qDHKo2Et7lKbzwxcW45
cvlOlrrekqzZ/UU47uf8W/iYEG0pZnaVEU5xr7MOCoOADO5MxrQ71RM5Y5DAR6Q8bcwhOrdLCj0o
c4zQddJUGti7e0BgGjoPf+g7AerRPvoOlWjB2wy107+pKVz3Lbtb/Dh3y3dFbE3OoVjAkcgjsh1z
o258NmU/5lwlhBgqoe7uSZtQbH6juewaklIhca5k/v3f2BFC4SsRldHGN4WuvGrYY0fomDTucIsZ
wTJwgTlZfUc/PtMu5iS4Gne7DVfJN7OzO16F5vaPg9/xQfKFj05sIemigrNjcSOf9BsoH4T18TS4
bMj9Jn2OafNJFacZ4Ws7IRWJt76Sr3QSlq6z+IzsSE7i/EkOwh/SEHgYPeBcwEw8x4fniChizxq5
P/yITCNPm5EWL3twIisgeURBgHucrePINjQye3Xx33ZopHcaSgOHkDgOb4KOXFDu7XI7R2uU891B
dhjhRdh03+YWwPSGm26YjnbywjNjFZCxzy+hbkPUjvCpce5jgo9Dffhqew6ZuybiAeICF+pmzIjo
CJzWMXgYLMCuASo4Ey9kOGNxNBIsFrhE1F6RIecmKlAqCX+Yo34SrT+Qyn0s47atG/wCLAb+/wNK
UE8jarOsnsExrH4xL7adsQ09tqX3tikXkUt4iGM031BMmQF71s1o7m94i/gHfGjuCf4qNIWG31gy
G1M21ikQA/aiq/O0nvY7wwGTaz7H7YbUGDKCPIZPnCuTBBmpOM526HVzFnk98ajzkY1O1uf98L7R
8Z8+0DCH+a2aZNYo2JpInq2Gr0MXEOb9ULjWliiDv9xgoFjTVFhmAEiIDEDV9UCwEZGENEarVtLv
0m3BnZzyetKIjbkIDktkTlzmSmLni0TM6AZWbPY0Yd/ssEjWfJl28YItZT+v2ogFXbI09k06Av+j
Mo2ddiKWgyB2yYF+h8qFZliZ3z/2eCXvfV3nI8brdKWfie7Vj0RIWXjnEICZEfjnLmumsPigcg2K
HPrSr/zWSBwzYVPM7z5x8ioWXBO2d7tOi9eYKM+1Z1s6rp6lEPilfUZQI8mCJlbQ80bOg9lB3huC
LzPBC+W2SmZH2mrco8vx5qpjVu4g7nXL8SGI4RqacbpmJUMrtUODxcr9r9X3q5EHLWmPSR84JMlc
rIm1fHqUJh6jI3Yjud9mcrRLzHG/H5p7jMXLbSuclDeXUAc/mubI0boH9HuzrJH/RxTb10YNWUr+
GUTqX7oRmtWUqbQRdeLboxJXvgq3haVq4ye6CbOw3UaytNrqqZg/gBqVTy7rJztX91J3kjLREcsg
cX94mQKtSTE5MQnLnazLsDUMS4zWULN7Ex3syfIXv+rrMfS+zSpTeik00bCC/cirEDx2zbJZ8MZT
7p76CeCdC/ahjY3VK+mEyWBC4Pq2AU1kspgVUfP+C48tJr48YcSNzCYgNJbwuQVeZd3iHMnBp2ae
//K4tLsMSqseFYBUFaI9AZT0rMTHvYsariTYbzlfonO/3NBB5E/zsoxsqh6/lStxZR04CaaDZJ4S
sEa0CmFasMFYFhRcXm5IbdB9D4BaKzDhGoUizGwQgTQMmQubqUwLWFQy5i2GxrKpDgKod31eo9V9
/wAxad6ea7gDoYMxb5A4Ew788uvzOXK1Mf6G4JopBHYTPLZCTWX7agZnTploYpuqciWGJI5+qaGg
L6SVr7EM5XrF+ELKG44pGzwU6gcgDxj7g2xVbm16GQYB3UaiJXvGcBk5nYLpJtzEYN2twOVWyVVA
Rb/emYMRUO1jliusbEakt+uJLJdrcKYdKn+WYxyBlN65vWs/ODFW08rHhH3XaHT3ZebfJ7LZYaIm
+SMCxVoi75Lxu36ApFvm9GhdExiGJX436K1Bbnz0ShzvMhrDv5uyxMCE5zHTlXd9+bcLBf8ccKfj
uY7vVRDvDA0OPuXHS5hdlRkXzoUlWcaVjzzfxKu2ngsvTZYEychO+BtrEGw7w72oKAbGr2v2KY8j
kOpLdraZhJ1eeqOk1U7sSffppad1hk0TuWvx188DV8wOvD3wbpX1/Pz+ZVa+M1uTt2fZo2BiAhzF
s5GM5Q8ccaEVlNhEY02HnhqzFzw/t+8JP0cHMSrmMHE+kUq1vViQt72YAcII/LYq9MFqGdoT7DpE
Hgc0cVX6AoF+0p3DDNh12ZCedekeYwQaH3LqJN8xk71U2luCyCuZxYpy6U88h5PrSw/T3mUNRqhZ
cbTOtsg4rGF0GyoPOUONG1t0a6a/PX+A+/5UG/Q2MskzvbToc9i//xVbcuSHIErzHz/0yvooxdzM
KwRlI2x2YroHnHfDRdwx42ryk00pCkt/ZZP3+i5VPeTFOPFw701NTl52jNPDcz+tBNQClqhWEFWJ
CcBVn0otszwD/g4mNWmM/WcLaJwDza2wk5eo2EZw07oUTgkuLYoTFlmJcVmPzuW5uLT+T1x8cCa5
gmi7diLV3sv+ksc1yML9ctk1V2wkaYL+9Aj92pixlf2ihE3rnfkv4QNHTT0NIcHzhzeIZ8//OLmL
PEOrvCNyR5bAsZ+yvqjqsd7H4yxZK4rO8Uki61H6/EEfroR8oz1cRk7idz4grbFz7Gu5LzsxPTNY
MEXyGcnm7q+DlMp+hU8ZtNBVOZ+7Kmn+zULGTu9NCzxujggqoNJPGMJjAt7ttbXNEQUxIwDexSC2
bBK1EXBHbpuleb7z0BzOJU9/gKex40znEVwJmFMXqZ0PvZtpBuouBtcHZyAvrk2Az9ni56MwsEcF
Ga2vwVRxxlMSGIHjoYVx4fOfZMtKd4eOY+/F3aVB9qaw1hoVtFiJsCovztD0dxdBKUnOCgdiGRdX
B9vJrusreumoAQg6OM3XFhSRYScnzvvEMDVCBR9Hd6pQn5F/C0+GWIharMpv4QIGPowzcFe05hu5
fmiWC7jK5zhHMZX2PABDbEhxjyx9HF5jMtKMcFT4K9MzqINnnlQCKxMJhQZeCzS1cqECs9zKyyr6
IrE5PoullpmdrCvxIw2TW82UWb3TzXN7gkUI2tv+kQVeVWCggeYwjyiHyoHOWLOYNHqsGIzDOuTL
K3DsnO8Uv/ECUJiGoaxiQEwUAl7CWAUzLEvkyz44QAVsFCSyRaRnu15/O+gWXRb5ODJXggykh7S2
dQsHO9z8BHTPIcgDoonefRefIc2V3B7eVpB3YuywZYD8FT6IHFMEScJFxm8uyZ5V9aMQoduiwsve
SU1ssageGKgzjFw+xrA0FRYMLxjQ3YDMXphUhw8V+nNxWkkJ/Zl3vnTiO9pWVaZzTe+za/lakKfq
m9pETWWs2R658jV4YN7y/VpWMc0upslvZaSo8s1JkzIHcxXgUmwl44f9w2k1mkibYtXJTMMPu0m5
EkWlCvNkLUOM1grSYHrJr0XLNB4G2NO2x207Vz+XebQwO/LQ2/1hmcJa6Tx2ZCZ1/EGC2ss2t6xY
Y2KGt0kD24CMXwAJbgyH0ygV9hOYiXTfLq1aZA75A9NWvE5Sccfu/GxFG0E7kkXYjx9K69k3zPPS
l0wSSD1okKEmBc4SeVY2qSJUmhhWo7nCRXThX4TxZPoJ2zdNZHZ7BQCWMfqpxhTPebJdPBSHM1Bi
YguKnMa/48HRbrXLrKcq1DoMpxHBRawGwcHxmpifTXa6sR9BaYy5FtA1Avu9z0CS2D3TXKceiR3P
sUsHpQxyPiT2DnPX6sbLRNOo+ecCen1Awk0EZuO8lkMq3QT9FJLMe9KhL9rSaBMRNfDcs8WaGGpV
PQuYQ2V2nKxz/8QJPpEvjC2xTRPi+u94EM1d4IRJm8rtx/xHQyU8eXltT+5tem4bLxS3enktoBh6
R4mKghp4Vl+PMq1lK44m94/UeWw9loKdT+zNsAbyOX9VllWS4F6dDcpYDWEjogXqrSHWI1eJQUhY
+Bu1cf/a4hbNWicrRzDuip1/NlsuAKK7EKmXzBm/Wuppe3mBOTlshbhPRY+BHX0FtPc3FwGq9sFU
d2jhMwp1Ln5uAJB4gkBiWOmUZPT5AFBWar0FhzN1GIpyJ2r6rQD3MzRY/KJWju6ISEgpJRf5Noxf
UYx6/zCIk7Fq307xNlTPMD8Vm27hYxs2LzRd5FAoTb7PxpWz6sR7XYgnO86Gx08r5y6++3F3BJ+d
OsJdkM64Nx8fB3AnH2eMFU7v6ZPMrNBM0Ni9DvYn21EwLsovHwl9eeii+6QYfM0GY++H85jSq8xf
5cTAkszhfSQPjwMMpZDEjwtYtfzp5WiYII45btXQlmtf/XYjhJ0DyX+cat+o+cGD+ZvWjBoIcYKu
4+8N+o+4euJD/g8snsNpNguxIDz6WQwBhNZAt2BcQpp/vG0dbTc4JWWb1jaCC8qcHM5OkLQQSaHE
uJ5pdBS44+YFz6kirwcNOnNSC+SLsXwF2t8DpUDlU0asoZWwiOGee27X7N2H4etSEqhlVG+m3rW0
DrfJOee88MS7W5RGEXo6EA8xaAAIIhglUNAHPVBwzQWzb39KWzGaGY28gvKCjvpHRphWIwFl0hHZ
gb6WL1uHYhGUumQKiK+SKmVMBeawndqIW2lEwFmqdtOmRtkvWNbLoOBoWgdy6dx4HI9W8o5hp+xn
U4YWZmls3u38x8oY2F8p32gB3iSqsjDwijhdWKdNTAQy1lCnX9B4Zb+uXI5OcW9Z5diMwAtbZJwF
YU5zyVnc15VPI1csP0cTbRAw7R6BsCT1v45xZYitM07CqXBeGnXHuHrN22iJOyVYM8MW2aaJPNcx
iuEpX1CXhv0UnXN9vqcOHI/lVoVtd55Rsge/bZtKjBEb0d57E2kjXkKzzLAt9EmfYxhQz5TPI8Nh
hzzn8V8VkrGGG+mDB6uzY9CmGOMyoHMDo/eD3GkktuTz0GhaisC45pDjdNi9yrEIUCL2lACN0uRW
qiYiz8dgLt31t8lqxTF+USQooqgwL2CNY4P5NsfcOIji2t/Lt2J4wg73CPtWwWnfin+3wKuCsAmK
SnEFUfPHBafvcVA2o8W3A0Kim/PmHpe3RYdmlHl6vlcBfeP7nZBu1tuISc9ea8M7MeFpRC2LJwFn
kVzcYLuspozXmp3kW+7AS4QIMHPSDkdC9bQz/rw+JYjTWUrwG/aXg8JoXwxbeUY9cY/MfHmV+4EA
jnp70CU9z5zIwXh1Jec6bwxggAAjWsUNFYtf0HzKvoJniU49TjR+7PG9a7hg+Rb4wVUTUR06q0GP
+sqgyfgjW9iHdBQShoLcv1uEg2JkUop9rbNXN0OBUGaesXbKoNRWhpEQgrrpLpvrlcaVPlGhd6gB
WnW56dgcGzocs4TO+Llx7WzYoYPkZ+kDVQKkoW9xgOb4XA+W4jkAMJihtjRTjpWEaxx2UXT6Via4
ZKXZnpCphH/7TwnOnYXyo9zXtWUNHwOugIA/k3VfHTmNdHyD4uIKaD13ukjkiCbEGBQRE7ihXinx
KQYdA9Xe0gxgKBEKQ/RMkikB0gFn0IuCYuSnhybfxbt4UiPkOAjsLIQRP+Z5u6e37YD4lAz/wDet
puHJiQBGI6SWh2iaLoVYq+sNsti1NrM30gl8ZkWeycWAkJLaz762EB1OzxY+74fWqqjtu6iJakhS
CUul90sTE5OW5mwR+DKW+XG/ISLAt1jeYVFvB9Avds8h8GTThqYEYiT36QjxpNAjQJ+7UH/jbjGQ
QrVjdjF5KfYlAI21lTLJGBDtOLwF+UDT6DDgHkSTl30Ng9L2l+dQ00Xjdt6Dnye0EOyIVhOaZf+G
cmWQ69CfKQgmiqlYcPDnOXguALxq13MSBHvw3IfgVrd2ZHteI64GgudCKxoM8ioUWQ3POgXksMHH
TluPk5v3cXxUTNPSsu7ai2xEFLGT4txzPdLKU0EgckirIpUcFij2OkhMGwA37s1pe4fWj9ief81g
B34lsl7uxOExJHzzEX/ryTXoMtPJ36Q/u4CQhZJUA62AbkYBGHs6Vr26Mdi4xJJz3N0PQUbHE51o
z1Yd5Zb1Otu/xEF0bZtq7tGYtzISKMyaEl/1IThZzubDCag0DJs/oa6xPFo/x3HmnV1c03lQUlCq
Sgs/HI+i1LrLElcoEwVytqNGwpbwo+P+HI6NaIXTKckzn5mAyjnI7YmYIHSlq6+ENr99G3frIvaK
YzZnnUOhdkLoRHAvhHFnhb0crUheKbMu4T/+v5QyFjj8H9kfMuedtzvrYjAUYFSuCZ7eb7h2z7jn
+fj4GYVMdnn7/Kq2hVj5y6X5UtXywjS22TNIceKm/IZOoWPviqIuUgULiUaYC0Ar0lbjGpB4QUnS
/NiU5aHNW++M3SVR3vOh/qBr2BjTGM87DXn5KaxVt0bgwCd1AnqY63VVDTzIZABY+AiAKsERC3rP
ovJX2CkomT4ivYqsjW3W12MTB115ze5dXz7LO0PxnxXP9eI7wIpaY2Cr42ch0NI4IMKgpQm1gD4l
rsDoRkg/L906M+9pU/UcK0jwJhQxZ5gtCtNBf2p/CFde+KNQaV72qIxuz7zSZiHznCTgGWpGP2Mi
5KpxJOrc5LeJXBiUTWXAlUSgnHo5uQUf2s0XrWgxB/B/v9ek+a6JxexVQEkBHvcpKnfan8VKbDSP
l1vljsO2Kj2Bw6VG9NGwSvRXp2xCQklqP2HD/S5aGfz2UBxj/sH9VEKF33EWoN+acToobHkC6zwr
jf1grsGXRpYk80HD3/jJD1UBqhXH5v82cjuG5DC9T4RpyJKWPEVTUFhEZvH2U7DThXEYOG4M7dCu
q98JE8nOzjFKkmLbLywXxnbJcv2A6vnXpK1Av39qKo4sxfMD8qNIlm8mpygPqB8oGdAr+l0xoOig
rp2WChPHy5/Kt+py59/Nvtvv0+UgO0UCTynbvpzJpLJt7gUWaOorau5iY+Ecsg2FGbN9gSAizHLk
tTNWe5JQHti2LpiFeVtq4PmgutdCV1DVKMljuz2VOa2S3BNNOLaK2a4EDBRuukpD6KsZzlOure6f
h5Vx0VDUdKctdTTXZy89J7UCkrdgSA0mQaThHHu3oYQjKpiY8YBrjT/nh+8T15yw4VNiLE4xdzKx
0NqpbeM1A/d40R/Pm5+/1DWjVbQMbROkg7WCUyKbfN2QiK8aqihY5OHQFYGMXP0rOv8quEjamwPO
jVljwTnYX3GRQWfAuAbrbc+5i4MqtXWmOSrtsrx3a2vXM5FswZoynH6Bn6JQBpV5OyvCI+US9477
S2zYXx+L9q0HT4maB+EYUCvmFUoPaObJlps0B1FEvfFkYAWjrAUqvD/GXE+ZqrBoSqTgDF/PYARm
L0E+KqEb+Or7R99yapvAsC3qxeqRSnTqoibYQ3SRSDvWunKT+3brovArwOnPjicfC2j3U20p7g4/
x3zEUE15jQ3xehuHb4dQ2pvS3jjpgrHj9yiNRMjTXdc+KgV6LLrZzHIabFmXxbXRqJRjNUaeH5w+
bqQG58cIbmic4YIQ3mtcG7lbAbtvYslx+63J/QpeZ3qCqdTY/XrYsxPK6t3f0iH6wTFRLmajMMZ5
gRqVALxZ2rKqAo4kfLQ/2a1fJ9xSeyEH+FklkuFL0wG5nz68/2YRsw40pE3kaQVyQV4+lVhfmgyk
C8vVkmRatlhA6qz0TY9yklQ8AeBa2ijCDBEITkVpGzypE3j0UHTCDy6JleKqDnHzqSRW9zun1CL4
ceZNYe0Hbbl5dpSKNQtYhIH5oEeYCorqKu/nf0tcvy+XLnpBBYMWryW1JetkFywYWzS0kHLyy3zf
Tsn2mq6mljyGlgG2DRjfXWdkBdKNRFbJwj9cJBcEV94ZY3nepXZ8+DCsoC/k5yAaJXtrliphCrGY
hRSwxSUh4pe5TmOtE6ZcfjEqpJri7skKgVSxwhB1z6g/lTYm2ru3xQy+8g6DlZ8+3N21HrUsMj2T
GowNSn6Yb+dg1HeJpmMp7uTqaRiRbtanZ0SmbJxCgaH+CMzBzzh6cLjMCm9AgOvNRMqlAL7KoyBL
ioDcg2pYDlBRXjpKfHnkpsJegOujGSqj8jCYndsHR12DE2FuAuZ+qy+c9nEfWZYCgIeIFtwm6RBk
HX4KYntg8xhract2PDHTM9CDYtZrtZiqfiZsl/oqYcZPW2v+EXXiq0aPutCxQ67o2q9oVXYvBT50
/FbX1qWZFpnmFs2qsu8Cn8aTu7pWiyCSjwDYa1Gl8XRMJAHtVLIlWtAjvgNwUYPRPrdn2CWdqdka
a0sRdklBc4YvyurC5vVrxXwD1rrvbh5agffq70lwAqzvne5bZaUlosbzvGwuXDEgNihkP4MzY1ar
+8NkltNvR4ot/cUCcEKRa3ITlJ7H5CxWe17eYkmTLh5/V+zw+XpJRAYK1UUgWYC595fPMStXwk6S
hjXbDs5NTU18SMK5fMU7Q1vV+LWoHXwCPJeIukvfTyDTkac2BCAonHLw4Lww8Yk4iESzM+tqflgX
j8HerwetwvrXwGxpiASGqyBmzkr7H8bCYADy+Ro+QdNj1VZVkDNN2YFYG03mpoMpFrpDeMn2M+uJ
lvhyt4Sgcpudp5AlSk1sLx6ZyIsayNsSKJrjvhazn4sUosShlolSCrZz/c8eE1Z4Mp/9kv9Pn+NQ
7aw7ilClkgodY9hGI+WcQEl+krHWfLYT8Pi5jEmDk+jEM15m/cFsOm0h2kSztKtGT9l9YDoHO0yA
IwiQi4eKIladHe4Rv1rovcoYycXJ4KZw7sYrkO97d0TgvWUKKusON1g6nRVXvnOmw1LKwtapOm7Z
17E4iFhg2JysnvQvIaXsHiy8VrSljv8TWhd2+YHjw6Orec83NAvt7c/BKutYfiHYGWqfIpgSZFfz
ycnWEWGfo6sZvfIjd2V5fKziJVIvZCAfNf9ekGHF8uscBnDMMKz6/v8XA0Rg1Vp8AwtzM0UexNxT
I9+lqyMgefvdRJM7lTfF+gb7I7HN5/l3EYVbYQr16Om8UBgmLLV9mRn8eAraMfm+MxMWGXE07LSX
AjZn+jl/oduBqOj/lr3PqKOsa5ypyo0zQtZ22prRyMivhPnlygXVBpfoxYK8+PdmsWLhKoXji0Kb
fSp+i7MHHecVG3ExO6DwEu5GU3tfKzTxcjdDhAD32YGBRZjoWNoZwds4I3kvcYGqtDLnVq1Z8sAg
1badsb5qnei2ar5oEhbqZM20Ej0yL2+0kPhOyzwb5UggCYhM3QJlQwZPD0rY3B9DjxOaYWzqEFHL
dv4MfjP+KTEFk31ni1JfGuw905yNnS9/+IPex1v6fc6v8VL2A7/tkGS0NNooL4kURZ+jIp5L9xaG
JzG8rgSnJENFkbj1dBHTAwE2zVXrAjrELpMJ3zhOr8XzA2YIpCn0tCMmzeu/xuXaJsMIdu0MELXy
/l8hl0Tx5FceiKCUwaalcY2nq/+N9A++/RuH8oiAsFwsP1W26rg43Nlq6OmSH+ITeSthYP6v6MYK
0rsDHof6Na69DTfIkgltCY1pyC8Qs+vfGXlPY9vMqKt7txY1lKVKmoowfDciXyTmmGOlYu9AL6yb
hzl8DBoe0UdHXJwor6umGcPWCIm/L79S8fsoICcATC0lMFtJRQW1Xcrd19mURXrMiVfnOQeNTsCo
hEziQoaro90JOi9eyz3CI57lFxWa/VKVyIfsAWgnzS/TPZIEHdPzjtaKv4XY4GoS5ITSPZyGZAYp
yOBtSeBP9g8nAGEKRsvpl0zA1jcGydYyjkV4rrjGiKVjbvDqBNEGtj6Ha5flwDCN7ay/IRop2YeI
LfD0OlZTgulCyG6wmUQraQJxtDDKi0aWEQOWi9ApMrQfqAf9Bph2JNUiyPvP80MGgpGSK1r2nlix
pa2arr2q+hEivNzdWJAD1z05VtAVnYDhAd+d86AfkQFsWaAgKrMk/zLz0Jj+a6waz6I0qYc3nKkP
IkGCzNt9ktoH4GTv0qgzZJbHsf/wXkeaj691KdXog15FKJHH8Ty259W+SNduXw06LlZbbCTKqlDb
Q9YpmMU/QWJQi9fvxtJQxRDqpVCC1VrIgNb3cAjYPA+cF0fWouFFF4AdZ3i6rGFJ4IY3E3eUVlxg
4OveAhYeZP+L3M/smJu6XXZLLIoQyWEn5NSlDuhUw4Ra3znK9SFRliG8np6zPe7bke094XtiaF+H
vPeypujHWQ0g3a2nlq4Xe+oihOQMEoqEux20P0HOGMzWT+bdyZbf/2PiQcdaQokt9Qsg9mB2x4EV
tKdJmLrpbvUBmVkJ3QsKOZ+doBjQwvgfXsaY9OFZbuQRLm5Xu6w13/bvctGsX1P+52h+APyKo7c0
IpT7mba975mvOnydlhl6fjJT1ZbiT5OXbz3jQi/A9u+5fRKbhSr1fw9Lhw27NCuZ9Jngj9cNXVte
o9SQNfN5PYD4i6Jn096HC4xu8XFkbOZY3y19vefZuQ27Ce9MOLw20pdxTPlKni5rYxEKGepSxc9z
tQc0g1F+2C+8pv9E3SfQ+HQPkOA22poOGV4aCRSBklXsnmO/6JypNCnLp3ZNeLP/UmH9+s5I+CNj
wX2bTI1v0ZIr5Oqp3JAv9Wy1xNUvyUeLMHJWGa2rSDpk4WbJBrVWXLW2yOg+LFLxcDWTwBIg4vsH
c67237MU3pb9CNnIARdCXllY+EAfi7LrH0060t3M2sir3XkCrZNNuPZDzykViELbJOLHP6FYZ+A+
24et0cPlgzzic3E8YHGQh9Nr5PXh/MK4XYKgFoJoBpD1yoBX/RxV0vEgf+loTIV+Iap1yfm014sF
63liAZQ7++vGdT2jOPSLbR+mk0wVk0r8BapSf/x03iNgH6FGp1T4tyiLHKfyu5s+mKYcO0relMSh
I7PRzVAj6kFN32d+/B7SLCY7lJXT2wWYRvKcnH8kZuNhnqGpULF57A0kTCm8T58szuVYovonKb82
bQ09Uw2EseGTOUpWQBaa+NK0WhRWFxbycNGIY1yK/h/QuBEMf3qdNzSWlbPy97DJUDb0cG+xl8iF
3vMcEA/anMLTW/JnZuSmcYQIFSpOMfgFfVCr1jxltcS31Km88JEzAb6McH7i0TpTSn2Im53Qp2bo
RenCzkR4+h8a/QNtE+cCFqtUEbnlYDfdBttcbvB0OS1fs5L65gK1DiRcOGFXFOOQmC6QQlBwqsnm
+mqQQlvzNfqYuGreCWVfrvIqFixaR8RVfBssv0y8tTjhcU6HdvQ8g3p2TnUydbDGnk9DxuAwnJBJ
/jNEKvDhckp4t3FV9XxaPPHxYSVc821fSJ8iHJx7P1XBjNa8w96JhLMdu7nnZxitNiOhIlcONcr9
o6JQrnyARORetX/FEEBI8AYlcr45O+ImJcQGHtTE7cn8JS34tkENFPmkj2pz94L/kyyEZ2HZTuIJ
ynHX/GaGJianfse1DRNcE8XDjLSGLeblDMvGksDJSnPPxwoCrdczZ6e6is6wWdHGeI4t6KQNj0D/
3LCszqFm+GHEmAzF5DZjREXb52bc7LktGOaPcGBqqXjHRJgoPFhRmhCnwCejgRdtCkEgMGyX8Yco
KhCAb93ZgcJXVaDHkMHD3SXQz5y2VYOMBwKTkqxKgj3RyHaoxZRH9EI68uIAQzBplmpfi8x0Dk3F
hwPxTfWbGcme/aJ5hVlZM32B6s89nvbkCQlgzZeK6aNKXWNCmRUGHZ1vxMua8mTfXKddY/Y/OkR4
eM86tr334Mv45Ioxa8yG6kXosumL4ko9Q7G8ss1CmzBkO4ei4IsthiOr6uBEhelJ5ClqrIYb9Jq+
0ejp8rrgFYigVJchT06C/wPcqP8s+xa2FzC8RSEgmHKTNnHiUfi7Q8i7iHfHEzzqHTb7YNTZS6RZ
lCav4XvonNrJsHNSzQostYmntoG9o2zLsDvsD9hWcGd0i5UXTm0djLidUbbuepE0Zby6Y6hPa360
f6efDA6H+M5UPPmdWm2mKJWUYPoE/h+fWT7o85a9fFPv+4PqhDqTFjjFdKIV3jskGPe9sutZqX2p
PxVvGrqurAeQZT1KWHPY6vN2vyNVyciNn+YjTxIG74AIrGm8SZb5iMJMdLnZbueK31wHdZuUJBPh
GUMZ7yTqCnrX+rWBAsX6WSyr8cJ2yXUvN3THFomE04zmVH9v42r5cIpAAHmIJzJyQdDvCq+aH9aH
dV5dT6KmJNROhxhdxWM2g9k8IKdTX4F9KJuM8Z+iiYBPJhnEqFNQZH16xVbCcfzWMPIIlwNGgSKa
4Y2cguQUV8u1lRWs1dB29NMcXghudClDlACOVmv7oUlXmH/YcVE08gnAN5tHQcKhyum2W6UjnCb0
V2VsuVVZJH8nsUg+/n4hoL8WHgTU1dhVLFhFXxyZe9Q/ESNNyqaCK2U4DEGhsn1bIw8NNcrJ/RsL
ZF6ULE5qU9FX8U58/beTNnEFBfXVBb6qvayVZ/xCJSA0uLufLn9PyrEeRm3f7ZfisH+nyd7AsKef
Ix8bGv4mT0F7uiPC6eO6jvf3lP0+jwhw+0eo2A/KxI88eB1L65txjKOJLqKrJfZfFmg3dVqFv2Fp
ow4QDSLBb2vI8PQcNwYM6aRY13OMZHorEV0r0nZYFfmPeW5lW/gZaUsE+Kzh8J8SYIaMAPorhQGo
pB97oO56xoGBrFbHNOUQcYikX2kWfnmhl/HRbHkskzRZFHBw6gjkIF1e0mG11uFnU5pVtWTE3WBS
sy6y89ouGHnFKuz+DSbjtAA/0zNrtZVGEwdRLs438tBOCvXMvxcCNQb2+5urG1f69H5cpP0R+1Zx
Q3sq3o0xjiG9G/0Dz2MZiydWeh9CrJyf6rd/EHKwYD06z812gNMV4O8QEALThXkvcQuO9Y082gNv
WoI5s6v2EB+bdtMGd4lQRXnx6fZ+KGY4ldg19AZcNUQ0+C+lSAUTgFwlHUaPI0CJA+o1xruLXg7D
w/Oxbye0rb9Phoqn3CPp0t4nADyDvAwj3MDJJoQVndZc5W4vsGVM2+acvTQ52NmXeMEp39JexGov
8nzinRkl2I3XN7HEEwPfrImvn6jfVzR1xkng7cvq8JZG5lCKOnljJMZXDiK9PRYgTtgzVojTpx7o
n3o4mFl8Eha+QdnjM2x8TlO2p6IyZyyHB9ZmrKwtIPdkbTLjQHVxUO3HG93Gd38DxnoQZsVZ+M4m
2EyAxju/IrO5fZPArBHqk429XRn3n4Iao4HFklfkz8aTOJe1+nJAKajIBd5S/DrY0FHyLFkcbIfW
ItObdXisKSm5nRKZKRdppxDmuhEyhGARbpSVEG1nvwsiYUydnKDOVwzQ6RUu2bUaTb7bgzPW3/8R
ZOzxVW3zwJTuedCpAfP+4YhygpZspbhG4RY5PYBo8lgE9ao+lcux6eVdOVBxXAemN195dnIbaBf9
NG96gwF0STuNXaJKWtImkSChQTjsLULOqYxzHZuZ7HBM9we3aE8Tpn+gW/CzP5PbpJU8rxs51flZ
jCOCmBvjYDaI4jrC0/RrwL0XmJ5h+OpyDr13MX9JjwF8VulXwqRLi6FOMujaFtro09aWDCOBg6FV
S38VmTTpf/Lf2UXc4wPqn1AvaafP4DLrmD9pgLdF2wnr3d8wMdTJorsBQRYSjYR7X0oj0q8FWUg9
AiRt5ielIWWeyoNtjxyKHgbPstsCpuCJDj08jCghvx93GaFI00PfBGXX1PkLafw7Ps7EoqCypaK4
QLbKAWmV75ABZOrdV1zwVlo09mH0qUrVSji6bqrOsCecyMrS1xi7V4haiM41O6fhXLsjDyGVJvkD
lyQHkJ1Me6Oew8A9UKga6jX2tnlQmwUQKjEx0i/XPakz/X0MLoGKWVYtKFtJGgqycM6N5vKnwHuf
BBqUrZsPSmXvIFiu43Fb12ZPJfJHGtAVTJKeOVcUEcGDNWHAd07KpSONvXTHQ53aaJPymhdPZAWK
lbYOnODUHaWvR47YamUcHj2maBtZxt0RGAOcgdpVtq6XXrqSCBk/CdvX44ul9luue+xosukCa5O+
AMxJe6AHrn6rtFHP5+0BvMV/KNNjvXxsMQoEJB1JnnqbaIRveGj6SjsBbp/9EbLSoPHyrCRUfZwT
UpwCFJ3miViOjHDvGtu4/B2V8v79OoKx2zvfqjeeW4f12LhxdDlwpNpLe7Bcr9FNIhgLHvqmwyBZ
R+WnaYdCfcKsnQxwm8NkzY193D2jpNDqWd6PSmJ1RPiDpGsXZW+xO4B2FPk64QD5KqMrV3ZA0kqh
L6pxRkSILPIA5oVDkzTR7Wq6L/5D6Fr0FLo56E9VsmOJShPbH0zfJwBndVIr+xQbsomsqdpM+2gS
5Fk0/2myGG0HILHd7xWZ5b36t5bCg3vPo3isgmfpDnBKkDdIThHPYxObnMohznk32SYnQSr73uzx
0wklAnUDpbzFDRM6LaUDAiDgvF6TpQnBOrgxrylx0dCRTtZuTmLXRQoWRQk2Aq3AtrfBef+SjnIo
bW4eZw43kkVLgzpmtMpX68UU82rEF07QVrxy/yu7NwzNRYpoz6AYKdqvkmoJsqlCjDur8txxEtU7
SgV5bDCo9p39Dl2wsdYFIFVuq6VduL+sS5mcWtjyG/VMSUe+IRrp0n/MLLia1JqfHK1VxgrvAqCl
fBZsQcf2l/6pARcAWifnKyA9c4Q8k4lhGEp/qjHHJGGzCiR9JA7el/WKvP3Zo2yeTawfDF2W1kG2
/9S/qd0WqaXZsfuakkY6FQ3JnuhIEGaBmecFgtFt+4bDTC7b+guYalEmgPDAaJV/FcRg7IWXH0vD
7qoxjcW3c6AoorIPB7t4KoNEGtIhBCD+/pixh5eROKT7ucRDWBTn/d24Ie2CEgf+GBAWWQV9idp9
lj+/yaDUmRybDP+Qy1Ck0LSSE+qm1X9i/J5USFTDHvrMcLIBSkhxb3Ke8pKysqaYVL5oATHwZM0t
BPvrxZja4c/9zEAOnB68ONT2DhB4vzhiKfZcQXtW264FmyjLCSUeExIb/nyOnJyJLHZFIq/uWSKB
xECn55Ef15s4Mo2MaIF7LcynGf01I3qOfMx1ImzKqI5l2BuGLmyEACA8YWvBhy5ciZ2LpUOkF6kI
VAkoZ8VYUtEaV07Qotl8ijp3IjWf50pF6EPFchbeoMqB0EynM0XCSaSnYA6ZEmxwRZ8uDF8bIT3H
5YX/Z771QglLrzQf+3UtanDli0fYfUxlep0K3F+xpBpq+v666nqvkykr+c0zRt6UPLB/BcNBcQVL
nScPP2lRZDudXTFVzYqK01uuBpMLSNS77vI+G90Dy2RqYgDdTCKbFwTGcPF6JTQAnwvQC7ESDX9T
jawO+JYTds2XBp+pPuVMcwVSJDlso/uZ2MTfeSqxAvI5BNzpILI+3eJ8+xgoeDOYG3kc2n9GELqp
9h1hJbPYsWSHrmZ7xKaevI0m5HORTNEoUWPKhWcLWAjYYwQdfDnyp0M4PSD2jY26mGpIQXlWR3CY
RQYJS5TResdTWKELRMKfRRwRilLC/5T4hXX5O7nUILlixaxESurxbpvtOhXXwep4lsN5MUCAwmVK
awNDzReY8PP5ScDVlSV1QfHPM4BnL+FjCtegLZUDlLMMOhdn2aDcBwwal5s9uqKAuBM5eQRylqzw
HDv8Xpew7EM/IBVf4I3qo9F/425G3lkybKF+N22In9vDIs9sDnVFKPtYd6BDQd2fXu+FyEo3w398
77RS69JftjYM2iiESM5YxZ5rFChOvdUsAHbzmqs9FgOmqhZtcwqN4BEk+eleMmHzNW10MyFNNs4e
PnKJr1i7lnx3mc0tlQwGwvDqBShnzrd94CtqBSP0QbdRf6clgSwyyY7Fv0owtoWbTgULGHHWqNxS
5ip7UYrRmMnWP9632NCkiYwUzcxNyK6JBiN1OyE4A5geWmT8Bn2bRmCAK8NDPiBdE+EikNKfcEyV
tK3VwHU2okTVOKwkeX5Oe71+1wvLj8BddZ/BnJxdznY76jMm3ITAOy0ftLd4W06rsYsO2RhFu34I
W/vFhtdWfAm60DTMhG6KPmBwk02pitWthKCXg4iUUMjfYImnzAyHt4GWi9QteRfTR+cq9nL2J303
Z6b5IaR14Zqb1rmqIPhukDfd+C/eecAE3VR1i1OPjFYL5ONyozpwdMqaZNi0meKynHVaqjSFynTm
KaUdObyOoAp6tw5K8NsexXFC0r1a5IC/hB0XAKEbCHHLvZUJSBE+HaSWtsF6oAj7o9jEbGUJeJIb
kQsv3sk3oFWXXRfLqwZYrO/S5nUNxvI/UYiWXkJldqdxUnYLxTXAbovNNCQp6gMLBE0YjCbQk0Al
V0dQlbmI3eidRarnovgKA9zA30fmYprkouKS7jT+V7Q8b8OlmhJdU72TM6Sh/L3cGKJ9FysMhKW9
2c3u7NlL5u67312fw7K1Cfuax6FE8jAhDTT2wLZP0qx7fmw8xwesL0tzoaXuTmNELHp+cyhIgPfn
0bOtPjWjGmQsTw7y4FinHSQ9po2cVvd8kAeVTbdK2fpbf6Y3ijLdlXzWU2DaAaCIIWW3MdbT92Xo
HVrMMIclwJ4p4X+tb7VTYI1L+KVyAWOOILRBdWOUInzbZZYHENfL7wT42FF73X7rJq+0G12XcbaU
QoWClPbVyRYMASmt1l1876uZJ/2YNTKm+vB2VxBomn3EO7yzqJlSZtwqGF7jILPKsG7c/WCrDi+r
lN0WIRpGFHAjSnP1I8THGwKOJfb3gLBNLhXs9ywdoYGZ66SX5tpaJGoWrwSEhcmhVA+aveUAwPF2
q5q70LFK/5r2D7ndSMUbokc3xU4+wCToUi9jhfxEAE+Smi0aQY5tnMGhVeRk92j+WlgmkY88ioOM
GTechotjhZX1D7B5km8QULkhNVzASFKoPPXrtc/n27Wy8eMHd1EXhRaJ19nB7B9h4Kx6Et/IjVxi
B1LB3BlwmFCOaCMyDBRsIDi530D2EudK3gqymfMEl8jhL4QQxos6FSVk4QNyiqZXWEbDinFDDPE3
yO9HYBiX4yPZfwVbYfG7V+jlNnL6Qg1y2S+GkngTpsNseFs5dnYWM7VHR5B2LknKeMoGtjRxmlnJ
D6DfKnVvxToqYKuOcJNeWpE2ucuTsTSDoLkXgWKT4SOiDXRxaHSJHeyj/GIqiH3oNPaJ9C2vyRnr
p8mZUyUvXyzw2cz8Vb3QNk4VSOO98I6KRDKsTHXYQ975/TuzqRKjwjGIr7bof98xwbpenV5fhglJ
qE7xpjXw+ppQqsohtDzU7BOrXY6Ryy+rrvO/3Av4GKlsbLQbdrPSMtmvR64toPn4Rxs6BmmF9pb6
5gO5wWEeY2BWFPzQ7gHPMyek9gi5UDiHB1zsaKAPvPtLoytPU2q3e6srF726fni7Vv2h9krrBSLY
YIDFHyKEXdD+TushCG8TO+rjHwQB5+jmjSvNPACOExl6jsBwcAyW1cLlMOCbbYMH+hJ5l5pXI4p9
Wmbht5FUsajKjx1mhF4lgxnfqoTAA4r9H2JiV4WQaosmBOHyhvzyi+cyckRj8U+n0NbDeCch6PBJ
QKijPfkjcOsC6DwxEb4ETyYI5HjKMf/huHPmY5MQZb96mQIsLYkI3v01J4R74YLZ/SZguuaYdPG8
hn6QKXf+aNpTCdw9qB+a7gcRHP2fWTAJgkULw2vv18nA/vfO/U8kOGKFONLPhcw2vNT9FtrSz7vy
WxEp2ZOrcv1HP/zWeaXkgTV44ykZdpn4K7AtzQ7/uA2qooeexABToBxhIaL82c+jzUZEX1MEYHAH
QrymGkRvwYa53RchR7D019ntpLpZ1Cd1D2p3q/Hmu2KZB3kgQT7LnyKncuRyBSp+qgO91V5vUwFW
A7kupPPnQfbriyqVzm5N21LJ+WlP8nfXb30g1xiDet+5CgC61Mz9NJ67IuO10Dv3y/rp2ygQDXoT
9eIrSsAD4ppFJun/7LMyJ/yvpL3DVs/iO5I/eRupChjtUMA29P0xnn06XL3mqEhZb6GGvs4Orbow
zzNu2yaTMDRM6vYJshL5pZ90CM14a+AYNJKbttPd/F8i7y1FQxe/6GkgJF/UbzuJQXXfTmmwQzJL
QIIAW3WmaVRj6zDRFxVk571Mkq2amEx/eU0DR7HjKEswr6G+LNuS3FolNr1FTwuJmrm64DeR+ejg
/5rSEHN1GhpUps2TmcPMPwYIYHlu89VTUIuMPzmiUGg+Jgs1dTXjiEPKNNsRJNFDvoj0dwZcrVq3
gdZ9JcetVYlC4+0iotFtvJ4TPrOJAsc6aL90fWpaTBwW2TR5fcFmvhHEmYdqmbrimmi6lSQkvpCH
jX7TnldZZkMM4/6locMoIgXb9QKC5MDj/i2YbiWuA728qAb1dRuiJEdRXDWC5KUO1jbYYP70arCv
k9pfBVmD7ioB6jQQMUvKEoqHBouQ72XHlewpQjMv+XoJ02Bf4QzZy8KqQhSMFcuhuS335ei+JMCv
P8Rlw0dVzcw4Nu7L7BqHyodMxmo+DLP25eQ35j9T+5bXuNqTH6Vf8DqpOCW/wDgkpZWVpk9oNL0n
toDefszNN6+ag9e3bPiS15MYjuj5URXwbcb3gmDMiGKPh4w/cQCm+nJTzuyn/DAvfPqZGUNVsFGU
a3R3AhWAHj1+DS4B7L6XqqsiHTAokbuM7Fs5nIiSMB9KJhnsD3ZOO9V6pW4cov64mVgn0dipwms4
lZyvTSd6UY6I9Xvj6PiOZS+f8O7taAcBNdri2fZhnGlxfTh6dGAlEGvXpzq0IZDjRBB2Mk7TAZIc
ZgQLEQ0GA1XS3FLTL9SUbrhcN2ljP17KEnhnheAM6w7u1XQxkTT2m2WpX9boBiL8fp4uhrwAhtWW
1YCI0sC+s4TeWzZZxqGQRe0/o4/QHXDdZVQIuetRgODHJ9+Xjio4N31WiL1LMSy6Ia8Bu1mRABZ5
8TO0nwbDouAvefw7aOWUNavH1eOrIrNnY+HojzTUylzaGCV2Qh9oVzLN4CcHCfQecMudkByrqHwz
p1dnzqKLl6h5yc6JDzdVmDrtzgv1RKhX20od6FIiSuOWkZqdhXDldUGYXJe1teAYPhAOAGOEAQB+
jYr5ghlKrHspEeHULed/pyuIpvsvkSPRDnX2MmP3xUB9pEGs6CnRV+PMqH9tIHbrFezF+kwzz0TT
z9xe+KyB5Y4rjlMM6uESgws0Fwp73cZqwdv3bLdi3aUEBW+huz1n6kDMfgU9yLO0fDQMnqKMRVl3
Q2RY2kAXrpYyzkcPkP8fvf9ByhrH6RaUkBukc6lo49OHD3tg9a+MVqB5DZwnfNMRrTzoE1Luteza
glBFlp3XoTNA0tS57Q4J9o4hd6+MgMDTj5RCmgdanA+HkHLicfhZtF8kX8pZlDjJ9U6G8pqYvPMn
tU3eJZ3BHwJrdZgRItLFkFjF3fkRUGz9d+f/igS2u1Q69YGVAi8Gm4Yrtme5IcbuF9tyZIN5o10i
7V7IzlmOtCh/MSqD1C3be7BgYjJ2zBpqcaVdQbEwR5mQIix4u7lr3JswV8dfgMWFfKvtiZm3r9Br
d6MNV6ovbzWSwBI2QqVuYJQaWxV3oNzf6iY38aHUYM11hqFXweSJA7DpEXH/vdvFa0Ue/zMa6b4T
OSL1IOUGNL/+zP74bS7rxFQIEx7l0B/o8oQ6ScWMQU/wKtNjSOqoyqtovBVw2SNpHFxOwx7Lcn7f
1Xa7FpnbNwska6DF76LQInFBRkEcWMavnfhRfQyCu3g7V/wk5Ws6ukBH8iDqZKGZGB5BNbt4jf2y
B3m/Bkr+uMpJv/9YxTAOBge9U6tyzvwGjyhF5P1v7tr7pot1vXO+A1PL0VOzWUQDvS3odIAJBw2B
XpENBT/uIu0MPoZUo02TezDX5deuL5bkg+vrebTx3Pr1StE0lGIWmnvxwBP2STqIsaRWuc34d5N4
KFwcuqJ1uy9GiMxed+BiCajvSC5Isfw7TQXwj1ApP978hJ2ZKVnQbeR2V34O6AjHwYdZx2GTnpIh
vMrke3kTwsEyI5bPTNl35+s35BUY+It48UAR9txdsltFBpjCUJSjl803eWcxLcEnWanIPc/Ya/9v
8+0zpteHrFtP15klObzgZfau2gzzwoIAT/fRrtP+DqZZ0zVYBrnSPuajVuMQZLDYPy1CedeOOXMo
TT1yo486JCpmHs1yJxakbaPNvBbP2Q2ZnE2buAxYpzUi6CvZX5oKKVcKsrJgubb59KsErmOtHQ23
w6JJNamxodXQV6YZk6YI4kAuNX4KnlN1Uya2nlwBUYd2B5ElZNuxql/oi83rGAOv3ArqQ/QASI3t
dn4QZxwcPPRHgUFVNMm3MjCN/lznELJN4ZDvcH7ULS2la8u02ut6IzTNDIgVbEX7nZHUUn0Sfbqn
DuscymfVZh6PPgwTr5ZgRGrWmrW0r1DsB/VFn/711h3C9JYbZbrDt1fpRZYFe5F9OxWRp0az4e0L
sDYNjmJaRNdp6jm3diMChGa6a9AcnSrpD/RnFKkZLRrO5ExYSeSriwMM/bxeJ0S+DU6N0LK8DAE5
df9WGkxgBHConOpn8e6MlnP+262Yu65WpiVz5kdOnBy2pQ+6D/z5hgXZ3C/ijaFrdtZrgMD7cltk
mmhNm8yYs+hGxpN/dEVZJrQcnpFPz8aXkkjf2IcOZ9XYDxUD1DCrsGiwU2tHJr4PPJ2GetoYGTwn
cHNq3k664vT4B00NENTWRzHqcA4+jdyBu86igJargmf6hNZOqVfZrl9yy+hV+Esw66OUkvCVkp4v
rugUEyN72H3XfrHVQUzVIBm0vaUmwHlfJA4lW0Xij0HqvqW2vYRiDqW8UPouWBX3M8ndyjeHk3PQ
S6Dn7ElTyAi47RJGKrVKg2b8n1wV/oS06HTntM83Ex406mFPQnSlbnacgM8p5GSWXPESMfChlDqu
2wPdhlSV+3Vf22x0LJktc+S8Hg2h6nqTF8jXogGGmSTvIrfEvACZq6ZzCT+V35AlPYLw64sGHDFL
VcZcve/S2KVXTxT21aCsffNoHo4AnmXq2+4GoBPMl/bcN1oxRbhMDCol0fgcWUQYpAbeWYZpVG1t
Bl22v6q64BUiR9ETaXhTaIexancJO4DFHTLQrCDjpxORWWlHt/1u6iidRtnR2gK2khrNMJGLrjpk
u1k3hZrC5GwnKPchv2/QrWZyD1yHXoI0cTgvY8Yqg+D3winC6ZxqsEzAwdui3/dHL7ABERcv/oas
4rzTxOHLGuJsWP2K8kowVA7lltxFvc0miIdKaOgqju7nvqXVALihG5L4E8vjYrQVPIhY3l94pZ0Z
W3anGqxc5QsW4KdzPIOG6u7Jk7K+R/R82/BXu/0OL/1AUTzfWqIlh6Bq+oWxOulNT2XQlCa6/2x4
4ktedKjvdiBfoI7v3qtD3ERG0awNlq6KozOPjPER60qcDbwsCyh78WH7pg2z+r3wlmWUd9wiGuF5
QqPh2aXr+6hR8GFE0eq/2+Y2a1EN0IRJaAb3x8+Y+kwz8BcBFP4AyTniXZBBJV/OPgeBmOViNFe9
GXr3m07SiqmDppt+UPPtk8DMIlx/vEg/nuK1P/hkQH6ZYXrui4VWFsNBopm8IbYynmjrkerzXMlc
6mjeSyoX0QxYS9lfacoVrNTTNkpgUYlkNYDEmwvu154MMm5nHQ9gFddhGw1JziLpBbOzcPL172IR
UsvMFL+MRsuV6I4FW75l0gYYAyleR/CCPTUsuROwnwNIv1oJVOFZ3pVT1IbuMwn8WpVmbqGHmE2T
k3v6XUkHt0a3s9jmc4XNH0SIrORjQatqVYr6SC94ASCofpdJw2df5/A95Db6U/6+/WSLoxRcGdJt
bGjn9CqqEtUto/0DmlMB8ysUG58Mj/TS6HEszq5tosEECz3oLq65jtEAfMDy4Ljc/wKURlfIqgsi
Hsy1zlvQzOclmz2CUy9Zwnrnircnj7p8e9YQTousAqhXFQ7QIU02WL9fp7wR6z5mEqF4sTgZpIw9
GqcG3AkSwIpndZSKWF7wstGPLzYlQMJE/RQ4cSUgQFeK1uOj9pIxONt6/cx0XLwoU8UUpK6jirVM
4Q7OEZFTPVDEfGR0KhrpI7tNsMXTd8fxHa6O7YNb+OKA3yoNgQaGWZxdSBUJQJa0MtEu3xxKeAEF
etT/YdNzUZbFOFaKjP8UlapSIBIzOWjCOYWINs2il6fQ7/jSFxTsn8gRu0Z21hut4rtoohtC8Nw6
LZmjJVJ8VsEZ5ta7+HdgxBpBJFhb4lEqxW2MIvFgD6v12rt1t5JIPPfwFCGBNtxeswlPPM0tFI1R
aLFwC2qKs+637V8//nMQwBj73LpC07mb4w5UT0PJe9qgeuzfNnhNaAeU+0WLmBByyq+kNz317JV6
TSVFz7NBDDfz9ttlC22Q+4Alkl/C/wx/bOiwQYH3B1NRhOgj6+GkaTCqsbTC61s+e3bG3Tu25t8W
kfrhy3SPX1m6mVi2AfYCbIJP8zeZwLRejgCPQ1LyXqnw6U4kba1vEIFycYn4K0BEWhnfjvYtr/D8
ywBwkFhY6BfzczJ1JBy4pixoPnt6FyPl3FreMcjg0ZcsQAOaAXhIVkD17X7uAVppqVH+ilN/Usho
K5Gs3MuSWFbND8NAf+TsQWV/N93pCx6WVmRHggz7OQPoECC9Ayuij6CgtfE6e6tswiiHK4HWyds7
NzXIuce7ZplC9anYrUnVHSyhNzrxW2dIfNElBBQujuhlZ8hwtvRtlFQAzJjSG3qBBk4N9yxdU/qD
RmhT4hb6zHD5hl2DbRuTLUifoXwCPk2n9/iV+X750qE/nmAMi765sKJfD0vsmVaHHHlokx6A6jmi
Hj1zamjjIZOFtIS8o2oVJeC/P4ZHG14RDMJmtnwlBOZxkDmH03pw2mo/9y9i09RZcfXH6WXZGs8s
GsQ80JSoYZEpAFgmE4uf9ScURIut3xCXo5I6FymHRlpQ7YojjNaEdzaRgsi462ivoItJIl24A9gS
CXzYC4YDvp6OL4UrxS5y+4Vihvg2Pjv2gaD2DnxVOps/oiFZIZrC3EUEv7CLtK2sHF0djCc7Uah3
4XLUUwBZu3GhRS5Zfw3+NpYLAnRHHdsqz/cBpFq3W44GJvxK2VWGHxgLW/3foEGiCXY1YjN5lCl0
QnANw5+pkOF/KmcFryTVs2N/fTeMjGzIGrThPms4fDQ2hy7YQNTAWnKMVtIpXJJbfvEnW0eq6Q2l
fG6QV6sAf2BIYCgQH30/S2GYb9ETZ06Wp/yd6n2njk4nfiXI0ASJH9s6NpQgTtQcr6X+ZpDU6QXb
lR41SrgR3K4x3X928PxqN0W34Ie1Fn9M9mTFl2XYCI9UAicZOamnU1TM564Ao6HPkQjqXLnuZLVb
UL+Dp0Jyy9KV0rIhRyN90JK6rz13tos5Zw5Q9uEaHzqdZ2TOuDg91ULAmXPHjE3NoySt9BCudBbR
40JxA5vibxpAldOqfn4OLZAXEH0cflx1nX4YT6WZK7YwlkJFML4iuZeQKvLNvCULrE8Ppatwv2CI
MgSgSwqAcqFdt/t2Ypstgz3X4jO+A4TM+JPOSUc32nLN//3YID9bRiISiIJ7ln3i4+gkE/ufp2IG
PnaHXPuUBZqf78h6nPUqv8EGridPOYMQrk4GBSnr2WNICdkgCmlLJsol+YJ3P6GqKcWSYBHWtSG9
UB35NqFv4rN3bDp38gpP8vCfGTkVCdTn1J3oQ5iNejslQDfKetv6WGyjXi9UDdJEv0oq0vZT3Se+
CLOPqsx3hp1M/7qzixsOOP0JV+vxtirYtKauOZM1L1sPXNrDCjipzBq13WEcstU1bk/1Vpa/R9X5
9E4gcSQto2wyrerFwKMsi9VfMpWt+LQxQKd5hy2pqSbhrToHYntxFiYeGtfLpaNDTlcrql/klAF9
Fyn0hedhtBm2DlDrSmZctzvR6PiC9Az9qvBHS+o9JMcuyjwZXMSUEv3NruT7tP4dQPgQ+gQTjrFD
IHx0NnhYSrjcrm8rUGEfEOAyw5+L0zR+axW2c7A49S920evbOp/rzjVn4T0vFQnYz2suMIc8gcfs
JBly1XN6xpI5PSp/IdoGkfK+tFxTolDQx37ZZ/IIbjGWVKqnyByvvChaUhxKJOgBJ6Vg9ruLmiQF
oMT0yUy+zGuTheWTyXOTZpjHlkLmffYC6VLjd/qGcxileudHek/PFWfwczqIScdlUkGX5TdY1gbT
LJLMw2w19NAqkJKUiIidQ6TT+nJhmU5pyByyD9O39ZY7DHsAk4upmJTR2r8eEyqi1JPiTlShF9Pe
TLL57W8Xdk7qkXU6wZ4Vc1iR0q2qQv4JPqKcAZcSZHkJnLvxl1qD6YB6jBEoh5UjVs3XbaNQSF70
uHmxlsN0m0NNnbvO43JCbS9agr7lJr2BWBYHpGpIXa39NSDGboF2+WWG/udQ55p4FkmvmH+aXtEy
H/g3uaxXepLPI2vS2ByFzAy1WyPIZiHIR09OkcxdKKp3HEy9ySTMjb9ygX+PHT7kovV8dscwIybK
Lf7EigBelCWE2QV9q6MWoqQAJ1UKBAhLyBa8GpRde7snSAxN9iDgx8iF1Q3HGZ2KxS2x8e8yLO6b
W6Tl7jW8cMkZUDWarF0bZY4NdXEwb46OwK1eMEdkHEe7zv1zRIv4oPtZAiDGiRiGjKydwa/den28
lQ53havtSZgsmaHcLMkXD7NhrbxWhs2ZTmwR5fS1YXfIGbfNrYy4g7fUFLaYIc7/cU2ZFyxRRQYB
lDGxdI+hNDk3M/mPFLtMBTwbrJGaabHVHqM1JQtmVYAxUhhIJnhWSaWI5/+3Gd7g3PQdSyC03M34
Ta/rGD41O8Q5bCyMJL0bZ1ihrYetOYK0clyb1JUcoQxU68iXGDEDyKVHI+RNmHuFoBrMOSOdgRmw
4ZTwtEQ4bkiN9dOa+6ERBk4OctFGhdvPWJHfcizARoZVOEHNRufuQXLIiVUTcCT3oKbdgZb7XM4Y
svwAR10ezLJkIIsAHxWlMQdJjvjnNGYYkHtXkiMvQzGTzNMutXxSzvXRtyt+5VXSeTkuGRO8h8+0
iTaaZPLWV9pOVz09X3iXLLIi8/TKMmARQazzYre3fN+HPYhq3zAh+tlJHF920kOqHbFYXNXFgdNy
UnhEjhglM8PBREWAzc7Jzfgh2vFsJFbh26p3POSZscmumYU6IF3P50f78lFJ/psyJmXrXjXf5sJg
utfmEFJzOfSywh0Sh5UT8TmFWsRwQBrNpGGJTa9rsQmhl9KwN/l12awqDyvUcMB8mzyQWAdoOrSa
1BLUY+DvbLX+6Dbisfu/Vm554TuZeDunJyiGKdAdLWoOhZ8qpy6hD1uZIpwOvPBmJHEtszdBXD/m
ZWS5PqR7uXoXW0efOUlxMWXkatRGtP3EzlpqWjRPoRxLN2pqlYeRlilw0IAM8FooYtHXNyAGKsY2
FsTKa4g9nFqCEa1xThTUuNfvbwpKDch88JDRWOxduXzmN8eaOHSqmr390uXZgAC7NRBQ8EXxVh9O
ZtjQcL6YWnI1Z0lBjy+safzH/J6HMoNqzI+IrwHcM0yMfZY7C6ip6TbmzjUhICAeiVEY+Z3eYXMr
/NdDmGFAEmsa21dy/UBNUIxU4M1DJPcMzU/HgG0EFuQAPNSqqS1Evx+v/+o/X0zYsuT0X6BbDkG0
wlDVkSYj713FxUlax0JnxTDkdmFM+1jYMm9jJ9nKl3a4oatTwBbCeNBa9clqkQVevn03riAu4gAq
czh6iHmO4oqk8Hu5885WXav7c/rKY41TazsOVi0gN68TG1gI5/S1aGaGzL2xTLGij5SzbKpHtmJD
/3lvs2Z8Otgnw3ekDOj+qZPZe9bsfMFhUSxIRIOOokJqM1MJ91lWJ6OuoaoLIA3UTSakn0NFbl4+
aHm9FrBJGvd1g/NmMwZoXOXzIj3W2aQHYYlQ30+pR8cNLqKCi8eys+ozSUlkvaiy8bRt/kj9BTiQ
7os3EYKXmcz8HeunhZ7KyRJfZ653uNUnPCukgarV0hX+jpncBn2k653i7uZKL54vjJeZnMpnrB3W
+hTETB0VVVYHwRy6aFwFkp00z4FyRdVugOrQrBedtfMPIyCsi+B7PkkSvzD0RcCM2jh+L9lKU3CW
RH/7Peh1V1kqUXyNo6XulXd0xFE1Ypligsn0S+nu3sOv6ObovtHFlqU029br7vDMw+QbFQuLT+ep
3YwN7wKVD0kSkgxkbUAr2I0Ec0EkMl1rYavyKmT3dy8oXJcRVnx/+wVVBELZYGy+fa9hZQ6D8k2A
qpR8Jdf+KwSozqT3GO8+1Z8HmgoHihpGVJ/L76o8BO4n7IYQ6X3xfLbw0wq437NzxczoFZrdqGae
GCtBK26UzBAGNq7qBJ3L+teIWR0C2Ihb0RFL+JS3d0rZr2VQYe3g30x/vuOgyHud03o9tyenNSF4
EnbWDGy5HSGi7t3Hb6hSZ/rRPqBYVJRb6NjdTwfGbP/ExjFi1o5bAxLgOH88Vjr8hz0rcQc7KyL5
/lLhaGtqBJGNf535KF8V9FE6LKJm3nkAeUrNcf+yISiphrGGeg/tVGt3SxKZn9pWbILm8Zo3shwr
3jZymVFfSFe7BOOOgGOcsJD69NmV3nsuMaib70oSeqLUhhwEZ4u2XiK7o+vUpv1YgbXNwjf8aLoX
DC7rpfluyp+3MbjmRVvAjXWFAPQ0Szsm3Q5KVmt6rPd9Zkyaf+hgzHNDVwhz7gppbrj5rGfmpACn
a3a9b7miyrmqOuOLacNmJzwCCp4JLA3JqvN9Nfw7rWzPQcpyLFdRR6gGmLhCBbv0CNk8NfnDcg/h
IIbaQa1rdzivs1hhN02SM2KPbgjwxMTSf3H9fVyQpltfbej03bSdzt1VK6iwJhyD4X39iJBMoQ1C
A30hH6WhOu+1WiXiCoKQRzz6IlhEtnnSAyGavRR9Og7gUCY5tlcNeRDYBEuZ3kbARNkA4D1G6GGq
0t7vzpkC9/JNMo8rWoDa4BJ5NMl8DBwjjZgpEstFgy7Ix3SoNbnR51irh2d4RPwaoZXafq+sksgJ
iPAtLnnPBGkJgDplzUarT8VkJRFUyEFRkEPKwZwSAXufyYz/gU3q7wowBB6mHTO0EQSCFvjsibAs
VA4D6B4jhQOwYW4YZElID8iKHSRK9yFigY+6Q8ic7GuA1jQzngHxouMgidSxknXx6H/TCo7JlWXJ
5f5ykOjKsBAmWnHCiSCLREVP+wITVnr6Wv8mJ+GvWDjP6ppgGxUpiE/2UaJ6qBwoP2uFefHyW4MA
BrNckyWp8kN+GlShbZy/6nQBQAEITYhDleZ/rzwNLhApnbXeFinwAxD8enm9TNUSp+nlCFzMPT6W
YQIGZix0rHKodyZfAeXrvlXfY/33Az3vR8Sw9s2E5kl8IB4JXd8QRF8l+V1wRedp38+6sIAG1dcK
Ml/GU0BXgcHND8h4twPh6DKQFXkrDMFuPxV41OHAnF9dDEIfflFaLiytwuT1uKP4XII7nuwWdIaQ
Zc3GU624j+NedPN9TGPM1mNfPc9WvbuCnx3QB8Yfea5lTQnQoIruplk6pPVArRbmMZ9FI6qOpuQ6
3EN9nY4yvKUMWlD2gJsJmOdPenOeWQ0gYf97CTj3jFfyKzCymHqpXoWPgTEWOH8z28uYBRa+bGrd
OxQI85r906Xmk+LWB40udt+EL6KcdZSQL7GWrFlzFlrzfh38x4NcM3SrObKqzhm+2y1wy24l/4l2
tQmqObqwYGm1FIkeKbbUFl3/k4dobQDCAVD0CTuztU24nrFtb+ZK6F39RhcIxow+n02vnK9cHQnJ
AhITvFToqGPyDy44RwOtDYYG2qWWpKawaSfhV7xVIJp9YIfszM6ybwqGKDYRTcoQ5GhD99149RGV
fXQwEGSHhE+n4BHZvSeChA73Tyjdqh519fRjHm1w/RhosRDeoZGZ6XMcmN1huN2NhqVX3Xm2mr0W
UljPcxM/oU4g2p3j1PhsU8kKzYOU4VhTGGqhsZ/TRtAOlWtO5AuXB4hEB1IPJzeSfYjatVOcrjf3
0wVKy9C36VWFZbqksCRfe7MuaBeyYGsI6zp1zb/TED39xB9xTAlJePGggPTo4A79HjOdhdrIrKCG
jFbMG3+03AQe0VN+VcbPk0eEPDLoHwRhpLrHwm237Zc90C7FEBH99eGCEg58XHtPHaFwBeONQwx2
Vh4UAc7WWI4AXOeqI4qwg5M6g7NN52qvlmBRSqYm4W/OQ0GDdb9JiByvxaYfw9BvKHspy7mNmNfT
QLAvkn5Pf9eQwcOsY1DUl/00u0xR6dBKRc9S/m1eeo7SvghOV+l0uWJUmLSQ39t/oDcp7gx/bV9e
4RB3fJDRRJ8DXrI9bcg+RbAZA+V3TwVPC9lVSvn9KLG/uGOce7ua3xF+TqUIiNf3nuqV8R/od+WC
O1Bp02LqUJwpVjVoVbCGaW9KqLKiiK6ToEGoQyz1YGHBuYb11v2tW2S5SNwbx3YTaROFmHjMDeiV
xezi3+k5Hn5hDWCTA/2iin/lPSiSZomnzoRw8fC1iJi9yclQ5jBkXrtLOAd3bHPHH2b013RTPdDU
fDRLmDn4UNPxdDKqGWfhX8r1+EMEz5rmSiFTqg94B8ghwFjWzODlYlQOirBSFOmw6TV7AhqdPW7p
CvcLcJBigyLiTkg8E+tkyqcPBt2+TIhXXZmPhlI3f+hPwyi7IJBe1pXjx/vLOm3jl32Bk6PDYxrU
MlAEWYMGQmYf7HOeo34ur/vcsuwczLWj0NIHjNAWgOrwv9I0arFznGqoixz4oP4xVdl72aGLSav2
WYq/7sC8wSLU5cU21JPZo4Dg1MczftcmSlJO3YVSTRFAqGnFdCRHCzhnw0ep1HHyWMj3TQ7d/37g
WCy4wUzTFd12NuBweAubYb6RfNM/99nGZxsTl8WBcJaMcrBldPhVPCGGtZbsltt6aay4xseLHnPF
GoqJrRrcdWXcYLQFsjdU2L6u5pV0F4XYngENcHbKuEnhiy7rFyhb49J95Mh8Vs0IynSS+eWLR0QN
CFo4ugNyyCQ7Ki3IQzA1TKOzLK+XWQOw6Yy9nTj2iqGbyB8nHCjW3wq79CbeEH0Ke6CZEQsZ/QBp
tjcvVQ/LpHbkxdm1t+rk6Pji9aIgMTp4yq3NyarDnITtHk2N9FvvPj173ivZL7Zwq8+slqmdJeEs
MiYBdmuWg0tEA6q6j03Mz/Aj/gHv/KyoMvRXUo+LLUlve2y6YKC0v/QsuMVXv27vJn50Ou2zH6Z3
62P4aPF8sFJ9HAHfe+P/hdCtl+dPElsKt0PPx3TY1kUZIt349Rk+PNToEWa0nmLMUaxKnqzO9kse
nMFbZCmab9EqiLNQEOA8HDPYcYndLPYNYZdC4vqSO9JTEW/6g5XM16f8JfjEO6Jw/FSMxmdp9V/b
zbu1pczSgV/x1MFVFGh3Gv9rBRDnyZXYxeM9N3+eLHPOHAGvYcoD3tCqJimuoEAxS3HUUCNQq3+M
NETEy0YIGjHVQk3+fuRksHDU8CZ9TsknCm/wlyAA4dEnWVmAKsyTrr5YvSUFjlhGjunQVOyF9y6c
sbDRHdY3yT6XVJ5Gmo4OtT9axlfME+JITkUcWWV8USACK7dDiMY7zyVAog+0vrVlH7q69QaoCI0X
DIjXFxrTaTJeVbdoZORbv6jyly6lrWEFB24SeMvyLxXfmrg7o6gN+obkDEta7J6iFOjaETtGuywu
G1KPthNljgfJRqBIyw9rlqYETrTmyhhpl4IA5Bx4d6GQyZ88Jq2j9UbsWEb7088RRpRyg66HadPM
CGAFmbuDIxb05I2SBakBuRoIUBjd9r4t3V6rK0NjJL8O95Xg9xStVNoCUXqiL2A5UxMeNtP2fb3e
b4uOkqMP/SfaIt/LLHWudUMxCz9jaySq8hBHvli1tHsrw8ifiKh54XYtj5Ba2Pr1rH6mmuQWx3nl
U7+qPivXJn2JGCjIOGDcef8XhcxxaCarjmdqJZlYiy8/WSMfHPLZec/D+ZDQnSvVaZHQ4+/xUrHm
BjZ5JeB5UoilAGxerksbTnFuIeLaRIS3SdG/iXj/kawWuj0Mu7h1OclYibGTQJoa3mGq2uL5F2AN
MeeH2s53AqsDs9nq7YcE8iT2y1AcC9C46jqWZd6DqPyPQrDFm92Nj9lSjQaGYO4a0ztN2gLHgvr2
mvUx1eD7X9nSUTWd/wEH6CMcRuiKdsVLUVbWz8QIjZ+8RzbZBTaYVMXW5G1MdsOqWDFhgr4gwsRX
kInMNi6ptraP9a1hmrrDnKy3Udyxv/0WnMNYCOdoOQLdm0gqUHRGAoiQZoLOtYvTSYyN3NkPMilk
uT9vBv35q3WTsr93nhGpW75Q/fe+ECJsWHjAOTToi+Fl22cnfvhIKxnwKHaJvoMgYwVqV7g9yMKY
HxSdRLoSZqjgGGr3BOFAMSupeVO2bP5CBgK6EdKZ157tR0ck/F00S122I15fDqqiWV2MmM8SBTZb
Esb/9CSVz5F9DKfIQr/Ckkf5BhNAUBa3B8KDJeZD818TLyNJT+MD3Msb/C5kkCTJcx17JzxODM7w
dtFFa1/FkvbWJBRmjltl77egw01bcOdCb9k/WHmTpw5HlAzQAG1+3quBJEK+yG0CyzK5t0Jv3m7N
qAYBcsFOUYIMhKyvoPABeEgwA5UyB/U2cbat0YY1oMtMwxPgDOt1NxqYbcApCo2pP73H89fBEX21
hBOGFI2YbcOWqHBG/oph8W6Qoft/JYOzGKn9CDMlvIXGjLq3aM/EDF2R0yKkgD36ZtVtoSFlqDMq
5oJ9VKlWMVyzxyKwEG9Cdy0kglDn1DNFyesN27nta7SrujBBVwP8Y+lQBXypr3esURmv8KW/93nF
qToAZfBuJb3yVGNNrRwpFX6kx1+27QU+yV5qHId08gwvvfqKkvpMk+UcnQinz/e0vIB4wg4jipXq
NT2sRftBIjoqkYTsyzOadA5Jzt6I+lK9PA+n7oXolfpTm1Su2t0lxpinVuv2+vnM0iJqqTJ2nstY
kTzHdVkfNg4i2sxxX9BHGeZZRJc9xcV2/E9JgYl2gpFTlL01IY/DeSr/3+1LkySY8Jse0TwT8/Wf
MPEabXKRJ7kx7prnjKgf8c6Bq/mBkqxcoVJU7ErFtUyQ37BHpgW8BKgsI2Skgz2o7eq1gPpWWjJS
YDzNvbVY8ReaP6ak9/x6jbEhdu3FlK5DrbWWNR6AotL/2Y8xoCXw/d6sHVtUsn90isJBdjVhaSTr
Y+XjJSj2z2hin11fOCCULO7Mhwo47fryQtxMwKCIx9CXuPp/luvTTNNc13YNMhVmZCotKwyt3dQ6
VTxuXfmkAGRn3Ec/KYTqRDWHFYVYLuGvLFAaJPWCgYJkA/q1PM9Rupxlex88GWiT1S9782DUeoZ7
iblaqhgJqfYf5PEElrLJvzJfpZpuWz1U7c9GXuMu4XPBM0GOBXbehii17PR/aiUtj7BE45ck23m9
Mql5cb5S9B2z5qg2NIJ1e6KSkbBz3YzdzcFjOyVHoCn0iSNV1koEZxfzFhAfXtWZRPT+FS2To3c7
aZVS5gJ+96wWfV1NchwKFDlK34cp2lG2MreWQ/dEgffCCPmnr0506cZb75q9iyZX5mJn5QY2ksVe
KqWoJJSX2Eb5PeU/TVYbNNvBkQkNjCZOh8tDZ7LJQi+8xfGMYcYGuHkQjjdrHb+yg7CWLPuN/f8z
aGijyQ3H0KkXiMo1YKcySM0gOR7qtfSKaf0ytY7SIfu3jGG7qKnIYXmbE4TUZaXScwnTVzcIzeaC
f/CsF+UVO1YHbX9sqpYV8OpZsdD6qo+fKjJsowYSoN/5NbLvtNdCHNCJvIiYa+8TYuDoBC77sb4o
RVWMilXwqctBTiESy2PTVJbMKH3/hFCdmuTB8469laBVXzwMyYyVJaBmlfxME2/dIW1TKtBfmS8B
/7PoZocJ3lP5Fy2t1yVphp7fpncXFk7JA6CG17aI7R8MBEVrI3vAZDSvwj2VxdnU0a8FyzgCTUih
i3+dxgMQHo/C/XKAYgHqQiPJMxQomINkk318FScPHyETBNKQMzIHKh75acjukBx30HIiY3/jRMBU
6JtAEEl+Prls641FiALxddKnPWB+PBDw2t2PA16RWsLtLr/3WoqAmaaJTsoOQDEM4FjFB3l6A4Q4
9DiB1QTJ32lNF/cPekbTq2MNN1r7p7o4w66aXxLffR2T1OllPlay13j5ggKPHJHSvJNXtfB3DocG
gXIlivpM9drCqt9Q5nSWNv++0UOjd0FTpEcOyHoKG7h6rpjiKPzPzHWi0DsVQQDO9eNLI8gzJYBc
J1E9DLl9PPl5LQetB70XIAx8znb2iN8MXskA8/GqL8fXRQwRt4hsjKABpL4uuuzDlzfZ2xL6vUQY
J2vGymdwRfHOZ0fOvctLkOCFUNhlgXyqIJTauYHbhpthX85xaHwmwJXwPOKQFChpp8y3zLQOoPxW
C6KelyhZJMM7fTPlZzSfM8Au51oRsN/byT3qXbJneqJLH1pnfdc7QAR66bTiEyge7FqBrL/97k07
gagaEvEbGZM/VsKAub8gnREcglXS6dbwj9tNRv7B8M82zZpqHh+LKwugNYobjmU8ImIAenHEkutZ
68nhBnW8aPM2myzJuD50c6HUkxiRoh5Dmac2VjTNGMmlNXyS1Cefv5mUEwuAsNbZif9TwT3DJgpQ
TBubGT3c7IbHTS4WJUu9RwInOYJy5lP5B1apXMGTl0gmN5/51Mj4uFKracqVq6/Rop+Slb/v3bXd
CbiCgedlYpGq8JbU4JJt+snze0MN0ztRb1Cj9Noh/YJ5qldB0StqbTXlzO4n6lfTe3eNX1Qrspwf
iwnwcKfktq+wOjLi+O/G+ksv94DqIoxQy+sKq2qnhyqzyH9oATYtg4X43FoWwQzbwPk7zV7+01/8
uhPQN24hlHSznrw3TAuqipRb5eP/zpecVXUxBo5gGl7PbYpvQvGMRjW+DhoGDnaIDIFRN1/gneKv
dsCpifYXdEfxHgr03G5Rn/EltOE25IoguoDRxKlxh1tl6Ug/uAOVPIU3JTFmPnJE6tBVf0t74Hua
Y6Lv8HHSJmaQzkzT2S+uaV9AJrZYZQgnUgv7lpthA3hSgmqqKYTQaWveX76hTCUE90l7vuMA35Zm
d+kUCBeq8k3db12Vz1yPruh7bUVg0QvLbzV6iiLJJdFrNUjKVYwY7Xywi92EN1GFc8dol3qm/0+E
aYCIcg855fHj2vIwEakdkZnP7vsm+4xVp4BOSVzE/fhytUGWBRnDtJCzl+wCg9CIuVPABjglpDar
FOmCOrqpcCLrdrTFL16aVZMLBdoE6crvxSwaM+R+S/kgQMvcAEl82O8d1XAorbsDpdCoHqcHHCaf
kKLVvWsQwtC8rd7YL5CDTpZ8Wh9BQSFkAb91+W5Mkr6WeK0Wb+bvqOoCm1mTMp1jaY2Xoshd0SpO
esFvXHd/iOS0POoqlSYM4aLMZYLvHxHJFen9803U+J544QNby4gXWEcy+sFRaAsb3Dlf0FkPMEdQ
7VcY3wqAD4X2XJziMX0i+ZGeE+IooVYpoYQS31oyu7RgRfM/5wI8FsJQp9gpWiHCPSfFTpZnHJnH
r4eST6DV+cUjQyb1xfcZOnk+jBWCpKzUj0pEx5lV1BcqRBwDgS3DIlMvXhcZvqkD2UjzUNeGXQxI
J70FxEsHu5iKtbxM8kZtQUR+HMIuUmMsGw9OU8lLQAZV8g2qqlBVf5nzaEhClobD9KIvTN76NiD7
0Z/I+lm4UyrJ9u3Ivktbj4PUZSWpv1C3Huaz1VMPVB2AwdnkCR8iimmPN2DBbbQ0NkV8cfqvNAEp
VuprUFt6nDu1w1z7Vyy8R2EcJ8uHQBBAXMJgL8OkHF517xWr2XNxSalFthA0lbcLk5vYAq6MRY/D
MPjQIjozBk+9eqvV9SzhtzyrZLGKa6yAZ6KQcurQAaG/hIlQtek2ljNEW7AqzAeyzXuQ7Gw7oCmV
6+eG0HUTRLgXQmn92ZyMGmruLueP6G3D3vR/I3weUP7WohGYjuytR7WTFZFwr+4CCSCimqpFHMUK
roRhL4WJblO+NHUu6ynKoxFTOqjeN/Qpr5yPBTZSmSkp4xXAAwcHojcBwGXPfoOpWePbnWQKF4K7
KB4UBN4uhiRvuwegDDUranG1hDsEtszmdjvsv4lbQCUSMTDq7mWDJhiHkeoJE7Aqz+953cXTWQSb
Paz7VCDW7dhV6ismHS6RVmsdGYaxESEDoXTPcHNDkVcBfgOnyoNSz3joHJMPEW5x5dTRgRxdHQ/T
ylRvRb9Wb3mAEj0Ib/7FWLWWDTUVZ/PwgzwXkBK4BXrl2dSEHMxq14zLHuyymU9N/2MDn4+kdnCX
s4JDDTHmbd5TkDSLjfU+M9wAtrRxZV8cQ4lZWlCfQJadKjVwGmgxU+NOJZyDMy4/tWAgiDElLrTa
g6SlkN6pBtdaDkMPDzdNFCcbx6zYiy35LEzEX5yAi4OcqHyU5BnNyNV5CaRngl4xI9sAEbuEIxoh
Kl/JJDS4dIOJEZX3lesZ0WJwi92LjgTe799BSweJXz06O+brwf3xX4zgjzf0flJzmZmUgOE8dgXp
XUWLDiTYLFApF4WtXYXG531OG8r0GL5HAmmZo0IzFH3pe6XCG4UOVJvMYlbTGo3V1YwcMbzk8+dr
s1SLlI/xS5aTaoK72QqsAA77r/pB/JBJnsX9bTnHTVZKknAHgH4BYPO6vC7fAF6wCrMG0rwXI68e
WduDzJSN1Vsy4j01oTIvznanXsLOQMWaTT1tVgVHQIvfFmTEMjMq3f8skclZzKTH7UER2WGqaNFj
2SSBlhH1u215CLMygIIblu62cEDBntGcdNKougATGMLWmsB6Q7k/2Zct7Wwv2uacVVOJzGvj0wyO
xgoIH/nQahyCN2SpZ+CdWwUX+crotYJ2C6PChk/QpV4WSLSv0BFOjn2cIAZQlOdvdVISliF/c7Nm
Jrq07EGs98yGxg6ZdizeQWryMtXm0aBOpi37E0+BIr2qoIv8lTQuJW6r1D+fP7MTyJp8b5woqVSX
cEUHrm997sOiQC1tYhyF2K6FEoz86zZi2nohIryN5LBzYz7KzXTk7PWDkxYZYbGm3dd4KkOA5IoR
krbrct8isXDsURklB2hCsTBQ8QMliCHcq+yXOqVpwBhJhx3g91h0tK6UR5tX+UVG2kyDwyLgs31Q
VRWF4Gda/JL9/RfLJlWb5fRGMIc0mMeNip1/gKMCfhoPBhwbar3qGDnw09uNNWEAgDvca8PLhAaY
ErUsl6n8kxogNJ5+i+zGVpuMxgCoZ6lTjv55YM4xzOMqJSdN9FfBq7Je4EmcjvORNoAMjLiqW4IH
17nm4W9TDFKdnezydaBZ5UyGJI37SOej5cDA3VINFaBu+lGrPK0zyQVcNu+QoRli1rNifuX1w05Z
qY0DJdFg8DpZIjZAwGNNEBBUU+fItAOEIN1RpAVBMpNzdjCssABKYXChY4kh2ApaaRsFhjaUBkh4
HcSHOj2qnSFt3Jatqd8xrkenigZE/8pONPIPeLJ8aXbgMg26kmlsUiA9rOiqetE4+QfygFrdH7Ge
BAaB/lzoLlDvjiyrgb2ZvAaTodQpqIu23+gp9kXJKR0sf6VOoV+KcJsC8AuTb/nWGKVv+mHSu+Ty
gfyEnJ7y9HN09aXIzZtRttoA27fi2oFyUARWr+gKvIhRGje6DiY3iRWD4HD63k7ZosyB3/8H/hLM
/8StML6xvEF64rz0xdWhZEtWEXLP/u49tueCNNVpYpykOpKS6vfz33yLkjU7vJOwuokRvPjCQqoF
4L7Gs5XkRzZSJyo/ZTQCkeSQeMH33niHHh3D5jxYmw4pktduvjHSEvFTMvbffrz9/sWclMITdwxA
ZWjilCsQ7U1L2AewyTLfPfqPJzDnLcy42nNhfL4I1VJ8stYHG3181R3rvTuB4375ExoDHW+Ja19F
TC25ME8fCPvLoI2I84RSJgRJTExeVQfPvVe+wb9d9pQTcWnmRfWEk7aFvfFNXvJ40mA4PkxcJkYs
vBfYJFDHa2CB1Xo+KYEAF528Jjevv4TMuONyo2M3v40ddEoOiwplr4PMN1CkkhJvInVy9Zt624c6
DJb7xGfwSpSuWHiyD+LmCT75dfTMo3CVomxDSyfH/49RnasafvhrHdBxzQASymI27Dww7dJtEmSv
KaXwzICGotZPd70NO2TodaFguo1h9AQQfEpfTC7/n3eKE0p2YPlnnLbYcPCvTBoCH/guiRiFwcd2
tojpG/B8Kb7MKdOvLQfhC6kh4H8hkfxUHpUpymAEM3fI5nClAlErKkIAaJMslFHIKl6bJ2CAJkDs
/pRMuGtUTOpLnZcmDFEvtMQmJMlEjC5Y+x1mxK+VYNL0KuXLAoeBxaNqbcR72HQ9e1DTXblsRym8
Hvidilgwnc+7RXdcNvLGo8vCPyLBq4F/KBz01cJfh14Ow+vP7ax7zkn7Z8Dy1MWylDCLm+k3BjQ3
81cEiBMeWVzHys4v+tMe81bkIKR7V7hvNOM9sn7rgq/bBq9f2wJwydXHTvX4LRnxZHnOTS8GpbY9
/ljvCPymV+7jYqXLa1QesiRPbNMuD9fmDi3adTvF6r0rFmuhzvFte54G2oPzvrUz9J/6JZl0NtE1
P75qDgyKZtiOj4/aVO92hdvQg6zhUB3aEAdsK6Lc7aNlAej2aJAjT9ueKYczP+2nWzk5CkYx0rRH
Reo97stR767pDa/Ie6o3OPuxDLDdexMbl3SZTDh5pQC7sxsjbwtAe+lqi4c6h2G4qMxH8zbJCEaC
5GDWD9VxE8pvdRqYgbX2Ntzf7gkHoe89szIferocw3AXbZIpluTocDFKfJIlNeD4b/PeFEWvpb+8
tQzTOhjrDzpQXjP3aKv6VHLn7MhWf1KxmV221FuqxQxO492QoBDzasRHWp9MncL1M+x8AIDeh/A2
StE9krxIHmrXzIIcC+d/PxduIWuL46O0y+U9n/CKqIj7w0B8eCP8quqOatFzXMoLo+xwkND1/ynh
oRdkIA+Xk7yJLGYg88ghScE2ijVxnd/YDqKRN+KiOZrxtFE1hH+SWb1sALRQmp2o9UQkIKlzEC/c
aX2G4/2IQEMwJ/GAdLG8p2Alfl/clec3A1oMRDc6g8JvvtjnIpvvLz/ZpgwvZK/YFjWv+lDJlJk5
46J521gmBTsdhXZHSYqyKmm57URhFJGeaHE2PM6nomX54+QR/9rlFLWmNXS9GZWobDo39GA8C4/g
C8isoBjivRz7O5NAaTmFwiHwEtghktVQsbekUNJIYdZeIOxzcuv9rpk32hz3cJMCKT9NWmSE0PAZ
H4jg8UY3RNGjQBGUWHdp5xUh0f5beFHeYvgTOoxsS2sXALH4r1RwyZFJuFCOcajbL7BXRpSKVybm
da/AOw1yjtxMIcmiD4NMFNf/DMfD/L6kbboJOC02E1TgvZJ6w27NRVa2c7ZUf2B1gWSh+vIsd+UA
UUCJW5Y7wGQBpas4ZvliUPPk/OY4ZWBjGjLJxhAf3dsG12StWIdfg1izIeaCTDOPZxduU6SV1ITc
UfWAS0nk2kV+TG5i+K8ox7klCawsJ1z43MKsuxLcYanl1nsepgB64R1lqfLl1/NpiU1AU60/DW0r
vDYN7/K/NSmTXR1mU553Qa2VRDZsgGBeMXRQVxVz+GIsrza/6mYt8EZgjUMYZmAdG9IY81AoSTku
k2fP5BYjUAR8VlaebL6f26yRi9A8SndREVu6stpe59UF8A5NsbkHGCrc6IQRrd0H4hCljg2PfcT0
deMwY0xYlOImXRWkyopI7IjgCXRyZmo0wdDjsOdvMt6OM8RpPtNHHscrT5wH0vhTP0Lh8YhO6llB
HRMMWLeP8K/KJG6J85WkkOQDz/Z1ty4iLAwv01940CeUlGJS+8eD2q7gu5KX4qN9j3h3vp0lrDYs
32MRyHhkTxId3cdiRPSREXxv15OGxREJe70M3szNq05U1YWecWhnTL5ZjHGJ1/GZewylHaOUziEn
K+ZrTsLQMwYjaV7fOlzdySzPnTMzW8LYUWRtBkxB86IcnhrsJiNv1seV8zUmbjxcOxAIj/uJmZ5q
/o3mMgiATZz0zWg1/aoq69sM7tSiWFB3Tb0ehlBvRBgW/jU/FZmasaINyRDwOu6m0RbWjaKvUjSb
JdeEeQ9mXghg14ThpFepJK9fFc5WZtAKWphkjNq4Hau+tCcp31AhSmjogxkrI1lF4gSefOsR+/o8
iNQXnF0j/HPynI24yuvoYlM73+oKox2eZeBGAzGrNzAXJTbF1MSLSxqqDixic4AZ3o4K4sJM1loG
q6KFflkPbH4k4OQiz/WSUr6EKGmsM6NIc9y+m7+/CVsJ7X/22vMwj6YHOrnnitpqQ+S6dLkiEaB3
ONmECQ/BpMuKlL2BbtAojKjIZwI5s+1pqAwCU5R8MPXAlaEiCVeM2j5thjPDbAh2r5BDT3Iur/C5
AdicQvA+LrFl2eGZF2QtAFffZrI2nC429t7jAsU4RZIQoAwf39YopoNg/LH+WIZ46el6zkqZhJ4U
DVrrvRRnjbvmIN50nOs0E9Kb/U9z+guPrdUPDWfMsimbpIYEgFj2Qcgya3flnRk6gLmf+8QsQOev
kfEqsWFfwUKlGiecZFYI5GMfEHbkKnkowiSWx9MCP7xgnSz+sl2E/nM8FdaBbcNCmaGl36nIAnVV
oPBNb2nj0gsk4zHgeYJNDW/sOFaxJRNs4BIytIWVLiwG7bV7jfzbkobsrt6+rloUEvN1i3lsXuBA
dJExaX5CcbM3ZMcd4rr45zOkuohFYXARYu2OeHHChaiInQgQWMP4LzbeHynmwXqoIZHz9Omu8bhR
FltokmMI1hmoiB+MgtTE0095YS5+uXe1OQ9p8PedqivRwoREdxkEGwhkP2Fs75W6bLuHYx9G++lj
8sHMBOK95xmrj6ccMnwqSRuQdLrqN4UEzSZjCK3FLAFfzZod6KDoensd/n+HTCwE3/ieDLWDJS/j
CqS1wers6oYYb5TYKwZtAIoZ8oSflE32Ze5dkz6nS1gY9pvcPr2aTTLvrXXMQ8rqlERulKjCSo8R
kwhsUCf9tLdX5I3yqOXPzxu1DjeDa1/BNeQgpTa0bl8svnCo5vqKTadofpsopbVpaT4L6lzwAojy
YyXZxEYKjblPT83jfnT2qOqNbQMmtNbZ1uWAKudDl6xnioby6RTaW/IjmUroRzPZOlxlf4PKFXSB
cfnOTBnwNd1xFi9RqIcN0AgKn62pqnWPVhCUvIg4+3A1bpJyB0vov3mH7wVWQKh/n+GMUTRLl/wu
DKxx38hiGFF8/O0epP7tX7r1EwpQA64qTLzYIwwN/A3xCvTVRYy4/97KriRx4d2eBniczxTROe9C
LyGzKZmSHxQkZ1vHpM0vBXuKnN5mhg2wxCwrCBtVnN8jotYJOArfZsGUtpzgccJ8vzCba7jWwvlt
1Wdp7vqoWo0TpaWhXrNK33TAEQKraOwzemt0RSuUZE9qNzeVh5LPlVhgvOQ6kNgAyddkYQCO++RS
1ep8rh7ouRKHXw68nF4jgIV9/Pqx//7RVHo3CLUi2wURmhOm0ot7ZyGJrPSgNgfZAXqvxb2O9H/B
z+tZ52KT3mo0+sGvRsXTJmZzSun93fHmqAXA5LyF/Q5gxMjGE3oo6Ho3uCx2Tadt7276BfcZ+H/H
haF9OtmtIhawU4NCxph0EZ0zL4oT/UObV7bPtknG2fpWS/d9lMLKVhKEta9R4jgIi3Ps73f9eXjA
GBTsGsbE2VoEA2AobYUOU2yvLgAWdf0d0ivlpawcAK0RP9eKjDA9HUsmEFeI7/qrOc/BQy2DVq2q
KN1UZBJs3rOxnF96WntKY0oBwAceie57J/8XXWvUGG/DqLTlJckOG2w3uIZi21fyQ1LnrahMF8SU
34s6izOAOIBIss348P/5Zb2Gbh/e00tBIYILmd9VQBL1crwC4HFsvJUwrUtvdTl/RohhewOS1asw
YZSQtm3QSWmDOrZz1LnQF2nYbaA20PRt1xUuNAQCzWeLC4iGLGBzF12Hj9yM7Sz52YNmtx0HvNLm
UPpyJCwbQmKYoIm5Zdwuznz+QD3shoxk5cG/PLzQXd4utujjXz+1qLYkvtUllLhhQPcz9jmkHDyu
0Dc9T3aE0/rhsR+jwUhjibyfch1r3X/bPxN1Io/xvN1gImuwi/TaoS36PXCV42sMQ4NaD4I0xHF0
FenR9WlkAh5apyXBnxkWgRSkm92X31GQdwSIuFek9UN7++pqO4568Pe6i7HU7m7emOKtgeVy/oAt
DUemFZBaQMzLi+uUVZeXaqZKUYueXwdeJWXmD9wirdR1oauJ8bKGlrWqOCr93hKDaeASlAncCPyl
KO/eKxNb8LC1I3JEc4iuAhaQVGw8T82lZ79dVoyAEK5g7GEuiZezCoedmWockus+tKEZE3VrfpqD
YdLwbCf2ERF7BxQt96TVDLYG5qVM5lD194QxfUxnAQ3c9YwLUzvU7kdL3pckwr+TQkRTpSgRvFuu
8tLDmKvvuWrtPEtvmEPiM01qjR6ocV8GFygHAHB2TOo0XBZmwNKpZdVbZHdxCq+Dssj3FLdtdy2h
byAB9h3nu93TnMvoT+uUeSj+nDv6jx9MnT0wWnIfGL/6CyxdJqtIExrd8TBJVfakiDJRZr4kONps
bVdJKVgCNeRUu8gC8E15yHFlZBFfqqV+ZvQOSobMta+6DgctvtOlzmGaz/SKc30hGMfnRwoLiVQs
KDitnbjMj/XNlCes4hxP0nn044/ebnWkvojOSOlSUtHpOpVGC8UB5hq4XoTTewEPOLfOmaC6Z7zW
9avAO+3mGeEEKptUf1XIeVpury2uyiMFcDNHWmRHDsc3GxWeoSq4QLPWpEPchXJ3FWIxO8ZljdHH
fqAqYutRMafzg3j/xutGG++rKt1+Nwm8uMRqFtOzLDWijGmuefcFwEp+1W9WjTbQtrwdEJI7za9G
OO5R+LE5javYMYdAHfJEINBNhOOJ1nhftXTB3mBnIqhXoMeSJsT7mM2im8Map3ZZLFwjd0T/iGTS
3xcRUvdYCrADMsmi1r5j6bpzMU4fYozbQRd8xzTSBjV4E20MtIot9RYs15ZVu5CakV7GoRWzJ9da
YjmzYZ4eWIIwE3qTUbbtksdPNR00aU9JxHAuOpPlrHzgwwkglkp/troo4KCGnHDlhgcAJ+oH7Vhp
06TnECfAsF85bUivGeVSRtO4K/ntNBipf1JGF97jhBLXgmiilKwhchzhGA7sjKdtJ0EYRMzgylym
rNQz90yICGqcWl1T0/C2AOukd2EOMfDdfpsbWjEvIrIdyRL3p/RxcdUY42M/mgqi9PwVldu5MJ0n
95bDpHhZRmVTMcABuD27OSPjFMzvkT0zv1gNeMtmVYcSwDwt/wJxs8Ou1/rs5xS2RRhV9TNCu2Qf
Gd7ENUvvx1lMLS+0zuA73eicFzFyYOw8r71S0VRUXc/aJTtwrVR55u5i1SnNjLOOAPVjsgwNcwvc
UF/7TYzXaa1iDmoNBRM5+PV6vZEuk0t7V6PmxcWjNrxcGh5uhuHgUjaIoGU4Q9Fd5YyRJ02g+ZG2
CJYGtPR4lHp/LqA5aZwLUyeUHwoyVbE9VJeHRFpuiXk9VGqz9c+x498lcPnv51lB/5WuOKAud709
T2QRy4V7cZkNGtZEwjqiCcXUk6R8xMhzsq3oJHdXzglnU9kVAW+aKS+NpdlEevEaomWAIVkcQt5j
BFsSlsUacGHFKsHmYAonrwbOk6dR29AcdqR27eWPIoMyuVzT2onYjZW5TYelLhKt1nALs9FLtBVa
d5HTNvvJg2Kmm/jAPZb6/44q27RJh64/UJEFZPJH/sy8aSwd4zVyBQCTU0POrVAFeWQRS72yzSam
BZcyjoMUdBVvcc/vXldnjxYBx9JHCM1KbIJPrx5gRu7ahn3/VCbhx7vg0sLFbHW+hOXul/yYxxgN
vZWF8RG/Lu5aVHxuFW5vJRV1dy4/HpSS3ZXkAZmAvOvjuXWXI4bY+v1RlRShLCz+hidjYItG2si6
jkCxGqx/gUBpVnNNYuZy2RI1JYj/oQk1oi4w+x+Zp/FZBXwjuHr0chGR6Ziopi30ouE1VyxHrbVs
i/CCUCcM2XnIywhWmBZJEC+P0tO1/23viPYkGnMVNlH/f3NExyl8Hwl3IIE22RbZfs3gvRtYy0iF
0VTWQsboBTOx829aOHXdC70fqSxUXSCKTlfOSClMNLki+DaboBYYjcUN36yqTtLWiwoUBF51RJ9i
u6jB7keb+pLawQHzkwSBWhJ8fTdNM67mVC7AG8nhFRdCSR318Lv7Y9LwlkJ08MLdGgd14VGwHCnQ
3r8C9rxBmUwc8KHbE0CXNGbakywR84/b/zQ+MdC/llTff8ff7dcvYniumhCCcRlSCmGD1nGls3k9
a/xOjeOPzAFjwwclM2RoKl3+NqMuQQw4yvd9P6a1+yYduy/lW8FJwDom3VkfE44GMKCUlhAum8NZ
DokPzfoXJ//ZYDf4d0NFk5PWlTtqP40ixYftOVSQbgBRkpKeHeXBLhfHloAlue/Anj/NSyK4YVPZ
G5h5aMVVrFIVBTzM5n3lmN7edVQftZDr47ywoRPMA6CtN/pupS5LaoA5YYrEhCzOJrKd6KmkEj5G
2PxhAvdUPohAcBWzx5Rd3Txps9AZry+VBmNCwDgfMhngC0X8KNfNEZlBoRKaSq/4Zjd4KMvYDmWd
FLF8BLU9FUAGEK9vfFqwp4lk+yoNEw3apca6v+wTOwYO
`protect end_protected
