`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
lpDxXkCw9L6rcpCJhcWegT8ffQAmMuLBLm2dM4ygDiV5xaID4ZjLvX1gzu2JtxIUgIwwo126DUrv
0Ne+AiNQkA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bI/N/TOD9DQj44ah2pqbNlWUTmcBHenKI4kuZsumOj22FBxyynctRM30nylXtXEFzmnuH/mKbDKR
zZoK/Gf9jizFGhlIThIcXkVA4BeNYQ0wbSNuruSl5QQkKk23LpdjmXoRWZZurr+LUa+KJ29Wn51S
u6ybbKEB35niWPa6qkI=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
epAd4ZL89OR6h1xlL+a8TbQQ68rgtmW1Z52i/8Jzl0H+afm4WE2PEN+8jT+fM/SfycIT3xlmwko3
osnh0nIAAbxFQDXmZ4zJfCrvwW7D7lH2fwurtmoFv3k3hDm5zw/IRtRWkn3dxveGo9Q5cuKLksAA
OsDgJ3QvtQvchFIOFAAfGoKqI7Q5ThBdCRly9HRzLqhNxFOx0FJE3ioJtYjbAG4Ux7wUCpqOhadM
Pp81FP/o/DGPDuKxkBQPxK8DGNabiJBR1x9qV8OeN+pE35kSEJnfIJ9VNwfdZusHOpsks04qCju3
RsADFGePEuEMar9He+ikTzODjqTtNnhdCzJORQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HRTLRZhpl+JkFQwu2nYH+CC+kBCGx9OoDOCgXaAFIa5SlGzFM+jPVC5EC4Q7mT/cinD1GM29xUjs
aTiQZwazBKIMcatYAChoA4sDMwzAiEIccofCp/ZbgxXa8Hr55zzpFp9Cz1Q5aMv6qKjFPtsOYiY5
gTeDLSBIZpUVg0Rm4lU=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cJqzMM6fIBtZ5r0Geyzk5Wawcol/+tlXKLGOPGGayGKwZRqLkoWm9cv0+h6a6w34tAZnlCFosNB7
L4KDQA5XKekRJX6q4LXJlX1GEf1pmP4BeuopY28HAlwtKMjjBkoAdhTIO0vh7hLWr6euhRbVR6cz
AvhstA8JBkl1KDYg0ennxLkHyHgNMRYt/a9WA01I8gqP1YceDCOi0TKf5/JFv1D5xQMHi1vx2gsC
bkzz76oEE9y1xoh8Dx/6lvaaUmcqoEkkvyYncu0QmrBDOljYJsDIez7e4u4NYQt2+yLnz8GGboZE
x15IVyzlInzszRQpO0JSNz0AjXUDKo68YufNjg==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DvDZCz3WiJB+XAZp05gtkTmzsa5eMzZcoF2JxyvIFWaj8L+uZ5frd3azdrYzY74Gn0ypHnKrPTYh
8IKpAYYy7x9TahJc1ccWByl5bLOER35ys8DiZYa0xngQyFSsf/xUYQ/smV4xFMTEJCbfEDtzERuo
ddsf8yi2Z86hkVZbxi6vVFyczCQcOrPTqQE9Dki8zTF2esx9Fc+injScf9767LPQ7ru3lOOobSHR
PMK88nG42T2u256Q6tu+HJG+0Pa6xF3/Gt5Niyf4cFE1qV0SQdIlth0ZaWNcg3ve3w6O/+GjwLlg
Xklus+Loc0D4rzd9Qb4AUioLPMhd5EwxFWpI5A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 637968)
`protect data_block
XV2JayWTzSZBAAAAAAAAAKsXji6nTpeu5c9UFlv2DqqMOzfNY23DDX6gc75+WVtbL95xrIZUhUPL
T0TKOq7P624SdV1Bfo/CItjqrHp341XobVtCtMF8DF3GX+b0yRdpdJpZwLzhfmz7IAuVYbYRkfY6
dugo4DgADUoOTj8DwKFrjBDUM6EK/68CG6T08w+HgXPevKZJ0hKj5k8KbTOyUxvPNtyJY7orXqct
AxCkfzM0InppdJC6mg8kDt6+jje7UUwt9jt23V+YaihAzkZ+p76QJmCGsqvhiSkr5atsGE1QIwvR
FJKKZEcRSRkclLl8ae9OOdVpzyujLZb8Pf45eXQl0z80LnsDsNdrEyyPZUbhQFY9H/wy4KIua/Op
R62av0u52U1bbD/+zbCd2uIS4pYTk51/NSlUcSfnO9A2/347G8EOuEiYsGz+BSxH66xvy5zv/2d1
SAGVvfUubkrnFy2a5kA6fhEzDVK6h7xgON/+uBe9w4INtaHXcQdxYXh/T6yJ55fesirL5enkbzzj
vf9FPimRKTdG2/t3MxyWtY6XUtQ3nzZprndjryjaCTucXuBuFcD7fI6UVpE5DddnWQeWwYbz8bxG
6ZjVzYia+03lbBWdDw3gSvXTawqUqmb3C0ruWWbQDFQz6SvxTdO+f0tAhff75v6TDx1/72H5WmYV
5pTlnnPCYY7M3YPrrDXRRA33BaaOmQDXAfcTeChrUdzjL6/kExPLJfUUinbcJC2b3bJKqAhB/Qjw
dSzLnGtOxrEES1qvDAyhxX6n0qNfMZmpi8dVPgC0qTkc8ldLcxjAnR4eekTPaI2MGffgyNs6Ke7O
aYogW9s/1tBfyRSZyyXXOIq1GcOj2OuOZ21EZeyXJipp45DW2UX8V3vHsMQChyUlp2C8auu8ht7A
uuXQkdWOQXzKp4mRFHq1SizzIum2Ntjdn323pJZyYWcf5m069bSNZ29A6Vt7p6esCRspBpoG5zI2
8qndnD6WdJI+wg9Ag4ri2eDIlzhqqqJ2JvGkJ8S8NJE8dwV+fDTxm0C5VpYUKoXpUu4r+Cw7jNJ5
ufeEncwdptNKLvbI6XygUNI5a3jVm1VbGBHa0JbjXgmR1EGbP2CbiLbQbHsM8kEHjqLdOe2IqvuS
w+9mtxWdB/OUAq7d109PzTCja2XmTvwFISfZei2+6InO1+LuDvHtTxuUi+g4xHJLY/bdlXpY+Fhf
9kal7GmNSWTWpVjN+lP/mRfixLapqSD5TuPbwa3GUAJ1Wu558x1dX5HvnV771diDU6TR4SWHGB7d
CSyaN7wlVxmBONlKXHmtEaaXscOZOrIqqOQcYer1kyObn4TDpyWyxWyzlBOred+o6VS/KIFla+KL
ATKhyBHgkOUDMRG03IMdJ9qlZ2COeLRYBhQVSApYYuqekFLd/H0ul+ikhf0GDW3kfRycihAjwjBR
q/0kus/b9hy5A7phANueNsJvar2Ghd12mFYy99bES3H3idfLW6Gzg326JSJaG9biBVtDJS/HkW/3
NgYdz36KLg9+VJiWJhUho43KC8fgfQjgqG2yXC3oZqK3O/CCIcDsqSHxDIEbPtCYeWmn/U+f9zxl
Fosln18zjoctIVGD98qFSE08fwUs7/tDwQKTG3/PtAMhCF21NrP+tU3iyflbFdPvdcr0RDv9x3bq
cBBW1FazdtVpKEvJdMWhBUxZ6TxEvRxnKW7kraXeqdjpf+SYM0JDJv2a6ouSr4p94R/qYSMqlDgG
Az7XJ5DP86cV76YTe5xnTPfERUkXA41VKpVhP/vlcJch0Ujmcm+4Rcrd/Zkh+k7GNXR8Qt+0T2LR
oO/E+0dfF7fHZZBX/0u9oHr3bTy1aaOXP0OAqfH3j7GSBBYt4OgpoZWGSWsYmIgW0wSYUhm8WWag
pUJpYLFaXeZLH2tpRB909RHEjyN7UNzm0QzWSOKtIzKmNwUdkhZ3Sm4H5pZgnaI+lbowkPQx7M5h
riRJ4PxX46qERabjzWxXrgrk2a6RcfrkQhhZ32V4cxHI6+8avsCkht5hRAZ1rq/fDvG/4RLmwN5T
GGdYopEKbYhJCfBNRiQYKn4bBdaLQwSoWJ5dURJbG3E6IprCmTyAJ90KB/L93pZgTQLAguxpkym4
pJdqHR66wxKVKCcocbJpW3lDsIm7lPePoC0mCOaqMR0bw0Z7tLEbjFZ3Mu7WvIEoEv0Dq71IMHkd
xglqr3SQU+W4Uv+MqspGXhLVKH4Rh2rqULDkQYY8I0qsMwcvjQ1NqIS16FRqN3cMdPWvtcpB4S5v
7rfj3ymfc62aR5N42Iy7OLUc86QfcL7J3ljo9zALMnfSGdfBUgPHBuvVeXo8z+ER0w7mbzpqKNiV
KYS7DQWBIfIQXgETNB2Gxhq/ZXP3l2DBgmPCNwQcP4N4gPJlViO5wD0RTNVAjcfMxPEqBRio3qWy
50aPLH4uzkAQhk/g+CtKH1qBRMyA24EgGuPGEO0dAAlf+xq2hLq6/xiCdFdjKaVgacs3Y5M5Vvxn
DXFBYHab2/Mtk5EgO0/hNDnCFOiJpqQjNd+bnVLTXLW/icolo0DHNqK2X1QY73Nq+5462LAWOfec
bJ09s8wYt9lowzGGYmToeeg0jW/TdQaEj9UyTxIj8Xz8Rp0FL2CPPy/ZlFiUIpr9iU/pCqV7roaU
Sazhz6gTr9t2WJtTyEUDAAaR/ZDnfsqlGggmhsECLD795CMKG/1NIPaV2MAdjNUOLbLdmDK45vyW
6eZjnd+RcpUMkrn9aRMWQWGV14WwnNm4kmnttCOlCUpZOu4oGoWVSp5imiq2D/LxroG4m7RwpOdl
mAkqvWboiyi3PdIHG8a4I9T8xSCxzDyi419WJipAcbAbQvb4z7jebO5Tt7nIiBPIvVm0J/0R07Iq
aBOwzPoNjJ9fjuh74f5/cqOoFpXJ7+EjkSpn3afqHnU3VupmsHrHGBYpwFVyPFkgJX0GcS4jyyzU
TOnJ/XD/c+PUP8DaXSECDuqfgaTYkgtS/KNDRlCi7nsr5giDdZtS9MZVF28xnhpvGLuWcSozUzc4
2/H9bRyWIGwiIxWEUfEPLd3xtxnj4jaAQW7OEGygm8YE8jAyvAVMHuTCemoWuHCKT4Fb4aE1aNkT
NxJgxFPjMBbu0kJPgHXNj4ulE014KaXC+QLIic2jOP5WNLtQdR2/QWhmr7lhgICUabs7oCBDdA/X
1Sej9iQJG2k/cHEss5p8LnpDCQKZQ+2FbAt2V3IWPp/7X4746L/Uhdq3EY0Fk9dbXzTvVAm4Zkhd
ib9gbhlUJA5oy+erFhDMomjsN+eqCPsLDY3+MR9z78pplUO+ZrRiLvt7kl6YnZN20g0PKzL5miLp
hykCHd0G0RvHiPZY2S0RnrFTylrdKOyoBxL5qEG6dZkAPvVZ3W1gFcULYDy50Vgcqss3JJS7UKvn
TkIf/8FMBYRJ+pj9AZG2PRZVi4GIrroO6pU+vwIOLZdXgJCY6OILrZkMleh7Hbl4z3vBNHv15HJS
AocHzFVDk3lGe385lprWifeznRZunnO6XbT/kzMABVPz8BGqfs//9wbZD5zC7Dh+GhoPnY/aUsw6
+fDXKk48buhqQuwZ7nR5BcKtyU048Kixyq5Q82mN4CaOAzyD5XNrNpYYQPF9rl6r7T7sx4neGNHU
wzSjXpU7PnT1NWmJR1awjJu3PYMZGo+a3OHExzf8JvmF643aYAZeLsb6vHIJei8OjH4qOBB0Zx4x
nAzrusKErsc7anoK4p7IvR5yGd26gfeCSs7nZf/PZOv5RtGeobH10G8c3g+lLEgrIy05P1g/upUB
lYR9FArgGKVwwHgUdMyZ9GIRBnTcSw1g0kD51swTBgBDjBOf4XKjGUt0YQENTXnA2v9SMbGbqblf
DgO/TbXyQuunuXqv0bXUa7zJZi/kSZmTem2l8oE4cisAZCQsHSG+iJmJbXLIZxGzNcwnWDQnsvdJ
KBnmQptJj4Fq4GRBPGrGoiLGdul/DBcfMEY6k+yE8HSKZWxLOarqWzq9NU1vyBiHsPzLDgi1g1mc
iMXRE2pARGl7g+C0yonAOkKrXH6579QfQlLrgn08atH+SrXYU/Xx/34CjYI3tMf1wCuLKmm4ONwm
BSfTpbfnkA+Sdcn9OIReb5LvVZmFvYQtwpyr2yk94mbuJbvW4oGQSRkrzIBGnn5la0haediW3pYL
nPqRWxAMBNwbDD/DvGOp/2Aa5h9SzyPcrlgB6A6lEGjq9pQuyJ0bHTpdrSw65eMubGzNoSZL6ewt
21eOHyoMmxdFQzB4dLQYxVgPwrMkJ0JuOq3I3SWEtd9Gur7IDCfrueS9Wqjm0nOFNqoqZEZ1LN2K
eXPvQLJVJIYl86EGWjkMNtk+njziRzuKGyVCpX+ltVMjkMuaf4S90UQoUvrGZb8EGFx0/NkDBHKn
lXq1r9eTCBhSjXUDcet9SlpWMRB50C8OmTJxe3brLxm/IsWBLPSQzUne4P8nIBPfuxPbnRhapjn+
LUE3gBxKWgzK/+gTepYI5wpU/cppJS4jnSFejD+3kB646xSmuRsspFpFjPKFgNIXOb+6ZYZgSpDm
pvzHXtS22EZ3118p95Jr5Ny1Ws3Ej4/l6w5y8q9pbz3W4Sg2K+4ShdA4Bsj+gpIKW1IquX+rLStf
8jwXWfzuuqUK/Uw9s101obpLZAEnC9v19t30d2oTta2KDg7boBzJLad5YgnDczSIVJMbDxIIqWcP
tKdtFihRfN9VsL+iGcsT5sc2eAQjDyvQRY/o0rrpIkeWJAAYH1f2QQ3eCdKZ3H3rpmOVoEKXiEbS
i8OeWEBAWrjQnmFKPJrjdBLfLXwaVPtLrOpGhyheAfKQR4ZP9K/mNz1DbrZgpHeahzNPFb2ecNQL
bqlYzOHtL6q08JiVe+BCybBTwHY7yvae/4bymYEpbqG59lITtdrL2R2Vs3+qSsgszp4z/wEu+Oj7
UKxR6pLYbRfIm3vzoXe8rvJvg8raEmVQ+w6ufAwBhZNjjlW6Pgq35J31NGD17Af4+1HVnwC2MRqL
z6Rw0bK+O9nLYc4jGGXa/WBMRpDeRyo34zErKwSqvdQMJ4qpYTkHp3/k/iELf8rw8n1lGfiWbKgT
4dZfcsxKVD86/StR0LFWCT9384xI/K9azJsujNpJglRLivthF0UHVibd7g+ahGWWF5wbCwuIEoSw
KUFZeFqrK8eYlVqbTyjSuVUTDOKvaIAXBDKCBJJxU9WpgPD8F8+v2z6Q8hlnPZewkF51/g/MK7B/
KSC6hzz6OOpfPOZEEpxpxpQUrzv0TuJHwsQe/kwbnlrWeuWu9dIMxlpLQkHPMKg76ujcxIeUj3cV
EgAdFGMo+24GtzCvSA4bhEOAAfq48paJVF/CX5NiAI2K//4IbAc9kPnNX41ki/+4GD4DBikqAj76
4X9WC/Ej9vfh8oOkBEK5vi6JhYxFMyIgSkuVF/w+d8yO+jkjTdUO+FCfsNW1tysmWz1nra0o6Ehd
EpTiPtZcchrxHIEa4kZ4bYQKUGw67gsSU2nKm+kF3Q40/VqRFAd7afw4phoQfUHiqZ4QXXULNxsH
OnKHkP9jIUHCknkoiIiMF6ynrkhTPo5wqWJwtxGGqHe5jbFXPp2G0/Ts04Jb6Dgk03MRyXidF/9F
2vPeLzIH9hUJ5rHFPqBqTT+S9VZVSkIeih2RaxdQ2WqRK/eR831xiEeTmuEklfvHBQkU5TSNmN1b
e3n72AO4yA8/tEf5MtSwRYfZljUjRZqRZEFAGoxrLNMB18SeXsTFFq/bzM59EmHqx1j5//W703fI
Vqpovnj8sG8/WEebKZQbnqpU7+kyZc6sVVqzaNfkPWAhbbL956G67WR9yRzmcmQT255aXZMc8qoY
CeayZKyKysPzim8/QacpBzH2dtPhAiCXprXYaY6fBExM2VRAJzEgvYh/Xg6n/FixpauKxLww90ho
kUVUJvzUaGxzNHgqRx3mpU8xkE8BCB0w+8ldeQFwPP3lsrsGs6YeL8iJeEfGEWu+EAWA9tWie26c
CP6wtLGYVmU9BeUCs7ohfJqTm4WK56Caf3Vz3h2yZPwPecAd8Q62VpYr4CLHJxP3x4P7uzpcFVSV
1UIzIGIHkShCDwaNMcWSjBsp8OGdLlBrk2cqpkjoiKkRQpvs+pOYeNjSt3z85ja55iVYUIWn44Ul
SV8ryReS4DP/WzTkdEkUvTdg5HCQxuuM/+TTy9tPqimppMQlLMl49uZhKZi+vi3F9Cwg+IozKqaP
xClq8R5CphC/AUgNloeOna38aCWfE5b/jklo0ER8uBLTu3wM/LMvoKtQSFX3uI7nA62qAd7Uax3q
r7jiEKCnBG0bgKVhx7NrIQmtrDusZjLUItgCqDYhaa+x2nqrCylNaxNeBz/f6SBbvT03mZOVeKMS
zkbwBn6aeM4iu5UoIjEg/PJYkGrujMDW6V/cnKUrMxRXQz8X3zUd09gr1hmPrmmzWzRu67IVtTKq
3joGzPwznXytnZJXMtHtNF126yAozKXMUtQ/2BUrcEWeWkGLdxQcNm/aPI1zUipyL53qoBTikNJV
xhghnkSqE5I0lzIKMCqK7DajpPSMpL5MzgwPTefT9Pz7zd1tAqOkfOAI552AlXMEFfmvmeGfHyZ8
x20VduqLmlRoT6G/xwz+aOu5zfvLdN2/cVLqsgUKWzhU1a3ta+7pUKEujc6dz/bXHXIdciPoauOQ
/viyOl/paKhVkb8gIHofl4U278UqlLMiYMGCbA654TsOp6NYGVwCA7NfKADxIdtxxlNj6L7+ofoj
hq/R/hkhKkAaOwylGTsPoEnVoe1e6qCFcPg1TbBsT6JVwz1dXU/hMNh/CISbBtQJFNf6QLEfbLtG
JmSegfQidph7txG3gX5jVFUTU0hP5F6hqSYwA79SfpMQVjW6++l9Icr+WcEpDgQ6F7vOOf79nWwa
iWa9fSYPdm0tJ04Wb8kxsfh0rz3LWE4Tydc2/aEYYCAfIB6w6y9Fk4THHJQmMiK8SafeJCdy+ttI
1Xj7/kBalQ5qgxpTETIrc2u7DHw8/LgBq9T7f2eApiZAHAxFzo4GkVrEzCucyBqWR7hLWhbVuy4Z
Za5AluZVkhpGC3gZCtHw3H9ENQItoSBoEfmlikr2d5KtRmm1Iyhv9bk07g0ziL08dGwtvMI65cYE
fRDz3AVSJmQcPIStnIbjg5SufESptQA6kjSJqeaHCGxGXXABXMMx1M2/dS62umQQaCTUMh+msZsE
4saX2cK36PO7Wnyb5I7iS2X1nFSduXA+qFu3GOztqciz3DF7GsWvv0V7fdAha+gCKPksdsx1ClUy
qXgXRcTjC+hMJqu8j9TWmNuBfEQFHTTjStSWegn6k1zOJpE4Chafzb2l+tohcBiAh6QqJQhosVOX
F4FCAtWVK5sJLdMfCVhwtLQipUpz5R11ERsZjKThsd0dMKzpW9L23xh3gY956Cm+qdTstfK+7mDr
VME+XJQ2HuG7JvaqatTE9xAoXXIONRSZUFXR3ZrVD+pylhW74/THkyg0rCtR8ejEtJ7iWEP4AMEw
ia+9McybvLcM1A9kx28HfnkuDGafdS08BIlA9FzQlDqVwqUcSgjKZ3ljxy1dZlKVGxhp4GGxmLQQ
LwLddqB19IG+Xrf6w0NV8IlN1pNU2znllEKoeYU+4aSAghC6JexZfHjo0bJAA/vLaAIL6zs8tMZo
NIxWOpzVq/O1yBDd9uNyxtKkRQfsvSFHV8jWha9tGkWTfDSnO1fkbSQPsTeifdSkobQACHF6kxRh
p/Vc1mwuZOaPGDTNhMeqeaozMWco7eR5HsU46FciaksKdKF5KZcIumjDBOMRnIXWvDMhquN1dVFY
HHKh4YjSP3uPqEW/2NjC8guJyO79fAasrSctHvrrhMVi6zxLMiU/TxP/9/qLqyL2M0WuaztoVYMZ
uQ6q1v95XXfygHrmJVhxatK1D68S0kdEyhyoke8YAXVPfG+Xdvv3Uk0USXz4EJJZ0xVkz9rGX5IS
DDzRY580cEpMAdAyHx/XcNPwA1RApJoewfbqK4cikA07Qehl/YGX5v8J+IT1YTJV+BMhO4SLW/EH
20jbQQLP7KeUEM4p423Uzyqhq9oXYZcUnaslk5RATqSzdJyl4G+IDTv3C3cQatVYnqCRmB8t1L3D
Oqq//YYGq1zR5YeHdE26G4yS6Clj8AcGYzC6ct9rdm3GX0CRm97GBZrHPNiOOF1sXrnvG/4f13Fb
OBYFOVlZl/XQI1a4ZDPpi0I9cCDNUfyN1AgDXQTv5dtFsNENxkgo8YNvjnRF3tmfmQvCIV8YDAZN
zzOYxeaGqWt+tukTPhhiLr+mvnrvxnorLsEEhoReGjiJGcyQeTcSi0AwxE0QfoGP2BW8np13NwtC
MurDQEg6+lxxhn1dEekrq+JBSliySeJ1NdTrCyiSWS6ZOFcW19O0cRGAUMWgnbRe9CZD41Z+69gq
k21ysxG7wpvhVYFtGC2JMvt2zavxhJ5axXtySfD6JKNoGlUG/KF8PR9sCkNMIHmve3s60NE7tqap
OD1ECxXQ46N7LhnP/rnaL6gmTZvZIBFPZG3o03OkjWLtAYOOfohUs/+CmqGIuSvPdCOkQeiaNXwM
HOk/XEegwkSBcFeRNsRtz3H7IYN8vXadVNaircENF4i3keIasqSynCzSw8Mg8RDX0pb26Jvulg+r
AsJy7D4RNd3cM5iMfPLO9m4xaG3BWQpelmJ0OSGtafnTkGyORs4M5vi4oojmUcHUFvsv6+/7grcT
ayBSldX3ufXihYoySaRvdlE8TohrEavsgHvnsda9mUKI4lTQ5qQMoRLBMdFK5JKwAouXX8rBRlaQ
slX9xx1og3JR+VpTWKR5XngXDVSd6bjNFYk+M6MXEJ2lnh9JQxdKsHx/KpjNXUJrfOoO4LYwvoPg
oIf2zI8YcCFFF1LemslfDUTLJLdvCUwjxCxxUFmkBbBDHH5FmvN158Rl4ZH3hShr/L5vXCDRBljk
ONOedNFXg8hmZ/vpX9+3U4JfTvs7GNRzhGVuTPk2UZNtSSyUKmqIqmSyYJ0onw79T3VEi+et8Fpo
xfBn2hzE4H/9Gnb4yQSUCR5Bn4/6HipYyXvSZ6v7lhF1tpaJorO4cehiwgxopLL7GylmScrTNEnm
8dnAUSOSQiS72FqXNmPtCChwAKoNXeGW+Y2/lNes2P5/FoCwnuLaBtOTPrkJCwh1QGv6l5cHzmk2
Ep9BTGPKbus2kARmFZdAY8+lBJ3ETyp1WcJLFQcNMFdK+QA7dBeG3RYRYhJ/IS0mBMyeZ5Zh7uzL
74h9log94LTRO9jeMBApyTgUJ1wuDErYaEVnN5NHqiXryuI+nLGbeEVOCKigTwjR38bDYn1xdXiI
vKAvf0avnLSoV10ntQfZLL8ZMDjoVbZ5ryGjsdmAim7NoiPzVramY5ya0Fv/joXgs1pzCq+7aOZU
lwXjsFPtF0PiSC3KpM68nORlRGNKvUIx2varDYHYhgvcsXs9ksRZfhbK3I+PZqo4zOOC6HigsUWo
wnokEzxjzCL0byknbuBUJX5FE02f1JCiUFAZJiZ/cfIyULj3KlzdLnHURtPGo1pAnxeUf20qmKrY
YPZziPbLshaWTI6ZSLv4z3NVaDxma9WNdeW548NIkRvAODenK7W3q4Mgns4eMYLLmQ8LtYW8XUsc
tV+8j495wU40OFitnyuBfi+3k1I9QNNIjHH3cqs1Asws+wxjPKGZ0SROklVc9EPHNwncsJYEZEN2
w+o5EFQzsD8bwTAfkDo0KN/rBNhvQaBfBoQh9C0KyIrnSTQ9Cj6FsKPHtv8r/9dEEtHMeHVAd1qK
ZDQmG3U4j9Tqug5tcHbO/4AfN9XL4LO42iP3V2syI2/SzfQ1iZhcCP6sLjL7OyDgYdhrqIcSPiMR
iDsG4mLjWrh2ndMlr/Ovc1IiXjTOZS7hZMqL1r7jfillYn/xwIlZZ4opnb/5PUWkmO5Vaffr0Ktc
Q7xtOY+Rg9q/x03Yegi7Ae6dhh89Pzai03Ys1Sf1uTRShZ/x+0vJgIruxJNAJLfJXmsfUDUWEce3
+tF43Tg7EbtdLQbrX8UEtAe1hsDZ6J6ViqcHk2ZqkE75AdUohEnvctsSLPsUDSTmwl+nzqROXshd
GpDuKQPQAMmXTDnodIu+g+aUDIOS3Ozeq6OUhp69PtGnoEMh9avbNQDyCteJxf6TP1+LHCwLQzbE
tXjwIA0P0cIqSMPuZMN6yTryIwQ7SKYUwCIimwgl3RA9gn9MdsjZcX4mCk+ie6agQlaeBL6vi0KW
URyS+Q7e86vZLKw/bSz+NCIP6A2MDKm+/zFzRvYb1GS/EkyVWG9TND9Ngnbm1jI9QGz4eF13vntj
sKk1F7yS7wZyTDDQYlNpqhh1UWJMOT+B3YeP2iM5j9jNG3UsBycjF/UDb+/g/JsfcS2nem0+SXBX
5YGIosIelqXfb1FaMEeC7Wo1SeEeP7P1/5xp0Ok72UfxWLKWxXTHIWDaYfgfN68DPj2gMFxlDn1l
Qn9phCtrsdh8V87U+0S4YXbser6CBqSSXDVZ9wFZxgG9bFYwzkAfKFQZNijj+D+oDP/dhb8AwgmQ
WXA+Dpw+9iATLdw/AGFVY12mYJ1ZQK0pneSE/52M9lUJw7PzILVT63a2hKkV1JVxLd9kQ5t/00UA
/7x0ck7l9jc7NCtg3Xo5gqYbxujEsTrNrDOOaW8J7VQzY28GjgXIfdT9vq4ISxX6fxlUGBlzXCz7
1O466AfYElHKnMNGjgGubiLUJGZwXMYL05azEWRfWEXMhvQqvXW2xvQn3zl5gcbvoZ4BLx2IE4Gt
Y0ehnId4bnyRDrqMoV7gr7HXm43A3RiPWr6pzcT9LFRiP2xJvC3TDFIHl4z05mgYAAF007ptDjL+
drigykuD6//Dn1L1s738xChm3Q5aHGv0RdSGJ85AhAckdn8pJnDdx/3sDGdZ0zSDyaIT463ME9ew
cpAexHibt7Z5JztcDNWAML7i2Bia+gitYhvU4yKIQya9idv/+EYHSnApK1cUk0BVwHB7ht3FstsN
vZvubR9I6/ZF3nsPCaQojgnfvLJ2yju99+IuQhFH7vj4a7DAzyYOVJFT3QwFDukua/zI1Ert6pyy
q71Fp3J7AYl4bI7GOrEqpmgdjO6LOJ0v8SrY+yUtAW6+3dLcMeB6soys1NC8FlWgv2CVkBWz3SfE
4J3zStgg14L+dYA+WnOpU530BQkitd1AGrRR3zlyK3YOTA7xQ25DmaP2bAoUzy9A+hc6wwYuESgr
F6c5sFa+jhpgqpgfg+7qrhc9Kno8vPhNg6UaQ9d1E3M+o11wZM7QUqEAmeMNQY/83MMRBnvVHYES
3NDvKx7H3CJNExStd12+IPH2RhNYhBe79MLHgftA3ZK2fymjQVHg3xcjXB/KKWGGnxAjvIPsnX6o
CxJ/U5Flaf/+mCRwrJqkHytl3mSTBs48pvpWHyVeOae1tjXrEZ7EVPPe8VBI0IuDnxysGECp3mUw
wDf83KvJbjJuI91zy4xOuFk5Fgygdzj2jgBDEnN8sqQce0gLsKU0iqwLpU6AXulNqiC9GzaeLWtg
x9SHp27Ze0NsIFPRTP3E+qVcOhXvq0MagiEGiPtNTiWv5EtsNgYZCX1GXVfzc004kD0NtmYXzsED
DyuTbKHNovrz0uypb3ToLOuaZZxKMCMlP/EfgngNAme0XmjO49Cxbzn0RPDD3tqYw1Nf2Gn/jLxk
YuiRQX1S0cFc3mmAk6Fma5OPuc93mkXqPfvxVPoKcqxKb1xLBqJtm0lrJqHAYfH9hOWj6Lk52t6p
WEDehV9Vrl7Fz20NvYboeii8BwaizmepRYhe6YTYg6vMY0KUlLzsklEDi6ZkYBWFTellWXzmwJUH
ZCh4KEifmLFvwLqBVKtKbU1kXwtYdGFpwbNGHgK3jbdMglAkL3wV96Fa5cttaulgOk86PsvKWjlW
ALbO4cwncIKDT+Y7HefM65B82op1afjC7kwhD0IJzwtLdliuSfDkrGkt18unTtNZzYHR4Y6MR/gh
YzKrXC6/VDrJm/mSC44IMyqTWy0LAV3STOuwDleXv/sI0Zzrt2BjCtfUFNinecFEIs0vCV8+4suY
WNjoF+5lbKR0J5udJYtsDc4i3aFzQzCJ5o9C18b6R82FKJGQEfRuHbG0T7PRn25/dT6qeTHEiUPC
bIctRCut5P7Nm/dtWJ6iH9bcOOd60Nt79Qh7K3n8/WoY4VOY7SNSyr2SJMtpBBZa5mp7nLHjJWxj
ONGfvqypgq7U4xWjkAbV83kTjI6KqSuXPRsi93ynAjZYWUMqxmw5bCRMNtJnnW/vgFDYVre4iGlj
sHdWuOaBDntSkHUO5TYxzLb0dtJwED+lwDNisxYhmcvClylG/s5JMZ0nd7v9ggR2BnRpzBnlL+Mh
05QVwnh6OkJ5iRqYyQAUAlpmfBTdUPyjg+OuhhqcvzcDQp+qVsbsrmNkbB+4HEzCUkbhoSTUvZGU
35lM/hSmmzGzlqP8+UBXjcP5P7oZP9i9UK2UTih1Hdfbbz6BTyN2c9lGyAJuKWceqq2z4eqgRZlc
o6/8OiO5+xChO+GAv6ktbHfRHZulAJUMtTx/vtUlIgfEbCizB8HUsH5tO2L2P05HiZ+5GiDZHXKq
RRizUctmRfSOGbXDpkXG/2KQivDV0IaUZ2d3pyfT46lm6FZMKVufTcldKRHEPbOlPb6exYtbZTm4
L6vzx0UvgNaRrU5Dfcwt2gchXikL4uZAStd8VNG4sBPwlA8mJEHHlTuWKnX+nm6Sv5vZPkblWrDL
TZHxJSHxn1YD7p6lOOyIoRBykQ+r4ChZvDUrjqDrpjWFasHqMywDpZt210umaBalkx/CmFa3/QJg
Hk1O/CeukX/iISXtIQfXzhAVdHQdRj/KBBLa91pwG1dCFyw49edAtBJHP+4iOORPnnTvRMhRhNSk
zSWLKCzHypKtrq8ZQ+s/xSWY6NUg43NmyKps/59I67OHEp9p70vsr1lO/w14j8Hg/yettcjfk2yG
pPBKset6rAKQhabulur1jNe+qATZ8e9VrR1w/zlfllQV7LC/lDs1Ci7RZGQXiKliA3oxjPbWC6K+
g1Xb/Gz6MGcKFKOhcGmxznowh58BwPt0AD6p2Aoyqo4TQlQ5agPk2/7uJfSAXdpao05j7xy7BVJn
QVts3pVXaPH4kDVmV2TJYcTsVNK+A8m2+toPy6n05BLH2hBoM0f6JBS4aeQ8ClGg3S3MTbw2+/+w
i5GAaeFcy6AL0I8lfHLG9TtUMWQ+hCAuLFnWY3iYnEcYQ3T9npHbWRVf76iikGH80muaC/TWrqO+
4R1qJSEws/xashpHxC05zXmpsCblmShlwe7Gu4pSZtzwZDVkh8lQbKQOP0d6Py2rUsqT6RmbII7l
payCkVSOuKrqQMJJ00xA4KlqQux/tOEshsYQmQDQ1zn6+CHIi4SuSyoG+ai6W/boH1F47y6PbJD0
7cfPD1+ihNsE9C6ZXe4yBltQCQbQC6emMjNqlJ6iSmfORf6CYAwjXbBLTcpn+RhwlbSqhOHXt3sF
klAGbN9GLAmcYgFfG+CgiI6aDdlh9AI+vwFdaSvP6uLj7Yy7sXtvumwEqSPuis7IQaOcBSW+/j9x
M1UXx+vtszs4SQBverO0unavnIdKq1LNxfKJ3ivk6VwtnRNSHLk3h0+5iDlSikEbNgu43H/mE+mu
sYGvDIuRiIJvWkRXbqgGesOzp2qcrFol9JyeM1hkjDwDFSz8zr6y/4/npaBKw/7QZpx4PwVf/TxN
B142SDAIcjDYFfP09HKNEgcScXp99Yu+Ft+2kSxjPi/jYeX5Ubbl2B7aV3GljZiCNcKf8gRjnDtf
oYmiOqKiu5s8LG/6VrxO17V5qggaBer4NPQxskaH64/XJ6jk6DvVC/04PEEMXB5redxuRmpt6jl5
cpN5eqmXlNoNurtXbKa4T8aVw8pSXrSIoif+syfB5D13yq4o1tBiP1MlWq5xu84571qJL28oo+Lp
dugR67UIKch4+xbHIxC9Dg0tUdNb/h4kAA6aY5X9bo/gxiB/kJ6jgDskIVK3LtXZbuCKHtMN3UAo
83W8IOkjJWIBMnvduPMDJ7TYZh9UBy4qayFbEKbfcGUW856MX/nmk+8Slu7fA1O/iNfpZST1wO9J
EgwCojD7Zr3z7ZPBF9/h6LDwiNn9y+7PpFlSuiomO2NrCAyax81FVg064NE7b2hDHXSB4fZI+4eW
7MGNrkoKeEkuUDeb7nct5vmB5jUgLUN4TT+8OAEnCsXBdm6pY+mRZVZVsbFtsR5WASa01+uqKzTl
p/68B4V6g3VQAGN4QRx3Hmy+af2Vv14bwcc6KmIFgPNC6vJMAumgs6Mtg3w+k90YSb4AiB4tktvR
cIbIMBTYb/KLOnhGbERGXZiNvkp53bb/B0Kl4+voUcPQk+LDwtqmh1+GV3JaYLWkTlINHnrmE6Eb
6cp46wZgT6YZaxbS5pMdBfSjmHTagQib7LTTlm/zHN7gJtTfSbFtThqKGNBvomet0vy5KrRYq5bR
sSbG8bhKVuLI2KoMAjqn+e46i7H6sAFO7OIs7z0ITQtwujUi4Qpf0iw2lzrIomQFuh9rm0EAgsIW
0GUSpWiR5c/G3azq0qhxnlV79oC2pDXpWrysUcpwDBWAXV1FtwOv+rGIa1JIbS93tLdhsLHbb4ls
jfg2Y8y6fj5Xx5/Q0/uvA4ndnXil3H9+QMlMMtNNdzqkaX1pVH3qhhtoLB14e1lgG0peZLiLh1K3
cIY/jPhjIsp+KWNavhuzdT1sQSv8ntvu55cfw/Utcoa8IROBezh9veauHR8zQbqUw/7xafZaNvQB
JUJtgAy2E2Pa5yjRM+r2wh22zbgRAP+iPIHIN4xlb+ncmYp9/QoOf5bjWj1ViK9ZMOmDPUn7T0gb
2L1Pc1gvYTCya4l7grnsXBjzkhCvafVJuODoW764O48kjCf835wzwNgobIiLJHkr3bImqW1LOFCN
CnllcW72e9qoIbJvnMuHCSHGubZwRll79L6eHgHpaH01TVRxKFkse5eiXe5megENQAacynxIN5eS
v4UnoxHD0BbG+tSfx3P45AlwDa3R2PHizky0UCm5ZJyXgx9NeQNaLRzrjtLvXeF8FRGCLfoK/67T
wQw79faON+v0Y3SX7AFLZMgtdJMpwFoKGb+/WN1hDXt0EUR+33rVeuOx+ic5g12nwmdCy8lsIfTo
iIl2y+/7/wuwWIptGrmqPx084XPuW3RZ7SBQiWiN+QxUZiK8eJLnHnyyYzMLt4Dls7wFH5F2PWJk
cr/jHmaXmjr/Avb2Po64TYuQg6dnOWNHdPUFeVJBNeS7JrIqVmDqa8+8m6ZOdXx4VEhg1uoIOgEq
liqxnPFgt+nZA9zLXYuRN2HC+AXiTs24xKgfbqoGS419jVVCMLxSeRj1zyQ2jVu4YX+51K77kd76
xn3i655xL/E+E+1pMwz4hSQJhpcMeQXjHj2BDc/zx269aasTz/FTk5o0pdgT6gnS3jkXtltmMgdw
hkQuvTDMuqIj0oRcAc+qOWXPWLiq1JbrqZaNT7zY/cWHwo54kqj2boHytPp2gf6ka6twoBveoqRX
wkE09cckyBjU5cuIJA/S8iAPaYahdy4dqaDihUHWZyJwzkNK8jQ7ctLv1nG8HRMlUHbAqZola8rv
xgXx5MAXMYDYmzRbCm7lDcAhj1rZpZhBeJKmraZ0yy8MfkeSZoGeZlMEciMKNfFB5E1OBNyW4yXH
gNTL5FqyWl/YVQ3hFIE3UNBIS4lDbIna30Gn0qnDE8eDAVONhLT2x5RjIM0DpgiTG1YBsgFs+1lQ
ivYVD4He37Si4sWFtpfO5B4Bdpf17TNyt5e9YcyNhpJyv6y6ejfeXcBB+0dKFmeAhRvpyMDnV3DQ
0rHawbz6ZnW1eC+yyUS1mYRxx0+cMVm6Tkbmc1GIjhz8BfoEB7USpqJkSCBQ9l/gaaPYBojnIP9l
6gg+Ew3B7dP99WIx/58Mt5pBB4DyRPNBEMFVgqOVV4VxdkPFyn0hoS5gGwjuC7HcNx6JOj9YgQLc
/7RNTd1UCXttw6V42wRh/gwHFOm1k6ri6FXV27MkFBJDn9SI7DGkYCsxq1IDeAvOSOO5OejReh+5
LB3CMywbZM/7VVmyGvzaKYt8L2MKDF6QOKiuuMvGildlUGq1nz3qxuygdz5iyQY09fdSMuKsMi7R
r/xMNuEHjizMvCoUr/jTFXcx9qyM5Ey7fzLcdok4LLmPNhWEx9qNRZhO+4Pmfkqi9Plu7JfFM93t
A29KVBRR4L1hQ7IXoQC5DSwNM3uyEB+lGIVwlzauxNmPdBLeiCbBmzCSUQjGQ352lU3uAPJtSUHc
7gUjhpP5EMRfIgCOX1qHiSXPJQTr3R8mFZ39GJfvpvgr8zR7BHLiI5/xRDhDPUuPyCswwXHReDST
3hM8tICEdrox8YEdeZWiCVF2tQZ3JqDbtlO1ZDZElQp3hWiM0XzzAjbg7yB0a/yx4qBd8hRyG7uA
tj5KbwBdJrqhfQTvF+hAigJvwilDkP38xNzq24ccaM9f5VA4JEwe4eynwFIaouG30ks/q9vnlUqR
9pcfPcJojasN1Vlwl1hg8VvoN2T7NtUnc1upMUDMpHDc2SX1JOWJCfWezNifZjsO56hiB0hFNwcw
kFy71yI3AaYvE8hekRc9BPg885rAk9AmiVqD5ZG6mWyRC8YCWhUIVIVcyW9PGkAeOHDyzPgnGBpo
EGcbNxC4m2gsM5cOr6e+fZbhOXoouyZD5gKUnbITfo4HtXoyMKJ1Nhd5ANLvnJtd0z/8+qF/8cdX
3JxxjdZLTPf8psLX0hlNLXXCEtILMuX2hlvDb6Exp60u/yA1ndifnJFdfanvFGX++pE1SQ0hSds4
WKZjNmUVe91Ns31a/1Ugw84aEZZt1ZuVMbmA/qBjLhoLPrgfmeOjfsqDmWtrJAVBhm0fg9UQxisq
mAFDIanKPlPfCn1IV9AzcS10MPfJ2Ura8fiUq86UBeXQ3x/ZgJ4lPY7F8Os6Qhp6pP+/SWbyuWFj
fFdGyEcud+rZku4kwpjgQHFmSC5px/Gx0PE6MuHnRZ9vyyMWVySiKW8UXR0s4nvYjUQQjivCRXZq
LFovPueqE9480VqeBBjbk8fXKiw1W1iSTn/jKckDelf43ymKHtVGF/VKf3h1KnQdxh7yQAB3MTiG
I2YsTQFyEOeMNPGwczsdqPAa5nhGZvOLBWget2ys8/wj+ASByQnsn6ayhoAS2em0jH7GHonSOomL
bPX5XCm+v+7dfHL1zG6Oy62kOil82Ao3xv5K0UvbhwWEqwWQhFAp3SXvlZ6pmJPe2jM7Nsak7yRn
x2pDvMSGL8agUntJMkf7JgLnBMWA7F3cwfGL3rGJL54QnKLrkpE0L/G8FyFIjQF9/NYm3RtlQqHS
gWnTzmXThCJBAPgax0LoiX4YclhWkz8fqQRQ1ly/JnY63spHTcNs5vUW9fIzmigTNPpTuIxrezcl
KJOqLQWx0fymMBcwxfZ3a0aw/XB9aHmXzuoUbtqQqhQcpBtNoy0jvnQPGQoFs+uPGLWdvmjib+EA
pytQvt2oNAPDkKkGZEhpmhy9g364PBbDg2sswgh+mj6i37jJfx5sZXpqxywUEDzIIPN/DPNcw1SV
2Gfe7BMJiM4XwaGZ1dXVrIP5PtYPcQBNruvoRKEmJrHyt8oOBEqoT6+aXIvCEb3+tjZEjkjQEX8A
9pnTYDxX231g8SSN+GoaYRJAKo8yCdJcRdHScdh8lzcezFbuRf3gxlcz0OOUfKhOu5GWs4pzto/s
4bMsGDfSn1o2XHimEC2geoQq79GZLV8PwmcA7uGZOqdw8LM189VaS5JwAoP+6Z8RTePhmob+lgNe
vfFmKiCrTnRvXZzka7g/EVPXoaRtpH/U5/2bH5A+l+4e5lS3xA2P6rK3OxpBgF39tCqHNYMs3bqb
msinGSV8cRL1EsLkerqpuVkMIti0GDmtnaY5fvWYR+biDqXeD3b+5QzfVHdqPObE4LPmYI3VBRTq
LVkTgOgcIOOW/Wliyvsz+ZPCkHnBI9wKoH9pOB2Wy1Lp/a5J12QawwMTIpPcaX2WGKPFHPB+U6QP
ignKlJHdfhVf50MWBHx+mXDhgN75CpBXRbqU53PBWlQCGXboouGwVXoUBnBY9EdlrF/6x/+EymKs
cJJBP5JttqmsdDNHzmT6sPMAEds1YPN88zczS6CK35VrjxxYVmlwWp5qdRVLHadsFqJsr5Vhh6xz
FJJ/dAEFcCRunXmnm3YAfUZ3gVqBsQI4IBZj6mbuqMA3RyawwR2nrxvMZIFIV4RrQY9aEyPVJLu/
39ao3KPUQZRl0IgCTlVKly3oaNeN+ckC34WqbDLdtHEYZawNDtecQS3X5fSeLCGmrjBBLCoHzGyZ
h5/hIJg2AQfDJNgOk43G8Isulh20N1a0cNg9I5KDmx8sK0RuBJlX7PWso86wO/RnuAp/s0L6+WEn
D9cFsn2XO0GG6GnvInSUq0eDzekueYMyI1a6y5gZ/bAg5eQhi7wmCV1ydW6EO1en+rtDvoaisWOo
cLukVC+Tewc49j8tbGD/P/4n55AWN6BNb3hM6EVwwChKdkyDGyWIZfvYi6aWtlc0ZjjWkI/NEyk9
s0KML8Z8DlVPGMaAGG7gMOXutKRYt7b5VyDvZXrLzeZXCb7orZa9WmrfU+Lf2p/Njdnqzdm0LChw
+jXoSe6J1yoqj6Q8I2jXeqPldRcMsMp00wxzA9xdeO1lJiTJf9WoBTBQ3KDq4VrkhBLnZMh8LzNo
mk6bLEsHXVPiTsoEcNDC1U5QtPkImITCFhewhf8xn9jpTT1hvPTsqlScyyYD50n0LsdJzDiFbF5r
nBfoC8O5yVIbeBPq6Ojk9KPykfXw9FO2KYZ3+Fi2ZnkCx402sf+YlAJ6PC/3FJyFlAMpQPQO2wFP
Yl+nYm/6k/9Cs5q9w4hRCCPgnnwu9XJVYM2a85WbF4GTa4+WZuzvNIHYY24hjkvLleKuqhdNAPPo
nEpC/bj22uhnYAbCtuh+0NKHc/Aahtthm18gOA/ZGCjIVCysIMmmtcrDo6mzcjiZoIALtKxySPwu
XDLV1wbwH/qYFCJnNai9FjTYAGcnskNGzbheCYdEVx5IXfFMuNS4Gpb8bkOeoh5nqCMepEYOZJLz
9AwQAIzXaym3g2wElOVeDfRybm5tfHd2NRqL7+owUKOJoIpGp20tysb0pnPhdSz7hgWhT2yJqk/c
hF5hqRfi0cVMztejeKZJ4JPiifxfUJfYLB5wMw9DsWPZ5LJpBNTSVUnElmMZCJPjQ+11XfNBu5ms
fwqYtq+OwhaMDCQcPdAaEL6D9QAZEiD9+GiZs3eRfMxWNNb0Azn3esNEnEL8B63ndJU7Spg/95CS
vv0UNL+spvPvMqyKoICcLBrK6Sjov1kNSv8VwGTKDaDb4nRwRufz9mru06My5XDwoXSex0u59kfE
qt0FHSkqcsDTYCEeusJIuNqduccnTDif30tfBzcXJmGzDWvI8TlAHja3Q+FnOmXZXPpmBBPzWfrT
a2CoJBAluCNinrfk6LRXJLIk+FYKzjZ2xF69W1F2JenljuVuRrmuIgzOIQVGiGo1L7turbFTAlqK
Aw3HJyYnNoWkdaa4dUrdaBknzlZXzFQ7RFruAbiXZz7IjiBrS+AtF6q0TLMVEY+G6mfO6B1awSI3
jniHTjVW3EzBOoysDZWwlsGhRcNoPG7dUwglEY/ovg1qcAnXxcBajZ7lQpqskONrUtO+7M1dG2CB
dDnstlk1fNQ/wxZsDCgOLrUiJpPJ+MwmnEgjgBttvghhIurC76RJ1mfepV+lV/z2yNF3ESYiGJhP
uAVXTCCmwhbo23VmbCHjIIY5pJLOmGVwZOuhjU2DIKz/7u6222MOVlkGAcjw/G7t3zAIN2/N8/fZ
2VEB58YB/VwQJan8VDd6xAfiX4ptBrXo+XTSw6j95ApkCeLdlPEq4pfFkFApUjEN6s/crJobODWR
6LfPP9iR/CttijJ31ECC+If0NB3xECMaS16R3d5mbfD9vkSQuHVPada7sXaTSdecWqQmk4psgV/g
aHh7YdL7wSsnAWDBd1Cy2oZPrrSFoDf9J0QS4sg7zq0S71qKAMpGtqckpBA3LgdEG8h7odUWedwR
hXBfwgSjmUmxfxklPTBEUYltaz+6PS3bRjmXw4ICeTUr4V/QNiLkEkNdgrxhR9BetZfX3RLcK4bv
+4d0wnrQE9B5i/4VQcO5M5VAzbKl8nDmZKVt7oec9AFXWEXm2TK/KM6sIEFS6xm0uYkmTCNEPgYs
ALLoVpj/L9pXyA5b38gMdzrUMolA7bFrNQcdOYKrbRfuK3zBlF4rF28QlzJj24gq8Z4inH2mi4rk
VaHcz6HqIGJijAuihtKmhAFUCN5G1BJk0e+Q0t0oLkaQGum7OTYr1rzaW7oFTTU2MWqxIarCllSP
Ud+oLxdtF2eIkuDy7liupOGM/DceXwtLeqIVNCO0Us6Kt02fFjCYXsifcbgfv76/fssAKUYfXwA2
7mdbCqWcEkc63v0tJM1Zzi7Swp8LY5ghNeKGUz/F6mR6g2c07lCx8NzJdwJ78diFoQOJ9dtw9Ml2
CsBMpiJ7jfAGeyBON5th4ZaPbB/8qNu/yvtNQauj5RgR5FwNUEaiR14y/HJjCe29LcGLTe1G4LZH
fWeb8S+NJHsKDR6oBxCb8J0ZV8PZDi5o3QLTGoXzN9G77kkbPcJUR3kOkQAPFXBSw+v/XK3w236W
Pr1MIHJtRow6Uqi7sxjIp15Wjhql8oq68ErZxHj9MndtF2SBHjOJ7b4Ob0KJlRq76qwQk1l6o8Sq
Qhp/VLaBxYAJ2YR3P9BVTaqv3mZGTelKNiMkk2KyHKBEI3UqrLyj1NIfaiR/HKF7disUpvkfW5lO
P1coG3wKfeQhrwE60a1+9HckxjKrMXRCRPSiJoPSG4qE4mCWvrKTF5ApFjI53UFwL/QOIA7O8rjg
Lf2SGtXSftdQuQI4fO6sKjNZ05FgCFLBgG/5latUPOIrVV4mE2MitklWmJk+YmCD5jpThiJ3gzkJ
PTUGoLxMCJTcwFJrheoftD1oUypteXXaXcqn2M2DlkVO03rNoyEKn5ABGvoEP46T7P0V8WjN49QZ
/kP4GdYt1TM2eCyd4ZnKKV1qpOJyXhVMEVHPAFwq4JeF8f2ZU3z5DM5nvYQTfsKJSJinzRT4XQhk
ocv2n8Mqp7KDzHCjSH/eUk4Bfov/s4qJlxUSW7yJpru0lvS5nwPHwJPLdIIzIPVCCSbVkBkunyNR
wMjoUFxp+WPQ7FCLlPrLt5xMqhi8aBGx1vx9gINYPeHjfp7tom4/zNH1kkQdlOn7IUV9yw8s2eU1
NaH70Ux3pFUB19dhZWijboW1AAem+Zs7z2HulBtjbyuZRE3MIy+13qvQa3+Kc2AQEPNEazQcLagE
c6DJAzIK3IRZr/9py+fwLqQB7hkDbkll9kh8e+gjYb1veDdaEZZjBXIEvR7Cu6qOzCe30dwtEN4o
fRmO8Dg/0qL57i9HlaDdIduLp34Dp9yQdffDLUkcNli2hkZImw4U7lGl+vloDVZDcZtSyveH8cUD
yzXT62pw3p9NWaCJ2Fat4pX+xM3IcXuEM9tvGOXoWEC5FpfgEyLwdcKE4XS/zqpyJmwci5Op0klQ
kILokX0xM637C79F4NfH3PmsuBjlD8FzrhtCBmL6w5J8GIseBBqoZNoBbnFSSiBffluRyS5/LgdT
AiL3/LFLN+Qn9xxYBEjdoqJ/mkW0hvMN5tCnUS2Tm2cLdSWmbHqtQbTdzWyNFdCf+C+qnCdhK2lx
JuQ6TgbHpKMtCxGjlhZbzeWxyGlY4UkF+6q0Vue5g1ZYg0uXh7teNG5waXKZLkqikxShmtC5gG30
MHcwJE9xuH2k1d+yPW3ASsdNtF1MTEnP2K5wdzzeP9DT4yKLAUDxXW7W9Rvh1clU0OdcPW9PAYyU
zvfjPnygdcBlDMa0jGKrc3UgWE8rGXJOsUvL699KWXWt3szIvcwNpZDVHttqCMrjTE8p8tA1bpyU
9a1NctD1KhAL3pZc8NWZ0Cz4AXGhdz2QfVrsuN/3X0XAoY7TlN8PiWyhn0A84O8q1jie9Fe7/k60
7eA8oUR4Gd9uMuj2AQNAi9UykG1SWk9wWKsoOW36yzpfRA2h6LJj8aOZHkwqcuXGuPWLtGNhKtSZ
UpbD5GLZOEw05hKwWJlfrBvsxJCs/F9jg7nFppEiQxm/OaW3fN+OQMNLeX5cY6sJiCJwjODPI/1x
Lbtb+4/U6PUF0B/1h9DwEFSC870geq592q5Jr3TRF0aiHHUW3DB2v0OJrAHYGx8UmuShYwJfbjKM
gupw5hldy1ovHIr5PlCsGpVq74ZTzlSfaTZFVJM2t0li+YOGaZqQgZP6gg23rIykLpienLET5XGs
Zvlui5R7lD+F0DruyMu2H1pNm2JLHxhl67q/yMl1cwD1FueZcl2Ldm48cS1oaxe2KueoAMBDQ5lz
RQuY9zlrunVEt/xYELmLbweT0wcwKLjrWczKNo0UtWWAt3NVQjDELURlgxP7dikCTmZuEcl+qHHm
Q5uZo2QZSEUptUszf9VntIHXswp0fivCDWdmE5cODE/+N3dR7liso+OUObwZvobQfUUOCpyw2kqC
WE3/yRQ7bCzdn8bsQFLlj9VyNQtA7sQaEDJHrSz4NmaEmpaR5S+A9yCvPggD9ZEyZPEHI//cHifd
It7bh/xpvYLreaca/oKVrNk+AYKbUZUETaRNInnHesdAunT/Cj3uO/a3De6zxGjOypx1u2YLIjv6
H20Z3eeIt2a7dnc8A9e9D5FGtntUpT9AdCQSmdasSzxoRB+nge8NKqvm+f087CgyeAsLWfgv+UWW
k7x+uFtUt2J27EjQEOkjEdxjDKUfRUPAkP18kM+MdpiWkRL7dv2qaoD2YDcs0LqYMhJC7BFE4UxM
9k4TXv4clBSXTctnNlz2QnYSBR0ZQgSxaNIlM+rQKTEDipKXNgR+nrWxc9SMuxxp8R0aRNw1BAt6
3nNqGXNKqJ6wVe6gI4lvAHw3r7ENCs6CmpGs35RAN/DhoWjjIuhZ1WHBJS95iyiugM+ju0CLV1PD
Q7xvzJPOvFby+RyxJ9pAszyd91y7cZrTZoSbPQnhtFh0kdTdj+gRBXTFybZDpVuOHrW4TwHkYIwe
YS931dRfBoiYyBfWxVjnmuCY3ngK75CC+2FPOk/DdisnwfaeBJZpF07RVE6QRCmgBQAJvFdvtM85
1Wqxh0bbitVbIsExZgGu/E6LeGBToYU6ciyjvmS7PSKw2Ca+JubZYMkn4Ru5bebTBLTB50ORWjQh
ldUIMK8Y0hdBDwFbUzPUuJab/zwOQQwkDapq9gyOAdWHxNNGC60uXmhUhQQW03+wCPW+inqBGdZB
B7yk5vkWf8ddsPWc9A5Z/dVEaRGgmwjwduFGSVySE174b6mjPRbd5jDZQ0k5DqbtoF9fazVyUiZz
e9dk3smoxdK50xCY+Dm5Igper6Eqa2HbjAP2z/RFwOXredfhT/jlP3ca+w2ahYfcydSZtcpn6r5U
Cbm4Xfm0uJZ55fdSWo9kYg8fgK7IL5JC8L9vrF9qyQYlHLLxWEl0T4h9w7zQx73dHampfnyPOLRA
5KpSWZVtiJC6A8mTDyjn/XxnxoVXU+381autbYmA0A/KNHmXxH0PwXRG7mue44D4W5TWI9JyTLTN
H/FbV+5Nvqg5A86nsVDltpt8P+0MCFbqRIiqGjYz8wnj8hErjFua5Eo4xUY9OKnw506+Oz/ZafLo
s6VSTpabSiYAK4XnzkfLt0AeVCv8KLLbz/+b8GDr4UY0fWEkjj4bfj4E7KKWQd50DjD9wd/WwfBb
Vq9f6ROQxzKRp7ZMOgfp1AL05h7pHCmEkk0JbN84O0HePSsMLrug+lE4FrRxX8L4K3NUW8Lk5Ruj
kN41h1eNbyTePUeBTz/NxsfORoMClcFyeCj8BjxGmbO7w2UtafzkUwWjhCqeihM00TNFZHh4PWeP
cYq8FVU/legFIWamoS7MG84aNOliJtrzJ/adDJZn2Fzi6wPjRqb3RrbzNkFsMSBtbRgALM94vd+n
3mtXoMCsS9T2e5JPmoza65AvGHS9pbX9esPRTn0C5PfW6R/Ge7+mRSQgm2YKQ5scdkr7yAJkyUpD
T80ezPmUO/+oqIAX2zv4laSkgze1tTwHlnsb6VWEVLg0gb3EkZZdUdX4OAXmyTYuynzamokD4hdB
UxXZKR5hvtOycYUTmNqoEPTPUNXEHefF8lh63hkv/iCF1+LBsqHPsn4P5uQJUu7V/9kYbnJ9Mdmx
clbFbKz2mmBemjAyip2xLSVjKIDSZOp3oOKyBH/gTn/j4A9xmGWeq+mSxNw4HvTrXHtfqb4gpTfb
78iN/lGiKROtPjZWi/5sHpFBFjlHOlsLsw5P+NtGX3Vao1+UALjK/sU95sG8IXYNuQz3SgLXwP1N
raiCD1sLPCH9QRYtu13Eq9AbOGPZel2doqJ9cs4UPCgCBWZsWS9DDhz0cakVyO5bz4ea0CmjYUcV
VsLlRNJN8wcw77kbw2cKCKp9Roi9sxzx4N0raJNzS3dUT2XW4N+hw5YsEcqq1i6QeUOlbNHSTSru
PH8hIyACoK5Zji7OhU9RAuHsN+h3b0jG/KB6NjxpLsFM+XFD9mwq3ELKSoXzm9zMQC7+QrzObNtZ
k4r8sXJfL/KKX/gLyt2ykh8yYtDEpdn+tFQ28Q8ohyI3KwnQfWpGTgMI5J0QmGh2NpPb3GnalTW3
czj2ZVw6Bcl5dcobpZzHlz5gwsYro5DpetOaP0LLZSZeMHsFcmzSpwRozoEzjjWvGqkjHicTXMAU
LRfL9aDWQU9eTSMARQAi6lyOh5532fblnvLUKs372ZU1nHA3ZboRoXkHEE1adI6APSTJBkNwRWdO
xZV9BlIjqqOsYCz4vrrt9akPDdMJwtR7XXEJHbPuBL/puSYytC6e1F47OQzs0PwHRHnU+6XCzAaJ
he796WxE+GWWHEGi1j9q5LbzA6jszEGP7m2nmYiTAS8mgHMK9nOTSFfhTEGU27Ci942WcHZ2Raih
VeruPFILmfksjSRgj/PldrCW3xWF52xxMXl0PXg53tRsEXOHM3CKCGWKN37TCoYp+jUVXBU9f4VN
zkdvOwlIRqio0dxK7qLPODMLBRw3ryd33PEiu62Ws83ZJcqJKomm+AM6c/I1hFdHI6sb83ekmgAJ
jNwi+ApU3RWra28SNjn5tP2gX1SpNlyjlrUPxQAucQFzoMlKsygYxjmXiup5Mq976+GIzC1rjrS8
Z8phJ+mjzfCd07bQmA+4F+C1pc5V2ZuAWQkHeFb16lx/VHAzQYgtsXk+/rBddNqfKJ/leLK2ySEE
Bvy/6lgGko8+TF9roS2/THN92J3WfqFrR4AVtVX3dklxW66QANnVVl0lJtL5g5yOBH+SWqnMXL6W
LJE4DtcHmTl/wia3zmyQkHQZnWERE0Jgyguaxjib9305865t57qoeXTFyMnsIrrYFEws6sxeO2hF
tr+qdhsuu9VFLeSuTeQpU2PWFkfkYjTOc1Ri3TG6OlYAsHgTolgYlvG5/6PTN7861kIuEG216uj8
SD6zNah/glcncnBYMPZ0D40EtY7YDtUI+vNKGjhauS7DjvlwvKFdeo3mB9hM4uRvYLNKQ3jiXGpy
LrIxTGkShdgZQ/okm2gVY2BGA+gGsETN/CRVT2ycQTXWNfwyIFjKolRHTG3kmfICKSlGIn4Vmjii
ADpfF76cJHiWUcttp2xtFztlGoG09tnF4fhEFVUaW77Z4jiEhU8Rf1WGD8QYLq5AGS2ZRK0jsA8/
TF40UE2b52d/qPactk/DXDqHkgkVzYul4iV+Qnf8cCmwo4NjlcZeDm+2tKE+lWPyu/qTMnlPtfdu
F36UOyVvAkkw3m0jahxuwLimIfSy1jA+j1WNDR4/Fmg2zVKC8Ml5fLa6olXxffrJECjFXGv/p8R6
t1e/UfU04x2DYSeL/AP4T3ulgMUYgqHORE2HHpRvs6O8Gc8x50Yinmw47nIcDdU5bPGIQ0ok7aB5
W2UhOyoq2x1w6wSNd+/R0KAHmdSYsvTqWLs+4fUYpKj1QPqTtdtgt37i8TJiegMJhmF3aoV8zxif
mnyxiyQuJlX3iJVPM3f4UXPDmwROy0+Ge9rJQGtyKqcEQc7FO1+xjc2oBnGhfSQ4oj+GdsrvS+cy
GzxeRrIWVvFoVPgZEA9TfB7Ii8IeG/dTuFxcl69eWz+OUoWRLweqoa2aB3OVyTDwmetZPfw3yDlX
A8KO9hF7ufvlAIw+Gr2+7jIYrH087lubbejmqWHZCJ+ZYHIwHEG8TK0TeNEP69ULgMnpNVkk/bbP
1hGY1og3L9S/gJEh2GFwPuie+O122bJhuc30bYDlnN37ue+/Jm1V6i4e6DEeX//5QwQ/RnhH02UZ
er+nXCaEIjHpg41GjFzhVz/soVhT0VXMzzQ/vcYTikj7OmOR2V5GrrdA3GMQHOno564a0//QyOMK
AdzV7knhtxmaxWxvqbtGq8eo1CCuXVxOBtx5rN0p/kM8SMV7fnFQ01CCd8J6TyafeFanGotMoMuO
SIl6GLJmee8MjdKL53QhS1p5UbrgksuQVlVK3xEZ4S7J3oPKOZX7f1jWvtU1Jd62tuQlkgkCkCj4
XWI0t48im8nz6cG5x8EmLSYJVeAM+bHSSdsgWlcno/y1zXnk29/4/KpxFzpKoSnRAIUx7l3RVsWw
FjtWu1SdXduudQ/z4pvFcBowek5343odgzJZWVXisxwQ06LX6Mpc+1z0vGH64IU5xtUWfa2eqgkB
XTGyu0wxQsjXwMbRt3QagzU0p4G5LYy+OpH7FbxayWMw+GL7FqDvP2aqZxvd4Mhv7bZdO0/nEVVN
n9HfjfW0BvoOSDCE6jaqnFTIUWfEBu0eCHyBsc70g3Mb4bf5z1MIXMyKDUGPA9QdD2Imo4s3rroO
Q3Uxt55GtlpuzUIL4sGPT7gbp9H2cob0IfP90BbgBgZGmCz7G7Mkc0To4lYx/sl6Ude/ASF2T5yb
qRfwGTzWrSrpgd5YC2Ti0CrS1QweQWQoVszq1ZxFlXNuohZ52UNDz2ss1dxfgGxdtI7ibShj3U6l
CfOzyj+x1H5iQoJ93ZSwqSSccWfvf0IbWhBEArMCtrOT/DhLmAgj6DrIZnjjtef33uQHG4iHkYd7
Hth9FBJ+GFm89lLMn8phpeJmKbSo0zwo+8CqyN2oePBqbK8bZPEBzU9iSWPA4IOOVfGDuFPkdX4X
R/8GKx0mXAhf7Bm50j1B5LALeT+050OklYdxmUlSGOmgP/8fRLMNzWJOEhcXVXul/ayV1m7rQ+J6
Q4+BSez60VDOTyMUFRHJebzykNPVH1Hs3TUaVU7v4UJHkLX0V/xdcWJREh3z8heXvdbAf+LSksBk
Gc/Wx/P7mWtS7VE8Y9r+ZYKKBaWIvG8xrGy2AZZVM2/ALoMgz0qG5Hz9BWjazMDBdD2PdDkGvXx8
ger46iHe7kosFkpELQqkMi/Z/iTHokw+uqLZ74dPOWa6JklbbolHcjwsOhNnXuaf42G1GWVljSFy
mcmxZoVCRWTEZEz2t8oW1EluExqW4szwTIxfw+dy3B8iEysjC/zje3vo7zwZE/ioCLsV2c59doUv
rAi7IIQWmSt1GX3TYNDhQQTSmEcj0efg/JqBnDQWHLh510cGhlbQ21gDHBrAfRR6Hg/BHiNTzAdU
tJafok6KoxH4b5ET4OBtVRQLgKbo4N1H9AEkJdVNrTyABJWbabdAaEjxJaDlbsX1R8XySeUBhN/j
/PkvqvZPQhMykbS2GrS5pTiKIXK95dOMbL/FUCAuAaF8uXsMq389ET8TVkBxqBMXaNSOMMQQlpEM
EX8+oAG7KUJv60f8mVmz3qTQI1J22iLvcufkNxnL1iEEFbZKm2ROkKthJvXuYrXvPouZz9fbD+6z
yMYzbe5REag/P/uIfYctXO0Rnpu886JCXVbHrx4JIgJVAu1qXxp6WizIzWvRJjHPShkKFW/rPfMu
Qr2yxOyNhy+5swYjUkDhT1EccCvXYN0o1FNB05m+LTqwr3qQFmAuWXTNNt0++Kz3UHFMzyfoYZV5
gjTihu3LgGsLRQZe+GRdmFpmcvy+lt4f9Eun/9+gzH9Huwj+lpfq7XhuUTShcylv7dIhoV6BGYo1
KmQLUIV726R4/2m907y6vp+hExswN66HNQunzOb454SZaJNDCOWqzdEiMSIIs70lPywB7dPTKU2e
vZZNDCg5/vrIC4VNITrIN1jTmSbO/bXOfyKSpQx+sDMJ7iHgAKVsu4WvqsKVKqU5vLd6SlU/mSna
Lg7UPlyI6Y/0RCKWAtdcwoxZWV2ajklcLDMbpxYp4kEY4n9SAvtFGUz9MVULRazSXqdPHme+mys9
XZ8r0wH7u7n1+PNjjLzRASONjJn3EE6OxjwpUJ1bKHR3riWg0X76gv2H5qVDTUjidzWkSi6uu7jN
PWOqiIZdWkGV14c3tmydp4s5hhn1G+D+wEULVcTlGmh7w7hLuqNHQkLDex3MHJpLGai65+DoEniO
6euj4cptSOpq/MNEzM5D8Jj+FL8IHGSIFDv3kexMVSheMntbQQ73y5b/50u0HyVpl7F8DYI3lIAa
eqJlwwCEbSqmNd3tJBxN8j+uTqOzqbMNe/xWTmtZHc2aOg4Q3fXDWx8n+hraTH8fgPvmSFtH+8wW
fnCxt3AXKdjAjdTRi4N51zNZ8RdVC3LSlg235R0qqE8XCIC9K6lJ0uHdHd/RRFgj7KUt5mg7QAz3
AtFs03zvcU23YoFGSNiNE25HdDmk747O+nyi/xrp+EdXbfCn4sNqVpX6pImWYaT/45LTJLxVwW8/
Nw23XC/Il1dXj9V+wsbHyJKT0ODSqCGsgiDx8VGqCge3n3WgMeUoeiUdk/zHff18yczWn5ORtA7S
MsdLfKmHcTebpGCNm8yOovPpyjwsVOCF2eGWaDtWfiqsSFgne5s/0VlwvyPyb6TuF5UeKrecZXvq
5GTtO5uLtvNcq64oxd2FOmnPN1C0aFB8ilx+HbQmt4NTOOzyV5Sac7FoZjrq7pRFXvdAOTa6lTTn
KlfOQuYujD1H1MwyTJf/4G3aQbgweWWtntzGE1cHL4bvKlV7wknLiuz7eUbLTCtRFsbPYMKvpjUo
dODFvW1Jx1DVmzBY1sLE5pw45UenvwjDhaHCsU6Ys6JfcOkC0u3w7Wbj3DwU6AfzXDSRpliBg1ej
hWzPFnxkN+AmW5WsdGhp59qlBZKhKjl54Ubc2wlWvigytSqbZYnbWW1Pul3Pz9W73y2+qMQlDL8j
Ndl4hS2oqM2BDRRPLGmWdAV0HK6W4VswXdEiM2Fkos2kVjZbT0zCiBaKYLfryvdSYHlaK7OmEHX3
1HR7hMiSC22k0tGcHlAgxxoJnLEE80YS+5fKV6T1thIivldeU5wMYs5x/os5JcrKnZQ4zkm6rijg
UEhsnp0Mn0xZE2dOsaAK/v5qSHL7Zv6L2f8LuCCNQgC6Dp0jBnEiL9OU4A7tGavjFkCzi7NViH33
SpfnbdV7NKgs1PRdL0ooeSxQaEgCm8v9/a3d3wVrslGGydOvSm1KqG/XGZA07HXTcF6fBlI4od7c
fOxMDfgu5H5p2PUGezXDIN5xS8xj5WmsHse/AFX2q7JpevQZI5h7CvUC/5wA9q9qZgsolsJ34WFQ
Xvj1+OsWbQfJlzrhcNguQhEoIUBzrkmGp4uhVTXLGPzxap2+S6bNv9wwDY7YXz7gyFGhNTRhcTqg
XA3cYRPCSwGd1pEfsTtbN1Gz3xlV+2PuFbP7tpe24ifD3s3zCmD8c6TExAjZS0PmVuZaU7nTgqeP
24g3coMyqPLBA5Kxm7QaN+jfcE9HTdfpr+3UpuFQZMjGekE13juN9fJmzp+1TbxkrmH9I2LPdVch
xcKZwUMiMyhISNOq/MIMxYIXqhYx6FxdVSFlrwFZS0vT5PxpBh9ZlBogQqjL44osMvIEBDZynaj8
GyxsIMqYriDMMgnOvThopg5E6wjMWMKgg6ViwGlrpmdK0gThoAu8kme/u2nHFJk4hpCjxXR6/Zvj
7pEYrqiZNPf7zXOGTedueiLNPvUSEKXEbrKSow3IVQQKAZiMl2GELqcb1t2+2iFhDHG5ar+kPekg
0A9VsueRs1iVxN4rL8h6/IJlR+uhJ6cZr7CEwxpodN9ZaLFT2D5B9kKl0ZckLRznN5I9wZEBBkvG
N2D4OMT8hKB11VA8CkeiaD5VAIO3D0nW0/NlVjY/h4T2vL8Q3ze2M5WDLcNDxy2VUUCPnL6avuYp
irklxKGPQvc6r94tV2BbWv922hbqV/lcHeVepgC9Cg05PEy2Ker3nnFBiJxAo1Er3wLvjsLI0Di+
lPt2ZfT2mcV47wpzEtolMDQfBSm4HoPVJr1A4pWH7VF876zOm+8XGveh8cBopfu+tqWNU4TOoLO0
9Gr/0nw/eluE3P7oe0qF+NPRJUGRxdjQ95X4HH5O3cqxjcPAOXRAfeY2HEzyidHcfxBnlE4WJknz
X5/q4fzpw/oj6kZt4jo/8uZOLy70JYnsOC6wFBDEzvrimxbetL7VHcffF932p/0+Tkf1w5wN1M+i
pq17Hyq2eIT5Dqu3PrsupLoWFR4S+MJPbu91DDGzJyl/rt+kBEqLM5/562zOKjnmoaWHO0ip5Rxn
+SPDcyIFOoyZFgL/8Ussxd6J2JfAf4Q/CXmzssWW5EbMnlO2DsbdB6AcXn0yAaR7zHqdu8y8gQnO
YNp251AXzvdJgh3gJC3t5WK26KSoxheEbjj1yGNyDg4ac+xh4vv7zWRZu0mFmaYEF8ETHpoLm/tz
9vb8TWNicfkV730zbdQ4IUOSiAERA7wr4APP8IJ4aTQwx0Kb13TVWqTYzBRH3pU/BdqpzlQtIsFK
H+0InM7se9XJhwPSuk4SqHmiGw+oGp1eyxtyy6j3yEwyQoHDYy9qMUlTwK2EUJOH0EsEuPuORdEm
vadg1sXmhjj0ZNSDM7gpEA1a8tfhvb91cXcEtekP2cvb5mEdaAy0E9L9apAJxtnxC8Ym9McUY1h9
7jlSQztw9kMr2gohAWKP1E1cXMGbCpWie6ubLRmOpRucFZ1zkkBRV/0oi6UyAR8NCQUVZX1DoLnd
A/mQ4MHRgiG/YMOux4kf7IOG+MgkhLfmkzhUA4qmh53eMG+K9yGfMUC+rj4D0gka5GZAOjDFF+Qs
L2cy3Kwg8dVSnhRtIeF2zFPSmBx8qDwaHlKyI91iVRTJXA19J4afUEuoywxiHDp1tRmq3O9YwtP4
QV2gUu3Xc9KH2wv4FW4/U5KFP1nUzpfvhtVOJRYzTQMpbI91Y1Zl5ZxcQ/eSq1vqyGEpFDr50xXu
KZpsw77UZwl7FOwk1b0TeGEglnRi0YqjD0ga/4un4kB3CDivUjs7DFtlS5uo5AfNXTDbknXLbGEf
z8h/xIr4eVVlRbk3EiFKzhYcUzCEOUco1JZrNtuDWPNkfGiqgQQGOqvKgKR02A/51nJPhyICAoAF
bLlPzcuoN7qkxPkJxDICX4ZvL7NoyEUv3QVP9vQs0Z2HHSpVdxhmm8gYrNqWaDo3eBa671N31vST
IsHLIsYEHyAMnNnL/JlESy34TeulxIRibnIG/+pT7095tL2iyHelveY7a15tpACCDMsGlNbvh7rn
+qAk52dX7FH5PboKfNX1eHMYAoFmWXulZYiHSswrWrZRbC2SjMc0n3cEl3YaVeHMIcHgCV4B027t
veD4sUiojF1ryMsXKlcvTttwdRq7kVrviLM3UeFbknnUATO/1hljuKevhyFrY+JNCOpzUJLydDp1
PeE71dFahfhb3dwTqt+0nIWxbjDLTj3FTF/OQcYObcOMuohjXk6rzqQ92vOt/+nTW4dVNl/7gBjB
9rOJTDDPYxt1M+L5lKG0ZjFBbKpQZn/6XwDr6Ghs0knWA5kZeO6LGAq0mSYFDTYg5bD/wIvwBFZP
yCxh6P50o6piFZKZz73+s98OEGpC2lgsJhHa91fB5mqhre9a1i7iWfXwSX7FCru8hTY7QdvpgmtA
LoMLIpk5cYaVVD+FUiWNqdvUXNvNxNS1g3IJf/JrEYsze2atL+199n6anqjVy5WUfJAS4/LThCJw
6hYdLtGhgxn7SlW0bSVQSz6y/x/e3Rq45N7TmIq1CKX1cvmi6GSuBp6lusBoXPzQhvcDt91K+Bd7
UVtRX1IvrP2ln3W76lpP7zntL7v1aLx2h4to3VERiSwEWNCAQRNsvyXYNW0gsr4vimdekh32kYbt
qpTNhGGSyRzI/k/klvr7GpvHDRaDLfI6pslcUcds7zDpHQ7AcFNHwZFKi1D0G9Vweip63n3GFyVY
DYXNh0kME9ho0RZB3kdH9iGNFcFisonvwOvSzcrOuiD6M+8QS2xgKFexywN4rmrSNnmYHG7URk0F
Hek12rjHsy+0eKVmSuIz1fktJH2xBShwCyjmUyWdPc9Ubhn0pM3KILjd0oRXju2gZAP4ia1SY47e
fwM5vyqFjAkWC2ztBEYEkbK8Q7aYyFtnZmLrG41K3bjFo/iuxOEWR54IpeiIAEz/tp8VmJbJMQQv
cgeBpOskiL+APdq0WEk8nev8nB3+OJELQTGsxFll45W5S+4DwxiPhWsYbk7MA6aGRbbWxwSwb9Ex
XtimN0xgdRW+bXAKDh2Ck/b5pjm8bF/OqjYIw1OvXa10Vnbv0o0G8dPxSq+S3gAPQJoSUDnPa+yD
mL14R5WtMeEQv2Hnzgwy7hi0KNA/CreiW2dLYWLTW/+dJr8wb2V3lcqIhyQ2ojSbPaGgKqJr764g
MEk1hV/u5Vws5Bkczdo53Cuo5cYXAL3JyVy/DhGeeOydl5kQQNzK6bZVJn6OODvA1B7SnwrUUir0
ULlqXZU6KmtwEoZFMAmYhzeqboJokBA3mwSXAq7tmRqfE3Zybd0akZty3df3skzw0r8SEzq7LydH
yufpO4H7IZi+szsqWLYUmNm2Pyt7vIlGzmWChmNrDOvcve0GPLMCWeDRSqr8N9R9fF43mGECn/O5
WCtd4iDCnAqtPHGnxAt9itlGK1NKMWPYwW0KCn9lsl9P1UiEm8Iin7S7CaDz4tCXUHOmWFy2hmOK
Gaguhfriz/pI/dgM2gzeqOMGGHKiutxmSqonyaNAoQtVkGhCeTBP8r6jyQq+p/3aO6dJHwAf2sB/
g8nX7Hr/tnDxOo2YxFSDvV8SFqGG3I08lYmzIZUaYtkclsz1D1K1YmKx3Q/oxk+19/tniB379GWt
fFjjK/20isAmBR+qVcCWBcdVAPFzOZn5VKcqjPJizzuCVe3C+u6yy6tjQgo3ZZVDR0Mv1fs8Aehs
ak9RT9LPVM4FxsRV7OogmvLlfpTHJWanCDDKdmGnRhxCaLzQPKcF6HvzC+ix3CKLsPFKLA562YUF
hpK1hEGUyFPDao4GraHlijwX4vvqv56KL4MuCVLKHFQCF/IUycz2e5h/A0MJwsSculPl9xFNQwNa
kjrJTv64TF89tgw9TMeZOFH2cvsRSLosazHczF5tftNiszaiKfm/No3L32kTVdv6ijDBRS0nTGYg
qy4VRHlwiFaH7XyLd72qbUWZ1NeEbZLw+4glJ27rTC/8BItkXR4oE/Cur8x/sdQHFLpMW0Xf83QM
uf9axEPR1MNBJpsjyZRG3fvxonxWiIuFKHJFDYNCPc8YgbhnFxu9qIQVA6r+soq6IiRCZGZX4eTe
mo4z4XIHZlmrJGXYA3GyqE0H1onyxEb0aDZVgkEZvxHlZZtauL8FLnvbA4LcI/rn4OWdPFEuNRkC
uyAb2BplAc3zdcvdusQ5K/h8mZABl5RsjFEfrSKbMwL7AZvRFg1JdjG1c/xu9rqLrI/B9pFgcaft
IE3xqOcsEM6NmB29gAE8z/Kg+memXv3q27X9BwySsdtPtM70mW5ilw1Kg4simTuFlH86J5GLckh+
+xtU3Rg3GCciryejYgylIcFX+TzCKhi8vZDqMX8EFiT/nwwW7ioH+CSu+NEQ7VMgO2+hiBAzQ5bF
Lt1YS1arL8N8mkQiRw/ADYM2zw5h+dda1c7h8HnGEMfoSwCXV9xva+fh5Qb59WQpzLQOrjy75U6i
CSvl9qos8BVLQwnE1NAeZR5/wMNwHMM8FqW12+1tTQ+p4qOZ6L01CsFcXEK1M/AXhcj3kL2TWwaK
m3Zb/TUpT3PgZS1yfEapsKoikDHs9XrUg1GQR8zHpY/OFWCN8e2+0XNsiyA60HcarH7Wa5Gfg/nv
EAqYJZNOofrTpyWk5YFo3XXS8AMyYDU6LG4Vg/dt9V6Tm8XsRXpi3E7HAbKEd2eEjqCw3qS/aB3E
5AS+0X4jNrmMTWX+dNjksxpkS3VXgza+MlD7XemHexrTx3nakKREhNZd1HcQliAyWxStgwadX+8U
Srn4y6hmp5VnEcKHBkyVH6uX1r4A31F1Tb7qe8fJcmJ424j0RT+wyQrXXld1typjNWi2ch73E2m+
hCZUyRsa4R6LYml+AOr6ViE48lZEZ/0g8qX1+Y3h6WZjoDuvV7087y0Y9IP5lzmoj6gOyqTABjyW
3ujneNiJ3yPx8O01mTJKsC2Kdc8qyScfXAv2MczixL4T/SYbFknFZHzWzj4Z+Nx50jeI63Lbr1LQ
330b1wPatRzcjoVq7v8tMXtPjX75BfmhQ1rrknEUcYuhOheVXf21wK7LCGjMsMRekQdTSMyhPbH9
jGutbRC3eJNbz7zRDtvtpdgivjwl0DmSNnyij1iPjgEwkRd57rDGGxSxjnwcPq6cH1kgepFjjYRO
TlUMuiwWg3Yf/KR14Vd/PkDUQhAh09kE2M55uigGTD/6CH4/oHdhP5P/FtrIbC8C2wS0RrP1SKnF
IrC4J5PmW8RCXYzL2PBem2CgzYCcdBXFjF7CpUJoDLeXtqdbAm1h+ANVfMpitU9kShxdz04/cAS/
PSz3geUXXrz5IgWBS2PYwX4kKVFPnoYvJ5rlIVphB1qAJ2tRNb3dVZbewvodd4giIfqy9T55bR0s
PNiosxmF0wtqZj2PumEl8uhpU6H7sG7RdaV2LEPwljdJS+4T9Ft5M6cvDYC3i4cRvs74IZm/6EXS
D5AxqQ4PSKRWsoInBdQH99o5U+Yq+3bHU5P8iZWSw0krGN3ylMlPfcxGpNzuHE65wSFW0caZWNRH
jWfABPf4YlXjfiETARDseHo3mU1WvJ26nDuNrXjrkrANxnNVbLSIzAVqC+yglEDDwFUoVBArkB0/
f2mUzzqtu2754Xd2Xr3PmLxHchtahpeKmrEp7YuyLnvfXXKN7D9tYrtGJ6Zzq+IHD+b/qnytEa9R
Mn+MMCTYg76U7zSAqgJwZBh8rRC1nw9kFUC9ea2Mu0cRAiynB7eh2t1rVG9Y4pmPWGbZpODgTErg
6pmof/NAwyEHSpI3/TcAFGEj+SxBDbo+m5vP1kISy3sMkem9aiNKkTciAOSJoAYTaIpZsIbj082v
8B8+EHuhW5ZhLMP9qrdGcUicbFFhGpx+F0Heka/tnCqIDXS1Vj0PWqlla/dAqrQvdIhwVdsdl1a9
kH1UEBKg2vM0F3GLf70F+elYYlS6/XS6/j3y1L1lf3m1xVd6wM7S4Kjyo91gtDgncgbGMs7M+KpR
2mBtKs9d09WWi7dq8AN9ST6RvgOPTSk/1vEOX+iGX7Dhv/j5ME1ts/kes3DSRcbQT47cpQo2ODCs
iIMqr0PYysnoym3jdqRVowtvDnUcvyt03mxJQJ/6xhDKQKqiUDo9cfnCRyCKosxqROxquK9otuhP
NZF3NbAP57OGOgPKWCFa42x0kMRr57SDm4HGOwLrtan9+hHiBpqBCSC5n5AUvryZpYtxoODOtzbb
KV93qA5Hnt6cGPV919ntkiLE44d8O8vrFeKhsxkZFtZtY9+mNojJotKLbWTtErWw/vm0dmp8EJ12
4AF6zO4rC0jLooO6NRRs9UNw67dPH7rw3fqn5HHYX509Vwyq0XF7mCXsw96teb2OhT9Klyj2EiO6
QG7fgwes4/IOtq7/OZ2FGEUHODjYRkrI+GBZ+wsiAjqAEwPvg0gslGtYE9U8UhA+g+uitCIyGQXB
87mHFkXBRAV6j9TbAvqVDfZ4ulvRa6aFh/Y+5qoSVXAL2HlHrcURJqA8b5NLyykanq/ZaHquasa6
XM8zqBIMwkUJ/GGs5ttxHaCe+JcQ+2xErLcwSSegAnVfRYbzhefIXR7t26kh7p8xpgzJq8K5Z0D6
0rVLK6DoxpLns2t0X613G/7Fq6FlP1dSoYMw/+E3/9mmLHP3cVm4C+g/ew/6R0XVK9zK6l4SDNEE
c6EhQIgWsaCH4nu1VsHmKpGpDFOXLO+geMUWDwM//R31D09KhtOSYu5aI5agtLp/xvPRDLNKD3ua
TEBApormhBrVIZhCuDWoXEWeXPXUiEsUOgPzQBAZHKCStX5DNKLy+VTeGskjy8jj+9Z+8gJLjlmK
fz3CGmO440QtEKxwj//BhdbMT7C9h2QbHMlx9Sv61VIsNzeB+aEY3x272Dvpp8YOZdk2MPEzRwJh
K0cH3tQvAQaEeYjdNtugV6n3xafaaGUi3/QdBuZwAS0Lv7u+CqXkjiJoOiJRaJb1IaJk3wWWC+5N
RFz4CX2z3vWEXbYJd3RgAPvyjF83Wxk5YkjFxhpgmrfkkIbJ08c48s9m2TP5yio5eA7UG+A8xUJo
PaZ/wSu0oFh6lXzc+kiHJ2JcdqbDHHzmvMjxyLPrTgucG2ElzG1jt3+WCq0OoTEVwQyKwIOQ5UIR
6ZkjeQ4R7sZ96DQUAgal2iGoBpg2LIzSBukxSqiY6bb1QbX8IKZ623XPhBzy6HpDWrGMUvs8/LFt
WksxScIYkjWVoSopGSpOvB+Xb81x1aCcxGqqqu+SUigZzhWP/Lgt7ETZkj1ClBy8Lw3dG9S8mevo
3CPjESDRGr2dGMuuKPeW2HJ6BgFqPuDPSMGedym/d2Ob37zx62pqKl02dSC1WvIzCHylXYEE4K/2
2CwVEVNLNlEMwHt89HkNX67TL9v+94ygz+ZSzeNvRUfC5PB8cfCto8Dx+G3WQQL4pDFB3kbZGzny
uj09hP1F+iJned9dEO/0exVSSA2PGjJB10/N0Z5i6HUua672Eqhx2o1ArPhnFFpa8IAdUpwM5EmP
QMq9qY81ccXa+Va7ZbC1Jz3UMvswHVGXuPnz7oL+QO7J8ghrx5QBctsLdxNNuLCGNJJ03jcqxS7U
4gkt/mVkU6MWQEL4d2vvvV564z8iArRzeyZ9zkQfDzrSdtDygYJNJ/Briptjs1zxsQzJtHDvJ/oB
X6PQmvvQreZ1Bzo9Bho+i3tHoRfF7pHRQtK48yYkuyx65IvyaiW9Ion+ba16nTnCcIo18OzSgfla
JFIZiDH1rgOXoRzvRiszeZGJL8fzmWxINSNhDCUmmUdNTmFxwaNDii92pYD+nCO2bJ0FvFK8+0DQ
1Ohe6z1+QrJE3gd5MGNr7DUlx5K47+szaZ3gmHuduw8RW2zgfiMCyWTo6MnDLmzzFiEEMT8LgNoC
Ijl0YNoyzY9VREyPBhMv4F5jN/Gdd6uKp5YHZrKiGU8qMcZ6kv//ehcAIu9+P4SATSj9i3eU54WM
mkM3sGXdD+TI4ckOU7dL9G1lzuqzVXuQsmUBIB2IiKWI+m59FXlR0++uJB2ujpXVkyn63oZuucW8
gA79RFq3E/ZkzEQu2VFmKjolRb13UG5aKoKNBOgyNVHIHit+xyDm1W7y8wpWINKsidJbXOa8kXxL
5iMRrDQ3xehkpZXiA3cQtvEAOkfNHcUsODR2AfMQtkvVYPnAmv51TcBiLBKnHxRZjhbodsnRtd5r
ohk4VOEjn2f7l+XVmbKxrEe1LYr3Gynd9ENP6ozU+q86yxozp2VxKmH9Vgr6lcFE1Sljb9frpmRB
qffAgeB4O610XuArO5Zy4qpVlqF8BLaMelJTRGAlbEWAWqCY1Ptzx5u592hTIl5gJ/oHCsa8FOg4
BVcDKbjvjtUfMgiY/EBVF6wT2PD5i+AY0/iVQaAr1TcsbO2pEcNlk8k4AQsC+gwqKStAk/HLbCws
LW5HVxZcruGDalSzYqDyhr0wIt79fyh0F8WpRlHSS2xiWLs34CaJKeGpWeTtirT+RsIW901GNcz9
5Dl90NhV4BUsnDkKuJ/lYkxG1rGva/h7//2aWMjGG6M9p+GYqDxDK7AIrnlkJpLgBud44OHeZpP4
z/hdtQ5mnYk/DqaDJWy089SziIU6D7ppQ1sPWXoEreK89lKMFH8YjE8JD57zNYryWUUHbQKGKeaG
DkQ52GwOLTBlmy9W02kA9smbPaKypZDsyeNG+eVw9F1B/zEMFddYf+DKTUNN32+9v3L8BmWwp3qD
aRK6or9s/s9FAAc0k7nDodcvQeE2h/4qUf266Bb8YqO+7eNbMeJ3t+lFYGJN6FGaw3+A4z/I4sNu
KCn7mYbKVelw1bB38CsevhcGVtQDAIV/V3BtaRHqkyOASGMpLOZYdKWn770YWztGivoDEmuuZkE0
LYdWEHi7gEZFhLGV2w6+UgjXJyPvRX7VB1AdctZMdH3s2y75y8ZmLyzOkWvhg6o+WDzqzbtkWaRa
B2HLxn5Hvica+d82xDOw5+6KXnuT8UY20z0gp221dgLt/ERpf5MQYFmS8BSVmgyuk2aCzqH2LZ8I
QD9Ak5CxxuS52hMwhAjg/4tzB7IvP2kzC7DXkCN5H+bb44WAWCQVk/TKAr6HAiGn20LW/qeq+Fb/
wI8YJgSfWRjUnDdXa+u+ZdfNNeUiZe82pcFSi8K9ayj1x+JCgqRHat8PubnEue4kD8Zurm2c/7W8
yeu6CTpqN8hbR6BaiwK1ry4KwuL70NGYnFbiLpuoX1hiYh1eGFqHeuv7ncclxz5z/NVjZs6kRUoU
uGIOMpuAP5Y/iEjfciOUKDBi1VOsD5BIYuFYP/7ir/BOhGs1Qk6hZNUx4Tiynw9NrV0fFfcBiNnB
ipzkiR9R7kRzoHN3g8miMNBb8VnHZuTfadsCKR8YyegqY8H3S76f5udtFIVEuoB+NCHPhllHCd8k
oPsxBdKx70r/HEbWqi3227vj5cnm7IJjTu5RAXfILs8HBb6k0NWhXgIkZb7Eno6dIwDHOptGDzDr
i1R0W6DI19ZuF03Qdl3WQdn8a0Vr71AMymi+NLYRzhFHpgw8ItSLZDpROP/pYgm9nfD0nCWmuYab
slgfNi911zxdyTMCNRbhfekDDRL9wlcgkaMvj72qAWGyCFTn15lWrmEvaRa4BYltdp+30YX+a8l8
pJei8zFPEIq0UFb/CZ3HTd9bCiCcJ/0euqEbt8lWRiFRgnDRZIkf6NrNPGOtcQHlS1gWbPN++/eo
ojVnyF3Ai5OvBjRrnX2CJUJPK56JJqgyPXlk9lGvPzm+GCeuRx1XuQoQV4km+9F6npq5TVr0F6/l
C4jfutJKXslPsFJx2/DTggq1clvTUTTQcR0+QpydT8gAt/kspR5X+PmiI0vHnhZxqTBU+Q2QcUAy
yVDuUHa/P7oqV/79YqOe4yyVqr6Kxe8amNklJMq3AztQxX8SB7cz8NvBeszmKajqAlaXB1bP7ae0
O5fVn7AjNbrcG3DQBfds503zsDleS+9hurQGlETzMTeh5sBv2pr4lUjvPPYcsQVCymGCY69p8qom
lOyM4jtb/eOf81ihrX/9O4xyOtejzX2MPj8IGxF76zACgLrFVR0dC/O5iHguZARetGhizIlZwGaR
jpJjLCmnqp8F8/5NfltCkIIul6wHbO0bnMyzK9V/LyUaEyxrcIBr06mXyKOxTtlD4X3pG6CfgENs
bSUsqCzLqQExOFhv0Badu4wSJczqFyHAX05FhjxyWRA3NiU8/d7+hoXU6phlxSWNx9QKiGAHMiJq
7JaC6lnRSuWjjKwG4/RAGESLq0nduVjszt0VnUxf2SMCADhbJ95Qmn5ln1LsvInLQqSa0go9hoT6
oSqn2bxS7KyxnP7H6eZGeBh0RAYF+ADx80XB3U3wM1asdtRHflBS54dt4dL/YgUhQ5MkhkV3X4Ix
esx/4VGx2dva2HvalqdsSfX2rcVHWaaiF+RqeR1dGl+aNN/T42cADTZpFb7vK48TejV14oOmFN7s
4ziMX8OEheUosoey749RYNLtbmMXQSCVK39GCqxBwvdWnjcTYOeyD9Ke43XkRRlPaIHxU8L/MGns
LT4jlf80UnZH2DAYa+EMLycw+++FxPI8VNa0yla+RkQZDN5NESiER5USKgEJHSSDsiDLRdq8U6Y/
9+xMfJ6hpIUJgtmlvykB89jqbSeB1RWuH+zUx5zGYRvy1cLzZoL85IUa710Bsi+Xk43danh/0MvP
MyUC9qXdcRsV7/qqqWGJ2FnG8Da67sJcA665sONtsuXyiUVuDvFWGIqaGNEfAilBUW84e0MGV8hA
2cY3sV/pi1xoVTdkfjWI/um3epU7HyTp3DP5dANCQQC7t6X++kxwXpHbf87MrXr7wSgV2bXwTAXt
IQNCktM1baZp3ePsfTbLDR+PqzrNTpMISbqfdlIIFmB78Elh7wJa7exi/NEPwGD0B4TwbnIvqyl7
2rZK4qOuqVXbWdaAKd4rV48SsvVfK09Vp4zIQblrI3h5tsGV6PIPWYzXSw7Ci8MTm7Pn3tb8+Sp+
9i8//xTSwh+eXlzmsLTFNJzeCjl9Lt6RFe71BFKj5NcJx+EeveIm6P0NJx9/yoYC/LYr7Rn7cJLM
AcwW20Co8bk0Hzx+CBsuJaobdovywSKDCFDI9g38CE3yfEmnuXz+zpel9w9e/XWSmJbG/L1vsumC
2xNziDT3jTIzLPS/1XLw6/kiitAWJGiI9dsKwEpr8ZXIxL7UA3fJJBdybyia5O6YhH/C+RcYppj2
3g7PYJSAzN7zw+KG6cufXS+TfOahmBLf8vEp1FK5UiYZRIrG4vnrMEtc3mHKXz7dE56Jy0WUzg66
Vac4ovoi+DLxIuWEb1my3h5vQ/2ebHDRk9IbuEAViXAIwI+TdTfAniMKcXxpFF+8K2T5lUvwT+wN
RzPsjpn3Qw5WLWu7fJAcS8KopO3qSrgOPXOL/i5YZWbZgyRDNifvIecztStXik1lGYWIM5QYujx/
lKFezhgYNNoihF34qaApVXP2t+7D3kfD2c34EMnMXcMUaLT9AwTilWDAWbdrpvrGaldUte0iaMWS
GMfR3Ldx+Izw/gDcmuQ0ygcVy+WH5+Q/5nuK4RJYwWMOnVSo1rrCo2pETNYwCinTZXm5JsWCnhWm
tZMuB3bTG1DB4YONgaNP2TB6KXG7DI10+Z+IPQ5iTqgx3G7m/vIuVUlW7elC7xY2s9pTMygVovPB
oOwDIgPaoTs0ujggFQIlv1oryVZm92CMg/2y5DM4sVvuSQ2HaMUoRCmz9oFMLVi2u1JMcxVCSG0C
3h/l1wSUEaJTOfUuSp6A1adSpx/Vhzprl6x+WeyjUa7TISWQQ50OqEGbIkNuZnTOufK8jgt1fDSb
zpvcK8nnVuwI2OfCvK4cqoXbQ9MbRHUcy4WSaM8l0AOIMQzLyRS0Ow/OVSsJmS+lSkyAgLv32P+n
n3t7q6rh8rkmsK8K3JA6SVz6jpN8QpTmBj4QSq+PRVSfTpkGgOUQpyr9gVauMo8LmDn4KTP0ePiQ
/U1fU2QR4Z3lCrnXOHx64oY3XsQ3Rt3+56hpZDy3/LK9YFH9Lh5nLZtBmsPwKOUHwteBSKUK15/C
wq7gmHnOfoXaeuEjfybnt7ZmoQ/Y+yjkl3IqIXMB78LuYLUv3dBr4w6LXbH7unDkO3PzmQdTBj3R
tgXTsnT0OInntNkvPp5DrSGyjZMJupuLphmp0aAglW6zsbumdMZ5mrf68ZGsQUs5wOuQnxYsQ4Ah
6gXaOcwjDYHuKO/dB74KhOoMHXCVSMqw7yR9zKP7foLk6mj8rAUvBzx/TVLS3EXFbUAjJEC8QgT7
BJyfkXDZniv1VOLZYV5IgrMRH4tfIZuIwEfwfXLX+ozdW9/E9XO2C2qGquiJtl0ZIaOEC0DmMyXb
zLsEqSqwcfrNmijyNcyO9vETFcBkeCkIRia71dcmbJZp2y0spS9kfZjCuhw3R8QR/2vU2bVVC5rR
hLpStCuA/7Q9Ji6Pnlkv25QUdY7GUORBKMjPN73t74GLROamqBes57FhrzwhcEAFMg9a/itfZ2UU
0nQ1n0EHesfNOLbJ9Fvc50AQtXyq6AWecYjyNmU2p2Mxq7hXwrRruciIkbPpcuSdYbdG3gPyqCkn
nRUwzPanoAi/pUiKAP3iBrmu8pfuLYAaEH5llqX5LzYzXnVT6Sm5RbYpQ8V6Vk+Zokde1d7yWIHl
4eawMoKU8udWIlejALJ8lDnNpgoDu5opfQaIc7fCtU8CNUGB1NZXPDqoHDu8D7/TNafUFEDreOXs
6UhNJMtwuVDh+SEnaaq0P6e9il0P39n52EQEWT2KFW6rYF9zakE6UiHeCW66qdDJ04diJX64HZYJ
zQPWPQ+T2HNuOIjCTxQf6XamblbTJl1zAbo1UCm9js3BeIdpWLRLjLDEaXEy64bAXsJhXZBrInLF
H7L6PoJakUddCLTVaYolOBS/6QwKFzbIAOEp2H1yQsPVB1jTjBXBbxpyzgCBbpcABSD/rYnc4qcM
FvF+TwlSM3ho4ymGTuZuu0SU29B09aKsMvNWwUOqzoams7N88/FI0kQrEjyjUleWHvB0dYNayJ13
6BSgrvNasuSxZ/WOmNIPctVShheh92KZZ0oBsD+etQVzJUR4RDRJX8wfI2FF7EB32+xo+KlKG1PL
De3tqAYN3BXz3w6cXgRs5CiP/katynv4pb5IxN+9daGtv/7g292NakuQ/lqCr6eA0yVZq5lS2bLI
GYpjUc6MTcq97P7WfQ6ibb35f52GsPMlL2Jgz4eP8bSUnS3M9HfG5hfHjNhVT3Fo280RbAuf/8gG
AsgbjOQdG3p//usgBlppiN10f8JlRLP5NWX0MY3B78SDrcwMU0FxlaIhoAReQR+h8nzuwVrftuhv
RdTAWRHDAMT6/tr1VNYJieIBtmMQ1+NJI8ujjgp/8AWIh5ePTto4RUnoYwS54g4Shmu+f53KRyG8
T8pbtFl6bgJLzCzsB2Pt83NJjU+1VplBT0ezJzRYrzixxg+9YLzi95hUs1+bLkHBXEpokRYMLgk7
+xO3H+852W2s1vBSoFzL958bt1EA9jyZ3nxJbxW/uGMKet/UusM/PBzdzM9SJLpGu32uBAzXD4Wj
Zi1eUKJFRIMTq2THBV/iwUcyzd1suJ++MTc5E6+R2YIQkhl0Bd06epbKp0uDBISBOS+oWl6N7yD3
gFumHtXnTM7HjgZAX92eBE5DpH4PD9jdjNI5lM6C13rAFYZolb/5EfxfCcXxAqP9u++4z2or3I9e
/rVp3JEN/vWB9/JcAdoq7TFKogYILP7yuSngWnHjigkmIGruq1mWmSpcixrq3UxQeJBXG9WJ0Yh7
8jjTKN6Cz+VurTAAxgPdx70IbRbMmw1uhcmeWIOjDobbzh8Qyx9jHdx0lQg6KDfobfx69MdUNFL+
xAo0rjhWocyfk3ETyjLJcrvlUQwOPTqbK6KUI3fSNNmHvgUHe5yat3Vc7FFIN+C2JTT3fbJgaYdH
7SvdMl2mGBqliatlHr92zRQ1qoGB5wAoetRIBpKLteX2eI7um84894lj/l4hrvX8SKp8bCRSKeYZ
WEANzOuY9shwbzNjkqFz/loO5pIpeCgBxBOU7T/I/gLY+NuAH7mJ+mFSzAADxvXR9W4ePcdA9cs3
I49ngnIrjqXW1utEe9MY3nYDevTIkSwbPn2iGiftaD9RoEaONps1VhhOQvpTOVvt5w6MVqkIG5m4
aJhrwzGxw/F1D9NHNIYukbWslVTTf7XJbxBcCbY8qHa7CjuX7a1gK4pnHzMlR/zBSJVpGkNXDE94
4SA847KAMYnrzfHrYqcDN6GltBw+GWqQuEPFXe9KUES23Wa4QOKbJEBHH8ePzgzr/PRWwHsBmg2z
C8YwX4yIsnYKVu02u54YP9uI1YE4Kq/voy/cn16JKMp92ChZq8sWVX+XA2IR9yxFq05s35w3iFQV
5nG/cfw2GnTjRCeGBWprQrwNnVMQIyQNlqXmBAbhI0/H1MzN6vonjXffL74DExdkqOVzBfVZlbN7
vam4wCqU9vLdmpI8anstUEibsPMssO65P4BMOJ49e3GAcQVQwDTixV72HoH0tQlPXTcfwXiEXUzw
TH4uggscspdZTImTtg1kAYXxT2Qx70MpMGrz9cAa0slCDy0EmZ/o9O5fKQYtNqdRb4zkerwMNJ9e
mP9Q8HD2SZ1teWVCSuCOhr3iyU/+VHQQz//ffpwZahpncGaDbAsp5if7vq9S5R/5iFQRheFViezU
Ai3wrjY6s9B3uokpZ5uh6b9EX1jrPE1ZZ1USCrau2+gJcorQv2+YbKxygtbGL484oyyjBAzzEWsw
M9uY/FYZ/PttBBOVcZt4dMz9lxacbxMJ6MYWjkKqDPJ/UZUDd6IoyVCScPdTriNnrc7YYqq+GEaz
wB3WGoUK5G7f8B4LX5fKAjJ2t4Vgm7Kru+W4wMwIB1iF39QvSj6kD/u1jWo84owxtX/sZb/O+cf9
gA/ePNoVa9IsWngufmv7Xz8YewTnWGgsOV4Y20BMtRm/1DE5AcOxcdoW9lJTgVyBU/sFVwciWDo8
VIBiSuFkRmEJzr6EkGwmneyfQhlXmrlo2R7l5zPUKfc2KOdlkbt3vJXHjTYFlYUHUP8G6xTkVytq
JZe4M9hrAtAC6weRVKQmStT+sPow1AnlLc4P7m8ltRTKKIbdh3wBcZX5yGngpTISEHX7wa7qfHAJ
meUjgtvP5Ru5uukXy73wCbBEiEETUozV52v/Fij7rONEvRFvxaQbV4S7bsgbmBt7GewcFxvm5bMD
kG/EpxxJu9AqVy70VVBxSJYZOhAoLv6egFVPBqcF4s1B8HIEAJ+BKTOx1bGBh/Ayytllxo8lg5LD
TOu23d6+G5vQNbv76HLbP+26PD5tyQYw932vss4XB9ba+2tSKb0LyfJ0hZ/lukEv0XIukIvjv49T
+mZfpaWcDlIfWASO5xk/CVlAugA6REHb/dvzzNugRPNIivoEuxylW7woTY8N4SxPleZPIvU3qTth
33ZDe3BqxP2bPmf4iBXqn/Tnzlxju6FLeqMebr+aBfbUwh+55Mr2jK8bR2Q5oEypAhhw+e92Ybu+
7kcfOETSgXYi8WPn4ZLxndKWbf+2mLOA5ESkW0pXxnI7sEGpe8Opi7mLZmrx9Kq7GVjFLx0oPDCV
ynZkLEbNnvYRCNm9r7GUrBePB04CBXm5D8/cUjLJJjpNJVViPwavLXhc6ZGzB+uIwnwu/FCKFXhY
L6wy0nxHtCq+d+j0bNuMw5nZ2cTQdzLWfugPJiUfX1+NMO7qpbW1umg+FtC0WUI562KAozYJ/qCa
a3xBKD2y7smPquzUih6YNbq6gr/XioTkW6/sCsL7qw2iD2el88GB5hIy91JoJsyJtKLxlUJHJiOf
QAuGpEi8p2UgKra/2BucIvUVd7pBJztR5uODqSTxHM2DyfPbjgFcMMWfJJav3a0A+0sbvKOJblA8
xcD1pNCRRjaTXVbJbwPURNpcPWqHh+GqDdG9UOPdUlPp3m2hJk/txl7LQAYcyW1WcyCdtCjXCzAj
kPN+7AdxBSEoDz/yzByltqR/rH+HWYhHDstDt9miHMEWZN87YwMnZCFICd5xOXorcLNa6xNg17yQ
+yMPFsTzmeg/w92wQjXU2e0MFoKL1/PpEzosBk7Qaa5cIcuMSS+2qX5kr9sWnwXy6Whiltcq3BbZ
wq+YArqwB0KGhCgXivvIpRLL4X9n0yEJ4RffARKYc145PM9Rbdc7Q8vfJW8X2gjlb5NFlpXr2kUI
XXZ7YB/18rUYXhsd3IBcPtu+P55kpj4osfNT4nKU36GxWlvTW2kLsipCnGl4XHg6Fgz20LDpnGpM
ejxjMe+vLtFQ+/mHl7GeZDtXeEUK3RBnPbw9fdmfQNMzVO6Vf6WL9cp3x/7FW6RrYxwj0xhzR23P
SzTsOgBQdILXsTy8jRYc+0MHO9/UW0hy7s1uhftfdklt43X7CUFu3wi5nSmqekU/BaR9f0bY6j4H
uEffoWk3iKJGwNNQD+FN4IDXWWm2VHfzI5AK5h727l9OZeTTQGeY/Btitee5HaiQ8NkNMQFOfwmz
Qb7JQP7LMmjyBxrpfnhc7NIqA/gKQWHiUNFymq56pSiCwPud0Jy1LhEUdwUabaCRZtLwTCVB1LMX
p1YIhe1/dWGksGGld4EmhDhsq9F4bGglMJLoFuClkd5U+iLJe1aT71tKjKrIP/D1/Qt1pa0YaYlU
MDp7i6lfa8DPKqreww23l4DiDP8i7vnO/yr5SjVoyE1NgIOEPWGRWrUAbFbTGTmEkFsuinA+qIuV
dwox5LktvhHDMpc2xi7EdPMOPGGpV7czXYfmqORk4W8FOo2HiOeQRc+SGyckCurch5dII91keLMI
bG+zYZWYYr/1fQYvJRIDwHvvtTUnoK6VznSw/K+RjmYYHFMXTehM4QdKbET24NmhSh4/y+aU5Jmw
Ax04W97W30QFGh4X7ZqRuGMd/3rNBVPheLfnKMZGCo8vRRuwy60yoRCd6DWNnmK4feKNFJOwEC85
A9yBOSVNr09xnYe2JJwzXx/B630+LqvLDqesssoBpqwpcofS37jj1uD1rP7kqmyi96x5Vy5Kj+s0
/a8hWUTApwGAnkorA6+CsB4nvcSlZcdD554TrQdQMyDVpBow3flwjspTHOTmiHDET+J35q/9yeQS
YYgndMjTyqyp7HQ9vVm5rZL9Vh/pwyZt0iSVPllzPBZFExvAh4k6vcJ3/I7TBVCvbclAX2L5ex47
s2mE8TrKahMgU3lAOYvNm90YZUbFVfVwepVvAD1uKre63MPuKRvPsCYz/T6bSuFqRsWr2fyg/OQF
7M6Y2drvF5smZNgQNtMKfuX4is28SRPoT0nP19fsMNM1/ZvGOHiA8EqX39vVKXCauKXBW0oJhdPU
IFvpD5ITptmGd0pz1FFu8SPm9OkZgS790Z6UXrtf7w9ork4tNOyhCf2qUKxBsB7BdeAe3QFHzSrT
xwgYbs57GLEBsrDfi60DY0P93Le15gefmjjuv54KT5EpwJtOQU88qoKkzAT8zesjyVeCIe672P6R
Qy0nSUxCwgkalUDloj5vCw6uw3c3QGzzk+2PgB4b+MsRKPPEg0h21eB1rAxM5OfYHUfAXsyriGpS
vhvHqr+ah1GKYMtzfG+nL/vcz4gr62Jd9IqZdApiIQ51danPzyXupfeFk5k3UXkN/qMCmlltj9of
oeD4NrVvxwv4b4MzF55rAwaoncVtRhweSGLoUwhQIlyE5xtcZEvLPGZI90fDg2o1Th3GBKXvQZQE
oSnp8wPqnE5uUnBm1+zyYlfPIqLq0Qbkvpc9XqHHkmcupswoTB4KUuFrDm+moN2CXGcTE0TLqRJo
h6RS4Tm4q06tsKMHd6YmxcXqmoHc4X1hXPRFAnd4Oo4zX1RFE3dNR8HsoARQGIUmPfqEkb3xoDTR
zzZsH8oi82K4oOhBJAmEaQALxnvnuhHLiNVb70TXJNVRux9AmYKZoLdIt24xqzX3C8lX6bhFVSAD
6dGhPtk0gThYNvX4FJ19Baja5DP10GxjFlDypOGw/389VQNzLzHlU8Y7+wt75xeeoWjmCvUq+XdX
Y3lVb0TQwL5IdIOfnok3nAzJgmDB2LKwuQNzM1gqIXQP9km2eXpK06uy6TcNts3u6Ix+SCdKT/gi
ACIG2O15YlBw4bhzRrGHv6EuIaIFHMnP3IiBN/4lbaYH3eVTWbgzoqauhd3jKaVN+wEx8yYffhXc
wNC6ovEaP/YuQYpZ3iYTjxNdRrVR2OF0vK2GBZD37JUbhSNEVz6sKtvr0SC58A93Y4lehDEfGLeC
I0Su8XY+Dx+Uit/PVIYldaCfdDRQ1Cj4WOPfaBOthpwkgHBARLujhaphaPW0poGw7I4RbB8vYX2D
DHOAEBXBBpRcWZ/ofm5SoTCD36bgkAw9A8hmKdTBcQcpG7grLOE7dPnKc02NciXmGXe5o8fVR/Rh
fNq8Plh0oyQMF3x+8XShLe6GAAHru9G6u1mQwDW3U0HX+v4ExTEXPq6CKI9xIEkMJcbBCgzZYSIX
ZxTqpcbW6uyfZs+/mklrh/+XUUuh/XzqJ684GBqWCbwuxDarheqIUF16Ppe3Ta2gdW6+b37EOSJJ
DZBOZL/HIpdjfai8uTkN8KIB1+0Q3McwecxiUKPt4iIhi54reVLgW4ZrCR8m1cYQmJbMmMa7smJA
UhkpzRNs/KtVStquSRco4GVvjxsbeasc5vbivRIocMzRZntkcANtNKSYGCRT7IykJdLJgTNMa1V+
8ZvM1J6fqGQzCwKj2n4fmB+lnA8fXIMqFlN3x/T1D3Nv3mJU++dLG974WbHBRwSlt9vyNyIP4TT2
pRcym5v8cb7hjWQwbdFpCZwHp0IEXUU8aZc039KtX0UpjF1d8CEa9u5hGmg6kABvc8KJsYgEn5TW
tjKnEPVvWiqO8vj4HpjK4j+BRly82BtNlSuDJPyY7t6g66AeHS1a4b2glqzXZQYahqhcAkvMFkKh
it0iwLoUwQQJBnJoj838usf/+boOJmlkkvZDpLcMG8pUAEKjUdmK+PHgf5Qz708eQ0Dho1iAeZqd
RG43okaKwXtvDoHD+gHV0vD+DMTNUcgZV+zxAxn/ZzjIIQBwsLSDKR4zVjDOSK84mDGr577TpKb+
Z/QnB8XMV0OKDtyXW+YqUbqc9vRGWPxDR0EckKPzz79ge6+8uTsmd2CfPlFJCoQNZ28hE6Wqj5V6
Z+L3qjG1t+fsFM6Y+NFn0GtgJy4QPnpT/W4IuX+8nqzCe63laxtFmIG8PW9HOIZel1/Deivae7Zh
F/TujJpPjImkveD3Osk9k30p7pQocMXfSKerDOYKWKS9wZvwYGdy5Jq8RfStNcRon3POTlmpT4CA
QN0Y9M8rXBRKxpX2PEBFXO2RePCC/O5GvxsHHpWeeL/J7gh4lO2giOfi77r9YLTIxvHhcfk1VhaI
6NFouxW1SiW+dUxgRFBxBSu0YLz9lGJ6O1Dc922G9USEiGBFEJbarqhNlxoHorm7gNsOXoz4l1ZS
oPySWVFge7F/QRatHV9DVXcjIgvrmDk/cMmZ/o44nKE/DSA9nhcVW/8EeiPDdFpVVifDf5944z1V
WzBH1Bj8myvB7pzQlTVq7TGlTotyWu5Bnaz8iBf8Ye8t1wMsL1WcDDvEdKJkOXR/E6RlXRJ0YDg1
/uRnyTvUw6xgs7j2DW1haJb8ySzbNy9VAS3YFFcY7UJ9NRpMWpQyTww7XxxCk8DYLzNLRwGtuB5z
PJhRdh9iJy6o63oA3s0VIVjkvS0YbKnjMS0z2GqNR+xGgAnuN7gSJ9mbEgqCo6K7QIxagy4/tB9H
XndkKnAqlMBj7pLgohBREATLx/m6alN14oTwfSXf+rhtE1q7rwsxMUrKk1b0JdtRZ59G+zmaaXiI
UI24pe78sf2RTWEZq8MXtHB7ux3Of4kTvJ02l2xm1IFztd2bKzZ43SSLD/SNHxH668jaD3mgq1dZ
51ed1PT5J4waEum1CASuTSW29uWHrE+5NsV/wAonFRj10rMZhBDaInm7Xitd6hlpw+Z5JKv8T79m
ShZ7m7gk7U7mPMbPovb6e4OH20cgl1tnyMHPy6giNCV7vk3xgPmSH+heCtdHgQFKf6FmHC8M9bB7
daFncWf6/j55i/BSPxjs66/CAxCjWfVejqidLcCdpcZ+Vsu2repuDWNXledbw9GNluMBP2xZbXUs
1Whh8LWPmXJkQ1e9ZHiPdI7OH/xeg0f/6tMTKR9BNCPxSMXgluYJ77YFb/e8eIbkfsI7QYMNF5Ux
3w3kxNN5lzjrWORuZ+WzqhibsGpUGymv84Dy68ydVpJLi4YQbo9rQfR40YhsumV/XRjkjo/pD8oF
qtttYxVwBrZGK4IjtjvjHb2bLWKSx1VxhgOF9uwbYLESiXAnJ+wQNwOzRiOpM18STsoB/mkVrBfA
/c0yMpP4vfTEwtWilG2dAsdJlFlFiWCeaxVPsBkHfT1zNtuJjtvAI3fIS9sR2pq+5tDAAnM+cdVr
xTDBjFc2VdhtFuT9KW9Z/25nEHblh1gOBqntBC7rsyMHfCaff4SldHNESoJCEAS9KxULnOvlyuIV
ZkU0iBWSFuMz5MxppZc0QwhqaOH2H3TyLMRN6rpXJ6xuVfKl9RlUKmJfcZau8hphEiYXtnqQKHAa
IjPdkk9kT7UxGbZqd0IcdFgkwD1eVA8CFAKrNS8ckTmsQ6/SQnrJ6YOWcnXEDE/BrKlpf+2/A/A4
fmNW7sVVUCfPVC/CuwSzRQX9Zs5OcGOg/CV70OaCW5t1nBMo7nCORN5eROiRpdxsnuayWLcDC9+k
JLWKrJ7qoOX9wDbeyugXksR6HY/KH8i/LrMkMaVwUMfpqsw65gLY1NYFQKkE5KBWC2QhT1WQRZys
cr3MKSKxUp+bff6jLUgN19mUOpyDtDIN3bFpq05rlqWOsNPjsRrDpOpK7tuDEGo6ZUj+RJgHiwCw
T7aKSRlUOnvvp+YAiO1dBjLbcD0qiUKOstW7QOGtFeiRm8Wh2LdsfajuQCI0rwwh9OeluC8rpnQU
9P82bqjcVg4Rd4YmYZxLtvP1nLfaK8CM0BS6wywd5wE7jH/pMQlophwiYWTiLqvsRg60gV1GA2VF
rvJa6mpuCg/9pEysrk5bz/pTnVONum6Gm8IIAmHwMTfTlboo3s2W9fJGlS+CG+RWaBsfbhBNe6P6
H/4gUVF05CenwMhYTQRGYgZwjx+le7wbQAsdxDrtWeEDwb2LWWX1FxHUhmE3JolOFdvt3JM5SbqW
/cZNX4SAOBwawX/zeLKSpnh1sWTzrCfDzL7Vv4dJ+5vLwVFC/X1UZNT3CgazU2+JpjS9GLrYRBdH
CbYPFtPumNzBgpw/xE1fgVcOihOwSOs/factt4dKoyBpqh6Qdyvv8mwZ9YGSvIGZ1Q/eX2Z38iNV
kDMMNOpB8hJI6GZgmEHCP6DQloyfcIlJD6tgbwlAdSvzs/jYfH/2c0/SqoKNwp88AhinjleNBHxo
K5bGq+D28tkEJ390xwBEsH9srr0kVufoTtnsvklRmUS0/FcsWKE2yqkDJeV1ttF7YkUuD7FcxISL
fgA1Wvu1W2w648h312+CmqfLoqrcYbwsMP1aAXk2hDCIFg7rWqSkAcS1dubRYL+DWD1CsH7ySszW
naDylpDzu/sd45lZp/rkXsjX36UpAQjVzC527/63L9UeCRmFmK63X0QqPDRcEpQBYR8ZC+MSy2kd
+JFfub8bcCN6anIDc9fhe2vNNRlxtZ+hoDwQcnyu13ZpUDoOOET3d+2zuNAG4UqHYqkfd42X0/ZQ
CxqRT+VBuezzAg1WhJA5dnOtJ/d5/8TkiNeearaB6Quq3BVGkq86Su/o9tstO38yi+rf2sryw2ff
lJB1gnNLWQUMd/Vd26swzNAhzbRIYBA2g8RR9x9Bo4HNokDnVjEixB/m6PplKj2occ51lYZ0v0aK
aX3kNGQPZR7AvZLgTI0rsV1KXsDq8O6A1p+jbkYueIOPMh2+XmKc3Bh54nYf1uJuOcHeVoscwzji
xb7Je5y8fyD3tz1TE4Madnl7NNFMhgFWniTjojEZY4fHrngZ40bshCVBhiNldgNs5kukQL4qdbB7
GzsJ2joCgIJ7vNKa7hUNbENqvLdka8jCNk0HZuVEDT6DfL7hVxPsKc5rNai2OScxM09NCed149VJ
RFlJpsnriIeLUo2R5sDRMl1me2Xf5Sp9KYIW0uc8Y3hyq0xv4ZFWyzROV40rPZSFquOCFKm9xmrZ
x2r1V8E/e8PexMu0L+XaW6NMxpt4nxXPHpJbSttXiD46KwzwGTOF9uEKL+ObhiLTRS5jaj1itO0P
U7KM1u1tEs8mfPuqtzgTcNU0hkKuUnKtlh3GMvIZ1NEqUgNo2gc6M1PdIIU9BduCUQxJO2wfckjx
V6D7/xSV21DMt8J68jnFdl7hUN4iAlQ7uOTkLMY9/tElMWciQwWRHxjS0oAxJFgTvYEX1/YX7HIL
ZiTPhF0V41S0NflUl++3Dki/6r3ZA43UcMG5I85zpVK8Wdq5HwMgcOrMiZpVwjOvarfuuhCPTXPn
BToq/9LsATsqdiymx6R9SHtGu9UNHDIRAd8aNXx5b3JYNK3+tkYSJk7lvTBU5WP2uR4l2TJT1w5j
GYf8HmBR806Q90fcgeYxJKMGxwqzhR+sg2vep737cna90jPBxZ8EJR9cmraAyBfyHr7gXZrLwEWx
bIs2aqYZrxKk07wtPY+KzrehvX2kEJWL+Gb+A8IPp6qoIte9R62gHfZOt9BtTNoP+h3Z2Ic0L/M0
tePXcFQODC/8eh+iOzpDXQj5G1nB7bB0FWQWFE9+Zeck/6E6eBcs+daSZwWNS0LviE+Vob8VjGoS
1jwqyr5PS6uTGl4zxD7G04dkT3Vozm50yh9WR4zdciZzk72b4bOnaq3I+YPOxk4b8PYg0QzoXAq/
Ak0yD8MC1if+oKgjt/291rZe45Kjiy5QxglLmjkwuDLD1H8avHffhSLQfM9ruS1azv4r1IV1NHdv
BxU3dWeda1klfMpuO0CSz7GE1uQ30RKA1JzuoKjZpZyRvHce2B9eas6sxe8sX6Wpm2sJzs9u+fao
N4YdmZ6YHP5BMY9EoaXZ0nucIHBkUfDupZBpBfpKdAuCJtva1eqRv1YU6++/g1SnthS5YbUAwAzH
GgAvPdaVz8dp14gCHgb0x5H70CbQmjzpX7e5Dxgc/gcichNZRiOcvwwYU1Ejpm7fe1e6v30//GAh
tzrTWK2XsWGNnc+wrqeoS2pjZKw5POZtoTjrGwRnypAE5xY4O9ZM9q20a75tQ13GRtFIhr2KUT9u
6t8EHqky6STz8x+rL9I7C1wfIMy1IEKF6M3Scgk2XHfTBdsr6xekjrzMKd9YHLNZUHdVKVIBQ1RN
pFjRQYQIMtOxQH1r1qdioy6LyhgYoAVE8/oytSCuOUb0fzCpyfqOa9BHzb7uT2FFRsjBu6z9UvVD
FKb8uhDUs9TJ+xlR5WZy9wcWs72vjT8M8UpOcDebV5YN6WpoHrtzjGMLDAoUZHVdg6Q7IVi64Mg8
06trngUMvMyB6NFit1ZuAo1dcWJiOiO9GAVd2SRrqO9POAfM9X5zWRZKF1flRaybGwbqQi7PrZvg
CVUGZseCNQF/9yyYVmNT75QiXjx727qg0l+3QiPHYbHlKFIHZYo3lucuA1p3UEN6vPTlR5pZuewy
I1PAh6S5C//vBFO69mq9EUjHCffbzKxkFhxJ2lmbS9K/eZbkh4Lg6XO5PHMwJiyjny+H9asTUnFJ
0VM23GSd4FSQNr22yFjvy4NMUHI/eQlmU1iqrKlEltbGHMHxQP8/IO/jinR6YVj9Vuy6mqpxu3LC
hvvgpveKYkn3AQ/cbnPZTCBItQtffQKjVSfSf8UeaoApWCCmYxD62FfNTC1xmIYfOl/7xxahjg/i
mJAZu9OYuK3SP40sCazFjoLstUf6X7Bb5Lbw01uloZmblV8QRElf1eYCWZqZ70C2Jh/xN/75XWoT
2fY6gvUCUgMI3LvfBPoXxW1VZM8WmGmGIDIohfadvhZ4LeTcJqzQfXEo1qkbplq04PYZWL9UpqWF
9rZEcCN7QcQUQmJYnJS7DfXUmqGddo4E0KFkVmvdQRvEu8Bzjkxa668xEP/3bFkc/mWA6nGENm1c
r/8sLE9iPWk2TkCv/GU7GP7p9fTilEn7LPdzFfxw/fNYI0caH/LrGLajH0ybc+BnHWC6KxfSOUqM
z8fa00Id4zbgb+3nc3dh71YkWORU74xSU+cXmhQYDWtif5S81p1VbCDVl8v9UlzgNaJgCUnMt1/5
uoNl5Ag5TfVk5o5YbU+m24I1HqGVJ6h/0hbNtHp265Q7bDNGNnCFKv6gGrW1qMi1igf4uncU0Oi1
RnrtJ/woz+cSN2YKWzPfaJbn8aqhLSsXgIRJ0E+6et1zBx/M4gZWGYhqpe7qQEjJy8md7MNztt0M
3YQKnM1fqicAhZx6WnKNHSDRPZp5+CNuDYO57yHXHCS6lopLFayeHhKeeXmzEVT4d7mO17wviY6e
YodK/japgLCW/hAhVLQVas32bcF9oSfG2aHBP8RyVeG4AtvJUrpNXsQy9pttNQbRvUemtN3opFM9
eUUrAl+QDJ2AzG2x4z+2+3Kl7L1iskNksVYUPl2Tgaav3n4WpNPil9jNUTums8BINVTSpl6XDKWX
3sNavDusJmSCyI8nE7kTBNFXF1ITx/KLAl1xCw8phZhUV0xgLLn7i2k+OBCjmtS8VHQTKagNvDVs
tfzjQjoCRpzQ0ZyXGApFc0W3Tko694qAxsug+59vG3hSzEpe3AsEwov6+7wu/qjkBZ8tAnlFfajj
qrd0ADj2uyn5QGw1vOf4g7Dldql7rgP1xMOfkigncETikOJ0KguOeFa034YcUafDM9NBQEm1FNhQ
h0FrQ2Qbho8ECMcNJxkA7XsKCRxjTQ3ijMDzQkvWNCYQd/5eXmnFzlECXgIbWJ4zBhmSm0BxZ2RV
58c/OV26nerbZ3Rhc7ckz5QcYkRcHwoSazGCk/W+RDazrk4vmYbIDSY01R3tPnplj58sIaUHRZgO
YJX3DJ/ucZ6IQ2nZyqrSDR9sY+ySueXFgtn+gPkRTuQp/ibeX6yFmg4evyOkJ2wsuyALRTQPMtNT
QZ9q2yJWKa5Qo7juXAH7OqWOMazKssRaVWT0CZtQQJVNnz4Vh/H5T5qgISQWgy2nrZuMXTdvqRWr
Tei5Z2SLm56cmSQ+zBgBdtty/RwHAJam4bLRUuDi766ikq1EPjXtpIdOJI4jpGIn/7VnJvUBeJ6p
miJPhTLTLUyez1/o/lumGgAhP2PPH1l/37ZxxgaJ08Y8azZ4+tpz5u8zpq/LsfdBNFE0Zp2QPZP8
87Ky2/0IVkGZncMQ8/hpEvCh6XOeTAl56yKV4uS01hW7Ed0jy6TQW4Q/oeBOXXnUGIA8DI4atU1c
xSiYepLXPIQVIhibGpBhKwjKjEbKfeKFUAnUU8PnQ7FGU3msAZjHtbCpKjGXkUU0P0pkANYHmnEt
L8BaQRXESPrZnuC26Kn4pEs+aOD4Nzds8+xZHRr9og2rBY1xUB6aYaarsqAD0G0zpqDdw8c25Rwy
b0fSg0Yox799350tjDVC/nfaV8MgIxQ3l3HNrZsjhKgyZdo9Px+dlws5Ey/xjiJbcF3Soo5TGrI8
dCApcOJ8XDAA/S627enlc7BiMBBIhOcRvx9oqQCeFPIwAalCNWcnkpKA0yrFwivINcBIoc1nSCbN
DZtXCk99D2nX7bLFdyjlIiZSBhv9LQ5DpdSi9G5c14euWdwzCCSeKXqZnms9Bf8RmqZDq//za6Jg
YSEf2wam4wWF97G+ux+zoMMDHv8iNgciL7kL9fLmn4NcK6vj5K5P0rWOb8RO/I+o6fIzYCPp3wFS
gsx5N/SFLLLjw+zDnhCbRvH9B0RK7uzl4ge3E2DzNcf+w+hPNrZrSjC6usQE6hkoP5cgexlK1rbc
xSGAuZ+GV2SGm829mep7z0/KbiPDRBTU7Lef++M3WorHMf9lY0T3TCwH6QdHyW20nRk2YxoszBox
uS4ssdLS/NUDVwUOhrl0DrquSVabKaWkgMHDGh1meBlNyQUrBMo38/ecbh5yC4ccAaelHGXtdAaY
ZtaUJ8rS4wiZxOibCnLjA+3XThCtuqDX5OrbEVYEVngDi7lQfNngtfu8+XxfMs7/s5FPSdFTsQiM
/Iv0eeozr2rkC6dDyQt+qpX34I8dmqtPvtowuGhU8D4d2XUTYCC5jq7A35uzpA4xmKzSdaXk5wns
iHxr/256qc7MxmUlUSXoQuPPe7G/6fht+eBumeDbyGtJR0QvKwnY04awK43X/jvKBj/nky6c+1OW
XxvYv34KzdpqE0gDKfO5wJbBXf4mAkwcWdRe/9jxPlDscKTDzY0QS5V7XKFUf5xCeVS0c3KUjNAT
mfxrxxG+2xfTZr/oRmqFE22POdQqwdM/iH2RmuEYjTjnXEJes+niopbbxWBof5lYflBkjVj/je1I
WK1dnZuiDkEL3VzE/KvnGSWIoN2WOW6v+U/HgNXYesGQupTnGX4d7PBMUYlfOguNiC2Vl/dVOJSE
3xWesMAxC3gvvUU/QblLZPS8ENcCJ/cVS3Hp/1En3DwJQuxBAQzBXAT49mcS1NIVQmKqY9KePtN8
HEwg/xBlFplptyqgvlCPji7N2V9ax5T4xOSAHiDbq5S/XNlD1mMmhfIft9z2k/yvhV8DvB9pNDIV
jld1DTVbWHvSlLftiogrlYx4Wj0h5cK/pfnlnh8CE5d6R1s2vN1lVEvURh/4z3f4zmJcIlDUB562
GaA4XpOQkA7LQ7d3JOkBTtajhrkJ4fo+dNlAj0nThyb9raglwag0cNjjO4b5/0eChEyB3vO6jroK
FtoCLruP/3K6iTgno0vdOs2cWopJUDettBMsO/wDmgtF4W207t9hoVcNF+vemFZHIHd28c8K1c+/
lUREN3hNBw0MFyO5QxPYS4qJfXJtwPs7gufPlJJIJgY0tQjYXL13fiPzooWO8/yogq/koLDlSrqa
uOg1BZsq4EX2NzMYqpU8Nceju9oOdGTxeURYNJ50x5EH+DB7jJNPyvNCiJSP+uv8c7JV0fcpTt94
AuVFxj96V1GowCE7RVCL7dxEMKFb2CpEVf3EgddSXbFmL1zP6wOo8+hkB2MefY1+yKnuFgGLwA8l
QLZbYgqx9Bln33/niArJzURgeiV3WFnsQOq4ORgxE0VnW+TPhECgNhtZcuqSKHZnN0OaFu4SclW8
aBGKi5uxTRU3A8VGCpRUUkiamxWWtMMB7lnUwm04EtS+PB0UK9CylnVagsi5jzqnktzZEfdm6rXr
kO5IYB9DUNWdEyNbhV8Skir2x1XqxrRCBYgNlNjfwfBmOVXgc7sHuSPFOg5rqyygPg3cL+k4jCbd
i3dR3rJQdlg/lEzcyddtrEKDvXDMVeZob35lzh92ah6UdB7IqAl1amHJU7re9ly4BPN3wrd7YgxU
rNV30AykPJv8hh5kIIuIcYWCWxn1cUOroepZFXdXUt5ispu3nYJQzB4Fywu2ovensu1uL9/J+TJ0
JaDcOrKLFY5f4HhrTqy/soMVTSvQ4o2JWa836crDsyhA4s86bu1bksSJCS62s5gHRzFAN62aKj96
zWYqlfrTdMaWMYC/ckG7lLszxwvYayDxSYK3L5LSnbEaPKaZpAfC0IXOpWBlxq9bZ1HpsMqWuKvG
lB+KhQu8CoAchMGc3kegzqhNLGrARsICJx+WeK29achOTPD4s52NER9q05woC1b15yQebIgKB2+4
5GSmfJLMso7oCuTX4zxbv22oU4c6HEBbMWv+8DjCf/ERNSELzwQSrexoexYGajRF+i4LTEJZstAP
26UPK3I3FU/+P2+dyFOJFJUmFx1tC/dQ8BIZzE2zGlWKOKehPDqioGCEV7OKHZSjeUxvDzHZDKta
XCMGLGfo508tbaEyHxjz9yJQccSocdPgeD2AZaQCdqSlo+o3xanZFZZ1FqcGbnyULEUYHIb9l+/i
4K330t2aWdR+vsrOJzbiEPV/4qpmsWCL/9SU2qTk0u1XXtwWtuDYttpjGGP9yyjI5IiZvZYeG5nR
ZtVJKyc/SD7QMc4aTjOx/oXlEBtEZBqPDThe4puKFlUHDQ8X2n9N4pW472Y8OZkvHWHFioEQ03wC
4g2FViGx1FXOJrfZE0ARK9skdS1wAKFZPeE44c9/eIBTD4Vunyo9WQbJ/qQ0oOglwqHqhRYKQJ0H
0tYRLlvfhnhdlkqmVBIPnIuYwWTKxp/ncnlPPV3KKVkI9oAAokvLLqVJVSHoKp1Rh69ELK2UkwQv
6xzK2P1Ku2DGnVCegNXILF/dEToHPOFfm17q0NMlLSJ2X9S5WFbxhm/66BedIspjN6kq+wbnSPEq
5P+GibWFaKVHbaqYMebeuo2IsW/na/ouyORhDxhybixUgt4G321A6caOeAqsy5Oh3SaXQs9vwbHM
hdPVClvt5CPwlTdoSnezkNuPSLZypS8e3mV/KoqAGAW5clLd//aKLTn4qFY4vGTNgbGhJM/TDi89
aF/4Dz5dhu02EXqJBKTUPVY6ToBtH6gwaTXIBBnlfN9wum9hYLOkB3BzYU9EKcfrxD0bVB5gw0qD
c/HkNZo14Jf4bJdiJRGYJXSDn5ujWIkWS/Pu1eNh8zP0HfaTp2vtGsdIrb7+T9rE6rrWD3Nc+xLc
sjIjTN28h3LmfdcC1k1QMnYly+J13YPrcBTqtpx4Efu3E5OnJjrjqxHQeizh9HaUViIoGL8sJ9z4
cr+seJJs6GMTXvLunh7FYp4c0IaQDrXDZO6P5/3c16JR1N3fmWRqEI6fLh7Z8MAL1lXxoGwdZBYF
wTHNoxL83wwFn15aLHfR4E+OhOS3xvP+ORsQ9krs2AA3lqOBduVyiQ8jG/sF+Ki4emOXS65TXiH3
JqWdFVow2XMJrigQqN1AOEqlJN08no7hM0xnoOruTHrTvoH/R1VOdWjSK0Cg/3hXvxDpJeot04Fv
GZ/G5pSwUnjZlIlI73ipWIjnWZCoTM7C9Q0ROh3eJsmQa1d7Zp9eEdQ4RbcaRnD6WTka/oNCQHEH
OXc54F/j3cMecldK/s7PmAgusOhqnae6X/eC1vvrZPYUgNH8+JS2qYxCLB71XV2aHpQscJEPY6bo
hVZ3gNYcBQQZzsg7g1/qKSNlNu6VvC25xl5al3O6IWs+S3Q92swfrXbGTIaQOHRdttbRBSpdptSL
nWMRCFghm5pwQUrWtRkonTUL+k0COJjZqOsa/JhgmrkrZ5F7p5GrZXw9X91HTxI9zYa5rBYM04b0
5SmNjEG4ot9ysFU/Rw74TJm4ESrpEm9ViWsh637gGvf8NVhSpfmB2L+taU0LrYSN5Iw+rG/YD/z9
gkIRvGDGfFCAParqT2dkzJZFdu1nfSMbrvYvs+PrzTICxv/xYUtqgwdq1PWF8ZWE20ThCUmOfFHY
WWqqONLayxpasRpnQ3AMXLl+D7NvRSsL9e2AzGSecGdcvJ81IQZSvNId4gCmtpGwfoBdGwykMjMP
hhgdHf1E42nG+4qGhJ/KDKP62Pt9trLIaYAIJ42XyvuZlKRN+ohfbSD7w4sOHE5PuV3SW5JQorYq
KIaDYVTuAl5C4K4taG2cYDdH7nzEp2Fqu1gPMxUfHUdAA9rZR5dFzGku97PG/kAnWDPIzrSNTtnB
tcEibZPP2g3hKhjFpsIZzM/sOX143PkB7DTJ8ldnfE9c7ZX7n912rrSx1v00zhm0prc8ddS4+xy9
OfVypJ3m4GYvah/IWhSAGNl+eQB65JgKEL8NqXudh7bpUpwD2b4Z218qRf+U7Dpzc+yEVg79cWqu
1rc9BuUebwd907JG/rtX4TOpBpfTjpMNxLZV51BPDdtpanNeSU/BAXIOM0VYlVY0h/XJtpeVta9k
KnkmVQ/i+a6d/fFdEEIZXFlSI/RU8QCFfXvxKHrt0dxbNX4O4tECWlp7KEvriFjxZs+Z3sYuWyKJ
buJf8OCGCP5KHiaQis3bHg8cgmef/LuThzNUqcwT/k4X12ZNBr+/RNfFDr2W1ZW0VU//lmfPi5Y5
vGQP+bVu4mD1i5ORQ8QDECBNojWMXwGmXAINYYm3pixj/ItQCFgxfWSgLr5p8t1YvNJVPdGMrDrO
JiwoRBNJ2PjqNnGxuOCVBmxeQm6UNwNtf0OEfuCJuCvMgrtScqVnlPPBkppYMIaNwxgfIbM31yMb
O1C+/8bO5A4rRWQ4G9s3a/T6+A3oaoUVU7LVTF9pSVOq7EDeN23jAdkuio145DKkIHnKrOrX+88M
SjQkz22ui+9kbT31guX22wKEZHvF5M1EyC82csZFIVf3iTB2FJqeNv5jJkmuPPWOt1W8eq6hUXPu
QhZ+Mbezip291rv/MUoO0KHCd24ia0qpa7wOmtaA6oZjOy4h6ld7GVMaebDJU0Vpl5mGKsqizzDw
+UfpjTsTh7V9aILz5PnbNis6LN+4t7GL8ACTm7zOkP14VViQvCfYnw+uDmTaDeeJ7qdvhGSbegvM
q0x7Yx+gz5t4fm8CYwU8yXKpyXI78rQRJCMkppVgUMYbrxGG7LsbjdoK9FYS9QiFQUfE6i3jfNcJ
BWKMoiRK1UzjjKUf5G9MP5M7TQ/o7dPiuwyBTyLryYCTGSAm7EEzwBAt6By1V0ypP4ENrLweT+DO
/sK5MsLeHvaBlu+lt48dNo6f2z5/ZVEminrJCN2JUYFSko53IFS0fe/VTtYiNOGltAulvf34LDYu
DeR3BOFbnupes5aNofcPAYAZ7WF6b6g74kbLe9kqVswZYliHKN82+EKsUZqiO3SXh6+ZBC3qiayA
cp3lxIzaE5Ig9Ri0qb5issUJd8lKeelaevP78gys1Mq5zeDuDY3XMDaRUDNltSXD5siTlX2sNWto
26x0llmbgmOH3/Ohwtbe01cz51IOAp9ZSj4wcxXT503FQHOROj+mtmKa3C5rHG/IvgEEOSVFroET
GysdA6lPBI4328vIP2N/RP0zzMXzLwK5gUv/QzSrCeKSLEKnkjhDHwTggOwtSgj555wZn3vLkHjA
+bpjEX4+zoelVw36OfRDHZvufl9yhx/N64pBG08RbFWajPqGY4KnOZpGNNL2u8boLCF6dcVMdDQF
JADTH1MOVeVS62K/hHhVgDcMKSG6DOZRv8z4Iw3F7vXkES70KzMTfV9YJpg8CCfP4Xz/j6cKvWQi
oYG23KqVLt6cZaoJDJnMELr+5Jmf20IxV7js9tDKqWaGtIZXBXJzzb8XyLeDyv9N/r5HIFpfP+6K
TdSTCZ473XGsmK535MUlBAGyZ+GFbLl3sqcn7CE9U4rfjcY9M7bS8kADDA9UcVRKY5ep36crZVHi
tbY97Eh4in7BlXtCcO2+u+qZNqCIX2/05KJ4jjLtlvyZqvJFouR1y9L9qwWucHJbK1Nl+ujQyEbk
M/vJWyUpvSn7A1P3IDGsOk0zc8/m04Lq0SyjK37WfThmmdz46unZy26AUEpZeBE6UCLEVQrbedJb
UeLHYBgwDquSajGgjvNLi7fc5QFWIWJe+WPEcBHxBu7tdvkYDCLKjuTp7Pi3+wmjSRiVIz7pjz0z
49LnvZoS0tiutLp6rrjZ7SSXzaGH6HaMo8lkEudWEeIdPnUnT9ypHaRYRj3TwuaqziZjaLmpBg57
5VJLeywo3rGAfKSPQIfKN9BU4ZEe6ePdg+1kglC1wIkemtrm/QS5bbNJFIipwC8M2ezpOPbrpbDh
KckzPNeId8nmfD6bfZlEZpfq0Iz9cqK5P3hA3/V1o4vOHNOIAOVHiJci/xfBRYvrDz0sKtEljnoy
hfqhaSRHhSBCWZ9kIgfFHIN00MzM5seuBCqXQiySq9Rn57mxN5Cdp9ce5xoH4z4dM/4iuobJXi+B
OFcNwGR19VrAX9V8ZgAcyWgI+vvM2ASK7h60fO3AWMKtljzNX/2Ure+csuI0ZpQXtFd4/GNn5sdm
YzIQP0w3x89FE9jVsOICldUavRQ9Y4goMsdoi5ad9VxKmid9Gy52gY4CCJgSKH0Z2UawqNzAJpL3
8sr5jVXe6Zk1qyzTc44/H7IVJ3I7Ugze7FxG79FjrvWn80bcaiXE5vDu9ZWcjSiD+vx3ehVZUbRv
e8Ce4xPlaNygQ9KZ4sZ0BNq7/0pMvmJV8SDtz4R95i0d0xaZRgjWbd+Q+aUM+EiGqiDBjLntKIbC
fp+3Qf5uhDbpmB/x7lhayTWsexOigwVklInfXqeWvVJpaAxrvbuYICzzAjSB/mCJJHiJU11a7H7U
PqKxTVQXoU5uDqDcf5KYg08TfVfOeb4LW4pGLTAX/l4Flj17eci34YRmw7d2cvpQt/aq0jLZGl6K
+SrSqjDlAwTBODlo9vLivIB/xfLA3o4wg7KkVG6W/l48Ybsa5rtF2zcYlkPSA57vfoly+vlxGxPl
xA7CYW5EEa2nsqtSTmpL5cvL1QgfZaOQNZn6H+4rnX4+//9K3/FPfP06o7cVmDtQHJfnqspX/G86
YuL+x03HvFd20Nd+YzzMDm+1bnr7tDdsWCyyF1EgLjr+lN7WFG5aj4v6HQy8it7g6HkSdK1Gajjc
yxg4QqJ0w3hTKXX+FqcN99VzfaKiDjEK5a3xLiq1a2nb/oAUEqBpZsNySL8N1uqEiZNncbsFzhkQ
vfk+i/2cCB7B6eOW5F6bFuef6VfIwDojUvJQpdEO5GaCTGVN7uHoB8teejnbOhABeha6aaag70c2
0g6dYJlLZbdii9vDsv1B1xm01cDn2bg3keZGHwry/bZ0AR26n8P7dwWmcyU9nDeP+mnZl48ItQgC
HMJmytL69JBeD4+50d18uD5SGVo2wEtUjCrZwNKSqm3SCmWJjvXb5QrgD+LaaV6jNivIshYtMm81
NYDRXm9sf+Wg/kJ2J/LdVW71NR9zXXXyfGN37MC29ypmA5uk4E/ueL2Kn0+Hh48r1NwZ1seE5f4V
cnt1IFos6NxLacIGyS9zA2laZQkkvtNKeLrLxU52UT9xvDxT3V4iQ9Nb67SCJ6tHe0ZMO6zicAkh
HTtJjoPyvCCoGQfKvXJjrY29wVfZEV+UCDE5w0sRncLplKkCSs+wj8VA45pYMjj3rpN9Px5qtaGM
pydxP0SXVwcgnHzNW+tmWwlgJU2Ex3xRiavnaO2ttil7IsOSuvIm/PfghfO+fZvTBwcpHazJ5SN+
bN2/o55987paxfIvhOx5imn6b53jpmjbmb7yxqkifkkqNxFKsh5egaMCD80uYJla//xTs+QbM9/a
M167kLgoZspUXpegGKo1EUEBthqQWrhoEjxUVPIE8aFMUQPJeS09hsuxCBvLAGsmJNl59+6rcx2n
5IOf/mcVuiZWpaCrTsIeuDf1Sjmv0XlvQAS45BMSm9JRFX6KSkRdEIm6ZI+kcOhDEXfveWsLuV7T
ZZ75i1nTXJL4ZyhAWHp1SWI+fgnbVIC5gDcWIqW9Mf+WzSoecw/OD0haM2b3oiRUzRxG+6+Gfm9U
1WzpUMx2Ox92jIzZmY6niiugERQRoiQLsvUFURAsHMg1DznN1Jjn30QYMH8z8B86nTT/Ok1bpLjX
SimKAfuB4GrA5ZBQzh5gm9Z5fUDLZyGC7jH3TCjV9VUjWFcGm1ATOfbcniVdGjYTRfUq0Fc5ojPr
S20zHlK2Wi0l2LskIU3BUnqA/IQZdUhh9lnDyvou6XwCiaCZ9H1W3Q1y0RAyrtWLG5JY4WPVjQaO
swFPIRbdwcMV8xQcF02twV+9FrhIsOKVqUxFqgj14b7AQgplU8vEOC/dxbIxsbX0lLloy2Wmso7g
G93L67tIiyNuAEydSJqnfZjx7wFOJE2BRHjuTxPYCD2wSN83HMa73LSw98jVIq5KWjM6IIDWDHTQ
OyZHwQs8jsq5NBwTp9MEdobBeRJp8ED52nvc9BhSlDnZ7V6ahSDj44FIy/bgWh3mmRyT4BbmJjGx
pouo07hThUpXI8uIbzg5vjyRqNf8khiVU8Nrtd8ryfTTTlOPacdQbrSzn3nhcSifN0QDTRUQVPg2
EIHjQsqKW4l63GDt55H9G0nKPo6FwUayCZCxTV0IPUII/k+YJw3BdqZgOGWRn2Iyt6E4WHC8FyUr
7qQGOdSjKK0W0u9hGrhWCcjPZzgAdOWD+2iDEF9/EKgblyNM6M3yLlFv2ll0vW7tvVIJ54urP0pl
oIMpT6TxIwc0k41rEju2TfKSh8wDzjrthLpKPJdz7GVH/uEIIW6o72gCTWKF8NAV+ziia84EQlYl
Co2K/3Kg4bOG6Vg0sfPrQ/GQsub+UJqAxe3UOh8TR1c+yXOKwG5ga0Db5VOL1lZF0ubnfKXD6o9M
+v1mIOj6e/UDRpkhjxh5YAFxvwXx0ydEzCGiHLIDg4LD7YCAkTXOmr3AV0om2g0OjGK6Al2+Y9vH
391qGuixtCCp6CY+tmdk2pvmbSFsrbPo3gRxBRTfoKcXKWvSwsbS6eCiy2gbRb91faPwyhfJHN0j
vzeJUzlMqV037X+KbcTxAIuR6ekZSOxZWkGjtOjWV5m2W7ImVM+VHj/BtUjAncazCGOpYouCGXXK
9h2ykWkUhfw/9ocNQ1kxl2mW3DMqU9q6mFP/7PD8Vy4vi61IHPGh06fvlFDDTj/8PPBPsOBH5eFQ
JDEo0aN6ldIvtcJ3AtbTs24irI5TE0Ti8qBKYsvJZEC4LolhLNxjiugKwTd8SRSasJNQrbzEiY+v
bQyUfvB3byR8ZVLPs3xlOTTIIQn8qH6ocwrWXx6UrVbKxkfYyvtEqGICfzjZFvt6v/XIYwPQAmEo
URtuPdN30hksNpY1awKSAl0TDlVj0TyZSed54vaL5R0l4uiU9/jTLmxPUkdswIaJ52XfkQZSzRU+
/E81A4RO/isuLro4F+eGChTm+y7NpOcFok7j0SvxPxSttTZ1PMZ0DMR0QHtt8660+MLBHjVymNE1
scTGebTu+G0cZ2ufI6nlxHtvSec8cDxPKXXIxfwPy+t/7i3SbX+pMgv0FhcujIFDA6fLDEkoUf3C
RmU2laWzgKGx0nSksGUeGvo4YiSMMRkv+jv+McSny7FKeuJNq+GkYTp9pA7woSdk+Pslu7oEUVxS
GBz7P7Ej1IoAiORj8WP8hioqMBdq5FGpvuQiJhhgv9HK6rF9cyzV9HIWpu1ib5SrPwHHT3ZBFyI8
uj9lckZBqZBTYMGpoupnzpxdh16jfu6uCNHthrHgsj+MpMDBSu3Qcs4SqCPNC6O53BYw8+Dv0yFW
zoA+UQcYmk6meOEuftjPzPI8KI4y6hfVFYFQUTFaIcjB0lFN0CkeIwI7l0bM3TAIXwvJd5CZ1lPD
rzPenGAVvJm036nQg+iQQPRzsdwsbiMOj5NFyOGrKbwdTEkZMz5eB61fu3/JfJ/yR9OfVFbEdbOf
ywkVwI6Wx5DKxlYGtP5kItfwD+COHhhg0ng8hqRz+feW6iSQ+Pt1HxyhQ66HQTVTxtKtLzWRcpWi
UcwinZ1Zn4Q+WOmOYuv4bFXp4LxHfx8pwXbkuqO+nFEx02/Qbi0zMyCu4VHkMOZ+hFCbUz+NaUSM
YkLeKOV/4WE2xcWX3LjLf+YaGIsXn98aqBdmcHDFq9myJAHYlpJL8LOkHfPHI8k8X6+dP9HYXtu6
cXpghEdM/CAG70KEIIDup9d5xhgXYNCgl2EJtjtgfNFt4Csxk2ncmgkfhgDQT3QiF0S2IvSaU06F
i3MKp/r1txuYdacO1r80Mp3ycsvKNNItfjWZYjvbe2tcHhYHuEIjB/Z83XFF4VzfgK3ejsMlE733
Elc6sY6QtX9lxnQf3c/6M+e3sxDo9cigJAHWdsDcco9DdcHUaz0jPHMI4HK01+NNHw0hojeJIc7K
vl2BhBx7tLEf3FJFtGbIFajq+oYKwX9EyPRVSTkdsQgC2qfM5sSf/gmhOHZBcCO0jffzHiHCIu2J
kXsBKcxmMth7/axO2YMWx9Gff8SNNnee7ocsP+kCT8LwbZ0uc8rfHvp2AXorNFlGci7AO2oLDsqB
neyM9hI40go92qlQvtWwC/qgSDUjgqt+mshzNXSGVnM7zj3zZMyGwpERPxzOHRcvpH8he8k1rQmL
Cab2Qu2flNWNoEaLncExpxfFGJSQI5T/eRKMFwaaT/pWjgHL+QAeecuNdGoCBF3Nuk9H8nSfQN2H
HJBKoOdtjk2VLJyvCxLXCDQ4Xk1HrS6xRGNhe2XXcP2Ffuph+OLTZSjjoW2Uw0t46Ob3mrCOOgql
V57COyxu2B0uykORwVhALj+Vzzvzv/Kf8s+Y35ssV9Zt0fL5Cfeq0Mg+KIiEBbaL8ZswcWkRSumJ
KfErd++sKLZwhBaZeYsJEuYjdVsJmUFpPffXqPxrM/aHpCC2AaiG60rauCvW0BYyGUcMSR5v1ELR
tLJHgtQn3sqOF1ZzU6gWbou+uALPVCyrWoBLq5X+KSYPve9Fe8YyVc5ibNV+96s4o6VwNv/61EWX
MOJRo+f//Kj8fKQp+y1xQ/qxoopPxNdfeE06zeyuCFYw6npKHKMcjXL1dXUYR24zmjDT/NB8vni7
HcIebjp8eg7A5Zee4k6Lsq0qG0tsObLeyYRqYeq0xAkPJk1N3aVKdsZGTyWKXKKtQYdC9kak557a
jO0Ji3Riy/jufRvyAqW5b+ZxAuZdc4/UfvGWWehVZd9mmYd24iFyBoWkXG+cG2+b+MTJIa3UT3UU
7lT+6C8d+I74OrUT4JikZYoOl/N+Wrblmae1JLMxtNrg5GUUjvERONJjkJxcVghobSbmNNIHFNsu
YLjAFsNyN/N/A9NI7nQeqVcq7P3WSL3ZUKzXtX5ulyeuo3rfb2msLkre6IGWQER0XQp7vzFy04mM
AOhlf7cNpDJQrqpk1jjjXer7GBdZzyQ0z4U3AWsKC4a0T4/bZ66kW3n7vUlq0izVYoSifUouxt7w
TVosH/qHA61LLN4n60mNv890AHvKKvL7n99aLiLzhAec9Jay61FkVVjvlpXJIyyfl5CNN0fDlK5L
BGK8Baty5uLumR65wfddbkQrUdymPLNjhzpy8U3SA7bLm+kFgov4v/XfZ9O/hQgqeN5B1lXGNe4U
1YaYVIqN1tWgk9e5qa6sBvmuNL5XtkwlWeARtNWGmScMbOA1hoOfrBM5O+StpYkf1rPPedPaONKD
f6g7AjxS5OkJex1UHguI2yD38zLp3jzrbzYFekIkefkrwo1gqf+Ab2r361kCJ88y0nvnDXRCFqtm
Xd9+hQxGmzQdmmFAHbCpZhYHtZX7tFVLnTyzHoJVYEhaES6XsWC4fv4bRLLzg2dXZw4ZLX0cT9Yb
XoTROJ5SrsDdMEkVMYJNBBVTKEZKvz0LMMria3s9+FeiziOMznH/URsDELDr9+QjRRPKEi6JrKXo
76LP00675mEOReh2eJzC4srORUGmoRDyoWdfLG3gZjjy4/lJ9ZYanrkAsqFClkQS8mBZDTt+s7Zc
/8oqvytMHV5+walRh4OQ3dh+sMFpuLRHykMGvq/VAS0jx41LM4AQ9zdgmoduNQPeP8abYrK7ZQLd
vzI1dA1f5uiB6FgN66jUYPndpIUU8eV8Bx2imRjAR2XqVQHk/oHqINqcptOJHqSuUU69GnebqjcH
Jhszj+Ly0HLZQqPA312kvHVPlGh+DpeNnECRm6MOzfJEvkVSqtlLO2CGtSG2SmZ45j678byIdlea
I//DVtj9/hL4a1Khvwdjczp6HnmeC98NIkRIK7/nSzipKc7tqwLStfBS6RYfL//FmWrDC3M6zXye
L2aAhFpfkPV71ahOG9C48MUG3K6rIXkaO9Zc243WJJHlmvzqmf5WkFr1vU2FAMyDNNNbPm/mdq51
Y8hEt6XhQcDkx4svYp9CjIHTvMeuU50e8kuFPGGWf0M0SHWm54T9Jk9QxDMDlrIhlN1H81KBoXzs
wka/yoq6ic+TWjbBE8oxDb28F4a4S6gBQ0SjTVodxzf1liTPD2ox7CfatwdnHrN+OG0TN4J0NJ2A
UnFte3Iv2Fi1z95YmAr10S9leiyHBMsP44fqyk5flTm6a81fw6zXr9RRMs8Xjac2Q77RjZb3yA+m
ay/3vSAUhRdzFMEX3b3jk6qyUD+G+rDz1f4L8TD9P85LX5OIptRl4QCFZLU9cU2cHE+W5lx4b0uT
CENONNIEWu1KX8NTncoT12g3L4n9eexfbkzRwLEs+8SQFFcrqkJGp7EUuKLSr8LnkOZQcVqZOSlh
g7s3cK/mCq2u2EqtFakD2wT7IdvqcxFDrp0hBSzgnOYbUY4gXbqljEIakoozRNg9j+KRoAKm6cSb
N5C8ho6Yoe9HjmtSM5tassI5o0pOUZN4SacafkDlVx02Ueae7zrnfDbWd81S3LY6oFUJRRqizCks
CMJqPepTYTO40WHSG3itHimzUHRed4ZqweLUViKkqOhWrmye55zBW+4wetniMYLrpkQs3cQWJoj5
FWFlPm1ewNvXuMIv0mz3rkmtw20AUbC28q5mG9MnMLbDcxgx2GCvkcXyv0YWFLE8OiX40Y8xbk92
ouRLWWCwJUG75AfyxuEu64uIT8RV/9S/pU1TEklUhoVfH6rl9c4vYpq+NlCw2zG0LkGukLwWK21t
YeSLpCKSzBqvnAPPf3YJTepyG7G+OOEq+UcJZk6Y+S8sB/wgzBlKecc+jtXY+AtQ/r4qoV7phIQ8
Av96qYmiPycUCcaVPH4m4csvJzfMfsUPUFtHfNhHOkv9JWmXJ1JHblyQi1hazHVNbj0vVLQz+1UV
MFFq3e++KYXXzF6ePwEdzRPviR3SqV8fU6LG5+Y9k9DhiiMXxkhZS67TrdlGxMgLOKcDr7eal1Op
HcOV8IIum4+TddtG1UhZQKHFcAM0cARCSX/88FbZ6ikOebUOGg9qd5+lXRKZ2DdRd18y7fusKxA+
72Utq2hJu79THxE77VVnguvZZAF/ih69rV1MEuBeIlvNJHcoDXnPAMjkaLsZw5kwXN9CIFGH84cZ
tTrvuU+y3ef3EdPAdNnBfmpLsBqiQSE8xgxEbvtJl7dCyrZXbXjBUj9AjAkSsl0WSYlvOLqMBMpk
6Tb3KMUAn/J937cUdjbLnmGBROPtA3lTwUJHmWdM63PyNGpJb+5dZkaF879CcAzcte1PszY311C0
/DwShdc1Ok4RKLkzle7OlhkPIaA7CKQhtaoKHcrK6EOa1FfBj/EOWCUgIUoXCg13NBJqhcZ+F05I
O5lCbgI9jyy2KiB1bO+On0L71MHWvUaX2G2xk7Sy/hEgElk4rwudTKHE+Irzs+xarrlQEjBhhEo3
0MJyjGW/0tsz1wrMEbZBhbLNT/LNIAY3i+w5Ca29TKyhA+yVwXO7N8e/xU1Nms/TanT4VsDK1T+4
J5ySmEg46uNxIBuZ/2StSjtF/dPed4N0N3Bhsb12bfvrzUKQUvxg4HaXL4vOVq26ODw1HoesA9Zr
GuDKkGzeR0ZXzKXBkF8Uf1teFx36lwAZ6BD9GOW3PoVvj1CYgu4a+aUAdAkXUeqJ8hRaJiJ18KCZ
gdTSLGG5P2bLT2QH7yoENs6zBGIX0Cu8RODTfSWbnps+Wna9U6WPm26G5WmsxwLV0WVcm3SWwBoz
s9zfVc3XpbKdY9oxe404xZwkXIGCj2XE7v5fC4kx6+gYI7NaYWki4Weovnr7wkxQsv6Xv66+I2n9
I8CXJLe88bEUXCofETEGYQ37gnSRxtAjKGX/yvwPFp8LxZPDlCycw5pzENpZh9LaKQKuQI5/RY22
0xP5ToAD4qj+3Gaax1srGH5MPkLwzgIMGMn45IdqB+Bw51Zp9JHF2rQ6QhHb8HO7a1XLt8kmLGwD
Lm17HCQ1bq4INMGZq3nqidCT9epf1g9AzOMlDzN0sbt1LufpgRUD9Qhr4yoJAp2Rm+a2WZi2PB43
1jJM+oJoMbrTZ+yRyj/cAX1rce9Pdv2rWhQIey0Pv+U8W94N2Br49SVKLuQ9SJTQPKW32zeY1C4J
6BvY9kHwS5/qTpeLQAOu9jz9EEHWRhtYqown5WD6CpZF4usK8FOcfP0FO2VREt2GJ/rQaeaJP3Do
66t5eM1xmfmsxb3bNOEEUt2D8BQZG+5wejR1479TMOh3iFzW1Ds+3wkMadLcufJ2CVFN29Wdnj8I
HjUU9w/6z6AMHbfdlK6URNAx6Z9lJ8L3MuHjkatRuyqRoulSsJoy2opaeDlfIos34zFVTc3zgeAD
18iuwb/yOOOjNtWvfA3iNuOiXtlPHf+SRX9caI/3miVG/ci+SwZbKkWCtUxr388EuGjRRO2XwL4n
+PXw2G29M40N2spFK8JyYgJGJ0eN+c3uWML3KcFO1ASwZbwAuNqAnF1awqP35PDhDVR7bXXAlhe5
NSdGG8fLD9a6M7NtznQfi6myZLOLN2otKM4yY0htjQv53+ZO7MPMu+h+WoMtYFXqzvmjjTNETGJ+
MyRspWxsLA+FGYGGXyjiflhSuyisbWMNqVK4vVz2GMMFaoXA4FS4wgQY13xmMleL2dfkS5NokOyu
/Qzx5aUJLvvmI0hygUymaPoqkQ/74XEIlNik/Dw2N43DUIobgxUoYc8szBYdv3lYTdIJzfjy7oKn
+x9py6CVW+gxXIP53Sq2eIEfkvdpb2AdTv7HQaYrtfBpH+votZMPjdSHo0a7FSFw9zaae/4vSdep
AuSZeIl38Lhj+vZB4o/ts4y3GRiTvocCSQYtUPqCbguo1ubEUxorDntF9eiTSlcwFXepYU/Lj+tW
G1cKLaW+EjEMHgYRQihqkiygAF2joMZOa0pqVNkywooG9Oxu9HzocH+8xUmc33ESHgpJjFQakoqB
ODed1th9KThtvQu0VFvtL32W347kVmLMjKvjkZM+KU1Tvv2vxm43aXpLbt6s1mN4gQ+jjMlJVT6r
byQNktrArH/MpK9iZzN7N7gt1rxhDihLrlsSP2+ikuEJ7k8A93nm9pXCGb0+HEcPPrCiFE1GtcD6
YjFQ7upujKDDF9syqr83qN0o+5cSBGRSW6GX4JgH82yyKabnJuIlJ8H0YEzxAVUYxtkroqNUsGwl
lfcD4Go989t8STca3AKE8XJDE7sa3BaR1p8VbDQrYrf1whgQofbBMnHiZFIikYxP13z2awb2NCEl
uVBbLpnMtU8jdLVoVYKzacCbOmN4HrHLQgUbi+w1Dsh0RBSgdJZs5zfTftOIlTJEPwUfzsgh9bIY
KjQV+G3/BNxG0c3RAaCAWLLWD9p0hbK4gn5GMo4Jbiea/jn22xF8vARWcNZjpPy1wRoPap/ye0Qw
hv4iiByGYGDfouikax6uFbGvHm0xfFVkGoSQtD/oLi4enuY2TDV/nGMe+PTpnB8C/qSRg4b2/MDI
q9Kfv4BpOt87gy9BTiR+uvEYqjhT8fmbSwV54fuBZrXJszDxRWhsfs9la5sfpCz5d7PmzGX7al9A
B7vwUyi1Wap7jrTNSBdGjvdstCmrQYALse4lETCsMpnDBolC1d1oGrh/5os8n5zsVoMpGrf3qKtn
MLfGikRvL/RIE2/z49CjoZ04N/lOWEy/7U5T5hq9kRpGvDhoCJ5HFtMjtrgwf7cIlVlKKPqiRkk8
hTZ3wLaTfso2pRJhHxxyfc49wXyF2xbB4zDG6cHD3opSR1cewGH9i0uAQHpopG6s4dJeDuar3xVW
EzhVmQmTxFK9k0c6Qh+RCiKcxvZPI6CEzWqg2Tm8HhVfzjgzDA0aSUE46my3C5Q/2eo0kB8P4vCD
W9ffrGnqoXtazceB7bHaU3oxHPYWmilo3WHuKD7eAg0QXmmTOcMlw6Ip/7Tb2euydkdQSa8RrSxk
dSBSW33Cj7gx3kc0o2JcIaz/0kL1h7vtXn92802axiphP7jac63MKJf/PMEV86HlTluJePTTXH5K
xNjo0lrZUgJFpEzLXpC0EH0sWj4+V3Qek5ZNG1asdHu7w7i/poVfsFVpa4pVxvs1qOAZNqc0F6DM
2f6RSMEqKhfB8FW6VHu6tRyiA0QZ1O5zPTcJHuonlh3m+Po7JMgDePK9l2NF4O8oowzcHhKsllpm
D1Ard+uESIm33D5QJFIw+ljU6HvwvDh2HMSe7GGkSmEmXlGE5LEBPjdBXVvQKqgVX3+1ISGvPmT0
pJeiyMhNENuvEIKFBwqZVLZoHDKHFKPuO3GatwnkSOO4BJUXesqJzHCWuFSsq6nYxmQ7WfPXMZ6j
iJsJbtVGxL/yog9i20dDbWRMAnyddg+VIgajJBcWG7vUl2YL37r8bKAHqG/Sc5G1mG34GrzOP0ST
2pBS+UvoSMPHoS0CYpKwU4EE1E8KAcJGozCc2u2I+jg7y5tpedxlIUHtvoRF0uDjZan4Zei5e6pn
07LwzdClJorvfvl4rrRMlnzuwQxh9UrnAMAgB6fG4fsAa9a6oqqHkZPhxFxJs9HXBHHRLeplcATG
1Q3nJEa16jQvNPWIJV1OncuaLia40V9cwzbg1WX9jfnzmRKIFZs/RwDBZCXDg9ApI8P6uDVld1Bx
vaXl8ADQZWuyVsKwk/+zUqv9pl19uVTGs3yNjoNKtwsqC29GEoUqeoPu38SIEwz3N/9zILI1FjFX
yOvIEFmQyzKryG1Kzn4UusTpzP19H+CMuU4yah87cA7gzEDTI0D1na3SyAmzu8qQ4iC5APEtzs8F
JBfRscQaOKHhaBBigeZUWmXMeTpV30vNDtpYiOy4MIHbZnndLhslMQHiw9W8R1HZGJEBb3jGTLw/
Jq7kMeEY+L41Bo2UzULn55MJjQviG6daHbJIcDBfWmXi0dMJt34qbHQvjOMJElfjIY5xyI7pjRhT
g06EM6EUfPQGlwA4jUaktBQwAjOu7UKb80jmrqGO82CZfMo2xC7l9TzIICAeMp2RosTVYoU/M2fL
teZv1CnCf31hU/BhUTsEQFDLNZK4C0GaV3aCNZ0NAPK/63B7anKqhNwC6k8mEqOA/xEDQZqoreiT
OEoUFjsAJRJsXrePKrcdgCCQElIZK5LvepORisUby0y+2CTZU7HKpzwzlgFmQx15PSa7uFfdEEBv
qqc7q8C1PK+82w/HJ4Y7Sd+MlzNsRBV7oYwYBk+W4z4pe6lF3C7eWQVzLyrh3B1XYG6gitjlnwpg
XnY3CwnHbFqEKzs0H+05DIeftS0N1CXVx9W8KyBRJPUFk5VwK9nDAULmDFFrw5Ptmp4iNkWTOd+9
Evv50n9+kypYmfOhVn6usGuJJP65nnHwt9SVgjpL/vLrfzsz5Ti8eSa6NMq660MHzg8Yu803kUJ4
AJToCe48qz95dTNrjgwTgxqFzHLaG+tpkyBRDfSUJiP567XHQx+dVAby1Q7cO2v4Y9BWX/zUxW7x
/2QLc+H/ReFO7WjFJ5BhxLUuD9DicfMWdMA/iK1BP8hllYnf/TNEv+uO2u0xckGGZ86JZHaerDLo
x+ery9CrCdQnG8eXb30p3/Nlgo2y1GyRVgo+7/yfSPjvpCvlnzA3/dl4/Cjad8+pngZDkaGDwqQY
RUv3mA+Jfozi99M6siAiamACeWaa723rVEUDGhQd+nCvzrMgZfzwG+31xEcs0dZwJiW4glKYTGTS
mJTqRDH67uDNxgoBWLQ9kNss11j6SXzTpwF4lj//ZeqowsoMq938F4io8xPPpA4zlc/L39rk0E32
5z0lncgmang78i1TZW/Fk0wnhFx4eq1dt6MdE2uhLmVGmI3PQKxjyxJ9UvLQvEHOIs0i3nyPkrqa
v026QiNROQoWY2dwIcdUHx88TZN//r4mIIB2kcAFKQtDNrXNE3kVqbLpulbDTAN/IuhnKJb4okxv
YyS3UGq5/308mEcTWpSotpxM4nzVU2xArHGHu3u7QKu3FJWJmpZ6g4owmUyw3j1iu7dn9TdcU7j7
n5MjiGVAvD7rl+FEOK5CMCbdmHMs6kQnx4oJdg7OobSdt8kVRaT7TZ7Wz8xW91R6lMfcg7C0O65K
za0BYWY/4bpBdZQOgr+rZYdw38phTQ119n11AVFSemYNzcdSBPzon6ZYhTq0J2LMGkg02LCN0rKP
sncgCG7IHbVG1O/MvfUZXji7SvrPJ/WfP3+u5GtP1CJ8Q7jX5/Ut52L80iAO0z1/U/1LbB1TF4SC
IjKAyo6cHyzJsTTxS7LScUL5wLMNGMtnIVoLlPJ8LYW/LIVsb9ByTMhWx80s7zKXzs6WR/RgSSaP
jwpzBAGicCXCGrDJHU0U28iNd6UlKapk9WR2KvGcQrTK4QoIkzAVIBnRbMAdTZzfRrX500jcBnDR
nPBxmC0NCLpEi9hCyBBoFbRrn3qG7KfYP5J3qbuwt6ndtrHhqWwZs7zjk3+mUQefi/4ppX3aO6fp
Dd2CNH2EwjmrURkuQ+lOqQ5PNaI8FyftWSHYqX3TPKnk4AEn7lofqhOdCYKd3eKeO2fjGcNSbRov
Kb15mXZ/WN864Zq8Yn1PURfTuvojWmspbUsrkacrsauHsBRZaeJzd5Xdq0YUvkscTfxd9Da8v2Be
lndqUBvK9dv0JlAinNGphRr6gby9YSOKbkPcdErb/XmTPzN5JjjM/uO2VFQGH7+sZPjff9Xo/ofy
RJhs2I3CFrQuxDFELenklfLG13DvuVuPvmKqmd68glzCZ1/39Y/YsNIzqZCE6rBtlZhSGankHJ0G
rA9Kh2G57Apt8Hnz/8ftnFnON5sY5HgVBlkREXmC2iAVuyv5eYy/grS2rPgLXEvNUCXwmdDHeRRN
sbAYTJbt9aCIzeQja5SEAjx0Rs9QcVh00Fg4MtWNQbFhF/agvU5ZDv5bieGrO/1Ey6/KtafDvIlU
KtdNXrP+UFrSQRzVTTpohVPQJiiYzhGGUTNwC4/yqpuXNuum1hYjVaX01/ugAeX/P/DFf5Zut39G
jGJ7mTUugosryUZ3jgrQNu6JTaOHJag8mlrWw6hQti4yeKF52+fOJB4wisGcGQLtg0nwDrjCB0wE
jM4RqrFSbO4xyLyvjoDmIRqL06wqHx9hjzs/r3HJ7T19PRqsTCNk4Ccrybm3ol4PALPUYkmdJJ7U
12gx9bMW07MYMlKNK3146xvIJs6eCRxdOc8wGeFXBLlSpwH5S53AMO6qlD6neypysK6VhseAdIok
/kFbKhz805vpGK4yd3pV2fbX4r/kELZWDx4SEcRe3CzNRD+YdURA/JrvR52nimLLrVM8I6QyR+1M
n992NoMmQsD/7fq1D6nD6yXv71lDUAD6m0WGRbpLg1TOJUUiE1I/7dPY9Av4yail/pg559XzDp5s
RXieJq11pLgGD9jTGeUPaeVOEx9jo+wFGKq9unCg3Tn+lcksezBgaORCs1clRdGq1m4CVx/9gmmH
Wj2JdKPNrd7/Mnb5QXL4p/zwZ8ibiNEJNZkIVoucFnZ7+15n8XsOjB+rJr6uZALllcrFx2f9EL6K
r8b9YrqsnPrjMawqb8xjgdLfXCfp5EotFCyZtF3CtHo2YjAL8quZRIgqrO9FTQUsUil2omS19gS6
6SDmGvWCJKX3lWrrpLCTYz8z4ACCVJrmjiilYzQv2ivywBrESaYyp06Hwfs3OqLNUs5V1cvYADNY
q/mw3IGnH9CmXJPxvt8HhCQeb7OlkCdiHHVlPcjOPNyzRnnz32WILcBEWUkwu1Vv8SrrTV1BzCMG
pFb537OzbYQ+QH6umPiIw2fIkf4qU1asoWcX9ToJKJygdcHUVHh14e03B0xD5XIPX/hZ+uNcVwz9
Ej3HvkrwKd1nJltMEfUv4GL45nhF+zWpSZChoFEfHgPQ/IF+Uy9YyYy2pPYIXBmg26IRiSGg63qV
qgDKdsroKqGc8oLFqtsYXw6JlxQQR/+kOQoz/tCF2P32tuz5em4IZTkAF1IUwOEUSw95hTJty07+
dP+lzLqaLUg3UOT5F0UCs+/ez3KmVR92wYBBLqavHe0zZnBXR5Uwxg3/VIATKfYXlnL0CrrBFOyi
tcFWUccu3awfDmGv9/Uht2BOYsrJZQunmR1mBizt730TDkdQh39WyQtFFfuv53p9lvRd0OdO5AX/
42B0ZL/4XXihbuT5iw2DuVAHa9c56UKYdUamfR3w1fdoqztTkCjBunEA5xQRPclxa8IMCyMo1ksd
hzBYpmVmoTR+KwEKjLimBONt3t/xx9wkuikfwKeyLQPlVfAMXkj9Y9ej3FUrxFUMaQhAxaqN3SGf
hVUh61WUpigOZPsnnzQ83ys10ThLJ5bJvyxkdnjtRrqyFeP9IVMc2R/97bU8s+EazOuQy6lj8WAw
KzT5veh9NPUSthEpqTCozdFuZf4RDurniXpoepT9mE9fGcxePPmaWrPkdADmoVXWbvkt2xh94OTO
ZEpXvyjuMVmN5U322Ey+nndLA5mLAPqChsaqqEuUq+V9q36ZqaVvVZfewxTpLfHqm50k4YEFnZzx
RWmd0+MrHhjTj8Jq4MLnMr5MbvnHkZXDluoKDIQVq0FNZUWY6NPZKr27/BLE+R3xeXZf7CaLX5Ya
1vrb8fzIqQGMVeopw3EIif4c7E5mXiD/fOc5WUKRRji55mWySkEna51gvpY61zeGV1Iq3vSUjFWr
tRvPPKFhr/nANeo5JVN1K7N6eGX+rpt4qoHBR7JU/bP4+K356TwBdyHr8P/poKDgZnPkyAPuguaJ
RcT+KD5vMjUxa7Bh8HF6tzwEITW/70eAOH3WUufcT1VB1fVjwo5H9DUBx1aKpp3rxfVdUJs5oDqt
l1o1wp3llmXJF/U+kAwJFxOoY+bsBLWqiWGkDtsy9HBzD/qLiibB5Npsr+cEcq/k3HhYQ4KVVA1Z
3j+yCg73fBnWqzsKvnpntNbdOfmglaUg6ygWT2d8eeuTdMfDaIq/oe/AF2RV5bawFJ1+MmernF/4
BmaevpDZmHMiXPBgkRejluOwa3cqaJQjS1bA7jbWO/QVe5HD++niDlLu0g9zFIHlzclyFu6E1diG
IIBBCGltg2syavB+5g+tR+EtefJaUe1/Mjhjys1asHL0ybZcPkF/W7qlWplQfB9hkwm7ZDnmPJyk
NqDccEP07+XaixhM5LLJViXqT2WW4MrJWSqe9/gEhF2JFnL6fY/1GyZfKLG0pOIiVqIYxXYDU6tf
dh+RNpkvHWj00Mo39Nnxmpi0DClPUrxbnTrq8JlNcY+jSOIXWa8YszU2hPn2PXWchttruQozqW7/
8iuFyTEQpCtI3WPJLEKvArJoRe/QjO4o4LPaKhNxsmaueMRydkRfEpMda5ikXC55cH5fOxgkySxY
aZcq1O7wgJOS1UsAuZdVFoUSVfUVWox4gTBpzV0QCD1U9QnQJsA/gjgZ3f8M8MHU+o6CqCF382wB
Cn0ky1HPbxU9wyM8pf2EV6QQtvivPD/DjwdysTzfy/7Gq7rR3fiiBwrRlPTG7/yJ0SG7xmczz6e3
zy6FgCTzYtYDZ3vniGppXRFXhRCchilgRO6r0fp811g6xaqCcthT70qqHHzGg2pudh80mZZ85sdm
vzf5D8LMWU62jep4uP7InNSiFg7HwxZ+aQcSEi1CjMkPH4RiBWr4gEWoYShXkO9533iTXqfY8xS4
+4JmC5oGGX/4tNSvsLQRYlhSPbaVkgQhphWEtV7rjPn7V5DikfX3WoRUMDI4dmll4OFASjnb8ZUH
7YC8Vk2O4ieilsy5LKAQ2VdWk/QaR44n+bIqotNJKdS3BJ9yLP7LEp3kC8B/eTN3orymCXsIJcDQ
x4CcDVl8XyKzqBsaXd+wd2tteYz/waFzcgIMDDwF+Fc4zqrc5HyRMJnu4iG4WTi9NK7eO6mMAaX8
MnC3mgKE0aKgudEdT8JkB5mlP6Lt2U1vl/K6agpLSdEyMWZG7tgz2Wwhx5Nxg5RxekgpJbsAdBcC
t1i+JfT6jGvYGrd/DQhqWKdYxwdHrpw+EKAMbWmrUbN/MetQf+4s7aCKOOtLa7rGA2py8fIRxSl3
XniKoEPBSAHEWAjzP4BBbuRv/A0sap8fTL2ObHNHOU8L00v9rlznG4WvLZ+oKRV8dvFpgmUpdYcw
6X4MXYd/NKZ5zg6HVJh1LjAJ0etm1WpagyF+bDWxbDNVlH512EtEe3nQY6EqFd73UZsZgv92a3cQ
Chqj2/zHvqK/e+swZ6UstYK5BKf8TgEo6QKDRyLFfe3gNMacjRQVxY009UsVHULYoFUQsQo0voC6
mTgNfj97xWRlqOuB8g8ADjpGQiBymGjaKLiE5bbM0q/k9kNSaCWBp7Pq/8KSBC9iLphj2AqwaqaD
7ZE9CpGbAy58oajm4/74XZMaGc/VS5vzz3q8FwY2+oK5SHLQ7lkeaoOmMbeU8quw8dtzONll+1ty
Ps0QmQfNfz4Z0LRcxtL7TDcUUuHL6g5OeV6AKQXexW5QCtBD9Rpuz+NbnUf9M42fjRqJ4SH+aqj1
Jbz8ST/FSXWACFBOBBTB/QFwR7/iQWZKaZodXub3P6iF3LWkLN29TTzlJcaV5Qkp3hK1otvfw46c
vu3iLpfGmOMz/oE9ZH2GkMkQn6e1enCvAP40pnshkFomZpwxtiTQ4L3W1X0HLDFm8aRTJY4lE+gV
JhcvL5mtuvFtds4/Ss02+fkwGbDskp3iTdaYoK8++wfnCDdxTjnB/lJFvibw0AaN5ilUL5tiXSqG
ikRPWiNmEgLLIpTxOoPC/p+EZdqKJbpF6dc7fhXjZose9ttaG9o3S3+UYRjxG3wFGzB/neYtiCBm
vpKu95PsVuhvJeLN5ZEMS5jmjwHxW1jL2VKz+r1xiCb7AmYDpXF+KAIDgU9oxOMWi+Ro7arlbE95
MWhUuCTuBelhJoDIaK1MDabMQ6w1+bg53upIrWFMHgXJM1qbnx3qvAYRjHsBWq46Y70m8ymayEdv
T3ct7Vzoi3vNoKhLcw343Bm/O+mI2NFa+WRfrz6c8Xn2ICTtgjGCIZzStSL7V13gTXasi9vnib7+
kTJ8xCKbsBU+bq0q3MbHzqgpPHvkMqWaZ8cPcISxVe8eKcD6+d48+eA1x3JDE/xppoyL7It5JE8L
R7pwstmuk9DBzOSOT9kmZ4r4Hux+MX5JNZClQ7yOlcDocZEEErDcHqjoqc2lph+5V64GqxI+5jPs
xKZtOyPuW3wOMa1uNT+Qib+VTUwXyDuPEPwQW0KsOqiEUZaN5uL8d1f0l6QSUrAr76ErbCeyn6te
xhlrYL6Khitlg7+f7DNjHhZdRY0IFK8jsxsecPCmuBmOnaB4qeR87jv5WIM5gQhof6nHTe2jP3JO
qN/ENnxCsN6B75UEK827XO5c5xaET1uPYozq13QtD465BJS2qFtcQUAg2MlspSGPJS/UDrn8eHw+
vk++odzo/aTyXjQaj5XL4PX3x9Rut3xiVm0WeIJ/51BsoyZLk7biPWIffjHbL6Tap+1QhjSz0ywf
4waGVrp2tjp/eCAMd6eiDIPSLg1x5yXYLFND+8MomVu5mmmoQ2+2GSNHCsTALMJ4JLAxJNBZ2iZo
0hbyTp6fORuOldRm0/m/FS17Jt5raEsEYSNBW4NvjPumQ1tbrwxPShjolQEvlG2Qng1jmcirmS6F
sxiCQSdsYWwsYi6OFGh5YvYTEHHdsKA0L5fsF7eZdKUmjk/809moXVEGdYdFz6sy32xAvkswCakb
ZdNB9ddvMhsr3xBXEnIPXGHqJRu49oEIeHNnp1mNoLNGzF+sI6FpMN8tfmoEH0IaqR1o3ovH+NeU
rAfVd/81lGS51bY+b+/XWkuAy5Jy25LBcv/shfnswui+9XzW0LZ7Glzy70FybcaSSCpDXfjoBYDT
J0UuV4mWIq6hFMRrRh2RDf5WqTZb6PV9BMQEmPZijxUjWVOy9BAg3F/djgQTVw9zEkBbRRgA7IDL
n29APnTRUeIpCYYPC4HrERqT6T0aA0sp7t05o7+yyAoyVKvjjyujzsknrXW4n0XnEqPcklByWT6/
ptWTPnwREvLlR7pdFpLK1GZjxxS9ZFhpo7W4jrKbHNEc/tBz+7oBWVkQDpqvowBR0sIBZLK4RvfS
RRhYGjAgn9i+/y2TuRv2Hsi0U/0k9Y1MGSlV3XQOWY+APRwD/w/yG4tajtwHBYV1iZ6dsz6YHBZs
tA2AG/SowmEHRbBDvKwZ5wVuaDmlw2AX5nFDfi483tGIBFm4ljQNxtohFfkznxIjuiwOGjy5zhWx
Ts17OjWmoLDHPC+ixGqOLRyuKc/tQjPOW/OV49yyBfLY47SrxLMcOvIHCFv/UQcXM0u4YWKsJ40D
cZ7isf5bUEdVMmwTxt4nk/LGgJW/72dbvmWs9PvZaOfyU02XpVG1t4SDqTwZBdVMYaAuQi35S6se
tPUGPuyNzCHPuXcPdLv2rWz8co4vZxwNEjwbsczR0VjKTFsYErKAPJQ8hRrPaUOD8jj6+wcMqT84
8RyX7Ipw7RsoLO24FwbR+JDVgKxak2OSAS/WvfUFEL1qQqqTi1e/hBaPndIo1Nth6vrRMevFngRq
gEm8iLrBDDiyP2lga9dig9to//UrsR4KL4hHH2nIg114qmcoEgvNdCfyLu2AdFrla5SivbEXs7x8
diIK52DwethB2PCxvDZBK7zpdSrsZTOZ+YcDZ282gWj87heE/wSR2auegqTLe7HLowZCVCsS07lK
dP4I+raUVQvO5RP/FgvV+aRJFXyHLss9kjoIxkp9M0MPxbSHdy9/h+V/xcvwx31sFHwmGwXEshEj
yt3v8rpfS6A7Tm+lrL8EXqA8Ke8HtJgEo7FMRo2qlkcIjY+jhl4t5g0k5ezj8tYcIvx9CkZyDbP7
VRQOzU5W0lmYG4xeGpK3yt2hafMWWry8EZEZBHOU/57+vCT/XtDBMTYpKrIv+l4rCxLX/jvWqiT/
Q1YkQoDlBn2oCw3w1pIujA8sfonx7GGgSPSdUa8A+OTIhCv5jmQdNqCFUMQveHNVPYSfKPYp1qH9
EumkKuiaE+9H99fEiCjEod63ssbZsvEEXs+Um5WqGci2nZpMEZp+t1/L3M8rTP8kmlT3DrZQBOG5
vjOPWWI6v38mZJ1aa8LbZu4ttY08/i21TMSQ/k/Gs0r10vCUnmxr7SOpTKE16XCst/PXkG/nVY0S
4eAsBjtVeGoggwLRqtUH5c22n0U/u2Dxo8kx7ucqdweAVEq/cF/Lfm+Soi8MdvkV0CllpMmE5/Ee
b/eye98Vr465i2R1tdRy7v+T1YQlfR6OW+X1x6DGU/wBk5ymtEvMqYS02Txc/CXYRsBGCYDnHQET
xykHiQKxVl3+fbcao0kVtW6jammcLLpdD1ByiASman8Y1xWEvau8pSbOaG5svmm0Dd4CKTFyon9a
pdgx3azUf1Mm+DvtNZN/4gXJgmiUIkRQmRZVZjnGLLkkeUzb6iJ5a2izaw7Xd5U+tQGwGnH3YIZt
WLrAIHOhLasmZdjLfsPOlKM8qP7utbTHuOO/U7LemMapsOkAABrbueK2l0rHwOhrb3T4nkSOP4zm
KGnBopAlqbSQC5Ohn0pvaBgeFN6ywBxDaSIShP/8AqbRmPYjcKN7xK7oOMkp5hlIGJXBnotiUU5r
3GeXVtVF1rjyG3veawhmqU/eNJr4Du+/vOKP8ti6JiMd/vpWIJCkkC/fKBydWistC0GwkTt/pxC/
blj/zcN5/Kd5UYIEJcqyLiMHDXQf0wCVGJX+S1iEvtdRDZqui8mZZvCUBoZUaP5Ohp1y4gnuntho
T5qjDVJWm9TIrhaNWRoQf8dgTZMm5diNuPyRxu7hur9QFu2MK16D5LvGfwboF/8WcW/WN0n9vpvC
8RPWiM+HkYNu4tv59D6YsFCkS3yO5SUKdRwxFd9doakQgIyv8itRQtaz32LsPvh8HS3KD2McQ+l9
HcUCMR597N1LRgnIsXm02OZlJFfSKJNU9kMBOqIOzqJONPS/7u1xfTJ0bMtbAvlwtMl0IN25RKQN
l4mEe7jPP8gPFoPPMJ+oEQxbi4k01zzPYGpkvL10kBoU0eGZwXzc8ddAnFqUPVStvHrm4CBguqah
pgB6VARgCneNuvfIjzQ3n7tX+NDz9tD3AYzebq7WXlrg7p/S3TjMGCn2GpWakbRdNku0ZirpMplp
x4JYNgGNuZR+mLEwP2Tv+T16hpaakxi48jqDOnrdKrHN2cWTrgna1td7l/5+/VQuUKaJbKlGtPGV
bomd5xAJ5tuuGjBrOeRmuOzDZzmSLNNhl8nP2lcUcALpynu0vYOYFmJRjRBD1c0X4+Uj/u/V/471
bybw0frbE8vc+9gfW1+qopq5/Xy9RaMK0WyRtUPPQzP1j3BaHQ5q9/0oTjKE75DIUYyXDmsPLKKo
HWCq2zTMmRKK4sOGPo20nAdIOWx1lINvKSMdR/3DOkuCT2EsrI6/TYk8y2JsX5DM7ZYroKYVGohb
CeYrLi5LsQ3BZWx72BOyJhjcM+s8MiojR85D+H4rvT6Qk4kH5kpbXZOhkSj+0DeKB4GvdvcHFqC2
57HUS5NnQlcGC51wQbHRYn9WAWKsT+4UzvPU4radS827VQIcoDBzhvtr1i+Ske2uMncqMzZcM4Cs
RxdPTJ4C/YObns5I8eiIN9wS16HXEi/ViPsDAYjN6urWla9qtZ0MIejwxyduftTZvOBuw3hNIStr
A3Mo7iobSEhNVcFxvdL2Mq9zJbNJIFAtp2nR+c1b/VT6OUgsONr1zulhy7IVh6MYrk11/jrRjIMW
LvHQEFqBnPRzCUdon8wUM9J8+0G9Ihy1kSbrq3T3JENF5jvBZRH7IkCjO3tD8RvRxh1TXMh8Y1GW
gzkGx3pbEOQm/qN1qzNLwceKYCrmL3E8vUmdQdbdjZEA6GjvdN9hU0fXXGr8Zm0oVM7uWKhy+opM
Ay7MEaXVMnp+QnewFYC/8tZe919WL1mQnPUPEvo0O7fd73hPQCkGq4gSM28oF14IaYoO0tkN81Gn
iVXpv10hR7un/qyQtqIqYJkzHYgdGqLS0OO+m3ZS4qzLxBoYUN3WH8g874efKjoc20w6OAZb5oeE
w/9+YyDMxUbnoR9HbBps5wBBOeAxoziXiXObAv5XrCytXTQfM0XGW2MP5+p773GQc+x9upV7NSCm
7ruUs7qjvnPRq9PpLmEVNHcm/J2IygLwFgZJ18+KAnl+bsoIIq0NexpjlK3U9cthsoYbrDeVVmlB
1/4PKEjM8cnDeZe07lFZk1riv5sSmICblHSJK7mcipkYTvT2OPsYrLUfLdkcGQKNAndvd4BOz9y9
MOzGImy4oI3hCMrm3zBPB3JvmIDfFl68X6iUuze/JyTHJtgNDpzPFGI2dBvqBFJQE6nHYHLdxPVu
RHi/8bEnk28PHQ0JtMLE1meGShmUPvRjaehnt2jXhWo9ugHrYydLVBfU3dYF125ODiLxUf6Z12fu
Pl0kPBDAgr7HHosES2FnRCYID2cr10bCWAjXvlQ/q0bZAFhcF0Bxgycx0BcZQriSNrr9TtinwHcb
b0KFgKP6XPTDIXW4V3jjzsxSfgb5wvMSXESLmNFgGwmToZpSym8U40uRXklN2R+2AzyUxBFL1ET4
0YLqfxGnX8EHcpFlK7by/Zv5aCEalRsCPz3LfaeLSGZwM0bZrMWkhav87May2+u4aX+iG2BrMai6
PBQKetExMvaGD7SMffHl6IszzmYrdWaD+ALkB/auAiWljcifMmJLW6lms6mRxe+OLoIE2qLnOFJh
Yy7IXTfWCrXKIxktNuXQMdtLuEJwZszjM7OgNQpIAKEhJsSnssxWgTKo3DsZhm27r7Jp1AbOH8rE
ZEK4YaLAfPVvEPXPkR2mtYRnUjwelQAMtJNIeKL6bvSiqcUrcdsb+4NImlRFHvsL0BKiB8JxcPUi
0zWZAp5mbucbjfwWr6TlLqEHOszOyGm1hBcFD51wxjL2CnKjWdwNs8G+NV1hnGT2L8i/MKx7YniQ
sBHl2D6zlEZhoACUewk0zfr5vvv1lIMtk7ZpwSPw2XwimeHeILAAGQyydE+HsSrq3LRs21zBI+46
O6x4NfrYsucwOU9T6N8T7fsvAn7u5ilC2wbpY/SNiL+s6+UeR0hkvBOVN/QGuBhSC3x4CwLzSu7x
gvbT11cuDr0amgXKy2Ofp9LcBME7lamZY5TW4Hzs6tNIsXudL5RxbuuY+H5Qnz4SvyMUQx7O8tiu
FnnyoeEuXXpcScQ+Ivucovm9VQAnuCTU2tQALC5hl62+Ir15NYiFlJ8nm+0dyTiSBz8DN209SQGP
UVzQG/b6YGO1QeY3frYEm1+aN7IzHP8v5zsXnQmD73w7mYg6DgGnL7JoRqersLq6WdVcvwcLUeGy
M6qZnDvr58l2WvgHMBqOr8eAyi5S0gR5JQEdMa1YV3ssgKTusH8XioZV3VvKF7ZM5UrD1vq1e676
3RkJMy+HtRqIQjxVOGCYJ+Zik2QoF3g4Ao6LENBaWXYx8YWpBz2GC2uR5K0dRwzHS0cjWQDcOn6c
PjTBl0xOEhgV00CVmlc43GQR4xOqVlG3s6zBrkdjrqaSp5lyb88b2nmahThdQ3rxLBsYCd8oaj9D
sI3Uzkfv7EiDC7lJxZcnD6w4BH4P2v5kt9Nh+Qy7jolxKToyLZf1FRAFnxmZgb4qpZ9xJfxTHgwu
yrpLoJFxMdB5z0pjq7W+8Jm+r5mpkgH0wEbESJ3jpA4lK9PZUMu5aNNDSIAakihnBeZ/myY+UgJJ
6bkDhL45xV3HkRYJBpZo1If191xjcvK14pPuCkM1cqgoLHGGXKsfi621Hb+n6Ru0oC1GwoW6KTrU
oBZESGXr20tWUKC5bQ/fcXkE0lBXo0WoDoTUmB1Htf1sKGvg/h2XLFnBxKVTi8xvS4G0aqJGnnJJ
U4AmOKB54yA/rTB9/Y9eln4bAuBPtwpcKku5vWyreEiW+7MSKbIFjLGa6N2tCijP6pzMsGr2zITC
ihjke4OYc0wYKAnJL8Sw1E4i/1cAc6zBMySvwTbQlFz/4UhHc5OFdJxb0JwmhKg7kgfLXmo7I9Kg
cS/i5BPYO7RFkVdLrPQt/S7zmBHJ55dYy1MLcYovpb5xdGLvpVISYlkXQpAenmSKlvmePOezyimM
PfiJ9Zs34oyzO5Bj4f8WKrRfaEw23PJGecsXAdap0rd9BQ56RwubzguEkS6SkBLseyeC5o0Q54D4
0+uIfNpoBxs8ViWlT+J1UIr7trEHcNN2TS1MJiRiGYsEGzHFnjSE9mqgZO9HnkZug7DCWGdEFaqp
N7uZ4/uYVsO746aFcXLvtTFke0tjTHnuHkl/3N+5f/cXYIDJJTovQ8ZrWQktfkwUnngZQIUPgZ3m
rmvpX8SxOGuYocA0Apm38aKBJR1DGO3CTAlDLobHpsEUpKaquO6kvbyK/SnsM0ByCIA5EA6qM5gt
QH8vwtBTdcubsrdxPHO+RSepxNNIw4NqYsCFnEY/juAcQbjpB3rDd0kgpebL8iP3HqrqQ2Hl5AW3
o64xDdOmC62qw5BI5xpO6iNApZE60rCnPjkr7FM8ff/Wu18aCr067IFt9nPr/CmAVEhKc5k9xAdU
Uyqbqg7+/9nvKIXTfyx24IIUgWRoAlE97S1Ozf1ouJzEE4w04UHGq708riGxbJ8z4nxTOiwRzlzq
ppNszbTMxZhs2zTc0nQJ31LM7D3J/WSDaXhuByUNeDKj68aXlCkSYS9WwyX7+AkTMBF1ZFT3OIFo
AzF4Qk7u1/LgWZbH27oDe6sdb/ZbDvvjMGcn87gob+Igfbb7eXnms7APYCqScS8F4omSGMTVke2i
DTCTnBpZeGHAzukv680zdiGl9J3VOFtBwd3rGnhYDqp41BZ1b2qSIQs4omjFLp2N6uEL+13tPppN
d5jPx7aKRg9GwUunALBWYMdBI7CnKH/ZmDTh/k9Tj2SWnffJuoBvqr/LqVMGEtiaFy0K1jDOeqHF
gxh9redhG3wxysJu8Q21nlhrcEGH8nc9nLvsuNfhOjh8uH46/H7GLIUDgx0s3LIBpfWdFIsbsOG8
LEvvTKR1ylDvagkSEylbsOJXoeEnl8qMuucz6XcrLPCcdGm8dhSNX//jTqXcvAkwMb/LAmpCKgHf
EShyCfahQKxo7qIroXxafS4IcLEgYLMt+ce33ixUl8dw3UPyKSd1rLPhx1M7y4XKeb1CuzSpfSGl
UocgiY2C1rBv7K0Kt60bL6/6K4NaRAICj05xPuMRdcJa5rfPAU2I+bPWUQfunvkTMMyfKA47Nz0L
ywagQ0uHE+cYK5lJ4SLQMxCXmAKvj9ECwH1aQNV8/eV6NCFXF0WcOBX+AeSnEnZfL0LlQZk/3/DF
CXMR3gOLvYVTZCO3vpMJnxuUbDnS+wbGOVg/lFcjcvRhlw71YeggHZS8OBA5NBZCxzqAnLLiYoNc
8/W5YEwpeR9Eb0+tqMsjge1V375qiWOZEMwzOg/t+bXrWvr55vIQ9BpFV+kOuUcO1hZufNEWeYCK
k/EnPq/SSDz1qVEMOND/y6Etgax3aB+IRov4InfbGxzMWRVKi4xJYHGoJokXfYclrhUQE9mTkxrM
IKXjlMhhT76IsE5JBRgwEEmqp7FfO7tZ8FOG9f4+qBj0PGvgmJDEEGBU9ZxFsb+dt0z5aXmhqTPN
Ss62qsWKcB0/sd4LLyY95x/Z4vQ/SZT8ox68oGp5vhuLE3/V/2Zg9ohjKjzU6iLIQT2sinUS+djJ
ftLyg1uSL7jYOCySduyM25spXQLdXNC7TFIBvfETovp18eT0P9ws0N7KBFTD/GGIXCtub43MNb0Y
VNP+OS5Rxwn9bfa+QWXViXn3NycpT/hC7AiLReKemg4HlAmzP7En8RwKB+ULT8Ysa3EiJZgPPq9+
709EXFKcTnZpFAhMTabKESIWlbqwuw9hPhzgscrZu5SqAjJRhL4a7BK8ea14GY6OUzMVTYF137D/
yQNScNXl1aNkDdd1m8ZhvOsKSyWyVGZhcAe30p3Cn4BNe6T4FJwu8DMITULU596eJV0twwpQNBm7
mCNCWvSpqFXtCtGHYRl21qxU7yW82QeG1S/FUSEIawBvAM3wnx0TievPkeQjGSI4Hp/s4cEVNXAS
5/QLeuc48spnYppCvow+FZxfOA5eUPxbs0Vit7xa7M8w06MZKO6YoTsY2a8B9x23m47XFDgLB3Bo
Xe4p2KaHjxNtiB2PQWoJoz1k7fKGlxZuLAKsnnTx7VMqOCtAnyMn4ZlHtbTZIMyHsJOlwLOyX5DV
YwrwlECi1DWEpluaOSoAp3JNuwBS6r4+XYLWE3iveEp+2Eis/op0J8WGuXc4e/K2mSzV/4vwHC8I
As0Zuf71oiWay40b5e7hpdKYGwlm5RwlGClBWjeTds06YwBQ20xzPpV3LfOAhpGeWigXkhin2aE0
r5dJL+cAJw1sbEsLkx2VS/hrwP6jvUGnan5uAouSLVlxOnioual5czcbfYImGl8BM7PS3jVNfr5J
343n3SC/ZOKaVXFj++gkBP4dCzTD72zIPrp4XdA6LWocak9WAzUQ59csKjyU73mPONmBo7rRY29g
OOsWcJDDS3ciLXq6dcuT+8uHfYnZVevKtDJUiT+Cm4dncosx6eV0rPYrXzgds3H4/gq8T7+hYtr6
V0BtnRoHlPrHzmzqr1NF4ngR1J9S4jHEN6VavyHXGGiR2PqnPwHd0SLA7LBenlyFwj02Ncq9PGZL
idsTkOgVsjyBCMixgBtWttzoeyKVO0KIgNu2UHP3QggL0vja6wOeLdKRO7uefs5FX9CBiJqI3oDC
uaBAa0DvcEmrizUFcU73g7iY8+o8QNIFb9MSGQLh3oR5vuFQ/LXm1eV7qQFBdEJd6GB96Nckdrhc
EFXJhQr9vrWMOxWXp8CxZYKQKZ6ppXSO6vAGXGv3nxGWHfsu/r6DcKX89q0a4mo9ehQuCpaOI80e
VI0GavG8XjDHAcLeba1dTJvedd2OCatavV3TKjyxST3IR/xDIP3xH8MG14tB2M/QJ0lryggx/+Sv
pidDE2ybVRL5EFV4mv3yEScwn7RN4osRCnp++OWaK/pik9D7+ipQ2xk5KyeQFfyZGugDPkkOLKbG
GZfYRnChAK02ipeuMjgCfaUheIVQ0kLRnXXvlX1FL6jF4B8RSISdbuXkVsqJeJfm88BynNFHYaw/
z+cUPqN5RIrkV8sswPf58sRNQNFnu6P00rMT7Tz5be0Q+HyAyoj1C9hM+GS3XwKFIOgpr6ws7kju
saGVjCkz9+UMgh6n947fbf7raY3YHevfB5roeBErYdZ1ezMJdmuCbAHqytBR5+fbjotEtAEefhKE
H8FArkIo9VHTPtacwQTcm0quoSKGPKZqL9NJp27RavIIUO7vYeN290XzB5g2Dfk22RL8SQyIFzla
RYnY8bG4ZTXQiJAfCc9jERQY5KywLXKDgLa2EYJSqDlvpSpV/MwkkD9FqDkFtIywXeIyPDnrngqg
6vUfLDyNcLIbzbXSD9Dngd4EKN0XnzEslmLEBd4Ou7Dw5VGtHBLxKOtWfQIRAL3vi7fcyp6yR0T2
oJASB2AdAKrb5r8KaErUXSx2G464H8cTBJbcUU7Rt5huwqLerwFhJAn3ZzqgBXHxIfWX5SjBoFBI
tv/ImG5IRCrh0UvYvXWCt3jIEVWjYYEP9+3WqS8epsKFONxJDN6Te6/9U3+/+X6AG6lGGKcCoQLQ
ILaZScxgbg8eS6rb4KqTEt8sGwuaNR++bDkea7Z6qMOeSlnLrYQ2Hbf9Tag1W2PfVjDzl0ZCxIns
dNWfpHIIzTr5sRigQmkGDO19kgtW2HkztCS6Vn3DjoUPukfRaa2tIKu9lRe6QqHvoYiRE1h9w33k
FlUxJ/rw/HiT+6YhYC35seTfzvG4XZaWiA68DBZY9lKGlitPgP5tH3PWdLUYDzUh5xGaGSmBczwL
B0Lg/C3SPvJOH57zUkyiObAjPO6s5gEe4uFZMN/0bWI9BgJ3YD8PwAwI5bW8F8FUibV2bfZADVzI
K8uN/pxK2vjy1Y1HJcoxLhyNE7o05GKH2SDN3+Ev/1fl9pj735Fw//t+r889krYqCznShpkLouio
mG2cW5eKtAPmM0F15wI/k1ZBtiv9ZbcMWlgVhVKatrKTauvPmgW4tBbcg6I/8Qq/6/roXsNuiBR5
SoF9VCl1JMybcgCTiG+gh2QzpGCwF6neLU+zmouWoK7MWaeO7n6ZcapRgM8DyGEZ0OaHhwHTkQT4
GVcVCNlVVIZe/OeSweY7tW7lqgkByp8sCVMmNruLd/mNOfo1Vh4/vzC4zfPZdbc8RoB3S8tnk0nT
fjljNtKHsadmDiY05Yk1Q+H4uPqaJxrZv/isdFUEbbzyj8tjOYLcDoQv5veYl5DfMw37TC6wCWwc
z9+wXHSNPqG0MW6MnYcF39j02K3E67ilrcRFXtjJg21UqV8icI71mX6a5yj+eHIOcOUJI7n1Z7nS
8e/YTT0HWJs9Q+Mx6KDLR/3Oqzdw/xGyuw+0z4JMmkc2kGeHpcO6dUMp5KlzYgDdy8nNGE9MHOwQ
JfX+cmOzCm7HQngfuqvipfYxqpyXyepBId4ERfBb9CIFWJt4q2Qnx2meuYg1mXnT0RwHAaFueeCU
TqTteZtDk+ekCPVeMrbEn3Pw6Ib+C4ywhuN4KAeWXvaxHVwwbzmMVg11VXgRiWa85zhxdHdNZqSh
t9QDuJdNm3IIkmYbgZMXxpYIfiXiOKCDbI4byis83t7z6GzqGwGggWHnJ4vM3cjgTZdhCPBpaAS+
moX5dTp71atxgBTr9r/qz4gxefMqQeAXgoaSv1NbW97VW3Y94/0UYRma54WAqsoaE7wcEft4etqq
sUYFkzwq5EY4/0d6RQqPiuZljUsm92gN8pfXH8eT7hUvvvu2nnDAORFgtFTv9P5YW6AIFhGDW4jW
RlJo75dFpkF9QUY75oXTcXVUWjRVNomPe7kxciKe8XVwQKyyVXvRDkak1uaY31rMmtP1KbS6GCsO
CsaMha9c7STCvhJ3vSKXqP97+Qf+/4qOyNNtRzpzPb80wWtCr8jBbZvaBiUIrcBrjvXgwySh8Qsz
AWmR/8LUtLU5jE9Cd1vxptp91B73Xg8xQ63hwkmItiy3LjmuSCou+3VRcMrqzqM4btZerEv9yPNZ
C4R+aLeSWgX0fu7eAFih4vqcbWaaiEOCumvovkuVVftkj8RBYkuCPv2kBcKW77Ov69Mai7pKXDYy
Co3P3qKB2DliFy1suuZeDCi8YvCTW8B70xNXf80mZ2lJ5OKOeoC9J47TWDsNTcrJbHV+C1IpMwdL
scOO6O+MePSfGofe9NcdTxyeACOli5BHzIxZ4X2ylh3wNtVetWzamDnOPs/QYeGsQtZx9CEjB5Jq
OMdAMw/6YnHXOgl44sbBKu0QatYDGQArTZ1lFhDhppyVINtSEH8ebYxXrnII+Rl4U7i3QugA2tx4
4g5AE4tW5LesfWlLfiId31r6hWWtvQEkQJyG0gRseImyfJgv8W4gbRlGghaz2AfbeiTKbhiGhTa+
xS0FkpCXhph2Sdb6CbkdTAeopIbi/3ec5pefgg/SuEIfux4Lwv/MatmJwBv9SV7f/jtun+JJrShU
GrYFtHwzbAI6xZzfqYFsP3uZnvKYRPl1JG8ubMk3cWcsHxNg8Usv5LFcui0chUtFGAqoHON/yv2z
njz2vBZ0+NkXrNQqfDqA/9tk/nWg2wlVShWQPhGU+NaMLve8YMvIBYvZoWUgDox64N7kh2OBKC57
0nvfMU6fpgUBfWJ0vqunDjfGPnCYhCKhxVdTohBM1ImRIuECYj45FqNoraHiGEgjf2TGyUngpQNn
GuEMuPc6427cM3Fs1+M5Z9jkSebMVAMazy5x7o7oD6L8cIW+5dZsDM4/VwxnKH4ictlYuOV4agpb
ZuTJ1grenid53H1yTAlKt6+UAzn8CmwJ0Fwwb0RvVY+bsfJWj9qd0R6JjSubLzm3r8jj8txn7DGh
eDkG5hmRl6eqoTalOyLmTw0Bn9uwxNmKFIguyevoGqK2xmuHupuGNjhXy9MEaSVIk2QAfNbgnlKy
Qy45/Nt/HEY4JmBA+gsOXa6+NYJfShoSGaE57ykMXYFSN6jsU5N+wHLcBL1Ivs+ojYUk3MSGxPZc
s6Y3Gc0fZKvhDi7C4KIc5f1KE/7Ulpua6XsW8fDXgAu+6wHsJ5XWG+8/Fm7DIOggt/tKvSzzaZbu
wuI40n4sIQBLY7ZqqCTCaMot5lwz6x0AWQ3xa1Xc0SoZwbhitA685GHjQXv/gYN+MA+hhIEc/EJz
q+4csP+S7Xzf+HZ6HqK1PhTznS5S3dCzAwqRKp8Puk8VnnATe4DinEdn6mXhLW/AYTQiID1Fl5dX
nUS7QkMjGuf/ZkO8xw5TvigtF88+4u28us/8xujjlhW9FayUfFTYwqlwdbqyd1oHnaDZCdPAhRnJ
Vj3OJasWpe22A1qXGXoQa46mBtQQs2cb+CL/StJ9/lL8fHFPPQici+FQeDt7NYtq0PPDJmV1CXLN
uGNwIf/u/xkFreXVfdc1aF8tfIi2vsQHHdgXuLw3tsAPiZJvYsksedNdJLQpbhpfPqC9zkWO1YkX
hJetaaUJ0tr3SQiE4cc77gbASBWJM7225SjhpRgxj0stUS6xqAmwMKgfgIpfT+LwZTjPcmBfy8Lz
wSSJ1MG9C3N+sVcLz8jH6CagW4rtyZau/FvbL2Bvl5k8heL2x2c5ujg+FjlgkxMcbN9MogJGTTiq
p1adHb72YbjFgjYpsv4OzqpoVYHjefg7rpHt+HIJ+NM6BL6SNOsH1r9r2WozmWtx+/h3J40QF9e2
e7HT/FeYqG3JdB9QIEVY9JMn9u0zM/Dt578FlCg/y9IG9KUWv/tB5nHOVEdVvYJDerqySkulTGQC
m8AOeGzpMMhSkXFifK/XW4wTRKDwHTlKhvv+PYk0rh2slnQggk0LJbux7is78iw4IEVHfVMZ4nmy
kByTqZTe/tw0XBzGEZlyWCH1w+nBU9P+MM+HaIexsBDsf7pXeZy/yLinUitYUeId1MpDh1WBxZr9
UiFXm1jC6eJxDTIoN2ZIysLf/EosHHt6u2f4IzVvNT+I9c2kdoOAeTVE2khIG1AqgdKGnOYqnV9A
Z7+W8TI0goxEjujqGtK+doYSljMDHZcMWxAhmbxZkYkB7D+3Ks2JZzcrTXUPhNQjNvy57IJn/t9G
QBaKqKO+ecTJGDC1wH4KCsxspTIiQeIl+XbY6RsOqHw5KhFPo36J8e5IgDdkWPTYsrPWdp9CQOYb
kJZm6ESJamX7wxAabqphpz0SCJZemEOpIZ+d5xD+f7rqgYQtVG8cr1Jtn7q+KjJc5ubTwJ/x3XSR
/SGgWFDG26rfpymKUrpmjoBCl+MlZ3QpfK8dzwPyYo5lm8oYoirMKgBsiwXn/QVoaRn4S0MRbAdj
V7KW6J7oWfrVATNIvQgDa2RkapwsIRJH4D24hFeLFmygoabDgc1d6cjUQhIF34ntgSNuAYAJ1MsJ
MmDER5DCbpxcGEUiCzODypEpcQzXt0fKADokkAo6yandAZgkPztEkiRbQdjBLyOAD6hLOWfl4PdD
opokmV6dxQk4lCOlUNuLDvQc4HnUIJo/7yKxCNg+cjJ4SJyHcGh8GExooOjX0LF0CqV7cmqrow+b
vgpo+c1+b2q71Km/AcdCReWJtqkCgsEhqmrCdEyrTZrxutDLzXkNA7/BNsudxnBqxzC05gwEO06W
KHNUbM2f4ucP8rploGUvX5zl2bi3ygzk64n4QEvJtb5HNQ5QAUq6eGAXvfxtVBzz/figNMlYQW7w
KOJCKgwtMgSnVoX8w0KLW6/+RjGLU+pLkVM2SR+1udtgbWRh+Su2X8bmVKjl3QWdYODAe8of0ASA
2MKtW7Y4UHo+PcHsvDCrL1m2B2rKAqsFUmFtp+seQOPRDmrYCV+MSFuSc3U3Dizq4IE0A8DICqvH
ThC10jBlMnTKdCb4uCqW4oJ6WHjuAJ0RzJ3tCswDyi2+jfzVvI3vN8j/YRmtCppi5a4uvm9wjimh
uR5JP0UN7W3kHktFsSVn1y1+iSqMENOrSu1AlgUHC9dRNU/aZXH/ft3+iKl+lRjhEyOkD60HAQCf
pNZB3Qyn871H/Y2wEKRE1WLdgIf5B2ChBoOcwJFIRRwa81WT/Sm6rJQSLeD4zoT7bDhCoBcg+eoE
NujtsuMLkrndHha0KxZKKuN590e4GQKcsT0SA7pRIkQzjsFVxoHVqiatTIehN38IKjhZFfB+qzwM
V2ZQqtFzX3ZYc2CDW9+QmYdS2mwIjwITFDp6elm1XpEO5A7Xoeyn4mBtvrf6KaDsA9FZ0koePtp3
MLRI15oqu/8pijeQLNahqzRgFta9Vd79NOnz6Ptn0a9LDtMOjZeoqehbvx8Mjy1O7JbkSJDSl7US
nbZLVrjaOFrJRrEVG5EEyGFy1Ckn6RdURUm3kAqEE0Yi/Oap5X6lgZY2lZCx6W23CPXsfTvZ62Xx
tG3sdiRUB4vvHBfH1Z6g9ZQCaytWbmb6Qp82FgE/hJLhHApcU1FbQHEWbjmKtKKIQdyG1+Ow5MyL
dnb6TgI7gQ3x3Ji4n4kNwrOh/XvxsK+noLNjb5GWZnuxBfTWrEQ4/TvR9bBNCjf3jOhPTEuojlZG
BohVzk8fPCA5SeDCxO4s+Obpo5ZJeGo5MH0Alm4Gl56sOjIfjLgNUCPIFBgWPVhtV5RcltBwigTC
xE1rc8i1VbMtnd/qPKl/qtc+cxW1iysVjhzY+naMaXqkxcs9F6EzcOBhgESjw3pzFMb0sO2dwrEu
ngEeZWAmgwado26keGhzdqZ5lSxKPlFlgsh6F6iHsFtPrNHIJjBL9mE0ZNB28EXCkqxOSbfRlPRr
a/yensUL/IiRw3gky3yzOHUoOvO+ThvD6EAC32JG7LaEX7zlcGV7RihxCMjfL/zFHby+lZzdVwVI
NSZPkyIw/f5nLUswNLRmGQtbvLmvYrQawpvIDuMw3Cwbqk4wPSyDC5SvicUSuveNZxhGLC+qwGUq
j33iGecnJSRlpQAM2xFHbjcqRnE/JK+xgoTI0Gz6/S37liwHDswE1CWNjvt4XcIzR/NJzO4m149F
puGzYwO7Bfkr3Hf8P5kmbDjJTT4BpIIslOtdz15hLjdUIgTTjTkPY4uC1LME9v8KD/DNMoH6NQVl
F770j7e8SvrmjDDs7uvBdHve8v3nVUVZECFYNvcMR7xO2DAo63FRtxEh9Q0lvsuOfqtq6IAUZa1q
CWNMxQ73znb+y0/oWnz4zUJ6lXO6J+/tgijhCVy5ynmNl4agr4gGzGDWO8Z3x/iEleFrs1tckoNg
ya28VkxBe5NbPCsCdnKayePY8HdECES5Vh7H3YP7Z2lFRnl3AUAHEzYP2IUBoB1h+AlJMAq/dmpA
Eq7PE3oqN5bzJM+R8ylkCBNHlUseUNekMz73M9vlRA/9xedqpzBEFSuxA+N6cwe36TaP/yyTH6XC
PUjxL1TEj6OwVfyLnR0oKqMSJ+FwNfmY4K4gaSO7pKmk9Fy4QKiNy1UiPLmhEeGm/uh3jMJifsT6
qUJMa3rgkMmF1kHiCStbSIA+ZtGfWhqhpQ+KN+z3VN98y3TIU3jLwrL+tnqFM3+vx0XjKXyjIvuc
lLBMDrfWTcNLJAzuxmQfaRqwMQDUp+VDY/KsgIqOI96yk/1C5/hcn9kiH1ai5ZA/aWxa/fwYgGPd
UR2yUfBQrA3yqO1qRVNuZzOGRr2og64HlgEtceQRv4O8C3hVT/PawluIa95S+cBjZprmKyhXj8cI
kTDfboDdb0DYf2wWvVeg0fTw5zxQXxZ0xQTrJ/HWT91Ne1RtEz72d6jCpc/xh6GPs1WIM8xty9CS
G6klFnzZNm5reUWjod4yPbjH50rOFgAc35viz2M+tgV5/KgJ/3ouVV2TyGEUh8CAGW1CZGaR2pDM
PTVmPc4qULwnYUmktZ89OqKj46zBNGS75y7x3Gqx3oL50cya/cYFNoQQixVb/SCl4vu3z+NTjE/8
clpn6yRL8wIgSjkytyYmVG2KUT6g/EBlXmMg1fDOZ/wa/h3Ofj2Ij8SR25mt79R9tm4FgEwlENoY
zYKZ9tX0zeTi5tPHvg6TxBGUeUQ4sOt/NugPjk+uw6M9qyrI4kfkBO4nn5E4j29as+GXswlJM/JN
iIovlSgFTnPSgSzMeoWAOP2mb1cBY8IXBa9M+UAkkz/o2uPz//+UNdzW444LL+JzgLo6/8hROpSQ
aOAn4jL0NVD7NfNqXOQG3f45pSAxtvxFCsFD+svw5nts+U0iW5IMMEAIYMWxPne9xoYJr0Db6fUm
elUbofkxUoAI+7yHltBPcuRpt2oB5GGjNPR0KmWNRmvNUBgB5HUS9q+0KPpq8BlmHW4VsCAhLd8h
EzddhaqBIL2efBteu7sjr/pQmFLk4be1SNR+GEHPhxpTCoBE6V8ACHA+3Tb8Cpfg54zjah3CI7oX
306DzqY7SVeegfxGRAmO/KGpYme8ZpvSA3SM0s9U1qTlV8zW9/7ZXvJTbH88rUAQzek2U5gcj6we
IU0EHDDOaM+N88JpevkCWskeo7mbZAkyRH+EN71nE9X3z2XDD+HOOfaet2LCRMXBG2PqtHJhVWRH
y7Kp8fsG9HaFNI46gwCrcp11BHG4W9ciotMquPsJJl247HQf9Ml7LIfs3bMlCiVQLhAeJNstV5Vp
IsUAs65Oj5IVhKAqfFH+ohghWyKdcqRm9fK9PBQgLeANYoLb5rjO9AWf6+vcfIntnJzFcgiRoy7q
bgOaj12j+0sesF2UESnvjcTo+A7BCK81cXNgXG+GJHByTrcm/03c/72xeX+fzvrI357W2zwQo26X
x1c8mBlVWYRLIRNWUWLk3xe2qF7YfoEBHYEfy7v5KyTfRqcpohURDGGvmQ0ocIra5fuJ7l3EcsPP
PIVXFSsl3MBpNreHACcy9wSfgLDP00eEXzhg9nrcKhYKYNoRLflfVzp+TbmwUVoC6GI/elH21B/P
2eaZCQKE/mm5KxIdrirRO06HKU+Ogd+F2fbmUsgWS07KEb2JtnauGem1XdvBh7vRDWkheAzLtqX1
RBR42d90IzkIBo4YmSLBl0pl4/1DPWB06p2YjipMUAo7w48ge8oB++S2dHRmNSbYUfQ9V/DVgcw2
CIIVmCbRbyHUIEmE2rDAbHeraR7N6WTOF4S4lPB5atn3dei6/TiHJiSTeHQhoXEAY5Mowfsx+xgS
a3ia2PUAgExfey0vOqTaYepFyqGESZzPMFOpqY5mz8b0fjsMNpdGaxcwHULPdDD/MvOqiBMhxthl
XorB5/Aj+cm92YK3t6WOh1VW1ClEVX07Ozx8sPbOm3dHUxl4TpuVznQsgV/CnXS1xjI3EcO1l/qR
1Asm7wzDdtJXEzcF8C0Ka+sxFR8T5yU9sNu5ueiacjDM24EITG+kYHU2l/W0QPZfkvdpQKzfQLlI
uheVD+/1ihR3F+GxNGXiTtrNVnG/JCpWEUsK7DjaiBKF6R0jy9sbFlhEUE6ykHtHYiOHZzDp7Rwt
u1EIzyBVMNKiUPk6lYlkkeiloiV1NOeZcAka1j+eFyJSmVjXArPhhnmvph6AbDy3z6cqHAktfAWM
hyJ22T9R1bNtQtegwERqPcLhHiuAyS4OrBaUT+yw3ui5wUg4jUo61bcXr1h5Dqu0ilCsGmwcM/M7
G8+x7KVwq4LtgpcBfDbl+pT5eK88jGaK5FUxKZ6WhITI5UmGeGQUlzXxpKLE4PWN++Q/mxlsyHh0
DTKbfHy2Nd+M9fG7e8e3hKY1vRn1zh5valQwlRcllW43eIlbkCWsaN15Zh4UOcgkn3E1JwRVpKaU
p1GIt9nn3aBeMw6HtkEGqzeXueeEyMqWV9yldMNtYwgHjkkABPFxd45gEt83LwrGQTTBfnyZfVUN
YmF45SM19533zMssc40y/j1uNzCH4akk3IsyA8rqRR4SVihVmqQZRSzweAqap52XwCddSgqXyxpN
pbAeXHcBITCLtL5tdD/KxhlywpLSxhz7yYUlThAnQ4B6jk0fHxZYgp5bGreJFmaT5X2/g+IdTGca
Q7N2ZYSBzNwSpY5BaKMxu2ZdlYzKnQF6AV1SeWJDheNomC40ET8zGjXi28cXpfQrnUSZCtYl+/W9
qAfQG0MGm444+adlIpM+rTrqZl1FqCsNIIqCzLeHlcseUeR06XoAShhr+2p6+J0GWS24OCFlgJ9O
I9/obt+hRgwDM9a3CkK2BlqWE0AbfAbBUlMSIIRq0blfDAaExEslTA5URXq9wAFErQJUBl0hQbKZ
PU3IwoCUSMyAySh1JSmnmpxypfyQYjItAkxgcdFBiCXS9eMsGCCx0bOEx3IL8UaWBYlgRMPJcpFZ
XgZdMsLbqnYsHWfEWumD0A8+0XGwa+qSyJ5Z1iBbfmUwLGPdNKEQmvEoX0mrDMnZrAR49r4QzCQo
k4dyoT2yU2t8TL3Jshsdct1ixn3l1W3OYD7IsDw3wK634ewf0wA1Bwznx5W8T536cP92vicVtYtW
oi4mcVPqvWscXPPbrFJS7YkZ2zlE+5mbwvAaI1V2Gc5yZgezTULVJcvsGV6a0KennZ7KB/7RM4dR
rp5WlrIofaFEoazczbwdQcMfD43uKIx/bHb6qpIOy3siiWnzqTofrN/lHDRjWuhONlgf09nTxb4O
Xs5H79xHMpzqUGWukiMPfH3hMCKp28N0Ohy60PRiryp6F9Niv82h2MKRDORHDQ7f+RoK+JbKdh+7
U4zmjFDs2v9pb6T49+8e4tX6q6u/7sZXui7H+BQRS/0iDF4HkXsfkuh8P8CmAP+dYOcOqJ0uCcjB
F/UsBVisFap9NZPX+qHe/w/mgonEQ3MSeb/6IPloasYwYOuZlZwh9BVfgrD4F2XV2LPvpAaI79oG
3BTkML4aLKIhlkV+wsRt2Fx4xCT02PM7vXhTZXxc0xV+UbJNdFBm4kD3fMXyFyk6bAWIzswPeEVS
aggDPWxggBjnMmHwR+2LvTTE4+2px4Ko2CV1f4HB/uOnVc04hWUMrZONDrJIulXCktmhCAiw0I3m
Ft3/8r4EFQIkYcZjfkM/lSLNiz1suTP4UobWgjEugZbCX45suDlcqwgibQ1/wq68UOYVS3Rx1ZBS
S7W6dcanxLnrsRC6XzsQmZKAmc5+MmVPlYPSwZ1K59ePzG7XBY7abPQ8jAnkXMerrEQgwBmH+YFK
POzuW/4Vl0HmXLc00P6pyUcFrTWeAJEJIOytvm8IBQTFzpmYTmsoCttDrGiJFeEXAgzqxZl4+ZZI
YQjwggmE5C6RiqG/fXIC1uqtIymUnXCLI+9gpFWn4hzw277FS/z/xIAJK65k3euqxKwpfHpeIvUt
Kn8FrRXPmgl48QmnP64NMbIcdJi7FohC4xKRhv+G5IMB8LpNeWbzhSP7O0ZJIfhOmK0hNm8eXJ8L
645lRRrFDZ6GcQW2YjZ/bITeXk3SVb6hBD8VRwGKbGh6/OYOSlmYDWLyq3f8/U89ZZ5vkYCq2YDb
DqsXiKNk9AbDG7PE03hq54YCPtfAihXPxXnZm57D1cjaPdLJG6LmqPK08wANAhq2EqUMciE0OU23
cd5zncd/aWWe8fb9HIwtlOI0kcv1narmnIjHgAjg8/q+Xg2+ugcZro+37dA86eoLlDt/liFrp6i7
ysDbnZpBrep2n+mRs5DhvJLZ4OgEfd9Ws4yKtTNJY4DAbRrBWDMplCixLYi/5nbOnY/CygeAyeWU
LkZI1ft8iGMcKJh/ff3YrS1uWC56rDTIwpRRgP2Ik+3+JHrD+ji5DsJprsWyQ5yzpUzrfw2dy/DB
NnuqhZjHS3OVUn6COazl5OBPfoD2ckqTMIScfVoWXQLQ4tE94+Du7eSY1HHMF+90/eMVyx4uV6s3
Mcp0OtiY+Q6YOHOq5RjF6+G7jUbNqX/ahmyp8TQISMUIy5O9hUttHmqkYixUCp9wMBl/eISV3meL
Rb/77jTZhTz4P1HJvk69fHywbRd28JY2DHGedfCotM4qw/JfO9ikyviZ/DYSXKTZ0iLmYjBKtqpz
iMWd4b5kP+cOHFOMZ94h6L3UUI6pnwLRxUEkRtXqzcfA4qqA4cd9NeNesE8lAWnYzSzk7TJqcUyc
/r9c5jFNXC2FJypl/+ioh72Q2zYaS91UTPJCLNizqKb7k9dB2FGfy1MKyb6U6vO3mSrXjJv07sOU
V1Vf1m7WUTg3LemNLziOt3/HaGVl8AD1U2n3qBHaZZ/zFLK9+XAUPCLzfLBl5HNQHuGQgmz+HTdX
j6gj76Q7L976xD2LIOInrX0kDYDvg2jdT7CfxIAT6iKrVzOSwd9pG0Usvj9K5sTkwG0XPIoHP1s0
SNdCSXrIJfP73tfRz8r+cbqQLbKRkOPLRtwe5ZXUwVy7vVTP68db1n+pyssvKf+tbN27f8RbEDqB
lcS/FR46A2yF+7Uf2VOzhyFn2cilerCFmcMFPZT4RPDo3Vt6KkBfS6RZpiYYgOA6LRiQnTR6oU/X
2r2uYGB9QT4lSdKVbO4sHSsdfG85NbKxRfNNxy7i4A3A45XrCo9K5ghraMzMCEjcY9FayOwcmD1t
LWRhEFEM5vQpBsKIFtDJJFKK96ZVxA0nxlWkjCf8yfAw4MXgE4a1BXuT7nan0UBc+RZfaJYZjLli
JVcy4nHK2AgE64DvjK2D8szeS5XYVy/YzCJNBoFvtY/NaLbvifU1Uj8B0O7nCZwUwIZojzuLnY3w
wdH5s3YkdqqB74Lx1hsGZdMOQkJaxhm+/+bjcA/JJst/bqta2OvsTSpsQvSy3BEAdiHHy2+mOcDc
CBTWT1CC/AC718zBqmRbrJlmzf5yKZ/AR2J9d8sGzV4DqMqO3Cn2KvbLLygF4Tko9niiNue/VGT5
xttpJXoZL2yi/U5/UejPWQWZOACGTR2AaZRGWZBbxRwrnbdCZ5PziaaJmQ7+IreB7zGmDUTdZBFC
s8GZCUs/oo37WZVFn/p9+fEu9zQKgkMAzVzfIIfCzcEPuW+fnB1GGceAtCuGUe3Nhqsm4pjaZzos
6VuOtL8W5NEznP+90RJKztT6CBN8wTj1jhKNPbSjN2GlTHHKyiwvECwO0eYdqtk7nia40qgCloC0
jDVhHqRN2U3CffinlD3XcVXLbsIjn2RD4exdxW+QZVE0QFyZt1nDEzCd15di3G0wFx+7Ik5KPAE7
bhTV7Dz9N3FHK22AVFubOYuNUDWlI2FKBXeY2HixLam51VyctClmoWxTyor0c1dgfFEeAiIw9Kkr
NzCy7pMMSu0SRUaTCtmcBsUtMOenII8EBYNJMHTxeI5ODtHm0x5yZGSkuHEjCbWm5h8jD38GXy10
I5sjIK3cqAd7Ssl3+OSvY0KNm7Og/7Tco3vGmPE6y4nB/l2AlFM5hDrjbGtuVbyZWCL46aBvCG47
OL5hnEHz4dmv7dhwpZXYNeSKqt8Wt6hrR7RVJ9842z78V5VkKIjZpyRulNfILBC0bLHNNRlU6jRx
t5/viyoyv8iEw81QS+WSC8GaUjZJkDOw5zdi3qB+X9e7ypCJkuNjo2qwxwouFEnIplh3v7HvHM1v
9PjTM26B8Hn+fyFdDDRByLU5IYGUGWqzRXGlMC4nVofqzs84MGTTxuk5RmEdmOpJCAiu7xKie9aD
aPo20bS+e6Iwov+enq/tU/EBFwUCpMuOzItGcSSg6N/F3Tnpx33iT3CgQiltSz5AyGWCQ8iuLPmZ
o6spgow9XScR4q7pahmRy2ZQqyVsonkGcWs6Sp34G/5Y9S3XGYSVPThDxKyfBomOnv7yLbOHAJem
YE9UY7DFJD4xU5NKYOwhfnBFeAft12DPGRdgOUXWcsjdC/+7uVE/Rx9tLar2OSswSLjLU2mg0ULA
SJPG+/5/j84gJq1kBVJW4mwCuO8NxHoLVWqoCSnIb4WypGaUnocQ8+Ma9SM7/5E5fmR0ALDO1P0f
SCQ8P46XFGKiqKpkq22mjaATp1RkP1rDVI7a/uQ9pIHA7EghX1LQfrHGTYqwm+OwJXBWIvki6E0Y
jCFcYowJd7d5nJi6XLtL7tjwv5cCcC2sdxZZRVi4ZzNdj08Eq7p+pRRCkXJUOjCbwCrFeBkoYbeh
VKI68fN0HXTQLDVgf3AiHkRDCcaVdtpgxzKo6up3NsFCd3Af6bu3BPV5xVoJue0hLgLuYEg4fs3f
JvNxnxhD/hoSl42CyG+3/UPn+ua3owFmBUAHpLpHJOiXzuf8Lbat97o11lvr2PAP+IjbXy7kmiA4
sa57uu0/RC9rHkCkawZvamrlFqP9/baKzFzMOW4t3u/u2mM1yUuT0BOQyClg47qB63cA5FzO6t3S
g1eyUWVM12hIHWXNeIlLeGKLhKDY3Pn1p9zTn14XAm0Q4dceAlt+iklJ9S6eHtbnCj+y/eT+hOHO
UJ8RqKtcMu4vl3+DrcMl6Xxo65k8U5Fr9NOXIl3thdrv41pLYt8oP2smJ6PHsPX+JeuY7cjlaQdf
eM+TnLkT4MyGkfVy6BjnFZk4ZTfv1O8KFhihuE2/fxBJ4CtLEniYVu6uWBb5/jcH5VAJcDDTyLy0
f/LYsG8dvQ+FF9jFl9EwI0CP+C2oPjmIQm3XM+Olol2W1cOV1EkVcfHxKed0xsqmEr1aN0HrlCms
BYX/RNuI7Fn+zCDgD5PcOkD/kTuZ9F7ceiNGWB2UpVLbGFJACOvoAIIs6xflrDjOvTE79YkcgJYW
oo2San7bTQ2TLrA7l9J/ivtJLDIC2Tc4ecL0zcotc/IqhKqVwAaFcltBupSU7AMIizcJrYYMOjB7
wPZUns3Gp46lkHx/hYp3sXxDecT9tDDAME3eLZT5livfxU4A9HFJsUlBgSJIyy53vKbKarYLyJN+
gXEVv4P86N0PkEPku4Dk/GLHWiHt6UzXgYKIxU7pjVsCRvsIIOFusThWtcv2eGlaESluZVFOYjnK
lYq+YTkrdapiK1nbVsOm5TZ5q02mHCW1TlBrAYMBAEdiBzr0ohIwAF1NJ/PLjOktJxxjFo67DJh6
8rJWrZdql8l7nB/Z2cD77VEFhLDwfQIy5TxVfs00EmRETS9emu31W2f2yDSOpB1wk3jWl8NUeqyI
nRhfSOWifCZQ1sdySTU1ETe1+zFSgv3grw1YFL/TD/Si+Fvyx1OYGEfnCHzfc4sRVDA5VrNAYiA9
SHx1e766yaiLOp+IyIWEC/wOG8wcVkLtZ9XBl5QTistY6OVTM/QuyPuavTxr2q3obJKrvhi8PBX+
rmLa1C2oW9cIwB2axZVpYTwKbmsTZFsuuP9xUC+T9xhw+HV0s43OE1CAz8gGXrbA9QcfoYyJB7qc
mNZpHU6Oh4ZrLArPMhJCkktqTTWf/Fk1zjyFmL4b6gkJp6srSqUhA/+aCDYMnyR890/FTRgTuRcX
mS20aw6zxJdp1dhkLWNLBKVe0334jKL2A40q/2kQwks2jXhzhWQkbuAUO2ELA3kj7nuaoFM4rWOs
3Ng2o+uH9KDa6Ftbgc+0jxbp+uz/18fyXtDigjAe6+H2P5uBL9exLoQifIdko0uoAXP1zywXO+wu
5SYf/yZAjNOXeW2NWEATq9xBk5JjIWITGXiPfzuDAVOl6nulKOtcTXUiPFpfbfnl7wjYIJuYeKh5
u15M3rs9UOzeCRqDmESTzGoadnYfPJwaQCpmc2NQqxIyQKbVLWMKc2nVoV62HV5vvROz1BUcvrpk
qMbfpoaBBeuBxOlJKUKz67YywPvBmIYSVDpeHGjPKlIYskj2u/zj7mcVgP1eyLhtY2GS4ScV3UiV
OzV9lJ4MfTqI+L0XhOC+Yvlsjt8uxhWuZIM/UcpxY9Dakb5+/BhyFUyJeC99xDOMlCrrB5GQZqZ5
3//M7TxQd8OWz07XQuM3srXXZLAoho8D6YedHIOC6vauscBC+7ivTOkRHMwnjlEvuQV6pjU6hUSL
OsYCmWYwHkabybs98qsbyv/iD7IVXcCV7lzacN4vK1r111VELeLOY4D6Z/PIm1BCn0szKfzH+ite
BmI33doYDg57PHsO0u2xF2bKZhZxsafT6fKBUnCTaq7G2RrVdYNG0UwruV+QXbaEBLV1H6bwrdX0
xue8OxDeRf4W7wc6IgelmlJ1YXISHSZbi3Znxn8DdkSHGywYUw8O2/V1WDH09FrT1Hdo1ZFzBgvh
86iN2K+qaa5Nk50On/5CqPeelFVgp05ZoIe/qYb6Y/uPq27x0IW4O82kVhYYEGzs3CP302XMeBuD
HHKcwxVysCW48MX8kPCERrzmnlbNmlcXqfPPjjjuLE5fAXNNPUQBVqRryrU6wHVwoo34QLm8OmUs
ax3uTK72fQ0MbaEKVimm8n5ZhSY7uzR7gQiDtInVsKZmnhP1rs58B5Hudd+taUV+PvJBp9WR+Q6f
zq0ROoKpEZkcrRHyWhdoBRkBwpGptQx1Rnief6BOGIgDtfCUsgDsk+nUi6unnsEvdoJl1hk+oSHS
Q7kpQL34sUMz/7esJrckv1L1fgHRM605f7d92XCzZI8pHrEA4MzTT0lYLCz3yE5+LJcmrwegUhtK
feQ51UscEF5JZ2fwSS64Astq+ieft9EkTs/W7id7Wmd/FTXUasltYLpJfkbmv+gkJ8SbtWS7wLKJ
ghpt2+c9KpZwT3m76TXtIPCLD8css+wp9gQFbURAoBx/TBs5dQ8IEHhEmL1W3BTDoX/6lhFf2YNY
KjB1E7rrjSCMvsO0XlUQCbnpz8o5iTFogqYW0Iac5bjtJWnJ0S3WDMulCJ1A7Ib/mBiJQyFnM+xG
pOZi0egDcHSlfi2aWzSZzaPHpReYwl4et35tWr0gEflJN4XuN3e8bcLTA4ar9AATfhYe5wCQn46c
N9Hg7ucowmp/0PMuAHNLV+7Ap4CiNDT5reWhqMcwp+ZP/gTLbGG8v6XDnvx8V8QoH2kfTLpSuwuU
Yv5rRNqG8jJ/IFhlTlv0jWQU4kd8EijCrMFoLT0raBtea6I0IsoBKP00GKQIJo20tJsbR7G893fG
pB0cU7UfWvbrRUclpYu4zO6rOwEPW+R8APinrDW8hlKBbe+91KjUbPK19C0if4JlhfX0TmRhnfIK
MQk0dwrpIVw98iMgzWJXm/uTQjt2mtsUqJPoTDfeg1DnQ/VX8MvVVaMfwtDC/nQnwKE5zlbnQ62C
j70agx3kyivsDw/juh7Vtdaz5BtTE9DUiB8Qej0nql4ILTSknD0UDudIae4PrLB2fKOKqvN9Fm5H
ISBHRquHr+Mwa764FoH8qzknsGFeHMbp1DiGfhDe1Jm0/7RTKfPry2xDmNMIuLg/gbu9g+2mzPxI
HZZwgd1RuAR9s01I+3er16E50gFJTDbDS3wOhSpGGdh2wwL6cutgpsHcTzWoTzfZwkXvjuaeckVP
V+IgR2HgCa2Ad891QQA5wVlt/h64hRQ41I064LSefYJU2hlkUmEzKuOfaRsi8OPRloA3saO/cJzE
jwQDxzDbsDtO3h37XdaJ1kLisudiXUU3mJBEcEXUdFmoL+R7cFR709iIfMnUNpg3a3YsMiR//w+K
Q/JvErcL8xD2xRm/oBHoOoTErS14Kdtv6r4KofVIWiMkfpJIK9mWhbSlN8pOcCcaftXpq+SIu1DA
FEiFHQBGhAiIuUdEn3XUkCXgTc5M2zI5qu83AZNZPqBwIqvwb19aj3+RX9UWS0+5LYs4wt/uUTZ/
N4Cij6rvRa0id/U5HBOsDAVGVUsJBZ9ANCz0LGzGCPoruEgFVfQ/oFTmycPuZB6jScfn1I4x6k2u
mG9xANQw2Z4mJnKjmkeqNnl1EkZYZVQoXS8SflkMY8AY0zQtOyYbI9aL5FK91R3IHabbBx24jjmz
LPTZQrqRyg/lDhWPNcyXGidk7brlAWjQTxYBBwlh3STB0eyk5AIU2zgHfRJ83hm54A8iwXNqGQ1y
V+PibWX0q5wB8w///xaP0dfUBYpnZf/e0y6kJeloWZQXGDOTeUKXztXaXuiTRA0mlxhMskOTc0vJ
Fkm4lLnkeobcRquRFX6NENbYOug86elHyg/QNfYl/lB8Q+XeByBzfK3OSqU0gPPGZFgfM2e6K+cS
MnOqmsoY31zfSuhRmBFbCJCdIolc4N1cxM18RVbP7xgkT412uFyzCShvBfArEuLXxK19Jhyi+3yn
CQGX3W9p28aBMqFpvZFzWLYLkaqc3P/cxcUlJedg3Ei9YQRCZrujnIUgsQoCqxQX6kLdy7JamI7V
VNvGjPW13350DYIQuVSrpfn5k+YEAJbfbpKhWRGjehjMvW03R61zuu0SNFxHxIaK25utCdUzGAG6
9nq9r1oEtLbDnsSUfDiagS7/yOoY9aABYP/X6b3OpM3nkLf++/FmF6XJQeCnOyqQZvhj8TbOneGm
J8ruA0IjgHgD6WWc4K1k/qMALsiv5+LApr0K6QFdoxraA0Zq4+Xvnwrr1KcUPYNJ7IV4i8t9boIy
xKszSMXyRWXohxBiEs9PD4ixcSbjkAVz3UbkIuFnDVCZD8hipHq3iHJ7l6bQsQ6AJrIayGX7rqUo
SFvdUYg2Asz51Gd+qMY+srQhxhXD1Bn405F4bSE/nrAsXZ9CTVp5o0DiD/x6jKqf4iqdCBsCQ5KR
/Hssost346CPZn+YOX38Bitd6QRrKWo+wrYGa8pmTecR+DZP7twQHFz7waEKSDPioe2WklXPLVZS
W/JwEZXxSFJT8oMaCQqWvxV/S+DyUFR1gR6K0LqHzdHav+1o6Hb+MMfh5p3KHW27GCV6dSc+VlxT
zFzGpoMhFu7DFdvSwvs09XNEKSYS63Gbpb/mBM/4FoAyvi96fE+c+CuB3sMqXhaYjPQixsCfAZOj
vIOTuNKZuTpe3RuySV6RHhF9Xb44oGx4QXJYQVXlcS7RG22puoY/0JwoSFeBTuzXIlyJhKlqShao
82aOiIsfck/yLZOu0FgW+kd0N7v0cATOSfV9uqOZMQZDecdho9tLBun8K4OXPtI0l3jSFZA0qMhT
OZAIc4m+moMEjwnXG5h9Qr7ehW6pouJtyTNgw7/PGfAXmNBKEb247lyAHnnDNNZHQ9ts2WNaCxC3
p5ydByI4RignMcALqq8jVSDkvjGUFNsNv6HBOl6XY7bQGIuCzovT+3zYYO+rp3rBVFSrCtEwSJis
ecOxrKLXRXWPHSd330dn82vo6kriLdKP3/350VzjI69w7WPGM4QlB8KAv5OAmJHb3qU2+/o1UOKx
cCVV+ojMEVx3AwS7elIJc1YknIB1J9+E27FPzhsKeikzW74Ey9iO3EVSZ4OTiSyG8u3fGzmq0PMX
a/IvIbYzO7CE6PIJ5YEaqkql6hoW5UcSC4y9VD9HLnRTFmNjKnPs9zz4LzTCUJ+On8oGbUMKjo83
aWPhCEspW7fr0OXFy8SqogZ677+b9lcJpBm9sUfRXUcgC06KTd+EaH7sR59jCK5JuzkdAKELfbge
qgnGWiU5A5Nx6kKtunIr5Gc7XZ0CMMTRKAkx2iTxK6sYlMYoOr0Z13904BZETikTMiIDYpGy+13J
E0bWw251/phguy/6hb54S5T7PT4ZLOD+TR9L9vEsoLw9UUvajXdiqKXT2XY7FEtvBIHPBBf3Iu6G
+ng2gEbJoTyn2ZAd8TnQPebLkFo/YnH739HBYMxbVnRrgvfT3NYw23b5dRNjlkf2GVpm9dnvtDhr
MH8ks90BvDc3MZ5m877r6S2xaxiq2c0ZdyvUulX2dZWbNc8MaBZaJmdc/Wft+MlX/IcEFgImc5ud
lZlATt+g2UJhC7b6SxMfHzgqPpVX0qyh7z4aQTnOD51dA1ksNE9a/+CMHbeHzOFD4prlWUsn8+r1
9rY1tri2hzteKss7Y3Ne2En5FbbY3rSs7Ov+xM+un3Q8VefCl2OmP4yXErqvdrX75keUxboBAcZJ
3CSlPDMm1mUHHS3hn4/5aByYoe1uBEBtT7sCHxWd7ge1ABUtIAFH8UsA3DIfa6ExkIPKcDV7AZMe
Cg9RnNHAO56yM1cLinPLIt2GlhPiMcrcgwHN5RETzt5BeqlHQfuN8wmTXCCMjUjikKp3kqVEi/q0
SDTvrbrmqtZ4Fre1kzgtqu98JzvH6BSVFX4V+HRIvbk2DGvFPUTXX0GIe7SY5ICS+cJX69FgbHkV
PIDIxvGXuQKuL/AW80IWdpFhJ1QP1qj05Uq0IknscbYHRnp8vqFzm6w76KTuzFbfLnYyyJmwz8Mp
b4k9WbDlKXCkufFf8gEribXuNIz91GvF9kicDt/poxvdxBqMII66fEkArIYfKPk/x/fKOt7jY0R0
BzE1o+vFs3vb4Oa9WRZLTEY96P68eEEAbbc31y/BYyuu421sj7jcL4ClV/rILayqFKDdU1K2re0z
0kz0S4aXpa6UX7gnxrBdFhxsbUyQDgNW2tHHG4GBnEbGml3KRqfFPY7yedmpx02i65BFmVA3iSrz
3LFxLsKPnbZVKlpNwtFN5pvo6f/xCc756EhQauw5CvspgUyEQrobB1MwO+xq0HXGrux9tzhLTUDG
bORdU4Oa0uGCDd9wfJ96+L+0IQEZ1g2hGZxJ+zloGF5V4oi/+8NxknERjHWI/WTsvgZHQ2I5GnZO
j3+l0zOGgOk7QV1TVNjwt/ODM4PUqUIQUCXEYauI27mYfM9EH9hkLHASxGxDPh48Ey395yGwaG8c
XMuPkkXdVtmjj3FyhtOe7cZyhenLB996Z73/q7z2c3Fk8AtHDA8q5BgxDyi+/ONFf7pSbNyNDMFy
q0UkKTeQdjLFsEVWlqnuyMeJmWH11+fKedi40ceHh3RROBMO9MEtk5WN3Tw/O8eIHXCH33wd/+H4
G1gmK/FlrLQ/h9fxtnWyQn+/53d4cRTOdeDobFPupdiIjvQmDa06hyA+PR+J7jy4NBenuR4o/pep
DUSG9v0HmJVj3rhbc1x0CjraDahRUUZNmGWb5zfz7ofpv+OkBzSyQeQPub+rw3oRfpBFvoMQPJt9
bSPVAfKm9PDC26lt6eEUHosvFHmAOcz20msSCigHkj6ueVQ3HA1+ST6H46gukQd0OFBw8RUlCaXd
ym+YTRPw6aG/TyX2fO3D0rVQ0L09fFUtkfXWjyBEzGkhSZL2DnJQ2aQbSP4QCEwTF14hzswCQRKX
S4B1reGgJQO5VZUdvEjAhACebZYhvolKRIOZXYwaSxHq8lTOXWMxAlsTgcqXIj2Kvid+nLYRcadl
uwIXn4F4rRUwe4g0y4+JhNea/J33f6/2pOQylLmbGAxL90ci0RLFwEKPFfJlNAvXaJn1tPk3e31k
Yt+/Y8f72cow0A3tykp+3krwSaWIMAJC65qIYSOwj0KXmKPMjQZwpSqQVLw1UN7KBLqNPdQwHG4P
6NnkdH7w0sl4CVPfyZceeXrtlCPGx/avEr6soVTrww2w1C/Lql6nsarQ5M8ZK3o3K2mzq08E98MO
L7OqUQsgd7dQdABZhXuIKOLWrcrqvOoJJJLsRtEfEiDgS2aMF7ycBdY9KXLHmupV+fLBOuDPBwzQ
XiC4WkY7cqFm3Yc4AjB6gTUIwHtxRBUpQ8D0oCpnL66d3DFi0rWzVrKt9OPkRdGgqT/puEab/Ad0
fgtPD/t7KNlFwswlBdHKig+RMBh3WOKqDVDDhFNUe2Jeg4ovwmXgQZ/2rnLUF1hqBxu6mZKFbGaX
KLny6JszIeSmXLSd11q3UqTjVQYhKakVnvQGXjKfyxbItmkuvsbQoruKsbDrbak5V+cxvMJ/I+Cu
2yPg5ByGdzMmPX5KOdtxyPvDIJPerzIicwQNpM0Hdzus3zYCiZM5k4Lj2QFvXrqrloPKr9UEh7J3
WYNVzny+Jb8SIYDVuf77tMuf95gGpXCRqblAJnBju2BsuZh252e/Bm+XZBxkUDcYA2VXNApM114j
mGRx1hO6kT44u9W0shZRK5NOlO+z+Kc8JFmHdViWtAHO/9we9KphlRe03LJgwKx9R/gotkv+ZAr2
Ll2/9uWO4LLP+DXzxppWy0he2UQe3rj5b1ElzKru3L4iNJvR2CVkSGICozU4GFRgzT90OtMht77c
h9vd1sQkZi/2i1bOmNfXnGEXTIEVSCqkABCWYTYBtwLacvwEx+wLjGJQFbUG611yuSGbcUP5koz4
6GdXwYWnQ2B9wtNFd1cU7aZB9qRUZ1LPR+48EQfd1k0B+OtutEvkmWBb6HVyMive0/SefqPO+TTC
ZtBjBqObPCJEFKfaftoWmy1YfYISkh/9W7kcaPgqxCCfzkIQEetBKCc1hghONqRcgwcrOo/pSNP1
lICV9+2K42rNWUTqn7PrMfo8Xad3+Al5gtzfPumwAWWpvChv3h8krm80tR1GKPHR/Il1cT4UgpIt
ZAA197xCEgXwQYa7mxmdTzmVtHCEGyi9bCqFH3S5PwwUONltbQBHMXt0PKP/gDAl34ra/rcDq2kg
tOgC7WD8Dl6pT6fFy+E+H7xIJuBRro0+H7F/LtqIiwJCOmkWC7SG3OR0IBClmAqJDYA/ndQMq0nq
uRfbuCzec8dR7pAMrpjqH7KLHHVxPXGrixXZPBmYEjdiwKhsPVSclSbDpaWcVL/qJseWw2nmoVWN
HNKXmZGM9esBkamLs4aS4GInMV3tQqX+d34QIHCu0AtihIWd0BnV4ZhoKF8E58CrWu4NwrmfqR69
E21JzEbIk6t0h6pGL2sEroljd/PS3UQ+GbMAmEJfF0OpKxlW67Oi3Hz9GXZ9QDS+CiP6BxuxmdbR
gnT1ED1p0uOt4IdNxq1o0TpYL/5Qs1vO1u9zombPCLHJz/Vfc9EeHYQ7hOEoEwlndzxSUAUKThtP
YP3heU43TreCeAfeORC7dThCGgR9VM0pewYLW1nz3h4BpuldBz8T8GUo/Uf3FA5pHTWVoZ5qv3Dd
D5IrjRa/zkZTjt5ghpa76HFXzvMEyOG/1H4kFldXyrQo2HQKIZkJ4ev2GcRtPIC4L0ZPO3C5gRT4
IrcnBw/7lYubpCXY1ikyMaLuCff45Ai0FABsy8GZeomVmPYcEU9/mpMfA+vAgUv/BhszbsrpHuZP
2eH35I8PrQnlIj9vvJAs5GWSWjPsAfE7jfqr5leWbu7BKsR5MoyqMNhnhYPHI5z7kuL+M4jZixww
JSOiHO1XH4p29HyL5pDaNL/AhLg60JK1DD9s3uNLkK/vmeWFbk5INh+5A/v1MGa6cwfhg4I+y7dD
t9qz56ImeOfC0UlYsIctyeVVddy9AP7ODyGkKWxqcpVn3hy/+rB/WgaWKQ3PSk0Xg2IN9pQ8WQx3
jruLYuKeTJBwGUx+BXiwZD12wlb1hym8WpW47Pq8naCAtoUYjMlxtVqeoHmpw/O1bBLEGphWwsUl
Vo04xGVOf81LQBMYDgXJc9OpdkHKCLrmjBoNGIuAgAmaAou4oSm5jqQy8EcQxeLBjM1cd0xes3GK
HrhwRO+dV/fbYZ9zj4KTvQa5X8M5MTCKNLa6u0GxvQo+8cUmPAzUVGjEKdDQetxIVWIDtOonXrdg
Wv67EDIDUQctCx/DV0XIQ6+pqbm5fEm8xfhDgPKaHL6hNqzQm04m5mucuT1RWkjnK4b4obQzpiwj
g3YVBRUXXdQVoEI/BHsCg5lM6ipMh9x8EV1c+tuxYb6URtUGOdxBP6JgRdpqoVSNlYJVaxqR9V67
2kF8uYTK6xidaS187fFCz5Xfwck3RkoAk+2rYCfMOh1bqlexjR4E07kN2TJX0cTqKZ11h6yAUxcY
nn/mVk6nsM8r1+/zvJoOXdO36R67EmIGPfgzJ5f8l9mS7IRiHaNK42+TH7wM0KYiWBBY9jnoT98q
rtVVJA/X33z0/6ScGz6uXdy3fLS3jo6UXtOF86BOQw2RQudsirP3XzBZO61E/GoWg7JLHnOT3rMV
bSd7OuWe/M8FmQDeLsxa4+VdmQop9AZ5xoj7Bo+x8/hjSgioTXqf4hQJUka/Sm0yuLO77S1dmik0
sbZWkP8ElEr2pLE0lZv68Ab9kL94iEyl4ES5PIatXsu1RkYQz8iWsogkaXj+OUn5u41a4oRIM8Ui
wKiX8SR5vdXwToBulrLP/9eYrFGT1AAcjWPRxBt66uCaW5zn8/rtH//bDi6PIsTA9tUN3HRSuMoL
Sw6Fol9NVNu6mQ+ZH2Np6ZxKmXtJt8Rz+jplJ0Szdc+dVqN3lp4wOaVNKR3FD4EF61CVt1cne83i
+hzV/BVyv3srN0ZWAbmeBX4BieRXUWbCkRjWUn20+9LzNyV7CUXjnhhFW1IeKrMVCOhuOonKcuKO
EvxiiI4RTEnEpBGXUu3G0cB5mzDI9dOmpNzwdcn0VudsF2GlVJmRegH5oPEmpTkqumuZrOOZUEAk
+QndbwA9ixjoJPdsFE2xw3Np3KsphWH2D7216BZajrW5ttpimdzFE+nrf7FgSXokiQedcq3mJAyv
Bloed7Ky6xUMSyRFRlQrxA+L2FYWygdR4DITZciNNvAS8c+aeFvp/eyvUxJxx/Y9ihmtrA35ioxE
h659Bb6gTnrISCBno3+YcQohVNAH+2ibqgr0VrXKS4RRl89dvgjZLmz3GdXtDicCpxzbdYTXqKm6
Ef1GC9yHhQrIACUMnC3K8kwlQKpBoztB6bgTY71gHHMNL6k5Mz7y+bbJrQ7Q+quLv20wsCf1EnVd
9sT0csQZ7SMpHxH/s4KU8peCjs+z6Etf0Eq4AI113/Co2No7oeTW9hma4cPIldujiCIv1HYrKoLl
AU++I64XPBxVBagu92KJpktcs82qcGX7kBd2vTgkgCWsX28+EJNlID2xS8WqFIyYgVKNgyfeTvjf
uI9y3cZkknu66Fw0Xq7FzKagxN9nBH1EVsa9xUOPN/PwyZ3Bcd133YtKgwVtep+KoH/d6hvAkis4
jKCwRYtQioWYfpIn2xecJsFQ+FwjzSZnMDYGE0HpuXiOtduaiUpeWiKC+SfqiOBOAEtiCMYdEHFo
4V3bqTiHJINto22MdJIuOIXHp/NnqUUrxW3KOR1dsmyFzx6qyVpOWFJXZ6TNR1A1rudsBLEoBN3h
PwQ95yHFAEZ4+2oBaTpTAgrDuxSm9eZLCw6Jvi05CjXXX+rG3m0fBuAcTw726/KjVD7Dn173xnt1
b4CVNI1zWoUu3mw5aNyVBm+XpbPX6srlRJftZ5yfiwM3NJgQ//114e4VYhSSS5VEpRFsAOS8iWq5
/4rd0z9MSDknzybNmbFz0o7o1zAN/Tiqhz2s9yLOttQ/2YDKAoQBWBWj9PYrI5OqL6XPJKS+Gn6U
dKHqi/r4FSsPNTuAyzny4XcXHxhchBXspgeDTCjtXD/YuG5acYtjJAuBqgqYcVKEvKlCWI40+VrZ
rwnYXTuznqo6Gg4DU9UTbfKXDEvXBAY4aA//55AkbVfxq0aVQGuLd5lzBLI8UNtS72gjVLVnakL2
m5x+QWe3PB4nsWD+aeMEUMOicbOvizYCC1v56r1MxPRWaYLYsgxvAqFxQpXr2W4LHSQqkNZC+S8e
DnAvEsNyBfI9zIWDPj0uyVAAlKlfAw+z/1X2ok/4+PZ5IWkVxDuEhc12bZEaXN2a6NzBTPrv4rje
uOxpJHOz+l2N9Ywhkb6n1d02eyAjF1kOoGWpFXcNLVnsELXe9pDhgC6GaypW+TzYS5QQWFVPloPv
VB5xleGNBCdvMJH9AO/eeTBUO/bddaU/0mk78NKnex4E2C/btOxHEfK1dabwz4bxE261yZfoMxHM
2CdTMZ1CBgWi2ugM/gpIgMnntnN6PfUITLHkQcEXvqV8N+t85uDSQ1N5YVK/Ppv+T4BzeVhz8XiK
TTmBXiRtFKxK9Ze+0CQoQ5ACOedyqffmcORv4WPxM6+pqGbmJkY/QmLpYTQtLyws7oNIJxvNm+oW
YvvMNKUz8mETgh74ung9IOFwa6HhelCGjp7lqVpcqDWnOFt86XQoqVoR72QqHX03gS8T+G81Xcgk
2FiPgNzt4gahal54LiL0+NenHGYu6tDd8bw0vUHGEgjbV9s2JISJ12H4yKSD0gH6GmPPBsDA62a9
hIu8Ry0BtZSzcZpSVl0PW/+Opc7zQbNmL0YwuG6V0iPmnWfpelYzxHKguDHYlJ69g+G9kGDL/gk7
Q0U8r9QXyCOXTp2rY3Je3/nENTMAxB8qbXM1pfPtwWBGJ4woJlDERob3J8bUDOPkTYeJTyKfgJ9W
FHBFaGqdhbhYDhfcv/fyZ4z5W2RsjV4/II/Hd6A7inOr58fuUPD8IfjiAbHfgL0lr794ZPtKuiGC
liADJyFqSrzm8SIe9Of994dsIBURESdMYSuy6vkM/1gJuJQTKCupR7oREnYwqN1iUR5UrDYScipa
Nn3uJ8EzSLXdEEMTeUpN2QlcBQfKRQDsCD4Z7/jGIU+UHS5iFuCFLiSSlm08+uqbRoyODFeyZUSR
tSGSC6Myjb3FN7wLPysmgQCL8cHVjc9w9GUxDadFFhQ7K9FBkDojbXaw11a5x0UdQiDzK9+jgzXY
fNCbSkFJVJXJgI9QbMXIK75zS7x/c2uHS4aX96gNTzOyLb8Qqz/Nl2EsQdNeFS/zyPYP7gI9ALzz
rPcrOAv40Ewl5SMqaAHcDV5EEHXjSbyopHXoJQnAItzciSZEkLCQH4w55uI2VNsXf8qv7p+XV6d/
v7ZIBijNTzwAiEYR5kEZp7P3M97Dxj3fL37OMBrNRRRYOvY/bgc6f0ByWJCO3mHOGZiOL+9YYlDh
LfVohrzvd8a9vpkIeaFW6kb92+wzVBqUomQvW6/ZdzNEo/ajpfb2s0X2/Zxlt9BvnSN+YZdk+mrH
nWPQgnaITu9rSV5FxMzTB3J2BWRqbkwfDy/ygCbRrbpEtxjb/ASx+ZjOvFuk2+5PtFKj6JPoPj/Z
7wBnVT/k81DsxtLtvHdDAjKc5CH8ATxPjn3tkQosiK9zBWvcjzMHwQ5e/6YuvnRq5cz4OnlHEdy3
y2EauorjjzDr8y+b5fO8+fg4l1rpMNu7UtRs4517ZyU514q9rlNt/kuvTuVQBac4nKVdFLUJs+hZ
O8EPYwMNuFEc2aRL9gAmL0obbhQTOsAg1D/UzBcOB58RlD0hyc8zNdGkwt1gsxHen5cEdSgykhec
bmA1CMtdlpaJZNIMJJJqBl8qeE7l+qwXpeCOQIocHQa5dwyYVVJ8+x0O1GYYEe8DpTyTRJdAC0F7
Is4zC0AgsfIEm91X+B4b7itgUrdqYUpECIs24QX25hWWWVKvLDUFLez7yTKf128dKG/LFovxQ8Uj
d9vL1+vOxT4d8s4OeTze1YzajkoXb9ATguVx7fBTJ/CcRT+UAaB3ByRxrfnoAk7trsc0DQbFyj3V
kJwtLcm7IbYjDambpXGeSPH7KKi1E3JzwJtclXom0oawIQMGwqOtJkCN3hFB2HjUyshLtR2OB4OV
YuoYiaOsSomFV5FH34aGgxmzkHx1ghvn/bGQ8BETdqzvdHOq5BHxyflFOBss2wGkefVQvSjMnJZu
1W0lyQH0R1U4sqwO4oA56XlEAeKG4oC4gWYNB3nYNTZxT58lupjVImODsniPtONm7jDR81GnYqpE
3dRqRRNBBmEqn2zhLX//FXb1619MJg4UBogCx9E4Lm22FVMNmxsoTuUNjWmB0he7P8ZZ+sQlVm7w
LXGOHzZxdS3xZK2lHMZjeA8s3cjYi0jIpnQSveC5xgwuv14QMW+4wTk5QN4gaGdkd6AlCkabrgII
3c+osPeSaAZFBskUY/2jPjLO9KCVoE2XbsIJ4AmhKiiu+onJJwZyOlaR8XRWjZVwHEXOLhm6qApY
qaLy4lYsm2fTL31lIW+y3ayUDARhm1kbShx3XiXl2tD+OTDdjf1jesVYvg3L4jturNLl48sZSR4E
aqM6RUqJIjb3BmkHqrhaHJsuY6ACumlBoSIfk6T8UwOdmnDKC761RrcOFkSOX/8fX7ZwwLeX5Gpp
jHcDMS0yL4coTD6nrJd5+RP3QLoh646SAaCr+hTAVwnK9I2Rby2fzNekDBtJxIzBGZOMDIevol5g
PEkCj5xBNRh4oGRtXOZ3eY5emx884ZtVpCGowQ7l7pW30aJxhsYceS9icgtiCPDe0NCtwzlaX/0X
RJXU2PMELwesi7RkwZCY4jnxuefJCjU7EETgIahgOy6dQKdx9h8248TDndQw90wjQXOMayOtKaBu
YekE7r7CbbTVyP26qkodYja80vL0WFDYNXbWz38IBuQFJV4CeJ3B/GauvVvSSUHkaOniDpl0zvzZ
bMcw0+L7wuc/2kmpE5SxdyPW6Ii3vvcvpE2DdACKrxMKIu7jDIufJtuLriINDexnA1Z4E9ULw6y3
Z8Pb2hYzJRtCM/Qt2MSs2F51olfx37UCCcquppAingPZfQNVooWd+sTQU5cAwRacu79x6f3eFsf9
NyGt7A+nQQ++XBGOOk5KN32IGz0fwrLrI1xmSBC21sJ5W/A/mq0ZDMSg34FIeoE0sFBU6hF63g+Y
Cy0JXTwmKpWDeIeZz87EE4tjSICZK560zT4G9QDOcjPzbSrY64xl/lO+VqsqFqBwIKt4adH6b1ov
HgR1P2Nj16cN+p8924ziu935zsjZ611L4ZTjW81Hoz/+PVvwehl+8t7J/XJ+5U9KFUG6sehilmqZ
xocjWDyYLBl36KYV+ejQPkzhaosIdkAgt+dYvOVonyiVdxF78EonwEoGtaNmo9Sc5mKf+k4zvq36
XWdP8kv+MffK0vRhG7Mono7NcD3wuayqsCBQ6z2SW/6Fga23U10gZbunfBvf95UKRoi0VqFTVfuc
xHAEO5vACGtJo9C47UstanTyCLfj6rNVXGUj7Z/u696rPSWuqBRhN86EcQwdAydc2BvJJ0ycK2TV
7dTdsA5G/XlcAR47vk88JYzoij0OW9irl+Ub74ZJacPmM6pydf/83QpuUwRq1xVgvq1ntrXz5/xB
esgoiIeQlmPofXl9W5iyPBMsqJ/Jt9xgm/lUYjPCWudeqFBqbLs6++VsytlmKQ7heC7CayEMCiml
Qlq7q8hyDMTK2fAQ+kaduFQK7BDyRdLSGuCkx7/OrklDDIEPO3aIulnue/S4Lm4uiW+NdeL2b8k4
siLjKCxE30Q2SUBaf+mhAUpv146fDRApdgLmHD6LtM2fAVDLAV0LNF8rMRZ5GlSHreg7wfRJM0mZ
hn7RU1pPO9sHiyHm77pXei+V8p+mt6n3rqqcdiajU9Ip0v86wr1eryeDSuZo5FsB4DAav5ZG7voz
jOV3qYJ+lM1lMokhpE7l0m5opNMOD1Dfj+UrqGXloqHmAA8Hvh8Gxx6QJFNUSckr3MwedMXzFycl
pswsZBrsaDyvq3bs+f5/l4RFRpWONOJ/1Fge86CQamgz6QF/l/i8OZtga2Qph1oVgrrGoEeLDKRg
8KNw27hAQwuXHS1wwOq93UxXlDbvjhswrwkQvHjlu41S+6ZuwVOiepDuTuBz7G3361ev1b4UQtSS
tafkXm7bVKXe+2lQI+IOMo2JO5XLag1UOvHFe+GY/KJHZgcFSp3EfJaX5lRHTw6Wgxa+pI2Jvsih
lirV0CuCEtU9S+Cz88hSm7hYjJlmiG8jz4Km+QOPy926PpPGbJ89snW9Iulxeg1ebFIagEFwSYIF
B1wIn0+7npnaEriB77DLcMR/+c1qvoCj9YGByHn4KeTShjZ+qf1KWHqXtjwbgkCBB5AlE5zRFHDs
adpNPT4OxzuBXDTvaW+E+pZS4RfZtonMy5BCbKF/9QYF3OIW1PRHCQYjr0R+7b6GhqeOreXdkPax
cWDbAyXJVgXIDue+2bSHcl7Y4Zr5NJGff5ufvYZseXWRF0795IgbZ7OKg1GZ/5lkJVCzJM51LM2z
KUcdfD87MbbS+eVcM0DQfHhbrl7v61VkQk9PUSqzpAd7GaM9oXXdjIjayWdG8uFy+Jxmfq7QiGcm
m+6JZYUuPP0ouHL+v4izW5uc+0pRxv+qTI6sZhXETKpnjNv580oaCqQj0Pc8S3cgzAyPiIQGUSIQ
h0qTs/JUTSnSDsYURjMoEqHO7d0jep9CPw0nh5nfYj6ruRSO1YMHSbfqXqjLwLSIuCdDS5/wNgAB
PDwXFl1J+kLbOWmwYgqZe56CNH7Cd66Oe+3NjgzOzRwanRZsVqupBzHYSx3K3JT3NzTdF4HGgjnp
/HdSadw8vN2LPD2Ao7i9dp7jaHdLMJhqZa1ePw++alBpILzBEaamrrYpKPaamasOqfJSQbgk91do
fvouKdSRm0oDXHDtv8U+tN/VOXemROUfwusdVyDuVxHODlB+CyXOr/wKLPFUlZgaCauGUnNVDWNd
7tfnunAjDOnEiNdevNzp3NxcqSSvxTxV5AHhYXMVr5/8iq2aoWRNwWJ715Pd6orzPfAudkd6E8T9
YeFmUVjH6QTch5DdbaXTaIH6xCAR60j+MAz4xXrg5Oy/nq97j2XihXcS1DemEHVcwCtDXKODMdt4
yOMIV01sCL5iVvSKjL3zF9kdK5wwl3FqYXhJVKcUBMsSg9tCkWy+Pnc/w/tPHwrH+haoMu7DAr+b
4g0RX74VKVlUjIHFY/BHBR3TlZX805ohyrmk4081xZWtQEVxIj6wL3Gf6fwsdBEB/H13h0UDDw6N
P0PgTv34VE3j6T/NNbnSiiTU+TMxlPkn1dZjQ6N65fp1abrQMacibpqJtQYop2sLsuSMJqtulTMf
PShPS3gfTqveIPZ3vmYZwOzL8H+rEULBhQ4QcyXXXLaP9W3c65oqzLAB/B8k836QwS46iWRk3I6+
ZrkJZcYbHE4BW6KcLTKJYN7+tOBQLqA/RmzXRsEpNMUUdPQoqn54wWm5HxRAu/ckIARnhyyrhNEf
QRuvT1uO53NRCpcxaqH1EMweSubPr88xSUD+ztEEAs1HEgaX6+/mHQL1cotK2yZF8HYBD9URpCZl
jWwLF6aOS7CNHmKcDv7RR3TdqvCt4K5QYzVSzU96g3B116eNKY7wxG9vbVcGVttnQw9AO/CavZyQ
h6KT4uqDCdpwZtEIrSOJHNwZ+gjkXzWzMDwJmAN7CgvtDABY8BS7MMtaPUDL4E+hEh1pD6drn4CI
duQwiRZuD9eLzMKwZNWakeRcXzTWb8kHMPMeAtOLw7gdZuP6LTSqVnovAFxPnc1wSFCimG0FqX8X
JYe9vh/GoZzjH7u/0TYs/7B9yvgTw9vreLZLUjCi1t45zaUSOhi0NyNgwWbEIzJwKjRXze/g/fBi
gh+hBxXZtd6TEuofiIWoRjBhugw3I6y7K/N3cWnM1NzZ7aoJxGWpLqQO8xupJ1q4dqySdaFGLs6y
didYZGJ2dh59+YVFdyw3wtjxb8jDoaHzXmdh20+rRiTZjNSW2Ewq+7ktkn21OfD3hAzaV3bxNMbR
UHd4Meu+QXvtxzawgD96g3tlTKZN4P7iuvLUixDsxc3ETfGQOnmFjD6Lba5eJlmldq9+KeN7JGIN
qjgSuN61YKCn+//MhpwuDZXTZ0QMAd72dCWU2cp2qKknWqXDTZtQLkW0pS9pkCw20phP0yWhWLaC
LgG9aVG2N23kI5h4LeTnJDrxPw47cyFOd0hugQ6WyGxm+2RQ6zpmMIgFUlM26/IA08M9ATEarJ1e
G5maAYgsBYl5T3auM1c6b4u09JC81i1Xudbb5dxx02ekVxakohgF4z37S5ey/otaHVF2yvsmO2yq
shmTKsA+p8vlnXPdyI/OdnDjbCXhm1HyW6/KM+woFJZYlT5ozvpy8AjiMwGO5U+aTGvgQZ87Aspk
peWIDYhnTBbR3NwYg+6KL9/1c/QbNB7z2dS/Fjg2HecawK6p+5tHTzcTrF2+wUZCKW633z2Hj3KY
oXxMWypNXqnG2TZWBZryxtgS+Cq9hKLkecINM2g9iXoq3wZ9DyCQ5tDS65KJR1u/k4AUCX+nbaUs
a97Psz8BHWl/0ngiiZuZXYCesT8MQrgBtxTDqZMNBLCqNPNJky6A1SX3QjV/C0B0SqfiA4keqCp9
58QEdt9pJjN/tTlLGKYcs7jX1FlG5WmGY/aACxkLQS/ByfqkxhZ/MA6oSJKESkSwGv4eHwX2dtGj
skqtqjpJ92C7+R2wdwv4fKeeaXhRH5chz8uKvz3P7/jcKQiGEzhd1u06pIuboItJJIjHMYmz7JJz
VJoKvirPBia9K6kK7rjRluBaTrprB1GjbKRNqygCn5v7TJnAhfC8bXeE3BWPPzxgRfCd/MdaLAs2
xYhQS8S+3U2s9XzALEaqL7tleyjlXEXZuh2gTvLVOKOm42ntpQezb1SvFLemac9bdocC4PISXxno
2dqhPDx/Sc8zqpDsLUU1fVtbpxgoJuSiWyTu4fbQ+AKVgjZ1oorMAGfqtwqMZbJPgfo7tIjO+rM/
xyTVfFeTI8GlzqZq1A6g47YyE8+s8420mubdqMuCjhZ7+Fk4tHtlqIoTrIpqiCFKHi0+h0Rxgx44
ao3bCEdvA+LZfpXNUUczBm2UMfBjg72EHQ7ZAVXri69K/yr1ypfO+bMo+ufAj5ICovm7TTx1sLMp
/envgQi4cCZmtOO5PgJ2goDeEbnGjs9le3CJbaqu48lIvPj8IMfT7z8XWPF9j3LsxbEd/loDqjoC
OsbT/U/AihVGFerezNfobJj+GEVMocZ9VTyassR24/seOGs96U0npHCinkf3ZgKStX/MRaGWTYE5
Fd8or7OnVkwpqfPYgp+dMfeV6ZeUegwkhXAbuYXgHzze9EWtKL5QRZmXSa5RihuHTdcF0Oc7Zv9E
hwltOdhvpTgG7/CeBYkkGyZ1eq/jnbmAPTUOKZvJ9kD/JGOTBVFhrY4sYk9ALT5GX9NAeSoKl2Sz
byZovaFgZeFeUeu3yiomIIgBS+sfCRKU0kOaHhTW39KC9CG3XCWqYJ9t5zstRTqY40O4LlALqV1D
cj+ctVy0v6wlXv0x7hIQZj5QVSUxEqJuqFVdopaC4Ig5jKiPp43enaEpSrdvSNNvb81kcLLJp/+N
KrKZYRu69tPY476jFuHTJtNl7MaJwmU6+55faWTLlPgamRKioUADYMRvfBf/8gwKnGvUpmGloPMS
lY9zgfmbsrcJ8bSTv75IgxQUlRZsqKoX0y/zbTWkpMwmMHSRPcmRYawY6tnnqOuL0OdO7Y6EEHC3
RB9VI+YFFiUYp18hMQu5WkkzF+o6xNYyZIVdviglpaCqKooYXOeJSswOhiqkoAaKkTFGhI85acI/
ftIkCGSFgdZbknIiRzAX5TvPm4CwUFUCTFoXkYWCBN7gAqtD4O6Fow23OLAQpFsZFkrFHAhnLzEq
jCp5oorF0AUKHeGC65bYJZHoFaIUeROVmEzD4zrUK/FLE9EnlHjz74vwdT9lD9wFrjOGXe0c60do
HpnKAxHwT78zWk9yMblg9qqHU/PsiqIwr5jMZk9TFLC3GLbEExpkSDIDGj21j24hQaWQDNYutmNZ
wQxpe6Ua4BEiNwRGpgCh96Fmfr2lMcU49iheaGphHqRBuQsF1zTkOnt6f+iyr2DiZoj7CgDbo/xw
IdF5c6UB0IPmYlOH6U9XJMkUljS1cj6oXbz38vbKUNsgqmoJW2YZ3sVuEIc6kpuNoJ8MK6J+wZHZ
TiHb3GwYqI/mm8P2e4Tpp84AKtksOW+Vte/OB8FJY1MoD3y0aHgwZvOeHvCuq30mTfFP1HOJ60Hh
ds1di8iYT972dlEqQvbNtswKt6qMqOxQzZHF28CycTPvcVYw7L0Wa74A8XwXVPI43t3s3Mb/H7HU
Z9GtQOgqQJb6CFNqHuHSI0nw/QVo8SuQlGkOTs/MEz2V1Dc/GH6I4X0j7gEkzpxpJP/LClPyy8ek
tLP0P72Eq2+5UOZYSGSRtoynxF76Aw5oR5iKX0k8XBhXz5/8uTP9HQfJqcpzdi+88Ft04lj5nbt7
X/mxlhZahgn2T5xrDc3paTps6GjbuKN/d8fnu5njG9M5o7clVTPXN2HIH4hUWGvMXvIe409sNupJ
c1Xv8tkgbbntxk1BM/QKpk3PFOHLx5rc68LwEdtqSvMtKR9e1kxRzxO63h05fgtW7QJr+9ftoADP
/7+ji1p8Ck/zFqK34tqJVX9r380mpekc37cubGt0C1QN6LTlCRS+8tHp3moZ/EICwYOsrr2zn70T
ACb1snpChfOhazEYD1jmSBFQitkk8jz2KegB2R97AB5+746a8sPcUUtktKNMOKC6j+DBLr4jx9OB
qJ9vu2w6PCjq2OvOWresaOmOq2dpbv6aGhdAibzXi/nwmhWHxdw1AFyJy9l8SRGMbz7HKNfS6P0Z
VTza9/MNJvlm2A8r8QhUz5nfTfAueeBAzy3Gyt5xdSJi7z1lk+uExZHsLksgsCvdBuIvlUItER5p
bBoLbc5Q/JcJOmYqg7XL8tLoop5I2+lboduIm2NaqZObfM4Wzr28+dkaBkO7xy2AN2ALU3BG3hEU
QuLUbt7PURJMmG0R/4PzlXLQzhRB42lPVKiuQ460iGhZYebHqg4x0PlFKBdX34r/KUzcS8e7xmF6
3gbjKc7BXq0DeezpHCQmKmTZUMt2CW4x61OPi1ChoWk3FGDloWq/moWWDiOUZwdeyp8YJhaq+Kd6
ztF91cm8vnHQe+1KW5e+wNmc+iJMzW+kLdTpenov50Qy05FUnfUh7rY4i9y3pcAZ5Nm14vx8S3GK
xlDxP2cbhFUehX9gMVNxF8AwecCkSmq6HFLZeTLFilrzoXZBlRm/n3kfImjhiscXYg3qOMFzUG8u
VQMs9b22r8QeDhhVwkf3LgN/ettsm6PzVC1M8VKylpA9HHK4W3RPr7ztKcXMCqjI7SnH5biXVZqX
qwtjonoDJV1oVNjYVHCYrXW65Az6oOaQAgzWtIzQtevQmXlQkMccJ3mT565y2LTXIfMMe1RhQFs7
YCgmbJJLoaeoq8+T8YU9GOst4/5BP5G7tkpa2CpGlHsI5Cw2nrQFkQUTrC4YAKstHIWd53FCvFVj
HOFE8AIbU4gbIdnA+dIybXEQkJiS1FUEDyG7DrHl99n+j1TR5giNe1iw3ahPE4d8qunUkQLjODpA
SB+P5wsZOzJr3PqaCQpigIPL+97eqWVtA35sfKrfJYF888j0yIRgZrp0PB2GHCrhOYbRceLt1RfW
gbOoVkTg6/o0zGMjXd233+pghBd42r7KD2aQye2Ljl9KxIsR4VPbwaU7HzGGzYp5ypAeJOCs5Np+
ZILgvsMD+xDezqv1/2rVEZ7h4Lsb/8RWu3qdkFRAR9ltOnxPeBDhbJvSBO34wSdTlq7xZ0PrdP1g
o0M9VCmOUj5pyU4Pg7c3Bjhe2E7lCtCwxDT5FxSHtyA+WB5wT2fH2HlsPuWKp//Gwyw9truXAg3C
g1/53xpxvCwdqnIijSQVzAqB2JlV+JN1Qn6s6ywmLDv3oV1Dahwksgt/uh3nHDpqkuh7JUte0RIo
5FxEyTAm9zbHGX6idMvPQChAHYA4hkjLPwA9Ygr2OH8PLCcuvf1b2yqt/ft2aBMYin5G+ONzvX64
7YwK529GZVxjuOUenRt8WcIB9T/eYrme5yPtzLX2y1U4krtbTVh/wpMi6yBXr9xoqTSQqR/3HAsm
mxf+uWvmkLBNkBTIgN9EFcLG29GiVhNENTRQFhiBgmjE6MKJ5GYc40Rq/HAfissecN6SB5IfxuUt
OBCc8Lh6LUPfALMUKndgoENqNP09RNgBH57aXB10QwGtN+2GRcOv0WYo/vTCndb3NhHF5diwc1Nv
bGDIeSwimsDYsIzqbyroP9EBdtFtpoqyLxV7aBVv5uh5gPqLQxOBYGkIpisQ4YYh/ZMa076WPsg8
nrr9tngZ9TfbFroTOynVRftAQi9LITYdycEXuOjr2amTPl/94UUO4W2YcE0PnBcr+FkaGPpYqbo7
eo23tvyQObcGluaG3Htgnx5JOl6M5e46mzJSNXx/b1IplkVMl8szeT55LRdI0wLAoZ8z8oZGy5TX
GabQeeSZeX0eqRoyYbWMu/NCeL9/plOtmfC3wCGJkKT1rCRMkh51bjvJN04eYnyqhf4VRLGYmBcc
7pe4iukI4nTzizHjSfs/W+hHJWYVNWrJT0s1hHDHlUcaOkKN6lr+7KtLZ+WkHGRVyGe3x1ULwwlo
hIQxlJ+GmiTyqtZ3bO9meYbMN5cs6BJdyw+4wDesj4lC68M4YJj68VuzR1/MnMGbZd9fmxJPQjTR
jLdwgnr8rc6DVPH4ID7Mik9tArw8fSS+eW7doi/yFO5cXE1kSTsCvByZWtdQtga14wa/ULA+sMDa
blk3EtQtN6Ak1qWGCVgfTJcfjJOcP5zJCglLk607dt2KNQImplKFR8hygzOPmocmuCpMBcip6HwO
4j09KHqcizNAMuap1nEM08dyfVL2bfqwswz6rRYHG32Rz9BfOU1hsO8dIa9TP4aSVH6JshCuFeaq
hIbVIevnZqx0HYt0omR+Q2zL/HMhUfCxmo8T5P98/SSQDhQdRzEsiRSErB1ZvOmFVDhw/hyWGjKn
2rUyPbsjgy8DpRMRzhI7hAaEU5CWeujdKw5j7Qc0e3uJJDWe524bugfCl91D4vSP4s4xhldb3XcY
fXYATIZhHYaqPrzDbmHeC9Wji2URlvhcG/bbPpZh8+smDfNlZ4r/SWk30NJsPRd1jseYKk+Q963e
Xd53E66YwZKNZvDeYnOZjoqbdOpQ9krrv8nRTUWWsPB9KtucEvmstqlceMn84qxOLKxZbC/O1kan
qxBm7Xfc13g/qtANx5hBEFI/uo27kXn810KssQLfAFOF3nt95bUwpDmw1TUlWvn2aWolgNjK0GNg
S2plkb2mgpq9grvFy2BtcNwoLDl1u2kftdFhSRFj+/ODYOkkPvj4DeneCKGxyGxdLz5oJWWRlRBn
cES6/ZO6rqVDfKcN30fhp2woJC+cLyLNgKcQ7KBCaFg/tQyxNl50m4mdf9esSWQDyDWxV/6AaVZ+
zgT6VHcLSHH1E0m49lo101LcLh3Z6fxfaDVDtpia6MaKjMFstonXA75VlcgbI/qku2RkKrJLbS2I
Sbz4qQZ5gPNcJdlVIdU3r21GPidtvkOHrj00TqnnY/qMNiFI8mLKs/vLevBW6SYzO8e8jc4QZJrr
hJDgQ6nWo5EuHrRP/olRBQDSATvTGeXjEnZ73ySgbq3988ric2/4r/Jo3BklJS9LauGWg8gvZChZ
2kL+d35j1Y49zPisSUT0WDCcj7pGDwUF/vf7UiZjpnX55h0ZgXir4nz4Jdh2w8WvUwe+oaTgzgzo
QhHmSZtqAX5ideFFYGuyS+asJgnTHVOfz0y2TyFijESwd9+86qGdojsuE4Yc/t/HcqRMrKWRrrEM
h00nVUl5WqxrLL6s3H3QqoUMWVUw3moIDKIdnuJx0bU4hXD6K5L3Y9k32xrQgDFUGkiiva+0jEzc
V6tGfnGvKE8C2LZ40JnR9EefDFiGNewp2epWWnIQb4SsfF6dZ1Uip9Tz7lgryCB7JP8GuL1zYVRk
P7kxc9QNuOxt9wD9G+KiEkHinr7RUvLJ7vPSLgYTBxRyxM8VTHzZZmjsqR4v10P7/kVz51XQmP8H
8bwcb6Jvk2CyVDeiw6XMU94mVHhuU3U5stRiQY8NlD1XgsJzTzye+t1iu+ZfM50rhqmLxweI6F/r
9H92EU+TSDW6Hay1jfVG+W/0GjotKYzGRofd1G4TPfPWVERYEqEt9uhqQsIqcnE9bvozOo2NyCfn
xj2XpFARc2KQWSPlveHOmSqh3qniEeMjVgQ9nSkTmUJePAqq354KhCpX9iC9aN0lVC0Sw++Czo7P
DK2CxK+ZkE4Made5P3IAapgDDbUrdTjzlbdOR0QmAH+WePzddByZbs2iGbBsPk76jLVM61LD4Hxz
o01qCFQoAv4uafvjYwrcByoN1UFjhAVXIQxdlB7l+fpiKlNHP6nPVUQYoGLuSTCL2BHHLPr1vcM7
eMszLRVMvT7jrgAdffAhGd9SFe00E7PadvzzjJ2f6FsdMmFwj8WVcFNT1BTFWwCm+lr/2xhrZSY/
jmQOo14XRQ1hn2zHz4m2QXoajCbNBwn6grryv70MQxIntHTY9VgDqcWqv9nfNd1VrCsmDpMrbeaO
SJB/j9+SqQBzHlZCkh6leEztfwt9HCb7rpUOG6oMgIQv/HlSFiOELyFXYHCfkVJd20e25KYq7zC/
CKPMTx8023UoZ0pdrNKWE+/UY3eTkbWFzunYSg8MT9VEXbiwUqEyK1hK7WtASHFWQVg3Blz08DaP
bkBUWRbJqzYmdGyIH3aP9SreA5I8Y6nHmvf1j2eTb4En9sADqvWowUW3kMOd9mmR5UQqgnL703Iu
IVmKJS4ShPwq9FwUMcH/5byYn9jjOmJoRYm0SOnswm2SUQOTnSoSE1SRbNqs36e+anbB+jUhtwyA
Efn6gKfgLxTIBjFArR3yjgy3KI9fqvndBSA0ysxusyp9bpchca/UaXWQSStL8Bkdw5kNCdtAGYBb
uqAzO4DFOHAp4k8FZr5aCTuMCfF3RUttyCA7rVSXWeZXycfEqwmL12/7mbBRkLNaRGvgvN36f9c9
uN4LnqUpmlK2+myE0jdfNjH2QQkjtaUrvP5zsG3I4fGhr/gO1lL567NEYvW6Kp8h/TnEFCvNVb8V
Wu1Vsw84MZYrjTgpc0AHnBd5bliXe5knSxh7nqfc6Aq3NVXtE5MFM4vXGCs2Ijs536SX5O08OQZ8
PluW34Ybu7Nm6gKulsHhJU/Z/fy/qdO1tg5/Q9r3/XWbNxTCj0fTg9o5+1Yq/lomhJYELCG7r+l4
p1calzcRysx2vZDW0nA5p+FqySrtY3imgs0yG4kUaiMPxhwN55PUktHbXD870oXr4MPHqY8EpEBg
rD1TJbYGlZPEcqozR7pN0dhCQW2LuhOI7zYyOrotUcofWvyEz3a9Spqpj4SohiBt+QdcBImkibb1
0ESjB4gUK42jXfi9+pSafUDT4qX1nhpZb54M+afaXeTvrtIUFKBLWWfujc/vtiWMG0hdfAizRQ2+
yrOF3Ez31FSLQsW+DB+IYtE01j/KAx0SzSfQpKSg93ikpVh4suauhxcvdAQqbyvS+ABXOdu8aK/v
xaeD6ANmox/PP1kpLH1xKJ/wi279uHF8sLXm8MjzrUbUuZdttVT2WN+rhbQkakTKTFuuhphEswFu
IzxvFd8cokL8oyZLihlL70A2BDGqVcwRdQr3MuPd9sCCIRxrXkeDpv0ycvXH0BjwENTwsWxWdYtL
Uf1AfFYmLiaWwIFBZkDMnOAW5QCVW+2G+c1BpHTph13sEn6+tu7Oy8Mo4beHTpD8ykIocNtXCqNn
4xMHcSSatX25Zrorh/Eml74KHoBd9YN8JqHFiXS5CFTpSgjdoFJ38Knr4qeW+TShwHSxG2h1fUfZ
WWMp2QxF2HLVYHhdBFGOQnv4dTaQk/RTTVdxCKXM0HPlDLnSPgqP/IsCDj4H83uuhgFXWttpA4ax
eVLebLtS7ojXfhg5veff7zUPz+5zD9mPCHDD9n1KDocY318cY1pLOocai8l5YXBSd6WEwHHYEXz/
PKd3FOGVmTX2o1GyKdnhtoI1f45lwWpZRfaef6umHsYsMdTH/NGN6kRiU7WTl8sTgn6c8XAh8ENj
9/Ov8QapALksWB+rZJz2pXyay+4IpsxP/cNUFgjecNQaoLpDGPdKRP7ha2GbzQsLMYmdd4ztAEHT
8IyCcHQh+F7e7L1hByC9WVkaWosa4OyyKVn80qIPiMyNdEo79QBTXlk/gWc62Jw2Oh8IIKhf5a2Z
e8O3dAj70aq/BGksDZUWFPyX0wcUiN+0mqVf+rPph2e87D14sW6jKKEKkjRQ5dlIxMOV5Suc4nCY
82db1HCnxcWyBk3r14mVkOap5DSpK+KLEXijSwQpJqbiOnkQXE98WUa4mP6Fy1OGtMYCGP+50hE2
TetxY5ejr0O0C0an84qlOWQcjDm5lwwHSVToaN1/A9oC+W5y8aTgAS/BBBSQq0lKyr2BI8Io59ZW
pLqmkGKXDtb8yV4YDv6uQ0BYvIkKfieBeHbRTAOfeJblycf2Gyn+0aYjQEUO4ghsc1gVPrw+VCpA
gk07QCzlSjjcY3V8fBIPqdlNRa6zEt3mitZF85Kk41LeUaVwOwmVYUCKKqifKL9+w1Sqx3c48Kkp
cQReN6YKIKQmr27tyMIAIOVwwNDsBnZlAS7qCMno0wsPfXYXsVzRofALERWsujLLxBfsLafPekmi
/+CpOpdH2JhyEfZVkrDHsu6XZqTNNNrN1oPoZPnMKhoppwUpvQ/zReX04Mgo4kiPVnWsdyVG7mhu
6sKPq2KyGez8OJXCSARrdwEKIttxFppyCy1m0MH8VIrg435UpRYCucsIn/Si1JmAHzd68oHzlIIb
4KjTTyu+n28JikuA+xnC6rjIn43qICW1BdD2sVo3HMVCN4oTIEmgq9miael4Zhzagzo+tJnHWQb4
/Mw7MAYCHy8lMGL7fTk+Of1xdXCXZTNbrPeQOf5edorncdbIa2zjHksnBEre40vE6lQHDtak2coQ
qXzHRoEHy+XhvmF+Ka0iYHYPn/t5T4lNC21oLoQqpw23ehJBQ1q0KaiqW4dNIEhNvhd5U0By4AOZ
rHbnYmgmE942YQ2o6XIqqrscHlvijUFi1UOAxY7qflnknQsdXh1g2Tdy8Stx1+wicOybbsDGY/ZL
VQSRyvxyFtdaUdfi6j3OT+YKKqd1Rgzh0IhR5xgs/CvLiFXy79vAQACP+vvwmKsqG47ieS+FO1gd
lHpVxfdcBy57M9BAT7mvXTfVG6zZE6rXCI+HgC7JFgSdPpOVWX7RePix5bIMFthd0s4nAsaJz29K
89DtsjND3GbVdFwPS0za4iNH/ozrkI2yCHpHAnZqpu0Npx33cZtU/vkuJr4eak7hd49ZagKu0Kn2
75YvpPCdfaN5dExVkxyytg1Ge4VGCJem/UAE+5yH6EoXslTW/LbJpICcUKgcQYGf6WCv7ZA/oOXj
DpZMnrJp30gBdFLt8b2/PfkJ/6xudDXfVkW7TD7CFclFDqOqFWXwFFay+7T+Y5WJ3QB88f7ouMvf
oaN8VT/Fxcqm+qJHDXXd4mqE17kW7PjAWE5iEdlhbzuQYln/GhcegW1FyASxv+DNo7KD6sJV7eXe
LGNpCF0UBLKXa4sW/CK/llJwRgCOJOkxsFt7XzDqpeC2kJ3Lb3hA9b2TJueM1Cf30t1mmHEi4Hf+
QJM4bfXBfkoc4zRbV/XbpBi3otuptPnSQLSFbDldxEnoYEOzeQ50MezYL/lBG+GaOUZ9ebvKqLGp
qpHjrLifwASB+ewzF8dWGuB+Dau71LF0dtNzLr4oEXi/PlgNhJuiNalpVPddmURO+A1CxG9oFeR5
tbStsNcRpQnxHMirR8PyVd5brZIaTOydnUr6QloFl75HUcEeVqyxwdAZfYHijr34+aLqXaPpai4Y
cefAkZN1WLlFU0RDtDLe1j+HHL3F2yqQHdmOv4AZ+ClxDDPFf3vWKTxj04EfDU5g9iNaSXziwv4/
DLvSoZ0nlIVd/mBx1NwZxKDplVbG0nKJlCnwnAyKNVlltJ00kFgJPxHpypmZAi7YS0+NTgphCQ/b
HlbOAHkwT6s566O2bKPTrkR9n2WOf/Mn/oCqsoL0ez6qTokD31YVSyXM1HAL7qeCOwGSuU/s6T0M
IDgQR+zKRsifw81jQVUqaMzPJLptWjOxcK79D4Qs1HD1CkHVZeugBFlEAnECzrWDXsyBkZVMbs+C
r6pe1ji0vWnodcFiOUw7ox1xs6Ivk8h1zg1/8iYKxd25H76XxZrwkcImRp6J6CvFwmuzOshLZ7Z/
MiXueZBWluSOicq2ba2XOpZTYsNS4Pdpglxtu3aplkBeO05qzp6bd7UrWZRiMFhebHXdSW1WEjC+
eE/ixxWdphdB9wqQRbSrh3uK6DVIWG06RTHm88duMreKUqRZqZk5ukPbGds5Fv7UU0sZoUZTBX4a
iMhfuuavoL/9Nz8kijdC5StQUu12dc5xloh+d2VzemEIzdNE3pcAHoPGzDmdSNW3RXkyD9bMi7ZC
oIU4f/4i4Jckt/d2a/DWDLXwpTWgtqexiJS8GGSblWJwyzEn9U5R6D596AtoWwoXFq5hArvVMQsq
ctYo8CvDZl1mHacDJo7PBtHj/RjMj7GarL0RBTrW4S7z/gym3vPTd83VkgF6subabnlbXhQguepQ
eMy/DLA9MeN7v7Phej1WBO9Lysc0nfk+JEBiQZnYMpOO2mRw1VFH0NF5rOxCRyEGcu17s3/3NsYb
yxm6hUDqgjDRFn5MsOgbuBtYMRaccBHbRLTgc6lNg7bjzq++u1v/sOf+D5tQ7hxLaFHeUOX+hwPb
4o+e3O4Z2A1L5F+j0ERw5oXEsqEjYN3ZGGV7L/DShXb3O+0iHvhBGKRk18qwWDPgCz3XpxGJTT+Q
hCeu3KNMYOkOHgJLQaDCicqnFWT25w8nTJaQDKvEj1H+FguRov9OANfvbDGZu6kPl0YP0U4661MT
q7p8eDWnO67NGMtQ3CfMVA0Y4qEyhQELMFEfzc4Ll63ocwRGfJ5KnLtykHiE0euC7wLplb1IbdYf
P0WkrlvfweXPHUclaogfIcipcvrp2PSR6ijQgnDzdaDpe3Ka54zRObxKJdH93aIFsKXLWr5twdBe
kfLEuIhTKWInWx3lKciopnNI0a9U/4GCOlxrBzRJzpj3qNisIo2SXOWt7z+DEOhdTNQQGXryXqPp
DrxM0OlgyaH4gqjB5251gN2Ljto0eqbtt3daJZgopepbLeVAluxg+/lMqa9HiaA910REB1HEdgEm
YVwooj1ImPvurIpRxSWD/6rqyqPebAixdHEwEENGDh8u3bLfYJrQtHioWfedjpOytJv+kaoQ53Y3
KFtDS1Jx65TkbTAKikQxUJDbW6E8ljy4IbV9SEygg4PkhQoJmZYrvJ65IE8VHGJmcMJpQfPb5PCK
4Kn1/X2KSDT4JqJUljT1WV/tIM8aFj8fQcfgN79QZ+bT5FuuO8CbLd8QTH2R+6tyubs/brhPxYbD
LAoarFJ60dGSwe/+0A5cs5r+euVb20/iOZVllo5e6Aaa6IdYtkQCd5idRP43AyaAFRcI/yKVnl6q
ES1Eg2Ajd1BUPPbhU0NG1Jbqg5G2foF4K8a8gVKOF1aICBwUKHtbpMRL5ZqFJ4AW12IVzaR0tbIE
1S0S4u9pKNoRZ3FZtQxgiVh41w2XYT1vZEREDlFEiynB+RuKdDC1F1NCuyxm/A87r2Rnv/E+BBYE
6BGPvOh0LMx6ZlI1g/OXgEHcG6kONVx3f40lJDC1PekGsQak7AZLFDSeLbYUcxTW+HV5vtaw8RUp
eWZ2PpV3yrPa/kToCrqKn/Qsx7sRJ3V4K5rb6Kas20/9hqYO2ZFV1radxrkkEaaMkiudh0FdpM3t
xUKfRrqxahG6LKzTuNjlMpqbQ6EnDUeN4D3MufNhtiWibrdhlRbNK463vj3G9+ISVSzBtRNU/EKK
5J+HhbqBC7P8mzLojrJE9UejlBOkUiOpGRhS+ItvHYbINu9JWN8n6MKsEYfCBAFYa1tgqmVVurZy
dCSnQiy09XX0nj2N8L/+mZ5A2Ea3UMJBFuw03mjoByXtfE2M4qlyoO6jyafOqizRE/GAYfQ304ou
PBdLUgsVNFvUKhBd6FlspNOu1yJr3xZZJ8m0//Y2gZ4dt3RqAEFFQIqmO/39AP3941rgGB6ldlUb
u0e/iQqHSFlUIaI3LDoSLmX4VwJTc03VsvvBJgQ37TOi8xMctOtoR3w7zhId1pPJ8gusqxNN3ZlB
TkLfCkPhn2IJu8+kEtEMjCMTDPbg9drkb4tNy8/cFDJEFdeDmOQDECcjcubdtcClZoVhIRz/mvKp
at4KA53GG5IU8e3tOWbckweewLbtpzTLJ15otSD4ompej27ZYNIXmKOL+ZTbyHe0o3tuYXAgi/eD
BNgb91pQtyF1jbKaCS4Y7zEW5nUfSgY5UcTC8FvqQBa3EuQugnLqvAr7KIYVGELyy9zXwtKfgURf
w1+Twhc0MAEsOvYVBFDey9dpfzZ2L43WfWJkreh+p/eCmbok1VDUx6pkVVk2GZgU46B3cF6zkNEK
QJptZTPfhujOmW9tSdiY9tU4yJudsccbWjBf+YrQxDNYGDvB+rkQ0XPOl2eF77AmV1Dm53Aoqz4r
f4v9dSYfXLxIr8vMcTkRhe5w95KuCfx7tsdM4PqVabc1KXJ2OeeXEWITfCYvZOgaOlVr/K25lko8
PKkME4VbAs4KIVuJjtxVRDAn8P/Vc/MFHxFPCYWYxc0JJEMNJGj2HQpQvnH+c0kIkRn5jOXyoY+l
wkMPsqhas4arwbp9AULr0WN1HE5FjZYvs22zAke3ozNnkE+ulTDHpMzGgeeriWh/fwRT1OQF6XrA
gOI0pgte53qkUrRQex54lBF99rdT7WlN94+aSXVv6018JJ6LI6wh8I69h3KlPDNpyv5xJ29zp+dw
ED3/Q8DwryjdLWyBgPjQnf33/cFB6k/8uyQVtf1NtjMmvuYWtknt9PPFQ3XJ60/trmnnUPplrZeq
YzU/TLWkPGRkZHBMPR4kxzV0A9ozXGKRp6lvkCwJivMf7to6X+CQ49sLiOCdXCw4mzoEPQG1tp8r
FZ/v23wFd3niLw5BIqSZxoEulfxqCRedscbevfCxAivDvX8tRHqb2Yz2VajxUXulDQdzqgC9MwnT
Iiok7ut8oY3RWuKy+45uBPmZzW+kjFHiad6RzovLXP+KPtrXQ+1RLPcnuWDTqPBLa1aAXCQ6TzEB
VbuDgQa4qUlJ1GAInFLudgablrlHBuHXGuK5aiVW8UpAg4KHtIVRvsuvgs3chv493i9Jvjth6Ha9
IRO9Ci1nlw1UpfRVgiCIwNxlT1S+IkNqck8FJAnoJXLM5+y++/6OLKpyU1rGpDU2EBNrxe/iOHhc
Mqv6N92uZwjEWVLxRScASKXLwCD1iV98Jjhm/gWw2VO9bD+qdGFxwILh/MNE55ZxA/cpaL/HeD9O
pAh8iEN2suux8xVy1ksFw+kXBmQOoVx+BszrKB05fSuXoXP2x5W6pn8bOR4t5M5izRQVFug8Bfkq
+GYJzA/NOEE554GnImJTLD8c532bI6MD21zxG1N+um6MPCt6OUszxf3SOQh2/IGbWe74ojIaOg2b
+PJyI3Dxn/tTKRpfhaYFZzfifuaHJNRWcXJ25N5a30Qt0FkKV2AogA0fCw4SJsMqhkvANpe5ZGeQ
NPDsB4q/wB7ZqHUkiG3lU/Xfjio4MI2hU1T1atau9cG5875pApZCsnOiB+HAJ3SKDiO9RH/Gn0Fu
QDKLTOllvW5R8W59nwhV0pkNoLiSJufQjAJwy0Z4woIYwJtpmKE1zsz9h2KvbEE3S52df8VVnLyM
RuQILsqf9s57sixMJ/yQYryydhD/pc9apiUYcbnj6g6vawGnz3fPbyTrDWu0+Qjqdar1CTW7D+6o
ainGTNJ0PL97znNiOOj22l9fPNvNhptQtNsesL2mQlOFQyqOSMHpT1TlCRAXDzbsBF3rYvJ5hr0w
5A8+ku0Zhbs9oJD4xLKd++lX/e3dD0m0A4i/mQSL5G0gQmsm1XJ6z4h/zYPKJPaC/3FUMUSL9RW0
ifL/hKpcZopWhIk+EbMVgT72kOFUqxE63IJkTlWgKQusvKK55WrgTsFFAW5FAivskxgk8uMUgpjR
rLxFrpyMBZroBOM28y91zNEDaRiF0rBw61F6hYEI0ZHJIp4KScyC/8g43nEk5hOUMZd4AP08AaiU
O5glqKBaji1WmWo/ZYoJBfG/pJRrTYFHRUr16pn4VRfG8sByQcqShTMUnC+70N99EBZayPoYEy0d
Lcb9W+bejKxpO/Rcr0jNCDHx4mzCeir7+d6CLEXxPW7EqQcl/g9IQWSmICYPnZqfe8ZtMKL4N9EA
uPFLe2vm5Zdj8yCwH556gZa61uA4tBWnNLru1DjDxpNR8bQgTfDD057eJngmLyfc7zLLIxC/yJXc
lz6qS+qkFK5/IV0H8TY5Poy2kOtjpf4zF/THtQoJ451AV7yAIuXGs3Lgb+Cy+LLgjcy/4Zq3y1PS
F3rrxbv8Qjg/dXNlr1QhkaltYCc4ix0ZysktJQnpwgQml0zV+KUcRZbUcE7sMdfO3KjcE/XSv/rV
QPy5ZDCjkD0DhTHR6/H7b646UnjVv8CYPw5EQlsvRuF2BiGaurI3AbWgLSpas7Z/hvuSSKY7TaEd
0l5FXwUPjpULlES7LXeVHOKFPK+UwXkOkL42K1m04qldEkGc+SBU5XPXtBBq1GE2RC1uaB1ywrM8
cRpPh0xZspdsSEiySrau1Do/klRKF0CAbZ1cCR7HsWSNkWbiKtubjtmYPIiQf1zklkGKe4hhvEzG
bwYBiSFeGl26P8ksey6CQBQTweMwSozoLmyBtv8ELGWZ5UBSN6UNxuhXpCRCtJDu8ADk2Gfooztv
SCIt13OqjsgH3eatBvkX2nvTMIedxtXEhDDOofoEJkfEaNnZdcH37+OQDGsxtg+bS6mYTLkMFJQr
FQQbthQjXVRqzUArmCEKmkSdReOdsOYxYwfkCGQOJo2s3/hDE6nsDvlotZ+i5FH+gHeIwMuWFRcN
xN/Bnyvuxgn/FBVLrv1EkcgFb+DBAbrFRkPc+mmV291Om2QB/qhdz6RIRm5gTIRs46ImKk3rdjtc
MJaDTzWEkJ8xRXGT2F2gKTicPeBka6UwR5PCDNFaM1mfbmYmvFyVUqCOGyUP6ljdjQ58sT8/mReg
gyHEETC2vYF11MZGsOvwjdC5C02MFuJSgIo9mUg812y8Z5hcrmQcbKsi4+SQWb6aZLAeEfiyyLrj
arS1TmY5LPXCE9OaBp8GDKRYhY1ifsCuM/lffjTPWMydMbvJqJv9FOaBUw6dcy644FuMsEHPLVAw
pU+iNBxqZBD0FPWGHVCQHXFe12L5P56DGonH9X/hvuuvsjQjc+4DHAY56b1sZnLTLCXsaC4mEj2D
YpTNKkm0UjO0RQdHyJqK8KfZQZaSB77aYWfjUaK60uMh3R0D86Jand4+cpwqtRBi7BcBNEBZLJu7
t4z3DnRxKboAIWd0oyQ8itObNvUm6APw6wXOabFQq+UHwA25nHUIJ0UyuMPENoTqjAajj9HTrxUY
QSMaEJO0wELgxAPbR1QJgjI8JFevCyeMCIdwtNmh1+zq3Xpb8pqCTsCFHsDKRkNTLDKjbIOXUOJJ
v/z/k2HBnTZVqEcQhUEctIgjrIb3DQy5Zq0cMFDCETm6wkBo8PHv4le4f/ULx0/5714zoj+5l7sU
bpJvZTe8rbmrpKOvBcTm42Eze9SUlNOFj39o3/Gggi8nrsUO65epc+eHWdSEcMk7AYXwsFomQQuj
SGL0xTt5PLuW6ao+cSv+Y9NqU+0woSXCloflEX6UhIn+ctZ5enuF3sTzFRi86KUltl5QtO+20sem
NLrz0KLPjbw5ZJL5s/HTiSVK7uqCumFNxRrjTMYBYrQOhzhtvvm27RzYnSx9uZw2tQvzaQ1XwVlX
X3FYPTwCVXxeOWEsRuCYmQkUUL6z7FQGO/YubG+loxDMsEH7V4lJQPV6HOwqugNvJAsdEQ7NAzGp
k0viyAMnzsNx35L1XHXgJqm8G24Hnz/hrOZSm8G2FIay4amns6vaJ/IKyD246CDwJNd8NGWPCbPp
ZjOgalNpaWaHDud6KqQfA4QSreCk4+K5rBKY1zjVy+RZ0GuiYO6EbVHBu7O7/+y3LTbwRgd3K7cQ
TkeR6pFUWeoDswi0GFPAPY3/cQUK4xqDFGPhPpD2QBYdQsm6Y+tbmyJ7XK+vYbuhDDa5kUfaiqWq
Y9h0KebUQRj6EhBpS3ayHXLYNENJGGY21a5KAl8P3urtyYQ97pMIOwHgfTrktYVwEaJVhvNO7Bgy
mwPb/u8b07FpHyPC6+htXL16np/UPL4y/2kN8PFxs9TMDcK97vpCbbQTcfCu8Gc3Q/eyJBiuJ3di
X0bjFaPg3W1Wa3ZHTVUI264X1KBYzRTHbkIh9buiZsfMgi0e3hFgkon2cP5lmCAFVS01vLqQ2c8I
l7B9cvdHYTURkE+XNPMVt8m+YfMjZC3qJwkCF2Jeeskv/euvOW3f0sK62+eBhmn1efwQCOgMy+sy
4lGKr5LjrOlb+7MTF07NnLIt4DRvKYauFDXkRpvNjpmZ2sbp2CNhsHScPYrqu4LFm0T3CXfUhIBv
Se9fcxIHfUjMHzCIUnX7QjDi2RedhrJrALJ6/mZ7NdDYA0ilGovgEgRWi7RHPZkqYxVtfIOpOdnq
jo4nyOeaX/u+yE82pqpeSplZ4XCoCS3Wjukfy6iHAHVK7OfFc5pjfNrOrwG5kKPqgB2d1Ypu/q0l
gFBX1WZJkOSX3DCFmg+PiEHNURVh0Qe78Ws1NkZOOg8jvip0VZLcBg5g1clXme6NOHmHvLy1Bxty
wAftAD4HW5lKbhMaty8I+9pOChCbRJpwomskLwKNrIO5vIrua/3dTfpa2+g/OYp3PZcXqA2HtabJ
HuMlJAGIKwDwPNvQCQ5njsNCuk9VwR0lhC3eh/r/rHmhY9Wpr9P3ErWoznjwrssYdFua62UwBRcF
K+zQRWPKCg30Ub7sndL24WC3pPX0kVMJ/H4d2eUdseWHd0o6P1AyNc09aoZXDC+qdpWsdYC7+U1K
3azEp1ZRRVOnEkvg65Zege0iGA8IrRoE8FMjT3vqAkVgizHZdNM7LLZln+TZQHoZp9YoOQWLrk+1
jhM3is9Wa2yGGoE3Tuo+sYlepGNefJeUR/t7y7JensxJHqdoufYTsA2oKJPu1qffUjxSQrvglOCR
n09qfCMuavixA87EY8pJDgE1fJ/wucUFN5j+Qbizova8HAtQk4O8E4HRWBUlLL3dPySQ9rnSQ/+8
nL98CEWlmR7sNaLv3vpOcuK4Wq5SPIfZX6eyTWCoKPZwZ5FensHqAF2fFOfjaVcRVoVtzjgneWpD
Th+ewiQu7GJuAWOX562GCy3ipzO9iMewKse35JxQpCLrnTex1ytjAPR8tZMIkAS30qKzYkudzpMf
9a6B6z51047KvAZMue7X1Jn1jg0/IUXa3e81Qz+8utplN9VSVKqOqYrKvFJ9mhG7e6sPOK1D8vhY
T8/nVXC7VH5SBlTbWpriuAd12x2+o3V/oTC2tbp48OHVaxLT7Avvx44g2C/bL8X3NihedrYeOxJw
TJT+jLZGhtRgk2WK6ZvtbxnT7fRv5CpoeuyWcts1RZOpEaHDWxZGixY4PLAOv0wJSK7rrSPC59bz
bUEuiOsPB62IzDgIhCqeiEnXHIHNPUxYT23/op8Xbf+oNDUkYLliyhrq1jo+vp0SlClnkzS6vHPh
acm3F9lPZdQANC9f755IMRaznbh4cH95oDH1hx14c7PcP377C2RItMtcx8UMBnpgPY/uqBV0HZdH
H437jus9bWOVQi03Vbqpxb1hNr3l3A5ft99V76GKyB5CL3IbyMWP4D77JGB1Mnavp2sWh2yND20f
Y85On4G+tf4Jr+dnPfCsDuWRPpVZVKeh1CaQmVIrDDC7ThNh8koR1UnhAKy1p5dOfrED+w5mnFsP
YRoY0igT8xFvvQYbF0nz5WrCuerpl9o8k6yYkLca04K/9XTNNU937IFGzW9a4tlgK7CBWmg5ALev
s5YObAFGGXuZbCHPg92fK1G4N1EEOa3p4JYW27GDfFXDoel5ckI5AW9YKD1dfZvEPztuqGp7P7xj
9WCh2BWJ6kkSs/jezDZ9QqN5Urd8x9vLQwhrHsqfWnRgjerbmwnnnY6DlG4ieO/+RZFk/OmK8BtQ
xhuWSjvcW6jvpQGfOMS6kVNVwafJeTJRpoUgABgNoT0vvw4bAgnW8UC9wo4Qh0nX10pKsnc2pDH9
2cpQmKX9rPfkwORX3oReG9PtIrKje7ecEPjjgLXNfS6HcUuXA1LNCKrXAGhRDhkPHJyYBJwxkaLz
cYCzWraF1iRYKVQ1MSqxSrT88cxXB46xtHpuBBGxYvRFPmyKmhBBZQ/rKD60VRlCPGlXM9LFnxRU
ib8YLD8J1iMV7HJoclwVmgnh+Rlpd6z8q0PDcBmS/KxNiCMsVXOJ/k8U/PM0bOqWZeVqm47vdYVP
fn2lZ7jmXv5q/SD+Pe4iaJOhBKd1o/HkmIL1r5b+JCTERYJpO931E5RipzpCWOkUhQJXCJqzuQvu
X+ziX1yFhIiKjMqCUqgUQTQ9TZ4LDISEx5YIbwH3i6MCXcJZxhhKiuJ2Ij+Q5b71Vd32Vl1jpnnj
J7QgKfkE73v4qWNBP4tnzirYzUFJCpi/h/2mjwf4rC8WUn96ipvO1isJhYfoQ2IRza8y8boH8B6m
Crh4GeemNa8KPvehTt5HWnBzXBXfZR5CDolpJ5noMb5bo7JlP4wGPM15Qp93qa6K89XSyfCV3b2i
CHCugpGhXYnTC5wIYB52D4FdhBSMv6n9ayWkOEu8zViGjxmNkaA60u8A+vnt/FO4XKCChmPwX5nR
NSzUcA8gq0Zv3z+cGOeynxXzLrWmYH1sov+wNtDRAwDxE5eY7E1unrCp6g46cbXPPC53TPRXUZxO
kXuIhEA+RIC1hiIyzXI8BXrlLn/djczYz/eJInE8ouzAyKp7i+2Mkxx0kxtobYHwsg3KZk+H2Ci/
T0eXBQWNWy15o7VeMe0rf9f2w34bZR7ajKUkDRoXrz3A48MJ4x0siSsB5AAbZtDjTubpP6VerG/k
c8AxdDNGUHboYhePTq5isvD8pX9xv3u7wwPu8fO52oB/Uqqg7Be5zpxu++DnIydtiDAdMDsauBYB
t7kCZ5Qti1tSJnCHBEuBs9jDOA5S3d99ko6mid7wNbw5S99U2e8LDT0uvE9aG3ZFZClnGskqAn5O
T6cBC/5TLXzc92s0NSfG+g1J9fsj7oeNU0YmMD2mUTLxQemAZOxvs2cvrUu81J3dQYLoDFmdn8Rq
PnTiDQm7nij5vbJGDm/BRUcQlYM26MhIwqGvoRZV1Iu9nqt3aQJ78fy/HmDDkDyLj4/bbI2gWg+Z
UwHlhzvkmbSt823cj9ZYAP3EKLc//r6xk9l2yIH7rbVz21Ap9754oIj8j8MCFxaff2NfMuNvfOoK
QxfK+xYJujlZs3pKfeJbwhvLLzTpfZG7r9jJRdcovnBPjF+9ad9SUI4eE58onGuerehvOmjkcAst
rTB38W2vsGLtjbTwoejtm6gqkADXX81go3j9nT+jFRi1DWJWQIkBlKEd4F6JUj9eG1FjpDGcSEtK
YFgnCKkvc6lwmtxxFjR2ewjmndQmPxdcY+GSy2Jwhuoz9omQ0WJtwAtVdhaPpnaDxGJrsBkrquZu
PnoMKtFSzlmPJsHtGfk5C3yr3x+6RSzjcOV+lZkIml7rEyqkrQw5014LNVW4CHHX8iL7RDSb8Uzd
lxLLWLNCBYWlktittn717A9o4dEst4e2/mD1/zeuX6KSbX0Pkp8Qnobc9LuaGkP2/YIjQqrBPLEx
l5mJFIDkFpVHnLTJE1XILXkGHzBj67w9WFz8P0pgsKse8fHfx8odl8Nu6Bm62897lTGXjyCTfhUd
Jw3OuvH1e/5AKnD8UeqO+6tvywwrtxp1lBwyRI5/f3yISvolu+2aoN4gK2p9OLObYUDcEmhV5Dhx
J37AuREOSBQSrddwjARU8eXLYl2UFudbITDLmJS+H/7IdnYrGR51f4K3BMh1DPNpVt5tppfLNDuq
3jUVhtxWqaQmuhxw5CU4Ux/NMs7/NyXFRyw3nawTcVuYY0e/ZhqQhO6XGckmDtKACD2/I8bSd99/
qrFJh+vlMWynlROvRVIq/8DQlPzAf/3C7E0CxS9WR5eosFyYw+seJyCz18SfPrU2rXnRPG6EEcYu
0gB15DOAiCvmOna9YH4/34f2W1t7bHsS4UGagaLLqBw/wOq/Ms/EOpID9MR+93p8gs/r1I0nbMHU
HyHIVjEm6BNl2FJaZKZsnq4Totb9H5DIqDYvIS3IBhbybraCCkX6nDkw9susTsblDLW+pUCtnUva
5KzvTQZ9107PMwXnkvcgFmhke2eSurWwG2AGzFQ9VaTwzYyZbxqEidqPlt4xGQWP95OSC5C2TawJ
yJpbm90DBfZg9C50WWonqLzueBYk5YLFbbhc3pTjhab5oYuqGtV8sSWT+HWKqJN+rg41HLPNaBzb
OlKgGi7rNaeOkQoBYieQkZsZS1/0tEcPACEyxw2YBoycjtF8y5XIAOeq8gC3d0hflZYW/p3xozQ0
/Jq1t0l/+M2uTwvtfKqu6Bd5DY//dtAAGW0qw2F2uzEbD7SzXqBFZTd11E0e2GtPntjp7p3J1s50
CaF3894ajnI2JCPc5Bb3vI/kgwNVpTIFi2ZwviMo1g8d3BrENlzXzGIEbl5Luy3rGpdumzMJzF7L
9ZNVC5PVRIsfbtARXrX05KQcRsR0muzIuG9zMMzU6xnCa4p9W6WoSHDXOq42KCwzfvmyAQ2FlvwU
JB/x29DutpBS0ySiucsWB1flzLZKVVs/XZZ3Hxt6cTDqMbwQ0qo42yKeSCgejH9fVeuJ8qkAF3WE
nqcX3C8x2FbI1Mu/JFmTdEs1lQm2rTUrEMrfNjbzx5JFNLmH327qeTT/D+3YAIBZuzhqb5t1X3FF
onXnzKJ9Y2UQQm+RYLJHpbD6FhUIclpdOtYXhkInJ9h2lx7UxMA9NFhx+KxlAKdpltxBPOAnTcuk
lRfXRZYD40GS6SYsEJv8kH1iqhRMQ/UuF5tNVK2mc9WcZLRC++OCOBsKHRrIkCw5sZW7OINBrxMv
x2IPllccqbckiuvnpgKSZoP619xoJh4Qy2RgQUgpvEQhIeWPEXBl4HQ+vpRrjVvMRQ20++dQcRU6
g1iJ6QRFJKnAEcIetMSamdorkPOoD+01HC7Qy3idQJjMXAYNlqPs42o8XerXKmJfYLQXJpIbQpgK
8Dx1DzsbYzrTz8rVXpeUZ34CY3hzW9s/EiP5wrnrK1IPINCCrkshAwY759+Sa4wpJEoA98LaI8GS
TXBseTkz47ZC+u4Q1DS4fYQA6CLfENv4JbrgL/BEOZXiKoRv5wH5TJS0cAifyhf05xB3eVMNA8ba
ARvsbKCcSWcwlGWNLnTidQkhJS+QjJ7uSuk1dgT7m9vWxrcjxuZ70taQLvpyyvVPU3Q1kjVX4y8A
RoQtP/WZ1NYyd4Fd3oXS6r+GHx0uML723V583vw/K7waA5CixB3CrZ7gvU4Xs4HY4DcjMccm12pF
xHYupRRYpZKFPwVCrB+w2ihkIQbAsvI11WW9hv41Iq5PrsZ7SHaGhhusyBHV2ihBMg/ytkmcsDn3
onpp7JbPZglD0sWNO7moVPnX1Ecmv7prw9Xb0fnPaC/OO//Or8mhmDGiBMjrg0K44X2l4FolK00e
XAYPq7un+a17FAwlx09mtQEkC5tbX7luSvaaMjTTt8YVJ4JEbYlUDN+Oq1i4IQyRgaJ/zQ0wZBxw
8oqtg8qPDoil3JNOuHrXY3eP6be9Fmu62p+X8P98RsBYvTwcYGqhryDsroruHV+GOxGgVVDJdcuW
WuaR7N8tHtfoVhpFe34AVzV1l/uEj5HdDD+Wd6n+IhxlTlP5eqv+Ppb5wBtg/2L/YKBDyNYXj9BI
7Zf0VA4atM5ZO7jPw4IGb+J3OAv9TB9LrAG8bmREvvAdgloW4i/P9znASIy153BZ9GaNnpAph+ZL
ysXkGD6gDr4A5/Q8C7Ag/ZHflRWtnnn4TsmfTwQO0ZLh9R3/yj8Wyam4B4AnYuDW0pP8KrIM6ndW
3TNMJyKXWD6mV4WYFMi5cQsqxaw0dtP5wM4NGuX2xaPXk8GoP85Gdxaa61xBqoAWxsu8IUKByHqo
mFdjhDtJz2TkjbVlKygda/o5L07Pfm5llU8jj874zTckynlI1EUbt76LmwtWmBxb8Jw1jP+2E3fY
jvOyout8pzBTJUgwnuxODPkoTS5+0qS5a4sxmIECSz1+ekFAifqA+lKMXEahHy1xJxrV7hhWkFut
nWCZ8mUpY4UV//ZDy/rHATy6WxZMxvL8aFMF3EjtMkV8OQGibvXsj4+UrjauG66Kbd2azkOHhxoP
a+mBhs+a5h5q6JvsDgPFA95xguvVyX54tbDReORH38oEOH+vaEAHBaRPl7x30AdV8X2Q3pG80s1U
1qRFSIpzATC68dzwaPmI1GzXEZB5EmoTett9iWDWTFxzFFNtB5z4AvT1CMHh1emdRX/Xb3tBtQc2
Li9z3rhd9ftsza9Olg8PPB527Vb6ucczstvb/Ag2g6jm1HUVvoFdHW/wckzh+0RZnT8aiEzgZmsG
s00vvBHnFtsVOlm0zl0feyrXKD9QFc9LaISw8dwcmVuPTtjvm4Ebd0TTfPnBzC61kMQ4qJaKz1iz
lJwxJyaglZdbTnM0HEvlfpElhxTvRGegZKlu1MBk6Ng0wwGS4dq3URX3UQEdFPz3t5b2KeoaGm2S
q3Tl7HEoJVBe2RPtuTWn+6rUQXCp6JtzrK+8dPto1ipdOvP+RKhUhVqBHpzjBFGpj8g/O89gofGW
ZpRji9anUm9FvKHgSWTwTCi5Chwo2cGkmCoCK8eKUUU2CNA7g8X7WOnilmKjpwNom86iVon7fi0A
z7qrkCSbDDj4otcUrxNIvbdCcwSyjJSwIPctsszKzvZ+6MEm2qqi/XX1iDJ5KKbVwPw+IKe2LTDT
DR7wYQTTeOACR+iG6pknmV/n5erXELtelqEKW2r2YeB6I1dKx/CBYb4YdLnnM2aY8lQgEuoiIL6Z
uWO19wZgPIjpW08S6HowwMgrKFUj++5Ys05fF/J8v5f3myA1wf3IT8wN5wXEZRnQtANzscnVHtVf
5Y8vxFksJr1Ufc9pZAI/+OyEkaFc8VcUtZ8e3OZkL8uvsamRxF8/gs+z1jyCJ+gielRwjxeSrpUO
y4rVviRcDtr9Jyue2pVLEbOTl0CDejgbHiiX4033Tjs9jorvdKexsOupCax+6Jg+VJ6LhHups7RG
OqgmkRgPV+XRwV6F5TPpDCoFMeay8P8Vue6hNt3ioafHqjlLi0FPFtMz3cfM830t1DAg+YGji+ei
MqY5BLj2IzjgfXpNZlSfSs7s86HjakBLCtp/q9lSaS0b8yH5U5wIOkTpdpOdwNzfeYwzGPOLnlT7
hWHgjyN9lP61l7mc25kIhl9rCjUx2g9bOZGNZ8H/SqAiSKNTyIifZyEq+n1ANtztGXL74A/viyzX
BzZhCI0+FbtBHUvgRw5MWNaDMN9SFAfhNk6NfJ6p0JXqD803/C09inEG0k+1M8MSNPSsVWEvM4KT
Z98ts+YgdCq9anydUjpBxWRc+Hk6rr1BEG1C5d6uZlB7ebdt6bvywJnEwCwF/eH4GvdaNjGvw8wD
p4WXbJs9nrf6pKpGlYzNOvz08ywFXMB7mIYEU5tK66GjEPWX4q23GbdVcqvdsZCLQ6PpDJyGLlAn
PTW2ZnO+K4SQY6jovPg5GFQALTeSOAwVDt+JAm1milKPriYFpAbJ4wi20kHChrzcMBVjlRudRN5T
4em8jFT14RGulP+hp9hm+wiXuQv1CeSvHVpl2Ca+NIkRMSdYnCNqm7k0UTZymPE0EX3Zr5KeAKW1
hhiOBrUtPKcUPajhhVOK1CYZJnSajCPV80N/mLTJAPTb1iJvADg0J+kzY9oW+rSNrXWZ8E9C4yGe
Lh1PdhF2j0FYEYdfhdFY0FFI/vad8iwjfY5Sda90Y2ueKizRFIlXBc9LBkuzEkipdmCrgdBuDsJP
qseFMDmgzGSIoX5Uom6fUNAtGfXXTvscyalY5GPqy2VD9/L7CqkC91WW476M+30IxM6RofwL+UWo
C6xdcSbSGPYUT+qVGpXbjZkaf0YbYpujK8Ka08h533IfZOdivSNTbJlW3ObyNwSy1+uN1VTiqnHV
HV9cEhztYgMD2JvvL6+PXPEoBwByL+I8TLAREoPY3YXOKq5FKKxpYvpWx7h5Y4fHw9DWd0xdVY+U
d0BVzt2NOdtLpyZLQlYf0y5zQSnFamSwqaZKDziJY+1TjqQQJxtoYREI7/fBknE81En4OL/wymCK
aj3tAky1Xqa5631CJFJn4RDWps5Vj0n96HI5TuHbperiBI9F2ytQjadUdyBMDMfNEzLDElkpgGN5
X8OkyvVn1pp6LvVaHDTN/4QPs6abmBwVbGC6fmNfavh1xUUfTBlB2kThSg5NYCdlwkZMO9IAaHxy
KwYEM4e0FUKHT9hN8KwGH4T62BKRgtBU91jxmwZukz1MGAfNnqf2mbKu0d9PeVD8s23xZN/Mwy+R
6PvzBq0TZVwAkxZhQkrQGESevuutA+h6KRthiB6EqxPzYChyzr/6TpM26XySjOtzCnsyMNj7UKpP
ICpAZnFRJioo0SpbS7Nyo17XNxwf72mGA8VYWIAtbWdifNonBagmik77rePLPI0UvVDVUVPYDb4p
xkQugEhu6i/zPa08AsTacY76fcpsO/KQj6n2I2dBuIlMMTKguZ/X6WLbuMLYy17aN53jxicpSYLM
ipZkZ7Th6qZy3Pqh7rHXAV0SZdAYXdxgCBBVbdDvRZBcAWhGThOUB+3Stwm49F4tgzROPlg74PSt
ntQMB6ftFATJADLM2WOWU9L0uHfCqEIGJ3ixtrr1JxvOsG4IZdoYUImuUMXm3whEpc2mm0SZJXhU
fHpPPlh+lSqJ+O8I8BoyikUw3G8oqKkKDu6eQjYFHbraxH3BVAXqIT+fu24+ylp+LlF1FyhvGAzh
ua2JPHGy2DkqsZ3ucUEbVPcUxu+L8M+tyUQgz3iHk1/PpkX9nGqvoRw29lh7vBxHhgNFgKBUXiC3
p8eomJDgUGAF+l21zLciLA63zpVEHvX8t9R9ybFS/K9/uruGbwHRNJR73N+7VJG83oEcl1oM7f9U
A1huIj5SJd9dL6WV6p/TDETAlHl1Bx0KLQRieK3JzzYrSt68mLnq4UxSnn2pUvZ12T707tU4WSxt
1NaZaW+T6EAusExFwYcgRNNlV85KtM3ITZYUVTplmzw1Ova0rD0uPL5iprW6+yb3l4g6r2UsS3Cm
NWK+VfO8cWIUoGAA0olBa3QAmZrhYCGkTjQivjySmoZ/QckPfgHJY5M9qx5xtOQ6aGNk/TTJMwNQ
R9Zxcj4uMmPVzYIuq4/j4nOF73kb6OG2aE8bo4jRSEUW7/g1ym8TIMzZMjRzmf33NlqbU2ZPQ7A2
8qgQc0J/Gkqb2zlIO2Y9FfHTRD+7eDqOizLq6W8r0MGdpfSUnNFkkkjF8A4KKREihWYZ1J2ACscG
D7cR0DRqqwdDqL8XKjggHIalwoO6QgstRf0IOLoy1LTR8JM3PZV99tbrQ/5iZO/o9Wl7IGGeaOx4
1UuLX7oegsCm1YI+kL9UAYYTM5OCHShL2JrDcPVpAXCLBNU+vGjwyXsslWwJBpZycfkYgpnzeVs1
S1xfJa7lCSZ3Ulp1yzze3tviQiJDCAEigWEdhVnE2TffMG2ScSu6EGX9dw6FXBelI56BZ+b3sGRD
+3yFR9Oxk4mIQGvog8b7bSlQUaGrI2BnEEAkPpHWHzpJHGuTV2XQ2Zyf9bZ9hdXeOlirBAdIf3bp
KqOhOQK5ozcd/iY0HT6QegLukrDL9znDnIXmo2LxwjAFv5BqnieO2jsbgsyc85PJXwz/po6kno9y
7/INbj0TxM26JWxik01XOlU37VnYQep6LnrmULD617T/IiANyZXx8SyVktFOn4VMtigqk/aUoopr
wzloHDpgtNIlMxcue7HOFEC+rtboFrrwb8B3e/DFmaY3/QKLBlbmYva6cOFGZQfXdyfbuKHggSnM
4KxM7mq8yT8Oz5gYFkeaTLHpRyfkZ/XCbdD6m25mm3pl1Jia8/t2Jfld5/jYCZJYA2XaN0PAbULn
8pZ17wO5iHr9JYgAUuEMjPZWL3RGS477GN7WeNp39xtl5kQ2CRgmnfCEeWA78Ykfuh64q3+gQdq8
sytGlAscTF1ZcwSHt2c2ESz+A1eR+8hK2nWNVzEY3x8jmj0VUNepUDV8NQgTacfvAX5J7KOZEryX
6iqEvrm6w0LS0rwWY/Djqqv+x5yqW5WoZQk1zfcJIxXn909rD8DppE/By32wE/p45ZHm8hTizmRW
gi6y/qMxfBIhoBO0PnIC7bqnMpSx2vnmw6daLj1ms0i13KyigMdjTp+poyBisZrJ1I7dwf0cNVh2
L2B9nVZEEdM65IdM3wWCJFJeLTfVxoWfanFwzLj6O50Az+g1aGdxpf3D2c+VNpb3lWTGyTu4u6j7
c6U4RGW7HwnxI7eK/lcHa/uVhvoA3cWcYUyTd6DXz6XXv0rioyDArmGx7dVPZ48fjBRzXH70QXxv
66zTwB9rtvhuo+JhrOWdMZC208ooEBuR4M+iky9z64SVncmSKXJQkuDCvx2aJJVSWrRxhtbcOkRZ
sc37n/6EbcC1ofEYhHfLHp9clUoSaL0zz3piRc3PMsDAOtCwNqbQUK6QudjWGBD+k+44Hr/ceCyN
hDyYn2WQRXjCAPIQ9Ddoz9wGxu6XgDjtmfUaMtqLrV/dBWcOiOCgUVhFxR1FkKsSXQtb+suwtOL2
0pRsQ42LCn9gvUX1BqePQQBPqOAU6t1tRj2tmT6kALuzn6SFJaRRN5Bd2XnAg+8dCMEaM4415RUJ
BF9n/tsqoJJ2/ikf6V86UZM16Y7Fvx6DhiDquENFauQA2xw+CVjfZqtsMoRtYEpL1BHonB7XcQTW
WlZ37ebXArvPRbFmlmzh2dLRVA9aQvkWcyxEdTmLwrsVL1hv6YZsWy63rnWBVrLcj02W5s8ARllf
mjZsDPy3bkXW9Ft5IU4RVIG+n91mVe24vNtG7STjv8fywx3RbyymQaCWyAw/qGoMCip3817WLZna
ZoQPRQ133PBSoAQUb37btoLeJZQdyB1Fhq25qr6m8A7HNcthBkzQK39Ho9ErRD2VxIlvB7/FyCp4
yKsNJiOSLmt7gKGxZhn/tNRr4Jl0zPM20tQmheoVvH1Wc/fUv/iZNXiwEbdQIIWOtf8vbrORjdE3
WKdfM6VEC4XaufGkr9IXxQN3iZTUutX9X0flPdtXY+6k1rDFg7h6fduT2g817WjlfuALfNWBa9zw
cEFlscOJrHeuaJyhmm8O0CMWWha60cSTqI+48elZzTJ+j0F+5z7DWwR6l/dBqv/lWJaaUrn2/SFi
I+GBo5unTK70EhKZb46rHEXnt9VIifv6SSv7OIm8cJeXI2z2K87PKRN5rOCiwK1yLstD5ymVPOSz
pi8lSbg9UucvyJtUt4ryGn/cPbgGtN4CQtiHavR2W7tpf8Bx0UOYqjuwtsQNOp/Pq1mE1/JvQgYy
DUUOB0L2bYixWZrjjSvsa7iGb9nc5r9ok/359FYs2w1Jtroy2YK8Ov4JMh1om+cTHSLive/OoUVg
Cou0fDApG8NlDHWj3JnxGSOAWKx3Ps6oT5lDnvhkwVCFyWJ9wE9Ixf00gbVag2qgJ2NRpvLXk7z0
NtLtbovdMXN2yLqNqm9pi6hzZLyd5Vo6eBJrnIJm4LO6GIQXT6ozdgeIiB9xiIwPT5vFNFHfUtPN
JKIjDq2Xt/Sz7nS6jUHHpIubPpui2RhYg4pRzOKHrv3B/a311gLxn+RfHEOEGsgBFqG9PwHdysgG
KmEbEqr/70lb5E0i/COZQyXwjiHUTRVc/K1/p3WxD1x2GlBCAEWxPFzAX6Bie/T8jIcuX2EiwJfN
FPX7iVXxUg/Zw4UZGRjuisHO3ipDSYypEfQyTo8ma8ACRhJI3Bg4jF5lpqrp5vvwRQSfB6OWrL0L
XNb0KKqRMDKk+dpLPI0fGOEITcDLUFn1oFmtFjgD1+CzIrJL98J8ComasLsPr8h3AgKCpZ9h4m7A
R45Uof29t0pD7VlBLQ49H+QaleXJ+rqK0Hdsv02QD2rn82ieTfxukIuEE6+VAv8JbqVkRg0TRC6q
PLSnRj/RmijnihjMn70YXwNeYCMieblTqQ1dZX/NPs6WIDgIapc1PMGxhipSJfTstPABFqBtFuAK
rqA2gCtQPtmtnxqGzubFmjiZF295bPBwFKZsL4WxUH5VcAAvDMtAkVphjSO2MXCTVnHaVjDsqu/u
dMS34LkDzwxTenQYKuMZS9SyO/GuXssl9awn5AimQzEHB5+q3IsXxAJYACz9kfMj3upPHXeSzxnO
OdTK0VOvFHd7ZXVlKEiA3KCWvawGQCR4gxEQQ9by2OtDTs3HZb2byi0NUW88dxX2PRA4EeC8N6b8
EyZZ63d2iMelERjeIsaUrdalF/saj5qH+j3WbckQbXohJedArW4bgWmbSMjC+sXLtIQiUBIeznOQ
KL62C6o0EXeqVBmo35XvSIJAadiwcxf+1uk0mVlfeTpN7Iwb/vjwIRd//rUFR0i1nc1tNohm5vCZ
VGx9TCqVhftMXYN13YQFTP+iCwG45EYxS3M9y10sDSj5qC9yfsxMHUEyk8PT+coQ3oeXv/zx70lG
wFbOHH2Bb3mSi5RsikCaLbNfW2WC0wvxOG8mB0ZGZ56oVy0tMNiBhZnhH7dcdmUWw+72nqorYa1j
ItsyA6+pfkC1/SdDg4X4dII9ey5DBe6YQaNlvIcHkKgTX4HaOFUqMHBmD3dmsSmOck3d7NVY85Mn
90X+iSN3+qaBIM6/BECiNKeGH0Dx/aRMe1XLk5Qas5stxurN1tgpYgJ8gq2iK7aDmR0GLgmxxWdO
67/U9KcjDLjsO3DcQRqHKkqknOFCgjNp/RHbT8ILeW7axP8w2K9Qo4GvG1hvUBblyA1hPa2r0T8v
kPq9FA53LfwQ6EKKtXFHtZ8UTSBMWyYGYI9ZUszftsuv7jEVBfEzat4IlBAEmEyzCRji8HioAFKj
UIbrg1g24vE1yvMnTNzZKAcbDL4UUCJjmDmoVZoCX3qGk5AskVvjqQg6G0ISvqKER9lJ40vfnrUu
rb7OsOh5w8rKT1/cRWQAbOr2xhyGUfJ81FyxsRGSeF3AUHRRliBLoSrS0E+Db1aDC+rnaApReRor
P0oSeN+j4ofvQOX3GRhFW0zUdNPAOvIj5CAXA4U7XRnZ7dQapa6YiRnp1F4mQrVzS/7LKiEqwlmD
i50lMg+ve33K/t91tal3Xg6QniZNiRhQK4jvPLuiguZbw18hXEPi4dXJpZouaaGEVW5cmQLrOgQa
Ltt2bAzF694lrxtR177fS0EGV3ut7mw2lZBEnoZNP1Y6/KYLZdwAGOhHiYzzE+hbXO3Rtk132ljz
pCSoPqCTnaEdJEg/49nRdY8xy/6oyL/tUEFoTDzFGLCpGmZbXQwUxrvOWpml4iKKokdtPyu9IFkv
XxhTx6LT55TGalrotVSfv1qJz3qQw1WYH3x+tIXAQejgoMsYOUVnds5uDQmiHIEqT1yW25orsVQl
LC831JfJukottXS+x1hf72lJ0MChGQvNN0Dz2+SpnPiYXmZ1wvKUDXqynGMUObSRv3DC7HwYFUhH
J5FhRGprqbMJbVCJI/L3QG1Qj3rvabiahGfiwG153g8NGNyxXFcI5pLItf4g04IwPM/0B2inX0iH
WBXSbPi61Bp6fH2h8f7e1+rUMi8BvAuf1KPTMnL6EKxipUyR5lCH4VPsc5jV7XWGER1zMN/40Dsb
OLtCMT5H3ge4AKI8wNLopVTabWJ5CTpU1Da5biTLAiC10oeQL34pKUsg1oU5UlTiwYgm2Rdc53Zf
gjDN4zc+C6n85uR/Yrjr7sXUd8+TM38OSb78oK7xxCt/juEWce4MaN2wUizDZOS4qjL0WCDpfs6x
pqSbjID1VR8HnWbv0YpsdGbzCDygDRC90Mxkj72dl6owDk2N/JAA1lOB672PCwbu5QIqYqrm58sx
r4L9fSoVm78sLkfEY5tvASjeg5Hg9XPCR5USeFJyUpiW0Ars802D3yOcrfE4Jdrqks8lfkhZ9cSA
TKbVT08fwheNb7gp/xzhkVrNMHcWhsgYbEIsyjyssa8nTMKT4LgBnXVixYTVU9GcI3q6hCwXpcrm
rqM1PUzzes9M9zi/3aTKTa+wRf2S0EZs0RybYheQbE1YngpbqHWuMbILmsUaBaj6C8f5GyhA1t4G
VCQBK7zusNg4pEOq6ClFMnNzFmSNO+8R3bTUneLo258mwsiY2aXmuM3V62DSTNRkXHpjAcV0TPrW
Y93QB3qE5j0gu37p/RpXOwNQxSRGfoBVc1Rpcgsj4pA5XuajU9rFVwdp0eg5VKhXW/QJ/CHyCayh
fc0wTIVegLLxrlPBwuQWc4Sm9xO0SwBy51Lg+dqLfFP1lGctBqSyVJSW9L4x9ZQep4EFjLyJ/r/B
EEm1i2O8ueN8oN20ECZqsveYaaH+3JALzMU5hIi97qjET5spdc/iu3Tmqk2ahoMPaREsBYqnnjcX
aURUorZy+0j7Yq972KVWssNiSvtHpzNB0LAiYVyJjhyo1K0EnuEk89f2/6j49N1NN7YZtPD+jK3j
sRNfm7v8Jv1HU084xXgzOqnbZ/cJaYo1+fNaUmjLRHgaqDW3hfddtYhjKZuZGr8WIliabnNsFZbR
alAFiTSphaCHvprj7+dv11BdMX2YNmhp9SUKM7nn0k2Ulmyb/pzFgqqvfV2Y3KsFNfjINsLX711A
Y174A8HLNM2iamLgD5+zah4uS3DEvaNZTWDG9REBjH1jfgiax90usTAiVkE80SfNWkvCeBVyFYcI
k/xuTbZuLGwwLuqEHAr+UYoUVxKOpJGcFRcpueKCSj4Jzc0ousJAW3hapn6mbNw3jTrMZLSagOqU
atop7SSg1ACBmpWSHqSJC1VVaDmnyyL4A7snEHKb7I9jkUQAHbvpvooECjeUaT/CAKezSNAWbwXE
fPtlWtamsJU5Nn2f8WkS5ZdDLmtvLvhp1W9H9qbyWFGAojRycLCYAQEZ73AcrvUnqv1bHOR5r5AE
AeXYTGRlW15RpWNuSdNsA7KITEne/FyjNG5JLmjpeMhYOlDwvEaUnYbrc36txMVtOnTpRo4y4nuV
yhd86udRfRCKRtq7/e8bRN0dgTz8mbp+cG2BvqwWBJWFS+/HcNNNs0+Tw67Tvsh465YhaORiunWw
Lzc6/+oljrKfigWM3wqXBKzQftJNh9TWkeolCLnjVtWiLQq8fDEM4813MyzS6yrrKlUi5orkm+NI
W06fGUMwAUXsZtz0r7s1exZZcT+Ebvxl5apzjNqVjjCIyeDQYcu2QN/VPCrj7/wUH1c27c4ikdFS
05Yo8LGQnig4aDfxn6GhIobT0EBKizszYZRjiExCqsjoClkviRmz3lUnWCbpWvj4W0MlfPidcW9I
LPAj9d929QI2LKjnp+kK17glNnNREkMKIKfp3IbgY1Bo5Y/8SsWgBcURveu+NuxHKmSWeYtfqUna
2xJBjMr+qvXDGxYbA2AswteVfX8TRtBg5kHnFai2fnNwt76Fa9r3GX03BPBlvVTQyKFVqe1lWHyD
BJWcCyo7LikNWy6xOS9ch8OpDvV2oiRxzd34ua7jsPKzxTc7ndyhfRaJ9ko7+WK5e5F+0fMl8e1e
YdhJL1qLwrlsrIVbxQmRZduxGxdVY0H1nfsvzXDcyUXB5zwJUAj17fP1Rd40Jl8GTFCxw8S7J5nv
FB0N/Fvt52WcJtk7scFQAE/pna2/W7VsUTfrOkHrFFxfBsW5zWaNO74xkXBgm5YpGYkSMWbizDmf
HixZ139ufEa7aO9v+5L7PLIFeykKV+PhfCOPGK928+GYu7J0nQPw4Prp7MhzrDEvpsAJ2hTca3Yr
K8Wcu8zwavL/9B0Y0YVQYTVwOCzFERywTXG2YMzUUcDiLYX3EWgLGvcYEQYntkao3z2q58670cy+
qTKZK/7j36z/kgankqgn6gKK9FjTjdpfZw9oeDoqmdKGARgyJBhLXQKAXBUL6YecMhqERa8Ql0FO
N2ppS0VNQo97ZG3Sr2DrCl17RFVZ3xwlaZuegQQX1KcTOsimjLnlK6IVoRkCMmJZpQSoou4Tzq4v
mE4k+g7KF7fSuUc91xR+RAajMMe0a7dTWSHfkNFJudXXu6zxvItSSYcUrPCqkeg8zktHEvyxWFL4
0aRQeQCEu6aQy+kxniGK8dZDQiP+Yb6S163Vzss1XfqNF52+0QjDpweCUQyFA+Jwi8Eicsf/LcEG
oRJD0d8SNj6Mo7kzvLi4Vnj3FY0o6JyhGh2gftXWDRzJayR3XrMjrXEDDD5CP93iZjMDWypXKv1r
7+uI2jsyVhRm6FJeUWlQwYkl8GnCitzwIhjNKp3zTGegQ2zxyBJ5bz9YaMcG93ejabzNaR6F0W37
kAzhytFALHZkPKO1cokSGHHZeMtvPbpxQJHKc5mc54ZeCyhnh2YYI9WuqexX/rHmqcAsZH9JJLG5
Se+NeK+sc1MMqZ20ncxgq1UZbX8xTcdXLEd3LuNsu7m9QGR98cFwTaw7HTqaJb4kD/WjFGqTMewE
sc4f445C4w557XVDptuD0wq5PBuojN20aLYe6xFeR3O0HRBb8DRtpWKj1nvjsVoRdovM7KxSu8wg
Wtg8ZwEinpvMXnbJFthCaUI7dA3ctZCdvjG00iCdksd5S66vEVyJxf1mTKQ8DMCJSzg4FpQr1Po5
iZ/hgEKlCJyvP3iSOqKmShQHDK0f7cP+lr8M5Ok6N7lTa2P38VSicNcLAmepK0HxbATGtkI8YEjW
U27p4kgCW0quGpuCpSvNqXY3oHQhxfonxMwStmjfdJsJt+bw3Q40VQhu22yCea2uj5ymjl50Xa36
ZQ/A/PEbCXNeqfBIfT8K1nJ9Xph2QftXos2iD60AaDX5XsL5bF+tzJsy0SiaL3LcFj/WlseB80FD
0TY4UcPsFxsUgLCkWsd2SCnAd11uze+jFAzFdGXZBs+2skX0M8UvAKaCU5i/V+U9ituth0g/vQzI
hFnscy11KXmTUZWK5cEmQcO294/TwVpigV6YldxjwU5nGEjek1vnhde+oRqs0h/YkSQkApfFWAS5
rZeILVfHYH8rhBVqHsDCLpNMr/PXmh1k49K0k9GHmTd+37Qe1ae/JmergleCnEHEyqgDPAih0TGF
VneVo40SMQuLOI/zrxUHX9qoQEhyHlnUCNV4I+50Jetqbowp13Z/J/0TliPd0HyiPRk1CCB008GL
a+OTwYLAxiW4GcI9MIdOyJZquVIQW8PZZLSIquyihiqq+JHsMEsZvLIn4EPaLgqFcaNHvmPFBPiA
rVMtge47CzYJ0wOrd/EJ6UXxViXfkD8nvKxA+YLwIqa9lW3RF+Nyy+1bDUhT4RBunYmuDVP8Xt9E
Hd/ERa2sonxExNlZawIjsdHCJMARwkQjur8uWZhjemijqlzxDWV5+b/bjAmmGIo8VPQ1L3WPkZDo
RgTVTeraJe5d+LEr3Nui9S6tyBVLNofHJ7QQ4k18482jgVtSP1gqnw2/wb86OrFzO8CwjDLtXwEf
7uorYEl9VFM58tVsK2pcf8Vjb0iZTWjStbdAXHkh/2UMBUNh//WNW75gKDxPhFSz9CLlkBhAQghE
gaOAT8p99APDCwapCkbF7z7ZZJ0Uh30BckMm91nGIsZGm7J+wWNUCU7xFrz6cefl2VE9N8q69Fdp
3+mzGYi8LTAMsYfhjla7kEPf7oKTKnWbL+vWC4OqlocNzfdmGQkYQOaZRqMJK/TgJxRhrAJVlD9o
DruQrEXVFjo6UBSSKiWPQsQLveUzes+WiIIRSJk6fL2CeB0rkRHP59bQ0RPs8BSfR1ElDJkf54eH
npfdDcJO5+0pJ4V1kDlmk1frvGQ0kslPiUvc6gnEXqcIJuaFPW3O8QRIbkzBprkCsvQ1JWRq1YGp
Zn2POaaJmnm6P/q6Gc75u55wZu7eslTQQbM27d1ki9GVxiAI8r7+dxP8rfin1BqDjRU86+xLjbJc
FDKX27VKWWn2/ARAHfK337r/v+e3MWyp+W4JhHbJZ5Nw6Qp+kNzsWmqsnAJcQQJqQffpPEERL1RH
0gLoXkZIjng/vKnq6STkRuHXeF1/UuhuqpTs/q1KJrH0wlVbB8N/baDzakw+tiQWIGBZrpBlcHqP
/b3GYlOR/o9A2BhmsslEX0O1myxnmFAOVZGAjCFIAHjg+e6LJ+ZdJ1q/WdyVDZeXUJzHAHhS8dwl
nR94a1Jy80WM+nL2jPLr9uJ+fznoB3DAkkYAiJqM1qupVoiysUlgth7kzlUHu7MBoKSnYg1TFdOO
p+T4FVs4LfwanPPjCzMcVsNDvk66xxQMuWFC9HnEze0BhDmw3rfrr9wK+cO/8h9g/XJ/VhNZasHH
WKgUki4FQOLKl5MocdT8IFuWtmGt9CMdsYR7A7BKlDu8tBb96Afgbejf2/nRFZjj0xcvXMQjMV7z
LCEIkCrKxUlUkAtSJ0vi4L3tyO6LVDGf78QYQpJ4lG0Nv7bnXAY9sZtadAC3OLV4GZsz+M/XSCvW
o+7KUVGHIx4PnTN9t5+kRu1n1rbkZ7k3e3dD/elNLJZd10xTjCItaSlQhgY8Dw2wPjDfUPC1KsNL
IkeVB1KDMIXP2x0dErxiEeu/jTckpQuLCekRkmHAEtg356HSsyCZTpjFXkFXx+X2Zab01L3WNrEF
s2Y9n4ddWotngeHgkgKM3Du2DRZ64L0LD83bdeNEOr1XpIkrN3cdnI+eVDCqLOMN0QhLmYgNlU2i
riTjXRxRzl6rlv399WQouKnledkSbfajeg/hKzQIrvSwCJpJyZ3yuzFXj/bqKcHxkDlvLJ91yZ61
lQjDZ3aPhRwYvE8lkph3hLCeuc0Y0S46gVrX5pgv7A5IiyliUsp+5mvkWvwoXePFLMfB7pB4B3R3
t0RfvVp7my9CQfb/rTHCrp0ndNyJlGugiVLvDu1nTM2uo9UAX0n+oVadpHO5U5lvPQ3KrdtcirlJ
NWyPSmhd0bVkxwLzxnac3YkjwdFrSrEM99idZ5vfqogwFtN0HBnyczLQBOCzgeHRH+qknnX8a/C7
F3XpCbsFUwT7JVvsYVM7tNgHGc76WT2REDiqGHmw0QeocBUhCEt1flrk3LWk9gu9QTXeQp+RLNIa
7ChdHNbi2NeoNrw8ZMW6eMrC8NCDdG1zY5P0YlY+xZO0vmQAnH189JLhB88bdpnfBi4X3N7Cseg5
4uRS8KH+dRGcTpaZTjFT1YCA8yN9L6VKuISeob9VXkrYLEXHDBsz05zPQzvWmysTabYbIPa2Jv/7
VHj6d5vr3sfxn01njRP/gJDU4kwyQciWEghZa2prGN0zPx/MOJzPRaWayFAOMJcDNMdA1xNnnxTH
rnBjgFiSD0nHXbGPKCGETZAwywXarLLPJ5aN7GwK7hdDnHF8RcMslXpgxRGyRz8OTEql6Bvq8+Tp
p70RpP/lvMYz3PBY0VneG/L3gXu83KYULMLQawWbVkFcaVGOVmQ/eMYTzcdLLNAh0T51j7TSkkBB
W+Ua1d5AlCENjOiHgAdn3Ao6x/cqMELKI7Llsm4GKkL9xsgWruvD2ngc/nF4UCRxFVqwyyvTmqUD
YbHykPt45v+9mX4fD4O7yxO7jn+iKQ4JzBNGVEisTfxmEB+kkYDQ4F3cBuztfZPw3s2nwBr+tYL/
SJ7VzCBsGAkzbHG3DHeoYYwKmsTQKBID4I74Y5/v6n3QTkXqPCSTYtFhZdZ1wn95lkW5DI/L52Ma
ZNfJk4ETcCtOGKVgP8DAD94BvptKp2caNvR0/yOELsdk1+jSDoQh+1OMjC/JienO0SLsYLk4s1PG
xK6QxgQTHDn50FtGhsPvHMZv6ILyxhpEIxw79WV8Zlfw3ocG1GUggb49/4M6se/NiVj9IXMalcnx
xseTTkbQtT5m/uH4ZvacdU44qVzXSd/m4+hr6AE13GUeKBKwOssSbLzIce0f3Qa51ikqoVuCN+x7
Kv1+/v49nGCMFCvDWi6SQgI7IkqH2U2zfCa/ilaMOFVsvfZkovuijXWBFnHBmm5zikJgDJNoIsyR
xEmNFeGn0f0GsqB7sNp8x8CasZNxvX3HuYkuehtYm3Oz2I7su6bENIXSu15a47Nq/Wyp1pGI2CY3
pHxgvJ+nne64wzpQ4pg4mZOzYStHoJi50u9Xy9G0Z8gbAf7/yZMX5v2WYkMCMBHrPHUtPZKBsWU8
3scGPh8AugN3sd8NXHFrcGDpy2MqjF8jYJsGwOJAbTBGy6ArP59iC4C7nKgasG5/kK8rSqa4CIC5
Bu9PoV5cWsrhvADQoBaMP+RaXrPTfaf20x8A5RwF59bf7pFAwVE74HBSd0dRrHO4IGcR0rrzJhdR
0lUeWgcWFZKyWX49XYlLb/YdVLmxi/MjiacoEHm9XpDXtKM0eX+oVJFOTVehEbToeYOG1AeN2nl+
o3HqsH6DnUzIanZj+UN5WZLWGQFdIhI/MYYbivXvKD6rYTHtOLysK+7VM2y1z5WP/X5x7zADvr5I
pw96yP2s4GIcb/qJ+IMNUZFtXOtyIff7CxrVbP1cJHMf2BvvYySn7oThsWe4xVK1Oj6zBKzY7aRf
bBd7pFIJPCPODgWt0baM9PrxKHHSOHDEAEs1E9Huzq//0MZehR13X+2el665HecLoS+neoCKjReX
hem3jLPG0EYh/ACj3+1x1rYQ4/G3U9MA3Q/CkwMFlzOV9D5Q2IVmTQACCcdp0WBrmTDKpY7LGTiX
dgkGxuhKhrFjrlirYbejXuZCTf14mAqZlhdQu8uROO8oaOoIMAoaXv4+aw8jiEtbZAc8QX9JKbQI
ZYn3xOd/7DQeI4jYrz8sqVRGhw6L0lsBOUgzE5dqITjna2u39cUuhLwOE05CvUxnKeSHuXOzuGHB
52v2w/cd6VBITOcXdi8/5yc3fBz1uXQ7U8o0mg94IgTX0euZZEIIYNCy4BuOZgA4B5QVDpv0jack
9ds+npYRDRxSqm6EVRB3PFA350rcSvDhijl4dlfm28mO9hCCHex2ZKgR+k6uCVjSYt1LUl5EJG2v
9TA5MFcGVw2gnSw1Q2td4X/GcvtLukEwVvzzMpYAAingqDdFQoxKI+WtPr610f5r8eeUrvY5N+IC
yDr4HllNWar/wMVAls+riBgsniZlEXUqr/2WYXulhZroPxdZ9bd1tiFI5qrLRuIX7yPytw108qtC
7lfFi+QaEMZHtHPtjWZ7sJUJxTB6W84q0werqBUWjl9K1RkHKFEXWi2dAnqIYSoDCbT594PMZdIF
7Qx02unA/CiC0ift10oO3DjDNjXq/I55rjd/3N+ZXOZLmZFoQOnuFtzejha+A6+kzK32aDwsa3oS
jvrcaLn0VukEdYff7t9fmEipC2N1ftAm25mmNgeVr3+kwmlDUrKS8SiRozDwCsLSEXUywjMXH4Cv
RSxmR1qUC+23gIrmbI1TlBgtkW7o8Pr3QP/mqwxZajyjLIxTfi0yFT+0j+RMyKNLbxCjQCsjenzW
GoQqIjb/2H724TZ+yR/lwTY0EZtn2Mi7qi1+Q+THdhhxkiy7R6cOzdGpot91y80yKJdtcy2VseVV
F8aLMTJ7iC5jfgZQKtTWzFQWiAOk6K4JnRb2o/3mVqTaGfLCdPUxB/2g90wxkc928sF114Es704/
mGiXIw2uTMkveDSHYdxxKaiWOR1IFPrZFg6YI8fTLdEIxedZfptLRpObKRV00fiIcMXFkwkLltA7
XzcDKBOBoydq6tPI5hZWGUMgpdQCTLm0+tieXgH42dyBCLPs5TbSRTjGMqjTSZttxjc6yjyLAOLe
qCyMoXvptuAJnUoFwMhg54R3cFcvz5x4x0jTU6mTVw+KuCLeORPwP3ah1Poy8jbECBckU6RXh/9p
Q/7W5g0l+I99NfHz/fZ3gJyrinZTW1JQ6eGX+NQI74bwIYbtOTYZt5A7386un9rIr0oQTGVLimY7
JIFTFa1WYxtx6qZqgzEd+a+yXiHowQ+2hGnyl/1HXrDixIdRmP8yn74ngpKNQMfVfwBgIYP5mJEG
MXT91S7AXhFIDjclnBxfIJ37chU7EklkFy9Ga7JoT5FXtTnTyf+5IrV8l3G1zJLdLVUD5HEtCNTg
JvmR6izOLQcDoRhbap72/JwA4pbyb/riIv3qksFIQuEz7zGQfkF2/7hjizUtNKPU0aVimNhGOcFW
+4ThoUv/nOr+B2LX/GLl/DyxvnBMBEb0sRlOslIGWX6IBOAzUjrrNeIrahcIN7dsEJaVi20ERLiv
C5iw5WzSR9tgZlyL19mK0NWSd6XDY7B0GEkfFEGDfMMqt4qV46HnDh9pyoha/CCoSOu8OrzSF+47
V92GKt0UI3T15tIAGhSAjOgJwgFjCZLdeg2vms9wnreAyg/bCbZL6gvyLF5LsvHRuPYE66Rq+V1j
NZYZ5QTxhpKygFa2W1EKQ4J0/1amipxH41Z7QVtEJ/GqwkgLmfmF0nSDTk8k+nLhxCwvXJbJp8NV
HSw03ee5K6EiyYMWt7xYy9DpOCfWHPjAvJrdyChwIAx2M6oPZxbbWCs6xIdJfHhkEZ8yjvcyZU0d
G0rpPRwpOYIbwV7s2Lw9w/S+I7a1/WB2KlgQw3maTDSFbt+ihczplAsKNJTifHLE9qfnfUiAzMa9
GUER/iTTcp7WGk3lKAqAUdSiOFGaknQwVzmuS2vr6m0VDc2OEcVZX6w+ufRWlVv/A0NeSk25MMMn
hX0NLtexcmBKeJ9ItDbafTutDuUCsc3FZe6Hr4tlNkzruxHIfIIz/jsCIriLz0+8IfSgTArj+h0N
xM92+SuAR02NBQ09pcLipOyPrCxP6HPBxrvuA9gh5JnrV/skAMSyLnPoRw6a3IQbpGywGH99dOUM
PYUb22OMOPb4qAyGqTE4W0rg1VfbKOIKsLjaya7xol3JWc34YeAk9/US7miMMv1ucLrfxXwbs6fJ
WimuYPZ3Jcg+kMT0b9ZFuLV3bYnHQctYkezJyE0JFooDTatiBGBiOP7tXDOs039flfVcwxOnF6oe
fFeweZeu01FBxaA0v7+8Vyxa21yIqqPRMqAO2xEsqBK4oraJKrVlZ37iH1Xqm3dLltwVtXK2Me/H
sDZ7UxztcImp/2uZhvnbgYUnzsmND+1wYBCS6chURjBuyQNSGu6Kf4LtUR1cQZJBX/KwAQxdcvKb
iWk8k+C7clVgtZQZPdh9enLR1wZ+11uRv3Tu/8T1eqn/IWQOqv4jHZQfBqUEcN+hluBZhmHkadHH
g8DNvNPRgRjpCiHChv5FQIoxTCJE841tEwyRza/ErcmtQDgU/ACFKfFsogehoOZtUq2CaIXpSvDW
lCZxnswSJASY1lmxRUYcQopUMtrXKVko7x6v+4P/BSgJdM3crPKAdOuVe8he58cITcUv/84El5h6
aSXcATl87OMEn/EEpootkXTt1ay8zJTWe2hWTVF33LV2JoyabCaman/Qu4d2JB4cpBLSdNckUZdz
rdF0bCi82Nbz42y1DwNNzTKXiM/g7iF8EHvo5RJkbbgVq5Tir4UPlC7BGFpwdlxcqQ+O9vTDi8jY
qbqmE+ASbEUrjsTDTnUWCq+bCBBRMk/7zGIZMhmMyBaLHbXkpLDSa49bX/6swVpc9C83ejuKnzqY
vUadn02zLueFQ8NvVaC97s1CEyKMvZJsW6j6dze1evz02edWOf8pR7HYNArL3ITDTgWuTa7dd+9n
+JY4DISAJPLB/C4Tj3YYgrBO0uhjARigXGTysHXsV/bi99NXjAHpNTfMyk8PLGKImDc7uR2wm28/
MAf886JdBbH4ESQou+xP3FMJaRT+Wtvq6cOiX7CDCbb8zLXiGdNbboQFufyir4VINcLnU/vvlghV
eMZIsUG+P68fkw3CUF+UHvGEPOgfGU/Wfy2FurXtLT7Z4lrU4ohSoN3kimRDZdejm1zkF2qnfSh4
lCdYhX7cdCbiaubeHha1s/43vEPt3od15PJro639GV9ZGuA4G932q3KK04qDB9rbzRNw4R3SpMzH
asaUeruF/tS/9AhvtJN+a+jZHQqiBUKJXcCkb6J8Cl8IRM4FTl51qAOm2ZoFNHppZipSR55pDW4W
LT/qbOtceqWIg7xhyNuGTuAboRGOMzfCHm85URXh1UOX5YlEJ13Z3WQdfnMi1RiI1T+dNpeur6qU
hUi6pZHA0TMXrWRmKzgQvC/I30lmfI6+uueUspILOxatnYViYDGQUAaWewgVZK0EErmEXXvwqruw
1KGbn/iCoMasmyIK0R8mO5kG12MpFS2ZK/7awUXZIUg15IaZ2aHm8nnV83b8zNxjJz/deQu2jPC0
4FUkuBM/CUkWObKg+oyRxScOKv23SgrEQDqchrCNal9keZa8Kqq3IiwfbLardemJchtKdGtNZHt+
OZS8RZyLIle85D9NJ+FkFilyklJKg82/Y1T7LYughu/9mYPcMioRf5pGBt7W6YB3DfwIL+X8MFuD
go46ZH882FAqX3YicVOpDmmEeWZ2Yi7JVNkImqH6ze0XmOWj5G3Qs2Z813+rUWNbaw4QPAVvxpRR
I7Mf9DUdeKOxA/YF2fdTQX9jZDlF+sZeWlrjfoTrdfYoqIda4BWYWQmZ0UJrev2vBQP4LE+DISLx
qFaz5wvDB+8M47Mqeo+GpmGMJ5P6F5WNDybdIFDvjg4B2TUU6wt42pd4U6ioECbPhZTeI8Rq2B32
+2qZIF3JciZAE9ReI4VMoQJ7k5Ypt6pL33+sjx0rNEuS//3H86eWf+77ySlr9/B0Alue5JfAp62z
hDdMxvmr44Ex5ftlpACez4oK4iVCdp4+7MFCf32N4Tcp8AXtxO2yXzk/0o0FyUFclhBrSqjyl7fC
hSqsBsv6N69vz0gjJ2Jh4nHw82c74DeHwPUce3nd83aMKAxUJfjwXlADrgJdsZFylZv1xshu367i
IgXCkR92Z7J718jCL3uxo5XUjPFvWZIne0s5xRbgFd3Y1U3eELPT7GRFPUtxva6eFHr3DFRcTgkQ
x1RKDYiyH5QYXp3cj+1X6NHLZ39yBicZ9Q/ubRb9N+xgtbEyqaLZF9w49Vlsh7Pf7Bs/EeAOaXyQ
XQDkh9fZ+SGOrZ0GM5yF4k++ccwwQ+mya0NxdxbHQ7TiuwKzDE9zM0CT3jjf/iTAXwmPlvtKdMiP
swcf5kuAb0w2WSmvCp4iXmS3l3nSVqjJsGqtbpYoGO4jYuJYH8IxdZdLgc2O1ayPuohGT/bhRLOK
iX+EyuTIHR8Jfnr8tti10s+w2TK0bAKBg7TrqggPRtgulNaGMD5iM1341oiG6yodZDfU1qUzQUJC
WKI5pT4PGZAiRCle4f6bQct0/6XkPr2pz5AEmVl27iL6WKe+sItoa5IbZxXLlfJ1AC7FjxdejB+6
qehc24e0gdSLyqtNK5hqE+Ow3zhGmra3jPnCLkcUbqRp5Icxg//eyKTxbhG9+M6Qy7uCByh4VTVw
BLUXZl82W2+fcr0bjwYKIABeMrkMlNjhgYDnFMadn3pGKrvzQbqaYLdgvII3FOw87Z2jRoTtI46A
HgK5iwqXHENzAigPRVhwMkmb4ohtXMCG+j826HsoX4ulT63pnDbuvsagAvTzsbeoIHGGMe/+HYlZ
M3aRQAu7R2vqoARVKU0JMGhbay3OVUhCZ6EhX2EGCS3GZHXfbJTmOt8tcHSnAD3lbT9Dy/IkHUEa
+miMV9m5Og9wFZSyYnMmU8YZa49uXfr5ezgcuyBGeQuDuxHi0KhJKib9CCwbeUXaKoRAteh9ErNw
7HCuH+tSJyGDDHjOXeNFEEPhbq8RzUCd+LXYWIVjKRtK4T6nY5WM74RnSnWRVOEA4/avVGFBhVbc
gQoA72CuFlyF8XaFm2O4W/wQKD+fhETVxkafRRrMz1zll21x/fAv8ILAJ7BL/TflkD5S8BHE2UlC
kotb01yykq0bNJZP35TMZzj6l7bO14x85hdmkP0yEFLEUTtO2tHpTPtdxIuWNvRBx7IzZEYFhJj0
PMERvy0tIePjXo3AK2ICgYhfS4mgDOcAA5HPWI3bDBMK2YHxJgIy3iiAl5I0PGoVW96H8m/onNMq
bJ2jABfe8nGRSDkcLArSelAC952fhDyCKExJZBQA5tXGGjO76BmZ8s2aKwgYevS9L3kuJpbiM1Q/
GQnKgRm7jynsHfDXxOLZnRUgpCBzbsbMOdRiB44sDlzEF4yTFgpGLEZ9MoCVAAOltzSQ4SNWUfW0
yPX1ij/Sc+4FnsB4Ck+img21hb2YRVHdfKbJ++wDu7SRo8zTiFkU5juZj4UnOd/kX51QeAfULhgs
qgODHWYSSFjcbBCQ0bCel/cSZXaj3eEUN6KPT8M79TY4VWwP2W4sE2XQtTsXAE9pxwB1kwx1In5q
ySFeOPPeU4u3pUZLDQsq2wvvRTzZyJXmfbQ3YBB80BRRRS6NOGAMn0/kPwc5nXavScHmKyw9+Jt4
DGe1/GF9lYomVti5k8q8tCYxtpkum9vBsou8AOrOlpeMEWMl4JHCcZqI37qxYcovh7M4rsHdzJvN
E+V1c5SpGbJCrakfJk34jmfRH9mPrFont+4J/w3bVlRsGONTni1HkIxYz7IPVqEObZDvGCFnpsXm
4jjOEwd5P98ZNjtXNMWHvCuFfeMwTTv3lvUtelsfwguIjP/Pc631r+kG0Yw/9rZQLufZdsB9441p
SDEaOd54pjG434zGoi/C/1UO83vBklw3aujqkrLsnF4/nV+wkmQbmTmWMZ2BmtXkx5g918U89HgW
ybY0TeKdDl8YWdLqYJ5EIMmR2J2+pNCihZXrWEDT48vADBbbjbGvLM1dajsBk9zuOB+pv2N8qf7s
DwEH7czNl2d3TKr33W/vbCIR6+no8eSr7VOCKMKoAD3UP6X365i+MtAJCP7SfHMewQtJ1Ecc+wjw
IAs8cjHSDECabgPTY+hHuFzJrwskTxT8jTWyCP+4bduwtk9p7lqF3eIv/fAgIdrkNK3pu14cc9W7
aQhjkhZ0C89Fne2eAc9WQDSi6Nwg2FEf2d3AL9TO2GgQGZHOfbO/f2hk+EFP80WThbdG9732kDUY
5vt1NSLYI0Qgk1jTOvxmxQCIU0j8AYsOsRjMWFqAjoiXJvCgPY5xFeljQzqh3F8W/wsbWH7/O0W/
r2BAX27Aql9Igmvc2yOc0+gKBwm3pJQarmee4EFtaTnHDqdgT87K0po8cD3+Fg1MElMlEdgrVEad
jI378/ydOlMEvK2HbcZX7IDWEGPuip3xjpdBpUIQSZkot5E08hX/vVFw/Xditghkm6BDa8eYBzbi
Q6lPQmOwUIrgqJTPcbvpZCxRIgg1nNDXvIoOHJUeF4MAnT1wlHc6DVTlQgzqInW1YxJ1Av77vswT
b3oc0mHPkSpqpoWKKRCtAthp7Y8X9Ma4jAYoQz91craxGDtFqQLL5vorYNGaCzsmiXRqd99HiaRc
KROLAwbe6ZheI4ERUcQhs7/CBGiiv/ovTrd7PKhBhHOSQ4A7JAi2arftYsdQ4pD38ik0OcBdEmaa
MJvrociqg/McuthxW/k+33JSQFGGQ6vmfPvuaPeKByHYVkqhY2mru+fUXXe/m4n9zLFc9gMmGY35
ZxShewtASpIGNNkAYRHbfmoeqCgEXnLNfzjnG9eWgqR4pgjKlWyvXOaG4SjFK/nlFUaYiLqhWDQG
mV3rwYJPkaSNfzcJ0d0xvp/rQI73tjHe6B8rWQI78Bs6C+yZjwjyQzDLEJC0VCho1uBeOFhD3q2u
+Ffe6rEZn7VABiPSgF81JTVveKQhKxMBfmNi/+Nz6C+cgr+4ACGI0aFjES+f/DfZwzdLN/8z4bFm
tnLRuetBwquhn0PSzdaaKVf3BazKqSIIzJLI3WhknqUK1JtI5CvjFiHjOMvmXWpo0b/1LjhwYs60
bV8bEwSpDvGQOXDC1CVueg8st+xQuhQwWCRQF2HlYNINaC3kyWjTVN8f732FbnSqIaLSxoMXVkHQ
a4s8jEEwO+Mhlq3JO3iuL5qszBoVlohxuDEr7mepz0bBIfvnB63GjHALQXZ6JWqiMJeJhulkpsvp
r4AXho7vxxBMVzzpaBX8lyqD7Y94qyo9e/uPi/in23d4+BTj6ZwoInZUoAjH1YRpwfCc9/KS6nYv
ibPUIIAZl7DiaySPlg0NuEVUoNXTIg9YlE4lOIpiQvjCsl00pkcZBxyqN4yO935Smr+FPyOskDaI
/n6bSl8weP5q/LQgWpTV5dL9V6WqjqY08Th9bKSv4cQYPuWrDaGE2d90aHKJkJKCct3Rc5/y2Fsk
wLLMRtWmXyfr2AR1wKPe/nHxW4LK7wUUJRQmVr/O4TJCpFUttDQ195YRDLiOd8p+E1hLJ2AnL0Nc
k4xZQl1+/sbH0PhuzY+v4Oml24cIqWA5aFPt+ivlrTUEhKK9nanMfDycJclPU1PFeqJFdKlyTEZv
RCHeZ8MFX8FllaRNPEzlu33ir6zpjcMFcf17Z9a6rjWsdKmoZGMfTQmzZSd4XYCzlVErN3jFClWM
x1KFptLM9u4lwZtY5xN41Tb5J4wRmjzWDd55CqQd5nwaYfeet/nhVf/rXeEOF9chJDJF6czQy9iF
5Ou/mENk0jw1v9B633a+HAgmCtrIyJdh0jrr6xQTMnmoJiUSEpN000qxUJoVvyeYiXp0w+ygzAsi
SZ2vt/ybmF2pdmfzbQscozKr1Cd0zvk5n/CAc+JNAF6/BsLZxF3fc/ZBmpGcFDB9rqC9S3YXHwVz
Cfs8czL/F5weELOFJ1C4Kv980AYlvo6exjT3BB7EtsTgEIONZZDY4gB/N7TYGhL/J79d7mH0DJET
wSR8p763b+ztMp4R4gFDMonLuFlzMyqHtXkG7FFMoyP4fBlNueIaqPNRi4e+kSLSSbndL6GkcarH
mm5S1jXdUg12cxPG3JeO4QjUaLMBp+gtczqmIfUFUbYjd4ILtEBkHD0uu5LWLmDnq7UKWRilF1hA
aG15WP5Bmb8K7e4Ho0vSQYrC75E0z+/dhgbvTAVW7L00IAvjSaqWgJzEulRXheiv9lMr4/Fabjb+
wD//SKSKSkYQYgk9/X5FY5+ZzFmwtq5lyz6YoJgiCFKOAIsBvQDUi1FSPD5XY+4nkSIz1h23wpr/
+WUbB0cx+J1+vIFUzGv8AJhfdlctbJWChfadnplgwJ6dKAXh2fRJ9rE5Z0Qqlsf9Uj3N+DiUUJUN
rfD0gwpFR9i1hVSSJ+6SXmx/dpkEYqq74ibx6aGByDAh+Xezr0mihE8r1Dm6QHYpuvKT9f2Em0it
sQKLuuKTVkJSIYoxUnCFR6g7q4DnJC4Wh1LLglD9JjbFUBydRptbBZB9O4gyrL8cEHxQeugQvqJF
Qhy9ohIViUB2iHT6cZmSauIGkMqWJ7bFouj3sMJvv42uMKncrFQaJ2bWaDEOhkPoZg8Kwxkfj9Q3
SeP4kcAE0OExDaBzu1SwllLACRrPyCNjoJDd/eNjnRuq63CnD604W6pFvSs8xJnuso09cxKsCYE6
YVMjdOcvK2ec/xzMxYyOEDfT+VY+vPfu7FeZ40QcCjcyHwMloX3sXBwfJCetuP8EEX1eBKka0yqc
u6dN+3sCL8BPCHIecQloagFeRDCbOZvaCuJAs+WesZaOfW82xXl4u3teec0sZL7LJUUFtjlBwn9V
+S0IFPnriwBjgUB0vC0DxWB3KaIhmu28cZ8wBVUS25nGFczCeR0KsaD/EivEnF8ZQn/OIiDwWEzI
sDb3NqPbp2tmGsuT5Ej2FCSMrbVJkGFeabhXI48I/ftkJecK0eHHwGSLpdqbFohxUT3JeHCvQ6T+
sHNjCYXeSr/unpC0ZGSNz1rT9/uXnOltF1yYIdKhtb1Y6WSXm+s92TGFeoLCT5zwrSaQLZkbxkhn
/IGaiP+n5CfzbwSzPBsB2sMIogcFIo+OnvxmBwgdRImXWAyLSYJg4RhhTrTHh+euPAlgXNIDpbZ2
Z2eRw/LXDlWk6OWsfHooJ1CdKCUcKB11ShW3P4H2yE1Rvhf3ZP+genpUxbFUMOu/eXbLOtPqErHF
qI5Rd0tbrWvTXVlsEbU58bhoYfZAsdBgAitc8uKIaDCEZ5g83aMXGuDJVYYaX0Q2zSVz4U2XAaVQ
yumSB8N4TwpGMrONz0IrRTHS6JV0sSXmzy+iXyBTHLaTCF6ocvD+5YibarPwBldUP3QJTa/m1StN
mPH9h9H6a8P0ooppqw6kZugYLn9hb/eKFq+nQhXOCuKp4wI1AqDtQsxRsttBPt7kMrEhJYBt9FT2
tPvaZ3q1flsIF15cBzw3NQ2jUAlBeDn8Gkr6sRiWOcTN6sdj7CAKSrvLw0ebn/UZKN0loHLDGDKX
3PY4jQ50T7KhD1EhbaUC4KbCnjiZttd7iQTW0hlZ6vs4haBXoz+z5ElLueR9XCISD6PtPBHueYWI
4BhQW697Ze7w8b/hw/+T3ZEY2nhaCAailZnyz6F2Y/Rmgu/ZSCsWbJGpbbwF3Rc3DzaCPEENAOKN
Obfg1DXA22p1od15gyBUyCjhiV9FQ7kV/ibrCnpN5mhX4f4tPhjSHUHz7nuBu4fvZ5it9tMwWvRn
UZd3EswhoyfGizKhRSL4Uv/5I6okWOyxCeEjo+nN6bGe5tbhC/g/QSn8LscUPajAKC4OzbQVqtYS
d+6cItIdpsAXqNkW0GZf33beDwV0026g1+PX75c6fBuK9NxmIsvbYkIRYAZxkkELkdj4HrP+nh4n
DNzvBnldTfQjtG9+gG+azkDlqFmAmhFuT9CtY6Q0qK+GyOm33xZEf9vpASXhg6ZSWWlh5oDoq0dr
V1zxrG4oHjh+4wB6qlLLFOWw1mKnChhS6xYyKCH2PabWS4/wTV5pG3yY5uCFkAx4zcWzaHsDIYSR
eWscuNhIF7rCjCIqKSObuffhDF7kq3mOTZTE7CnvlZGMn6ws10UvlxutzAhFvtZykmWoSWJvlX07
ewFfSPEwittqFXI1SJJ30AoTkZvLAHUGHXNaI1M+U9Ak0HVrHYBzzoxDi37Jbmcbu48T09IZMeoY
wgiZERidYLto5llTjKWHRW8zKVXBGSZnbYY/j6RaJEnuNhEpzDVkJwJOvoyS22KV3IIrabjA/JfK
QnIKXM0AY4ox4TrpHYRC+a4l/OqtyiDKAfKhaeV1KpWKPr+oJVAGaY/0eDgm20M47MVc71sZJbKn
alDyG3tevIPNEqKRnigjrohmfuqWcQZdfrK0KGDojSXO4c/ft/bPurKw9ggyQg+TUMKk28mvGw0h
de5ofovu8bfijnXxTgI3Jx+53D96nH3NBgcGrdbuSZJPwRTa0tQGJr2MM025ZtHivTUohnAR37qr
0P7rvyolBEbxx6iuTaHuLvKeQUbEC7EyYnaHzFexXMGLMmbkvSx17ncjLx0dnp+KNIk9VMWI4/UL
FTzcUylnsXeKWiaGxQEnqwZhGwtkf7SaSyAzEch7xid016lVPf+NUQ5LCm+MUBoXggAwtmqZbxg0
HvcK/4YWthCUJMwaPCjS8wbGfV2XcS2pWW1jkzivaZ7q1hCMe2EfgRM+xz4JfIn78NorQUmxrdb6
kMP4QxrITEetGd2yMGOeBEKJXeHXBXNpaHdWj3toZJYCLwWckvFKJFRKHgM/CKTdnVw3j0uXxxiR
3fWjj46RWRKxeesLlUfaWzkAdwWZAn0j71hzJURBLD2n/c9oJmXFZgGdSJHqFowSYleCByrOQ7jB
J6kiqUCGwv3ahOPaA+W8ZCIYoRyAljWN9lgjDrwkMaMidpxzxH6sbbBq0MiC8wvV2aHq5eS17Oal
D1m0ooVvfsitPljOLDki5T0+ncc7miM3B0vmhRSYtnjKBPQSNrN7Q43sB8H0PMsaHrVkP9UOn2P2
mFdgYT4iqrHJXygjJQJdkB4ZgacAGb3oIhRklJx+hcVZUQDWMUc1RzojRmH+DqJXgIziVQfOlWHK
b806p42dt+yfrvPiXAtaLfk2x5HVzZXHrjHgB+BgKhMeSig9mjUcEi3Y74lfCr+BLLi/YZ+iLkBf
AnoHFUJursELtW9AVtEqlkA/O62R56RgTybcEUdaXZwbNUQR0iy+1KNC7b43mjUy2OrowaJuF0eG
tJ67Hvwbv7w/5tVXzwAXq2lsBkV2/0fnqhj3B8HYNOa/kqk7yZniZAhjpNJ9jfV7jByW838xJ+kQ
vYMgLcs89yrvCBliJ72ixrqPrW8Ont4YTy7sYcSQjFPdlhzIeb6LY2mtuAJGm7dS0M5lIuM/FY/J
dND26h82+9XcQULilVraOIEumbxjBiUaecZemq+zvsNJRDXf2souVz9CMpptXjQDIS9IDjJZrV8Q
Ng7Dr/XJmfGpOE86dH5WqubaQo5KXXrb8ZkV30lBPbOvgs2eTCGZhNgx9guKY88+r3IMIDwRRpTe
w/s7rqhIHwfA8DGTe6cl8N9LEjP6wwfqP1Y5XdsOlDf2isdawDZtJIOXlWJ9sFxkud1tR4+Mt2TF
8XH4rRw6mChKyQCpamcCuAYFR5F5pC+gjTAX+wFqyXMkFkH1pAQtS9L/6Y97iFrThFUhAN3xMlNw
mQ6hXX2EelxwUOcevJSvIKllSds84hn7ucCTJ+CEsjbg1rvkYWBfUJC2tmvaokyFiEWHnZ/N24Dc
F4eiukyuWYXqUwoN/SftxEceVUDM+nPCURwIANyP18yO+7Q/hfvpbXnwrHcE221skWi9UCw99sFy
TQqicNa5Zikz9BKfC0Te9ThioRfbb7bVuJVkcD8WO/JvA3Vv3gueB+hcCYpI/hR89mKr5xJVdGI9
EM484lqfA6URtiT/tGF+zyBRlg1qXs1dYBB3A1cbNe+rFQTIFl17xhHp8ZyzRG0Y1lwep39opT76
9qeSqXdOKaWIDdiOAC49PwH+udn3Hk188jPrHlJNdJCJiRIfENZJFvgyRim+HZmPRXugI1kU7x2t
iIENLAJu3vs7MiTJOgIVcc713KV01eUwPVO/wHcC8PjDLN6CwOkgmctxzMXurmgCySBsHr1UNIhA
mwuxM1fZCT3RpKS1Kx/eftKyUku4BA/HzCzQqIDoZWoMU4y9fXB9ijir/Pf4FNktdYFKG1EQHu9V
Jxg6kOOtMX8onmf6JYIqjVpKLhxkY6K/85LYZcprozkoIcNKHYQoimCGk8ooAq7KBI/T2M7RJxuW
q5/8fu8AlAL0DoGLdeVj4ImzW/qDjVMxFiNSvUbq4LHhGQ2PX8velQUpgur4A9hhfaifQpLjBllC
NwEF2WU0/jwuspWeo43RpDfe58wtyAGgC0643VcM0sTSsNV4qVwUelqpi4UF1gXr4AhUyclFArPS
D4z1UH6bLTM8qk3XjpYAvTQFVw2qALCL9WaJ1Xp9EJfqDrtE3pefe1v16k3ic4zXb6Q8cxlwzbOv
MbqiL6eb7SbNpVQW4a4KvN/xoZ6gf8HQlIQiZsuFU+MU46iJvfMDJWLm8VGcGpspf/ocUk+CKhlh
qdtPKxgfoHTeBcezfIOzXxdCKsMU6Gi4wqOrxS47fGCUpWLV5kMXZ1GoPVYbPxMlSebthewlwzLh
odQ6stMyh3r9h56/OwwPL9T/l39QhQj0aNPq1FS+tKyrTx3jnsqfPSteuu14JtGmdc+WWKLWQYiR
COzjHSKzU7P/fK2q9Yz1H715XqRCQVg7glrJpSqdErfjRCxwFtrbQI/YxLUY4quXp6JaweNGEQA4
ZzJ+T+nHrp7aAjzbBvCJGUjnJOL1Dz7m+SXG0OBeRORpitFkD+/Rf3Dqxbir9lZcKpzsdk/GPdmM
DI0s+bRIm5R0zc+HMyW2bii8n+OS9eSZ9IbFtsF0mIQ7bttPE5Crgb/BiRAeRGKX0ZphhdGsWgaW
tp4b0rqJGygPcTWE6AOnCQRSdPl0hXv6YRJ4wBGr0stOCUO5dc+UY71aw6N9K5QYVkg+UKJZZRes
53Lq0gN0X7ch2yE/5LdsqQVkgMDgQN1qsk7VKFayXq8eQuN7CL1T4jas74bM4nfboha7aiB1WXg+
op7XzhpvMLdLLEMfnjP44Fse+4OLQ7DkLDNtteQnRKNADopxkKzY8VhqwaYmLD45aIbH4eA0yLha
8Et1iNnm5I13dbvDcD9wrl7iyHo6qvVSCBMcFDckyFfjLe4elyqagbMK9TimK7u0xJRMqLcDE5SU
upwrfGIUOClwEUtGIJYHk2sppfT5YeAkfH0Qd2h5kuJcgTNXP5n2CWQacMHhhNhxe9dcIDZEC5m4
Re82KECTz19fp1etUX0zFEKfU4mjhGIX2DqM4Hz0MziqlLPsiaiOBDYIbqYf02uPttxkejKuEc1s
pZ4+5MzmA5q+dHoymKPAaGYS4oE33oEvNkn2Ejqt7LKV/PhHKUg7Do/lh6+03lS6wvhmUTdlsA5Q
qveaCYBb9p4cj7Xcr3X7dUAME7o/S5NAOsi9rT9z2X8saACM/S8SrKzZft09ThZgm417VdCmvbQN
BFYCeXpOyOklevoEbJn16/Y5oIirnQaxNlTT317CN/EBdkrAyZ5g2pVfcKrLynJLxC7TxT+ODQQT
nxh+7E4hDJi0FQapbMSgVj0ivnEkbimxIboeHAm8FbBk3XoIJI4DkbWIkHyDgnWnJ28Sajtn+OWL
QRh/uN9Riq9QTt6ZrsrMVVEa99qWCqu7QUcWDJynNSTNQgytAfpewHRQBCg1BepB/q6y6yapvPuh
N0mefEhDvBMFRuCBVsr+xRRTzHLyI58+K0xVhwbUSDGvn3ZRETT0jI5CvXIjiroptXDmS+ptvyUL
SKUpvO2/5qHOYGpBQQnsM86yWO6z29CibZN8FYavj7iMnMC2CQ/bXzo3hVkWLdhLM7Np7j/VzAhx
gCWerxUnZBaPI53IC63J2ESYKQlZMJ+nok5qlGZScqBH1QIC5hdV+AiXODcZdf0ZaXR69ZzRjvq/
pm5Qno/KLXnkjWn0rSul2cAM4zj8MXWSNUMmMIk6k1u/20AaHMjDIEXpAII7vVzS3ui71NKkvEUu
5/mpJ7osZKaeu4fvL0O56MJwQacDniKEGCTpD1Jgmg+NYAFDsf7rwNcG1fe8LXdlqOy4iaeJ6oRX
1EkSvKQuAhEHLBEPm/zXCLIdyJqtvQq3FNBHrnCWvpxwZ/RJip+rTU63XsyGy0CjEDENYOBKPtcz
gs5Bif9DxhEUS1XKpQGAkmUG/dM3DwAwICQQQBkLaRCx7d/ecylESAKmQGII9tVl1aNjSIqwEaQe
qdCIC84GPBuHPhXP7LCoS3AeKzVlV6izZ1r8JULk30hUxk8x4pcUg42O3qtEO49s6Lm8pg/aeePu
umqiKmwkB3lfa0MxsybZirw75cIldYbxGgBs3vA9GrYsIxHY6DHf+gYstyJ6PBioSU5TyCEI+rii
5DN+yYrSvJY+H9/iNpQvdV1RZZrZpa2jecTOCKnuG8YxSsoEY63w4NohRjRScZ2N1z5ItYUUQ/w4
ag0gbKVhz8lAEFO0lG/QAIXtjT2UNC75RkZF09RqwSqQz56+DpwClw+1V72wHjgY+/VFs7gRStA7
Gj5aBEzfNnA78x6M3rSeHv/xNuzdgvO3QH01nJEfojgnRlhytYUnZo7Ra9LJOWuXf05633Dmm5cm
Jm8EcZZKID1XbtRQdH0t7bg+KfVK1Fjp+Ov/Rzpz+vJ4urYM5tQPZbeGeyKuJEfDFGy8dUTUSOx4
+3JRu9leUa7VOoiLiPCBImR8HkH32rHUXl5616ql/IPqo4SjzxNK2IsJINUSwup9jLCzUlr6DhrQ
q/j3KCLj/1/0YHe1rKdMjXhHil8/EgcE0qutbNFe08qL3PJPuzDsMJG4ijQH/vjS+iF5+klfD8rm
ncY8GpGivSqJJUXPOhky6/Pbmw4sLrikX4DmI4RPazP6nF9pNJsVbKO+LoZMpSTox1C8NYDCiNRT
kpjDxh0YFpGMsXpNVYBeGf0H/duHfsIRaByiWRhZT5vgv3xegsPCCPhYpQubpxdZJ692ZJ9Aq4IK
c+g9gNDAA3CvjX5E2zmRZ+wHYwXot0Hx3nppAttCpXepMr+to6Z1TBLC05Ay6x4cNvXlv5YF52aH
k7frBAQxHIog1L3DM5p3G57N/CySJR1zlpHR9CEBkVsd0SE5OjoyUrGMK42aE/1imd7Q0UdkB7kq
Kf6uraWF1YjZ+IhSy3+No1bnWn3gGXgGfr71xqCCmEnslgjawWd5B47+VzzaeyBr1QU6zbffDDCM
RPKKNBcE4i+zCIWo8UG8S8Ton3KYK3TA9P46fkHsMZdYJxrZCknPelcz5kxMhFWUo9GGsKnoF/D2
442F9cu9g8KoGoEnlPvZ2ZJIKwcDntFgKj3xhzyWLXU2uXORV3ZrREc3iORyBXTaS1eo1AYvxf3S
InrTmj6KK+haGpwzYP67w6oPLi1pvSWPtJGIHYRl/niK/JFiwinnGI+Y8Vi+QZR5xUKvt6B1FAyF
C71mDBxnkJEsXZx5zIR7unqpOxNQd1RJiYE5B7gUwhj9ume70pexLMgcq3pzzDACkDPVEUTuTp/E
ZetXrGDs+Hxxb/XiNu+PrgLch51Np7iaICLpxMJ7NQq1LUgw0LdSO6F7XmhSWKD4+6pgCHpQhaMK
kLFzO6QV0LkBhV2jcGnbkLmDGvTZusPNLW4t0HbB3Xof0xxIYwdCoAalL4zSttHbDmfgJFz59LLC
Bday6vDqN/wT+qF11yeOaNEekAXjSzzEcx1A0nvnNdD/k3P8DneptDEb951v8qmd7zj2Jc+VCQb/
4X6HArrdmZSoZuepU214HlhIsBRDNQ6Nh8ElFI/z7/vskI86wFjQtKVw0u+iSAMYFFrImeeC5YsG
2nLVIRtN6LKyj00W+acfZU0URsygZOQHOs4R1gYGLuXNIqXkhgFTMr/+ILLbEDvIuFeQHQMBcSH+
FyiKi343Mu7jHDnfN1ke2bP69Eib1azFnlmE16E7Z5+zrDQNrne8iKWfj3aZBIozUH4WffGmYCjq
xYkI5vWTUbIve2luCxXbYiFu28xz/H4VtLcgEaiOZI+LIJ7aBkDJOTdVaC+9iwqAJTr7DJJNDFUa
udEv8re41UTdJIjuIY5PFklrWBREYeclDwd2Pef2JEBn+L9W+x1E3oU6+F8nxxUb8WCeJInY38IH
zdutnODHs12EmVc3lh2LObJCJDPEGPPsuSgMYnY/BFEQwVORB9wfsx19XSjOaY9x7voaEqkIpMQz
VSuQjAvGnGPNcsKPJOmG6gQ3gufj709vXez4wEu4vFv7VBhDqyOjoCIaMcmstkzpYYlqm9/WpP5M
RJqXpjFIjId2wSgfdjrz5VzPYOY56GcYdtnbNQy4yatnruDELvwuAuwlEhc3vsYCb+NMavYbUaBk
D+LjAVwXKnJGtJQ7avJSp/sLtnT9TyEDXeCotN4rfn5sYo3xrKb8j81dRx+SSfiVXBDtsyKZP9Mu
oFM7RNJhEWPqWItpI4h9LUUqw3k25IstC0NFJyt4tlMAuJqKtB3sKi81keDMaUbAGplVAHjCvdmJ
0YNLztTToP2SMWwpI9lGCYv3/1lDEZbI6lvkf5w7uE7HvZF4UzY87dceTqOQmTuERgOHGwhKklmC
Fqb3LfLprFxJAt4tanHhvQJzMA3cq2VoHxcQ1oGmRVQCj7CDK3ranyrIwUXAEQ6WPcH+qggxsvZW
C6aQdWl6mXaKcT2qVbvG/IWKHEYUaA2EyqAzslvvkBo7sjdJ1fzcHSOwhWGSL+rV4vKl1MOrCd4v
WG6MBd/cmyt91HaTRvCjwGvOJyDm3OCdKkXI5tyiwEQHQehE7xgiffzB6Ehi+9g4CHSju9tUJqYV
vlPpPWYna8Do59jD+3cLQHVxNdeuUsCVxXlC1r40quPh3iy/E7fGZMgDtLLD7lrfBkAMEvKFDxsc
rlgDIoUI/KSkIGgL3QRhy2XZOD8BIUcfyvPbNtcpRnoDQ07oqjDhWyDCSdi+Kyieccq2qHd75HGO
RF/PUni/cJoj2Qwc/XzWqrEbznQ/oOc/wGFeNU1T5ECdj2TKiQ17bXDd7DBfhhpqj28E4sLK8xfg
x6U8Pe4fat01a4LYevTB0l6nim4GkmvuWQSJI+MpLOSos2iHI+7EVmgvY6CjhxRT2ScB057KISvb
kQluHV5/VUwxhh/gEG2ZV105jSlL2LN9EF8sUVisqEzvCkuavKowjsG6yx2QXxysxMrx0lJa7+l4
rer1D+smj6gp+DYK3WdIfTAvnxH8efxOwCUMP/wC5xcp59yibm9mvTj+GA+8R0WKpPh9v/2GwF8p
NDX4lc4/6tisCzVhhy3kryuYs08AIKmp47S5Ut1AECRX7XEUuhGzSrHPYFwc6aGlVyryE56kEYI0
Pya3oC+Xsa9miLc0cqLuVsjukcG+r95MUHYqAX2bnskQRlF7GTyTG89MnCQbkWQBp+IyIHeBc92Q
6EEsKFuUOv+hjXFk8gWp+au717/N59VZ0ies/WvJZx0M4cpkRDxXP6EiNrf9P2wdsM7rd14nYF0U
77R5wRP2wFZB8POVVKlCzYJ3/iIzkuRP/UBgs0qF9LFiB7hda/jkZIDOktqfqqGdOKkYBULEVs97
yqwatm+h+q+D+hvT6gajoBj3NjMWuMeT5nhErHn4MwIaLG6vemfpNVqoJPf6IYvKvoLFeRf9I59K
ih/Kxe5FEEOTJ+ccckYG7VmDJ6ISQkv12z0xUN4s1phHjz8KRy8qJBfjuAkwNp/paCVqaKvPFw7O
PrHR6UWK5g2cegeGT8lfZUnVEEC1FNrxB93QFk9Hm9hLfAtldW8eQP4TdOqS8PGNTECzEXBtTsGV
mAQQF0QyCDigQvLtLXMzTz1J8ar7joHVi/5lOou/7rOGKoVAJK7flzP/8mx8yIJwCdC2Oalkdsaf
LUbmsTHJ7tV/sK04AnFHDL43DfZZGizS6r2cOikRW67wiePtpP/eR/YAdbyylA6HTlQRdvPvN22B
uIWwygISwKKppTS47fDJbeuaoZxV7uKOUY2KDY6PMm2/pcK3idFszVV1+ENFSYNsC9IOZxgt49vD
BDqH1WxzTknjmCmofTR9CCxuXQeaQ9cb2UDVCfdXbdhc0KvkyotQAMX4ytZ9/lKonu7uC886gbee
waqyRuVgZ4dquKmleOLQWzxHnV755eikAhEFrWd+unKNO9s+8jOuwqb5Hb+czLG/zOj4BLe63I1X
og1GDk3Aq9pJJT7ENbBCDgxg40498ngvnBmq7bBHcKfd0TWpLL1Eh3C26vz5akmwXuosu3t8cEDh
ADIgFQZtkTCrC1BKHP6Y/DlMqfgSKohnsch9EMTLX3io8wxktTC7C/0ixTrrZ7c9l1G1jX9fyF8j
xui6xBo4rrVVdjSBXuyUn42aoYOcw48VQq2c/f6ik35+DuMFxooFzcLZNwCe5QaeFiG0Ns3TTbp8
yycFobUxRzGV/DiOHgdQNpeB94eZa/GEuXdZEkivb73tlUZeQqEDBOYSYH2OC2AjcbDAepmSL8RQ
F7uAHWWXARedOOZf+HsgavfcuhyfsFwzPJs1nugZ3bqa5RhbTT+qiy40BuI42rqdkBeczKrFiEjK
7KDhCLT3PO7UmaIszGD8wK92qyhjuraMaT/4R3s1LvQWLhcYRxD+gaOGhB18+VQ+nLFK2NhcMmJT
/x+uaU+j3bj0eSLBsofgWAq9e4PSaboL0C1hcNffrBMztA3FCTSxBrg5XRafWdEbKl8prfnzib8j
M2RUsJyF1f4T9qPjpEwGoFOQYjDIpYYZgrQVn2npeJKDO/nkc/dGytAC2zMuYVYshI5W8iy1AEfX
NwSsYHapenguLJ1/B7Ym7sfH4HUTqO3KbWarx/t1A2BPvlPBEvWbKTNkx7L8cS/j8XOV4F6/uwp5
Dj/+a4nXJmSHTzy4Ln3mWJrkm43y0YRU3Ei9/AoEvRNMfEH8LAfxTr1Vv4V7/x+F+njMxtS5EHTq
XGzX9XZj6e2XNB2oWcM3bcjGbaYc9qkToIoFF/ykFRn1HssKerAVHdzezKui6GwQbWEpv95qJs6r
hmzQiee8cqTFRkAdxXN43dAPt8N49weUbeW/lEj0z/FDx6Eq6xtPp5reDdaOFkbaJgDSduNuvwlz
JYYRDmkIMrIku6xnWsCGbPNDAkUAw2De7VdUEwephbNahHB4L8ogKbSCYZ8Nwr0sS+z9HYa//MH1
8ZE+8SFzdgsKDqcQzrnR76q73p3X0g6+LAmZxjOTBULH5cdroAKtXAt/yjwlux6spUF47dmOcBCC
NPU3+GvW/EyVCdzExobBUUfCI/oi6b4S278XMJjYhgNa6/K05hPqpEXC3sA8mzE9lBS/vCOtFALa
Eca84WvgF8RuSqRUQEte0yH02C9u47jzKmruuKbweeKer/J1ZV0WvPTSTRREyRkklJPKcVSVqvgB
XQu+UZF6YIYW8QkCMzLotK6d8GtZn5zSGR7u0H2kPVXApQZE3ogkV3pIeIYviElgiSqo0DAmAyC0
ZwY0QlCV9V84R2DdDQO4OHv+1GkI29OzhAzoHiBzcbkC4GNyuBZ8E/FZkgVb0JhPbqRKC7GfvvXi
EP8mN9psUe9a+84jEFSd5LfvQrDdY/0WfZjqWC/VWehIot7FhdiD3HFeKc/HpfvwJP92cHgdw93H
ZyigEa16qaAmO2dxwgPsnS/gnYZqd8Sf7Wvw/ibmMmXKnGoHhZC8aw2NtN6vgGwnvpOQ3FLeAkff
IN8P3Be93DdTv8S6MB1WBWguw5EiDCwxvabPbxgwhx0rNsFwKDVfUvlqxfWaGEvBXAby31a7rvII
aRxmxiGDhXvB1hNJOKcflk3UD6JjJSoQ+hSUO/y13c+2ZNYeI9VVBImrVAmBumDPRl6NoMGMJpu2
b8S1g7zO96YaHQ23uybBlolx9XIjh7+re4TvvNFXZHZp2adf6xc09I5Y96Lv+lv7jRAvGE6UpJ4t
9vrPJgeiDq5vdQRmWIipUFRdPnegnzub3sJ1SpH1iSH0+rgUmXK6wMYuw9pB8gjiPYZpm0zl+lps
Af7Cgs+WHONp0MciCYFd/x/yuiNwTo0/9J3wWVXZJj1WXq7CDbaUP9UBtPmje+gnY0GvGBtDkT+t
3XB87RqpP5Tmk0mX13fWmhLPRZ1le7PdFYe7LQvVgyw0ws0QnclZSFWG+02/VWaVv2DoAzvGhND4
tnmWy4Vg5dkl/OPeZS91JaPlpHrhprTkQTb4VMnUZfeXxMzNZePoOnxcwFaSw2yrz89UI0xJCWVE
1w7d61zG9Sw9P71nSRX5QvT5fSU1VV0gYAZ+SaovS5jCM8PhiZILeFdpP4tahJhaMmvIuFkxIM2L
rqUeR400J4mFSgDUPvdSBTSdsCEbMeBRoxdFiBnsH1cIyfNqZ11m7oPAC8LY21sVFf5484Klivsb
fd3R1KfA+kZ78a65f5YQWh+A8m2sRuo27+sH1aAtsDYcyHKAAST2bngMgGLpBqX4Ng9t12SCIS1i
0EFmElUsihY4duQvfH086C7mK2RBffLNLGr7qbQbQSGITEd5/llJiwlDuSoZOqIocWY6UQCOlJh5
EgohueS4py5ZqINLGN+Kr0fny0aERc48wbukpuuv0/rYKTruZIoW1Exnot6zODHTLcl16A79fjpS
CoXWsCnxmt5bvW3RLsc25uh6dKfW4HCgMhROCc6KLCTm7i76rgk+GTbZie/Zku2Be9hjWQx8g8E8
MgsVy2p0TK0oxRBHWoWKhkFNVhxWlAv19AWcNriqdGB0XE95XjIb3yGt0wfNjvNbaP9iM6+HMWqB
b7ZsJet9t6p0YUxhIHjW9PQT0iMYDuh02Q1eqWrfDisfG3DIOjOW9F9+jgObwnwd7bN134+3j1k4
YvdJa3lOtHt2cfdaXSeOfoS+KQ64az7Shv1IDdaz6SU/x74lPJN/MESwqsj+JJrnsajC6oiivWKX
Vxn6/bhvG2oDQG9dSXZ+Ixgz39xFOze0uBq250rPTUkyha1YHhs7ug2xJt+6B0ybtQFpUIs5OMZ3
GYXmA1it+KaLNJYb1lbWPU1bruK+d+nBtJlO3iRDRRX/4QDw1iTL5ApHE8FWya8Y0fQBWdDAQnAb
bn7kH32Qt1Nv8NISbqMjB2QLMjEL0uD7IxBNBwrqo9hPCmd0DD3XrITiW2IJKfalhGeQ42McWRbH
JoThiTs/UZPOaOwbIZTQh9r3nuFEXkPsZipsEa47ZI/0G2Oup0ePqcgJWdIetqfHfhUWrkqv6bRx
63StCMjC8P2PcCIt+AsJLpewPt9fnGoyT8JQXo5mrxMRCItam1rtEElwlW/5uWrSeLwDcEnjfYCL
32v6i2Gqr91o2+R3IJIABCdyryImDiQdsU4zS3Lwp+ZNAKA8SQw0mgJlWWooK/T4r75sYWkVQGrv
W4wvH4zUSEN1PMm4CvDDVpu0bqKvnQkxQKbdahe6YC2+6zLhkL7tJfdd7XyzMsScoIl0DLDrzqme
Woqvjd3e2Y0W9qa7ocmSvQAFRt/hRj4N44vhv7hQFnT24P+LN0bN9yWeXcRxCwl9rNwtLfcfg25E
1XR3SSEm5DyMQwxs4PwNQBR2yMxW4VjXMlU2vQaJjpevnd4snZoPu+7pLdB5BQ0F/9E0skuvdiTK
IlnEYr5WF7Io8770jSObmJ1wgLSgoPPxqDVm1CSbSpKW8ufd51JMvVkix1x2IR3CC5Ipj1+00Tyl
YM3bNYS4v+b/WX0dDdYvjUg9kk+80hBzpXxivJv05P5bWhIOkwYWPbTsZbU+6LvPBNcAr+ountw9
SRRIcJJZJJPGfMVJKJDMnj4qPsDxmKgm6fSGrsSt3dGD9OSDkCsKs41Ux+SeugODuMFNPgjT+J+p
uvGBI1IBUQKZsNhGaqy+ShJ5AcHjyFY3r5NcS7x+werQkGOk5aUz3HM31biNY06XeEedJEe229Ov
MwNZOCVXuM1sqmbVru4sjlSUZrZEcw3fjo7+yJLCdysGUe3ZSL3Zi7eeJ/PwmFAvRxxmV1/xubpJ
MzGx2mcr7lkKRR65HnpoDg0lrGEVm8ldi3KXGsPXZU/aJWwTzG4ioK258jQILKvj0fMUjEhx5oxD
j7Kk+BBxzleXKfkEaDB623hpLlAMh7Li3hNhjEnlfXHZkw2Wy8ZtvmQpJShkijzbv0AUe5xP3pLo
ScG0BjtOh33KqF35GAMm/UnMt4KJXbIWm9URqdt/ZUpf3anOCUHgCIK3KL/4EXIcE5gDEIBGgP8I
W4VykDLeXyn1l2AJqCsm8yxocWIZxa5GeugePS3K0MlvLuT5N/YXtCuVK4DLb8z1+2w/rYjhEZsr
+gtLVOXwYlpeOnmACoVMNqlL9txPtHN4677ddCe/CVO3jGeGyZFcRLWUPm+EBnviQol3Eccvrlfq
mHrjxYg8OW8y/b2WowTRaDk9aKN3Wo71tTUe4AXZs1KEYR6dMjjFGAKbDf1UjWrZgZMH0v5n31Zi
XkFjXN+BFkifShsrDjUV6vl1de7bKi0z7LoxoIKQ3SrLqZD01WAcKaoDSdeIO8G5HF7SpAnHJ66m
9dW32JsTgaSIYPvL3Ks/7lhKDUdvlzDQb3N6W5Enz3vE6NDY1wZbmUQR7tpr13+/+FcjM7anoKwU
t7xXB5T3KLoaVNkasWfg7OQ67++l8tJU079JNRtC8+9SjuQfA0gOAYON1iAJ2aW6HMu5FmfJXDUT
JMDOt1QN4XR9fsHX5JoTz8BjmNeUMlxTUWeSVQg0orEWWbQNEr2zb/0J+7yq8xUkuUyx8n1IZPYz
lGUuNilmH3qr+B4jLognIGdnGDvxchEqnRnfOV9Uv4/f417PJ9a5uFh7F4ZKypOz9LPSDX8zmk4g
s/SwlXVfo/9DsopwZrlpSV1hB+SxZ6ffytz3ehd6TevDrX9soLwD5WD6R1tKVWhbbs0K9olav/b0
3zYdRtTfFBOjZkLPDaNg6lBFS9LLLvxpA/uUNlCRh2ydWQVj4ybg7r7EWaHLuAiem4cCN9lDzLQR
QvfSuabKLa/unreP8spsUpMF/z0QZFCi8SJeyCtNe0dkZDosRiEiIm8KFOuX1bHHe6vVpCm2iNR1
EKpHEBq3p11gPhQDtzaVbkj0idhdt4zjNAjCnQJcRhK4uvgVd0pIPaYZhNUYM3CA2dJfSvRNuaX0
BSnlCsYflGeg+QpwbgET9LfUt7aGYNnTOac9+uRrRM8+p8mbY0xa4Gc4IPADisWy4bBP4byGtZxV
ByqApDQ9p9GJWxpzePbj0WnQoTkc/aIy0NI8rmpwlrqoi6B9uR2nCJ4yhQ3HW2G7SnbybllUXO7J
aLzY1iB9Vg5gFox78beOCZOg6t2xTn9A1vMyAUgOyyxGfjWOYbNvGf9/Dd6OrJmqYhsDI06eP2KE
hlElqXac3kg3SwvojMCCSDFWVwbZeGKDj3GW4QhOTW4pj0YnzacYJyrq/Qf2PzVDvLRWFwtV4oL+
profwdhAj7FoFI/VySKhnbAokc/F8Jb8aakLAw3H/s14FIKMBtd/zhgrfeV/5We+mWOCBBzKWSax
W3k0xx0T+1GoAtOv7IuOZojdnyMwpKtOKZsjSeXA3SAuuPERd9oeqsGCbX2uDA2EeFdJljisd2jS
ynbrpR+XSymIs2FyjtDxEwbgqo0kYOkoBPhybqTu1JXEzExqRjbqmG0DTzx7MYHZQ/lYWN6nFhxR
4YBXWdRiPki3278dGa7JFTI5n2+ZcwWIM23x4VRwQRDWj1A9JmuDSMqTX8idYRarlCL5gk7QCQn9
cfajkZVpRdkXmNuM34hUghxiBr2qhFIofPrkUErIEvtuNCYW8MdYaVmq2FOZDD5W/OvD08su33Ke
nwNXETcE8GuPNBT+Hf6A2pVzetaeLn7skpQLiLzp47eMZ+rVXW4TOEe6dBGCYMfZNnWyoPJ3dr4A
v3HJS4K1xYR2FAn9sCkNuPPUib1VgADTMTP1lEK+/8Me67lUZ8NQ/j8y7Nus8Ntc1ucalbVuaxeD
Twzq9j8BnKDvTWVRNHE3dJb2Js3EN+yExHlqADET7uMJqMWs2+6uA4Sa5y4bF0B3WzJOIk/8edgo
8lQSuaLxS+m1O8fG90Tf4jjQER/1aabU2kuwoTxRspkpFzMAVSgvWXfAiOu+Hzzv4aOxZI5+AQ3k
8zg8Mmte/RYc0wQacwttslLwQ4oAHJ+aeAft8CK5mxPEjtYVpNEvd0lAyQBPx3QIRvWInqBtcvKk
pgdaaPCDpLVtBKSA1j4Djh4N+nwiOQ/d6T/5zgifc5hX8+Il/5wB2t8L1F9VSqd+aj6LyrzZQS/w
xv0MM2EEVJqyQlx1dhffAkLFTjKK1kIbUUSBeIXmL+6+ViUrRzm7SwnzNRGNjCLCDN2HMx2uEw76
h3J5wNtmLK/vJcb6cbOhHAXbAFyKgKzN5N4j2R3eEGON19MQ/hWxGDeDLgbexUGv6srFFye5LbpO
3Pt7WAS3veb1q+2dAZM2+KtoOqLzNSQW38pyST0wRA/0Avj4e7CQfE0aLIKoC+1H1Zezsyhmhy7w
vj1UQJm8ZkTFZmGF3Y27H+IHOsfzlv23j4/QMaYtNdjzg6th+JWp1N0Eb6VcsX2PEgkUYwN3Kws3
G1iJoU5/bJrYXhDTUI98LTawpzxMdl5ZDzhdJSSG4196LaDkeBqV1xgGR5PlXdUePa6s3JbYI2/7
p0avJtoyQuK5H6GHL36CU4iEVHXe75734YzEHY3/M61SWpHgA0gGVLvqejFi08a8NAY4NaGEaoEt
9dbUG8wVJuiAgN+rPd6gvpnKSdBvKg2ocxK55X1YIHjpAsz7RzVjs/adqIwlXqwuYRaPM1P/jC8A
sDIXvJA/ZVzxJm6x/DPBwz1F3QHr7q/rcw0H5XyxAsjtgbaRhdxPImh35XgDlSs6SV3UjsKKqwk0
Lha1yWPbSuekBX5NJ7QW3MzA2FTLkHU+Y2PrALp+zHtt7PjxMAFXBdis13A/KfiXSEiHhIYk6Jnx
ufgbl1DxVNMRrnoj5X63UYOYUteUz3iegs2cVfVtVEv04f2Hj8DFUETGoWFpKk5ROqFZZ8H3cPdr
PuqhZUSS8m3t/WmN2Zs30HEoAkb0CADuTqmfqIXuUKpwnXVF1UZomTdfwI54T+sP5QubP8yW4w6W
Utl68zyGcNGhj0zVvBwUbqmw2mm+v2FN72bXePpkB3o0VfvNs9dFoet5giwzkvU1v5ISAL1DDGHd
eCZh9bDAD7Mfe/bYzKtyy4vWvutTmmwhuLGYp4Gkiq2zcOzVzdqloMbELLmIK/SoVV9O199AEMwa
M801LEuY68NvgXnWOgdllvqlb7TnLoRJqbPCFpdY6Ku8psaJy82oRx74UflalT7v2VEVn4RmBgW/
ZugziMjwnT7jzu8O2ArqjU5TFnDD6TPebNJInWjNjNkRhxu//IhdQ3TVbnPyjw/iX6g37A+U7gCY
P8kd+ivI7fwF7lCm2Vn6xd+ZncSE0n/lSWHDVGkb7/TIHnUMKkLA4IDeud41kF6j3sAOoKL1yzOC
QjhT6asod+AG2U8qvCrO88jPfAz4RbBzXDIiB5Xfk2GuzW4gdM48pbnEa0L4x2nTTmMGQrxG6ABX
PrIQnBFrR22ohWbuT/Qdv9CBp5dqMB730cPZFbU/TzmuvddlSu0Y6WdKHXIcajJuJ9+wJdClRjJF
lTP7q0pqFy4aGqDwPYDawvQGo+n3f9G0angK+onjMo2F/5NdvVBlzEA9vuVhEV9rSBlLvPyfTQjC
tua0/k1d/NXoFDW/0KuRUTMbAPpTH5IEbeg8hPVamrM0Ll+gzwil/GSyyNnXfI6We0s/pewlp/ST
/oh+pqt+pXoLgAEIHgg2DirwSI4YU0muxHHYLfovScfmm0aNHUhVG5ws1LqHYveKkyE9g0mklalx
Eo2g91bYXRmSBI2dRCHhQZE9oxOKdpwrG2zgIN+BZeflWsNaI2/hSPIrDfNbMm8rZ8zSU+dBoc5x
4wMgL7VoQ2R/OoZApz7DmhdPBK+R514B9wzlA0dn8C8U8pk9bdHn4WY+7vjw91dHNb5QKcJ3ErvY
dVaoKrIUSaKovheccirRs4kxYsK/GEIh7Gq0CWcU1Q/Cb2l6haQuI2/OLArP8POfi3L+f9TnOwCo
z3ODc+91iLWr773cBWZfi15bwWH2bUucCLQL9diLdXzqyVUnJ+S3Akvr42LsAIJtInXxFd2SPDCV
ESe9AZagrCxf8nAVEK2tyC7OtygvUDKTSWYtHp/UWjZn5mlfsTsuSC3y4bK8SiapbdWEccvCdclF
9Vo3qK0W4RTnijYQqLuPktGJrhlrUphEu+AzqytbWWZ+SQPU1mUrOk8TK3clnD5QN7GHdM8I+nBE
b3+tDSoU1oxEfhvLvnVRgQ/rokkU4uCXwx2VmaOsmrsx0xL0aMOkufSHeWnRAOyW1G5lu8PeelUO
rd8p87E/aEzbMXtYcBaxgEPi6LZUjmzdbBxnvuLr8Jp6K21pBnwU5oqgNBgXFYeiFahEOGmxtkyf
vAwP84jCcVxsF6dwHt8yF0yRtQfP//3FHLB97K5FzRdTfeDCtTKCkuR+9SBHfu10xmNnKa6Qp9D7
kIr270yNkfKbO9D2QoU+HEr+eH+9o4Wrx/FddkIcRf/AiudgBWmAFy4Ewm55qkYmUqnKaco+KjHr
w4mBWBPS9q7lRzxVJyr76X5pNeQlZPJm3Mu2JFwYRG5g+iY88N/dMELbf4jszppYewO8aC4Ibnlb
NN3xYX+jCEVUP6sYM76wG1ZJZv61YJdoHNksdABbfEoY33UiaiOem6F2aDaTmv+ZYIUvzADa8ORq
IOrgr9iJKITWd1uLcw27PgGLzsNO8mMvHVq8dd6zsAHoh6NHNY5XoIPwALY+ZbiXBKkTf8jbzcy6
uC0en/RGp6PFZyzASYDxmnK0SvlKfHgyCUBic2EoT9/t36NkMAmo9a1lPPOcHLLiXTnmhYMA1+Fs
4diy3P4dQm4pLyXGpHTdYx9LPzFXyLxSJ/DeX+Ocn9DTBAFqKN0xxY54IczOig/pc+kQJibOs7gH
SlPt9xse+SjoNWAYzdBnbHq1CrBln1kZNwpqWR5+yrATCtE9h2o1NBKZTKaqFMniJUtlCQrTnkTy
R9K/ljmdpQ/BDCmpTMLD61HZnKCj18jD9eAURmhLuPDxINOsnMdo/8gxyCWA0Om0q0T4YSfN1oFI
oIlzouT9FIQ+kIfOvqgCxIqPyjY0Gky0Ln6v4sq9lMprxW98Sp1QI0bFwRJAIm/jcR14uu6HJYB/
FKCiWt+eMuU0cjUw+/UDDnx2q2xmwdFXBWVRhM7oECOwftxkydgZn147gJC1cahkYyfna/G2ZE8H
bbhfOKFdg+MoRv/Mq8+YzAqIjVeyl/PQ1tuiPeIMzU+VQ3PkDiMwM/pzHVgQgTaisWV4T3t7W+nA
uw3sFHkQLgEYSi0OZT+/jaet2K2eNI2dINzWD5t4RP45W/6EIxW5N72ucZr+oY4gtte7ijszXmvz
9NjS/Z9nx7GeBe/qHgr6Dwnbq+SIeObhVUnKdK268AJn1eYvbHTGMsFUCASS6LxImLayGHLhhPa0
CwrA1Lab+lQmtGOYOLQmDFcQuAyhItYQ9bg8Oyo7J1CZSG78Bkq9ok/0bhaxJLTeLW0/hiwN5Wz2
XU1HeqHa07HmgB9VKXp/9hAYJQ9jwfCqLg/B94ULdvfphcX3F9Sim0uZbOE8/AtZaRT8zvj8AiQy
mnm6bDeNED/rYugLxDXozKHPQ+gec9wmCjhRb8miBWN+3qoNODsXgf9Qij82FF6qYV1++RGm5Sbp
oP5KOWDe63Y6ZwRXEw/7mJlnel90A20ZtFirI2OKvUuMfcZCfrcYOuG1pHFEl375jqzxo/KEhnMZ
fkbOvLpyyKOYv+ZJtb4r6a/WnBv+rsJvKlWcVLlBqElHWH4wqsxQWr9it7LMS8MaH8IuWjIPlGOR
5Nit8Za0xVfIzJslG9MR0xjHgeiG5XbzHqVVTHbLw6myGOyAEKoNxCPfhGhVGWgzYDzBXoTKzrP6
y6rRroZsY8QpQs+hB4Kghi+J/ynNpGbGMI81FFOTSy0hVCPlMPXjvYMG8SEo5d4YRBKUJzkRlASN
viJUJz7nu1YE7zJf6+UdrqPUdQ2dNHhkEbD0SPk/LQGoi+LkU7Rs26WB4+yQfe9x6ssXNLtlLGmM
nhkFB1whzcIkiwqez9k8T+62u43RCeQebS8CReJ9QtTkh1XaTnpdiYflddYKQXIkYGB05+wXiPrs
NpuNU7ZHEglkVoslh0vAY5uz2nIeCo1/tOzkkw/qgCzTqatcjCaI28FMhzqOBdYSm4ttlfNgKkRA
j+iskCXEB54RXXF6ti2JpYlMYDrHLyl4z6iLpc6yUiy+kpSFvGpSpcDp6yD0RxFmpoQkXZmpcNFJ
W0AK+1sib46gg7vB0vm0lubBWj02PycV59UbcROKDn4SdOwlO9hSiF1U3qdFLPmCMmxQ/TOvvtTV
ol/3gbUGEPpgQeJruRmERpHUzzULp7e727e+1iOv3tPauGaY7IJVxjc5fSlYL8QQKhbJM8pwK08f
I9tBWHJf7tI/HuZZLD1t6DPW/gS4qHudVXbS/xvaHXLA4YfUVB5r2/J4SI0UvpfQkk39Ubn16TII
NAW4F0K0ljuzlVLosRF8Wnhr8s6K1+VeFbe4+wvof/AZaKArisKyLvjl8ieSAaRPZIz2R5HLWmZ/
nipKFJFU6jUXiPMEGh/h4S5GcZ133yE/mHboHi9qtyqM6WyogM1uZmaXzJTPCnqgyliBLZbPmZBE
XMWEclfYY23rwjse2NCc7gxoUl9zm3Z4b8IeDILSLa0XERlvhO90g/YwLIa+yBYk3hEp2UQrTsI1
hxK8/I+/F7BiwyQvzDdtxYT2e5vfnSs7Km2dKsgDFT3XCSBE7hvz9LAR+KGc3kvOZmJgtgBaexgm
Y9ABvpcSmoju9PD20tQjHGO3iJP7Cyozz62j3bmCymkyOKl2BpV3/4NdVm8bTuMucnpR3NjbErJ8
sXAxLcU5HR83BsKGAnlC3FXcHoCZT7HUNuc4BqFEFPqUm0I6DUAcNYWjHVTytIXIHX8Dz6Evohaz
C/kGAbm/1FkzQOMFeIElJS8GUCptvIXMqbATUEeL62H3D1zXUjRRZcl5wkwlaaqGVbvWtQS08Ztk
dnoqq3KqVB9LXC9DriLpwqeUVjifNUL93Pd8dPIebxJtMJqScMr/4VNtfTSgJaFD5Sl1kMXgoo9D
Vi5Q1vLz+o5OB7lwJeDIhb97+AlLNgCkphluLPbb/NE2xE8lj31H57xRLbYmBNbmPliZU0OEZ8T5
mST5cNY6xWzgo6oW3CqhbV4qdRmkBzKFaF/6D9BDKv+vBamkgbDQNakEfPsL5gRVPcELuXPj4XqS
vb6mJyPH6c9TuS1Jt8ZxLNzFQuUZ8qG7ukKPZpSZXnkAzkvcIomkxkHyvF+I4LZYI8FhT/hxlha+
kPVtpEjuNsj+O3oBdFAfVtJG95ap4Oboug4hZPpxF/hZOWSKjLfVkmHyLgvPB+O4iK6RUHqvnyjm
ZckMLsaBpSXl9+sAtoBuyJvUUGGvOsQusvr5Sj46NUP3o2iZeafpSNVXmRjckMM+QITKUkd+Alk2
V76uABm3Az1aZNkKtqcEUUqzw232mSaU+8xV6FahUN1ZmP4FRqF5EKYD0YhZC7IcXNySOAzbpZaX
ZW5GQIloi/HCBV4APy/hxZprIihQq/xhudt5ls8tL9jnjD1k2tEpaEd+spiw5Lhj/ybIxUVyduLg
adFi3qEbNQxaD/jXfqIcSEpgkDV2EmzLEArVaHO0wC6C4s0tNcWBDDRbtHUBaQ+xkX9Zq6mIbBm2
//gyeAFVEpoy2bg9JF2M7duFCKPZr0wfF3R8WdfsSjw/wlWb/QNTB/cAV6UfKNJJ80+Xk5pWYQfw
bn7mKij4139vCwrpe3LRxhD4O/Avy7uTkLmVu94bbZniFGRkXk/JtAcEQponn9U1eL1/16igOTeD
fB16o5b576L1MjPniDUiqXCPJYabOXkAMQNpaDICavcXPk05905NDfVhyDa0KD9nqZioZN4SYJrS
jdn+UMNjnbMKSUHVWxHWu6UquFZF6EMfJB7/n5hdin3EAFA6yAVkiF4frLe335tkwHVniFIIz5Ec
+KMWSZvZ1i/cJknzAD7b08SpadjK1B8oGlCAknjifs3wvzdrsHlIU0zMID4qsYcAysH6mVUceLpc
sK8REm1pv9t0athLhE46awM7LaHTWd5bWq0hHy95iO3jBq8TqJvwNsAiim9NY5+rT5Me28g5Dfbj
xx2ntJRHGo0FaWTsvQhY5D4WIE/bqz83I1BrM/Ia+5YCpiZSCdW03fzuPyvIkv7PCVBjDUOpkxLy
/k+GqHcR91HYrYECL9Y5AbjN5mr2dCAZJ1kjhl9Z/0NZxwl+ap0++DzvntIAgDV3mtqhv21+nFkE
mciZ6X7ZkYvfYL7c7LRX/xNrD5SP945qTpPcH2gmDCP1X0hdWzhs35I4iwjQ5ebxoqNWk4xKA8LV
Q0OUlEh2Ir4dnM0Q7SbcRreK5mva241bW97Dfsa3wC1fssHMTOrLzv4C3TQyRYeYiFn39gR8C+nS
JdnUgYuyYEGf+T1kTGOnDZwtBjK1CSpmNnTzMPZpWAbaUsv5cBdn4CByi6rEBM0lNyyLGah/8/EJ
CuLLNMuTeNK7k1xDUl3jXMFmt+K2wUy9XZaAYQcrVEX8T6l6Mbq4Iu7bg2mWsIZOJEvkqAJY99Ph
D7AQtd813AkQ2npoCJB+M7sdBH2Nq8U4WZHoMsy6qYU3BQtLbAcwBBUGgP8MWTCNT1PK1IvfdJm7
ZNii3Jv3IZzV8HKNY1+rCZYyBSM6FFLWy1kH3WUkyPVmh1HIbRlqjwCFuNQ/vq2OA+BEEUV/ykGI
23M+sE+/d3p9hJRC/UAP9j+ziJp70qQDA2l6zzcr+zwPWxR7DXjt+rI6J0l9C+ltRr4KQmWAmgZ8
BJROvjkrArhvR9Eq5uskND4PvXHn0I54LgmK3yGs9XPQJ2e2h8Tu4fLdchIQkh/jMzqjIApXgomt
jdYgLcvl3I3ybIN5Wtgq5tI5pj0qNaFT6blQEoYd/yqwGIQdMeiwUO1bbw9yIm83K4umLuWVVMLE
XS34hU/oX07UPGehER5qHrJWEDuzmVyelefMcOsYAo9Dn7oavD93J9NrQzpAgrT67RLtr2AwzWc1
q19xzz1fcDZiWO4NpEQK3ytYicnvhBrkjnvay+ZGXKbDkpYNsyvOXd16in0EVbhZNrNDrHU6onSJ
B+FjXjhTGQI4Zb6b66XoLK+L1R3o7lM2OO24cicHY61kF01QtrhXE1xoIEH6bQckmDBXPauoCo4b
hIZiS4M1Q68+9pHOH1AnmclH/c1z9wiQNoTSMvwMqTQ7i1YsOcLju8xqvKgyZpdCXWruK0D4C6vU
oFQYwH0hYJbaAPe4RYDt5JMkP389mIcZ9XWXRuPl5/7cTrgLHtsahQX9OIV90kpIzH6Vj/opNW2m
X7LaeGkFbSJ77mYoTGGTuf9L0p4RCg8xiCzKjfEW5JOPjEVisP/8DZOHCQybAkeCaaxTcILq3ny2
Pty+w2bL2psLfq7q++hEb0vzbO3EyAlBvyvAGNFZ1KyVaNBwUrwvwcZBnqXNaacL7nByaefUNPwx
x8b02ipUIsy6igszZSrMe34Kr24K8xVzM6nenaUDxZ4n4XUTQvaHoixJLOeWY5LMGfiuOpDAFELP
7XOx8vGGh6Bi4H9oU4WNQI+IhaRHgT+pxp0svAfCLs5bpjI2fe1+XxbMJHV+HGejIxcL/eSSyS4K
SGXg5iHlTCFRHA0WtR7zUYXMpxy7i9mNYqQ+D4DW5kOy5vMmv3YFEA2s5DHURisIsh0IpaT8Bze5
CO/c3mlm5qJKTwEE7g/COANi3CWDhDTSAg9OPc2DMg9uYRdIKATOoEuMCJlURfqJ1VRnLsv9ftGB
ZOSblSYAosNTvG4WX8+3xaJgg0s4nUzpfVHR55TQntCRrCGaKNFPgUDxdF1aui4H/rAefYTvc8SJ
Xz5Edbnd1/w2OTuFPy4Mj2R1Qqc/5ydDr11/aUMRxAuC/6O9MJLQGzO4LCIyahvi+u3rLrrPdYzr
uQKbw7aAqbalTpC1FCzOMAv7dpYGper//qMCtCzYHTGE81+vqBDKulfkrjD4q9mwreYpXzBRklUt
5/r7MimfKO4r7hlIbrMrMK7fM+FwFy26tpIr7A/jKlCoxG7CKwCVbzXt9h9MCMvkrSMuuoxUsMEj
pbZSSzFoUeo41Xel/T+CVNy/u4esO5nBCzS3mgv8RGFf2vFAEf5yBByXTX90WwJJrUdyhlocxl9Y
0pfvx/38WDBn32nCnI7yfwBD+s+u2cGBu8cxJxCySjXdrIqzj0wNza18AUI796UWZeXn4GHYUvF4
qjLHLliCJNQ4R5HTlQXKZzJoxCiVb1dR4P39/gn2CfTU9jcGRwGOBNIzirjJioisOVSTR4tFwgwN
zEwL+L8AnTdFIea4Cx80cC/w8tD+EAv7hxKBljUIQBGaggu2FTaVyHeZTfOeqLyoesSrzQH7av8c
DRRbMX6fLNabI/5gHA2S3iYz5cRZ3HnPPXLM2PiQMWNAWfp+FXJRd5sGxdByC73LFtWknRnt0Z3A
8ZsY3Bu8nR0NNFMrZkCSJxxaemOX1iPc6hnNow0AwQ//NlmY2fTwYrjybwBI7n9Qf4NoCdWLg4fO
S9s6zYv5Srbf16vvhx41fWAZaWa9fpVFjBnz9xKo0Th/dwolnMiG4q9swQC9HRwOtSDYn+SLf7ha
IBsQKUCcCmyKsxyAae1k2pyKF7u80t/q4XSZheM6r81dlg5WMtLRkdvm4YEA9ISA2IvemhxjMOsp
Zo9p2IvG/+ssQR3maXt2jOj7URVCAtEEsYLbteq1VQy8mOB+itf2GCOsDOTt3uHP4BOL39UHvBDa
hV7MIxZqHcQqdw5DHo3bxSw8vTKNtAnV2SCkPFH+KjHp3hgXLzEWhzgiw48bbneKqCAKg+/syWhO
8dgp7SXmtMa8DaFqPGYXHf3JHIJaN3vKXEUM23JgqhbfS+9/XlFfPbZSZqW772rRNNYcLlkRF4VL
bM2gT0fJ3dxPSmOSKTu9GLV/fT6KptR3RdlWDt6ZzcqLN/gJijg+WigSD0wUDvWWQIDvODqD39py
nrS2hcH3+TrxgcqyJ/lwNiJ3TdoqHhlLMwZl1SrQYMTwl7IIJDq04IR0rajZxZu1Ai0zXqwEKTXP
zjqeaKJeSEOKxisXirAF8DY5FVJx8E8oX1UNdK13DclqZKhp4qLo1qozl/Xnh0RjVuqaQxulsyN6
DEsUjzuf7ZwXh7d7XwC6syBvVWreP+clfxhh5isavuBNRwBYK30NtPbUVRWZX/TZI0u9/uKrs30U
jGtzk3ng9AJ3LkLXi2w1phkRVpu/vyPR2xefbKbPHfJLeZYbhsdPMykRK89jJlH+GsC42Exypazv
whiaETaWpvvS4oqIuMKq91TnAlhgfeN/DikO8janyqtHbAqbCXTZWr3XrFil1XEL0MBZzdsQJRSv
yTD1bKJRO17fQfik4lXbWUwuBeyBh3oZYSaSPXQZT+NZb9XxbVYvD6rL6JxoBwaoTqU1VqN9u89H
kP83+hdUOBZA38p3WChMrj7LRdHxnBKcidWO1s6c4KfD1gGF9NZNIKtJT47pOScXdGi9narrcBSZ
UyIgW27S1Nj48ZfZB30qV01eVTjSKO6NaG43wZn5vZBYolbcml11VifAO39zoHMh8jfviurVRCTs
XYW3RcFawI7B/9bJRmwy0/ggjIIcb6tU+/2oPSa8tFQogVHb4bGti01VGQy2uWmBTpTR18xN14aj
fXnE0YeyQwIU6kIgckJ9Wj6CYV6hndxPbfhQVKWyOp/M/HYWB2mt9p9VFn+3OITGXBRJt2c2II/+
vyjPMO3T9GRGHVHZFDzEp0XSNt/bJRuUF48U5I6H+mgvF0AZKeG03gGXGVg1hLG/zZ15kmSPi0My
PvnhNNo2iFFujIIWryLoUv9Tvk5q9kJEmGDM3xF8LsvHAoJ4TxS92Pcg7n4CTT9jRGyIxI37rDCb
ahRHPrIEnQYexIG6Eaj4R7Qlhu/Dp3XEl2JrVy8kg7WtWiNhsX1hzeSrEvdqeDH+HdJ4nFAjcciD
TGjdESOSw58TPo02Y6iisXicjoOKIgBzAEQ4OMbdo+yBzaRRmol0Y7F3/qZrkFeUwkZYvEtK85vB
94lR08DcGzeNr+iDCTQWfOhGRKA6wFW3VdAPB80y21E/nmxqewmeHZkifCEgvnH3JJBlVNRilFNm
JFwt1ApuqzTAgd+S/PqRFdcMfG7pEx0naIQj8RdJ98RdUil4C6uxe2tK7flLwAWO1EQLV844Derw
5TfRk24lAkuXtX5nw0RoyYw6eh7WDOTS9NW5LqXwyXdyMo7dEHHXi+i2dB56O66CRv6eaAPmQCX0
6SsmWH0l03MeyedtrVp8sEqIbIVPp6huYB3hoim6axLJWYjDaYQfHwAqj7O87Do4llgsqDIVwsFQ
JVJhDd+vhymKacgsub0OfEBZUvpyw0NM1TxYOJxVfrGe1wK5iTIDQO8nyev4ELLgA9s0quLsGT3O
j/+jQPnneUoRMgEOajOmgwTbRVt2EqzCTz45J9IxjkPKnej+99e1neTO1/PLPEa+NJrHixCeQ3jH
A+k9oIf9Suy2Gd4JvOs/ynEGlMUJyrEZ+iVBPQNUwOaTPT4me+FX5XB1HnvQzs+zCvxF5dDRAd/1
NyWaupNoIqrOQaqAyRSbP3aKm2bwMlFto6LxkGBZ9XzIyZZZjNheGn3EpjAzt/JfTe6GAGthuTOp
qdJ4TBhSMxyypWO/HqnEmDFfetICsC5rOF+7K3FoTstW2oMxwRQPu5loCIsHNhvQGqKwN3LwUSYI
He4duUM8cew3ob4+ZClbpKUB9Rgw5ivrK2mxCFLxWmFWz/5FHNXVfzJRQrTv/fsRmkX+AXfV5SCs
7z7dqm//UdA/E4F0AWsOMs6zzWMEMi/BYF7J37aNR0+Zf7moIaNc9LOdLzdhzv2Q77gnQ470I/J1
l/W38A10aASKJbrAi323kqGkJros0iYna3JlX3Z3VL4RJSRvThWb9gqHfpB0c1Rt8rZHsaIME5h6
V9y5J2R90gqMuatIx15YmXBlNYY2zBBAY9RPJoid2CHepvcD/MfMgoZu/lv332cVVnwF+dPTb/Jl
0uQ8rx/40cqVuoUcBaMECQ8NQbMCHK5qsOpahH/12yBNa5m5EQSpmtUdTd1frvN0lxlVDwswERdT
9dQGwERdR5zogTFFz9l7oH+jkVODn3JPdjng4ymYKgKISygnVtPNNgwe+PtH5x9MxKaIwZu/K47J
J91Yu3UYKa4YWMDPQVFNTGC6orDU5IX/JGu8LzBTWrQmFZH9tdIRwYDMkIYxYv05/ordv/XpYieN
7vUQXWvbnucANW0mgKAPWbNRltxxkK+L7NgsWroDtXEtFoR5SLtIIci33Yp1zyvxRhDyp+do/U3U
kCq1hVHhE6HUt2orff72rrABcY47SGJkcmMeb3ptWwYwmcsfiBezFXy8mC5LQWU3QPLKyjY5nV4S
N542ej4VUjNEzWGfoFxh4vpmTyvkSw1Wna4EIb3C4wWYJ/Q0eNQdN8vuVeMu5tSdqpjIM+tLrUzh
SUT12+eIEqrwGuFTYkpnYX96X7s493AkvT4noNkjXRO/FAvzfhBfhtKkrHPwDzdHt+X5yeX70+f5
eOMKDRamFgbgIzRWzqyywBH/SsWjzDDCkvUC6RFyRV4UPfSHW5JvHNTDtf7lzw2hhnsOJeYrg3UV
dsRcz+umtqAU/+EADVGnnfbSj4eSS5gHQCC5gz2H0MkAlGGX6y/eaV2Tfs79xMp+Op6pIdfHgog3
qisOrlIZWtr8/u9OYoKndeTeQgCQbzRag+j1suW2h7azz02jlsOWpNHkxN2vlq8jraoY6wC6VFyZ
6zZ01WN1Wiui3RVXamAAGSNBmeMiY3qsBCqujwPEBtKC6yieSjuAjAD4h+mDkWqnU9agJdfGBRLA
xhQGfkzMmOUwYIFXgSjBHIgU8uC8Y7u2JVd4xLjbWLTSL9+gVCqMfwOCboP6Yp4pAQcklH44qKkP
tcsKLqtXmcMt2c6AUCRa+nCmPaf1Kv8U5PUwcIVcNwNqnaFVBKxGRqJfrur/YPJbQR8oYGZzpHfX
UGMdK0/aYOPKxCArp/yA1slMQLCUz45Zs2tQt3oLluHfTkxD99kEL44wz9RXzBkVYgA/oQoBJ7M4
64OUPbLJrcGLaDgbwHDd5BOi3KnEpyTRfMFiXCLSnbdTVRXg6Y68Fi9J+IL3Z4ZNmBv4IfqYZc7E
RnQYR1nxRdvCOEd8eOX4EMSi7U8AcUqY4RZLPmWkq/3bZtON4TBZtfOgXQcuKTOAtc+1dv4PyR6S
/H+dDNEjjZKSgxBpivjGAfJRANMRonpnFvpHf6PVdWtin24EP49dbmITkKayuCF8qEN3uCwg6PeP
q5Lp7SrZw+KBQSfXEWho7oc7woneLkmkTe6dV/i2DVGCrn5w+UBabaQIGpE29DuDNwVWbgNeu3Es
wVM7U7btrYaWxvN/xFxzJDnOyBqBgtOTbvGlUlViy2xCy5nW8+0b4t9uacyU7PPi5gXtQBVJ3arm
pZW1CRMYqqmbCP72dqejPtZ4a4huWE5lzkvuruBfAIiXKl+lPaJhmYIYYlJnn7fphYjrR25SnsXn
rAB9xIRu2j8tV6nH2CnWgYosYyJ57A/QYDuI5DtVQYdb60n59NGbuuEKHshx4o+UkOGHsgw4zTZc
+9EWRMjINu7HN+Wi7rD4zSlLEVgl+zzblKXAxevHuudPFcZEJpDPB+p5cU+rMf8SRAn7CIxqjwWK
2FuOTFrcm9XOwodVPSwwP0E1JSWDvnh9Lrz7K0xY9ySwYC7P1dOaY9uJnDevljvjeh3iJavRtLqG
H0YPaUkvmh38Ox5ZBfiHMOqP6UDmMYppXMGnPUd9QwLOquRdKJPREQtNVuR3LhLnEqpvPmLGYthN
jLiq8DIp5aUBDJ4WMHgLVGCY5J6TXnDG0qHEUqES6byfG4/4IRS73TOVJmgQz0SDLY0RVyrNSPl0
Wv7JUOrmiV3fBdXmvhrZWwE0jNkkdX+Sq/TV3pGi1jbKgYUldVZSgiFkXe6T6sSp8HL0cAtfJ/iX
f0C195jCygYkECMxI87JkScswPhWUd6HZaCbQh7Wscg0t+Z5AbUQp73tD1qj7T9MWSUnUFRt3xAT
uwxHx6M6z+QBZAHLC0IrW7cZMCvW19hbJbCVTRIHC4hxvrHfE1u0K43cZDHG9vjfnBoG3U2I2Lj5
QYNNX1a3F+224RduMgvPYysG3pobMsJQv5uNGcYeTal1I5x0s5uoz9n7jQ0nIEUxChdVTqVREoGo
TvynKrmoT4yap+CMvpD8pPxMQUhBFp9+zTqPyr5KxrSUpx9eKZkkp7kLt4LlxkQFU7MH0e+Ngks4
JIpUkaHPjx40AWpsyyDzCGPuPGRnin/g12z9CDXo6u+Q8Y+JK1XPTmjASvu6gGOGjudVMcIHf88c
gzR3ujR364EhOG+OyVk3WO6QXV4+ajfbyM1BBCDgDux4RCQ5fUFxsQsebKgCqgK9TozAcGfZ9vU0
VdmygAzcA33o3SGamgSyUInR0YwXFdai0GIbzTnAhLfDpwmCR4JFVWDMtYcMEdcrOJEL1wtPe3B4
wrSn+AK6sdtTqJhmrVyAxn6W5xBSy5QckFOMJTvw31ZvStNExzzKf/TJIoF2j1vx+01E+2pe4kmR
0nbos6ws9qnk+KP7hiP9/SQ5AiA3pNVPp4UEwkZoLiJm98E6HYGLnRYFCBpvzaREAwYW/l+BjrMG
gWgdcJnxL2I7PoKrr6iE0WkgYLdVTVZp5O3IXaZvvfc+m7O3ousX+iOMXieWL0YiFhHsoa2yjH8o
AR/lcI/2/WVAO5lpp+N9cgWwwc/9B1GI6pk/+M8E8/WSE0lR/Z96+ABquoaZsDvFXW0AjWHPCVuR
OH9EI9yVEJYbl9R97AdxEfIR9V0kzGnKSYmbucFbjxXaXGsFd0FjQ2PMhBlk9nvIagV114VWV1F6
xx7VQGj97InY1j8Cmap3GiJwn18jzgK+4qxHMlAv2wdu5h5VMJ1V5P+S8z9YsY8GwAX8ewTabmcW
hJmd6hJZL3WAFiMwlKhreEFOXmOzm7TM8dh6rhsavBuJY2ixZpreaJIsK+9RxKEwxchM8UzAgeAJ
YOWz4G9Ry8TXaKyRqmZdpi956UgTGDPkYvMchS6B3dRG9nH3kw9+2Vpa8n9gURE8D1oIT9LtLOlH
JJJfr/W/m8pPTpKVxhFcijDep3c1eKhdcsE/v+1C99PyMeE7HVfFuTnQaH9N5noS9STNml9aEm2a
3OlKJQCsDFlXKqsYdr+oQrmD3LXk2lTNXl0M37SIQyGWJSigxMuBqJK7wR92FgBgEvJJvP5g5tvy
thav6hrGfH1PLHPvpl6OkSs9CexDSTBxS+kfC/74/bV2/dOgRK6a64MZR19Ul+sACA2/ljlrqCyO
ICipNb7ncYXFcyCCmJfLenIcyqLWHgr0jn32SXLsonTt+uORe/EKkFBC/kCymMFcq8449WjH0Z5b
ishoavnKr6FPVru/O5iv4RRtJPE514gdl9o+jLKI8UErKQiOvSI0HNdmyUqArx3c38WRh4DInReX
njhT49lDyMxkE9wp/ZyeeGMT9eLqbAOg+lHAO0VzPkUjmRCtD4fuUk2BLZ5D587+toM2BMMdsrmD
emruZFekatTMsFIqUu7vzTCr+NIEXkouLflx7SS7eAezRqNwAOGHY6LO6HvbSGJXKIb9bvfady3/
DkdE+KhugFiXehKrqT/P5IAsU83vTKdvt/iodfh6qPliTHzkIDkD2S/d149Ldjdtrb2aXDTu7Vzs
DujXnP8WBdnikneMxAYAO8fEAtCjdpo5X2j9on/xCHGbzq54l9oAIMMQQQi2BgCx9YWcp53Cs2vS
mfUE7u/nONj9vMkRo2fKR55NbsCp9f/CpZgz+SMlyeS/+ufLFBuFFjmbE+IxCnsPQ02xgrUUjVud
PbqrALC1d02D65SZzl+aSwjCYmPFVlQjB9+0JbCifr2K8d49OaVEVbBXC/WM1rCtL0qFWk1PZj2a
eXOVq2ithrENoMM9LX7EzLTTt8GpbvN0lMVZAF1I7C/NnLQHt+xdZe7fdDy3zdEmEIRrG/5zfPPv
Qinha/Njp0+eaVdGCqpkyiQTbnnwEwwxOilzbKaFIa7Y4OsGWqzQOmHfbANVAhAmIU9eOo+DkfzI
tklpD1FOMb5KMGUNAgCbrHV71rVrpSbWXja70BmkJ2BGMg4Go3M0AbSrw3Z29wHCnjwDOWlGTi/3
aYPaSMYvMkk5WwdPXXFjLMXMajlbqrqA1/gSVvF0I4BujbHOkM4A59fD+3lprPsT1CnZhQ6+s9yg
w9s0vvOOkAh2x/C0tRtEdO4Elbw+8LBtbd4vhdV423vke2mXfQbmsPUHlvoh0yHA/kf9IJ6SSAt1
qReufW0sWaBdfu6c7CgZMv5dJ2Y4E4ZrpBDuLSJvdnjB1bQgTrcyZYKNVIjjatkAO1H5i23jtcQR
lEj2hAOIOckJGqvkj87QW4Zb3+42JIDZvzYI/Rcngc8MWlRVYA/vOUg8T4oTL/otLXzpkB3Nzem8
xUFoWUFI7sC1/S8DUhuHur9nAm3Rrij5QFhMPeV1njXaH+xRywnxBdTUiZqt+mzSZFkJ2I3sCr3z
oEa6Gn+nZcCVMIc8Eadn4iWE2wxCS+18Rz1jEz+d+6QmdtTMPGXC36tCKl27svN6SFW8Jcil6k5V
U3jv/cFBqpC4ioVg/5+YmC2GcA94VAXYgthz86MVg17kn85rzeKKvg3j+sZcujZ8PybDj5ty70ej
M7tJYUFJ74oXvc2+5h2is5yA2cPOIY9J4ErB8Z8YVQW2IvSh2fKo+Cs9e5kb2SWiAk+YqulU+MvX
gpfy7fPOYuV0LbPFZb7m/R4yP64f3JrbzQC+v+jHPDCa4DiV/swHHO8U6oS4mzp1SPKiZpTC2usN
cW8GFKcbRVslVKbi/sTDdIxBDpotbqEvsWZUTCXh0FmRkyiSzkD5nDJnR2xSuQ7CMESjShb5Hjfg
AmruekPxSFcYXmUyc5YmygAx1T/iac195V5Xn78B8uq6FpWO1A8bFL5Kixo2yn3lebvxZ7huVJ3X
jOENrZOC6KEflY5mNtUQrbPV+pkHn/4O0sHRaX8AREqoO/TOdvWuOgt5gdVsz0cT2u7DO778N/3/
bh3OBMa6gi4MmAIGqtmpQAwN1KveJzanRlKG2WWPPhfes8Z92sKgkXlQnNNlk+5leL+QGFACHlx4
7ekzjCrJXf29L7zMHRrbKtkF4l7awWNyRHfItjH/LLpxX3HC8gPmHEnJCoq4YB0FCDW/mrExbOqc
NMIhkS14zqb7DoOLEZ9Eb+VaoaqoelguvUs2Ctv2ZCdZMKK3JC9T4uceWkSvr62SkfyMLtoud8Ot
usEuGn/rFoTJiOcO5uwbAs+HOS3meMs/YXnRtz7VEoU+7cB4kxDEB+LtBu+DFgNHvUl6PT0mXg2V
12SjXJkRiSGXJCTh0X8soQI1+/1S+s4pIfHE0e2PMRfGVIi34fnR2RgBbhKXc3tw69VoTVvEePbM
NsLSdyVHRnpTtO9G4hZoaTy5S2eeQiak6bdD63Hvk6ZLTjFTj9RPduEkdlJFXs5cgRFeej7Ve2x/
MarEuYYl9H2eS2tyFId/jqmku2uz3QzFw/6NmPmD0QDHR2fCCa7qELmxy/5bzWW4kEIt9RP+4FLJ
TCYjNxCZY3kDwFUN94LNtpjTc7EGCJDnjs+pE4t01Oa5k9F2A1p7lZnmjsTMOJFEyEQBuaCGJ7zH
CzblLA83W13HsbGURWQ6Sb4hsPR5thyicUAJce9d7a4PxMTRdoOthuKS4fa1g/C4yrifP6nYm58b
2dLbGjR/965ZVVbz31PONxw1oZPFMY8Bt8iW6xTxvNEiSsHhWXGiZWjSTEpAguVlhMGGguu+iCi2
PK+fQOhER1rWiGAa5Z+4BkUk0rCFxCMXa4P0i7qkKe5V/7fvZhTrj7HJKW8mceXw4qUBJjxWbyvz
rizuoXfvwGDxqQRM2VmElIb3SdzGJrxMTf0Vg/H02Hb124/oRAOdbUIxgV3oh44YhUZeC0YadrmB
PPbp8n7DkkQ3OQwP3CBGxJu7Xbv2qTsO9RU8Ze0KotV2Ekn6Ix4LtzZHEALXvXW7F1cVQwJnRRqu
xS5ik/eCjxcPAGw3rbhBzmtnu5EEFi4oeX1jCYBlSnPgmM1KzLBykZ2Cu3dm+MPDZuR0mmWU+v50
xU37UUTNbJ/sQq0oQ+whJagCNXt9GMbd38QvLKk3FCU4NGsA2xaLDfly4uOBVoNH5vtS0n1DCNts
yuli2k/Q63lcXAOLLzvBQfNBuWJBGOl6KYsbHQaWR6fer7oW6t+vUHOmQ/+W+rYl0qu97MHL9Luf
WTk6cy8LcSsn9f7owZbYK/h651RkCmQiP7SfeBkDsbyYYtgvq/niuf+x61PidJDHH0QzxEhKBfUu
+1FC5CnE8mTWMj9CryCzQKuOtLHeDiAx6wqSrpoocw4PVEd5YL+IFmZNys4QuVZl6TyUt05t22h5
XVE0V/Yupjt8FkwWZzk5a883R/KB4hY2EpGOJKhILDGWYXE58O5SO+/ZXVGByWxPLWYQYLFiJk57
3eLUZ3Bl0j7bhiYsKiigAq1OBX7myeQSscBaODg4GvBJEjIULjt8ADhx0IvGeyv0uCcCl5bQ9cfD
LkPkIJOdCsc8QPgzbwYBzNk7vxlLybtv9UEv5EZb9jAakI2oUkXGuRbcqABID7PdBGF70BvLzAc8
ENEBNbcn3H97/41xCnXV12mQKYg0EB+wq+6aavO9QZQ7NeGfNWAxjcboRWEBZrS+iRR6JSFnPY8h
BY3/RyM5Q8g6XlrfuFJz5xVxTTOXgsCKxWj479yaPXmRjFSGE8/RdCJIi7TX9liz4yH1P0ucOnbL
Luwh+u6rvUw72ujrmz84LgclWkFUGFbct1OQUkzutTMeMxLwKZjpDh4YmJbNoQLhOPkMjYd0NRhk
AiLmkGlb/swwRJvbFNlH58vZLGfrqEpytxtWNKgqarRmMHSvQ4ADD0m0tZ6T9LSOVVpjEJJ8VQPC
wgSeceeoByquYhITfe+lwRWt0fQfZ7+9H+2IpdsIriyZgy0D1JJ0vNvYoPHNNdmWyuxAezhiuEbl
MquM2UCHKVFs74QqpaHNfnrY4OtXpZoEFHvNgd3/H/YlcHqjbFcg+EzHkVcu+Xu7JvahYVvc/Yk5
H63YF0MithXDeODaZXKwasTtbgvnRD49stoYCxk7fKDZKBPQHraO3oXOEXgPzie0/lNy57AIcZri
qgAQStV3smOJ37aBEu5uZpICwY2/5KYmuwa2pkOuo1V0ckIFHOz6J0/Xsu9i4IXe78mOkIwivdTN
uRzoS/ctWo/Noy1HAmfkQIRbRTpryB5l4rH0lXyDVFqyeXTW8FGsr4KyROEE6fNedxdyUss4f1B6
72z7WuxWTa665GAnzHs3G49GdFRCoSU66yb6HUqOtOI1bxtPGcmhtPCHJXezPEmVtZYszycYtlca
NeIlQNoN3jY9elcwW7FSMBHlSu2uMUbEUJ9ZPZxzUvQHZrOY8usAwb/8IQCxG9DHnDKnEX+dyLid
4vOb3gpbXimrytA8ikSHPzNeqscn3vZXHyEX+RFCboimEpJzrZCKRt+n2Ylb2/RgDmPrl/pOMmPU
mUqDBhaNcOoUdEWxptU1fLsBxLWLX3jwh2njiEfagnkBjg457KnppRqDhQofvkQUmxCnqWUwT/Br
ZWYQhbW0Qi7zlGBWWhcPTF9ROEiaNsl/BBQpiQFlbxcJMa/U0CZ9pKKmZT31kerwspQE1U9z1Ysx
ojR/IMCmx6UbkEMpdRi9rnO+Y4Tr34AMHBjbtLc49kWddNPA+Yb+z/j2LWcBaviuG1agzYnktnAW
XxjwCQP/GzxUa179Lgg3R/A3AK0a4bdKoTC30pK0hno4jh8gle0v80MeDMdCUxv/NwHYF5/NfCZ7
aKoXbQDnKAQK36r/ARa7vhJPv7LeYd01w+NUmttB/U0R9slwZbx6QOUuwWhGlUJE5b+LY9526TBx
Hb9324lZKozUUu1JDTri0yAwWxhPVV34pwUyjQ5TsD9l4iKYpviqMkSZIMBGbtzL1NwDZGzXLSlZ
R2lYgBEGcKe/oqg0zQdA9lSEkFyIQrkiFiNnCDpOwl3og1NHM5EWIF2E1Y3c2mcE4M/go2hzVqfW
1J/JjMcDtkaV/6zBYMjY3GUzLAOU9EUn0A/Bhu3kXrDUIq81pdy6fEwG2yll1dYOGCG84X5Sbzyx
I8J2JmcYD+AwNxfutIzmr/11J2U9TMrGoUJ5HlvyQiev6Wzo/P7SrkgxPd3jbqoxuFRb3p/uuZhq
Mf0oAJzm1fYuL8HutJiFUY7jdiTke+nTESR+5XiMu5kLlj0grSwpxrEXLKYNH9IrLstY7epSu9T5
YKpmv4jRNWo3yas1yj8Tnn1siNhZXxKAocEo/i4bJKZ97h/5wds9EpxyZzkrBX5J4glYFznAeqmF
BbMUG6r+yBaRKGSWMCb5Ti4sC5LgAGWiBQd3QbWuB3e3/m/6ZBeutGEiC94ZaZafvyroiv+9pYWW
I7IqhxqVfP1AgpRY3zLXU22s/xJeKTBd2IeQkKEpwNhijy8wP2/njRAjm7S6YGbqTx7ZrkKrm5G2
S9an4/asaUVcosfJAJvO66kqS73v7n3MSt8U+NHcOpVi2bqCAJxSN/sc56AM+jzZF8Qu+ZRZU6nE
g/KilSKrZ9EwuIfbEfeBj+ymoOQD3Ruf0zo/3XaX6+bNs/x0nx64fw01LZ+eNwKTFweRd5R0kIJ4
PX23zROnpjEWuTuHvdQQqjSOIgYsdTCfurG3EYIc0GteQnM8AsZEKG3D6xGzFwq+EKpzHyiJpe6s
b14ZgUDPmiupyKBIIl+VdPB3yh8VU4DiLiB8wSjbFGhvd5mA4iSAY+X2TuaTagDvorqMAMnBJaK6
kJoA9lGgP68k/3vbrH5FOqnsRMpBuATMjJy0kvWjxLNDM0ryay1wF6h2Is+qcvTdchehRwdRP1lS
WJiJ8yiabo/vB/4H0OsRUi5amrN6uP8qb8NzTWJb3BgwTZ2RAd+kB51zT+66K8mEFFG5LBsW5tpJ
OJsYP9e4Jv5Dfmggn2TOk91j/0Xj0zsIqkvKPy7e7CUyd2EsUGYcN5zHKBy0oADGlMEak0rkvybJ
GyD6Wm+BfSrQrEkRiJ9ERm1N4rS5BnST2sDVChme7O2i6aJEukS8bQufMMbuVpfRzPJK9mPdboPo
P5kqAs/zoSNqHAHq+IvR/YTI1jfaE0QPTsAXjPiUm8bjqBBKijGe0V+qXVyPEfAIsBUvewPANKRi
vR7gwsuwSsQnczHqag6EwOl9HJDo7Q3QYXEKgp5zeBb9UR9fT0VYnYGstSeUdr3vJLBUGTFL13dD
kvRGPsddr5Ok/ulQpHuRbzVHnkcDxJy7MqzKG48YgPPE7v+EJ/vLxEIV4Smzkji0B0Fr/h9awc9U
lxjQ7sY4tKaQLn3FIr8olFuioozlISRNTgaNTXaBaJ1loPw2buwq+WLuumKLzU+uveAJxZCY5Ymq
ulnNHHPHrdqLosR+SIJ3Oxn9dzn/W+ybFQKJaRWhvxddBGCiUhgo0GcOL7wAYO6mNZbcFT4U4hig
UchbvYSX8Z9YTcfgh08yPha8fIOapoyE6bXaoHXvQs4m6q/mygzaIbD4lWNxuYO3LDp5Un/+gO0Y
95Q/jPFrjCLXnEd0zMbxJ6x7z7SAJsrCs05QgSSc1u2nAFdPanct3T3p4MYe40SAlTnEWD7ZNUQO
vv8I6lEaL1nEOMkDB9tckn26fLBVoeDOdmjPE66K3KHwEKIsZ2nw0T24xOsptqeE7DyxkovV5nVF
7X08Wl6NC4EdRoNkLQTd+kUdim39CVHt6fSACi6iVlKEY2WDqKKK2Fsh4b6vjSlz+vpeuPfbjLZE
nNyVLzZGK9v1Xh01AhTMXUFO+QN2Mxu0sd2nbhMR2MluMAr9Hr9SeJStLjNgRDb2PHntvfRcFvfY
ct7ys766RX1OL7hP9eLrDBBFWMNoQg02+k6clStrVQdPX8+nTEU4xfNNWqbBlySAlw76cc3qUE8K
c7b+SGDhinV/5+t4K9jUHZM1fqAeCUi07klXzhto6XTF9ptrHhPknqL5HZ6uXu54INdlL1/lUmsR
3wDIo7m5da/c/7XONr+H3+7XYFN1bcKs6BamGdA3SZtBYjoJs0S3m6flRk2n9psMAOEnw9lYSesl
PmwsM69GKcmtBDuzEHWW+cHKd2MUbWG9ZfK2m+b8NN9aLawGcSIUQzymfOyIrxMBgWCI1f5ma57G
JngsjbWVlupbXiwfSI8OWucuCqPd76VZgYZ+Uxr7m2h8rwgptpuzOQn4fbhWNOhQZAlo+K7dAKUE
vWfj6X5XRbMpHTgUaTUCwiUOJeDhAOTpS9XKI8Q0xII1JRaaGsKePGdfr4cQ+WMzBSvclepovEy4
PucGnmj+z6PwYNcZwxGD3S3YnBcklF8HnxvlwDTeO5cNT9+m614jcYRNTQpdv/8J+5qs9v1lL1Gx
Vq5NwsiAXHor6iJWS5VNWyN5ILfSe0OuglDe2RlVagWLn+V583aw+im3O+bvBH1awqRlil/Us78d
S4HxsJTwbpfBMOBdXZ0cVQZ9pAoxDdL4zKx2L5sqPB5YArz/Rl9WNupLHvp2mZWE+7AbULnVaNyQ
gl/cpa95kV9e60Oq7TDqrCSv7Fb3xih9j32v0yF+werHWGSDnu9Tok4zSTM3TlLAvIPAFF4Y78qu
8Bpe/VTZZQtrk8H1Ij5bJyHoDyGN0kTkTwwObjVfsMEnEK4KAqRV/h7m81mIlojKIJLKqrOfex1d
zUs/YA25RQTwEa6dhFeBf4q+ZUpK5+bz+ap8oREVKHuwIYbh2L7cJ4eJlknd8ZAnocAdyeLqKZGr
xTfKfvSXEnuX2SFLJd+W85QAYfCxJCYEd+5Z73APkGY4Cl1JXCU08lpXlBmJ21fQBhiUQYiR9Qh0
0SqRVZUge15lpJONXv5jZsB2Umxh8icSBBlQLX0NJTItRG/gWcBwEGAHdpZsFBjxSWT1tC4xkgKY
SIKI1/R+mRadJRYodDDodeXWcIdo0i9SCsiJM7Llr3yBXjmgCHHh3+IcsL7EbkAeECHnPNW7fpRp
K0C2KWuI+tak7wvUzPWEextSu2Pk1EKjWvinX4GIBFOSVO4/psZ7ZQjSUbMiPJD7zHpYUWyYVS3/
A70FKGGu3AVAzt5L5zTA8qJoQWLi3Q20evnFWyYnlyLp4IBCKeFTOlacCeEvIoIkbIsURKuNJIP+
8QB6PRNX09sJsD/sI1Zmn6mn8pH865yac3/3VaXlYixk1nlj5U7ekUJ2gqxZx98mdJnEF5O2AW1E
Oc77J+KEkg6CrSWmd0HKxz4L0MnjvYcJC04UXAAFIuve23LYW1Ya6m7mQpGUv+CXQZ46CADPG7z4
V2gweDKWnBeMgcOVI0j+PJH89ce4ilXq5iebjKmkFqnsifemYPHs2Q6vjP+MJO6OPUdN/lhl8Fol
oGV0pfU8L2xJsVeho+8CkumqdofYofN12sAfRql6tts2Mcr3Gt0iVCnBHfiJWCFEPmFGB7HyMyHN
n8bZpYwhNmGztediCscI40gSTgwcpe9R/+usJh8dvJaSMS/YSKaT0Q0Dk5/JxTL/GnAD9IqEkB6N
YxDbSRtEAtHY3WYi5zaoZZcWhb38C6IEm9jPcnPF4C4Rk2JiGnjYzcgidvP9Iz/xOXcg+oxqotj2
MuGaPfvaEigOFrsA2Nn8WV23KV1JBFtGIoB3DHRnSGmTrXHJtnuweWgUmUuc4l0PY187ClO1W35L
D/OdvreO9S1cklR1S5BJ2BG7DX+6mMt5v6zN4EEAKWFCoMuE0ng2NVvX2oWpt3wnYXzQunnQRupx
CH9duZ00P2qWrBJLPvJ6RQvrr/T/DKhiWCVm9+kBL9kmCLlyQx0RxCIVdujlWyz/CsRhwTX1m/uJ
mSCbd1dLt/6R/f0EJcPPyaqWx3mU1RWtpxHpTzPIw6OFzNatpHYSqvtk9n5fKzU17QImgkDJhEhB
EZiZZvySYZjMM+ojPizFmZB7yWMTHPSYRdogC/9hNEiddYBP4RZ0ErYonpm0kWB1V+Tdza+2tjXG
44c1e4ZurX7qWKH6eK/VmV1zvHdFf6Z0GGI1h/j4cNinAUJ6RRlWBy20rXhRXOYzziUcovg5zivS
Fy59qV41iO0RQQVUeYn8pkpG4p7Ftenkl43aJUCvyY0VYq0VtaNnumhCyFvfLcK++7luDaBqanv5
Oq0P54elu3oH0rLFOVDK7iM+WBsu0QgNhUcR1u0mcCz/4YX/J0ba3/WjbeSUzmfAlBBHJnYrn83W
EELyNZBdRCGR8nCOo3vOFxG3djz+bQjQc3WsK9hE5CV+e+EUyZeGzRo8/TC/UXe3tI5q7BRpomv5
896027nZGib5zvYOnXV2DcTbSEOeuhXFD2zqM7AC+HZTp/fMZBJX9pvZ1RNUjcToCU2QC5Jp/Os1
GTy7YFPRh6lvq7cd1aJnFgA6NDAtOIxKLVi/0TFZy7oYvPh+J0HJnLeUElr3rH9wCFDJI/qsiw7K
38r7XwIKz+D6wQPg7SLnE4lz4P3ecgL4FI9Eb7UbJ3hWneXAWBwMQNtMzsHqJv6zAgUQe9zQQgeL
b17xAwNgyGdi7qaGN/5Hx3T8z5Rlm9wW3avFmReXXvtlFjaglQvfCgNnHPRVsjbo2TjFbJIejFCH
9OBqS27GDV9KsGmVO/yEE5A9kkIKX3SkGZ1c8fAgM98o+T/1kT7jl1IgX5JLK4NVyOr8/h4fgAhv
HxkO/TlOR5Gy7GOB2ZcZTWTE9/hzu6ZqQ54B5bk+wqQt5ikOb2ddT2ef7VUfwD2m2KVm74CwlAnS
HfoHXS54b3PSycYNCMz7dT1CXNYvlkAL0zGxzUO6Bu0c1kXvO+Mfrk+5lzL1bAC9sRBYQ6VOvDjj
Su1XFwETNpG8HM5mQxKWggiDg88ltMfAbHTQFxA7+OwyFNGZ2wveeDOWtC2Y3y4SA4FwjR8MgdEN
V5TdGYCTiAuryXIk/PcWcJcXkqRTxv/UIW32/c9w1DcAE967ysgJX90i14VuqGRqiEhXPe3iD5qw
VQmgqdyOGxmkzsRRtasPrCof3qdOSpmqDXmySdnp1MvwRQB+TAtyKA6DfDSlpf+m/oPUg7gLEHx2
5VsKhWCdl5zaS21F3/dUh5ccsvHXjPRVnBtt3pr611RI8+bXxeguhex0s3IAt0wyEUCE7+V4yxm1
2+dTIoYE1oHPakgf6FgwEiDBu5JvwX/jeONpU6ZkB5RikCqogXA8+H6pA3R93JEkW959vpwfAks/
yJxNkE8CwAoG16JBCaRgcod3vitXcqEnlmSQR+S9hSe1AaYoRJ0+cB3BXAjOek98WCHt9Rcs65WC
VPh8yoDc6aB1cmXemiQVu2u2t21jEXurjlk0xkGdgDuXpv4AtfdV5sSy8iJopXmeT++ToOS+ctUW
E0t0ab48Xv6exSWcb2qDA8rtd3VuaLwt4jeQyMgudh6i1V+oqj/69V/Att6I7ayHH7dW0YX8efwv
Gv2PRGKf8tojR2vYSwzx8Rc6pi7TOiJKTKgkl1V7iyTp+Gw7Kp9k2is2J/NKzpaq/kZu6DpUgbzV
WR0s8IZOvsnBmCyOJsF7JRZjwhdMgKBXGskKBlKE+Zfyxp7kwOYLPPGcpg+VdJIB7fyiEdhtXXDU
aF9XDv7AgUG6EoWhmwvanivg9yv9Jbe2mb/J+OjlCpjkYbc2Uy1pXG3R9PEeiX2KaKEuSrpDOSGy
EoceCX+XGYePcknYtxZ28fNSNPZJwH+W4jRBTRG+CanJDdusFUYCJjZMPEKWZMDKrEFk8Q5HQ3iJ
JuxZlRr5UmsXlsRmqxqenIa/D58WekOROSgN9CGSUtfCcWi+ETDVzDQclO/4AUsXFF0jrL2DJ9QS
hsowdgmEo/T3FPIzPeqX5tbe4mWp2u+mD37aslpLor6ZFDgvi/jW+kr4pp7GB7UdoxMGphcA52/G
YsxGvzHwmo+y1SPMuv2BjHgL0FjEfZYbY4SAcLQer2+SRmUNFCJSwIzptZ9IVueF4Qvx5x1OMGMW
u2aI+fmUUWBvWTp2UYLYfY2ijo4x/pdGEOXUB1JYVNuZ0+Hdu6XsTHkIcS00i1VjFkeYrSAhEFtz
StqhQ7Q9jooLcNMYa3iwQc2VZISED4Z0H/01DVKXi5A8Vb8Jd8m8AkbVVEwlJHgSkSjDDb1INm1/
QErEByvPjrjk3bmCCR2+v9EKyBW1RR/XRynqYB2HnEZSznAwZtCfu3HppiaoZxzHjpTNhaVS6sxK
iYFbka7/cJpB+EjdCmvyJpDagpVdppxUNu+mrZUa2XP9NZkDwMeQF+Xy2EiWWYbUmXWSdaryeIv8
QvRPHxcqZdDvut/Yj2ZwqG8KBSP/9KtgBY3O3+7fiX7kBR5Y70nz59YHcXx1GUpuwDwZmnCO3DCJ
boBIy3jJps8szMBCge+IOkBVRtFLUtlkPWqvDNW3ep57VzkqAkMXa3SLR6G0juQqhrasfNkFfi3y
0WRGl55y1VGmOePHQzGmEpvbMZUOTJbElbm91TjCEQJ1FMgfvEzcJ1x4+U5yMM7EvWPOwgulDKro
8cHdR1bOBNwPXqhqHoOdRo+u/kSJiwth54Uf0v0FQN9mfYl3SAGgQeieBs+XKAeAJkm5sAdPWeOi
iCPqfp6eFzCL3PCbJJ8hbK5XxtMQinws1Odeid1eyY+NHYF+KfPFANsyuTG0bl7Pmsw/CO4gDzRP
ZYbytgfVWw2iZnGUAxpIwB4Q2bhIxgk7uw73asQBIKWrXYzysJROJ0E65aJorB4EIY9riaeBSl1m
0+5FgNxki9QTU1Dm19vtALFcsDpNxRoDeOPZQ+9dq5ptrop6pQjj2bav5C7jan3Lv8T/XGNUU/Vz
wTJyfKQSlv4mVrVltpaAZVM2cBeR+1oTRYskKPWUksCjK7mlFnzn9AslKq8d9cQ0Gf1juAFbv1Fl
G4G2PeshjzUlvbPz/ekpCY9f0YRGphhVMSQD1vtPdhg16Q0aReJqGU0EdxkNiy1H7dbT3K2nqV55
CLbQs8u9tUcweYWSdnrHgtGhq1ZocyPyuf/jJ5Uf935GKyyIgp1YbeT4fK0ZsE9m4H70/OObuNZf
I7g7mBCd/yruXbiFdgpLTU9PLGY+4Dk5rodSz2sbs++POKCaOf8xk2Y5YsMYPX275bV0biyHJluJ
1hKL2sW+atHUWC9zmIeGZTZlMqzKJgkZyEPWwtSPNVFYYzd8TUoXUTLD96+XXBw2uaeVPd6PytU6
hpyk7cJcHJF+CWLJVzJka0ZiPR95BJIk2uAfOMRGLkx624v2o56Y9/sydXrCP7f4u3/5+fiOptck
ehfBpYns4UK+Af0NRh/G8gCX53PVs0Lhz/Sp4qoFuxjsqq4d7OS6h4+LH/aVjmB2LxuDP/vmUbiq
Oa5Yy8J0Mv73fFDKAxLKscZYjv7uTOrly2BXHYLA5Q4oMRHC+6Bc83zFT1WzFkHNABQqYd88cCqR
FTVvbxg3fYXERpYqONeF0hillD9jT9R2EIQwiRwCmKMKpBQumfdgxXCmlm8RwSp/J2EZn2lFOga+
7TBVDdWpJa7VbYFGwpbS7XAbz4rnSmQvuak/aAwuug/bkR2xDQsaTz5nL0U/2bWo4h8QkrMm/HqS
wOK7wdvXufoGvfPjiZXUPDB3mRY47VkqOqJQ4hIFSQeRqfFpL6ciL5XTypLoF42bG1FH1zCQvQf0
f8Xne4xzEQoPYvIWGk1v9vJxWAbIoPQP5QUKWogN2kPsCZdzsevZln+RVQaNLsr8c9/Ebuz/Umc6
Yur3ILMrqThPB8UZBat4dpsTLKJVMsqlh1fQoHDprVsO4Z9O6jaGc8Md50sCWE3hdXYtD3GY99sr
9eqtKeewwpx6BubQYTENGhdLuLT+gGJPSvkLn/bJx/YV2Z+o4RI3Ekdl70nXD4qZm6MIXvzkngCc
J6yPpTDD15pw48Xb0453HHRCNPgB5tLyFiqPd7aHgrlgwR3fyM5OfYM3UUOxsI3JDymv4YtxPzyR
WceYhZEzpZ6WvEkqUEPr2B2BcWL59F0pKJ6buMmfZaIV4EOjlVMaG7dTbSYuzxQRn4cjoSou5PL9
zkcLjp2+bYg7rt6uidkZQ5cZyAX7qi2OgEoQdjCAikv6NIT8owaHkR7xcTpK1A7RGl1AseuXwGbc
mm4W5VtF5zGz2TP5NUSmvpWKrM1M4hOw9TKq7Fc3iWPDJjzc6hV2WQZC+5YzznC7Kay2FljR2gu2
4r14PTyHbcmR1/oGyqDaiQOcNLYBEYGiXxAZnTZu8E6kTlgLuQbLjc5fI1D8zpL1w4txQ5xCyL6r
IcFTfENXxWlHgUt/QHJeIn7Xb+AmDbaBnDlMQ0vIKZn58/4CqtSCwot2gT0wDiw4xYOARdYJ+H2r
ZJz6Ak4saGmiWf5kKA9ASEhTK0Yhq6E1peXOXPLZqmzPnAX2QCC0jeQPKOQFJKIPTfPSitBD1ieg
9v1+pemraBAiUkpi8i19EyLlv9vwDgNuFK7RZXpur61ui8JLgpxOZuAh56DSszk91gjy6nkQv4uh
WNLTUqrkTxC3LJDzlTPdjIUNkDiWsArxYUlC0+hjTm7Wvbt1NoSKdk5/kIgWXyRnQtKQMBFmmctT
en3gJvKKw+dqcsZCTXyG3bKZ2X3vtWnr8odlidMaeAotzxCHgQ78Cf3QHP/Ttfw9NX39qfF1XnMP
Eu8m4SljOd4yciDcymY8Wv6FNczf7zCHL/m5S90Hu0AfVbRpL8nCRxty2NpwrjfFjUucNKFooV1W
aWbEGsBeYyS5USFFJhOTh6C/xRA5k73Dvrl7JFr2dAb/1Z8/DoBaAHD5GWK8R75EBtN9HwRLt2Zj
iIMypz4YICFc1HkYuhgVqCoRbpggJ496YdSyHG4ik0i/qO5OWQwTU1Jzp5c4W+983YKOQKONB0Yo
J3Hi5xyLJlU+8am12rL0Eca16rYph3KxFFGx5/ftkNBKIyhHH782G2/gu9Ksb13PpCtGNvzAA4qE
Sz6tf4dxSJDVt3c2c5uDaE0LCZd/2FeKcT8Z5sWZzY9Tx4PtXCloSCoShGDro2jZLW0WcZHQ9xz1
KuoDPqAOygbV7N5Y1SZ8DyoAJJh65hndhv+4ZuJURRi3kJK+qIb090ReMXtIcY5fmZ08zayW93e/
WUlNHRfv+YDf14I1BT3wD6K+BpkptoRT9GD+jkm97k0AZa1/oLroodL5CjmCNl0IDUwxSmb4f90h
I+sVN0+APHaD4QDfh2zYkopsm0rtYrfKxx22zDcHwfxBs0b01IgL9PtInEIa7dpFPnyug35hg01X
QhHFWXzIXdSDQqwQBuTq4zM1xUVZJY7al/ZF0PFzyIV8S6V0jFbuwlrCyvfFvmaPv2gO3XUtaLvw
gXjHAYBGunerg8QRblpCs7lhalDKwOEYEJk5YcfNEJOLeeZvTOsc+GdMpYaydlv1vvYnQ+ky1cFe
mI1apQ4GIu8cXMK+V+DDWSQpm1DQGcAS9l8Sdv+APtQtFFzU/WlhH7xFN0e5aNIk5AlYCLbfmzii
+kHKw8nUX6pZYqNlgaDK81rNSZsKe31+SOKO8rjVn25uwtuhHZoCAT3M//yyIFZIZd0iFa8lWJhY
J8WW2/wLxSy/ze9QIvB/BOyXM/w976Ep1s4TL6tKK5vdTc/hzJez/5nw0KiGK8AEqrFqu9aFb7ZT
GgcMh4UkVYhJcox3U9jy5F3AgyzyHQ1seXjx2x15qRMwW464zCKc0ieXgb/QoBdS+ySDHVk+rGo1
WV47pHV1/ie9auQV7bTiz1TeTgsshI7x0hXKZAQBwnFYLc6n4gXKYLiRIijtgpHX65SWgJFghRIV
XothvaEwDLDrNTliOYLxqZr0Ki3lJrYtIROkIEngsuhDL0730/GDILcvlsVwVBu2xqmdnhYTFc0w
8gjb+7KLTzPfREIJwAwd5ZonPpbHU3b6MbJN+IN5prEwoS8mIcmvgBJY6AglVXe0/JdZhuzzmzbc
AByAEhROe6noeGDT+0wXfgqMQCHfravkg1HXkLbog+RTUnAOOo7scSWEbAKI70EUkU/f34yMhwor
yzM+zVYmdpfYMsS9c/rz/Hzvn4owh+GGz12cnCosHk3fkDCQ4whkpkQ1rJdWsHPvmkVYU/aXsJd0
YoVk4cX0oPdLK6d0UD+gcDlnq+TUuspQ/d6j2MKybD1gk4VWAY3AR8/Uc4AUlnt2ejqnZ5LLNRiC
+cVWnO5fCBuu/kcEpq1hUme7bYL6FcHZ5FECbDYTVlpvZHUlErvMaelj+gD5RxNMs4djtBSLTnfn
yHuKJS92E71s0NacRcMk87fb283pUWA7IEQSoMbgdZ4rzXfbRw3kzdLpLyA0GxZQWsxEuNB8D8lk
lcv/S5FW2xKjZ16RnW1qQR0JvCWBawSk3BUHVJDEENoqLWEbdf141O8Yg5xH9bOu/4fh/zQy2gm8
ew10ALghu/lfaI69snCl40AfusHzR9WTF25VTOO7B6wDpcqIGiOhuOQ2rr50jrZFkEh+DCOiGUgf
XhIYNSyoUfFcTn+CF3ZrPqXSbd5BJ4GypM+TEFH8djBnaOmWZXKeaXiBZjXckpR3F5iH8vjNyfWs
TceHe5c8IReRS16sWJFePRx3xvkLR5/14EPLyacwoYRBk7uvSDKDpWgnKauLm1r3rYf9J7vVLc+U
pipsJwvzleubGfcrSw+BokvALLgtEu2gr/nvWfvCNxh/BlKcFvGcqLUchBYJydgNpkallceAkcc/
WWNucXKFmkZMLGDzoRFjQVQItMQM1cHqo/CIYw7C5VrwqQF9JXHPsP2xBRtUC9SaUzxKKBIdRmoP
XFDollOtg+61cIWhTpQmIxYr6KkrShEva9U07gQd/GS3EuaLbhmwIceLPsXzdZ1LDXLcRC8BbAlS
rML2ACPV+jOJbbLX3BGQFxHAJhRoMK3ZSuzAiQJj5BOv7O9WvVQk0P31o36rrjCWEFdzjASo0ep6
Y4cFT/JpPex7VSP8SqbjZkuau+xpJlLmFp5XTHzWWyYnzL4SEjvlmuauuo8uyFmDjxs11AskhQRX
HJD65cO1sneV0wyV/oD8lAHi1Itm3P8jwxmZpKuMV2jjRVUcPhZ20kvyaxlxKDOPWAiT4PJvdpk2
+Cf64b+ymBdNPAtEQAIcgOnIwJaSRe2KveX1FlhGybsepzA13uYrr/g8Y5xjK4mS7F4SEcgOPqCY
EaA6G2dqkLeufOqxHrSHZh54d7fjUj9izSqYlmBa9QDJiCK/QTNYkzKpEN2hXF5NMfMpD36QNf3e
jgouJe2WL4rlvXbYvpgijl4OcMNMg9HLBroCgAMuNJhkj/0GNf4VK4a6j+cx1BTKADSscXqf7rQq
anURHjFbaLWS0guzpwSvKtZkbmZBD5yIgagedoqLC55EVFpnwc2jE2e3sKYt7IQNujI+ZjghNL2L
A1Tpi51nCa5SzyMNjGMJ02sKaZmp0oweXb+vIQaYJrnm/hTNKXyY+WHeabF5y6BNuFIo+tMr3CYF
ODgUgnmtyTyX4rT8JuPg9eCmTA4yrgFnqlrH4bOugYqrYciU+K22eew9Gv+yli8yXdadEFOLR60H
sbnTrDjXVMdKC5hBw20NuEomJzpmoWgaJ+C0bj5GLethpS9miBrEF6okaGbL4t2qT9zkYMAstcy1
ZPzCsFVCcfv6k/JzQEsEmP8hjDUJjppJqenysJI/ZXukyODAnllrYmjE/FG/YXJDIeAwO8fpF150
Zk5JFTRe7ivevn994bPsztFghbuLJ6JfRkSeGtL5uKkQ2zxL/3BQOrStWKV7ZfpZ480DNGGfIouA
mmieey+Y52A9oCE6uLZUBh+6eWsdfs86PWjEARJSHr2Q1Y2Szbed7AXGg1Hr1vc5vJ7PuEFNK1cq
B2gXAg5IqRibZ8REv9joge0dz4gco5/Z4TWVr0kSNvrV2y1qsR2xMLcbd6UdVTFdTYVkjQpILa2v
3qviC2dBDWjfLCSkcDYkcAgzB+YG8ngPZ/aHlqTVjYeuS4ZFqkeo1obqrOtt2+K5zH2BKKRFcV3p
WtTuJnr8Tai38nrVpxRnjv0YFxmZ3m899rf8LYxzkzK5nvcihPdSXPkuioKWJ05jsi73nuupJw7H
SjHqMY18IQ+AoWXPdyQHW5QcLiirLfcjNkbkfGlMB5gGYpfHoHFxF1Rk1KsAPNvBIyBtYOsXaMxa
YyxSxn7zYjrT+b7AyVKMNd1W7ij+aCrazZ8XxG0HBZ8rAgiJ4u5L3e16p1HE4JMYi8t4A0/hRLqU
1L6pRicpVsDdSRI/GT9R+KEVQYkiV5ss9vX9fLj3ZCr5N379KaCnvSveEo1WcMghj8rxYPgEQwUq
MW/RzTMqJDOSJIG/7hUNKWt4kYx2ffrhhh6JCHoFxU5SuZrbIw1b8NWqhUbCM0XNeGPv1qUDVD+Q
5hzhKLFEV695R5gmiU6epOugYw6N0vbvCiE1lat1vNtWJgJwcuLywswvbQd+OsoPfinlbcMIC3eG
VZSG9jC+MTvqrEoSoeXzVAbpw7QGAh6+citJyQMxBmHdajVbfG+vBBtKGmC55iTcud9VLW0wHA/r
rk+IptEwDdjWLUEBUGcgK1TRtufzKe5HxEJrt1L0xZpbgXWQcgzXWPLO+E8vAkwQaXzlqJ2VcbFH
HHOSNHyIcC3zKo5de7QDnrIq0wzg9aOd+Xeuj5ldHbfPH1F/9PEgx1ElmDsIMsfJreIwdY3V4bBW
1AKCqAMlSMPVZhDOXDiO1lqoDwD1oaQC2571/PUuX5vfFvCE8whorwqwjG8uX9rMSyz9VQVKXsa6
jn+qqAxn4dKImEmLYcnNrn5pC7SKxJ+sStSexmVnJKVbeKHn6+Q7kDi40PU8ghaR5p6Z7JEMPTiQ
YPu4jwbjaRCqc/26uT368c54QHpiechEvYCCicXzn5oVU/6RtkfUy2izMDbMSGYBvHf0rsBk0j5M
AyJ8G/M7QJsaJRyVgjM0zEwTljK0pOaLfYMDl3V18t5ZdiVoYHRydO7a++qUQ0sTKL9K94VHapd9
23f3Rg7DHVo5qYy7E3gF4muw8g2dqEkoLAFUolKhITD+E5R1kalLXbc9TJ4XuUahWu3s22CuE9NT
SOnuHvoCjuXVxtWiedcUbSArPhehnEVbdDjz+gkkrJrSHulpY+goi25wN0wfVK6s/fG9yD5Zuirn
fcIA5iJUeUwcWnZBIASpbtzJN5sNiORzHygo20OqJPrA/cqXqI+iKCi1Xy3SBi7/0isYQ+oZrXhU
BtwADLX6iCjWjv5S0SR2Z/afsrEo7PvHeXdvLKZR+oeupVnWpWCE8+lCgZhzUd73CrVUZBIzMi35
Q3yiG0b15+fN81u1CNjoeIZFXat+3nuUh89RJqCqwutZoWU2zykaq3vnBlnUBechVGD1F5VGs8+8
MQRnEJgi9umX1ERSbartO0vO6kQE5q5AAVC01vmr5gA6nvCvegUDeVsCn2Ql7nDnXj3bFE7oXxgZ
Pb7wpAsibZhLk3X63XbsZ1+jJmXj4VpE7LzLx2ArmpR3YuTmIZezlT830cJzioidrjNjm+BMR+1E
GBkJ65bgfOw4sjHEI9ELmkmKJV6YXIy+EsARPq9JofIsM+J4bqVAdAEwAVQa6BHsD58ljh6qnCYG
2lbFmFD2bmNEjeUJ6KVw1V+qAUeumMS3HI2VbI0rdscdQD2BVY6jodfd6LADOJbAEDsnhK0BNEO5
rXTOCb1x/xUVDnmSxQg8a/njh9zWHwdb3NH145Azxjdy0VyiT8/Xi0ZVT4xIDT9/bft9UWpFiyvG
WI49IWhaIN/xz9Hbc5FHPy8Kd8XmUQvXCmt9uW8XByanHYabPgC+x9MUBJu/pkXnhhnbpX8TDWCw
6dj1vBhSxv0rG8Kb33b/9l7j+soOhMimFH7B4b8wDrbW2RWfY77Hd6X9oJIf8hR/r1KW9GITbWiH
dctxr0JBlnar5cE3yOSiB8npAypVybyELUCAdMwj0hT2h+yMiHrvAriXK4UpFOcQP2g51mknQQTx
oU0QYWzeMPz+2qhvdgUerkOq/Z8wFEnZJvCsrFtIa2pAW6PfLAuIUN5TdVq8cXdb5o8BCmvkP+ey
Pryjp3DZHFg5jpK1QeVDRVHt/QAR5Ul0c0Fc8RwOOP2GCHo0iEm48cvvNqbOVLV57Xp0wuiYBafL
GQA3d7T3/pK7E0S4BVKX+3sp6IcBouNfebC/es20BYmDhY3l/zG2iOLXGi9EHJtavyqA3kXnS0Mw
awJ/nkUyxnv7pXk1S2jqiPCYhpQJ2mZNirQdR8wGdFAkUcufAVwNh31I/nvQuGpFnyJTVK7tHN6e
PtUCejfUqnXUEL9n2op8BgZXCIdFoGkq0V+53ZQNxhoaV+qaqBozQUmtBKsLVn3DVw1QylvuGTwb
vYUWBY4Ccd6IpSLa835suEh26HEN9jEulWlqrs0Pl3rJF4N+xA21uTGNzDifOkzLB5ICITaRPTh5
qrD/22jU64fQXy2/vXdcijcJj/mIDmgtRYybDrrVzUiBYF1UqOq//Q6hX+CBsrWndkBpfmDJw38T
6sUcSEE3jHGX2QqpMMzejafpBZtP6kLw10Zn2KQ2Jx3Q+bwMp0NYrryNwcAdLfls10P/9TD+awLf
k2t3Mc7DAaFj1PuoPR/sRCgfeSMqqq/tIFk/RTK1UTx0URFAerh8GNfht0vRMO2UtQO7tN6w2cf7
szls+Z9BobrLlejcZVg9IwKKZkPkG5Q+7Ve1BMs4dJZ2q0LZDFdctuHyia8pAZpH1EM7U+Rmz54J
0gItd+EkZe0C00AW9iCh7t/Lrje9Bx+M2NKkizOedNtnLDAd3bWjTwr8Qhy7Nqf7GktA1q39DD8B
SSdTimJJFqN6mB9nlhx/hxm6WtMRrrlpZkFVrIR7wQNYyzpjnRUE4954SOC6IG25DXwFB/5Vg0ot
oQ7hz2DuGKAHSkUK0lSvvR6hIE2uzPV1kme9SljXJQq4zBWCp8KHFzHaDMJL2Ehfv+LG3ELI5goj
ugI5sqHmqFxbrYDJne1SxoQrjg3LYM2pnrT6efcy6244A8OmmvmeCotA1wqRoDi4Xx2MkYV6twtL
dc1gQFf3VnTUkFiaG9EQLp5WvEf80y7yiu66o/MkpOxKBykrUEO2pXhRiroXgzT8isfMitlYibtU
q0TY+BG0sG6BN+vMRMcE/JEEXXdy/e1i2CreJAdPWE5u1pKwJUcHuOj6VBZ1FnEeb5hVTKhDufnw
RKWlQOxHc//NoSJ3KJmz5248+oNmSYRE8hkSxdZw+p0fEea54OPqyJ6jGnRme845rpDCli3soMn8
cwbiSzrtCsszOrxR0M7KxCsejxygUlLGE2M04wmB0lq2QWsYsGA5TV/BdMR9y/+HGuk84oUkNHpT
r1mupTZM2Rn/CrkqQKC6TDS4TEiXFcA9n9wUJ7ZuaE7Zix/HO29CPra2fB6VhMouRGOdYAQFYhUC
OQ8ePMZd6aKyUOngUOOJPCBMlRdlmJhWE8nBcOTVziC7L8Ouwfz2lu8EDTskVCvbunsvU50fCJTw
3AXIeJfEiO8vyl/3k35iEzJ2KPYCDL8Eo/rVxcS9LR7sTRfYE8wMJqu2DnxfP6Asf0SnqdisdrxT
ZW8KERMJw+O3AHfZVDjlQpns1fMLi1r4yHjupX8npefJXt1OSBQAzQjIIbewCbzBBsfBCNKQvkfC
4zF6bDSzv7CMA90Tdu3sqfh5YomKzxTAvsRPw+hbQaCmbYIVTQlX/qVDOqDL8m+jWnH/TZRyEMJA
mqOlsdVA3SJnuthmmMSoMOkEqtm2Mj0XGqZnHFOO534AxbN+JBU4dxWTvkQzEgfjfZFaM134omvH
7f0pklmnq9SXOOOhfkoogH2bhKaBWjL1q4Yqapoc52CQtKV73cqPVslvg7S3+XXxsyVqyDK1/wMv
TsSOpMxLkkT5XEZfkBwmuI+r5E1vl8B9mMFlyx74Po5nKROUxR25nhZ7mn6fA9AgAxQFvuv3aLnL
P0M4Q8r10ed1yAM/qp8rNrhMVDBtUs7ALXTD9WxLgJlbLyAEjQrZw0Ry/v9LP9l+rcBJMknw0RJq
tf04e7u4em0X3Sb1cN6AzsyS/IB8nirVyFnDQ1y0HPbnIxRdkkquNgrSXeYZTZ7TzotdmifJK5dy
RWW7LeZbyB34jZ2QcLgnKxSPpf1gDbBwMeBLy0YrbxgozLGN4S3+5p1Z2KjfyyPb07Uub0lipQP3
CyT3chsaSGN6tvu7V3ZrKMbr4MjxNvsXRsPLzesb47LSDeDthr1VkPMe615UN6o8IMw6MYklX0l6
b5U3dGmSWIofxxB+lQouoByq/8p3xq/2JJxnDgxh+TNLeegPDouPGMV1g4xr3+tN3RdqglssmcaI
hTW8Ef1jZwhN4TMv3xdNS3Q8AiriYe8l8WcMZ8mi3S6ocXuxJiSzIhdCAFwC0JoVSmGrkOcVQsha
mGGXBkj7tP5EzjmElv3kiQXRPAdgWRAtzRrzJetdRHjCR/O50747wQRN8+JgpyWzl8MC/UuNRo3M
F+bB5eEKscrDnR3/J5J10mCmBKvQ3Qb4F56NLCZH1QAvdEZkvGDFkifcdxLRlL+bGdl05+W0d61c
z1A3+rLpGXMjym4rKEoikZ/MyXJ8vpjMLF/BRz6etnK2RJOfh/7AutEPgxRP2O1ppgOqP2R2+weT
r0IE7uAy20kf5LPv7CcpJbHntgcMocoqsgnrhll7PlzHkZziEXPOCCZBkBQNLd8xzmaqOWgM1Qc8
FGFdNA4+XIHB37XuUYFk5raErS0xoUmp+BZ8TvAT81CRJz5EaNE6llPtPX05GmTBBo4OjB52+FJ+
5i0MghNdpImJg+BMROI06ZXRQGqNoiMnR4IKdlnrHReCngdYuoN8XN+1M2h5r1/4Yz+k1K795U64
1xCwUJKEa2pTPZjKAAg+XNenKd8vERS7VRqQEDRITJ/QGpJzXWTKAB5dZxKoyWjFmm5LONoNcQ7R
Vxzlv9V6TQQE+Xky5lw5MFgaFVY60PZKa8GZNfnU5lJ6Le7Ra3ulRnsm2rA9McyG4uvVICaGRTAh
rUnNGCQMxN7IySDS8/7NAyyzd9d3kniYa+LvFCg14dpEPQ2KrGXsEXby/nlOnfjRgX5gx5M/JFf0
+vwgH+gBMVpiKYurLL+B9FK2jOuaQhX1aU/zUmR1kdF8RI1qDzlSFG9z475T8PJYgNiMMvqfR0lN
ihd0AoiIwnrejs7v3B83AlhOUe2GWSR+z61GxSH1fCOmU82TDOZMi4idxmM1tazlgeRCoNOVPM6B
14MTrVUA/DkUSw+LgG9QRojjr1RgsFtHueHt4U8UtRuK7qNzWEjLGwQ6hGY2xv44HE4an5Z0w1mp
FvsicEhtP0KM3pGBfLNl9AXiVav6gMhltFZZktrFu0/D8dk2sJgOvwVITuJ/onf8R2rqGCbfPHLE
gcXmZ9jdJaLqCpqXDFSmkb45jQ0N7v4SLMPERJBHOjPXEORPMaisImtESgsAFLwnoerfYtE8nJW0
4Nj7K+kBdMC7C1Vb2aSl5+j2V7VQELLxwMPV22LA+8QT3lbjIoeTA3Rr0rvgHm5oxr9x+X0iJupV
fSbDziGSxiY4s4fvWwDbgnXqMR7qB2IgBTdwLc6feHf9HcqgbnZiV/xGg8a2tcQHQ/jRfzcfNry3
bcK3COUAK575CVkaGo++J/nlaJgM7ea6M8V1drzP+TNp769BHM9hLbDuXN6BwD8KisivSJ9fb3M3
nZ/lJ4dYWcHgSLfL0zcRby4+3L7mdr4nxpsNOzst5VoaYig3b/UmD3lJXs9BQlM9v0fXHLEqF5UN
R1YMfRrEz6w/awbQizf9+E9DPBq7t1gWms0WHZZnOiIfssPBnaJPwDc67Qu07HagVtkJseNBSePS
mPPhwx0cxpCawv3vHuFcMj1L9TPPFj9uJKJDYkc8g0UDzKODDbUS2X1NbtxE76fhretx7HhUnv2z
K9EEe3pfKZ4+cDMrkkV0SxJccOWYrhUXuV9lY/fFxBcfcmdJEzfNkUb9D7nJ7T68SAPIgSKIBwfx
3rB2nA+i5jhls+EV8/0y2T35/cmYvKl21/YP1sqKaNtSZxCxMrNitm2WpgoZoLXiXDP5cWdFRBrK
+drqirnHyUYij/lBxZnnXk+6m3VGu2rrXUqKEMaPmI3GeKlacseh+dgCJrLPKxTK1XN9hSUrfz0k
ZJK0GLMqsdXbxOia40DPZX3dl27EfaWcA60N5IxeCsRl2kYuNX18+p80KHV0P6JtFK2F7uKdMr2F
cljH3ciwscPWLhGY+uG8MoS7DA1IyCN7YduXXguKZisIJYtMLUpGxd3Sbv6E/kxKZZSkVs/zKWB1
swWVbCbXsxJtoOCxVc+R5+pdw0KyqBaK3N/DJv8q1d9Dyk4kJf+VJVChn9EY6KPZQQ0AIcMT75Xn
2ACZeN6e3lz7jL5Pyf9xo5ov6sWkGeEFiuXCOv8XZey9soWlcdQzeF/VUMANVY0Len4sFlOuv7R7
SxAbpm526mV0d/6vW4XCygoeLP0HjFWWuBD56Rhmp8yoQj3BHL71/sn7PzEcPaEhqtOyljaaZaP0
IkG4D5T72QFPw3l8AbtVQpSEWqjiBEtbsh1Gw2X3rduAYjQFwwlqlkxcrggz6+dE5PdxjwddnaZr
cRbsPOfEBb1OJK0svt6wg5TK1pbMHgOl+y+m8D+8dBzg5Tv+tbAvqaXCF5cOb2+7xMzXOymv+yJl
l3zxmOO0OQmooXooIi7NmBOLRGI7MZ85FLSBudm9+/guzJMkrT/8N0MhlfccGehNpt7h3epwoS33
QpnSIOSo3JikB66qDOOMe9NK+Wuy8a2zhMOFHYH+0F/slfpr0LwkHOeJ4JucrJ09zLCUPPSmzOi4
kfNvBGl4tsv/JxZkK/Kio72vehbEZRCt2rrjgfyveQGkIoY097hQe6TK0Mqbm44rY7uE6UXtQOVU
XusdrCyfoyc2UmEg+thshWbMkEIAYYdjZvtTgkahbZB0xm9upEsQ0GPTg2GJI14c5AetyezuIsZ7
30eDj9Xn5DDYRFxTyBpK/jXCzcSXQVSqTne34IzdCQzJ/ORiSt4v81irkVSq5PX5u5g6SmQSYVKS
UUzpPJH6vrBBu7gyov3rd6eQu0pGoQPNVfxGeeGHIAHz7GzfE2f/2DquTh1oHT1TmWQv3bCVlAlQ
WTySYZNVUWBvUoo+r7JwsdjxzPYjwA6VMZNiHpvjCCkMV+cirix1V8tNNXE1Kj/JtiY2LSSAnJJu
iRvds6ETPCm+QaJSZrzdDWRSqY9l/zjwUV8lw6FGBUe1yLDhdW/HWjoesaMcGgCwcxrkQHvKGChU
v3646vPKFTkvQwAVbvUoHRytIokqmHFQpSzSElHSw81KPDI3FChiVjYYUqLsfPUESc+onD2KcSHR
mZrpW9JpWuu3OcRNXiAm3+KzAUdHjVKU6sdyVVZkbb03UuTjAa7N5h3CGo/ZqRw+0wQpb9aXe97M
csZuAiYroE7VqdDxPvBVT7heDwymQlq+xewXQStdNsG42OvS9l9CZuiR4cLsBC8IpS9O8gVmzt1B
hHUoC/tYv3TPtgfcmQO+2fAlcLEhkIhP7NIh3jTUBi6hkSSRZd+Aa2A67B07enm3FVuXISNUzl56
0AziO9HqBTHQUQTrmwM9oWZX/47kJaRVrNkrFPG7HEjLAf9wg/xMD9nDNWtQSwwTnbvyOw87F64R
DaUINYKNfKL1y/bKxS8lThepxYPpv1iMIqd8J09ekdKJyNF8wQopUU/BmQIKVIsFMy/5d0TL4HnN
SSfqClK9M/GagZ7uFxspGAqE5zMYc3D8L4GEJeEN+iZymiZi6JD+LhTP/vQDXWygMDl87iodplYb
F47MHTgq7ot+K9PzuWgP/0itr7uO57WBQlND5trNmbYwrocM3IZ+mjrpVL7Ch6q5rE4pekaEWSWT
fX4NDw3NKmM3r/xQeaA28kDi15VQednYN7BSBFvAylaFCM/nCo31epJyr6vSeI2R+MJavLmnWvp+
OQYM8seDyuIiAxOgrnqbHCphwlm+po4vpfrLoS/9Uml9+7T8M+yf3cEh8GALQ/voSLHVyCD45GKF
fCu/HqNtDFFyZm567F7KdUqI3fhpgMBJ8JXpNH6YMg6blMZxT/7fTlTHQujP3tiDIpqku79ewpPa
nyo9bKK3MO8NooRdekN8QtEgPQFDnvWgdl2u3n2h/1SS+At4Z1JS1iQm6zXBoWlo0O1aV5v1ICF9
KgtMsqLODus9L9eel+riZYZohoR04E/z9ciTyw/r1dCzM/XS/GL2ql8M5nG+csLMqEhZZu+hPp7s
s6KmLAgwPyBe7yH2/JADe06SetL7JIK6abH5xBCff61207o73ZqQIp8J1X8+NitqPZoQlQoQB/Gd
L6RIKnZGdOPSGgWN9J0zFpf+OH0xE/hFfGsYE6DZP1kjlgnd9Ol22wWKASs93nlogJlTaXZ+dwoU
v4Gi6cssrmT+sm05X5wKRQF4eBEHl/9CMyYFan3GzpuNDHLOHZY8bTC+S+sMjSK/lisLBVMYOyoR
i/nKOflEjX4kx+K6L4HrXNIkmA9qaC3xsUfUBAzOjQwD+o7AfWwxcboGjjpFtElQzzUTYHJ+OPQd
3nbqnJNfI6trX3k+TIKr+oGUK8ELwiIumZ9T2DiW252NILH2I2hgnl9YCXf/mOSMDRLNdDVa9B3u
AnEswOFamqL49fQiz3P1iplczlL4z9hbjLGgHa8cjupD+jZHq9UyI/dIyNaPAe1Y/K8N/MwmsB5Y
4akrnP2tO/eDOc8HpOB1peWqMrBq+yZ8BUxLWy8KvYC2sPthx2dTq/iXhUNtzfDOf/1CB0MsRJe8
6At+FAefiBfphYoLZSxB3vWNfbEJhk4b3yGRUsr+KvBPQG6mVGHi0K6xre1EWX6rF2E+Uauu21tx
hRbw2cKgVt6yUNcw1DiKVec/Y2VR8MXebQ90VY51uakyiYJ5F2JASw3TvBe857XumJQ1yXAHFHtf
bnSY1J+w6ZoELa3Ooeqof4b+tpn6EZCnMac+6q4D6ZTPN/BCFONacc4RIHK8hB/jdMNmV8FVxxqW
0cEbbuXLo/3Viv9BdPzWkxoAXaiuPvECBKLfnd+aA5Vp8Coi67ErEyUXVc4vvBCDrQOsTbYOBIed
Cgi18DkrPpUXq2UNaHg7k6zoHuOOhQucSV3eLP3CM5Jlv297mgooqJIbuh5IBTNK2sfLRHBGq1Qq
1fn/oNRmpz748rv8EZmhSBm4PKn9JOARDOKNRFhFSVbdPeQ8XxxH2HdqPcKAKAcATxlNjlfpu3qp
rSiY37UynxJH+S63YXy4FczmedJ9hFtQ8Sr2wEXKSzA6EHfOv65hYg/Qe3RsVkFHuFtcjZ2dS/SW
14RuqbRuGG5ZSB/EPhhmyHVaYZLa19QeCg7p56qSCvgCGkGWhXAnLF+gsFUSNe33vEVMu15KKyn3
Uf/+FUqODw81nPmywiwzb1Emxj0mp+iqJWVWYBIT0ZKp0HvDM6IPN23DRGVmoue3eK/G2xswYk4s
v6A4G1RXxyzcDEi6kVQ5yrZ8rPjGmatS+gH//4AmCXzzxBQti3DugQFjX1nfZtwNPAC3UUeCiI1B
QKybaPcUZ7CAZw97jo2S1/nUKR50FcYOEC/pXxKGTW9XEV3a6NJCJO/PtADDXf8xLjRcUmEITMGP
tgYfyucI89PYQc145u5PjsNnGsoOEiawCa6MXL6eB6q14MoRQkrvXftlkWkzihlD+lfwvsWda9Xa
9kXhSVxgm49+9rqs1SCe41GaJ8wTY673fSqmRgo6qzFi3GL4aQ5WjBnvz8RKWZTR1+m+7945r2lg
lR2maaHnlkVclmsyDGAr0lcJQvjs/Aw5eH8/aQSGVMJHo++au6m01PfzBdHkKTRulmh5ZdqlvHG5
oc6lOr95NW02Xp2GniFaWVMspGhkitiZBnXBL5JNgICoTOup3bF4P8ZrmXYIViP/Z5vpVetFYaDT
0KoHim6uv3B8y1cTrgffcWUlwgBqknx+pZGqA2w/GtrMsi0NPCIQ5/lHq+sr/ORKg1BUtfEmmuZ5
lajTdOpRTAuA4S+bK+1XH6UnZ4nen8h2tBsROe+7iQHELogamAbL4xsOCXtqIBUDCFE2QcVhJON+
vmJDmgQ7F8uzBOZQZl4uxv2f0ef2S4fnu9P9hzKSA5j+t6XkgPO2XXsVNjahOkTqubojVpd+P56P
G3IQ7LkpqK1XRlfM1IeQjEvfuxdoVSW2pK0wTGPWhGA3RZLrBz+QbSIQTqGgepltJQC7jiPQpyJ3
bnsjTBaOsOpdcucOYyo4dLwUJEdprQhRLDwGoLkKMphe9g31GImKDl2gMOJBLIl61qm6f8fmN834
KbilZ3pIQqK2SuLWD/BclWixPCf1fuUAGTr00oWYv/jdCBZw06hDhRpN3aYWK0lD+n9o7Be9SZ/y
Pu/gfG/oj14WYgui8kgJSrgjYwrpu8wfcRMZmQdQpe+FcnIZgtC7G40EDvGVx4cchx9SmnyE7SZM
4Ok57bn/aS37dQ5X3tOTFu4rm7tQlJyu0Eaqc3tP/gx21UBpfc+xwWlPj5nU60tw4xgvUuBDVUVX
QTffu2jKovruAjls8BfWi1of3YN+08rFcyqJxErpwPuNyTnX7LLyFBoe6+We7Kz+EToTfr6U1Am3
CKEDUF05GF4EnKCwOh0JQ2doP3GU52Uv+S64RuqzRJ8oQ002qGRcQbhFZNdsj/kB0qT3YEQp1hEk
nHCowQNNBisuk9PrFWe6aLcwUo/wUmRCDHhTddmg5Dls+Mcxb5ILyIsmP75lz3zdcI8fxzJcIN7/
XsKcF2A02nK9il9DGPTDzInR/Xd4v/FN4P9QtxoPfNdBkBmWR5IfrEwxehywcGFZLOb0YbUrhwzt
I8dU4Kcz25Adp7YcxXZy80oOgWCp3NKzsmYDhfIxwgQsXMINOvMWqM4bixdbYQYaPJDozLRwWoGc
2Xyd90cuXi8P0h1/Irb641MH3Ms6LBv4P+7Ejwgf0ozXnBCEy0DlOLoYCVGfp6F3306IRuCGIj58
ZCItIJChgrm9QZQy6IwTCBaKQCGe6ka+qJRzUnYpTS1Pe4HbwDzEnf+AGECpKg/OikwM1eNjbr5x
hmvbeMWrctBHtgBxlTlfgxZpT7bS5vA6C6Pk8Gs/DVAZ3by9wegki2ztAzLsHWfXJkGBMLlGXC8d
Io8raCiZU70vLPF2/7jwC95oLEECNlXfybhblWEBXMG2maJo+urteZ7ZaN4bQ0RJtob8jjVOwert
SBsqVyGGNVBZ2KYVlM/CZpu5pM4R5fJm7Zb4Ha7GE/pUf1ZkigSM08DFKCU0MpqjG7hbOZAEVtxK
uKesaSwU15hoLXcnGFlffWGOqsbBrjTdWWE/9StdiAfxNtDxpeIosjiIsMFxcD6M1MknEhlBtJxF
Hub/HkZZo/zR2FrilvuCHHQj0DU82zDJYSZNEXpPiQVrGnn/9K3AEQZv1rRUwMq5SGjwWnujd2ET
0PLVgqwHwr7LAuTaQTKfk6IF7gRcQKjx/D7WssyGrMWLRnPEaixeIW3auGFKXKeaWRRrgAhBh9oR
QW5Xq8vJUsISY+ErFKQRE/xx47k5dkFVztbnNKRmOYZv27hew4OW9EFEpf4vIMQ2vtntyfR/fgrn
CT4RlOXjI5jrrZhahBDwP9VPMNpYVMaTUBTGEFWFOz/ADGPJZNlNpLqWy1T7zb1TZp2OBM3rSzet
RtHnvpKZZFrgWeGoPVtqGB3MbRdhAU/FJOV3QYzGXyfWCQcv9kONZBNgpbh2oJOBuMuQXRCMA72w
Xp5xDbhgbEW5M4G2pZvmFHNwBbe/ZRAstKOdaOio1Sh91uYWfzvZ0tbM0O5IYaORiUuxHIOQhlxB
v936ZuU37rjE5Rxq3M9/dBT9IODfHs3V2v++CHy0xy2GHL/8reHaICq1UZZKyD9EiLxTs7kY2+Vs
l/Oe/jQM7oTWIHz5PaBUkldjnjHlVX2ErpOMXoxVw/52unoigu7dBLhS7hhuxI4zfChWpf5XPQzr
27b6LoRa/Q2nwsVxA3h1DjKb7J6ZuSOW7PFEE9G5YK/Msmn6N8XEXHJ0AQVTJqHghwg55dy5y2vI
0DcecKRLZFO7Wozg+1+MOU0Eh/WqthhAgyCfOZyfXAaWBriqQk0q9dr9mD1fwWDrNazoG2WBPZMU
zY+q/GgYSDDbCWX/EtXvb6ssgM0i6OjiHsx8rK5y7MpCKWosna2WtrwR76DuS79CSYNJaOBpPmOb
5ynwil9NBr0V9Lp7x1rWzxCIAY3ZVpfuMhC5n9rKqwseJv5Q3Gr3ddQVyuqyachl3IdI85LGL8+M
DHBYWw9HdPxVxiCcWsc3gjjybmxX4nqZRV8KVmXplTZvxg0e6qhhliBcjceZQjMJ401sV/9ZCllt
iDp3eTeAREM9ILTpvoJzUbrOrIY3t6hqdOqzpgFeRYdan9HdZ58tY2i9PdNqWDIo6C48HWRDJFhy
bJ3pSP1ykwjdLjU7CtqVrZnaX6j7+cKekAzVoLOcJmxS7dwOY5X7AdgQZWk7BNy4uC9kxjXzraWI
LlPTfYgJZq+HIHaTCJLKZW7+hKDAE4J6icCKSqoOXeeBcnoR1rnWJfa+Z1tDsmmlih4ye9RbaUMG
rgoBqwHVUJSl9NWnhdtKy3axWWQH5jcw/mdWO7TFCLlOK/64+jzBO/9V8aVuwfMWpxFivjWApu9m
EozVLlhvQQIr421/xQzBUivgjlt9+HjAS2sqYwOlkoxnFJnOap+STfk4ZKHcuDownSkIhnk8eWRi
YrvxP94UV1l12aYcvqYLgLe/tUQI/J6+MSjtI4CjSgEfUb2caFECOmf9w8xExk+s6Txu65q+bDjv
ZX4TE0wLYFbeHpckfm/x4FNYTd/G8jYdKz8yeql/IM9nPvYFUWQ5EPxinTnd5bFaAM6ey2iDYrzc
lbhypGdmmgyta48rqlft68kIcgu4ONVFCnEqTzwHbszRbdASPdaPFuazEKWNdBXM35j9Gpc9VEqT
KFKPtCG1DQbZEqkzBtnvdcJ9fI2RyoKHGp7GJ/2L4z4+u4RzsOLqlBtwwX0BnfqbOal4Z62BDHSo
wSF5fGJrxVvSmaW4bebphJsOl//K0NIL+4ay7YbXwF9XitFTMaasxlY3fyJQcmbatmRX6R8UmT2t
kASSORhfIfpL2OqsxR+5NjADCDJX9Ss6nWoR4AYdD58JhSxISqd7bIH2M7Ru3mOyiw1KmLwCIK/j
6ihAcmV3fk0S/7sqZIMqM2ZYWVH1Pcq2vLAA8sF98wNW0A3QZ1S6WvHNCUrX6WRAYjaJqAvhMArm
fasnF29hbtdMbOBbTM4BFQFZNHHNE6t73vvykZfG4pNkgwqzjmSZ3E76bOdjnSRU48QzG1OkeHNF
I3VEu4LtGlqnM1vho/NKBrmXlcSnuxuUskqwFIwwyts8fowoSPMfgxeX8Txf1WwWPwhQ5uE4oSrw
R5ALFFQ5eYVs8HQOHzcNmsKQOe4mlSWkzPoZwUQOszThv3p7kV4Jy5Hw7Wjoi1VWXfmGM6jJ9NXm
iD6HCL5fINl/uZwTxDmEYNgx5Fh7Xl2LwLDpqo6zp4DNU4tKRd1mC5P4GcUPFnCaud08xdAw6VKU
5M8fMXwD+csjUHLReQHMkyPE5PoKvO2Jo4M5LuSyUaXKdpRK5VnWYKdK71tkPWc9HRqe54QZR0db
jGoRWbvOwkV22kV5X05FW2iXxgC4/eMhXDNoOmFy4pm2BRVRijoaxvM2PF/5K07F8xYDVTS5cLBx
Nysfj5IILWoQX9bDxGt0r/rcQL6GKpTBoUbGOzP3dnt1h5CGFxb+RIifzxgzcCUxSlwZwWu+8mhQ
CwE/0n+jaJ/SnoDUuagNY/MRLM/1C46d5C+zKAkfuWBUoQo67r9YKhDXH/Ll+K9WRuSS2UZA5FmI
GjqPlA9trQI8TvFhfqUOkCnE2Gz2Ut3bMUloo1zuVchcPEy19J8dkldVL/E0eE6+TZOrBMPq3L19
1NBy5+c1EZtWytfdXOA+VQ/GeV5ClKW4aMQuj7t3T+5+UzLXzki9ZYkEu34RoMDjndUc5oaCyx3K
ZdVGKy4XMdQjIXSbjCbALmZmGKVFBil9PW2CVEa7ZF/S6PFSiSQ/YtQtlIDsVfKb+DwzAvYdezjQ
sPYLBIP4aDMc7jA4SgeH7oHs553wQXg0F8azNQF3seOs/I2EBkLiAIg/bS4DEiNFNyVGKtlSpUqU
3lW26eWO/wr25yv8RUBMpxVO7knBvGqLU5zdG86VuSeji4zkyB0U2YpblkuB99ZXIG5ewerKKA6w
l1JW1jSJJ3a5zfY0dhsIA2wcdb3D+X4dnkQ8j33qkNOv79XC+uY4D3X+eNp0WbkYDgHDz20q5shE
c3nqg5hhNMzORTA5iSqZyMExSGtj3NoHzT9vfE9GWzu879P6BcX1p5nX60ygTKCIm+QvhD0J/vDl
D+rNcDPq1Ay2SK+hTYvo2RzdM603tEjJ+nqVzhZd89lBRRl7q2ZEDPqyR2CGav+QlwkEaY0jP5+j
4GqHVvPgy5LS7pJBjqNG5u86BAg8j4oSLAN7wEemNNLcABM3JUF0EyfLQ3sxhFrvpN20G1Sdh7A0
JZrYrqRdKEjsEjssV5FvFINm3da+GGaOZgWTf486pn82ek9ooRs7x8qPZAvTUV9PS4rAbeZYO/lH
E9proTBBgN2WIpcVl2Z5jZqUKmY8WRRCqFgibGOQ2JEn7mvIMk0usvUynsO/ZXtw24DFKryzlA9L
vQocMeHrKk5NQecBhKKM7LxoucP4VjCQIaCiI8I5eMSwwFK6PdY4FWQyPzlTqD0N3JZQ9cwZRY5B
d8dfs80D6ljBw0aGJyWmgyyB6rTDtu8m2u5JD/G7lwBBn5WVPKK1AgLHpA50/V2Vqp+OGSU0DOxT
8MrLZNxnctffXlkcdffEwft6IrnJakFvhogdkJJbkKfD4MrnhOQUYxw34Lz2cUxdp565QWxjHe8/
hoTBAQwuEDxyr0MYl4CTtBr7/b5vLXfsOr5LAXRpTFfct67qVtb1zkuoMqOsr+FmRf16wtVOoBlB
ZSeZY3oPQoA52a5DTzGO09hrevTRDZBNoNjsiV8OXNjWkiedEt3u34nihP0YpB3ZJTKDT+DuryRb
wv2j75KzGRRtwiSmfqpKmUBPBG3vT28gBCTiAzF8iptqrknJO0Pciqjk5M9iUi+QuTD3RjbFVYxm
e5UtCIqVWB161WqaXQBvHexPZqGPm6gXsIpw1/9HYcj38yRlwiigA1AqNW2MB7isri9YkNxKmwBI
FM62SrYAFig08d4Kb5J6BqnLefgRl7TIz1ssoJqdR+bPX29m+Tz9y1K1aLDOYMfHY7DNmJ2jz1yO
HClmVTy9RuOhzgmqNQhpcH1by8x2otPZOo89NmTxgg7sSWWAW1f39ZpUTBKSEvdLDhehIrVjSjTy
GeDMVX6au8HnJ/qbph+KJymWjmQqBdXWxNDIkFnxYJQrfKyX13ADUYfGCIKFG+cY+FQZN3Rv9fON
VQkC+qz1mMUTHLubzquKO23hrYQjIPOqBnRmWa6TdlditHs0KFMG424iwIkxmOLPrKXnoartlUmv
BUo63yJmc1q2PMI28w6P0tq95ZikPxbVKNTJPMBW/SaW2mMT9U+ovhLWz0PldbXLPDhdQnV7adUJ
1ayc0VobMQncHXg30Kl8kWWN3nTC7IsYyB9DNqKLJeu2oslwqYe+qCtMbUViUgiEvloiciFz0fNi
Pe7Sf1+oTkuUpPLmkeky19ijcdX/CD+rETIiwD8j/RL78PobAiy1I6iyX6wK7oRHA0x60IHi5Dp2
1YbNqNkpNqPETvXSXG8zkUdBwVVnK7GkQvLI0y2djfd/3sLk7mL5XNoh5lAjjENcDryJuqv9b4L3
wwR4Kp6YZQeQU0V2YgXwrEBVi+csO3ftRG3kGnJdIsFklWW6HY4wlprC1WWVeJtsTvHZgTFc4Lok
3upAcMfVjF/OvD2MJUURr7UKo2rZRF9pj0Mdryfhle4AGoqcOm1AFx7uvrF+u+pNErJeXSM7i6/m
PVXNz8tiGgWJjZuWnlDdCV7yDBWytthB5Z3gVEosCgv3ObbYImJlP5gqrBaz9Dj6BHiY6tl6wXZd
v4DYOc/1NNfPy+T71gCfmTA4sC6XVkNXZHVw8tT+jMI3UOn9Zo0HH7CoPxOs2sYTrTuMwyCIpIto
dXT0b/KfqyRZWTh+LpPvVYrhOZcbFAvWLBKfoQD/olKMt4eufNxDJBK7pz0zEwkZn7LtWSNK1BVo
KkDedxROLQMHGPMKw8XLTCKTMevAiH2nq4dgadcxcj0YUzldj70l2mhxNJS3D2qT0tGzWFYFod+n
jdc98xWp94rSjbbSDl1NqYOGUb2zPNQXw9TOc09JzexGAF1fXAH2OdVS7lR25jcrdehAlC5SaFLc
liFhQylFjwhFW1JROn8Pu5NFSN+d9h9s6E6r/50eb43+VdJVFe54iapl7P5MU37+rcrKyvMerM1T
W3SVWx/4UJkUx3xkLNLE+RzlmaFkqJgMl63NUV8U8ThtBZBgpkr/64Z6W76xYy38OMsvJhRpmr0C
dlUA548Jc67WN7OJAcxdVzDNx4KJjqdy278ixSEAlZKesMU+NS7ARpykhgd3dKE1LE4ef+8+9iIe
me0yAfUX3LP5F/sjG+CMEzFUVXt/4JtTb0L/DXJ+PPkAdhiKQVSFNegw/286rswfVaSLkSUCl6lC
o6GvEJNnaKzlyjCtsBXkKJPAV56FIOdGlm/RDQt35Bpdt03Do/cPWE8L7rp1OYvdqOyF7HNgvl58
UwmPlBfdKKriBLvvF5Uv0m9YygOYgkNWVjVT8L1tmLbl187mbcQgS3oB6nCOfmGKEPzvm4wJnXjl
k6YTrOLHMoE9oMd7kzZ0i3Xjblxgw8OUrg1ER30q5FtkcDrwxr7ZosT3vzuaZQGN7CYhev+aHeLB
97rLvOc1TcnkiXbkF92SYxSdSJOxypna7epSCmXTnOPg2sa/dNW9vXrG7pOVqePuNOqlwTRccIj2
nVj9Ts+ZIwJ97XzcqxtGT0PPAobqatTCQhrOql5FMSZxvrstjGxwVal9O69t1ihp036bfdOlbkUx
FMMcJK+2fq3da6P1k5mY9In6ZirreUjFRpmuyar9Bh5Auc6mmQAIJuj44eTOTCy65h2Wc88WT5jI
i0vwW3gGEBDZ4x2H2I2QAtbZRx59I7R+42yQpfhSTLHnvKB+5P3UAOBkQ5r4ewXTrKI20Ef0vLzj
aFqB5Iehc9AjcxLBipbySwmayEycFXNTq+/krE+PELrXk4QsFIxyMeWBXkRQaBxXCWo6Tw4IQq2L
NMrmWR3qQ7Tn1JlCvzfxRG9wr2cBUOEMKPZtqwil+wDR6qVo2rg+IvEWLV0IxuMWtxR9HIVHe5sB
mUJlBYRPLTo3DHM7lMPZJmDx5mlZmOUVtC/F/GRgVM4s3VmvDdEHmd4uG5OWMZzkiJ6Vjy1ePou9
590aG2BelLqlmLr4YqTRANoodyHAj0+9d1e8Rs0yTkPBu0xJmxgTP+0YzxdkaId4AihRUDVzwV66
0zvZt/CEu/lgt/Ytm1kT9Ru6kpHJV+YA2o7J3lJrlBixWhCyNIwCHikYUdDXFGQJ9Ht7WBB+sHB2
2PhWqsFH0owVhAMiviE0YP3vCjXyLayCTm64NOmrfpR54vWhwm5DbuY8bhv4rqM/xx1sOLvfgvVX
Lbkkj3rm5iCBUx99l1te2Ibr5BNXfQgAiALFK5CyYryJq8gzzKikrwsuUH7Ko0/vWEsYyu7fDoDn
GfFnaKPYIKM7rugtgz1KIk+TJaIoa2lF9GyEN7bdJ4eNxMI7P2oNRKYL4bqZiCxfsLMD26n3YgdN
KyKgXcHDx3X9cvEUCUw67uiMDsRq+LWrpQOlOBJAs4Fs3pRVveZNE1i2jAJ623444gC7CpPpDPtp
0qdYnCGOBY8S/tDGOjlnQxAmzC2AoC1FnOXgwf+GRvXat2qfBD2DSvD+xydsDFFoVQT785GzyVKE
eLppbzKron5ib0cm8D0zixejScwXT5j/81nsNMabCPB4Gf21+TBFDfPzJM4fpNTnLCHWbYaLaq/m
8lfC0MK22AF8wZqOUr+3GVwZcrR+InDND3Lrr8MtQfABFkdq6mNy7FScPx2RkdMH7rGprxvB2fbn
AOtaH+HpxtfPi9y6ZLTMIjIiHNCD4kY003KKoG0TGMnpki4oVWTMQFtGxBgU53mhEfTe86mwehr0
t8xuetLRDIqTupVGCHmX3HcAt8mfU7tEbVv1nJ2IQTS9ErAPktnAGajdbA8QO2eWtM5xu5+UHRTN
gj58TrCfQQk+nzUCQRXeBRdRX+u3zKr86pIl0sVYXjFi33O/uBn0d/mU5U4Lny/JWg5G7HAYZOfi
8aRTHLH1MpZhTfyOeB97otHgkX/gNBUZo1zz/WirtcM2z97f3aqzv62w+zrH700vglXaP/tlj+L2
TkoUhz7xFjBrQCu8tfoGE9zDhOr9zrOOEuOsmvGs775s9vcq+K3OKgtiNtITOgcfk+veK5atvZLg
FqGdKDiOLTiCwMQVO5Th3ko9ZlDAVqChy7AGvSl7EXCnNklfSg3qw6PW15kDc9kTOInONXFtSIKb
6fRhQIHbku3yz9vD5LiJppD/MUbcz3SS/70fwBxvukUNKhchXwf+f2amk0BlRfgh9GRcTltxgDlS
1rNk9hF+xhCAm1NTh+HSuIpZ5ElAUtU++kwH9UJT7JHBM472Wj+7Vd07nOtS83PwLZaK9A2V6pDY
6igVvtNyMrtB0UOxCth/bBSrcc6MQtmHuDlNSP03ugipgktI41DPbUrt25BelKvKyd+tKYDjajkY
Q0+ezgGFNR5HWvwBxGJeyuX2FEw5bch7EY9YWT+i3Yc+bo2IwzP1LO6f8LAqc63mnmU8XmakVH30
l302WLglNtFTkPRdkwndCQ+/cYO0rwe6RY4RXhAdIk9PSS6tDWzdrdybIb8Ctc0SG7C7yGnOqQGH
gS6bkkNBHtyQq/2x4wMjwk+uPigmG9G9/eWoPn0wN8DaieYhm04BojT2ooFIl2SLjOCDJPUUbSVr
P1U6YU/8aBqh6jH4tZ9JWy0Hjwb1ZMhk/ajCNuD7fPb8UxzsSKo0I/t/mQKZwbByw32GX9opTNOt
YQSGmF9shzdeNjjKbbROcdniYakAaW6lptQSkl1SPJws4JlmAzxwPekbJW8vuRopKDcbPA2JqXnu
f1xCSvIkULz/XxHa3sJB4hhWRiE6Sb86GjhHjx2GA2Kg0/VMWN2BTzqSorWmgt2TWvgjRRM9wNam
NFl4PXLVAoxXgIOLmOzoL3Da8FdTzyUyH2Zr87op6oggOPNmr1R8qNhJDDLMotStLc2/6b4Q+0SL
y7Elyv72+ZbmExe9zZWQM0WL1Yl/BhHg8h8dHEJokk473rQBiMbnSjldJAz16pMt1EZ6NGGBZw06
iEya9iSAwUlrj0lsnxDvZVYqSKZ1QRHlbyxMyP+cIpJzzcV7ZfQ5umAo1/DHLOcARZKBisnvODwg
t/jtSIci79FseLTTCqSnpYv2HoFB7gYUD4hi4jKNsENEqNUEaxAa57DMP7s7aa+Wnmo/2QeKJh83
+H17ZL8F1k22TIMGuoTKBWJZUoEDaeKrCFXAJ3gE13x7lPkiwZDB3OkGKY52bG+W7bfCP9w4gD17
mfhgsYCUVOsoniisZ4FcgPUjex7YeUhNTc4d/C6Jqztct5Ya4dtBxAZxqu6EsSrd6G3/v88+Prcy
RLlRgE0lc0PhutEOJPhRhoNJf5he3qERQMyS6PliO5cdJdu88hPbHKqJPoa/PsDnuZ8ghuk9w6bj
wfST3ztgnFVCj6pxnJ2ggLvWzMA44tIu0tPGnCWKljUDg1yVtjuQb/mnllwxBg/jdhoy6Hds0+ii
ga9Tf4npmYWpMNDSO0zuk/NN+AqPFYaFX1jcqgiUl4rPTB+Xs0OAGcKxMlq/JrVAwqCEbBxQuGTq
UNNBVk/0Qzrqxy6mUhZmlT/jsXQGh03r51Xu9dv/9pUj+1F2mzXQWfy94smUKFY8iXXQAWuT9qeu
iysgTzKpwvgAvvq/NqgnMGI5+dT1Gn/fXMGrxmL5PT0K9E9GWKLOe1rj7RcyUIj1TAxMlurr97lf
ausvAU3n1P3c64sm2mt2I2Ei1tJJvEKcn/pHChV3e/6in4TGFQ2shnyWX8LSn3tPpQU/imVdi05x
RTFPYn3z2XBw6FvS3J7LAM7aJWS1Qj7AZnF+IK9nVgcGVeNBhI/BEaSdbBf4PbIUYjxKlBvSrypl
grc+1biAtWopU/Zm9Q4hxJghBRpNmscrKyVAivJvMr6QJ5jKlhrfDE/FWuUrbZg8omCydS6covTb
TAGqSWaRM1DVBL3AFxSn10qEwH0laSBbTQOEK8KAjHe2vlEJCyMZzNVwRD2Jeb+xUpYlwKsgbfgZ
CBGuWiruZI5pLZWHmrNjY2pC0BhXXvKIbu2KpopvC1gpmh7IvnT6ZoOwo6+tjH404o1RdDshUinQ
FmNmvksWYuerTv0wKDQivD/5p6zRSuHU9fhS2wByqecNEyVInjvDfPjXZXp8E64Toe2FkIJ01wZv
oouW+8/1Q3RikhgjIrAvyY63Ej3kst1IAD1UDFuIhp8f0fCOM0iXLVIKorM4IoUPg5nwBSt3uHfd
LeT/ivnz77MFa5cmajzFaubL5nasvY2gMbEaI3hrmB11uURQL2A+sPFZXbUliQA80zh8ouCzxCaK
pRCpO9jfilDvd3+fInKV2Zsl6SIjuGJQf3X5xtCO7uKzJMVyEMtoLEb2M5+OX1xV5GLhTsnwP3TR
MwtpCTfFmnXEd4tc76RtUPqX9x8Kp90d5JjLhqmNbEnhuZKQknNd6Z2EJYnjBGtPwqf4dBk7Ko8n
O+LLEz8mPGOehNkmuzYTHbRZpX9N19RVrO4mIRP61I1LP8+QHQTXMigmmM80sgQm1IxgAYy6Lo7B
Xy3EgKQyLWgr2LyAS35vGIzhrc18ZDIdW1F1aqWXQVJDENWaFqFOnVVmuL0AIHeJv40K7Vklqk9/
bMhL/7cNQgPTNiAQskw3NCd9Rq+xagR1CuRYaY0vvXAp4mUIp1ET+dfJWP7ouU08/GEzkTPsqbv+
74IOZzFBGXUhfLfowdpJXez1jCviEiBAS+KFk3HX8+of6hMhFSA5VCKbZSf4q9lh5pDZyFbGrBSs
xZ9LiNyWGNOiI2IKsyZtEw9xf//Ja2A8J2LZ2zRdxQfW8nZbekCMgY87dnQuRkw0oKl77Xd1/7OU
YhKuPi7XpQtZsbjA17D5ahq98twJTj2QNcaxtq65j49sKyhyuARDGG36EkEaDSp3RL4agU7LOQ0q
GA8Zhvt4+ojioPJsmKDlZCUNhaJgEZcgzBJAOsFXWsn5Uis1g3gSjm/WD7j0zTdG3lmCNgOmun7j
9/eN8FWrNfYgQUYK5laKcXnVcSipA5vJTHkzFi+J0iP8LUsDPfGCyjNsQkbIsFWBvNMmgQ1iMIMn
Fo5yDUhZ3V74o/tPXuCURy/ncVGeu3twQZsH1JwMzY0kScnjQwiha+1S5GowQWBbydmgLhtgoEwl
DC14TotzeZqZND+otlxbXSNKG6VQ7IjZJmhBMvh5zqMaPscJiPYxvsPl2QXVGvowiNOIB16xRp+9
TFsiSz/JPXaViDYoLk+Yq68sqzpS/K8IRqiTZuw7Lb36wps8eZdf1cP1LWU5eDyLQgbQ5te4hU6/
Qatj06lpthLZCHqFRwMOr38V8kU+7iLO0GABBkXayOmgyI6asJ9zwNqPfx9BUR1fm/ASEJ7UQWDk
0BQJ7Xll/u0Vhz9NIBB++1HdGFifiAE9klQ6bbGPkXwHx84aCShu+W6kFKSXJbbwJXJ2wz21Uc34
65hwUViLxWqB73Cb3EfMDIO+5Vs7+t0XeYCDTBw/RPg8Nhikgn2ZBkUmoLxq+yXgkYxQOEPWX3AM
gSZ70LdWwgWsnIPd3ep2gPXTaSU6L3X4wpYnKsJ6E+/L9FqR1cZorOQJjW3pEHOhMHQWKDgtgQl5
+TTgoC77tCK+xmeAVzg1qfEt3PWmT5PkrnMyBYsC0Y42+ssavbY5KbcvlYFAKn5+GG0Lyp82j7rc
Vc4EujS6UClQPQkwvMFiyqNkIAztw+a4oy08w37yF9Od82lyNjVXcsnsWHaXCrPS7XGsK5qN/FID
U4OYHLEXcic+5DYeDKxw+WRnIEoJvtYOpShQUltDs+iJLPhRVN7T6EV8uCM9dBy4+9k96xh6jwt0
jCw7U+mCNv0bXor2iyByhMgBU6aE7CaPneeovnF+s3eHDq4sUbExvURyo4W5EIpnB7o+wK1cJi/a
pHklONd/r9mCllofO4CpApgYzlnJEKbYkBaw7WEjYN8C2IMKrO0WrkeuRQ7pTAYiwMk4tx4qAus7
UpZ070pQyR5Yc6UmmFg88VMxoh3FG3gctrq2hGEceu38xu4TNHElISfgJcNs/Zui9xATa3VQxucm
1iKOIrgXU9pW2RsNujgHqvngfNUIL/An/KSnZiXyQgV+IPzw5wCq2Nr3dmkRwot/PYsEAfEcIMwR
5kvNj8IjWOtR0XfU71PYFU/D7oFU0HyWh5GPiiOujZ0Qs//AbQBaZuwIk1McAA4kQYIimADqaX17
WJoS8f9jCVMDpndMcDcsW+IrlKagw2qH3ZWzYwCrBjYwOnu/ZnF2LVonbzfoUH5N4HyT5PD18vwb
Wz+Duw3C8oRYSS7HSQriFODnuo6uc/ZhhgsCJYzYcPO7+MsZplbs2rjqcRyiYO7k0jAvHxnvOT4T
ifEziy/gsg3rZ+xDUXgJg7RACdFXudP9C+A/t64ieV+m/05XjHU6edHMxKmi/tgJWCgqejqQbYCw
8buTDi/VPYhKumPwBIxnkMAKkgdyVHVT50OG/4aYLqT79Hg5sl6VBW7UjHwWJeHBY2CZUDwNP4M2
AKhGgAkpMY2iAebmZNX0uo1VZU6Ff1OOV2rbqygaZLuCoRbMcNU6ZOXx1ij9qm/MTUB1BjOI7syu
Aj0fikpSnPaED6fLEbHOlyLuvpDJZ2KSRyrX38lzuqpfejRZGrbIBLu3G92I3Ha+J5vzyRfbS2lw
54Dh/QfI8IS663F0ZIa+RvxMdmKsszj4pAR1FYZyXqxjdPYv9PQJLFlrm3845sAPfg/ct7JBVCac
Jpx6qE3GkGNYRGJLWeHL4/esDEwUDRfTWi+Cg6Hc5ZEBfyBXB3cJDO3jDFkkHST3VtWNLDHqYPrJ
T9i6DdpYc1SETCsuqomNnh0nBaItWooVqjnUxOGjv23hm619GZPAeDV1juLudtwBiUnIDn57h/rR
sRiUFr5SRzHv633ZbxUftGwT5DFTMyCRGiuIlxgsOvFHgNwmmAqNud/5peUE68eoaz8gU60BRx0X
fgy3jvGNTw6XaIcTM8pPtPBLVB2E9KQEK+UzpvFpdZTWj+12gb/YLrsi+9V43K4jT7j9VKQFqfyE
NGBKUZez6JyNNZzxFBRcnBv/lD9yKDkUhdGT6GwRxQjmwZ575vGD1suqClyo94s+waZEAQZG5D1w
HUh1zMMT8SB/9PUykPnqspLwNXqu+eWweryF/qSUsDYdEGXpsaZ4KEJObBNoq6jgaDYemyr6rSUh
V4wsaRnDoNUNPhhVZ6cbktREfraCKk/qfBt0Eh8LzqYBEds8rVH+8MM2AY8Q6zSr3EpTVUMYI49A
NdS7XvlgHXKamHg39kQUz5BaxSi0W24kL0cuJkBLmLXfRtd/tHsSvs1pB+76x3UQ3QcL6TgI8zQe
Hy9Yqwbjey2usYCwCP1rsd4h1yrziKdptVuTV2zgVashy6p8OY9QSGcpXFx+nbAPNoxjQbU4ZEdb
agvWdER5i6uam7GKaCpoSOqtz4hmYjzizB45r3jxJ0D7g/tOM7MVLB35o87e233lfZyi/5DkX6xx
JdIn2ydJqoM2RMtJo7Oz6T6vDP0DebKQ6CfTcRgMUn0t8XqYaFPcwV3qqKPfY8TPLxXznI6ZA9NG
Qm1NHxV7HfC7DyMBOv6mbjkO9k1Jr2NDork4R9MMw3F0Y5Xtqp2LSWaZkL+M4ImY75glKIzcMCmJ
aXq4r7u47gVbn5DTQoSlGPHSusEr5KlmQwBYGAkNThPG8wzOK89rFNCRXT0eutoRcBbsYqMgp7u6
vpzpC48p9LhAjzPWrq8mPgbxsR4Nlpd/BwSqse3lgNQO16j40xu6pluwMOWQ/u5f70vQeOckacl6
wCqSku6WZ0Y9ebRqRJJt6VgoUG2phVzy2o1ORpB3ufqoUkKjGTEeFd3QZxBwqLoD+Ke6Sy1fROXL
KMMvy9zSdwnhvPj2IOU1f7MG3m3NEaQhXzpGDNWxVuntr/QgHnDdhsTfdZovWL1Lpyyl60Lvh7Xk
tBPxUjbrI9QDPo8siktxNtMDoAxCn9TB+DVeovFerJSI6AN4wTewHZ/m2IQIV12fcYlbVQzkMwWq
OwMw9D4WgJ7RvmzRpGWL92jvEXPFxtnYUqd5dBmRzG70Q4GrFwtiKNTsnzrRFhSDUInQBOWS+sNO
aI1j6MFV303PT1ZkvyDWqA3UtSeOA4lc5nhrV0Spqj47sSEB30VeSKDjhVYix4rZGhwpx+KCxL+S
+0t1WteeOxaGrKw3KbLzkWXq+20saIBhNaz4l80gh1X59zM4RtwnjaZgMYreLHNyOLi8bo8lkIXy
WmYIm0qkzfDu+NJZRDkJiSRX/mnPqmYgQAr/XbajJjc2WbkPKXlMHE2aUvUip9mejwS10BMOvrpA
wsFlGEO5hujHxYjDgMouxGTP1qR4fU3IVn3DdLVuioAx6nKpW0kpmf3Me4mwVJxCZgH3Cb2LALDr
7H38jZJApl8OQ5bUuS82Qr9YoOxRapsBKThn+mL5PfDLmzqv/dm/Ro5ZNrtolGtlYnfSuAvMJt+I
p5lPeNsmpMFrDibU154LUDmSvsmocdlE4EnNMvmySmZ4d1Z37kUW0o0ZBEiNMp73neaFC/7YciDJ
W6VsYL5YB5uzu+m4K88Y/twKLb9CH5pMnQ6VFWpQuvs5NwNbHr8Z9QYK2QeejB3LJ2lGh/G80xqs
0zmAKXC/S+p1HFljkdE4PUSfvod0X9qCqBQp2n9WLlIoPBEIg5B1DMTcnovSObmdil62Z1r/a/z6
HhnOw75ZHcpdzrl8OREStqV0e3rUcmm+ntz7rT0oPriCmlMw3WqTBvymMR+B8B9qHyA7LMve4Q0T
2jvazQdgL7tIDXC6MtMKoGfAnMUpmhlezO4AyzVMGzZBxZJfPwzxXIhEouERzm3XFbRr816A9LZq
eqj8SlW3WSWFNmTCbyoICiL4tgmGZADKk996HNlCEKyQgydZHseLj0re5jWZUs8bR8L91QosG/0r
ojOynrJ2SyIUHvvQZny+CR6ZIWOVjEzM85V7N3j7dLWopj05WrIdpGhNatoneLjtBnygFQCwXV/B
YSqykMVfzPiVZj+EVnXO/oJnMFvr/LvDV+HUB7uV6Qd4aSBxWQPExh7NV7z/fH7O5f+28fpNQlX/
jXK6ZK6e3qwSf+quB8+XOuips1uMONr1ndgm8PKSo2ifkS5cD1SfAp5GNmFiHuj79pwkW67d0D+H
0q44ZCMmkEeNlxDYm0nWCW4Z8gc3Y5jqLjYLstllj6YG3yqKEomG9MMFrhpdAfEqk1yKLIxbXSWi
vxnkxnLdfU72VVrfF+Tc3Oml/d4R8GnYVCvAYFgUMbav6ee5M6oqouHdjHi8wFnwNnogdzhVdv0t
qoFuGtekS1HTh3t1Tb8kJwOunlFaJWOxSVl+Emtz+byy/6rIjoqocYAaqfvHYSRIYss4mkAcE60G
/uDlAX8EMVavM/L/MaZ1u/5rEU7rjCRGlFfO3HVA8YT8gWvDTW96dW+48sH+AjiCNuara1yDqGkr
kO9PinavDhccD97MlR5zLfoldFhD6G1g+e11Ml9SSEwJAzrAZ/y0++xvHUITSTDlRbow0xzhfbZk
mFV+6l3pJIPPzkg2WaI61x+fjJYg03xbWQvWBm4nnciCChOkJVU6m631m8uGrDmvDvR3ObOTImKm
AXxMKjOkDluApsxZpYkwm/7UGme8+7qFVOiQmDXc7icl1taDYAG4JXTVwMOxY3KFk/1V4Q2+IW3P
xgXicd19T5bxXcKW0+mDh4G0ODSGQoXCzpFqVfB05SD/JQRxKFpo+vVL/Dho9N1H6Yqst2HneK/z
mrpORzw8ui3MdI41y//2XiACPld3zeNwZc0gZ0hZn1pDBU33L4iaOTq6UQJiaG6vsIHQcwwVAa8r
qaoxltE5j85UR+jGWk3Jx4TfjJACn7xITn4sRkaT9UJ0YVv3NZz+mGwBiGq+rIxnhYT2+tgYzea4
FGfA4ySxcQBEJErnWutpyjRxC6HeAYLTdgUoJCITKzpDTiUwv96wtYNtqiljdEWH8Tx3AtSsBrVb
OABw/5W+z0F64nxen2oukk5TG6EoNGVBfcfmDaJAWK/YfBy3sNWJGLR6KVItV0OyHvgfyEXNels1
fGgyZsdaYudb5UyeiH8URRoAijNOaMHVFKiL4bgp0gl3Nq05oah/0z2sABMQo8ezi6bUL3hI0as4
ImETpj9RoUrrtvcx0T2YF7UJT2Eva0C1dtnt6jys5pUVcm4p6BlE0LyDqMF0/2joq0jwdX1p7Nhj
Wvzk0OMylPpjnfUZtZX7y2l2O0EZxvnkNnysAHFkKzg9o3dqg7XNkyBz+b2iviG7DKejJdRqYG7v
N0hy45bKV/VJukz/y7Hfoq2/cuMxFI5tt//c3RKSSZAcJcusJSyNr9Ik9PcfcBKYSAyeBknirVbV
AvnvTK0Wk42Sg7cQ9X+d070sdkpGAQULbB7nCOJdYRO+b/DR+gAL8eipo/V+91wz5tUkfsYzwtuJ
oRS1MnZTsJ0KS8cc6yISElW3SBjsM0c5WiVCJ1cARN4KraNJjsAphcFpG6SaBlGy7wdcPCBdmUa3
LNKQ5GGR4jPm/AtYS6QsgcNEXbG3X4BVAlVWQB1q38LuYw5boGBVl++SQiLrJmdqxdmV35qUfahC
eAX8Uv89mNzE2yPjvlX8b28SzeU5PCiPHbS2ENOLPt+DQUKYXFTC21Xz/GxWSjzy6/l+OXTPJ4E7
qTy6JZjMHfGEasNK5V4UQ6gixajyPgVCF66eCf84Wz6gaAMcdnTbqQNTzKerfAwWDaOIJpkYJNQV
TxOJGjtKPmx5E4h/l8aqjlmiUKES/wNDFPHZ77UOIZapycouYG0fpul4h+kTpEMjQRi65aQuyMLq
mBS++FApTlTePsc4V7h2C8JKg4Q5B7zAHaGbh4nrkXTho/VmiUN17leitvSDl05RXTvShz0+mbH1
YTlhmRe3KCGTDkV7eCwDaa3uZvkw0v11mBdWH/LJjDiWZ7Fln80g9e1xojjdULQWYYpULKgMa5ns
bWzm8IGVgVQ44C1Zm6GQy5TgAPPNYjAGigYG5UCw9OgnQpl7dyoGqQpirhCzy0If7UI3RbRw9Fw/
rdYaztS32QAXo3lxarGuUghC5FUWADafAJ6DVYLXOCyliC76UH4/PLcswwRe0GeIc+mXK+pXKsez
IrW78Naj7LAUvidp9UxthyOJObhaJpBD0FocsOBRWB4Y/5Tfd9SFF3XWkV10bGeRJJ/+BnMlf+iT
jIfV7RhV++IbMUWEbvgz+6ty7biToXrBDirpF5kqjNTy7WyvBJbwIrCZ5GW2qiNcQc2+10R9L4cV
7CiqcFjm6n6nNpfrG5Vupob9sckx18GyrwilybUvqi8DZ7/iTgiDGtnpk6BAdoMEx7GUGvsZAlRV
qmtTrOi3/cHFmqOUTRHpB6EthbpHWCRZMWgQlvPev8fqpxCngk1czwmX1DHjHSdhzmjIPY3swaxm
toxd4dmqCm9xdZv0XKQHwRDPmw6lr0fnmgzJyyehWF2pydG8zCDczEkXQ83JsMjj4LZErj90sn+4
6ICCx1t/pt3/ZJZRAVRseuT+yIbW5GqrvrPr9FLwN4WPiw+NKgCMig6VV5YTc7VI2KEMzh3wf/OG
2FeMaP+Rjy1msiznfhSEh1bf3e/Gc/mrzcMfFqDxf74mBFRZgzSJpvsmKj1OgIf177QBt6RDcElS
rTNFFs7HyIdLtXaWsq24kiWW6PZb4eGcuUO31NNEVQ8i3QxJnDbQefB5oOYZSVdjTef5GZoEbJ4Q
5cEo34R7/ZAJJG0/qYU6sgVhvIy1WZMeDrhNxzkoAD8Jr5GoeQk1B9ptkfwyBW23eQnAAnBFd2M2
/xaZo3Xqj1KuJdHM9/Pnf1IRaW2jt03lyOgPxqwnCVzR5dRu4j3efWfiiOjuJUHPK+5L4NliFLIf
8U313AFGd5gSCS5tFlyyiDrOaeIRCHfimIRdMNlFByzwyqyHEb0b+Yk+Ibct7kbAjG0epy0mjjhE
LtGJe4q4hRfXlGnyVPqj9zqMuWHn1+USaMvhIZt+Dq5t95Z9BrwoLICWYWsAjPhUqgFyKHD5GEUZ
NTfpPH4FhNfemKxe5/ik+XNEi3K7lKS2FPdBtz4z+PNstzp+sngwkih24w+jb4lVxTaqK19VgJzL
fW26FFjnE3RWb1ljuc3nuegddmkkRERvTN2LWpwV4InWYLL1o+Zgnj0kiQpl1svf8s07C/+tZd5I
LLSF+KND6d+QbLulUg97o9ufdqurtz6EwfPXuUAOt30Ay08ahxhzDPE2MYIEI95nMUVlqoKCn8jb
DYATNPQb//kKo+vyr5GYmsWdyYjHjuVxlx1pXCnX+gxIfPvs8sbcHQnjWW6qfZ2FaDDV1fpVZ6eI
Fut+zKEYUtG+Dyh+KZPe/l44fNkjK/m/SXlHpMqodFe+tk/1KwcQ/KOSrrN3h68TOa9LvFWBhww3
gqd/eFUXqlwplsCnpsGtrfRwS/oHqh1BTQQ76xxfX03KWjNZsWhI20sFeX17ETBe/+vzAgN6Cub7
oymI4c3as0xViIj0NJqI2TlYiFqvdjUY0YgtGA3PedhznkzpTdW+xDcOVxrbjyXcFc0XtQdZdPOH
b2DrAqH5rkiRxC2Rci6RWTLWWMKcQW3HoozqC9Oy++vIS0z7ImuGTeNMVTZxhwH8VXtPeTYqyU89
At8xuQOwd2NlbjaObEUop1e/S7PqNDfXSuv3MY7p8tpU+haHyzMsfuycdD80hWVJfm0jdKc2/PsP
anPwcRipDo3v1If+vu4kLsDzZmOTcy0Wa6F9L0ppMx2X48gm+GGNzEv1qnyjhlC8CIXkF4kESlnK
EfP/LjuiVBcvEms8IjgUuapqjcbk26T3rfttmNKW8EgOwn2ln/XGVdrkW8OovQRgpXOYioT5jhec
XlAu/k+Y8Zr8LZJgT67bkXWfZijCA7JUSzi7j/f+5H0jNJVC1RbBsdl+0i/uwbhNdie5vCNVJOrw
5SYJ9oxMmQkkBaSyEdeC2MaY+P4hzM0KoNgCiEQoEWOBspGbo+z98MPVyobuoLmVqVSTFEg1xkex
4CpDzgDLG2+olHPCgWM/P6FuaqIlONfxTNE+HN1YIa/DQoRzk5J1zNQEIMw3HvhRC6s49oB0Yyvf
M057c+RoBBFJQ9H6WSwcLJwC7ajUTpTJ7WKOX1hYx8CGZq8N6mJu27KZK+xK/2qAFa665ahhAeDh
9izK9iu1OtVUTIR9cNAVggDXwN3jw7/Sr8yMl6xxrfgqSfvirzNIYv5gyH4wZ52gaSg6nVBIuHjD
LiDd0aH5p9FIKQWd9YAQs80+tAtcUqJZd/Ccprz7tJKtdd91ZjHuR591KNtz63YlZrsfbMTzw2Hr
mGquhbB8njMWYF9sBhpx9eEDc03qKmWq8Rg+vRVHvZQsqf8c5HpZ/louvxstqD/BD+UHHQMxureJ
bPdZgpzYvopqSdIVWOqvlGEuM6WRRHVAN6qiXMaNBOaidyZsHVMhZeeK4BqfcZBQMkFKapi/A6tZ
w0fyWIJJB323WH93gjwP1hUdopEcxPb+NSXjbGhobpXF9b+k/KdHdpeNI0mXdlQHM0yXHh8sgtDL
XdSE2VNMfMZgaUK6DSu9WFEz6xWQDuflsE0b5rHn86eHOs19RBcjCzsg9WnZewwpy+7G+4PQ7N4c
zc8Joybtv4uvsEsu/10p10uyAtkrK3voVUnNrYYP+sNIGgFhsddBQC4HQAvXl+ZHtTfERN8RGT1/
bspXyvqMnEJGX8BQ97Df8tXRk5P5mj6TUBTE2MMznvwtLQA1eZJbyHkdDmRxSgFe4e9TMCDtBKnH
2sAfzwH2SrVXZwN4rKcMPXE1qx2kfur4mT1Um8xArIUZy/Xua1jKhgw8AP2UbWtyyFPImzcaWNIY
pTnsNL8WIxaq1mHtJIrVrjhuvOUc3eFoyhy2hMz2vNd6x1auC8w+w74NqTPZYCDWAKgqnL61olU1
VFSZAngYXJMe38JQXLNxGy8lr1aX2DXqGuOO20CADe6e5OnOngidJ0AgHkR3T4Oke4ei4ioGjH+/
HiCE1huMSQCBLoLDe+q/Ebxf9SRrGozTtSezNtcNsoC5Av5ZsK4idAzrUc1BYcaP6zVjjYVlZuXR
viS33MqnvOzZsbHSXXEQrYb2pbPPF1/OSzsfZUpMojROb5w0Tn2YDQQ0U5JeP+X//8l1D5YeDggy
vaNxfpazUsnOEmQR52RRrju/KQjkw8xSW950p4HGjvhW72bBfuffvtaGPuBtNlJ7svlM0zNMIdYS
FRsV8jLIBDCc7976mH4tJj0KyseCsehK2OU/42K92CJGTLGVBfmlTFqYoGSrrjnp4IQNGbbAYR4x
jLWArRM+YZT9bMqFm7/tRF122kKgjb+w9idix6mHXZaH4LlmajirTrLUKvJT2dGyAZZjoWIF7gR+
pnAycqBS/1D3RrVBV2DEITh5KUP+wlaDGhlEFjADMMPblKzyzMCGaltkUqq/BaD4+0K+IG+TwX0i
CN4kh4r9okeVVC4sk9IjjEvn1h0wx70j2qLx97x9bG9YAFq08izmx28bxI/Y0sAtuiJRkLOdV1Qd
njTP44eZZEydpmZ+a3pERwBAbkzfOsjA7dwVIXgTMY815ZRqtNk3p0GingE0ol0cSMZTBYtXd+HS
6UK2Hxak63U55I9g9MegAbaZSX4HkozmBiQpKQmRmv9nBnR2la0EQZPlE4N4o1qTypsdHf0kNQ6Y
TB1AIRSm8xowUTiPxgHegjDUpTgTF75/68OwML66fLXU98bNNMCMhxq2FOjvmgGi+TsLKE2NDgTI
AAU6TkWhO/kI3Tim59PdeRidCDkBzAYtzKWx1+EUFycLSoDX7VoI7wCJNyGb6LzBtTdDF6iqEZ5X
xuUpkXeXonkyEYWIwJenYHLjAZ2kH2Mefa9U7hLerCAiGopd6bqTHmtmWDO5nvGBE2I98FlHZLxO
shv1aXlDf5slQVgSnWLOr1+iAkrjUrbeJBOx2HziK+cj7H/OwBHlU23D+ORoXYBDjvD4q5nlA66s
Zlk0zm+24dCmaUL1H1ASdlLNMvPv0nB1N5R0h6VpnhCxkKGTXKApcU13DLOvHG3DihWJJzIb7DOC
5ySPXJScvY1ZiJHXV09/Wma1gh4Q0v3sCj5N5yOZYwQC7sGY+0pjuTcwgSk5VeKqqOI6rDGm/dn/
9oo9M2+ExeXPiJleN2wbBIxU6FU5myCmhuq6eNwFV/pIz1dy25vduWajG5RUEZJUkquRzrj1aluY
jbhRh+gp6cfozTVN/kH70t6/c2E6LnGeh8aMHL9R5s+ggYb7KIkiceSxwnHG2ckkVNkBdozZC8nq
CiAbaLXJXiPngyOMjUE05Pp/wXW8EeH2k5Sb2mixhtl6JoUyVtMO8dVqSfIho8ZmwNQfsI0oS1Ir
s0zmFuNHrvWwTXKyadjxEoWoF/9TXK/XITRv+MPCMbCKC8pJsU+XqMAMa+Rrg3FQKSkeejit0eZG
Ysou03k4M43nSbIPkMfyvZ7t7bw7mt9L+Hxs3LhVpWtwzfRxV6MKx6fKMuCZewMk/r46FkKyXGlf
SImwQvbobYR7MouQWi8GLMPrJUQ2ezyd6SIob4zBnWlGnbBkhy7BQhw95t9XDUeX00ZlN5Ax3v2b
SDKQT20APYNabXPkwCkQ5nGUOd8Ie+whJ2p3xuQyl5SHjvDFpjVu9xDUzOPlGgXyXiZq+F20wEtj
XfcLWUsoMh/mA7m+tc+hBn8WxZpEATSKhVFQtvpEEmF/8KC9ipjpa4HHIYK6MoNVhfqCRGj6VgWw
85LN1GC2J9JQXRLkLZfCGvlhMEKl+gr8Rc3ZL668OtasVV7f1mlKWShFS3/DI/FvGyJSySxhRz5D
Up1Z5Fx6J9tCPjVsTAHcmJUsmuVSyF35Q+qbheJoKln3a81QbKp0MFYzENQyc80kK2Oo+djYvfrs
/6exJO9n5Bgw4m40w55aaMQEO3Co0oTLtk7l5ncUi2pNNPAFx2pzW5FS0UG+AEy3JQhVz74/LT8a
nSVCcARtKOqiDUwYLyWFEG1skcZTo3XT6FfViTlTyY9DE4gUDgHD99Pcn8o9R7ywteT6C4b4ek2W
poya5C432NtQn20v4XeF1EfDuOMUkcTw4slMf8m0/8cC8J+Yhs8O5K2uodZ99vGRP99b1LhFTBHK
wi3RrHK+1rzk8lEb8yQo5oC89WjGUMxv7W9KJ6yK1prJnUg8162bm/6Ryvw7UgoL7ZUJIu3YjhYt
ybn3FhPgTucoa3n7I0nk6NkPx0giIYsoHv7+ZOysDhpbZ6iF+4QXmgi8wyzaBRfEDK8HrJRpO4Bn
n1J/+F9SpPuBKDoV0/wFKFel/9YDHeUaZPJ7/Gm/s4VRQySqkzeX3A/edIkqHuCIJIcbIoiMg4UI
VxWqDVNd1cqZa+9o3kBuEAlYmttxnuudJKnuZa0CVmTaXgJCBg2brbJpS1lgOErAbbVP6XRSHd9R
JsnkQvQdMsr9lDjqk6+V8fUqn3I26lJznnPBoH+oBeNg8bbxE2MlYPv+vqo+QF1oFUBF1QNSS/2j
hAh1E2VohEBTYaf+oGlDn7tjrAvGHJBS4wQf6Ze6NMBrUOtcVMT2FhK/ae+0abUqxD2H5sa7SmkN
bCL0xsg5Ua5tpEAn3efyGIw2o8IjVrjgBo4loFHnRfaZoyvxpMteAQW4FkA9SjIlvU/mHV8IWZF9
vQvBWMysYetAmRt51ukKzM+BHUGczrbMEZ7aZ7AAsO1/71/ILqh8UeUzu3OkVOphAG356VelDQcu
TexxNqXTfOZovqvUFA2T3QZU8lYT7Qbau283OZrDrOPsdudu91juPwoINPvK5FG6goLrcPLYMvhf
6bqnP9HJyI1khC2P3Ry0Y6qjcMRwdchRWMINpt+CYPiUyrclH3INifi/YXyjOhSrSrDF7RWgUZyj
d/5/Dee2AUDt9i3Ygq+hdkkH6kjMge1zOaYVDUstaae56kXcyJIWdVdUhorMxiKA7SkADW6Oq5VT
/WrcoZPigR9LU1kgovM61a6TLSEeIZFW4NoBeloGGN5GKJYXUYuOIKSjn+g5HEi72xl+plUrArke
N30gKrvhK2h3DDd4bWfUCFT/gtunwE9B8pF0W5zi30AnEIvZkaEnDJet0BPiTQVDvLQQhipZDkWS
o1z2ucAy4hWOINZXD1yDQ/qihhdKOxaXsDtraZmyJl9pIjQLjDjNX76vW2sS3dFYJUgcKdybLng8
FhwNVkPkMRoW1cfnM2TikCyeej7K3FJXUe4FSweqsFpc0stzQqu9hM1dWOW360saiwJsAzTWVFtp
OlCxBGgPNbAmUgohy/QlUhtvjRUGHSDOMA+5QvnaRwaVP5qFSVxv1FBJmxk4QFZ3+i0Wz/jAoVgB
KClcxgxVhc1lg/ihHukQiuORzvOYCwOeYyf3Aowv58XIV0LUZqu/KRTkOV4/o9BndtBe9PPzgWKH
4mG7IZ+nrRKE6j19wID/5e+7sfUvdzol9NaFCSYTCTn9/lXmPNwfiMsHxH4b2Z24KFeGb9OzaPkR
gKfEXZAHVSEDt9Lz74FslW5C/TqdjU8xnqk69V2n4rk27+pdcbdnsLn1xFYZQeFf9OGf6MrMgzAO
Msmzfi38A5JNsxHbKD/kML+QQc2Kk9ZzEXkAMY/+s4tnfnICa+NARTJJ2eNPXf1chP9qu/xM4jpj
aNuAgEqrezn3eXT6u5Kg1RAZHv9LHsPyNhAsV1yIuHpEA3UgxJsczN9qWNttWHductxA8i0Asjb9
aPcr6DlCW+ZVZ6xf2eyppPCRQ8D9OCY+98h7jG+0ctq48EcFaDKJXub+JSeK5x08OI4cYu1fVw8z
o6f6krets9dPtz7Zpgx28V+dC/2jDclYBHVUynoOu8mAMozSR7xYFlBy06j5ZUP/HWddnUbedzkc
wD9Ub13JjpWFQPpE/uME0hYGNX3HRt35IeHGa03WnXo2zt7EB2nakoO1qIlTDSonmDeMoHOqn6e8
AASATRYVGvMhwvFfiKGCI7JsJV2lDVhyCYK+0VIC8/8VCAenWQwjF01m++95NW+TnaN8wrjP4qRr
uEY/LKaQD7YxcRpkAePQTJj117h82EfRTPzvuW2VhRGndPDq9lUlQEtz1+b/uNvslbSHaU49SOze
KL15sMnk2jv0wYtvW8FK0SSkIqAb0Yti8IfqpO0xzuKCXct3OEt6O9/8Azwc9fqcDQMTYv+lsEYe
hLnD1fXzNmi4npW0GwCgeDyIoBXATOLRSCTNVc9QsST2/UjlM4jS4Vzq80W71G7Zz8eeUAEJyqIh
OZ8WNQWIwQXayhpMsWUrcSwnyIrMbsvCNsmdt6WskPm/FVQkzC3/TXroN1WRu8uEJ1F+NyP7aexc
h3YKkRLVsylpSNq/SEvAcmmkftYhLP1n9nEpkXiRNb3p6uCvL+SjIKoe4ryXFUMEnMHaiiiYb6OF
5Vs9KGMeUWzXmrmOmP0WqpbOT6L9PrpBBlNubvok4yXOYwdllQRGI9F8Th4gXBY0GW9qU9YK+l/I
XJtFFNao/3Q7Mp/MERffQIfVAG6zJLOS3FzWTWhRWprE3bXhqAjGjGbhk5KUDoTLzjpA5x47ru2y
W2yFgR1yFuNlk1hxzJjRcqe26/uSruv1DXXhl19hUItInbUSMLxpyUQhTNme2MRetAjDYr/2D2oN
hWGUXPttJAZkGKCub2zamsSXrjwynox1iHxV/Zr+vsU1H2BO2uaDrU5zYiPPNjwvKquCv0jEYRk0
GAP75rcbaDONRjY5GmbDFhqkSXuXJ/Gz6hSl1BnjQI6iS6XagDuhCeSs1ZmMLJ+1l+GgLn3UnALM
Y2zglfjJC6EePyVMwQqfbDgGadFDIPo8caRrpgHqbGpiR5vjilJ+dte4w7zoWTca4r/Q/azUxAFM
pFhXyCA+kaxLPlEsAlJlhwqj6pU9IcMAlOaAaBKN48s3qDfgMvYFhKdXBcozhBSLOjD2NBqNLGtF
oVxBueKRU44epqDQ1xfrqxnYTZxzRDG29i5Fpm/yImJt4XKwPYz9FRjiCPSpqAyDT6Y/dZJVDHmB
hVcwserAco+XvCkOwsLcFTsMs0B7nlZCeXrlZmwtqWZQjC6Vqv4l+lkEGJvxlFDEetvWcJzbXaX9
ycaF8sJvLBmimnW4qoyQHzwbEIJFn8WdXT9GvavQ3ENNtI3RU5TuNNPIk/0vCUSg07gCFppAkhxO
acdHAyIefrmmUnt/csqYUKYTAIcqsECz5Yj0jiMQSfNY41G9ZyLuf4pZohz4GI17B0TIitZby2i7
ajaRvoJUAQNg3tYVJ+ti5kxc/pcGq6+wThDubdYr8wTX/v1i4lS6irm9BnxoIuPovrshxx96DzT2
P3UfTp4E/ZP/QTnU3Jeqe6NLQcF7icdGbtX+sZyn6Jdgjk5YqkJNAB42QGKc/yX3k+JosL+jt3m+
Er04WEG+JvX2y6Dfe0YmJiSzoPUU5HcyNx6oEZ2UQ7GPxBt6sauBIEfBqABKzIHd/cyD7D3qZNa0
PpbZ1ziCe1MxYYfGpgi6SF3Uol2J/h/BOEkTnYU5iGj3fYsEYJ7mcedkDTwzikwakysax/Qyykj/
BrX1U3GCEmkQ3FrGlENjbtvVEeyhS8qYG3k6vvbX6ZfdBMduqnu+siNsGce327ibhAa8RVEPGXKY
EPuT7nZq6RzoNl8eRTXPBJ3qHzXt9DkQIDE9pb+2cgyi/MvkEnRYtBfKjIz6T4I2c0i7UqNBawJC
6wn0PhLLh5dQbxWk1E56hUfDJvo8gYDmJPoMNmUukR+LJ6+bddBDDYl+amBpJKKXR1P+IzWa/DCR
5eX/LLu/5OgLp/7oDMB5lXEuHkXIG5LOwh6DGFLQa9ku0OVQOPAeKEZEh6RCs9wmSyCDEuVcnYWw
xiDUzI6CZS3cGByHzwQB4dCVYoNhohWgfvfZk3yVCIxaKkZnxmBzCgTV0kLFaF6HSoK9+huRfZs0
TLzVud0lZ1gW4hXB0rWWwup34sqYHKhfMtk6+cKTl1A6MtMyR6ggIpGLknbnhXvkZjG50grjUUO9
qeFmvMP0rmyTlfyPXcR1rfvd5BhmN/jDSg1uQzjL6D+C7g8wNLX/abVPzxu+5A0LinIyFqQx8s7K
/WTQ0BXtWClXmmhi09XTOd4yH5bx1OEnNz/2JrkDx55+qq90yu5T8X1kx4Crs/cvSFEdYgE/WfNI
tnzc2+qPQRYTcsCe0VyomNcElcMLQ8vzTtPfi1HBTbtH1de7vLsOyPurdVDjDsJItW0MNOeSsqag
xe4dbgCB2tCuSytZg4SK7leSJ4g6xdJ7weNqJZ4t5OppKRW9P2pOkMhMHK+gywy4bGrSKnoPdFVG
tew1X5/AQG4FSTZ56FnghtG8sCPdhP1tywwTAtdLyRPh4S3fu2JU6uUEbEpRHRT7b7FqY0F66mt4
In73vW3wwDYKePPtPIojnqkmW1i3nPOHSxI1ADnTQfKdmkbJOsrYctRERAlQRSmMgOGBs30mRLTE
EgLT+vcfTSsVfsIFAH+TjExgQst2dY/okDDn7D2NCjYrzftiEfTvIOe5YV7vY9ZC5ROHSNYUn2wU
zgk+r2hYQSsMan2xdv2LP5rEocCOGRumUgT/c2QdQPehJ5R1lm5naB6jDxvGpBdeHf9Tj84e2eAA
aSyRCIFNOTemJCl3Hz6himLHOZoawkwsl1pEVJVPazd3Rxy1FRYgd0SPIczTFC9/dUyLPOKeKklS
Z6k5tCFqCOnj3V2QW9u31EWQe4LYdMPuPIPcjiR2ve3xfXB0uPvOBzar/hVWs+EbXVHs7JH3nkp5
X0DHoWxqWZYB5NyAw9wPGgRloHI2sTwuGWehEY7e6TYIkQkyo0fHPTJhG/4NjzebcBmrcvThGURz
jQ1Ipd/o6nEbvCheRMMAGV1WzH6miyjvmSOvIaaFm2BOe/x3c4dXDqKWdd8jXM7OyQ/UkW3HXSFy
T1kP3hpiSeCyWR4tdgD3rvtJL0lva5bahHV+ho3yDsSpeiBn0uGmlRGbyH+pWZDnlhvVbfsk3GV4
YvUvfOS+5O9eldkdcriLp5AUrhw3pwFc9zaj/GGyuJ3t9J39aL2qGnkFliaBPHjrL3Lt4xjXEINY
C/npCRvDBahN23DIX1EHn+VFxtQbcUoBFpYqUGKZ8Z68Sot6k6vY+9ReH95eGB/vY2EEsnY3+KCR
9XiLuy+oZdFK+TXhWBOYitSQ7UnvefRwA91eDU9IELSD/2YxBsd5Gi1jE+URcGPSLVcME6l9Y3h5
mMz2FOzJE7IskrkwK5xWZTIuRJRgJMZnTghWcVMU7+xSwSg5eclP3ZhX5A2mil6DwRHULlWBN88Z
5SWjrMnLU6+ZLLfZnvyda3ChineJOfkdN4AJ/xLe7nhDQKyzAZRDUwbfn9cIkq+kg4AWOPPhk1pj
TPMxduAU9RUX1A5ic4oJNR0BEJOG+dyJQwpiQkNJsBhzHcBNud1Ta5PzuEtTWba9dNYTbSlAvqZT
XSIa5jRAGWldEzaSAoxVgxJaX84JbgfMZFPQ33GS2rFqcrLxK4WUvUClX85rbCjtihWTRSXKLBay
uX2MD18uxSk0M5uc1HrQY3m/qWzbuGY1JLarwwekAH7j40feWV+KdOSjkQxIlsQgQJIRfIH9jXnz
qXIO6kGz4OTntNqUiI19k08yv8IWcB5Y5pBrhr3EePVz4W0qFg6QSei37iqTP5EBJWf7YmZtI8pR
q0QHfFciKUV4fwHDQ+WGdnRLcxMA78ufX5iPVN5LgNq+Ac821CYhlfqyuU2mXM+phtCjIdCE6CPj
3Aw3rxAe2s6n66DguhGzm3f7EGailR49wWFjonq5zBkKIV79enPo/dmcSohUbpXRPKZ+a1e8I0wa
TfZuNAtuXDVpFVLSSclFXMOP8zqUGlOwK5xq79Oy5q4Irkwplj/DXf2GEFKLKk6PK6uZQqjiis7z
yrR3sxWfrkeeaowpY4YI1xxrBmYBD16jftLjjHlSH3nlNBQ9GCqg2Fo9YxSZi1gKQXpUBJfa2qXy
k4OdWpQ/dOpYAIz7/BbXA0AlqQGot+PbI/6ujvXX2nFEIw2QDVPEeptoRecnQppLzqFWNr+giJVG
n0FPREy1iQJQUJIBi6xp8LdMpd/owl/m6oWL3HyPs+t6g9Tfk2eSrqRBpIEK8gELgwXgywFBm/L2
1RJFiazADfC+tB/QLWJR6vwIOZlxtX0ZBDYzLXMDIYoW8oAQz6/s9mrJbJlkpDfPod44KU/3Yec9
OSzg2JPhyX41nm1wxuP7pKhf+rbsQq3n/TiSBG4cAYlmHf558AhQ/SMWA8muK10rgHGSD6j4umcR
3s/LvQZkT5O842dSyNffuPlHk3cPfXbxsp7jSlqt7dvlj7r51Oik03wHYyQS5POt+LXxQvQgutwl
AqIwSqe63T/qy447h6DPJn9w/9SDwwxSO5h8MUVqVJziofcTnTZvUtEddNJ5tl6zOB5LQsdxxOEW
UnFEB/vttoPO1IYJOoq8d91h3/qo6VxMxpnQQSFC+9oesETG7fXDNc0+5RxHjhI09eS32SB6I7Et
xl1R0DYmm2CGYTNrpeFV3lVkSMIc8/DhZcANMrPAH9asj9kJPmgeS/CYME1Wk5tMF92X4W/0UqRt
X3x+kqTFYwRq0HAMCVEDbEWCOtHGL2GA0BH3qz9HkuXo81HxZL/426066yLRSnj5NfAdlSaZLrJw
cmzcBxpZzD5YwMx+vYvBieli3PYLO90MN+Iz4vkqSdyEaVtNKREkBMpZfaEjPr3IRfEDzRu6uSfl
Ilvu1+6PHZtJq4wKP4zziKCgkzYkywLj20aZteBCT7duWR8G0g4WlhjqbsRFo5rpYHYuqTvC/9BO
tXtQq/3cSqijhEGQPmI2ELYvE0dn0zRdyw0AMs6U7q1ULDziXVvba5i9S17eEkf1I4Su1TxsNTBL
M+l9mANT6+IW+3nJaJnD8oHjziyucMvgyzmezy4yRWfVZwyB/Gc3kyzCcxNkP+x0ZE8sCJTeEbL9
ZrzJc57u16wFcdPftAhQNTISeJ40VfwclYHoH+wx7RyUxM9fdz8rSGzkQ8UxHq0TgJn9cFS1d5nX
qKGYahsfpcXfxNmL9DWcEo647OpE79hkhLjf65b4AGKiownOz4miAuuKc3nJWfts79dqaIJaBvj/
4F64dbBYTL8mrovBoxCqQLlGi0LHSRATOGYD5CozckdyAt1rZiT3X3GgX5kdtbExZA3YTFZQEeTv
ZItoxtBhlQ24iX8leFdkNrQ/40MbWcRIoOW8EjcEwCB+UsvNZEDnii4sPjpTyxsb0lovL/LdTC7b
LTe/Z0y+Jru6pxgJkLPIGv8piCdyPg4lVQj+DAaZ7M2O7usTfsC2sCZtsLxlBTbYAueGWr+pNluh
66CjBXouossi0vrWytkeuJD+InQVX5Za7xKZNGPbOt/LxQck+LctXFlTs735ZWDO8j+n9TV7OCM/
hUTxelCBLIcZLFSicgghuIfjOmH7qT8xOdnDBJDv4pEZwfYv3GjA9rQn72QkF7aZN4Q8z52I/tZ7
G1QJviRNnEMpoknTr2x/gI4nufbgWDIZ2kj8Tx3hQnaBZ2dypv1fMtrNqM+we7EYVTuHVAUOpC6e
Fwz/DySVb0sLmrgmoza0Sv2LGYDN7V9RCK91OF6eTY4COKn+VgZKkVg2/fvSdSS2kxErRh5dRvFq
ZWZ5SHKC8gDeH2t49oWdr0c8k6uFGpX1NocPa/BNa1b5hBL7bcBjQPU+BH675ST8LF53IaVzgbTF
OTuNDGqBN8u9Q/y5ank8jdhfF6hjJ2RnfTIwF7fh94F08fU4Hbk8zPesw0LbxLHaoslQGKotI9lw
J0wKCL7qTS5ShtLPFx1of/qgmfwY1v+4FrvWyBwZBYv11WHXh+C6rHfNdQ6E4o3Tb9UhLffeo8IO
1AhXuFyysbt5UEv/LMlddTMTCb+cmOex81XTkJSk0B77h0i4DgxapwSo5MKtJUmfKPBZf3ktOCFN
Pd1rv3V/AFi9AuEbKiORVhI+dF2n6Nb3PI192HpaNaiREgv0GpJzMOhd/d2rezWlojXKOzlBXAR5
MF6XGyu0Fi3O4pGUUPupnwPE+uKSF18ZHW0F24PLrW1NUyJim78qQC2HdYqcNaEgpgCUL4jsIjx6
Pj+U/f7MZiLtBSCV+TC091zLmyrysTUbp1SoJZPSBRf5JvGzmPcQ2Kg5IdY20LGnzwnhsgEIonjY
0n0FZMrL53OZuIkXzyIXu2p94UcDwU4GwG/Ua1/4wZaTVH6d/rHnDi2xM7MSe2YWzxgC/Ilf+3yh
Y/uLKfhS87EE3z6c5nc2D25efl+kk3qHYoPahux4AUHMC7WVz23WEfKpTuuCF9RLEl2cp3XLqes8
FbIDdWDJOG4mgcF/k18bSkXj5RDRc7ys4gKyk+IIyeRObUuBSi5USLej4yl7sZTQtSYyBZMQzmlZ
jN4H1xB9Soxl6m+d8hecj8o+2sTy2RxS2T/fj2JCMblGxzmjlxBOvSZ7GwiMVCe2pGb611JK1lxE
aLOXXvN17G4NaLA+WZRnAd5qBLZOl0SZ5naXHQNvWefASX65pXwZpIauAQWqHomjQxtYNnAEVTgS
jl6+lRtMpPwP2RG0S152TK+QJut+IT4EYLTJQnrOx1aPdnvXLK114Oi74dWRo4G1box1K/b5402D
2u5Q2NHThAunWCFZqCyZ9Sz21Ow//u2c7MNXf0HgS1pDeUNrqALq3W/NHukuycEF/xkT3Pr5dSSK
gpbKV2I7T0YXQET6EgNKzvLwMVdHvcl5ySuCr5XZLaXPW9XHo9OqB+ErkXiBSpVa0n7UsDpANv7V
NVt4lt3+kYDb9J/b5m8HvzIV3ynTqJcaV7v7itCK11dsFn7QREVf+ax2z0bfbuFTUzi+dusJvuU8
KrYaGDu7UHZOp1Zpg59A0Wxg0IyY0YBXfl9l1EseNNeiuNoIZHetmMudwoNmswxVHwLLkoAnSFwa
9Jo3D1/n7rCzbrVQiNsuXGuPIHAKnM7iOZ1P6faJIGTFcVfD835uEec6b0donpJjM7IITckBu3eo
D9qG+0p3WCO3kCI5V9tYdTB88kMU0Tut3uJRADK+s5lQAtqfEZVtaEyfvSNQXq9kj6+M0twBUwnP
bG30sGDnZF/Y7PCU84K8viVHeSgDz1Z+kMh11jSybtEn7GY2ZwaoBMvdxvkU13n0ZRWysJsavRSI
pbRRneY64Hs0NlR2WenmiF8oYk6x9ZwNEj7xH4SfLmRLueO08HykBMZ5iwaXnR/t+6LtyD6umrn9
2YGNe7E6sB42iXEectUFGq5GJaPKsuJ0Xkyzy7VoCzKC/50BLbKeo0ytV+WIG9HvmURYOCJtE4In
YSbipEpGr60ItLWLBstn+3lPRFAUBJ30cVO5IrCX96P3XfdkFuBHHH22Xe6SK80awzKcbF+AeHps
Yed/8iM6RwORZq/PWPwTqdbqvHur8jbuBPOnBl4M0ghaKz9CvGIh9v/K3QPe8PuwiyokRWyrn4lk
yFxI3KQJx98vfMfRLduUZXRIdsvRWDzgk4xsYDngttm+thFka+WYIeIjXIq/xQS7WLp608RUDAVo
zqBnvh88ot/mEmZAMpbgLAQpeML5gYyNVQ8I5i+FwnMBpor+WaHPYjkLrS/3+9CeshaLz+xdC37+
RAqq5NU2VL9tTizOKv8vE/fxmsUWJE6WtyznQKktlLpqp3PG33mPoVU5GnMCJUu4VaVeCPq79yQr
LjaI/B4BJZNnwKmg7Ixr2d/eU0uUaRiqEPYkNg+ZukUnUvbt/WlBBXFSvpCCazx/cBZmYEleHHHx
jjN/1+fjDRV0HEx1BXG5XxiKLt/HyDDrgoZ+E8yQGdeTuy0oHCA22HUsPFNqHGtTdZacPds7BfC7
2SEKM3cASmm7B6EJNgoPLDcrfqerjfs3xt/Tbx0XeqExDfzhbGKQiTvuTsgXC8WU2WS+Pv8wIL5o
abbLqQayrjln6hQnpaBDN5R2f03DBiFhG+7uhdldpSzpEQzVwTSMCDWRTMIqnKqmmJ7BHbQ3DHSn
mI3R3X0fKvmuf+laL4y6w01gBnweLh6XxuCOPBq9mTYc2/XUO++GQoGC2Cp/yt2FqIEUqD8DmDqw
oyELC17N6Ca3xuqyL2XWZpYrzuhKcfOcBo9x7MX5njPiVM/hYkdsu1Q6u+CT+R51MTsAEo+W8Mix
SNoMXPruCG8fcRmvPPZsnHfDvazx8XjpGDPQFH5SMoWO5TPbo27CgMU2lPoSVlmWFTpkBZUweFJP
utJ6b8iQFnfJiauA0FyznNZRfKHC0ggVBXc6vqyz5S5i0ANi8pOClBvX8IK8KkFuQSIlfV/dTguL
/4PYp6guO7bXKpVW9K4KW5Ud/gIpUIaJdG1wPhQrzEO5D4Sq1NJcdo1xngMImrcq64QyiS6z3IwJ
FrMK6dDtvnpoEk313yFc+t/qiQ/hebgaRs1vv+lpiSS/l8gKUseaaLe45xWcmjB7B/W0o4aIql45
MWIbd03wfrkAp3mqE4pAToVSc/l5DEimqQuhoa5MRKWTMjKOU/DKSJv7T4cVWLdyj9XUnLxFWpL8
avMkJ0FiEKhdSKlQStywaCdmO0zOeUNRjZ+Pj4kj2u3sXRPsJa4QsbbnNY0aAbIp+60G2c6jN8ln
RmltUkncdAPUc1wOMzcKvmlpXtA3YbPtO0WisSXb61TnTQzgky6KT1hNd0T3O45YYPj0e0URb3hP
/bkUusQNxKMHov2qEbQMMVp78EjScN58ZWbB4vXkSnJAXV3DVeUKuDwcX9KkyxZeTbTDUjx37fu6
cQclh3A43Y1abdCdqmP82RDE7XG+b/5spHp/u7AsrDCuZOLd5bOjX2DiBhAiYH91L0gb38qHoYxn
U6iXqZfRL29GfXHM9rqJccK8Yf+Uy1pN2OaHiK9dfFsnbDkLE9oElTbdmnzgRCmcU8uenerrXpNz
VBaC3X72Pp2zRZ60Ur9xFq+x7R8oOdXsy/XfopE5ElZdu4MsclsoUjK91k83HGLvdO1/H6KW/YLX
QIeKjkKx/wLRA/WRsD+v5Euz8NHdvTaIN+XkFkpv+yJQCPL4wFcBfX/lIpMv90U+2Y9+pq9KNNNX
jN/Q7WD9IMmL52nc3YcjAYYYFuSN15N4IxizA99qeu7/uP0qgTfn5pl5Ab4sqUFViuSGxt688ar3
pyqFp/6gkNCk8pKeX7NIFzUnbJOZe8J0UpOiNhybCgI4AFLljp/BKB2VhfGgPw/y4tV131VGkjOx
gZmIQjOl5DILY7F8Aqj9qNTa12rbFkW3u2duE4mHSrYCM6slfwXr+OhOBSi6aU7GK8HgvOfFVbBD
rV7u8BY1WpWMc9UAJrUN5fuAAD05sg6+Rfasv3BGeVrMYhRqRDB3+i6tXBDkxzTID/0xfFQnZOfY
4LKeHfCyjc1hALjxhw0vnxZK8QeZsj0/W+kUyu906gIH1D6iUgVcS1U71N+IiBaXFdGKE/oG5gco
tCDVBJWsZX9amuQOWsnuUyWo8qgk6dC02GwipE0CAw0ibJWNgltAO8MNAxw3fQH09OqI4jvoR3Fp
xikqmg/3w+5F8x2grgVYL1Nr4dTzIFV3zeFhNrRh+7M5LUCevzcie1MH5wjhPpnXk4Yz7OUe9LBw
VhYgQmICYm+t/t0W+OxeS1Q8dChVa3/HTxeksVriw4LK9j5cHuM1OtZ5NRTI8eFMKaob7kc7dD+9
4B4fzmdVM+1FDIrbZdDORL+Dd8wXe7gtoZqUUezDDz8ZfIVvBTFPizbqYMucKY9fmldMIJOwNteB
haQatGGlvy4CTGYUSVQHbPluI60QJJOeayoGarhqyjGFsKHh2Q7+3H4tzAYGyM798fVNTQUOay2n
SJnA0emR3mVmxkvGq0P8tNOIMwXbWMyzNtZtJteiSWcYvwcQPSLr1vf2QC2IbNRa5cKA8WS9vet+
3/Mf/BvuIh/hHXZig0LU3B51kNeO5cX7TGaclaABbj+z8ZQGpBZk3yy/1GCrxwpLzgseOEcDeNTF
cY7Wwh6adSrnyHDex8EkS5oBFmhOHTavSEDGmWtvA7Q8+69sOvwJHCmB7iDZw4nm3R8W8Go6T0hu
F9ymramvEmRfC9lJlU/EpH/SJNN4+k1blMNuTGdaqri85LgOUsyD3DMnCrIlkwNByrPCL88RBZWN
+9TQ6xBB5u0bAyjbKFFlAOmPXgpiw+nsIvIOLvZRXKvkhOqgEssd+P43RfGqpl7AHLoy62El+Yo8
SDsopiX/BUe9vpXPdcF7KAWJ1zMt9NtVY/JIShq7/OUc46TXgng3Y6D7xKCgOPPM6ctqUQfaYkZb
U1lp1Ts/x6RYtYTufN8LmJ4EkUG3HOUEhH+CAAJECmLWab7jUggAFRjUBlbKOhbooCsogX5VDrIE
h5/oUq1e4K/eXTXLnOTwsR/5Laz+xYh4INDgyVV7RynKUb18Ib5QxAq6sNaVl7lCuVxwCsqPc3S1
LM91lcrXPdFHZKYOP9FLFuJHR+OyZjguPBKJbpFLPKCb5TyxbFo5ipYeIXj/dKq/uEb9oEYlbakJ
R3XI2MncTNKrVR+CjfsEig/xF4w6/3MqdXSzBLHfchsbRV6LKdSJl7uz4MeOhiZJ4daem4jR+GGc
fOF5EZVMFjgyp3qKykQvzZt+xX5/PmFuSgX6K2ZY3r6Mbo3wX9Go8C8zwyELk0tIpLilYWgZc2Xe
BwR9iWDUMqsin5tPU8YsNRz/uGB4Kxw4XhGt3Fuw27cDBgCES/JLXrTJcIZMn+Ofy3Z4jO7xgznC
Je0xBjOHvkFv3MzEJcvRSUKwbkD0iNLYBSwNDpoSHt9qXEePQANJEBxvfubk/D5J1eBIN3DRgVnT
n5WGzhtqjiSn+wjbScsHNhNsqwFh+IEx6MldgO8wOfPsqJ+BxPydBQOhdTunREpiI+erzoh1FhGc
49A/M4Lhk0jHsO+DTFUTvHBB7+BELt9A/ig7NlCj7EkTsPjsxrcrdn4NOKEWdMYoXByNeFeC/ypB
BRvPNg1cJFMCq09tUXOVZeJ1EwatxqPKEFTKPWOUIKguP92e5IaRe/07Ry3/yp/Jo8MJ8zqbvHtJ
3gryhefm5Xg/RVByiip841CL2LzoP3+FoRBHfX3sFQLZkW20xHOQKtdkmrNeVhBzMV/Hm8KttAR7
mH8bTDIjpVuHpSsXr+ppo7uBfNYDfRWzSsxzUxe3Z4V15cutlQ8L1XLtshyPEBCqHO/WGnDLXDwz
+DFElweTOioJJud/XscwRj8EPSxLEXSumXhqs4+ym0V3tnPiPo2EwY3XjHQaoB2tixjjyVrJRm7Z
87TxYCsp73vRyOdwK2vs5V1IKR0cLOHJTFz3UEiN5QiTN8yQWUsBTOAN1xiXpGnKQiB2S0zbkNJv
lykTKs3nt4fih37GnuH51alFIQizIw4v282/HcuuyvnxSZYbu8i07XzEb7vszmjfRbzGuY+Xfzig
OAt1bkbqWvT8rBYdE1pipaY7C5OzI81ynXdXshCr8ksPqTL5TuLQxO2JOlKdnRuUYt/w7ptwpzwH
b11fpJtunqNKizmW5BLdNhZpY60NMn4rQIPTFfvoi7xit0k2+XL3nlGLPFoCI2BJB8L5EAJ0sn8m
t8l1mD/p+nfbEVpmWJmpenmedvh9tV6mesOM2LvAoWct7F2zHXea814yNcvp1+CJFitWLQgxRa8p
zWWzi+hjENoFTZxhB/tpWQUlDSQu00bZZUWLIMeNawRP4ZwdNdr18L/0tziHRO5EZopiEyMROcho
hSrAFE2NPU+Ia/ULwU0I22eZF4rdrBfNLih2FhCFk6z+3kgzYhaI+Mi9oxhECzaBteL5VT2iUKyz
PaMnYMZZMnQMSPIFllrZTDYROEG6X1E3fq209Sa1Kkoe7AbUh2RjKZQxuXxZ6w+N8zjY0/eITIiW
BMhakyJsfoz61zL59lb7Az0cfEKYmrcKPKI1hNRFAwKntREeHtB9f2ukOHHz3iJYFSZOviYD610X
GlIPC5VsxxbgWP/POnzNKVEOOAC12EfEAJzjTyUNEpT7begt8XA48B1VwrWIu4VqgkoL78sZfESe
KeXjYQDB5Ycdlqlw1IiL4MtwI1Gn68PkwL+8jJ3cSwn3qW1LB/mF35tf+zS5qItgo8bMwmy+rgPC
VEQFSdzPO6TzP+oWv9pOndJYojK7AG2gvz7XZwq3y6vBpDypgC7OFxwnmmCGPBFAj+u4/1Zxdwr5
L+N1PHgqsOLaTF0ucmLqePyp1TlBhUiakyEepGBwXr2FJOnTvjlpv3OK+YuUx3C5qBgIIif0hxCr
qJiQfPTC/OR7mQWYUJyV/CyyhrbpEpqkHbHETpprzlFcVbmywowFUtF3GsIullMQ4NJS4fUB0JdV
QKxTqBabmNgg3hYBeZADj+FbreMKRPx2YFyYvlt5CekwgmsXwvx6mbcoGmRoqyATCQKp+qXV66Pn
ZfwjqwR7ALh0mawfYr+kAMQzT+/WT1kmXcc3g0TPGH9X+nRE/h83JntjxOu9JEt4sy5jw3sNwcJs
DLVPc42KotBN9Tm8Ifin1elXwhWbbnVnd3ActqE3FK1B9pBqiINdHXtHiU+eTzFFGnGUq1DdQy8p
phs19Tk9TW9guOYjyZu5Be+jlfXbDP+7xjm1aHyij/YWlUNYlkA/0O/OcS5waN42JQukfY6km1/V
E6golzlPLpnyGlPvqmmM5KHM/UQLvPZttbT8e7m6o4+2TyLvAfhuFMWDvD6sMdIAeezE/y1j/S88
JrlsBIr+tDRXUu5RYAL1l71PTXE2wBhLBqw84ma1/caK8PUnsSNbDIFnV13qV4g+LSk54UWy0/ZL
ALSBxK8CaazWOWSxpQC1IOPHGIMOpSvx4DKfYlPC5gD5gYnaqgkYR2FSOJuSwPi4CUpC69tDWrSf
b0DZ9+PvCiRDdu3FgkJGzKbBVwUWzrWFo0B1bb+DAqQfIDg0PiMhOWgztYE5F/6TpzGb7MBhWCHE
0Qn/QqtC4wx1Rkf0xXx8ZEIK0PwIoxlpA2ibkmQqekEiJw6Iv2qw1ATe6uU6j83vY8mnSCkj+KH+
tJCMv7WENoFbAkOYEykDL/tlSMSdzvDFTCSJPm205sqen6+T5jWxRyHVTTRHxN+so/qRieTIZ/Z6
3wrnV/6+/iRHCOH95QKU1U1sgmwfcRYf0Qrp07ItGfnQKeMDI5oiWXxtjsk3gQxLjqeqCAzY0tb9
uNBsogdnHn1TYw7QdeJjPJ/fYeeXU8aK7xaB/s6mvpwDrucGbBsYdATwYeX5MwFqOfPkOS/bldDn
vF687Iv3Xf1+UC63q9Sdxu1xwtmARYU0Wjxptu81lHpTwtlCva9yy2Pvm1p52W0kWAjNRuY0wxXr
qZXNmNCBmm3z/CckT0GnvW+fZtP/yjGC6uUMzIJFIhWDiLj2t3Ln0JN5JQuYSFmzhM+iYuj8gAHx
J2W0cqXQCv+jI7ylxXgpiKOb0WsYksAJgAW6TB6qLXEdRZs7PFqDndeXjljYf6hziH74fhXq91Sp
jjC6l7Z7AHCCDXvxuPb49Ms1ZgKDlHU/lZmHCvC12bldXCu1/yQX6v5Nmv29L4e9Us8IG+0zc2RQ
VH4Ix/W4ncngUBa4EEZRWsMXP/rNnmnWGAit8u3HDiiYiXcGCX3+7WkN2IimaxDljFrJeu47LyUV
uSIAqfmp6lMUcsPWMfENrrbzFjNo5SzDqs6Emntuo+xzeBEkYhotRyNmzns+GTGhXMkIhIAtzlwf
Wcj8bE3ifkpxRZt0TckYAAXyiFLZws7kOnea7Y/TfZTDpLpDucEWus2rDtdmDA+cj8+3gHmPDI72
IKjvcVTwPisd7/YywKkJQE7rgRsW+WurjGufbH9PMHMh+lPx0IAacgdwatwaf7M1oqNNfBmJgVax
Fi3+lWh2N/Nn2JxBhuP+2wvpQNo79T8ODp/I46zPIhVX0YQLQmNxp+9c52aMSCuzA/OnXj26G6tI
OTIUnLs/56lwefxLj1H8+utdzTjJd9n8lxnLQ/XsOZ3pvTa46RN77nh+ffkVUxVIoVuG2bW0Xc+B
qpmuZ8fIcNfyNuCoKUZftqmGfnQTo9ESgNPdR4dUosjGCY7QdFprQPk2Atrq1a3eP9gt+KW8Igdz
BCO0ft1wgKH7metE9sLrC/vAK7Tw+upWrj6JXB/hZDz9FzV61je7F5hAhtaS+XizuyNTUaw7msJ2
9Om2+cwQPGGX9Ye0Q4zDlVnkMi4mOw/RpACP4Zk0TIEDqKG2ocJxDLODrbfAy6Cg8vDnbMHx/n1A
7scR89tWZqlf7KayNlntctQN/DhkEJlFB0wUentNNa7R6E+mIMVU3AvfbXwz7oRCg/evZ6dtIBjQ
PIYRETCSQPtTSZ6PvxyWWFiiSxqURovjVHQfhE7PjaDjE/rUHv7jYtSkvawv62akq1MFb/oIk6N3
9y0oNq8E2YPDvI7kIk2ykAxxeKCQyLoJR+/BmIHWQv9Lr9EmxgF4lRWuy4NHj4tiQ7jOp/iQ2z/z
fotbqWUnABxuRIb23Xw5IgZCBRmpb1UYoVtZ/WIvf+nVgEh1jriu2sChgUNE9DP7WasCtEXhvE0k
6awiGR0BmBVSJoaycMBXnkuG6vCTbUAipWuK4nfVj9eym2eys2eiiuL+DTd7xXr+ZW0xmPQTeqiI
rnt/RsRNXoddFGKftFeujhXAtWW/bZ+jFx0b2Ut7lLhCq9tdaptNsqvxoRZ4lL1yaZCX68NPPpCJ
nGRHiHSgC9aJ2AfIXzrAkxtLe+esXSzVWzFI5ePMVKPnRYMT98XsJgzdzqjzM/68YpbkUBej3Bl5
aaERheJmcB29/kugjHe05d2aqDmtpqlBKcD2DCVNFCzjK1Kq/03Lk8In5HhR5bCtxvVOTmmAOTKd
vJvTFADOlww1XWqbSKcjaLqlAInXWM3KxYMnTpZ6jLqQPn/4+Y9+d2AAc045+P1UaH90B7f7Trtw
q497VVxG3HRFL7/T9AIobnCVzXwFqx4O/YHziQfcxr8eeaDhpo9WOG2lVh/MyVbkZK4W5ocoyQCE
TQ2m/RgNnG6Rw8PbQwN8rbvYdYKto/Fc2KII7tO7/R/R2NR2SU64Y8yONt77Wrtw8XhPT0esZUcS
rc7B0li8tFZdxBFGEhy8P/V7zl6VtlE7pq46R1waI7wP4987nrAHsK4MHAePu92Mg69SG2ldtXLB
JE1qt3g3EDeVWgcrRA24y3thVyre4KnArREBRUYM2HvEbBQkAjQRd8+C0TTnE0tPNzWIj5JndRLA
hC8wWc+0TvS2yldZFGoFXAdLw87S1DtAGz0DOETkd/6nPadfQgI0HfR4jBpdXOoPNcBegdE1ZpTU
qfNTFOYwIjQfVACmDyT9tCoxzHLx1m305pB+20iWer7rl4NE43AF4jUeb15AVXck3WUktymRcGza
KqQdIpx5tmKmzksO7Oh3vkX8L4G09Wxx1C2hKJ8Rq92jLt+v+mJMeF9ySjSn81oVv2Xp7okhVZUR
38yO2knAPhF+mr6pyhaW54dxF4LB66BGfcex+cFJIJDnTkPm1YI7/JuOtoAwbbVlqGZOP6gDpS8A
lwkxO1juJhd64lMiUScKn2L3QeUmhH4lsVY9dewJpW6nQSjuDwrOXoW1aSLk2pG1nTThjaw8lzHa
Hg9GhSpFQUzYlljKO1SIx16iSUVojBiIJBXyCD9OyU7jc/6C8mzJJ3XE6Wu6yPMl2Dq3XAjMJusi
+MqAOUbkiC2PSlQvMeIcuR/mWw9aBJ9PBh4BBlhVqdbdDpAvUnfqzz+HbGZOdhgRYxc5Vn0x1hlR
L1JnPQtamo26rvzI3eoSWprIIYWfkWzKCHucQWgW6kztQqcF/AaWqdiVk9ke0OlcThkx4DgCQctC
S7dRHpRuirGsmaHA8/6tDlnDiQmKhugAAk/bzlwUJV1UktaCxrkpFfe/OL157olNje2QELgAWJFX
Tu9A/QlH2NlWeGDFNF7MWJTzNES0YMOFEH51PJIeN6GBd6aRxaYSjGuhhBq8K3XTgN38eRYImMxl
KNYvZCyzvEtUWmBOkAQ6FPNkOnq9Fu7sKp+h7PMdmExdkEDqrE48r5O7Gjc9BGxFW0BNaG3DyfYq
4hFGvAF9BS+tpMRyHGe1sdSakXbi1yFi0J/JxrjFUSho7pL7zk/ld+EsSno2VJ5kosOZXkVqjObi
CiKY8K39X7Y9x7KoSr0lYEveba/+c+WxbnPryFWltDWPi4myi+ZbWJ5SR7sKtdFNcPRRZfJBAjqz
uOXKO50mMw55rBjbGgRAN2PONKqzab/ekva07VmnKDlaeaG+yE4T72HmKPpryru8MyowbofsJs9I
rt9d70Ys9HTSArpouhzTPtSRqjN0dReg2ZOmxF3vmajaLeY7jmCnUjm2noQD7LFxb6jFYGVridfu
7A2XV3SqhiYXIP+Sh2tt6jnDpf5a/1kkcosbeJ6nlVM/mHmPaYvFMabOnwdaN6o/uhWbOLyDgqpx
koqc1KH/4lmHnniVBeOsZhumXPpG2Q3lrpGEcdIV0EjKO6EdDtHkkY86PJ2SWgp/DGnuVbAJ0q55
YyDNifO0XOK5CYAVZ1P1GQaKtE+/hLEdccIm7CN/gQqgKWwHmg+8EATSgtQnbli8YW19YAExqlrN
+IShGk1ra3uCu7QaP2+1Vo3faRbUUflmF8gcLkpGw5PR+ZCbMxW76zWeDMHGhKui8ScpQfDVgU4+
HulABjtipQDlcA51vfAUGXTxHmzd9PkKft6WwrCF0QD204Ebtnn7BbxxUrw2dweVqHyfzS7r2HYq
B9srWG1DbEmI+MfMySSsmCzCRugiOlGVnjFwbg6W64Z4Iw96+SRSX0HzlekeDmcLarJpFgs+9QmI
Mx2ddWVv8s5m+tVxXUaCuPCFvlLZEiQN4nZUG2eWOk1tbOzOYWg/8ck+pZPrgls1jKE7p4UHd/xT
JtsFsPE4vD9+kCM53ToURcb06TPhXBhLSvWx4L1rdCnMiuIgboObvffdkTto+RYp2UKUyWN3qJWM
GdcawEEpCsRL8GKbtzA3HjEwujr9okJp4XbeOe96jOl4srZbA8ocRD0G4CQ6ioJlhqWArameW0mr
vXerT2okTMLTGRc408auUF1NJl4w6f7Zm7VTzivvS1Z0AIW4p1f1vKSDjewt8y551VAtOhq/YA4h
Kt5VEh80PlANyefnkDKJ0Wb0+F802mvGcCGgmLXLnIxAM9U0pe3DkOFgcd0nd4SJ2im6T0W0LDMH
7d2seOTa+Iudodx7zmTCynDvEa2LNdHWyHEhkk9pho+JsSLlVh3PbdrVVyEFD6JwEdfwOdWZbr89
i0oNIQfTDF6i1L7ixbac4Y7lp6Rx7eWnHmlbV3lbDXpqhj+xE7XK2UBdtnlJuWNG01+F4ebZKQpB
f0YtsWRbYkZ4fYP1UCVjBjLhjqTdD0v3QCkEbgEUPpPNnxcSz7/qjNmtU5JKGDGgbFPIpUqc/cr6
i+bJY7m1Wlhiv7S3KsPVqJCTTGDyHjCysZl8e6RunmYB/cSaPp46vUN5mcdAsPtCD63zVmh461v7
ZTv+mt6LucUpXbvSgfWgx9hNcX7/lvxwPd28EKCuebreYfxPd02mqjttfaYIBCILWK7ZbuVLwa2J
PtscKLrwg1+pMuCZyRlSfJ0EtR1PdvPU3U/uZcYKu22p4PkQdKIDd1XOHWHea0qWkcpHvCbfmNaB
Y3Z9wboVXFzhvpfbvSpG0wobjuGcnHzyjqp0dZT3/HDJYYXy1bpTEW8hbaJ5sVHNc9i0LOhXeTa5
1hIPsLEf/G2gHG2XAyKODAQhILBTdL7jyRB2uVlXAne01anOPW/H9KYzfyTnbfcVbzKOFhwtjKX2
iUJPqVLuZ9m7LpdQ+36TxxTOH08v9g4R9jstBPvfoMpD86QkOFHeMrdgGu4esyMWoVSe3cNdySqY
Oi+bJnk8BmK4i3YZqqEXd/lk1H0FBDjEl5kViCVQZArLZI4rcRIyfaxCjL8CzVz/9iQicQxN1G9F
t01uxA4n1QNGz/nMMcWgVCp1Lddymz8MhzX1De/y0qepnsO4atgSTqBDIUMJkbqxnvVOf4Ptjd/P
zVTURPtwuOpmM16MHgg0WRTkfldb8n8fV3uXEdXh/UedNiMWZywZJkDM/K8863FpGn17dh8rRaiJ
Ut6pDaMs5tKHsEO2GLL0aAJp4G0dqCZhTwIEnjF5nWgZgcG0bR/yhjOI2bfG769TPoyRo/MsvIMk
D+g3VpvuZOFBMPfkm0LajNqC45TdwIGKUuwSalo1XF3QNCiCrkYZHv6cffesLCyyHiTtUu7Mm0JO
ba4Dv7qG1AHX5X9eytM0ITv/QQMVKn4VZJ5F2RSGe6rw4Y2LZFZOhM/aCKuC+PeiPfrA3ksTTfR8
2L7ioz6EeVEw073B3CmInJf+vDFXSI1yGQHCpLvlC+y4G3OAWdkyRTD+8grXuamKK7JEiii5GyDX
KioPaWrueSi97bRtA1jvwLOc9pqQ+EEc70yOjD205TWaVvbsXTDq2ysa4poLYDO57ojlW8488BT2
XJFQWEzBbwWPtZ11LGBPi7oF0JhA/Rn/SUKZYiz30ctuvSxVTL8LXQIp5CVvn7GCHqKtZvIPp4gl
RQNQs2APzeRqND/E+jDZtX4tT3rp6V9I/I3Lx+lEPNSKTAIgUKoNkq4jResfH0x/jqa9iVojc8DN
cFD3WhC16kbZwcca6jFwT6ddr/EFpl+gxh+jPMbAkxetvKUmljiNdoDo0p+L7jK0q+zBdyrAjS5c
aDKb5MAPFimz8Z1i/NXpshlo7X9H0nbfqSs8TrhI3VrbN8Wv9RY9UKrZjVGcgowG8ky0zafLnsTm
1gfxSuFt7ctT7dI728fMtqudIcbt3qAMVMzFgBU2xVF4LNCqORRBwYaK4GvD5abIm25FB2GPOPFO
JGRx2gt22smdDiFxEirjgjRmXn7sXy31Svvap4lQOPWtRnQPn4f19L8YXsjRBgTXl2SxJkR8HCGQ
7qQ38QKpvs8xeo39hMSvGiEMM7PvCKP+sCXrD1AxHWi10bJAmA+ByV6vsuq8NtUByXSXfihOFxW0
Ox7bVABQEhWgqlFPnaFUDgildJnuQypNFyeQwNGGNMJiBZny8Y3IBbhmNmOcitSC5J7XqCo3u1TX
A5wHmIYXTGP2H7SJ2rFGxfrsyXA69wOd2R5GqNDbRF/irxp5RKS9QN5hXn40CR9iV7f6FyulUgcF
p8WRKt+6r2AQoUAO1j4FrEgRQ40emVRKt/5KNDjSQ22oXA4BcN/A6PYDTwkQ1by8ucNtY/JRKXmI
CIErNel247E/AxeSKMhyLrACxuX0Ur3haBLRz54HbTx00rrf+QAYfVhsgtpbCIP7ffcS5BBkVtJS
Yf2kXfO/Aq4TYJbutdTStyfRCiF6Ged5GYLkOCwR8nPA9O2WfRKy87HDGrFTDhduP1eeIChai1m2
ZggJeJnJffvk5Ia0G+pRIugrZBZenY9oCmZ1f40MeA8gFGjNONat6tVcCC1l5zBnuNBCd0YrWX6Z
tVJDyi9iQT6g7l6WEVPfBmfiSyqWFF6QOT2Pfa1SKBmzYhTr1AdwUF45lWxmoDQE+F4T7CfUS2PQ
m9uMfDSkWT7UWL1CuFl4ZpfuCHUNHA4WsbV6KuaBeKnvIIsLQ7OYhwWh1BhXikqE5G6e0kqtKkv8
UvI54JrAM/xxTUK9FTLDNFNB0Hrqk9pYlNigpUgbkuhy4qaFIyupUaewrLNi5OCzV9ZSP/sEFVpD
YVWdSz48PQx9tlkSFoZbWRDrYADL31/Mt/9i7VdS3Ydsd1o5n8nQLCRuzi7q43Oaqx9JtGCn2cBI
mSVXvhMz714bVLbWsT2bYPxiMf5Q4E65h95pZ0rVI2c+eA+VPbMW87FSoRmF8slgvsGwsOJPBpXD
QY3T1OBCCu+sovDG6pB70+W3WPRtw4XgXpd18qdNK7nVucDj4lm4HVQDCyGys9tkOJfkvHGqz9ZF
SyCgCn9UFTcR404F107E0f85Z8ZSg+ujIKxeoJ4knCZOc6IH4YnMXzIbJpii0ZMmNCPgOOPaXUXL
I1XOxD8bMk5qXTmKolxiVrAbPBVL1eH115HqEZK8yj31W1c6a5UHfmLBpj+r6cXuHO4dkP0xe4E5
ehiKoPSiq/M3UJjjsrhG9Z15yn4QrE2UwMXqU1CiiRRSmZ+s7i11jURW4D5cT3wwQCMbMRz9jQ9a
XW3SqO031o8lOOJMutqbPGTZdmn59PVyIp/sd99ykG4cixEOW/K0SYM/uo2KkgAsRBcZidoy3qr0
L3K4stS8huUs9ha7tGFFiWqZ2VSZF3rv4KRJfyrv/rkX+/Vut2Q/uQpL/6HCajghlLDCdDDJHAmp
xEEfqwduW1nwdTyYEPKZgwzKlwUolVLdr2m+kGoSxAVu9EOsRmxD6lOsaqOKmLag7geBNgqzbe87
xXKducwVay9Eb1elBl9QagnDt8cRIRmHlWsTXuyGlp2M5gYlDexAx1qNa1YA03OX5mYFYYr222GR
lk9dw+9FsD1LWAX6YhemrS9ijB608pUzI+M5bSczvyal5ZTD1Q462tXzIplr7e9JcOjGz4vm/g6m
onEGd+tJ1JBJ+2wtBBVSRC56xw5Z3ms23ZF5IYcpcYFFA/2vquwdbWjx5RF+j1fp4WniV7lkmout
90PLzAPKWZpFs3VqTixZwFROIN25KMnzSJqzkbEpvwApw3+4boK2fNydle5BJ15a+Uw1cCyBkNzo
QNa5/iPOQ6OYoPxkemvpEy/cxaVXEKc+B0NqdslswHW8kto5kJdcd1peBJ4ZwL45SZXGNDjWRENi
5USf3cgTdtzqMgbbKgfieoEcXdNUve7o1FfTGMrK/NUW4R07UWsF2egv9C/B8hcaxAkeXkDdb9XV
tSm72xL9nvNCSSiSMZVN0V6dWVwFvDeaWzRsBenQDuVFHKvApQlkK71f5ZV/RLUEHOgn2ToBpNb/
Q3KcBktEcldzVGJBlJdxkzGEylT9RlgTjyV77r7R1/8ElTWDMOMZCc5cmKdJuC8oUj5uQuI+gHkQ
ejEQ5RZWEI1nTGl6lj7rr/3f7/BoNamQ7iRLvruhnjjcRYqiUvdILfutE6HyQvTOllpWRAqEJfvH
IKRuQ4R7MiTkQ3kvWefUhDgEQQeL+7rD3QDvVXVBjK1RcZVUWQ09ycxoNDo0sdB3lHMHImXATJiA
B/LoYnd1ILTmEkxKK3reVtotoP78EEn6k+fEU2nvWWAXuzWT370HFSeysljAUj7ngirfoT1mhJSj
6+NUwX888FoPE/9uq7uiTI+W0R0nMyImOw71zsDGCF4LZBQOUEvEdYzkZKNEmBokeP7xzAmS2XSo
vl6NmH1Ik09KpnSRV+pydBhpoP6dZIbPTc238d2A73qXHDY73vtmlH6RR1a5wTJZ8SOOyI+r5jB4
BAP8gvfk0cOcejY2GN4v0hzwLFipu0Xg4QTR7vI27W9ug2v8WF9f+mpzEAM5TjyZ4cnUo+Nczioq
XG7WgK7N47BNvqBsd5hx/+kSbdALJtJX0NWXdgFjQCrl17XKNUKDHxIw4OIKd9qRNAUyt2znJFI+
lb3FTLjqpU6djbHrOd4up189an3hIeetzDf89b3E/f/TW3wtHK1ZxUq+zTzKF7qQpZFNtyf5Za8n
lFhaL+7/+D/igtVeKZ4quZzLeUz4W4a/vOeCiRi5OAEvXbCT7HViHKPdki2TAd0m8vvukE8+ZuAM
MOXvuAwrP0tmo0FO8jsxjhQpxF4AV6lWYco7o/vJNS+lrsJUyhKnbonOO4zks5YtfUK5zeupkPC7
xxwCk7uGLXGMwEy3ByQbSVKq6A6lNII0N3c24WQviVzL/WzOnc6Iztfsfya4TLioiTp50Q1OPvmQ
6zk9VM1pI+yFGOzzHjS02K9HW9dSd6WcbF2V6p6j/x/WkvY8BrQU/MUVGCVg+18HaE7qAkoaOBZS
MACIAHBCOx9Qe3gWUDYu32Plx6aGul5DWyqnAfzin7SMulpOgjRA7myo+uy3vtebE+fj0kSHkIol
4mXyuqqw7XqEZtQ9mLRP5JuWTMkNSzHkWAS9SrpE455RSP30kaem43TaE5UL5MoP1zMUNL5Ruchf
WuvadVOBHld0o+XFCHLRB9aqN49hsevCyznZMWKjxD78zr1TLNLeA8IUYZZWEA/tBEMZfnrkocDh
0+CHy+t9p8Q5aYOqYcy9j2YM0Ts/6lVMXoFMM5Y8Qw3cRp6E3JmSJwp55IXl7jXkdQh009BEx5I0
s0JAreXXA1ZKijHlA5MZAV2wI2MKd/0Yl9VJu4CZtZZK5Nm8cV39zNl5I4XT03y+BYkthWkLc0Xz
JEBYPrzWl+I6Z8hQmh+n8kSgxoOTOzJGNbJnM4oAjQtWylZd8iTxDqwOB1LG5sbUunax+nlFzpza
Gi/i/BZXH+PIouQTADmPr89j9ZF54FfFGimH7fZFVPPy2OPBiaX6skTam48dA8/DGFuQPs7iI8KE
YIq2VAYM5FiG9lRRnOm/mHplNmhNAp9TD90dZx8Ph4Yp7czoP4TlRAZtqRV2YnB9qc9Zlv2Lx8Q4
bO3wkNdTuY4ACWpDYsTQFe7ZlGyIWGsiazX0MEkQiqGNXtCQ5hV3L8pbM7UteTaQ/PES7M4+1BuE
cksp3ZS0EIoHydPBeiHbrBXr7NvB51IHUdxYisNPDJbmH+228tGR8U2OUGHQhBScDaNQGbUD52Pu
zFSEAsDsBVhEC3aZieL9HlhWWX4N7eDkUr2bdRQcAPqbALumttLUqFRoP30ukSw+022dZYadTg4c
rDaekPJqD+WExSQiMJlHV4nutyPB6zh3U8J/PmZvw48j0euBpo4bhDg0kKR0C/8qzxltBDtCeJM2
32x773BvZe7+TmfgflOZqLtGyir8qJCSBhMVoFOm+oynBBl+DC8BmOQ+kGRX12wgMqaQcCkIBbGA
5MAoVBwlbC531EJIFTZnC4Dv4pUAeOn/vmGqCyYcUjWird4TyIS9gRJgbiTlie4TiVuW6e7QlhAx
cIXjpw3etI4FIVI4RMHeVtDlPEhYZ+hmprk2ZYV0JY5iCrULrkkIuyuWGWj9HVkQ9gWnuHMIB3TR
SASsb7pUT4opGeZX0ajXF+9Xj9XlR0ThJBwep0gIjHJqilrLyihyvmoDuyscVTWyLXZEHdGnjkBC
HPsjPDJ3YmC2Nd9/BtP+MN7BO7XpdrdR2aZaTIs5cSCGfzgZX6isBLU40yKPiRuwV2SGLonwdKuh
1mP88ML5fg9gk73hiHD0z8S0PRWpP2u9eVHQ7FPDdhOUwPec5P3i08IqXlg70mvdCrFxsUX1cbrN
2o4owi08Z3haMh/AtUV09Mn2wT+AsIxqPtzG1KkTuh0G9WD3lL8Wf8Y3xE9+KsBmrwNC0WMpZgQo
gE/Y9LUbyp9JlzfcBa9lKgQX+e+G7oo9BvwqaOlCWfXzp9hHCNJ/D0heRuy4+/VSOzZakowua4If
BIHKzw99Q9FAN4jN8AC1Ri1khem/Mk6fG0VjxvBF+rKemhoDjMDSW2lcUbNUxq2LxOIXWNse4R4W
A3XpDvQVFzhyZcTMpAJOqhAxVxeCFYZ6r+KEx62L1sHWEqdjMjtjfQp3XWXKwlk7O6Qp1AkDtf/a
XpgPFW3qFNmty1xIqM09TNfjUjrsL0EgA2tt/h9w+McdysM6VdFZEcrnWuOIoITBSETsLi3kuGnz
Qh3TpUf67TBNXzS+Z/o8psBljc4qWpNuK98BjVNDPgijiJhKxx0iN7Tg7d6g0c1+84FA+2TYzMmF
IrS57YWF02NIHY8KBTFRzhuKD3f2H4d7n1JoAfO8t97fBFJX1beD2v7VPXUVN/g5J5fTahJOlXaf
/FKJYbYsT/2IfaqJsFsrMta8znwNCNKImfkUQeUNClBLalee37UrT9Zww/mre+5yowLhMc4B6PTA
rhH3EBPP9ynCIgZ/UsMaXdQqnS8Kk8cLG1TbmWKu9cDR6I6FByueJutzOgFVQ9ZA6okjRg6GCTlE
XNZksxwq8dFIREq7B3KzZXnzQ6ABmuYOibULwp8RjSzirm2oZACcCR00pB8Om87u0+lw1IE26Zwd
UsojhKsKq28ynkGKEwu58xCnUh3huo4RHC5Zoyq5R/VVDMWXOc/HI0VrF6BQyF6ejxyulFiQWG2H
dut05BSbAMOjyoc5EJnIwtxdSH+N/ErSDWNaG6xAhksJ3Fy6JWgpgtmgl5NI1yW+NueqwRC0uaO+
j0IGEldq90duQjQfyD0YlrD4ooOVAAjsbnvQkjXaXWnlHGXH5rr/jbnJFpPQiDyBp5bU8m7UXCpf
v7ILx/xsyiJbo7+MWzM5QI+8qYanmPzLVFiqvKwaLKxRIAMb1mSJhw8UUFF06SrCtTqjH3iYP0Xk
7rWfRM/QHJeN9DodsXfZF5DbLQj9nTQxlBsULicdHR7unF7EamA+w2/ibQaIqfmIgCOk8gQDADHr
bw7daDB2LUxAVFiF/JzyJeVajlv8OeBHaMU8Y/P/QrM8U05u8MCA5YCAmkazvlSdEGsoDfAh5V19
FOpgtHATGZu4udK7rNbgIfQ+HxB4IeL04qQ4zg2s49HUHxNV3Tt7iCytnfHUAFf26agY/cAzXAxf
NbtLwqMtBwYxAt2JpBNm17aj1LYw2xTCGoXSmNphXFq2hOUZ1sG9KxpPFKXByQygoBTLPYvMO1Mv
3GPiTmp28gp7TJC2+4+IFL5DBTePvkcm3YHdpvSyKtaq6e0zDUTWZ8BATWCd18ydf+HK2YowzoQ9
2/rcEqkvYyH+P74J5vbEjaTiuN+15OSF2da0tSqmiTWEUHDJ1XPRQhYMRAWUWXH+4STukJKcuC8U
4nU3ordUwTSGGYvGIrBHKX+fVA26W/dI+Hitc9j2uio9L5lXBcXNL5J42AJKw8HYfBaHZOQeHOE5
WRE5EBKUaieLG7TMWZkE8uyt+CTEk7J0e3h2gbIlZZtBVa8PYq3Vm7rO6c6Zj48PIVkJrplNmVDy
xdBCMnZJf7PN1p0OYv58L+Aq20N0TtADk668sm3nEKBuAyWQEZMX/8938dWKkUGvlHI4epM1/P4e
6AB/BQ0EST5GBy/sOYawKHaXHzdF4+w+DrEtT/0EUGFSXbd1IReTI2egEfgm+uqmbFvh0xlj1mGy
3oAKLu5tfazZQ6CUnOrmtcn+iGvsuck274evSQ0JQZfFank6PTB20lckwNB383f6JMkZ2nkPeXrb
rsf+hCvRzyWz2TXYFWJq3ZDVa+VZgAgANbaU9ilWoYD2ZKdk/Ma+pIxC0mI76zfGGTuWOyAxEUF2
UiPN4hHDCWUIPLYgXHzBCK+9BW+foW2Lle1bv0GxUDwv1Vnl0ymWy0XxJb5hP4m8I7KCzcWxGVQZ
tU72blCVa7VKFgcHVfTP/Y9fzn58H0oDfAdR9k9rOot+XeOMcTk4ujFlK9+Pe07EJixnEDCtauqp
Jg3E0NU5RynWEL6xyU+XRs4Y6z74e4yU+DR9oK+B30kVOMlJYbCte5EXQh6oDY3Rm8bNIfQsUpFK
DIwjHqTdgR5qJ+7IqcH74oJ0kJ/dh+xKjVkAQSdhamSGjZXEaR9dISyinjNlwdr7QJSsSoN8Y2e0
39H838NIAfR221mkwidqCUFrPz08gouTRfLQaNDakWH/MUOUc2zH9dTitCakgvLlGHoREabHsPv8
1a0RU2G6qKrimHsQzGqf4PbCX4HdNiMIcQ4WYp/CwIKLeKOV+LPLHO1ScVEAxJP+ncFuRfrWAuhE
wCw8Yfie4wIMsx8u9aKNvgdmOhwmnZ+pGSYHIun05wSbNjTP8yFkTIB5NKOeWZreeIPvbsYb4KLR
2GbrX+lODiQ2Nao/l9Uw//KhFXUQTgQBGFR38F9pH0Ea1B1uNmaAxl25EA861tywCqK5z/Yt8GnP
u1O+uuNmuLaDpP9YAezol6cErEqiPc5XstErYD2ue8X2DZ3dz0+A8JK50BQeguQ2WwjbAUwW7bNa
ZFiV6IuV9y9Z3qs7uh6qXm0z2RMl5BpFEhyW70YF0H0iHIPFuPpzY6kH03HUMzHSSB4BH7LTQD6e
TscfVKb/Q+6g0kNVMgUp96IynV6wUuMF69zLdXYYIvwKXBs5WPFOVeSahpGIoeUNDIPAxsW5WQs0
Di9CySRxLCrRR0Ko44ACxUZOf2NMaWBt7pXZOVm+nrdr3Nh1im0qcySekMrh2ego7JTMYerBTEns
UCdS40/5R3Dh2WHrkJ+7jGlscdjZJUw9e7UrcNQ1tgNH+KzUPz20tic/YcTQYUbUHKjn5m96Z8E0
/IDiwVbxHvMapHg7mIGO4R/flKLZ11DNCGn5/+5MdRAOnemYZYhjrAgUBFTMYoI/hqdGsbYeI+qU
C0d1bg+HIFQZt2wn77J9cBN7seLDFFCxdN1lIz5YB8o84Y47W8ekChuukdP2+kS5mZAK6fGPrHdM
OsepJiBS4gwohptjoiPcxO3jQagw53p8iZIs4+14C04FyiWqagm6uWCHU5kD07OhjMPP5ov3qe5B
pDD3ChhHF1ylBjeLYRgfBtlDbk8wP9vVXhWAvTNzrclpaSdHGHDSeNWwr4um6yf8B7UFWG0Cb+wW
Lbsnvz5j1DjrWTxHIXcPXrGLYtB8Nt2sE9ANEgsIFPD001a3UbwB3JJZVJBSViAeAVMoPYNFfcha
ebl7gtUsyHR8EyJ/v2KDm+QchYHilqJDGNaSCA0D5dSLTQhiV0YHF6LhWy5RZLI38rWNDRuk4gyA
sChexSW/b9Aj3NApC/zCC3tmYdQJBBdTIW/IJBFWxRLlKhBLeaZtQ5WowgqFllRowGjHyctVY3Io
B7wO90+orzYlG3iTxTCn3adWMfDd+1iJo2slhR0iYwYuz/sR5ulK+KgsfTVtp6jmzW0ULqhMkrGD
ZYsJaIQAQRYkdwBuXbHEJbh6DrhDtdz5FPMxiyJAyRC+RuKsneTJlmHlH76ENFfEjkpZ6Qj9z9Aj
vcWkI2s5IK1+D9vAbPZ3CjCUvAUGj1g2p5SdtAmbCUzKHy4Ns+7O3lJ4yr7rbYscaxm4if3uhzw7
F8DD/4Pxr5mRrj1njeUHRBpMfwhQcAWfUhsSmbZX036A5aCppywrNiyUWcJt03FM8fuvNX+hjhBo
bi3ScFbjHFyGS9ITTIQBwu2PQv2Vw4pmvx93zdU+VbASodrBlgmQMMpr1LUp+RFSIqxPYMUMwhF4
pqPKxSIZxx9wUooJr3inFW8BTAGdvRkHOja4UZwG4XGYoLChITClvPXrToDktpfL6+77dDyuEk5M
kcSfwmqzEHApPLH0PeJvaJLcY8La1p4yOF7x6agZ8C24HzZ7HVeZMZzBl2GqKWsrFsC7G6MMpID2
tZzLINxArwFyPrytwmPxJuOayF9ckcBnAd5LLyvR1qfZMELqgEj+Cj4MZ+Bn65w6CSFuD68tDfNV
1vjwH3hfXwZzw0FxMBeogA6y0rpoOVbQEXdQga1Do2wBRVuAhvQ8h+9kN894OdBCtsBPwGYGpYTb
N3TeWIA38GnA3aRZbzqmEoWvRs4g70++Rvg3uyKrsVIugxXX3V3HgTbPkdDK802W5v8RfmfRkTFK
PJUoG/IZABQ63zsMMmcCWoKzl/jU+BbqMMdVkQ7TdoGe48WxhqTpOptBn6oOjuNQguZeDYppHlcQ
BsvSM+4M2QDvk8DixJwMeWMAjpisUxBJXTDQZGtLM1HIpMJVlZkQTr8uDvb3khgVZA6hs1hMAOE3
7c6IlZJO7JDDn6aVBnfhC6N5uNjMxfP89UEcqEYjpUYof+ZWEdQpqtSUGjT/kLbZM4tEWO9dDbVg
63cRhI0J/Q7uDfLzqU0vxAYfpbcYcV+dcV/n0uyVaWRZF/W5b805VoUdXhklcpNPjKFk/ke5M42A
lE7c2bgpTGd5NcaYGLxctr5Y/O0XZ8FJ/5MbVTAbJaZEycJpnQuAy1wwN5cyZtcSvGhYF+eU0YaS
2zH2zRR2ykqLvb1fZncqK8gt1mnzrIMRz3Ktv5E5RnG4jRQz3yWYmEPamB4N3A9fhqzdAxLmNvpR
rMfvkkg4KTvmqNLjw8h+ndmOcDqmz810NkhbjeGUkwKHo7NoudiBFd3FnXVrw7eY7tuKWvS0mp/a
y+VVMt0uk+Evf3ta26fhyeRUeVQHGStnrN/nDhhbGkH40CBjOJUqL/KxgjaX1iiOJ6qxl7sDf8F+
sDN8kWoHJJ+I/k1sNbF679J2qIeTWcX74WlHuG31Xb39WRHRjI7sxKHjozWzXAN5GcXGl8BFSAM3
h1hM9/0DZQ1CUiDPJNyY9r/Md5PxvSvHpypvGsDnAex9xiGViBqRPIDa5Lh+G1o0Eo9HCYRykoiB
jqFG1PDRu1tO57PDqG6Tly6oBij5UEbs++nB7dQOUgGSzOXpINtbQIzkK4wmhlK/85PztRfjr4u5
EsWhCGC2znyWypiDB1GVMMDYHMLsl79huF4sj8igNZp84fhoZ6p6ZSrxJVdVTii5tkHDf2320z19
Ilgm0bIQHjPuXHHPUgHQfCuurisg67O8fnnxlOzJ+W//86aPrz5gP6I+YpJno2L84V8QaZjMlsEB
qGqkjDPeNzPqKbB1DCZVgLaGhcpCqGjXJqynVYctjQtrKLIhgg3aYoz1XPNt03Edj+v/RFJL9pAw
I3bA7GN6CX4E6wcZME+JrYd7NB+XFRppfY3nN0KDdwIUuwp02geMsoCHGjVUG+sQpKP4EbazfpN1
oF0pVytX+R8ye0Op318ul+i5bHAL+7OnPxwxvOeCXSrJ2h8X9hC1CTZNsE5+thotogZ6HXqJQ3Ud
IxNr+Y0lX3iqX2YgnwgqNFT9ohLUl0C3JReqf0wFgFHOoOezZAijaaUVDUmO7OMUbzNabhZkcWCT
TeAwtuI5/ar96zH1XRwoQWEjzG8jd46kchw6F3y5/SkeC5//I7d6dP2wjtgR3F1UtlF4AVK/WSHE
Cj1xLYAnxrkO6EUpVib6GDO2WYda8NotcJaryGaUcTHauixvgdYQgHoo6pvGL6IWJMiSZT4pwNOb
fBXnpP1mc4EDUpxT4YEpPDbn68CHv6xN2wJL5xRmwJy1H2DRR4odhhsG2SPePkJYLd/9GaLwqu2N
aveI3dmyQwR222Sz2f3nmdny8FkJGXFn+03RY6UUinBidXGulqTVcIqUWGz0vbL4Ld3tT8H7cpYb
L8uz4yiOunfUjRkTFOsJ7IeS9fW6V8Cqnt59yCgmuNkYDlxzlWfFhNcWeIg+8S/SSnD8vjPBBbaQ
hGYNUzCT3AhTFyINaoxi8Kq2EXKt0VgAIgN5BLOKUJRfTf4LC9dmRS/KuJ+TQ3Bze/0ejli6N621
ewyRPAGyu4Lc4oynOHAbUey9yT5WtJ7sqg9wQX1iY49EtY9ydzpVdQ5o5mUjnIVrevhDF7FITh9H
cAbil/xDiX2aynt/UNNGakp+B36lP6a8+BRBxbq4UClldIwIrc06Bt53McWn/MA3dDrVwJOJjmYe
n2VGjjHWJ/cLimRqjmm5+qposk5Zgbm8r7kgkff2HocMySTnH823ISFfOL4LtjPgwXBSqLkaVhQH
9IR38yKx7a9p0jK8KRpMQjCDCbANBPv1lvR62nz8eFsawZ4ROvFNERnedwclWIJrAvVVRvnHTK8U
wue/rqaltl+gWMt9zEHns7Nk6dTl8ZeqTO4/uI/g2F1irctNenrxm5UbzrNreK9CfMEyyFIy1jHe
pb+rFFVZqZlI1v81hWJ+7xS3YkWYbjcEbgpMw3IG0BwZQh/dHVCS8JUmOBP8co25s+XXS77eDzrX
paM1hK8brU9i6wRV+NixTtvJOUrebnMB5DswE6tUZNxIqs1RNeyW8oktje6CVIq3/pq82BW5ik9w
CyQVUIWf6X1J/wXsKzMH3MPJqDYk09ll6bNKeOpiGtgt+hlzoS2MAEVlW2qFPLduTujGK81+m8ZO
F9+b6PGjuW2/Y6Y1Bt8nyO8RD1Qa2Sg5iYi1pBcqW0EQNAwHwlhij9Vzt6V0rDpQFduN4wd1elbx
l1oA+O7GVAM4lHGdoAJo3wX+mYF+681bR2+QFiXAyRkU8kTA8VWict7NRrYCel2Z1mLfqqWFVKsa
FsHqKAiZwCuYEfaiklPbyIZHRTxOpQSG3DOg7kKYGQtnhCyDQOijlbd6b4pRSWsdLYgsmLj5fUYh
biGPfPLg79wztGikM6SFAQ874sdbGP0SWnijZt8D81CyMqX8fs+ur/MFVdBLVpxfIIgKcXVxmBKB
YzRZZTiwBWMviABb01cNF3QathMYnfNFpiSqpI8iXWklgwReUn8EYRrgXW8/mSwPbbgi6wlVQ6Wv
mTI7VSPvvyW5hPN3+Mo/Dwjtts1w7BKGzbZzPfFQOBCJh57dF9ymiuf6RnQntK/S2w1SBUoqCgLG
/9HwtkI/th04/HCK5hWoqWbIk96XHPpVkwOtPs3nG9uATnGwBZQ5GdWnCf9erQ0iq3Npn2b08L9M
hT5thiSuFYe7Oki68eWSi8gQGkmjg32+FLYjh0E1MvhpR3Z6ZVQq7hJtkxdhECnBVTUqP1GvcQV3
JuO03t1Kxh0J1h8AipUw9srZpMPmMDBo7AClQK/pxV+fNL3ghR+tuzAHt9QYndq/HhC7Neupu8Cr
s4WMwNq8ZIbVz2ybzpwFW5I+OnDzY+Mew8cAdDsvK2nBNjcA4CcPOVtEzanubsnmyRPG0J7E/nW2
fA4x/rydx9YHsaTRqj1rlMeTNNSdVSgWyeUlUyIoAGHtOzdwmIOTcDAsoLLCG8gDX92C2Db0GNJ4
jtxoitQ4ejpmK7sJgzIdxYSYC9VIlzjVKjWqs2btlr0d//SSCEhLKVJKOzVrDN9TEH61mQzkh9yy
ifx9hdcgER1KaHpnpsf0tpgUMbBlovK4GOBNDT/oSYpw9Kpkbk0jsQ2nK8ft+8XUIpDhMHwk2WAC
7gdQzvrtUMqqHtl3b4sxS7aKrkPdtNZM32DxqXruHEN6Avp+aFQs+XgG/XhiXNu4+Y0nkoDoAgyJ
Pwn4A5tCGOEw2srV1SzfVYZTMcpomZqj44BrSnHLYEkj7ksnLm/9ZAYPIWCpg/ZhUZrMHO9WfaND
PEZUkKD9N35N3Kc2oz32FiSSusb3RQD+dTlbfcAejCR2P1mhrgSk/Kxc1oXomaMTYGBD6PBHA8x3
ZQqgtmroVRWZufTqvfqJpN0rLbp3UBTI3pJw/yVqw7g/pbx9eqzSGTe9oyC3yvMuiiMjm9BODk0a
GFNWK9fzsAOAcJvRVLBleP0XzY1kUnpx7BpcQT9ugSkLVhBVMbBor9V4+4ht0fQRdyLQ/Si3lkpr
OgNp90c6yz5n9z0K1L+dCRsLOori1Xsss0wjr6Zyd1KaW4/OlTdXzj0mzSsNk0QKLjy5Pxf5TE71
q+gZNCx8bv8nOchra7K77jSy70qRBULN65rWotCn4Y6s8u0qgTVQ5EF1yMw9gJaEXry2u8SYUUMt
YrbHAhP6v8VYV9NQosdtqDIiloTuoXnQfZ2Ji4Eh9tvzkX/w3u/ZAFXdJ7Me2pssxpHWm6vcP8w3
XnVtk1XYZnHjakqcgTJQ84jhWKl9BK2tAume/SgZpdClny7ln7TUGkBmkjHtEvdfiWCE+9Che5xx
MEg+En/nyfIcjOe459C8gn+lKCXvrYeMlF9AA+SmOVx/R/norRBv8LWCeKs8uivx8rhpbUlpwGFq
8jaSMlUU64l3lgxd7Z30HdOfSVq8B+GCDvxR53MRTFw5Po+K8O/iOWZ4jar9Eh+N1oH2UQYIwp18
jPRw+wX3y8bS3l1Z/uBnTYK/ctx6MbPrcGZZFOUmMXI7ewESt8ctP3mMkpIJz776muZT03t+bp/C
1UDjkObc+gVizg//9njSnAEZTLLU4JghmDmSN5Fb6lrOfEgMEqCe/FTjVJO1UedzWtS69x70R/EF
w2sGFPBYFwb04qzXa0NEazmvRI7PQPF/7WOYKswcKKbBRaI3a0w9bg/laZ9iOkTWFwNgEzOQPQ7P
s38zak6hmnjKX9Ffh1L3R6Q7blxn4jlbxN6ZD+is9ASljmeeDcWkJhKByikRjDRauWzPFeiWwsi1
DcMaI9H+aTmi8SJUJUtgFLwGCAr1vjRYNiL7T6zlEETKRj2hsv8LWK558lUoz4pLVs8GeuIbaV1u
Ibsv62jRz0LTwWZyh/kC96ltT2vZP2PyKD+k+edGyQ2aJRZqzvBpm8TqaGMEx+LgK2Odl9OV7k6J
hRIQI587o1LmzOnCjFA9zBuyG+kyqHY+n5q/xIZn9N3pkVPSLPqovNxMtgoi/SNcak0lKxwXOxma
v+KKKWiav7xEIZ5WRFtbeAvn+IuKNcHkK11M1zRBa7pq9XqzFXnsPiuKNIhaIdo2hVM5hREhGAD8
WzK2y1uOtJ1h1jQjtv/PDQCn+4PRklebPyoCRYRV+OrkmkTKpRc+zmVMfPy69wg+QqyNtFdAaa4R
R7rGqUa9yLH/2LGGL49LfTXKIYGlwBxEP7CEQtov1mgwdgcSaBwdQOtJsIRJx4v5qPlaU7KjhJXa
Rs6D+HQMeyZnlx9ZN4D3RwJd1bj1+ZqMyBnaVSLEciNHqY77bv7mmUgZJttN1Ij3MXBOfi19TwsY
ldat0DY0CvcrkPtS7i+BCom5OB8lF8xXmcDZZdgRDuu+XWFBPdYGnySWGTyKL795qsdRS0oSR2j8
0gbtyZIsYSECUIfONBOdHH3N1c+6BbIw35lYlff5SBhjJ9tGxGdGoFDJB8GgwhCIdoiTpdY/qjuI
ORsOixilTQyyNJGL3FAYWB/gQ8q+quMskbuDqaL+pJE0Gil6gt8Bjfb6t3IKbCGNgpoqsjgl8xDP
CWiENZIQhjOIf+QD+/2C6vJwww4LnzR7RbFJMIjTNQXoM2XvM1ZWGrXgeMKJzxQVdhzeKy/O9QpE
xcrxJoiB6oojgn+0hYvAUH59UwG5VB0+5Qu5vgMafcTHDMOibmVcO5sr/EeUubp5OooGksG3Gbuk
5t8Aoo+TA3exCbeBlLK1dCMFZOTe4O9GUyhGTQZR0FsuYQkjNqR0f4zDok7Cw/t/EBoK9WXVXLCw
UASHkW4EnM85MrlvFqWhZSrGlbkGcQMGh0etHI7jsATilsIPZ0IigsS03z++hse1VBPOln2dc+Tt
91nS8pSVWjHWAm4nyd1W71HzeSqFUzTcxnY7MV5xNu3ctb1hu1rr9MNS549GeEBJFH+tZkQbEohO
pPK6GWLBadN2gzLPwpM6wPAHAnQIQEG/peu6Ij2oXqJ6EtLukQjfSjmK969kJbZRC7rXhNhVZeHr
McrVLA9irPt72wzJTohN8wGlOVt2VfngbsXC3qLFkcEs2DKyZAupkCcAc0mKSL1oIajTwAhQbqYL
TF1Szn6BVdmuvoWg6IxGP6NBvjo2s7uJ4TGskbMyKBy79XRn0RgY7+FuwOk7NvbdXHrSudfC3vVg
mAAUiltIlLAeME1bM4p7foU83APnAReCAw4g0kFlBvjrZCXxtbFeQLuwYsHkDwLZ/RNm/S/8AAPB
NoIAA8qnR1VvKxLPxrAU+Y1e5nrU5aq4l+gVUTV5XtL7zcj9PBqXdkNeXLw57VZ0CZfvW87INssB
WCxO1CanXVXRUKHyePIJKBmC9AbMslxc6K6lQ4tp5/aCEIoaOMlTlLCyuUvVDJTj94JS2xHjg/fe
y/SRRlTLJ87k4Ar9j1N9rTxLvY5w3/Pp5Q3yPwdgwaTZVr08jHk9lQesgBBmg5T96mMOlSrnxCOy
A6czjiSUwuqR+P5Asq5CNpNoXRJzpNpOm4EuNb2DUmv5ugUlg8/oOj2xNQSOHCyDjwXZhDirzIih
eIwQ5l+QVbs/2k3zyPa3oVJwwLy0fydS8dz4uINXL9J0UAhXAhUCFaIICYbczcuzyGK8IM1HOzdQ
hBfyvjoQu2jVTgMe0G+cueq4R9ap0y0a8o9Gd/cQg/SVQXHYbx/98LGPzrKIC869QQPBYVHu3DmO
lfgvT/O6syUNRNqzP4WqH1j3worDvNTzrcZPnavaYkEscK1C1nTek27+6USo6dAe95uEtE8UjZQo
V09Nl+wSlAdq9P02YqKSj5PtGKmt2w+innm5u8y9wvZZq3glM3JVf2V9B1fLV5tFh2F/np6Ka/AL
sZTQfsRwEOJUzwaMuyipIJSFqmpjoMlCARSXkqNE9HnfhsVu99RfN0Ve5TXSDG3Upm13C3zuHeP/
qeCtwSoa1BAE0dS2B4qF/gLF2j00gXONeheK4FwNva/d9qnBaC3gtsvsMSngxDNvgmir2E8pS6HT
hQb/OE2UjXZqCpEqZg5dF5+BBt9ZMKbpJCkLO7/r4F5eOWPgdIDLgA4UaqD4vueI1HXGgIf7Xg0j
7aRI6Gus3Skz57W8fp+RE0Lbz3jsswrYKyHAa4r3hYQSz0NGupuCjUttd4CXKKchHe8pBOm/DBN1
25XpNVI3BOqA1fYwb9Dz2XucYKAQ6DkIVeCG1r9mulCLFpGzOWXlgC1zE7mU6toXT53HClNPM3XW
AMlA0AMLjsXAySdURLb5n/nV4/2FMydBCp7JolVIIqFxvT3t8RnWB8x6xz10hHJnn70E29MYbJLN
R8c7s6rKtmFvR0CtFLV2Rjt1hZpTnIav3GJPtWLl78Ixw/JSyvPWsgnsHYELkVmMg/EZghnip0bq
libIudhb48yVlBCQcf0vQ0Vn4cDQgPYDN0RpbRuWeY2yQaqzcfrHeidjcGrIx6d51j/YabIfqWMp
FYzcZT7vtyBUoVEp6qpnHue/9UXxFPC6q8YwbOtp9fo3vxJdWIAGEA6cuxEONck6KAEDCF/LT6XF
nQ3jVUtn0BZYt7bMNZM/Qig8TJECFJEix7CJcJdGL+BDicUR+hdQ8SUL3Gcjy7pGQLKsb9bVU5K7
bV+SkIbydiKDW0rmq2S397vehGmGnmupnkUjxytZWSn5NjSvIxhfRs83eLKvOXAvOtVGaUkDMBLg
gmU8In0uVFDJIh40ecizgeEurFfDABaKgzne+YQMczRZF4xQTOKEIM4/+h42A8ft1bFhcV/IX7n6
jq5zwy8UaLler/MVqBVYi6XsNXea0YghlIEEMgYhNLvKX/g5mbRxPadiqj7XpTk4VpObbhwJzudA
8xpqpm6vgBiEBa2q2zxQdeImY37LBHTm4xz+WM4q0LBM/m0POMWmMHk6a5i+kbVLpxWUtLiCa+QL
iXOhgGDv2u1+hRbjopF9McVzBalQF/ZTftoc7Mg6LpGc4dCPAU/vrFo48VChr7SboUg+pbWhR9bS
PN3cUI9lzNbWyeH4q4PgsmYvgkB6c06z/mQ+bZ9WKXg0GxRuNlLpi99wSrGR6FkDiAbIgTGDF0KV
HDnHU6yas2uKzG6fn3w9pVgXWFTg6C7MC7+z/geXK8O5OAVaS/NVDXNtMbgXPQBkxCHZbdI/O+Cl
Y/er0+l+9Y1U5tD/eybZ2cDyXeVLnjjx9jWfsyR3xZ+IGePEHeukcbdoN47qdM7V+rBOp/0Pprzi
soV6Y5AwVnz+K4yT7/1OJ/mWh6/twmiVLBH50YOPNucvLJQbQTSO58OQpifJtqY0JYrxDH8OZq7W
NPa/g+KlpORYnMMwjaaqFapBWH/c0eMKg2ACt/3J5Kawb6DftvPh8uU1AKeohjjT3bouyEq8rW6D
HhhKDQgcWJI7FW8qtAFpUG8VtGcTnUs3xFbiP/Rr4dqoXfpUIoYW5uSO6v10H1w5FOS3s1cy8UpZ
fRip5NHPUX+DVt4jDMqf22HAsqEyQ8d0m3ePH4QfluKlbDOfcf+GF9haxK6S4LHKQ4/XXWgvqgxU
l02KgXqQo+/bibVuz+n6P1dpQo/nXFFzV2QpeAtai10aCVE6sgyKLrIbuc6gI7DiyAW6YQGdVthl
DEJ3d0G2FJcpoprawEqx7+UxmTtmuw6WPYM+O0wrqnPITehvmShKjjxrzj50HRIozROEK13Y3Bb+
uivLl0pWBTUm4k0NszzCIo6ASZqnXMsK7dBqLgKAAkkrsX/X/Oauv39Z71Ly9Itmrvi4/7bWlZmR
4CTaGwyka9bcpQLOR8mU2HP+uoQ30uGtdsn5Fi+eol8N9OGRUVvilMytuxOqIVek8OrvG2wxWdtb
RjVsnhlWOGOA/vW4Gw0LsX8Vzyw2c12WqW/8ppAvXec7SXD6DRvpKoWmlis3w36l0WuZKMqJp3y/
QcqM9KeXQqQfJHYWvaCsQFwU/Si4DZHAwc9uM0gx5VfJUTJQmh/uZQucAic9cnmEWUd0xMJ4NtfE
PAl0zzk7k4rAqVZrZ7pFKwzmX69pFrNyk8GiaBay+yjTGNSvV/ca6TRpTt1gabcj5rEFdGEa96He
zA7uuuiI9ZIWQ42DPvYU6/pywVZMLL1RW5VhKbLvRC6+mreqjRfZ21pFWVJbgsi60qYAWlNEQxad
YgbktxnWxYuotDFekoUsx36TH2sRFxTnq04jAKro3J8LHWu7OKfyjz2vnE+cYTnmoRr1tVUpmIaq
DoYQ2r+83ekKUHbVuAyzRfrw36l56T+HKqVVL94kbL+WV0MP9S3W+lEuGxZRk3bLS/qSR5H2yHTg
GB5bu6+owENVm+H1ba5FSRMGX8ZFN8i9P3OuE7CE51Ou3gRKjxUCfyWXsJ/yEpRP+e/PGiZV4woJ
SL+9PiRsSE2Jyhyl67/nvz4Oxk+EnMgWANUa4zcMhBMBGXMld9pq3aBiNWsCIB5e0vBnlVNxueHN
Ws43CJnqvTjClGd2dOjQhJvlRTEiRv7wal4iZWeD7aEz0WaBzLtNIBydLn0n1b/xlIaXAtMB/lBl
yxvR/HmibbSja3ZB386dhGY+OUykXRqFj6gsRqtBrLnk2mKB8ORS1tcRQfByPAbBhEuz1hMyUCU+
lK+mERaMrX0N1p2k6B1qNZPNrvWjB5u3NZ+Vt0TaFY4Q/3QpSLb+/99fMvuRWXVmdlOtI4q/KtIW
kE+9qT06KOvRASKzFn6zIh6seMjiOmaE7OEw2EZu14WUOCULJzjRrGmr+FNgvaFHP+SdXUFlOK+n
CVEw7vmRC1gfT34T1U8OyRsGbcQyxE5xd2aeDIuWkSzkjML8/CXl88MeAuLvDY823RslH6FkgoR+
j8tfVjUq/k6jUUaXzTcarJdCCVVZ9JcyxwhgSV7XSEBIjeETNd9fZqP3Hg7WSOELglRARCV5G+rQ
/xner+mDAgS+LuwxOXt/RT/nUt5g8hBDnowdEggaTESYUT5mI2T8+0+aHu1DGMYXj6D6DpDSMiVn
ilW3KcpXtCnS7GRWo5nYsin9nz9W42nkV9deUL9+VC7IlbWFHp01BFPnCAI4Y1AAgCiSlvFWgwch
BahnM2hYmiApMLDZZuC1O9sHMQICyNdLHwGPezY3tV+a7RBzKWmtcXb/tutCL4dd7HLYzTeoUz17
lf6OKHUkPvuD/rZpGsjqImNaaR0x9n27qqny4VCFQ0guzRmhVufjUjhlXBO1eCLIbjzrLVNtb/z2
3DqO4uq9LreHYjBfsiob/2MKXwpUv5mETUsmZdKHU2UM3hl1u9UMHuur9rLWirp1P7Gu6hEXhpLg
F9QoAi7y/Q/dJU8kJ4AhH6NMAO3EYDS6Jxdgrh1NK/tjiB4HID1+hauvI1dCLYWcfwMOSwNNkOwi
e/t6K3OaSok90nVcbDl0hTmAAj9uDBfXtuYPpZPTfPXwGFknhUg02Hx3ncpybJ2v+MiQocZMzb9p
E9D+mG2ZuNdokq7KgPLKT6wpfdV/Y6XNfwrWLMF06K9W1e1L6DA+edTsD/vwkllN2n/i5RGDm0MQ
vFKhzlNucNv4usa5dhnqsjeV49XIgQbMEC6tmnL9EFOQuy8iQ/E63jiOILKrMj8oFvBzBsle9KqA
7jB9XghFouPbWHFSqjyatErDiat54E2fiYZMxu/jv7os92hyP4M/Tw+ihvIZA53UvMoH2bUldUyq
ve155eGvTRFVNaToGja/iWSccFlfu+ciV+xN2e7Ox/K2YrBG6vAJrjVCvbxGAioqUKDlky2QoucU
XNsXKsA5ZFhviEsCoyYhWC6OQoGUOPwzTxe1C1tDATlcnMIF3H0kaEbuu3MTkHoHuOXQEyLcv4cA
otG/wk0NOTH4Jw+26wZCiWwxNvEbWDfqlc7d97JIk0BsAzvS6HaBK9togAdfr31jdkPB5gwJW2di
yMpJiWlfXLND7o+Iysm59DqBPMbL/DvU1DheXvZZK2FzABD1VyvWzz+4i5euTx7GradsnUCdjZht
/4TgqTts01Ja32ElFlCXorveWDug71MJXhHDOT6VSmnC0mHVylC53ydbnj0GakgnK7U6QheBP0Po
8w3blltqgF1OFkpVKXVlVWoIAiIQz5YO+0QQBMWs6hghG68I7L9EA+kC78s3nkVSjb+xrbepZOif
aipGc0sEFidNZyOKyLxuDYGLlfjMtqoA+WOlTb0Sy24xjc96o3eXmQU3Y7aHKhKVNNRp+rOaNsfp
ZjHYiNiDaEAFm+BWs7V6JcE3WOYUMJrUEJhCaOa8WJv1VeLvf8hwMGD/3FkqY7zgEbRDcweJS23Q
VtNG+2u540JRZB4b+Y82G6TFuCWE1SiBQIY1oa1hCL/hq5eLPundt0eQuvP0aBuUwtT9v6krgOXD
x2zKmL4Xl+Uv3LIsnWKNmsGNFmTD+muCX94YeEwlJD95n86SL53oz9hqA7W8yQsXN/gPespuZfZt
hcN0mvp/j+uTODHCJses7pOw7iLn6wKjADGU83/BKdjivydSwSWV2QSVNWLmj34y+0ZeMF+Ug6lQ
40hRn0V4I/F/ipFPpKJ2LLzPwAdL7pUo4U487uOsVgrhwZskVcXbzFcZqbJ9PwKoWaQfBK6EYcct
2LrD8icwbggXsYhwv1uYQT3pJPs8fm5qutCjswuLrbm4Y25dM1HtVlu/afOLQu/ri4Vp6tYez4cq
02r9RyevohM/5lNRfsJuabLI4SfRKLwFLfsSQfMXscWV2VwYvQLILwb/44esNUUVm6o0o0m1XUiI
GzwYI9ayZ4iYzVxiv6VLVWV0NLMlrvq2Mu1iVMyloKltqwffgwNxQjfw6sp/9EY4RJ5hjOOOmk3s
vxJSbpLjePcI+dZ+xvbwLEl6c6iIfAGZ08a99JtVBkX9o3HGpp54qsC7L5CKWShK7XL4sgiN7xde
3QiV+x+ZJRctnPKeTiaCaUJPxawg2StyPqZ4Long7S9z+BK3YgzreYGa+h2p90BMKFnJITgW8I04
C6BdNM0GWBzWwGRjPA22fjsnZ7HZVpXHJ6FES/tFMTVTpUFQcNivirRi4TP8clZ/yVVPS7dPfuUG
VaNlrwNibZMpIl037b785uglQ/Q0ZhkW+4MggRCNEtEQlTczD6p3wt1iPd8cD6MZyOpnIZl6uo9/
r8UO542U9BjeNcLuXuiMvh1XrluJ0h9lC4jsDZpraWYd7/edvbxDSwrM3/FuaVpRZgWoGQXamOW6
EnACKdeS+wvhrdGJe6XJN86iXzjdiyfvoijq/iCkMosjHXCaWHQnNXm9bya+IoE+Qs34hiVFS/rk
0B0Q64I36HP299y9Gn0FTXp0kgfUfKCv8TSwuszyjgOcOuvwDkcEjL0FMsxJmery1EdhVrFug5GJ
xbLKMvpbcbr5TA0HsCAid3uUJvYD5/H0ILMFqv2uQwRQ099b0eoX1T9Iw74kR5xrnKP3y9SlnMXo
V0ofUAu64UOC1vW6i/l9rXmYJplBQGfMu8EGqlXywZSdwFVzf2neGmEvvP4fDxfqNDQ3x6FTBvBQ
JhnguA4kGYgGihEQX2MkWnYYfy2Be+jScYUt5usVRPA/mtxmIhCINDfukQZQILJHpVaJYohSQj6M
Gc4LWH2KSnOkWfpqAxF9ij0RHke7n9uVravIwMaAtdtGoMygH1qiGOTcWnLol1HDcN74apij9YFf
1m8zpKO5nlyuMqA1g1AxLuSZfKcDWiUPaQ0bCb/b6BfwDgBA2Y4xigXTgOxEW6juCWpab1kPbWZL
+F+ZOlNcXT3lcRLc4P93iy5ls4kxoLD1l8d46JKR82cbag4lcEb9OhlXiKetx7OA5tuW/GkJ5Qs9
/FOXNHDIOF31klIasY2uCRaF2T3rPeT1vsgLCBcj6zvQOEnFWpu4q83qbMzTOMxA9s+Su/qeMnhK
xxVBv3UzNgjJrlQv6vLRUjsKjEc7N7uMuOPzMd66m7TehckTHOQfDk6HUJl9Ucpem4S+9imDlEkB
+codXmCINLlH+kTyc1YhsPMjifFAuVGcu+ilACPb9XPVlxYCP82qbvPmHeEw+oNq8vO1Vq+Ev4+a
B012KGC+TYtjeOv2LN6ZgfXEcsEwNu1L3h0KF1/Ku8XS4yhOh+yVTqNww/eXxNdZOebTvWvOWs/s
SBxRPPNccJ8risbCunSg9uT1M/A8z3FXaUyY2lBXwLDaNFdYXrbdSbzSJzw1L9v9T8wXgcGRVfKN
IKU2thx/QIZroDDhok9DB0Z+nWRLHMnWquatiX1Etn/7jnEhtiXQhvYcaVo4bnbuU9Y8Wr+gzgwh
gIpkPHe2Rre/hTsNujlYK4ul7Gbjpx0iVb7S8nBjsEyPljb8xQG49xJaTH3iOLc2UvlwjmxnzaWN
/AuvM0lAr/zlb36PB2IcGjacFWZnXmLYcIR1fM70DyT288V57z223NLVAVxnWd5IrazyG2AEDzFf
fYUY+s63lbHiVnTnybkwcQAYQe1V9ryLuGDIUltm+mEHqEQzgZfYsEej6D1j8ykEJDQ1SYaHxvco
uWBkQHi3tz9/nUxnplz7eQJui+TnSgoZN38/TmPmaxlU9BlQPy448vTURKWY0WvE5v8fJW8lCURT
V56yJHkEmMAvxtkzEYZVOOTtxUU7G8QTLhxkQE8W+5XNkXeFYfZWLuloQoSeMydceT7001aqbij1
fBORRfM1ruT4o81NZ8t1PQEb1tUTJshAkDvqaFsvNMBD4Qsxxkvk6umpsvHua77xBNw1/rMjVBwD
7frLhOBXFH+7GkiL6+n0oHiEq72+d/ADrw3efc5WQMimIG5ecFp3Ml8KrO9/I91LYwRzkyLCz9R8
iuP9HTCUv8EzsU4EIkFhFkzOCxtYvA2HkMDmx3h9xWSntNtlrVyDO44uOFplLm/kWNADxlGguVkE
sSFNl4LzeB16kwJVxwRayPORpfEsOUr7F0P54FHRSc7WLqgvI1lwmLveEYPvvsShz71aHgSRWToq
U8sFjqMgtnzDsc5k62iNI5ovMGZakhj/RcR6KzwrSr03n+KLIFj3dXCG+l0/0ML2S4O2vltKRohk
m9UGle2UwTHxX4Q+To/hSaX8QL/iUzZQ6kkU5hF+XdTxxhvF9JXqNianPHdT7ksFqxG9U2ltXP5X
4asDIVShFDoZJjrp5qYXWM+VWlABRKGFQq8McQsPO280cbSzWpUNKMUv18FxWObZwZwTBwDGDKQr
sex+hLSAwFevz2lFii8SWUxRsFpBhEiEP9ixhSeWZXAUlNWew+hhYzQ4wwlzXDi6gxODO5wDA3Th
ylCP2YcG1gdE/htTdgB1O4pH0BaHu0XZYkD9PBN9VfVNNY4o+yKTLXYRzSXzgAdL9qzyuJ7xuLPP
lInQLAYVDtq6UG+C/5klOyJVZLMrY7PUkPjSA6qJUvM8l9qNl/hl/7War7acKv+TpV0hyAygjPBv
/psdbqVQyqr4Jse3byafchiK5VROTJv9Bl33v8aeRjJemtfhkAGYqEHS5CbTI2oRZLtFb/2nz/8O
kruBq0y8h8rOWIXf6TdVjAhGtmmr544+EdiuIr/SSIr9mX10X1coyF5ECxPTFXX940HO4e7wLTIo
g3L739o5FjARgT08UWwQ6NTt0hRFIO0RLRFpKkcXiIxXQePLk/R3r8bJOzEcmp25DxP8O61wju5K
lQaHT11rUJMJ2ukdghHiNhqnG1HKX+dIpwEfJEeX5OCPDmWG7s3hjbB5AG3LnT0kgQsWYWAuxjsE
nqLt1JeIAhVatOQyzadd+ZtN46sGkotS8FgSxhK6E+90vCAucO7SqP/6l5i8IZEEO5z2bZlErtYQ
Yn4QPvbtcqpOJBlwFlA2agHjHFK8r9m4AKl9Htayw0zH3giAeqo5Ev3ZxIGcnlleYMciJ+uUKIKW
0x6VHd0jndytJbmElzZjQ82/RWM6J00IFfyqZxCaG/eldlwyO2gkwOHa7I6EDTP3fMqc66FtF+u0
4Jda8Gmw6x7Ihq7DpYqdrZ1L8QKDtI/kKa9h9VZ3B3/kVSgFlBDd8j2XTPt8/kMvjxRV2uYnBs+3
55LcV1Kx35U9GEiOJ3Pgt1yKmGbNhg2Sea1aBr5+03fqXoW80ZkAVjQoczfIattfbIhMQFJ9OlrM
jYqdrKPcxBuPxRyqWmghinWK9UyeRG+989j9gfjHXdLIzxkV0FbMpu1IBsuibVmLr253EZfMb4yK
s+qgnLdB20rO8LHbCAd20KZ3qRUNPd/I+8Ccd4wJbt3GE8I1PIJNdW6TuDxBqRLaeEzVywMO1bxQ
r6pykOVCUvF9ufoQ4/69th+ZYfVvB3D6K37ViFydzdELy1CCxSpbyDYIEoOkRDevNkcWFRpdAiz7
UTmFb61nrUaZSRm7MtLAUa7ypZ4teepVv/idqjsz08160AjQGcsE1Eq0/TWzzujUHBFDrh/Qk0N/
Y9nEp7vR14EiW5K8Gol+Dh0H9WQVUZN6SN7Kn7upOOUn7R8TzYsrYLKNfaD6YQscNVEiWU5UKaoc
a9qMiW4CFujx4P4h2OniPTOG8A5UhDAOe7bIzAXWy8qiDBLCNQdpcFpk8hLfwuT4bFIfg9ZLfW2o
BqJsaTMO3U8teIbKGi5FhaGirMNFi95FSbFETwXmoXlm8ZDNLv2WSiNUuL5wo8ISiSLSxkhYXKyN
TIHUfqiePxlgGg/HAuJTxPRXJgYhTLlO0NuhjOpz6SR/xZ5PE1kHEK8nC62gk3/dCTJb1LWMMtfF
ddPBPDUAMGG34GFBE1xM+fB6QEoIl2l+ZzmoQ3foha1NNxynHm2PA1C/QFtuFU4j9a64N2rE9iiq
YJi4VNO4fBRwR9wOwNhfIh4qzXvTEWq8ZaYFJGTVup8lX0hxiFpcX/aodnEEKo0jNLLZkKKrl0Th
8qiDbiRsgFPN/J6YvDHy51dt9q62+TMgSfOqrBNM2SPPFtJq9DkJOaBxsr7MVf9/RImiKK5Gl0dB
if3+JlBH2inrirlV3dLMy1NDjFSvsNeTNIdd9ZtotMuDE6am1z+e3QLk8wLMnhZ4Q9+OCxwZwDPF
QxIgjhQtY0r82od0AeyziCnMoeQHJnm/gLOtk4OP7x4vBM3PCdrPWVpvu/z9fTXQBqMcoZssJ4yd
miY52P4mm/NXhFUwL+bTXa4+7eNqxf5io/wpm2L+pflxUbQ2PRLLSCxcjFdK5uu/oFSCC/u2+ZOd
mRa5a5/GkWqeCi5J1A2FxtcpZS+1clMsG/3lGANzCvACEfdZUedLuz/V5FgHLECtut077bB/di4g
88Ng073kpTsxRyPbyZ2r1uaaHOEOX+awbUloIy+JN2q8RcdiKythfoPIB9XF3hAw1F/ujWXUt51k
AdjJSIOPbhcOXooYRvuywcBHbMQ3funaEFPYYGSEIA9YMZTUTCNuPzTzF+eqDqUCEbCniySa/r5E
Y0Q9Iprc45l6Y210FMFI1N6zh86vMzesZwMcS3Cuw8cO6z/hZWU6YpWlMV4E2bvx3liU5RK69V5Y
wvSxHsCIn4trMEQhxS8JaghacSn+onAFz0dJCG31utftA54+qMOgQXVb1vS9SpBXpXEqDBdaB3KO
iByJ9hUPppXSMiMoZXgTLJd9Jm+S0wY+nWUFh4hvraItwiW0Dl8wTL89327ZMC7qY07KJBuZjozw
007EM5mZlI6JufjmaoUXLZic5gB/s10l7ty1cS5zYhJGyya/KDSTeAwUXGUIof6ecrmMIAuRt+sq
n0NSw+rPg9EziS/O+mmECZp0wdaprO8p7+oJOyrdSSAM+7B1l9UGBhUXcb7XuXn9OKztNC6Y3z89
D2tYFsWExBEbkEba9rRuA4T8n/baCz9BW6nj+1MlVSQoFzW11FIkB0wIEh07FfGKpdEOR6oh7ZU6
U56dOGNMkH7OoB4ZVuYkgQMGAME3Arp4f1mrM4m88/8moB7LT7D5ZGB/B94h0XZsrqci4fLmuDL6
hkO8PRlmY5GX4HDRGHWFIcBScvA6CgojLs1LM4DprNmEMF/mSVyYhlj/LnF0dj1dmiq6hSxT+2ru
Ek4Nndlty+uq0gK37oBGmQVjJn1ukeLgkRMnwMvcGT+60zUVZTMtRRnqsp1m/OKPG8OOW5/4nubf
Xgblce3hn/ojA4iwYjHrJflAy+5rRnfSMQN6DND3YNVOKP2TPMqUwjoAFqb4iWwVi0+hjiQ8i8D/
DT09wQHCuWmQhHZyWzYklmX7EqCAWCJSnL1Yp57rlE6aicRVmY2IC73avWt8vs4qaVrSGqcS9TEz
NNrpVThyjE81oGTj0getni/LyOo9apGO/vfC1Y9iOq2PLKDA1G/A4LMw+Wmxpn/ie9RRUa85wiBf
2rggN0vP8dX9uUFEvsSPdBTABL3zUTTark6OyWvwaOrdC4CLmvXI4lNj7yQRBXAMjSAXBfrOHhLz
3ScS/ZiZZX46Zj27o8uwr977pHS9Y+y7T5Ae9XhOFuKye9qwSkIpXfXb2wQHAigtHiGxoSomVWw6
2vx/heiVZyUtB2aVUMLUnII4cyUbJc6yRiDXEi4hVBhL4vI/Z6rvkmv08/Fj4S6mEW+/C28PvKTe
Bv6FajT64TfiGOkhBfWJkEJ3WpQ1X8h8uZDbJx83F4Wj87Nvvd/46ixKCHifxBgrNViDn2k/7hE1
RaPlt2o7xRlRzZ5+39u2zvUrn7bBO9syNvAqx6xMqLEJGzMciC/WWJMI7QnZ1uCDa41aH8vetgyd
fv+R+X8hgjYUdqCbGgpAx3eIMQxjk7QXz9wCQV3PHFpgPmPhnCwZZdMa4KhIlBMa45hZ8W13sUEZ
UkEPb+ZAD2sKwLQ4k0jRR9b8MGquKDKutxfwy84xKn1qn2Rv4a5ojFbih1QPle2cFECJWiF0Q36k
zm2XkRRIT68z3rXWtIAM+75PDbuC/eLgDxY5bFnAC8HpL/4c5SdrbA4+N9OC0FTAa3043jPwg0gk
uWuW7s6S/tWJIs6kmfLjYo86VuJAm2UbCXzFvmow8eyaQab2sNEsLvyie76XjLX7lRx6dwnK6+90
oayadWQsjOo4bd31QGLk0UQpBPaP+43XTtvpJ53ocgq1qId/bK7Hc7thOO7hm35yeslbKTKOYAjy
SEjAWsaecyRRKJklTOY2Fgku4OldYSHX8vAVcDNR9BSXQuEyMa/yXn5ttiYr+90Cn6Uh4MQS9KyW
mAhQQ6a7H4NkYV5FI7nVlDk2/RXprKiHBGY/Ff/bWUErsOlcqap0EgQkP35lnYrCjwPs+ZE59nHc
BauoxMuTbr1tZE/lnZeRFTKeBn4YTqWVlZ+lkQs74kXtDYdpBR/erDRFkBG51EctOI02jSxAaZ3e
2F/lkw1Ex2BuRN/NUaZ4CYjr8n0EqxlfRq91QLNX+P9XzkFRP56dHJdaDZ3n2TQQDMF/cRKJ4GbA
4T7MjoMsDQzCRQ/PoWYFZfIudmiNbBIsuSU5aPSexpAHq/a40Pg4QHl8y+SH4FOo2j1QhityqDCl
FqiXGz+ohOUZaLa3o/Re9xXPjDK1M6ucViIaUlSNrwN6lc3pl1uNyylW+CtttBvtm+EZmwz4KTPF
Q2t34EvFWPbVOgg5idHFF78WCfsbBuhFniy2/UtPkBoteSVlwYnm+1DRRFRQFfUpIIJlPclFaomV
y8V4ZRb8GFTaMn0ubQ1l9Lj34dIGeIN9icnGSovLXV+I+iqrlyGZ+EgNfcBYRDDiRJOGhJ4/AkQt
/QA0cMH+6rkAhKjYkH8TjIk/q2u1StrQQKBlBVM8J0/CUuP0R4zZn7fMjjgrIz7A2rRKMpVQA+Yh
bt0DFauf4bRPu2rLcSCCIc8sddsiZddK68CCgjkbYMPLQJfS/l3m8b+kTekFzUT4SDv3/ZydWd+8
zYz0runkzGHD1mh3MK+n8qCRnWBCC/q3SxM5az67sssSO0AmF7bRIpcjMEil41nNpY/9Xov7Q/Dc
ITMsssyokXZeEvglOYZ2ynmHRGIWniG83QpRXsOkUuOSTiFR++anyQ7wCLyG3cQAd1pYpgVXDhJF
rLWIGL4iP2iLDwPxct1Wr3w4xFvWlWiZS+Zp8FBr0gSz8efZsEO2WgKrzJFbA7Zvhw4q5cWXtASN
NfCweYzFfTCHZK9usY3oTOFMmxepo77Yw9gdSe6VoutrZ7LRAVBjQ4dCSRQgeG0Dl1YsymISFO7j
aVI3O69CR9daZGp0/pKEIU1hZzY5DbqQye8uETKX4H3SFEhLnRSPtz0qSkhpr3hfcAkHFguBLagF
bcobPzJs1IiZ8KpXDkAe2ly4NAgFA9lKEKzQEp0p4/LH8z+Xr9BrmkiYM0/lWXBooe2uIXLtTJVv
ooUXA8WRk5XiOyAMT9eF5dw6PMq1D1AuOFrYgvp0aaMcEdVeibPj4ndutmv6C2bu5oabAbx/QgFS
6ie9oH+uLPcluHi7sYWyLsKSqNq2sY/UxZNg+sizXspOfdL5Y6h18frV9XpWvpUbOzwwc4P4kJ0Y
f1cJbAOzeQmMkrvgtAokVmfhJ2hvyF94sxEElvOc48uwdmxsXTE4k4k1VSC76yNqVSAl9GBvsTFC
nkxmZ77h82XKakyHHeD8acPnKnCa2TN7N8y3A98EWMH1nMUH/A8RFte+KZiDUfgdnGuu+vAAqytk
VXwLw7QNAmdp1t7Nnsu6GEmy/a1Fzkr7MUeIm+g5fE/b6tzr42rkJiJhlzObcmuzV14hBNjnQFsL
WWgf5zlMuMQM4SrUvT0UJcYZj0AfdvJJq5o0oid0trADOQxFjFKEfJSyM1HJ2vZRHYByK2fWHTUj
Gbxg4nHTnwTOUX07Q7oeBf0UT7aMW3F83A4hxkQDzP7wp/daMJqcSKLZ+Y3n01n7pDL2F+Kk3x5b
MfA7ox2ppgY42RLMk8f/gB8qiI/cyHRQ5oXV+Bx8ANWEu0eh7DczYUhduwBYUg6j767qilk0sg/O
sqpgT9givjAYosItuP4O6yfNzCQvw9cdL7eoClYUyniMfxATwXfznRqe+XkCekhj70ABOutweGvs
NrJ1F1YYz2vvVb4Oa1YnzphAgV1KZuNWZdhqhGfMifI7eqfXvlYn7fmfmOxCV3G3TgVdhpMZ9R5R
3cmR2DMHGCh1/2qaMDPmwhU5JkT4hR0ufftAwTveyq5YfDESwu3OEdJDYdhdqgCKGH96f2WKq0iJ
ia0ecIVERVlKnkfhtP4sc2o00piPbVrq9eTpWmioEGTs2MHmlXECizR9c4CZnDxzbgcrsq1/sG4q
wy/wAa5FYwkGxsgpG0SpSd6cHEClvjKy8svjfBGRiRgfhfBQ+Se+iYFEAS/8tRl2bM348mBGdE3I
0lAmD/W1KO1DhvC+nq2tqqr5rrqK0yjWQ7VMmTlWz9bbmDyfYhr22rUw5IIMU55UUTh5tO86zDr5
2aHwDCC3/AD6TqMkHkYpV3FxgMAm2RnLqU/sL2ptIZxyDfnZE0Fixp5cG6vVmJYYrnEXhmW8J8sQ
sw6mS+vxtK2Fh6Gi13MQHyFsEhelAo0hMa8ZduoD6BmWgITFoVXC1qFv3jMQOWPdhy1cIi/elYHn
phOTQUa3dhJNhhIu7QtVUltXRT1ii0DSmuLZqS0l6Xb6NhyQKIANIPuU6fJnPsAeaTzBJ8lEOcv9
Af5lmzYuhXu+9jmV/3d+iGbJJHcilxspCInYL7me8shyMXCiPqWmNdukMK+Qa4AAHNVwgYWxKAV8
wHA+Ttv8DfrDUwD5qicxz0EkXEh+oVKJy/HdoZo2lYTs4LKljBpMSyz6ZAVNQI1oR6ASt82hKRb6
Q77gThvCwbjtt7uHSOXrbYxWBwzX8HxfETwGp7bDDEcIr3HdWCQtFwHna9i2yio/9iuhS9k9UYjn
ibcpOuqr5wQN1iswK4whzNNbuq2CaLYOa2K+WOtc4mR2yorkE/u5tGtZZUw/wshQfNHBpadT76ca
dvWNtAmmQuDqApV71tAPuzNDP6swT+QTrXWMCRJPBQAP8IO13PPTMvGn6ZHB6a8u9QHvWTGjTrbm
uBO7rr/RO+wBXrPE+EvSxq1dOu4oM9BNcAJAzgeXP6u4FwPt3UOWd8fnueedV2nePENg4i85roz5
Ehxolt4GnJdneG9s5rQtstd8QckEpeAP3fqbrCWmhSeYNRmbHZl9X+iZHG5xLdrL4vEuZz1OrWKX
eu0fCPddffEareUG0tm0uicrIJDic+qVWaBmQxb+yFJpdOtswk71YwHtMgDCTGC0PyBTn0g/HfZ6
023wKgpUvVz/492KXrxg33oGb/l01YzWj5PEcvfIRL9FloGF4yEpuuMPbRmSV8W2aYYacOIehQOo
PvycoiSW+XQampPY0NTPX1qCKDG+OwRxm8Trlg7FvnyAx8xjKxO5vAbivd2EQuBietzSDLt6JbvX
dpLVescLOo+invyas6uDq68JhORuzpaIMrsTJUUGx3NOotY4ToGhqI3UMy+WXsQ9NhNlHk5iLbIT
r5h3zlU8gNo0Ubn879L/YfYYc7bO6eRnWkIomAPNFvEqLEAYqTKDXyEZVYoJpBsv09LimUrUvRm9
7XAuEvWR2Co/dqY49kGg6aFFCfBW/v2rW5scHGjwSjtvCdRVJpOam69dtopyCaSAHoUz/KDrX5bO
UpWBCzpCfsoR+OOv1lWoM8DhD7PK9H6Z8G0yw9wRZ2pL9ZSnkdPbRmh3NrCd206a/Nx3dKqAeyHj
/7o/IX49JavXAd6I5pYqomUl1KeMZbbprzVCXOWaZF8uAut6w5DsOnDhi+vf+umxPAq/jYbA58kl
Y7KtizDE01tuVniiYiscsYbiwKj8kA1Nzc5a4/Gk7cBGoq1Y9H5PDiT2CUF2M7ZOjp0LPW/HSi2T
LQReZfbPY9TE47R9fWs6veYSmoBDudExihKqc6cenS928shft1GCQcKlPFZx2/4P9q0l5w+RiiIq
qGIl8/1C3ylAP+Y6R9kkjleSH6WZ0HDrjtACh4tH/kb/TMTFlmTXrujBRLv2FYaopj6FTm561EFc
uE9p/T9sYx3dR52oh3drFzb+ucUUg5O1Nm88vt7CBo8YLEaGwKJBD0a/swoPI3qZN52Kvgcc+GQ1
A36JvkLIAOZV09vPwelOALzpP0eKi3g5cxFyTdXVuIJNIHf6AHhJFPG/Z7Wl6dH1BQn2YXhyAKFd
mGWHOknKHASk1C1FkyaN0SQmN5J7kK7aXK5LDLQWtOmVT8AzFjCNpBL2NMNoZdSmd3+c25JPTlvD
J22Vjct/Iy3scQuqrgkOiyNlWUlIkMCw13dzenM6Hy/fRzpw02MjzPtQFrjlGDon99uPzQPwNTcB
t68eviND+1p8SRM5UycCNjBSHRSd57ko5GjgHwe2FGm4cVD7hgWUi1DKjW1g5j6MfjHVjFKOw72D
Il06CAyriXISo4tiM0HQDqforej6NuIzGqnqEwCKuEa+C58NWBeBu68o3t9WrHveaBqyLSkQTO3o
lH9Yy+sRV0RKsRecvDEEqGtmdrpqZ5rRQy9nvXQNS2yScFP/K4JQTd29sXi45/cjM6Tg83A05yCG
dkbZ2Debid/KIMb5UBMagA2qPXOTXKLfUgMGnFWKOByhgT4jOuHOvnTPZ8TzAP7NdAfyVMYR+518
4oZLNjZXmFnwUnUNR2bhmheD3gn0ozSGznTrtBJIPZc8zQugDes91aSy8GN3tcBK0fhjcLEZ2SMz
LElJ921teowRyyuDn0idiOxLaRvo/PPteHkPZHQvxUsM70eQ8WOWWxRT8njUKUbmi9/DNOybI/q1
riFQ0Jo28tKT59S+gnOaUm3cvlFDvkhW9IZ/N4ZL7XJeayMkCWXEBu3vtnD9gAb5UvJpDUNTU42N
I2kRil3FBrpQSA5NHaz50dpV3XgeZmRDbNBk7jGxBReCkS5gwvMqY6r/mzxShlj6CZIVVoiDlVX2
jRGWco2qW69tpzADZsZ9PqphPMs7KdyVyud7kELy5dXn5S9MeEz241nlkbdO5g/XxG5KNleoRcAk
u0+auPUWYETjyh4dKryQJPmvJ0JVtc87ISqS/28rL0PC3EwFntQInM9jtPnvP8muH7AFQliCB4ix
kYWZfde2p0Wz9IIDARDtS7NPgMhezuncvCZ7CHurMrFbndep9glKkZfRoH1Gn0ZPMyQaj9jzXxQq
gmEB+brvuAeZPAz+uhdimV91lxTXE67rl4WzUctQfwMrMlIL/ZTL3Cfmxkrpu2RnV95KGxdsy8EG
Mc/RZ3A2GB8KDiBRAmPz239xpYhGMH5hYaOBmido41skdX0C+GsIRWu5va6OUGPyQSEwJ7NiHsSo
Y7GaulEEQslPAHJ15FK8RO+RgYCXrWfH9N6Cjg8q6VSl6yl0tUUjfkjR6hLMKACvehnw4WiZsyC/
b7K8xuw6Mym72Mwh/gEBXf6QAjXInNb94L0EW27mwX9f/zqGkfvoJaOwfydaKYaB3rxKKzl0Lw5n
iR7Ec1bkzi5Qo2/8RDrzjah88eLoOgLKcE+1zJ0+T88iYCD30ozcC+j9IXAARs9JrgaKsJJ9K4xi
/FfP3uMQGR0Lfgqwcau021H5zKGRyEELDud18A4lYdwvGpU695jgWvZR1uVAZ+P6PV3WnQCxu7fF
edMG9OtnM4hIxfAw1T9p+9LKIqPJVxIR07sQDWrHDdO87iG7FjInac8XeItQoKIGeQ7yx1LbB2jq
h++t0WuBOZGrTGeDOGHW+pIVYA+9uZRbh/otnFRFBDlp4C4oyJLWBRs4Iiuuvnk+Urxp5Tng6xNO
3w8F2rgS2AgFtUpSIcKDilNDcBcO3GkB2DvnN9EWdm9c/y0LfKFeyqNvCMWh5XWBnnBrRp4G0jqW
JbaKgOYk/R/fGeUJ1Y75PtomhOxzXXrCx8+ThNBs57C6SpAKnTosIgoIf06OhG8sjLLhVg8NtzjH
fOoGsepL2YphAr9FjXqm1lf4rJjRfE8TdvIS9YJL2YxUh11BqcrQetTyEeWrWTY0luqCr5zaubiM
VXW37abUO9wGlPqj2TbfelYywMi1zzKnqLTixFYLTZI2pD7Z/VXoWlDHZeg7unHBPATxM0XGrQKQ
7VteCL25/HAzY0tOkRVUTgSCOcxBvvoG8hGNwbNazYnD9KfIx0iSnZW8YFaJ0Keo/AJYMLZid4po
Skzw9qefaJkctOSt7/+Hkz0hlXVUhpVYEQJFjCJ3WvbbY0oznoqDWa9JYYc4OLJvpdbV4TEQlu9R
41ODWeIK17emSzTvD/UivkjOcLtOCM6sKEEqJhI3Yp1wMWW+lKXwT4KeekMigz1mqqoYEs+wL6nO
5q6gYUdFG/SHrl6NggziPt2n0oXDHhGu2aCbeVlCBPawXTDTxkMb4hBQ4kKo3XsgGVXzRsasbJ9S
igUT1mvYuDe88q1rQnr/tFEmranJ974yFhk43Bby1V+eov8uG+ctvN5FAoGq+wx4ChllXQ01bOWv
moL8uWHlSIPRD1DqIkFjRkIeXwO/Pe+JUshtXpPOUelNXyVPj9JD75iOG/zfGJMgsh2yxlLE9LUb
YoFO/OfAhp3/zZyMpWKwSfRRRE9CUSIP8lE7UZzru8kpm8mngi4zv6T14n8eZyGQTO8SDUXhMpJA
7by2qQ6Uxd6nd87Yk8CeJ+XGaV5COtkSNIK1z1+FIFSRRh3ymZCCwHZLCtdtMRbc6XljXgdAYDNe
uFAYOVkvXneo5SVl0umtsmbH2WuxWvDZE988r/ktGeLhvHO0+tGuEm1qAEMO3/G586STUugUzX7A
OuRGNEZSFPGS06Kzn/l6PZuyXsbE4YVxWtk/rzXwRayQ7NYZ9DMhOIeE55LhZO3f8u+YIF2X34zT
etHgpQc0+f6CTPpqcSig7hD5GY2ibxPo6ZSUiLDPg+vKu1SKivjJRjd7mL8VVCVQLQ6MD8BAr/Bq
LZS+7uwz9fcPZmFf8qCjCubcp3fVfgRYVR/J5/PSEPm4o6ld2yRTXvdyAIZuOoACCARV4pKjSW1J
Lk+yYyKHjXt+/FUPllQ5e/aEdUumBNKArI7hkTV7bDXMU/UWQuikAGtJl4t5S15t5JlxJ9bI/qmy
qjirj8/r+0xRDsxzWd3CRCrmR2lknRhbHmDHQd5FI5EfU5BG6XG6vzXtTSt6gxZCryF3EOWiy2jV
IjFDPNqq23DlKAK0yj5s8n2RwJzjD0WCZazUc3jWEtfA4tHBa88j0KJzLzoXwEn3NPuF22CCEpBj
2KiU++5bQ3dgcRIPmmry96R9oKDKjcuQ1EOeoMeyIcU24qfiCeeWnqd6GdTeZfzSghVNlo/DKc5y
NJCSxJ7ShTvEGNtUyuwBv7VsHq/+0NEnCD4SqfJ6mMcH3Luo1VqrwMuq1MAK9jq6aY3OYGAwVvUj
xWWIGmkF+5EoHDmv9PU97Ia3/au2xXJZu99qsxyEB/nih55hXa6cQKkI6IdIw20YsKnK1c7XGGmh
YsUBvZqAsdw9kxuLJcoouRNC+lC7fjr3gdeOYuXxkJS9kH5JrgEmy+gZpF7QUR/TqdW/qNypyHMN
cglA0pAvR8ey5AI+nfscFTkCnMhdJMqjlLagJFsmLOHFvYcVc0EX84x1bApauFsIHBTBncibuIBy
0OwLXR8VBJuE0zoNQUSarqs5qs6DbHv1x6ZQfLZwUSTJ4DZKi9nAEhJZrUVHkwZzU9CxuGMdMI0Z
4Wrb2NbiPcsHi/1zyR6IuDxA3ltzHxcyNEX9mb72pzhzHp2MyDbNHUrQO7BxhcvbHBsR9uLGA62y
adAV2lfJjX7dm8Z3bPOAYE/cfneGA7HHXTItUi41LDxCXQMIWMM3ZRmBqKCFWN+mdw+an9imjUX1
sJY/M1R3WNWIKlKKgY5rb9AGDjmndY7i1phmhbACB6kQtraS0H34ZDP4PSl9rPbAu0I/g3juRkrR
KXT4ZAMytAsqtlSdmvGw+ulV4uKPniF9OSjgzXfexGvGXbTDosYcTY7P5vW1OggVOj2f+fZCbZIM
GHJLO6LB+oALg3rJwoPxsE0S+cvoxNBvQn8uZ5nLFa3bxEgmKihTrf7fYo9jfOymPK9CXym5doZJ
iyPmU7CVmeLXtQ5f/OoufHhs8LO8jUL5qqr4Gu787rMjmuQKiznuKX78l748n/BrGLrkzWwjzL0o
TmR85WgdbeN8dpaOWU7OOXllNQJ1QlHvtdzu341S/bRgWNIEfjedBJKcmiRs5/9uJEzYInWBepSv
yUVj1zK1iY/RxE44M/dqOoLwxHEIEmz9F4M5RaIZSSgSgtmdc9rpO/R7N5wlwzkWQ7zrHrYHupWI
akBcwseCqFpcK2C/IVRwscWD/S9huwZNtrJeurUstfVQuZwbULPXbx/PuXc2O09NXfV9AgNZ7EYF
nfWGOq/8X/MKcG8N5dw76fANMoLzpK/u4vUJgz0gBoYbT5ACKPj19VRYOjVF0B2M1w+sqNRI+gvq
h9MUla278PhfYoipOIYtoVtGX4QkN/Sq3BkEskT4TvoWtghjNOi0lKRpvVnfnq+7jF5grhRBut55
7K0xksk+1g31nZTuALNUyE9+P4sJOrpnnn8trljfXpma3i+v78wMSWZE0Nkl6Nr/2skYT3lYWrCC
YsYGAnqfu964z4tCr1QBsf2Cfg3BdvYB27fGeSn2t+r+UqQoDnI3I+VX2o9lSakjVBvANZWW/AYh
xqnm/ICobZBvfkQe55e9pFJUrQfgyyHudjJ7udaFfzC2uSMgXn4UZlVAdnUMo9b6IX+0zZOwl4L4
d45RsmesTH9Kg9I8SndjOz8SMWjIpTLyxH9qvYO+IkkIuIFplIjLrnjWZicpyGaGzSX4ppCcZXB/
dokLHiyszoRTd8JqHy3dS8NbVQVXUnSqXV05qAXLpqGKiSj1UcYTH/UFV+KWjRrzUxOhiT19/r1o
HdWae1ty2VrhHpYJuSZbWIGZC+EJmElDvoZLKfNZNZUtKkT0y8gtu8B7kOAy1AnIhY5TBCV8cVcM
vnGMiEPjHalJdHU+ziuPz6aktpUHlwQ1TDBfPmB8XbEH7/0WrNjVvEd8vPL7uWP1Uung7/TqevBs
yzkGVsoT3u2u8HLS8+SSWjHtBgftPTbO6oRRW0qukr4PxpsAE39qnSgrKM3HDHUl7+BFmTeU8CyO
3aY59SX4QSw4X5frBvg/z6HzUOlGTVUAoRrZhUuJKo9vkIXHA1CvKUWrvFeGfgyJ6iStMH02HXWl
Gn+B9zwYJScmDO6q3P6WEG5EGwNYJKHZre4iw4aAZDcrDs+CKD7MAqdOPl3DNOCxsLWgkKkBrrrh
hWQAetCPk/KVJ1187VjEyAy4sddzR2zz+vIbEuGeENgvgD5iHXxOPu10haD9H2PcIjwbBdcGQr/w
aJMC50fGSVB2aqnn45AFRGb1i4KPQE4nLTf9c3O+EOksBeIOgcic3E5HwzL7x9wBcb0tJYNaxdjs
pvtfRN1DlH2mZGZG3kDoJ7J2i1macQmgszX7iKztowSSRRGjdTms3+L4Xolh+rR//c496O8QEmfy
0CUvorFEhn9nut+jCZoVI2poMEDKj0WyD9a7lZJJvaeRbD/Z6764hVr/AOl4meCXuG1fyJSGV4NA
RfYSYiQDQalQhmIcBn/cJyGs4TGuD/ceL9mmFwLA8ZIa8C9BxFRYcB70nTjjCUegnrMMdGhwjH3E
seJEMUKjm0HVd0zstQeKHNn2bhSt3qrC7L0jyyhnIcHqyspTWkZfURHN+lfO5lIzijyTHZSFQC2P
fJA9ycM+F3jQN/Tclrl5mfS2B9TSYVM4MSZVGyV+A3jV6vsszxAJQyGTd4y7d3DAK9lNwdnixgYr
tgfH4dzTfvRS9+yHu9J+kgkY2zrDtwp39xB6kpoSIOsnEcVTGReNFaQLebsnbJ9jAQ1mLHR4WO+6
lO2arYNZ/ChTP73gfSu2UTDcTGJ/ghn10Pn0orJNVZdOXZ+IETGqyatXxUDVioGwb1R9Jj3R6Xef
Xl78bLFkH6PCFi3Bq64Uw/l26rVJ81c2cp9vt/3OC/kG8ovfhMbRzZMKnH30meazGpiyEhXnQBwk
LKu6ho8dltCMr6emYvKAn+E0856A9e/0oHI4y1eWN+2GPnqW9NnNKDCseZC3CDxtjG9K9z2r+sni
hNmF5UvrqkVHrBnhp+ogiDweImHXh0rtx97lSVm8/JPEvI4D2ZgrhJ1O+9N1DKUbiKDiwTT0PjnQ
tmpBUzxUUygGaE2xiZBKZNdZzaWd6ocErtYN2L98AAcKp4RwdOKcVYsUFfNnQgpnijdzluxtlD0l
f+AzGopx0qId+43UzqNFwLc1dJr25/g4zIlC2xL3winE3pIxpLv7wlhyiaDIRSDbVLICSh5HtKHr
faTW5IH349dKO6CibkhIwCBtlNowj/RgYdyYT4Cd17XHI1fNZU/jR/n4MTDZCCYkVovjQ6+cL9iu
cC5uQPkALovEMyQR/eCjjEIsrQmNPXeMOM1xSaEVKTb9Ef+4k9/0Jvs8mMThvAhNIy6zh6gf9ye2
l6YI3TDSF/Le5ztUnzVEB+vmJTlGMs1DMOvGbMHxe21slg4jbXzJoLIdC3gSSs43TD7IUVYJIpsL
YRsaoQ5f1mVS5J9ujhklfT2lzsReFLpeEDNSWGFhknY2p+hkRzZXhNZEewogdfjp3PRr4seH7hAy
C71oWs0yYy7u07E+2Po19MazK84sxfxGSv+Y6VzMTnhmlWuaOUws5c3jWILk7+jVS/0L5SNb2N8B
MtTsS2OS4IvAHCROXOq8GNTf+C21UVulxybIV7buQ6aXYVIVTKLdt5EhzMl8h90K1Hrbj1n9Bz8d
J4PijwhArll3ZqnpZacdKcz0TCCUaZ6QIlQKuCNswHqfPnDipAoWI7izHPv5cue7Yw9AzrKE8vW7
YS8zO4UYo3NiIReBp755NJOa8/4ODucgN+bKWWcaYlMOC3zvbhdzidNsEFGpM5cHBtHhoqVleFgX
OfLCNuxvvWTGcWLR9N2DT7QOlLHC0nzS4cvWWya1BniAOgMtFx5AjzhGFsMr6rrENqwqHXyIlIdc
rF/DaZW0ABb33luznfSzz3GRgnUykSI/ni57y81WmV+O3mK1jNRjg4BGhte3pHp0/z1xbcUQ1Dib
zKieYGxnr4/X7gc3dLYKNekSQ2MaUUFgXNpL9TGMS06DTbXbKkBzzIR9GFWOtan7fx3L3n8UNV4Q
9fVW81pYvRFVepMlYOHeVY/RVFFUWjYXp/O85YUyGDolLKOqKMIS9GMzdcAQYa3uB9cc8Er9yZ1J
gfLthZOvPdy6oIX+7UnmhFTCyDLjCCPjIV/MaVVWZ4WaKJBRhI1ym13DDrwF+nLxt+RdeHpw+ymO
Kxmo5qdo+8+fV8CRwGfC9AC/g3v0itfAHeIfVIZl5LDjn0SRNypk8cWdhNxIb347PBloJ0WfBsZF
8lWd9tu6fQAw97VbyAVM3NFVuYBYxU7Cm4yghEqW9AHdtGhB+85dNQLxSfjd3PGVtN8IRASFdPKc
hLA4dpH2vrY1L9Q+dN6H9zOdi4hB72fClH8zjVGo6vsCK8XHcvsEgAfOBCIZzrPdE18Bg88PBF5R
qmzpt1F4aP9EdEKC4HBbccVKcrpd1WT+0oSxdz21zLG5vRqZAAnD4fT/v8st0B8J2fruvcEbOV6d
rW+woiFGL94mmTrOA2iIuE+dN2IQxgzT26U4gUNUoJrr2ng6xJbMIDbxjQ5gV/Br5AA3UstCN9hV
/GaXA6Z9KD8ts8xfSIy+t3X+I9t+qORpOaof8A4jW9a10QuLA+OSPPwrFtwjQ47hxqajInLR/fj8
bKcXBbzSiMX3VJLEJXQNHJ4GI8opOLsWBr5qGS3V91HGyzxFx9LzkBi6ihh1vMOUNmkBg6sNbC2W
sXe5MRRoBdlzqjsii9GlJ3vMr1uZ3kgh2Ti/LU1/acfYYCpjPUPRpJjBQVCwMQkXh+AvkTdnio6G
jhsiFgIVCcIHBmfmYlmb+jOz3Q/9rBtGNtSgsZfsd1bCOQENng1kwfgtFYctvDP+qfIfmPHCZ125
Mmpv295iAr4TVgVLExtkBCcD1aOo50/EeaTAbsosAe1k13Qc6Gv2TzKWLbGodi49W3lop9/ryLLp
MxpOCAotpjVb/X7nzqTfrsMrRfRShiWvql12QB87UOD2vFbnVuFOnk4+1Ddi3RzBQ7OCpoBKWZW4
phFhzpOjciiG/pNn3d6gGIe7zFt3LzSATK/zlSTQPwBHPLXeW5KXbG9egOwOvhgfPYsfb65noNFl
L2NWQTyOdErq33cfswv+jEb67MHxxIj20tuNF/kSzLzR3K6KDGd65Ft3IppWNpbcs/1esatSaCQu
Bj1WIfReegOk71e3yeI5Ce14DBR0cFz0xlAC4nW9z8R6WsDpC1S+9viGdtFf/XTxRPfQobx2c+xf
WKufLdaXmeKiv6ALf4Mrf4WUPZeNByKz/dzXI2WXbbYCS/YS10Pbw4XTDtQqM0pU3JiIhwHzAHnh
gEXdp1lW2DhEf6MMlIrLHstbx6g8oFLZhkK7MhDcmfrQXaWXfwvOZsWQL+/h/p2J3bRsz1wLDXwW
ofTeZnWIBiP4u2irKVhyZDP0uMiZ/oglNTT2EKne/n5btSbTFU0B0wRK4UAIO3CY4A9UBxn17XR0
pItpEjFK8epwxXdBRKPxeEoZbCfuxMqxeRHpcdjGFTWh/Wr+3LlvwwlBboUPaIBirqugdTMf1Z4U
Yf0myC0qwup4hZDLUl05OvZG14Q74ig/mitdZn4pCzN94kDXS7UqGBjJZBZ3Qj+GUvPZZn1hbLZJ
BTbGtJ0pnld9Qch0pqzebNeYn3ty9HncyyJ2W0dkbzPku1oO7lzLs8Sw6mEHOo7Tcpn33/rtrK9Z
fq9ZvgYHvlYDgirVtB8Yy+l43F+kblq4HYyzZmCjLNg6ECZ0p0EehsMZeV8Ctv0E8ZMJkMkJa8tJ
hWhEBVP+7zYr/5phLdFtJATtGpF9dL3u7gXJ1vAsMXXueR0KGTu5I0x3C/geRrloU3RSORXwcBV/
0XINzU3neXWbRMZLvVAIKemm9/13xtIng0OjtYAe/mChr8D57vWwrfLEeCHA8ive07v4spApVBsT
sJUcF/FqGaelXwnuHrRZt6/1zsgH+AGqJW01a3AiuttWp6P7YYrD81AVkqecWTt0KYdVUIZrEZVn
nWDDOlTbqv9TJkh2mAeUmWGIn6YsVxkS1W9Sl5zaueEObn/BFfJj8K7M9PnK6wpgU+izDXkGRoEd
vk+m85AaAt9U3RLNztxrj4WG5T7tJfYiICOUeTFvYq89gYcyTG308VjugXnCOXkQlu0GJyk6MInq
8q0QkeYKGOhuaVEY3sdivkerc665Kpm6oFFZg7PNOfFUmNVglQVtfR/6rQwSULZUN1Kyn3j7c35U
wXB7eDwx/j8xQOfZuQww4e13Ab1FU/hoKstRsEFjuGsiTaxE1RLoN81LFfcISZv9DNseMBRiEnay
XIK1Lhup2/MwBvCR7TcnL1phUBY3W/qp+WraQXcAwDXJ19fVRS+/iADWR7R8RpVJ8hscM5WzMi/n
ZmrwCzh8jwiA4m3yL7y06p1ZiTGk6bBeBL5l21UrKEP8WD8pR03kQ986Lth0WR6FHVUheXUwcuAt
LjW5dObxGyqdedfLvXmJNQNDOFbLBChIGj1wNgmZ4XKmz6wwQ7JRvlbP06GMv/93HC1jMl5Sf7cM
lQ4FfNIUgFHu2hiWLBaGB/YU04Vyl9qummHbV77glB4mcexkn3vzOHP3aXl8lSXd40fKZHOg/n6O
XfoMnU8Kp8RsnvKWMLGYuwQlLUQe/x1U0N/K201rQ3R1gud3WHk47Dxnlat9b9a8YYPKVxpa41vS
v488LZ1BpuDs+fKaOHFoKqn2i47Rmx4ZyFQqXkfzQXlCgcWpiAFMapwuidub/Rbnl34x85mFM8PI
tKa3HOlvp77lnC/sxlLtOWe2JaP2Of0qPN9FWIig7PuWtYyMTsYupxTLvi84p0Ecp6BH4E4pKk8t
yke7Cy1jR0Jmq8ucgg0LZELVkXWblKSRCsV+x2alEPCdH6Km5PcoEIanx0YfNmUf/ugkFOmuRItM
Vac9RAtgnxXbSFtFhcFtgxMtI6Hv9KgIL/shnwgFyAXyMQlqfCMSvq+TBuwAvYMtZ4MRSZVL54FI
S9O1Mvbhk4LIIsnopP2V5Ng2+J4WdfZLPDYEsT+Wrdy5lEEKYCJbrwlIGO4qItN5s732q8gxkupe
w6mCoXRfVWNbt7Fn17bW2SXqFnTjzHglHvS/eSL97mk2DFiS/AWgjf9Eh4UWYtNlZ3wuwWSzb3Wg
xGUm2PcBsZ7S64z7UHLdMawSPePgCMH16Dmpm7yNFqXDD3pJtK4TO9XFvK88fFM/tzEuiUboe/Qq
zEzVTCAb3jR4NLMakXFsOgu5uOzPlI3+LqJc+5hRKo+k5M9vb8c1lgqqOT1HAh5E/qi4Q3l07JUj
VK+NkuAjsGPMZjTeBO8RVv5LBsp9dBF+dDzgepMsLZHDQseaaReqXiepP4k0xVhbm4CmM34LDOQM
2D4t+ArEp/b2mtYwphui9ka0onNkF5hitSm204Gj2UxjC48j/Xe/PAsDKtusoK41dDA5itbgOG1w
oOq06KKol3LGbr9a2VHxAIL6KV7C8m77xRNBCvifzGyrawGtTCZf4BvI/OZB1ksnvs7bKlK939vL
reyB+aqET5el7QYhvX0vwMQ6TBvIAUtYK5rUTPvfEbl6Iqq7dGBrIuXyT5SdP92CnccXGLLEYZZ2
hlSGFC+UZLdKsKVXQlTynbotPCCXCzOLLsNe/YtJoxZte21ALCOZ5eseAP2DLHnxg/KjXTb6HpsR
c1Q6UHjHE0ZvwD22gTHEbI1Ki1Bcc2olgJ85pJ/D+YeytafCykmaGe2Ok4/XU67F2tcfDcg8NN0M
jjHvO7hX9wUAym4X9TGMMxFyiA7UIQx5CLBq0h75bU/MkaQyhbC5u6/TM3Bx3J0nl0IUJ9QSy3hg
lFyLFUJSU16Y+x3SllOh5qcsw47jJMZYW9yissLtaT70YLm+o8d9qhjY+nZzCM3lUcSo0jI2vJvF
fr+IE7wVgffKb/5XIFuTL8FkJJxlZJs23UUpWiMwkKDHgfbTz12wiUm5VaBDr29HG53r3axJDrUX
tG1RuEQvVXrRXc2YnI6gRj5wdguO3oF4uirlpM53V+PNC9sSfyjcsb1hZqvMQ5wl6jYjYV/Ujeg0
FtYdfVpB0HYZxXaJ+Df8pE4f3QzWP4S0BGa/bfy5+sm01BuacNYYTSo8EJrqwS5CEEt9TFTc4RS3
L3vE3mWjabZMBWaZJTBxA7VIY3H7diehZXuPnpR8sfoJlKx3oRSgtiyuOL+J66clsDIJWOwoh2QI
ANW1ls5TOmPpkxlAOkMt+gWoF/MVHDKR+uXWyj4n/Ng2BQZJJEzrfHKB63/GrmwIOQ1yn5j2lcQo
IDZmrGZqBYqaL4LcaI86zrfN4+3+g48WQHUTri/P2thWyl3kv5yh84vOkP2CcuLSZbUoYCzvJtqp
kgnX8jxyHhjXwszVLD8JHlldiU2YgMLw0mBBz0JdfAT5FAYvyCX638MCyxzslnWhkFSqFk/xfAcC
F0WQUh7MNHXFMqN07VZmVWqzUARUdMMLQO1KVg4B3SIlTEBBoCZmWn452fzf6x3skVps2wPYs/78
6ErurFBniim/8ZbhHJJCB2bKVx30rlCAMURj4yImZ0kANng7vtpKKJy/YQgmm9UVr+QawhLCcbuH
QwF/EldEpk7LhvDDToCErdEOTTWEHKQXhgfjWmhjRFt0eaCG1L2/1Wcj0I98R3bHGVG3CBjRdHWX
dCg2glr0g9bjfnZA7+8hC6b+IOxIhhbdXJAguZGN3B0/Fue3DvnQan4VjHZu0YnYBBuUWcv3WK0h
FhWEkoyRhXnOx4wdDlnBaGIfoqmjzIvmQdPWPa9vHhAowVQmVnYZ8ec2/s1YO7SKnNrtJgT1CfYW
bZAtrAFxaQ27Osmn6/FaJfr5CNXAgq6I6faEG1FjG7/UH2aAYOXYyJcbRxhF3qDXh+Z2C1kfqmyA
xUr20zR1rM8g3WCib6i0LiKnkEoh9Vwr11lWHdzY43zgHwQHmJiDS0QdemK+MoKiD21z3PI9jEhe
2fbiVW2Nv7o3hySACTJVhRJUPQALBLwBpAJoAIEqEcvCr9tpYzL5GKrhV5ZcLaZQGlaVvI7w+SO2
b/n8jwiTKgsh7InUJRdj6f9B6dCKBArt8vSqmWFNhGPiAYtBJKZTKSNS0HcdysaSXqa8668YPTWZ
UdJEQR6Wg9j2DUNlsDXot+/+Xa8TgaRVe6ftlHwECKygP/ekpRMmXv7vBM66kIjoGbbPZPR6TMxx
QZtNCSpxDW3vq0CBQjfkh+9XEvdadSEDwBf4GoQnglWbqqu+r225Fvs4y5t39+J0PvsDJJT3DCin
+iud6yN5BcGEmg872ExXMFn1/uIivmqS2ny39EPCBzj+vTDNGco0Up4kAoDpr4xJW6wp3c+JWQyF
97KPzl/Wvu0jN/9vCR3QmKS3ok9lIkFUCVRJ/XuFSJKj0PjfMU1DzgBHuDF2jNxodKV4VVZ8nNwI
AFFZrTvXTw625zMSWgWXQQeSMuJ/M535DZfQUNRCyJuyfvs40D78I0S1zv7cxIMgdYxuJlG8/Zzv
5R9SCD7ojAjWaGffm3cHP+UdBCq5FN3B9yBZPUCLoCHjlDx1TWLlB+52YhoovC4e6tDiMnSnnIdP
Dqb8o9HXguYMogr5hWQAzxrWqXREWF+KO3qdjTj739cyLa5N7HsplA4yUOREgZFiI0rdfiayns+p
OLTYmHcY7MDnrwUOovSlKX9i5RWOljRpCsbQUmSV2DS1eEFaCkH2NDUrDXPVHbFrDr7lyeuHzAvu
yS4aH+laPGsxnGkZVedAHEYHKd3a6wSx/pPP7Z0Lny24eoOV8tJn83jZfzOJ8a4bGWKgivHR0xZr
ji3q+9vheYNl5lntAmnr/j2HuXb4oDs0LsMvCk8A1WK6GeLZPOPRwYT2xSHXeubH7yU2BbQkL+V8
48M3YTn1V+RCGkDZiYXMZ5jgCNX5DWOGNjMb4TmrMSDufxSpoyJ/i5Fc+rduacZqSO55ySgsxDwd
IKv9veradZENqn9uFj87QzZvuAy4fspni05lcYsLMVtXKeUauF74sCeREZA2OoF4k+NHLxCe5Ds4
GirV/rD4DRMPK/WsiJhw03QbiIPg3eBAISW6PWAHDkFiFKLdxkqeE2J/kM9gl64ys1tzqOhbx3+K
JC4ZjvIoVVOzS1wi1r4/b8ta5/F5QutFYtwZO+C8YYd8f7Af49gMKDl5NDtMHe9AA8IXwP3ENqbk
fgd11fsMbJIa1sEeZt5z3lWhBKU2FN2Agtw26cTsb2Ad084H/hHjzJY/RWe5e9fOkigrSUOdl7ZA
HjyAKADHKXNJ+XKNjhH8s81tfvSMk1dEFdQIgY50t2efrf9v7D+iR4PZ3XxavEWSiI9PLXpxR0bK
DJyB6NI4YdChBC9PPZ/dOM8DcTh+I4Pb0qu3GSInVZjwtcQsEPVQ5x3JYFTgbvb+HpgFLEO6xIT5
HGEFBhTTppUnxORb0OBzP+E42lvERLnMKPQyEzg/h9gULcDl0qshhMexOS6MXqHSaks5iSdXmxRX
qxNCC9uLtqsIaq3hQdNhmJs1eFZN0uD21vJxA9yTybiMxHyhh0Xb2G6BRZSbqPSLtlI5dmbSavjB
9ir2QJn+th+c/FtjjlvggviqzhLE7HDIpzHyyjK7+vH3tZdIbmttBuec0JZbJou90b9G7ajsmAQ8
l1PZnjSehPY0dYZjxgsxsB+jSkdk44L/olNvTx9c2B/RH6dbuSMOpsvVsdTws1gbMHAnee+Jy2Yh
rO8dpSQLX3Sti84RhVdPP0NpGyUFqp4P/PriPBGks3lHfXNnYCbly0oh0VpnNBx5TjLdfTavXNxC
qdq8D+Dg4idMK5yHL/8hw/3t678xGyWE0QNJypL213OYoHHYmpcI5QoJI+h3aeMOPqfnqFGRXajM
h7VtR7ZojEJzyO7KWTT2VdjZZzPKaQm9Q3xvoeYZ9IiMsxxaRGaikHd33z/PCca6u5zhi34UIl0D
nugi/31wsqwkwM7FkdZGGCSpg0mf26cx4vC4f1vf0zFbateuK6odIBmgG+QvMTW6B/eM5/xKCWyV
0kUOZVqm0w6z4SPh882k4aDYefoPorbh/P+ZC4LqEGyklvPnFEVtZMXOFwTymujgczHYGMWOzRbF
yLYQkUVx9K0w90DNM2RnscJfj8rTGk9KNgIfvTDDmkflnrmvT2+CYN77i2uR3znqh7J95kgUblcF
P5L/KhCreTqaS7LJxOzjWD6obhJ91ckwQFmIXvzjS6vsjV/TuR/62jtasbVdjiNkVVL7UL8vPoYO
4ahIj5freZozgHOH4GOsRifS4Wp8UilIc3Gtluzdw9rK60u7WQUEyLin4iPt7dpr9Z5pqjjs+QiG
MwbcCM+QAVqq2oraYM5WYjyIBTfjiAlKIui9IAwJCWgp/MZh1KEBA7+aL0TFbkrGYOXyFsL5SWfC
nXA0bbssSD16SY/JC/umFleDsNLedgTSoJIgwxNsNeoHUDLU/UpqgB3L17YoNj93k56Ur4bDnpI0
66WefF6TkaXDsdMmyi6gEg9ZFhgHO/u1lpqcii5OHq9k8eS5phmWOOJ19Vkmeqgalsw5KsJok3S8
RfSzqUhZRzDVrgwzo9gRLUCJYWd3LWN0Z8G4wlKfDpwUr/2+orZxS77tMvoqSZGTRU2CnIakqk3+
ZAR9bSBtLXQXA26h5xRpQyxMXCWubfx7WEsjP2cUr6aGEYgCUYk0/MCBncsUDzr/kfRxwxyqvvLt
jcrkibkjBj1hbEXdbFY3Jr+giJ1BIQPeNqLa8uatRBKY059IoC10hIl9ZPbs166d0E3cbXL6B7db
zgeZsV8MwCPkFhYRQ3fhhoLeQzP8ELcTeBGC8eQTkoV2XOquNNqNYxrDJhvH+BwMnh3dn7kOC8g9
aIDa0pJbfg6/xKehxU3aiZaTLmBer1eu0xpU96a50OqXnjtRfmwbqseI/QnRnvmPVb+ZU1t5JJJN
ByyvOU/sdkqoeQVJjREF1o6f9NmISZsfXN2kSNJtPKmfUtiwAnM0TemmdeqYmBSNaj4ri3jvpr0A
T43rxJo8O4vPyrMhsHXXInLqEJXl+1ZbjwK/e/b31zCz2KsL+XGO5zXxYFZY3ezJs+MXj7psiF+2
WfWid+8pyXmayIsxeOnmLAQqM5x+LbxvOAuJAVvUxF1XyF+V2UpKiYLwVL2TUrl1/rDFCoUG2I/Z
GgLSW4+VCi99Ty0pI+4KZTNzTEsMAYy0ZRE3Jvo37QLbt8GsdXDH7APrJTWNK6Qb31rfsPOw1PE5
WO4II+g4EkbQH61NH0FPNoFStJwmrP6fPMNqIMe2ZXhkjQao3pPqTRPmko/P7xvHN98YosJDEVwI
2Z2l2NXmrKZkF4ee3tQGqjI76BuboYbX23PP0oSb5K+CboN75hGkL3vAcWwQ/k3gR7kKtdzfL3HB
tMpZvtzfeo6tMOH9p+EIB4oBUqKs6aLJTpDqV2o4okn0i9JxyP64Kp6j57ARWPvdkOv+cQ2Vpe+u
y9fIST/+1uIJyh7/T8KDfhBGWrKYtWYIPdek5c/a9n+MI8XnaL5FnzOwRG6nP5Ar7hQX5tKgoGIf
vl0VeThheKGxLqcTbaYKREsmKzLFlUwROJs4X1OznR10SoiHzOPPCYzwmUGkM384Jh8wrjhQxlBk
mDcoN9vLup9+xSufKgRaq9USbZ9TGr3KsHuAYNqj5aYL3igQKuMX3OB36r495maQ3sRfu+UJX8rd
xBpdpt6Lr+sQGMahmp16wsWaxw/JmfvpBkNZvF9m5f8vDOvhK6Cn/nPlAV8O0MGivHHdu2p48USQ
57cy1nuECGbwyhH+rUU3eKbYarhSpXX5t2GMAnxhFhkW6/i0+7tepqmhTD4Kn/uWsmTGuIJ6Dk7y
bwOwyMTbJsZZ6gws3MT6bfbTGHqE3aDb6OcgmQ2UKgp0BbtNsUBGfpfXs+KsB6LjLSIdlgcu8K5S
DvLWAD/zOxEvDGNIe2lhCKonMTTU802p9CH7qNsn+e0k5PZ35YL1+yAHuNMIVPXtehSgLChWSdXz
wsecEi8G6uTpRcj9QLtvufnc30qOTOI4iTN098xqdXKHWYZZVP/SF6IT4KT/TlPiLSGbmMMVBtre
+LcxN70jC/2pdiftFc9ATCQdNYz7yVJ0oLg54JJfsu1XI/lfXORDelLmAKQobA+zuUn/GgjAdKbI
BPteiFytTkv7xXxrwPjTI8ls9S8y6v9Rmhbf0OOXea+t7rCxHi/NLGNRDj2NrGvS1PI8QYDrqkk+
OqGaul1Ucnyzi+YqfCLbUj4Znqi2YFB5o3uW8ijmIszqG+Sa+Tdi7BlLE69AhyiIpKq+b3e7ZGyr
k/k/+zhcA6/nnY1O/mY1B7d2n31IaO/qgc1pSvGTnRCm21mwFRhKhkh2TzAlA6cSNZVbR3tYq1II
N862IH3MzFSjLFkSXQN8N5tX6Sux0JEqcCIdCqoKooP9crt+FOUsF9cwUIvxbUoKEtK3goGarJwg
tUu3KN0t+nLh8NWu8qLVM+OqSqmv9i2XL2EvkT6P5fUr3g52IR5u78xLnqoEU/k0DqWxMaXUbL3j
BGvpcbY9JpewVnIrmmKWTmfiNfia2Po7GhtBoNIaS139YwnY84h0cJHpEVd+0HFqq1QhzmRjb9If
QCvYuaWTFroVMtdJnClarz0TcNo8DJYQpDT3gkT3LUzeCA/KQxEuBz8EDhCLBrb1OC+CzLoFGq+M
/cJBUeVwfS+vXZKwsOV38nSkYujvnCT25iP8NX7HAXPGVx7ozFsBOwte9ZokoYqfBarPdxRTxOIf
NO+HUI9nafxFsmFGH+y6xu+9FFhp3AIXdH2ngjoAP9a8eMSwTU6RBgYK6K4KeQsrH9PedVzlVvGq
PJ7RGSDreVjs6DHqFUeiagjEcUiF4XvdXcW9/OUpYKHzhi3WtpQtVLAMd7aBIJAPMNYuRoNvastm
WV4DFfm/D3K72QOBbsUh0nCrj3vae6qRfZjcMlRJT0lsWN47cifXNT3o+JXisMTxE9BXYc0W14O+
Ew8fhHIuimhi1RfEtcZSpUPhaUGAyBLUfLOIkTgqbKU/bw5AHZRsqLCO+UywjkNfoWbP6kIq304Y
PB8apEtHw4kYRW4zsBBaUFz+AbO/rYBSmBAIBQDBg1HVZdKwrAzFvzVdI0nZyPdjzBVyhrYrKISF
MRGaI423PMiK4hu3y0U6NcaXYYVd+xZliwDAJwnYVlFfJpIQWPpK9xrUzPswrrf+ZRK7Hb2zTjfS
qO5cQieD7VSkp9qQ7IaXpX/LdbTUf5z4Jz8ahlkobsTT5xxWJt0elXdGiYP9OJ0xs3EzGKW4tz48
PBJa/LZl64M4W2E8PYJrtjUcldd8aJ6oEtMXq98QzD9a8f8g41A1Q+HHDvVXB1IYljkIgHUZ2rRv
vJ45GbekTS1AcuuHAhueovBpXb6D8utPlUmmml2+GnPCOOz6Qup58uhkS4J8UrYSJLQ9pBfJPvuR
xDjT+6PdVcYl3WaBQJoM58ThiI3F9QKcwBM8i3L0M5X12qwdf8jNfYoain4OAtt/gtVUuqn5s1qF
BUiiLfAxl3fBYX7gMVCKK3ooQpdLTEMqKKRSLbniGzhsYXjuFiv3bmgifwNNuS/STW6bv+DB/dlx
53uwXXisJaScpDorDCgd6TtFx+ikerIc8YfFo6O4aubsJhFlEkW++0SwVvRjE4O5SJ9ZZnnLnoX3
KSxsUC8Nr460xbVOMIq0O8Jb55vHdG6qoM2oWA2BzaROclEtU0yVqqNNUHZWQgokK3zPOZQ9NJi2
RB5FIbQ6ZdDZ+9+GVMra9nDkP3PFjKNkA9hWgs/S2EZ7xtEoBz2zSF9A4dqh0y0hpJeedcwdMGUx
RkDhUCDF+v50VyawYOKgFCGK22Kf7A+HBKdIrzIYWNnk4slDpInLA/loC+2att6jmR1/UE9A2eJ5
yCSFhFiZsNtCuZQ1tYUid/vFvrTp4bUgEhP6AwFFHBj/CuylETwugiARu56dSzFatjos7YDbix4P
Df+8vM3sdkomwPObectSp11+BYuMFXB/VtF1e4HMwnAFYOU/IXwZJTwXXZt19JQVIv1thHlwyCjV
7S/hAG56z11Knjz4iOnxUr1yRDGnPCEq/5aMr5OG7MWkH4JNtAqBpBnJuPByNZpxVciFpKyfoRvc
bhFBoKbQTHsugOMY8sBXboFXacnLUnnmr0S7QuQQg/isQ3r3gvb5xMhcZJgghIPvhCnbTzON2Imi
lfrLZPXdYoGUIAQZcQbyOz1S/BSqJ/bmkj9uYm+n5g0dUK2Z5AFzOrJFvNhwtQNGds5jo76RLbQy
GERgPH+3v8DxXZE8La/rAa123XSjlM+59baz6EoZik4dHWdfY0IpyI3d89YKJDTqjIrJCwFjOgaL
qhkG8hHa7VSzXn7Qr2A+/E/gGpvXr+vdGgUyJsNj0ScK+rQTO1S94dkMsYd/tJAMJKotZT5uAAnY
EFGxQ7BEPf0MxZIk+t1UU0aYkMO/sw6jFCGV2a3x7/dN/dAkQd5SGWnIjE+F+YYOld01mjUsh7tP
ZBlVgDUSLph2ahvEsqgyFII2yeZY0hB+OmF1Me7xZ/14bX1jVGqiqGQu9+164H3ZN/ozBtQSvprU
ItJYGraQj87DIF23zk3u93hfCgUylONgmHSHWhQbFMpFX5jygAjpNRguy0mYQNQjeu4SiR2wsqth
kbfVmSEhzW2ogaWxk55xoSnUck/oHPHBJjcjZdnq1INQrpxmzdc2x4L4/gz4MUthkmrG9skxuzh/
Uo0n2ZRDPTh19zF7T4nMsIBqu6k5HHsansntJ2HiquI5eOUjwGNwUv2jwON0lqo3OYOyR/O6Fm59
TLZ6R0iwtmPNwIwmWyDzMAsknnOK76qno3Fox810kCa7yjzWKcOSSkf5O7nKHQGqbNBP+SEzLYVh
VAKYzR/2CIYWXEbwAtSZdDE1Aov7EARStKIdO5zb0FNsfF9h+X/fhNB10BSWK2Ru9TeFSImU9Szx
0KCUvaKxS29D6KUYOqj14QsELpPqZamG3VguX5FogvtaQEY1l0UtxWox8z2wx6ZkIcph+RRBPpNW
BxsKtyfcuLeH1XYvYwdlLo9u1PoDjyVdMY1yb17d2AiIEotASvBxArdjtshPB2hJRSt8pKdUnF7J
NoxxWuOTRJA5wvd3DsyEOK0+prifdW+KC5/Di6HfHiupqs1rl24bjcwoxDeXPr9o5aDhQye93bfY
137jICV5TFcok/cwsE0omcGP4etoGpAItYb9Aysr/NixKh4juweEXLlTNl2foQc24CNakzHLYf+6
g6VinkvACNQpoyZBy5z7g+mqMo4G+cqJ6NfCQ5YD5ipKKy/6FcY0KHKGnSO+fGkxMMWLDxRPXBFA
vpOQUlZ4I1mug9kN2BO5zm24kWhCEa4R8z9NLYltGwCk8EJRQ1MvXEcK9Z6ls8t3tYjZeQE0kgtr
jWnTq2SlRthiHzvxT6BNWCSLwRhf0YUgE8OGlqKxszJ/GQ//VcN8/lPo2sXV/wqamztrEJOxWoAg
dt3BySjAUCp3XIZi0ETGSWVEgd95IgRN7/tqt9uG7thb/r4unx++axa67WEU3SfM62lCPJ7+WWo1
quvCXCXOEZvPAR3TLAwABYobBab2WDv02x19CagYqkZddUeDYPwkaHjlzyvuqpyoemp2W3IfNbnD
Dc/jT5a5PjGQswh8yGVf5wUDDNdCOJ+zjyKfkWUo47ntSKK6GVJaJjCjiHcVpbyhQpipeE0EsSqj
HiVzasO7hJi2HmfFkY7VQ7ac+84Xry0RWW++xu98NOrziWEd7PSa6kKewJSts0GOvyU/I785NyMc
4gLHYqb1MLLNH+/Iktj0r3X0m2ixHA4tWOxhLI7flKMUuqfZB7dKGCiWCRwZ85qUeiqhCxpWIsJU
R4GR6Z9743/JEjlSj6tJQd0JK7/dCln5FlNdppKiRdLy4aph8p620VOPnivC7PnnqdY4PPuH2QsG
rllscAjbZ2EqmC/2BTxA21Ao8lHPV1NqO+ca45skaqyi8/1/nRq0VXTH7jZF51RBzGoBaI5C3kK3
d3oZMTWYu+z3n+Xr66r01dtfarmCLsbTdsqJ+JHJL06Dp9H1yNakRD199bHKaWD0IxuuND9pwv7R
2c2fJvVHV/QVKB4jkbncgq5//MnTuj64iRV1P/a2RRSV4x2LX4GrPzt8XAn3zoW0IsX+eaDfdkZ6
bofrULnCwfUtpz9YMY5m9nJgOqkr+7+s85Bbuy0ExGNumHRgpkTzZf8Avvu++YpOxKkNdqhKcyBO
QEfPj3B3Yhem+L9HzRXhMB1oWScV+6XpBLC8pixra5X06eiw9eKH9gIz1m7pFsCKhyOqShgPw5Hv
+38ZICYwY9ybcARsQ9yVuVaGCoMskynyXrxIGIG+N98IlaIGZrj+LL6Z7QOZWLSR/DgwBpL4VULJ
FC227618o9IH8iq99/DXXEMluYAMc0jumwy3pEO4wAbLnOrV7zm62dm5KB3PfvlTmJmpZtABKU4D
yWufYHAH8VVhztVJWTDnH1pTRWEX9sz6luPQLdGoQyVWqZY/IATpB19UKa8wBubmbrHNyPVETLyj
dbzlUCEJZSC08CF8Tk8OTHJG1acpT9YTeFw7IP64BgnwcWhFPTCl6ajCWTPwXMIkD2F1FuQUvAVM
AYsfW4xhLj8/gAa7HUkRSRu8mYxz1A7BcQemjE8+e/tbSeoQA94hN/fYommA4GigIp2iyw6btz0D
RC4ZkOPxt8s/U3bz4yJ0JSwAn00RSPb5gnWqFUnH0INsPhgJnh9v4Z+BjWSheyLZvGT95DqclI1u
bMEbOtxA6c9KqJxrhvIND2WWbx2hyx+BzRi/pZETHdT/0OCiLEfLtdIDBB+4DL3M//YD/yhDK8CV
kMhULGmxaDnzt49nhB2InhGbp6U4DRUqn/wsmoMt1sw1J2iO9Fg7552xOIjGLFYXJ4qqh61/X2f7
WTVS+Gay25waaL1e0dy0/QxhwknmBtQqCZAtuJKMqH9UtSecbQyoZMkl0/GLaOVAtdTbKZqZQwPB
fzBan2lzX4B9tc5vX+DQdqn7G/VUn0pypAr1lLUdPDEqtIO8uVGCfVDZ4/DLByYe5bJAPPvBo8kx
BkPDlvbkR1HJNNUbRO11hWr2rKPfO8QEfNY30q+SnQNgdYiy5CIyCsE+sp2iEhvVtmHr7ME6uxaf
LSEQE1IK+p/IUxjboU3v8EFURqdLcTJs4TMOH2tqOhMxD6br1RuI08SCfCXNECjBqYe4/UYSogJA
NXIgUyR5KNYPZZiXEHar8cDUpJf9II4wz10gXxA+cSC/IsrGWm2xnaedNiWmlQdtuLWwFLU738X1
VFvlvuz1GOfWgiaKvOVHU0igV5UkPHWD5crHeWd4z2EmoIA1TJtcEDbFPd7lNuwW/ZAIOrMrriiE
8xeMfoCeE7E2l2lUuC3nQrbK4pW4JaTN2q+qIRdUubh4FPlFr2u7lHHaYlB3CcLtDmyUMORe9Po0
IM5asZFaDsuTeHlUvW/lJi01fyOIKUUS3400qFo/FlLY8tQSd5Mp4F9JCR+rAWcVGnl2yH5vPu46
GAM6uEpbZr5Ah8gUdMxhu8GYUZ3oDcHYpjA0dOPjwl4IH7izsrE+3sS89BG7kWs2Sa0H6MCZI7Qf
GBvrHwYPh8+CoOaeNDdlSq6li3FQ9OurSyV39+F2Zt6omSvB/A5EGedK8vzmQYJP+c0HSwi6OwrD
x0SxJnfbgilMc+l6ZHxXfXaESaECxNhjLqxowhuyp0SVi17PhxySURhpGWJ0JEjM4Ndt15glzM67
6jrGsPBJfDS/+0PhwKXD/ac+Jdl/NXISSaLE+VK4PAb/AqfTVOnaRyIFGAtAAI8FrvzY2mYei+6D
+Lg7IviVU+JmlG/vn93hxCYoHT3hB01D0g3R+usgG7qRRZPXu1rUL3sq9eqAy3Js6+twYDdxPs10
ogk4gq1Pq3IQ5SxGMp5Lftr82P/U5SG3KVc+dKiayfZJ4HrONeT7X3LZ+sWA9N1TxspsY2sVT0hL
4JZo17nXABKYYXfjqF89uMbt+aIO29DRLNV1K4qzRYZ3YKeSM27U/uh5e6R3yzliagVmdAP4afPt
xkpiMQN8cvlHQezme4CP77AvcuY7SnTqJVFqRRNk0Qt+R35rxJxA1kZqmhlOXl4eQORC2zVtLIIA
AWKc6PiVszWVPMGZf3tWR+wllpEMI1tX8TkWODU4zKFOdVFzGLwpVggmSVJF8WF4WDm8BckXB2s3
N3A6tXr+nilr+/KcqS5bCW9qCGZhMpxPC2gneOEbrrAXQLmnsE3FLinIupAu1XPgL0hkgOYFeEec
3PRLEwXK4kJ9lXz9pBLAGX2aiLB1uNLq6GnhQS95YEtLIcGJfe7hE6a9hPuP7MhzlI1L5XQwlmah
lkuHCvjwIGfELQqeIJZAiOTisoaFHInQBpcenq4isJKctP6afq+PYqhMm8bGH4Hw2Uyl86pK9Me2
h2uxD7Hj64jTJwaJJt9ZsIOAvIwgCqzHsdPzVbYs4bv+6XmVDUqVD9Qkv5b0301Eca0/35WjpcGl
EsNDf2cWIk5Wn+JSCdBN0hPl0zwUH4C7ALdmr1CzpjefCqz6hUF/6kr999UC/lgnMYWS+rYHI03V
3x0FMI6hk0p1l7cq2Eme6ucYxKS0/hMjsbfs4hnvoZ6/GrWwN2f7WnHKZZ5GF8PePxKxP8so+pps
/hLrCDUt0v2Y95KWRDBqkxFQlkDg8gVZpbUKFjImTbTlmZ+A/+YolCl4rcJkxnx2UNWGzRdEg42A
08TEwn2m770/+2NNHFqNwPJQnQWe+1i2pbVQuwD9gNAglsm26p4TnWdOruILz+7jLJ8Vt3zAmwNt
VUXXb3cPLB8bvC35oKxnNGYK/MRmRXkCptRc5uK6oVlTPiwg59AE7OpMO1Up8pKV7sFswqEjkk4V
wQa17h/C3c0av5vV4Qy1sEhjubJSvksNDu48/aDPj3dHKeTdZNJF8rqUlU7n74d2Y7IsNP8eIU4B
2WWz3c5WpuAIDOkoqezqLUuRy3lCTcL8SKRoq0yRyqC9qa8Qz12WVBRsTlLYnnxEJOKwdCJO/TGz
h6x2eeOahrGz2DEtwQ+0TKbWbYAiqkorZPxuSXasOT8fjpcqUaEJUHwJfIQJYpvRwIx9C7t0iVon
0gZcgjnR/v/OEvvD+nR2aIOgfAft87JkTAYgFQYDjQ1y58Ur/gvu4jJbssutYvjQp8YtyT/GT8JP
0+M268vgJKwPnclOkdZApgzzPmSGn6EdE8ZixBEpcpXxoMrsPZaOoyUG0Dch9zxQwK7/eieX0rLK
yHQStljcSsZmNz9aHZ1CzA9M3mZb/vYKTHN3vzIFl/YvbGqYUbf+2vA22PrmFEVCQyX5zaWmaRY9
P7TwuAe1AdZwFlZIavzJKQbHot5ecpTwcNoCvOoS2kkRIbPTUDrWE4hf6p6XA6ivWqViNsyyGpLf
7yCXzmPxWrMmFME+rp3VYXTr7ZTLv5ooMw55x+0HnCmYi+OYpiabRltxipr8m99uakOh8zZ7cX56
82GPeYX9BqlUQAh7LDqYU1+Wtt20xNZ3fhemEkQhZc5TOgHoa73u0Az3OX0T045y/dnJ1ibhOPze
qc2ZtA0je0XoIdldRpkuk6z8SHkmdqFqeIIWjB7gCje1cKqgCXo1Si2EX10VPuFw2nYT+ulV8wlY
4FD1q8RRei8Ehsd4KCABRVv29twNvSiBmxwh1r/DA7jjK9hN6/vNddg2WcrcNV9LfCVByirtTDNr
Hyf6sVp4XJcgqD9+4AjnLB/Gx3Smcd/p+e3QaoQYDYq/AqPp9bJq8vCwuiL+hG2zvVa+ZXmYDUAt
z9WhdDK3WuQkxovreYqdo9/clOxabolquB4w/AtzJeLcSWgM9jaNscC3IwoJ1BYAeLuvann8wrZj
31hmRfwiFHdHwfC8H0gYS/aqp4WVk772VYKpSEqqn0KgMJ1z9LZCnLwC8TBE+5m2VRKTwwZZ6m9j
yhM8k9Vt30QW83YxXWiJ8gg0dFjqWnNd68cmce6GSN/7SlB9UMRIFccjBZki4r+ouGAyJJSUiXa1
xob7tZsWCaelQZnkgPB4EGTorSKJP33yhLazHDvdxOn2tsF3SSkmVVAOa9ndK5OcuudzC4vQfJQJ
B6se1TKxYEVexX+e+Zf+mVBvGGSWuGmO0RSFWbxuInOCnzpKg+CzDtJtW6tHyh37dlm4WAducr97
JfjvmPC2vdn5HqRdogqjmsin43pPkEezh6jz1c2jdao9fLWSQRcwvxM4GmzwkZFUC9mm4ilvhX12
Cs08389LuD3IYjqA6C9Wdz51XF1Y9i7iDLv7Io8WPffQT4vU758459Rms+F6AdatbRvwPF+cAzEJ
wuMDNby5Dw9UUOIqCNAOZMLZFGkw8iOmpEdKtGA18QIGIHBwCOoKZ7aEjIFPDnitLTKtDOLc5alb
KbWTf67fgfB6cBzZH5gICL5enCNAGVjVWZmD330dcyD83GT6p1GxcUB6qwopmjcESknlAZ9KDRrI
H3j5ykROPfm2A4Ip9OvcBjzrauNHZX8SMUitu2tbZqP4SxW3+K/EzuhS005ZGFwS1FVODcBgoRn/
XzNwrSC2yyh9ksEg/elDyOEpwa4zNVHGz3yZoy9k0k8JP5OrV9eFM2grETyN2/ZG8bR+IVwMrUj1
EAI/8CB+5t3EDz409/eJ6Y+MboiXL/R6ZOQkTckh9JEYDm8LRWuDZkgVfUqaQcnbTnf8mTYdJRw2
rCxH5BovXBywv8pkJZ2ZWriRWVxn2WYthN4QxFpNosqxrctT3aIvnQTWUac/74d9ZemWFHuUb3xh
SUBTLt0zVTjunRYgSQBcHT3v1EMlIgh35wLVvjqIuzSTBT8m82HOL38pPBFWIUfTyyS5DNNQe3Ob
QT1tn3dWRw8jKE9chCsZaIBM+bQVwobtYA1e3tSbH9iGHxI/I5iScj1bzsuqp6XKWQjOfAfiR9Kw
N/ZECcU27xoeCCKpGxxhHyiU0tnx5IVYFcXfnKpHgJIoVgGgi0oOe84Rudp6mRTcAErUg4ENOZAX
A9kNJ2wypwSZotAUBo8KjCUGxYGLNNb1g0qXbcN5L1itfQGG1sAN6tp75Ozlv9EtVALkMqunvj7u
jo7xmKlT7kkL4JbEPnOOF+OWnn5Hoz/r3RN5z56tDaqmAOYKmURBneuz4IZ2pshFB0Jnh32Dvitp
+1IQI/qxzSCSyGED9QlAlqxzw4DH8krOhOOauuVtrt+V2CXvhN/8h2Rp4eWDkGCO2oCykZaI1fMB
y8LEzK1PNT6Ne+26+kU6KDC03nc+7InSa0VkHTHSzBqRYTlorjY2ocGZXPY0WRYAm21qxCcLyWrQ
0jt8p2wXF9TD1+ay6MEQTEK8KPXCi7gsSAd69eI2xaGwLuN4x7wtkgQTp5usKXXJu0fsilznn43M
E9TQSLBpegCmQHmJFme31BxFu6ugG5GAOOHNaToahHHDSjp/NeSxaeiu9AMRJDZ5eI2XlwzZSAvH
WHGeow1fbxB/SgUy4gqLALX4mF8DJ0K/kA/uGw1pAUL6VD4bL9ue7W9SDjEAqdQLrVjytFXEWSgD
/ycj/fGccmwjxskKINMarXmj684KmHcpRrB03giL0rYHSxokLgq8nJ26GV8vlULKta7kF6kzLiyH
5NjK1cO+5cA1Qyz+cYH8I5UCQA3U69lqk9HtlU3yun25C0pcVcrE5+UHs587c7zkJfYu8C4Zimh9
GYxni4Q9evF5S4DNmp+DuzMjAvikl5ZtrJRePWBbMm3kWTllyDZRVsmvZKG3BNFYEzlCLeOIG75k
SmuM2nEnf+NVWGq1bUHasbcO9rBVR++jMtCQEtPml8x0w1NWlgL3GQtefb5jEjWP/NuQv1nX4c6E
IKyWisgoujGQdi8Q4UirFsG6JFsoapZP4g9BLZEZiIP8ff3Oidgx7ajqhziUfwb9K78LawFNK7H3
JF9fSAWWn8ceCAwU1kSxro1ASO65B/PtWGB17xlq6EwWcdSH3+UvvIGvhhkV/2G9c4HB3bSnObEn
bl/WaxuJe/UAy4e35DbY3rs3AOXJWZYjLb8v7H/OdIKgqZFrwKTp/OKKR2xbmJgSBqGVkoqKO0YZ
zdaeyqGCRxvg+2qu7nQMWRnSSseFZybfMSYUkbX+sszkU+JAF2AVSRww2wmvH71R1pBr0Q071Itl
+0XPPKXWVyfpUalj82rmJ7vC9rVOQdOv/cya9GG7qQVIYkNsLT9qtxj3DBITRhN+96mtBO1ES25Y
ZLgFTCnDnNku82vHbU0yC8/Oj1PnhKnvuAVR/EEDH1qoVFFH8pMFqTfs+CrMvJ8iYVm06bKV5tBl
miJbGid/kWevj239+ATaWQnbyi6xsjTmUFsOqOdYQVrhM4Cw9EiWX406dy5KcaejgA3W/obRB996
bwndmbi0dD6K6sm5SIuJaKy/ZkyAhwc3NruB5hJFxN7N5y7uI6bwBGprs6+xvfc23AmtpzizIdsA
6qdP/GIq3/Nj5UfGOomexHUezuve4iflhUo6fP08IVyx3YsacTReZZCIvw7ZoLJ9BzrP5Su80fsj
oRZmJGemqbR82jGNeGwI2wYfLf9lV/F/iV1L5yfu9jQiY0OcnSbc7uloYHcJOCjdzcVLWIM0QeWA
SGVNvKvwKdsU58Kq+F2BbWhgAc/TaZ98Ea3LAumc/d/+WXeKQfsxMtEQ+qtWaYDmv3x0QSLAaaWw
KKV4KoJ0s4/qxQguqyevvWdJlbZKfzcdGqtAzL9cJPpZMDedqScUX86meweEJNz2YkTo1SOXv+Ql
DlNkCjiT3nRwQ/hEgVzRMorUSjFIRILN4mZvpK5hEDWjx+1A+1oXvqPpIjggidMNNYRLqce3xcaR
CKCi+XE2wookmG+UdbVlL6ZF0EbLOm1G8Lzfn6phnWCd+BDJ5rc7XCSIeaRF7svo7K7HxX/yM7XM
ksB3XU4FH9ycaUUg766Nbrk5czFv5Xe/XE14bQobeJem7C9ul/5k4Qr8A3tmXBJeIYuogQPFoJFS
sDtrBeyYqv0e8S+cjTaucq/dRkQN0rpIXiTjv6UCPHrfDstI7tvuRNN4pwaxp88B3LF2UeC/IhZn
c5T4zKUvqUDy93teuBFMGISKCVS2atKVCB4WYNVXgjUBoFyAZ/l2hdcyRoMABQdlnGMwtC1ZJ42l
Y5UWteBgpembFFNeEdFsvy+BzBk2S6wtIxT3gg6DlEzP6hxGay9BKJpwxhd65ZSCSQfECIqNlXdg
Pq/cDWkXGP4ydjm5gBr5LBDiCQw8BNJ1ZxID8K5iNsqeKEOz+AvxWHFOq5gyugXPnU1A8iZ03Imm
s0j5uKTa3n4U7d54TRh4+ISCeJ3poxL32XsFlPORgHH6tka1PBCrYv80wEl8VTIiV8pLNzR/e9mU
/KqiIWF8K32gg0Xbr1Ew1L4tNxFWHs7mRFKMOHXnJGgISuRFWFg0CqW/r+vUd9OwB8nOTeT/shB7
VTIpp+QT4RscFz30xC+JYuweG8ggWTa23pHh9RnAFO3wpopyY/hNC3XQaCVQzRjqbT4q24tjTJzJ
BlDuybTwDRbWiWkfJpjRNkL3zjfcvCFCqpBA5gsP4/rjpFBz2Jo510uCUUgHJAC2hdHQKvKJax35
9KSgHUivMnUpSy4cFvSuicLe87/UApiWn2M9B5Z+6oUuDwYAVIJR9I1591Z8iqLgFtDLVIi29yaZ
lpvLGeW0EcekzdTqm5Famv2aYPY5XqHDpCR3bWUGbZm/TdWneMYNXdxsjn4PoQQ8frd33Z71UggU
qnMqg1g6rZxOKB2s5spvDAmDeFsl0aJDk9rAFyKbMoFFCS+9d8pVMNSC3jeXdupKMhOHVRl8fgUV
eAVI946IfRsV4JoCWr3XytLbKqsuLnmHYS/+TsKdEeuZ+99X/bbWA/GzmWml9RCVe3pq5aCfKDay
YyOH1MiTexg2xWjFlcbZ1iKRfmGlAI6T68BvW5merONBhCPic8Pl3V5TeW1rMncHc3CWEPfAjOap
e4BXJaj87mgOfuB4/Nb5t9hqxj8erhDZhGEz0iPRqdl6jbDYAt0qKN4/uvTJrBjkJC8Wp2pM2FBn
hfIs2bdYoPXMyMDqpTvXd7EYk91F3zYFDnT+8rIIEzQBXooBYoN+3ks5D0Gof0MlaIG77UpA0E32
nBkLlFyTnjcKDn3hWj89x9SgK3HvD0GYfwaU/cGhpnHjddqSwx8nhK0+lKegBbsYJAsTqAq9F0Kg
4UfAng3dp0/uRSx82hQvGfK3aV1PEMAKyVJmGZ7CYZr8roYQ5a9wwp/kmcPY1cQvLYkmCTP8/Srt
cnBR18nJ0sRNh8Cx6sUkdrpPU/NNbC3hg0gYog6GqBFX91fOrJkYqYANMsrHz6U/BYsFNJuQYj8A
YHHnMRgRdw0ODsc03Na+h+mkT98/yROhVGAEF7GsXxiFAkfFGGBDbiwlU3rIwIsts/xsKEFo7jUs
btsjfTSK7gyxYwmEU5ygKoOwh3eNhBkWYnk5M8g732EW+NQCt7Pr3+uGc7WajxsvpdOlIRB1lUPq
+NORhHkArve9nRSlmOk1dzymi00yHAmb20lWYlwqe4zq6LGuzKkf4g+ZROgaX9w0MpGn4Z8fMEGx
Ff11pf0f7kXsEpofjJD3pKARjVtECvCBJW2IwKs2PNTIXr6Z60G+nF6ZCgRiNXtgyBE9i1ZwvXel
HT73t2CY9bBKgWUMn+AdAHJuNww3foBXtM5tyOLTzgD63Kwpz9I+/ylFlRo+vnj9R5LcBm+vAtFq
1v6xC8cpbIdPwWBNttp3D+qAj/vgfFjauUoSdurIOIFmD6jZ33tR6DDFVtseGxq7S1IRD713dzAE
Dx+1VeuTl79CFGthw01GU4vUyKTCH5SkAhok4Vf3hynIRwkrpwtGCMpsSWCxpBr4vfS0Hc6qwo4r
ZbVpmPu6LKVbIh+eyR9lOTApuoazoG7WhW3bKXSndwMsMptsw/xRvxOhk+NO8iEIqH7bRbfKIAIz
NL6W6i/0jfHH0fyd+YKLvlRMutDCaFv4gw9ZIhgrEPLYXx0XbOGljpPbBlSFLxSyNtXd0y/N83OC
xRoFmzsB5wajwQGGSgdYeXo7wHIxkX289J47YnQhePIEBISOvs2ivXLEDELwECTRP8Clf6pj5+J7
kcO50mONDxezrjYhAuHDjZ11n61FNWWwiwC5uDKlNO6eM/R1/oHNG/S87oQcUIdC1XkERIZkzedb
gOTS0hVbfndG/bEDEfWaDJSFEBoAeXyWxUvGr6quA34vG9gop/etq7UY1t3NuwQoOE3OhycMmvFi
WxKJqUHPgaIuykswhoz4UPVrn0HKk2m7KzvBUbux1FV2Tx6bx2OWRE9lkQdtdAqd68a5atdny9sx
CWI1Ouqf090lQYJh0WSR0MASjsvguP/R7lz6aswRtU3qRsD8Bkhm1SHU1mzacwfRAfzXwg/GhdHH
1YESJa8Q9/bw9/RC3MNZ3rk0oRWt7EPNEebp9H5luZgF4t9ch2j/QlgWCotKJ3uhhfHTchoANNMp
vV51rMLG5b0oH6ahiw2ZfOOI2DsRwtZZvL37fu9EnpH+gmRYGwTpB3vvV5zhgZyloXgdJCQzDByz
OvJii7w9fvS/jmtK8bmRPlUtSocO5OChG3/uSSPzP+COtrHt6GmIb1FtZfcmqQzWw4+/tDl2QXhL
Y/hsxLINhBzFweOYHqTsNe5/ie5On3TsqdmfnnffR3HadCEHjqhr7KIGkZRWwVvklYPH6BNtGak4
UJoIRCizobV+27nMy95OEVM3ZL9ZoxFtw2vJ2eHu719c7EkfeUin5CEhvR3k1vVoZFUZgp+pU0i6
fecWKJNzhsmdhN0ExXRKqKdHdspNWPq1FGVcXJViCAS5OHhgEu2jr8eQ7ERDCsNyb0TuFv4WlTIt
EQkFpqOC+EzwL5srom1vOuQD6D/w/zSPDFkeIgU9DXOJdrH8z7v/yARWIR+4D+5CHQR0yldjQIgg
ewRrEMLNi37qnvsoXUI7+WIX+qnZrYzK5vd4QWDc/8IcBKx7Du/NbebLWCUg4KsVDaC/XtOZrFvk
TNZT33lf/hSYXr5Kz80lAbqpx2Euht4MONyRnVuFwpXGImnFCTkFv1r25u7LNg7CfYrY5lMZ5O2M
TzO0/Sarj5Fcd1xwcC5xArtHqAFUfn2gtG9aRDzGf+H2LDXoTwY2r70qQzaPObygntDYINFAKXfT
t2fuIB135DWtYrMIM54WmMpxTdVwCCNBpPhlR+oNYNs56W27p4qPVefOjQIamrLa543h9TBLTJ37
258VLR1X4zy+vT0KTy14Rk9W8U0qgezeaiZFlOoFm9YC1ueTRzjDhC6EAHDibrXOiZNIvYMQOOq3
G4Q5X2Lb9xqxe54IieU/4CzT2doyWbWHjz9IOJ7zGvBF2whJqeq1Ox5uSTq7ixn5uiVKjYcQAH+y
KkOQF7JAsiag/pzBRMkPB7ctkSXKzY6lU5711ztNuO/0I6rRE00VlvcWjaEB2z9xjMQUv0qjiDXT
X3SnvIKtXxnxCrdyyRkjzz0Er5LHLZemFA1fp5ib/e9B8U/uC1OAqRNLbsci7Cgxi97SA7SX8chV
1439ZRGO5XQ+kbCeBHwhz3pNq0z1r4v2WX9L8aesWgiOdmTK0KXLwm+9CQjBq0dxcYq4FXUhQhZC
S3pW5Nj3P+Y8L9ooC2no7XIz6+YIT/RYPsVmwWw8fAdtsxJ0J06so4uXM7Gy0+9MidupMxVkfUIn
XvtuEc2BezEoDMaXvk3DgzvGK1C/E2JBLBtlZ57xlh7Z/P/nrJUt1kQ1KJPkw2rSivtct3uA/8Ix
+lhuyiKK251pwtpja0eGb1+nPIsfgi9/hnyRdZFql04U1n/Wq3PXVVPi3R192cVohq/n+WzStIf4
XY+xSqlVYVQ5QwGunfikzMvCyFG3Sqzoe7kBZFVnylxHss8hKnKU3Jl5+OQ2AhnXglbCdt5IX6kr
c8qTHm9Zyq6LX+jA9ABXZ8gBXXdnJ7ZyUesulru9ywEdw0FJIsbXpybrkIreCFeunnlC7KZrMsp6
vuTK/j8g4+ROfcm7D4ZPEqzDYWxtCConnx03WifT3u4MLWFlQAjbHhZB1IeN7Kx/qALfJrLA79Ks
UVn3ZH0g1nKMXtQmT8FmrF9+C/wAXtxwmQQBQLqqGgEfU/YSduoi6Mqf0mdKKCEbliDCJaWd0oyz
AK1GX4F3CdFkyZMC0vuQBn6tKwptxLnrCnxtASFyhhMgVF4EMwmH8bUzfdFK3+s7M4NMZNuasUG4
3jXl90QEMb+iIJKGziNlWpJJPUAkYiWF3a9CLEqk47xtP70MlTppOTvC5t0nxJTI1StejKp5kX3X
mJaLoyHTziGwr66stwQwK4Lc7IeTU4B64JM3eZVD6EcUFGQufP0iKUgGjCGCKxQupZXTX6M+sf/S
0gyFM6Ez6LcE58dng0ySsDk1390KYLNPbMEaGA9QrHAKSWK8/OGmEzHuyGYtchL5jHFTGlaCfFQQ
fxH0V49i/JcDEngLNNYnLwouWJFCMFM191iYgCVR5wI+/9zXaZxBF0tXCN3PmTbqmJFG8t2lzdCn
XELAXWI3FM+JQ1jmuOK/hn59YtlFElQ3QI5Nkp9rW2d9juy0qfNnB6BCLc+GpJPyGW3WZheMKHly
/OXfFlr2Ps+zLtqwav9FqsINHQ0UyJ2B3gtfQy2dCwJfi5v1/viGBYZSwdnNJdcer5aNLJb35qVa
mS2FW7L+hQ6HYQHVI3K+l82SCGaFggRrWxSEFZOcr2Tv4xnDTSKr1vmcyl5b6seDW/1VGTEWM9FC
c79Fiu+aFr4MA6OlAV/6qjbndpVf0SfZ6B5BoUTd6ypKYBoA6DbcIGd5to8f+SlbawzkTJ32LfHa
A8bkMMO5ShZgGACUeTBOoHVu9zBSqqOjv1gufu/icistHKTj9UeMVrgnajBV/ReWt4SsyS+77i9E
5cOMjSht1IQq6ZZU2+437Ra5S9oHcmrSTlxbJ3qMDP6RPNJvNAzoV60Ky5i48YxL4jt8vlEVW0X2
LGAiFnFoz/wdkotxFr/H5Dd1oUO0Rb1Z0Xu24yoHEMIGVqSgarACdl+i2LYSysgbN54ebUzrXBQu
LXT2LdsqoiONZsnavQKY+PqCxRp7waBJtanfIKsQTb5NtDLmlI1Ur6VBkMKWXekWI1HGDiD4TRt/
NatgSuxcwL4zJCt+dUXYUHN1nBn5CQ2st9yWIM5lXPX3xHjF9egZzOryfCEmuNIMKW7uyDr+EiEB
gpTrgPyN17+fGZhYNOQQIXC70Pggkda2BE/TFZ0vy/i/9g/Xa+LDACWv5ld4/5+OTQdYadYoXwPQ
T1wRkviFFpcW/VFOmehO8te5KaUugOCwm57VLXOcIS6t3foqsS3gWO3hLjyuO9MLN0kch/fKRyLG
LJwSM9vZkPiUofOiLifvKJw8aRlf5B/mrFmNFk9mmwMmZTxzQLoaAPLDbbPtsFvJULKNzhtKSDDn
uBw6RjoR3QwoNsC4BrPin+gWk/84LmUffJYF51dR8Xbb7f2PX67yXtg2a3zPnWk6pd1eeahk+Qxc
DsqWz/fVXVBQ3Nswu6v217LAKQ+zgRX6aD9YICc+AG9Ng3QbJSVCcLqRLkh/mmifjR0S95/3hld8
ZTPMFoQul52eVphKMUwZFwPLGjNaoROlxX/rjCFHs3x6yUG0SL5tdvuB4+91R30G5pjIn3eM8bZE
kws11tfjT11kS3I/Q6Ti8D5cM9fQd7JeDT4Eends3AYmy1Dt+fyUlGuYXqKwQ6YMQrqrADGXfceD
H4ciGcnKX/a3hXxSIWy4WRrgE0wHvjVwX6NfcpEhOO4pFYVuNOedbhRFDEcJKqlztaG8BtqwHRz6
Q17SfnJ06HcsxoK446f+VoJUX+ONbrDinBtouspfmhIXxIIzo0IFflNyzzcXtcDVIAQQmewkY8X5
7qTTFF/AyrszaTtpeLZaZSkSvyHPbZPp/YqjHQ53RkaqxzR6yIodHTFdRD29/jW/B7wnewq1mJRD
KV6UF6p+q+OaHVIgwP8gr4oInjbmjyYQRzSyZFuJSmMR14rjwxkEcGf3FZjgFeRG0I0EUCWaP2Ps
rJ5S4n8tFiBJVQR6bUldY7F6ysJZ3+ripDQISSYuW1izTuinNxJ/hvikVWmHbMa1rdd7z1TdpNTV
bigppAGgnf4LUv4m5eSVLctNHeHePKIyL+BloYUw2cnsESgd+3QoHcW7q8m0+Svh1V9MIZp07yFU
5P1pGOShXd8hY88eJaoId+kfE/S3aq59qZ69Qnn09GmeITa+62erOCkFvluOVipS3Ja9GU7grc62
ecBrth8vA8w7HHgGoWTtNbvC72gflj2utzCoSaW4sOS26F8Ylrd12jRRvpVSU9Wzj6FbBiK7H4TS
AipiSuZTURd+NmyMKBiVO2lK/C2NFPZV4FfQ+PpdOLvgPnZYIMwUUs8IHG+K+o/fuNsigJk764Cx
A/MrqOTyGAB+EiY7971ncaBjI/fdXrVvvnoo3eDrrByW620Mvc30l6HomQ2BvV1E5oLU3874HDwy
mQMIfgcpmLC4uaqGFHGagEswFyQZkvv4Mg3bS/4G0nH4Yd4ZgUPQ32l+hpl/aD7ATf2+b1yvLWt9
+Ao26Ve2geKXFMYDwpORjwUqzkn6aSa1rUgi0M+N42fFWZUWsdbp0IhO4+c4E0DanOvk+8xA/1iT
7Azqf8vzZTRdhv11MwzXVQO6frALRpbMfbynPSitQv0hBtaVw34sdBDjrRJiuqnhHcrJewJylVEE
51gP33ipW1TXBk/nUXtviF6CuY1w0AbX0KDBe/uR039wTpUjrAmuXTfI+9kezV4eQozCZ0WE93DX
+oFHsvjUJ0HF7eZ1KpkYOKYkDTDk3bIhNgeZpcL+7S2AAyYkaTW9Rp7CqNnHIdu1dzoLN0obv9b2
pQXj1b6Lf95eBAdKMioyfO0NPTdP5aNBNXeBGL0Y9eAYdHnJnWq5k15HRwCxh9h6/I14OntHts6k
tc4bXgQLVBuzX6R745nzaSVNvRz1e3Bct0BlKADzMsqUK/3K+LTvCjYDFowNI+4dE/bMhU+TLxCM
2PM1qMgZVKpKh+zvNqkTA75jzsV0Hkh4CT13UQ3cu+WjnG1FunKG0UlpxgU8t8tYxA+U/Yyokl8c
Ly7TCvgL/6dCdm8O1gc7a+e8W+WAQ5gXO/wACtaJGLZtdX8/A9yXCMWVCbgJhk2jw6WO97Yi+GgW
xFrVcYysm1+eUdmgoKrVpkQlOAVR7CkZcr0LfhcG23cWC+QuM0mXXgJotF0MqKPq6Z6w/dgnS2+s
NwtO8gt/nKr7Hvqjwp0ztXpnUMzgn9o8kRzeLefxq/qaN5idtidrbrR+PAumNxrIGucmywLpp/0x
tuZGdjZcGWsQUqszU/YtcIJZtZjSatBThJsoZgwNcv8jIdIAihbgX8BU16n02w0Voul5wWxJbHwa
Sccicwro8k1337YVBLaJc7XWJxNC7AisjYE19LYe+h6vJWIbQ0ON9k0pE4tCYCEfJCmyT55p0S6+
Th3ZTO8CDtT3/n2L0i/paluWJEDDMfRq8eQHhkmcWiYI0rZeZyJHKuZFhawhGSjOWOYFR4LNqumv
nxVVtcfx/CI8J0tRiwcqPDVLTQywi03g4VGonZGUKeFjPpE8Nlz6pdjnfQJAheAN6YQwGQHKy4nm
DLLbuWBawz1ZC2FH/WxVXxN4FtUoMPAXU9Ob4b9iX1NrwSGv7Cc9O5rsFeQtxxnSAkCVMQFVbEgI
q4jYzjnKh9UZiCTMzr1Bm3yEps7UhBxujRwZjzCSLgw21S3wMeUQ0XgdptQl2zl/VfM2f/1jYTTW
0aqXnTKV4er5PhogT/zNBRqIzTLYN/3UEGnat070DCELsbyr2GtQtAGUsf9Yq3EZ5P15uaafarMA
QhsuFXrwRgT/y1H2rWR6W2lc7pqEPciWcgqBlfS2x9GcnKoRAD4dD4Xjs85Ph6P5ZpUVDLi06150
LGtQyW1fN9y38z8c4CPHm+4IFK0hHjBz1Bw48fl7RjrBPRImwBwxNMKlMulUBURiSUu4KnTnKWQN
CqVlRdQTeA7Jy0KXMWBGVPYtOd7mk2MmSRdVmaiqtU6K6k3RI4n839nZYf0jywBz6wuTrbayB1qE
CZGNp5g9qwL11bS8aZbnlsTaIMIsdqUOCu56GTTlA6AO8zwZyNfI8JdKPkndjm6YKrv6gARf3p8t
rlcNi03Lqo71r0PjB3EQ5Kgou41ZvQLFWa0M6sTuPKSsEho7k+gV5c7T285QIJjzxCujA7VPA56H
P1Pkcjb5vmWTQiMjBGxDbPE2+xG13t4dsRL0q9IALns7fC9Lf9leOkLALQ5deNnLp0hCXAFdtHOf
R4rpvlcIHjF9mqCBWOYZ9ewJ9lRa/WPP7/ay9LM4AKcxefTE+458B5njI4lZ+ghjo+SGtykmABL8
TnrXWcHT4CfYU2CoqxApzRu9n1xTpiuBvnjGo6L7rGzv15R2w6EBJJJYQfesZinG+6nZOIoL28KQ
/f5UxWXeThFO86js1yv2tA0j8ds+QFf8ZdSnRTILWzPOsUg1zf+szkZg+sfieErhYem5vuKYvC1g
4CVy2ut8KcOufd1V76xXLTK10t5uMp0ieqbEgXNAuC0QtPXeOBrhiBUP3CLLDNUesW3MXsSrEpjw
2UD7Esg/T4fLC/2U8BA70n+txgafCg7BXFzIW+AmIvm4N1HVAsufEh2hAkYxD4eqtg4Fdcyxw91m
nCIHEYK7/MMh6BvsAl2p7qC0F/rAiuofcmfn7dggtuwC5zLTunBLNj1NO5VTFfqHs++l9JkLOgIT
UispeWEwNwpmT0Wp0/3ZFZxDRnDE7UsxEq/WV9SqLAz4PAt0BcF/dJozj9DyOjnyuhYsdBk+yDFA
I5RqccuhNN8TDYEzp1nJzlPv0OAJQppyjWATgLm8qsMeCeXjOs74UUanYJRcOfRzVLgPIPojfMjI
2IcGPDYw+ifMDTkFhenMb9+sLCKjzyTJQBNLz/4iGI+ryaO6ur2dZl3PTBSGQbjB6BJkEF5YIkKB
UDvqFyw3VDlYRz/q2t5c7JDQ8e1NRDrr4UoVHLUeSbkQCkOh7TEyutqIxG6vK67tkAoNQbQs29GX
Czo/X7GjxyPuOEUXC833KmmZ+EV56Q1mDEx8n/qzO29ZeQIAoVHoTzpTNwcc0MK4O8fZnkofn6Bl
bz8m0JHnCzCYZssj35LNu+KSBtyWnYS0RZQz6O/kc+3aPAv2yeRvYKuDy/sX+jHJrW6xO/6JBnze
4F9W/WhxjD/yuXMGKdzofXSfu6AY8gfwIDvkc2gx3A/BwD8sYt1cauIDDAW6P0PauGIGIinviBeV
ailhBn5RoDL7nmjQkCHH/b8MM5XaNzNCq2+kq+i6ulIBW7pD3VBTrE24lkXuYZ7BZOdlyMXRf9qs
TIRkw8P8HlxDcCvwe6cRWjZNH95lTBe+ZhLzOsxsafMHIc5hj34IqI34a22CnEdgsFhy/wwZKE7O
+vsw3F3DY4qcvg6M4XThhwvi8qaK8SAQM69MEU4fczN6LHm6ZTyVgZH3TOTaPdpycHwsf62eqJMR
0lkkZ3sfrfqhVHBtTuwe8S5xTI1HbYBCFQMK3iDz2HgQmtmUm2t5aNdjQ47pOt4MJ/rkpqd/LUnU
h0RoCCWA1sl0Mji3QZmvOq6jPGPKi4tuAfR8lI84JKhm1C4cR6Wvd+xXJSfHiaxL1qOsdDAMHZEy
80FThYlYj7zmuvdcN8uV0T1cJmoZZX3AIRO/JnD3MGq54A69GCFfLYvWGiVW5YXiRWNlpjfmY35D
2F6i57cKm+eFx2ibzpuDEBs/Gh97sZg5mVhsrz7I8BHPCKbYX1snP8T5YRyIujqBCF5qXGKGy3GS
K5p5I7y5NupEwdTrrkXoG6VFvAq638oYIwyyTn/1X5qGnIIElWnFOTx5hJ6vz+Vkn1VM4Ury/XhO
WR2YjrQ84Bn48PlLb63z2/pj6aBEWaUnon593v4YPWesmI/qeSPWKaEHNUVked0OfGW+l/w60jm0
dHF+PNUTMNbaoEFHws1X2HxUPsrw5feWNQ+qKF+y8gR/dGi8qfqoJ1xRyCDq7oWfcDSwg1E2CK3R
td3RWyCeFnH6H0OKtf1P2gLeVXHTUpoAxFyIGKpmYWGtsNQg6OJoqvroQhv9mKMHt8QY/rGnUygc
wgSp4a4y5SgHceBiXJFT1hF8fQMn+4XbS07noVtrd3fcdzx52JBlUaaymjV1zCIw3UQD0GQWPMDR
6RIhiqz3lnWyOu9sIhOAlHLK7LJXdN4TEa0KmvtuzOOvbF3hTD0xqN4NVCMT7KbuzJK01ITUnCjN
W6u5L+a6tO2Vh1D6ILh+6SvfeCGGhnEZelkMsR++Nqg2hOR5v/4rqNDKEX9wndVs3iVhpfW+rF5U
u6LYqFTSublGNxEFlfmnEv0WxrCn4C44Y+DqczsO/f2oO0N4vUIYCUs0gNKZyGg/XQBh0zNQckzG
SnQuwK+L94klKqGV7kMqgGCwVv/7kME4NIEOpCW6aGuQvzUnDxjSc0ogkA9FCBWEQ83qA9BfaWwW
gZREgSKeB7RSWHQ5Yy5pfn/uOKiKPLDGRCdxsdliH4+PlKhtpjLkrjMcI4SnQYmNEF2cFzw5BZGG
QpDJOZ4TZVeh2iD4mnlQ64Ub0hDW8HkbBYqdVCPxEqXh1nlit55XyN7hPPSf72Zub4ilpV0nYS1I
I0YW/haCS75ibQpL7PMuKGQoD16/yzu9LRYOeDDH2mN1T3UZp/5a+4NiRMgPz4Ak9tS4X0m3u5gt
qC5QwxyDVcUudpzx/yXZkLLH7QdTRNQBN5shyU5tsMWrta3YMNiNebPXjuqjD5kJilpRt0bvqMzv
drSer/OKzGjiE5DSe50Mxd32a8TIq/lTSP9wOzT/i3+DbQWYV2FjbJvvx6Vss2BHilLc4Z52Qt3b
nTDrreqRFUYCetms/kHC9r9nG3aHXQ4ES1bGPHMeyq79E2zCoXVZcFcZU54BDln1gZRGYzODa9K9
O01GusDMrC/wE4oS0w62mjMY0Z2gxNfBz+ScSYvz0hWw4ttvvdyB6XvK6takg5Ro6VBW+rHqEh/D
4/j1CpDdpBMXPk5WOeCn97z9175j3RdaRAUMYB+dAT+/c95Q3e3RuAaEP9iwPhvhtxIHPTVaOdKQ
c0l5uiYr2Xpv7GHby2UVhVXDqQLVaLX14kCkmNO0roNLzytGsEj1QgVQb5V3dqPQ7Am70k9iiqIX
0Jqku9HBsNZu5bKJAyMNljsjkroXh26alXbxsjpH1NUd0OwP5MJDrjWhmHDWhiyUo45s5nL4gxud
BjtbE0r1DE9umKDsUhIcobdBuITuedVn0tL/tm6lngKRv3ajpPyd8LxweeXrz8AFwwsST5DMZkwO
gHci21DdEBWzEbL2d/9995R7jZ1JXCtIoFK0b+bJAPzFDZ6WIKJp22kU5uUaDUMQIhyMWSHL7bBs
cljnK2q2Am7IANg8uYb/yb7LNAwsDWqVL7JRzT5nHkppVv9enZWY5GWnVjALO1GcSgkuKGSsW0FK
BAVPDvySS/BUrylrXuFSPwlGfD5Enr/cI6QxWpV2pgXAj6N+XiHOwLIHHecnDp9LlQKHbIj9q+8N
AdinR55ATFDF4scwgyiEQ24ep8R01y+lCsRE3i1Sjv6XslatLV8wEF5mtKSkpI2kmWryAYm3N5jC
o+vWBojgX6leNC/LG9EXL1vp8l1DFUMMMrC/4W7ZjAG0IAm8ENMU7/TbCALOnQXFfqSkiH3eKIyc
jds2hGOFLKYtopxvMM5TXltHryyOxV+7j2opez5WMVZXIBWJcc32XxsAM4NWp8v4y9SvZm7gvpe6
6/SsJRyOYziX0G+X+ZnSOtni18KxhpumOa7kfzJWsjpvTtdYrBabEi9qKGneqrRgBYOlAGy0eXg9
FgeXBjDWX3ReOgpU42s6oRd+iw60/25x6v/e3f806/o7XFJDNQjjnt+9bnkYmlQNjXja4Y/uzG6Y
bxyC3Kq/vwAL9DEzZdcrlVEtx16b3+J2wbCcdcBnql8iNK4NYG7dft15NxamVd2dahzxj4371lsT
s+QWDtSwyHObYVGTgiON2rG/t8ioiC/JrkCs7xtje6FrKTGIyuCHNOZ7iMRMoA9IvmfCCo549h0e
qyj9Je1wDv5kP+w4BvJqwQ+9mopahhl5NmFYwINMYD3f4079XKqie3q9CUY4gcRz1QMa/6sN6mF/
EkwnqsOgo4fJ1gRTFtIY6mkGTQbuZmA7y4zVOb1mnNIYRs74vAUTLnfi6HH0RwzYupQgMsh5Fah1
mn01cllf5uWdhAO25ZOz6VAVq+Y+gnxRkwGynPTu0Jbh3NdGzeeCIQdaoUySyKHE5mh1TX/VhTp0
ErffR8CTww9k2bXc+36UbA3VNfw79GJ+OZXpafoPgDezcme76bK0+V2XOv1jy2SDF83VWBfE+tI1
3N9t6qSxDtNIQj09iscXG2HMXisr417iwA+7+NghC9HZ96iUVzSsQq3NnZRF2/riPuQ2ifn57Bpy
54aL/6RCNeSpHxoLyfkxI7efZEJXM6IgHzYdUTWPGPOerXvDwFndtJhfclJLM9ls1gaE7kc0U0dj
NRSCMfHxjPDFHf6xW77zXsWg6JCV2HyupaCKIG946iocLEKLzr6DjvEeKPWD/IVYaURrluGdWlja
eLcWDw3TpXu3PencBe+mN+JLWPZYVnyODqsaeXXfc6QsJea59y3PMjlAgfzkAReX4ttyI7ls9WTZ
J6qgNtPnJ8iYsoBzGAYSYXK8crGNcLxFrvM3dFYg+cMETEZWYlgIx732mt/wBmAmtD5zjmgpgxpH
kl4vw0mTko2ap+2we0gOw0SdhSNLEwNIDg35CWKIM5328LZxR3gmxU1PGzVNsze8oGtPmg5/7Csz
ygNKzt8UFwgvVkYARZUMeAzgM7SE4fFUlyc6XYtBfLqGpouao+b0j8oNtrIIgJSPAPkSGzALXMzz
KQMlzeU9AU1ngJYCWS82dIWOdTWJqYXCPl2PEOxKhzXuXjCWFFZ1rINrvpjvyJkCY4ghQ61E3qpd
yLrFpAVKOszZYiOAzklsvEXPm3COMuE6kHpDMbbYCvZ/D3r8yjv9t3wKxmPZA0TkvS6mY8Nv7xvh
JkZN/+a85enoxsFkOORyVwgRWEfSe8z1v8NVtcBbgbn+p65g4YnRKRCF+HvjXuwf4lbQO6hhys1T
C4KJepLKlflIMVA5j4+DKOfCwudlC6LKDfUB38gaSn79bdxNj1q3o1/f1keWEEA3oeQ9rrFQxPJm
WtaE7cavg07gRL3URFpivYPbYs5gMbgS3d3BIau8ffCOwIArqdS6ubi8A0Wv/Ve4qcJ+aMJU+rnY
KsTAL5Bv7ImoAMB7qoP1rfvY5jtJKMw55dzaoxKKzkeElmFO9ubVpOg3noLN6IJYU59wTB4XMU7F
DYW+/tdgo1Nh/RMy4vo7z7ilUGYoF9ShRf2Gbo4DQBVMi3sbpTZ9jxR5wKK++xCYi8qgH6503sXU
yZEjfGUgivJZu9pe+b0k2q2QYq8XDOFFgobMXeLaLMsuxYuPy8X5EHyGq+cJuchTyTUneJTk81Uh
ies0485WfarY9FeiSAinxmsZnoMY0sNNxxgbjd8tNp7rkmO5sj9R9a4Pbb7Mm9ls7J7rynEpX/Qq
5kwWuxGDWnWhTXynUFFhu1HBJV7Gu9lPt/YB2v1R2u/QqtyFEEJTlVJwNM/a7q1QVPUdW1drk4Ov
b7q40tPxxx2xwjDOL6kHhWJzIQl/9fKAEgp80jgXVjzOLF1fRVXumaNV3fUBMEKPBDfVObkVfOnD
Bq+A4kikisAxKZrWWHdmKJo3wvOzMwyZu/7AlWn+4hXaBFWBbKfZmtTaLZBR/WdUV2uWravfBT3F
tZ4OgZ3hlpizdQ7bNUknQMJCdcj1DvBZng86SG6fO2qcoMpwk6VMgyw4W4RCxP0z7PaSv1RlBGPn
JT7kmdZYV51hRp4pvlmc9+CPOXHN9bLYt+rcett2tQv86zW+Pn/lXvyZhll5huI3UzzJOqoiAkRM
rtu+5wUhCT1pchcvZDqlQw72loAN5FRBSvPYlQnpv67N4RUTYi+Zo6L7hXTn/AWbY3AZgD9BD0Ns
RwwnNU2vHg9W/P2S8rwck0+fPTnosNZy41s6txJODDPMJj356LKIS4ELUF8JfrUcReLZQuDV6c60
texBrJnAqq9HL7skoLkFAXEkk0jvAXb1vAF2/AO6TlwMn/WQ0y7SienHnsSc75CfZ9XPKk2vzv46
OuHOHK9J058AGQrLrvpxgN0vcjUHxgZkl2k3+iRlZ/Xjs1EM8riHJofyj0Xza8jpEqFpGzRTnkIT
WA9aCpEPS2JwDpFGoY4aEMeVWIAq7Xt/W7BioiLOgKunGjB3UnRmZ3jh0+/9dPVvIFbd/Dt1N4j2
2FBcy6ga3+rr/6dY3Ssw4IoWN6XkRlidh4zgcAc92XWQo/sFDJ9XdE6EP6AxEUTdlE7H345odJoX
IaYkwdHycbxssJeuz1IO8gbXOoq6HXwbGkhMzzLa8vREjDKX1NQheTD7efE0r8D4O2tNiaIm+4yO
abVV94UXA/ZXCBMBRR4xUv9ZPXlN5xs0MnMkbGBI1hohvZNDlru9/5alScqxgpddAF85tqJMSNLb
OsOylrkx/ilqksjAvLHlVU4dPjW0CsRegyoI6Jt82dU3FSWdQ/weyapw9b3kg49N+c3VJ+Vp9JTA
+l5Qp503yo3SgdjrZaKgxkk4m2vZAPnXmTiJ56jQcBpcIzp958UOR83DZJmRNEjAanWxqQOBvgQA
c/lzAKRUDdjhzpJqTx50Ztx2NKADTJli5RFumQbEQCeVJQuK8ZStW4A+90r29ZQ5asyn7GmnqOan
2LyWC82qflZfOf2tQt4sILlwzg1+uSRKVBkbB2IONvaUH8MXSWaQMb6D0PyIkQMCx7h+Pz8nXN4y
A7cEoprUeu8PE05vdsOgLMCLCSQ+t4qSZyyBJhVSIV0oghRijolYF3EpIwLzId5nnDGeSbD1bMr2
80pAIviJr9Y/TWrRQkAeG3t16m/oTfaMKsX3VLIt+3+qBfOQfuxD3uxwaHqRHJ+8Hv9xOOIWI5ax
Kc/vgTJ9Umbzg9Rspuz6odFr2kyVZE/McZy7Dk94T4Fq0q4Y0y0RknwOXVU6ssb9ODC4vbqyTKKy
GEZUyqn81ZQGiOfPTlx4fDanKe6Y8qv0FqZcOTXzLx4VmWKKOFTHsh2r8xovk1xDWlelG40dOGoo
6ErgKgGaPF4QDXu83hvzQjMDNHi1dVK3VPaNbN+DODddT7pJUuPcSUVSJ+X40b6T1aHe9s3mIOe/
VGEU83/bmwvfLsu2oqFpRomhBinYxSU+l4F7wLHChnXu6DoHQdSoX1GRnfSL6+DiLjz9lH0q8ZYk
4VsZDFPNZjXWeeCFkwqAFJIQs6BU1zA7DxKVFBQTNd6Qe5YiXvu1xzECvEyIzQhtnLB8F6TdIa9U
AA3y0Pa192eTbUPhcSZngGh1+0uXXjaDBxV41xX7OPx7ObncK+qaqvOmk7q/hAnx1CsWjUPilkMq
wQJKQxwy4pbBUgRq6iD4XpmFCxh1BVC7JekUnOS9MsuK1T7s2qKM6qhJMzM7hWR7KFZcMbd38pTC
V6LytKSfTRvt74ucYWQ56UIemW2u5U1VokZBK1svLkcEj7yy81f/CJyC/WblBY9NQxDETzajJ+e3
d8HlF4sdwAcojuPAC3rX8/haE78RfSM/dPSVM6eFAlSmIXqLuD8r5E9SQy0Yyk3LIT1d+KJU5tMV
75UeQqmw87Xz4umZQplbEYVDzyQZGY6Q1laYhBYrckDHBk84goqWTWLQsc2p4yOJaorViKLB6F5z
2mHOhHeil5WXZjoi6Li8zidWZ+JuPLenXX0r9Jj2ZMtn0QBPENlPlnjsVt/rJZ1GSovl9FV/olHD
4InZq9rhjwRFaClAn70dQ0Z0g3nWSOb8aeHpQERnz6iDRVsrc+oBdB1LMszhVpheKuN6SB1M9CYl
6kj7maUphlGIZSIGaJbhbJiwyJcPwXzM7ML+gsietCRDFWFo4ZqOCNsSGIUkX0CKmvj5D4amI60c
A2Q2ndtRsc58hpUUXT5En+5tNCA2QFrYJ7+4yEer7j1rZQcyJ9CHHkNANZoVeG0s+nydLrRm0sBt
kV8D//OynREyhx82xH3hUwy++sicvkq7ZIOrMjg7f4FQQo6RtoZPgRHhDy0ubvwb90uq97M7z1B+
Ae6Sl7J7KOwJlqAjHy/3o63YmNf0ad5ZTIuyX3hwnkLfrAKt8DrPegw6qEDZUAPOHIg/AUG1gFf8
OYr2qMNR3wmmJxgs812/Mq9OMpnU6sAUWKwIhz+ep0V5K0iC3TKRX95tfSphxpO1nhIVAj+a5/d4
ro395/hafUL/+/1ELNyyG0vWvgcRSGp6OYtCj3OPvLgP36IpFf4PVej5pFDr6lpSkUHORbXEc2SP
NRp2YO6Sxckiael2u7zCgmo6nzK/bui+256ggnWVKuxF0/tKUfgZwBPK2GsAnCDqx33lSi86nF23
HiGj277qkSNPAyC430c6rbiRq2qm7PAVjBovNbV8bIspl1fESJO/XQnddTxT628gxPYbfGgT82GO
TvoT5GWQ0pjz22xthURp6bXk6VrzY1cQVcylDSQyqPqWrqN7/etXdCcRIqq/s3V+FWuqEMN2j2Ko
Sf8wCztYjna6m/AGAoVYfBAKEyZkh+3vA6Abg1vfwRLgvmnwWKr4oT0gcfBIcJgNzUsQL2e9JTqY
xdQmg+/d2LLAMDsyhxbiEClWSnM+f9xPTG6RQFHby7D3RGEq++IhHASJpMIE2ghkE4ifBaZhCIMM
IM5Iazf6K6h94gUj9dASmsq3su0MElYbJPDugoUTAZv32je94mncSGhGYcI68tzkq27gS9tP53t9
+vRjkXK8qQDbeOp2rGTkbp0B/zf12bTSi7w6zY8Gk/Jt8oOm4cv7IRmdAXGG8EiPJ9s1wrIC2un2
aZ6m1W7jwkJCH7W2ISBC0lWRL+t1HzQzCEyCeL4TxvK1/1ltWPMAS7fAW/ClCzHZ0UgoucCgZQwz
QTDrnEk98NAmWKetm3WfNGlqFgyxZrHhmNODKlL5m9NjBohf5uHlgEoOaAg4MHmx8gmLLyZcb4ZN
30722f+6lhbovyptwk9ODyfc0y5wSGfSvekYovfvEzLEMp20n7vSCMhK/p08wxt+pzF91V3rbeUE
fwbO5HC4rmURbme8tolHtF7IOaRNcKbM7ljIzk9ldGBkBEPJcz46FVYiYJ+5tRKs3TnxomtAIV2k
YsHJowONgaoC9TpBul/VEYG20sxnMc178DJUyP/+s9ii5PmSilHd7k5+beAaSKoCcswklInkzrJD
mMUPFRFs2lcGKg22kOYBNA4KvlucczNKNFmaW/vTCA5SHTNz09QXd7YIIMqyN+PUobF4kOunVWdv
myJBd1C16GdnHbwPrYBp43jTSDjmFM78U4Pwg7novq8skrRhcFwcRij8D4Ol4jzcnjfRy2ITZ0yP
XLMBw7HUKTVauTvd9kH1KCafNF+DTHi7qummBp9J4rCI3nsYljKfZan7JJk8CedHmS6jdaRVMw+A
XuF7Zp3WWIjPJhViSWWkpDb7v3/f9UpJEnmvJuD5qwo+flWd7uQYjAvU42A7afEF8tmbB0XnH9Et
80eou8x8BnC9LStlWwK6RvbjvS3ayJWBAwzX5/fNYqtb5LaVSHWbj/1FXp8+j5aY+ZZGO0InDepL
qdtXwKkAk4Jki8zMm1F3aIYSpcNkBZkOHDXefjmj8OuF98vk8f+YzlP6JvYOlAarW+cO71Uyoup3
Ipg6rVCc5L0TOjX8B7l9TJLpGOPACNoeE8poa0ZvJoTaW1wJVO7/OQyYUddf+sFgqTCSVL/vapi4
LH4PMDg0yftMGhqGw3n2dB8U86dQ6vSCAg4GjUa9+pq8p5FbQwOEbbPYl4qfTRikDr/ZqRLYpQ1L
iyNSuhA6t40Fo+xiG9DW7mF+YI0B89U98oUI0ZF+nLOlB4HyFZfNF/oaAW4GgTiNbvy3z4rZhRlS
cPdumvtXrUS1H+YPwinLmQkGbdi0WHMFGNXjS+3c0SOV2bSRKD4SMy8HP4ZkvG17XMpe80RrUkUy
RJN9/SLgRTTsAifONNEyU9ERY+7IWXZXWYZBXC2WDCL4HwxxRDJQPjKGbE5a6EeUeXzgKN+kEkJe
nb+b8VvBcWpcy0g7IMEEgYcaHNGzL0c1uGjWJLBTA+AFaDFi4DOLb95YF5mtxCxq4ge1v8WwH7lT
p+QwZgCBrAsgCKLSzkDHPOQGTbDS3BDP0qTUKnOsxsCK4J23UQ/wV8qi3XoeBnkkfQA9sUOmBlom
2lZQauWqz3n9N4nKsXPCkYRpl/wO9OsRu4aeNH2fVJMFCLZdNjhuw3P2+DXPH39D8f0Df0HU0+ee
FILsw04ko0ATbzJQrI52hSC6fSx1PAfHaS9pFLyTtNJUIg4eHJFrcbXcsnvOSQLLpywUELrPTFTl
++xlDBms8uZLOeAyuy7sR7d8v/UBWu5SCXZdubbafQ4F/ck1ZIZZcBWsd74vxT1S1x8ZLjvnumjW
FXutufdFP9Y+CUJz4yKzBwTU+s3wE2R1yKiInIREyLFxcyMIQOLlCHIHh72d2n8h6MDF6yqBaKhU
MITHCBAKFPQvSI88G6Inr28BdctQ5JxkkLVYWrTwL7cELIcMXftEkOWWZ/tFPJvZgoOJBVlsICAk
4LXV6WUC56glEgpOAltSynDmB0qm9HD6FXDBpt3fCArO4mdot2IZYuBMOp995yec9NE3k54jIpSt
J9+EKEJhRh5j/P32N3zS5aBW47+d+cWbCRN4iREuqyyIycI2NE9lLYpSunbdTKfDDgvneqf/Mi3t
Ws3RQIT26jY6lnEkSwc5CMyEiOET/OkW5Kgbsuufp20J69AnuJ7VNQpcRqnPTvoS8NiCFgQ/0MzW
EuIytr1kBmcHtZyzVFULkSipprG/q+JP/nI7zPM4d9o04t02ERef48lx0cdwgA92BK025lWlxFpK
+k81LVvLQqaqYyyRAk8Th9/oU/wwarKFOtLw0T/kbp176YrfIYSLzIsJQ4i4DvkjMFoxZC4ZSWzu
BvSaSvL9BdQrAByCH+Kv2XHHMEKHo9TlV09D+ftOd7kc+BcJXVpC/a+DUZ9i54GGfqstl4BnS2Qr
Lf4Fp20PDz29Px0+Ta1wUG6gX8kzyiBxrApitjpCFCGEffp2CmShUt05vZ3JXrfGMzSMPonOO5Rf
vaJt7eInwheE50+pkr3l4gKZDUBNXDxrklIm/Fa+FXcnb6h35524vfJTYqmABnsHXnQn95sQISB3
fcMuYNGlJrAZT9mN/brXE1SsXY8rFzG8egLrh1fKO9axsasNoYRCvuKB0lpsM+Xnnrqz8kGpLt82
y8ge2XZ9tbmR7kl55umjidK60W7Obs92VV/9NNl/sg433KWKgs93BOd2Jn1Dwcq9/0rnp6pSLv6w
dq/ZfUpK2qTVft+W9N8/JdbNnVnhXDFh5O1DJunQqscLYL4uKhkIJyaoSOc6KRUIHCBOM8fk8/0e
jNypNbz9s9zG9i1wXySXseNZDUueA4o/qCV0/ngZsSB10c6W3qEB+HWE+c03oW1CNVfDworHWqgA
HCHyhmtj1JQPoG6L5JNNb1pKd39ZaagPLE8V5IKVjRnk6FIfLs7ctT5PJ+Rf4BflNj5XRteUEqKs
Cd/K9H8dii7Jteu41SSXEILgs5Kw76LXyYpWQaziO9qQjh6w5Ph3dzqkHZBpLpLcj2tkeWdLELCu
73rIqbHcIoFprv5nrETjNUB5P8c7wOkRt47O4RUoS28NyoB6XUDV+6Z+XXYacMBlim0pQbdSNLQw
K9cZbXam+C9XkPoh+DqtkQgEAihW+to97EZc8mu9SCmORtG/wXYDu8oEzsHQa5ypPyZKA7DO+Yu2
G2cKHaEAUWjIwFbw9pPcJ/NAisjzc71EXaBY9fGVgaZvi/G+ySODcU/703ZAy2TABFpknH3fku1b
FFH9AZo/ss6Uq3zJ0Y/bedM8m/Hm7quIeB0plTcyKmaX9rK5FOKJh04Hoo8iXWd4tH6763Par64x
jSuRFRtNAc6XpD249f6Ghz55OLaGnQjPYT0cfKk61vpJVOEsMzHOSOVMwUDqWhnryt1FyDRlaYER
nhsJiIjnGx+yjYz6ftFr8Ei9OLOaTpdSwijO+lK2SEU6cxeQeUSFhd5yFiL+ncnTwAAjj0zPUKGu
VghR+biEdaLslHFDYR/vrubP2P12cIreN6pWv+oePkoa5AUUeQ2v7L9DT0loS0ftVtSyED44hdkW
IOlw+uI+ppjyK2Bt3WYI0pq1XpdfC3V7wbdZcvhB0UJrxC12ADL54zvsGMxfXxY5FNuwPI264A9x
X9SQ/W9gCAVefgwwyaNrDF5INpc5cUGD6IT0GJXOvgLA6vhfw2a1XQ9Wz8bki5ME8CW41FfybXCa
QtgJdpxVA7GeioGjfD6nVK4CuiRpIms2oac4bFts8+6UgY7ovm3PvD9lz2Fee9eWRtT4JASyt+ok
SLTdZBKfhRWAEx5T7tDWgZAb67dtBHnajvcumzSdrgVmYmUIVrN5swiP4m031LDogNRfZCfZRC4Q
c2EmBcqc6Yg4zTgteElC2bb/8QCm6q6iuwFeKyzDvCyUy0FKmqz8UDcqJOXYxGIa2EiyIcNTsG5M
gP11FY8FF4F7px+WEhC5xLTkz5qh3q9O7CWrMjZXIjldM7dE267RhEYcBcQtwSKYE6KL6QPTlb7/
1/1XyJ+L/EaCVDC3gXeaCe5SK9SCZkG5xGTnAixAF4K77cYIB/mdzT5V2HK215XWrI0uKjWbydAD
m/vg5abr2vVR5ORaSGbS7JWVgKCafwb3zkZtn7GssHEGh9LI/5HTbrlUK3bCLZm2HP1cqGroYFw5
NAhNfBXM8yLps34vpQ4aVhKoXywVV/g0+L9XvdXgAWI5CMZvJY8Pw5aFVfxkFC8XX2q5bOFwCzO6
juux/cX3k60iVdSmHrhAol8zETWtKkaw8PmMNUDjhpE8xIo25AjYwQNQW+A+hXZD+AKGOXXpIKnq
dhZFI1wHKjA6wdClfLF5pN9qHkokuGYI3PT7t+X2ls5Y0xYsHY+Bsru4YIenHzZIHHjI0e8TeNzS
wxShmPn+evROT+VpDW4ZtJjUmYWPGO2UopFmrTN4bL/6364O6cdgNk7RM+Vpz8wmGvGwjFINu6v5
KTUAVr0umapIPtWx/VcuWNfguNIempPxBc2eYfg+b/GD89nXEEYrzlXllwE+n68vemZhFPtqnW++
Zm0TQiomAWAVcf2yxIny/0hO+y/KRCcx6ARS1g+FHd8PDG45Hujv2iKZtxUrgOtXKZD88p1kAez6
W0S9hIn9FVg7e3Cgw8qwty5mTa2k49xjMp6dpGMktL80huwBdoQaAc20OaZKC2vBW/k+6WhUOisx
/UaaCs16DM7+ruAqYkDWGQPQcP5BsE/XcNaEm80DgIjzs5Iw1MgoKJOOwI4Q6OWqil+sV0hG+k2S
/KRj2R+P5j9qmGMJ2PVbMjiwKsjul1nHpZcuPvKqzqvBszQs+9HjfPGQ9IKtaZqqmZpysHkdVBwX
1hU34dayMKAJsOfPRXv1zWz/ny7kyuiYfnnyGo34O6a7dYc4207mTKcn6OgKuSNilIuU/e8EP+hY
oHe9ZBPJacZvW+xX6/KTBaKsgXwvwMdvqAibtk+3dQlxhsU4VJ3PvYnrVOosiVmJc5hvh9ESSQ9J
GCwDM4iqLbzqdh+Ma91b6w7l83+A8lo2lIBk0Ep4E6xfZH5IVc8QmERRSzG3k/3x2rftuTq/cNF+
AhHvMoVlISQd2lOrzR5/XGdQ8MHIM2Q8sN7VKAGgmoYN24J2X7o5hUNnT1i5FOaPmqo3tz15HvvL
PJgjM3+J9qpL4LhP3HkZjc9kiedz/pjNOmzM8tVl8R5a1b8VebI6mufLum0FZwwsSPr12UUsv6Z8
v21pSmie9LQ4yc4OyJ9B1bQjly8lU31aJWc3nBpAp/oC9JMEPkyfoU9NTC7h1IhzSIvSwFaruKKo
Dmmw2lYlVEXAzQlMMBpKzQne35LLRWU+eRf7ZIgxAVSdd6Z3BnqNoW5IXR4HSUFKhtL5g5m6PS2x
AYwjiV5BZBcrap3T8gqmBmDM6MGwnYkce239nKus/I/bcTGvdp73wdMDxw5MZCTz/Wsh4ls4PS78
koUPkzNKgUGQxwqqAzeE0tcYwyuR6/lSN+wYYZ2frzRISMGl19dt1WHDEaUAJ2JAm1x6twSDBKJ/
dm4wvHjiCUEGMo8xqIEXGibgYGRbo+IZK4Uoz3VWCbJAd/ZIbdqTJpVZfM9kOSB8+M/ov3YCJO8y
gnMbn39n6UTWnZQEGzDBomFwnIXg8av2dnlD09vuKe9WlL46MiBCpgGc34T1YnaDtr5PijIF1lno
xNfIdcMw50R4wHeYfUKwAPSUD8BzZBYAHrpajvcHway6tuimlUr8vXBdVHc9/cCl2HSrDNFjBgik
9dNgemgEUSOIjW+kjn636XkCx1IcgxXGt1RKF2he1nercGvrnURNleuMNqqBjfcbSZEWCdTSacy5
pwU98y5TRize6W0B0SGU9C98ph8kufuAsxo2Z5hKPrRKgMC3nl2YrlYVlyacjFkQa51d6WY39hgb
Fpqg2bFleEKG/GvOec2/6lVS5i4pkgbeEbwpAPaME14yIkQAlk32MuqEzav2I9NDje+SvgTjCCVZ
ztm48BxYZTlymlEwwWD6n9keOCvgxVmv3Ddl+vudlb6geU6KGphJx4olKwnN5oPoC4hmEhC8aW/0
OSPC2KpbQ4YgB+XSW/IEvmULAu/dbf5qSvJMHuPyesAbexhU2QR974Q2IVaQf8Dk90KNzIIx5Qo8
3Ty3GGKymZPvmjoojVmY/8QEnP7HWTqRiQJTA9+faw+ZGTNKfZDIbLaMOX95/PXMP8c9GVxPo7Uk
k6HNTz9laQzBc9bQ2VzDCMaWdRrVK2CsuJPFEU9/uFP/h0mIeQzjAecK5qdsfdD8gNVuU/B+NqLF
jndocIE7cbP4lhBkeOEJl8YPQzoGaImntbcw6vCbR4FdW2J2myE2VbF80O03mBCHSGLkobKIbO0P
I9Hb/e2hsD1wr2FJ6uS4fgJFam2JJbFqLOauPddRfmfSs9NQRY4nRpkZs6mTFTiMaXjKo27G5vDD
8rU0R59Gck8Ib+KqPCa1K0bhxW7Xe0a3un8K3SS8ZvOj9DX1Q/TQt8EFh7cp+qWam175afG2OXIj
v8ISEI2uFCVy6nEmK9y7Fm2DLljrRHLari/VIOai8ffirFKQ4GAWaDAXwqA2F/CAuzVAOfGYpmYr
ZLAcNZn+77SueFe6K0mIz3eLWHgVcWeWgujwP9bH7ZL2GbbXtwm4yILuXZbpN6qVwH6aj1T0S32A
v784ODAqRONYHLS764xenE/Hhdr+S6yCMerzyRPmSlW2bIlaH/5ud1AfGBV3L0DCr9tJDZnDikWC
R6wyi5tQ7eEjSYl8h5fYwfAYX7/Eo2ajmMlUcsoZq8dwEcJdGBh7QaLuS1kHDACDDvR9CEonNlY1
WvI+VgkZxTcGsUL+FxVkB20E6kUyo2Y7wyxB/bihwTQPt9zoipdNlI0FDl4z1krBVGNkc8Jgc89K
W+iX2zD7haX/gQ/uKXjmtPqCzF1dC1ZyDrjs1YjM6XJcRU66qp4IMTuxKrumbUpCLfhcQZ8g/R5E
j4TMeo/3nc1bvJbJY5gQcD5w4DY7IN3Th7LwS8h9T3Ni9PjdgjxI2jV08+hB1vdbSUnRUYrM2jnq
r5ZIUbZt3V5Zxkf4k6hMHfToXi1tapocMwykM28RFuOIm3V7ki01bc624ZEH7lYoQWdnwF5jpjpw
N5pQZ4DySUZsu7LUfA8HKdsvdsjQmp/wo+Cyjp2gr6Qyn+Y/ynA463wtONLeE/Kljf4Pj43g5/td
qBjUVZtZLoxYpqVm6QnAtTcjT2kX6roROMWRQIEuwlcR/tAswonVH8ZmDFnVD1oIsftGCEEHUF4J
bJm5WiuKRFe9WUI8uZvZwPKO4FxyMNtuFk11T5xusLrBoEZtauG9oRBVLEGe7QnL4FSWHEwyVW6B
pLXNJQmYUOcTTFizt1Fn2DED/QRhv6Cyd8BgQhv2NPr16AnJwAH0R0daLje69SWW8HZyeWK4YVEJ
sap9LV1xQIHr1f+LVsuCUAc/nnS7oAaNYvlVEar32cdimKnOnJfHtQRBRn5i5bzYb/KiXVSY2V3V
bLJtrk/Ke25m2hL6HR2E0bA5wTcu4tDCkOJvTDxwOT/HvesTKzZGc9CiDyqm264jMDfVzCWe0YAQ
ekioFAikyazlW0cbOYNRTJubnKsSi03OzcYFpamPeYzQOImyV5W9BLPfYZIqc4Vh8Etnu5Ixnik6
8qYk6JynbwAOvhii4WOV5rpYW8/cyoWoD0oxK2NkTSErSJVQlBmMSSfhEDCdhTg/jjIylSChnJ5S
Y8/OELyTAu+5nLZVnrJ/yK1vTsJzxP5Gc05gG7wFZeRl5RRzhPrnUJ0TMlz74GMazs8830QPjzLC
+THvM6EdUs3R5PxupeezhKnay2gJ7b31phN8nMjCyoaAvJl21G6Dy1cNmt0M2zSjCM2AtuzVsdZm
MGlMFCbyUpsvmTSjUZRl0AADv5J6wr+2fiCax17vuU8o3lwlOKrQ1WzUUowDBzeomkOueHishWSA
Sweg06WMkVIYUbKwHpR47am0t8PxfWU1yLMqnWBtRDVvwFP/lG7qwLLJ4k44+MmnZrK5qE5WZ2M9
cH5lBREayasr8wYWV8g4X5MRCOiyZEYKD70/rhVX7gEys/6n03s/ZCQKspqwWjY+JL+yWB0HKYaS
EOXCg/p5+wPoM54Vy6Rhj7h1q3iPL+Jmn0Vx1dzEceu15A+jFcMh8VesZy6DHxuCHbcFlGsIyFj7
DGA+7ipjc+UP/jflnYSLzcsXqqJIHjTebFYseFOONF3tAXtc9GY6mb3MclQ79PcWCjPeN72bOV+z
WzuY8hloA7CHQ16y11QyKNs0LsVv22aN7EajiXj/4LikWwn7I+pvNeMxPnKJlpylYu+CQEM3cm8K
OB5hEHYwQUS0u6roogl06Shz03ws7p+N1xjs1e1za96rZIwpXPry6x40tkziP3hObapV1mWs8wcZ
JnPNj6ablgYkXGAfLp5Ub0AUmI6P1REPHmLBdGTcD2gj6vvAyYrUwMGbG5KvYqbrtCV0cRKK5aQd
K+W3D/5UL6rKLnTiCSiXFjLI6j58LoZDZFxjWW+gjLa17GzBSYcq7JyIeeH6l8a0keol3YzRpaaj
oPZdhu8YP9GjuleYbezf7SRPPC82XQ6XtPucsCOzKhqFXmtJl8q2FCQsO9tdrPEK3+Vg+02WGRT2
vfnIPCIhTkvb3k84Gp52k70LiaCKfznb0g/ZD1kAara5jBvhOTNMccwvqsFbV8jvc259yX195gkp
3mVcJHYA0XOaZQH3ooDu+Y6v2DYiBQnp6XurqamgLdH9CInX+9Q8tL4OiMfPkOkgDUapfw/Bojme
diLiAeAL/Wzd+7Z8yCVz7QCgdmkRjZbzsDmArtoiFc1/QqXVnOdpiKx4UBC1ZFd+wu/3dokvVxo4
6tjOjdzdw8eYe7hnirdkClQIeYZcv/VE1Td55/pBN55yUzhYdeR9d2YxeT8pApx1MkEl8CFXkXqj
QyD4dY+IPOVnXMs9zbxPxOgFn2XwIg/IR7u6E/yAhzl6W0MqsyAZeocA0qbeekLXnCWb+JNhNwYI
DJ4tzh2HHRB0d/9eSvcYyUoeQ1zhlc0s2SPx2Mtujf5XtoyDjpE8iRPM0rzvamZfBWsd6mSz+qkM
c14VzUFgJiapXheY5vWaSB1uYJdd8oZbTuQs5kt7FaIj8ku4Govul8h0y9byoY3JqYn52dkPeHUw
nDvfDU0P9kXy3NxspXgwS7seDeZpfcL/bj0spWy0zuUcAByHcvv5+q+Jb2g1f3qJX+An5wZp6jbx
TEmWbVlU+UYUmI9PvQ/DKy07njpgEXxgtw+sBONrOTlN6r4nsHMqGD8Cf2fiQ1dYJzBVcIThtM4D
WZFZEdesqbO7IdGV1IP9duFNWLrm8EHt3aDWWXZCtdwcKJPvBrK/W0hGdUp6H7rgk+UjrPSe7y0Q
UvHt3XDP37ZIykYXWTtPggCfpss8xfhloHO7hhbya0q0bMrR/ukFpyFLp42kTQUrKUT6IFmAFbqf
8bukrXFPyX3ldhPfffPgNsdIhdehNfkmHJgChGCTm3FFubrKDNKwOo8pO6xyGCVaEucvz13pcw2G
2rpO8h2/E7Uz42BAxgVcYrOX4dPDY2rj95tj+rGvvZJGNG2K8Ig989d943ozS+e0T5Uf10dfOu6a
uMTGdcLKEEGywrZV+ilVR9Xb+fbWjgA8MHpb3SQ3TPQIeAT1qiy3cjiekLETZ+HgkMnquXFhtZ8E
32vIW+Q+yi0gHBfUpb0QWRJV5TeYb+CmMA6qz3Iljpvakc3K0nwioJddKU0X6dm0xQmnP4YE+PKz
KRUYoRGwBVCv4rmjYrqEh0tKvobk76okDP4rt/to+Au0rOy0hGpYsmZck2MZKtWJx63MWo8eBvqt
phWvHsGiIF+GADCkobVrNOqUTyMLokBP8UT2QhSIXntLQlLMrKvPN6oiN2vEKcRv/9Q31IkSCBZJ
SOsj2+Ea95NYvCSFOH9632C2tSLVIFwmyXEhb9QcxFptAfhheLdkclxV7xOG3OTcSsvNNaR2kwzs
9UkIn+QLVLBGbczpGh0WuY9ynzgB7y+rTYfyOpDWxZFPWoEdegx7EwH6bYTUXH3eyXy77Gz4I7Xs
1hwIasB9kd6gEJXPE0K+54GtmaSeKfChSr2xxwCHofUQMlWZYxDU3K4851HJAkH3A06Y63QOFLPf
my8kRFwCJcm2UfcDGBtgm8walhuSgVV5dLoAut6sDQdZ7BOsHzs2yNgMG6qjS9zPs7P08XeOnDZe
lFfDLpiXc0E1uDKzv/SYcI3zYnBIBlFm3bGquWoGD8VpK6RziZ6Hl2S02l4d8zIxESfBHmvvSyGS
APLsU3QvGAB/quYMHwD3ndBal6Zop97YwP91t1cD4+BbWseOJ7yIZJwrK1hiNwar14snwAcOML/g
SRF0oKSfMykLvYaoihgzAlOmZklWg8cn+yzW/xoUqsFJmtGPvrZCZ4jMr8toan0hvuSz666ZiPr7
sTW9rNITMCRXfhER6BY8DaFJzFCH9/CMOSINBRIUbL4XdZSqC3UTPAlOQWhEeWofcZPEkdz2OTTk
zwhShuL5/iF1ilL7PLhnIWbXPLnGTkPEd5yaNWOOCeqMUYJXm+hGMJnWYzRHiHi3gG0I9ag2HBfT
CXRXqlO/9RD2ToXJVQjdEEKCRJHWK0whh6s1Kz8uD8EQhbBEkCuKr8wactBkzPL1pF9i9ma/at7i
7JlsZgyXEYmCqlWFGhdDGioYNL+AENtjkSYnwj00MhXElK+QY8uWiLdg+cYTiMleQcTiS57x3LTR
98FxE3putKdCTtIDBErSQFGXvkQ+dlZPmCzRSsS6ispjMlF+JBEIVzRoJoTEJ08EdR0ri1eHbSse
JhGMl8foNWiB4Nmg0D78S5NjG+TyUwbXfDnIHQc5ouQzHBJCDaUxoYrJM97LImbXizg3Ink1lmBk
T3D1putXCv7gWsUsimsv3lPkHdvv8PilQJgoc8NT8DT/9wk7lf+lpQ5CecrEPXTZNO+tDWLjM+ep
5EDK8qFYX8PVG6M3a6OlItdk7vYImUDblAMfMlYkO/lzG0Mlk5nteGBovnsUnGHtj2kcCJgXjoGl
LiiJb0HLkE004JeXSyK1e6a/ahQvFMFrggjW/M6fxBP6Dd+XZRFS6rprStfjDAwLQFbj3CIbRZN8
rhVs+udAw+E+Wi4DxuKx+4fjRUNhXs09r0ysdFAgjLi0nfTUQdg4uJoDkFsaAouOFAzOX3xPFXs7
LIRKhG+EoZnOXELmFvW5Nlh/AwdGvyfGsCPhyGq2XjPvU2HNc0rnEWY2p2ZqvsqB0PATXDLRYOnQ
fefPCR76Sw8POALAY7B5CRzgkltf6B5A0/9o/jH07m2PIMUaTEIvAshnHQfQx6AQB3Ujq+J4vE55
W/vt+sOrOu2pkCFwEFm9vFo6WlskdZBnZpic1eU3czMAvYaf/XIyMQ716mEzpg3R0oDdY5Fo8PdN
XznrX55XtuZEYhZMfGkl6TJXd/eRZT0t4pm+PfKIRHPTgcanGlQ1KfwdzXNq2dKy2LuUjHUwjxmE
OF1c7GO2TTPhV8KxsPaMa+vdxVKX60SbZx3wSdrLJbe6V6z2aXglapXXLjnKtl75WVCzy1e2OVO3
UKmlz+RIFTtdNv0O94vCdCJDF/JzW9EXP5q0GjLEzWla2hO1zRiAs4QtQLKs3BxjXOqE/CzKDPMo
Y8KQGGGHuPnLCb8M4lD0T7B/DpZjeuhxk9HInAW2yPVlomYYicFneZ696vbqmz/yGZELl17bODQw
rfuoM8O11a1Kfsys/Qb1ZeF6sVGwOTvACMWYtyFzhVmVrzExx1WfZZK0AjMvjMP1Vqep3UW1Ojzo
/5wmUm7T503zmWJ/EzHJXgbO2hRXvuN8qCTgjihUuFyGtTE2pGHj7laYh0EPDelrkwh4a9sGgRL9
VcH2jJvSnM/Opiplv8rNXRi0t3xVf4ZwY8vGm58mUStLV6RxLEt7CzR2GXsGy+sHFvA2CPsprmMw
8aBTBIQ/uM0LBtybxqGPpJnrzjrkf1X+7fyxgTPwSPKuyi0z452Dz+eja1iCUrKw2v1TAANz8Gdt
wHhvFdh7EYq7ss7vWvzmp6vQQYwEn73OHg4mhTE/ou1/M0muRAYAOfG0XCaycqSg1tQkTpgAvwyF
6XeOaLbDgAzLGKoxysbpZeuSjudpKClFWoOZKOMtgsnlNpyCm7+/4WGzMX3H2+O+Fn4B06jjML4O
Dhx6P8nuSLlz4vvi+YpBj2RgF0boFqHK0K+mnG9Zy7yAKnjSzo9pEcbXfs+y0HtGzvK8RXcRPTB2
yL/AWsDD2wECPmI+rTCBAWTgOiPeAZnXxhyGtkEF6akwrEL/JcjeNv5t/rLT0lRJS5YAu0APsYbz
8sIcc03AD3DI0ZXP2X4Qdft8qkXqLARBZEZeE2GLMf40I15tR9FKTywF6qSq1hJYPWCp4UBuOR8I
bqhMAOobEvdn8QRSBC3nNDDRw3mb/jSTo5E7mEk2L9ZtdXWKTa/bLxwfc8hKK0NhwL0yIDOGmivr
WcLo3r9DqTw+OjI+Hzqjb+d4MzN/rlYZNPVD+ctkVxpDJcEIM+XsAmNOvpfK6yN6dGP4q8xJgVlf
TVVEoho8ca4lVypUm/T9InKBZoT7D398QzdshJPV3n1ATagoAOoxHRrCLlEhZaUprhMamj6Owly5
bzwsmTFHlDbEEfJU58B6Ch+eCe/5EgUlLrCAytsyu3/JNXZBANsXm/YvrPNykT/8Q0qsFz1+Dyja
F6Y95niZWTmEUnDrfWHicoFjM+NOfYYZnW26IaK14GpsIWi1PAG8UHZWzyrj4DqDXwtH3sFVOZ/m
aBO+CxkrOcZL9ziTve91J6UDhJLSU/Y9NzkYzctqx0aviAYyMHInAjlj8/Xohmot/HiwYS2svJM4
EPb3e4vUKWtLmlk+V/SBEGs9qmB2jnAT/NV+qz6CHnTVwkAeZfsQlbyINcF3elA1NTdjqQ4xB4w+
lWP44JyplLwxuRJYeVUG7qko1X1ltkgL4wiqtEx2mb9MbTdoekK9NXts/zvLnZdygQLs9DbtqnIu
u2XThA8G9IIw2lIPHX4JknkQq3nsfkCnFjqPuoDwwFwJxVoWlNqwDVZuTnngbdOTck/NWiLaHPi1
L7s9PNmEpo0oQx9Whh8tHGFEqNc2nWk+c/vo71XA7m1Xa5zWwFKVUFFAhF1Fs8UjJW54nIlsl0AL
EIG7yAWE5/lQklUlJamcL5IZkDoVZze93m7X/SGb3jkozc5jPjDeJSe/3BUqMhP5wJNIZILvvCgP
qiwDMXCWJJ8SVrZmX2qb11VtWq6aKUutIB8UzheC7FO1GgdzFrt2PmKnJKTtqyatIZSVCcFsdKnP
Attz9aeiDEHs+5tTEFpKqeeV0+W9ZWZ2zm/SQdTu8F/XwN9ifUgG7/V41SyyneJkbPRrtTpkCZgj
WiBzP8NHnqdsSjSMaWkDxbL1lbXgrYuW2RUTeRIYvXmq+O/vEeKI9EZD13bKk+WlB5tWg7p+OtEH
+pT53O8iv7VGrYka0VwP4XtazMpEtj8LZ1PQL/XBpcYAVjheVoEXGV2e/AqiGj73Chd3b3JaZGOB
3Nb41+/7Kc+q4d0q/1lhLO7g0G6ZQxmxf9B4mZM2YDI+yMr6UdHPQdbjmEDk0zCnEGeNaOUlhqc1
oJHqOf5bAcJ6xcA+eyAVOYTMX/IbvL+TxM/PSir9K6Qtb0NCqkZLYaz6PqwdHoZNI2NleBS7ngc7
Pxe2camhPXdWl79zGQ9uNF2U1KJK+mVxr0yiQDok9aWUz6eIxFG9a5amCz9izxTgT2AHw4JXvx2s
8gSaS7fjWTgDa+rdaISS1AnYcQZmkihvCB2kgUaXYYX5Onk1OpZnLr4YWVGEc4LRU0GGdQP2C0v7
gHa3AP3K5RbH2EphzTvQbJNwgG9Hp/TtQOayFKBkrYiufFJHzfXNbqvXBc9lpxPH6tmEIMJSgRvw
tO6bD7ZmX/9jzAVsUS+nEwroWU6vM+sf0/7veCRuAnpbNqhPOe4ixOH9/4A4eRkE8qBJwnJQWU2H
7VNcyRN4PbuR9ScDWdNTw4n/XkpP4ulzyD4pAFltfD6hNsGq04ty7tDu2g3Y26yXrRFTfwjRfibD
fAYIZLiXO59LfRJQZYfy8rXFMSMUp/UMRSrKV7wGa+jJgIXmRxnsfJL/2eZAR2ttkuQKoWicy8qg
r40gFlwj04FJ978GMLV1mJyucuOu8an8suNRDQYg6Ciovmsnw8ILjFk3Mxq/+GbDWVtSRzVkCkSE
sT7P/e0mTFjwVn/QOPKs8UdItWPnLEJo4czq8DAVwWCCp7lIYaCgK/HzE3HIExlnWc3ghwbo+A2Y
WtBhPpjlMxgNDSauQiqMEV8cfJkzZ56++Qz5ouDAHkzmizqLDZW2ee85hpbzAdgkmAFjabstzZUY
VQf6Ohi+rvjNOds0vdVgbp7WS32SHIR9iNV6bryV3KadAG3hobjg52j0FEyzongeVF5Pd+YrJ1pV
HY9RPiZt7cvPkTze86M8SXh8KYZT9FCj3LDQaVRtKevdFbhc2Dpiu3nnSXIrwFCsoP03bQmvgGx9
tERbgQ9AjZgFp06MZljnqHpq6gyt2D7hSpjbh4Uf+0bcfnWO6t07gLMR8A8/00UCsFnoDO+rrx7j
X6GfEtzX4LSs6v+NjfO4cbR/Y2w04OFy1vhtlqsMWJlNQLgIJXiacTJ3J3tRdBOUAF9saOzdMddV
PGZpV2fraqSBiSUhOBL82fiVm/9qbXdeDyCB2uF3mOHU2X9Md/uaTbYIrZeZhKCySE2ShgZxa5v3
Uyt5lEOpux2MeCMESqhGeosHPZKBEmeJCdIMHsLONm4RvcB8rfSqAV+lqpwtCSRJ/geDI65oJKXZ
lWab6Du1auL7LGMT7d4J1xSk09kVZodjRROeycGu2WnUuRXJJYJjUIvvhpLWgQTirhceN04yy3v4
RJplROZ5xKkakX4vebDrGqMcEW/cB6O3PU6UC1le/bqQeyHESF+y+rtEULFF0a2Of9Bud0aAzpPI
W8Su0e/b+tasL7GpF0xLF7FratR2T2xmnHDGo4EitcwtHFmJ3RZblyi2WV0dqEyB0T4moUpZ3Giw
s2z/K0qu6PsoXVay6AMJJoevYV0sYDuLxYL0We+tNG5v/ehaIH81KZgFv/N36Idv3bnlO7VAJJp5
WI7DoTxSkscsPq2CdWtEG1Axro1zD3Pmqus910A6UHKCFckXczurHqJbo7FyH5s9lQUh5cUchECY
qs3pLAGYorTO7AFVlGACOc+Tl8+RmUGrz8qAcOhACveOx6ZdLDI6GYDn0Xis3mvd0iXOLwYcGaWi
YdGWIavn6CJTLozFQuP2m54uwOkHY4Ca6SOTmn2YS9W3pVFMKi4ALDnPUJP6cMRj6NERFka1Recz
QYW2QaQVdBke2K3XSa3JWWFi0MvXnEP2cNsbwwc2Rz5e5ONLD63yd0mhdHvV7nc4kyFlpTne0yGy
EtvAIt2qcQpw3moNT0Ozb0c/ZcM1jPqNJG8KXr0qSHsxSOziZTfQx7YPkkeK2JoHTHLHqrwpH42+
W6LDDXjfWffyVj6GgSskGly8oIXOaVqqJ4rCi2LhGmzaxLflQ1ssnngAkAFQ0HtMQczHFJIVBrUc
ygQIJM/XCUIrjePTiI2hikLWPbR8aWhH4n4w7eltTWS000mYuGarRI0u72DqF9KimDruFNEG2+f0
Ad9oNd5WJb8xpZF4Fdp+aHXRsOWz58CCE5zpRObYZeJ8x4RUY8HUyQN8eD+OiR1znT8VkEHUeI5F
ymDHWnQlBoy5ezvgJcrLX3qcvkzp0/BABt/do4FXR54cIaUFF26mq09ARHrm9hlu5JU7BmHSrGJ/
UNQj+cO4yQiwmoAgNVpMQCVBxhs2485Cl26OXk34mq0MOakSWQBo+Ir3cyMirHNJJ7U5A5FDv5x0
B6Zl1F8VgVUFWf0X4/EeJWDBfw5imsGmZZxnhpuz3KfwM3bWGBTXm203ppwXD5of8yMWBjGIMhLI
NVr12sXQfn2V7+AHM3syDuNDrezkACVy0/k1tOXO4af3Wytt+iqPM0NQhn6FpZJ8J3R0hZiib0X/
WKpeLl1j00YrYlEHo8FL1AS8E3VbZBNTrNPinnv86PHBbiHCZDKR+96K7MvBDIkct3RhNSTT1G1Q
tZRpyS/WUsslnSQ6RAFw1dZXT6RHDr/YzTDTW7Wq5STGXB96AEBkqR92fT1vXayRHbRbwQRjLeRV
FbB0dexf+bKv8YAjA4AQBdjQPXwBkcWILe/7Py7iNHBhDoAmgZz/RSgPrzENmRPUUpuVGT6tjiOf
Rl/69yWeh9FxITdaCfUVYsIK1786D7xwmYr+vkEVxrljjTFcIUjAvxnxsOgc/HwGkUaKpridaK5D
N4ygTL4fPPK3kKC3IEM5k+qnYzWPsFFr0ltNTdiz6PcveqOwBH7GT6fqaZGFei3vuLy3AaqVrA8v
AQFi7PnqSxGlJPzI+qe8PaeFbEQHruBwaD1qdxhAmayPh75Md+m78g6jB9Gd3CRkO4PBi4G5/Bno
iB89C+QMwAHmwIXQ8I3XsPAgkV4Rj//S2WoMGrxBtoreNtiktBwgiic2MOLjeDDtCqyrCMiMbEEM
gxCl/IljKg7f3CT4/DC1S84Bv74jgGRD9t0m8UKjjsdtjCeFOJ2sXKPsZhcXnpFQqGLtXkiGGQfM
Ie2IDn81oPSDlhzWe8VwlyJZh8earX24EftZMqxnbq48RG6kV/qg3O0RfzmSZh3Jkn2oSuycaqOX
KS+RuKSe3669HQWO6f/STLqyztLlG1zBx77i0AaBtomtuNCugdLMHGuCyj6HmllrdioDFAKkj9rm
dv/TWmqmi371+vSp3A5Zz5biHL1Sq2JUMR4R7LaVluiLqWZWcVqcd3rfJqep4GpAIemRhMJ80wvl
I35xtrpTEWtM4Xt0OHYlaXAhTi929wlg3X1BRs6yz8tD/g7uWJoPdhdmx8w+h6+mv70/g5cb9Qzy
yj3ItjYjNxQ22MaZB06Yrl1IRClu2OjaozhkZfGhIziwxu6/NY5qVMwR9cwm8bcYYFfGreUsupyv
+x7R9lvUbIBOWxvwDg5k05vd8Wvt6OeAehYblWXNJBeujPTMT9IA1G6xflerqUlmJBQzN18MOu9a
aBVRcLrx7AFUxBdJX3m3LiDeQTuERrOo16WrnRfpZcdcwPA8m5Lm8jJfMtK60KxrjdwDrDuMWIhH
NmF423VndmHj+xryyxhixkoCvNBXEjXCh2moNqAEcS32ILxnLBn4gLAnn51HEn+ACAMfjEa9Xh/O
HJvftCwrQP6Rpf9NE6J3gMszWC2mcA6EQeHSPX295AvtfNW5zVcpuS3IgW3gTy0W5Hcv3CJ4yuqO
wp4w+BOIDcLE0FFSjvV/6JUai2eRqLpraSSVlYPNdNEPxSDi3xH2pPLqntaEyYABc//uGzNjcwB2
xABpq2BQCeMpd4MkM4ADjSAZZcTcoMPa3gSFErJW7wLNNtKB2btaR1pDgbJBJtBtR9ieqB51Yw1S
yHz+QXjgpj77a8Aq+ISzLONk53RxwatrbzWnfIrHQpwGQrHZL4Ks8Kw4AWNmXDYNwXEo7JqsLjt3
lsl0JkDTRcwxoAbz3Sf1O7rTG94BYMP5nUwos+tU1ON2V5cM3oOMu0pSDnggcmd9ogYPkt5IMDGt
7anc+QC7UZ8IDaWPO5SIclpLf3CSzhV2YqEfc6Ll7RXnuuJy6jyZzj7g3/XFFdRk0M0n9P6NK54I
vGX2DboxdMFCRtU36vHdr6FFHH+iaf3yB+ohkPfz8Cattw8hBqVXxB9OgDXuFIl1QdPhRdwj/Fot
VannZf/hEl+rP5PbvYRF+/KHXtN3fb4Faf5OF80ev6b63gL3Z2rxTmeJxX6e2gOd7bbW/VA0RuXL
OZZScFD7rSh2QVuwPhcvgVWRJ0WEQ9SRJBGhHM0FY3WWMjwdocFRCpxutWYTsV55Oe3rVQ0Sq981
xw+Wf0S+Wzr7Nks/4/7aZpcHiolRzjcAElnTVq4RXyNrOY6CLc0ZX9IhA5zYUoZMBveG/X9WvJw8
fSGLPk9SabbTF/J2R/1JWHDwivNSijsMt6B+DX6B0hB0wDCrkR8swlaQkIdFhMYZCedV/NJFrTvl
BVIW+luLfeYe19XlAI1uq4CK/2NnWJcAnC96MyouppyIxYxRt3KypU7U1IbItnFWlkl1/9WtQFfq
MikF60iNyt0qE8hwftqBAGnEfLoEbXl+X8WlBBZSnnsik4WmfcQOOp7s9EN5y6EOmoZUqqQAW9HK
ejUR0LQmW7ode8obdtMaxAUTQ9lmuObgSYB4lEYynNZh4PM1uY0QbkjWzq0wx0u+s+4lrquERLO4
3Qz3UgiLW/9MEcjL4QwtmseGvxbJd0I2xam8qQ2cmwU9RM/yoLiSEx3mBgjKGi1YwBb7nlUsuNVH
p7vUht5o72ZRE62RMM4X0qCUWmEyATdTgFUF4GTAk5hn7MOGzfFzw7+UJ0Gae5J+nkW/ayTyGC52
HIQ86/g3u9WbUGxK3Z4RcOupZRcy14lIomBYiRCIgnuWHTwcY9ojMAQ/ppu7276Bht1qi/um+pMc
gd7M0pMRW1bdi4c/unr3FNP+Y5apzw0oz+e07NCfuZW2+MIp9Y4pV3EeIMVv49hXjR9k1/u9hjOl
XqV8Cn//JJmvQuOXOqAIn2313MJqvMWyWM3Veh7/IxKWr5T5hXHuUvVWvLzBj3XkyQRrmrAD7LVR
UT1tsI6ApTVIyR1UKxRpZ8EyrjAMJx36cVVlJzvWLTlHiT4DaPoij+buRtCol182mrl4KmVwfRdy
NaWa3CipMhHwLwlqr+uR74S5b7cgHM9cAo8QG+apZA0RD3cwxytdvaJpHbWB413fL0TYPtIQMFXz
PTPFOCDecwcu1B1KwkgAIY5Sn1ZPs77/vU4CcwG3PZbysEnDv+e8mNqqIcrWX6z6lyH/zCbwlMDw
DsDaofwDjsXWEb+mHMkwU0oROmCxlt9+unysyRDyRiX2ZDyzHmYQeBD4ZiLnb/aiqU8XXuEq2G8Y
yBcKINR2izYeGUnhS+dEaAtDoqzAiMjJ8QvT1pUO3I+JVWThHPdnbz0IQkbkS3HbE8Oa1Rs1C1wA
Gmiox6QmaerrsZlYZz6Nn3pnpbSQNfiW56O/iWaMBQuYW1evtpU1zgj538H4dp7FoLY0ZJ5VJXRG
v+A4mThS2p053f0uua8kDkgUa34hPR1TI7SmgV+TlILSx7rKt/FgFJB3geHTTqMHOT68w7jHqDvb
K0GIY2Z+a5TyR1k0oPxHaBUV02SP/5epWUFM2UqdaDVCiKYum/SCvfsUWwXAI5jKhwg8Hwv+EF+h
w+sZAzygCdSvuM2csD1/XbEdX5LOEF5QL9XeVaZrcTXTAZH/u6KPyFsNYT2UU4baiyUwBiKhYFq1
yU7DU/DCeI3BdGZvvArDDCAzf0MTU+CzlXNxTuODMYqK9cFQWhbpLu2XNSZ6I8Rd58tYnl2S30PS
1n28gBcunFlFlxiaarlbacClNJuyAbJLEjPUR+f7OL05meViIM2rLs7p4bBh4lXA5otS/Ne3DM3g
8usrKE/kiGYL5i91FQ6uNPt+iXD5poQWf6xkhUO/IrGExoSeCQ2nPmEhzo8VYkdzRPowUGBRlG47
nyx1jbNS2yw2xMS/P693k8KBoxO6PgFFKoVkw5R1KQ82pFzKwcUod8YWmFoyqLX8NScOVBBlksjK
EEzhQpkgyZo/DpHg7cPVibYe4gFHiLjPrpjFESDhX9MhhdmqfXd2a7cWFL2tHO3PKmPtKin5L+4Z
CIFULVtaVVx0Ffl/bSx5eSantpyg1WPX216SPALr3LVBN8HaKNzetzHguvXJNG2G4jV445Mxm/Ad
LfODyQXAoUVaG4SMcbmCmuxaHrlbdxAEre37dDsOmZElHdYEJDnpprdWq8/dtf4lBqzWc2Sjm2mb
WJfcTHR7ARZWCzfr8FdWX5TrTQMIOEsGGfwRRz09i9WkAbQonteKkOYUcEOZE0hIkBIn6jxiLdqa
T+zV4yo/5B2n9PqpNxC6EUOtRGXqsBsO0Ah4moq1waIZ+Hq999D8X16IukUDEogRhk0edmErDEk+
F+LJnK/u+n3mblOn7YOYsWcvPkGRhsX7qdz38WT7GgEoilI0ihUnRib9pAlvyHtA5CmJETh39aG+
NRX0ZQEifru041R7/4KnXuYnBZAMhj9NiEnMSvphtV6vVH/7nJCj5AYZhqiAlHnRa6bGQuEhZF11
DCR4ISaCCOdwZHEo42Va7/pxvfWUr7kUxvN5dE9vKU3H2e7nbpi2b5kS98J8q6mdc+5ZaiC4Ypjx
lDh64HUrceMBlQ0JkUGyduwr1ZwjBlU508wvC5y5X3qw0GLXG4LNbVfE5+MaInHHjixE/7nyMPOt
EiqiQjL2rxt+VTr3xLlzmjGCzKiMI3QBo+eOVeOqBQ3NY0Lq0695nGNC5rlQTPIE5WtWG01L0bJZ
mS3mZnOuIixJGZOX23YovHXDjZ9ilcXyptJuPidHgjcMK7Pk2Q1Puk8VgiFNstDerqdrTqPH7r2b
42WaTUlV0p2xzJjCZwaAhNx+KDzEm940Xvzl84IS5JWcHLcK7QVMcfYz5DZH7SE2bfn9d0nRIc3o
W5RBsmohF2WoU2iWh3TWNsOu3CmUrQCeJSiyCC0Cwkqvb1IuibJHYw+ZjwORGxzDn4DZ+m3qSamS
3uWMXiljcllhXeNvce7mPh+aFL6PaFho6WBhhrt/j04M5N8hLtJ+PMjrrRyMuJb24RnTYme76IeK
lpqq5Pzl6dt15neVocH4+JmjHZ9qBypg/IhowAtnnC8FhyzmKZlHU94QJCJ/o7khMz8NbCKsBvOK
GezRRE6cqgIFbwhUhGPnpzCCFeJlJ/tsrlXKpT+qeKBePl+EJHYfmcxhqsMik7s8ST85G2YtQfhi
agCih3gqkQCOBYlZGInWzIDqmUdMTfme7f6+V0XyGT7H16MqTGaWmCNIAVpxOJydG1ZcDRSqtwN2
BN/+NKRquDgtwcP+Yj1QdyKd8/TdDhzgyPrs/vno9eli6hjHKrQRAa82T4pSypVCl7RlPKtV3zW2
xz2mb2fJAZ1/DQLxuDgAmkMzVf1J4XZcULJtMeTcuO9NSfEFvCGnpyG8Se3MnNqyiuqqaYAuJUcv
cajpmiCQ8blt/eCL/y5KvWDolpdcvi+lwMvTo7tVUGvjj2dKmH63H7tZdLYQyKghmOpGPRrOlFnx
/9tU9ewMEfQRB0FkgwaQIFKITgBsrrgk3c+Y3IcBbqy9XgRsAjH3vUPaJOy302yuHzvnlOMs/Pc2
1sSYlCjNtp6bvrU1yCa4E5zhggQ35i5Dg0GwzX6hjS7LjOJsj7kyUlXee6mpuWht+BHCzqtIA1sP
xSlTQXTPSjGIKxdXvrFj1mi3hCR5JXwQuv0IMmREgi6e3dYmTW8Gtq/Z4jf7pZHoqvOJrpLeMIhS
pnCXNQ5D37DQctAhIBJVZvsYxNYxD1ykm8wdTTcR9pQiI9Jsj6OXE1iU7iXely+/9EC8+VgHHCOx
tz/GU3Zd8ggLlrY0jKtsBFj05OX+PGe7pr57VJe5YLG9PgK/gNtM6Z98oVd2ffu7nS+lYvsIqU2C
xJZcsAsRcXi4Hum0Kn6ypf73Iw/fgl5pGpdmCsJUd5x/puXH0lPXnT6FsywA5UUw23qvFqFYlZYr
Uwu0jifNT9X1TmKmS7MnzdLHkwYaHXLkxS9vHuVD921EJA1XSgetr+ag7tPVb86rYr+XEybvg+6w
ckIcv34iZzM+B938jp4uRNEVO//BwztStSrc0LC8Nf28OpDEQx9CNezs4x0gBPqTESQOEqU1O1Wm
+2CGc/Wh1Eh0ZMRa6U1CAUlcd3/vLIf/iXIozJg5Nk323POmcKVYoBuUBiCMywD31p8IPkmJbl6h
NmdUT3SLNDrfjmCIAFpkUPqd2Cx812k6WvNqbhRuTBtN6BUua3Cy5QyyPo3HvGbZwVBRwbkaB/ZD
aiEXux0nOnuzYpJnpSazQ7PaIMl/VXGLTSz2bzY9vRpnJN40v6YET7GsI6rf/ciUn+MXQYIvvuFq
c6qRsPGi9SSw0fMh/mTOU7KUjDsW7hkjxiNq3mLxpHH5Lgw/cUgS5NykhETFLgJfDJJ/a7zOLAsK
NXisx5gkJu1Q6yHPKaL5uVUBc1GsLUHHqUGwAeYz5FS0auA7qnbUfr8iq82wmLku55doQgyYhPi8
F+Nd7S4gMMnTsosnnRdvuujHdr1h+axgJsXnhjRd+yu0Xu4a18Olq1GiKf+m41kWU6x3DgKrz/ql
P+X1WUekLa/QwrGWeo/8sG88PzvZ/6EpK3uuECylIXmKphVuFy4FY1v9+zT1ekNBIE6kZBq/uZX7
L5OXA6wOprm4KKl5muJxxCBUCGEiZ8hDyDMJU66ix/Kn4UNu2Q81TsPW6PJlu+GuyrbU0S/ivYU+
IdDIGhRtFPukEPrrGxFh7+6WwlxOWnG02JAXwheLz0nXYT2Zx2NvLx9qbsnodmRkldn/KWAXO9NR
CK0rD1CmT993B1zQGY0wxxvd4dy53X63yMZlJSGTCSO1DZZEabQ75ppq+nJQAfcn+bA5izey/IoD
LhgU5NcSNtjpdV9+YMpMjazkVbmo1edVWc0UcCkEDIV/gtvuYKhrO1Zg6niBzN39S9iocoTOD/ed
9douKyzIqJc7vIcesnvEtLASaj6k14Mda4rWn0qejTTCjZbSvBloGZLeGRVvXlgxqwCGRGLXIhru
S7Y94KXax5qwsjm2JXdzI0HDMab0HVsJACcj+Cmsgk4r31Tw+6aJ+RDx2AMZN8l0Xm/T8HbtgEQX
ZgUhV3/H+pwDL5C9/shRno+exNO10A5AvZlUtXCHrW5fdnpozer5ChevxAWN2nluWYyh4OWmO5U2
N1f3Af1K5UEsPBhmIU2jUeDrw0XU7xtiKXc6A0WKLs8JIooiIplhOnz3XVrIceQXAsKl3gJSj+QD
YSphtzFiHAfG6i9vaeZGghi8L2ypXuWvFC7Dnu/iVtmpoTLYQ2GfnBQ/m5SGXkb5I3GCwuwqRRef
nNN6ZzQAWxdHftt/nVprGmqJ6sxzj28hIlfYsjX3cQmTkt3Eo3FZc8k7hvK/DezmzHrPUasX1vk/
DpuTUyEbWTARrZQOejjCNMEyrhImLFgYfnqAfkEAOb9133b5HgnsQ/1ji6V8/ugPjJ5YY70SyHMS
0SEHN8hKARPhsVUPKJ2PDwb+wo2NEu4srHEz7yGBUUisxwaBYA7MAvcqDoKbtOZFRuJE6SKZkgxV
2twz9ANxpGMtLAvPuNnnZ7IJG1VaIpBxFvXnmgoe8NZp8bhp0X0g7dqzx6JURPz8VSPXfJisBbSl
kTjILG/Y8TO+tec4FyTC9wK1xdUVMTNlunip/hkDPapzU6yY55V+HNoV0QJBa+sl2duJaLb+60OG
SJnjF77KnryH6+Fw8TnH7POR59j6DOjZeqdROVqMNRNzlkQ9oEUNYv5NEwomlc5McIZjuHtcqNUN
RY2m7oocHFqGeGceuwWXVlM0njerS9t0rBMwISZC6DXcOS0n3P1OrswsuAVFHBHEViCZsuZQqqCs
o/UyA3AkLXgOgcdgK0jh53aHiDitxNFFvlexmAoJiQzxei8PzG/ZLwZk3D2SaJbIcHsFyLXIcrWH
7N8LfSW4x7But6I/rsmrn1u1MAyoL0Aao4rl13ZcPk2gkId2fKGWZrPM4akv0IPzujPwfdEfVvAT
vaKJWeJC0uJXoqZM1yExDht1t47nL+fNQQFXcVkeCogj7Yp1x3hfSfqJMBb3zR6zdzpPjzOx12Qs
6GRAE8av6iOxVviKAl8ZFRsLt7xKLqPy7ebrZOd6JvasJrA4WUvmx0pTUSQaQD2Of1bowIoXjyXE
JnWkjJiYffEUfhQOawJ7hu/N/IR0OLR5Z/w6ZtuWQsoOAggA5O+YP5tI3ZylwPn9AVdHqHfZftbX
AKHrDmFgpTJTc4rRX3lEyDAhLxweIsRWjmo+h3LTeWZPWcakn8HUZ/0awNaY0FywhgTfesxeMdzs
zYcQQQ4H4B6Oqi0QO/CabXW1UNdziZjHPEpL83r7bgl0zG7GRrnhAgjYcgsCoxFHrCfpcE5NSBQ7
1zS/P6LkwuC1+avhOUg3aCDvj2XXh3NEWkp3c7mWNSd/4+EafrsMua0ZVBAZ90W7ZJy58xgdn7y1
bfuq/1hp5XiTxW1bBFO0CLC91mXnSQHI/8pLJ6HmDTIIblAaRizH0RsibruK3jORpHztdOkMTGaS
6sHnF/RzjzJXD0D8HTKZHifDlkXBCO1KGMDZX6qpz3+WNdjQTaHsxX6W5xUPVpH+V3j9cm3a2J3r
rOudjPIgBbSDuXjDSWDbTXQs1XFbnL9siYO9Ih8tsXeC3ekMJHjTtDapy8XEew6ojnAlhYvIhBLb
FPZekSy9HxCXjziiKdtCzjkvlqEe1dqhK/IDnurExlDvGf5G5aAG8PRKeDvifHGglwqjhkVMWQMs
pdink/Jz5RzhPvmEUal80u5fDvZH9tJIpJHHGGkrX5iS/2myk5Vml5iIOa6O7EImLki2VZpTCdb6
6WRk6BxBWAyUHimAbDeTRaZxdTPFJwV5Xn08iU6YmjV+Hqgf3QYcjRbaRAHFB85o2RtP2IPE4mRL
BrLgTx1shTmlPyAogRlPGa8e2YWR0CeAjzJJDb4AlIYkiG8Ld8MYC+9qj/3T5ubUhMwgkkdfW5LW
3wnmDpGMjWZaBzAgldh+X74EfEDY3vA5mH7a3Z2IoZmrPC+vG5x08OfVB0dkmkv9eNj/lzKZBB5H
5FVG/342bon2yo5ynm6jgsnmFaIEtJV1tc3TkJYiTMe8ItdKSwzlPZyIeM8TNURRXZGqIiZuDY2A
QQimq/IsIX2sPh89LKaSE1yFQWVURFDMkI/0DEMJdnWrtub38T+rfZI6J4nhGXo+xkar6Y9eeAEP
HHmhlbGOgy74dkhBs9OkOiDnLQ6zl87Ez+ydnHl61UWWAQ00LiFIr+gKl9E9MaTDFL8KGYZgQd0K
CBw9Zy/93Z304nDPkEcIiu6I2q6gG7dGteuNF3m6PbEvw75rWHHQ40yIQ3khbySJ943L+04vQi6J
f3tRyf8mRkm9IiPzG4Q4rGlZlmqZ2Lrs09eXyROpEaVDhYA9fWoiCk0WV52gxD+WCBQTMkhrYnG3
X44QXnsE1x57m2TuO5ttlpOG5EzVdU9L1M0l7vu/TjSwAbkrQauZ3bJb++mQdxV7wGzvI4Zvnh6E
OODG2vM26pzcbWmMPefojLQw5RXDA/PJOSKiXT/BPri9aMJu08P3oLyJWu/xJMcQxOv8GloehNbG
ICCTthtlm5bsyxI1kXHhgdrKqfduX1pdDpQ/edD1kErqBUGO1Vd9eh7EPWIDd0loChBz4jDX554R
i2HbKbRQGFtyeAtHtYuxBcOpssedUoeQ+poyTFx4MJTAIe+Nm/LP6oahqddgDz9vF55ogS/bCKFM
hFOFEeDe4wSvwDzcAjTnIKhqQ90hv5ZALKpr1zIpCCKuDrK7hZw9rsxdLglr1yC9WpUrXCIxHarm
nVktS7zFvSiIWDfqcRGh7HEZTb3uUAdLmAxc7fS89J/2pzuC8pt9Lqpsdlj4R2jW3yNfgj2sPrxz
uNG/FuN+bJ6HosPUwKFwBDx6ONVO8ZEJnCk8OdR17unqJ1kW8+MFEkHUnzqc1M+0JxRKMPeqKbEw
JT2jdYuvk3GWjCjBnLT3M/CBi2cILA7w38XdbrNcPizje07GPT5PuHUTGxIykyfNWSIe/bCyG3Wb
8TNiJEyIfmMI+ehCy/mLfkq/uv9Dkl4m1t2OGBhqJKezLWI4sOtGVE8rqVwA3GnpOMS4oWmhsIMp
j0yHHYduVmYZNvqaqrGNAtd5bpefr4pXiVWNwzj5hP0uEaRRJALwiiGxJOk8rrKfY92w2XdzaHv3
XADRLKg821kZCzmv/dQaubW3TffrWEtfTPrLx06qjfSBSCMZvLc6Ya3WtCU12dHLd22j0tMZD5io
pQvuBkCtBECyxG6rl7SHaQXyhFuJE+bP2ZDcTCDtoYMk33LAjHP1yBItx5RbJYw141iNnoos0gPB
qKezrj5Zm6p/UggtZDf7aRx6Rrhqj2zH5BW7fjN899ulsEqebOtWnrddt/PPoJ1hu8uMGCYKcetQ
VkSF1rCze8/pOntq2bs+l/14sPj6oJ4IdCsTlw0ZLVe/GqoviTqu9cA9Y+zzAM/cDzduIVBjXOqs
sPn5r6feRpdTkYWh6mubl6xJbialix7Sw6+I7fHYHgGYmQpA/OCcyh8Sm/JmjU85qLfHZJbJU4do
Zic1AAuNHQEzxK8NGezvH2Z0IDZzclG6LpBSVLG/ej9Rpq1X5sr859iIygBgJul9gbS5dazmWkfO
+DPT2da0P0Tq+3eJq4RuPIgpOKDYHdL/gpqYKh/nu5OgHYdvL86upGW536im48KVEoKK4DZ8hk0C
yNodcWSTyGFQuT4zvLFZ6EpRUjIFGJwjJJ7TbfE3I0ahQFkBuI08jVhco1nKRF/klGSlEHBxR47W
YRCMWyIfRImnrS0xhkRoYFkQOBwSWrNGaR1iYeam5mt7Qz6UuIEmD4kWz+Is22e4ojILKNdPiARi
O7LOk58iH5P9LetnSIOgp+AjjFB7sZD0BhNLSjlJq2fAWNxF3QMs7dYB3p68p6PuxTdWhSChE01J
sdS+awhg62kvJzPPgoNcWckmgy66/PxFaqBpBfQ9nbv5SYiix4hryyqnYym1R7Z93871CzvJY4kV
yW+9mt4fWYjijEao3IIJW6/5CNyIaXAAzBtwR7aIkxCFPYZgwWdzuSZYcNXG3HF9aZYKpBolcEXw
V1S1muHemwyjsdblKBLhTaP6GVAjj2WPHQpN/svOWFMNqlTu30cPFbUe0t0Z0HunrgiNAyrZr70y
UeboLcGYXRw2CYIQ5foYZw34HR37htrcUCXv5NAJ3NERfBL6NqFdHTjxtkO+tSgUrEyDC9Gi6y2e
FCx9gSmKK0ga8EUeLOdZtda+LqBBZBBTLnHSWZIVsfMHsHyavY+y6otgDafM9aL1zxBIu7mpW53U
+VEfJ9VOXyXnZFBa8LIYPlIw4oswu91roi8BwfHIg4gOqYNHcVx3ajL7dJ43o2nDxZe45bgq6XBH
uKwZWiBqpNsYQBSd4vu51ILDD8d0tv615VVXP139mWhc+xh7EylvigLtAjJyeFMjAzE62FXlUhsZ
HRoJpytl2iU0/zSifvbxyCw6Z5H58QkpfOx9QhYHSNG7LwlIvy3OX7OKVjuAHbk8lBm2KmkdoMDa
gAUDds5xmUcGY0KqG3Azah/xRmIbUBr08DCd+4jcahklFG93AgY/oLtzxZcnY5+tAmFWU8iHPhLg
WPusyOuremuw5lbFbyo/gqNUxCSRgkLeAfwtCYrgNllKg0Tx2bJ4YjQCIZwrNHOCFnLcu5r4bb3z
CKwWa1N0vmbrPYAaOOq2y235N/5uFtJ0tU0uGbGH8qPBQe4UI7E+0Keikdsxb59K2l5U2nSIWHC3
ILXbAFab+ETJgUlNgooypXzrjcxfaAR0uTvIYVbOvchV6w0UMcsaPzMAxBw1QCvtyVm0Fd4lLTaU
MCS6cq5m+SayXYQ7CPE3mgtWgqzNmiZ/L1xh/pVlJKJ2ANC3pq+5UFQE0nJ0c5jl3l9IrLxdBiQ4
+c8ct1yD74kihae3YJZdlgWKYWbUeJ3H7dpgDuDo+dxTXggQDetFFpAFn3WnC/vV6WXmSK6VOyQX
nyL7w0aEZgr+kt0SoTJKDKTyqDbZrA5NlQTXIBEOJ+uHcNl4XLTui3K+AZMtyRcq2CkAMRyHws5f
XgiPWN6BV0C7uZi7LlfG8nkT1BsmT9O6zwCjaaKX6IhgQ/wV00zfOj8/up/DKOaPTkyNzTM42yil
JHXVi8dHPzxJ0Af+STzMaXvZQ6jTss9qhnZCWu7mGQ3OKIg2xLFvNvq3CODfUp8pfGEQEOtbKKqz
xgFbtCTREfabwlkJquPR6HMqxCSP5dOygVTfL3oUeU8oZycY/sq4KssxpaBO3Jqq2D9mo7GV9WKo
z7R5XYegHcmyiqBbtE8kpT8YzwONsHaxSPwfnpdSeKzAQBmY+1FicyDJzee98A04Psfw8D3FKs2K
1kMjQjvl44mhVYlzcACcHX2m5eaboxxq9fQudrHGnBYCNcLCty9PxqHjuLuShebn4vb6KfKYDcxA
mDv/wz6UWUL6q5RXYL0IJgSzSiMZikHznv0AzVmQlM0+1PEW90YuV/gYje94oDPy6+v9j2A4m81b
YDD4lt478+owxyZnbmq5ikzDfnDGWwgReUh08RsO30Q2q//UrS7GZXFqZV3pj5XwXh4CSIJCbKXO
s7r/zbMcjmS1JsjGnl5fkvQq5mqUp8b8/JHjZtOyDd7Hlis0MWV2+tqUJwPvr+x9kSUgRLmM9PHe
xjX9EGKBq6sgdePe3coxgnbI/br4dAWAFTdWFmgt/92ZnPDrt7SpeqmlNhPra4NYyBPtIDEUhfIY
Zq00zsL2SWPI7Qon7+537ogeOT4KTkBJ2IImScz2PPY4KGXw5PJph4aRdCXrNRcCdBT1zWF2bf4M
vuRu8x4mg3biw/Anj5CHtTISqThYH39P1v7Thb2a5v3qovGdSG3wCZq0ubhWZS0IB5RIhGCF2dDX
SMxuNk0jonCJ+VZcbRhnrOoSEpbMHOxMXwhFsJnfCLJwjOknWnGkhTakaVFiP6tjC7eAM52GvT2F
bj+i6h1VOfFC7bLsatMryPPsnxrJ59uCKdE2ZQVgdZSgrnPejUG1uIe8PmJpUAh/Clp123x+ujmC
CNmRBqq6Cj4r/2lVmuqACpUv40VCQt3ET621JvFPFlaZA3tQ3MXRCiwdcjnajO7jXhuNjdGENPua
mNVCAVCn7zZclHMXM5ZuHCJ+t2e/d29bzbhCn9osP2PI/h7s8KKwXfl/BxyWcio9PRC4CCUjJ1Fj
NHEnDTXvbmAaFevaDV1YN+j55TEsu2fxZt3yQHjgidvEYMUbU9OHqXpn+n0fQubXr598f7/z6uJV
VdR8gZn04+44bok1xf51+joCQwZmvBJPJ0csn7d2OhiOsv7uVE52IjhWM+Rn/pr9046ASBNOHuA2
Ko2SCXN/QQyPkXezSpRPOfIzblTxhYkRezh6bHcRi4NJ2x/Ty92S6qhro/cGOaaie0oIg9nr52cz
Ns5DddG86T2fNrv7tNFbO/XlmEtEF9aGCSdQ0FipzPbsKFVqhkT4IqkyEcDzmEfznF9xDscA4/97
VlIfJcXN1/eTrWLER+F/dWA5NyhYJJFaPh6HGofyVtRpeMdFELkKMk1+8XGrphFcDRxSaCAdbAbx
6mixkca8Fp/dbeOMvXYgfeO6hor7o0XDVb0+0rNhrQ96zEyzB5AWNjTyZj+Ln91JHsUtW7OoxfOm
fiXMii4ShBcLbMm8oOfALHMT6W4lAZQUf6BxnCujer0ft6bbrxDuRvddv04m5gN6cKuhc41ZW/OW
+Q2liNNDEM2EaNmE58tsrwNCITPi+o5HpPrdCLVol4MovqQxTXoYvt+an4avunGsdQeE1TJrrlU/
mObqQuyxZp+VCsPJlFUL44UGpAXZsfOpqBe2HuDKXUzOO/a7/LaH2bp4w4HQShT/qO/DmaFjZpm+
C3u5+wCJ22O+zOHGzau29A80FxWMHjIh9lPq5152NILs8sExhzgQ1Ul8DTe6xCIyWiZFk+/Hodpn
ASI3yunzWwMnPo4Y7dljy2DRBippbrE8KDnD/8XOb4PIwvcYYxfVVo456Kk5n/zo4KbKaaflc6Ox
7EQPkWaeovI5BVvMtLClHgoF2v25i2bHRgWfi3Pc4ew0sTcQbDQTD1OH33WL/rKkyX3abatLHlj0
aZg0s+dicFl3xx86YE74JRAfxzaPlX5IvgDI9RUAQimGeJEJDTKoD2TCYF6p/O+p43aWkV9lHL3B
spPb048wyWSIG7zGcHykKXYqxf2u+cPytUGEitSH1Ey8fubNMfWRwFDfX/fsMm+h0PCczqw+XF7T
gdO3YeiosWpR/lKyUs/lnir/RNLzNY7gbskvBVpZhA0CcivNpH7As909okylhA17L/oto9a6FhRF
6/rWMupGuVvhbkApTGZ3DQLIw5Alw2wxkXKvb5qFr4pGA3LvlYt2V6hSA+5Ub7aPBoeWfleKr4sY
ZtkczbI8f/iDyexQw0Urkq8YLT7qULiY5642kps5cZvgwIfwBTIqUoCyV1+EDgzgn5wYPOKz5rht
OlFbAX4Q2YFqQtocHwDILkRA/G2h7/JWZhkNQ6Qu+9nQmJi1vAtYuEz3fCny9SLEqhtI2C//hOW+
dimJ5f5qY8XX5WBw+S3hVDexh+xEvqpe89GZavDEddV48g1NpT5/hbr7yK8FgqP+At8MKH/7GPrD
v/6MB70fvKWbMND7tLZHoYNN8R891eEUc1q/6TYUVpurR0FFXSz8XZOX/6Bqr5qVDk0rwBQ8OU3r
xUC3cG1uLr6arQSpnrDjOnpI8R4fNyXS/udzf62RC/LPYW3qum1XMbnwHSYsQnziaN2WPrMQrons
kV66Mcq8T4Jy2B2qojQUkz9vKdkEBhIQOofhGHzd4XELNaQYnK1KznxIc68u31WziF4dSYyejL+y
jwOpze/sOM1sFpy0pysWYuQEHheYYiczFdGRnnsr/D1dIe/Vk26NxbGDwjAx1kDBJ9BBZROBRzEi
iv+62aO5xIaLWORquCHmEOMt+fuSBcjl+RBRy3hNdikaOoPFeXwqCaUNOHCxQmY3vUu2oPHl6V+P
2USvrzEWAfOIa7XvsAok47LymCYAaqA+R0zkEzu2KbFSRgMvkCWUO8a7JFDrKoxBXs15TRrviAEL
m1hEldJ7y+OIeXo88v5X6m0dogWh+Upv/TmcZ0gKAOOE+/DTuk3bdqY1VV3DEQhJxr/ON54Oincb
ccExPut/r8tLcyUF/iTcu4q3PbspHE/25hDaT5jwtUwgP0v6pvwIxYpA251o4FnfTAFMxuRn8+Iy
uAQEWlcVynx82dZYH8dTpuHKzZsbMQLV7hIpXmMfcwgjnftY5YQ+lmnDfI3CxjvxzT1/krxhwDS1
roSARQasDMGYs0TZE93G2XWmuAOY8LsXGV8zmbGvKiTjU/BC6Gy/M1ISYpCTjCDZe+PtG/Oy2tkD
N89k0mdZr/ivQptW48pk6gjD01YZctcHet061s9IGn+6AqiVn7GqTOEggI115NhRAS//npl/QIWq
JSVmp93fzISZfcRvIZOeHjEDJh8Sf1j1zbgxp0/0kDw6F+3sKOAi0vk7LqKyT6cZvVGoaTnRxJDX
Yw3ToPKuAGDsv65i8l7rSbPiopXcI+iwMPgH17bRycLC+WHGjNVKoVa+IEQcfMWTx82ZbcvGAB8x
kCDsYneK5vSRecbgdBC4EkEIzgYVNDAbYZcxIQurSVA4MsFrJFs4xN4dZzcdg9nL38iZNreHKCcK
sQxB7R19Ej17cL0k4BUjpVI+/CgGAp9P//wK+++3slF7Q19ZVR8zvPHKsxsnwSVT7vu2gQz3A7CG
EeenJEGr+fymSshnvC+1py3CnctI37P17Rue2B1RnYuCedIeQnuvC6G7haF0E4HCrN9ytHN0Vo23
RjFt5f0m8oCrjNNNDkrz6cgXWfxUyIoKE6oT0E3+1m2iRlR0dPlqXWNBj0Avg7BWCO9Xycl4ejyk
wW69/QX11qccHzBUjANtXADZlow/AGeXBFZ05+dffSv3rZ0O6eGO+butstUITTLwFBjZIi61LUKO
Q475iFyYjFDjkBKncUBopstJmqgGEHGivhUbezhxY+oyGMNcSuh/9L8K7Nh/z7syno2+XGgtBt0E
XKVZ5CL4wYfbgi53QNIjf3zYzGlaKt1P0z4sf+g7/L84pcOPpsy4nmBWFsT5Mlb/58h9IHsdVkNa
pdjRbskbw/LH4K3Kv/tBfOWYXLhoTN+/byVYz22kaJTgh7bpLWVPPfx6XWPZ3GQphy9UR6pEOul1
rP7LgCUROSW8WQ+Ty3LPRj4Zcvj3BLHjiac/GuYbF0ZbJt3Djlh9p2Rw9XTZEUXVhtmRuOQV88yg
c/kMQgNDAKToqQIfAyfvpphK0X8fHUwVrJ1DKiz4bAEvu5Gqsco13XgiWZLq58jdqBP2HyQ0I6IO
uA2pMabYn8HuiVvU2r+LoHqkxz9TBDnxec3WEOGEKHTQlZyXKzra1gEuMz42rcSAD5fu74N0eLdr
NZscOALhoOAlcR9yQUX5w/dsNyV7lzTM4/rbAlpVI3q1PjKs2Y9B1WGk1JdaMsm/qYb6sKXnY8z7
dPt3bhvbLDOBGHEdVTyb4KNzbKxG9y4NZFmHdbs/W54HXxNhnkerZtWHdQqRnOXly7Np1k11Us7D
ykLXOB1iZA4H9Hv6nhEw2rRDcluOuNL3GFL21G3wkIdXh5x0iWpKfK/6NKpaB+VrqBxvSDB6xJmk
4zlLT+JfWfj7I7aNNqiJWNVWUMFGkqt0E6k38aDpf9C+ZdCbOMmrch5fWRMHBif4OY+KpKorjZpx
Q2oKSnVRJLin/ziEJ6EeA3rgaexU5avo/8vx4jgWUDqro00clDhSQTI4r+W6DGVd2wFgm+hhH6Fr
0gYkbgdsHfL2Ct9X0gK14bbl+DH58o1k4a0tCTHgv6jpZmhVCK6P70CpylTQZiIJbWlxH+JX+UH7
sb/PD0wYdR2bmHo+nciyeJUd9689ypZY8ePvyEfiKt5RUPx4ugQRrpvVj7xmM+nqsNBrM8Ph9kOy
JTYvfFwKPKiTct0TtlvTx3Lj66TatblsrxTCAsEi0rv6jFTUAOg33UxxF5kWs5lYTzEteNr+Lvco
GSkSKWjROVtHEg6OJehE9TndvlMpgBns58cI2jwYXuRSV6h8+jzd/xCTI9oFWKkSEIUThU4MBhLa
KYcE7bTtxijVf600Ilhd2teQiC6DqgoqBjBc3hvfxyv2+gLS1W8UFdCtoQRsJ4o6EdowNo70bNts
rfr2B3vLX2xyc81EAswBphU3VMB5q+aknnFanVdlxYmry3xBF6t56Pyh51bR1RoEFTnyGHhdu7Za
OXwwVStuQx3XG0BF3RFf3v2jiq/G49rTxxfWM+F0u7J91LkOzil9ynWCtFYaTmuqXZzY7A3uFplO
6eU1GppnV7cMLM6p55mPg64RVxuDA9vzwFqvuEIOSA3ZtnjltKxHp1EXq36UUPHlQMvd7KY3gd0X
GGEpXzW6GOxOewTrIlZhB5ci8nNcw+Kt9cUcwItM5XLhYHFRwVh4AyRDuallkYRfH1JdJD+PvEIl
Y0jPBODNiyflpiwbCVNLMf0vComfX/kX4wqon6/GZuqtbW67DsGy8hTofwg4cavPF6YfxhN3FhVD
krmS45NYgGtTqG5vDNUF1h6GnHdEDJa14sO09uW1i0zMG2pioEUphGSJI6lHOUYn4bESJPtt4Fkc
bB1yp9Ewbb9yB+dAGY2X4l73sKguodG9GGew16W+qlCLPKfftBsWK8cd7o/8imy/ym2r8Oa5BefR
UPU6+pET0Md9zNdEiBgonAmDHJgZiCnzzLqDTRWY4FxFN2KqmJe5HjP6aqTOXSynoV/Tpp2dgqZK
2hgOdzV1sZs4s3K1sjkTe1p9hJcJ2qXO2fHS8OiTVBeSZsyW30XK9OyPUQjEQur03SV8VUOOQhgK
fDR5YGglBLa7/BInX19oySnyORv3NFHukWPhI8zhG8WknozwgjCVHTcxV67PAYHUFZiMvrup9IMR
LlRIGAxCZ2S7koiek1VCMk7UYqYF4SAAUEwk5h1DLM6aYhTZSMt6LSZhl6F2kok8wJ9LQT7FAc/R
n+WzagBMXiW3LT9mTAUvXiucehh/oEy666qDfKUfCkBmuhjC2GaD3AWR7Nb79u4kmERWIQSOCa7t
5OWyrbM/yUDWXRulHDhTL7DyxkZ+fV1OKx7NcQPQADidS4cl+qJxyu8WMG9/cG6NtpFCN5nhwf0Y
TKLm+qJ9hrAa+Q0YQztpRGWe77a/crlZHVVeshLaSplS2EFY96LCjCDgb2msoS2LyX3w0kmv5Trr
fPGp9gq5vF8LXwyfPUO2PbJwbEwxnEia5eKf3lkm2x3/3qAqknLDsXzKWUDdXpaXFyDZw+GsaK3K
bcnJ10Ur6NVuu8abBXh7i1X/OFBE01d/66+eTk701cwdGly6iQr1ZiB026WLkBDThczxcHv5d7g0
cTu/lUjcf5dHSfAE4aipTfQXz/Eq1uKvowpwzBcMLaFti99S0lQwLvAXdpwjaYltNK44rcaPHbca
hxIQFHH8uxqLnBYvf17RQ0cC5r33+SiCGIDdr8iCdJ792XGFKC6YPCU4PGLCPKOanEYDgN/0uzpe
qmoaD6eB2PxNhHxuqd6ta1dkvjtq8EeK2rqV07Z5B1CpFKvXikHJbJlJ7AXuXO5DrOcvABDYhMpS
yOp9DY8+a1des0wUia99las8DQiqYKiOa5t4AUYxQVColrI9afgztk3ozv3BGBEhTkOSGy2NVDOy
5RMUD8AB3quO58WRsyDEv4dSSK9oT9QvN8y4N/A7ucd24Buin91MyrDgqtx5w12P0TI7GBc15t3o
u21WVUM/PXwQ7UaBxaqDRpz238TUaED4nQ+EduS2KEgzBSZPw2zS3s5uTCR2p5wX5TnluEQTCJRV
zqjrqmF+9BLH+q5d0g2zZTcAO6+UoCvfy86Sn10gvkyk+qll/J7exh2L0jR55cZV11nz0g9kKiz2
Jxb8uDp5SHJFDEiDVF6+jd/id4a9Dt8g5/D+Z6iXQRCJjCPPu4T2KK3pmw+l0Rxg8PXmVxC7z+JA
okxscvEYHMqiybfviYB+Ax2Nctuo9f7m7BPSpKlP62FuXqlEiMkxTzyaANY/P9VvrAMhN9nMXdjq
2ArIC3pDyGDsl+A9dBSd6AWbT0RTaphWKbr7rSXzdRKNOBewzTkAEYq3jhwLd+hpkBPhh36WKJyZ
BVZGPOMaKZYpwIKW7LqRW/KMLLCroPBNSoK8GXGE9gThD8MTkL/pLgAF0RInLoe/jBafI93vHcas
xf/LUWfC8USOz+z9UvExENL5tQoZUODTNiExLtDdd2PqlsgY9Xh/ljzGeMJc2g5ayS0DUXnTJi28
0l4XKpMavwxJGqY2hWJ0k50clFVezo/YA00b2Ye/Q7d7TQ0e4/jU+wOLsTTpL1Z9tFMLSFUAFZ3Q
GdrHDrz/GSBy1a1qtQl4MTxDEjdXKCAJUkUpI5GhzlmsfuQi4oPKefHkub+iMHVpHVtH4R8VWl1r
NjFeXVNGhK35fIjfrfQwxaURerON8oTZpPS69RMX6KqR/9jHddE/JuV+aZPFheuI1T748ea+63c9
Qxvmq84e/5MAG5lusaKZQafUUNFoI6gcyNqHNfF3WgbkcZtTD5DRH44z1XwqTsZDXsLiGJ14qrxy
gj2UREErHWQaopN67Cmg4BWCj7RPvAq1+FZEhJxunVmK9/5ZKwLfDs7oYgAdANYiHHghfTEWnFfB
WMtk9tw5+YROjLVgECKCwKJupqZtZf7ESsLpBC5DP2Zl5EImvoA2yqLCIT6Nwml9gKM7kXpsjnuO
iPuLAOL+dWsimpjfPUejrmGZjixTCGUEuJUiYZDBlYgaNjnKTdZ+vSRJgK4AFvXG4FmbH+fuDpaP
iybX9GOcBlOwH4XYx9Y+ZnlF5vyZPslSaU5xDRfdkEeJWOAznftcKQB8RsdVUnn/ywO8K8Hsh/4l
W//ne7icybp6HCYMAkgNf0IFeKIRi8Km3DCZF4itzT98N6yTirzWDqBEGKEWEFKTxskG9k+8M5kp
Hbb6PldmxXM8jRK9Kg3olu09w2LDVNGZCmJs8EV/zIJwkrg57dHdt739iVPRH7d/S5QWhG7TGRTb
YvIzDmwerfVsr4bBie+YXKlDlMsIQGAAFjvpD8zecmRXQVSXU7/dqu3kDgWSgGKF5duqjlGx1m8d
+KKgkTowQUC7uuEdVWlVHebVc7hG/dvSop1+y42Q1gLNBuz6MommA1AxC8/hdHlufuxM4QPgLH6V
qHheBrZAD0r3nJ7AL3WJPOPPcN0KWw4Y5aOum52h3q5O9iiN93lroRcR1rHqzXdmLDStAooqOlbU
zYWIq2fFBDqP+lzFBd9JUttdeAUmZBXAfuQPgwyVGmON5INfV9lGNeB+aXqbVgTvQXbSJh76LGZS
52166Aot87N3gXwqLkpI4sgis3AFHiRL3yshPlrR/1La/TP9ABEtTKfNFbp2EHEm0AU59DKc9ls0
3cg0oM9kbh0qc21ttxs1DEDO8DRkl8nC613lPg7G91+UEO7PQhAk8D+WBpX1mE24gSz7E0pap5qL
DUTZQTO1rTiZ44IgjTk3eMWlbJ2PfrRVZhV+XnkgZU4Dlz1H8EkljOmdo8pkk1FrzXxfgIs3azOj
64u7rELm/7W6cFKiHcMg+CM9bqMWswxIWv9P5SqmWqdX/I2fDZqzGYoXyhpyo11bsaR73qx2if0m
Q2GILdYkz9w2mcUwemEHoKL91NqzOcSAIk52hdPpWoOxy0tpB1I4naJAfoFQkxOKrI/Fi01+lqQ5
TGUs5ZRQuh4lDe2TQ7iaqbHkcmO69Lz/7rau1nXHCK6HB37YatUL5D5btynRJ3tYGehDfeoRIUoI
PJ0KDhCYuF3WOuRhfxvFcZRwB759Ta0v3lg4f0awuAqycFjg0auPq0AIDP7FdINl0FCt9QE34lcA
Z1/INx6uA0r9liK3XE5ugFiSH9t7c2Wy/nD+/nH5ATOUOaR6jUmSzs/lZt3uZBOZTjQku3r7LQ09
WWf0SMXtz6gwt9/mxRxYWpYFpx7ffhYUycIDhSodOOIgGzjwkHSd+AqvnPuQPoUK+6sZm7+zW7pv
N9ixMqySFwLhRdrxT2alxMDEWspQHFdOqGkX6DuL646NDFokIg30tp9i0cpaRSjjjkZB5byqzej2
KAb0rJzzetjgm4wO1Set3RSPNm/u11aQDiuDJs/k4UMyRNxrOZPOLrtH7Ziwf4rZzUuvEj+cUPNn
Rki/OBd1VTJAaNnBkOSB/ILG7+TnMjYK/nowszY3R4Re0voP/9gezxPdtYp8obgzui75EtqB66py
2Fq2rR3cz3eg8/PKTiyPuSNpffzS7MkDPLCCEkpZLEMItlWTuRMquYk0tkDatIOoC9b3UNQ5C0ye
sCJNJ96Htc+V/VEMkOC6GmZESbR2Qo/8/72IaThjATmXbH8KidUloZpv45TJl2q9PZkmr73FACSk
R/3yNPje+56ApIlcGOn5PBvWUDx0CWH71dt6Wo6TTQYEQp9xYxuZyGW6ZF5PQGi6Q4ecd1I4TKn6
lTiFWDdVQaOGqOq+0bInTPDRhGUCBqKG04jTzZYXJcAh9yGyPUpxlE7StjTxRxK7f68D2DYkX2YD
323UKJTjlck7Y3I0bFXDU+mkLBzpzvTvFi3WdFmhsbAVnX2JYhw5WzInWZk3BNEyhAK5qWWbh/WA
o3rj6eCoKIayP/zoNdf3Ii/F3sVZkAjwrQBiEselAUOpnVXon+i8rxmq7mjUYmalTQKcws/7YkA5
k6/3HndklhnrHWb6xWty+aD3q0eFtLm3mTnO3R4nkPaxA5IcDRTxxnbv/lz8JBA1rX4pf+dZAHjH
qXNVgS1Ti6zANBD/FajC35/AdznU19rz9X8sgmVO6pZXWTPSz8qqWNKmUDRINln6eIUHVEyjMQ70
1CFN+AOOkd4oImGrlgTpR7u3nwl4GVSfxDGl5SYQ+6mqKMqtnSS7X7GTQarUXLxHXOWHJMZBuI7O
FZ1orXk+usuYardIGCijS6wiesXoF1ivBjFqgva5mYCytA1+eN/5p2uNfEpZnSpqYPJaMaiUVxEx
9+mlJ7fEWVyplQ/kLG4jVO9/SIwUpmlFX3Hsrg+eB9cknjIrPg0ZUHp1tbBL8KP9XJZcu/dRqeUr
pd/Cjm6j7LREx0DC00JprKAvH8OVlRwahJNktAL8Y1fdlOogb/T9V3RaaqgOUVPWx/EO4Ce/rfu9
SDzSWA2hhmzl4FVYKNE6dBRRtT1+oCsqB5H6hmLpysFPVOgs8MHHtZcZpQyO8HOCTkUnjTeXZYkk
KIcHSeitbFdYmMC5w8Vu6Hbj2dx/XKTL+qwVsUi/wP9RmLRsjGBIQgY1C8eCNplwmfTuY1cP5Gbp
NNbCxRv37NwxzEnO302FDMKnYOflmHDEV5VPmV6iHg8ZiOz+rHZx4blCKrwpwovtj7vHq3IpEW8c
cEhlMk9O25uTgMPjAYtv0V1mChzotViydqW1LXIh0rx170v8IYooOQEm0eWovjK2GanqRsuSlcHl
2tDwyVCUHHkxeifM1XE+NloaqPJscPDLxr5OH3sdqqDVlINkyisRolpuWPCThUaibnHmr7q6/ALg
b70aJ2mDGXxEt4IlEsJE76XtWsWQNeVeMbrwbp0fldGPkko1GL4qow0VMUGqIICyBExYI2L3+CLY
SwEw7SHuGbfwtatfbvvMaBbuQlYT3z4j6g9edrbjY1vm3GOcIoK6Y5XD+0/ljEJvuUDjLa5lhpl2
HpCWL5E2S8mIg/IQin5amA6RqUL8CcHj5eQggJ7VpnnNKjIu/+tljGlkBXctLKaIKXgJFfMrZFbR
FcYw2Q0c5AhXwqxwtx+CKggf2l4QlIRG/SBVLDuTBHlaQKxuFOkYq6OBywsz0G1h1F6xt2qX0eXG
tavoiUMzgq1oMqjAoRN16izIVJEKPMpg5/1mqDhFigfkVCQwfLDteqF6hXRGIx2pfELzylHZzkU+
ip5sKJR08+ErT2aXUWXqk4GDse1iqDYM94i6d1bkfvaHuCorEmczPBdbLyv7/AY3BIFlX0KCeccU
ornslfGblMSpFjaj/MaX0rv2NvZM3So0+aTHWh/aQY/Lg02dp2pGFBDdhu/GMTOa3wrRMJF0aX6h
j5hAwXU5Knmkrfy6D2sAAtxCKC2ebMFQVwfi9yXJkc3ryEyadTkIqkKzuWKliZKeWVtX4CEGpG8g
20VbE0A4QkDJ2qjPUm2IuhU+BcMCOisBJ833g33sgywZNpUu7Fb6B1R8X25rmOILAgMEchzYXh+w
iBWRloX+BGVWUneT5vP9nbmmqrnm94LglRkkpwVdG06heNW2zCWWDPz5jD5qsxY2BV8crjcJeVrU
V1gVyP/UF04mMo/44HsIBZZqY0SdPjXEbpL19u9HxhYn0EV4xWq4/+DrSmzWtRX6VTLSD9e5vfCj
2XvuFuS9XrlNXW823vKYzkxZpsVZPhTo4RIi04aDtmzvrIMuNMCEAN1rohc8F+JJLhBnDFmGslYm
Ox5PFASvEy055sTp3ZZRe+xSoP9gm0nZp57bAfBBlJS4j5p4wj2NwHNeMfqhLu/pqv/1k9jI4C/2
5iS/JDW1r+PMbZlFH1Lpn58wUe11GB7Ws2voBB1kCA/osAu5TUmbdmeXPfnFGWH4Nv4945QdaJhz
YQymkbL8FvdxFePkIJCyqufVV4WoQ3fHsXyxYIZGzCNPWSTNS+U0Cf+Qax8zvFL1ClY9PkQF+7ss
Bh5eYVB5eIWy4HNg8KawtTl+O7MMjXp5UR8KavvFH189e/WtUv8mY2qtCouUz6xL05xkVKAM6p0v
xuyqFlsM1fboMtw52ajAawpUEV+sLU4OacnU5YY2l2Z42C5Q8PJnUU4I80drrazGsFY3UzVkKhOI
O6zc7WUzkVWtKyIXkM3XOeKNTpu0JBISOsAbHGZVosNqG9dQuyVSq4FcIX1ElPSMG1bV2JehDOco
a2kcElumUtsSmCHAT0glkz6qYj2zmFD4ikv7G6SQT5ElRPN9ig4RNMxeu1y0rAPXUZhWXgGFEvaH
k42I9iFHF4yFyDwiMi2JS7noEOKSlmGjRJHlSbDf9sNaHdPbVqM4Doeh6EvK94QwIqX65DzfcMq8
tt9vJkNEYXDnS4lluIyxMuP9YvPqGCVET6cI+9T7qzfJZalX5jHZ7n6PghRLicrPfj1obwNDpvhf
Aduk7KhT09zxLlY5lW9YB+6oJ7/nlyKp+H67nEkkLDV2OhqsVOfF4Pzaqp+vggt6q73T6ll91hiz
msp+shofsKrzQyddohH+c8vP7d5YL3NZz5iNXen6taAJW/awXk63+zsgO2bZrfRo0zEQFVErsByJ
OpeC1mFCXBZUGQumqaJ9L9Sq+1SGfw8iQNMV3RKQ4Y5P6qWlFPkBJlIPA8haYeRCF9LHznwh/XVn
4ff2OdYGkZE3J3fq2UGxgd1JdVaNFuMPVbMQQh9OnQ7zT/cENARMU+UbVuDRMqKgT+S6ZyxJcpsI
cypDWDlillDU6V/r7JJS9y3/dG7nflpb7QRgdanEE/TQVRU5SgKTDC8u+fFS7zj2DdWEdzbiYzEm
rzi5hbFKdbjYdi1t6X2kV17vRdTgs8lA97Nj4XgilBDyUiEZAFODXLmgTRy3RSgkLD66/Sk0CY+E
l249w43N7OWdVMD2r+UHHoKQJX/Ajt982dVqwAZ8QDXxj2F0lkBo+n6z3sqqSut7EsXKQ+jxym3y
LLXHsX8fjMpwE1CKMhCbIzOSO5lrhzHjzOgrl50Q8oUkcJ6ymvAsBQZtCnR0aA0BmCMz1M3W2dGH
07qz/7gloU+x3dapswwrwR9Gm6S8R3qkLyWJ948lg2XEoVihK08P59SVJKNX/m9+I43WzCF2AYbt
ay9CXV8HSOFCXweie6/TwH44/0YIAyjQBhxybHIgsvPIhC2mkfyQj08D7/xIOi5alRbdIegbFEAW
5iAacbckGxcNnL9aZuGuC6xehGFEpI+1AfcLRB6+WIlsX179Q3JNhXh61KbS7xt6Mq4tnVW9AV9a
qkXj7vj/wMzPbA03Z/r4+kzPFErFONjG6kzdDOpp+HXxVOMs5wT/MvtQ4kNZO1Mq0ENqqovI+lsg
PdENnDApsB/mimVWNn2MxD5Pq1n3W+sJvt37IC5hvlqvqPt3Po0O3HKIGozlAX43k+OU4QguQbdC
Zob0DT3V+cBXsDyOQRvWudTN2eROEanutHBQJSizUGPX4AOtX5DM+zwGqLc/Fr18BvCauvMrYkI5
aRRkzrZErMY75T6DTta01xYFwchgtPwfLXeUhHbwkKpxu90M6iAaIUH9p3aHX7v3z2To72tfQWJB
vnX2A3u4zOue85S9JwN/EB+06NSXLM9azzNfKp4zUn0Dgu8IfU/GV84ZwC4Ro+mTLZFtgoDAZnKu
F11kC2DfhIu7nhqb1naw2iz9TOV8akERBXva9h0oohs7u6zOYovxJ0u8XCIKNNOyTqiThP5vkjME
6QTGa6dvssbGjz7UPz9xqFKbK5jtSMNAC6HEbuFs8dZfYeiID7huW9RhIn0+6rD47jh/55krlZPe
7Q9McGUK+GLxXP0kJa1MguPICVKKrx2a6VRFI7KYeFV2gFEW1OAxeo/gfEgT7dP8L3KHRhuuLl31
/BxK7AxRuMpRhiOPicX4viQTv2L0rC6M18J6TRc1vfUTlBnypS/EueFpgGQlnzgJb6teIu82Qvoh
ci/LorLxqENQ2JeWC+znlv4OBoigTFR1udHHPvIhX3Y9zMZY6aM9gRRFSplvPJxjVCyuM9hvnNjk
kpthKKzzqrH/ISMK+QhDGyi4ggrBYPZmj4PaVGrtM2u5FtXaLgw4eQ+zFWdw5Iqiu7MX6RxZWWN8
azT9XKx3QXC6OmJJ5dQUEeHITwrbFPlfLkPNycEnQA5lxjs9Rx8U1rnJDxrRotl5nwDXIF2esX4d
xBTFDQI++tv6xLhGaCjtmlc5YX3Q1DjQO6uPm0XdWm54TH5VHx8YEJ+JzrDpSrFx2IEt5308wWk/
ritnnXdmUC/7Q9Wa+aAAPy+1J1FbSEib4E77+G/jkpExqENvWDFiuEzdKq6dzg9jklTWFWwOW+dV
eeaKFeCd3ukrXSO8UAJAhxHFF21ZFuKI8o/XjWmzVdbH0j3Eb9h02GLr9CtFfqHIvCX/00Rqm/zU
IcJ070fYMwtN+JBm+LarBZgfncp59yWpxY0S53LgZryDGstKx/bhwb1XYU68u23nzommhkQ4pInr
c1nzMzPGTp5hh2cuPRFF0Hm4zVV0+U5QRLl1iYhCcZqp3yuvfBtK72pGPpI+SCr6Mk4oM4O2DxwX
we5AiA85L4PNlRuVNel05n41N1vmCNmbOIXuOXfTcuhBKeXu/gJxEe+4dLNtIPpGkDHSq9QurvZG
oz9LdCY8nuT+bj9ucox71+4j13mYhIjQN0jsQte8n92JdPKoR0MfOPjOpA11sUQjeilVB4brcLCS
Tja1iDJ/9odkC5uBj/wL11r7+ohZNoA1Pc/HRymOgHzEJ4d0+HEROhYVsS9Wed8N4hvUkjr+pGHc
pxAZPfrfwbmNkF/9oFbxtmoREWFQniAI2dSQeJ8agajLM4DV2EHiCTXE5E5oUjQVuFNTND5vbFVa
fJ4gE69snZCnw/WJckSN88q+kNqcXC8Epl3So5YOGQ+XNV2VpXt+YPjn3alGzIV0unkIbFJ/uOry
xeOH4ukL7dmFOqC67XCbV/ijJzG4IYXKNEyy7ycSBeg+yOsbeMIEyrgFeGNPGqRyi8XDh2ZO9dlj
knlmOZ3TFrKR2+M0klP4+QBLJU1Y8YB7Pc8BBdN5PPgFio+0mkFPJoBqqSNvCWkrni3pruyeEUyu
sByBBEWw5y/BcnMFxhMIh0VcwsqDzbPmOBWGaEPggiKhdP8ocIT/brFzQrOe6k9dBY16Qn8HqTPw
h0HReybuHI45EdApadoSD4fFKG+T2IG/uaVvOVdJo9J8hGmYk9Ft2ouZng4H/a1gGrjfJ+74dYX/
D+dG8E+66rSU7VOhVjbUxnkR/phg8Ccw5UkcyjIOR9aD+7VpPGGRJFzWsvtd9cVwtfIAzPvAqpGf
2bRnrisw3nSOncnra1GNiKjBASDNWWxuRdy0UUYaPn/ZoIKE+h5oTgTchz7EgCLgKDuGg4w3fRER
cmUibf1OkQjsNR9/CZm1uFIYfJ615xU/JAmtzUtsRBxeEilgnbnXD09cexaZGElCqzIayCoo6L1r
fPp82ar0QCwnir52zfgJ7cKmTNqVb6VU51qEyG0aElgGGyPu8EI/1ufyG4ekDhBuU0f+4TzNddxN
5Jy/H9nRnkwQwwU9kf7V5jO4qSQJ3jdhG5DsYHMv6qKuUwpAQUUMrnN545snH0CniIt8HLTmPncE
plnJQlpY+5y84ZGlXwU3VW3wBgCeL71MTQ5M17Fp0aqU9sqUEgni/HFYOdjhLI4ZsZSAt+ZDk8dK
lxxwjQoDq8NNs3zKsAeOgit84dRp0hbULeabM2HcvSVAA66g7zG4jMDOj+rAl5TDyx6sMu2ve814
qfRMn6d/jeAaVTkAevPKaWUVpLVGkHJ3G/+W8yke/VDf5tC8DK6d1sWgemE3gqUancQjHqtv26/V
N/lVkV83Ad965GGRhQisj53kktV4Qk6Q2hBWBhLS4wtBIN7kf1QghEltwHUj5bMqlWSMQ1Eunxp4
K1cppXjt6LjAQmCEH1N2ZXKvm91Jr3ffTdEG29Kg8Jn6au/XHH4AVyXh4w5MJ0HzWxoTIFJAcyaV
6bU6NiPXvZtZkzAOYv7j1U8Z6FD/BdQka5mdQcDucCBmbxsa3DmZ1QwU/8DUo5VSf9IKA/qL+dWW
91ktUcep9cJSgaBouWn20uxfXjDaVF0V586D22edSNxRYBQ3pJlP3m/2xK0YcX8t0NnsLkwY6BwR
Nb1bvzB/dp1mReZxCpT4lzEv9bjHT81ZJ5w65S09PeMme3vuZ8IGzHIhIoDH4QcB/jQcfumC6g1X
64SAJyD09/i0cPlqgltcN5UFR4jyzfT5ldd7RPkOGWYJCk5eP347ua3R69Tj3vYIRhifov354Tl4
N7xO427Y/MeynJvAJNboEslCYuTRaHl2ifOQac9FGr9Jh3OC8oc/wqZuJhk8UlAtAEZerWPbTs1M
jkqy1X6pI+jbHyffh7fwtoRtd2ip+cJAiXnbsnu6t9WzOCOQ/hX9VVyG1hxlDIQvk86au134tTau
y/0zwjVEbnVCLJnFrqV6nYqU809NBmoNWEu/QrbRBBcnFXAb2uFIf0OSg22Shu8n0U9YmATlsFwM
bMHZ+KTuzW+YeBItKimJbqr3qx42MazZFbpEax+HIGv2xdYAa40N1Az6fumwjKBsIikeR3uHrvWm
sl3aI/3OdrhJ2ISuOPrq5d/uyYnu/EPw3Qcmr1nrqE9M9BzaSPsc60Yk9D20shJqiQbL67SGbKJc
EJOE70yhyOLaoRha3Vcl0+MsDFZyCXQZTpW2iUqiKx7KxPyTa5kLcp0Rv3SdYoROm1CE/OSaZLHt
VzN1by5nml73T1i0/lzkcn+GH8JNeazQOGhBb8jXcxvL1F4jgTNO6OxaU7+9ToQGC9p1zxONpHSq
0EG9xO8KXhcJrW+gSzBgcQq6snFRCHghIe8hPh7vIfWP2ec0b3+ihF7AKAmdscpYPuWP4Yp2OuPY
qYlNniHpUx0ik+1G0tblyLGTSkV+/1P+FtF4p3WHoEiNokEVm/8eOx6QuHe5Bc6W5z5IZfU08RlH
6Q2LnXJmvOAJDpn4ywrDQG5d1oyku7wmcDsoCoLS8H/fyay8YSfeGQ4i2974d241noWuXSeGBRNY
TNfOYFFg/aIlW4XLrkVvn5AjxBa4qV9aMBeqb8XlaZKvbk2PPgsrqPFGsMbBrQ/h3y6bOjcN5Brm
hFQFhSUWRpigdx26tbWolwf2bYzFRMlNAqqPRcf06svZuusIeXzlc7qcGBiA3FWAFAFPPH1IhNKQ
nZEWISug6C4oCyphx3jxrYbu6ihTfzle1do1n3C9jyG6QWxXUkOSJFNTFwOfWZKmBFP3eiH4b7FI
OYEynrcdQ3kmwPIKoitkoxxrEKTmpRQUvvWaBvgReIfJgcsZyxiwJzGHzsck/3NAjeBgRK5bfxa8
Q6kC1g85rB/tNEnVOnNGpYQi9q6FgHDzC/d4Y7yRWHpsVq2o53QHaNf/M+avEvF13LyGLHIBD9Md
flso3ysdM3PtP0OEyylvRfaxC9w1+RJPXhxKxZ3blYPVel3W8WG/lTcDndJD5gjVqOXYYLvSuQr3
IGIm3qtHndkD50cvLyCUeDh9NdCMb4GRAXlMIMwtGpuqS5LZSMX/CW2J+du7PZ9O5iZQ0JuVd/Q9
uxcI19x+fNLTuv6aqPwZmyRYQVeTob11q6NqXsfhW2JxMdE5eORiULanjf4hWUtwZMH9MO6W4Nd2
wlmBOrZciFQ6w4zfx/lYN4RNyBnLLxBVxcrQSCAJ37gKpzWXQ/JYIzUZur/p6S8+MgrJCO3NN60r
m+FUNDUOD0tS3P0nmiwIEXmESeCSXG4osz5RkQQtdz4PoSXFUd5rSfNUb4dLTJ4shBOH7C40xRdr
zP7AgfYe0+qfYWuLF57sLHAm9IzRcZkiHUy58Du/pjo0xOxlHXgbbJwKMyfdGSbCfBLPlOjGyvCM
j5B8ojuTCE/zfQNwrzKHRWllOiFMWMwVOw+4nfXSane9GIkWbDB1AV6OQ47QrQvhuOyYA4TJSdgz
+CuNDyDWaMxKXj8TvVW49ZfxpZIJ914z5mzwDMpu2OEQt0YjV7IL/rC8qpyxa7SWuuI7VUl1NXS5
fP72X8MCmS1dcY+Pi7AISGMzLoA0B10w3JAOyasJKXlyT9YF3i9YSLpWxsMalL/ywLT9ZSHKp2xK
pILAXc4sWSnT50wRU0SUqsxESaDcYrlWCtfKmfI0VtnbFBaFC2D0W5/GqB2Fwunt0eJibbJ4N7M+
wzvDIDoUIBSw1WyYUtjYkWaAqYlCA/9w2cyXCzYkoNCMpjtydgd49j50T+BRM26IsISaQFIPD9hI
IvSEtw/gGa85bxGkycsT8xcO0B/XGiUl1CwRhuVSBQEzl6IqDKE38nJYqr59UpsUQ8IEJ/K+3LPj
g5q1hdtOFpmdJ9BGzook6TI3bAoFrpkOfcId7u9vMbZ+6sNqYMcz8f86v1E0PwhSzuy1Hmgfx9eQ
UvyJFHubWwecmptw3hwZRjCEh0/OamOesArIb9wQONZY4r+sgDbs6LFb3KDtL7M5/tTZAwTxs6WY
nspDAWpH642EcY/j1E6hfLjBtrOXXtv+vKSSpkzlAqw4hLp9r3dXiNvx3+7CUDQAaonNTL5j7K4u
Vp+MS00T2Ojf8NyhNwe3nQVMVqgHeL4W5kDblxrauj7aN5CDVLcjjve1WevhE5yZzsLCHQums9+H
GouHjWjg01A65HL/5FoyG9FoQdlwVJZJCjrF2hR3Rc0qXs0tSPRh2vL9TYrxTBnhOM2eBOrjC04o
rAHJv5BPiBs3d9v6qyRz2GFYTcQXKieR8qCHbBeBndAMK1PRsMFe1UWXUKPiZGuIUVQB9+9W0y0B
8aU04EQX0RD8OUs68HnTaoVLlyws7w50JA0jEcSS8RmrF6Rxoi9MHpgsrY4O/cYn+tYzaaeVt5j5
P2E8YXYGOap7qklgEXAyXRJF7lRRWyU9cRMXbL5eNfSI91jfQ25hnaArl6mTWYAAL4KwyVWCShWK
0CnndFeNj6Kzv0ESy3NXIjKzg418Wxc/QTVaHPSzhy6Pmt62U5V9/ZB1bbYKgE2V3sY4Q1u5wFCA
1+4OfKw2bb1A/H5LQZO+xvmHNg7cmgAmeOOz+NAd/L/f4+IZHu17hab/r0ehkHxIdEqd4ABHRaHI
6Dga/YNVf8E/vLRC2IlhmwnLHhbqn9uk2WujRz1QSLYtBZlOXz8P0zcveAMZemFJ0j4HMyyKMz/8
VajQxmmUveiypbCdKhzoCjM3rWycfpPahmJ0SUL/2rNKD+u9/sW+sOfNOUWbigppNbciAp3haqGM
FsTcZhZr33YaHh0+we0KDlFg+Fketocvb0kT9BrgzW1H9ZBZNRCbYlsN6ovTWIUOC6LO31k6Gss0
Lxm9L7jOuUF46u5ljpcPxjVfLAIiAlDpZfiKuj6cPOj/GI14NFVbbvWyLQuuanCLQTebDRV9sl6C
nLvt8Wrl8uhzGvoV1dVaYSVch2KhN7xL9GRszBgl1uXAv4EqbN+2/HR/duLvuXh7etg8WSCwBKLr
jYwoE9IKWYceODjKFrrZs9WP5Jry/fgAK263PdeNaHdkjP+s6kCMescoZ6dh3YpO08t+aHeJyX45
TO5cazOBMFWh5sMZos5+XOzAP8OXbLfHZwbujMjMlRan2aGutS7QTy8QtXfq8J1QxfiIQNPmWB3q
urs6779uBRJVTaaGWUOOCJUTXGMos28SP+JqxQ6o7gs1lpD3gk2hVzb5+g9V1/Y1fJ2OkUxwoEa9
JJh2arcTFIV1SwZ0FXWQHChlF6co070m6KdsahiPiAEviuusiXUEANcoOLJe+AXkLPng22ejG6Sb
Gdw+CoK8Hwnmgrf9tGNsw2ZcJK6yW2p4D71BnQO/DMsl4gKBKRvVTG9Eix/Gnp9Hj2Ib7CNKhJ3i
wESCTwE8oXzSo35BuyxnQgEP37NDt1/V1P7iTtg4+kKikv6XePFH+RcfIzU8y73HzFPfXPGx45Rt
UVG6zsIsL8E5yKEVn/znf2KM1qPXnP5UHPtkptPmttW4T/37b/IkQDKNcM3mDxXPSy2oSiNeS8BY
IluyL0JAxkfCWbC+SDMXqNWlHYuSQGB1LDDb1XgxYZddvh6ogzdtrP3CFEB/iPYhmNlGZXOjqCf1
0hiQtY8mXXTVgh79E8Ft2pT2bTV0I+8/LP20r870Qq5pqIRMrrHeCXMmvisfXEd2usGkuuWMdryd
8OtFvJy5EIP34gbkTwxB+GiKiPdERx9El2xVhzyM408qwc3TxnprZkhxncHZrZmGGvPMGXFgJ5Ks
HWNDE8OdfyNu5487ToHRwvT1TshgaN4SPxy5tYvQI5SORRORUFHAmxjAjAkaUKyjmId64f2Ppqxl
rqvlO5HznudKdd56PB+STrCKukY0+bp3/ag7Is3p2cAWIiAW4G6F/n0heq+R+rzXNybCNSbVONzj
9K05G/H7nUO3iqsUkJMFOeOOxGn7skskBKIhnyILM5N5eaCoC+44LYHntgP9U3Sv7BvUVM0Eanhf
T7HzjZS+01Xox6GMWi83spdLzy4agZShp8yVqq02GbiiR+Jl9VJcZYhLkKbmaj5AErddMUNsuRIf
7Jf67bokARm7eywbJOy3LkjAFsLmPbGeUIAy4ZVzR48lN1j+wzacIfcHqapjC8m05u0+YDGazeWi
9+8slcibioarXp4VVjyFpLlN3Wud9uLKCaiXWBw6oY+lo7pSsicPlhdWwrXjBahIGluRvMKeN+oC
5hlOr8+fAnic+Ydp3kVyHioUwE4R31jSUbNtLQrS9tXdu9782Nu6ZSt6piXY7PO5xbzYOU6s7G73
IdRyFI0xyKfzj++X7eDx1F5mCVGVi747M+GmEIIowbmM4ymWS1XUtzX993AqjcNjLgjVer2M8oWm
65kVNXA3Z+6HocPpuEht7bhgTJo/rPCpwoMRdS0Q+3FH+Sm8P16ddVH7M74g6UrNNumEc26wZ8qR
Cp+1ApgDkg/BbPcOX+cq/f3B3qvINU0v5efDV6zKigv2JFfG1QhoCulvsaGN99n1RbrCA972s+u0
GGQK7sG5HiChnTQbtjDNqJJg9muTozHSTYLzzla6qGLIe5bMprKxyaXi/8QDK0SaBx1lYhVrHpl0
KUdsO4wpfklYeLbgH02Lqs/SNs88Mxnc9n+464wvYyduwb6MQhmuVTC7aXRzB9nQeNPjs5EHheN4
AwIflbGwltgm6GLHbMWPEbFtg1/OueYl7nsxtFO3jeWz57sGNOA7r/SGrB1dVLqROi6E483zZ3Gi
ANruBFfE2KmlXRCmVG6SVSHQ6d1wqR6ZKsO00LRMwwmw+oE6NX4i7AURphdRWu92pI1YH/V1rZAb
J0wlmxgEgW+DM1xvK8lmy1bQiqtDJVHezI6VrtTtmtL3Tu6AO8URg+xXX3N8NrI03T8LSG2/rFGv
/3IpnwnHPa9XOH1nWHjtCuITyNZnv+r4UgQ/Y6kahMR6xlEZb7gMvCd+QJVkB+w1x9bOYYjH/8cK
jUZfSNDEyyeYMu0Dz37GH87t1xqxl1kG6qOvnyxJhESIX9s0Y53bSZgoCJuvgTJgnA9kPsFy+Gtc
dfc75OcGuv8gKtn20gxpoRkX8mVk8xjVOfcr2uuizQsVSB2dsvg+X1DVQ9602r8KbbJPT6tPImZK
6N+TQJOa0Am5ePAPqcGmT3jKAhkQNL0rBnOaMgZphcOTf14XlLSZKwBzB9Rw903a1C7krhXvnPFb
0wRWJ7UiCsGd+8zp8V+Gbl4oqMRGL5Uke4Pz2cw6THsrz71/cATUGw8Gn+81V2ux+IPmOla12NO/
KVWc2s8/spfSK1zSKmSSAhqHPVcZacLr1NRNBW7jC2QNI5hgXETRsQQZ641S0FyrMue0vTBexo81
ZNBf9m7oajYiEIvdI09M06snaN38YjDOFqmQy3E+R6hHoQBr014Quy5AzVAbP1m8FS8R8+OBhdFm
lJN/yGL4i9oul6fQfF9Q+W3UbrjJhuAqYDSauTF6/OMSUYFC7C1Yzu4X1dOOSfHih0pRHCbjQCWc
PvcjnDOCkpJ/dLX0l36chFbmqfBV2bHw0eoEWVgmPQZxPepazHDDHLJUBxqKGziuu9/3Il2ljHNi
f5yd6eFSZQzjFxYp26z8mPQsC/xGugN9k0xd+MYIOCgdzqc74ADfJB+8YTjT8I3sRk32OVHEXB8i
YCk5nlDCaGMtnDnSbD++pCynU9uTzjDNLGdeU/QcLXZPQR8Vgpf/X+NMNzFiOl6K7Io6LhVBlulP
52pnCazZh/xPUwkTvSRuBRtbDZjjO190WDtL7l4BTvomAvTCKPIqFO+nqYM1i7wIKS98fYQcW7o6
ygexgkKWsJl465z64KmvYrL4UwA3hgnpopLYjmKYcUetKJGBkVtuh1rcdov7uSxfRh5n4u5Pfhjl
zcKokWdrXv2rKdsnse0ZmD9pJI86g4ydlk7r4N6wqqC3BAZ2+N9HbSsYFL4UXJzESMkV+CouFvY5
DmkVzzahH7UVthX+rdruLcMHZCIUyHqeJQ8d/kTLVKiPfvxZ1tZLrDFxPdKE4RbwPO4ZESiQLnpC
+FEKXAji5g4+qjDXBGAnvfdWf48hzWLG5RYDkv8HIL9MZT1fUEk4Bs/u1VJG2g/wNpeUQTfcETD2
Bivu6qL4HO6kYkFO6LHu0rzb/B62L0nBBtH3TQkfGE84wyqGpiOd5Eg0ssbdXtORbk1lJXuEMeeG
Rsc1Gi1J0dhLseY68efU1VIj4mipPeclLAf0ZYgjhG2GykgbDvxUKO2mxiRnHyce4B1zgapytr+a
jqIWnNmxlZ81u1Mj8GD9XPsDXk1urciP6htApiYVoFxDFGKIw4mYhWI0qgFFyH49WM+TExEoZyuI
yfNd7w4C363M1u3ORq9gIYGxxeiI7vKW0FpNYNDiLhHXbs47GrmBwf9gx/6RaxldpPYmSg+duYVo
ZRg5KlC1Lia37F8XmYl8pg4i8isY2EnDb4S+O4FRXuzfDHskrA3B8ijsCA49XMPP/JkZwW2wXvZ4
6spC80HBSr64YSb/3woMPN5XXaTKRM91LYh7ClOSxA542ZWVk2NXSfadWponnOlbjYXxU5Ckqukc
T6lNnZaimVqHAHy1wNNrQlwlIDKueQgNtOvunT1mCUwnGi5nTKleonrKMvna5OKZQgtqgIGAVAi7
U0I0sJd+9v+FJBmVipLavJwS0eB6KdgfDyiPTdjaehaSmg3ntNSAwBRSiweya3LFIBHODHtGG+Nv
YzcE5oqoVbDU1lgpRXNp2UM2QFinAYk6kROkH+utL+9JiPNr9S3ea3SED5NIhmOUToKi7/alJ+iM
yEgdRzdEoFXnWsaedt6zjF7IagWPdU3ljlHNAyaT7neMjg2CzTA0EL7KoEo27hblrbAAU6BLHDlR
X0iF8RmraRkl1x+ySMx0F+V03BTfvl2Kqbakk99yAHfrfRLlOcMCPdHs6MC3B8Wg/MpncH/bG2ve
sHabdz4uxSVb+jxRG3PReBXzQlhthOWk+27RKxgHIIvhE7Nv2wQknPRlAvd35mmBYyOcYd0IpABO
xyX66NdK3XNWiqzdeeoRpZ9dCfVmV1e6BUmCCZHxFvR090P2R/WpWpankCprFG3aHM86ocn25Xse
NnNyireWpliQOJKi3oufTbXRpDGvZM//jozXlKkG+hZJD3makjKjBlCeCFN1tAC0vxxHxMMcfN4t
RYsP9tiNsdq6X/Itm2dQMSKFAlAnVB2WQekP5D0Eg1wAlnQulP0LEpvxaidwCAlUOZcfJexMBeWd
AbFNeIk2qwzBx1KBV+kFfMFd4VUkOU1ioWwH1xPs70NiP5VsRY6qGDnz0Br6mWI92B4MmMSfE8Rx
V+dW4roRWvRM4ZnEWWxZvfwBDvWyAhtES1nFrBeqBcQBBz7/50sZaKpgVHEWC306VG+WCTRcsvVp
u6FiIygkFUpJMsVGHcp78DmN4HAmHQ6s4Ucjur1kPbi/vNzwbtYtQhof7noPTNaUhF9w8tPHdFlz
PVblKUt/VJ4UD6nWEB7IFeRGkeDoR5vC6qjbz6SP9Lsuuph43hyby94ea2QWLuFDjn2mhHbpmpNs
de/441dT6MPOhOKGgN4m3zpC3I5107J0q3+cdykcOxs8DVZlp/EhcdvOzPipgR3oA7DUhJuNJ0qi
0zijK9jFKaCMyUV73ASw53FQkYoRFzYvyVzlWhxQHxkMqzFmleHGjZp0OHrNTcoB0IK1NdxCx5o8
DBwAI5U0u+H3Pt4DJig0eBmIXsOpabkGMdVLAKi6JS8/wp3AAjvyYp93SegetYtpgsuuBi44QPho
DiraSDH4K0toIl465zaP64Kp9zz/3pW+tLM0LmLnTYMgrsqON3vz+Zumw/GUpdR8Hn6TRAt34s7k
aor3jhmFUWaXcvqoUB7zQheLjed9gXFnaK5wng5kPBVgnGjrPRgXh7TApIfmlOCHbxLafzEf0YEG
IqhWODJxF1Pc95+hj8rmaLXos1ch+0KH4DnKZuT4a9kx/lFY2D24PGtDLiVPt0EzfVd4aC/zm4C8
HYvxJkaGHB9rjQv0HeUs1n2GOjkzso77NgsWQhEwFvICyOXsMH8+i2aCsCmEsrNSd+XGY6HYqNtP
sVzWX08aZ9zYmtPpor7VEHfetCRPTszVU2IqS8547aeLwt5P+7GY9XakV7dK1bqQAWVqaSCLJCLd
S2Lu5iDVKBgkinJx9yAH59sv4LU+P7Jc5THejxrjnnjPEHKuFNIcmA1kZzGOYNanYe9uPOjJ+RwT
kmvCt2S2tTu8qdEJZQcqMYzIKmUAzyRvJz/GUY0mB3oz3wKii/BZpZbgPUcTGsHhs0/Zv2mzVsEQ
ppv9wltCqscmADci0B6FIzdybGeoS4jDaDyx14AyYemNCnZONxkokZfCEFElkRc0TD4/4OaBaha+
T6iq2gjXS11iOE03EXmh7/r92vHK9jsi7RTdrr/28wui4NGWBQ8U/mdJCze4TbwKdqT0S7G54/ea
Kj0qQPEW5s4dJB+AZc/xZIDXQSX3mDVxMXH+I8Rvl2ZPiIQ6Seb9CLzrUaZ+O/lb9VWMoCBr9nDi
a/HyWPuqkaDE6O+OtLmRkdhTmS6iDD2aUvxji2oKbA3sdOUNEKZz0iUn97n+JYvlk02bcMCWu6Eb
KKItwo7wx0vAYYzzU0Gl53aHztOVCeTQ3tRhr0lN26X39skZ3cLzcGFhQrRIDUkCJuPzo1osYMK6
698Rz7QeXh9Jlu6eigd/v7+ghqS5MGvz2Tap1CKVPlK02cNwSL+jpkhbvzNvm9OnbWCqlbbPIibp
AAtcVmLc0aCOIKvwHrXAdIcVXYxXEWNV+sOaKCWBCDORytkPjzlVTNz+ZXyZ9QwJh0UEDvvWC9eJ
xsNOxd1YlZiMtoNRoj9yxzvnHi5F2zUyn1UrjwyrgNu2eBVExCwG+9PFw5nKv3WWDFxQBJ9bWDWK
JKJCOADRuYrw97qNmIylEFH+eiUe+ynsx68A1j2PhyprYmXFoHASvjxCXoUxjkjigaA23KbW0KJa
+2BIyBxSUR3yK93ElOnMzqAHuWxfzfW1/AnMo37MaSNviYdldOHOi9Wzp7vTsbUJSWxkYmFo/p7e
7B1kGSkwcr+7+G9h78bC/+Fhnr8MM6DqECKuJPqCGWskYHlE8/5MVp7Ajpeug25ZthrhSBBik3NG
UBPVMSZVK/ir0pUKiTKgaUKyWdPniclYTeNnc57VHf/qrg9I7CPKPmnrW2qUOoF3XZEFfGTKB64I
ezCr8cu0cXTk9VJOX/Z0n48tN0QA0xjTOClPxBHSPY1gXohFXdiKaI+zvsEJj3oyWsaeb/CaRkCC
nspqYAEGqnycEopqyx6iNEf878GlFjUDlHUDpG5hcIMHW821mFoBo8Zd0uBZtnowexviI+J5HMCl
cd6bXxAG03P22BEk07KnAn6IHKMUYrcnfD6InZMgXhFLE31ndpvSRBIBgQlitsglB7An3jNz2xx7
NKm08U3l5HMftn8NRRpoF1Frgy5jLeBz9dlgvnjlJ87fkIri/HhVOxx0JNwBa6FnJfL5plny1q8r
wRExPxHagH9n5wdDoxjLurm36zlGTTB3GNREsccV9Iy42HirUB6nDTGIsia9VqBs0MvRfgyYFJ7Z
C0eJiiszzKRN9hjrvsI9hdPde9Lk3xLUbvkHAoIOKCLGBGFtyAzDu4J9uce0QQJ6L7qpgnWnOvqO
GPonIDffultWCgzu2Ds7PMp8bc822PcbF3knyzieMMrJFtgZPAWyZnpehc2wfrIjsN9m0LWMw03a
8NVYrTeQf5kUlYQpj7/ri4JZdQMAHaqvFOy0DYmuba3DTTypoR6qOHwLjh7EYO5QSjAGcemJFtMl
BNDemRKuek6ct2tT6NsPmh+ym+cKzEUd01Gg87kUFkDjlO33rNtpFlYPiTJJGc7L0YyuoK7GQ0mz
ocMQ8NVetQVx226lT/BYCTEFQqCghlIG2fum+Y38qi/LbY3WC3CoBoHpfKGXtg3s2Fr0ldvq0g7O
38ERtLyV9FGlVg2HguAos9AMmn+jLpCanBRG4pjdSiLuFMVuA0VqebRABtirt71+tSPCMuxoQKtt
wAc0BhBOLmauM0n6FiLpYH4Fka4PoZ6DelHmAhSSR25N7kKwre2q/LCssLWMOtyal1laf+/XVQug
+etwQLLKcdYHm2uDktAm16FEwWoUSx4nBOzMGEbhHb2fcqhMqfWU9bPZDx3KApnEBxBH+zBO2KI0
OLRwF9ZImrkUVT5/P/KYOxysz0wUQtYFaM4kiP7z0zFPoIHMGjE337nkJueFQlbk+Sey7ze2CZOi
Q8XkL+jqcsit6AOGcrvibmAJ3Y+EoJoTo3LliO+srGrTMZNozPIr8Gm2TV2pB3DE56X0Gk9q+9Q+
V1TC2wvR/O8VG4SKrx6pX/IYtpDE35LIynIkBgwC8O0vrWdR6BQqsHGSnUVWRGTNWZ3xqbBAT1ae
28N/gEVroRspHG9ZDgwsvEEKRA4yrfMhCZjQSwpvkauaSRnW2vAMrbA4scQmbBriFvoKvSjIZACf
pzAh7JbRW0e+RzxkUZlLTFWU+v670Cpz3Qqslc3MxTAxzNDaql7f8efcQCFRWVxSLtp+0q/QH3sq
p8YpUIxerRt15bvsrx377uFITCmgQ3QIvwp/4CSOp3+nunT/21xzIiEcGtPWpcWQAnRKlNvjRKkc
9s4pkcVICFDaGK7oUMfIe5kGxeRq7XqomLomfWFIg/njFBxz+xMLs7unz/umtsenk76qud40xwhB
xkQ8uVJRH24Ks/9LqzjSEEEDNx5J2S6EYDvztiror6bDcNEufKOovQkAh8o6aq5oWvXP/6vNrFDr
QwQErYpaNhzpraabMK9m1ml85knyOt2/LgFlFjQbwHkZ79QfdV/D4HGZs9mj62sciQ8+a9yUadsw
IaFgYK4gRqLiGcOBiyFx2vGq0gcRmT9wYMNtFrmvVRUtTCGZ/eBS0th3J1mPuenukSfDRt+GB5mH
exdj6eNwire1+EHAmhMyU+6EKbFkkL7v15qVwd1OXw4C80UyybvCFEezdXmBr3ZwEs904aBlaY5s
sT1GsPFuABhDK4aK4jQjZybjOkKvZG7UdQT4vUIZRpYF9Bo4L2RicywJLOEfkCDBH2GAOUVvyG9j
273GGFMaRVeH+8iEDYIC6hd0n8Kywy03qYcIlxOlo13EQjwJMauMYSobKbAaMWPDhme4iehWb9o6
XYWkCE5rEyDqEUrzGH9amkY3LnZ6IRiyFyqfviYnvyrK5guP/cTxwa9Fy0UEP911slTlRS9MJEoc
D0e1yJA4G7qsDsHJFgxWAtyL0dMplpN8stzYH6snxkKAiqCWtpvdqHbQXla7qbfOCsDck7LVLjUm
715H4fMnDpOV2wzkKLOp3pbAdLBz1BZtfM+MgFFEmZN8kh3ekE58dr7wBfP/cPDq1c8fSVFw8VZN
jWlt+7MTEp70kNF0pzUcM6ssCCJztcMht7Z4IBRYNAb1mDNb6k4TPhgFqFR4usU6i2O+XaR5Ai8X
I+9AU/9gptPOLJCN8NYkK1hStxPfkYb18VXKTNQbsQ0/fOUmCOo0/EY3LNwvltSfLez4YWDIT2vx
xYwFj0KB6I72w2OZHJvm187OW3WJOYhOrlQ7t5r8luPtFH8VJuSG9vKyUpXp8qwvpt0Z/U5fy4Lt
Axzrx0RP1iy9sBNn8EmQ8FCvzivcgB0pUsh313Aa77UrwHSEj+rEu4+jb3hqWuAnWcfij7f8pRma
Llvtj884M65uJaAk7aWuhA7GWuuPM5fPITOH0JDvZF7heRxYowPDnaI1xjWJ+6TFGXC0Xx24dYyD
lvov4FPHp6vhDUNj/d1p5eXUBKWDyjBHa7sogqZ1fd9G3E2cdrK43/MKE5wBcspxouMCKecUxOS6
wMzOU1rNMJE0/qbfqbXZscQyTOQ8Rlo0ftNWWc1MxhqAVNfbIZtzbjGqVidzB5P0PAk9mgMQttiN
IMfMawvNJzkl5XyqatChNX/Vd7L5CdPx+/bmBfqDTwv+xEizkcFU2fsvuadn+sFHc011HD9eTnsI
NYSxnpMQEluBiDwDjXrfGDaGItzOK/OCevA2dZfZPyIogsGgRiuF7Z+Q/HxZ1zffLHAOBEZbigbV
hsZHuKCmZii5nz8rbdiMvF+xbBwAAKAubJY8w60f9kIePercX6RfQSYw2TVi4Gwk6nX//NXrv1VQ
FxFytEd9azVFzCrKpEV2+BjMWlAn6rEAMHp86Cx52nJBYbaLdzdvjsDmiIaD+x96l2XnY6dk784t
4NOnA+Aeh4Y0w1zC4FsD3chT6mRpu+aci7cXH0Cv6q6ts/bAHKM5/0nPodt7cDY2lwojnVNVm+Q0
JnQib9gQT0KKB5D3ihRlFPJgkPUlEa2c90LtHrH55kb/AkOWVdncV5DPeDw0+IDGgNHz55sURvVA
Xip09nBo/Np7KQp929svkLg4Y6kilGZippG6S4FdTzgbcy31BAY0vuJtKCJdl6t5/hizXYtuAp24
TpAg14ocx6KTGugEvkXdIP8NpP4A3rAARAXOYwxhranS4gZ6q8779Ll6lj7ygaFT5s4M/cWOsdrQ
aP/pqkbsMycz1R5hUPmGjUJoxMI8LkmsdxUmKbXzc5OruNnoeqW0LnvA9TeHEwr9uXBk7KMtc2XA
VlW4iWCTJBrx2S2PkFrmG9Ffy8z463hFFy3sJ8+3+IbymR5+l5Xz+aqGxI6Ze10Q5/YxVoWDXjv1
ww2f2SXxFLormd/rKi09rs8FFQg1C5uDNfnB6BfW037/c2qsbJLMX0QM4xOp8PGDgMk/+D//4bc2
LLzMgoUFFvspEeAzeLmX+jJIWNB04SqhifKunx0W7qcHriLoxGZdd+k4AjSGrrYP6+0ZsRou/kf/
lNDqZbcWH5USqItpTe2cA0JD+vWXFxRO4fU/Nze3L9MSYA0jYPr1rs/xVCYe7H4t2Cmmzd6lMe6j
urUn6MsJVOwzYw/CLTCBvrjBXTEroiM/N8s/al/XkjF0sjt3Dzqfei4rAxE9FN3EAz8u8brIkeyr
gRj/zNuT+WLPoC9YlraWH+aL6R2PoFkhEJd4dL8DlHX9BvqCW8G9B0FuimQDC6K4sqSNVVkyA92k
OpTS0HAh0mSJ1eqzI0/ZuJ/CKztRdBYCQxq4zCCrJBgxhUgZugO5o8BtbZoUi/G45bpjJ12M12Wj
1rlr1LlohR7X+jaFttfiBhvA6Y7aAjXHsOgHfYqxtNrlYDrIzlEdmbokvcw2QUiIvb1uT1zIncNo
WQ7xnOVshY/wt8gUVqFqtvtQcVIkNUqk4WjkXacWncJ30+eKwQ3ktbjq+L0CJBo5hhklaqQLHaTl
N1w4rk8KP4bxd61+5HW2QcR+4zNK6+oPtesE8rIpbJWYcNtNRs2FyXO2rMceSIO7cUe/jlzPks+0
KnPOVDiCLwFsh398+TtZscdrUks/rS0YRyfwh1lnyDj/OoP2uhiGlKq7/yintqFRZecZQFZusYA8
oxc+2VWTa9/HqvyxCOWQIQ+pRbUpOLcBx25NQpruCcmxnOuCe3YoTjbrQpsQh9DTi8gJDzdF4179
rUpUSabYM7W6QZxNFRrqgSYXUTrg+cmMW3xvoinXMe4NwYhP7jYbwELeOIVQm42dv8wxXiT6eglL
zC1e/dmJ9YOhQxOFJg7JKMnxUaO9NE8EloXT/3ok+lrlcmw4RB4mTknPA0XZzV0u2ZJxNY1az5/2
oUwtjvcWRg3p0OjdYyN8IJiAvotPuH7vtB3YS1S33mcYKpAsEw0E31Dvqxt+/dwOVSJ+sdUrOT/X
x7JzDtN6CjpBDdc4HCc1mP5NTWrfiNYaaETbvmlmKMuqQ+E250w+k7fZsQo7LqGDoT2t69Uu1O1E
5bC4PFXLmgGYntiVYVcHAiKpgT8YLDf6/hCVfc8hXyV9U09Bc2R8hXoGjGIfABTISTDHvs5N2ihV
F18gtC7aPLI2nq521seCxppgr0NueSsZNLPhnrAjAJDboM6pjhSsMgdiuRTobstURy/N46jBaIBf
4CN/zDNjGpyVXyxVV+LWJWxiWqoRCQB3Uf4B5WYOl56l5rWcpEupsXXbxd31xLnZhBihY/yi6pP4
2k0gvRxNnFEL+clOvVKGzlUPZ7tHvuM/Wurj+zbvTUPcvcjNlKR5nGHE8RU4NFZJfZlPICorQ8o1
41/aSud0g2ZuTN+C8iEoPzxrSl/FPm1kGwzf/OxT+IE+W/Y7Npd3rVgGSHXqF2GfX+xDg/kLcazj
ua9Fsfn68+y/qTPEYYxlNEanfQYhAuiZ/ip3VNinUst2BCMdAKanaCkl+Qg6OsbbiXmPHTBUPmw3
zkkXRrJ+hnc8T5eQwSbPmkWP+s8fgz7vOXjH6+YizU5xzcGY3x/cffkfPkaQcuts9yu2Q/yLNPYt
Fin5BJjusgFOWfK9dPY4JC+zG5TZhK/mezAdE0IIG3XnyU1RTph3Gqzmz8+u72TerYALhOpm1m/V
Bp8hdWoBng0e4VmsavplvQVlUDQ+WZ3v99onDj1QHa7DSkxXPwlLGw+HHQUzHfLpn6mluv2XmnjX
ntT1/OdNgO0L1f1ntNcTrWcvrVMNVUoqVEFl2YMRf0o9VqA3uYxaQEhRZwldSbvkqNc5DZUxQ96e
zmTwjqvF2Qq+o4Qlebu1O4VWvoSLrgIZiLlGXABiP7qMCp6rQyf0IzcIz7no3URqdPVo/SYtq7wh
KSUw9E+mkRgQygxSk9xu5KQ0lk41xs0qCdsAXcICYem416GrsBM8X59dYO7TDIesLaxlaljm1jVV
oZ7XH5UQW9q3GgCdfJsD4lXRi5rGULCohQoR3fZq6stnMJ9DTOFCIsUEUo2bfVC6Ax45T6JTia4g
OuPOcpABQwLhePeP2efWazAm4ayeEVeEID/kBhGVpkjCdscGuCY43dsHLZy1CkYUV4wFGiX52Ufd
EXaT8h0OJHooxEMZK2Onul37/diOZSwkblNKlryb69X6XkyjnmvIC7ClfsBN33g2/jHgWP9N4UaK
wX4VAHPdrf40MCDupzRiJpc61p3+8Oasb6cMA86KllO4Xr7uTAYv5JcXsrY2TF8spKieMbz4nL0+
z1p1wUI3CWuu5TD8BGFc6ed6rmU9kFV1HZpAdLfnO/s1TgUQd3aEVTuEK7OvPnCgImx4OyhmlNxC
fIlvUauqO45U1w5w11JinL9uLHQRrf3XUlcBcP5+N6sngU3nxfnc56X685uYMnPO1I1LR0A6WGbH
FTdsNqTPwawpT7CaiLvDQDyOXFPVhUmg/0+EEk95bdO6AdlBD/nT9SAfw6Cebj13Ac2G0pH6ZtLy
3nxoul6/tHD3MQyz0vQNAfPlHrGxhLc7NvcOXhcdPZuIHKeau4W8vm2FbBQ5EikVHjOiE5hoyO5H
OlE0i8+UnPOVBDaJUncymXmkj9FTGdgOPN+T/eGL9zDPox8+6K/CNJuh48GIF6XlczPOoaKxAgK8
iZHOfFLuqrOlLG1AimYobfWspXVMYATFDn4YhoX9I3fXT+flkpxEgS4emRTSP9qcicomZXq6S6DF
BwTl+JNrSkYvnEz6fTpwptk6/x/tSDDI5O1cxges9qsS2apxjfpQXxag/38ozhk+D4cR3IEMt/Uu
/qAkBXx8LAeCgc1Ii/jek1IzLmyylF7cYBpcF7Lf3tOs4zmnULGiA1CBEyGpCLoPZYMfjuhSroGu
PQBuGcXKxPT/GB9c3zRIbMmL3QpmnULpp8peNK36f72gks1e2ZnY7foHrfeGCzIwxbexm+zb4DEl
wL5wVawfJ5iRGz6u0tZWhgouFKQa0yE9CoOMCh9KKdm6XQWG9UMEYX/r/DACg8moPAfxH0hWROU9
gKZQUxzYRXzzA3iuBpVM/j02EJEfIcyGWt7FL7tdqmGRiNsUNYa6XSFQZOEQ6Cr/v8WUGPqSi9/8
e+NPQm74S4Ml17VzD2ma3srodrVO70/dA+Qmh2SL2oYwgh0jcdjLYckLKvbQjueTSxEY3Fk4m8TW
xYWN3IHXaq4AR8n13yPKkBV4lLY2701mOxROMDTLNIZ0BHRIJxXGPcLEAHyrOhrgeVI/0JZ7/L2X
YdwucE4l6ZdtzmEnYWhluqkKHqADGBcwyqKaoIbZar4XwJUttG/oultInqlnUpxenapH11M02vlf
AapWiUGCAmSEjtKkfr6sdola0v8ZCGZlE5iDAAP1Pa/eU89Ll31gZAnFWpkU5c6b1wRaAy1NDMZ5
PReW+V13yJpN05RQdVjX5AA3VNo3mLpsbvL5Y1q2KoCGRTL+0h6WCJ3hYnRmSxhLVkdWN79tElvJ
Rzf4VheRyCufnWLYKWh4ofIl+QLS6oQRTHsDyWaY20eNqPTylcaeQHZ0nKsuCwZzAwCJoDNvXXSc
wnmtcNKtA7iur5We2VYJkB6DsZSEkHJO3uXqvt7aP/zcAeMDQ3Ji00e2PnCTIPcXJnftmywLuQTQ
BnJQv5NSUTYClM1CZo6Nl1aUcLYFJG+sZsVDpLVw2AXKR695rd/0CDDD6zEulsJT8ojWUE0au3Eb
U9mQp9TlSd1EhY/gmVYnNWFX+q5r/p6GfUBok4BLitFDyC1VZ1MylJpHwqKR8EvQiHG1PmTD9Skc
vMCgdlIgPAJSawOiBxuFdz9RqXYnpkK5BYwDfsPrAoLHULtP73R8uJtEU/dRRKQQga/5YE37GnXm
wE6fD0EA0J5OKc6iUQ8+XLQw2f/s4LDjCpsCnk6mWo1z+O0g9rnqzrXBtbbaeK66DQeNxyE9XCSR
dbvV8aq75RH2xOkVujgZQuWl4bALJ09vIGcrPkJxjB32toSJwwJ7KXo3Qgjv23dQJIFDOS1pLrbK
dEhN2xYFbXXELX2gcJrvJwMcWUbz7tsJxM3Sb+VWpC94taB38gwFUHBfS7qjkY4iZmQPZykUvE0k
JbsZm5zuqAYbuX+dX3YEW9Mlj3WMr8KYHOYgI1wCh6vlxNxq+DmVdj5lCmxzrv5Hyggovuedwlmz
hg0SYy9pda95Sp+u5e0x9spW3NIe+/XoMa9kBDcBmJIbR/IiR+PdyxgVEMPQlyJ6SKOlvb9s5Grj
Gs6P/+DYSEPq3owqETOL67yNol360ANAmEFRQUzWAMWuz1WO/ZhbilJ7lnGMl5OJxnRWTkSmMTgY
J/fXgpjgyD1abW7ykLaLShSH2TodhA2O4pGBh4AFRRzFez7VhpK3+7LtdJDsLxgj5fxPBNT+PjfO
1IyYOa1omRKkue5T5D5vW4rkc3u8vu4TeMt7Ogezo+JudZsxXNA6fEYbP6jz3dwWrNDtwQDs/DOc
ceSGdlTEi1XB/GEUhpR610LHHhUiTLODqcdY/q0e52HsXdcaPzAGBUgYKlFyUK9goyWE0A/OBpvI
rVoORctqIcS3fDm8C4XTu1v5DhRH+9ls64dCSRh/zSo3fgv4ObUikpXPzQw2cpRFYmEWH65UJ2Vr
Ttqmadw3eMwPMlZzcGexBEkphgVUp9nSzyrWt9JuX2nADL5tQNVrpfIGVRsMPN99hkBtSM7lggpl
U+VUwNNH1WpP3WEgt7I+xCQdDHZSLtYDIUkXHrKhzMaNfyUzroqzg/wc8hbh21du+noIsvRrcVjb
30mkyUODgxA/cbIQMHsB78G4iomQ5FNOiDXhZ/Nr3aVhR5bQAJBgN5zNsTmgkMWUTmFZbtLXMJfm
s5twECVuUO6X8eMmVzq5zsCjN2fT+ofVS7EBzJO5rw+JBHD5cOLCu8LA1T65zSAYhS/NPE+faIj4
x1IG5Ho3S25r7kjG74kYXt7lXGSYFzBxOs4inxgWJ8qPseQcHf+Alwi2YC1s4RwfietuD91bZQg4
GoDhvu8DOKxOfYnxBbDdP5GT/HLUAkOo7DFnLX7uxfnXwr4Vmcg+mk+v+Ol6wwNnkIbLCfr4jTPs
jByzUuZxavA91DG0ZxEQiS3UaZV75II1bzvHPVoOD2Ol9bXi0Z/4dJ01h9bpn3mV1qY63NwuVDCB
tvDyPXC4PrKSYqP+o9aLMRoX3trKLPzr5WAMxKoLul50GeLyn5cNNFp2y/8hMd3ebzbbQUEhaU2Q
qI9fS47zxaz5IEQ/DX6cPCxI2V+WWAj+tbQaPOcjYzfwcna43nSAoMrZwlG/RFl2hgv9zYWXPSCb
pwSA/cEPHD/HYBr9osiX0IGfD7af75WuI2PbfjhXuEXFwNHSVvkz/8R8dRNgd3zDoehYrdJ4qujI
1Rb+yUIARQRvwK8PWKx4KMsJ67hLwHYMwVWgJ6h2DTOsixHoW5MOUQu8Y8sNxSArwfJYSFkTCO2s
0eUk4nscUtSeVdOWL0lJBu/2d3yVuyuKbVYMn+FtdvrJyswGI0OUpO4yTwzaVRNLcUSvLBqurynX
ZgaeKQfM36AA/mWpoTS1pPopKKDpcFFWkce+ykLzxSimRDCuowba1Ntu9cDjnI6kzZWq3ErO02Cx
pS23jiDMgLcld18PQQrn/gi1w1GLm8sl3Kvyztz96l4yb9e2JVkRUEQBIJwuRoHFD+UOA67AZbiD
htG3xgr45k9V4rc98J18ocsAgcfWiXmbDaK3apAN5RiFAq/jecsHMz4chy1/93R1qJxngKVpt8A2
D5CyKov3i5TKoqQyamQOPLIGqM0oIYIznPyYT6Z4l3HnECOX386+orylz/NcV//70qLheXJ8V0Rb
3qIPv7+TEJgHlfL4R13WmpKiMVq1W39bGUnADHazF2IbX/hVIl/8lmclVR7D+f6M9uFY81r9nRgz
iqUYvYhju5CLdam3gGIbvyZ30CQbYSwfhT86n5VlL7UBTh6/yxCesAfaZjh/IMQ+fwIb2aln31uk
hCP1gPeDN4O0/CyzXxfLnz+NcAJdtnJzwO5eqYkd5fUhFuSUxB0BmlMynI1iszC2z0JB+YbbphHC
fuL0wbzQDvpYXcc24QmYvA+X7g3tlKfYFDqRPg6KVYsFohLFjGeWMaXqH3oTWfX9qdXxvDGfSbTp
mJRXKtJ02UQoCQltamESKRtJ9RIpmzs7TLPAYkxBgLG+FssFNpCPlsY25e3HvULlCaGMW2jbCbUy
CVaNyDkXRBU8m40JvPHIgFLRyfKE04nq8CfMH+QvDx4iumoh8sb0c3LlpaUHVb3bWI5RE/yz3NNV
fViVR/G5k7ik11NMJc4q4X6lUSuBJDrNmB3BEOcGXz4qM+ah2URgKvldIJ3JrNSUZSFehNvwzo7V
InC0bofh5MJ3l5V9LxaTOUyonylGUpy21wHn1wvAjTY2/y/RVOe/+DEb9vAX1XsjhLm7f68w+rmn
ZwjdoMn1f9w8pZWSnhZlyLjUN0W3pO3QEJMepk6QD6NClQGIXr+yONOC38+SbxZVAKCKTKJ5teV7
DDLBi6tIRE0ACU6U7DknDYM0TY8LtszNpiroAiiMBPp0klH0VkttquWJa6Clyh/z30k30HTRAA7t
j1IjQ2LcJwVTWtfBthOQfA9ypyldaFG2qEQuBKQAS29ht0mCfeigwT0mw76MZI/IsMYkd3+7Dedb
jzTwQm9P3KDH8igGhTDCjjbE5893td+upC2HRK6A0zf4b3MZEqDJfSQlt+C0IN1ZXT2fdPvzfBjq
FJaOe5RWF1VbeeE+h8EUUZGWEtpZZrZ3Z46s+QpMhAduJ605vBe8a88AqCQZof2TkeAIuTKW5Slk
S8coqsm4NmY0s9cz3oTQ0tdhXzOfUtLT3dy4WpIeJ2mGHiKAaBIOi5DBNSEeooJmTp6O6OaDyei+
D3TfdmJuCFRQ4KbBjt1BMIW+QnDeRhqwV8iaUuLsIK1cqz96PBtYxoZHcDGWxXkfE3+kMKFirp5M
5blNkm/xepRrNFmANBZAvLAtaNe4n6UPq7lzz/Rqo9QQ2f+JxzhmQ2AZm7GC/M8yAYzUYWMk0HhG
tqzOJzJtn6uvLpcorsFyNcCI6qf5yjxvc9YtGcgHWA9diebevu+yG316QLDcVW2dgla3hR0TbgBn
AA+K/I62ma05GYAY6FmBZIoS4y4NV5aBMMD2cveOcrqHjry7RxtH2E6XNLyarOmryHZvOQnc9phJ
tqAiTPoxZ2Caf+QXLEfGs0DaHMogE1qMS/BFe4pDCbbnJJZxzCHzKj2uTD0FAy6fbT6n7ebHteJY
oYwhaKFOHhnlFbpFwwu/5M09iEhORXM27n+6tFhOaxKrlLBNyYMZpf4/7hu0Y/nxFx/CYXRh6blF
+8smP5I4Nhqinr0lqRvXLKMK6NEjry6RWT61ZcqaXqU0tsMg9So82NlVG503Ub/N3u9saJCogS3K
kH93+7dtVyRGENtnYcInA5nJY96DOwaoy9k0P3z3h/hjnZ02FQc7bSZoeDknRFV6FMRhcg+4ZfzQ
tPPSrk3aeoe1jLbzNa0wNACo143wiqrRsI5exAJOU1gZgwhw1udOFirlwgS3pe4RJPrae1Te+A/9
kUm9LO7bkNCLkhsOBAHkcovBXlErTZ/gvJt7OyHHh9rLpy3Dv/SPsCCYQxhw5f/ZqzfVGaBI6R12
sBC7VWR4ao6RMo7VKXjuFGCnh4KL9DbPY1nyJZttatI74CFSx6VJToyMMus+k05kKWLCBcSVhgI/
ZqxNGc2BN1iHw0+YKEz3CtxY72Z4remW773cTLDeNSIetrWiSP1EARRNtpxzhm8uXkraBKInUybq
CmLKK4AmgxlAWivQGVo28oEka8fDhxzG0FCvBSXE5k10m9jO+8p4FvQ4meQDdyLn5wnqP1x831sE
M2V4yLUpRgXlGWR/nuAdoJt6GVZDHw/NTqNA90TcZ92UyWagzZcTunDKLla5cWNOetch4tKPg5FH
0rgdtVqwv3RSlclczr6bUCQAVMw12FCEc10b49P7yUkGxhCBr/PhNuanKTgv/E/ftBzW5TIiTkch
5dmLXkmnFl+cSTA3Qe8vu60fKHfBAWuPsJLtly17GN+r5HplVzugLf6HfUBDS9LkhJqvxVFhTjhJ
AK4L7PBgrlYyZdHC/XFcER/4a6EJAmHbD2PSgEKlDKi+74aqaLQ5jc+5F4v1jrcYiJKpgGsguqIj
VAbIRc94qYibx+uOtVHZVoDR0tk/4mz1dCKzuTyqzhQ5mv3p+S2U1d3e2snbFQpZSKX8PYU8WFYP
IIfkd4urdiPNpu5LgKaggGVg0UUtHLNZsZ8a3N40QYJartfYvlFs97Vvl3msBsjeTgJ7+gxcT5yt
S8IZf4jCatcJ74fW+JthbEh2dLN/zDK5ob6ZeBRH/AgJ8jGBFeLNI6gs4vJo6pEHmm3EyEqky+gv
Auf94GUcds/bDNzUXETg7EDagTAABfDz+oI7D84a2ldF7i956LrtatEntgaO2Z8dh0tCJjzsyPSN
1Ev0ar54Zn1blBP3IMTBVzvz5QPT3X3Qw1afnj2x9ufFu0Gkk0xrumdmUirLeN79RXnUJP01fBj7
mwOyf/eeHDrML4PKGK95V+q/wqryLhJokTZKoeFPPGlH9VdFf/6r+9kLiKdrORZQ2zd9ajUSoM4u
/7RA5nSofp86K8EF5aF0Cvpfdo1mG+Wjygb/EnOpNy9Mu7qufRZwrX7Hm/kPxlA0RrcC2J966Ean
l4lWyFyEwZ6uFDJx+zCMhcvvHyTbgGR5Hd3qHrE3l9id1//Ua5mgEDAYycsPYHAjvldzhkldrN6L
KyauWLzeI2QsSNp/+kqDBo73dRaqMq6NlDivHj/h8InhFgDLIbxRg49Ds9/UtS4gIt4C2edhnTe4
FFbOWFJ8lT9yTQtjYysafZTuawWVTcr9u7vbXsSIPzcKkOunogU3c/S4PBdatTNv0WnX8xuz+hpZ
45xWViUbac4uHW9p6gWIW+pY8hRyldC6fTE7X6Zp8nrGMhQLwsZjnG1wbtihDGVrbDa+YQ+rd57o
Y3KYsy1skbqq2Cczhazq5o2RvpGU18TL+9LnKiaXbiC4iNiNP5yOto5eRtAEvWqDCqSZyY6GSz0f
1OrQuxAls+r209TSqZObokD9gxXu2hYk7c+3VCVI7wN8FeqIPrdlOsL82npfDcQk0oIfLrTHmKoZ
R5f5MYf1261NT2iNN/HSGvdRqB70DTDPVhy5iVdU3ivkv1hAZHeOqKBbiQ+ML10LaqekK87h+4Qp
exXAxnX3oEWwqvt05eZ77c1RMzqG20imzFnfZbuRtxKWuDzy0RCcP7/yFwmL4dBL3q2DmIPcCkHE
FxDcOjfRk3kt/DcHwsHeDTUqkcILLrsCaLQmMGEjgsCTrfWJVATFNdWm1jTaArk/cKVWKMNwYQQP
I4/MkikGb7/ydiIm7UFsji5vgITKLaH/rpG624FHHP44byc+R5oqESzJ4ECePjSbEalNAo8MArih
HCropcPZDgYD7YbnaBqGIOiz64W3NFEpKAvNFOT6ZVx9Hudw7U55MB5edYEnglO8Jzw8MF5Hqm4K
zJxDdY0I2nz6Iq+8J3JvNR4LggLdilRs1UcM9Yvzrj+fv6bEgVo7QC1MdXKEIDUVVVq4t/nLQAzs
9+JYHStZ6L156MXmjxffj1+PtSprS+51XUyZG89soXbzk2PHi5jHsKs7yO0AUy18E4sASe3AV0cS
Shxb9b2R9xd8jGwpnDDQyz4jm8MWcFrIPB7G0FP+YtsIMCYNDtMtgkJSFlyEhpnV3mnFko08rXGj
gGe6PrKjITwX+Ab9jx063C9MP+6HBodn4T2t8GE6eueTqzvpMlC0EBjXz8UVJn5eMMgLAXdx65Zi
SnoJfvoLN9qN8bHyQFE2d0r2m39gEVz6uHN/g4ZRAATeYznKnXb0czPGGaZPj8wjMAo8Jv9yWmZR
BFH13P2B639uHxmZwqC2b4BaBE573yUS+w/fb9eklg+l8p0C8Fys03+OXqZnvkHBhNoCd45fGVOI
PRwkLcrXoNPrGQZk/6fWdsEDpgXgDvjvhtZkDyn8hqtHBPtsCBJuD9cWCj6mG3quz7rxQmCbPKLt
ZxYCXkRnQ7CRJxSqo+u7ydyh6GNOe5jtpDY1BemlGKhPi/m/aVsF/yPv1NKZEJT0pIGs0ugV1lEF
JkLotPLa6Y2ASbtdjmL0XNCakmXGYAK61SOvqCKHKU6iloIRAQ5OKdo08U57hWWl/2cDq3sP7ywc
duXi6/sU8uHMml4X336rciMjqUK5ni+s585MVlmV3MY+WG20DuIe/Kkmn923NGpKPESss11qaJgS
Qt0oYTZT9moTaaNWBqtyffmZL4l+Vlc8Gx7aZLsPMJ8FWRlxdlxAPXSjPpUhRF9t3pZFMJ+PeIoE
1uF07xdc1UDs2D+8xChv9gepGvfWzmkrjweqvyJg49e+sliXCrpKmRMD46qJFj5ZEPJBXPHNU1sG
x+yJ/y+bu8drz00hhX0SpdSVXIrJqx1AAhW0PfB0di9HDKH04+Dsgv9s3wkCzEk1jMF+Ypcg3EhP
nZyyBD71zIwhIQrc4vSGv9U8iqyEEeb0NYvjiZv75dKSxO1jky5VP2ie1kCfKnDFERGn15vvo7Ti
6Ru72O4Zk3idbH7rG6hn+6Fo5LAAjylF8OP3tuBewPuE/sePY9AQ1f5kefh2Qdxjf6N6X8HNsUHk
5fuwYWujesqgnj19RiR6QjGcash0NkQBqgtlheoIWgnR/LGesmPCx+nnxXrjvMXsqTQWqM6rUNwq
e41SRJnoEy4Yq4MLiD/4NtwMaCKOWfH/G+nYDg/mtxhNa5qYJF8GxocvP6o0nXZM58TzCml5njxD
2BClAjYQWXRqNacWJBHjlaH68mT+0vUmxoyNBWOs2I1f5nsVhA9l1Bp/922rncTw41BpWc67oiSU
/c0DsyDU2xL+m99t3/mnrHLylQWH1OaOo8fYirppr4pTQW0idvUE38ZG5Hk3+86g5byHes9bOnfY
UsZ+68sccDnQqK8nZDfZQd7AbCjvFjvGETR6eobEnmhhcTXylf/iiimnSYFUcGryBXV5RISbwiAo
V/eUoavBEs/CjF79iB+MwGrIPdc/POqkVDzX1qV5FEzxEKM1lsDP5TEhM+DA9Cos1TRCDw6Ti38M
sYE//1ytA+UAumsGZAq9iMDTy8o4igSyI+1pU0hyufAQNHJr2SaCgwQsOenxA+3u66kW+ztYjOdr
EPjCYvit8UbPwZnbc0R62f/kixo3fWlklYE+e7SWdTyGfm6Aoh1UPCmM5Vrxd+Gv47CVB1jjvj01
dpwfov6kXC9jh8bzAeP1MNBnf5e0kiNBmamE0MJYVOQ4PfACeyubVl5O1SgOA2Yd76WJgvNkdQQP
IzgEdTTVFnHGJLnPlgTJY11WnvyXjdQSd6OUn0tlNkdTjsY1bhlQZoEQuS1EvwFuQS/qMC0tEIRO
o4gyPt0tR8SHJiWT2RkozojvbdEmLy7NwpzvSYrrzpSJALkLEqKLnGmOCAdJXRIBOefdkbkCHUVm
6MLHIT3csudRTaxjwOiYdvoO8OQuktg+5ttgEZ94ap4OtlZekPJHV8M1mNR3PTHj1T0J9LPmjJnA
iH1uUAdFpZXe4C5g1ivT7WjkondsXlGytRz01VU4qf71wCZfiRQaS5MSJjUtzGSsxoVfUPC/4lEI
HKphoA5DRRKVvRxBMdfBxpR2nMafr5I6cxGNTq62QdVopGO3SvMTLJELH4Oud/5i13TEWFhgtaie
a6s2OgtDgtMF4tSlnNZAAk/4HROC8CJj3P0MAyltAyzjKnkrCVVoShD09TsXZ/mYqR9QEIAdDoFq
Tq2Oen949+myP2W5K4Ek4qFS5BhSFycK6MU7cSKeJnyy/i2dc3Q0AMdbMwEqgOHS9nm9slM5AD2I
a6MLFyZRIx6M+PFMEBQDEXTWnw3JDHBaGdbC5NK1Rpwx7x98dP/Rx69RuCs2JSkbzahGtKNyD79O
0DRwKwk08ie5MUXPU0X9YdasNBTfgsXXyQbObIld4VuK8d3mWDrhqrTyZF5MX9w05FjTuHJ/Dl4I
a4KjyrZLoMQUKvZnIUu08QXDZPf2f9OtQNCeOaFZqbkjrHvWqP6G3yZHwWltmzjTtnRaxv3Rssts
nRPmCdyrOk62YOVsUwjlB19lUeKLsS7YTaGlSmjtKzgPB1q2Ght4Ve9NCfTYu6B26R9BP031fMqp
cfq7YfEWF6JVURvYfIv9e158ZWcLvj0YuwiPIBN3n7NpGFALIvqL8OZqAT3e1R9FBusrierX2Z6L
My5pO6QQlXLwLlfb8vWjv5MBub5ZAt1kxLUAM9zaSDz/xd6IcFfwPzH97zfVcVW7h5Eaz4ooJXXl
3CcKg4lfssSJ9TxnIGXh0JFKe7oTlCswgZaRYgN3CFns4CpT5Z2WQyKkkEJTC4ugH/dAyfhiw9KQ
WcS16kBeREuU/8QPQAs6J6ii+a5tn66DMiyIhcJ+Rf/NkG8YB3u1xMEx/82G9C7/9a5n1EZ3zp4R
nEC52v5T6Rq5kAxlxK/2aCFU2r9YaRw9b4zvKYi7Nq/qSO4NDhb1SMwYIJIUXYC/lhXrNDwE3BbU
uJMiqdP5dD2d34Z3GobKiyrVsg4a5XGcbHbOrWR9sQBjccUs6Bj6Kr3dOCblUOTDujaHlJ20Pxmn
QBWeyWMfS+9JPOBUMOMSYHgnWhuW866039LzFdkjLRnq8zUNDlphFJtIcEu6WWz5IfWWo2CguuTT
Qzaa8XXBKgv4A7W15acBpAM09+ARbZDo99tEEwMGl+emYjmnsShvixV322/mtoYcKRvSRV/0Ugsl
qc8OQeEMw8J8reqWG2QW8ubNv1kiW4P+AjZhuLQrqVILzsJshWBDv09U2vRTZzQvxJDxvEMUyXlx
Po72CDacIGnKmmn5T6g9kwPp50jSwREeuJ7YYGidXNqFnX8ZzL6ueyFgrD146weFc735yCux9pXU
oYbkaPyYLuametxgA6tKxzbfAK70yr7Is6XIgLX3fGVKHKsoAyByW2hkiuqDuPUOGx3vM0+YVnOG
I6ecEcI2taQyHshsnswpMYObsbD3JMwYw2e/9sbrDIqsWHZ/n34FlImnDFUNch9zyRzM/iOhIEMx
RC/E8FWgu1kpWfbb14PMe0B13NLpwDrTR5JnX/RbcsxbImtzHS8mkrIWpHIkh7cRsiZUPEsYv1Yu
bVUKMmZQquEKeIaXr7EQiEAeJINjNdPt7cVl6pBu1gTbcPUSnSM94pxJ1jFSMmE9JQnNpmwKMN61
U6RSRLU4tud6KkuqnVFZcfvCrHMnt3i9iRNQJoeiVbRPidzddwfC1VWItXDcFPgu+hMALFBEn9cI
U/51ZQruFQVIJvQjVp+sbidgEbxIAbPwhzTRgGAmmsLcixCFhJFyGwRqiKy1/cifsl3d8gdhx9Sx
Zd9ZHZZqBNKNnNEzz3tHqRZiBKtmhzNxNUmiXD850eLE9UWN0f3gsPfIS9P+R8F892eRzNS/dZkh
tKzYuzMi5m/1HzyWO6cI8NnybRKHH65VcU59yf+tLeYE0MlT3H9cZES9dB3qmBBOrm6NnoHSpVb+
ayBza7wPQJwfY0yX5BcBkN0VQvQfNn9QPg2RdJEsq75emF0/BGCyPZJBO33vWhoBGy7YVRGG2k3b
+wvkWoW054znF+1j6Pa2/WQPO0fV5DkiGzUmUu/tSukr7G5RvbV6cD/uaF7uQX5ByjiIyeQprRS/
o/1FID/3OGTMdtHSC6wmc2LrLLj2DIm9dFVH7tK94mn4VvzxzW4iaJuT3lTEeu95RBtwnyof9gCC
YsnHtCPgSEK5df+m9DZyLysS1vMJiAoalrqqjYWgaVF+cksdO3i/iWo05Tv4RDhqyUhxKY9SeDTY
fqXnWmeL5LNlR//w58ZMZI+l7czycZwrZXZUkUpY9kQX2R+V8AjoGTj9D576i7I/OfTB3O/XQNI+
M8VpoXjmVoQuwXkftq3i8r7sQ8XdEMDigB7D9azCpZel7d0f6JHN6EZ3S1KvuXYsxcJ58kZ8bZhI
R09prZwLXYnhQl7V3jegjItWK4YwNM5ptRFuktIwZq2qYITa5vwKROWYNuTHkhv8tceQUkNUZwpd
z+sbUQ2LO+e5QAmbrM+xrb0vyilVfejUbue4Y34IJjNz6r4mtVV/y84h72lP2rze+z5w5Gi95SOx
Bof+lQd5UFz2QqeQKbj6+bdYq/02UTriI3i+DJ+JzXcjjZaLsZiO3EfDcq010zl9bAS4l3d90fp9
nqvwu3/uknMykR7+rN+rF0pcX7HQir4uaw4ihlZRoF3kru02EnNPQ/S2K8y95rOPpK/VuHxHMwno
2B7CU8IZIBLKagMyKGVdOELT2iFyFT0WpvyyOXFbWJBMaUHlhUD9sZ5KQXMwW0xosiSrAeY+QEEm
yPby5dRl15OMnSVQMF/2k/98Ph9H8T2zjJ58HdHrrmb/5OGRkPM6U5K5Ki6slJaN03v+sxKybwbW
M+ysnDPzk9b0uqlvwzsQXXkbzLXiF/MtScNdc/mEvO5J890nTcycoTUUqnUA44ZNyFQVozQTf8HY
z4C+Lww/7sBcoab4yY2X5eM9/LcBjpemmXtqRQz2Scz8ChoeV79eKTutiJadpQepXX/CInd4MG0O
Pzs529LBElzZfGwmgM0ZA0F+htmraiGV1JyIv00dbnQPiLO07vgLM0GpF6d2OfUL0eKIDLRGW9A4
WLhEQLIZGXfnWmB5JB2vD4zlrconFWvi6AWc9Hh4pUYZkmpnKfQoN3F7Qchevzpglt6Atnj1cs8h
Y5QaHHqy0knuqchSkmMBUmT3rE+Ec7Bf0KhGLlyThdY1QvjPWvc8YIALuKkWPsHFWRNHDI7Sau4k
AiYCLxxsgKn0sypjVMuDzb8EVhLgpB2WtNvmBrZ0c4zQPUh5li7+Nsd/Zh4WJRM9vbQdR1CdkhkO
Ob581SfXfn5mBoTwK+jMvpR5e0ufLylc2/Z1u9zTdKZ9fpeWkGf8EFUy/tSsZHB/gwykMLsWlezD
RfqLiCCJUM76iczbWAJSBXTMIHnThtz9ym6akQUKm1RHYNMtZKi4/koRUTL5BQQBbWKr/4F0oCbQ
mWppZ2TD3xm4wubllBGvCiPPooUyo1vTD+VHA145y4B30G0DpKikRtodNDzAHkXTzZqUqV9d/GP6
IxiuzvUq8Hc4PBRHY8tQlrJL7aVvZACo1CMbxqoXybbrqIZ7wnoYOAHUN5YyoRvactvrS1oJiehO
RKuk3G4O9Qg7TAn4AU3bvlIbuX9YiUsgXQZKNibngI+HaV9m516+DR929FwGrA01JhTZZ12BkYtm
GBDecYChdF8Nv4NCA42jwc82O+nFUgyMlxw0mj+h+1/oL2AJcESaonqwz3dknUN858dSuYSMf3RE
Z3M4xgWGuvugtt9aoruz9CtED8T1FyPCRmEzNAByCULo6aTSTNQVYIgFJrFayDw1UrGyvnwE+Qyq
j4+WFwdgYKVu9+96P+RsADD81HVs9UWME1TpACtkShSqOqWB1+cbLRQnvruWX8ERZkNbuJeRWs1k
o3ay7KJuSQWQuRabbM87/uQSfFBBf+tFnfla9bqtU/9GxEBE+l5LCayPhVLu4TZBwtrVCmC2ju7d
BTJANJLlSbwGpVyrKEVvXVEELWykiXGfTE373MQ0/VkFXlGfLxwrN0492GVj36PytYQJaHuQiptz
6sWRnSLW/xVYEUHpFGP8/WhlpeRQSgcrHc5Y2leE1vd8e990kYcSrxQLReZUtO2Y1THVWxASnax5
WWDDGQl6Qr4fury1moVJ+AJg9yccL9vrdrihX+2aFxEokxFMAGKdPOAjhDBIYLKMV68vtI/iQiuR
zztYWaYSC+P+3tJKekCAn8tExIYh1RnzucJ3pd6NS1TLqqW9chfQGhz06b/JNfT85dvKhfZPAbGi
assnAgU+AotM1Ql2x59k4auoDZSiFMsUYfzEDCIIv9TMnY4zTZzlv+tulk/2G7bFJPh/MDaKq0CD
z5iY3u6MLvLdY+uzbrqTNPMtjQNxDCEVZotZsj9vlLr1VtikypqVJF2S/VOzb6kw6bigll4dTOWY
uIdDzITb6g36E60xACCAq+tdJ0C60CyPsUJXSyOjYo3bUzY0swJIo4hMezlPNFrVCnicEe+nQbgJ
zY2BaHkNE0j5ddh8iiWAp1qj0auD2FnUKeVnj60TYjn2gLptvnImNc5UetGWzmCCGPOuOK2giG+w
HLXntHXj4SNfeM5locuZb+3GNOd7MhFZvXbdrWVoFU3/wdMsOZEnTWSpDvVdZBbEuScbGxxCPjJM
oKC+I6w3PsXS13/IoU7S0b/EN7AHcUia8iN5WWoVUGtTU/92VZ8Ne5MWLc/XzB33F0Ak1kCt3jO4
VTUFL7RfUutjQBZmL8RAY5DINJp9LNtld1367eTvB2ckNP3TJtnqPu+z7hs4BHTIrn2bRCqcEYzC
Q30qbIj/Tsf0nZ6D4be+ss9Q+nH8Wby8K6+aN9h9GP8RcTBdj9iz5dfjt7p8d3WLODyZ/MtEsQWN
/GUM2Z5iiTa/quwDeENl8v461A45g5cVUFQXDWLLIhsIyz42aS+l5CIGLyZzcrbbMV5X3VizwMG8
UqdiMsW2mKm1izzhxKmByPVVMKRybherPsadzr1ppV6OX1pR3UlLIth5KR3fsp8nkVM5vJzYCs4A
7U9BksPuckE83nYB8WG3mYQptcqBNalH46hOoNXOaLwge6Me3HZvDyC6H0VDQnNChUsBBu89+nfL
p66I9LB4adaWhQA+Ew6OnmkmiRBnxRbcae1q+rqNS7xITuUxIu6o3oVJhcgPthfMKGiuonLAbNue
5egE7D939qjyUa9Y23Z7sglPq2YpYarnGzhfZUXUZY/oupYjs/IrpNt2wQXDpKioOzlWUFf7rp1N
pB45eZVExvlXntScv60WgqWJcvyrUl5TN9fZ5wrXgkp9WWBeu8d75lvKlPpwO4P8Ja2jQkDAAvL3
C45+1C+9j76BiO/TvFR+ERjI33Up8ZHjRyGVXDnheQydF/dAwA9r4HveP6ttIWSbj3qOo9dmvBHy
ujuWaHizVRcSK4Vc2qHGwmxFvhUrtKsxwbNBzaSUx5c4sZzFs/IH2X3gBC9UONxAQhAXm4TEOgZ3
5jFwoqVXeGHf8dLGBdRojyPSIh/KrvAa+SMVL5qPlQS+MQ24iu14KVVt2cC3dk32I2iasLyTPkcT
OU6hY5QKG2Elh5FXqN3YADzDAMymmVtXml2TgORyuI1FFq5QZOevyAPG4gvi8s3gCFhgR+/foKan
fK6PfREeexbi+TbnyU/pzP4f6HiEhMUAGRhlFuyjntihSnmjtufR8UrJlH5uyHKzlzr/ItneLchG
ssJF4PQ515izZgI2AeYti41rR57IefsjHGZt04kM35vXFtrl6FGU0wuISsmHmWt52l8bctFPxIFJ
U5G+jIMwSWRiBPCe3wkusJXFrV2dFqgYDAYz3JuVSHYinsoAJ9MaramMgz1EvDQW+SznbPMRI7nl
1egidqNnOGRE3luLJRUoejkXaKqrrO4mZcWq08jDI/CtdnkOlaqeq4Cr1f+rKDCYz0UBTautG7yo
CVXPB75I/H4t8uTVW6Qmfuj0H83xH3gcabdXRhkffnJBZQu68rwPKvDWXudSsuyL9AVxR2TlYn3S
7cMuDy/KIxJWkrgR5u4lZ8kMyZ85V1ruzjkZ47dQ0w1jm/GP4V5NVH1JxSmvETolpoh98HiRBC6i
IVYGTM+K+5bEctPRYFqxDRip29zNJ2R5q3UrBc0tkSk46jj/Ay+K5rO5GGDvEOZd7kTgqGkyijxX
0e+w1lJ0tsWjkOHoN1vwXtopY1jumsa7pyURMNxacNg5aBW1GTLDXply1gTS7NDKRuYiZmu+8qNj
r0RwAz7HDkVrjq4SAl4u4acHaAwfVDFGilSV/YnU1QPz/qrVAUmDmI6c+9lueHZsNBZJ7hdUckOV
DIDtU1EjWhYeOMBR5O7gJ6243nurYywp1+TOa7hKM4Ttbqr4hFoZ4wOBgUGUzu1siswCkFilpsgC
Qj0GEUURkY1hSboucCBCeguVsO0HcaBWZOFoEyAW/2aw04naH2lCc1jB/OIY5OPPQhcGFsoyHXYO
qVUuvBPQKM6B3amikPFZZTFoLHd7msnMPwgH5IzcyBm+mnbsGhgqWIYl+00McPANiNls90SIreDl
3y95ja1JB/vsSmstIQ14L5joKKUzmwCOg+4oX+G/HglNT1DDBP5SVXxbmJT+Z8uDebzFH2/R457C
0FKV0pNwtpbn1Fd0WoKyNeQuNH39kdGmEE6iV/kelz1Cv69TKGEARHQMhgDVReQIg3b5u08nctvB
d8Kqy/HX60gV69o+zRJBw9t2/KaqFwBL9oYUlcTmvqV6dXU2p93CpP5PbYiLtXNWnQjj/s5J5LOM
2c4ALP5tQtB0yBqsRNMF9U8ZBTx55zsHp7dU/PpUXU7DjMQgfRN/IdID3iwCIxnHZQtpTq09+ELN
4jzFnPO4kXNEQScpHXW7tGg3DqLhIRVHlpJ7jTGsr7ax3G+pZ8Q633S6yInCz1zlTw6pNFimk50Y
O9+CD+IW4KNJGTNDy2p5fJO+ffa1KwKVbOAMT+eRRvlEoobe8sphhOWFINIZrfV1riiKFnFiu4PH
fPfm41KXLzRG5ILD4M9Yarcog0Q2usVo+iEpOiXRWIse5OfbsEuLJY3Cqr6oOW9okDkLwnmuTcIf
zpqiBZUlqozwDfGBSNr1mk4buYzd6mxYnfRxLFksCucmZ29d9tHs2OZSWskyjDbRSqwMzoYLmcJq
j8riEva752mNonALcekseOdKtKUKM9YiqpF3Q/dZlHJyk9egmrPIoaCpq9fwMRXIxyO5M9Gv9zlH
Dw4iFk6Hn48EMoDsSSN0cZS1bLH1jU4O7e0Iu573T8heA43XJGQ42tA+RyTBb35RwjhpdN6JfxsB
+d/eynJx8KydI/bSl1Me+6kmYkSMCDyR3lRWP7uvikgQoMvFR25fxAETwKRqSEzTzH43UmjfceUT
ucaHdUVnhw9EbLwem9rKdYjgRP4I4RCD0M/9znGz5vcRfEDgaF6mYH8DZW70QvjznANvUMWMGLTA
pGxolTPM8LBlKV4OXGeXu00jdkM5v7FX9Ik2peueeiCK1wuRsTADatSv0iM2Lm0cOBNZFettBeMN
kkhIUleK0yaBdM0cH3ypBr5AJ9AOjaw+h8WkcoPj9af1yC6VeVIxN+hjvC//BveqTJIbXuH0zz3m
J1DBkBe+KkElsTT/ZhJuIPw60w2r+I5ibfK/tRvr465kUDh435AxnNFFLiWU4zCkSkgyJ1YLKEHU
4iZhJX2hO4HlzxO6ObiD557y0oOzv3BD49qPweva4ZDv6ZFzMN7++Z7cRa3s0BsJB9sU+9rAKxJU
bYX36IauMCIU5pP+kLlP75aaBUfnvShJVb4l4ix2gBztN0uAqhhZjBSbVc4nBcBRBpeFbWMpQmiZ
8yr4/r75Crl+B1I4iU2crUGea3b9hyH0gcUPduJLo7YPYa/3q/djmqWUmEerSCSGz9tdfI93jCdj
PnPjoLZzcYS8aAQfy0ZX7AworH1Rm+lgF5LuYxOntNe9sNFJ8bwNyfgablRJOcn+NBxhFQD53qoI
dRsIxwS8Gp2G4/5mKYTWAUgqQOSIm+jdnFKO5dIIxuycFZ+M/CaI3mzo4Qbt2sXsRfDBKj1Tj0Zi
Q/By9JVFplyCxgUg3wt+62ENEVv4Q9EUDbxEB77m8iKy3W9PQ4T5/0bERQ/GF1bqU0EIUNfR5hPZ
MlXeV0Xy6ynmbteBu7n1KFlUMLU76e2VTf47Sjv/E+IF1ku7NNwgiQgIejYw9q4DgpWngvWZdFU9
wa/mdXg77c+Y+KzTk7GoCOlVyBzbPnNB8UuM6rS2a1NWn6dWe1tDIXSvrChL/7a1NqiM3/3xLqeZ
qt88SP2nuYMhlO3kDHHtt3E+mW70u3flsDBUyeAYgP97mvNH8T1NNZoD02Jz9T3eIORPIkvYPnAy
4ckBV7voRjwp/N/q8+R2yGVUr1LpOfzp20nBRAmm6HAKPkeB6urgv+0rd77UdumSyiMCybxy58sg
NzFN6+bV+y0C1PAJ+GdFdGdLEP0ZeYtiXKE3nIOOVwFrxnXZC2cUdvvch2EVwP2gxqIEOU/ARjSD
mrs8Vs+hdLtlpgdqy6EsSnRiVz/cm5O1Cy29hAmhaPTLo/X9Nl79xUhk9fin33DprrcPqRoYj7Oy
0HQ4KS/nkDM3LKmvp29Faxq9CmhUBuOHBnHYo8CGmgnAGWo2oHd1CSjqYUG812RL1nIA/27YGOL2
KQ6BT3Zzlg6bRnKr6JK/l9cRbcZbiz0aH6aMpmOTZF71SjuzOCLNfGwOk8V0Ql574DI4n4Uw8ZQ3
Lm1HEcMd4JjRHr0dCoq6x4yk4s1iaMDh2fVGtQyu/IYiZruGcB7q106IFXCoU6QbdB7LLAMdO3du
bf1viSFmARdCvptQlwtKd0k3/Z86bulY4xnP65IYm5O3LQY/3EMbwzev1uz03MqEtYKW08PTq+4V
eH68lq4I+y8V0A40tY9IOSUI/AEQ2RFev49vnVV8LbYsxroX2YlPEOGDZAMvfcnOYXtyP8ZsFNaY
2W8dh3Mptqzn+w4jdGsDVX+ZjZwrK1qnR6/osk0ySi0VlRLVWCfv9KeLlTH6fPZkFFSEpa3U65tM
1/WHw97dXeIv3bAqzJyCATAU/yS/Xcwsg4rHon6M3uIHuHN2eZ/VqkTxbLEBVofWsZcs1rXwbVkt
Qj5rc8+OLu6U/0tRYQxBDanlbwJ4Qi+3atHEpQ3cXhN9XV2EyGMgYyO2mSnICeDcrrBnLnPmT0bz
eNugVAer8eSE/9vO7eMOdJmbcX1fTs+DlDsXlUsQQyQF58Mq2eBYWrzD4r84ovN8HAsIL04Qi1SA
XzvUdRXhmdwJv7Uf4U4KyGAk6lKU6FErHabOjzuxH98aXs+2J2FtSX5vrv6ynf97a3vjbn686Y3H
0h3YdvxNQdcIZKXpGcsXVqVFm+PtJHYpHNHjXeI9dr/4CaxOTWllef0u+HtMMwrdPMBLDYD10w64
Z5oa8N3/ZsREk6aRvY2fw1vA0IDlE4Gno47WFRK0mSt1/Vsglq9y1JmZHxTVyeVyHd4AfLk+9Fsf
KBpxVsM61Trz9HBdq5PcLzWCBk+K2RNFkO1eDJLvw7NGgx1lOuaOq3BqhI/Y1u6b9FSDguwC51fo
UJknRnxWH+vmGRloapgYDDWYpv3ECDyGa2+ftI2auKUIV4ioq1BNZop4NoMtHoeJScs4wrzkNtw9
JdclxeifIPRpE9FM9EGcefK8geUj7PkLsB1atMZDtAIDep2PpmYOcIEvDWtnD5iiUjnM6ZvfqeIc
zsXZEcE/7uHBXkP1S9D4WiReuaVFGPcKq0B7yZL1nWtSSOmtmR4XBLvDBIrl7YB3QScdycWlxCMC
Kxovq0BmB0ax6QCyDgjJJ+DBasyTppqnTtRKddV+skdqtYd/Uq08eBQgFoxUpsOi0yyRoumtozlX
dYhlDN+LqJH+8IF/NKRrEZe6t8LiwLZ6ePb+0+t85ofwN8SzfRI3CdBoHz+R0G/1dip+Av9R7DRA
t+KHfyQ4HFxol9NRisUpN1WgEU1FRLX+SomaDPOVunc2gbpe9yZxuZBGpvIC9bnSTkxHUqf+WN+2
MbHWn/bv5hp5LiF52uxNaldbL+NTkLwM25W3feTC4MXBmpI8r8K9ziJlls6fcOlr3lWqXFm7s02R
nXlZFbl7pdzVwytSacYZkTWCTf8f2ny4NSzOUzXOMrX8+2qCdXPamVvISwr1WxZ/e43bEbAuFILn
GRg25E4LnMnQz4x3zbfPQhZ/X6v9xhDlEYgBW9hME6MDtKhbe7cWOtwmErIRglIClRADKp4rRklj
PX38l6p0sA+ZioQ7iU8/phDnnHV+AmiVuDX3J9Ro3OyWuDoC8gZjFs9/bcg1mlmtYydfr47I8Rhl
YXXLj+LA2xai1k1ckQoRTnG2XhcNCCmw3Nll5vP8jyXyjFXHrgXJcPehGW1oNqWFHIc655W+fa/F
FEpg3btaMegP3gNy3uFmTYgZ2DX2nbwd578gl6urnIaKchFQPcUJBvQrDz1+gAa3jQz225x7YC6P
7Y23P+YF2q5DyZebiHAZZn9E7W8B0jOXRuGgtqfjxloc+E7VrC+eCpFEAQbsc62lUgoQK1N3Z570
0YYPOAiF2X8TI5uel/HwGZ0Ka80NUBKVcr+kn1TZkehVHKrXHdzMJ308RQCm5jw/uwwuZCNesmJW
A3mbs6uO6v4+0SRQ9gUqU7NIIhQ4hMRTME30c0f/sYtGvsG28t+7PjrcFThevAwRQ559ih+RcN26
tjVPjaJR+38u8ELAP+IzHq+thlqcvH0TF0h4RBu13LE1ZResg3EslDkHjfUXyj4aNfl8NvcSPMwI
Ge6rw2Ibs0JM+xAHuHigvJ3FoQNc85AUndee3qChhrPictB94tIxgcxt5SuWFCnZnQYqFpa1eMTR
NzTSBJewnjpsK9irkliRd1JZQx2LAwL09VrH8f9UOcb6p+4dy9M2M5FXcz6sgEVhUUo1CrWQGUcq
4TSMlAk7XD7q0SfRpnR9rJCcf59tozR4wzK0EdGVSeEslJsINWk6/a9oYnvCEnbJFt23chI7yoJz
mvWPefb3Q8B6jyvoZkOm5DscMPH5J/AF8MC9YC9OWkqN7yVG3/hqPbNC5UNKLLAbL7iiLpx1WbQI
vHBHYyV2XnCJI/tCDWtaTHPWFN+I1juMEwC5AtBidbBfB5F61d7yKobbTy9h+4ROPl/ChkoJNg++
JP0sB5KClo+W5j9aTPmPeFKEBQW294RBiVGhcuMq8SEagH86gnA6M+2KxmwJv9LNHPXEb0kvEw2M
BwyYFJi4QK7fHVKFf7sWNMmluluT65Pg6+gMKHaDRKvqZt/380Ug0cVMMiuTeJd+Gskd3BVm4OhJ
Lankc5OwV+P5Gc7wAs5RGhnJfIgizeQg6C+ysLAVBIjDPGH2g1J+EM8ExHnrjfphWWgnUGe2i2mO
w8A+KQzGBcw51JIrWz/0GJDoQmYGEiTeBb3PrLn8OfeWQCvo0UhvcaOWhqdar7sLvjdHk0tKeLY/
GQyJZ93hMdSYHJgsCgyUI72LpQCJrg2ag469MoatDSp+VYGUyWUrbvtfloK8VgHPIAWDMUBO4q4r
CIRDN+ikDeA6QHNabwrA5cPf9AA9wRgPx1GQARCW+in+2HoTuQeuPxI5NWhlzCDuAVk9IDKlMDWR
WjsYTJb2ZCkGaNRwWqmDLEyUvOSrDkhd4tcHQmz7LTDEZxQNdeHCCGIFBiDyHya41dxIq2+/At+u
ITFqfLWnAVgqt3TiCwkY/CuLEsd8jw7ADSBVMYQbzEZLlThHbtkHSL54OsAUWqtTegMIaO3IUpeh
5F+/FT8A1rEpPzebtF9Yc5Eg3uN8vaPVDwvXa46LsURcrwkwLYuGm2lhwLq2TLE8Z1EUeDZEcML0
1Uq5UGAEvCrNZDYVpVYkKxBZ/buIL6Z8gkcvVqLvGTgjCmSJN1QoaBRFDSRSCaNjgPvUVo7BtyCa
PkD9Dju96H6jjKez1Tqdxs4Nx8q+rfYTI9+b39xxhAmux46GOu1zUrelPP7A4sOY1QVwrzDVsErZ
Zee9V+ajlFvPyQAI6pEk2ql/p4i93pOI+hVe3sUyNsMLEE+jue5MuBy0XpQuUX3ZBZYpFH/XNWoy
57fnNKjaJQxBeF5nxBnSeZrx2jfcTGOVaDySwFeMVsb72GNzscwcFGeLFTezQ1ItAtIkCt+6iGvB
yD0JyiCIKebZYh5E3ooSCuheuwOU8LR6988XNzI5kA28aNgetptz1LgB+RH2WUHOC4OcqZwK8/3i
fW0ugm5XEb5lZq2MQbbWHilrxJhQrAyE+1d/w4YER3iUBzvJMc/jCAk9x0aFB74WxC+isiQRW+2B
WKWV6Qp5EUcK972uiq4sK9clU4ZIQ44VZBigQX7piZZDr/6fuHoc9RzOivHtctlK5/COO0kd0fiB
2ft3oxQmqpoxv0e24yCq0FOt2MxelxT00tUqn6HYUGEjVni81wJFF0IzlNGpOQ7Joem8InCfBADu
SklgEkUzIYrv7WQY24J8fNXtx9fbScNPRIPOB1dZT+q1SoAAY93+ncHV6D6fXg+SMxmO4QHpOHFX
VZU/r8C/7RaqR9D1RY4Igr0dC27XefzuUdjsWIQfXusSLOo9G1hmN9qd68M86b7lUdzzqyeShybe
pjMsXSSp9Oj/E6Dn3R77j3BcqAOhXxne10tuKsPm+sRAoLjpDbcMdB3TedyQc+YrKJuJHQ2yEIir
liLjn/eTVl3tdtmAOjxKAtnne6p94DwN4htqrQkOY7hCyKhWK505b1TpY6kdjku9T6M6z6AH7yHU
zwDvsD8o/0g4qJX0Stylpl7aL3nz0UIgYGQWhXVeDcMBCAN2aXmj0Z/2/B4tUsYGnIKNb8FrGizD
M/RAm0hJZHd2gefnzAmnlbTz2mZUMBMTzt02ZqnhCMEOH/bGfSfmPwzoa3+i1/DYhXjCd0HK9rx5
0sep6QatLcCwSwkZ5I+DKJobJ7vtiPqJqeU2GSAn1u8MUN+wZpNBQ1XquEQae2objPViqJ18Hzi/
brOgThg78/tvTBt8XbJWKQNhVPGdyKW2a9N2ZuSzmGU5oRvXnAFK8xLEVMYuCscCSL3a8sToSrMT
/Focs43m9LrIyCad7R+eI4EQ8G5RHrWxgrHR91QYZcedgwd7zHKw28R6e3386glvE/8FLtq9h6Fj
RsdfW6pJfwCWKuaM+FxoG3hK/XCWY3+4hAI6S0Ejti8QPJgq0YTbIpABTAT/OcYmmjBt9naDOExs
fzZib6jucOE5tw5VejSvbQMITk3j/i4hQD6xhora2539piKt9874T12kU0MBwTQjCNFTEYJKNElJ
sOkWaAWjLSoK7CdJng5v43hl126kaNhvJLqJ0TIHThNHcdD7VTNM7thxf7reKdvXIBH6Ict8pkvd
bmxkLIw5ARE51L8HTETIBrJQldsbTNqzb9lHwp7bDJLmbZKoJI011ixjaJmkOjYW1Rw2UZDiRSn2
CX/hr6nksQUCm8gCEIKMMJEiDVCQHKtJcmY/6tESfkt3EFRMil1Z0lSskXJNLgqa5SRfBA7b0HqS
0fPbwFEdSMJNFv7OGjVKaoRtOBPJfnmngFGNIA/1Li8kkZy9xY82Mt1ulw+ou0wqsvZ3sgGlf748
sXOf1dE6E9ErloyujDVTtzO8nTrfBoktrBtZp+2y7inlXWQK6RTex/pccRugvevr1s7BjX7DV1Ps
QWjgl/Y33/DP9nOCxSZqG+c8w2uWc+KuFOrab1rWT+rmqg6fGGCsuuZggM3Guf2HIfZzpWyY883d
Dnrz7UnUeOCBfkhl4+YFLAWWYc3eJZRnuMQMKEdQuCdc/WwsvM4LJBWNeakfO1lmzc0N331ppZQF
Yov6BJjzgKMRoHPMjb1Vm1DTCr7iMzfFSa+KP+fg8r6Lly2idSNfh3icG9TBRErKCliWFnN/Kd6r
6mLEi9KgxFYFfuDK56ifmMuE9OT22j9DFbenN9gN6bsZ3h1GmE1oeCuc3AexI3BbLsF4JIIKQrGI
3FckYAzJjNeatryT+ETWV4JH3mDOorh6s0tLPBpq/AsHqVI8f1Ri+imMev8wA+sBvzOg9n22EA+l
b5OvY5P5CyUPyY1+MBoJ21CGjLyZJjfEQnApXOyyAdxl9MmPeDIxc+aVrwtsTAo02LsXKJFBNZS6
qxGBdgiZeqTKcCH5zNog2RwC2yi7BVI7EiLBhfzT7BQl6UaikWpYc7xDEqrwIW39y4n2eYWZNZqy
+OMS4UT/qvfgCxK7DYyulvHHQ5Z8jFuIib3K8SphPMZuix6rZNhXpynzbxPVdOKHwASgXZ+bR6ol
RM6sAJ21gruea8cPDCkCRzVN+4ZKipFl5Ra6mCj4CqCKj8K8ZnDGo3cfdOxoBPYZE0rZwiR4mh6G
6r0a4Zxcs+KW3YKnBM2T0LjzTGXjYP3Oul0jXvAM3bnmphvqcqTT4ucWjH5eMFZZrGtlh5tvpzXU
0lCPRsN2qIlEI4d7mQAYHLboaDsUgiO5Bo/ZvD0Q9mNVFEEcJ7iatsXL87+GI8VrnT5g3rO9x/ky
HoRUUUq4TH8atOSTQmfYipG2L6halICI3dYXM+tKZuer78nuAv6e58es4N0mq6f3uy0HHR8yyG1n
f6d8YVh9CYupsVNDoA7BmLs0NIREfObiELZ5r5c3zwOWlUxJPrY1U3JdlCyJkzdMiBecREecB3lf
qGWiEOTq+dPDMiyjyiKgn2hlJ1cDXbvgCYaaK9s4zVbJm8JbJZ+JNnKTNiUNOCDn+hF4k/d+O90d
6MBIxvYk2OU19hn8iLRSQwaW5WUqJGzGY6efW4dIYWCDm3p1RxwtUySPbUMCVSWzBLV6TndxcsyK
FpyG6QIA8cwHRx8g74effVA2cpPwzpURcfXo2fbAq0tdZOj7uQqXrVh89NWRMsvC+MN0JJ5niFxE
6MCtXul9GSMdcPI83PDdoc9AqBaGDvWgKNFTG18POVTCtplQqr0wDCvVyKR/7Ksomi56Ki0xAe1c
ju7tm8c3dbpjpoBG9zVvcMaCeeOjbk/UceujhM29dnrw249F/Kzbipg15EpbxBqe44e+JR3Eq7+t
XE4bK9jqfww09y/Ei9eV+akvrtmOPIhM25DULBGgc5AphbsJSEUWKGWb/oV8VkRztvFHi7MvWXf5
sA9mCuzWeMHeJm0/zaNNLb0anJj+0fDWunJt8hMbHEyPnqnVeXbkN5UZSNoCDVqQO6Q2E5m4CUIP
zHqITyNJt5YheezO/FNQo7g54sXJyqtEMvxrno7WaNiOZ4+dtwsDbhjDU9INesPpBUVBt12oUjbF
JxPX3faNvC53w6d/t9md2ZikRpvYd3zj0UgJvTdCJNU2nkqmqCO6SbRHAMmyWFmsj8YdPF4pvUsE
eqWjQ4du1DBXTpqUUEsVWeAzd/RMn8COqyz+bjVw8nI5RM6nBpS2uP5pTzIhafqQszPNZ99UDpdf
hte/LhaR1aQQJnEvqOKe1gRnepcA+Kp9ixz5TOPHLFqLFfoeLKT4qrXnwhMy4u5X1ru3UC1bpNoz
Zgkc18kIEQzP/i8wyjjyn5+qDVqXLfOCVayU7na8Ajz5v+40ZLFdA/sUVcvZ7Nlkd8rIxC6Bchp6
65i6Wd/7NnJWp2XrB4p8bPaRpnl2u1lqRv07ZlHxVobAiAYtMkkjH+fULxr6hL6Wu27ZBJeTRSr3
jA5Cx5CURvqscYkCHIHJPLEmpFlcgME3+jCiU8qsbAyIlpZsK2ADnIsyyBqE742kUQbi9mxRQ4Cm
t0ASm9iQPm+XNsXrXNebbbnmm9cLuDDYY0Sm3bo0TRFrJt98350uxK1tdhd13Qnh1uNn+HLdkcg3
2mgNlhMmr5yHXCJv1gcYc7dTlS348f8DDJchhJJLz8cGVroKGL/ibj4cL6BgvT8spn7DCH6D6rCf
uEaknPLltxZ0uqZVATdS/EgdUFuZgHkLBwEAzvwj79dLT8r2j0YVdMOAx/xqln4+mFD8GDpFAReo
ijioPsSLJJpV8qXfVkQOLMdxt+BvaxgeMdMxwaQrRKruKcOwk3dn45hkNEW4Z03/hA2uu3SC6WbS
6/x9E9dyRMQyWIkw79LYURFHFe3Bs6pN5qrUMoe+UFU9aSqkiyuRkTmxQ9FPrKZPF93dOdO8oofb
1NmL4lDwxPtTj+L7ezWTbHUangAq93RNiiZEFA1Dko/MiVFYR5LK292OEPbFkTdE0akGy1sz8pEe
u/p60FGziRwKf1BlES4wQFjTzVgZmTxuuXnyODF6f23rzq49C+DofNZzHFaN3+9C/JHl66mjKHCO
fZ4I9oSnmuIoCjIyE3U26363nyUHtSWCcRJHlZa8f3e8JU0r+ZZ8Dl4QOPSKDvW9zI93CVT4/FzA
53o99QnjVraKtyDQx3dB57B+fmbrtIfXpA4sUm+jx9UYMr1xtp7Wok8wZd1uAsO7mj4WeuFNGsFw
USMgnF35STz24AZfZa9yrbMRGRpevtDUyruWfpUU8sMyAO8QtaRLuzHDNKGAc/dPUHr6boLhGmwS
oBujM6qtg12fJowWDICPin8mXcKU0jHFURuRDsSFCyacNAilGLynt6N7+8ndB/DtiAdZyct5vszq
jM6OWVVloDfs/ILilrIY45GDc9PU1s4OWwS68AbZwMqwXWv8r4FpuUEx1/YK7P2WlRDwperhRbwC
dQEPxGMLZ38YlCFseK/lvdaeGjzxa4yd58ranoTx1CfGDgkmQtSgmqTrXLKNJKkacUZhz6wzQuMb
HP8Tur7gKatR+ihCwgzu0zuYgyep40NxbF1HDGUfxhfjh99oT6dWrxEg5+NCekqAK1WDLz8ZqiHI
yNY3TMRvxWLaT0Bs7k2F6xjfn+qZa+B5aSNFHp6XhHbjgUB/Nt+v6XgeS83FgdZ0GqvseT7OTdxi
82Q5/xGbXywEfEUVOJbMcY4gv7/jKdktxF6/Sf4creQFMLnwP1H84irqvP2B3zHrI23EWlilVxue
NqpDAw7WBgjrm3Df0e1laFYYSJ3eQGR1xJmQ3Npp/zno4L92invF4e+2iYT9HFoyjJ8Kldd6fgU4
wkRLx98r4klYUdVUutGUBF5RcPfAt9W8axFkSzNKgSq/1mp+bqHME4BzhyIUMHzSVB2FhvxUNerZ
N+1BMohkqGGfNmekdF/TvGZQTZvAGEDrA17yBl9n4AApwc41Mbmq+TCs0j5SSfVIJKm16noZOrdp
DtTm+32ddntrpOws0BZHS8Iwqj/agYT+DPxS3J5umJOR00RkQksRdexdGRgg56SzE+4Pxirctnwh
ceRXsRvNkMMquQBxoxA+7HxyVEGXSWkRgsl9+WvI6aVMGosN5UruPONzuwvePrW2QMIJt7K7FePf
LudPx/10wBoT60I1t822I0IjIUoCw7cpMWlkk/yOfCOAcSvgmSqdag3tg/1UUnNKHmmXKj15zmSs
OUDbleQ2yg17Qixz5vv5yu++4hODfGPBPXHXaCHO+WuGGwUlerelF0nXdQaMG2OWeMkbFoCydLdC
fCzWQsDKZU5oz+Iu7CaV2qv3XF5QDQg2noAzyhXc3KFNQ5farr3wqnDz9oAFAMA3PMm7QGTCDybf
AgYp4R1CjCdpjTaW9Z+14+keDFXRCQxQYmYj+WfRG1cQ9+Q1WkOA7H0P3Y5WzpT37cM+Jf0nYxgT
32DO17slzWhg2Znb4AeBzJT89wCjPKjbpaY49YbYrPUTmTBPzIkcZgtDrgEHnKQ6qNHBrqxF40Ya
q3b/Q2XO+8nMtkyTKSsdhDhSghy9VgMzZZBb+RFSrCYqL7tYWgrcKOh47F1kFWoyb5/zUImhhP9y
1ewbeDy8v7VcpWlSMF81zB6tRqQv0kEVYENQDQ+O3vyiZLypdgCP9KmnF86qFXkwEIOQXqR+oVpT
fplfg5WGaInDoLJe5UiFQYJzelH1EXY+iD3XB/14mvFexi0VkNn0zfXrd2vlNFay0glT+9ngg6+z
LZoQr+Ha2U/jnz4JjZbTiX3YpfXNTwYFoH/MzBuyxdsvdRivA6itfpaPp7vFT/Fdwmop32vlQ1NH
yBGOstxp0rfzdlbC31SZiSOTgibOehdECFcg7vPgTv0N1CGSyhaVla+mzsU/uRuNg+WPQ6ORDISK
hlxanA+E65/mmjO2pSq+rAIt0NXSSt6A113N9Xd/v+cpeLBfED1iZ/PAA3IeWmVymfoEqj6YjKH2
cRcxetUgAohiXoTiI8xs78M9t7urOUyI2x+mjMhgBvvWRMXVz2Mi6JrbGUUAyg3HcAk28H/KsVyL
RF9F5zj2KLEtqL/41Hk3FMlnMkbC0wwwlBH8YO1XbRrDUvJPUGAQTAiM9J41b7AWYhbK7Rr8gMUn
bloc7PV291ELF08nEGTEaK4ZuQpC+rGKBopbkU3UUi4ZpPOAgW3Ry5V70CQ0avaR7+wBD1e79Xmg
1mangmYly2zAL0eh1Z2FuTSGhYs0pe35LKSFzqEB8KL+MxgvLMCu+K8nfiCj8TssNHSDlEhEDiKQ
VxsqAuW9ixAQ5VnFevhWTot5eDg2LLIL0wKhL7EuoHZRibv8GGBPSPtwbCwDeTC6ke31yy6pbRIx
u4MEuXIdiz1o9MWrqMyQIblydv8kkdRFBnAaWLnal6bn+66HOnmzhpX/JgOnNPVUlYAct5wqm/lG
TKiMRYbIeuCUFjIflHXAT05A1S+9PkY1XQx92ujt4RKE1JB4946FAY1QpjFamrZVBRG0qF8N4J02
sAORmixeiiDZtvAC+h85vexEJUEkXhyU2FRoG0HWJ6ZWjUkgyyn6S6HIVvbgdhoB9p07mjQcnfLC
ZYXifG+Wy2WAW6aFeb1uLkqzmoRxKbQazdy+Q0W20aUY7zmS+D3euC0sPaUqKTw6Awu4pmnRGCfn
1nvHx3udVMGVt3OZCgNj+ta2Qo3hPgy/ApM3qYHDGMyHb/dDEqv3BWFudG0/9/h+/GBTGHgtOsp7
Wksl0OGp/mnUEoMaVk+rAMGdy/YFRYn5PbeIwmth+VihKNQIW8pXmJ7MeWabKpsboufaIK/FOxgX
4HQTrKXyqenXJjavtfXObZaTfAjKzh4yJQuExdh9wMVR3seNSl+U2KrnUIXTOoYK2MYrg+8ljNvG
KMnsJVS9SYV18XsEPy/T+i/XFoHAQVWH84vufyuvV9WcSqcb0LDMixFrV6EBfaBB1AJda6k23OfS
dufO7nuwSG23+NwSBGidI4jDjqTo36lp35ca5Fd0ANH87m87uR2su+A6bbV5VSCyOGaFMgaDosRa
F2IaKjEBYvBKOZDxIRSGAk91iTOg4J9EzK6AxOsd9xu6m/YYykcXyeeSjsQ9kJCIc/pTKeLjlkFI
21HmlYQZg1pGRHi1y+bq4XYNGZe3Lq1cGB9dBiShYs3NYKPfbMDtyIpjDap91F0NZetd3QmImJWC
h5OLDeJ1ZLUOEgR39+E7wWq95SSFtD1INYZ6+UUfIrciUdCKCrJtEZStgsWiRnzEnGM2vT4XeGAW
bycx7CANLKtn719/eCSsAwEsGHcXsHZd07aMI+cXH6XIsnuNbhz+SVKOiV6UPE/uerGBv95M3R8u
jSxD0Z/6zOGnE+N2JtIQFZy4gJQ1H8z7JCJR06Rpt+Ze4KhV7pQJjjoAXGu2apGvhEbdBwxlnrx2
ngGz/Fs+wYuBpGVyP8PlLPRhSubA+GsDPTGXM5Q8I5Vw3OPyJGydWkHkL1TPcPIRvg+CoGCKw92A
HbF5y8Fy+KqG+6c2QcYLN/n0CUQp3xPjov6kBk+NpqLdlJddLux9cfx2bwb7do0WW03BEVC8bT5l
XwE/yu/uDSqQjIlx51OU8PjF3J9MoHtqHGM2Cjp7KqTPKfbPNA8MlwCxTNEdL8IvkT2IPQ6b4QNp
0D9KDMMfSIOmuSF+8G0BMy6inbsNhG7EVVu6xy215TnVL+3ZnAOzQP2nZ94dgz7CxLFdep47TFw9
rM2fbtQzqmIzhtX72QZkQS7wuR0NO8lsbPoiv3oPprQ2oqFDju1LIc+P6YmyngxT0Fzv8V0ITbqp
DsAipUG4hjA/Ozwaj0AjehkwXB3oeVmRE/ZP7bUGedFXtwlNYSGH85QiJn0MbNjtx+gY8XbBL68o
8ZlXfeTzpzzC4P+hOwd++C5IswSnv3XlRFPzU/QfK0oB09WCZekm5EYz2TRMvdBrHqgg/jQdPfgv
ZoxRBCt9BSMytFPmAgqt0j5RZH+FXFaip8P3REZwHOxWljjVa8bjmT5cbcvMU1lha+yIM4HLG3QP
SCSX1bc1MevaKdS5aZdvvmy/LHb2fdtQhjh0kkwpbiLw7J726Jo1MARog1MkyLsqL/ryDCA/fluj
TBDRVZko3wQ1GfMdhBpmXD3oN8/0In8tiQCLd3QY1Mzr05/7037rXlp4omuWg/n7RJX5gzLVoc6I
+Zg23ssen5MSLjaq+Ku7RF6qw+UdQBI+LVpnl56yP4+EkGLxMZLh+twDgAIxPO7Q+XHo+1NcABxa
CW2snbgb9y6JHwunDI2nf3yOvqmL5pv9DTaX09zXIxqnXVIwgYoxO5Vwn6zcYU3YWB96qjpTFGUC
QDUHc7YtU1FTLyqDgI3myfbVxZzce1oTLAv6r6Oxv0+aJltYrzo8NSMjqRdjuUDnG7dr4qn/i88s
htQYPlf/U2BApekWT2VOvErTmYoD0e5X4YvpFZqGytU7KpZQ5FlFuH93bNoPwEDAP1YeGEaUBhcw
nKO6U+ms9mguq8fMT8lAKd3Rx7G5UPghLBan6iaJM9TUKAwUbt2CTY3C+IULM6Q8xLMaRmXSxP3P
020tcRFcgWiz3XKohCPhoYlCpkEy08xYWR2Ww3SbfQ49pu8SsC7qUqdaAnh2oY8gHE0C0EKmCMmA
TrNoZIuQUq/sNdfFh3wCxTVnhG1WdM43Bfv/oI5YcUENO38a/8r+HcPwF7pJHR4V8I25PoK4cTrr
MYvMVmXMwJDGuYz/d8UqURF23ekXr8H03O2Iv9ulg6vMLUMEZaKADh/PSWW06t15IlEznzuJbEZe
wa9t7O2xbmiFos4rugZWh/LMbO04P6qhxG6hg1vzuK1TkCivenFiAF6SS+WAFz6d5gcx0+lpkdP+
KNgez5qAwNs0xdv/rhMWoOcsc264XuRj1J4VgeT4sLk1rxMgra3LQaHgBmXQ0cwg1e+mydPzNvyU
TxWg1FGhEnadBO79nUnMFaIG5Y1FXkLsaOKawJjNfjqOF+cMRSPo5Or4K31WIdew0798jX5J5TN0
58Ek/QqmTd6iP/t7SpHQKJ8P3ANNrN55m9byuoVTHsZMQQigEPghsyEgugVrvhaHetQ/h8nDO6KV
flOC2RV36R+mux44IMB7T81w6TiaWstEUVglb7/s7t3A4uo0/QAxATE4Wllnab9Wkpi0PTZNZGlv
k0YdrG6H2swO/luhYjMmL3Mpl1lUc+sLgBB4FXVAHAd2x8unzTh87VxvIWrLxhSjL/t3Ep/Ny7oI
dqXH/P3GNOK5FzyBpphL7V1Rg23eUloFqxeZFXUHtmTdTEDfpuks1SdHaztKsEhp2kGPIkVltI+m
SZBLxnjxf8jXmBMRV0pir3/OCxx4tb/wENMgwlY3U9JhUuHk9kwyMM/a3MhmOl4TpxQJzbyif/2I
N/JgW7SMhYpc5gPRBQ3btfh55r4YxbFyqW18gTbs167OOVRt/IwPAKDYFi4iwvB6rxgjvT4IHEMk
aU0L3Lfs7TpVIINC743z8wuBn7sRmPO4TgwoidsbGs3t2+WBsNLbJU9nqcOeX6m+JPectvqnR7oE
VXTXFr3UsrlfygaE1nDmosQfWzaKJpoS2vfauVtrzrMzrQSD6R5W/pHMRQSRN0PZcG8CY/LxjrsO
SAJcwnPrONBCozTC9u0OJEBGikqFd8CunLHz54FqMoRvmZQhsBDPoiu2w79ep8i8UN0axfOliFYw
Ds54rdqp1SVsb9AG95xLBCmtArcFWpOgjXb2Ws0eH2bPg1wFWuK9wR1QZgl1LNGuAoPNgXbxAsYx
CFyjPhTA3yFndBZ6WvPYhzyd845wYDcFwFOuUh6r92tsM8FJL7ry+i9idmRmDVNhJBTwkEbV2t5M
8H9WlOFNeydG2FGAvPzXCHZKhxZCr4t79hxqlCQuFQ1tm7bsa+IFdkz6dcWqcANi2IUjK81f+eY6
sSJZ1qzmLbgNG1Db7r9SuLYt7jo9C2joAuepaYRJoH7faq29CAKn7u2mLQO45j5tBH+/kTI+8/XL
n7vf7Oguc/rxPL/XmFs+XZB4CSsLqOUXAJSVta8qCdHyPMzNCo/2potsfU9JhnwrTVFcqylggwy/
fC9+hAn9dGHF+h8Z8PmKbAQ+2fWiSdlvwbWM088hKTDzDTgcx6wrv3nLtUVxliK72bkgQVon+HzL
cDpWCbNhvOUWGkgfOnW1EACiGumtRQ6m+ot1T+oACVTbaRJUAwuy4XuW3oBsuDtCqna16lJXodeK
vsdh9dv4wsOwd68SeMBv8Y4BWO3j6Fy5lpYUdBR2QBPvn7S+iK+1I+fh2Y0PdqhOu1hh3q1s6Bhk
cz+Ul4zfc6k2dmHrYCbsV+KVq4hw2YcotQKSn7NrwbGhhBPFLQqU8F3pWe9pKQsgaOXPXEbsnBws
nMhYIM1Mf2ox1JEXITXr9xetpIHvJp2PWx/+wJ7JpC05Hj4L4SwY25Uz4uNCAqsK/Y8AX+sPMAYy
vbhlRlbz+f/Zoa6ByLJKdT8n65V4kyaZHRkyPxXuRuW+HGebELTy6C7ac6llqO/sWKrbtPpysZor
4PcRTXFPPj8phzoPhzDeCxtiItr6rpYd1cmdNpdQIIinXrCCRp/cEi1CGu0R02Me6SVnGUGT/+zK
yFni2mLg3nAn9hyfJAaDUh2CNoL0MnMyK79/Myr8POPAuhNSCOxLAHU9W+L/2Z7nMSQ4VtLg4Ca1
rLxtiCREBtlaNj583Agt1l2RmkqLnHhQKSrph0Pfcl9pzA4DecvEtI4qwYQ7UiwB2OL+WUzM9NA5
7xtJwYRxlyAnYZ9ki+ebxi3IXUMJ9/UvOYYLVv9wPN+fE37k0kwOO8QQrvTxJux5CQMfMwvosCRd
F1gcegO7JSTRdm3yhr+1tIOcG+R7O7QZE5Khxwyz6eqGYu7860pFt7WlHcae7J90kq3jNp2EhRGo
s6bIVIAZsg0mkwt2zm4rKPxi1wbHVEzKQ9FcC8mHNdTlb06eIIoRnSzgq/yWaspnyoL/RLTvzqW8
iMjbFxhQuyJwWzXTA+SYkUWBqANJtfi6ILl1tLid36ZDhA7vc9ivaQ+/zekZuEQ/nK/TA2wVApiq
UY/cEz1IXOLKSrDTcAk8ieKP5CzXOfiM+9JkyiGgHxZCzVWQlRMAMYtRzWlQG8wsgzTc0wwUHXcY
0HNggjXQDbW0atEaJ0Rj4bBmRcxbVFEXNtxxhi7IsjnXHxG0o2RRdJvkNLvH+RuEafva95F8gdxU
yvmA/7KujF3ocFxKac62lviexvZ66cZ96L9klyDV5mVQ8iYgphqBwsHGEzqsQIx8QoJi6ZWH7STl
HxkxUMHPwJDwKXG0WTQmaPrS8lihVDXHSYidS3QKMafhwC9uVYeXU/Uc8h3+f/1Xbxnc7jDb1Hem
IkubKZ7vtHFh4xPGpq6i8CyQ1fQBzLtqm9gV5RvtorXMV7vvbehZT3uv6zpgud6r6rRf2izS3Q7D
epd7cyQAIhkvgkpXrNexK03Zq+17NztGg52R+WNQB/fRm8xjk06JOC2NyM1RFXqQQv9fVlQkiDaQ
yd6y5m6r1/MqocCS+4cYTjMqazjXhvCmIfIX3bHgfB17K8TQjGE8jmDXdIJFJauNBbIYKlCHAX5j
cRURk+UE0bZ+XYjt3q2c2hVZNNHS0Yf8nxMpLY4ljhZ6ikLWjzsPP5D8F39+3UyJD7jxl2Er6/xN
9TWTx70UrnEmklR+2dAPOqEvKzRCbeeURd2X7hUcjXSLbJN/MpxGA1dI4jlcEbfcpyPOpaUUlOAz
q/1aiouwJLZpfDeWUUxEk+cMg/q+w62dBo3y99+9psbDCdAE4vlh7nhsj/Q449BPcEGFFSnstYwo
DDft3bVMeFJNjDOpxVfLU/CraN9lEWt8iNhP/eccPQ8naZqMI9bD0me9Od8zkLA77bzy6iKA+bey
zf/bIwC0siD30UNvzvP5BrY8Yaml3Zz3MyAaJiicFbgtRsQTOLpPACsMhSht8B+q5NnGEQdWIvEJ
mTNT+XEFMiiGILEW4YovZm7iGlkNagm7SxTTs1mWK8AxptuRVEOFXZm8njQ9YFdz3FCQDPOHZZO/
ef3B1eg3zbvxTXtplRdOGC8oycWxZUsLdi3MCeLKCvxtp8j8FDqE2Q8GkZ3y/td5dbCbPlLKNfqM
LDXdN5EBxVR3wPnyvCuOcWl7V91xG8TfsHydFLslonujuYdpCaSHtHu21LUVHv6vae/aLATyH6an
cur32EsbNegHXNNWh5Pd95EgSt82wO9IeCBJ7IFt4NkYGwwKStoCgR9zDqE8Q5iZwPIm8PmrG1Ul
nZCo3fu3Vl+rmpmm1HtS97A6STgzhSdklzbh2b+KZwu24iq/ibtc5fc+xmpsYHP5xoVZTzAzfWAX
r9UMjc16fqKVcTZRHJQR9wLWvp5hUs08DNLLewsFsDRF+T4cof9mZES7elC1NhTu3IUNAF/7+R/b
sm5MHz/Z0dg2d+d5/FMpxOH/i4b2oQa88UAZUaPBSL9sYbe68bfoYCXNQUKcYo6XptG29u6gPyud
w8/3uS+/zqTWFyk3HCzyTs8mnhsPmvWRY76V36O/K0Bv51WtVx91cs3aFx0sPZvFFWHMeDsm1RQZ
qVtmJlegLZK29VAI3Fp2s6jXDlsiOCbkwpCPnUh58xvcKbOgHvifpCwzslzl6e7GnWh06OP9QXjK
pV9nUY8Mclbx2tNRg6X0ZVOCqQKN+z8F8Fs6Bj/2A3b7Nk/vnqtIs2hFM9CoP3vmujSl7S/sMXDF
ffNnWCqTqwwywLp9aHaMI2xkEhM3Nci4i2pBAf7+jptQmp5HIBzfJyrJe2tkKemiBulhaixtDDZl
toJdmxu2Znl27o2B0glyeU/lrwfO4njJ9hXvKq/2/f7l8O4LQX2C9cT2Ocj2ttvvJeNrFm49kFV9
zV5kQXiZo7K/uvz/O2i4+OK2U9vRpn6gZ/eoEilzRL6zgDQ85hxUQo4YQDlvM34uV1gg9U6/nDNm
IcGHGbv0sSLV8xV4/nk9oJkRq13TEDfdc8FT5ZBASEJdRTfZA8lO7re2EkrBI6DZMw+ba9EHXWjG
luAVpb9uO/kfFGz3oMBGY1waJTNv/pCxppdynnJ67SjEj8fE+Sa1TDgczOqyGRN++W98mUsbl9+H
TTVJOKjwgWfWW1gfyQhHwNhUbTwKLyd5k+9XBg4sIUNtLEU5yu950NcXrvoO95sjwfZWqJ3Yif98
yfHDvOL2jqzhs5IkOKg3hLA6iMKYB3BCknpyGbMn2eN8wCw43V27ibBh4v410HuxfcTQGXZk/lq3
ZpErzgsPA6cVGX6QhgFo9GpA+LN7BXYLq4JE0CGQ2WZGLDjV6521FtwBquY2iVYtaeBeEwNRjVnf
VoHTGEpEdg6LaM4dbQSbBZNPqlVkbt/rX2tN4+Wt2In5EJkWbHb7dLVBiAj66lSGU+RKunh9y8aN
bi7AmRcYtObQz0VsOqT42aw+DCbAzV/GryT+Tzz0mX/1G+igVyQrDa+3ttWOdXxcfzu4ioyUL0Hc
zMWQFbpgwj7u9YD2cOekt0fGl1Wgo9IaHuwT645hovhcfWsfVRq3piK1RYFvDsvK4q1GkEaJp8nH
zlgqk8pywn22HtVxr7BXGzo5wt08JMY9Zm9g8X3f86tT/mONcIASN+ZSmcbNgJNd8LuxgqbTfLJ7
JdPSGGDvMF4J8wYI621xn/h0VjR9/EJcCjn+5lNejkKKPn8cpE+p7flwdCdTZClrlLqE6bUEzUtT
wXDWffv0w6N33dj96pTckY6FAa8s2IKXKkwPJR0jdx9+PIUFDmDyZAKfAaB4akSF6QL8V2dPlFPZ
DsCouKJ8IZIcb9g1z+VotXtVezLedCZRqJPrY6HXXMZCN0/0+ocy4QgguDX0G5T2aghWRHZfLUfr
GR9f9zK0p7qdh1ycIvN5rwKxLM2p04I6p5VUUT6+8PymE4WGb3ywwpdgtrpium+rDSVW4dxtAzs+
fbAT5G/ZWHjbow8M19xOx4eB7WjkBx0gvgHAdWwKuS+6HqbmYAeopWBoCiPLG+rHyr1UYbYKnupG
Lifa1Xpi6RtumnEnkMhJBYP76G3OaUfnJNT3iuFymwV+fb1Eb3s4GrFhQGbLHg18kB42FO8Y2YZi
cSxMtZMQks2rhYwccWYZyQ2AfLLXXvGzgTvvRZarePWZB8X8WJjlS1zAL/Bms4B3gn+GN1p439qW
7tICaA3QPp5kYWEeWfKBujzGNqsqyFJDqL93DqeZrIWjf48A/P9IgXdGoCfvJXaVGj3B9MmXep9o
Kh8ESsHo2S8rCOU5593p6l7ow3JpczFcaRknxiv+fdqnOel3hLSmumnsHPVtAriVWmb/+Fpp1fbf
yqVYYRuM6kABXYk8TAw+olvMASh8/05rLczGMG/viwdPPU6tPzf55KjJlDmezMkW48rInBdJce2E
X7V87+U+s/aGHREmilb6GxvxVBZdhGyUcaSTHy61p9UCvfN/boWAcgSM2XYMhy9JrGlPAJo4yYCl
ANMQQrdWfxfCbC27Mq/EYX5+7lRiEJq9QJSSG3kcNvze4ibPunMvHYc7wCefBBfLJJHFnYhp1KzJ
rvBDgTV4zsfDAQwcQ2Qe6bmyr0bhV/bLrfXoom9nXSglxNM3qoRAm/c2mlWflMpWVRWhsG667OqT
ZaxwFq9x1Oaa/5iTm3yVc/BoIWakirfLzsxypBQ+HUv3QsH3kdplfyMZxqYwji2ZDvfGIc5WFxDR
KNgpO/oY4yueuZKN93WI6HbCb8Z7j0zoTzrXQ1zAMzQhjGw42AHNBM0sAvYBn14vCzithUhMFtmA
9rWMMR+z5O5sPalzzv6WyjQB8vNUuet5kLk4qsC7YZUOjS/IBPkBM0syTkpEMJkLjur2UrSqPMPI
XMVoonhdDV820qRUZIslSi+Z+RCN8SWip1CrMKwR9rI8+0towA94UQoauoQLX3S2TgARrC33q9ey
tryhwxc/wW7A1wcMFfZXtnsZzOv78q39HpgICJk+9T7bNHwoXXr8xwyGV5oRi23v80SbDZFI1UB4
iK2KqKyQ1II12lSPgMEb7cRr/n/GSnOpfay1M0yr/wiMV2YHP9v3sakYeU+JYCy5MTCGsgDwk6lx
KfMhRrnRMM5qQxnXomeA0sKwGBQV7R+5uQh2QjHkvXtCmjW3ogWxRYi9t8rxUT9h55bo2h5+JZAk
hyczUwymyxF835iLm7k15KydWgRrXH6AN5xLF29lRiq2cuRUb4DwSFPuyM+JclQsKkMjJTSeTyaK
GfaSZ0zETkRCmahhDLyPbmMf5YRK8qUESdMlG/5cC+OVmPDDr+DS3BfC8SlpR0YmNdvrS7m9IJLk
C9dLIdOkWTiDn5vgQhX5DgMUMNmz6lcCPjPNYI7ro9Eg6kva2CpvtwppfzQeXYUse1UTvXFtWwPT
MS7dc+APO4aEFkRb/0lCNnJk6aLg1lnBjYDlncEZ0VG368jccsQx0UAf6VaJhJ/pAqaDYWxGx3Co
S4wxCSapQFR7p3ocIdw2yjL/g+5ZWCO+qYQP/8o//zDKT6SVlp5oH5Bt95uW/bpV9pp8gg227wKi
5JrtIAGrEFBl8G6iejLUpD0SRS+mj4l6gCXOftHlTtmkrP3nDRcGNtDn4BcK6ptyLtEwiXdZDXvK
MFXdASWcdn32BhQO4dv+MEjLWuaWyHOIOMJp12FDVtffpfGkju99ScwpASH9uJYRxUJwuuMQ24vZ
0ucAzyanVXjC1dIx1AcVv5C8Btfnqlc7QL0cgnvjBplT2OXIQ3VCKStIf6mrZgtvmzEN9SWv4UhH
2VpkvAdpHObvRM4AbOOZNr01XT7q6judP+AVLdE6zLCwXPQr7ZfznMZ73m/1pP5pMZJ/U63JFkzh
/cTvZcvrvG0ad4DqGBNJDnFp0VJqGS0vBKLESIjtOvU//OhLP+FEyuZMnuOz6gCPIVn/3n3/hNF1
rhRUsMRfEc/ULqMVONoNCJpoEaW8xxJ8ehGYCbNlF7ip6i5jgarZVw/uyHkZi6shi3gbehUPEmyN
rfYfX4HDHynmCp72vPKoSKo6WaniBgq/NgBIOUE2Gd+/dRTznN0NK84EzvfM7Zrw1ACBPGB/YbT+
RBbMbinuKhnrGlj7Cl3mzFBvVEei447FWrBVvFGa5+E8UTDuBVr8TFq84ep0uaN+3FKbHTqLKAD9
MsK7XVfAFbgNB/dGDi2uZVjIWFt9yx+bEzmAB053vlYjRf9CZ1+DCFRgyRqwsDOHv/iY/Ab09ILF
av255MWA9jI56dNVQ83TqAzhysTZEjyfcQMg6b+iQNXEBPZE+tz5IaWJ8n31lZQzzBw54/cEHVCU
HTF6LiffRcdx6XhWVJuxqGxR6xAkyNVh9fd1tbAQ4HzfzTuIQ+7OWIA+N0B0LzKMCq+H7cShdmD9
D/+MMsyuq/Lzr5/Rfoz2b8Wn5cQP40/2vNvsWUjqBXJFpjj0WaURX636fGpmrlfqWLW46Q53F70J
hFiDNJkLaqZL1fROYIM3drB+HgkyP9Oe1jvsOYgeIGT42wUPgqyYompOKHlY7KyG9XE9lySXtnP3
isNQzZl+EB1MKEw8oTx9OZyYsgWyCkN2A9amkmChq0AR2qnWhkemNHdQI8SUtm+iiHkhAvmdfda0
DXbkqPpdLBsM9LuSQfZsXgzvl3NeugoYezXc2T+thgcXcOl655GZcFukjg6IWmskacLNcJzBOZKY
d5dUxgNFreb6CZLqX7eAcNYsQCxGcWcxOide490XRQVlNqvVB8r3WL2nXuKVUuBCQ0B61bqEZGLK
6rW+1YpLoX8R3tnvh8LIYT+0Zg5rOIxYK5065xG/lG6FJnHmowCHLSrkClE67GewmRIUfDcU8tPg
OV88oneEgWzD7VNybn+i/l612UJ99d7gK6WuH3Y4dighrTN/LRnSR0TBXw4wns1knMRcqU7uxeFm
yXhHk+ZxWUiA/HJJpT77ccrgs48jYb8hNwuP9u0/G9vg7/qj8H5SDpsu6Q/C/i+Nq5jszFsHdWjY
IBYOlVOZyyeAlN3lkmTb/oa9AZxqwtsVYxLZXwnI1X+s7yXdOTirWkFAdgpFV4piajmvdUSj0Sx8
zN3ajYeMrKayx4dDtzDsO+hq7fgJNXUxMuHP8/K2TuoPnnY0ZoSWvP3h2RCvhjoVUuRTUS6GDnvj
jh2AYVQ5DCM5PL/gBfxTlU4P43jtxQBOs//VMoTtDatCE2rQTvxvlbYB2D3BsGOccqTQaZ2YjQ2N
BXnw3dAcc8PUteeKjqB1R/lIKks898lLINpcCyfgyHW2wqmdK/bWQSRvZQxz/cqyfFjtRDc806bL
898AvEgImWbSYnwl/I19vPbpXKDnlQKF+gPmzROTtjjLIlRvSeYDJGzE4Dv1ny75JOpc3FDQYY0g
uBSOMnWyDUJq4yMxhxS34W4mbzE54+9zmMCa9XaYYt1yty6SWGKZzMc/WKfeW93TfyXiUfNVyTO0
Vw2uu8jsci7ZdToN5dbgI8eaeEYl8MeQ10jGdSaRpX/1hj0AU6nIE5HhM8qIJAq0Lp9AFblw5gRN
IDkFZcveqlqGtxgfA8sEFhM/5FGR+j28VZ0EfqBZfb+SwQkJ8V+bwyaS5it0Ep817oL8yiWziW+y
s8kfsdrU8MGKY4CsCIS2Cu8nTOkIiaCBTKoQ+K4fuISnJynDZgMTbbxoj5Z71o96tUi/gCR2PpIw
dOMkKp+zXSWFfx0K9He8VOeC6A1uYlb/dhSJvHU9KGyj4h0OF/BrNZj0kMEHaDCpkIK+YvgExm2g
7uYE3Q8O8M/hFA/RTz1EPh2H/f275Dk8dteiV9e8Kbgew2heo5eXipKExTwh+7+yF3lqiBNHVeJ1
N6y3cQtA9R1Y6kEhDDRzywKwHUjI/s8zjmvsbUa/7OjPFmYw8o7bL4VQo7i8roYkBEXkEsR2qtwd
QelTTiwd6e4vKVFSY4feAblys/yj5cHARs29Tpxj7w0NghVlOr5a1o+336dfHrYx0eOvYag0DkVS
bbbYu+G8xKGipmEQHETjaOEgnhji3DFJA6fHExWJqEkAH318CF9kVwhSvYhlexyheHqPU3fGTYW4
csw3S0P1PmSygDrFu3GFNnuCAPHDLj6kqrth7pg664siYMlp94Cegsy4VRaign9QeX9BBdhLY4AZ
Odg7efvY+uF7RoH9iQFAvDKt9pJOsvt+M7jhuBeIXoaFpgR/BINFHEcT73PfRqvHVUp1/eK0RbHB
1jG2uzGC757JdgVkq+DY8pghQnxbr3wWZfwZTXYq6LPZ9r/OeXUudQdxgdpQZcjWAI0sUQYEPtm8
YVzfHNVd7ZIcvMRnAOk6UDqEorNumNIPyAT9NQyvYqPNKrPMS0kr5d0R6oICH0Rji7p5ERzpe9DO
GiSMnykW7xcwCNznKbDCLvQ/jcwV8d23ntpnLJLoJLXaJJnKV6Gh+6ICBoRCQFxsj7a+tZOFsE+P
yVHHFEUGSR7Mec/9iD7bsP0sREgAlsj0CbTm00JB4fTfqGq+uN7BXxThO3B7rxPyro9eqphk3x4r
DlSx6fAmTILWxnW2FhZSqh0sL+SDFVd4IDvSLrgW8TqHsFM4s+1FRhy3IrUQwWcmGrA4rELzwfYT
Z8F+ykZO1am9eZxlNSjnqUQbbfhWymM6IKukZIp/2OZMinCdpNkN80SqEV565UbntCIUdv9uhlsN
Aux+BVUuwqog7I+Ri/TMOEpLFlQzZW1UM/r5AbViy80/SlR2VknXJO6yl9k4I86svz3OFapOIee3
M2lQg8XUsIwhO/EHpvFb1gOPUPHKF6upxtZYH4cAZVZot+xcnidABp1xkmIxinj/T1lxe6a0LsOo
xxHvwD7gTY8U9gTBSZCN8pgJlCxaR9kufkD8TBH0PevCGajCj8DfmTiHFRqnz8ug4MD2DUj3l7XD
ubE6hRVcqQgwVw/tW8oCiNcTkXcIui0aOZ70zLxUaZv5O1LdK425l0ZJS3jVfmRAPvkF2vKR7RQy
Tx3VrgVimVXX1lo3PRoIkK4CeUhhp71eACki+uzB8pjsBzLYmfCfxhSHLU2QpZCrVIqNpR08MyRk
EeHiCY2YBWfENlg98RWOJf/fMrAOPjX2YuPPKo6Mgh388ff/9uj/TMIzmkAPP9uGQnv/s8Y+38nX
Tv+cQBmz7YVaB0Z61Xd+l20+Y6krZhNPbQdja2H65EfNV+H1VpIa/k2LTa+eXfC6eUis1fSYzhVB
mX5ieHkba63StD9/E870b+CbdT38NQsxeVIYRzn52KCgdUMy/gfKqrkaK62g5lLoU5DiODsRuWgr
nS+rDBFW8vWAZOPqPHT0og4d6wAP6Kf3KI4izpB/RK645LTLk6+mzvpIX06NkAKZ/nZfDxqArDgh
pOMBJakhWmRUcIAQlWt2PpxEgEgHmcCV+7qQKkrYDodomjvsM0bhiRymBX1au518kEK9f2JXtfNY
B/XgTgexMAEodz5qDUxxu4hRKtoFuGf02i5ycQsPnnzMi5Z/CDn5Odlx42tkK7Ddz/kg+530QdbP
EscznMwI1i6v8IgqEQ0GuS2iZDZFdqae5RS/+ZX1lTQ+wHZeDEQbElJ1nrULXwtM9ychNDF971bA
p7ny7bIG9T+6nGouyNHMuPTiZUSaBJ5pEU9qghcQAdQkx1BhYnA0HCxX1OQEYeFyCqPstuGsVWe+
Q3E2EqdjveRqkmZ+VIw67BkucrN4JdaB/vSt4AYuslLEEZPEE4oAtn0RdvE1qbgVjDRDC1jpbkMP
GVfzmcm6Ve3uyC/o3zaj8BtVuhKcjmWgi28sqvHnWXSF45aHOQBfq0HN8zPsdnO03vyVRG4/ouJv
Qcodpi0KoFENyB2B0MC8N2NOxMTlCXe20t/jc2bz2FuUxxIdm5tDHEE/GMtrguqyhDE71hg37I1Y
MjxZjFZNKZ/r2fV+N2E4GaRl1DxAVHXZWynw1sG28hUiynhe9erExkR270G4U1HnmVH+zK+4flsr
8j3wPY/E1H19AL/THLYSIy4vr685QoXdJP0RLGBYfR0dYZWwqAftGO0akgDDGJDlu7kqII8oLb9C
Xpyg2gEmL1xqcgo50cBpErJmY7hw8cCr2Z7wKA/NW+HW0wibiiU1gyHoXEAh/X61ZLtFbHml4SyJ
CJcG6lyTEuh1GVnTG9nYs3KArbNDZjKl9jyhu16V69iYh62GXRJdOyKlv1lQHEWFyHLzNB+9qFEY
EOohD1eiVPzS+TWkUUN55mj+lnwuzL2lKEkLbg23I5KrlArZz3rbxpkYQaKmkY9MfVawzepm3D7R
5gJDNL7ciGDiQb48gJYLuudief42NF4FqMCc+R02LpF6J3Yxyo2oXFvVtk0eOOq13Ep+yBw6M4cI
6LdtY4OvW6ch8z16xhvZwqpC7AidMuQ4X1BHM8wpPyaHAeTXGKnKyQuUenqWz7gZTPgGouky+FeI
szl+cAD68ThKF4u1THsKxMp0G2OuXOCQ3XjHFPFY7ek86/KQETr1nKLKGJ9LLOqaL1KPxjB921GE
sE0eagPDQnAqU6Ugs6EuJRd79mJgfZ6X0rY4dydBoqIGeaEgdSzsm1aBVWgfyYHtrpa6CB29sVZu
XgUOR6q67qn4Ay6JbihMhoPlQ/0vQI9lDLpdOtIlUcHR+/RpKMUikViWkTEjOkQxdPaHk9feog+1
hDH5SXYGjxGLtEY1Uie37uYAburg6ZYlwyFGb7KXN2w1yDOQpf0cXOR8FUiGjBArs80hmccfqAg1
ultmDRPT4ZxBE7rEGVcvzQR7wxemCySJAO8Ncmc5xZ6WNWd1whM6h04/Zatzb8Ho3xWy6PeNCZOy
xWvD3usGJMXDRe2aSqWzasHC1mQKGwZPaHBt6qRYwsO5Eda8GpcUeQHFOyLwhn8Hni6pIxhMlzbl
BeaFPakCKJoUj+RmzIMaRimyxcg8kLuYxt/LaFo/pwgo4DffvFV97Hk0XLZ6qYVktuaoqrEVO597
onoSrVGtJlWuMOfDmTfhdsktBDVyn0xG+4tCgp2VAe9AQ4W94tVpSBzn71nECcwL3RJO1lVwsrT3
62zXtdyP+tkXDToxslFuXz9z7Xbvomz7Z42Vi8a+gbAAKrmFlOsQXwbQ5jyBaFu/b/DYC/GEUGeF
MKZI/xWKWASDt8ZxxaAoUGfv84eBFEgd4IVlGIe+nh56UA03k9mbfLUSpwg8Mum0nrJj4GsC6rRo
MYf/hkrDCDGe8imC0bwRjxtUWm/PAGvWtIKNbLL5xBiEHnjnG/kGny+OL0nSeY+/nNXQE/csV4qY
5uSK91tciHvu8XLmRY2GVnrfW3m308qQ0u2uEMt2sIq4bb1Wm1G1lYvy13whnjcmn0r35RlRXBmT
Ksg5xos2qlTFMLCy0sKIVYoIQTjqbx0M4FvKwB/nT795hn1mCa1CQguTHHpx6RgD/p92cWVoGKQP
0uRiiQV0Uiz1HU4WQZSKyunbxSOd0W5pgqKttBoTG+G8qn8J7a54q6MzM8TNIqQN1wO0bGTiKfU8
3Q0/4ku9lUxUqKFwhANpi7JVAMGsQ8KAlFNdubn6xaqTrYDrOIe1kPVvXyhR/22ebUESy62kkJUZ
vxWNhxX3uSRfLCctioacHamjkOyj+ZZAbzWjOX8BNG4G3czmqaFuTkQ66jhP2Xrl4zDPogfZIJmz
VNSIcwVJpLEQ7SFI8yHB8Q2oKG6aJXnnzyVq+6yUVdLB9pz9zjbW0Ev2rJju1ISdJ8rs4OSvL47s
0x+olPccPtB8txu1plOStBoAgI63OONk2Rrtxf+bH6iUVrYPuo1gBCSE1BmpIxJO4gfagpdKdQJL
8vu0xs860R3hZWa3pwcNj/Be8gu3YrBvTcKDOKK60VWkQxXyb7CEKdXb8fDUrZxJ4cvr08WnO1Ig
OWz7siGxfChTe7/zmRo6pKn4jd3930KIqDNEoi3555kxNZMaZq/i1MVMvq/Pjgy1u1NOK6j6Dg9l
Uygk1wSQe+enbUN+nmgfRR6Qity0l5hfGfnc7VV2oa1kGjgS4jM0mKTgsPRp6aFjZcZomAaqhD0j
avIdMuzGTb7+u/F/xi/vOwm63iJvOZ7sRvWuo/wrkXq+H8Ci94qAPoSyqtxanOLCr9Ao9RsbdnEK
hk4/p+w74Q3tcqoECpZI6MSmt1xqs4uxBAyuWd9kjwMHr/VQszLm2XrKDG9+ZYkA2qevZPvWLSy+
3WP1DiNq+EX4BxelmFoXIR68s8N03CdviUaOzA15gn1HE8vGE0ghHt6tsubIHh7t82oJ9+3G0Lp9
cgxvxxyDYQMXTu7s/dES6FHhtQNde1Qa7L2R2CcIw13cxttZZC4kmLnhwsOt4OcaiUmL3+oh52bO
ifVB+zHYJ2IR8+U2SZ57kvfOjiL5t9AUMiGrvIby/yPAfNonUdy3WQbjt4qxmWzpLhPiGeWW9gdg
FF4iyW7k6Tru350VWu533LlKfEJEUd/Ac8SKIKcKipDGcczjbbMxF2zY2yuVbefPZpURsb3kY2rB
TJldRdhWj0EArhdRzAihxJl9HbVNcH8w6PQsqZPc/WLd9RuSBhcsVeGvqK2++bMmkVchqJOLPJLb
7MACFlCXUp6oX7DYkHdmZkE4XShL9bLTKxS2LvbOq0x2VtAXJx1Py7JtphquUg6QDxiURFKaH3M3
CZON8cQP7bqFwoxVWApO2VATmOdrQEN6mCDdJUd2wCdcEL0nxsBqkVIFXu9B6qiXsQdjudPTrZBA
VakXer68lP+XfxQjGOT0Siz7M/Z/uIRZQBumC86yWjuMokF9/J2QvSS8Z/13Cp5C140aRIDFxNDG
OJOCMT61/dfbtMTd9z0K8QcA771Yx25A7m7knsMnMzfI09iCqN866ZDt4onJi20F0INxk4lUhWrh
PHYUjf2jL8jeGz01ToauXY6SKqpeyLVzNr7ajUyCK/c4a8grErd+fbZeGebZ0E2uvWwiFRZr2VI2
66RD4dICCMI0py/OEuGs8ONc2H2RnOjegPGms4p8w9NllBimAGkQAACaH3Sjcvq5bw0pC3o+CC9N
gLMvEDwGs9TbcZw9yH4YDgMhAAcw9o17IlA03TJ8SRPMgFyL1n+gPHwX9vpF7rwXuO8R9DTsBpu8
+gvefZSnd4IEQe4/vnzf6p7Lu2WAQPC7y1hcQFDG8Uo/DNZWcZVaJe2DQe9DM4K7RzSU8hdHXh7m
HhGwGfDWrLg6y+VSaahu5UY4spC+umndx4B0XW093Hk5nO/GwJf/Fs7RdsvhPn/tE6dL0Ld2eUMn
IfZx+82khAyuxxMAXWIgNz+oQ2N+7CyWvt153MMhBeup22pjxI3Bb1C737RooGovaWXqX+Ce1XLa
mxsCmOxH3XeR0m3bE+cWcjmCSVXKJCLlLdMqscsgYPG+UX31Tz01Y1OfcDzdXonm/MN/N5bC8JX/
VG7P8yGaANgO/45vDu+l+fH1UpkmF+b+bxVI7bUuWpx1A6Rl8A42Uvjt+NDF6NZwNhyLdx0egaFe
VHidLDQmkAng+0ZRVKO9pfdBz2hAVop9JOh8zuguL90wH0lG9HncRjWRMPW9FHgZm9y4BspGXALC
tLODBDWKsN7bQcWd9cOnfG+XDODLVimywEy2kLdJJpkDXfUm4oAVrRKS1t1hdD27rj3B8IH9NTLQ
QEnLoL5H4nofYur+U3E5lTtcHIxzJvLykqLnTKpdhnh7KUnizOZ0w2qwPNr/qCv+UahUijSwqM6e
fkKv92MWlAvFOg178slzk5ArpWviEPGAEVIceYPJlCdoX5/lLWCbpQBXZBLtXLU6IqB0ae9fK1vF
FDzOImi0JZUH0lUQ4Vmi367ioUZ41Lw0JFBJ1y07dngm1HRtCG6iSf2NsKOpHCkLwXiXuc416ITx
0ozMK4RR3UZNytUDldLre+oRapcXjAYwxQ0aOAPrdFeQD6JF0jGElOAUvmbs06n4nV02AoBR8s9Z
NLvshDkiz7YpjUl1LszVx5cWY+gH2pIUyKkx419yzH+6TrkKyRnwiOmCqElZ3+gexuL4yzKM50mT
CHUMyH2qWEPefyh6EysEYjYg0Tf6novHScyLFR6grQf75SYL7KY1vIZ8JR4dH3aG7zF6PFIy8Kq1
0fF91i+Qtp4757z5cqTgIb1hT1SdOMP8tYkb646kkfMwe2insbW2fSoA/ZuzNkmeuC4X0vyvhGoe
+Wz019oEF5yAylRNbNS6bP4P36Sx60+6lUCSK9s6iFNESYXYvng6IOlt0PR7N2j0K8heFNnRcy4z
/iS5c5oyxrKGAk6PtnMj3+zMHJBf0sr7R+Yc5nNFRh3i9t+RewtyRW3acQZs163VZd+gDm+40ZjO
6pvyF+SCq2w2mGBKPsFXnQlZFgNsuXcEjCPtm+4z9AG3J2Wq6U1tRlSUvzosT3lTpkWsVOced9J4
kETVd3TefWNQR+n2Yryl1qXWrzPNziXSqYXiQ6uIKyVobv6xXzcDIUWc1GG+b4/wVKrUOsz0T/7e
K7myAf6ijjx/9wZWMJmYBdCTqzM5PUmWSpcgODl+pMySK1KrDY/H2zHAlHbFaYOFnp+pn7bR0Dt5
IkxIQWnuD/Veq6ZRNx0oueFzzCtB9Mf7n2eQuywzc2RnCBcqiSQQUEk0FAgOKrB+FX0hMNx/DDQe
vbDdKWASQdMNsq27OoJRgPhQofJT6Rs4X/NtvGdvz8R9y6tT3XuaCxsSy7sDEZHTQCRQ28/na7Gl
wLuu97yv6Km4hYxxwY5LCMfGlts8YMD09ZwV2Rnl/Lu8Rc8FQ4hzrK3c/hbDrcV4jOO//EpY51FI
5Y4g2QB38bZld6yAJq0HGxu2Vk8CFvHpmydUf5Ri1Zj9RWZpe2o3eTtlOUaE+Q9EqrxoEfS3wD2z
QILa9HVXzlsoNx5zeFsms8T2AYyZvXmeOiQCT8nsYWZg1rVFELGDRHUm5btFPcf+7or9gqhbxbrd
yn8aGLbHG7YgyGd54IOTMX/sk3gKOQymfy+z/YbmgO1WQd4rXGrl7TF1Jn2vwWN55mgN5rsp3ad9
xRXd5l1ITXhYhegyaVNaNX+ZFVMziBSj0krqTpVEPA14OytkKdymmjJJqpSrFBXTSq2v+t8rhB/5
+zSsuAKsEPYupR9tiRcUB65geuthrkcdk1DLJkHq2eALifixeHaEqGxxGIb40Y/xbMC9veURoLSz
Fx4T9pHn/6b1IwUoi+r5vTQT5ksLGU/uYpb7Gl45n3iJz/5Z7kXrAOH8cnja6CF7RClITEO11d2n
krUFtLw6X7zKOVsZYF9/3jRsOZkCXBLtemm4w8FKYQR4CvDQ9TjQy1uoQ/IxYqCi12OO8RUvMaTd
651OLgf5auHOkgYHZ/jaMgzZz0Ed2+c/PmuYCvcV9PYHtpiNX0XJLJDbi8oM7Tabvmi6XuvE/B+7
+jPKryeL1qEvRL2O0EZ5OIjfkJ8TDtMNBESChe8gPoADBsLA88JFrgNbubEdS9N5rxc1RfCEOuPa
j77k65yBtJ56mXhohiCIR5cBcwHckUYeGJqeWoPYjnWeDlBy53lIHe12uBmF5tYvOkUvonsyyNnN
Al60Ef9mgsyG7oo8GOsy7HYFAezkqNqv2YmCKeblabRtJzvV+ayfl6vTDBpOgLqmvAZkOl9edQVM
e7y58ge8R1acFKfE822ReCy9m/WI1T/+NSHdMgNsa6II6BGPqAg7erAv7Mq+A8hmp/Dwhsxbemej
jB3AE5I5CHs0V2N8/zNOaTOM03A/sd7cpCJdaKBFT187wpTJIrAKBQn5jiOeMeRgXY1ylat2i7ru
PUt6wjYVqMhOTQqoEpc19zOWE/XwBUIs+CzArhmeJM5/NVOg3011CDj5RlyWCbVjjEzOODf7suck
znZU9dseGf8BZdUJpM4yckD064R8a2pDP2T1BedQtPNyXv6qUOZuQF+i58PiHMxgeBHWPrhPZFwB
Ng9am6oVyEhLYIznpbsAu/zEQCvWwirA4ii8klfaPzhB/Rb/bCh3SbDD9JAJeYCfX2nDJ+daYEU0
db7FQcdJgzOFeiAACAoho0E9DAxfixccn8Hq+Uj319rn7BYMKN2H0vXtadmILeoUElSDS+B86gmR
cj1ssjVwE2qlIq+UhvCHGJ1YAb3rOnz92JSasGVR+AuvjkAHLqPW/ccvCUczPaQvRAH+CWX6z4b3
S5/JFN5TvUW/8uFJoBERXl1yjBg3KHbFnhZRhYNWplhRyXQTicORlEN4SK0NWhUPZXDiky+iTDqJ
hGhXhAUJQik1Xflw/rU2RVDGAT6iJX0IUzDKD7JNgY+74tx223u7kervbTFlJH4/4dxDF0UF3STF
nWi5hGcfIiNzLcL2c56KoyRFEeRJIxZYfEay5tWGEZmzNJnzS9Bko5TnGT1ZhWeYmPtYkXkyunaP
Qsq0vJKWaLp6IxJWk3H6VLLlWSvvz3i96QmIkOdOtMSNviIMG4+Faj/YMyrFTLymbsc7q/P1y2yH
s0qGjGNDMotudeoZ4Xxx8kh3nmwrN4+UOJx06NADmC3rhxPT64GUxDV28tS/NeMK0lJ0ySF43OPV
U+lrToz0pfCEX4XPIFkJ8X0Q9YLEozT2iKhvGM1i0K2c+9uS1+fnpCM6gYM+Idfyuq1uYt1zWsKH
R/iytcE+D0I2eU9iZEQeqwtITYLKhZiPhIgmR3emarpG1Zb53lj2ITBCiSm32j5aT1qEUYn1qdc5
gnB/wjpxQ4Vw9fcDnIyvLxNOtGCeIw/clL9HndcTutShZDdYUq0PUtq5HV+VsVs6DI/AYFnXLdjE
qmM6apPi/PgdLPYkmznfx3gWv7e3uhtKSjlPnKh6l+yFIc1FO/APIGEkStkUCdOgBAJdJihHa5el
sUgombmLPMdZhDZI20bqhuPUGDxBi+zM9ASgevRu6MWQxjZ1izqB2j1t0DoC/bps5TtwyP11ObAK
xkdlPzZS82LBu4TPSXeEDzR5aSCvBbUEWFe9ESpVANpz72SXBNVzaqEjVo1GlYh67s27AQVaS5wF
+jdztx6ap4dVOHjd3o2g/S1SvEREiodqzvvyEzs0K4pKb8bhR8O4lyZtQln+AcOmaD1Pap+sm4Fa
95Hc/+ce8aD4jlTL7JnvuVAQl5zrkcj7Km+F/R67Bhs+GvvQvL7BNbnQuduJI7Kjxzri9+4s+YgE
bsrfBCOqJz2230uX4tfY/qRH5Cm76ah3KuzUrDqyVGZd9aiIwbGPrtwt/ZeKVP8RA30s8DLaf9ny
WWaH3IktsPPOcHaWGX1DgYoACRsimqY5tBCTOJXdrhn9GPwzLCWSlUtMFyxNcyK/HX6bVvs3BaXz
zAM9SSFY9htIMQb90nYK1KeOVAWzyjEZHrFWQEvPrOW/lpRM+TTATZ/VWtpuM0ZDv7Xx1P0cVpHw
1jTXeIbgSI7jyZ0itoQpjrUIJtpq5+epDGzGNaNplzbFttZzlJYLsWjeykqV7iTLjVODLytC2RAk
zifSgK5wrOWNSPsRyZMWWqEj5gTdWq6uuHqw1fVYxXv8UErqatEG7GYue3wrf+uM3yYQkxB5z6mh
q6rT4ysN3LNbznHYYi4sg2UgzNhzo/EBsh7d7z6AspKHpq/XfY7GJOBIX76DFT/L/nhacOKl9HXp
I/YjXrATfWFxsR1urZmcpuLjPIGWcFgs+gOIU26M0nU7+zMo4VH2X944Txw4ip3j9N/3NT5MojB0
MCK6DnQFMhbVGwSdTQKM9TwjdbuOHNvEbBLQqmI3TdrwpCroRH9HPyAovpXWExphG12YvEvUAWT/
51lGIEJGVSJ17aH6CoqbQdvT1utsdK04K9OCCgsPT8LZvUilJYZbYF9lpHnE10NK44PyslEue4L8
8jLIoj4PzYT7rFd7rY7JaisgbDxSQRtUrbZjsB9tgUCirzcxkjamwIb3YK5hxl7jrYrbSv/hmK7c
Brq8aP/sZ96gO0r5M4TJlw0R0gggbA11j47Ue0FHXV7im6T6y5G/i5764RHnmTmzpB+hBq/Ddhlx
ctgzZoYEA3nnlKPU+B5AYb5rfUtjITy1GgnrKRT+D9IA8sHsXbGrkEiEFbImr2OpM2Wi0LYuLgr8
G/BB83xM9HC3M3J3Jyaj98Dr6Z6KCp02jCGWtZvabNMljulXzWQXF9cRdOJjl4+aHnLsBBVwp04c
kl/mQCp5SBbd4FmDSySIfoWrfMaOuOaMJdNKYkpiGjDYlJopg1OSkyC6Gu88hg2Lug/qlUsFnyrH
J5uorixd8o0ccKjsLG52olkgXuvrsd8chSLDo6EfQ8qJDUR6lgYg2RyOOaGgiSjf3Kc7bPbEqZam
RmM2gX1q0BaQmzG/pFd/lSH3/FEI/TGMlLGpj0+oXIel+bvsL6w6d1fOSMNK7RUkIRN0bG8H+fuo
dFIB6d9N5BqslPOQX7hsEoKbSA1Sc1GEIE77GQ0qrN4AkHaK5EICttFCsN4JTROboJA6WubQ36rr
/CLgZkeUqaAtMM+uG+hmTEy+PdlucTu5oMzcD6FW4qO5rKeJ2Dv0yXsTgzJcXXuvBCw3+CWDX/ub
DPRfJLMNq1J32VDF+Y/AasbmAi7RwVJSb6hckPi5Dsj2IH9elugKAuX84lPlX5ITU4I7mQ6vT8qr
rpcuuQg0UPjm9X4tNOptq9yhjF3dlxrXWiRgSZHujYDpVlwC7HL4TvK8k4M5NxKNRPB1Sw2tz/jG
ZiGOQEDufLq2Jf2Kzrmngi819UlFb6+dloLV6lHr0D9OhXIENsqqVUejYp2I63mN37IQMJTa23r4
mJTJPXSMqpFJv12HdeFLx6n5YlLC/KvcpXsXi2a9MJ65Ip3rfB4DVbz0xdtgIT5GEuqgokP1UgXO
YqC1R6gb0LhEa18+zeFHIgFOXOg3WLd1mW4OR/OFrtXMY/Ykl2sODDtrkurO8vypAzmOFLtLy6CG
Mgof6Clzl5VKDikMOHEqfveWzNCHNxIdWGOIINq9dDppHI2mZBTirZVNVKpF2NFcLWZUjO94GMx0
JPNyJMtx4b9fVj+xPQOehuy80jg9UmLzYyD9F+3hKIrA9cwXNouZ7a5k7r6rd3D+zsyWcx4xdTbM
Gc/nA/pUv1AJ+A81RPwkH+vr0du31lhcH5rcDW7H8iktAsS4jruqeI9+/hJaIWLwIEmqd1YwEkAP
bgROoY0xwt9mf1zQtBrj52FsP1PrAKrxom65WetI8eS/+qI9cgFWGb1KBCrHB20MnmLUzegvUWHf
BtUczkVhxIj0bG96V2ovR9/OaZGF6ApbReSz1Unkyxjl30PNBx1/+gjcj2i0QChzAte/yY0xtlNE
i08n7t6ML4BkBlVJpPSsvMEaQKAxbZlTv6AKsok1p6tk8fqPm68KDL1ZOc0DpU5z/ldUwfYkBbPJ
Wee6GLuy57+3iKFTKsWZz3QyF4vkkdnu6JIYR+f9IOCq2gRzkmgqKzSimP2WsfoRrbCPNhDWOT0u
ZyDP9cUYVzmxqAnAdSd4NGj9LnE9BPg74nqT2idCIzT5RbzhVzTrvXEZjAl7esM6wfiRoGYQIaUm
NEUjcqkU2myPwq9i+V62fBjLrh8eZn7xrxRvx04JzwrgtuYQkigVzbs42emfPkZ5dtx8K03dU5a5
MBcHEwWSBFlKCPSqQGzX294y0Sal8Qhiqe7oMkCfgiqHdtl0JFqIFNQt4LIYVpFm4uap9tgTa3G6
avKQDKrTRXULMOTZdABkEQ0dKLAaIAAPK6PGucB9XmhN0qXm2j/n7Ul8RtDsF3SAtGeEFiCxL1yM
JK/zCO5AvuMxBeLFjcSo+S7lODQwyd1IbEjFmanHF1l9bKZoFxgZX/UZNDCbQzQElTwa+oPrBOWn
M+mwnRYbZP5NDRSN7lJFc8HfSIUcwst1l3KgUvd6nYXjP75DZKIs8tMSG4ciaFpmJE0tyqMgmkzl
SfWQQ50mzHBsrNPLkVdMxaeh8y18zJ9hDe03JT4aXo0qhswbr4ojLqJSIVWxGnucC3Qe2WLGLMzA
lIzhxnzmowwT1VZoYH0AEn3Qo5q46SqzC21CvcRkgl8j+hx1CDduLG8tI5SttpG/g2n8YKKDo4eu
tRbYZKiH0Cx7mN8GEBR/1R6D+Djs6yvPNUjb27LSQlLUi3dFicCBuVdFEBPiuW+VFVfr75BKZk0w
8ZVVvwF8J6aGT/vxLzOrLVw+aAwTD4pEvUYYEONr2BlfUWhodtMDXhk0C7A1gzJC1Nm8Ww4fBQ07
Y6u6jxQ0B5oatFhIjuHrYwC0BWlN2cOIRoF1JeR+ZRwt0SgXcT62zpbM+CuqjHG4/ehjbvErVKua
FYTrx6ZKXUaRVPhZ6njCXpiPnOKiss/QBcCYP6NQbFDB/q1PRUGWmPkX+WqsJx1m1MgXcza3a8fy
n8lbczzqHaF7L5JtOUPEbeRr+YstKBMDv8UTNcZFaCr3wa4PzpF7WXeIAAFRtlFMsre88m0ebMCh
cCiy4Xb/2Dit+43j0A6Q+UkyAwOa2F6O0y0xsbT/Gh9eKlITmQR/JodqVofRNUXHqKM4aqKpouVq
eE0YTdDOhuUfLaecAnUA1Ajp0B50gdahru90bqCl5YfRn+CFFfSnL/gssqFLPkfWnvwqy45d5oBP
C8XoSyVGNtXCnxTTmMhQcAR35R5IZiYhlVUU4AYtEUUCLt835fUGIvjEA2hrFgUXlmjUew2+7Y3y
tWh5XFBp5kxXfuUJjx/i9JS1kEgZpmRDk89oUN+k+cKWW1CrA/WzU3mXWG1tXSUFteFpYuNUrQqn
gjJGrHfT8mUbp9hMC13750HEMYJ3NZkoJXaQxbkzr3rXs/LH43WVBj5O7Feo1XcRlXososCe2/4t
AR4X0xIsHLV5et7AfWTKGcvUjMF8cRl5NAQtERAwlMX0dkU7VwIqrxFbPg0tuyw4yIkK4jR0vYsa
TucJ58YsgvxR/bl4vwJAwFjsDcP1yrINu9LoB0GSTYjdpMDRPwlXrA2Cmc7B71v6wTHITJKMoPyF
M86M8RPFVeddupV/sED1eXPCysV1bkEI0hl17pLh/tjFSLngQJsTmd9+rD04MZ4Z/mYceIDUQdLu
4kSj4hupHQMfQQIZs7pyfr33lFOz8UUTSqBFpbqPcUSWg+hmCZ6bXxWIuCJqEanTMHTSh7MSDr0R
QeOp0K3TmmIbnGYv1P7z28Iw8a4iydpSxTcFeXm2xc+XlbHsj8R+8KuwrHfKF8NHjeKl4qJAY3qE
YWzWx3TkTM7DMwqNhowtQC9qRFQuty6sWzyiF4PdCt+IZzkRrpg6JqjOdJTnTDU1OQVJg7Kus8xN
qKKJgHxKdDCBmAB+3TqU5trx1MeqxNWraVyaqkby2MH/nKeRjPq8vNGP0Fom+9zrbxqwSgBppksJ
rEGXpoalVjtqKsMTDZbSMVgJScM7ZQppo+FuykWjy2HPIb++BIfZlmTQAluHjOZWJg/07YbSS4Dg
Z+h9nc8yj1K1MkrssljhgG3Ch1XZznUVC5StZXBXmh84wkuHDwtul6Z/IR2Dv8g1laqGnptJHTn8
tprvdXEGKJZotYVwOECShuVF/nujKmROnYfqUMB+/QwSv73huIRXhzH4+4ssdtIs/qOiEQI4JMOe
YBaG3XJiYyjVWVOQukAz0nMqS4Xd+evMW8DF+hfZJFAxgtqMq76ieh7XEGT1q80TiKlYn9Bumq7d
y6Jj3tF39CEGCLoYDHCCHkEJxGmMFgpdVN4SiwM3RsKZLIEb/HSE8NzqHNcmqaFldnJb6BGRXHmw
govuP38+/CuoTSQbDYvbbl7cz5iW/wrXF1Qbitzgn26up2oaPyjtvXcBwVfpseI2DrUyzv/dKJ9+
neT9GPHnWSWQRw4F/yp2t1V/PVIc1r9d7C89DEMR8BXCJ4t0iEZydfCfGDHFsOlHpmEtQHFujtnn
GzUE4h0lM2/GbT+kmCGKLuVfWoxMA7HUWLGQqGzB/3x+Q74+S5zNlJeoQJlfOJo1M7x11JghB8qH
b/AkqWNdWC8XU5iTFvCQP2EB5SwQYsxhZ0dGOidI2OORTXTjTOZdm4rkFl5J2uqKsBxxS3M6kipr
9ht56Dxex49u5tz/RRP0VX9V0iI0y9izkJrVQPKjyV9+4E0IPTQ792+RtiX3JoZe0VG9HmqPkoX2
Kvqa2wx9bUAvBLZN5J/FeqMMKq9wjMmHa4YCJ3lCRei/M9DxoHXOFx1F6EZ2eP59h9MIYHNm93Gq
q5kH9E7nxAaByCIYQE9FF1HBE4WXhY9PZJKJM3NaswS/FD3lNh12+ZLDnJgEIvP60FBAZpAohGmg
jRl8jIzeH9P4fl+J8V0/Lr9Csqkj3Z12/0KMa/GJ+th3C3MIgEosPmzFdqRumqYtLh2S5FkVEkcZ
MMOi0ZNXgbwqBRjw/uoUuDPAzmpVqmB719mEPYm9k1kUtlZS4IMD1fEjz3hS8OgHoWtYaaBoIeMm
qjoYI2YQ3gSYyuzAeZqikN3Aud+P5gTAGtMwELcCqjMoDYU5t8oQh4nLf8nn4LLUBEtMzvQrwF+Z
xX3oxRjcuvyKWXzovxDyGQ9m+knIMOcnvAuxmZW/e8susM29hsv27H7fQ2hOxblwkDBsh39slcBO
j7G9gqhfX03C5Rp66uKh/QNBqkJWdqGucB0xmKLPs5oH3DGOLhG6zTBT0dlPhMROs68FMrPSFBMJ
yDehfWzX496JpvNwzYyWdNJTq20hdUfm3Rup4v/28SJcPL+CIMqhC8DW5IFI9XDOCUeB9rVxWSMN
elQr2OHVurYix8ANWa7+uRysCYskbW5yvWJhCTNwnfoBkRtTSLa0WGE5Fb0MkLhNUkMk5CzWyqwM
SbWFYuXSqZD8AAoZmHgH+BbsVVHEHzk3rcekwr2QPoHzRDwZEgEPKHmzQRTFfbeLgfS9YVfn3MxT
uU0HBg+KwKqeuQeq3RbtoZfeNSNLs7dYmpkotlmW2KwQ2SF66yuAbIeK+45vAEdSy4WlQHbbrOJ4
DRYIU9f4Jq6cD/d0tWXFY4wAeunhXlp+h/hfK6yq28NakvcsjRmoWgDnKaZsOPIb7WGqMnPOGcow
Gu/9VHCPFOvyNkMHIRq7uRE0x/XkvvziGWObp9ijhOldYeUGIaRHQmrzZpsLAj9aAW+BHX6adiQJ
tvB+lu2hozOyuZ1mUv4w635H699d5RUgMWmekiLpPiVBTn02NjmXOyOnO+3/4zRDBkn1AF+wHAZq
MeEF79/1lK+y1WvwXx6FStzUPmmfot/wjDcWaniPR84PoXoQK15zgbeY39bRqMltKLZ4dfqDeWTc
rnnsk2FblbxQGD7whc4HrIpvB7MKaV7CaZ4H5+r+L3O7GvpQvTjjUiz8M9c9o4LngXwa8jJUfbkl
U4tHntu4sx/9H7El00oIjj8Rikl87tWfsrKhmbIncEhWMfU0pjmRHD92/SJtqGawwZxhBvVQG391
jFhZtgj/Jq6Dn2fqhGN+y+hYwKBnMbElQkmsJq9f3EIB0NEl8xNc4sLaKoosRyAfqbDV9l3F/nhH
3UYYuiaLkXcfX9N9S9Wv6NQM/ocijs8AzG9ChYQ1oVlj6yqPA26VkUOHe5VEFT3+6j26QBKnWMGQ
YXwdd72aqIGuklPJuoMHT5h7hQBBAyNnVx24+4LQZT4lYR//om+8WoQzxOtD11HEC/e89pMdK/Zb
Gjv0f1PVVK67nYY3iqF2rm7Y1+Y7oEXELfwV05mvjbVENVY6O6W5/tu+qzr0vpjf4Ozd4aHxtbtE
KFtzZ2wWF1iu7E/VjMfPopLmhOv+lVZx58NMhCPXD56s7YGpgRvLP4Z0U3lK4ukJx1fk6ot5mN9W
vTtM5OjrfnogkUVCNzugzB4YnCz077aX3CqpTOKzHcTPZ5D5V1NuZIfl/ia98WEi0qk3SvYAwiiM
tlZ9SuHiyLf6RWSwy78wAgI9OOdW8Y1yiCyPIFD03lYpUoAKvxyJ2SDb1071uu66Aay9xuLmoirm
3W+prEYOn+GjYhu/JEWkPsmC1ctk5hEKHO1hvr3va29zvU+i0G9ItyvDfvxrCPKvY8Q9PgcoQ9o3
1+j5ZED9kRBS8CbHpwUFfMb+GUoQqi5kf9OOIA5pUx/T4ybn+WkIk6HDQIhdlyP71rS/0XFV6N0W
fPx6lD+qzMZ4y71bgdc2bR6utuWv7IazE+W82TJ8TJAl0ELq9QaS8HGDU72JNAp2XnXAAdj9OECM
at0TXfF2izCVC3egZupHyGXyzKZJpzhTO+ttySkHFsApO+JwwxyoN3li3H1+OWrl2kaMvZyql1K3
HGgQQP+TUl1Y6kmWH3R4n/2L8NxBNFRxdJuasXiNyyCJcf9+YayV5GT+lEWLrYND9PA8SE+FvG9o
2XNzXYuqHQw6dDko4mnkRvRFpZgu21JWlq/6FkrM71zAnq88JRZquMTtaI8ykLkgxXQ1o5E7dey7
xLK8CyttlCYrvh7YbLdQuAS2sS6c12LFIHSUNIH9YDIsIUc3Hlxd48PKRdY1bJA+WpN8cr4/xUZS
nRP+aNHA3QpkYEYlvw1BsgWp3CHyv/Gv/yEX9f+jc9jvtc4QGS9uKtu6HfX/VnGp/xme3ZBvwKW3
qgCygKs6q1fbZCLWXBv4mqmyAkYay8oYI57cN5ZWmFS+5egyC4jm907F/c6PJ4L5WmidNNYmmvHd
ol3Hb2/Kem9gXnenwi4CK8paHz55U+JmIFyoNTx+zZMpyw00RcBncYVChUZwCVli1G8WgBWWbCuc
+AXxXxGtH+nJgoRuvdunvmW3f6XzuVk/xcwX9xREPQgwF/zAOARbXzt+Y1/CeNE4LnIKRyxgsbSq
9xxT5aCjh6ZDiE9NJX5VWLVDvhEDRvjiUjoY9YyO+aOFFHi/JI8jUV3QAOTt511QJPnONm24gxbP
pWETnd7L/cXfypGBEe2fWjjWPl4lVks5GsnTqWIZ2OlciOTD4pTn9akWK/lMK8bRsGE5w0UoUqsg
26a13wcjpl1By1X/Lh8/MUeZMTX8XH0Zy164YPj4Oj1CSHfOBPwI3UeLBGfsG7ig4152ffx29cja
clLGOx56AWr/ij0OOvo8+qn7+VUlAMukYEuWU01jC+jXwuM7LFbE70c+FVMua/RTRtBifse5Wivb
ek6GdBu3/Pz2V4FoU90WT+CZtbnaFcYyW4UKyO/BrfccEtB325Tb/WNDAOp4eRRKBeCk9pc8ZJx7
AWMaXF8iSyXAiy69W/IxvAOqMhWCoWJRwI+Mu/jHyKolXFFeWkMVC3dd24XzrcYiPDgZ8mXLcuNT
bc0ObzR1HWjVjZtlZYeNm2R6hCo2GVETAQPftyIcgnlQHx59qdlpP7Tfy2rucHyUUwUhomFXHaST
ufLIj9Xux6SFfDRbNk7CalqerTGZ29sDKd4FIlWyR/IfqdMW3rZyL5CxJSGlsJJv+8VLashsG4zr
qKXtztfa6unudaCqsO+us7rVrQuVHJLb9ozbDWYk0wRRJH5FgAWb6YACYzzcmsg3aw8+3CaOn7OF
dS/HvmSDj3sUMcQcWPpaTNnOtBLieB7oYig/q4EkibLE+dBkdtwuQq3kfs/Z1VBPAsG4HeztwgZg
Mje9X9+x84T13CEOgQ8N/g8SLuh1k8bDTEDA1LKl6PeNy8Pu5RWwOk1wL+tap077cv+1/MJLFfv1
YgmbiCaXuIfA6SOi7gkMw3iDCP3a0l0ubX7/2ZYPxOBDiiwJFKG78KrfO+fkiX02OG/PsYp/AxRf
CHSNKxR/s/cgC6XS41n5vOnILO9tNdVLC0L8ofYXl8GBggHYYsW+8Cvbs3hA9pSrZh69wbWXLjmo
fmbrjjRUlrA4yilF9NMhbM7Q6e6u5z9M6pWyhAbDByCOAchn3zOV2H8OE5tPqwOzpo/3bUC0Ndwl
hhyLm0bat6z117B5IWgijleKGoaK9fhR/ysy5ST9146JK6mSN3KZ93HnZAE/wR9FPZNqODF0+kCs
iyDAYZufxfZLILq9bsVR+3bRMxVR1BnZEkewhEOmvRPtvJsPSBRdtkDdA0L3A2yl9kIS+NtPFykG
kVFfGcrg+bmkFqUuJrTXy2HmRa77dW2+SIT5peGSGrLiXcBOjqn5KdgXwBLglrOBaNHxPQ4gPXRJ
6iXTrTlWveML3nXgvcaLkLRyUo2AxOoWOj/T0+YllBPr3FqSMM9lMh4/DSaTLtiBhEFhHagjw+CP
LotPl9Xz6MLxACFX+HeOWenJSBd/q7qWWobgf21ZCF9ZCsb96LULYOHvCj+2aLMheDbc8a9aqfkH
7Mp7CQ7VDOq9XGLLjnqjDvGNaOgqR9/F9XhXCmdufZu5lYEV42+8oZA8jzB2OZiEhwmR7Qi0yDJc
MT9heNKyheeFweUMF/2XqGlOSQ5clQs61jbtENUTAVwA43mLOTniB2CV0foWIOPLbLuRfqnbprCG
8Cgmv5izEhZ95Iz4hFI1J6A4NHPK3YinFe1UCkSt6jaYwpMewY74O6P7cOAyAnMWPBCeTWstZuQo
L36il24JPnLaA4zOs1wnjpVRsjd4O2dOxI85vSRga/Y+L6pCUCzEFNRISXEYfmJKC6s7YwazWg1C
URxWZlo+A+6qRlJD4Geby85Od1eT7YVJp86lhK23eW+ttHhcHVioKGIqwmMlNYb2hURaSOkSGaeG
DMYZL0QWZ1ybe0DwN1I/ki9XPJgnOUcEQlkb4IOaCWlVUheG5kX8oITxo8Nyu6HG0Pl2ceSB+HNN
1Ra5hx9KdODpQxLlg6ZLkje08+Tyx1gUmE0JYmh3QZ/0kC0Rvp1lXpM042ln28PiGDYWG23Ph3NX
jwte1ELinIVKY8Td3whVuRUDXkpjOGbsqCaj4UDwS24W3fbdQAZDJaQk2M7crCAi+/k+fZVEv3+0
5N3E6X1DtcXpFMlQCn7R3mp/dQbAZqKTyqTqa+JhsWrs+vAhSrC1ryNLpn65vJP/gAvcwrhDN4Ow
kjD4cHXROP0/n3GzMYL50BKWouGidnGr8og26RAJGBDY/0j33D6R7BdjhWgTNjI37G17i9cBd8jz
RUI3M8Hv8DZyoMgEvY0K17ctYvQSTzdPnKHmC/+6Q32ERZpGbHfbzEeob7R8nyhAlPlWtUHSYYoC
DdUyPxkLmLhS9l3f908ZA7excqf+mLJL+XlK4VqTQeWUv8dfmFq4y1P59BqSzVSVf4SgsIwgUuE9
fMhqCQdctryme+PvWkTNikriBeQhoUmZOpm7WWy0C5DttPoTftYKX1zagoQTKvUQ7aT8FDr7lbSz
YAVpYWF4BeWB/fv9bZAr3jzPjcIxie7EiP9z+8g3F7Yq1NbY1gAJ0/kmv5xA8hLVbV4JKhvKl7s7
I4q/1qFHeaFyP8fxdWXeHQGmqV6pZjJjOhpCWT+iBRpr9GNPuWCYJPJQ2buIf206cZxsdQFGPAmp
Aewnq8t2s8DAMaBuioFPw+6weCjNxu8wshVmrgoJC+fA4gspQ53sZLy+VYv6ZfA9o8M+EGdUjwlf
qG7RMB+NCIJW4AAVEo/ZeiWQ+L37SFyDK25ABjd/sQzww7EANKGb84IISDi7PsY9IWHxGe1TYsvp
Q8r4N7bvvAZx0kzEVFzZiVo47Ut/SYIEu/1GnQhScDr4Y4LGtRe0ZSphSxUauFWoJDuNirzjPUZl
xDyT7EAUOxNoX78rFYDFSMw72xTZVT6FCAluSgiK242cp27yEmDcmt016AfGMJS2/gJAnKEMLlZf
rXC1r60ah0XxQEs6OoB/GD2jZXA70Ik24cbMmXVQU0wsA4bdCcWQF9Bj2i9tAmZozNBkXjF2RLSm
sOo6lYcP0FtJyA+vUGUQtDXorUmdBvDA6z/U8YWMlboi/dx+vIAyNFng1eryH3zYfgecydSOUpxx
+frEh8fgr6xP3UJVRhyMIRoct6cmIfsGlgoUNP0KhrSpgCP0BQ1DQW3vXFq1P8ZVV+rlWZsv/jHX
AYity5tlcE0LYZQ2ofSeDdhXn9wL47AKrbi6R8umpci6R6yol1kQ2SK58i/1gRbsuJ7Dwbjp59gv
o/iMI8gI8jlUYrNogvKvp9miNNrSju1JECFK93P4xRwxe0S4oXMCOis+IxB9YjdgAOBa3dw+I7hx
4Tr8F4QetanqbrygtGprlB94JmBqn6AlflLItQixYQ+18hsuvS9uE/ghY49xE68cB98CAypqE8GI
3i1vbtkqbKHfz1HENEd/vQnLW6ePTD/uubjSRtByzOHYBrUGQdnoHxcozaCd2k0VI5IidLE+qR6t
k+qbj784xXvnGfCqEKcNWrzwvl984E/8+amSYosv1Nd7yk7puE+v0jCcaHhtBZ/Wkgn5ZxWMJjE6
8TOLhLgbtH1RFsP0TPkn1qXe5fxAO0JZWUYUDaU/9U1T5LzMbfOjbGWfhW2SfEnHDWGaRGTuj1sP
K31gFF/nHv00ajljPp2l0j+hytumCrgv/Qw5KI/eFmYfXXygP42K1Vggy9mE8WkkAbLfdAh7D2Q+
qAu36lWOzRXix5vEb+OrDBD3SdiQzGaXtb3dW8hGKAbV6jRqs/AkO1K7waFpI1XJ5IwDLKm0GGhZ
D8OGSWp08mejBEg/tWlx+WOAfRwntJY6Y23hw01J3Ye5OuNYWPke+jX6GkfYciFXYl0azfcWtMP5
vgEodA03xVreI0zLx3ydFVgziCYAIk+RBypeaBONasM6m2hS9qzUS0Gfk5Ki7w3cNp2hStL9X6vJ
arD7sy7AK/tj33ZIl0X8TrxZfQsxlv95fsBzqJDbU7JQfR+GpVTMYrARTxdDlmFS66jNm+9/IU4u
cbuiuaSbkm4wrFgE8XD0ZXfkTfHG+D9hkjSyTm+i4QES+H2mXC1udIOVI5PSni+9ftXw+2+jcyh+
cMooO7rRnl41wQ8+AvdWk5jlv41XuBs0SWlb//0AI+I8OutzZOcpCbRzKkXaiMICmgbHZcRa69FM
ZsFh2oxlCiSR7zGczOAh8rvHzs36QDdPu9B4mUFvACsEpJduj0Pllkh1uAulKmZwTEo9ReVduxrJ
rM+sbnEqZLhcuBXACs24K/bSTJ5uSOzcuny4EZ3HP4sfSGIvIk2LNrjVK46+MlR1+3zOEZNztRws
mvWT+FK4C7s3Ko/tZNLiOls7uXzKpkNB8bL52F/gJVVuar7ogO+PwNxbEo8Palyj4VHItDS5Oq48
S/PtziKqWeZ9pOwbcGlufzNlblhbvrPX/14WOAEdSJrBBR19FwITkFcv5vF/wqBlkZgkkRTaKmHG
3iXi7OlhEKc9moosoe9jhxzZl/B1Wz5ysGc0Kfr0jJ5xJeUpkjTkVOr72Ppr5Z5NzH5i0+V13Vlj
7YfdTwHvDQ3vY0Sia8Nx0qvcRoXeiy6Xo0nw5rMqPrDGOyjb/DEk1dINmbHFOcs1NDjm9SnqJYL4
t0iOUED+V5sfByTiddBwrrSYly7gaFgNk1avh4SZgDHryhvxRL6CZ48dOYNRUv/g7gbhoKjsnwJF
mobohGQ2IcaAOZZyuhHYHX/qeHrRhNH6IV6vQ1loqvcePdQmJAH2af/TKR8ha0EWu73r3kSRM2v7
Gm/SbX0WzvhpXUy6VQUH/DludlSHNFR5MZYplKItPMQkpiRmchSsUTs/gCBkHpH0TcegUYGzPsXN
hE/Y7pSGPIzqOoTLe8DCvuMXdDq+seysdlPM8T6MBVDL8ovB5g837Rg9xfHTOgxjQp+0wu2wiKuO
yWRuMTwOARlZayI8WgRdc8lXwNG7TBU8pUhBP8qzygo1ABafu7KyHanptq5/dA1CC3sGbg3wQ21b
2w6G7XDTJKq6trcU5VMYwsGkwMCLrIWnOTk17Xuq5x8BJRXpx8ZrpVjIWhkHq2xa6QxPYrOvYtPZ
x4vIofMgeiEgigAQLVODS46j7l+RZ8eqJZXQFCZ7cOHRt6M+5c2keraq2BVHBhBOjAPQ/16isORx
nf1ZPz65exqnO+c/pFMNVnDWe8OsNVWDGP+K3xFenOkZG9mo7mHHCzqoaK7NMBcr7uBhcZ4N0Nw5
dHl4B7gK71Z0tDlHbPJsb268NnPAanhE4qD2uWf/d08awSc0JYw9kl4yhhZ4r1yRkPl48z86wpMl
mJjfFA5NxGaCc/3cM/6m7DyuxvZ7znOqzgiGeB+dRZdnuvWNmSjS/MOn2MTb3Jiw47oXGWUnY8v7
3MOQPuDelQt5z02FpxFM0wY11RiOE/ikoTN788GdEKJ+eHGxO2ZhVYykuGGrsmXu67S32VTTmnRI
exgucEDcOVTVan+8Vc/DazahORFrQJRaW4hWztmftKmHlQkwkqPaW0llGFJ2/ervtojJXSBv70bk
5rbJVkhZffWbay3JQD5bTiKpeFnqTi7ETBYNfiFjkDGfjQdrHY8cQm4C/eigzskXiDgu2Gw1qzeF
gIEUuERYkshLTGq5/udjVC67vNN6FoiRReMv+D/jyp+c5J6C800bVvw9wp1zamCK3L4GhfnnR+Sx
Kor4gyGu0H7QM/bGhailDrc43eLfLUaHKIuTsXr1O1VUno6gbFHnuoQZidsVbwcehsSG3nfE444X
ck9eJQ19HQPTNxZDnwsE5bGldUHIeSCGtbbbhLsZKBH9cvp8wipy0zgtlcvjh4gunDfiQViEwcfj
KL2cQs+pQ4+NM+dxNgmBdtfFNPbD/1ycOBVPRd2hRuIVtFpwRjQKfhc8sDVC3LK9RndysWwHtQaj
lRSC/S6lco68sb3BCTV+hIP04fm2X6WGzTKst0nALJicSjCjwm8myCgdhwvF7DS6WONqpNapZGCh
Kqwiaqomn9uFrYodkjAEOLhMA4NPMLJc2OSgnBb0ocfO23xXBcrSZ4mTj4dTXCOlWbLO9Q0i+g5/
SyLdR/3ObdgElrQHKn/SzQZh+iS5ydMz8d1im9gvHfjwuMPmWyi6MxXUVSKrPuB8WVyHmdLXcm/R
7rzxCJ2DByLUpKhEQoQ4HnIqXoelo1La3ANNSYMCb8ELml9gZ25k0rMzfH7Q3MnC3+9uTW9I1y9i
ynniK6FR/poKIkCf3SjrSzZW70YSwwZ23JiLVPTB809Tu04GJzZNVsIApb1O8vRcRPUc8/s4hwSx
WipZ2he5tnht2p+cD/Kb4ix9lrXslWO0wtPqPYtsvyeo9TUWiVkfCroWY6VVbTYGRbl4NgKAqjv+
NeHAIDDQpZSCvHXB2+1HRh4/f0eajXMAXfhMDnnBaKK/XbSWk/q0pOXflBzUMUB3dsUuJTVHh6co
JJjhIgMhdB4e2Hoc9orsAhX26ncsH2Guu6DcNa/ypMR/35ck8IxIX0TxHDVl6RssbQgzGNdQcABZ
kPH1mS4hqUdg+gD6JoBsOx1itMdzd6OIkSEFqErJE9Tcx4knRVSjGDvesb7nmhvwHdtVJo8QovRM
0A+UdBUm5Z3Kw528JtGSfIz1i7Cg2OP1C5w4HnRhR+Fc+NjGpnsdqQogsLQX6/cBg7m3pptxbCkm
Mdqqm6uXqsovt82VRz2X4mYjjTJqy1JCAtEroRYR00T6XtWk3VAguSfD6Q0fbnf4+8Ebnqg290DD
H2iU0J7s9jSQRLIMxF/N/0Fjg5ngK6OadAO7CtrtXuUxuzxX6Wp78ohP0T+3nBevFr02X/judyIB
TpWR1/fx8vC++YcXLDvLYww0tCDos0VaKnaqGECe8S3jYW3lyuA+wrUUhLbcMaWd3h5AzAku0kcL
eQd13YrgUCCjd4NTSGGEtAM9BLIga2KOLkt+atq3hKnbLyZ31mH6QP4VT44qCtnvmThX+8aiN1bA
ys2xd9ofj+UOwPIIPYbRf6DwArhwhHfGqx8X95DaLCx+5XpNjrnVWYiwVDv937OeKItO52BNgjPs
juyg5pDNgR/vv9WAkC2n5u30/B+FacLqu8+P81I3l+2cCA9I0EejqDXz/fyAwoWOkuTHmb21HAxc
dvZUrppBtPSle6Ydu/Ce2srETUsRhxzkvFZezGCFUKjfzBwVV2L0kZ0/8vjk8j4iQfTQ5ehD5PGw
pm/Lc0JztZUBwHRssTTjbkL3Q/CvqGWrl16l5OEVyo84f4zwuCV3rVYl0VRaBN1EyWsr+KYnbFn1
knlyIxu6EkvnCYo5c25kxNVopTIV1UDEQB0TLEk2rbPlJZirswqTjMYhvd+ADsKuBCy4QXjLy9Jq
EgzHqDlCFzunwHp3XT+AM9a5+e7iYwDYdzh6ipfbeP7SftWy0D/x9b1xowaH2MUz2B/imIBEPSQp
/j1BgyKeRFREjwoNvMPg/RkjthKzuTBS5FAhm6qDq2EoKWi/1CXs7lBChkVnIHIW2YjWg/YRpcxc
QxnQbIrES9uucS6MQlKn4p5b8JZhaqJupSTxlfer/yijdq9m1Yrl782jW630SwlZ74iYjsyj02fn
cXmtcyy21/Y4R4EAwhNPseli4RGrq9vHAkWcfuYaOE2JLaJuqlCf7AA+a7mczngSGHZy4WP9Mg4/
HSJTZTIsqHP/5IXvBuZ61K+DK1aFHv/AsA+2JQqnJkzjkNn3xlUZj3mgEe8I/fgJv440sKp5TXv1
cCAkASLfb5gvGuXvVrM13pnNef212T4YeUXg2OXC6RoYmK6vg7N1ZwvmjI3BJ+k2HQHLBXOaRup7
HfCMa4I4ozftJedPXuzrOk1XGBkvO8VXxuKiTW6IG3borwylkVQCU59Vcdms6GKhOcEbhtc7WTHY
xry7AmgKHNWqzhZWathmBTPf4kDM+8fbRnCV0rifcHk8pWcOEQt7jEYmVv/mX08uxmkfNy5vrmQp
JMigjilqTPZgflVgwJz6532HnD3mev59eGSkrkrHBEB7MlKmvJXdtzgtai2iHBfcSY45HcT3ln5p
K9KAyZVylJ2PssQTeLqkxGl/PIdOh19EMxGVpmJHHk/zhrG/GiRQBz2+BQl9fvQJjV1xbLlxU2zm
RDiZAfFjDeJCGICKp+iBEPz1MymaHPRFgT9FFbTW/aW0NBWJ3j5AUvYjgkIWl9ibJ1QtrX87/JNj
2k5nloZgu8JdlVdFbLjLt5ilKcAAEORd4vB+8VTCY9hbMm9GGTEBpbifwKt8Hl4HqBy/qPGt+Iat
txC9NzWgI9v2CRvVgny19xqJn1fYC92ec9XeyiGSeZNdJeY4vYkRgQvCWQYcyM2mshK6kb3qFH1c
eB+VzYXKKATXhXReZUDkPyt1MQLy++qfkI+0M36I9JOOpIl1Unw6VfYNe3Lz4btoA83q3FAD6UaZ
4QIMpMoAqvzl5PVkOy0TgCf9WshtEkePkW60RBvcf9PpCcahs364417SWd6gmIVLjYsJCY35kPJ/
uTckm3e2GB1QNMCfwk1cH4mo/dVoz4QJja041IbIJLLuhLoi+sXATdTWPXIhn+ZwXjS878mTcY4D
pREQV/PUV/P/YuD11qAbYX2d7DD9kkmCf15kbLBfR1H0hNNhyi0B5Dw00DcABnPwTDMAMYsaMSXz
3+/XM0yYSt75lgUBA7SrTjBQaaSO0sjdkjbJktySkjMIkM6z/szkX9xKYbKV1FNE3Lmg5qdj+Jvf
u/4nc76YFKgF0I8BCNync4zAbdaBNQwns9b8we6A/KV4TxBah5Tr7wVDCXO0yDeoI//NPmzO0J31
h0F556uWWjHFTBy7uhAIpAWK51eq/WWCs6sh4ySm/8ALHD/J3enYwT+lZYhnxuGxkluTDz1vn+KM
Jgt1C0QQig7FWY2MWu7C4EtfJ52tgiKwy1Vmv7Nvvr7TV5ORmdnVaFAX2FDlTJxEQomn5cXctOv4
aGbRS1ywz4CieSOC4AKW1vPgVUti29iZ6ks4wSoluo0ve/gYfVcf55OSk8yiZzk0V4MF347YngaX
4kWwvQbs4jUVvpE/TvOFSfoFxmCwztNy0ioTN2VkE5BS5tqVsmX/h+YC31tVspvcXfrmG/JMKUOI
gGdUGeMEsq5fL1ByhPZ/eR8Y2gee63mL8PwppNq0e3Q6nndEA1BEJGxHZEaDjO2DG9IW1w+GJpLh
nlFummEtlTZ+4Y4Mq4AuXJZwN18lRe2pOqeJaShiLFfwk67NqIZCU9da4myuyJkCwcr6wqytMtAr
vbMK0fxKh/uURh1z815AgvAkzRabcSGS42ocD2ZfkZWjYkAJybKdWCOdiLSyJepHbZP2EkYeRS7T
tbdwf/bo93f/F8PHJ8TCAAhofa045O1J2pKj+nkdl5kKm6/ljv9PFuqmAf0AUNBTg3PuzY+VFZ8q
EWSXmYX1clZvoJqJwIncdWF4GvCaHlKEp+CRXvPu/Mzvrx5QiZ9NdVMLJg54Aja+l5/Gw629VSj6
mmwu+6KeITNzru6VscSm4dcCOJoogjTB1SKw7hhvnwWk8U5w60/Kk62w1iymWkFwT+dWlP8BDafO
sUSqJzPo8uedIeQwvh8Wv0FM/T/7e5WPHbCyXaS4s+kbg0PB7xBu0xSYKtPc2oykbFJOiH7+NFi3
NNa1VwuXHxfdZRZNRHxYxApYgOt+G4ONzIsWpGQdZtC+5aK/fhBgWYG4BuQgE8OLXaDOywUw5scq
3haRQa89Iz93H4dbh8tWMXmC2fcnFNrToV5mmAL1ml8V48sZhz1npF4pc0HHXbf53LIcyM64OfWw
d4pNOrH+FVK85+i6LoijqWHrz/m0P/7fn6uS0L6KaqRy2Dzn3Hx8l2ZHhVmHWm5ztRLewPjSL2b/
EJorqdl2pNejTwcmF7O/MyaQ5bmSLVuU7+pGShpReQUCBzsiShPtvccFT6VLuxG8/2RyCACjt4Ja
1IZelZmirSZxT/cSt2yhgovCTcaJf2jj1WtzZqmJ4QjeOg+Q/N0nFjEv0r/01ovamwQ1wyajh4vU
aeoFw7z9kBChYrsj8UX5g9yXihJ/0lEzHCEGcjepP/TWaO6MmlU5YdvmHnsXn0vLssKbFksNdosO
6oKpPAEaXYNuJvD1Mq/mUByt28KrVJUN9aJjRM32SHoRt93OYBT5x1cJCEGOV0zcB1FDRc9IwGAR
tamcPzzQWSEyIHAjasO4mMeo+rz+K7khDM0GWHySmOd68+XJnkLOrF8HnofniG798wMm12FjPxfm
nuqyCHCp9GY9fiXPrASk0RmRyH0X1NiU5HHrjPL3fbYpE8VJkRdNq0oPjaFM81F623W2jdWznWTz
mAt5UmVin0fFfPd9fPOMxNqrE8kWMcGBQ3LJPc8I6ttu5VB1dFiWT601fHo6DgwIRwLiIpV8mirF
YoFlH7ldgMnOhCe8g5xmmtmE6PM99ugt9hsU6tRGLkaiviA7QCWwGlJXgtXVBn0LthdlctKzZ27C
ZWnalGoBzjsViK0ZJOwxnZFpsHxiZgH7Jh+itSUts3NOko+8xIPRZSTUqRsO8H+xtTs83O5L30cr
MiRgdI3ptO1/YeNz5TCW5am6jvyd/6KpAAcE7NQ6A8LsF1EEkiHRBoAYhlOwh5MtUp5N8GRkIJUO
etrjlcgUMKxP2XW6mVB1TMbnD65gQ+kInbVTgSDUmpzPpcvYxk49BHUvnsj9a5ToBnY5+2pExkyj
qA1JRNg+EyGeFnpYM1U+u9CGMGosZpFRUixBUZigqXZ0jJazZgVR2iK5J15duCVQifmKMsA9s7RK
WVPZJvB2zKIR2STg276pA4Ok9ZvdJ+iKvmcPzByQbJVJSAdQX0Omu7+F25W0AhUBpUN/frdpQTMA
w9+kIbkISKV6qdQ/QeuETzVNoKKm1TnwRCrGrOb7M5HnpiKEwGrEG85k/tG/HasyQGOBC5ecf+x9
j//8dWqXXfbl3V6meHZqP62a05MP6pXdcH66pDMdCwztCvefaNXIHeIbOFbK+j97k7Ioxp3TW4Pn
BcGfiG0CvcjJ0OQ/3+v8YBQ27sS6rnTMvMlfvMwv1CkG18aizNgv41xkagYy+lF/+ZUavxwMSZTp
Z6xAf6uIUH7C4kKIXGNeTPvK+FUous3pGxL/a9Vcaf9LV7VjbIsAlEY3zHo2Dr3zZAByJmKa0pFB
iGD6U1EIdU34x2tNcv5Vp6HjwBSeCxNC/Jsx2dK/9WKhEuN1GiftwOe3NxCZ5Tsc2E6eZgambyCc
ywSTPcZHS2t8ork5yWSLLRIQOT9J96iIoqW5LHeEdGl7WEfCVoZv9suFMMBCzEu5uh4zCTMK9beq
ReNGT821KhNCZPwsLTHZxYDEJWo965t45RomihSyoQtumKk6vZ30Pau9S7JPHGzOW72yogGcsxEy
PqRrmugsxBR2ZGOmGGKLH3dWFCELmDGMAjwxGS0t36q8jeZ7T6mgYCT7/Y6bGgkGFTtC2PyduBOZ
jor9gm0T8uLEHmRhbf2gP3guFjKB9GzmvOXPjSQIHvphQbu51l2rxQYo40pwU0cWXSNhfjSjl2Zl
o8PpMWAwGt5YzRDuuu+7B7JoU7rKco/fWPKI4Yzv4vgicjtpn769ERPOxvPdWuFcQ/rIa/86C2fN
FajQpmWBxPbgCXKXerOOZ/K3eZCLixCPGEktA9PgawDPCZ7OP5wIIc8hNQS0rVOwU/xhyI5SDh2H
/Ot5PDJafD9oSPXv4zkHtNAFfZYg2s+T0Os/X0qCWpLg5vzo7cosIjpqzRXPK6t7IvrmzxeZKl/r
yIABK+qaH4ey1W2oy0hSCAYkyz2SHkXiBhy9BRyqLEZx8IGapiHyMz/nI+V12Gw7iu5fiRWFnbEi
yBb3K7elJ1YFthEuJgzCMhRLaU6RGgG2VjyUI9tO5QDj6WHXNcAp9ABJ7Tg0aMOYDq2Yxb4hIes7
ILYrNURt5jjFbQuDXEzHDlXcXwjztNW+GkAXQ1w2AwMu5eF+5DsTqkluSW8q1xCjChGtRQyCQ5iF
cAwcmiJVbucjnfBU7MSkDuSdGAbiSpB42ODBFY0IU7EkBTtCoSF74ianbxQDSPvtkghOF06DMcaS
OTJ0FQPqvp8ZxDGH5d44m6uXhwDnNMNLx8PwHblAzw98GGvahWly0pDU25G6FqGHfUv92tB0OmJI
7YK4ZUOlri9kQ6xOlhCp9C6g8y5ECzvi0EzYCCjrfiIFOk6poWyauAZ7UgPiDxGmwuGPZ+bufPD+
vKPMHm7C7c/GTQcuPYXCF4cso5eFWOzU4R/lvssk6SPe8X/+5oCSRROaD7arTgPlM6JJH3SmtsUQ
mZ5t37RYGyV+EX1ZhXz01+22vel5js+MCQBCN8xID4sqz+XQ+Five4ddWG5NbDl4y1vUsXMLbHjc
vKARdo6QkV5+jMr+WOv23UD5NXf0O7CEUC58iaHQeaO62dTwabzAePL9OWIerGeBpCMKCoBh8oMr
4ZTTLxZ3gY70PG4zolL/fp8Ta5VTLdJ+7JuoFBrSh58p1r/K889T/pyv6pmDgissemwSe/rpU5Lh
69X/MCQxTUsLJLyaeV7vmJsfQhnBtb35vyB6vFod2w+rZ9OcP2cT3ZYKjovW7hY2LxGa0NInQRjq
K913FkihyGIV0iynXDZaDAReEFDNqaWOmYQcaT5muBwoqS3YQJ6PqlK9tI6M7FKl64hVcmaFlyGc
c5RsOn6Xn1tI09wFgGP+vbkZMFx6aGflz9tCCOOONU4PMXJDdnJzMjiY6AQQ82Ka+0V+rl1HF2Bv
6xLmjrLAP+dGU/RQiuU1EbfzgGTJP5NLYJRkIZulYJd3lsIZ5XGE76xwmHBMHpYaslh+4GI0V3Ta
lfFqSOcBBfkf03LJAAZxGo0rYemdS2JB0xjVrOkPe/+gfcVExnVOUm3R3/KNPLtFc/4dlOHYWrJi
36xLfiAd6Abzl7jZHdvm2VkzukOXmJADMyIk0OIhHsAjr8K+KPwVZC46nGhCtexupx4QnyPIDiMH
2qNZ1gVCScLpHfT3wLQue292k1MJAli596CO2LTzIrp8oyZcJgpZe+ZxAS0MxN/w88Ee/UT4t+Za
Hhvika5Uz2PqGnW1XVpKuXn4Cv6AvSRv7CJN8jFT6EHjwVM3z8a/dczgMJ5XvRt5ajkmwEx/BdgY
v2sXIph99gYv1+h8OSkcxxMKNxFNjtUbwbXwXqqme7jyikYUdaY+KBKZ1Juh0kctNzwD16yUSCyk
Qi1j+5G3G3TL2e7JN9j39HL/n1KtlSmYLNP8tMu6QminSyJeLnb+k3F3f+zavALCYIwh4aQjH3bn
U6jTTgVTfTV3vf+HVvYM/MqNtSWYD0U0u4T2F9A6aM5X5WEEU7UokqjFnfSQvfLVXxX9F4nuviHe
76seuV30L2CZQRizoCegAqVnM4B4hvZaOpSI2zguUNpHFSWWrsq8kq5vuwiL9hjUztQEr97aPYXH
tYPGaaOvGuhUUnGgCI04RvQRFuii/PwTFn4tEVt/aSl3ARrM61ELq/AEDy6DT+1uFik54voDd8lt
SJWYR/ORBHfZ9eocKyG91cXximEZrAHvUna1jh5azs5P9uDh1TXDurAK04CFw6KgqY9tLGyYr73M
6+vIp3uqU2HiNb4EMTmq5h4a/vnTM8ZAE7sJqUijHvtvxPWECjHeT9eQbELaJlmNOQyB1K9K/x9o
GMAlKwOQShkuKW0Ai2gjkXif9agWc6rmMTm2U2tEfJFn8OTWEJ9+wMj6baEArLWxUetWodRwOBbv
l+btwOshddyt2C+j5X9Ympn3d8Iz/DxPHgNpNQDfnSEWcbMCQr4v/TMnzZgAGhcOT9mxTqhcqp2o
v7wgXFnEaCUXYs/abBGA92VT6b8l6HRW575pXclqlPKEYQs+viZcJzjN/Z0P40ie2ZETROWje7ax
bz2V7/JjQNgn1Gxhq1i6ETzkG3eB8RSOFT/P/uK5zHrs4YrK5k43GsOhcppqboQcCvZMsEK9Gs69
mGGl79UZW/udo/ZH9KgbiRq+Z5lE4V7bTRPTNDnjxsWoSPTh5YGoHsRD1ssHIdggEC+p0xTyuLUe
zwyH1i0nGby34zGtcUyU6IlAaPEm6raAFcfGxeIEKNr/yyX1QULjCFjkqEQDSyZH/wBBOeUDNYSp
t5epzIKm/UwLCX1LN9twdpLmb3viPVLTXAVCTWGnSrWGPo+fSfcI+48wlje4uMqGf7swaGQqfDcn
zDNzh7aLk2jGRf0zgln/mulhQwVadsGJgYDQmzpGbc4tZtYSdjYtk7m/R385AVbP30YjOAMw1Kcs
mxQwQEcBxiy/YPBpYRo8DMiKihd7Bk6mZ0DIwrcWumK7q942w09/mFlwl6FZQVf3IenxVuqxNREN
aYGUK82P8mJjlJSLCBXDqqP76SGvwVwEVOMAfZ2H7fn4DPE25MMVEEFGEBgJo0B1Hd6BGXibFxe4
7bLN0n45qN4QOX4FXCUNJ8FvUWwRbOQbKruJMm5jxB2kBJ2UDA2vjpCuxaLKRJ9AaF2+f7ZvHSEY
beFRCAtkFPd0wftA3pP5TcZXA8Itcd9LuY8DctIZoai5EvLEbEzZiZKr/KfDxhi2jXN/fYP7rc4u
LXcQYgFRGWeSshZxNwfJOV9sWblyn7enC3JAf7+ckfIijhY718rzC2GFVh5N/wIIsr7VgLl3g5D0
rrojXFdeuKuFWJgpL+QcGPBNzdWqHZb34NbMEF7GwI1izAZAkt47npqhmyZKS2bIfxiEitqx7Rk2
ZmMhTmh9YwT8YhAFlcANGS6SppG29y5ADeJ5/vGHhu8j11mXtDiiwRV/kqDdz3PfrTt42iFpoiE7
EzbxNBi847cHHSa/6UbLcWdgvav6ZcTy513begyPa6pJ/cM03eW4sR4dlaf8Pl9Upw2myV0+IhD7
dHHaYNSUr2dd5lZpAEDAcuTKTmeW0uniVSdZivs6oYYRJUEHVMz5kymfg1uJ/rAH9GgIq6VX5E/P
2iPOTtKT2yy4woEMIxpwUzaHR096DIJ/Wq/hEew+bMCcdLg1bGBJ8YPeLlaOWZ03lrFd6tDHiUKd
5AOb46NK1WV9dLGhCgrhVP0dS+qrHkwcmeZhlQWaMLdV0vI7yelEhjO7PzcYDMwxpKILiK+z/E5M
WG2BYf/YwZh4/Of/8TjRF/r0ONl5bGKKaxeozQEwFWWmYPFi96HB/r2t9OuVHe38USvUY8x8jF8c
KiB43icPrF82HHvD8BGDHrZeOoTDLQ8uwvNj/1bHPD0h81go6tAMc8/+LUXvsG4z7ZhP+z1zDE81
kGDSgtYR/SCv1MnDyLxQFTNrKotwFCzDcQYmbf1vDsETqOhXoHn5EDZUCfu9ljznDy/m3V3bQJNL
sfoDjAaxBmvYZ1jPowZK0rT5NXCFCDFw114UvyB5y6eU2Z9cdvbSAkR29aXyNxfU6mVWQNQUaCZk
rgkSyiTOso+U+Z9YdML7uje34JEtfHKKxgDB5All/U1Vnmi+qwZMepfRIvN/k5x9P7/g+1aKazmg
x/qddkij0dLSx5I9W0lFRNyaQfwEWWktOtD7FZdaRwk6Gu/CUYdaVh0/Gqxe13r1y4vQ6yen3K3X
ZelgKEcYkw5V4mLjJZ1b4xzm4AgAyF/s05iiPmC89pfk0oNCtgkssXNqm67K6/vjpC0uDYnFppxf
RdEpJiagh3LGWgBv2RKPhS5tFJP/ydlNy/pFtzD6VI/G3O/uDCa2wWz9xlrSVqxgo0BEyoGNAbE6
sWnnA3jOCoxwtV4pdpYyGWkolU4Yii8/yq2bTNd5yQCARBO6fxOvSLzOvis6sxWxMyh7hc0kUn+6
Tfi4plnXXsouGrYe4qEugl+PkbbKIlTCM3R6/D7y4cLcvODb0kcPKFVXM4wM92ldWAEoJ4O08vUR
nWJBxHh37pbeCfNbXcwS3koAjcr1VRip0GtAzpPrmCBkEnjp/Wq0zSh8EUhBzWQC4/qRbpeOLo+v
fycLO6MyR+FX22C0L2J9C7ObX6yQLWnJRHmBwhHLmTDmPfUvwEGB5xV11uAn8xJXC0N+JZNgflaZ
oztpuuSn3XBdQKwk5ccx60BPlLys4iZX6NH3GZ7KY55y4RZyvZXTVCbCNEatgnTg/QXEmbGC2yuS
dLCXhyHL0/bWbDo7i/8mO9O2NoYirE/vzV+vw1uvwmwkaQTTOV+jBCvrnjGXAHNSm7QuThfhqGt8
SVX23UlpFqSs8J5743jIA6YvWlvKhhscph+B3PMxZOOIlyJJb12H4HtE0Ne7rD+bZXOrIGLii38S
Uw7I2sCAzBmiScK3wal75Qo5u2hGa4zTV5a5YCJ5E51OIT1rOQXMwq0QZ8K2sK0tscfsgPxCNsI4
pQ21E6LK8DUtMCvl8SFqwVrST9WNs0mdVUBop7A9JBylEtRj46UOnzBSVuh/xZqNYPBCp0HpgXmV
MKkOI/oZxMqa8TdXRobr7Sfyg7GEtOd8Yl4BMNJ9xqrDCCG68ATIgRQo6dICzV1kNa7NNNnqTm21
jjkQwNxmAD8hsWh+u9MDc5TipESFPAXl49lnh+sQ/EkyV/JteYGGU5SaA9wtx3F10yiF+0LscdDb
ofeuDMBxsLe0jM7bOPS/8HLXopo4ucvFZExD2g4x9gUDRlLeK2QF4n8fRiYAj1ebheMiy3FrFXws
b3vHD7VhT9JD2xGPm7Wbxua1WomCM66Hez3FenIOAgzWG7wuhoaCGviw8YcN02JOLswYBDtca7OX
w+9SVw5qskhqgFv0ts077FneMqulTxzkEmmHSYXJu6+vLd421yV6SBxrWxWNyw/7DKoVby9ASLAJ
JHkrwr4cAxRc9X+yH2GNSDVTdwKdtNG7XPxthTYAk6vibdNm8zbdgXKY6aGp1dNRje0K1XTGQppv
l7JCK2CLHXa5t90U5yuMNmyycxJhfEBOezvtUFxS8Tjiz/T3AQN69S3cuNyfMTByrQuVVB0Zrqn5
ephY88ktuDTPw/bzsDEK07qL8FhjmAYwLBw87TAKP3nCOZycoCM7DojTaKJbA3XEAWhPnK9qRYM5
kgUPt4nikQaSutHSaVHYJWjC35IoCmAQfj/mDYv+WH8Y8uk/IWOt2y4tWwVURYlqL4an7EfnWT/J
L8TRI55p2OQWqd/kNgWZcAjnruPRG4k4au5ZWaJ5qB7HXxHizhBsZ4r4tMwJCQN2xdNzq9SV8SYv
XU3hdSXG7woFPt4xjKYYZetbtL4LgPNYDc3DUBPV+Sx34FAySuzr90xuujZnmKLMDNmrtMWcT/VZ
B0o7IA25S0gZOloZBeh9G82/IaJK04tEbnwzTMKJzP3cZKecRa8fZkz7hoLg1oah/81mdzXIdZOm
WnSNE8OLkER1TWkRj12ZAxefBjDgV5awWWltUcFPsFNdW/y19gVKwqF7+kqZ+rDbZYD827dxxuDy
gGa3utYkE7dbS/AMdcIR03nsNKzW0Jl/W8+FA7nj7tRRRZER/lOPF4KCjixkW4FkaRYEIIgjCq1o
ax7wesE+pxsLAqQP2f0l7fgoYqvvPVXSxCLafHEdGreUKVlvD6ARUHJZMmCi2BG/WeM+A3wTUhlb
ZTxfFO9VGab0LUrE9okmqWgW92wKxMuFJEnDAJ5VyjcEcGjSUH1O46w9oecKmmRmLjSvlwigv8Jm
QOoN2f4Ana6e4phuMgdmCjo03BsW83qEcio0Z9YWvUEgWnUWx6itR+bGOAvyzfeu/pIN56UTBAp2
Ij6kJHP+RT5H66ZSKrikXQ0fEtbU5KBmbBy081RID+yMASM6zh5IWxMpDrFZ78sDa7egoDtWCbNU
xct4Gu5TQE52uieIJRN1yXlqlDOtU4gP9lQyp9Yx96nlA8mHyrE8LwAl98ExzO7JRyLF5PsEB05J
HRFtPx/vRO2wQIH3aNtKy2IWQOeLiXTIvue38RmkzwpUtT0rdQdEaz66G062oiNcLr/iSyNIPRKR
Vx6KI1iSNu4ApZTNdxNS0Uu6v2VRQVxdViRHk1wRtKolW4Eir56uq1iPrppqnZ9e+YkGDT79CxUH
lZ9gCv8OYL6X5tEZ1CTG/5th/OodSmrasVEN7aoznuHkkl72ZlUWXQ56envr680Eg0JvZYTtMoQj
sR/5PDeztRz04Uc0RuHoiyVEL53qhQijtpCWnXIlAiWgrTbr0IESiQGwGyaXppaNou/TGlDFqxh8
WYOlZCP7RVJbl+WRX6THzvI1Aoy5JK3p4yUAbjDS54/phjEi+SS+lP5J9MWzP+vOGF2/M5tYM2P5
twUdrVSjKoauA2ItIyBV5CB98C7EQC6248rjBz6X+zq9YatXYEWgCsz0zEc9FDSiHuRyDoLlMMWY
gRDDXzdjQF08GpFbojrlNWiRRK5VWdxxrr3zUBV6oGh6d5Mym9590V7xDdVLN1eGcaKxdAnfvcNN
OVpaLr0NrLQ4PShEofKMxMU4NIWIrgAqX+FnChb6ygqTaMGloYz02f0RV7O8ck4JF37wH9v8A9lT
pdDbGzp6ulwgN91wqZuB51MYF7onaBaDlamfjADAQguCbzlMIWO8bzhocfejOFwZWpuQ1FnNoNb3
m3jl9SpimcVff7nhoJYAt7I9HCHuxXcXBrBryjfSRcBbunu7wS314evsS7kUph47doluQD4HSm6Q
kM/B+JaCpsdG7GrcdcipsvZWybKa1Py9asBo4Z/YvRYn3ciw8z6JFfvdcSbyEXl2khpu8UdGjG6W
o1aiqqtJE7PFaEPBiVsJedKpCeS7xRtSN3g0aT0IZl00tSfUAESGCQuOMpKD597uRuyMaf7YgvDh
RGZhA0/Jy8wGmJ9dWZT1jUo/o/jSzGxOZBUICe+INyDgsUVm/yb/vU047OQ78BdJwFQdi2yfXJU3
OpTdEn8CTVl/AAW+yKCPJUAJLoBqnK8DGYqZCNJ+iXdCDY47FVh9Z1hvm744J9BzCxMas25/xWjl
+Rupi9CCfMl+E6Mi3OFBmZt3x+DsBUgNIiQP51cJBGlxCN6zU27M0plV54cYeP7TZ1SWIXjGWWEP
RGF4eCm6Vd9FcbS1MwAbs2qRHcr286T4XH88dqj0LHtFU+iBldphrCZ+oA2SL7RIsICF3FAswbcR
7KoexvCETKGDIwEzczBAo5dWtMJqnYe8eG84Tv3mUdmFhZspuzA3OiH4+gndxF+PCg9BtsuFv7NU
hMrg2jRmeCztXWzOH0JU9Gfan2ncsUcJTwCO1oZRvKwhcUSGom7RqmdfO1EfTPa9mDfpkR4SKDbT
Twtu9akC8eTZ4xXiHzezZM4HcyjwsuFb8J166LhxxSdEILlhAsj9DVSEUpC1bC4mxzAuRFmzylba
NwPlvRSdNFbvCnk/9RR5R00Ov/Kfziov6wvCXBz5aTKbywt7oZPlJZWFKWAZaBTn/cmOxVllyqCS
C54Qts9eoPjTuyyhkXXrsLiFXxXrfXwaXFt6OMszig/dguZJnS6lW4LXEYPLqMZiCEZ2aEFqEjkq
nEsisiA33lxrX6anM0y5ZrtvCB3PVkE4NgbWhfXBPDgJbRRcETIrve5kvi9Y/XHuH+65+FPoe397
624jHnxsKj6bwnLLgWwGhShON6VwVMskuoCIR8ub65ml09uvtxRf9LYbK0GtRBC+hDDGtGTf2ANy
aFb44tM14DYySYutMzuM6xNdQPPqjfE+WCAW9A1WnLWvtrbkSSh6wGMaQb3vLYlTMfcRMrcD8ADL
N76ek6x4W4ZCZjIiIrzt5uFWLjIY2hwQWHWkFUjdFsiaWGwY5wvsAwGrtvfqbUHgYtqnoflyXUvF
NQVy3v/EmLeb7Aupcv3SpnLbNdkddHOWS+3FwdpoA/2S7dst8VsCL0yo3obd0mJvILX07/jc2FSh
2HMYrAZediTetZ2EpZqUq+PwtoC1RSx1VsZY5NVmKpZHE1y95UYZVTo01tSMN57Qj2Zc4xaytUZr
HoIBE0OJt/3KTLRjRrXu5oYYYlMZUwL7A6xD5MQ00RQdrACNjgKXNyyULvhuYeyh+5PJHzZch6Zn
7vC0Gcg2rCPHXlS/fR1HvRZU2+lfsFUeAJaml5hlW/+xjxycNGk/Uf7XfdIvRfCTFpOF4vAVYknw
SmrAyQiE6PPzgy/9/yjZOYT+pXM1hDJXy+IMImptevr99EqF6AuuWP5iYiSqMe9W6yFJGqTGDeGh
6LQB4DX3ejr+9QUxB8KhagsF5kYOJIO562lvTfch0vFiKUM+AaSlEOofJs+k61Srj3XJZlJ2I9kj
utLrjbVi1JwghxGJguED0fVlCjc8++sa6QtcGwnJLD7Ms8Hhjjip+lwt6N1P3Wls8HJjb6rkSEi9
DU6Yvgbffq/JW7awnX9nBfU1cn+xG+SBMbgfXKq0JkQ6TwgmuXwya163lEc9hYHpqp7KEjbsGkXi
ExTgQDmRrmSz5HjlYQUNMPZZebMriAsdy6jhtQQddbXKfQxNM9PIqArpBhL2MAg2l3O5EXsXuAWQ
eioUr2bw0NJhLZenLSBhSVRzNy7Z3NATMTi4GA9Mq8TgikX1UUNbCDIZOxf6Yr6Xl9hZU2GmAPPr
fkZkB/3G/PJDJmMSHzBTQVtgWzu/Xic0efUkzdLxRSLuHE/ue8RAC5I2lNGngRrhYZuDwRvAQ0+c
roC/bf2CTcXxhflKuHRMLpmI+EJU8tRRSAbRD1guMaKGUj4Yj0Kob/xLFDTgjSo4lsZKrtOrqeAD
Cwg/fK4vT+8YYPamjUEIxSxwryrPMG89p1NA9XoVlc1B9jd8MxlFt4chgpVQjHGaybemxE9f8ebz
Xfb3CcZy6Oza4o4SZHpr9wlnjbiHxg0Pm90MgyFKHOJp4+M6GZAKJe8dyYAZB1pMcCD2u5XiUiKF
irgswxQRMiexO5vY6RLd/tW149c6+iIN87XJEKR9QPIgQjqmLuJnTyPECVe6f00iLQk9kBpnBkXk
J4wzxI4AJ6z1viiLa8UxTCXPbHscFx6O0ZO1qrMrDKmcP5FskADlP+ULtYPaixFeO/Lpm7O7TBfa
arfhfRUoTH7g0lSVQEaMjwddUlD9EcPGw9gwcMXCiaWcrci9/Z4QYv2vllquzmkltwCOonT7xiqP
2433oXOInR0AWjv6R0X3pWnpO7ol3JaAyXLxw+x9FdXCrXe6yIU5CiiJ9AtBjs77LDAaRSafgpY5
gzVJjFLnPg/1aYWJDSUnIJQmZl+OFq1ONFe5G2SqyrEB5/PM3pHBoBcnsX+kPVBqCWR+cvkMN4NR
kRAz2Eno1tp0/98awi3hGx3D9b2DNOmiFAwiu6okJFmSKNGwn3GcgLj5O6GvyzH6uDf0EVhdDvQE
a3LCtZonTUVSQejTTkLNMM5BTNXO6TcYUi4CuNa3oFqiyeDNEPY7yI5Fl5lYygWvoRlO12vVbOAK
KSUSy2QiKDc2zdVjTQhpeEKx0WrS1ASuM3kbBGaWOegxZdLkN9bKDzdRvFP0zsA4Do0vjjoIsDC6
YmIqucdJBoIWrrhoZXTcRTHgh7kEz43z1ek43IrOC8uiq9qr5pC90W/VAvSao5b4T9fANsAvtWXh
EOKwNrnKv+4evUv4VpceXAUnbjqZ4IeAHECF21pW42bYRz+2ZVITvhlX08Rwf70nGMjmS6AmZWqn
XoWvcH3BycQO57ZosW1N5OBnCUxEP7nLgpNz+zhnnKS/p6hcf65NHQ0WHFs8N7AbQxWeVThXCiFQ
mdQvoLVLYjS0WMpSipEIDqazpJg3nSqH3Jb/kHj/7qasosbbMmZx1iK+GqLfP2UL7n7zSmiUsIIB
PJ0W+jiqOC+QyU1+jmZ2nyTOHKn2iY8ryIDM7IGDlrVgxyUQuWNZrJXjYTdPcskybVakSmFGQYFc
lmnJ/j+GCdm0ZoPqfYDLjVTSDcm/7qP6ghWx94CaACUoks9v2O5NDW7ggbdVgMZZbY/HUWMtOJ96
JGqsjG0rSkSeEJC1WrWWHJZdY9UETij8KGvf6RSWO8ipuCQMXbpWmVKGLflI+o8kOkinti52Ty3B
zEvsU65jPyoRnwM7UIWeM1TgkoYiFwG9g1KcGP740X9wVXaED+etxV0BTVDV6a523I0pbJqdE1BK
Hw0CAG1jby7TQuxoeJgPlc5mUShiIwPbcvBeS6ZaFoyAZZwK7aBzaXbdmucv3A38QC914mnMfvme
W5n1LJU/J0G++fkfmKDGq7YEWtSGm/SdCiSwTgHVF+B4jX2DUWW/DwcMirH1OvusKuh257wta8vt
dt8fUNRPFEGfI4mxSDCIQIiyY+OtyM9iVsQyXa+Ig2KlJJCEuR6GmFikcdXCBqfkKfA7NquQnuPO
IP7xVoWFjK72ZVnrsOpBaD/1R1CevlHvpEXGALVqlxJBiCVJxD5VKsKFjA7c+lMHMDc8yBXutEF9
YW5ryYB4sRMuVezwXoeBgsMcpCDaeZTzu1Bpt3427npWqMFyju7CHtuKWVBvJIJFdkghUQxn1XIq
imj9llONNDNlRzTV0lDYDSehZlI5+6IJcPzvyJGwYFIOFcj4o/EVZbLHtrjYdMf649uJsPjkj01v
XV0EexswhuursZZimvL/IY1XdbbGiGGJ7I4joQJaXB35aniIP1svDrkWilAtjR+gphtvByvbJ+UG
WltcN+byejUismLsjA0uwymrQx285emwZoNVP5qeyVOVhZ/nf9z2xamGeNkD4iYrgHqLOMGDqyz4
WjeAKgUC4MlpQztoEFtDt+3ilRJnC/Dpc9hLMZHq99qN2jP21Z+7R/7YUF+Em8xCyjKpoBcoQ+2h
MBEiqcdLsVQs8uIWBp/mQ4vizlZhZ/WEOM3tQiBlsICl4PBTmYgwqoDvV1rRaQ3RjknGk+4CTLjz
vgNnwSo4ryT5oGdRL6o5SFOhKgpvHS9NnDtk/wxNKJPawuAUaJsZ6C5k8i8clHmaNZxKBbsAZA58
68fHkfZ4d68Fan44JDfw5aDzmgwZlfwD5y79HSzLflVMWCshecZAeT0gV9Yx+EIs41z0+MaDgTZK
wdE4Zc/TjdAsWKHc1s8CbGBoiaaBaXsPgTWawVhRGfk7HvoLrXAsOIfrD/cmbb3Z/8NlN72eMwnP
PS/wDsPss7NVp3SfGAKA8jOFxZwhYYlL2SJwt/syaIBrs8tYO5T0k8xHa/M40rHfHIjpEekm4sXH
UO+WylvVvurPJGrMnpSY/l9ISlwfJkFLkVjEFwdzBVt57XhFfWeBFcUH9LaUW9txNm/5ykMrZlFy
SaZ0f3G/OQOuhHuAKtdAWamfzNEaZr+biSJjdPvsXmwMb/4QIgSo6y70bgnyJUyBHQmbVrwH9ApV
c52Oh7IQMMIV33B4gdDC3FYhet5Lu7hM85/SatDsnMldjThllZhm9h8xQHwVLQdmCKP1KdxghYpv
M/oo5x2rO5QJDcWVZAP27dhdQYCwVna+dl/HH3l18q1JabAtwtko/pbgIVFr4IGsxOpWw5pzR+3a
SkJvh+oKn70Anuc1Nb51PiaUyHMb4aGw0kI8116YwY/wmgFjSud0KuvKDmYH1Ypxf/2RelaROaBg
L/njXZ49Wz01tNpQwGBbPOD/nkjod0zsC0o360ibTM2xsnK7jnNXTR+1UkmVijpVL8u1ck1Qsox1
VS1TtZfwYHnYQOg7j/R9lp7gMyjxzDwy9HhQ6h8EgevAVLuqL23M9m/op9JoYf1sUApEJA/nlukb
xbakAKlm0uNnKVZ0bsGAQdaesftriM/xzuMtiqOnmId7bz1HaXgvgVh/nxOXvM9Bg8LwxFsVQb09
BaLh7Mne70Xsidu3U5yzqe/LYJF+97MiFjbIcmPhFW7E/ns8LXCjhBGw9kIY2/KeiJcoELRlT/N9
TPYxL7TR5Pd1rO44Hb9he4Xd/9rCvg2+0ORvL1FKuYKkvd5PyPPm2vmqNM7yCMSpl8f9P8q/Zuz3
5WIZXJbBV+gle8eRjwQJ3u9ZLg7zWsYqlEYMsfgoYS6cqczXKK303/v9CEeAAlE06NB4PFtES6Af
jXZV9XqslahvvG9KmYF2/F0SChPdkoua9DQHsWD2dMdQO5pnvnqdaXU1t1JJFWT+PayKdQ4NDC34
8uRID0HYEHMUW7GTzB7otKGgjlsGXAMIEY2wksjBIconWfL1rOB1fLK2ydfQMEq/A7dZh+GEJo/9
PJ4mmw5532KXALo4Axpjr2R5FZ+eC8nkjSPJiYRzEpl0yZg84wzKlu2dZJuSkKfxO1mcpQ7DK4dd
9nB6jSz3blPDHzxl93M2n1Tc+APQJB8daQyiv8HqOtHYhJvEaSQWE3hVbNpAHsIUEuoN5e8vQhEq
kpSYdrwEqJV/Y3yxMzEW9nuBSgZGoNGWz9myMm/kWFE0OFv3hJNOKU1qyDVPt8eSg971yeCup/66
cvb62Ip7w8cq+fvgSzim1zS4pIcESUM5+1CulV6Sff97VBPF9xITkY2LaY0qR97yugU5uXADNjAw
+xwXt5mQ+pPaddLwwm42rXa3JLdmSZU55xMAvWf2TtuZmXgkU3Hb16wT1mbAAgHb3AceFAGvUQ9u
VyHge372W0TAuSGu01e7W1GxrovZg58xRka6TNLuqegfXPohtL8lhA25cXuyeYe+hJ/mMNqDLT4+
ZGxB0rMeTinOhMSBHcSJH2Ygsz81YLjGwmd535zwL16BjUn/uUQ5khk3KInHolQ/nLwDRydqmUMI
W/7R1p3ZYU+KHTlTjNWBmT/Qf5zgE/SMDS8f3bWBJTku06kYdz8WAeXA3OOXbTCYZkFKvyxKlhjK
3JbEk4Fx60b3MQbOsOHpuLTG+svuvqkXgNR35ouVIk3KGJiXJgBX4K6GpBdRyYYAR5nT+VkhohIt
lpJrT3WJyNhdHmKPHf3kmMpRzs69mzE9BuyKjYjiuoYQgR2FtIdCUrwT6PBYQTFECCnuGj/n5DJU
pOHjhP4n989JcluWh6TsJhpwtMpLDX4CmLMvhJiuk4oeXArFJz5RKVEhkNmULGlQt9UDGljkqH9G
SL3mpDlI+JkLkaZRiMncrUzlqXKrLoJQSnBKSKwxER09dYi36klsXn+BJTcEKKDFq2hZ+QN7sALw
rraqe3OA19iODjgrIZRZdMYAYd5/wXW67yTJau+oJGe5DGK1yj9nv5KVdkqG3pX5ew+Snz0xDzr6
y12aKXCVJt6I4z0/fMZLzA63gMKdm+rVLDjrNsbubch2P1QLxVBkbbOC/bARUh8x8/2PCpOlPvn5
4v+nRp3NjXDp8fm7oZYR+OIZl+O/+eYC+0s9dwTGcLtjQ1zcR5HElZnoI5ru/PGvD30UyO3eH3gS
x6z2NtIX87aTh494Vb2AXOvdlggqhdMXY/kj7/S1Zz0dVwj9LYAILuzw7UJc68q7i/XVsDO0M7SK
pQJX/k1mePSN8jH702/RyYcwIufuYfFut5HQf7BVM03uAYxyB/YBR/bVeu/y0ma/kSlp/EBkyF86
pBhu6ikINzeZHsEPpSzrX1TnrjZHtJ21J2pdnNko8bOmG+S3fLnaEIfMb8TGkDKrgT814+vDnGY6
Ifr8WBSjtOghOC0MogLFCN+xAyEk2gdOMyroKkhuEts3AJkECLbWmaN0L3igDpn1PJl6WQCdKl6R
Dr1Ya9BYZ0xRFQtJNHRAepBfjOJa8ayh24ZUdmTu9tVUDYcgQUqk6XgZjtSncjYDaEppdyIYLoD9
LP/rA0MdWs4NMPZ6JVDIkNhZvE4duewgNPM5L5CAuZWsaVZDImE9r3p9mCMlJFWdd8ae/uvCeiWR
IB4y+C5woW0Nela9Ne/Q4a/LrqLZVxuooN2ZfXYpj6z9i1M8JFEOrsbv1PKqC0pVk/COauG/dr4E
YtPfDtwJYpIpLYc67QE6TdjKfJXMlTWExUZlwbeiU7ad6Kg+eLtXp6RTciAJhsQyVRS3C7O5geX2
6TVAF4U1sweR30oXJbvqYVR9zLPnulJtxC+nSuX2pYrPMHI9WcszkpNhuiX+YqMD+sT/kMjgmXX6
H6bnY8hJ7RTIM3zJTVSEXLhKn38qRwcy7SpXHBqfdsgNK047vna5sh/Kw+wBtaU++rQPtmIXBWXp
mhb+vr4R2rAObu5LxijHf5J5GXLawci2THCaYj72kXAP+3ECMZljOU7cWzk14goEtODgk+pKSMS3
9beA+ysRRZCZrDB14jhOhq0BCR/+aEkfPEbMCMY3LDfjkrudf7Q1J3+1lgoUxGPvsSfuz6K3Ccvf
DJymcHJ/subOiUEe5MfrOg0MkOGA4c0Ucf1av9P8tMldREsH8KHY9nvbB8WtIsz4mYEKBoLg2loV
/C8L35O+xI6YBZgz3DBQM2FHKfDmKCbFly34LMQu6WjmE2/JiK+CxOiJbBcCWk551PtwXbYBSjSK
mhGpZah+L50SxSA4tnGgvNrkaiYWcv0YYcAiaiTbLJslIDW3q1UEbHWdOBx3W7rGYN+LMORMjEfG
5GwbZen4nQ59ap2guKBUenNKQoP+UbGZyQ9mBvytMVsYctimZH+HPGiXhuHdl1vqxNnTY3YQi1QB
ROD/8dTuy0mMdaZZbQaop12Esttalbrusw8BSg/CxcfzkCq+bbu0D/j37CkiHtBZsnUfZ3V6xyb1
cUoQkSTBF1Xt7A+iAFi71tNyxdbt1XLka7BACEkqgpNYz0MTQD9Jr/TFaKt3gr7dzozQ8u8q+PSm
zxi51djTgMHa/RT90jGMVM9HOM8MiqUQObZluVGhqv/+HLL/QcGRPdW4zARaiQVaGF9TPz2PkhZb
2jBcH1JESFl4eGA7HsKhwKxXv47Q4QIWpTYP2IzeHYtSWDNAhvh9865hK2ysRSWzHC2OE03g5DKo
9sQb1F//CwtPrrMow+E3fovTCAMlm5XOfhQguM8QwhDJLJflzzkguKzoKgOvDRp6OTMSkG9xeyN7
IVobqM9f2xf+O3ORgOferjfZP1vc6AWIhMnbSCKCjp1TZp8aIZP/0W5xVkN0cZ9TjfoIDW3UM6pV
piX4dk3aS6bAC81SRqiyPK4vyTCN2wZLE3JI0CDQGujjzojdUxrZoAjbOgTXPMrTeTMxL08d70eC
KWGP2MvAZeOoq7SZLmjf5yNrJ0A2Dg9yKff4QYypcs8vJyD24c7Tl5tam58CLWhP7/wARBfXplMi
eESWZoUAhUWbut5S7fQ3OqBSguRMf/0oq3sdhJSj+26eM8FJqjukpfrggE6wzAmjCYNJnXyy6a+r
xPyisnex6V9SetCBhjBYzc+l6lh28OpITM7xiyRYhUN46J7Fa4UWRp4/wguJRvUdNoCSBWgRB1I6
wTSDTw+3CdKeKHHGu2a12heunn14jOuJb5yzJk5qnUZjLxNCnuJJG1Ph9P857w73uYVeTGCP3mfB
ZS/0CMJg/gczA/tA0DmvYx+8vMwz0tRpjQoClx2VdnSx4BkhaqbUidcUPz7acsyf7fsMz/CyQ5Qg
CQNBDNoM3ehZuSj/cDlBv/LmlF6EI1n3+NI4UZEW9p1+atF/01Z8K4u9Fz5JW+SXh18Gl5Kg0Hfy
WBkLg+fTCNBlRPpuonO7RKS4C/zmEovlMQSx7ms1KRPcGuV3Vozq1p8mltqXYj3Rg5WYm+cUoftl
Jwt8OaFBqZDY3ABWyjCFFhaRtU+cImjfS7ws9bw+PNFRIFceywGU34BMkudCYRITZSy/X3qK02OK
4YYF6hRhpfCNiJoWrmQ/ezySHUe6W5wJQBKoUttYpnT0Q0BEH5/0e8CuJksYCC8EoTf4qfvyg4Uk
cp8PMEuIHPtiAHwobFpOOSIyDEz0NUVJTYr2mGMrMAOoEldO2fbAUypPa6pwxGP9qyNYqT8uhEX9
UHInyAXASRYhxca5LpWBgyVW8oyZ3Mhn4mlbDo12PIlnzCiC73Y14NVK6C1a0B48T7P4yyqo1jln
roAAyk5XT0IIizz6TUdwAjMpeXxlx8ws3xCsWoWzjVsQ1d438CmbDO3ZFY0xI7E1jC/pHv0NjQ5k
DRcMaVMWfTivp4H3wiLCgUOJykTXLAYkq21rfNLe3KB3DcPwsDXhSzU4Tfdipntekoxv/PRSQBzz
DGqdQCVs1nmycVGq4J8ja9nlj/njjnMrlqMZw+3TdHeqEyX9IOxqodBiX0oWG3JwLettfSVv3q5b
aroluQUPqZent060ApyAvQacO2U2yYO8GjrXzl6VDkA7F+sfEx50BgJ3Pz2pZ3z/+36CqN/y/Ve/
bYAuLGArUSFzYC+nyotz+0sbr0S0EUIK6ouNhBp6JL1JE3I6Esf+4/ZpwkfgEIuXRG9WR4n+z5j5
kU8MipCgG5F11Kxyhvlut9fHC3dsq76vM0fksoewVm93q7iY9X/4gGTf26dZcpSWwt7QPH6BQ6TY
hf30zqs8vS3pT8qfYKmUL4pUWWup5zYFP5hsHSYCX4i/giiFYis3rW0lnXJtanOO2ZZP6TPfcHPD
/FdJTA+kKf3c9/qhz8LBDQ90Aqt2UZKLv95aKV4kkoyGfUdF9dBCdchoh8Jl+ebLrd8UQDpqNgBH
oVJiQWBDkxtCBBlJ88tdU7Z02C7YxfFEEOKbsHDIvjs9gfQytziweyUBcXAeLdK4WYhtru2DIjHh
vbBEo278lKAIyMq21tNob4F1bBqvC0awJhdy6PhiDyk8cW+kfx6PgrIVh8z63ebGkGRhTdtrXBQC
L5ue/HC3yhhdOjUYD9CwE+p2qdxvYyfHFGbY5F+wx1ULDuoy3lLs83Wzxii+QLt5A4Pz4KahFn1E
PtewkYAPDGW/YY/PZ/S36ykjT8lwOt4S8GRm/N7C7cV6L6Da1XA9sf/WUVB+LmwXRC4tE0SJEkDr
nvROMsPYu5BJFDQRRBuaBWXE+4gYPukItyCNFDQjDmolNM8wPA7FsGdOY0plKxXBRGNapKLkN8Cp
t/7leqHBMIPmYntpNDx3roEeFtEgyGl0pFC4mmCUt12HP/VEGJGVUH4guLwQ126IQvdoqaEOLy3L
1R+n1loiPPZtvkJSOSpqFr+uufLvCuNoiaOI9NQll3aRaY154qyeoMl1CqRCnC0NBu+6UROeeKHr
KCyZQ8lT3R4SI7e1/Dtuf+c1ikFp00SS86MPgfUVDsH7rFT6oxAh0xVSdagA7ZP3NZXpXcBQEIFT
Q9GfQEW7zAF4Ut4W/vPCUyHKXyE+xXiVMNvhjMJmTu9mks1iEL4RUt5hYbEqYCp0OnHK7e9Zjiu3
j+W6ACHxiD/cvhSBdquKlVCR5uZwjmWMQ0P7HShhY3PXkwr4KCCtDr6mph33KeCZjT8nR0c2D5dP
IF4ToTLK20vrJ8M0dreURy8lj/n2HH/PykoHa27OnbBDsBb1kcgxoCOx3N/w+RKG9A439e2BI3J+
FQONcq5z30oyE+sQQaWDExEw9s8hKb1HMYNXSN5ewFHSw6kmY2u1IBfqF9fsle/TdlaDBqIrzVvu
P3UU9AdSsSMnn+38sj/QfL2HI8pCCAOuOXiqW8lBPKsrHJTbwQvofgLXcJ5vXnZc9Kcuz8K6T1ij
trF7bAltVVQzAaKgYApXP+bckA08nawOFjFUaE823doYpd1BWR8b9VG2QDbKC/DqiiSwh/r76R2D
TeqymasHuaapR3btTJNmoOKrcfBOIyBq8XesNLWW6PqcQkC3jrGa1XLNzdNUBJX6Ime6QVBVRICG
uj1LisJf9csdIMQsE7VZtx/KW92fp7pjCTS29XgfidlBHZq2Q3IfbaN22im3UjMuCX0RqNeZLrLw
MPdWkjDQv/3G1SxxeOoaNp53I50C3NvvpD32oSnk7Yt3J38Ucno8X4Dhj0J8EbgPTpP5co+YWqum
FUAx3o0m1PNzAaPljptCR+Bsfy64OOxbPWRA+d42Jl0BHN6j0cCe/ouTuLE34fOSLm+Nmf+os2RK
Ncv0g46RBwr5KKVmkSUtM5Tgo06YkgC3SV8Zb0UvQzKtjPu7IN3A2qvzYuI/5ML40MGzky/5Hzu4
oCoZHfKLB62LfodLE7vrBxEnxjy0hGjuf9lZx2ExKt4OITHSZEdxVaWvRAGI1e3LiF/g+KRs4xul
Q8RV+6rlV5i8vtEVaT94uNEDB6eAPERiZAu6H1fmDNaNVqMo+dHQuFIaYqNeCj/pqwFbshfO/Ov4
tU7wf7505UEuttsLg2eTF+R9X87IFQCJnhPd9WFYeBxmsF1xWdPIxCMl34Vul8qcHEKVITeO8VjK
Na4f5g5ozgFhqza1UrtHHLdRV7OgkJw5QahCOPwcofJvNoMgPZ7Pt1kE32EB0csBhZYDVgEmUrCy
wSo9A0ePkWMLeMgX6D/2Wq+Vmwwtr4SppNZT/qQ+Ip+Ats8q1BjExc9eB+RiUYUvYsAAI6OL2QzZ
/m2+aQvRibd0KVkgUeHiQKxNnEnwoi+Ro/UMjhQ3Vidoh1PDnVAPwmhB+vV+m8lo9ad1y8gyT2d+
PQpcGe1Jam2HDDlTQ2MXXmtK4/3xhYRNXaF5eBELqpAn8rMIzBzBm4S0cNh+uVPqiKr7kHn/HrRd
qSwdjpk+EeB82DASFiJ5o8sJBs0WJ+BffuAEDXrYMowmu5/U59bFDYn/sZnuiFbyhCsg8v62NZa5
qv97mQQT+p5Xy0QpTNP3HBfoQmQEu5ejPqKTDrLsHxTiW1p0UyHZLq6Q1xnoqV2VzQ4xynIdcds0
1W/xJHZnxdG+VfYTSwJcLxo1S19m4+yWD8brVqYmtp3fOS5jhl9U2jh2QF6ET0W7iOkZkJfFj3C3
KHW1KejrSOXotuHGg1s5s3Rp70q2G1pcyj7kAIYx9bpBgbKeRebJq6EHdp/IjtcQxfhxxkxYHqT1
ilDl74HzhKhXs6b/80/oFHbNUHg5zRXY6xonHoIp+PjTF6eK5+7mP6iMkLAEZkJwHSpng0/NQbBt
/sddcnhjOYPUGSuMzNIAMf2/QaYCciuiGs69s7wHl/cGO+VjpmzLmOCcvtYN7XedGYsFNJTpBkrS
DbhHABhHWAMDd2jIbj6W5pnwNmaTq8KjUBrLyLKvV+uEqYTkgkc4YzwIQHyBpnsONJQsRf98cIQx
MqLVt+8SvOhbde7lUCWYhZZNWQoXIrBpBRpJbEx6YZqaQ9RTRvSZABi2dghAl+xrzqlOH3wDYZIX
iD+d/uOA9Z0cPV7viYd3J0fT8YbNp2AjQZ9frZuLIbtoEOj9eguRjqpp2EJmCCgUYt4JCPBEzY2+
7gAjoIhZ85eLJafPGMNpfDiFGPWdSWVTU6zA6w1W3ptyzEQxgMstbQs1fzwrrzvVmDltP974cIX7
Ahsr72feBdwIt39Nv6e2VhxVxSsUJgVb4G7ABbQuIKgoYqUXwSCp4yxUglUoTSTGRfv//A7Qx9WX
rvg5PEIdO14bwtTQeewa94+nfA0pTA8AxnkhLnngbpwLBCDO//2Mylw7KmAHE0aPvR2nWr3LekBN
ZSP1rzz0pjpnkRJtgnZALDzEnxfaw5Zl4omA2eQfbxR3xppEFa2l/WF+JIMazN40L6fHBOaWm7ua
WHudgtsOemv8tKIHgKscOO6BFNcWDVyY+4vu+tr3MHyldJic2EBFDN8OaqM4J9+mitErTnVGZHFt
3pgdlNBQEzENYVaGkGXX1Qpn8smWAU3TbiePOJqNSqm7N2rW88M/b2ou5BlsMS9H+jHb+S9/FhLL
jWZbLkAMXqkkJyLUKDJINVaXYCnakn8curjVuHqSpld6cl2wA9v7B5lo2TfZ3wPiPc2yPgUfL2GY
zNskcR36JrRsKovdj/uni+I0mwKnCmNgjlcrMljQgtgArZA+wipwGQOdfVRqW7lsSbC32IkfreV6
yyFv37P9tC68/yumuafREfe5pFa665EzNiudUqfYJg1xvlMyYupbQlbQsV9DqXBFOQvTHaA09tNG
d3Sjvh4KAPNZAkQq4eZhs52LiLRfQOyvvwrk50l5RmPy4lRkLgSd5UuQnM62qmL+lyGfvEksUdwo
FESKWQAlXQkgFcE3D1qZaVgA68C88QwotnH+ctaw1dDpOo2qUMppO3HPnUYOMprab8f42OcZm+QY
pBKCdA6+IvLnDnFU+TXF/8cNexLaI0SUViqNHICjTNtXhg2Zpy5xWLGVKrlmgauwyQNh2ykZrSLw
PAjj+Z6M9qX5mOE3AEx4biZ7XEufRAFcjDwJacH6VO4hty+7AdHFxLeFEg14iLRbEEUfUMSMIgdf
QvKlqyEHTcmrbMWVmrR7NgAMdPb0zisaWCI5MnZzrQHcoO+mDf5IH9vlsBIjm3svpohG6DlnZj6X
bvfJOjpCGTHqiGce70PJHzaQKsbx4bdRvpLT/7pC17siNBPd4ZDeKsWcLPFie7CgItNifZvhmFFb
zcoW1/UP6xt0g8ockvozImZ+RRpg2M2I/AeT7CSiitVldM84h7uQHBJwpkcBKDGARWVscu9VMgVa
ER5LMAdKgYFBSSJ9tbwTyC+DcbrOWOjaw0NRN7ijinak8xXpLExsVBzSz2XdIUMUpD8KESnfYbRS
rw5966C3lok4jUoIfOH9Mry93wLQW2cSy6cjT9mGTzmc18TsYiengCEDAf2uajqlqMldmtJXMcKf
8ptLN9ogoTbQvK6UclpK2hiUTsZy2yQveNgdb2QxPNgTIPUj2MkNakwaccgwyGJVaDxO54gkkSCF
GHkfd0h4EwQ9zb2FaH4CFFn0NdcPNI4GIrADJrjy6I09MO0bkl3XFlEpj+oRarZ4w6v1gmH9sPE0
kKJUj4OY0+oPTRYKkJsv7bDuBZeV5F8R/RnjDXStEFma9cBsP6DlsgShNDuvirdud24DlEder3Hq
mI5OO4htVkkWpwD5pMeZ8dejbrSApMRpVRbE4eZGi8BvaDvh9ISEthJLfmX4rYMgPIT633VSXZYp
FdgqOM84UpMYPGZr88XSHAJ2MKEgBQb3RxcZ1XOKTmRrxhz08vBEWbvc6/be8IuzRkATtuacJCzI
uJavJOS5t8k3f8AUA7iE90fKqhF4O5A9lrrSk23QPsroIp8io/MlMuQ9Os8zevNWSRtMYhvG7G0d
aBSXnw77dm63F2On67Q9RZUcsXIMwcYkRbmDge9OqzPsFWb9rb8aIQACXV/XyKDzSC/fmkZXzxax
vZDDW/3wc70NEUzfl0B1qBGuobFWHjTiQiwQcb4nB8rWghE9kA0QSU0JVII0cBRl0kBKip+lQL6P
rIwHJQeNcyL8HKirktkMTbxnQtFtj6KIQnt0kpk3LO7M3Zzcqh9dCyY2EdStvRf4AG76yTQP4QBh
3UL10wBqlytALa9NiVfDAdDrhr9uaP5sya9z16tFIWSlvuXPdHvWKOMkgy1EOXgxQ/lfjyQKK+qw
JpNJXbuUc8/AHkjzVtdEyoPjuEnn1448mYX30MaYpFDhsLbV2+coeEZgf+4upTvopksLssFrpkty
E47vgm0I8D8Jwsd1QSpgfVUAZ6sy8p/PxZpV3OXR6uKKr4mqf/Cluap1ANQ+++KByI/mHxA7pWGV
xy8tK59up+FcCanrpu9H9V1JkjCeK/ITBWm6mwbKPvwYKg3sZPz37Rh2fnRC46L050AlspPOdaHd
Kr1EFVlcqgen7k6rCXdW5vnjQEu8r4WQFP5Wfo7Cqkx831I1YA7yroUrece+JybA9fTwaDGnSU+D
vf0SpG9AANuPbvRnY5ehWoLB6y2OQPO1oaYnO11lvtx9Y/v1ZWuKUHZCMbFoGW+08+wygK3t7AlN
dTKuTT77e9W9cgub++M2dW0KEwS8/fL8ElQG4fKuP/yaVL31TcpoAYA1bGP1ghxJuISctXGgKJ7T
cc8nCPvjsu1/bw3qBe1HNY3lW/Dc9ZjmFc000mziU8rhq+GOpwWEEuqaCk3NZKav3awQrUuCtdCU
V0TDQ1g+xlKW/oe7Wr8mkTboxlH1XabVfDo/8u/EnIjUpB/ZiDZkOEq5XIWmXmo/zi2pU2DPHApp
y2pbgsuRhR3Hi/CiiM2IgnHXCrfghyT3gG/lZRL5WDOPDp/vohVM2kOd/Fjpwkn1TjoIw3K96JVJ
WBvnMFbf6M42Zn79yrH3sMKJl4ERYY5LAVb8owCvh3YQtCj+6t9vEUyM2SdMkKtCT/iZRZ/z4gVN
NRp7oZtz45C6OdP9IwclCULxMAeEROkSNJwELCjEnHg7OCgegfSp3SegyyJtMQgSpeyjFIU7KEYj
7IGKQ0NSJshssTnglOPhLVvAMajO0QM8t0I2OWUlGLPH9m9OO0b2FUksp6UUoUHdhcmwp8NQymP+
ZVtL0ZW38gu3NXWatZx+gFrQ6smX64kvg2Zh6HwRUp3QUUUr4bFhfq10RgK9sDVqskbmArKfQgd3
LtT+TeefM1onTQ74El/FZas8erqZ09HC+JhrZhhDznG9QNEkI8mmVCMvgYMouHymwOlwjDJfj02C
0ZGefy6jXnwW0m1zjxCaqoRLdsTDWzIWyiO1N2Fjp5cFHJFxGmoPOoAHMQomnuuWPTbEY3vuaZfl
KEsSs3X5hDGlzzuR7CoXAoAEfvJSQJjlaOx35WGUjuQc8UKF5WNij2/crQs7tEKkhSqVCnXWZwPG
h+vqTutX9cMoJgpell7GvyFBPckP0zWhgbBaL7P3m3GoXuWuQQQVYW49nVjhnPaVYbt4Rc3tOHA9
2/4viQSiabV9RfmIKT+bjxYXU0SpqKF4xe2Q2K5bu3T+GlrxKHGMznjIHQmXXKoApu+Npr9pjjFV
uF8xjIpoeUFwoGWRVL/ZHtOz74vQ8WXNB+D54TL7KqqVOD5+r/Q4Jae/LWf7STUhMtMKK8SEp0WS
kNeDOkIDHNNFDAVwfw+wUDAboj1OYQ6K17fVBg7nXJin4VyvXfAYH2rXMyeJ4286WqgiZgIUC1kY
FVUavCO9whiWxLTNag0Ay7FWyb7pmylhnu9OMx30tuO2HfV6mx1NZkckL63MMP4dKnuPKFg/EaNP
X+lJYvP9fve9VpHx8ma5mncFus2F4F/HIu8ezeoK2WWmHkGKQlEvsFXk7PjbXdk/HVn4MarBqwJS
tzfg6vRK4JoTty6pAZm8BUiFrnYjxMkbFbz0l2lSGVT04//llyn6BnHleRHGt++5ngxYHpzQ4nhH
48ZIDGNeXIp5HDtmHzxjbswTzzY9eSa+V0WaIZNQ6zUiUzJvXu/s2k+NCorh8P79vVy6feyUr1Oj
PZ7piFALFH7Cgp5HzlX8p1rpLHMxfn8zXuPH8Bm9v4jjjTIwMTwGReFzXIsX77RM0dvOxi3HFNgK
djXp6xmfFEJA7NxpXwFruitoqOAWUKsdHwEZz1VzOz2BzUJ2pSb6Qp1cZNivAZ1M2aCMTOwglkiz
hUzoGeQXVGsvGJSwxp5QPT2haSYnvAfr+Lltt1+M9xyDnS3NPTeKRPCObiQyrYgdQ4aNjJG31jzO
b/ReLcMfQ1/67j0IiYRAORiYM1I2EtgCgSB4snSqajSf4isnKctDLXHk9MeUyhfHPS1oTywag4Iq
1kNBz7VQiFqSYqXedx5+9mA1gmXHu70MDGG2sEAuOsEhUH4LaSSOQGrH5xvEn5J2bLwyZAF8YGER
eFQ2eNAKeNue0qwEzZeg4Y04PMF8SlukEF33ltaga09a0klBU4g6I0LeDyaD0WD77mEZN9VTyLUe
lC2MHbt1XK6HaKftT/q4cSqIFJnW16ikzAe5YNgjxDhRjgbeqDPvShMAXzVrx6Df34OrLZL4WXCi
y5BamJH3vWiouO2xOv4YwOBpPFGUdzRhStHejF7GyFjEuUFxKmFUhOvguUSeeqL4qN+kQ6l6ivMd
7qJ40rdnslrtpnXD2Sku/OMw3txIcNKfDu7X5lUstrON9SKL2mqKfp6IX7iNYYBmK8lJrTMH/Wsf
IXi/ve4aFAoMQEa0lKayRVZg/8K2/BaxM9VWi+gg+Vd98+LJ1z4D0k1hxKQ2WonbCAY4PER+xrJv
3TyxvW64Qhe8+ftRUCQoWAb56w5ZcxMI8Jt6joD9sDVvsG9JkhDK0znE5SGbyPGwgbtiVPh3r4Zy
pLTi8PzQ9aKsKiGWxTewW1/gFrRNOws/x6zU1yyqFLNzd6lWVjAVrwX7HuRkfT/NaEjJbiFRclN8
AzFrzXnRKf8O7/7HLnY+gIk2jtJ7Ok9J9+PCZcv6GUSuBLmEwWEium54Lvma+OnXBeSgenL6XIB9
31mtXSHGKVM6QtP6fhYWmbrl9l8+8ia5h02a7zl1Wrg808/3qFANP7jfpsRjcSvYWxWFr3MICn8Z
EMkJPbR40ctLxcnCAseY5BAL/W/gIVABMhxqIHtEuu/QwOyaztTrsosA/mDQMusuEWF7Dxp/NYcA
5NcCVS7uujfv1pAXF46Yu3JEGl+OnMQz2z1N0mGxQ+4OH8nGWo22GmfHkmOZEmBoKxWDAYIdCn6p
vxWhuqI5mp7lRxzfAdQc+hd+l2+RDP2+awjUBUdaRZl/T64rORdvDyCvU+9AjZsz0ZLMNHQFEpAz
5wJ64TWy3c15O4HywzD1YXCy97WAwCc12jPAYEDzfc4jvP7R2efJ0YlxEcdMEAG7MFp0N5XO7pJ6
hkscpTqBXmg2kKOOrPbSG34tsninMh3KZkqGbq1pd8CR5905cJT8ZsPS7jyZxrYoEXCJTlxWav59
7IpskEXkURpse3WmWuf58ddaVR9oSIFEbqZT49FLOYHEuInOkAOh+6REBAlNKmeNJCI/eDC2X7zj
yJdBcjSUzLbj8gr8UGn7sken1+uAQtH17ioYKNEXrq81CsiZDSLEgjgZm5GRyR1TY9p8/dQ+5RGp
OR2KEwT775OwoZ4jLPgTwQE4WY6vlT7xNBdYRYqvT+3syTTEfrbGeXr/x1eJLPQyhvciVbsSjlVN
PG6qaFRwiShX4ZZ5GnEhVmZDl5DUIJyvA7B8H0kgE3c1oWUJvrevcTsDbX9Fi9FvN/wesLWP2ESe
6f3UmZTiPCTuzWATdyyq67IgHK7fktS746xIGqUeJw+mOsJYPBhS1WtEXoKAD28Yam7JHYL/tvRf
4POeFDJTNLOxeIeH0OEloR9VAiok34v38iv+BFFTUUqe/euL+exm5PIIWPU2Dw612HkRp4uTZL6A
zQxdK7lX8BNJZ1YUl6YgKA3TRNqr6KmXzbgktVblaQ1XN4ATfWUfov9wqSoaVZLUcnwlovEqXkyF
evRtvWwVgb9mbnkfyblLPmIG3NSOsz79H8SUS8STeOWJvKnmv1fSs52U8lha/NVB9oeLGR7KxCET
OyUeiuS+Hee/6F6vA/XIqDXYKo/mCqNSfhBBWN0+V0GjY0pRC1UQ9T9B83E8CARx3VoRf/Qkzj/L
q1H0JLdYj+Qq0MzRkyfXz1IQBMenZJjFNpr+fNo5XLdMY2nQXeb5IbKTKB438ShWO4JcnMz/dSia
lCj1076VwT5zE82qvNIs1d4GIqsXfajxK9pT/7Sw5/ZaiQHRpRw3pX5N5BLwAEpn1UX2nzvOuGql
AghB+Dk1DqVIqsHoOMjXJrd/eC9Kb09C+KSe5PrecLT4F4JbgeUoVhlR9Yb88iHOxA+2+QyH/98D
9wyg47sFrzHLH0ByueYpDQHQInSgCMIE+Pc9Q/93VGqIk9PUHD2S3A6A+79LOdztFFUkBSKykmKH
Y8bU3rGnib2fBxlHySViz0aa5Xqfe4Zt58oHfQJxnI/yP5RzdA4+YYv8fGHDDcsaHWcUtbkQYjUP
ef0Yw4026fRkBmIEsy9Cf377qQY2VP+rhrhpvrjnZYx1mb1DNGLZjNp4A4mGpZ+rFNiYrXNdoSFO
m1H3MEYQFcZ/FtDAmgxlU3S07rHso4insSBYN3SQLaqd09B49KkAV1XQNfvPqmPqqV/yAh9QRtAq
CV2Z/jgz1rymqj2f1u5bxffskCtCjEgRihitbGJ1D2B2wGEK2LnMtttKfnuNgzpqgktfo6cJClKa
583Fs1UA/+g8n67JWde7zRu1r+zcdUlOgQUXPiqTobNUXX6NKsOpFc7SOJA+fjReWxOnPDMdUiVZ
/GL2xJOH0q9ve/j+GCjHYPTO2eW/CIweq3KiZ+OXICgVoqXcLh8YShQZBh1ydj+ogZz+/cVBWEwG
umfoFx6kSB0kudj59e5G4U2/Cl691IdftetjNnFFEJ5m9ST3WpvZj+QCDUIC7a7HInKf5buqydiM
m5PksJgCQdv36+Kz4y0iaoO/cHQCB2FJIFYJ5coVfO9Y/bNC26z6/qCyy+crbQji0H4GZsfRmvZQ
LXuYDsdNzuxsDIGC9aYmz8n3ITdxNYjp6E48AJAYr16C+6Y7B55BZ/VxL87phn/fmcXZupnNzvx+
Gl14tMqHFS3Pv2WB/Oywnv5ziWAUxj0FHiHSRGYlXw+c9ERyukPNXYOx5uKfmJvLEhF48lIVkSE+
rFOkEIj352uQu5Tx59Oc/FkMRvL3kUKREGqM6uFJXdCSF6Zy7z+uuV6JuyQPixsPMwv95GwE/vxc
p82FxaeKg3VbLGfDhar2hvk3xCa5KJxdFq0zVv/NjCSLWA3c5xRKNQM9uqsvgAy8Tj/bJMpAVW4e
Ij3ps950S7m5D3HIBaoOGBeJ13WXSuEw0WCQz6EeA/qvY59eE5jHCAiPus2tNw/9yebVG7ZJbSzJ
Wb9Zbo94GUqkDYBTV9a6n3ZpgU1OCwUrSwdqMTJ70t8zPJKDqbeBwynPH3OLAQBCl6oo+TbtUIWb
FiFAjkx+cXZ6U5T54WZOU4GoZiRddvVN8Ray6Xia7nU3IDGRJQDYPXmJcJJayBwWBTM3NnYTc7T2
5Uti6Bca1toQ7a/Qy/T5O5Ukp700PcGGBvSgmjelta0FTzRv6M/aCbMWVjXrKUjpceQVnC3P0sBY
34BdGAyxkL7Lhwr43sLWiCgbMNffCsNT7VD1VQmPe1DZetw6HWGpPXYQncnM0q5aIroDHhTmMty3
qGsQZZGNSzLdLzWSGBF9RHBfxPy/VLaWh4NKPafz5hEKvQs4/k89Oz9XMd7+UbQ3etT3HwlsqOiO
UuUEDxC78Lq1f66GTWBKfzKJ1/ksSBmME30X8yYjkzIkEkPh/FIZ+7DCPDC1JiCi2xh/xXHZGP6H
XgGrRJUbtkf3bSd9OkKj23i/Tws6k2Kz2YLR/c5JYVWc3HjVODc5oLnMKfIJj7/vc99kWUtb9ewg
aD2EVUJgB2/TEE94GzMqlYYSnaxSLh9cpRCz60fQFtt+Dg/sgmIvs1GPEDvs2MvhfLX7I6YpNgeM
jUb+AsgDVSspXjkMGTDzUJ6SgbofpfIfaloGLZkfAxqZq0JSI3SX52WawgVYhD2Xscysgj6hWTqN
YyBbmvc0SG7g9fhfNXljHepgAUk20PmX1C8MgI2AfsotZKPpa8a5E200AQW3UG3rVBOftj6Yzmrq
ZmiWBOl3fPTWoEVMmLBephgp9mmFK11JFpVNz0vtgo774W1sPAF/9ZiwCH7tzGG0Qz3xga7w/duG
tVjRdTJe5U8bAzbStF0uBLSRYJ7CSHzg/wyedceo0HFc9QxiA/ZpHTtHf6r56bLLgn52Sh4bcCZM
dtmcGycYhqHvUCwcXgqbTpB43JnBxYwE0+GX4uOFz2vgnrUwJfTI5neWWJBjX2+SgZJRnKwrpgMz
UZfXuOllOsypiWXhr/N07UtPqtTdBklizlFyS4092AYQMwu2rCPcJesS7tf4R/lCi8Fq/q4RX8Z6
nq1DMESnS3TtzWDwP26/B+bL+Ls6gmSVeaLNxkR7R8D8DIWmnwUIPMe9zakwPyuzovxztGJJSgXe
rn6K/ONNR41HD4RzZui5oFxbm+D2iXzOXFb86U4w3VHE/WZ784hfUXDGcMzz9iRK7KC/rZ0EMN++
An7qje+hwFlTZPV5hXOvyTHAxrAn7yOxPvTlL0dqRodXpVXhvKbKdHooMET2PMWzldW0SbrGd+IV
/sHZleJvN+T1P/vrwq6jltwvTuoOqXuVw25dq509/Fl27y8123E6b9NR5pmQDgkFjoA9qHeOY9AP
nUN7+lYfncHOexVDZONF6TU6QVfHhV5hpQ8chy4ViQ5aLTg5Q7H8xihUjV2Vt3VoNYP9F8duHgqp
R/rKzWkBmnnDntUW0wEzvZfITBPPv8986mFo3/gjKuLiG8Q0bv1OJvWoytm8LaZh/ifK27j1OktN
aluCa3ynqWSbUSwBIY5pdul/v8IYg72qY8SeGtWDFpuKKPasSfsmQHlRxY9dWCck8uN9eax8fIH1
SYxmQmgVxVo67bPgO9XedYW34M1XEE64blnDmBopkA+a7qhilTozbDJcsr4ClBBROTw80wHxj3CN
LsvTH+9TRmwfNO2xq5gZuuhBGujSXTcv/Z6sLjv2nOXeaX4g/MLkz+00cwJlkBi6K76cvWWKpHI3
gg9KAgMzuvM6g98DLjUDERc878JhK8MLSwSmX2wXOHbPaxXvpf725frUu14z49LUXmShrqVnIXAG
lalx/Wl6j0DbqxZQXY4YrTbFf+1kfZwQsbNVLmKb3S5pBfpQgK/Dpg2iBHi4TN8HnP8ZilSt17+C
rFTId5T4jCR7fu43r82zr4Sp22RLyb0iUmwRfMYsHpF108ahO87/k6jUKE/QmfDh7XIn1qvwih1h
6iAmBS2esNoofDz08eiLBw6A3R00iyk/mKoK1kw3VtSm7qP8gisZKF/0Sr+SeCa7BNH4bVhcvmiu
Ck5+FkTMMYn5/clm0XN/ZbPGlp3QHGeVWOHHfE8xzqVOS33tYfdi9vrJFVdmAA513FaTqSy/n8oX
5mkKSHmO2AOBcyionaFG8QQxt2pSEMyc04X0ipaTv1ErKqcdZudF++6SA5nNfkTUs/zG+MQYkC2x
V0L1wU8kS1VX2czX0+W1gpK8VM9lGLFLYTj6jSWAh970NuxDiqfxTcHj0dGby5qOdaHDMnHmPU0n
Q7+KZDFSOqG9ArOZPezUBKiXdIzfYTGgZOzHajN/XhYHYUwvwyZNM+/E+ecHx90Stb3H0VUYS0lX
9JzcTgf8X+VCnbdTFMhrNyy+iwyfI80qMOs4YORmNn88/1+R3a5qJqidWfO1xZyT0Xt4pF9fndNF
lYKywyrraNf5zhMYV+iArdEsoMrf9QhaCRcNGaFvIkC8J5nCnCz6BLJKduYi878aw4XpnQm7uonI
wYkfTg0MRNE/J3CYpM0nZe8wzWOj3NTc3Ej5G/Rfsu7a/IYmTxMh3ss73RjOZ4pXLe06r5Z0ZriA
2ChhICAnCmaJTOAB9h0wA4F2IcKMOl6rCllRtUYgG3AziKv5GQg7cBiiywgYovjyJsRxWtOBfcGh
h4ZioWKVnWon2EWyFXIJMtGDpuq6bcq0AC1UZt2v9+6An/kqGWfXdArJFy9BdLHjDi6wx5Ic2Bez
X10ZgjiYYnti3KafTEPpqqEWY38cD70XPuEWnuPLjaZckgeWI+E08uBJ5fSMP2/tAwiS/Jr0+Z3s
zkYP3ISv2m5Xs5xNSsqaqsURPnV/p+ahpj5+ajW4GlbDwg6FnVaPC3TqUFn6xMOUFd159O3267UD
jWJtvJaMrV+Ef80ePo947L5EBEaYq8rk2OqBNS0GaRsZupU5/85zS9uy3zCZTsfJUZfOamvtfajn
PusPqf23Gb+EVvIja52hIrSXx+enqIaLQcJavG/gVdvcnC9NTfhKz4Yb7DEMzAUkQ3q18Ypdi2Yx
2//XIKruZ2x7zfdovUiNT250xjzt/XG2z82/lFG4LJx2h9nCo3Kul0ZLi5dmdoRJGnEsQziUBFy5
x41hDUs4NE5o8KM95eFDmZZc+vajnJwyNJu1i9Rjx9lGk4yGX7TGkjMGNiVaTlGd5wJfd2cfmtQ8
0Ekq0uEXFwjjPx3xzywfgplLQeC71K3URGYy+u2Ddl9PQpEIwNtcAlJSzAQv5PTyq8XrUjFi9aNv
0zeyt+Hg0WJlkYdsP25b2P5DaYOWWFoV9teLTnOOGrjbpFPJMtSSpzLem/z01uxFELpwYHLDPu5A
olPupDsJFfH85KmGRU7TLE7k0yFMm1hyo8mrLy8/BOKRvBruVEgf8t8NDJYgsYdvYgetUFuPWyO9
rmDmUVf1TZtUXDxnDPU/t7ZTvAQPFchGlCEtB351MN2mTrbDR1U4eEIGCYtsc3PiahWkqfG2zczN
eeCFGVuhUnojUDYj89rHHLyv3vnFeCXIGnvHM49buGUonf4Lu8eJFX6+WuvO9CughHHSwQEgC4mw
IolHtSR64xM0+w4NwiVktpDncjFHwfSts5DOKuKDs0ma9g0hYF1TtsHcPU5rvuRtmu12hELwYYVN
ZUoEL7d0H3hX0NZf60IzkgFoMdEjLj806w2nd1rephkWL85rczher3L/PZ7/qnGbNzIykXd5S2xs
V+ghkWhUf1RlEfCWwRX1Dv/h4dyZMP3t0e/wkz9WyNKmIFhSNgff6dAm0ok52Gynzcryct3eFlBz
6cqCKv+q827AdOF4PDfz3c9uTbslh3o8dRzUU7R520bL2PQi8WNcRCwgtVSonTOdGK8FUlMg+ONr
p78M6/+ejbhGW+gCdag+dDyItn04Sut8LPBDSqjRdP4WNkRwflds5ZpnLDlTdxthGhcPLoh1QYv7
ZotVFNroe4cgvE7kDVBpCB8PHZ8na0ehBK0Nkv0XsxrFL4LyddAYy4EB7dN6NrlBxzmh5cChlQb1
90v1zsYFuzVHhnmEEhasyvYXHtBH/XJxjKTTuVlqj+g/6Erx66jBmuwEvv5J+SNZR1C4M5oYputi
3oSKMQdxPeT0P/JTx89HAJcmFaUOenlZao6UPRvmLDU/LO5fZS71zwiaBK+5UvKDAZO462iGMveY
Rkr4o8mWrcIoV7Qu8AO8RP3MCjnl9tWSOGa0wDa5nQQoTmjJibichvDzoDCOQ8UyCofnMzd1C443
0CkXo5bzOx65HJMHQlEIgzAsYesm2NIXDvAxwBkK4wkEQ7oZi2wM89UfyGfdXAeg3iq1izGwakCP
k9rnEfwUKyKCJUbYx9FWdi29RZRsCwDFuloN10WGLDJst+peaWxgcCl2mTbK+lM4GrVIbKuAn9eI
K70kv9xG3OKQgtgmqpDYkSogjuv8iDZ6odgMInlXmauSTgwhKd1oPKlCncbCgdX7ItTJ9k+ySKLA
0oNwtAQV/zMbZEIA/L29XX+Dms/9x8fCzLp0G/1FqRq2Z0klSf3anpeccKp6Nr998kwEtneUDCAY
RLubs9poi7LPdeoSBFceCSZCva3Z0L24nQSkPvMt3pdNc4ALBxChoyJWOt5A6xHXWnXAgdWSTXWj
jAZuemp25S8umkKfu1UlfHL87crYDyz8z2q8Xx5F0o4UyQqnleN3tuY0cl3UCDXcFfesBY+XFqNA
v2yzVyXsoGjGPgH40cIK5rBd+vW+nwl0Gz5GIhBB2rz3mQtXfY2F4gL7vFWSHRsDq2hAMzd8rnmB
tZEn/1VqCymcug8b4UU3twrPyz041gGmJcjnmO5Uq0umBa9vuXFX6sYNBmGXdkST8SUnFyIKt0l9
J3pu8aA66z96J3dBwCJHID91mLjhMgwEU5s1WyozH4qKyJ50lKSy0cJL0nKdSh4ZiGgIrxkezItm
fJgbqgmESxHAnw0fWEV54iBCWtX1POXB5RCfctySUHIUWZWKLhGtWI1WsVa0CdGTD9c4zfF+iDn/
UjHo0zt/rBPIMFel8ajkMNhUlrCwVG5V4TxoCO11K4MvO2uPTjnytiHH0Pi9/gjF66EUJODm92mS
nBOR+AXM2EkGhhcazKkWtcoHuqYQNOIH/pZhalN1uLquF0D2ErFD2PePnnTV2zyqKTdASg/kbIiW
d4qN6IsPCB3ZUR047BGZRCYziFstH6JL4KAWj75L6GCaZnQ9gkWhOmepz+XzJ+oDyqyt4pllHyTy
llfMG2t00RYtqGGBvHJyVt1W2n5aMx4ODRPn2fmjjaukg2HsuA7oZdwyGrRRLkJCChB2Eh3+8B6t
ziAPRgDB6UpVrfDXhkZNYhR8ElFaCfOw8bul29vvHd6w14ky12MPHTUbTMDdnGotfMwnf+MdYGmZ
SDydClUMIJVkdCbSWrfM26pFTc4ftP0zZL8pC6lYbWnLI1ityccJ2HSwc7hNU/HRF4RJYtESA8vo
g+uUW0qoATw/me9dKt48vcTg5helGHPTada/sVa5GReQf86XwSHcRY2ZDavU1LhExH/XbhDdaEIg
pjHa3K20ZslwEN3xbHIl6NEjzcx0LvWujX4mlBZFYZYx2lGGsRF5AHtBi22NW/dU8BEI+GJkrM5U
pS79eZTLraQMx2JCxJR2rlsQRucSz0U4zHJX0iWusASLyq5o8h5YlZYuxn9uWmc9zyA9mzvKBUAu
17nxZC4MnE11EQ2k174h/nyudb+JtySzlu3pNUMYNokWDxTm4SFXyPl3qTWfKThdrDu7Gq9lS9cT
SOuiQ07d2dbszrn3eyGzZeL6AZDGC4rZmtdpbTgYGG6WkDmUNY4awKKSNMwvzWpiqwPhjKgWUcCJ
Urp6hICVJTz2ySk81EyXm2ulS747kq/QF8pIOKNpUCb4jwp8ioD2TolWdppKbpgYaP3P8EhSv6h5
VwD2FP0sfW4yWOdETVGQTfYOsBpaK/oullOc3y91Nk9UgD3bqU4LcE6fE51rrUeWRWEPk5s1WB2A
Gi9+cpxuYzhtu00rBoGZ7y+arK/yyCFwjgNUec8EvHLo3FVQDUZLvTzGGUyjtw0Q7fnKm1Au+LGZ
PZZyVnJ+wgA+t2GTp+X9Qa+w3T0RBq1hiyR0Zd1sYeLjlct9SnJGHJzWKLxzp7mj7Y4BvSjiKLlN
v+5+L4p+4DliD1WVUo1v9FZNJln6gH65imcv2SzFN31LB3M0rV/Z+z/S4CN5Qz9h5W7T88TYdLiv
zrKw1Oc34LvIwaYFxEs+1mMT9oFUdpTFEHZIYFvvGtgNlUjE9TEeoUKUTMbT21ukOg3jEDsoaoKQ
W4WQOTgg4thwwC9bm9rHSPXPo+NUjWfIIRFmuOkKXdNrdXMvOoTEG+hG/SbOgdVCELDiFORyvWoL
1WL41ozsVooJaLg9ZNS+QI5fh5pqEsT4xoWArP7whPfLthWxyl0QHkqjyMXF9L8bFmGyikM7lKSu
gLJPmwp9rnNG2FqmxYo6RlO+2QZMRzv6Cvds/BkD/YuM3ZDlVcdP1gmKgEKYxqdSLD5/id28M+Pi
8ljpyYh/jry6e8jnNI4c+SEhxv4BJ+y3ozm59J13loJZE4sSJ38vlY3GWCGK5TsTTn7FDB/1E0ns
SQm5EMeTI9vd88Io2e+wN6DBqGrOJc51DfzGO8zOYT9IPOj7EQMbXCUCD772FHdWEJz+zwia9UDs
5fZ3hLox30gdkX2HptZzsoUlNAghsd7M/GHBo6JGiIE/voYvJV6eSxGja2xkoe5OobLu3bG6EbO+
hALSshlq8Dc8R9EpalabO0xVeLoGDHvYnEscbRRgSUFSlwOe6hTmSmIBXWSeYJ2lTeY6NOQ/0syb
67KmznfDoT9sZQ799K4WHSp6HgWKUdDso/5ZhyQQtY5o4b3duiy0zck5qSABvNAuWFQn24CpYiDZ
XIoz5YM+OWku+Sf4+am6wLCvZQoVfR+iazILPJyDS2q4RjYWubbu5Rm6SRykfyPtAMFqdSVQVFgC
oMCOooOWJ9XVXUI0P7hB1u8zS44k9BQfhvV2dANK006GScgDAOEtDHvlVOeybr7A+km4xNfHSBfi
T8MnTmGwF4fPROEnmGFHzu+Dg1e1PIM9u2/pqQ/Bx8V4jzzmA7LOCate6uYkDy4nMUSd4afhc/cf
FpR3gpCo8XDr7r50dT4LWQODPWSUOv8xnu6LGvt33WKhd7op1K3tyzUFGGet8yayOXBIq9yhppMh
9XH9nPjiT1n5rSxD6pcjtIEzOYY+s6HPDJh0nu3pmFfEPqhB+dTzdobK5qspvgMgwIGuOpBwxvmD
m37saSLkuhM3lC96UXGEDRaDD8ApYD+HRIUOHoYbdHlUUzO/ykH6ibV8CI9+KOuj8swJuhT9QPcH
TOxcQN8QaWxgXo/+fjchDVChKZQNHYW4SykiRJ7bogHduMl+p04icbTZANFZul+MpJfPTF2/TV5u
Pv4VWsXi2MMcN6/VQgCvw7WbKtoeaaZsmXM8uFYNdUYKNJkhYS3HTmy7c666JodHFutKhCUEhZDD
GPVJ+bb0VQZaGtAXLN9CbpVJ1PT6uUYbQBIa/IUo7lVjfODpha78V8xVGQAf9BA1OUCXx9fMT/d/
Ak9J6p/BUUbqbQj6y8Zv+tVmSfH3CV5KUS3Asqfd++dkWQeAMsBxcKUYZjFfp5lo0AL7gjVvocBv
0k6DiGAw0PDB+U/ToYdYCd/9l3jEi0atwN8cENhPd2YidDPS7K8g5vl/vpyT8ij4sRe9NFqOUBHF
6AelSNM1A7rMzVxT3VZRAjr0Kj64gnNwRZxZhYetAbZ9+2vbzIl7zfk5ZVmkVtkKQZTSyGHgNf8+
hcvJaDhbMwAAA9QnzimhNXRWdqzXvPCaaJsNhTwdWUy+cOIrxQdpO/Rwt3QJWf2OiIwV6dy5Wb/6
OANfU1XB6U5ZWcAsYbTWUONcCXzFiAsCD3pWnFGeujbPjt9MSqpc1jtMs9OlsGxruUzaxFwsJ1BX
B9ra0ZjtTm8+AZyC4EijPAaEl9x1mOMdHHzByPXRUjLHF50WCT8Jr1GfxmvS4A5qTlHq9aRTCh6v
gXbAuAvp2675BqEjPO9oZf5JDyvXeqLYNVHf2tCEL53+uvbuem0W7V0zYT4vR1qlTW63IlJ75sJ6
GzvP8x4mcVSOyHiHnZ6cF/gL9Vt1i11bhB7FGRcbO68bwPOG2DL2gSwyIweVcCUwj3qrz11vMLbn
iL7r2TO52YuNqjFrm0pYDn+mf9Q/fqSoXr7PVRrbTRunINB0ClDOcxjtBvgOgtD+u38U06qXFOYA
Br+L28+PIi0xyGQvsci6+8lNK4DU3W6KmcH/kWZzVYXiqI9kFOxO21obZMrtfTD62IBl3v57KrL8
l5HE2LWKAf3Pj3tBYW/uK6UUNVVABpOxysdzPv/23gznRzbIj7gcuosqWPttVLJROIzrXByjV/ul
LX9KFi9ToWpvlL19w5Bn7Zv4xv7PQ45zdtIabgQ6mwRRSG0AOwutuc0U/6bHw3WCBpF6ljrSpviU
XeBDSJx7z7RbAx9k5ZDxbzVqK1YuA1wMEW3RGp1zSE8WFALZzeoQYiPOpq/PrKcyb+87EXeyPwRf
3yCgBMIEOcA1MWOBKBk248jvLPQCFPtwMSXllh4kSM8X7YQNvh0WD1+PNnH0ZDZZO06dc2bvrLq1
77xHscRPZlWMcdHAiG6I/nAeRLBZL2zF13wuBdr2Y+EHaKpw9HqFwddp5e2b/B65TJDwMMa27ECL
tdanc0eoAuPA7Dsvkxg5cc3FmbO+Z7ZG8EavAwqpUid0vz524D9zjOd6qAvhZ0Giqp1MvpKw4obf
vYc9gkMEJqssRqNU8GNbovdd5OvWjRgyjKnNW2Dm+0aKVAMGBX+48pqLFz7okJo/yQ9BYnaPK4ky
Y7FfygqoY9PC1NDHYMUV3j8mLkqmHHMxW5Vg9OoJKv+wJppOVMlNezPko/ohS+fgUFC/shvX0J0K
fA13QOJN+wgDFT/b+LW4uxn/6y3PD6NlHYG5Ff1d1pbBJ7HrK5t011NheWRVuiwOb0ouZJKbpbso
Vlx+v/U1gX0F/pyKkakRtb04BS0Wr2auDiS0a95Ly4UGpa0IQmOPCfopdvMmkJocjl1/Rr7G9IQH
vLD1sgjFsKMmCDJP/tKenkfGmHTMJPgBwPhS0HmRECfGumwQqWYV8Ncd+/L3XTAeuIclSB64kdNn
D02it2c1beVWjjhrWpO0yiN47YwpfFdGJy13/RBjH8klZ5v5W0hEYpHgebzYC07ysxFB82BLTHQG
YYdYgPKp8W7/utg614aD3BH9Dkh45ciakT4g5O7akQQGaY1wNcHRLnVDuuz97gm2ukxm/X9Bb5Rh
42OsxEV/6aogJxRe1oO5v08Scya7+QHLyr/1zUDy9g26xt2YqGDqRFaMfhOiR6RRTuaX6YafhB4d
uC7rLSUGATI73VL2wQ+ytlOR9A3Sc+/9PiH8dwoMNFyw2OnczDjz3VQ/6sn5SJicbuF4a6kFDt/H
V7K/1PfFuNaKS5oE0G1SYepLUpKcIP1n/nkX2g1M4IyoRiOeQiJAyq/VQVx88HAhJjHQybZZgwCF
3gSwJ/bgR7JVCYHQIXOHzdFDyK6QBSC0dsZxKg71xAfe9xrKDJqvG73DAyQ7m10jvIDXzoioD3BL
VE8vx80v+HMOrabkNKmCIkSp24V8/P3SuntPyOAekbx6EEdAGlntT+vUc5vIvP0h3SMOmIuNE4/q
Ri2MHJNihcKl0ioG/T1HnEdnT16WfEMcJ7gdBWEFH+QWm5T2vn2FUnfYKpiha/mfl+DZgmZRQMjC
O61MUMRnmHGW8Xd+AmmSeqsFYOfKtfhgo75EW2Kf9MTkAgfuT7MRYjFakuG63ah4/SqVbqoJ/cU1
UKD1algC2bS8JIUFr2vS1DMO9CDU4lrj7uU31x4y1wEQK2Sc56w8GO+mORuSCWrJrD2FO10RW8Bt
DiNDXeCyAQ5Mq2yEtC3URNqtX4KeTIXhOXVK09HFetv1jTW7FJ1E1AqhogH78J8pufVUP5mcqo7X
R4s9Q1i1Xyw5mXG1M17TksWnClmLThGSbv//0WZwqp4xlg4FCG+BXM1h97pigt9hu06/rjAUiHQ2
SWl1dNeKe0kaxaiSiT832+loW4nzMncEB7grclgFZ1ZW5/WRtTyQvYstmXWQoqli1nsvGQsM8APM
m6p5SQ1Bketx+WcO0JdTilRjGEx0BGFomYQ4Anefs42MAhontVTS7i8i2X9jM03aTImVL8esdfHE
SbAMH67oCFbqufS1xKFn3mCohq4nuVr9hw3sd1sa1+Ppm5EIsOY5RqPcjhnYY7GR3GBr58gXmy9k
48T6bNy4lFufuETMlqXrL7ooeL67A+uf0K8b/hW9k++2YEicP6gMUCiO22uh1+sYSa8/B+LV4rln
+yyCSBb9QnAFh/MhUH+6hwTyaY/fvCWcaZMR36uslP4VUoSM/oBuZprk4HDqJHGMJ3mG0lk4nlHP
felAf/Fz5VtDP1/5TwtTt0VOynk/IQAeXt3UWaatr2Ibt+BDCLqL6+pPcP1gmNOUNrqjDa3g0UmO
YEY7fcMdpWw7mof/k0d6ZKaQlE21ej73+3i9da45M1srwNHd3F73BFAmmtw8coXIhfZIaPkquQ8J
Zhe6quxxGl6WY9amY3vDLS8G534pebko1Ng23mj3IG2r8kjorIWJy97nyoKvNWRZ7IhSdb/Yz/RX
6oVY/7wk7+4K828vA50WqE66pTCWcFHDUh+ycAAkZo8/3Nj+1uZ5gh+ewsh06WioWb02K+7ytEDA
OPwiYnyTSRFpi1+PHGMUqxG6lRgOQ3S38Dlwhc80MEeQDRJHxVKNWDtXEuQdbg7khyHBUszXL3jK
jsRZH7lMqOs/TuzLCHQaLMeGu7JimCEM+2kSCxcVm7euI4Mrtk31MA/i+r4iYzhNnHtl2hXEv6PV
tyiWRDHAG0PcVux/nnymN30Kpg33WxNU3ztwLs/LmjwtcdDQMDnRE4oxzvv/i9bwF8E/b9wG6bTl
vbBYFGBlQN+Nz3xCjaVvnlz4EXgbRSsDXAHAyLx1teUwzy8E2t/4u5uZYzX0nHgxgtLOtYnBiYWl
x51791JJa2ZIaBRzkJ5roWSqOJ6WeWIpohuMTkcKyQeVLbXgOEUmoEBldq6r39iuie9xLIf7h6M3
Jun3wQGmhKSScc4EgnD/JpPxK1VogsPKupdEGJHcmj+hR6Bq2Ymseq9HFpWUG3gCoqYPI30JPs62
6hVaggoSr7j9p+9nOatNiC8WYDeq8KIbsf9nKpIfW/2mkThhq5kL2YQQvJwnxuX8S4Y24Pr4wpUu
pcXbwrEgg/IFQ5v5EmOw2fhacKLtDNitLwsroX9BqLmQ+10BYeQSbhs+Rw6/a7wu0z22MCSzogf0
ofJHkaQnUdCtEg7pUcpgecBvhc5GUd8LH8bkKJSHlWF45kHu3uUAS/tYWQAupivjcWtWTBr1fEtV
K76S3JRrY5zxFqHahR3943ODOyqet4IZR1FZ1lwuwDnT/sk75xBHPkbQOnS7Qa12ydmPTeh/bhwO
4/x0adPULZwXlK4fSiZuqFZ07NFwqDJAu+4Rh0riX4Uh2JT/ZlCjyJkCJmKY6/oiKLlAB/MDzU3P
7NBE9lp/WYD6QnQhJb0fYCOkE0yloWCQOjE5b7FR4iW35tFjvDSP03iYH7SS+gOonl2/5Lt+f8Ck
MlCy6GHgzWYTYL5UoNeTymr0CWILwHbkVtw4B+Fm4xxhCUsSry/8akLPF+eMSTAimnxp3X9xKfe/
H/pQtjJN7Z+5jrH7DiaWOQ0KkYv3P/mCm17oELosvktx7hZCOaofXw1r+Motw5AtbPt8M9iWWtnj
Tn9+JbkXsyBO+pkwM0VYAGAcWbxFb/f/B738cHoqS9mC1+y140IacvaJ5tsi6Gabswi/z7pamsRo
gFLOKuqgUHR1v1bF9+waW9rNbGXSiY8zXqYQZL/Yn8J/hBQ+Y1NJrJu8q4xkZgY8H06M9MBm8QCg
Ji2dpPFVBi5uaZhMbHdQONc74PxfkfCnpWxmgI4BqZ+FkIuVRAC188zJQPibtpyG1W/nmwTTkRCm
X55Qd42FJbIJSxiWmfsxZ3WeEfjknBkGbUFhQzn1L8+EvbNvm9r2n72Utd8V5upBYA4SEV8bpIlv
Y2XyHX2cTIiCqHqUFQI5Z4Lq6uV9HGn0XRZg5tWCW9PHdrz/wctg1S4T3id/yhgZS3EZPmLlDzWj
J2PhKPEFWJ5VDs4fgaIlhKulstSXDih6hGcbs2clQcsCK0Q3pRuILEqimMXg4xLen1lULNCP3yEc
wdgvatviacC66siyfAYODTugb6mWudlbsqEtC02O5rrSuSm9YINmzAKMReo/ibdv6niCl39fhSea
KHx2JI4+HbBDCMa0MnoVph4u6mQQHyajHGuCi897zF3MPXH4W0Yf23NIwMOU15F1Eo78nBBHw8u1
EtWNpaNkmfEMrsqOPKwali95t6Crh6lcdu7pxxUzckObZxQ0dDoXjbkzn8woR8jkMQJXaRE0g9Af
dJ+/kBtIzV3P+KTfagRSC+0DgwCA3pZ5YmywUUtrBNE7LEePvIVRGHrKFM+7SjoA65JH++ON+MJy
XwgvmmJc6ZqEfphNaGCSblSADIHEuPFsr/h2jfcAwyVTVOYploDyKu3aY/KYU4ly/mUiIDansEfw
2eV2VzhPFeicZeZHQuLqIV+AfY42jl4u4A7dfZVgvFpqd8M8wXMMfGO0214ld3yPRvv5r4Eje4rv
GOgKazxLCLn0SQJ5anoXI+CrPGDZnUdze2dc1/dS8QI3ekFgIqLngsdySC5G1hRsVRo4eygmb9XQ
d9Wrik5a9SJHHOZlpUzWkQzegYo6Ns8ottZtKhF5741THs5YRZi0jssasM3dOy5Cg+nK1ByN33F4
Hh9YadmFdJqDdaSpWJq4tNaohwCQN2XcK25304rnZjjWy/HzSaC+hoJWHdZW+u5m4hoCb0xaNsCj
3sI2OkZ6JDgrp74/K2+LEhUTpfOXh/TFuPvhqHxJAJCYoxIblPrgw8V7GTwgsdnM6w3GbMEqv7u4
wJb0KlPuwahbN1DoQ3tC5+s6YDlkvMmdOxYMcQ/YTF4AtTqydTJg9rTTBMRCKeW7K4WweT4APQO0
zcXcmme1SZCNxZibkC/gzUVqmHQfz3HJkCw4/ShsMyMQnybQmczOThED0t38C0YcxWGJja/ef6Xw
7fOQposG0ab2LL5+oSJ807rIHGCJKoJa0OjFdZudBbvCeXVwTdx1/TxcNMsw1smtwIykgyF1jn3N
eY4M5Vj6jSV5T5Lz2dcqSuuCGkLe2FWpIrM23NfpVJNlHtvDRsUBOY0mNbYVHlvbXJZD8sG3MT8+
kQZvXnMGg1PJUUY7cF8f6cHijY71k//J4qNS7xtOYSIYLqDVEtFag9WVldAgTe8NJGznGSMhYrgI
RCa/1MwVkl7rIHWkFdCXXxuQEs0/kUmwR8udV59/NuDuarrtZAKwEEZZZFr4kRABm3oWVHT9jhpk
LuC9uTqYCQF6v44xG8PX9DXA/SQ5QYQuLC/2lYfdDSoR9pvj6KRIScYqRT4UT444lUPFoR6/+Lq6
FIEx0cV/wbMmpcJC7Rgou5hgIecGQsanBzSj9MNPTNyxVf8tDkVcy0OO0kny0Sn7M21lbUh0pUm8
RpSoFnHKcrK85QWxyLYeovdxbBMww6g6e5MenqRDNIk1fYYROTv+BTx3cZeDla/IdgF2Pjgy3AyW
Gxjwc8ovnjhGpzHvbPiU9GJ4PKsjkxkPAPdHeBviJDLnqiQHXSAwvjgn2WxD4+ntcxLU6B9L1MCi
OhgROv0s/xDPcRJb+lQz0i25DN98Sp7Uzp9GFXGohL8e+RLaKJn77akFhVjwZJojWmaSq2OIw+eg
7qLStKayPfIv60CMcUlT6rcCUD/1TZKXdOuXJVZS5mDHv3wULqsOTiwX+rbkp0+K1dLQsQvQ0YPq
5tlxboCYRudonglqch4pBPDnQwdT8cJkVA7UtLJ7gJSz9X6x5NqtzeIs8wnKszet1xvwmjHFEaYU
FSh3ez/6GDn24XY1hWhzHlHauz26zVONHjqA18o2tKd8JeTzFOapjr1WydpbWM0g1MoRt1KPVaRD
+8DsJ8MLDzn0fXw5gaObNMnz1IpuneDRSEnNSsSegIcLaZ6BWiWQdMfzSmipa8Q0jGnIEIz+pdrA
gSDLa6RYBr52zS4/GOV7rEzCnWmcE5gRgD3tm5txQycMGuk3VC/Oe1MTR07qktj2XFj0mVTQNVT6
N88aEmpj+4z13eCP3bfURwGgfgrU9MCcKmB+xrjT0f1F67Ep8kx6Hutq8jVTvIo2XRYgjRoZiIj4
kHqHjuSDP6ogLO8S4vhtp57rkZeNtqz/eqbyh9BiyICFsvXk3dDQMbKwRL3M7esO3SlIsxKXWJYN
VYBc2YR4tJ9fXKVSuMHv3XP6SrlNDsUSnt6l1DHA4wXsvfK68nxkiLGEqPbNDBWdT2iJVFuwnZ5x
XFakYuLejp43UMOlYdY1fT7uzHzLVjZNLRVnvUAhRZi8Cyz2HIIKj2cmwZDeo5w0cUjakehHeiCp
W/Pk5dS4fqT2Z39z8ly2QqigyOPc648uVHwWgJXgJFXEfjpHLOldtILjoe09yRTVkG8A2th8RtfC
Jfv6/dGk/vqRcGX7gnwte+qF5PtVmV+2FTXAiVOXVgDHJyvXPK2INn8bYbup5cmfcSye1YUdlHD5
/ViMdP4GKbz0Jr8vR17A2vheNrLEcvN63N6SGVuFt2ZwaCE8rsMnK95C7JrtYa2LGIVakxhOkWFL
Eni5VSQNsqZipQ+zPeYzp7dF0kAdkDmI/TlXQEobXfMl9O2d5MzHw/CdA8TNnjrKuI8aGr4zag1E
UPgcBpZehPUr4Ug9N3OOzc/e5YGkvX0RB9ESceRnZA5OR3UT++CyDay2HdqQwbl+uRoEOIqw+ZZl
yZQoL5ryXpsx34Gs9ILcKtqTk8vJGxs2ZbhknF/rd9EpwDksXqbGNhD25wy/wFoV1n21liFyhW0D
+0JJcbHMskwYw0aJ41OGvl08W7VOYTgVbyHHLQolweKpx9xJKHWkdmjB2AnMW05ByOs3cdgeszmv
mCO6f3E8R8yMGUXQdiafTjMNj9/EQQV9XL80qaxJRDt0/+d6eSkE81IJKveFImdz7N/rIT06iJLo
AlrDmfpyA2Pi1nkThFxTqiYgyUHB2vpRxkdoz2VI9rGf7qV2WpxEFhzu2gg1m/98/bF4MpK5t2i1
YBSNJpcH80dzaCqFt3zKpnbd8cq7JKRSClJ2L1xAwNmAWB19uItkCcCefS2OqNC4zoVSxHkf01QD
cbyfwckFd/p5AVPwHhcHNjtwM9OGaYfcmLWryAbIJzAYzO588Z6GDl1AwAj8uAWg/gxZdWEme8so
bWdT1ETyGLAm0jkZE25aYMiIcNdDQQ4yuC7NoF/NyGHzK9tDluvuVTduTTX8uS+S4OUSGRr02NIN
arYRgseJBchTlibMIDzJ4yjzWVScfRrw9om2b8G3/v8w+z9QxBONEtsmljVfUCqGHxJ5Mos8jQtb
5oFCrYBJTGFKjHUNENHSltyoueD5YmZaF1LYbME6rFmzzsFbPHwK14Dgin7KSF2h8SsbkvUouHhb
d5jXTGKzTzfljKqILwLsUdaEIVEfusK4Rw07jt4xo4ZuBHgoe6JxcNrnFEfwUM0CS/lT1ZupeHeI
gJXl5+/EXCrmea+pjSdey+f+dO5XANnfi7fSPcOD/gDnDq4WQ0UOycGXFjBecfmR0G971KuaY0WM
gdL+LJxQ6VXVzA285wKqFvgjGWCoo6be1rZXfn3OcAPz3610W7+B3XUUS53yJ4TJyiPNZUrNs+oH
A9E4csjTcOBJEC3vNnzvhLbKXZy4Kb/ODEcmLAKzlG5NuZ3v1XYbMpErCUC/ULalYBE+Qf2oenEn
KZLOTsXcDw632cYRaAICbcr7N8g9JDmZCQy8BJDOZmoUoYb9nwmzC7Jko0QSTMHDnRgWBuHVPFej
Jm52UGBIiDSmWZDGmi7fTNfsXnld5LwBoRArCjwDgBUythI/SqQcfr39JvB7sxwU4X/A7qS9NqeL
EK2RylokBkYnauNkdcXCT9265tUCQLPmwD7qAB3DyzfArZLrhD+Mwk23BiRH0yem9h3z0CmT3Tvx
Xlus4VF1opDwwHdU++QJDpg4OV0YLDFkQ0PoNNdXd3BhhhYhArG9z3iC8lxFdNcDdjohX1Q3Sbdm
stLuSce6xx1iV+8tJ+FJyysyKUD+lG8PB2TODz8E1Owyqp2DtAcp5QhGKw8s/ufKQxzjH+sT0Ti+
svswdvs++WbsffyotCXp3U9iWGrDv/Q9qHLm18TU6O61r+l9bB97KdAkrHzYev8AscBb6WOQuQA0
W9xi8FZVeaL9BG3asRgWV6cQbcnoGdhji/X3bcd8LU+mhN7nFrd2vdX4wxrtG62PGlXgo1fKzcdC
qXc9qdC4vFvVE9+E5z+BfwOt5csA8pXzMhShKYzJgQ+NAu9butp76vvxaPMuWeEOhUig8OHlBfHU
upe4AEM6kpBqnhasS6Wc5Ne+qpBz77ITTwpl4/7slgTMYtc2NFpsrJGBLZd+uyDPLmFR3tb3P5d5
aH3/gy48dRGvfLZ9hZ+4+4sBXgK6K4YMrgOvK0EykGQP3z5mJsXacLmfRs4ct8NiU0WRZ6eK0N+b
Tbm+7U8eHQmRr9kvHppZOn/upVguvUpd53TRsL+MnJ9fqTAMMvmYgUM0k4Dn59ALuKiMnApEsbVt
Y0mdcaUmg+G2zHD1qoHhMhEdnm0y4hfbP/IsvpQ2SF+HhRHX37bm2+mof/zabouyju0c2W1Pt+U8
Xw/GKD99mGjhtrT9dTsK2zv7o8Yxmz4ZhyPGBaX5UNaJECX6YukYfsXuUZ5BZ5neyRXl+/9ziHiK
4jenLZDYsd0gFKyXE+csdb2Lh55+x2gvKXSagDUtRBTIhizTm96h4AlSN5MZUWp9jB9CbN1CRyGX
Mj+WBdLr3yByTSQLLFH9NXVix/CPkEdsQP7f6ykPo3nNbmeJThQ+rDNk0aeK/BvltNrh2Pc+FPxD
9WS4546lDXvlukD7KQaipnYFMvrF01d98GnVhkajN2ZW6V4CezyjFekj+GByy0gwd5GHrI+zCvZ+
kXGrBQql6+YsuZsw06PqnSSyQa0w2KtDxHfdilPGqHsGZnNtFqMNJQHGKNqA90Z27Z2mFfPXqr+E
jLzUbHHp/5a7JqNb1fZ5AogCcY9JLAbvWf3Nqp96zJDYelN9tUJkn6r6WOW1YrqSIrPp8erasFY+
JYFI9a/b6liDH6KuiaMu3Ao3PX2DQm8siMQpVSr4C8S/umFwCQtWf2pyKottJrUfrgKwTpevG57w
QLcDoRafDPxXKuAuk4Odc6E2QKb3OJ7k95q0o0MnUnumeG3/k1TnOTu5sesHSD7dGezpLDwZhghy
BAt/UXtWyHug0VcXRYX/q71gZSHLKLp0pTIsMR6HKdiwLdXgiSgqqnwkTXBIFBssA5benrfRZOGW
ZQXZGUW3cgESJH18KfaoVE27wDELIaC8yDSBrB+VlStFPZXdXucolsj9RxX7mc9CqLkMuZ3MzV9K
BGQPnQ+8JgP9fF2yarbNijZuuKXBG7eXGzCPFcAQoX1T9EdnL48Hrg0wGprFhkzlZQMK8Agnoi0y
PRwJkmASxfsYFqOgXviFWgmve4oaQlEVItBm5t0r41yIFtxmd+VcCX9zSYd09keQJxgTnO653OD7
0XpX7r3mo1+amIq0WURf7/x/IYBE0Lj97U+nxOy8R9UbSclpOM9K51krWMMDkoYjj3CEUqod1a9f
T77YHeCiwT7kVt0NsZwJUcxby2Yb4oCkp98vbTBJJQ3tHU8QCE581AAO//1c/a+iAXmhcHZcQH9E
gWCzN/XaL4+GC6qDGkJcvdGqUOIKlBXJop5WbGmyHRAgqX6P03eT2Fbnn/MSMuCfflHU520H97Dc
UtQpi66A4lKBBXiCnmf3md32eEhiW/j99hKUPcDwNPXxXF1ibqFVTBOwSI25zmJZXoHDty0L++tR
d4mZKyxsHiN0VUH4gREY/+0PDfPqA1tPWFjdaqfdvSeGZLP/1XDE5e4Rreh5VR8bISGo4FGcq3FO
5LoN1mGStZ6EkKrpivSbtgWtxa6PtIeYT13MilUJpubRdG2D2Ak6jYwrNYkroH38C5JOLP2ZHV6j
VJBHtYvmw1i46xDWM5d5DkV0uNCsQclW6SLGg4ew4++MlX/wFpN35eQJbMEpaePAa/jy0CJ+lLhU
UL6ySgZLbxAMgw1EPlATI224Y2QIW4ta8OpGOr4iX3MApJdmrZuKtGCQRBakf+OXlUkTTjfRERd1
+JgycLClpCxxQbUL5ovP1bmDAqjkUp1rhubktgD4HZl6jwtpRDoZGflPWVgQ5Hx1yJtif3c15G93
flDLGb3jOktiJhkvBSXMWDQKrdMSnnM/Ompkx6kfd6RyOhLYgS1/Bz+a8ecbrW3FwWPv9XE2hMcr
vTDulcKgu/OdnPqT/H42Bg2vxOi560Q7ROKvoNI+qF86ZLOeEmpBWK+rgawgJklNGd2yMHMyKcGc
ktHL179lE65ym/VtLWEJKjUqiAyMgb+iIFycgLTS5w3rvHee6n4nP7tiOUxYzhGmdHJcv4fs3LBS
uC2KgKyWj1yEQLYvuGdGUaq6ajcWHacni+CQRhoXH0EyCy/uaAtNhlNcWwZSmlVsf9ZXMT1n/qcU
V5MLNcfveRuaPihbe30mPKierCc9mTcinbz89FjjKSfPpGAdyc73dYKwkXGkiSpXnFdxcc1b1YIV
EOrUnrOHMoYEa1Dl+/RmvTDTgcdCxKRM6edXi5fs8VI7V2KZ/A6+GX/2ACTrB5smPaYa7proKhSg
Voi5vdIzW1m4H1gdl1eLVSmiBfZasHORQed262v5H3Zq9sfqeaIS0pbJVB6y4XwNp+CqoTJeQrPt
zk8dnx+NCpU+vlH8PnJZAdg8zCPsxbRjN4w7ZJvyyRMMj0h7OWFWmb76paTVrF8Oum0xHK5+uIY1
QXXeNFC+dgQ82PsOE1TBucZd31IFkwy7MwVpXsx6eD3DVugDI74XblLkg0Us8GW6ES3bhwbTDQ53
fOven+3yvlKfuc6Tega6sfeNNazn2ExM8afT12dAM8ll/Nq8Hz/1/FOg5yNtxXJWU56ehOUE2tAf
5HL6T4SsyWYfa215yMdIB8rzCUmroWXMjRR94wPcRlmzAPhN2gAXdfD5GL28SzafupTAiJUK9KfY
Wp8Q+xelp4UajZ2qDhoY6wMsfTNcRfiC6cMeE8wLJwO51pfXKaosEyaOpoXKbuc3UNOfvj0ppdbH
6RvkWXJ73xKm/kzYMcz5smaeQpIJahV8WanKuRIIJ2ssZrpcXMOvpPeN6PMFZ8r0sVqstpXvrySG
8FHm2YQ8Kg5UTqhon+AAFIfET4Ma0VvFFumwoH9NcFZz0GsnVe15FRWKZmy5iOB5bNVTUaEjF4Oc
zX2JuazuFFB0TifM6DRVvB9LaIFpDFwFWoDHKxxOEFheX4Ihdvxltwwkzu2iO5y/w3DQYGFpAckm
lYVW/QwCYSkFBvlBTKZjP3pKdQJoqGENKBVoGDDz2faDrRI0b+0MbPJNjEgZV2v8y1Mbt4XuoXyy
agjTIn3s1rFbodYnF4d87J1Tm3wsTPLtINad+ghI/M4pWOB8+b36O4Sund59OUw+1IWXakgp7H3S
vu9SJ2knp6jy3z3YbwWvg1q7cIlkSDasL8xYHHnrTlF174VrR2u+EYNKCJaEIga7xk/fkN5QCsZF
WkeU7H6s3xN2gqKJmxORRJp7050gVs5XcT1yZMYrhSL5AAi7ztYUzBIrJJT2uWGaRlXG3pxbAyAz
K8Z+fPdQ9oALIyvu2dPP5AO8qF+7Q+nV+K0LhhOEZX/+MnbGRm+wCjcwkoJLJd9l/OUuObJlmFoe
tCyvXdAe/i5uUuP3dLUrrzBTj0IlG8OdlY7nlTHRsu9QbPCyeN10MItUY54EqcREBwpYzOSEFnjV
l2/jZUKIYVmGULZu9hlnvP223rMVz2vzVuUBrny5Tl4NT08CjsqlA+NODak3g4Ur4qalz5mDfxir
qWQZSdHVhWMznxaI7T5PLEI2gPBh2vyHVSiWHGhFkJps3+Ykd7Mtm6Ne64dIYlHG6ZaEa6TVQFZS
QS+MqYis9TA752/k4QCULbQ7YXSdT+/k2ZYW8fH8eXzYh0CbmlT0euJblEu4BhPzCTdCXHfXSRkY
lPXVErjw6xf6fFxJrll+RmiaxOjLM5qHTNcUo/iA1kIARkH6MWLVK4AGzsW702aJhAOxrDFwAOsq
P1HjMkdQl00EZfF2g7yKiP87Xo16RWlgQSy2Pq6kv/gb/M57UQUeeBLhRrhdsY2GMtJX0ZikqLbv
uKi/HdertCaxAHk/cFiEF9A8yiclKAtF/WG8YU8ws9hXermX8HLpXSph4MrvFdMI+juXNq1d2GxV
g01EQt18u6jk73be5Sw2h9S74wJ0PmIiUoHhUo9svtqjXK3opCNJnQRFz3UB0/kibKRXmbdVuffx
O724gLqjGEaZS14YC7IIHyoie+qyMO5Jh3/0M/tfOK+5xSe4F8jwttn1ir5r3W82W5+IJeTeMbHa
bQMyKflbJm4cjy2zQW6Y/p/AZEKiuVUcnYIE+EmHVhiquI48xEaW5fRHQI9a8DgdbgIlk9/X5vz/
NhiNL9uwMYTt+G88k1k9BPvMUgRhMQVzaLEtOOSNw5Xwl1gAXpKqhUS0ZOhAaK9F3d3F1yE2iy5l
OM1be4lLnMSl2I+rVFfeue36sDok4+spm89Y0UawWDaSE5oghUQhQDdp30+hFnEBirOD2cEBAysf
zBxKjCDooEwTvbbeqaT7XHYv2QzlOmDB6VStS4FtgzHLHr74YyY81M8dtptGcl7IhEH5SnFnx/uv
i8qOCYvdyELVz+IN5kvTyw8ViRvoJcyyxcGqoyE7xTh0HTSzvi0SBbRvf7/waemsZKBv/0CiYja9
8cF6Vst+ajihjTKRRU2Z/rwYz8F+XNhQrerj9ScNE5C2MBGpG3LJ5WhidJgVyWvC+7IFj3uYaG+9
PztGQMoCKFIGBOGmuegsEIRLSBMqc0bbNJLJOKLhngjcgp9QXeugz8psjLQjjWLCiXY3ZYvdL/Gm
pv8pUOah1Hpw1g/UDHCJoDxN4+TPyv5Uib0+4cwIOODQpfEMUEcezUdtB/Zx/vPpywvHbNb0oF/J
9B7ovqDsKxWLQQhT2NuZ7BR3QaTuykxbRor8MSJdzIl0DM7Ps++DKFm5hsKFSZ8ZY/avljf2S7BS
/2aXbjoSe4EqzK+35Ra7R6sOr6VzHnvvgi0O7Ej8Poka8S6qdA/9sGA3PSe9qNBobddJz10dYAdV
gQUyRHyaSNWa6fC+RDm84EYndmLc4Ucu19B1KGu8wRQgDLvV5MffehtrF865NxF/0DXi8ikzSPQE
fmrlHe1sI52LXP1nVKBOpvIfl/CCmA/vMi6vI5KGKGHffys0RvNSRJymxCYaiu80nNB3b/V8qQ3f
pWZ8Qg9QlvU+6NpYEzKJAyBDOwdu767vneL0VI3XGh+jugDQTASGjULnWt9KW4jejzHYnURg0/LE
0JSbma1CRxdS5spusIrhrZxv6VqiidM9BGrSIY3P/h4oP/SDcKYscnBj7iN3yyjyps1CglhFwmoo
Gs/EQT4iTAluhC3gbBhcRGDoNJm5rA5v532VjhtjL5o3FtF4hpGlCfsXZLTyLZgevykVKEb2VdRO
tN91+DxEz5SbQ1Z1Zxs4PFh5+4gExRqjl8rJcoxxHw4OHUmrBxyG087QtszqnsGHuY54W/0HOoUU
S1d2WrKv9YzIjkFL5R/xUFLbHxtsZ9TPebK4nD/52E5mIubJtcs+LbUQVey4lRhJbyH7wwADfnkS
v9nzpXYfqlSVu7gk6xzO7Eshgkhvyg8BwkXy/wbviphSOpXc3A1xnVPW+zMEj/HfQfBG/1tal/Nj
4ewepQEgdWOiMQ28Rffm+zVcNUqI3hHZICxQ9E6Y5CNiGuIHKrpmpiouhP17EnnMgjRjmgeZeADu
jZs0N85cKPzS87NsKGqOBybaAMW3XyrEz8jgEUtHhF7fyOvY17BwpzzDuAFpFfb6uE/OJ9jk62z/
VwImgCyHrJoQbKcSYPhE5le46d5qZy925+6W7d0prxu77VmtvwZ42+3XbPipWbQGQvwMTewAojT5
LTkzwBRBXynBlFei2wnfrEno5ZDthiLWJTtsoeJ8nc0YiYaQZRBrTQXsbYaqlkbpMW1a6N9jDwEd
Sgu97FZM1UmuPI2CL0JpHZl7yz+IuBDqPd3YZNymIlEnnC1GQ5VebqFtCFYSLpKXxefmzZR9oaTZ
E/rIxCiyfsNRik6jli3sv5FgvPIVJFTPPaBr8MABIGzMlVrF24NMOwkZ316M/jG38nig9KlyrPt0
cpG9lOIJG3TeJDR4mfbW/OpiFjePu1agrK2a1Obup8PO/m6+OL0yhIpChzymJPyOWGQB4vJH2+sK
pDN4z+4AIi/dojbshNeVUhiRE9uCwV19JcUuttubAwFMj1kiyiU6t+cIx+YHICscdYxtQca4Q1w+
AiDLHkkW4LpALwkmmf9VY/agYi7V2fKz701ijwX9otJSAjy1+RTZwLvnWo+w/Ov/Gm5qNmOeWJpo
YfzNtYbPAub6isVtKArnNCNpzOsYRyDC3FssPskfOwC8AKVT8OUWW9H2BjCeTR8j/RF0Z1Gjt8AN
38wdJ3H7o+ftPskRWPb81uogcbAZ9sbSFph13zfswqXYKG11Nyo7bv1Fz9bzfHqbLqlZxZEN4TXO
4b04WnkGtNR6CtivpKhqNroxNiYR38HBW3JvPw+mpk56NbQOL8xtwws6zSLTFaerE9zds6Czuprj
gODbnGIQVhfuKXHfNzH01+M4t7px0HzhGYabh92Y7R8fvkI9vuXeGwgFPCeCrvFPN2r9GOXA8nlY
HWVYZF4WO320ddEF4Ibqb5OfIf78WxuvT2W2gKTfd3VAHsA/TAs9siMMQbFEUpcHjdFevlH5QyfD
KJipYbrz8YBKX63au/M25Jwk4JQV9kNyM9QTOmFl4NX6T9dcplnsU/4EHDJFWwDiZFfBIp5Ahp6x
tzUiPo7hek8iSeDGpDR/b1aHsUESSF17qC3cGjFnXlWWy3QcTO7wtTLfzfa1nqRmqnpRRVt4aULb
jqZ1juET+QBDfmi7Y24x3xg36GV5MB19Jf17uY/+XYmYxoV2PRqGzYcPELyhWhpnwgRXZRZMLZ9P
HeULDtTzaQOiDG4HRxlk7dVGBDpSDN11ABFWqkOJ8bWgEx+oMFzV1tiKeKsfF85HIbF7W+gbwzNR
Cl923sZ5YvX4v0sK6zysAaRVqrlHzCrIkyNOQT3/vrsf+O6lEFE3KSRyiCqPwHKWAlLjQT2UqSZP
mcl9rXPFVfrvpako9xp8YWrpZ9SQyd22c4A3T5/YUtuRVA9pB1FIV0kLzp9+bgQViWyGYfiJy6xT
8ePU7csMY7BJba4KwMm4kng8LCM5+JiPpKYYzLEzI4remFA5yINmG9o6pEP6Rz5+2r4f1ENe2K2M
VRctS5ffE3C0ZBZk1Ed7EUORINYgU5qgDp5zH6qk9M8jWAOqqtV1XKAdvsZq9fobwJ7lbo3MoRmr
Ejteh/DZ3xkJnhBuZJvOku8YM3wIr4Lm3O8Pmn/50YCDLfJ5T/2fKWNZVvdL/GNuqJQexgDG9swx
T/jJ4IHywUml9HFb8jQ+QXGvY31FheQVzPP6P8b12PL+F7YZDLOAmioEJx4KFoPhUt5LxxTH20l+
Vy8dczU4UTCXF4WTNbJICc2g8t66LTknLnZQCh2KttLv9516pQctaA6pldWA9YaGvjOj5OEustvO
dLAR+TM/EWS3Yq5FR8/oY2ZLXKGpSfO1YDPDlbVqxZuuU292yw35VYtMAGb4gBKMQYhJCAXE4MvG
sBsLjUuFICH4d8HNY/6/l1ICB7PQ02+h6cFU77JcYPloNyovm7nvznK28TG8Cn5wgaIHeUD49dSk
wpxnTATh5+ac8/esudbTXOxpKo3QF1p6/qkNv3M4IQZob/ASLkJRai/HGvY1WKGTWbmyyfw1AQnn
Moggvd4q+KqHi99oax3zW3hOJgzlP1MbZB6vnoX7L+dQJH54UPUXcYTbjZAoyUSfhl2kSzLF/So9
OslC9/Q9awi5a0h0hdC4SmKfk6uynL5FlnZ5Zq08IDy8iKAUO10ZyyFtSLii/eB8agnKBd6cVVkZ
fa/gFWBjnhSQlsaBdTobys5lB8iycCfILWE3vTIwu11rMeBa7U6CEcfZYYqeWvL6Fo06SEBFVuKZ
PT5Fidv2eIaqV/TOmrBTYJudlauOszQTekB3IsESoR9b1OKlhpKX5J57awWWRxad/w4e+hyn9sGz
ILI5JhSxS4xIOVtKCgouFDxNEb29ovk/qry2ClWfnvjvhKH+BXUlwo6kAQcmoXNFq0/ybGcazL7R
ik2A0ENwpYj+cCXRDPDRjWblfb5PNtjwm2s7O4LUB52YJAoU2ba4eB1+4CdRfeE7u5etI1LIFwoF
Y1aFDvSjJddx7V4I3lwl1Jggapay9XT87n6fv73uExkul/f9wRrDJHFvBO0PDtqqKirY+3D74Dyg
RRpHppmFnjgSiO+qsMuOhV3CXc6q7Pczxk3Ex+8zj9X4R7X6HA7wmuluAaRYc6qYpe653BX36aHc
OrCEFCHXcqlpMZFwUJ5yc1TKlZJHbPovP8iW0tEi0R3SSLfMEoMzJBGOql41eU0jAFRsY0S159t8
eGHrsM+hnHM3iO3VgQdvi+UKkMM+9pdda0eWarsmlITK5tJcNZkt2kboH3XqP+ueFCJPWOACXR6D
lFBFrNt7wVWjmghZ9qOZzNu3No94RyxTnkqLn1QvAiN9zxnQxzhxSXAZ3UjHgbSYItQRLsDlQN1p
/l80VQq75B1cGZzw2jokFH3MEyrjZ1B9+nqID5DL7k3XmqD8M8nxpLJKJ4JxeEYwL4xFRmUgeZPK
L4fpON5o+3WwvRcSpWDNI1pcFdMLjbzhHEZm/rugUoIwldAlNyqbE7Wd1Zn8ZVU2ZtrBSZinyNc5
tygJZ/nIj0qGAlFhPOEvnp1TN5o7So0nC0cDN71Xe49m+q60zn52m5f2EJIRI4O0EzMlFqYb+j9I
eCjAYnDZYFIqyjb3OYSKvikRlDTWGyOytA0s5P2muAO0sCJ1dTmdyELJPYKJr1W0GtwUKeYvIKSI
9DG3noYppCdSIhFg7/0Cvti0xwkJ0p0YP93TQNCoLxZON9J0ry5AX+hCntAUbN67ekgD30CbXnmR
s/nIdG9PSyAe0vqcNWiuq1MkVviJLjJ7JlAYbfPpSb49n6ERJ6kFb9ACsZW9GqgqVlry8FuWw4qL
Nu7zPbImmczxxPWex8qn5jY2AvWrnP5Bd0qhrabmdvzrQBpUdE8Ao8yxxCpKNlQzwRStfU5P1VRY
cW9nSSncxPwuC7HexO3Yzwrpkt/1760cL0K6KX4xYDwnGf+oJa2vSRO6sU+6xTQpWbz9nnhCOkFd
EQs5nGdSL+mZgBAXOT5M1degBowFWPmk0vt3+7l1b5rUUazDg0+MKXOm06XywB7t7gqL/6CwwEV9
lt8dY0ixuPGyAWvfe8ADC/1YFHHdRnhNsvhbBAJe8Ij7EQJCkqzS2vCJKxLHgne7XNNSKE9RwkIN
YYg4QbmZck4d5L2vqGsTl3aIK7WVTJARpiXzqJ0wgkZWl7QfA50JqwiMX6FF/R1rsocnduTXGnNt
Qw2B5dDL8ouL4UhCcLY2pn6u9/dGG/dcUVHxwKpK+sdIdNBddLNgPBxughJZ97GDxcctcQaw4IC/
3LSASwnoancUF/Ca1p7hpSGVIlW+bTnhwKfR/3f9bKVPEIKQpjkXEIQl44fQIZsN39PjuQ6a0wDW
i8Uu4fVqmM0+jzAwUYlOagP95mZebgLzIMLq3w/fynvQn2KOpVukjrl1jBtgfJlKWkvniBeumw3v
+9FK91xJ1f0SGVoQK8+gsYunu12k0lbDPVYqdGcgVQfUi9A6k3U3LBhEPnMr3eWlp03EKsmzknIk
f3S4t0R1pXBHbWuRWQwcrHLUDYk78Wmxb6/CNu21hdJkocABQl3ZbggGCRfwB6RBIZh1zBiZZYXs
KJ8B2CKD07vvn6fSxTR9df78DLhYuxQgC5j7bAes8iH6nVPd+DIXs53+Aub2aDX4siy3tMpFhyTt
GVE9tu4ptEbe+dnWgmSKThZXTaf/xLyVlis1d4rjol2XWxS3CRtmAYT37bm76f5+hzzksBNnItSU
XwwRzUawcVfiWywOYHt6hiJgDIxmg7W/RXoQV2Rm43RbV66qneLS+818kZmCd1Oq1p/r3H/KV6TZ
F3ombtV+5ayBOzieTKCSZXu5lLNDhiYlYjVVqsS/dopKLAmHeLhI5HBYs2Aza7g9NwsO+9IrkyPV
BV+1+jc5Hzi83sMEBKoOAuCR2CWgLks+L028VSRHxbccInFVbEFeqeOv8/CdcTUiZ++0fZf6j757
VqyFgKu+V/EsfbdT6z5tQHJTUSUWzVTM2gmfYI4aQNWzGn8xiVsgwKxACiJTBBv5cwDBQ/tTZroE
ddfDiQBctwiYJhECG7PTcI5+EGkXgY5ioTBCUri9i6y775S1A880BEn9bAquOcq6zzB9ZwpGiDPH
xe5ZrVpCYTkqMCNpq9q2e5JNSMRb/dIjY6Fx2k/vOaJ438vTInZfcMeNpWVTKgVFhS+ioSgcmLJS
VoYbpMXIDYkRZOwjlG+cV/l9UJK1IoSpsJHSySztsnC7EWfkzhDhu7c+emN/9LFwRKBFr6v4FPJ+
mX2hEb4chsgZRjIR18cq8wZcwyHIa4fv5HoX2UOa9u0jfj91Hvp10kyP0GpfOt+qzyBgl2dag0jO
+spwoeePl5lWf+6hdc2PoHIKbhDbKsZRDf8in731G5hGrO8cvSD59TpOAk08bZO7a1jQqjSElmAV
W60CrQiaz6dWVDvOgwaUvh+E/d7dybd4t3clRP4n5uDBVmUeLter68YTbdA+NqTG6VFLWTCSRytd
WEqARgsk9fxjp/boJNUayUTvF2ZNoIPJYmqLiSQkmNPgR4gJPzmJLzyOa52PwWWzGiycS3tVPHSh
/ucb3JkmTvY+OwPtdbZwRnLGs6fWKCs5UV+l98475ikDXmWrmHWla2Nd1eBeG9BuU059gDGW+T/M
wrmw5ONRiePFf3/0s9URrYydQJ8YNVBP6GmnSfELCE1hp1gVBkUX2eQuIGP0dOFWWZ2ZFrvSyMDN
AU36DC30Bwb+Vz1Y6guEkfpycsCDPlzsSwBNiq/95t60xDInP1OSyLlRAOR46Mxr/If81pHtEa6/
w2F09/CtZsTkLuGSV+yRNlg6Yfsdpbh5i85Uw9SXYIx3hit9n5bY1HzgTnuBbz2dpIQfJ6yipNnW
dtNbuTvyFsLSOJYBRA/MlBvmHRRKW9AeKUghft1nYNt6PKCudjJFMzTjkF6BvEaV8ozYR8Yg/3DH
N2BjrqIjGB7gwk/hAbhyv9OJ3VYtDZFTyVGYuDkmR/erwEqJgJ02hEoB62ugpEtMGLR8sMPggiQC
C7JJyoFb3xBFjteN7yPDbIRpxU9L7gY/ME4W6JF+l4L2qaanKdkr3QEmUZo46eZVEXzwFL1wVfNJ
QG+kUH5fHFvxOSQmjbV0ZvCX0hmsLxlRsRRYKsK9BNtZwdQkWMjKaMuxgcXDtGSsl+9LSwxEPri1
SPpRywV2P7LPLBSPTE79PCDxaPZryYv2SmV3kfcsa8c9ZImEOZ7EFpOwGGGj6jt8rYK1Ay3irXwP
u1nt5MXEsTfHyyzVp8nuMG5HLE/nWqDtFOJWYARwIVP2hlNXaAJ+7vVg0nA7UIEEx158bJgufIwT
xa4990XYghT8iFW+hfH/j72YVSQBwKb1lt8wBqCBTjn/7ocjnoauv9B7ksq2uSr9pSJMXphO2hFK
BWugbLWTpHozSbaTKzGRipZsIUrCMbXNKnbGSxJfwXywCmEdoF+AiEgHAwYJH0fTfA7YHXRuXZff
DV+WJh1cJ3rLx6pGDRx2l/2i2+frLiktd1cXeTP3o7f1Awvxu1ztVMhu5iJUSMxWaOMMqrXduAwO
3iWTEr993mj/Df2DbuDR2w0sCTbf7MHxmTNODd02XmpLa7Ked/ZlawftW020GJsirPauAXQ7lZQe
s2uyoP25Wb11zKI/YVy5uS6S5FOp3TjIfj+7nQclDq0F+ETVKqCHDdKMheAtU8t4pMwX10lzDQIV
gzf1YAizu32McYPmFhWxfww8KumMkfwoQiSjfp+4tWSFIkE7p49+/X05Z+/zghTW5oBHkvQDCEaS
kAhnW/wV4AKw6sNUuFaMnN98NG/XTVi0B8g7ywfFt2ctahRvnwgPbf2qNuirQhZ6sIjkfHT8YyRo
/yBvyHfhePxvpfYgyUJlZTCmhRwRgLkeWzXHHKUrdu05gvGpxln/wI5DH2opfpPmkggJqPTIuluV
aCvPqZR/Q9BMnYe6ep3+AItyK3NLnNJVPZyx2rCXS8BXOI8bGBb6RUL/LwIOhX5cvJngXl5yzQQy
e+UH+FwK0TvAlwxuIypXT96jG/8H2Hz5AMHddIxR1i+XCaql8aQMHhcuSLDFevRR+jWWL6F7f7Tk
wqrdJsTvlVeG6bPkzci+TKrS2fOixfK4C6mnv0UJLZhEvdF3ejsUK0Bd9gfUZBPlyOnpD8e3QoP2
FRCJx/8ocJxW2Msoh7ynhZppVNu0tHfMBzi2AM6JSp98ccAg1N5vi5okPhKRzdfDzcXLdul1pWAm
iFTggABLF6Ng6DNANpNansKCblt87d+YWWL1Ybtt09H5qFyoJEDcQpLFcOnCQu1EsI9JnRSqXGRm
0Us3kyGAher5QrTcZ1QvaFyVlWGhXcXqL6jRQkuooA5CSSl7Qc7M59eFYIpjXN0c6QX7A3XyzwS4
gWQfIEGoEC2YCqBEYT4zyav0/lSLFa2Vs18Ut6oJwqP9WKhTz/Wik5ojY+DOfT7apwrOAUgJWL7j
CqfWbpO8DsDu60fkEroydpZcZxfjOFXyAZtPoT7hZoF11pz7tMISo7eAQ/plXm+agtzbYl5u4+U8
MUpFsCn9GrVpXLknfMUHRbShpgPi5MI5NZT6PDO0UqVvFdLuKoulXPgu8H2drhs/3D/YhjaoDiz0
HXNRKi+6YjhA2wOcE2L6WN0s4XuYSJVvcqmGq4l1bf4VK5PRIY25gdILeAioFDnKu39IwZtxEOoB
UyKm3gRJ3rToo8s6juNPe4Pdwf3WNvjHzpTySXgdpbep++0USimyvYkq330vFRzwGdJxZOZKFRKS
t4+z9WhmUAdN6UFeLttoGlIdgwIs3rURZT3C8+GMk3o5MfHpJUwtwhJ2luJimiGhh+piWbvPtyfg
iuVXMhOAbC/7p7YT92tA4BD2w5S783b7hfevHVUBsxbFmjSvw/le1jDClZXyyExRJFrjwTsBOZWZ
65W5CwYgxbcJ4q+iPQ/QVjL2QJkepmUXrI1Hzk1vnuEMEAxljzA6ocozZlV049sRY32xeTjF+9/h
KD0jfkU5jFIzGDJbOWqAYJ5jnruVtN2tIbPlikdimD1Vwu5ebxrNchuoLIn5o0GAv4Lz4W22A5al
iqgZQD/64iUjzagzQ5ER8dHvmAtyGL6P0XgmE4fXM2enljo+PQVuA+xfVpBqvNnVm6+VyBv/w/Dg
fEeB9oG6Y0oRX1CVu1EiylDSyyaMYsWRwA3rLZWT1ozChTjvqCTU0sVmCEg9Cboql1qkxjceJtPw
nLdedg36Ek+rvWqIK6QWg/n8mXz5Bj4NtoJMP+71arRaHVh/m+LfzXCnjazeUUSNuap/1d3SOnVg
y6G6VFiYYhDqhRIVaad6SyfEYvuevryFKNsfq5ln4KH1PKgo7tXKG0jmrw4RNXmcZHN+N0ieuD8d
JO7x4wyKVI2gnko3nT6XQxTvLSOVYmy7CttTNV9OYB1dGwseQkXJ+gRhA1Eiye3K0/Nf5R2Jj69D
eE2ITXxlv1VESiGTbMXeGFs5MHJhF5DZSNOHlDEzufzqIthX3ecyiimy4i0raI5/fBu69kkzyqFL
1uD0rtDIHbqb1NLmafnVtkVEYprFSz/9VX6duY84V+0uZeRoTJf9DtzlUzH1WSTAkpf1V8SXZw3l
7b8U2Lo7t5Tzn90LYUSe197ody9tnViVaYk0iduSzgqsIz9JDg71LUji7KwsvpTNMm1xSHFkDRRp
0oxUNKFUKnBRVN2YYoALDNYRHD3kh97e6BKLd/aag9OQxSW0jTIPFr8i9neXy+ymHFvvldIGmnye
pN0DtxY3MK8OzkaeiHv8GdIXYXnX1YARLwPeVHenhq7892avg88VHt8m4ERruvhGlxlRfhUDMoBR
bC1CbJ9NucnLpYWPNg3ism29+scSlDqoQ76UdAE6vjDeW8jDjdSyepfCNKL5Qu4XO20EEDJ+m2dh
ciiXs/BjKV/E3kNMCDY7Lt4m1QqeasWL9XoQuozOHXNGMr9/4OXq8AAuhEIg0tMkVpDTLGyxHYYY
gWyrIaakXtKwX7dwEV+CVbm9mkY810M89h+eOSl04n7ZQh7RLU0jK5ssuI4FDMiReap/GROPFpfC
YcGd9/DEmEqbLZsnXP0qqpan6suqTGEPsSMHjLY1fwD/tApwdy9sh585cTHOVjZHsF0RyH8qD0CS
+d4XZd/JAkZOAbpejDqysaiS3YrZbIGzrv4FeOJZLpguqMw68wrd3dSaK2B7eVeEkQlMJR2zvwVo
Ft0gQbGU/hi7X6b21VoAi8rV/N0waUf9S3HuQtecnkg6R9Nad4kpyNRS6qruXi18oaTbsNSM1IoP
EipzrymJ1wMsGrhYtvVPrBuleAgVP1k5WGVVOXOVkak6Mn6RHK3+dDC7xhdfao8qCeYi7rpJ0Y+x
D5PS4eRm+pPKk5MfMzXZ10p431uDwX/cMulEM2cbwod5e3Aa//tsMmU85bvVeqjeuoks2DyI7eaJ
iWEFSinKYpFaTrv20rLg4NJ9mQMtg/uqhWt0vdw0KIOctZcc+inadd1fO/PKQE0bMOq2rrMW0ARo
wFcG+mSJsnpZgDuP0YXIeaxEhJAgGJCKbW1re0i9YjfYZT3GbIsRpQKJqB57o8wt0oxPTZrgz99R
QPJ9OqhDLepgoVtcHmR+7r+eg5d6pAZrxtCeKhLG0Q5vAc4vytOD2meGvRGuVlKAKVuBoXUgEvjZ
6RLL5lb06Kp8sUsmxsh6g2S3xqgAPE0f6OgISMjaO3LzIVIDFesPLw8U2EEcXzvuDqjiFr3QZ4GC
rJxnDqifwoTSqQTgdmBWIWIFeJHMBnc0iuSWXEX8FyzcoYxQZ01QeXY2yy2ct3+i8hqomRbqKgSi
K+nHERrNNtIIBtqeNRSAdykVMzKOvaeGw5bjO2XDSv3z9sTjZhydx/nWED/gfg2CmFWH0xKfFFsn
cZ6Xx/fyY+R1Br0fgm9SEhzcoyKX/mlQX2JcU3xHj2COpezauGhAu09ziZR4JwjfweccRAKmiiRb
Xdh+hAX8XYs/E/Jaq8Z1xOyMJ7E20uW7VYXNMzIVaxd14lOnxqhBYASYFOtJMFez/TKA/caZPGHm
s2Tf42wBBOpHRDkBLNp2zHS8RLyNwXruQa4MQuwg7y5dm/4kIcfNtqUPjmnJGS2+3M2b7HOEsGjO
TPqF6MnTK9oBtTguZaGZcUPBQRa7tPCedaKf9VD/yXh2bct/1TpawhlE48DQ0Y/AuCAFkbcBvNXc
PcruUWHlxhezVrNXb0/gilpRbnWf8gZjv8LMpO6RgPaTR8BA3sadMB+8yhhbAL7bVi+NXmUmniAa
zqQ9L2PZ/ilLP/m+6Rxvi3gOr0zJEg4SDuj4aD5kteVoPWaBnxANfa6WzNtGGLgYShklxW6rQ1ol
uFWbXrBBwU4V4hv8ig5IQZ52hw+z2+P7JrGZPzvKIALhaUNF9LIl/wH6zseo/ZDdpZmuB4ljWLT5
+DIvLFsBbD5csLu2PkCTSTAlnWW8Da8FALmky5lPq7y2azG2Rxt9n7GmbGBWBU5qqxNB7QQnmca+
We+e7/+kLlmWLNEGUUTobUb5jIkhLhijDnFaDgmN3dhova6g/lLXFLrXvEfXKETi2gHS6mONnqEg
cJTwLWV5DQy/IeDRsV9QLzI6rIlrmSED71+7YHKVTSsxDRJQwDsIDivlKL0+WeN7WKsv14k1CTWT
SAJSrTYqfLxJxX6Bl4OMpMuHAWT7+qnzj48WsFkZGhmis7GllHq99MlwEagawu5w1K3iak9Aceti
OavOXXHGTYHf3T1mGdtyt9C+j80xrv4qlrDlFkdyL305DpaGMNyRaf3TdvlAoHKnOd2RRg7B3/+8
JHeJoR5JIhYzhIRn9b7gW9rBJLqVqdsNiUwmi4jHkBqRcRAGXsaKRdOjapnYuUP0nHxeixl9s5m0
FykkQy3QNAr90NZsQHrwyO5wOdd98mlbHx4GfFxTmLSE4Q2gk7umeSbNviUxlCffhROLpi5Ajm/j
S+SdJKubn6lSdasz8UKLQadzwkcWtiD3PQ4G8/p7LiGbCCpOSteAWbr0LZcodCZ8lRaK1JAk8Lt1
kpqLiD8ack407ccmyyEG1OYUTy0KcUEwo06n+748vDATOyjpkHVhEvZZzcBjnCAK3JWgHer4Prqc
gaj8kw41UpvtOSuLfsEU2m4trqEFSlAt8hRtuySAiVAewDjVw2mhRTzP6ulN8rJry0YljswfBdG6
Dl5kJ8e7ZWnqfjNQREzXF3aZCUeJi5PlCt5X8SAmLOpf+3pJIhfMRN2Lbms9ymmyxlKs4Jm6yr+s
4J1V4nDH/cXsTNku9EWfk9tRpe2ykn2AMv4mEGM7R/1AZ6ktv54un0wY0E3Pd5nZ3/ZxqdHAVxoO
YaORlIzvbjWK4EoPhShNLQbmK9bhEMpwPtgLdN5heqb7j5QHwCkwFXsTKz981PiZWjOeLSnuAptV
yS51gDfwDMoDQn1KhF/Dm0ih4uOXEWqjnIC4qkp5y4jwEJBd/Gb0xgFwlx8T+YIRTMogWgO3AgsK
x1WRHfN0IVidS/KJaL430VpKsjZTTRN/mAlkusR/6C/RbHBHA6rF52bbOJ/p1SpHHJ/nLDmP6EkW
gGbAC062xxVhx1LcWo07e1ut0g5mMfVaKCrHbTrJgppsnApVIMhsqSz1YUzlwwpsAfwz62TpX4gd
bhClSTmePA587uHY7qu3OvrQqTTEN2/cDuiSVxTepkLn+QJ6TzZ6HEPJDISX7CmmWNYpi65iaf/w
awBeAMMi+8FkcMX1vJOWltNDd7+Shy14aO8RMQDTC8ftq8n/TFuh5Zu59ldAbY604vVE/hGbRsg6
GNefN8WJX7B5qL3JelPUBx6xHla5EyEbb1YbhALj69HP+1EwRZy1faetgAvfi2TQAoT2xdqHqDSr
C0H/ydjGDhdTlFcwZnVL292+YdLI6ZPv8HKe2VbY3pxAAWmqHvJQs4VACVV79edI71Pj4wznbroK
fEG9j25tb/mD2W9FLgMDdPoTHdZwo74Lk0vKyRMI9JHNvPJNeu8JtpsTav/UjT+H5yXDRH5gKO15
i8Ef91Dpz5rYf6X/A5azPkPk+ArnFMLuXJ3zOpDtf7uq5h72OlqRr9TpR8l9eK8FgZoLcLPNAT3b
2663IB9vbsoaMgKPl3T5DhbXqC4oXHvd+wcKJXQMVp8BJUrfxxE5iN5F53RUrpFAgNmX7K7wRcTi
nJMj5A6yeVvq6Ur1Q0S37sBDUakGH0Z7eJA7URfXLPN2b9vU5uIZTHILCpJX4LD7qAuWqJ96lc3h
kWd71S8fDTAHSeFNN38H7q1/08ZCb9RMGwG8qZqMVe82erNp/7iTaKd6pfm5IR/AZj3B1k1DPoPc
GQeIoL21NMmpYFjfmsfKxQoNKDfKNG/Pjzf386hVkUbXOFqvys3ecYWsBSN9X/x62obkIAnlpR/+
oG9xrssxWGqv0IegLVEwlnNTEt4c+AoLOJ5w4RiQrx18Pg1cdiMAE1slmyx9jQ9VuFChxU2teeze
RDYv4AH5YR1UDAfGbK+709jk9GQMIuqHOkyO30GSDSAux3DxQ9yjJb8qPoW75i9ijsJ+sDoqd5AL
oxtObeXQeexdHgi5pv8UYtW71kEH34JitOBt1gn6a16Pl99B2vkxq8RFyJUfLVYe+hlKqftf+F7j
UTQNB/SSnaBp0NGZubmMdM+nGdcOcDvaJS7pOILB9xEZ0TthUWB3/HNFcjMUbsBkpLTwM+DG5ubw
QXB9y/P9aorw2hW7tHvaMG/5iBqbez/e78pA+yGYZJJJia4TSRR5yPQiepwXJuH7bKUWorjvjcuQ
Hx5XBuNW9vvj3e6aySO6Jr9p688BghEVGlZxzBpHwCBaAK7xwnkFxPVi5jC6CFawzljCq6AcelzS
0NN2C39pgR41wNZczwS4Ht9+eNvOXOCUj9MfVoBat2N/qZ/AJqQ5Udt7AwVh07j6UiUpTtZmerKQ
0OWHeoxRxupw6HyVcaXs/zGa6AmqlrvbwmLrEgsSCaXwNo91ZTtlf2TzBnkKNk4Gv5apFd4mMI1Q
OOdWw/BZVdGcQJUlYL//dV9L0UALwyKxqjQaGMrFOvO0iJIyf2cVW3h0OgKw2bKDeHK21EManLym
9LZjvsMM0QP6jRnkLpyMDUitTU4K9eKKTKeuxVOH3fhrUdgEdDXK5i2rz/GGWuK1fd9MFk9l6Nxj
kajVePZjGSLQJ5FrUVO7wA667QmeaE/M1Ve1j1K9894evbNnKpVr6cL/iE5Tep+R1LXV4/fQZ14X
a88ykN1lc5KLvCI4LALxUtRtwm+Mw6n48yTTNA+ySMr2tlouSE6kuOo2I6yjZpZCJTgQ3E4rKKtH
jLpSGHrjhZwnTQIAHbgYDYXHp+9qMzL6hZfJ6J0AVW0G0WetfTbvIXk2t5KfW8yL6WebxNYUesTP
0N5epx76vI4hh3av+DHsmqYa5nMxxtOS4R1sFJl8GAdcerXgbeCZtnwTGfWjd8QhrU+3sKdTj1fX
0TzVDnaXOC/XOiud/onJCMNgyMwKVmyzvbruORWqh4wn2YaVMIjL4upB/k4ojuDco363+FdjYnsi
LGpF7l/pYxFUM2fvWnCYUIVJhvQHzo5HZT2c+7AH8J0pRhDXE7mpmh6coMpsQJHsOCIsxeHlP8C+
u6UHxgKy3LpzsDBrskBgfhZQ9MGC7VF51JH/Gef9KwxWa99pndRPbiKSvpVKD/IElY2+9XKlYYgW
2bEJws/xWmnPkrf6E6OhOCrt4+Y1+tccbo97Wf/1AftkaLTBKAPc0uAA3yGFG0iohLFWaix3R5pd
1WlUFLcKoNNL2FrNlV6/mJg/kJc3nbreLRpxIiDn4phvGYmfsCYBheRSuKfKpLDsmWkrZsB16U2+
P8VqsZzaSWRP9lTsJ3aHOvbWoeEwHK1dLho4XRYRoZ9lZ7PcZYyyD18jgfqTJqK8mmFjBA39c3Ni
vYjzlWeJSTPEGZJsAGw7s8noxsqggsoD9KlP6m9rdYkF235rL4GbCUiBozCaTNw/jOvWMqHulQfl
xXbhzyd9Oyyotcozwu+ZMIMYohjlQuL2jDJWhXAikyrILeQKm40wxUU++LFMzxLQbZ6eTKKCmuGb
ksMMvoXNtgz8MqPUUz9K4JCDd9K5bTNY0D+sFkD3fj1xop7s6doEOgGGh3idO+9AirixXvxIYb+0
pwZdHT27vqboNsif9RhY9n3Q64DRYo6Tth/xig/6rCvqv9Zx9N7suG1Mv7YA1UBs2FCF3PVpJWGd
uVSjcPRnPxrLBB/+f1Ug3H0Mb3LGKrXV2KiZQev/dfrhQnXjH1+wFqZWclTIJyDGp8PAo0vf29MJ
pzLkz3a+c65Fv8Ou+wSvf75gQn8HY6+gzyiI4Os/iPADjqPqYUb0ZxfpS5yoawiHlkG769NMyiAh
XRxCdxZMGLrPwADgUTPPWmerpXT0CnxBHytUs6yfwOV/LmceBzsDhrtkwbbAyjPK95151wUpg8Db
QSUpQONMoOO6I6l71tRgPPO/3s7DJHmS7lBT71Ch0J4m+ePdasI+KRSmZKdkbWob92rwk1b+78Su
IapsccY3DQs7d+CRge9MVLEJe2X87cgnW7/tJltATptn6465Ip0Co2MoiT7bB00tmo9wO33jlO7B
Dh6scJpcQ5js3/XuHqQKUQZcsx2gbbYFjM1GKLHHRwGZe0mgM2bZ/WWGUwebmXKPI2PDuCwErnRq
cjmPl7hEcahe54i9TCmVaTHCXeSgy61GBm9D1wiLN6y0ihnLPTHVf9jaEN5Ee0Pv6NHVLLGwRYQt
GQAKKOPabC6cOU56HOw1qIt3efI8CgTR3RfeZDqljBShi8UXNUieHWp5wQqtoLgXherpHFxeo0NN
+xTUCYBSPmrdjpQzipv7zO8lwxKgparfCrYE7LIGtC76cxeCrCn9taoAm3EzMdqBIlU258whyWkD
tjOSoOJli0u9eYBElR5By2oPdmiTihdyXLlUu876UNPVb043TvzHV/fRLeaLvNIqiufutBJ9vUK6
/Dh4m1+20JI0DdoEdCvU8tiQDe8pIZWEIe8lf3Bm0Z1nTXNgdNFNxFpI0hbLvzXo9+2L2p6rZlDC
XFmivBQ11lM+8vecTG+ntMlyI+w+ucMmIMi2DaY8tNUnweo8Ochhq0QIGQZG9tuXGpqVMF+kxbS2
XVFlmhNHjv3OePc2QF3JKhbcZwQ1XspNsg7IEu2+s9Oolr+loCVSKGx6hmDlRtXXWRb/N/yr+YF9
9sbSAxOhrDAkLY/gV5baxPxVsuyGbeRTNiglWAQsHREfLT9t+e4boPh3V6FC5hp0Ny2Uy0kqR72O
yS0Pw+wtLvkXyM6OZpKs0uWXBhTJtI76yzwbtGimA9Lqq5b0xWsb6zc9JJtmOTtKkAeNjYjgeB14
3dyTqeIIo5DCPkuDLPpPn7rZw63M/sd3O80wRmyuq4y+EOgLaNE1kAGZB70ZlM/NtmIsoCjjGJIT
znHOSDBrHHV7SIGgJvHJRacXyONj0CCeNSoFWGYYLcjNBa/pZAWPCC5qW9EhfjtBHIqjXASOwSF1
WVN1RW+wPseuWj4T0ixzZP2kCMOVhmJmF7QOnNV1g/Ze7bLRxJsBuLqKV2HjV+YNK7yivjNoI7+S
0V/UXoq+OddW1hCLOIBlJxmMHZFMniHHuuO0bzQLoxBzD6w+s5/dMi90BOmhlg1YDt+Wx50bil32
0yWN2Cu/g1WyovDwIGi09tsAEw+klxDYoPdh3No4y/UFOCLWHealmZdNcaS+tO1x8Gi89MDzYpuk
ODYUOUXOikWTtkU8VFl+5W/y8Epx1FtQHVYUFiKiudGUOFw74Mw/ZLVEed/QzpTjs/BlJKB4gcD+
jIFjdm2taUqJ1oacxJZKQa/eEfoscDaZ00jEXSD35m6kzJCKRKexxz8aeGB0Xhwk6JufWMMdPjHK
ZRQANpzPVxexlD4vYzNL6Po8j8BuXi1hh8zxq6LkJ72hVv3wyqj/p7D8MJ1YJj4noTva779QSxjS
wlDXqyZ5EAHUc1eE0To3kIczTP1mlEQqMUv1y5UgQe+pa4ptuXSP1/VCz2/h1s9ot8UyyOxbsLkW
+XNpxh1RX2z0hnltcWCF1oe+1Sj4pq+PzpfuDkxinmfOgkEX0gLYMrPVe94WHce+dbcFoNEBH+aN
plvuqFQi1M4vKud17vZVK/C0QDG6Y60eKQTkx8dAVL1JUrUG9rTs6+3pduBC8P/KnThIeT3K/x1i
IpI2RUkbBkp/FdF3sqH6aHd/IRwnpNW3AxUjPRiaLSzEHaBASXaXiDLhUbCTv9fRrQwEQVaT5yOp
N4f/XDn8MUNS4I/OHwLjRIqPlOGgbx30cWwG+e3JmwWnqVoasuQk15QrRJr7CqvFdD5oA/SxgU5f
BlVEfmvtGviWMoxOHbV26hiLXT1iSHeLrRqxSxqgQCjO0e9NZNo9TmDcfRuoOMDpcO/yuZ5IY3Hb
GsSN3x5tj8GoNPMa1x6vOJIIJ1qhEEymk8e2kAC7zGAsGsrbLsHqLZUrURBc9XFdfiLOAQXk+ZLr
+ArOcXIUaXuzGZentZCVi8sOdnJwX92451sa8NVkgTEcTZm9urPVFdu5tuGPp4TsSI0XA96obh6F
WSKtQkfKfCs4re+2Y/Lh7z3nWCfWebboOIPtozTqoOUSZgZe683dazccCjqE0Bpaifvag0AfTC3R
QSsS7lgnVU/LBvdBfl21be8cKc3XCARdz/NZPfTD5PHfNcfxpOat+1vkCz3P/mNi+o/ha7MeIKpR
2JF0mFQdmVOns2wBThqx4GrC/lLzuCzZ63eMoUImJdnEIAKvoEjjDRHQxY27EHMANMYVppfQG8/b
TohDYAYQKuzTR6MRcU0rXwRWH1GlNE0P8trDdh/oydIfh+b/gt/W9riNmhxz1M9MeJTXwLtQ9oF9
JtoEqX7KQAmoFLfGM+yHiBA0tq9H6ztRf6VTKlTSczTVeeDjAvO4auj79ydx9kFi5blpiXjKsNf4
UlSH/XUqPybcxrqPPGXEDxZiq8tMXfVYEE5foe/MRoYk/LtLIjEOerbjphc27huQcsFYwQmjpACh
MqcH8RvpWnm0yTqU4ml+C7fLUU3V/2/IuJRWsxfgF9QxqGzcV/0KZgeAHyclB5W8Rc0I6nCk4RGJ
JdGa78tBQ5LMdl8905GsPPBgFIznZAxMTBgX0Ffq8b8QVR0/fygh1rxPx0fdgBcvXlDpXnRELwWt
snKAJF+0qUVOtBejqGnzVdveYiusfCtDrHc5Y6WK6r8wURrOhAbO+potHjJXqn56VeD4nMdAf7Dm
/3wErUCKwptB5924XhqSXmzRKFZqOyeDzChD/AGTR0xVYcVQFzKm5tYroPG+66VjWvYSAWU2y+Am
65TDYrckUtS9Hp+OxiQh5FEc0i80SZ3XvckbUUup30ubk2gZYJ2K4oTAOwndEk6reNe0qEnyqPen
2Fwd4WqpRY3LGQYLQUj69NotZuHicYCRorWVWPCwbPXQRQIa0zd/UyE9XFYsMH0jQhS3J1BQtMB4
QCYV7hkpM+s/rgz4EInMaHr7IT3pPX+Vyp8rfbx8Ju7SxiSWZtE54VejHWxVdqbc/waScI4SCvp7
hHBfhyrRJ1lLbKYROkoSx7OeVxj+gA4Dh+5VValnX/9kCqFmfw1cg969laawUILzyx306AVvlfVr
pjpO/+qBhXWk6k+SqKAwDxfkL2LCC0+wEh57q8cEmCD5JD+gP9wME5G+H7HpcIOXs50izbLSOrsu
0TiTTUzyW/h/a2kr8Hq2rFovE+1lubiNN/bOdcY4pAHQRcN8BTsGXwvHlSeQED+z3BKcBJQmtSci
Aeuj/cKLENqi5R2O+QcnpSLh+zhszInh/LsdFAIPCilVeCA3uT+2wKDvtxoVe05w6oiGeAi48c5j
pusy2KRMPWc2+F00b3IgEzgX6feicVxEKa4RMLOiyP5oiZVRPyNdiwM0eE8pRf4KBqiUokmtI+VT
+n7XUA0Yv5YEF3nH5zczOM7hV5ncGrfD72rVkRZOW3cBB+HrJPO5VGdRzXnXNMmzMswMOpN5G89o
McYOGng6Bhf7xYRCBt6vfWNYfgEbq9IOEEy7KHoIvIAMQzWjmfvDQzs8MbfM4E6hXuLMD80kON4J
rlJjbqPWXhIAp9ERYrH7pgoVXTmnbbpwDc5aqBopGNF/haR7AQjJXb3oV5Bo1cE7zvpvniw4HLn9
Mxk9EgwxI0+Nx5VxKYWlXaNFiEQSkE9iAL08AKv3sJHO/wqatKUDJQmSVH/gF2v/RGmJpQdXw7am
qrI1/5zRzMxPmXJ8cVzSzw0Qxsl01GV9pSDyAQ0hpk14qvke45w2IJAdn0nUFm9d0h6k2T33Qqqz
gBJKf3j6BXDNPxiSWbaCr/tpQFniBGb9R4abGZ1OnL73OVBsDWNGHmxR3FOVt256Y99VA2tZtu5s
FaFLpX58kIDySM/Q4T/kvCvKDnlSmTK8V+CjFfRQA62XDzK5jPo17+TO36xaXmysZUlkHhj+IZ0T
zDYaesr2M3I50wexztCa/dJ994EwouWER1b+hermbjN/FN+lqXc4F996ZBUCtEarzlpcs5vYKTyF
pj7/rQrffCXPvcD8Lbq7HlWF6iFEARJ49AHYslCGmqZryjkhDTgbQgBPB27jgOd8aAjIFDkRp3Fl
jeuMBZfgpnWRQChP7uMIs6rAnbT+Z9GFllgqFRfYUy10GBnARgb2lUr+JKgcF2eWr5pb3NpkCOU1
7hi3uIqgzNSzmVQ6bETGTJtm0T1sRHfTpFGNM05epD1x0v3PmDcdzCByHswvl4N4RVZvmV97ZqXp
9BA1NmRFcZa00d0Zkrg7u5doOtXdJrR6U5U328TE7DQs80yyl3fqK4nl0/02KQjieXK79TjEpmVw
EL6khZpodNR+R3qCAjz3lqDx0JJVnKz9X6cpRqfWvljsZ94zMSfAqhVuotflQn0NHUT9M7Kir8Gm
mx2lOUqwKb9E5L1rVpPW1kNTfR/FDrX6mEfh35alhnzwCSchIzI73N3GMcytlx85jfBCQ8kNLBI/
w2lbDTwr3myUPhO5j8fUVMPFJXn7g4UfiAXeBYW4ANYr8oMEJxXwOJbwpMLJw+hCU10HrUBJV5Hs
5rsQZMuFFItlShYzm7oECUdYZgZ50n8+s9TCXXCxp7YdHoJifD8EydP9kFpvEjc+YI34vZHmK5JH
BT7k6K27lpLGHE8kJu+clKvXDWRUA6lEDlYiLwbkmwB3ZR8sjkay7NbsNEY38xsqXyr0c36rdJNH
6jb2X/PCROqDp7PGDHEF4ogpOSYF8BtSilcOkmsWZTK6H5CJjQ4MEt/uHj8UiqPeAGhR6l+hFNj/
R2SNiUVJVpznaDrvbX5nErFS1XB/lPEAHCvy97tmtBk0iSqZqm2jMTe4zdTIoxAHew2zFYwTg6O5
CZT9IqKEKgOB/lBLpFBOtNjIzfustbz+Cmx9j3+10ssbWwL5Xj5ApZsodt07AeEvsPr4ac+WIwVC
l4Vw3AKtSV5r0jld/0skl+iek5OGdJ/oapd9ZA7XuZKPWgUW6/1vIlz031cU7GquBzqyEcwY0wCF
P/yRNGUE0mZtKPZL6M8w1yVVnxq2XLex2daq8125AsCcq/eTRoRZUpo8bCNHi5mzq2w4+uklrAVq
hjvPEEwIg+VYFnT3x4YSsatKFJWqHq8ze5i5NVOvvfP5Os02CUcRMULw+1vIVMpTHFmeLb2BfDaE
2ZWPjGwydbjW4NnqYRd5sOfSI2wLQeE86QkIQKGjUUxxM7nDjsKy/TaROkPTTh/eXcSRyC548/au
PGOBZ+xkHDStCwovFkTLuB2f/L4bicotYJLn8JJKUgjcXJGD6cNGZbhy5pQgbOnyruaMzeWnnJyO
b3olzCLN+hFchpMlmeZZ4w2Mv6BfB3DF9V2fGKenSBPUO5qIjKSmlWCiR7VjlfGqX8aAvlOrSfSt
uBfyhTh/8RFNrxciqmQ/OC5A7bEUCtnM5PfWWqK8jF2/7Cv4S+Kk3DfR3tgJ4+c/YWAXB7qR2pmu
bNimr2U6OkeX0pOb+CYSAps9LFXeFiKVNmbEnvbVG81RbeGYy1vFFoKS3lZx65P5t3Yrae7vkBwt
hFJte04/3ov0b04DmUVc8YbApgbS9KGcZaydfqzny7h7mobnmdbenE5bOa4+Kcbj001GKOFkiBpP
1wmgL9PMv3HTqr3vIG02rY8Z1y13swPzfWQz442ebJGRB/XvH8oJCfhU6ZW7xjYlLukgnUPmNdQk
X6F/pxcavrF6bdYfOrUp/5BQhQAfneB9iieBldHg1HlapxHLfXXZlYGid3M0c/aAO8VbQ/M6wyBW
g/aqO+/58WBBjM+xEvuxAgK8tVGz6HBPf1KVWwpkm0jM9y+kjA3+murJxmnDu+RSAzyki9Z4u1S1
6yosIMebAhHHt/I3G5z6V3hUdWVO4AXk8iLes0IfPfAtAUQHx0MlN/qmF2kxh3hfBQhOJ1WovXMq
TgVVoPT8Yim1XSVDatCb0XTLk2yj9e1Tvwso2Y9vjGmqQt83QHiJ7oLVCHvbU6K6HL1JV7DdPWEC
AEnqm9mh60ty80XxLaHyaYJqzDX393PF0n70jrMh7JoN2q69DVcAYcIg2Oj0OiaMSyHgAsFVY7/y
9Wq5pNjjDlxauScJzfl6LsQ4cooxLOEBXqMNfGRg7vbSNW2pvKlmzkVv+UlptVfDsaCmqPYefmdn
J74FRoDIcZDpmBCTZxAmBHAw3TH1f0n0fMFJSkUVCTBD3ymhSBolGDqEnVpI6jSpSIDOLEu+XH3E
WoZT9VIAj6yn/vjuo/tJGMvuJZ+prRD40PwOYQnbjjvKZj+CBFgZ1gtod9EbJyVxx9Aos1N34fe7
+LIhzFglRI0nas7e/RvHICsikhLOuu5BXTbOMyXrPnuxpFG+EcUqct+hyRupT7MAdK150Fv1bKu/
dXj7y3W2agF+ftHQuQuv7cTi4P+B48u0QmzokZuKHBcXBJuyBP99E+hlvKCCWWouVqhrQpAn6Zmc
btIO1BGyZLdSOCPKZHP83mNliScWBJN1Gi8X2X1b5m3u90N/zXlXrQtBKFGp4bkHnOMXUKXLKe3F
RDrKrK62cZMt6pw124gJawOfPK/0BpX7kQRm0+G0KJN2kxzF77t2fnbjoAIVWZt9BM513uATxmIN
a8xMMtpcts4CmeyZvkEvkVq3Z0f1Mw6eJr1SEyo1cMUyV951jAjY9Y98w7JbnFl7DIRk6skBNHpt
wNts9CDuML90iIsNyaQhn2WvZ1msj5ZcIlIjAiQ8l0AIuT/0kDVTnkBtRR9gzVM3dp6Mt64BnQVX
AReTyiy5XSjS5hbp4YS5DkuJBZCkEXi7JIseoNdDeWDOZ+TJ3pZ8ImH3KehG7d9ukAQszccdCXX9
bYwTW50ZjypWCVki7MD00/AvdfxDoHjML6Z7O5aYhx/ddb6I9VamLjp3fEAvKw4ZFQ1ilIpNp+0L
FHU/EwAPpv/MvV2Rdzx0uAJwsiOOdpF1bFaLOt0Z+2vCvhxVwKgMNhW0r/WZFe4QnEQVZZF+jNVh
ER6UOm4bU9V280KqUzmFoxLONzmhiKRobQtd8BWF6gh7MPfc0Hbz4MOWLuEwSUR/iQHLraN5uvYP
/PV2gj4ZA6+qkokdGSFaq80bAbWCwLn70BtmggJ5cGowfSqn9vzp4Z5/ZZeWuD4UBbX5Zzx9D+fw
wOvXDdH6F59tl9WRfW7XUdOe+sz9fFtw2h17nM27KurHC4TKcwyqr/yeSxJD87Kn3zOswWXDKavQ
V+6DUvTn2VPxwtQZOSt1MfBfRMdpmqpvlMxiouGbuHaM3b8xvn8LLiU7SA8Ak+gCljHLM+hAFvks
9GL1d16VKFBK2yUnsDO5NEetidzdy9X39/pqcXbzVteUKTa9ZbQSZSnfk9xqMpmDe/VMDmkI66IW
bn49ixtd2hgYE6blvSh5xdhnS34f+Tkc4ncs5aW4ENlY1FlTM0zUJGpUmuaTZcGMASDzieqqDC9V
gDaG1kK577x0LvyWHWbfU8G/BNGIpR3V4Nf8yrNdrTA+6/Iv9rPIOyZa3TOabzKYcMip7yW8JFLA
3us6rUhmqm1BYmm1TsDthp27j7HbIuUniGK1GCAyW3fI5fkRQ/PGtpcUKodI02bx51jlJBGHjrgs
Sb/DNeCOtjIX6b7BniRECW0NT1U/AuaJALTQ91gb7g608fJn6j8s6emq6+j7FklK9HUV6in2ETgM
NpdU+Lg3uHIeh3rqWVwlxgR8lH/H2Z8GDNM6zoys+clg16hrjSfOkFGubzbswXHVZk8vtnPBaBLu
1DrtLDMuQ4gXzT5kigzCaJUyoFL01+8vfrAZF4QizVYkQpLTRnpzfVmBkMs63mG+HaY00O6gQ8im
MgXUq98Yb2ne9cBFl6XYd8BkoxisizuXohzH9EjuNAWJuOxUKeQ+qgjuP88lJxZCEiDOOmdZlx3z
1WmSZcB8OkEWAKFejI3x6rCOUsSh9UbgfkcT6op+Vx+AHoR+vTU6Sxc03dZNWyOM71Rn/660DBxs
oF4fYv/hiQ1JDMpMDWORScR+h1DXADXOWIXjcFQ5bO4m+SUZ//x+u1kT8eolDztC16ky7UB6u8Xv
iYf/HpsfsSmRXTF6aGnpCCFjD1WCwsPA+ltQlczQdjp4WFfW6zV6D7aEvItc4ifMVvUvx/k5mnBi
5NDEE0d0Gc0GHaOaY75vZBsViRjlUsHRB0xFsLm65zYhkhWdNOJXfrY/azNDXv0YRSeLTd/bVTuO
60Rcw+AirCRg1Yr5lyv0qXZaiTTWqxYydxQEnhKaj1PgedCXcCsDI4Wb0oTXol2tGGOnrM2oprwJ
WOL43njkW7kgFkSwRCJuaEBkNwF+ScxR+lfwP/CozRYenV2BICQC3ClXTEQPg7kZmy3NDF5vxqN2
FMcYnNN8ZCU804IZ8Xy9jrNr/2W4uhaJ9g8WPwSFvsLPrSROoBLayNuxtH0PQB/BJ1NQ9Sdtcw11
2ZdZI/fHexhTEa7uyaLa6reh8Nh6T0jzZInrC4H+g6e1NBo3XNJSr0RzOCrQjikSxXWHeEqnXON9
5nJozqZSXTC63tK/JBzQZGUHtLftaahSbvdI6w28OqS5kczi0p5MtmGzAbm4/iU065UMUyATvXoE
kjmPyIyFT7jQUroIBwqlPq/M48qoFHSlHseylGvMFRG1ynJqzhW8RYADaLr0uGKzJOS43cy97Bo/
IhG8lIYZdCCCn0md6IKwb9sWBlvL/yeVHhaLFsyVbAk8qEuHE08BaQq15H3jJuewe9iiaKG5Dxl1
GFhE/+9UjZStBnW4lup5EihtWkVNMyOqcVqq1uiH5SqA6GNqyWtNAVwmdHMwjJ1d80DoNbCktuvH
nXQRh4ir70mqkw2Emw7LssRhh7PPDp1F83ahzroc6S69gLxH9Egxgy6XYyiwCNoIqHAT78MCNyBL
xxW50TaIXbKKx4cmkSU4Te/zi9FGcSK1olKUnil4/17Vx8IrH5MJw6Ozhhg+FMrnhZoWCh2kMn2i
9CwFJlvm4L5c6Xos+QbkYLLQnQ9weju82QErmw2TW1/kbL/kIQERuHC09qNJbnzGzr2qJ7QBR/qJ
jBcUIeBFCJ2dhGUn00IAr0i1jZTrZ/YpilPTOPUz4d99fWtqpPVo3kIDtr8X5H4McBQ6aAAY4o8B
AJWRfd4b8OArgbADfF9Qaqfp5fv31C6wNoBN3MwqjFBPxvQiHHIMNhmUenWHfnDRoGijq1phInS5
5TuKcGIlETY29gZjW/8Vyt/oEYTN/82uZe3ZD+qT3EDaHkK/o9Tr7m+cXoCOeDypZBiNw2nk8jvb
pndriHAi2dGd8wWvolruJHBaeZiYSZlkt/v2n8sv7Q4ruSu9uWTCnhgEdLWvHhWFUsSEc3Op/2lf
5rPYnDNAFAGj8ZIBt3oR1NL0R2LBDGR4bYseZJYDvDLNdSFCXaXC7WZxkwyMrbVdMVK/fZOH3Ogr
E+rljhtqoS9CzJyRyn5Je9Oqmw/+b+OpLwCDM9FegJm8iFFexKeOVq9OY3+/fh4sL9i24okEZxfx
htT5R0sM0bWykMGk3HfnHuGQrUb8TqMeUyK0q5IH3HWkC4aGK7JYRixWiM6ObgzAdrl7FbSTj0Xv
UVt8ZwkygOlngKaDCQ/GXAT/VnsFHNXUGyTRLnboEQdkKKLNdzxbwoMMqPzc1T2JjWBtrHNlR5eR
UHSX8zr4zd0xRPoOL4wQ2O97jXFQLLZripuIlT/glPx7GG+Fh3kqgSUu0H5yGdy+5wmNzQgDS/o8
Eco3mQXiwV0scxG+cHZMaxZLGLPr+gFs6+ASm+deLFHsAJFlsbhVQoUmExYA0L05TIjtBYvpvwxN
V4+mR33ZyFe0IwQespxBUGsRDY6lr9pDNpz+IW2nv8EfcyhrrSFft+sCPhZwxPPmxJNTsHtnyyAn
UpnMlKbzG5yd8XKtWtPME6S6Lewl6wLUqMOlVNqZl/oZdP3yIK6UKTz01rpluSvSm4+SsY/4SOG3
jkp0btA4dq6sZU+ipT9xs3miUp3Hx/zwZwROGta8eWpcL2BPlC8v9zHjq073qxFEDfEKuvy2OXLg
qJ/fX28U9RjzGQAnYD6SPL0I+DiUyoRbv97NdTFb2ExHXjYSWhMH6VVYLo986mI2oXXTppNN1Bl2
L0JhS6GK8BlAZZv+TRj938bFkJ3gGZb02LFkyRLDlN2+22W5BioB06sFjZnAgPL8i6n6LamSUMNF
H9tDryk9o7aFqqhsC7j2hAuOfGVUkELEsBp9jBYCByFIsJADcTH/yhD6VSQuPLO1bZff+moaJZMN
MY8EFz7VJRt00vlLitjTom3FIfy9i6LLzOBOqVp49jTuTV/b6LYovaCSt4B6xtIrVTO81YWym3yn
tyvqf9POxvI7MMfiwoqg6fn7uyjEdFiYeIbxdDzEsOPb5VqVlG5C3aHiFhG876/if6IsHhui6O8X
NPopJZPjIM0HO6BiJffuPWEOfI0Wic3hqIFbkndtLLMClxQHxw3WaZNawLg0FRtPnSRmDinXR66Y
vxGwjYj4d7iihfoTmeVL7rA6bk4qwMPKBsDVn1u3P36VqQNHV8JH/6uM5cmzvVioHUbBGJUYtbde
AYuad/5q3C4Jw78SY3RA/77uM12nPnhvZC5hGGYbhfA2JiAjWj/lguCjp2I8tDuOqJgPwFFRo3uM
l9hSiEiFBsKZ5L1+8tJoVkC+RC1QGt9pqtg8F6IeG97HqxtzZqfSgHJvkl2CW2ggc8B26sS0qwNF
5hiBHFe8yjbN+WMICfwLbh0KFcf/9vQ9HwGq+2oGmDPX4JY+OEC8rRgi8uRJQ/wCiW0aYZv3ze12
7p5sgWZ5jS+qQAMhp6SaFShEQt0wSvNJ7s4sSKd473tVkALNZv98GM87gTvDUFlqTkPNXjjeqbTx
k2heg2sZTSETfAqNtlAGoQJjXWW8J2bkNa4f4MWR/GDPPkiToTxA+LJVnCrAdW4CLIl83NNaTcNU
ad/4LoIi1as6dMex3NSUuQOV8EdoZapq8sPRVf78IJ4nGAuS5JLpc+LWufKZ1tYneg+aflX3SJRC
oxPsm0QDYdWesTQ0eA9M37YzR85DH2K/w/7S/iTNbOzKxohBkBvtb7BhPFdWbp94GGY0NCvIx5MX
w9jBmVVFJmKXNfGOPH0x8M8R8s6P+BhugT5FTR4/1uj0d9eknaNOjz99wF4fqOA29/y6CNlPRdMb
YOKCOlh9RC+7dxJ8DsKei+9xww+V5acwIy/KTcYEemJLwbVCh81eAhcZXIa0PS60ridErhU9006m
x4daD5Bb1N1D0xjl+OoxGO5IJinbfJlo88Hr88orgDASu+EESdwHJ6SRZLg9h8zDTrD0F7CPB1NY
DMJDCAselFXa828Oh9NwuJVCe2GH6i1FX+qoN/YbRlEUpYfUatE9oO0q0gq4JVUB9dd/XD7OnEO6
hFTidf5IiV7cV9oKoP0OobHXVnWggDVwISSk3oOwsa27HT4elDIm6Hw5LHsLmCaewNFz5Iy817BK
1WtKA5URTuU7qbZ8FegCybGT0tuFU73OV93ebCWzdrYSWSPXt5hr+HiL/OJ99fAOge0VHdDZ1QlI
vPeD+ucpgFnfcVxAGQaKqaC7R8UpsZU9cTyjTRy7HkK3NLcK8179Bx2nsUXX3PVyznOq6eEHzGA5
epUtme79AJGKBi3R68pZjfMxxxsL67bt4phaCf8mGcBmOMrVDrWYEaCnBwO4KOqCqkXSBmTes21K
hKP7ttSKtfQVqn52zSGbuHTolWaB2lFE3W9axhfJqIBTI/A5tTJxnpsvbIZa8FnaCr4mpXluRS76
skvldO/DHC26aGVsgjASItPBdYHlCfDnxrDCwI1YJaZLS8VprvQD6cyLBM5NRaxoHm/1uhVyepk2
eHmeipPA2VnIo8az0nPIrVYaVr4ef+SsfPYiWaEyMcCTm5RPOshuHadUfm2m8v+iqkcwmxX8KJBD
F7+28TEcAAA50KJ44wBtVw7Wz62yL8WwRWZR+wd0onMZCY9po7AnCJ9gD1cT0zuJLoHkYTCWi32R
dGJdky4KzufWo/2tMAIi148wLaGugLHYWwCIvtin3LHMfwx1i8TcBzmDzyv1GW0QTs/GpbVwfMzA
bmoHpHwYD8twMMhnhYwmsaBXUhgVV/kcwLLS9W4HA9cAe+lGGezISDAyKBGYZheeMNOClo3vFG02
Ccjn246w+4SdO5+eghTvTf4hUq6JEmQQQJ1I0yGcbMGDIdNi6nowUzDFwP5U8eDiG3sysuREaadu
TfLPN0bjhTc71P7HIIKxaWAJ6rRQ1lCXHU94HuSvu7dnJMeJRLaYX/HUhL4iEH+v1xsiVOttdTfo
aZBcr3hrKmdV65SfaTxqHCf62bOzfglRN1EA4xdhzvO4pnhyPrU+WBxZkzpUVSVN0eorY/ZL51l0
i6OXiYhzpaR5FYNAXNRXMEdZq7ja/suXyRRJVRYfHOYri8dWadHLkjLHH8CB0tLFVgT5tDTGEcbu
kbCx6fnhzJnVeWpDboLwCOr2dfOnckuZl+ebsh15GX4blyI6X51Wh5D4Bj0RjDbuZvsJ3thW7iFI
vO3o+jQ1Nab3B3dpsiMmxLj6MMhsI1X64VsGA2ZZ8zDgsi/+m5GgtvMDLrEtJVrx4Y9RVbd0b8Ie
zWc0jt92XD4iKWtpivfC1YSRZzon/nN6fJA5sxHsJmBfqA1+KaZQw7WcUlRS6P1hnB6Qp0WnKijO
H9XwR6AO1WksCeKk265Z/BWiCnHiXGPQTe2f2Qt2NY8rQ3/aCeNsuZT9dpho2np7mG2QJYbgKmIR
aioCjH0qaOU5P0FllT/Fw0Ry7pRNfNzWEbuumxJIjW7MOEGz257sOPxI5RIHT1bixe41BVvKjRK1
YM5HG6U4ygJSozlXgiihB+KT3WsQXcCrfH20hNTGkqcWvZgz3Boyzm73lG7Pg28YhSyAhkekKYJK
yeW6fIPhvOBBO/KlbpiDx0P0QA5QYxUVHwogLAUgg9GgvvjbmY4t7+WGMJOpVl0p6mhrFx7IQ19L
uTVXgxxVTpkrSjJMhgXREeOvOk3WiETY1aSEwl5es3HaohEpnm1XBePV0lZ3DLoXn67v1pdueWpl
OjjbfhBJzB391IwQHFXOv1bNcVxfLTM78QcT1RQ9pvpfs41eLR4/2Qu+BcKJHyiFbaYOi9OxbuXl
52aZ6awjVoazX461XfF/MOQpiiXGsPcSQ93K3U3K87oa18H9YkCZTzjM0w6WN5D2qf8PJK++FxWs
SQsC2gYucQQgXKOrB6uYRwZsnc7ICRPj6I9R7+6zEFYKzrdFhV3/zddcOpl6lpw0QFrIJMycZEz7
i7xacpKBywPwz2ATA1VMvVWp2LgkLt2adGLFQ2nTALXFOzA1DNPXrroJ8eA29+PLuXWz9PowzXhS
WaKtgSQKhsXI+p6JBMSN/UIYJhQjKsjlN9tG5A/pCCbPhJH+y9q9A/vgE2TyJrSYEO/iYo9qBc7P
I/FgSuWuO5s2cdRL2qER4WjaoLP9V78c2GgJhd26tEqg02rwFfcWKzr47oLpLtv/X7MtskfeB8t7
yR9btKBMMoTku/qwv2I2ceziVmtpLnnUXlyBVPQdGsK3Y4mjhJ6XPs/JD7SZ57Hsd1P5wb6EjcNd
aT1bjPIj+0ELiAMeTq8IAyrX80SR8UI+v8RUxc8h4itrIWLYD6h04HEy4HzF6d6we97mSil/Mvl3
sZGMiQGs82D6htNurQtggExsECzcqO0jC3Eb5eTnhFGB3u7ofRISeDjRovcj7N5oea4ZWPMOJ/1f
CLgadH62oznpL6Vr6rJ64+W5moBdSNnnioPLEEtkbsJ3wIHtp3REOanFkuXJkOLgY6QWlTVrbAl3
l4/rEhErgrP/WWtpFLsND+TFkk4fbyWY6nPpl7ZFcrU+7eWejcbB+rQzJUH37NZPdAtlU+X5irOw
X1auFcglyf5jw94pM6FOgfBiBqyasYhf4EMfJvsvi31AljV6hnk2yNVplpE1GtVuGa1PHJYT1Eth
oVMlwE5c1jmtIjvbq9wPF0XMBIIELISLSE5kpkrCeytRKA3LxIgqhncPWgxMy11o90ilYxV0Fmm0
CtIWlIuiq7cAbEXgfJ/98sqrIw9vktFjZX1IcO41Lr4ZpuW2WA44RnIvRawG3AA7Dpvn/9Gfjz2u
4G46uG0GanVLD48w/PD9QzgluVtpR6zLYq7Ry8SARDHAlJGWyrywkRrgrJKs7NUn7vl+b5r+aw/e
uRSBmT2GS+gMqH5OpgPdx0rADBH5AoidqhqfX8R1e6QsG4f/gmLSPHkRJGXV7cq9NSV22GREPhQQ
jqXYlcDNAICFZF6a6AS1FSWsR7j8I+463NbithdjaXASzJtCZzKsyft4HG1P7o2EKXgTiNDki4m4
T3N0hSUF5SI76ydZtMB0R1T6z/RAf15kI3cNx22ZAPP9CUqzOqaCSr/MGRil/L4wfPyjxo2XPw55
tTBtI5Ow3R9NYScyjwY+KH9ddz7SIFQYRYYkWsYPyBD3pJNDnnluNXCi8g4QngPaCTK/ijNskh8j
dxnbZ7EWxSfritvrBVdwB7gvIOa7ytRZAU5kt06CELkaX8pMe13YqJ/7dqTj9/PB7nTGwR8Axlui
WPAZp2VxUbQIloE8hFGBULJ59xT2xx9N2v3ImwwN61DeOJp50JfzSzLyppJCILTqddOs/CQPtJ1s
suev1f853NuL9IiKJqQlb79ut0DfCTx9ZDsVZnM1kQ4gpKp2uxaKSSl1Ol66xRTpeBbLBa53QRHC
QGmMqYKL/ns6/L1lfebpeCU6VhtuHXYmvLPmNiBu0cyk3MIEcOWd4cHxFucWSit3GMkUCiUhAtWR
Z42J3ZnGNHl7o7CFsaAHyZJZNr/YeKJI6t561YSZutxv1jmL8HVICthKU4wbRVMh0TiMENkkHeUt
k14ynffADYOwQ/UEYlC5c6p2XJYFt2xYm+wfNKzPDjeJWqzneKvLLvPZig+anh3K75xmfaeO7rFW
QCEosIsV+i/1SpRTYch7sNXgtHISuoaAAqQQme/tKakrJrI/eyu2cnYhFY9VYun3S+KG6r9wfWOJ
/j2LfdgkRERSCyCWVyslpgsfE2EbKw0yzGBy/qmtIBuC0GHvuX/8OpWolGBuf5gOZ3dniYDqKxyD
6SfSq55l8DR/v62U2ZbwiIr4MGPBS1/EYdHzIG973KXhC5nnX8PgjUCPSVMiJPt2P3icGY9gs7tP
A3a0BzXGr17CiVnfcvRgNbB+cVfRhy1eVOUtQWu1TGgJCjt2rfpQgpmj4P9996r1xm3oraBGD1Nj
dcdPN3+RLZs6tVk2HS0s3eqmOzCN7s/A16Gk3Y/w6DsGOpVzuzteyyBwrVgw1+gx2Z/0A2o4n1PL
cZrOuVt8ptxrdH288y5jtiuhxgasw7QjcoafdLcEROx1v6du+nXFF/ngw9SK3+Z3UjD5UH2rDrTf
tEMVojnbuVwMvRmwywu+qdzWt5mtfiKQGH+aTNh3OdIp0thmaYh7QGtt8/u3/Qljh6NQPp07rHlk
KdpqFGJ/z1FfKLfWh9+7Q2E2h619GKR6DmAVWsbqSn3bNRAYDzgVQunV92mMwtRyqppLcGhPWeLf
gM8wG9TMAd/IE8JxD4c6dQtUIqYjNgClercVp1Q9yylbppwcddkwnOJ9A36YwLUyajEgM+Lo8mBS
asGK30B+OJ2xpeoFjPJ7JdbcjfkbDVVtrM2OAhzdD32nynZJEEZdqty3oy5+bGh08oICEra0EW5z
P1O/IhTN/p3PTfftalitqEEekSAR5rYCm82RZsk932sn7cVCj+KqxWC2Xupyr90hov1zBmMJI5zO
xVjLczvmnvQbq4NM7FzgE9EUEDZyLaNazXpxfes+bBW/sgaIdszHkP6O5wKxLV4cJqIf3T4UWE7k
7RoMF56c7BrxjS/keXlEa9AJtpjFzceLJa7wNp+dVoj0fPrqt8DjV5LXNHY2tzBsBGNTXS9eIM8E
nHuHZ9Mu46YSVYtapWvDj738kq5aKiwUaibI5UCRVJsWMk4+B/QKkDxWTnysBf97fH6PUYzYD19R
qGehXvR1WJSY5fnfyCe9s3g3/imm6bPkLV3RRNqPZl+X/5h6IP8WCCCmRCcgvdF1JkmcFtu/s7P0
Q+tSODfhsP4HuXJDgbhySQczt+R98/5sE8j9B0mEZq8Qiqf2ntiSocvEsZBF+fgqXY8DBLUBwPOw
oSz8rONoHuNh5D5STG9Ax5EEhoiNip3WE/lSKsMgv7As+WeJ/XeVyQHaR/q29jXR5tDpCI1pHniq
jCvtLSfzl0dFGaG2tnyq7yhnLxtnbECbqF5Kq+YlAariokFK/8QVhKVUpwCgkD7gPYeIbfmrrm6u
LIcx2LjiBmqo01+//rb/lnlthvUkjc89CAnbM3G000mfhhvIFh2+dTezCfRvWSEykSMH0zUwxIqg
hm9RRlb23P/ieI+c1cBZSVUxNaoWQh6XTctjQ9H8fm+yVfdqLJcYKIFz9tkBiT4V8VcCBGzQVYEu
qWIXBWAdjJw9zko2BkO6q2eBfpA5KUd2DMpUU56kEbWgrksvzvyKFqDueLt7sNTEgxAvtnYCDF/m
TqWwDwKxytbnDDMnZHg35M3VqNEXKe33PRcryvzqUnzAj7CtEHX+hYVH9msvTdPG7Ws3HFqYgMxL
eJT1U+WXIrlHiDA4jVEOmKxf9laBcRNdJ50LQgHwKzhhVFwhV96Zdwbw8e81LZ6uS8lOiyTiFNrB
NrcyMUMY86gahdTTUC2YUpDmT+DSgkH8sTrlaLVWcmpmG1YryUKJGVXfRl32OkMV4DZWWW5CTFsS
8uhMv0MsJ7F8ZmQooIiKH6ck8q6Rr2mQMXwk6EUKj3ingyyPQJn0PeU33PL3BMScERuwK+85eNlN
mIekhrXZpgnBMi3F/ugNMXZ5isSKZp6IagyiNwIYcRc2ZdAn0vVIDcu7OG7jUz0ZO64oQUIucHgg
WML780lqhuXFkEbKqyBdKEvePp2ae1cnexZgKODIOJ7aM5BjvOijMJNcA0DPcGhnIwcBG/MEBFcl
/a/a5VeRJXoyx7oPHFYmOkG8ta/OhjIvC5s1OWRGMNlxckL6yfFr19PSN+hrLkBVdCjJw24obuCS
aCikfNQt+C/egWKv2IjrFHd1etocVycBQM8dvQWHSHX0YVyiHa85AXtQCVkM6bd5QqL0pT8AThDh
NmK7OLssMWFxZ7UQRGGfIHl5tp8V5fBssw4J8Kg6WQroi9PWib2p5ix43qHFFfSjAcqJZsgq1OeC
Hh4+r6jX2cmUgZ2MmIyA5Eyl14PXYLW73aExVrm8Dkd1vUip2iTFYvx8foZoTOGO87K5tsYf99DR
RXl5GB/Ve9cF5WHudsqfFrB/XIawxLaxicB/XRJr2U/bZHyIBkMlwMyZLWcqodVTldFVWSPrKtRL
y7ZS+AIK0X8LxXJuU7RyMXGidRJODhFzvSbfngC+8Eyae/0hoUgenu7JMT4qmRhNIlff7J8BA2ub
UNAd0tiXVNjwTaas+ww4Y/4CzdAeKVHsQLHl2IrLsOEHlVaR0/Ktj4LLwJ6vfCyLceiKCOynm2S/
cMBZXy4DLbm2BQPIs9Z+QYJTUYD5rXeRd6dJDjUZhAsuLNzCkwXaD+KaRNWRQAT8Lewc7ZFD5P/V
mq8621RSXGeS+3SE2n4gQ0+DYduDzYItvTE4zi27Nk6s/ErUXLPzoKQ87mFCCzsVokqVQGg5GMtR
GnyRzL5ZSE905lPxtJn1zm09MNWuwm6GcNoxS3idSM8gIGpcT5Sw/0FMQNJ0jaT8ByKHtLqLtgoh
x2SQCDXumyIkYI88HFvxWKIMDTtPWbjyo6bBtrXWtBdssGQ7kuXNqP1ufN7DTIZaND35ZOfnqo3+
KurBgUiomzwjaEiFy7R48mlx+X12uTndQ7ZQLVRZVjutU4iY9lMjwpm1k4TrQgxBDbXL2eicJKT2
c6NSz+KXK2uMSXCpdVVobx112nGIMykrPBDvSLt76WwaEN/Wz0sOg07QaSGPMaeQIS6dqIEGUNMZ
xbAZjKfNI7pgawhNTa6Lun18ymj4XB+iS4rImVLWtGfwJRkqvC0qaNW3opzECXhb7PVSwNbiXpJ/
wHABun4+tE20bs8QqlPOb9UEEY6hO+61OFIeonnRpBpR1TynF1bM06e4c6uy5VVJU9LhxsY7hAV7
zQ/PltKkfzGy/XurH+OWnl75MUxDl4NQeohkQ2eXYT9rJ+4cE+FYX1xBfHtnfkruQDnCIZ8eCHkJ
gp5E+vxZP7l2XMa+AxKXzG+lAs3XapZQGNyhc0gtHrVpnno46dN7rfJET5Y53Z4pqB1fAmAliZGD
CYYdTlVfRlKmpMeQIPnfkE3gwEPLq5NsMa8ETG8EFKIm79CvWyQxdyUwYywUs7RN/M1VKO4au2WG
9/jLSDHEVOa6a7rbLxgR0gqbBML9Hx+DYr1648hCZIL5wZwbQrMyNuwkPAypTfafUH/pQ8lz8OBh
G6tsun3+9MNmAzHRlIzcAmpkXMq4GyOyE6v/ybsf9OboYC8IjrL/5sOKuy/yRzAlVzUiuE+4jZwE
9rm23gTZX/quYUH4Pih+VltQQpZDRVc6qsaUhVmVZSATkfAJd51dCZT0oLuTxylaa2CyQZCVDQ4/
DRx3r5PgwODEqptLmnNOcm+l5vRKu1FcOeaGcrvh8v+FHRGL6OH6XH0HegDhtBUmYCSF+0WyYd0x
UZ5sepykWYweUBY+nKq7DOYeaLoUIXIgaHtgC6+5+gJB1vcpiNY0eEkIlrWjg4vT5Xe3SxjiixI6
Qs3RKaRZMcusfam/ZDvsY96fLJECCFhCD/Vg94H2Xk/4A6Mm0KVr/kPyIwN4U8b89yuI9rIrnYEq
DJoZTTHS76WoTKIqGbYOmj8894HVpJAJ/j3BIryrfTCar0NTdCjOMO8GSqO5DBEIQUOTJti33Dq3
xKZBRRy3miTgRC/TK6C2dxo5f27SgkmO1V9uuQSHsrXLASJQW3dcAmq24IuZF3FstnRKfdSAnKVC
uFN1sZZyp/VNdGXT0wZI7Q/0wDMR1Emd3PPFdEhvgfuo0DyBHc0nPhGH5PVnnB9k3vs4/Zc1eGTZ
XVqGlBQ2lIPUNe9l9lfMrT7rQ3U2cH5vPE0tKmedhXdBTRLECdxSXecYtZbh1EYW3G4Dde9j7Ed+
asOmuEP0Ugc0OQX+lC0LWRUbj3eyoiDo4JbLnon4tI06lCcQHj3eODw5YIMEnw7SY/NYaiA8iWVL
zEeZgY7zqTmBFzKVRFhHnp0ssualqaA2M5oNyDrugu5wNvhon4T2ZXAmE02BZHqqkqql36T0Ayc+
d/EknSB7xYphIV5iEKPPVUakMiSval70BKNDl5RLyOLtWjuUhU1Bk5cmsncj7m0OY26nh55w1PQ6
oFkZCArmmXV1z2n+bu91s1AzxunbtKnkcGlv7hlJJWQsrIFyc0puoJF/KViwAEK9erq3TYIjTXgx
i1dAwjgJpy2Do6435tLqN4NONTPPL1x4REIy24Gaac6y4H0FE+HoDFNQm7fGf23S7wLVeDXjtaKR
RK3GBVmR2buxY90t2SIuW3VEohKCRqB6OLHjbc0MoqKPByiX7tT8qdP3a/s6VEe+R8csDAcbNB5w
/GdRojOV8Zr3XmV0DPvFBM1LQRH4pjqXpo9U8HXZdFTeKcHU5Rd7Yh3oWRcchi44szpowKC2Qp8p
7r/FU7ibRv13xGQzH54eUM6oAi59Ej9J3CB4fXIQFk3cvMqMd0S0DgeTN+WJNshYeAfCcddTwkvI
CvtATR/Tt3X//frI0I/7B6SFz4ZQkpwQsVA02IwHAel8r/mqmCxkO1O9hctxQdvgjhjJYpn862Sn
n10oqnsX3ARgGlDW8V46t8p0Bj3xy8n3lmSlXntlQBzBkYRjXAR007GEC1t+K5bIkmoFJcy/2L6d
ivH+skjzFbeIuUs0Kmy9PvL+kPQ74jy7JQuWtfklhQsjDtzKZYshgSmMXC9vvS1flGUWBwlKzHFM
AAo7Xbm6QoSa9JwVEKiHFeHJozH5Rj8VdHYjOrpi2G7LlYeC8aDG1S1HeyDYQVBmIamY2Dn/N3JK
W/atovj2oBDo0c2LthiDZlzFTt2SKl2WMztSDNEd6+lAMX2eowNYS/S64pLycxFR7yZ//TWcS8Ou
I9i8dJB68PFda/pSD39C18Zcpkp5AalM9sIIo4zU3FQhQPFpJc4wgGo6CLlbKDzO6B69vdp0rvmW
SPyjlaqNJbt/YL8M009837pL3sWbM3tHst/q5SeSPTYW3NVrtYZi1BJBqCTZJxODtJP3uVmhK7gI
GaWUKspRC+N+UdhXhESnOaGcgqDZn4Da3i1lFO2fPi0omojX695FHijpcaVVAO0KqzNQvhBlQhnn
zmWjCODA8J9JNgSyQ+a6H7/XlrNrk6j9bBKc4I45m0qakRVA1hUP4qancbm8uZWc7bCA2xZeml1N
sNRbR71qw41Fdsat0w9mZaFKEDCtjqVWCtx2oMCXCFwElxuAM/kWmjGzJoOL2FPhccvfY5kcghJd
drNNtI/ykOHjcMXq7CUYYXUdqpvVpLJxHX/cmj3eSGWh8SrksDtLS4Mu+T7vjjnIJPLgucrXHQ++
V+ssxWw6M9kQhcyIA5muwtH/+0ml/IQWixU39H2SVFHX4hjsCRTdYhFua/Wu0ktXthTIQ7tlS42p
P2NmSxb6PNhHv9y8BfpchY2jxi0om3YaN8ASPht1eWPnP+eSBN2Jd64ZiGqdFwvnnNGJzI1orKxH
dSDkk2IfqFet/9cpUozvi/o9N3kB9YVMu12JwWaLFGmVyDWdXs1x7y77Kp7T/kHn/K6rWh/A2j2C
0tROjds97x0K+5txlt02ky131XB+fd7Pg0ulbxBFF5WLgoY+hON9yIQFKoW2+XdKsShmzUGD/R+I
2YBvwZfZ/EtM3QALFJqI6UEy4+fCfm1pnX/ajXjUKQxF0/0RQ6OBK5R3mMV63D0F8fjMbbATFD6E
02Dg6KUaNvLzFMuJwEuu8IW0/M54LGFvdEuVy8MyHfALb7obruXFOXdf2dloqFpnEjoDqJWiRXHZ
7LALbmDxu37hK4LsA0NQIod7Qvsa2bIqeclgj8OWwjbxUfwHy7I7puxUWQ5J5R2ELF7yUKZHAFcf
vt3ZLnG5NxPvN1hbjDt9bzpq+NRicVUKKT7xAs0Bq6UQnEUV1fM17budYrsPLIzgu7dtKG/9rImS
fBsLPY15PUqFx3sF95m8WsHzJECO+ZRL3hcfr9xfwSostlcAqejS0qfgQoEDo/QcMsq7XXIJ3ZzB
r3v4lCf4cLsWpuCciNUBlZKvp8zB1ptRTqi7maGlcrkFC9lDJACQODwnGnD4EoizvwV2nDmjXXVq
ATwRuHN3OeD90qPdZ2gszy791YqCUOUTFJWBKJ39mu6t9gvVeixhPDZVvlXNs3rRHmdb1i556rfP
dM8V4YtFBlbUwJB6oMwkBg2QFQUqqqBPkr0GW2B/enrr1f2xzotBr5MNE36RQ+PLKlK5RCQDGMx3
aWags41pvrL8/OtAT7mx8ajVu5kvyQ+O4OMdRv9EScEJhu0gL1xEWip8di5tmlEOkCfKRY/nAptJ
1bivG6MJ9kAWTrmqhrqt5qojkLfXqWZVdg8mnzUvXGBisf0t8Ap6OSCSInuxS61N4ym0gQwXuaji
YB17kMMuZLo96WY8meCYSzek2YDenBSDtKh8opJkyNOwSs4onSaHJB60c/hBZlMoLY+NrLEb6UmA
vVJhrKFY9z0fXYmVL8/aEZqNFTEtwmorLg5mE/Cd10mGNsS0yGp9E3HKTFEWSmad9hNxGf7oDqRN
uvRWatJr5ZCClkBb3Stj0DA3hYciYKB6s2p1xrkFvkf2394WboUrBro08dy6XNMm8NWJYxp+QCCc
y34JzdlTxJqOePBkopnwEdbCe+IUigzD4qnfN4+C4UScO0Zl3fXTF0muVhIwZ6GSZaN5myYtamSg
FNwRKqwn3FC9bl9uogJJzlBB3Kc91JrunEkN7VKhCPNNSO44FfDrzPSUShlxQwgfRknT0WSSjjDM
6pHjsTKNA/jcq5QU7YjFsF+5EoXWCrrp1/wnVUf7t/c4QKjl4x79tiOgV9XnX2A3kKcMmRJReQk5
BOWXNjRML2niZbHzcAkHWdJ3mbZaZt0rY1OYCet//2kkn9ZMhWLCajfPyiHxwVFMjeuOExUAGtup
eRk2uLV3Ru7lSC2M2cIqaLInIZsdx4v2C/4eTqKo5I8vH9xrm+vCn99946G7pu6SB9nYiTILr9Az
51EkD311c9GEs7o8k6LHySbrygWLyf2CMj5D25BLNgU/A/fYVU1Jz2I3f1otBFHhq1ZpTT4vx6jF
+pNO+qoNW0h13CbeQOfxR+kZpssYUG/2J+dG71NzL3T4LFF/HVFm7/Ip2iJhtQ4NMjhn7O67Q6T8
zkm3DJuRxAdJd2GZ/oUAiHHfwm4SM8ugfOBdfZD1TbrNGfkJ+zrra6/FnfYWvBZ+tZRSa+3EhbCG
jqp+k+qNMpOuoBiWp+bWnzk2/FTXikznnnRdHLZLhFSf1v9DmpyoQFL8P/4OlFBoEuYs5XSO+Gsb
kTbGC19CuWF/5t/130ICtwtec9uSQt4GSX2P8krdFjNuO4BAkUhlwEuIsBQk3hubYa/h4E3EYqvD
X+aZ7hSToLEORFdgCMm7aUSRtkuBNwzYDzAYWxgiT1yngSOVqqjgCL/9SAuJpRsgvesNQgYiKIkd
Jp/gLAVBhJPeNK5oyCWUjoJ9g9iETvIptT3NdEOJXymzDxkq0WkIh+pW29I3k1ut8j0YXHTKxj6z
rQ3fXVTBgfzVnPT7lPmGP706fldHyTUadlIpiKMpw34G8FBcCTF4IhuScz+ryQ5bu/8xzCQRO9J8
VVZzNKZUp+069nHvmPzk4qeJ0b/YoxjQ/q1NukLqERgOybXV6WFSP4B0tACE/vEYbytqTuqgHe4s
j+jDVon783ySyjIKJtYTZ62QNp5N2UhWsbq4m4D7+9pc7+kJZMzljodWhpnvu1C4B3fM+Y+Qwu82
JhkKhr2cjEs7D5Weop23MIXV82hEwuHy+dtCkcQJlnGjSykourkU61h+FEyWIq73Jw3aY42P475n
eOOhrSnWG95uRnOUKg/RfqmS07SnAhOkTF7ZKQCh75pLbEwqXGgZoZOCquqsn2+5xAA6LalRN6Pl
JMBxE43y1HuBLtcnIvexe9RqGKNkBlvv6L8ytK+kRfK1d4XpDpaNwDDBeMpeaxy6RkAD2XMvoRvW
sDrMNcJ+bKtOGbo3FXOmZYHJY00IVLI1zWvuhpx28ETKJqQd98kXMpX8YPqCHsdDIYwnvCLiFkFA
jb4zLFuc5nv9gdlqXrA/ckXSzebbLfT+AIXXFx/Me9jLhnLJr1fzjiVrrNVlCJuEX7ryuV4ujMQG
5piFpiYwmGuCsdZu6UE+zqnFOwoc6Bxz5uqduWWEe7VuO2aapJA2goxLAiZvtk4+xg/iAjxkyDR0
ErcMS4bfbzwdZZjuPNqIGtAh4VZVXKSYDM9BPgllJK80PSLW6cCxbzNCnhL8YbtDdCNYOV6ltyXP
4jtBJvsRt6DBqRzPBUreMkCns078XuQimzBPU9ShHOFw46VQJlUPv9lmWXxyryjJWqw+QM5fkybJ
GTOSKQy8MrDKWdcCBl972nLW1SmoDwnw746989V0EoFCzftsEWgTm6sfSd7Thdji6Auj/+82Msuk
lW4xbASmOMNQm8Is/MborDT27TBffYakoQYIGTE2lZfptCUBiNtZxodG50nQi/W5A6D8q+L+ttq9
yixrI6/Z2VM56YxYkW75IEuOawpdHCIMaN5kOuvOdLhBzohyykhX1aK2kIhBv7piw35n9+RXSVTl
TIkkwZRU7W4p+r8NbhSPKJDv75upVxOlBLnPYmhBdOlfgysp7+QXZ9wd+5gZRWysi1627zDTJAL/
zOusURqE8RsOSuE/N+cJxGO4+zUz+LINuzgWjLFi5KUW/HLPdBNw1khCarzIcScFaF37kvrJxlIh
5NTj6rEb00XaAeQ7qtYT3xy8ktaVogDRYTPkxElahu+xhq+QZ8/m9dP9U6owqJ9/O6ve8YacVez9
E6Gkswgir3MIYmQU3WpEa7vLd9ztJnpNI/eiGZTi50DEeR72FOc0+wLALuA4X2qc80kEozzJYv2+
AwN/4QzqrA8Vc4vQ1XooVosfzKLSbHnJ6V0JCUiHWBJjpNuIfIyj4jfq5z7AVNV3Z1Wc8h/zdugR
H+dpQK1c7clBy1KcjuPrsrRwcDFnhAPq4Pd2ScDvsxtfVfMTwUm4y65ZvFnVviPk99VLMkpAYROP
O6bPcYZ+EWssBbRd55Qf+oRqs+5yOAeulIVLX622Al1haptwbV2gLh/K8U/2Tcn1iv6dhWOeuGpi
sRmFEaQpKI6PsFjgyP3jRjT9s1k/fMlt4kcc+lkOhWarU51iFbuwM3av6r2QgEO3sro0HAKEx6sB
Jd3VaXCCNaWDl41jMUlyDFFsb6sVycOBsQrHUvqX5Ktlike/DhtgItuUHHmKQr4lLqoiSVtkHdEJ
ucPnrxy2Jbz61231U1ZL5J/LxWmQUxqVZGgKmV0hCcrSQHfUjWpPlGAs2DGAH2nb4uy6BO68jC3S
ufxUXKgPMrEIU1NRb775+gBO/LoBn4yAc3r2FQbSSIv1D0mcR6aRNPV+IsPxbdBoFr3Qj4FOugEW
ZlNOALVo74UHftU7K+PA9gTsWMyiTnYsFT08xUhBgznQSt8mpk3EO0O71vg8HrfKTDjA7oOp1BK1
6UHcPLLjUPRCq20RMjm43yKgZXApV35a3myi1+S7R/AgI6cs3R2doUL+rcH548zAb7IuPF57v5BT
U6AFD5VT8AUXmSwojtPNFNIDDCF9uUFraxGybcYIr+rTNsYtAxLbqi9gD/ZhWK9wl3oT2G8S6TMb
HDP4OEypC32IAQSADbBms77ABAguaa4xVMtDOUygm48mOb5fP87b1lT4pg+j45nkjg4TUWVrOHGy
ONb8QKOdp08Ivm8zIpD1bZSBG5bDQTNAMziKKQ/j6Bw4/oCXuLYuGemi6leIhF+DRsS8qgvFQVNE
nlAv4v2n472sjXNOak1snKtf2bL3wt79nOoTHmy60Q5XwnUapi7rRljVeymhAhQH5Mtal0WFYqxp
/D8mjADRjLO8Iep36/aFjH1Dv2+JR2UiVG0ry4DAvQFHy+M0i/KK7HpSBRIxYWxZe7LwOO0FvzjB
UnYgQ4w+AQNgnHZfUEjpPTNSE06UiKkzrI64dAPSy33NxEe5H0+d+h/XqkigJHliDphv2l/GmISy
EZH90RPgUZ2LbEBvpNBXMQzoA7NjFyHTrnyfuf7oekUGdygzgzGW21aMNAqEUPoh6BSohOibYnmJ
egax1F6QStjDUsGaaqlB9WXrnofWJeBIuAP3dPPECM0jT/pwfBH5jzoYVEnE+wKXT3r+0x/gTl0Y
StoAMj9eeb31z8yfozEmlylC0rxNwrm5+cXjKpFxi8nnimJa43GaR29FIz4mgLwE4mNSOYYfg6oM
Y02R6+5w9abHtSQ25XX22IRToBji4C0kX3Lh/96fCfSrHcs/VE1XMg6glj4RfpmCEnv7VPVBTiw2
46SEj0fnn1Lm8jDSdwb4jRlwsTSX1WXguLK+DSu7XsqdHXd/aGkOFIRyqTkSaJ8IK9FG0qss7J1B
ymPkv9zURvwzIPUY2Ri45UFI98emnqIkU2ZLTj+E2QOmBvCZc4Xs8NgDq4rG+TbcWmNZar2oqwiP
AEc5lXM48Iqp5JHcfkofi93JxCklIRRSwxXDtEBxe8ZlE+Xf9SV7kKS2jlUpozlpCnFliwe7alrK
yfDHq76gPJHJ9dRF2iSVvmurrUwu1bumXe1ky5vQW9AE2wshz70F+J7lsxnepsLjKDFrE8hPSOFX
4ftusvWy26IxYTapj1EmX4iZBQma2MdtiIVeItiohCVpfIKQhGZZ/OTQx+bN75lNY0inCDf+IX5W
Yhnd1Zvvdl44lE0go+tsmIiBLOD4YpMQxYF2UnsiQ7XA/T7y4NFGUMxq5POrXjSAkBkCjhVnR4Kl
LKuP4SnHxno9JwTcYCZgc/Ogt2rDmvTNt8/alRCnQXP3GwnJ+3m+HDM+LIBmYFle9LxSLNKVEmh/
CdIka0O4Af4nIwCqboaecDQAYrla8foNF9yI6Htgwsz2R4Q+ll48ZWod8BM9ob6bfwvkeUJZoEZk
jph2aIJ/wujMSEr9L0MRa60SP50847zaqkPpLcUbKXnQOm6do3mEM+o3AVuaSxktSBjzh7L1wJYx
dFZRq8sWTdvy08Wt2FlU9ukKh+hkXhl+veVk5Hgtp5sMTFIkqhpq6bDwDbrHoyGdG9go8eMgkNXM
xplmu9iWAG1nNzA7Q8FpqUBmvi1ogzXRGMiv5x4txThn81VPEQKuUTBprYbZMLXpYV8kU0aZGsEw
j9EC8sr/eQMd22xtZEQJ9991Ymtvo44basHM7cGyrVn75CQc6ffgNBByAfH0PPagVtTCOB4fjNN4
npUcXl5iJW3i/skOdhr5+iXMP8w2V7VX+zd51P/BoHk8ItyngujElvHCzlvdt8zF1HHNmu0690bs
zWjGY1aNEzjtEsV4p4hNO/lab8f1gK+//to8yLWQKrlWzYswwX+j/LYZcQqwSU4McOaKTI69gPQi
3Y9G9uFCtv6vfPT+PatkWzmy1PwB3I/69aJbs3WhKycBdnXHfVgihGxSVOo35Mx1L7iyCu2l4Bii
04fDOHJ8ezOpTcTSB63rXu31vLzeCYO+7yMG3bS3KQkO4gLgPB6X76XckamLFt0YCacX+CvVU6x3
qyRtE0Q3BHautIOLE2HJPfcaLLhtenzqyFz3dAFLB09myk20uUnCLxdL10gWPUt8D6gokOOTEHel
JdgzzLeyjS4MTr9Hfg913U0wcOhK8p/WANLM/kBTsJQJPG+IJ5R1v6DlLNft0bc1XC8e83Jwx0JF
nV1bSeikJ+IC+g298F98SpdCZmtYjHe7XiAMpyhott4Igv8qev9iYof1sQ72TxFzEYcemkGtTcLw
i+b/6UlWhiRvqkdnIR+rfbLbL165Qd7wffO62fZraOHdIlmfoJdKP0EZka808ILx7em04MWVLdil
9D61WIvhmxr79ub6Bu42dnHMZUuCSLILQrP+tuY7zLZjD91XJHjaq5T+QBtsMYYWzQZvddr41xgH
/ATjNb49vPob+PyUp6jVLxHpgUTv15dZxYkFJqB3ageZLyg+VkwEIlhiMMOl8Db3RN6ryPuUga1e
YjxUXcJRE5DdD671UHhBpMYF2UwjfFM7AxpBq+F40PbTUHLLTvZzLAb6dIRIt5ARYqKGP0WJBVxG
jF8lD2sLJeOXBjuB69y7S/KHsA/CAn63XEVWrku4A0qnvbdSNpxZdhpip2QDjwHKhDk6G3tLmHoj
IOR69uma0I3bD2r/ft47uV47m5XGJl4IjmoCU0ruCbrAkye2STELoLclhfdvtme+UroPD3CUFidL
2DMV7H2E1/ZY/FUniSc1TLmYkq3QY54GZ1N0WLJi5kE+T1n4ZargbcA1Dd5tjbR+FfnZYcUudcQ5
tuH5VrN28qyyPKnxxoROhW3Ui3F+RKQOZdBjz9lE0G8/iMFCGlHmb5IJMYchsZi6V0+LsTPfKOV0
w0ko1lg0XKtdoWNONYhmTMQwLOQHmAv+UouFrFV6LiXfpfK6bWy3Z4LmTSSyrG3UtdG6jrAYgm7c
GIPU/tRfMvUf0DzXMvnvVyhyUWZ1LeczpYWUgGec0d+CToeY+JH4obhvI3uy+pqbuyif4mVQNs1X
wNby1iY43KP1bVSTthYtgeWoc3rtHIxsNnaHIwIzobojUCqxdQdinsQMLCJNynm0VwHMUaoN+BgP
7T1dkQacsWehXnis2fduhEZJv52u7NAuSFyDyiUfLy/Lk7hFMe3IsvimzTBWtrl+VUPX3JtuPlbL
GUEAqyJDIqBih46pheC6MXo1q10/A5EaHOHw/0fUqptQfM9jlPnO7TZ8Hhqe3irYOj92bPQvaoC1
ETzZckEmYeuqtL5e9Xg0zIj6hGo4eBDmmQpVz6VfIjI3zzey/x53ejRXzeueuc5vnQKRQYTWWc+q
NH9WocimUlwcku9EkQ+1/mTHXQVh/LoWYMYfoAfzpghqoy35FiIl+RQyzI5SySqKZA4N9TYjwKiP
mYDnnEsAb9gxBf0uHTeX3KuEDTRa0nW8iyzmkst6YG8Z4VeKVWj7YaXjH/qeEfIO2pRK3q0tQw2j
ND8JRiDzHvicKRKx6gIX7aP2RfF0MzwXJSDeq6Xm5FdRzSiZQap6FcCDUrYNbPq+3SVKKazo9WeJ
Ghsf3eIyNvek4I3e0/lWKmGhc/Z5oEVcMZWRsjFrzYsDGywgMoOXpqWztVfI2WCt7tqOt50cjqfj
n63iB8bdVWTe1QmvE42bFKwAV4aJTdX/2i6nt5q5u6FRp4IAdnmUKG/8tGroAYRm40GEvX75TLde
V04PVAiSU/uQFuENFRoQATOKBw0yZmoeWz7JgKxqkGgjkxVBBeh77XBnFHbMTYC83QTKjWCqQ88K
tma7E+XgjVoH8o1iwRDIgfzs6znRdB25eG0Xvm/F993W2otB+2G5SNsBbG/82t1dWXs1sp3jTnW/
odpLBrvehQsq1a6uAaDyRknMD2MtOANpYxQ5nG22+PKdkV/CmqCvRgQ1yRve4RfWXvKts+0Vf0Bn
bRdbNTn3abu/DX62SEw2wFmgGVVrG+4dntVgwyxbAxaKMlScaEsd8RmGJA9FxI1d0/RxvMkZukum
5NhoN1x7/htzoujWijdEUBN9C6G/VJf/Hdsh0G4nTI7gYhKhzn2kKIjOflBob4h4nvITnComF+hm
Bb5GyeH2ziYJ0rFE4fyNUxE3aTa19eMyVu+wvditsEaRP1o0aJyc5LOcr3mky8Fdiy/fhSEsHETA
ebxzPX+H7l0bRFn7UIHHRMw6SpiMpMQR2ST+HyTe+zbwV49YuR+OCFhzrS1TU8LfJZVqmbZ/KWHh
XL7rBTmAvJnta4Ga1W3QrrRfJH2JhYZxxAt+c06SxO9AELgChKM4UtASYkPiwaAkRGjnvE02U2tI
GVnKw9pY72vmeJ2SRiV+Zs8t/Yhg38LHhEE2EyrUO5Faywryroo/mA5vqQpnggk3PQ6X4dyM6wH3
md6gA5OmOCvNLS1iAL+vY+wSK6CBewH49Jvi/q2llqERWTc07OwdkJpffe3kSxF0cel8DfQMrEaj
FPdGMCuEuCn9jOSg26gY+dlZSjqpLtxMwI5w0gNX+O4mwUB4i+RhBBspDg+9lS+HUW65yMFIrk8r
/eJdJyz/j9lsQVNQ+LjkkyNQUHxtiwi81wd+uf7xJpLggmHlHMGIvGqeK9ag76FsnD/IWgPBRaYW
tJgLmxLsddhS58VVuNXRp6aL5CGnn14/RYMvMaRzPFDNjNE7sC0yhzFfklCZ308wQK3T3MUCyZn9
8g1InqVqJPB5ODOqSj+8rAskZok2rs5NgxQIYiZoq6ovvUo6KYT6mWWvUhms3AIOWiiiexrKCEn2
P7lEdUzDJtLZv6TybFOFD/F4GBhuwk+HcoG9nsg1mFtjLAlhfKvD3Yq4nYfLtI9/YkCUoZkyQkHr
3wcJONDfw3fvo0X+yOhK9c7U/ghhHaCpOn/79Qzjqvaggaoilcg6zU2/Gn3qgfHv+s3etj4qEBm3
i4T54N3Q6vxoh1GYM3Cmd6vH60FPxJ0Q29D3TkE8wkbhC4UiWhnFqr+KRpN2/Tkzm0ByOlIHpmfu
niafcBIBuc9qUE/ex2l384/qEGytGt5pvuVqFtxGfQR/6klKFiKYf+6oi16X8wIUMXnvxjRZ/4wo
DrvtE57KeM3C2mDgCPDpMqXf0f/kS2ikGbuZzarGHfrfmddquIFtSZLQf/VZgnE/qSWW9UUROaMm
0aJRXj0winVOdVc+I2vImqxpEUAn9i6oePT1oS8WVuouA3MixaYa001bdt+S5ZyLuoEHMtkVutqx
DW6tRt6qxMVJG8GHpwws/3rd3Wmnwv2T8bdfpRW7ETJDRSjA8OEhIWLjvrnRSBKoeDMnjq3A0G1c
w7PenmwWSqYhcQ5u6hcmSmdvh8f5HwUA+GgWRDst7gxyn1KSMF3DW3qKZQ15Ntakhieinpu0IOEI
jD1tFU/JxQUfGz7kMo007kwuwJl48dSfqH6VNQuWhpRx7SxUExePBkPrWLUDU/YYUNTbOx5Io6O8
yb9c2HLMmvsPqDZOXObuWhGRQ4ydMptKObi5X3hsROxX4gF59259DlBFGlT5+PMtlUR6R1II8TpV
MrhEYTSx/3UtbhNHTFh4CRz35ke4kE/HXLcR3UZ2H9up6TRCUUGQ3DD5pQ97zF8kr9r/rcrNb684
KT7pXOX9JGi1DFKe/2MwVgoJS2PoMUUbHKPnjDJFSgiLBvv8vdAbGyg3PENKn1NOYjrHasoWn8Pi
Uhq3OJEmyQI7ALXsel52hqc/VtbVQofwYWaSRtB/OsBqJ3xWuTM7SZPEC4d2dyZ6zrwf8Gd7VPBN
/pedNLBH9CeBtNesX6V5AkVw2a334wP1Gcfzd0qHGTJk7jiTc6AT/PvXo2JEPa0ij1sbk39MNVLg
QS4rzgUNiEwVuqgqPZw22SovD7LKk8KIrFk+ZykNCF6WGnCoOtSJOtNP9RU2/h0X67KvZm8AwiMG
2TmRjoFgjc/5HKExpx46845ZOIc8KJtRRUwr9bmUjj4/FHmFaHmivUDP6IjkDmw92y5i7DoMvMTl
aMuCfallCBzzGoGHvLJ58UE35Ix2XzhwK+m3zyVsXHP7CIzHMXk8il6SMGeyu4BnkWWQuhPT3VAg
/tqkYIgoxAolwugg/YDhLK44F2ftwUo4pcaTBttKwbaPl6pihP7jVrFpIaDGf28SDHtVJXVYnP1o
NAScdm1YnmMmKT3e36ZmOrzydtdAVlXaEOz5GXqKCT5Z746QSPbvz+aGV24B0D29vedYcYE1ZVSB
KSDJkELyUOO+0Abtd9lfkyOopQVYVIgMbEI4/Tl491/RP9yDc9dRItfqPjBufRket1AE5LHQXdwX
m566w595xJg8jqjNNq1wQ7H6E+zGRkOZ3T0G516fo7PCs4uCxwSNrVZcXfClP9KWEIHN4KyoJ/Dz
H/rPU4IfhG/qmeA62YQnzHel1dKHo/Iak+hAasRQI9rbi2Ln4BgxbSVCjW0kolWswbvBTPk9MyIQ
3grurBINmqbv1nSdKupH1II5DXaDlFS/ZYQVP1L5c2EhJzNkC6ORrTxnaCZHN9oX2ntcYYVZ5OwX
haRFWNZfPHq1cbozVv+SGNP4aZT9H9wFCPtuP3ZFFbOtFV0pUFJw9Dg7vcFBsayPKCbZq5slHntC
a404i0GedB88rqbj/mPXQrpHKBnPpmiTU8Qbyn0lKpe0BvQTDlU93SedYnlesL0hCo6kqnUsou/e
drjbA+2jmNzew6J3YWwMHbBQ4lZO2mRMXa+qfuCew0K4CEUBw8goaQNpxQZQrPEaPKc38DT/p+ar
kzuzp6/dSSeT5StuR7p357b+xSpZiquvFiqMdLZK7re1M4Gv1S5zKPt6qwSXRsRNAzGEszyIiG7/
w00JBpufDVH2GkzcTPp+r6zwUhET5EoSIHPXISAjDzsY3twAZqoD/BnCo/2kcY6j7xikH5wngSVD
fMJ7VI5HVM6cOaGaLDY1tlA/aa1DAcqfZq0lx1YCLgvgvAtgK7ZjCUoeUe4LswkecN3KBbYXaRfA
zDg3hUNZQYtzw6GdIlrYgs3Dt3x37zUSa7HxSmiaxvRhIhz49dssGWA0skH8QK8rzRCWiQrihDr+
Z8Zn4vEyA25qCUH5P2lhAx+4rYMYrmBZgo0O9xptN0cacLblX4ewmAMzLBpe9MLYQpIrS+dDF4/r
0VPCCRwyGsDo1s9aaNggPZaSBfOaWJJ/aO8EG9Op3Kw6gXJgFWgN1kDbzXhoI0V8unIp2oKlrWv0
GO+hnBVx5jWAYZPw2q9u6qwHo8w0HocI3f0dU8eAM8VbcqzOcS5q9ZfN/NVxP/zWjUouPQ0J0f0o
d3FabPj/y89DlM3LstiEneP0XnOQKxyGFEtGmr/1KGH/pg+Jf93Azed714quLkeo1TwNY1IXvPHb
NIsn0TmvL+Hq4La2Ffw1/AqzoLmkzgRyy0VAFpuoukTCwAFvBjrDwSq7xfWwVHRuqv4aVuzKaZSz
6m/CxOSOcmyZ2RIS2m6zCAuiEGBzWUAvT7NhnYYfRJA+pu7nMSR66pC+LEJurQ/A3EoinlOCFUMa
R/HzYsDw1YJjM6D3LRSu16FvRn9P90FbJOEerdTivIwdMn4P/4usGcUCyX9noRVY4QanqXoKJYie
eAwy59xW6cQIyGw3B+cl9wpakUjD63Q7WAlT8kJa06bO80XCzIr5eE9uGEQoMI3teM2waq5pWFr7
yTCUe6DN+ekmqt+B6asUF79WiXQAkcjP8wfZS/op4oLR3iKbJu8MHvRzCCAZEef9xW+MP8nehGnm
/t7FB1GAJCIwFE/aLZiNcylTZ7BY66Wan6nZ9KXEO0BIG4BJW9dHPEByCtHHIcBK8X5MbRgUxIzQ
no3peCD4IA1pLnPdCln6+52zjsegR+8gCn2fbMTfDcePqORDV62sRXzT6dCpfjbMTreyoUUdYxxb
UGYa+roHI2EwIDb/ofd50pGA8QLNa371n1Knw8hl9Fxed5X55bVK6yFfssOtZ3326DBdqVfmUCjr
5rMba8E9+yxvISDh3DPBpGJg8cemj9sP+Yqg8m1xelQD648DS5sD3i2TKWbmM+OkTQ9VZ5x+OrIi
PrRv6gjyLcWGIRB7avHElBfyO1Z8/Uw7H3YUaPJgDVygqlaEByxiwvfP4Gf9mfbw6gu2VZ+t1krQ
10tRnP901KCLbJqUEOfXno8Hx4cgJUJLiNLj4zWsO3yM0y0X3cgODoZO2acbtlqaIxm5ZJ6+z2he
Rfezqbx9fNqgXg+6mzTyyGWF6IrP6XFSLbF5s3/F85h53/FdmCaLdv/EaIW5oG9rapEzZSqy3rHi
VLiUUqHtZdsJY+PZOkOw/OrCwWi5Phj9xu95K3z/FoEWvctfgpOSn15vNpc3VMeE3M81sWSICZXP
2Mrbxr+XxjaWfUxY7jMuTMken/DEBdsaBIywUphPNruVYWHG+as95qIjLORKmViDub5jQCZ4Bu5a
jr2N+OLEf+GW+TiI5MUrZywZxaeac2qpZeuYC3c+uh4mmh48S2pJ3L6w6jNbWTZk+hI1K9J5tSgZ
GkpkgIzFWRN8d47+nwHG1Yy5xYefvvv4Wq7JOCULlTofvFgkUbJDxpC71tYnz+kfMTvmykko6lJ2
5HnSUtlSY0J8/PDgYmneZ8pfNC6ezXZwvvzvhOGua/GwVTUfgaK5YeyezyQyL1IGO4cRdFQHMZ+/
K1atGad0SqonqwrDaFS28wwsfPiybjbdF8MCV5Ost9iNt/lu92tYTcP9X6RjY6N4b9iwO601h5Nc
coYJvH63aCbnLE3wKni8pn54PsFGZ4s2oeoQgHvnBtRINT+8jMcEFZUeAv4vZm0Rpvha38mixN70
ANPzbrs8WOuUFBHiFQJRmrUjAeyuWRXw0VtR4fAMnV7qLuKnXpAACneF6mbjMi7+wVswQZ0hlbDX
mk02CRKMKxH5Sn5JuiZZlzoElIoZ1mxcF5SGmh1OkmTK9u5mEEwEuBqZ+E5umG07IDvr/zgMlEjy
rvOosHhdCSdMRf198ZaMMiZNtB6nteQERvfWkFxV+pemo9yth45GTEM0201SWWtx8VaQx8ySC+pC
cgRdYGtyRqW9sqda8usexyQafsnn526pheitT728daht6Qu0qK0JqcyglnNEieS/QwIrhnLjM8TW
7afrQvUoLVjm9ceoXYpbG4HsW2BagWvpDFkMxZUpDatYntlLeBXqnOuca/huJQ7fWuiWsDWYhdW1
9NU5kaEs1u4K5BWoWGQbtAUtIHNA4jZaIDq7qVxk9vAlM9EYxgZutQpAUL5DnIo7dUgRK0K3LLJ6
6hP94sEWHoX5x8aZJ1vTv4/aOiTa3Is9slyiN9+hS0zRBhCiDNjnGjkjFo/Uzn8fz7ua7FwA9lzg
47Mp5yxfse9vrlUGt5I6PwCZv0cuyh5O9iGfmH5J/GkwmBUbA5M2fVl42sA54oiTelrOPnXG3syS
JJ8KQE2/Eb/xllssRV0mtpDIgOyaH6GD9RwrKt1olQbYxVsLLWuqlPeCajsLORwspYdAQ7xKd3sZ
gqcEV3pCv2BcS9Q+ptPA2oCH8N80sZkximsBFEqLRtRAdE8sdmkDott2ptLE0xkrt8ZzeaYJomcL
bZt25z+ZZtXJSwPtEoIend4dhQ89djLDEGZyYw/Cq/fkzfSd/L24jpb6chGBbsCgP/cofMHDGv9v
KdYEkrUiMN+75hKNiP+2KsxJs7zeDgn+F8LbrG8VuXiej3hlgRkQtLkpDxOG9Ef4ABu4tXPg1uUw
Nzxow6n4IM1CBnXk/bLQtCNPmQZw7bEGvIwa35DYyR1MW391DdAg52LtFfZ33PP8KmTZXnDfkd4d
qmpbePYrx/SCNoSbYpGdo6hla/R/DSoksPsDRx5QSSnBs5X27ejh2BmO6ptY1NmwaCXHy/XU0RRn
cxxx7El562QvRkmxEZcpzZuFRLJ+ASjYl9qcQPNgJp56tZrg4L+4/rqLPDU+qZ8Mcu1yM7p67f0y
h3GglawXcjET7KBkRhCI/QqWSv/6pB7pNknZIRUh+qz5ulM3N10+BWLu4wsr/chDQTxYZYI+I85Z
24A9fXkwil63siFjNRo08ah+1A/mESvRAVflwwNcKB7VFyQ7KrRbHQ+ck2x+JOoOpAUqcGBlG0PK
oO4tnjFb+dbMfHkuEWeSpkcxLsVUdJFC5DYzLf2cM9wZ+LwekzIY/gU7BEMUSlSt9Zatkj96o/zU
KDdf60/sCMJGAb9jPKHx1sHzOEMJGqpcDJVDJjuSxW5YYb/gTIKemWcx5Qv0671/ITLWH2TNrL4c
E/F76WRn90gQWL2bVyvhe0RXonVZojp0uz1MYVMg8Zi5I7ikoZXU++crTxcEMXneTkgRgmF9z/dm
FUYEaWDR318VBpWlIO22dre6XJ5VJVd0gwlUjA7NBKaZZCJ0mcmbZYqtG1aW8iJT8dbtE4SsFQG6
9A2Ojy+4tJqm08u6yXJbyCrdb5KLI4Y/W0S3Ok3clXfRCo3i+BlwKPEca73xWdJtGJw0GUipsTWB
0sZVsYj+UeHLQjgZZ/vJmYhB4WxAbIojbuVbv41OKtcHtLif53+z1ctaN28dGv14cAK+I2l9W0n+
qfxxef9huHnKUmUcunEFNcSiDZRF/LkqCCzuSsb/yjD1sxpNooMMYnfMsWV8fSc5toDJB2FmNL78
WfMZTeLrpJlJ+m4tj/pYzCRH12GJyO9Oa8kTlE42oOS6zThktGxr5O6/8gzlpr2xsxtK28BaQbRT
vkIxXEigasbMuZDNmg6jdFZnS30oobx0fmSQZfEbB9+bEuP1/rmrtcj5nQmI0+76O1YmXw2jaVlC
Q6s49KiYvZ0SM0FtEejtPLVbRmX2Xr0dh2QRiERkxi2fReTcS0xi7YwsjVNVhHHDr4XvmKnwc+BU
789A8WzQ5RqPBVz3wBRCPaX/9zsxVpFArcPzTusJrSxTNNY1eZmws80l4j0XvElJcy1n+cRLmHRV
9qs6CMHelSuVnULNDHdgiJ2qaAMgD2pQVlQHhWLqeDSehDz2qevjv0agGvEBVbQNx3qKPXDCyEh4
8+5mKDuO8qgDfwCrNOWVvaOr2F0bAx7ThQi6NuU/KjmrKTcTlJNq0Vx3nSYdag7cFlu1vx0d9B+e
A91vKZ5cn9o0fX9C9sHvohBfhXG+O5iJLnO99xZBMD1X2lwbWeIl1QgPIM2eNER7+F7DhzTt7tdt
B82aLxO8TN6Bu/Ayy+xRMIRAUWaqATR2PitEpNDYzQp0PIPbstiAScSOyD6f2r+8pRobVHGQYSHl
Pr/sn/sFmEZjK1zJLAHhn5ZH0Q4ZFiOA9oCJA+UZbn0wP9bGYVjsVgao6dCSSjAdVI7AO5d+3gLi
aqA9SF4NoPepGatDtUkD88BSuRDEljdcU0CaJ18HhDvPz8GkjroDgKOkuf8qMo9028mRx7a4tRqg
CGVhxLooXP3RKZblssi34GO8RkuBibGB87gwq/XRH2US/TjQMr8pyw/GAtaf1kpFt54FiKcfO5/s
Egxd0fSWKP9Yy6yJ1XI1B+eKsb8QCqxiueDQNVlz6lLNnfi6mHvhszpUHz8h7DsBDc+aBAJhxLSC
y3PhBr/eemnR+0HM7ujG0M41mvAG9lJKTnadRlTwbHp+6j0E1VrZzQ2eVMlDRMf83cJqLPBpG4Oy
doBLA2VHAD18C+wRH11kIqEijySTCA4qLjExU0yZYYPc3esumLfUC8VWWi6sJcsfn2xQ3qB8e9jh
HzAuMa4lwo7DfYU5GfPxiioI4/Y8d52UNsJ/6FmHigseLd/npKpMwa21hD9ne0TRxjWi7twKJ58R
Hq9JEa5Ji42Qwiy8684xSJ/F4VBmtimiHn2dYHljrh8CMndoK+2gSiPu9dPedgYWDvEhdo96fiZu
CCawdpfbfpILr39ZXsfNqifoQhR+J+WCAt1pZ0mHCiTups9e2XvNijVQTJcRRww5rp8AjYrH0pSc
FjurZJXc1z50Njh8kd+nqblAGRKn8g5KDuWP32H2MW57S3XsXFJtVcPQokuKyjvTPPNyMEfybumO
HCI+O+QFCK1vLGlmhv/HXu7J3gi0YXQksDGmqgWhiAin+sbWPpoVR8Er/JRp1SDL1R+JfD+aqswD
YtdJmmKelJcPCPVN1e+MN5/R8vRN87aNHFO9fY4IYdIkrHuz0LrWM0zcMMBLQZUlIq8CSB6dAP0X
jE1kRi19/MEH4UaRuN043VvNmVKKnSHNyBv0DlXJot9WcdCkvIcpGpvTPpd8EjVkezyUz4GSw7eI
zEkkCSBO7PL6qAs3UJ/GBQoIl3EEBr4fOCtD/7az5yYMoiAov196uXWwEZXOFSbgOfwx9XtxEs7U
4gZpZGi5njx75lQuRnsVS/gpRfhWeDeezgXsQUeTsd5mdtFgczBVzyvTrYi0VtpIk7qtH/KqKV6l
usjrUFAUIU9sdK2XibX6gITNhfD0WfTY/cADBSBbuPxUe0/oy6mb0DuvDUlG8ZsMzmwxttDbvNoI
MJIjXoEeKoBsDuosYk+nNVJ18/9LxucNckC48aN27H7CrBxxlsI89OOIOMXjc/s9Cr6+7RGwTT7L
PiQlR68HtTFjEDA1uD/eJri5+joG4scDerTG4WQXxoY9L/4ljo9ggPbMOKg5MWs8P/PYAjf3yWX8
4nL7F4wFDWxVFXCfIduBWhuvrrRCTeqxLuVm3GxxuxiFhlWSUR2Km2GMEEYEaKKX4ojTZYo1EDV4
D7i5OBwDkkTIEDYqy7jrzGQINR87NfPweychvCj3MwnYqDjwsF23jPJA19GjgJq3Wc3o0aZJnbjQ
eFWoXa4U8/y0jXGhEDegeWjBLR5S1PF7yT3zj8QbHggBR2nA5zqaeerAaFGEf3lPz+Sp9myhWIai
VJOQgIxZspnDrMjvO8O14QTMAsSWaawR7r8Vrz0LniCUpyLlXUpHqfDaMlEsEJc4+3uFDTbok+lP
OLOUrTn4hbtLjJatK84033ErsF6YuSL1M2EjKiGFkvuOYokXc25c1fALWEV7sfb+MAzGVvXpYOSi
Ohb4D/V/VA+VpgsgCGx/kFoMhpmjHxOLQRn4KJfGYxoKau9qr8RYbR85S1MW6PNAJwAUONXHMrJF
/E5HC60NQLYjq2X3tv3+h7WvSTAJ9jSYB7XWudeAc52yBy8AXwF8wbznzqXHrW3Vp7ddP7//IPHK
UUMzYxpmFCsyHT2qbpzugD7SWBklxpIBzElUfYcgftgcz6yv8UpQ0cuaw6W2nQSEyM9todU/pzrq
5PlcyD9vPXXMgVnQTReQPnlJkIeBeyskcr22Uy6mt0+TrN7UFm7V5FLqvmFu45EBeXV4MR2XmPaR
iAaO7PLw6Rw1N6Bbkfa4li+g/PIoKwbM5nSpWOsCXY9rct+4OJYzuEXxq2dNI7llWT1qFiJMwWcP
N3+OcWAbvnY5et0VxaeqDNOsjMUIRzayoWsf4jgDBmc5j8A+P8MHvYm8lOT/gHSqcK9WYnTrRhZC
AlR76FfSoKcPiWCVG5stDO+FekHriu9Ku6vt2jxC6Levy7Cht2K+LdxqukCWsG/SrNUmbkOpF9KD
qEQM4ix83HxUp3s5RSgrYDddnzvyqAgGsecSY7b50lLK/2nyMkh6zsFmwlhblEZEJA61dcsxc8C+
wGexZLek0LDspY6q0I2vnNKAeIHYmGEfd2NS8/MTQJiqfTUdAxapwqVX3Jx9ZLmfhma3yMccwhHU
kw97r/18PJNAxqqQQRnUT0wIuMp/O9IQvuteowj+0pVPnGa4tm+ZAhtapPnuiZGo7kKgIRRidral
AW64f93FzpfKf6DCyHyjTUV+QOmryxd+ewlZ1cSsAdJjattoWbPbQ+uA8bM0AcOoV/4UDQbtJdPj
58tpmVR9Z5bIlfOJ7/Kh/KmquxNDG0P3tlezgGsc1rrosOwu+nGYONwb+m6Cfm63rxvb4UsMh4sJ
HoxeINRuxRqYU7nErMUF+QC3Ro3SJ5ktR+n+XPmWJ2DBTopi0p1oOckkm3jZhKo4J38i+FjOzT75
8Y7BRQpVsr0pNwcSQetkqLX6oSAPx7F4YRZl2qlqcHZzpd98tWvqcovB5QcyGheiDJVvN2BCgGeF
bm7hL6ecYXt11JtENyKBF0hzXLEK3o31QAzY251WqOzWqyLYyJf5J48ZzNK43WUkrAnZJZ1cnVn7
mxsPfy7XvzhUCWqfRtzX8CCD6wYCid3BWhWUkNB37AyCNIBEqRDj1CTlkflkMhNV4dOtZMCEISeA
72Fk7TRZomXiX0aY7iXZvpdEPtUGeOfNCfJaj+BMcY5poDHC5NaNB1D2+VNAGd9xGFr6fvDuab46
ArLr1AE2oBOE8Zn2hv6DrZRFF/XSB0tIePYrczwTOm/qGpEbgkD2BOjltUGfG48LKRkd6B9AN+rY
iRH0BnOXCcQ0br999oGjfzFAhY59Ep7sAHY8tvx6ifDMNVSve/FaurSIHiFoEHjqzAvY8fOGbi5O
hDnY9753M2nCLaruyL6F/IeGnOwQfKJ5w8m1aDEzSXb/P6SN3t5KW6NfGQAeANNKIvsuy3DSunuY
WTwDctwwR66qwB0AbCPoKOumJx7ZuFpXiUG4vdZGg0nQbvkwvKC8hZ5bESrLcPdkLI/2Cmh7jDOo
CQ0V2WWYFFtVnUFpp+ZQTraBrkSQgLbb4rkT2QXxPJ9y/laTklRYVf+gs2/eeunaWdQHprpSQ05G
ZgDNHU4kFZSs1QWTYFRDhkzhve/HgE0x/+lN1O95lFs0DcSsk/hI+1ntDJQrq9MnoL2+Ocjl88iE
0FOuD3WBF2o231sxnbR5l6Xrxjbupbt0RBJgLaZqBODZIFaSQLeONVQco7kpebwtt+jnZnpaNX5L
smWpwUu5A7xYoF72M5M4xAtKYAe92ZfkoqFCEkTNDljdkPa5go1n8NuxT44GpzM7/y1JuYydYgJX
xFIC52L1uEOhNA0TqrJnPl6VBWH2eIOXFQr7E9v8t5Z4CH8j4+093KjEJPml6lPYQig48VbAPLwU
Hz1lUZ2UxpdXki0Spaqjsrzx4HCEQOmyw/tS8NLXsKHw8sWQ1xLJ6h19rBYZJmKpv8irUzJE95lx
/rDibSaWC8dCkQav1sA6rDnDkXifiznQBxTD3/rLvYET07I2lYMb6IUIAs/MwxokqD57Se8CrD8o
oFXYGrD1/mHhHgQQHPvNrj0F6JejHzRAghhUVVwayFnWoR23RQRDHADvIuWfX2nomTibZtVU0QXH
aEbgCXnSh2L1XKWwWN636YrRr6GiGtnqbSpA7W6aym9UZHYtg8eYD8ah/EfKjXNTziVZioDMi12z
1O/t3j/46VNQq4S14mJ0aA0mo03Za/lWr+f+nhs/gaz1TmtIeb/q4AdDlyBrX27125CO7XYxFWIy
nraZzNMEAw2Gb378RS1XoSokRuAmoQmuLPbD/p+6At0RNbaSr/ImQ1K6h2JSwVe18oxHOuCq2S4I
FMcOCVtKXcT+ettbWeIf8DF25HY68uCO2TF5qg2+6ZkuvPkfjO9s+5nHJFFJS2OtL3nlfNoLEQiI
H0piNQvj7wn7MrmgTfOtpBfxxzQNMMed0xTuwQTQvS1ACno3re0X/Bsp0KGG0cV2wTj461lFm9HI
64xpEV2oJjeacwlK3/OLCv8uSq8eTOT7JecNke6Jvplpr+fgsd7y3/yuCcJUJmSyUBG9coHY3uvj
Iddo27CXmnH00wsZUO5FnzRHm6KYz+J02bQ7eT2ZZba0iTJeYCfT7k6Z3TGaAfDsF32SGqyXUkrE
VSpeAgqpSahgoP+z7SSR8L8GjtBYWTU2+GJezaMgfkWAr37elgWHwIMR3OqNfqNlcp+1nHCti1V3
VQcqp4kqTIZnXOKsCqnvx7D/j7E4mDuVX/bUz/qMDk/H0EbKzCmWhRH12A7g/bU3KjhbccqNTHs5
zk7/z5aQyp4qv6RAZiG+EPuNQOWZPznEmtYOXwVIanRtZgTXopg6CiWm54tgT6URf4jBj4mR9Vda
sTYmAVd3XyxW1aYC0nMv9s94ze+uXgIZ42XtBPh2Q/WpZiKAEU3YfeL5uZTT/pMa8g+c3ttmcnO5
sO3ydyvsyE5/ObB+fC3cu0Gm+wJvx0TShPjV3t8nqNfugxAvG7iskYwOF4cVX9slG8ThvV/tuWmg
KsoFJ4RPalCJUogvm3sSVc8vDLkzNnAWpo8J1SILrxdLR3Fa0Q9TBvou69m2NtWoep0to1o4OSDU
foHRCYJItmIjMq1sTfny9cOlSmjGjhgjx4RiO1DASBNzUUo7A/HPXDo0DnUh1LAtzMCTfCGTRaTs
tDAV0epxiH4FgSObN4OPB669e5DuxvX/q/ffGZskf5t5eVMFIFrZAXHBRjsheQXC6WgoCO7n43Yd
Ge4tyF/1yajPe7GYKGAQ9oMyNCAYkagOJ1tFOKcz5xBTnfpKuTytmfoUK8xT86EpZtsmtD8ChZzV
/JyHnBVtWZPmILXK6gpLedhL5d6xeV1oQHrn2tfnBn5eDS49l/feYuqB/qBzt8QSI1op3Oec2pPj
3ALGdj+ygtrZydH/YxMhgPKbc9uxp2hCXpSw4LU9/XbXp1UvzeUGnhWopMMx+oGGtRM6X4l9tuoq
DNLRcqs4P93wNRt9DT9chCTHluxs5nvHFeuVKc8ipaUP82uaHDdePaIMHZqNH6/fusgXAGp1t/UP
VNC6Sy3sTV1N/KghvNVZTVgPMAz2IiKnrRQuSjLdwgd0FkcfD98E0rkxmwr2rVT7Qt4gVNkEFASI
/zM23/iQvdksLeNLd3tdcgbRfvZGDayN2b8EHGDnbJOEi4Xntp0bQEp6cAaCb1Rf+ZdLfDVgsxgu
WqoWO6EGw5SiypDDD2bFYIyhZSY22RGmSKSudpRmZVHI4z5LkfJRchTO92//DiQEC3e/sVcAAh8r
gXUWsUhtu4vnVRqEU+UWBVhqDV9tJEqtYdaNEiTuTYxdw9BzleliWu7YaZ8SSHVzyyG2gR0ifvt8
fBpdM3Ga+vT/fTEBNKX3UaDX4ZZsHiSZR3cG8Jozp0bHA29kERBwuOOgFfOuwVzABWCd5RRzKYr/
ZIsHbqN3iQGhsoR8KdeXAfuLp7DTBhaRDadv2QYl3YFfBKuV9P88iX4uf+7BovxBtnNuzAc2dOxQ
dGm/Es5d5c3vfoJIDaGXkVdA+WRYGsFZZSjZIs70sKXGz0Hiq0rb3pCyBq4bW9c0wkx932J3L/Av
StprTMbj8JWibUlQsfhfa/HWdNw+nXIzxseokc7rHrtaJ9v6vFW8vBikiQofoatS87J2S3bfzK+1
RFxfSDRETdu4qyENLwSnHVucSnG04uUIGldFE+uXlLct56LqXjNR6/zRnGaOiCSLw91NYJOSZyWs
Lzuq/AfkG5avL2u12LcE+Mai65VGJtV5hpXO11A50ZCGDFpl2BPmHDJBA6ZIXlLJlDfLe1+vx/9v
yqYN7vRjNh/w0eL1Rqh4aep+cYYp5T3/SeVz59hyxWvc9afr1R+vcyUkkhxynxx8nXM53i0QIpf/
alr6FCfthas0bih+/wnrAKmgTmp0732bxinr008DH027ItlDjQCG+UmohcxYwKr9kHhqU93cM6nA
bPFEVk8wkK5vnMLigJKM9RGgmoqIpBWjhkR5crsQkqScOyOVf0bCA8lL0hhRcyTlkDyMlb7lyZPk
DLjiysfsG30oOUfezAzPZq9SdNTV3n0B6/Lcn5ts6B7N1CxUM2aCNtT2KExPhs5911ZnXcDHTiES
0T8QL0yk6p6MQ6Jtc1hBqLid/My+yIKApufWqw8yNAgLJocAdp0eWb7aGByIsERMTYLOY6HQY8tP
XAu4uDUpHkP9k0I4zaqgPcTBIE2RosGRzHQST9tCr6DEZX2CSNHCOXNry1DDgOI7A3CXeCsqnITK
czui+eGrI6APWKxQ130HzlOwDnVYOEEXUNp3mX1uAffhTaFq5qRcAoPTIB4WSMc6d2rK8LAE0S4j
NemCdAXZphhkuXjcgPVk8VtAm2vuTGghKXQaD6cFtRjtF8kLAjQsUo+ePNvfRrUlvuNyxCKf6kps
BpNVgeTS4dJKJ+DWb8KrSBV+x7eZD2QtBcuy8AYJKPn20nZm7StuCfvnOAm3bxx1kQNPwfQ9W6Y9
oEbZwsgpcGSCv+ulyzIxWKiGJM0MFdxBgwMouJbdR5seylhjcfofmAg2daoBxi44Oq4IRW97fWok
JSDqwgI91dZ2cj005+W0FH80hjDDDlGgWkZymt42dDVILdDFJ34tc0K+8F1CSsM1jsYBERQtlV/c
LKYk9xXm0oU+hglJ/oKhgMdp+MI5J+/S6n3waLjfHhjfUayppjKG1fcH+2WG2A+ovNcrJfA03g9P
c5OYt7gXrtQbDzmWZV5BbBdt8VkYjQ8ZsuWUfQknBHDIN1w7zdpkyZRDWbXsTWC4b30BsVqMOd3Q
WDhCcGUdr2iesed0JZF99pwso93Si0y+okSJM6OifoCX5PXZJ2F1IY7vznqq7FxRYV8x6Yc+yiSP
OmCwRRsRgLi8yTbbBYz13EwW7Y7YpyN3hNohlIQhhe2BF6/Xc2QyFR9nBYQhE2J/LoaRt5VLiogC
cDxuMXo4spmB45Zbu5EvAqGcCsPcv04FzSCPUfCJDep//zplEe4nl2v89R74W4V+0Aw6hauZ37G1
IAfOFoOTil4Yp4NVQFLqgJwsM2J+MhD357GmWZTqv7rqBSUpkad63uF1VTbFn5XNM+QhCpZW2QQL
KtIdupKAAf2JBkMurSmX8N1vq34QvBCc7HZe3LUZgKoZjgQPHtYE4KpbJ7/1P+jOE2VNifhf7Q3L
eY7pfPmmjuvxyYuwtmHQJbvqh1YolEC0l/tO6CQHzlG1/bdzFzK5/BQdCL91gE2Rhc/dZdTZFdgt
XKerwuAHQUkogXMq2W3rn5+A5K4TRAdhw7ImbdXULbEAn3YwbyyA0ij/85RisoCXIkbaXd+zE95t
doeh+rKZjCzldXw+LtLzvFi4pNu4e6Qwe0iprOCY9o6S3CAwZPfEVXoT3IQD/NPoh8ygS7/PX3e5
XvmW5InjdfWWtaHjR9XAkH2zY2hZa4Qpu5uWZ9k4Y185PU124diuwdx/bz1ZsMKSHOSwgvoAt7hu
681bvDgGPp9quNCbgZyx/bfZKKe9ZnTHPI9tZPPMK4H2Ozu9QHLYjcou2XrfYztWS1n0kFGJlPjS
NO1CKZtTXqOGBAy3dT+46oOtCzE64uFvs8d26le59DthtH/qhGIH2fjB4tWsSQ0viH7AmDHFPZDZ
8g0cyN9CDUn3h/K5rpIyrajv2h8YPeqN924Bn5UKuZqDNwXzx74K5yQBV59cCKl606ptXRc3S54z
f9aYOdes33S3KlRp/jjgPcn6bPjiEUPHDiNB0hr/dZn8MdVbIeuDeZmGFOQ7QppLBLOLW/Dv2Lks
IWWF3JGwxzgjLKaKHKqIeWXWXyY3soqVTVxPawpYry/BbhXvSzkwRqJ9K35BHNL/lEsqRgxDchQv
QmE1bf4r1xNsuxgSZmyFYJZ2G1HR95tl8JM7OeGmL07QQNbxcx7gIPq3jP6YcjwieSgtLox3mKqG
n8UfULfpeWOXjYJrdwJGf/OYluseacu7eS3VJQSaF77QD3ZvmPnF94jsPaSGZe9KyNAKk0sXzCDM
QRrowBCar/5Us40Mr5kXVx7Ge6IxtR/J6O7luDW0LfydnbOc/k5FEQoxq761M22XOdnRGXx5q5Vn
p6DKSBXU+nvgywHr/HApnK3YbXGeq9j232uf/QRC2fx0XN8LKAoMvRZy+pIh/RWHtRV1H9z0iH2m
gXtc6okBjm+zhvja6rUfQoY4Ya4wwPHEpAGhVlQFRaNXqBmNDSY9zbkKadBrxyhRGoKbKidmu4uj
bSQ4Q/Cima80CsAc166X7XIPp00yreBw8cs8R6hx2u1PI8PQP+d+6OKRd9AdbxNGXxct2swH25Kq
utmklsYdUDNycDWycnqRsVU3PgQ+gL2MhWA6LqCFxDuDVudYDdmgivy4D+qhDyHBcHVtJ3H01gls
Kyafe5kncBlc4jgJm4KxaUsmnJCRnVmqRlhZyY2ew236sHX1w80pHc/idMxFrDnjQG5NUy8Gt9iC
DMkjtBsSAMRizC4vszGWI1F7cmHl4tQoJlLtqvmtmhXOdZsh+JsviSYHOHDbKonBoHJcA145CBzB
CsXkd3KLNTbyJ02OTvyyfDTb0fwAG/GYJtPJyfN6rpura4mZtEwbmMkcw/RgeUWLaELi1xjUI9x4
8v3QmtsK08zc48XdaTwS4u+o4y0ko+1ZupU6spuJR5RupCdh4ThIp2CWZpIHKzADqo3oZ6yMRRTg
99XWYVIKiMaipQmV2iY8zH7fVhwLGVMk2cVCHMeganhtgBXNURDDi7JQwXjqnZ10UozPCEbw2ZLJ
+gsQtZ+OYdrBYt26SP8Ox+L+MgzjZ4/Z/69jUAt+lFxdPDG0hPSde+6VqxWTZSQuzIgpUO7ItjXq
Ow3YXu1y7OkJheojvcIvfZhWhAqNaqnvjbeA6cxdRLMUNWd1aQYWSP6pkLdWPW2t76vf5JquM/L3
8NPOOo4JsToJ089q1PnJwuplOp6aLT5epBe7n58v8HboVewTap9ECiTINBMSxDavvQaT3avDwhhy
V7mf1MI4DrhmLCGB0KjOHWDMMT0Uj/j3fGGUOxlS8TVrlL2yFi1gJMnzwxr3CVMR24ubjtJPOUXv
zRijCe1wtgti70m7huvWqCYS9YmXa3TAsEh6ekQLON6NyKO0C5gnkp2wKAbtvkkeS4C8iKRPglXK
Y1UTaFPyaX9IiQQQlGmfl66iurH2Z+99AJad9w36iMNjVxobyJRRmj4kG2LYgN8UAUBpjV6A3qKd
osuhSZe6Q3voct0Z2itTJ4AQ0gmwsFm0ce+PjLwKIQdrOpkGCfnaiPCn7p7W9/taUWAA1fja0FbX
DK/gZcTPvX730/BbsC2z/09B4qKGhf+PON+cXVmzaVc0EBUQTXKvJj6CwzQtEbOy+XtUsWrR8d5h
qzLYh66lPE6EQXwJtHdXSssq+8Hmc2L1lOpsh4kCb//Si7Ia7IHAsoYeo7QinvRn+V2f8CJ3YdWH
A0rksWHiWjjZezViUjYIKNfEE5NOu6ScNGLaUO4Cavvm/PU35NWmizLFLDfj8zm2nq6mA5I0R78F
UPKj5mWwMOz4tqFcJumwEtYXt3/40MlS9Z9CvPIiy5nNP45LNkR7c18CgkH60n5TB+sJu4Ebzrvd
xYYUWKQqypExv1gHLGAcBhY8ORIr4JMiHOawv8+K4StgpcVhaCk5hkEQ7XSl3mq7WsdUJFWpCVlY
ziwBQaVMHrCSZhX1K1KD841mhe41jebYzEWB5sRQFSwULRw0k97uVSgRJCQq8cyCx7sweJD6a0ap
ZmpDU+4WGOoa7vrSGASM3oI+bWQSY6rkUoR5LdwRNqjiy9LBJKUjYrP5YoRH/6rkHpkeHO7w5uFk
NzmKMzqHVBsa+JaF001sdvO5CXy3pHc2EJzi0kQO4LzuyBnbIfz+CQtZrerpJwGg2HhD3tfDCDPh
2+MCFbj3GrsyT6ArH+BWHgoDNCfgwt1Q2kxXqZ8sacSVzTJL/N6OIUHe6DDYQCZwHEmkGZNoGHQ1
NF42K7WC8szJkYIJxenPZDkBlUKgRinUDvLVmkD45k0cOK+Cft94zz09dg4cJwQ/7gXjZV9CEVfv
TrV59DWNgfmzVIPU4/62y1WxcusYzxm7PxFLSkX7tJ8VuyxtqPQUTRUEgj/m/G5A4O5TDoK1m7E5
x06W7Aj7wBfL6DM4c/Bs3wHFaPHKWRJCN2YLKh63/SIo5zqNKoguzSmM1WrXwD9DA8j31ipFZ2PZ
oBVXc9KWGKoNUjno06kJdYaSfJCRMuia46CYyqY9jRNThoI9f3TsJgg0kufFG9YHFidc3kf+dFmk
vWhrcT8ygdOWgtP61npYw6kKPVWLBursuEbuLnwO4A0t/WkMfOA82VdxQJR0jK9TIlSyKDmxqi4z
uNott8yV4r66oSG2/OHPhcIQ2Yrv1H2zM0kQlSeUxo7+4qQj9ENrCxv9PK3qmRHnUKnvdYuKIRUF
J5HKXgnyC2QnRKKGNJi23XctRsQx/4Jeci4fc9ZMsaJm284rhyDwRdTSe25nTUEjUJ9tzefYUQgO
4GbGUly0sUPYvJcBj46L7VtGm/Sl7/ybhUcP41nDkedHv4b92rIczMz99ceYQKyjAQRDCrfKi+zI
bBfmzRiMFkc3MQysvy8z3ViEfhomQlljJlzh1eaHt80wkctfp4ZCiwqOJCWpuOlDZqqLAraiH/eq
IZVR3z1YHllseQMoIYstBb/f3xh7U0dJdW1nCBc94LxlQbPMQz5EZnHDJcPLUW1CmylLyuPaAReu
oBjfWK+EnYhANU7rj45kfGg47HsdjE6XVMisjA8JYDadWomuR/Jtjhzkc+hz0pq92mAt34Tt+4rM
hlZrCtmPp8YkuiR51mnHm4iJ+Oaj2pOBDzF8t6osJuz/itAls0BMBtrgdR9azYdebRMmQ95i4u/E
qKFVzSHJf5i75gSVieIZ1Cydh7AT0M5dZ4B98Dj4leIClaZDRZT6SdCYDUXPVMZU8nABjfPMn4N+
ptcI9a71PM77vmtBRNNfydK9XWKWfRlPlETGinkuaFfmw44ejFpxTt383ZPvNLsRCcedawhmEXUY
/ektPjy3ElZxiuFS/xJY3zE94sLaXMMUbq5YsMqOmJdJvT1DXOW9YBDD2Tuk4jvT8lCWCropZmf8
Xai4+2e2RPVgfBA87S0VNK764e7AJfVxvIoSBjOoeeydEbqzwvo9NsLqQ0mP9YTLrIYFU789nGks
rNF/FAg/R/hUX4O6d7ioNb5fuxcMl967/kd8sChFh+xJK4Wlm/341p6czXYj+3SApO1QlxwWSReZ
AQkIW7Tjm5NYxKLdwgvFqXD2HWtq3UReNxGJFkJtvLxZS3Uj2gDT8nFSufbd0eRagmPUKcNWREKL
f89/q9FtRnGukXyw0IFgNbNBBOWq2X+HTg5geoDCbynQ8WgP9NfU1Ttlkq8Diy01MTmbq8BZCD63
6lVq1CSvNn0cmrw9HVvlc5SaRLSZaQz9yyHQLQKUHVh+8TraSDg93sItLQBhAAZRdptn1RvkXwP+
d0vgvEtG9MyFxmij27/IrEbF24VC//03BL1f1+w+N8J9eSDaH8P9eRhgKLkCTAvi2TQce/1HYxsV
yF1HrGWx3lGqUyYHNK5AZgvai7QIqLQFre1iaY/ZgCLPdPYxoJAsP8lnIixzRLUl3pgIMivd7Q6W
5jJZ43EOLkpb4F+idJLa4TK18aNHrotbSBCUtuG+9rLultEIdNF3En675tuei2/FFMWqGF6QHNdC
o0slNZLLm6ex6eAclJRIGsUXlWReSDNI6SZ79fQ3Zu6DBXKJl8qUc0YR+vJmFVqKgUanrwPLbTK0
e8N6qm20OycNqOa28e92o8/FR5bbYMku2WfkpeSsERuLrAhkJ+wgwrvqbOeUsqyrN97o93ksqHrM
nyHJ7zwdILti30sooeKAh6Nd/lV38gqRwqjsau/CAAeb2CoWDfVTsxbI9erHEjtmHTTXNX5y2lEj
CCLGJFQqyyImvVNwlPvOOrUONuJC1KB/rF2Ms2LWP6716lyNkHegpyAx6AfBO8sVN746aVawyHIU
6+2q/WNjLGSphUccNYAvryjD5Da3O1pPmDeHHetOq2/SVdjQb3F4K5t4w69pm4r4y3/ptCozEFd+
La+AK3Nkks8D61dOqyDihaDUC+ZJyMM4tUnRdaeXmWhPP4MAQZHf1iH19a9JjhL3jk8gV3x++K7g
5mDk08ryofNtNnrXdJS5ayLlBMT88JqtsIaoWjd6h4o3lW7PGeKgD5RQyIaErL463ISuk+URemB8
Ler9c7YRYf0C2vuF9LB5+Q57htludxRYMKc3YH7cwTzYEfx1zXv2TKcxwec1H59KkUoVMeTvSbch
WFUZ8XaOHbM4za323Lat5HZfiAhEa1HDAqezKkbkWGm7qHZRCgaDflCVdJPNr7JMY0hPITintsD3
HQtwzN+mXZnrhyxMUNzy5N1TNsZKtR90nXfhTYKoVPnKF/YWAdAGDnt1soLvaN2I/T0DhItBETQZ
/dkU4garlzBGeLRXJydX9SPdVfaKnGGe4WW0+z3rfbE58fJqnZfK/LflsIV90fsYplIlwCG7Ub/H
ZfCMepFCKvrGh/L7iqUgpACJD/V5hnitMLIA4Ymn/qfkEZ5KJsZ/UHyJwzuXla8zsURADxYL6D/D
xLD0jVmgEFWVLP7xgILdiE+E5hHGpCabZvqkKkp94Jkf0Ayeq5sr/oe27Dq5FDRgH300gsPJ0pfB
7wE7afC9ctQD0pj5IdcTQFqhFabcEALUvV/fSENqk79MGPziYZTlOBxPtLhyQ6k+jb6zF7e5PfZq
xKO9fi9geCjHwvphavxlfgtHpoueCYYDiFFOc8Muy2viu1k7HfhinSEzokm7EcGIl6+UJ5fuxrgu
tJxB/J16y+vkoajRBILHUSN7sSdqCAACzSuhjfAPIpiURY6hj64Y0gct1vdXoUPt9HRhcEpnpYSJ
72Vi+OqAX7/kWUKunQOIjiEIK3XNAT6aQpN5rzY5YWr6UIi/990jh7rwpfm+R6ekIAa5GhYrNPdr
2UORf4EmOL3HvqFxI/PAw+FbOjdMGrlKmC7jUWv/aNlr4u9kOFjzV57vudoRpRVoJQdBzQfhjNZj
Qw4/E6B8RXXZSjkhlNUqPvAr02ApFOcd2NPVc4ZdWco1YrPXe7h6YKO+jv+3/1eeycWV1wkJi6cV
8PonQpC8s8wfD9/Jln9TRhTZEkIQ4ER3WAGjkOAsL/9H5F6ZNWv/vdZ4QaN2n9BXJvKP6bQfzeax
WL3AZ28rrLaSspg0O7cSEoGHtl5MXZx2DuS/cyx81U5GVGwRXjZ0XLnNkOf4LzMO1EHb4CzvjE2a
tZK/JXc5+V0rIJKJssWUIcOaVTrpdauyT+gu50Rf1TddiC/XSep+1inGSt/4zaMSnyVi1QnquQgI
zAsTs/iiYiMsIv4W72ul0PjfYgwyFVWUvj2x3Xednm6BrjdFHmgFrYW+2dxYdCEJutUxsA+bkVja
SRW6gQ0q31byjF6M/iXBtJZ1XfjmXNm+faxFOAYMAQsSm1SoYxJxotdCzV52dCHKnfNfWkqupSSf
F7QJhIOkqKrV05e4dT4yvNsH6rPlCmwBpDdim1Wglmkmk7BBluKAPh4h4PU5h40uO6on32y+6M38
sNn4sRw2A8UWAbNC8Pr5KZZSJ23XRRclWFYVtetlql5vnYqH9dlbXcGOl5BpRS0JeZo5BwbcWBOq
s0Js/oeou9in9yVPK053ZFmWB/CsqM3ojjnxzVyko3G+40JfXF01wSRX7nIFF66/FdeEC769Fyf6
WOByk8XbY1PBWA11pMvQbz/EAPa0cmNYs8M/qnAfCXuV9k3RUFMEzdXYMHzXfmD7+Du+wedQWFbs
cA1d7gUxmr8bt8lX7SVBmHYqyVZemOtRKTiDKg9QL4FaDSPU/SOmLZREn69afg2i/6EgrgMddytb
U8YRgU90qkxukDdQUaFOhGmvyI8IimsCDVh81BiRbsKznD3+8e17WZ1wSJCvivozdRu5J4t4LWn3
kafIpWmUBedgNRCV9QCciR6Q8OXYRvt5v+CgjsqUOI2qexndmT6cznlrW8BtwIDlSambzK8A8fJt
XlD6nmstjSgqtel33VBej9mpOoTly0n0qI1mNHm7C7zbnYD62BTp6KJXXd1J8emHatKr6w1xFgX2
2oqNv11ovplilz/M3G4CKB1DlIC091/iFBuRADgmZo1gxhNbYhj5RN2C20NrBkYDSAG4By6KJULw
C08Q0meu8YsZoAuYBswJ/ofZf+2wKg1nelbbTOewJFm53APEFPSFk7cnMrWBET8xDbicZCy35IHe
EmAEJ8DVBQdWOnnyPMzXlC3aSoHecdacuvxZjLoXvbn520tH/5EmTev1AA8ogn1f6qUgoHnUQTjt
kvECdhrbjaJJUTWVOmcUkWfG6K3/6RrxjrBjQk0bY/Mj+eQek34lBMw9VOYVz+DAnNqrsukEus82
2QHtDeQFKY9AqBYTXYlHDylNFwG+lXyeRxNyMe19rGNHrZNE/4TrrLOZw54XLhMep3d5BT9wqTD1
6vYFWfQPyohXUd9ErG9vvuvqYcR98QyVO8ylBjJ9JTGZlnXrC/bDlO0REf+1a1yTOSaW+KhmQc/g
3WRj3L3z5KZaUMdS6jOy+ydswT/hOmvVSgxn42zy/hH50NOGcBMuTNdSpthXuCmEl+S509BT0NeL
/zbQ/tOwQVyPWiBUxJ9ZBW+0axZAUiMGLyd9yKX36LKEqTJa8YF88ErCpU8Dw6pVl5SLB95I2PB4
GoxW39e6N2pdZjpDXlpDPlorYFH5eyE9LIJWfs3l3VoJObCAbFSwx7fVA/ocd46JxksbRNaLL4QC
pfB+rISQE1kocwJ2Bh3spzku7IdTePGGKv578SwEIbXA84boncGeZTmE2Z9YKZ8DlAQ/xzHUlBsA
L3ksWzieCYI0kuJDdYkdwWQrWwtfFrqooEvBnP1sunfUZYBhY5Oy5GF1y6k2Al1dTF5DNww2UNC7
KDCBWTlVoU7AaUt9HD3TW91mP5B53P9Wtm4WLaRPlV2Y78dYreLf4iNSrfbZOe45h2cFSygyHD/T
Z0+6ZSGe39VV/8VKwLDEBPBDPFyPzP8tyQL8NaWTZkm8KPM/nrsWYZ9K15G0Q1eNNTuB/rxNc8dA
lbVS7dvAwpWg/Bbpxpln2RO42qZbhMSHf6VnZtGZupbH4AyYEZlhjdBLPvRN711jDpsgccXwmy61
1tSqgafFoMcdSCsF2oW0X1Ma5LI0wK8hn1OSTTOlsruOZPUKjes5BrB8prykywcVrv6ibEyg8nJD
ceBb7H6+K13djYJCs6UOcao0G4TLYwVohygVOgIOn1PkMHMIRBFHpSmJOSed3erAAGEYc8LmADLZ
DzWnS6DK+/R4PCykdPKH92T9HBEEM9C7ydieuvAgWGGPkLikzZ9NPlklgVXCoNTWDYK6ZAN9MVKQ
gl3/w8CVL2lbeNK4LWEXSoDoqYHm7ER3sPS34iOJFqHLUdkx1G1zqOherJjjI/SeV4VzFJrjlqYX
SVFDP2a6MK6XMLiPlj2+9x5f/mWwjoUUAaTgtnyxCtYXbCeX0zGpGj4bZABDmcsedy7XHUuyM9nf
jerymO+07mslQDcSrtyNxbx+1Z9o96SQWj/ePQ47iFoUvG9/T8XMHxhUCvlvvFaevHM5yWOI2Rh1
1D5CXi54sJldXrd1ChKdwVEhLIRt0eSQ2j7xXv1TsqUXtVRSfYLOGl5gBBBItlIxOq6VKNt+MM8f
2/T2FMVxeDs/rLh3JmQ6ie0FbOkYygym8yYOrjRuUTJwtpEr/6F3gwp8CRY+e/VvMI2sC8uKGB7F
bHIPzntTvLYAc0AnADqpktqae8BccGPdgSOPVBuhliLZYJxNDQopnqIqO9YjBp7BK8Y2OExMEeIk
ADMwwUcKa45iazP1xk1dEP3jBqacsnjW8dHIb9WvW8srkKACZ674VFxLcxqpaZUBgJtN3j0ud3ks
+JfhTCVZdwNaftFysTsrCr8y5txTyh5ytwzSKNdlgp3U7Xk8G1mkst+5FX3+arlihkFYR8nNqr1T
79tLDTDCMdo6WsXey3x1it3ye9ewuN/sQ+cVhr4bftwDU1I5z5jRX0UVANuCDKf5NzwrKiRg/ugx
9o3ZNKC931qbJ0lBRmFR3w+pi715TTk6kI8Q2JRv7mmHmoMtbxxCKhBzp1p9dG3Vb7nlJPdH0yOY
8B5lTjzWn4dForBhU0btJaNCX9XIoyOtyOs9EOtWfJeDPjLskhUkBBwwyebFFttbOET6+6z+5IAY
Z7t0LCgk1jfpRc5fttKfU7tL9Jzv3+xrUlZjVKtOfPj2S8sGG39P1iRJjRZv09xuwldZDTgAuTS3
V/S9lshEPNWCK4SMS8j2NuFAZ9UC9l3DY2Es5Sae44RVw7663l/p2kO+qt7vlYsCxFSRFSOpslgp
g7yjUqzidGi6gzzyqxaNmh0jFE6WEHNMhfizix719/WyN+5CC7/l0xyyOO+wXJNMJkonIh4DRyTO
tsJM330tm4aYvq0CwIU8AdMoQdQxU+7aEDTBEkbph3DKQVAG5Gkoquy35pYc8NeQX956tfHoUMp5
jageAAD7PYQsxx92AVMrfAZEuGwq6fBwQAd7bOEIh7GclnsH9xodRgyNYb/gDcORD9e3ymxNiX1U
yYbqYaf3T3m7CDklxc197mMOu3rwrAl0hAkQD+HIZU9AfBPNxKQ2l0ns/5QatfBn56lq70EXZnsW
EAKOPO9Tn08Fcfwav1Kkhe5s3HrqIs0Bzml8mdGmO63X3H1L1FnQ8IQ07kHxbmT5nB/2W47cqfrG
BGVPTQVMRcG2zmw5bCAb7osyU5tIpgVaJsrKbIy4tm0q2kUW3zGYuuF72BZVHjI4Je1UwA7gQmSV
gUUP2ZReISObqr58KS9En5Q/dikyje4ZJFcp10sve2UgUkDwhBe+oUY1aDDOZyJTJa665sLV0Rhq
5Gc3tnWwtbOJwCfPryqd69SiELwyQ+u0GpedbU20lM0E93BGR7KXMbb9c57KE7XE9sgYRE88qEN1
FaOvCWMZrdvz0GXACaG4w5csT2bXM81kcBkCcRTlYrfTvl57F1GVu6lKTOFpTxLQJPIao1PbaKcC
285RxkcNMXNaWgI2imQdgj7BOkinPSY5bOjrgARauYjmtXHZRIIIiAyTkXPw39r0B4Qyt29ce8iZ
mOclOs3ZNZOh7JrHHhWctcmhxQnpYw47cDbQnBPxrWerLqnZrf/zy4nx2VCUWorZryMm/MNtuIBK
K2kpGXAOWom3HbWmVmePafdZAf6BodiN51j7g2NEOajvqOrWkhueEmqRGPIu2As6+IRZmIGJVcvB
MK83yGq+34wUHAi3+4uoSYDyM+hymTRBRWqAgjfGIeq+34/btXKLnyhwkpv/eu5iL/mZYdcxlYPI
b6BN37Mtsne5Xia9UY2/t67BwI2vsFEYOXU5ZPOSBgA25y5n07w8FzJ4W/4o/YUxaDtsIj39CCgC
vuXgLkkhIj4IcH/kiKa+usGNDi/SY/UJ8EJV6HW0j6UqASPHCcjGZ4QNhUE4RCyMO97AO8u1Rkez
di8kUCnGuKLMFXq1JkBz0sh0cVJnejR7kkssTa54tr6daz24EpPwI/AIER2R+aW9adBWfsUSkEbW
BYntn16xeePv/xqXCnQyhsHwdmMnBH+Nb+Q+t3yCykZoIJKEEmkldawNF2q0X/D5Nlo5JSd4CVMn
DEhEMCRbjyqR1h18vbGMZCU+zkb76zi99U6OciXVD3s9cwS7xj0l141trwzzXSsCR98M+ty8Ah6v
s/gksdPT4pA40lJsXX6G5raxJLZFYkP1frWdWRfHOmh4tZae2gJeLQ2R01YBqeBQAvvTPHqLo4rc
/N8pLdSnNZ4SEAL2RKZP5usljefo3JJfn2KQ0dbweVwI3XrN3fUT0mDavYDnj5AoqlFhX4c6c9p8
5Um7IpIw4gi0ONjsyjXP/7QVxpXJ9qi7UFp8A4Zc57Pfyy99um79At2wTvhi73aqb428R0tI70jV
CONmXJV0jkaxjEfGvPKgJvhSq+PrPHiqrqPWL0B8sGPCnHDatxFicJqRBbBDHWs+xIfizk3mpHiG
h4+sjJdxRYCeu7ghggFecSLWKsV9NSvMUt9pIgqdHn0Et7DW4SQZ9FYgtaHFQcAJG2w+r5EPvMFp
1MuJMCbXFl7ux+WsF8zGwCZkP2jAq6F6AT5e2lDNVaNnGsZilBoqXYKih3x+xbyxzxmYgHP6bOO8
+nnsz91QRXh49o8UXcEqxCyEkDQJ/6uca1T1VtoDmL6gZa/1a+mVI0dvQAJX8HkfSFPNxZOoS32B
6NSK0keak2u6fR/vmnlFAN6KGZ4m7UWMG2LF1XIQftAlle+MnymJrHje+ujfMbXrWJasYFj5Ikol
1AA35J5MU7EmpoY80Gw4sxIYU/L816BceJx6lEhbda7tR5xfYEXZOgRLalsmVYKRsK4aULlRUPcB
aqugMyrByLueWoTdDnchfoJ2k6HTX+J5zr2LlN5muLLUVk/HbKd/JZrOC7TupqKPtjMGqVoNjqyS
ItlLrIzC48vmnBuMDl9c5F1FzmI9rPRricntNbP4JEaQU6DkhAiAr5YHMxH/6kxr0UWun2l+iXbl
aJvme8BDVkXmIjUtcG3vTAE0LKrf+b71gUeHL+cnnWp0IiGRfNmKfFNMXCt4ZEjNjZo1I5hI75Hs
vS7HEbEsGeKDDG+2u0K2mlz6j4lUC3T0SPDrnLegF8+N5owKDsXuFSUm6jZdgmpIczRG9yPkEoD5
KdbgFzrkL5dOcNU4ymfQOPhE1nxxft5walyzWUaOpXNl4SL3q4fM2X7byA43G0Mozuuvb7uhcYjX
oryOpSieLWFx6vVAL63se5NeKoWF39rVunCfbqOCumlOxo1BM7CFlmrL56yJ5oC7KzCzFkTzEq2O
uYz4z0HO66ZaipOIWij6K3C7JbYphBgnDZPcQi/Kq1VyRtElidpvQ1QZS8mDcDdEDCI2h/verx9h
PjnoyHFfK4xY2jgdf0syc2WEj08/tauoHzRCrVLpcF0BMvvWI2szfiMfPP5RBJyxvRdO8hzPN4Uh
MoGpz7LCyC3vQb19MeVAR142ExCJUdNYN5ycP30fzChXVRZo0SPfzjH9dM7WJsI5qWbJUQVtximQ
fX5aT2gMHX0HDZMDERaSDXQUbLfi8XBLM036rpoAH7jLui3oLpuBN3585r+LZW4Zb7zhFS8lvoJl
rWXgHcvWeS6Z9TZF1xZ2id49L4AZE4+wjuSk7bPRnc6CVyW5grHiOYTLTPkcErcPCLTI8VPiJZle
BOe9lIT6/vJTewWKEdTFrIt9HJj30GoIw34m2rABqPAoBsN7KhlKRww0Tc2jRhZRNubLUZxdf0Du
AdBGPsnYU1d3+vdbc0ixu76JG71sJ6w48fGBb7rEhR97/F3gqyWj6OtEbGM6vO/iCKdspLJE5yMz
lTgCAUF5o+cSK5+43SjLfoBx6QJ8k0v3LuE3o/sRHFihEzSnZvc9GpEUUOtR7DDL7Ox+i39pMYqF
EraFEQr0Bu6G+BonM+bSKv3vGHnnDy5aMtO2oRaokelqeZesXS4Q8k06A+QWN0nMGVruL0rV/VRa
Y0OvxfNl+o5CqBaALvbkDyMU1IlvroDN/iwkC3NC1UUBCbdXfOayVO+QNfSm3Y6laIR20rSGa8UT
SiRtXC5prAiXR3atQIb+SutzATlzn9ZCklUOxhnGI9t2ibRwVXlgEEG2ID0RSjUtklNUWqaSKHAG
+gQVIJCcgTxgRUKE2Hfb+KtHZAnfzEeV8Iz995cEntxsG8LHTmStJkEFWHDfr5ERuBEKdjtb/a0g
WpjxlofCtLoycFgJbVPWzyhzsrILZL+d0lMM+AwDVRXjJravbfs2rW20HXZbflfb7OjUimdpR6ZN
nJmwJRKFEKLhTmGOjaE4VXMlY7/2GkI5Av3sYR9drf2oZghOt/8ivi+MpyeGa2NTmbbrbObWmNm/
cdr6mFLZZgM4DHI/XAytAUBuUV78T7PQLnjGYV3bQJn2WpOmhAViicFgvil5jNDF/Tr8gv2mhvp9
vtBgXBYgJ5gdpf/BPCyz/ZGesvUMN20IbHpZKkfbjnynkpGDcl8u01rpES6/ih52pNZbUMI+t+ug
n8JexOaAHPqB6sMZWW2PZoeky4aX2CLpXpQnum5gKoY7v7lfE01u9GnhkVJ/iCZHnfbfGT57ydNS
gwzR9mLqStR8RZ8EaRvbKlagGJ/dsJCBWLQyW6bHx8Bcl9G7Fn/s1tb/e1N6TR4zQz+CJtOlZRhO
PXSffK6Uo6JsloLg0btcmj8CVPJykk08MYznE/92PiAitkDrrXY0HDYPH7n5PgupG5BTMkAa6yPo
yNaOGRfRg3Bmg2NRtXmGOHlQGrnilx57A0GJKPKT0w9cv0YwpipVSH2fiTXE3hT5NgKDtj9BYcXD
lB4j4JYFJEUJJTGMFjCQ3WgQ8kniOObFhjqbY6O++W/ROEq3TpxTZwtyhisfvPvq4AdgRzyRMo2o
xvhSOhhE0TmgRqDUUfdZ2K5VQfL96MZOT6GbRU4O5Rts54vETaaUawADlyGqqnNdx9cyHGqpl5o9
PKVIxL7UPavZuujDwLHskM28EBhjXAnzyQvz6+9DK/sSXWwfJiIGmMubOq2+iR6+kRK5DWqHFlSA
UZ/fegGwYo+YtB1JcpvDwXNd5p9IIT0UIRvTUQ7vqa7efEv557AdACRlPdMmHVegEln7RJ6uMy89
2LU7InjvQR8VQJ4QYEtTcId/Ti8TfQHMQTdtDsf3/bh6MWdkahgLRJHotpZX3HaJv2uVIvz54wNU
f1m29n4pL9HOMlEhIW/DO2/e1V010EWmd1GBoiZngG8MCdFThvwOuqjvB6N1vyqkkgS9ABYzUIaR
HOU6ZJFhSxxZ2Y+Jh82Bh0I1l0CzmGQj5lXddofbe7tdpz6t/SEwwj5jaB502icSpS3y+YFjjA4j
o9Ytswfpx0sX7gFKkmNElM3C9d6HNjGZra/N4pSAyZ2GutgtbaH1Ki8DwGYkU2uRpYF+tEh67tzD
lKLHc703Wy8EfqMWd41p08SfmtqoaQ1oPjUsQgnpBY5ueNoSDhrxUQcWjj4JGM7z0lX7IRyyZu0I
WFYoeVKiyNaOCFWvbzKZt9cFzuATemhV2Cdr7KzviHBzrnmc18PIlh7n1mfGxGdkeyKwWQpIUaO6
Q07+k/oh+gb/a2zCNGZaNx/PCL84eOjMwrF44yMitxf9Z2eW6bhO8SKx7dv7B0deSm7EHOcst6eY
IzLrMgNeWZVGUnwSeYD4VHymH2TsuL12tniGlEmMArdO0T9ST3kdjBalKgxlLh1taw0LWNqftro9
WvrtOhTA+SsKC08ZGl1z+Q4luZgrYRNyAj8oBxi1ykL0U0t2xiUXd3+5yamFjhG2JYI3fMiPqjPz
os8C9taOiGQ7t/x0qyI0MN4IwV8GTJNRreb2nB3xdRDxaPhzeXjRvTLtj+nFp0EN3b+uk8L8U7s7
LyxxeA8+bz7tY1jHqS6zFO3VDdof4awbv5TWsPjygeGYaXmQ0Rt9bp54SGBIZce4ZDJzJ52ZoYNq
Y/EvwAqigdmBh6eBH2xHab2JH14p4FavqiAGNfh6cW5dYpWQocVlLlzWh1y1Y31zPPfmW8Yu/OOE
OBT87GDbEd8Y4c9hQPQ5lgGtHNaQpr0zWa+ffIBsH9FE0CyvsuzSeMyhFtKuOeDqXiRjvRy+EN+v
5yaWv5gcXsOK71JEdKfOfZt66Zk+XvBkJZAS8tMiops4HU+4HYaXhPh0dk7TDUDFzm4XUPiRPauT
qKpXvmSd0DYzTaEpR52ihpjqLylMehGBTFPtTe+eoEcRVSTwJGpbyqrsWJVY7JgPn49duwLSH9Bw
C3A82bWZnEzjd+BVxD+M0VoMSgCHYYF9FedRUGWHXWNi68mldOmrjy6hZAPDjUZNnguc4uJQYb+b
asp3zmEbpFsS41EkDr9TRf/trpIkMxnFedZdfIjLh4HechzH/Dq/i4MnIWYnlxq8joHBsywWSBrA
XTJ2VHliUzEZV1J7mLr/hU8JauspWYTEm8QWXC1vljFkD8n5xsfBJxEkTQ2NM1reH+kSOzGVNd35
frQXUIuBIGRIPrVTziK4Lh909UU+e9iHQ0aBeL/MVc6vMmVTf9WlwJOO7RmcxF6deTNzMtmP3god
7LBXj04Dk8W1bi/qacyOVJjSmGhNMe9fvdp6ED+3VBlx0lQdDomQGnnyOkp48NWOP9waWMKvUkT6
fn81vIMqA1BMtALjaP/eonhEnn2B4ioEYa+4oYxlG7RzOm93GIyCf9pPOlivDm0GWXcdf0tU95Cv
dF79M/7Ci9gnW75CkaBbJej8PrWOrY9e1OtKn/8BngjefGxXfGI6q/Mz41/31GNvIXQkRn1iTbgJ
Wr47By6BwrTevAX925dfDfUq0PyBlgonryBZcvu7U351tbzHSgizQpx+qBceI8uQieMN0gjNXg1m
yaYV7UVMhcr+a1mAW/hlrZxJXdBnYTu1O2VMqcysFJrmIz9GTM8EgLQRRo5c4GzFWR50S1uDdEzY
BfLURjFc8YRJqAr7FiwxN5mWZ+5uQP2DZb5YuBb62WJIOi42AXCDHc+z+aFM4qCfgC1meEargx/b
BCP9dIAQ0Im1EaIv6YHBLtNSqMDU4uHCTB2RyV2yM2st+DkPpxBpeTFNWEQqpT3JIF+QfuRPE0ta
cmuxWJYm9US+SCXuh/q3wzQ34vS3imq1N+Xb01v9xRzbIzZV0leNVJbzQQ7/F1TSZVzY00vQLxVA
K6dsimnscyWMGohBicS/vhFG/OvfzHGA2Rtq9iYUQy3LGOqBnb1eIZj7JEeXbhuKYITTDMHHfdIe
XZKacOqbvl/1kDUnXdb+40Zocy+wMnh+7xGwD0Ir/Vp9gmOj2UQvvio9+5DaMu0KcA1kiiyJxNwd
Mmu9respPd06ehOlRRjTfS3WN7GhcKQ7ST53caOsmyr8gJvV0jFm3JkA6uPrn6PoXXkeuAd4EGNN
GW5/UwagqbaDTFSf+JwLXOlNRnAz8AXWj0lI1AxhKSZka6vJ2C+7k3BdmVrvByKhY4kKxGPg2/6v
wRroUZsJ3+/HKx/aYyug7NzFqht56NEA5zMZ+qRwuG0vfAD0GHRhWdM3x2RlIthbOmY0P3gbjCx+
L6n6AA4pjrvg9bJia2FqbUlIeUGfOS66eUULlYBYPM7uuo/GZRd0JJYYgaKZ5pdkmzluxCTOYxgp
awxvfWHj49E4PWBJfY5f10ThTTD3EipzGPaXdrD8EsKqjffk1sFL9iH3E9nVxD1+ZfaygfLux/fX
k2DRDfy9CGr96R5zrmBURntc/+WsUTAc1q0JgTrUc+N1J7QaFKrT8Ef+0ZXr/JdVG+qbEAA6QwAg
ycgxhliehjp15WI4+v75HTEhcrN9qVLucJlkJYvqYH1cHGuRomAEnkq2Z07Fsq6bAtn3oCWF8uAk
0T5h78OEgCfSjSR6lm1Gxzb9Qn1AHerTntl2Aaa7BPBXIg1TJxWPciS/A7xfjqtrvBCJ7voadp0K
V7xVO/pvnYhsoFnjQ23cqWodx0qV3R0XFOVbbX5vIafkJGxLEgT0uorp7rEJxtoDCqvpWFA6xXtA
DkKqdtGsnoyHsX9KcS7yNFFmpCRrZ5GL+x0e4R4SiwVj5ufJVlVUFZWaFWO5pVdpyujjf3FJb8tJ
vFgJsJ7stCLjYs81JUpZb6U+btRCFgIKJjgzbIk8+8bTKfM6r1RVvrNyAUg+dJ1y6IyYfOFy2r53
s6NjLwIfAKbnV8zFdozsRoosxUF65pf723EtJJL2nan5HOxJtSWlLteTAcfW7rUGlbcdOkoUhKcR
gdKpSi+f0Q7zmP5Ks0JCh8GLurRZiqorvTNdoVl/5by2geFgXgm/qWPkjQIuDVcSJpImekbTKU/P
ChTug+UUOqLJq8FHmcwVXtoDhwglkJtWvBEOWRJQRRkhyyURGpHtvIkkIRSYly2XPEBQ3FjQIG8W
Vu0/7mOu7LsiDr3j+woU41cAJ0DlJsclTS9lPMWbwS11a47AX9P9e9ZNdlO2C4pt6ZnLet2+CxWM
Oi1DtjqXr57yEcbp+FwyEvPo4MOIWkmXaircBiTrhwXAD272h+p0CiDrNE3mTSdeMurgxTiPEXrp
r7QD8A8/np9MwGFxcnFuZgF/npGk8JLwbrvORR5QeC+iVBP64NViO/Enj+GcMrXfPYCCCArl684t
GrAmEFHVllaNnZpYbkCoc1Zoobwd9VAS2xyya+KPwRdyXVepw4SrPC0PGcO8tEPhw+H8gg1fwoH/
8UYwe5zPcEodFlWDedbuPkQsVWwmFQBy0T44sdKZJNOcQkws60QqThm+Di7gxn6giQvRTPdGbRvr
OIh2k5ttS41p4TGQ9F7oay4rnX3KNJI2JsoMRCy3rMmC7+1CSxSdN4WnqQFlFb71BQqIlmq4a1s5
bKU3cA+WEJPWY6cM01uPbkuzubmdPxtZpAmaYY5bALKmE25qmLwEl9TuCtCDYjpLaRT8arSu2g6n
D3UrUWcMBpJf94L359gRxELDR2kPLSsHtNbOLmZuwHBIaZbgl3w3rRdxrci+SSwTZh3TFY5DLy3h
eCMsABrqDl8MOKWZzeU1Drpwv0kGVTV/EgL6IlQgtyaaYAyTRoOY+vqUVAo53AwGfl/SB0bcRkqo
hX+ABoKl7sd8yJZBA2JrK51ndqHBgL/VcZDqpuf8r2EE+jmJvDiRC53QWE12Hq2OG5qIyRA4qhZf
XcMTbsI0h2Ks+/CaUKu6L1jQOVRsNTTiOSgF6oKWr7HsXwjIV7iUVlANkhgGLIBKubrkFd8gc8aX
+xqI2aVqf3PFwY7lcglbTupL2oAufGbFE/r3ryVhUddAipEVZHH4mXyuE5JoOdoHHCD0y7Tut7IE
lEZy8hebrYwqt3r+DTTQEymnHEfxqBk8Ix+0IMOz7gyqHJp5W6eb57DesxL5FdTaz67cIsVQC6aq
o+QmEBRiN53hzfAblAN7BrKzXpQz4KpOsRxPoRvUpFPkkmpJkOr0GkcC8pPa8CJNBrXTfzI+zHLV
LENFYq5EZJ7VkShvOWG0cG9iTTc/OTqh3BLpBes/AapQ8r43v60EspMSJr6e+DjdxtR+QaaGgPbs
kxs8VYE8AaimnOqCD9ZvuhMyOtf+eKDw5H4mor7ksiIw5/xVq7c4Umz36O4udPwcfKsdMc1aJB35
N2VtYR49kKsbN1ZuABoMZi0Zqmbvm6jKFzsCjcC4l50tkFJQjou71VFYUIy3nEE01ifErAh5KGnU
7tEnQ0IKzpvimAjCVvwm1xkGqOGlbeupuTVDZ3cCL8ofM9tqg7xVprsL7NmIXCM/+mmKbsqCrIQW
Ox+ju8eHLxvV+QFS7VJmY6+AIrvJgB1DzOqso36/doR+AWwyXfYhdb6rH94Zkkmo+RVEfePXyTxO
ERBHkKzvH1TipnDiRpNzTIpoD0J1UONBuh97OECW7eVelRjPrTwXWWTBF/rO8LfmOHK3uUgWJCBR
fK9MSaDnPwXD8XCGxiyJ7RTqPM54Rr1fUtRXn8T7w0XWGFXS/zDC13qW0sUrWffV9dgkPpxe5a2U
6x5KUPQ0gt9YTGHr0GkwBJAA8pRulsqgqTZqbXdXhIeU9wFmkLEe1RBRYDle/fcs0sYa46Z/3e4L
lnxynm6OmDuZMBcPYKrp3jrMUG3VYqwOKzhTBji8ufaI/3vsnNZnlCJL/T7hTy2uIFNzRqdDx5xI
xn3/eh+uLpdSs9Xtyl/d3HLbYkO3Q88VPJH6JybA9zbI40MOzm4Oty/C6s29vb/HdnCFuS/IwZ/c
5j2jtYbGNxPUG5mkb8Ey56eh1EiWTs8oJ+hg6hdxhr+/pnZ+2vdmGfmHyLsk/wRsaFjyJFowEXqS
mvry6SKbbFtaB52qm0NVln9XU1ASns2HQXjgsqJLn0tnPssu78KDNwmFQpYG2N84epwweonISNPJ
mlW/v8Xdy1ubBThKnjDXIf2zlwJSZzn9EE2VMueA11cjzlrvtC/zbvT/3cJqFIDJ6hEkLV5PYAVL
9iPWUv2RhPFfvMn/zxpVIuJ0+0CkUSZcs0cLsbJoDmoDqnyMG88Vh/9l288G8wK7xuVLs6oMKM+b
nz+9jEWxiI/Mubt594S5qC7CiaAYfstnteYkjT8BzLTGuil98dNGFv1o31TODWiuAIvh6uOpM00j
53U7EZTVNuVn3qOXUZ10dUrsc+pZtjfu6OGju2XVQ5ClTR1d+tBdTvT5EC9h1JDjRKyrt1P4oNn2
+12IgSOBrgC9hyRxJh6sUvr3N8b0Tjd+z4QCr3CIDOQfeEcYv7wk6GirsHOXs8UwUWc5nPze8FdL
g239r5sZ33tuc32Vooh1KygTFUMds5qaZL0mGhHClG6E4g5k12kqQaAz3P6v1QoAFGsbrVtFLPFz
EqR/EbSYjuhIgTaf8Ay2JLpcdOF5W7LgHBsuw7yNAeRkqX5EAayESW1EFukgOUn2i6FVLzeQAtUf
PSe1ozI2Mx+GERt7zyQQun3QpKC6AVoF1zpsYBQ1cGKm+CYmTxxNrWbIne66B4waU1V74QXlEG+K
hZ3HNABrqKk5qNOLCb6P59+Lll03cXwNxTmruqAbp3JyRTol7aKyG1Okis9njlnzzfrkI18lqCMh
2wPI7wmLyK2PYuQnWmkVDu7XYVjs2CGG7JTSPI1YRVvu2xJQ3KLh4O8QRBnYNRKIqQPww0MgY4sE
sdjsMGZyfZuco08MPJPsSSL4iygTkATg13p9T6p4/BQBJWmdHgaH0yr4furuDfh/bbaNpXpoI7Ne
3uZJ+xykMZwi/2Grx3ANFb3bjdfc6xzUOOypapKf37gm7dXisktNUmsBsoirMIsrYBKQKOH2IPRG
43wAta/DlLL/bPYGzRlnJghIRuRNwSmpekkao8lozmlEFlEfvtJG76F90QOSPcp7DdMY91C4yjTo
vkysFApHWXXe4VL2Yza6DQtVWuYVxwVY+2MExUSwx9uetJnq+o0MWVyJ+9zr2YGo4YMBwg7NsNqy
bY2DoUppkpSswJPRLdUO0/idu3xJvInpem45kKkC+q/JvXpzzlqrdmUPZUU1To9vfodDHGERIin2
zNWeZauulKrShfTt6hPq8+PvfDUJ3a15dIbb35BxuiFxW5Xga5S/ZB0kuvOdayvGRo5NiLBHQNAn
BU6MCoMG3fu4JOCIf/8t1LniFngEdAjcZO3SF4iOAJKpiBekcQeu9QiYvjkV/GbG4qBNKcGNqCnh
yCkuk012SPM56nWnkfJWngkKwGYH4lUImMSGkzwXD5/lHoG2i8mNeUpf1CJkoEat7t3PxLR0hjJG
aCIGEgiQJYni9A3YwMnnfMRW86+GUA4innFNh1u8KMOrtMZ4ucrM1nIdiM/AquBF/DeYTg1BC5am
EQd6Vcl6Fzwuqlk345q3Bzuf0pxKDPRFs+ZuYhQmk/PlNXFxOlXw7DOWsO/DtxhUxAYXnqjbTWiU
TUcBRXy7yymUkHvurRL3rMyr4K2bmqeF1wZvevPY3sa8uR5c0WljGzp+jWHBBk0Q9j8xYIWlpViA
lC997B+0ScX6zbgC8q+hDxFSqi37MF6h+YssZ2GUD62jJBxtBEUUxvwV/EupinWVRa22BhkTuZul
6lvRuNVucAAZ5LYOz+xvuHqEI0uCHdsZwRhyoGMsjX0nrIu1OZ+VSgfB8El6P+FO/nykUFF9LsCx
0AkxLVH/poEKB7vnzpwnDf7FH0/P7sLuIdUzUSDOyYHMU/ejhaTsu9rXiOEcVAV3T13RjzfIug4v
LLiybbucZ9nJCjt6Swu0YsUmd5V3Am+dScekNwvGGDl9HycTkHc+03u5Liis81oeI2IafDEU1Agq
roIHpOwcpJo/I/P8Pf++PqEPsz/a/68LvlymrK+fewbAInI6JkD3IfjUHB72BjbAn25L7qXT/TEI
wRoVJXdsZT94QYc3FNDem8+jwoevD/5I6cfsKN7dkEsSI3r+UfOc8D33NVpPCfy3uaIOrVlp6NAq
QibjPqZcDUO+FU7z9HdZm7u7xCSBdKAoqTWbywa/x6xDEnhK/UYafyi5okWMHz9McrghcqnBhX2x
8eS7RbRVejZP8qmeqIL3kvqCp6Id8c2fA+xi1O4ZzfQw/p8KqC/IlUH+YggBtdcuqDHexRl8gt+5
UIEZUoYWa/pm0rX1AzgBO9jmpvk5CO0plo4FjLNPOjj3Vg16qAmnaVS9eZWVeHzeiHXyEyN4QuWM
Xz2rLP+auLNIGFIKQt7T7or9urVTWfuZrD+R4w87q0FKEaf+zMJ0dXx0HT2kvyXPKRqIBfx3mjwg
foc2fA+4S3UJFkoi2i3TK8UHIhWVSI5wXf/hJt9nFnPf/BstAKAHUF5tkxmdwGvFvdcvpApHEkrw
IPb9iO0OYlshtzSqEXgXBksuoNdkNHHj5c9xmPiMRJxuzSJlFcSKpybsXAvcSoxGn5ZFRlaVadg/
UqsOen8zVIPuwIUDn5OcQSmMJngDUy56O5LSxcpU1+b6Xa5nb68GguzVbFi/otkPxRbHD75IfTFr
nmNRMS1Ij0ad1g9KIvQoTwtxzcfjqdLAGPkXq4o8sis8j7nUA1tojjKhrgCBwY8TYUAC63F3gUYB
xY4fo4Obx7oWpBsLYYuXhkgSYoOYH/9ShTwUeZLUK2dM/6f3WKfVXTjbFLNKExy5Sx8QCLmOzwgx
qAca2koG/O5dhQK0rj9DdHjeazVk2AEnhz2w0hiX+1rWBwIUvfPXG4EoVBl5LVRYkcrimXfwmjeq
ffWicJYJefKN4lRmSe46aK64gRB1OfADGtjVM22zmel+80qmO+L60JH1D8HO73+apmgXXCm6alH1
s03PKLxmamcEJva8pg9grmHrMZOjxyvJTE9UOtgSZVfGN9O1h1JPyIr6WDQOGP5MIR1glW1vk9Xu
Uum3fcMsLfcLefOJtJY5KZwbYHWw4zJNa1BLT6Hau2DwnAINuZGS2dkT477BUVbvkf58PhniX/7X
DEKCB0SYLwSHQpOLSGcwhHhsERPLSm3JVB/VV375EciFI1UCa5g2IzK6jlgi3rp7X3DP712h3HqK
2+iExPdJqZ1734UI12zoXvVDOdB5N1kmC97lr/zXRUsbQXK+DEcDwu88FjyGBhEUThCq58ORj+k1
xIxUgp81SSq5rIyNijQhagbBLVhWoDteXDK1Kke129kWdPnP18wx6+zDIeLFjrGTPDBFUrrWR5Xb
7QTuYn4OOo2Pezs+mEl7VKb+FTS5nsEYAEMvohf9luVSE20ElwR9GojodwyNs/x0z6fIUgIcEPrJ
r7wWnFLk4GRYUyfe1zud+CTNcNbn+CZRG4BiUslbTA30q4BK5sZaUOoNrRnsIxcSWJyZv5KyaSil
wM8JKrxeBo7XLsdSq7T1eaxxoLKewSrR1USIhkXAT9AYs9QIgBRjURRCt761tKNI5xkVuXHVBIt9
Bd+NEN1vpuH/sDEDHFPbE2hHCK2+qETkcbzUq6QOAqFa+A+8ZBNcNi7DwY9yjCMmC5Yud4ve4z4D
h9WVvZx2Fv2790+e/8pQySez3eqeKQN0qKYjdSdGvpDDitJ061flAl9+z58u+1xMvhf0ATCYtb5d
3XIeMd2MrZyQjtPM63aGyXZEV9WDS8y9bSXgYQEu9qvzVm3E0aVLqKIa6Zp+Qyo8DR7mA1b6puSM
gClrcN7yxHmj+PEvBzoE8TuWDs3j0vKnaUDdE5BTyRuPfe5EPTZ++3o80gNwq2twYgFf6IsqA7Gi
EvGs4lUSmmUBkCvqoCl164AeCp9h+tpOxNMPjSN0r7H60vEhfYDVANPVsj/449UO5Q9k9hF7vBlr
xTPsbkKBiHTNLM1qibtuoLy7n2SVuwIdbzm8x0U6a44y3UTmGRMEJ4xyygEeqUGqUMUK+YvWDV/3
JonDsaq58LfQda9OSV5hWh2F0lNzuBKHUMKeFNQpyPfZHA3kBkinKEySKFHMDD0sz/67hgVaBfns
s9cXV0RGFntDHmNgIcmeH4CVgABFgTvoOtyJDvJd4DqpM7QfPMmnjKGjd7VgPV3WE9V6K+6eEbR6
zuphoZH0P0MGr787PWeJD8BL3ZoNZvVaoK6JTAO3vHwfRmmKNrIVchUCUTwWMvK9ESxz0BSELob1
tXrppQfFy6Mx+hpfS4kIQbhH82gATmEwCwcVqrA8AUXVZg6zbv6FopyJeYfeouCwekW0LtLN6GjK
pPuZVNvPHyuT3YQCKZI06/NZymP2qkOPJR8vp/g6qoPwVsje3zHRAXggDeL87yWZ8zTA6vZtgKD0
I0YRYJ3ZtgcNyDDAHwTkHoDK3kAUH7jEox0EWQvl/0tuiOf6aeDjMCYWO+bhjYIgwJ1hhZW+iFvq
0MrJ+jxXrZKn4UbiTFowAKpuYWXbDGAJXrU5VKOMI1BcC81xIlZ2vFufr6B+Z0K2/5wfSaGqmVys
yVwFLFB90rFh0yorcV+hnnOCDFFgdEAW6XfOdrtvogjdf23KPaoPVmE+sAJHAsrLqOecMxZR5YwH
IUsLw5WsF4js0SFn4f3xg8OHuWAr8/MyJma3mWrSEOcVcUYKg3f/6NbERGX+iiTPL6Uq2JyxPAuq
0r7m++gSr7dzAnCNbs2McVgOC2XZOXGo24qYMsgAtlVJ192Mm6TCiodKrbcAfu25NlwqXZBRwEqy
WFTShfi+b6p5XO/4MObGH+ytB/JaTGFoUHgJv9SSG+iV4g3CyH17aQNXSKWSFbJLYh9pMAw977gE
vO1umkR/NYY2uI6tSOM0IwA8ituMUEFex6wuCbuLXyeXlO/ix7T1/N/aznUtkRSvaeS0d2/XT4f5
qRTXStVFuF+BeI5bXLZaPN7Fh8BJfVoQm8xGjOERPmbQXblNWYQg8qvMCGuoDVH7qA/BcBmxvqUk
dkIKQDcczP6FD8ZLpME/k4Vqd4JUXSY+wxx2vvuDyioREoVZ77VjHq1OZ+nlOBG+xeDOgqZ7W5FD
9WE9rBQCHHDLy+VDXyXo69QA84nCiBQjBVumS8NT4cCRanWbvVzqFg42/u3monCXFogX4yeyhPVb
EPDs3z9c5e0plSOmD3bRT3fZwZf5nQc+j0VDUyn7yu1uYW+y27eUkKE+nwflA7xom08Dfq5PBjdN
XeN3ZFQWMh/kmHm9YwULML0I2NZBxdDaI9eEOg+UP+UKXj3K5RFco6o8+ytAPhwsFLYMR7IqMhAm
RXv0p4XV248oZZfb4yXzfrp2qwJ2/QtB/EJ5+pmGvfp/orfp/l9hvr0xHIvTBvHOAaoN2+0+iXMs
saFAckkel0WGYcLTIXeeHOearGr8dxEXWVICK9Cisj54YMaZFgDQnSqf/v4Q8qoJDKLOv40sM26X
zGxNxQIC3Rxpcnp7DCi9UYr5QHtA2ytbZslhO119v/txmsYrHiPzpbrjhSfuHy0xYskDuAC8a9hO
40qE2aMM1eDBD89uCQaww9U1qJ0fFOJV/s2E4DFuSx0KOPe7zPw2Df2P557ZdywhzHcWiudbSzHR
iu7yH236NccxLzjk6mYvt9zljc/9xgJibGeg81R23OcnyUaf12Y3QcK9XBA/MoU8nc+Vwir0574q
EYSVAqJJW1zRgvFwiN91IshTkKZwFtWb+/a3Jareh0MrkwyQo5sOSKa/5FMCrdP6I7XLdlvljoD5
7ldRT1uKmsBBqi463gfwgYryh3mdEjqt6ctKdAoeWCvoubExMncTUSdS1JXricPOh1nD5lzdj6Lh
eAiN9vjxCMC1rZdoEmzv+SI8dA7+KFfE3Am9/FqPnO6sG/NNj9Bv3wS8IkP850HRyuojKp0C8QTN
6T/n34+leC28Vj6iyadP+El2TIdrFvbKdKkR5hFwreHEb6XT1bnmMqB/MBq9DNU0M31ent+lHwok
lHLhRjwTpdvONjhmlGxg84n+NgomSFr1eroQbFL37yxyFHPKAZiX8WLpMuO/+VnaSA4inGKkREgU
VUn8zDBgF8TsjulpMEv0oj+SYrSZrWpK06lpEri4lZSYWzeUEUYJjiTuNpvHd7ZiYjnszs2HAIBt
1+yDtKsoYMSYhAszUMBwLEoZAUK2uWxtSi61BVhUSxLTaawegam6jmgNmMnhcVurWFcQFZG1CQ1R
PsoyA9q7EDfI1/Nb99Ryw0ZVNTqHqlUdne9y4nhzdWWO1bRNKJfsvW1EfYdkpZ6/fuLq0Qs+aUtA
tX1/6KMI+4BEwrB0pdHF1PIa6ybmHB8GLsg4c/p40uTUAc7d7NeJ5BYPo27DzpnOuPpO6moi5zLD
/vGoJTr+enLqCkvI1ai/9B5gJ3ODCHiEMG06JS5MPEokEq1rhC6fLJ4EynXZf9oKgZ2xdzn0aoUH
QXs8m+Y/GES9WG5XOTvATQ7Befzj3n8cE1B6h86emRa3b8CQEF6Jq/Uv4zvMSAK8+87k/zZ7239p
rjo81VJ3arpb45AwtsRnEnkoV/urL/clkKcJs5W9A+/XJSUh27KA39RHy6rrGwyB4DGRGS8TmtLM
tVtcbHyQm1eEUL+dNEt6vJtJgRa+bxHJffJ3gZjBwp771C6x9wte8gYP46taAGOkjO91q4acJSDc
Zy/HVD9nl5Ma/v6TYcaDUjCobn2ptj34ZwxAwZnxbU2h3dqNYDIs0s5Mw+OH/buDD/J7r2rY6Ivo
FP4z1BkxcAQ6hK7x3959zkoTMyCLI+86VFFrtDLYARuV+LwbjGL9hr8XUo06gXvx1ZS40wbpbl4E
AvSJlvBwlPFmQ6vrn3iC2Jlc7yhkTIGX1aV9RSQq2LUepLL/wg5TBhI+tMO+cCpILsk8tHJVfbxc
zK+DJ/LfJWI5sfY+diCSVmqw1jeU+0X8mzrwpnnEhRgnJvI4Cj+FPklpzUrtBOwATu07LRTkAy/0
BsZKL5IWlsUuFemXJt1vdPahcbvLmLW2RlMX3HNKnWGPa5+Xk0/wV6OeQqFZ96uo/jcagEYTBIuA
ySJDiAANiocmgENVWg1Jcct6Y/PO2DqScRQb4dUrqaqo5m0M76XH36q5UxoS/3ee5z5XrfNx65UI
9fJW7xPr/RMo/5cJ+KuEqJ1/9ubsD1xhG7IcRmfUyl4BR2kpihN2Pr/zCgaoHBdV2dvEfKApJMis
lI7LVxsb9iAKpP8/72VC2pPGbc+6fU6//3yOZoOw8fRMELQcKApC4XJHd9XvhqzX7Zj3bSy3iTj+
JdG8WEM/biP+wz8t9Fm79EGan1uGiXVhr3RRHDo0ngaEg944X0c/IWrGIGTLRa0xCA3QdVO24sTm
n7k/sRwHxFFk0DZnjQFCSthX0zMm5bzpoDMbq0xzW7Vfsw6hC2GDS3KcGpV6ZPiwvl2PRvPq9ezh
AV5l0DF/tLZOPk1V92xLqVrtfGuofkMwteRqC3YdAZl0Vi8Mbq9k3R10rd7G2wFihdAOqq5prsh+
j18B/RyNdlLNIGEUKjVvivcCFcwv6fLKJC/py4R8CzcECkf8TrMcfl3C0m/Z7V2hdGPJ7gNPSKGf
kBHz3PxkLJEfQlvur68ACu+zqyeptQ09zxQQXsU6GLulvnnexUAHrpFo62v9gc1P5iVNCQT8AuW3
zmSHPjNXzbFGu/qpY8zUWezQV/xY7YqSM/2wns/TmuXCJpUdxohANexnwnesWnRayWqeb1GkEpx1
NzY5MsKuZEDJyEp0/Z5B1PlstMz4xCeoA5GJgk0JK9JbmHgE/Q4w5gHzG3/xHw527WbAKMyxZDEh
nnUXsGLk9VlyOHvDQl+TYa7dkChu2hbb5Yqq/SvcEk1RB9ppynhQ6fr2n/Y/ubFGkXN3RYVHzEX8
EgDQ2LVjxEgAEwg8aHa1K+TnxgbtfU8r5kJgbESsch2K4OB/wogsn6y1ZClRSgyRlX2JFZMRT9cG
fiCeWwCEfiJjoPmqPnX4E1rvsT2FhY2qFIlc1+ITc4LkS2tcPaB2vDU7G2XvCLTJtGZ417ZHtd1X
ft+3FjPKfWns1h6bPUuRt9SpvkACfoIeTfjgxVjSwKYM2OOGHZlXLu2vNJ0SB62xYhxALl22aO6Z
EIBx7d5tdMHfBcz3MihUKm4DwMDvtVDEwfL8iRv2DbTcDLedas38xEJQ7gmsKIhfuYHoNY3YK9XF
I6zalEoXjhuncAfhV5bqCxMTzY39w+SAytZZzLvM/I9Q4EKP9+q5kE397aJtUOb2ckY+84/WHfCP
Qe0PD6vdrEaUfIGGsVswvFoyXJsnfDJJ4a5smREdnsy/SGoFjbs6n4dQqmvpyf96eCRd2ZIsTN+0
APErAyAvbmiegxWx9auAUNHVbd2xmdnNDJz1LPSJndX2g/F7VJwpyC1D+6cdCLP1KOYdfmRy81vH
MN9bSwGt+0p+PY/FpDi+yLHzdoCQhsbI77NbMcHOg+JO/qSNkRu1Ahicy09KmtgG1ca3CKER8xX2
yo2Hxi7BpIsDf3sGcQUm7usG2rtM45Tg45tZzzN3X7CTpgQjKQYQ55eKdD/Hjg7CNqrMNe5FP4dM
cwHVJDB/ZQUiVj4S5G2yTzETFQmb1XeoCWOwF1/7ps/X8cU4DC8XQ7odAazrOVtQXbgmvuOhEZqG
XC1SE5E/kseO7nDhed2VsEcFmtGqpc2PH2FyBEyPYxHLhIctWklwpROwZCsLlr1TJ+kDdDp41869
o++bGxQZW2GwsNjHuTZgBQr7VwT2fQyZmYvTMF2yNn/AzKz8/lCeibXmFRnwAteYJbuFXgogugua
MPKIM8mSlkaxYwwIcl2DptI57M0FooK1rT3BZKXqw1VJaK9QnFJASgeVTe3xeiA13jUQVz4Ld8IH
PY/uf1VqiCRePsHGa7dWZuMXlCqi27fvOJGHnwWuSM/yfs/Dy85gFlgReLMGbuK/FvHMPMwO5b1v
6a40vjH2Z6m28mw3wqVDnzftU+iMXOHXAVQ6GyKO3X43NdaSobI9HWyF9koQzKfejtjcA1v1vugp
jjo8mWy262SYTXAYHpibnNFCk8wsn/gHTDsoTJUZLl2Y1c9g/AZcNy1jdYdLKrTueV1OyMHaBEfl
DmSoVdRJWuJKobj6wl29+DYiWt1SSHf3EUrX7e+6V4bJUQ/nppISxJbGZRRECMTbBRoYoFjIxjs8
b4oU/eKLt1XKEbUNJa7uYwEB1j9TM1K3RLc1Ct+StPLjPaerMcJrtHGqs85LdCbmRUVqSBJ0VJy0
JW/Lum9RBjY3goztgr10apqkNdnLytt3aqcTgwnK0mErjl4cbFc+plxEevIHt6LuRkuidjtNpdnW
cJeIUbZKkWYiPk10+d8yT9Xrd2PKUAA/KpEHon9N6N/Y8UXp4h/B4W307DlBhAVmOvaa78+erG9u
Vbm2+TAneBGljT48gDBvHAMh0wxBkKWqjtnVhygRVXCqDu1Yw8CsaLZ4mrzCJ3yVmRxViJ6O1ZZl
7sO6Gk2u+n4SGEPJT41KVU6ZTp972PHVi7HQttUYMu8hm/NJgHMGB+c1iSPOmSv+75iD9VtncVe+
5pR380cGJUYD75a2dckMVfSkxizorig4iBTPW23uOk1j8j9gP0BDJQs7UcOdOQchUWJYNaOskp38
0WxpbYmYDq3X7EP17yx14ait347N9UBvuxlUAlR7nfxOZf2lQhszGd6QSjMG7vCppcQNzq4jABu/
7sFMxpRdYAXJSnTFpx2FRYU7pG5eUIC8YABLeVQxDVLIcMYtfmRROmump12nb89g218p9Ljmep+A
6gbUuz+e1T0a/l1GWLF58Pwop3wCFUklTDaF4Bwl8sdzVQQgeLTGmNae/ztlbGd2WBuVgCI88slC
0MVH4+O5wdZTUouw/aS3f4GJ1+WcTMjJHf5hSlky68MQstzo/LiiC6mKBiZdlIoPaYJ430LU+PmU
lRZHxHuHQJYBYQa+5v2udfuRa6LdMm2tbTVQAI3jx4Sga9vXh5BynMCkjY6wl7w4tRl7lgER6iGV
mjw9zK/ToKgGeQXtlFynxEeCRgLGWguQuLgS+0SXFq/5bcH7XcEF+MALqu6KWBfdYQmNtLPEQlbw
s6YzS3YxeBlxMoj9KsALlxtn+WNvHEaImDThMHiN7/EgZheL/lIQ+Mf0mEVxvZHs8Tqk/kj4WvjU
VDXgYMSTZMaDeLDNg/+jAN9SReVxyv/eEeUObBf663Zeahgjtb+AHAXX38d7uEE7lDgnqQG0OzFE
xFOm2ShXUnLuJODtAQ/5DsNA6QzW9Q0Wmphjb0EmSgeORt5y3XjWVOl5ASsGNeA05xN3p3r/M4v3
28pvTxkPFDu5+VACK8LIfBZ9IgTr/xkwKpdm6U/fjXQYoIaKYaFgwwdjGk3GUPZtspt9vBFgCDO5
Gka5R1WzX5EAgKELittB6w57Hao1Ldh24DclgEg2JtJWeq8KCPwdiLpb3RAT/jjRt/nyQM7JlHY2
DlEAxxltolupJhWf9PG5ISERov9NR1swzBONhLiVR/BVgup4qylqUDzPFolox7YkBENV6Vzkhfai
80OmRFiGa9xHmftp5IggmrW+ibmqMiyyJDdfXeM7KSHY4SOtlSGy0sULMXO1D7TdjTr+COWweq1M
jYBwhepxolZz8VdmHy2yK1tdPbMLs0EdS41eXf86ntGqxTrMitPYs3Y7AyEZwoVC4jseILOtunvF
cWFS8fdJvfz4RFQycwFmaN80dqZXCCTaTDnK7S1bKEvWQr5qrDPIlpplmIJJubjfLhVV62I8xb1Z
QYHb10BFSRAu35c55gmWhUwo6RSzML7f7W3dOGR1oKdFZXUGY1Ho+2pQke6RJHgH70l/rtToI6qh
K8FpMweRBELBQDhB6Meq2+XnNMLnWLo+w9c+qVJ+nmtszrckE+98sLyV35I2UJfdwiKQaKI4WFYt
uGFzDGE4sNzJf9EBBG4RGYYRtkW7eetlWRNz+LDhw7QqeHC58bRNvwOvsbwF2uVfkbCbafq60RTu
0e3BiJxfHTzS32EEGAGgw5j6A85bG52Uc3svjG2VLBvHQEa2b1FOnZ7idCIX01xeAARdymh5XU8f
YkUYxUlwnGwDeOK+NY7HUMHhE/Zmh1wkSkwFj2ArolwlOkcWo5tiJd4tQ6LzDKsHC2qcrWXNTf5x
kPDLmfPif1EmOhvscP1HjRrV8cCaoF+ClHsaLvr3MUwQiYZylqMD7N4mzrY191Taj79cCr0PPp12
fU/BEaUZDaunuW8BZGbWkP+6r5dY1AU9NU1ncbYCO/eOBU4xCbN8Ex2vzurZ4EX72i4K6ohYuiUO
xWoA3D7Hde/MGpOUNIzCUV62jSpQ7RugJKtXG7r7xd59IRjkeudMnzWnKxUhEHpLsUL+jiOkcP2o
rpbL4mooTUujnhRqdWDJupy6pgXyeriw7rTooeQ22sBfwe4LRF0LqgNJAkTjbFIlqZnXAIe9x/Yk
YxbBuqMo4ZR/T02Jm0+JQdBrPx1xfUtCq5KUBynNb0xShLGNXWyitlEYcH/AM4SCmKl3O1tGLFVN
K9axQSherKQ316v9JSabArI8enizlT6YqEK9JJr8yVuSZM6D5d5Hxh7IE1CFxu/ApgASz9w1j+88
nJd5eZofkrTN0XX3X526GPzMPk7S1eCgolbZcgAPO61xMTZxD0oA/5svMyQ8Z+aiTmajobceGYK9
9cUZQy9ctij9BaGjpfqtIfancXlI2Uar4oG6/raqsumaDlTYM50NZankmG9GobikxvbbXNqYA8Y3
v9i0gaYLEe3ZbZ/qFCO7iEGMxdtfyTpAKnEoTf2B5cBEisp+2azh/0j8V5UQ8y74bYf28W4lJ23u
h4ggDrnPRtlKd1tAA0feAAi7zBYkIdyuV5NTWc0wj1KcOTCSHOzB8hYkPSEWnSF8sUAVg+6EgCWf
UuEBMJN9S5+i9+05Kp+0a6CWTcAW8pOsQU4B90tEtNcp0KZyR4prI8WLzJDmYzEw5SJMDvcXqIcO
jngEprg6flNKumo+h7S7laA76Q1C07Ddm4O3abd9z5HWSkcBZPP7gsvp/Acxssdr+PsKe/2bKfIj
NESRlkOiOuBqsoOaJbW//Ok5UKozj8gvpg29qmn6gBVXFj6q8lvZz29RwHHm2qZt/B1sGM24peuk
VYgKXkTbLc8y9f1SGCEIKgcA6VP+eMJ9Q83P4WR+ChPY5D+SUmagIscIsA8EP5RabmPr04Sqcy0j
5iobeFxq9/v4lZ+yyPzloFbWzMCHWoVEbT0q6FsLoor6TacDn2bglgTYatn26CtM/FkrLKu7EIA5
2isTQovoNDUPWMxLB9Nlq7LPV8NodYLJ5Ckb35+4bGg5/ygfbHmc4TQ8s5JzdaZAf/4f5W5xW/ro
ERewZoELeJuZp0OVpkFH6JMgpRYJ/d7q3WFllUKHsR2VxblwVGaA8t2UZzQTo1ARfrTd6Bc/WMXS
jESeceGhCgZ9Jv5cvHuSe5E6D4CMXSqZQ+24m/D4GOUd0gbT9NmWEsnQgtRruoAlvxuNujbzjYZq
4598Xf221TjTY+rKRIZDqMKoUbsjAxH9Lm6yw0mmXXyFNyAMACKIV7eQGkmnEC1aoFoTIfHrQOpL
iA0Rdiu+fr/B1SnCHNFvNbMdyDGuywum910CamJ2dWmKBGj9c1bcUmxUqd3pQi8gBgEMM2GrWMh2
pg/xdW+3KNdkUrWebGu9VlwTMmIUyq/ZvT1FqBw4P8cst8vnfS96Kbz/uTjae+Ef5bM9XETq+839
2OFVi/CCZvW1sF+49/eOUEZdLN6KTjk73Meq2MMSqDyWbg1cYXgIhyZphFE3YCH61q6d+leoQwd0
I1lB6CXDDB9y/dtqV+SMPwHumrspIeMMDbV7xD5//nRWYxO7idts7GvRmPZCZNBstJfZNDwRHi2r
zwScTChYecuo60ZgCwuXg46cnrT8LNeQdaLr7hkHOsxXfLyRP/6UzROJaQK2QCIscYe5Q3dlYfj/
mLF4+qp9Wfdb1Bhqx3t8i6ddKCLr53G6ESoO0wPKN1etL5vxmYFHble6jURetOcNLjgBm5dEfMJ+
V4AEn+Gs0tkwkuTofFuGz4mPNB/t5RQnogduPuZ84A2PxIVEDjSMRI1A5bUin1OPc7+wD1eagFTr
+uN8vLLaYGGcVs5wwASbk3m+3MXOHOpPnJ2ngVh7Kihsuj/EnovoGXxCNRIz8TML5HNhWVcPbLCj
J8TZYc93YfyB54EThWPEq1c+SfdU/bAywzvrO0SgyBuKEYGCCJdV1GKEsUE+GZhwgYVL1b+Md1JV
AE8mQxIOzKDmXcwOxL8eBC8/1SumK6gTxntyFNtVOKRlJXqb+TBbie8FnxgqZqHVPoFjYscnHv3L
dVB/RXVFvQ9nMqm6ppxHQZHCOy9gKGJ/oho/6PWDu4M0A/WWKKN9XmDs7sirN76tFs7fIAnVG5G1
KQRQwWK8aDgZg+2pEaUwqA9rRyx1ZUlioQSdO1c/oDdizomYF4K3RYnvbrzMGGcJZEtOpoKnpFpS
bjxOHJUZoFO9EERi++sUr15U2b5fMwDPLrMarnE8X21gz/xigjuCHY6MX2k06oGyNeLi0IymDsoC
eJFKpoNo09PdCWpCod5qomv5NbfALfG0a0SaqImxqcDqAvBc444XuUC3IHSzXqJjInC0NvU5GUY3
7zG2JTlXf3uDaeiKrtJw7rajnrfoAmtZ/4APZqziMnnLKxu3s4NxqBdclbVKcLWpV6F0wzkIhAjU
fcVdc10ysDEUnlTQTHhPVlFsV8k6mLALvgnT47JTY+6y5d3fgHVb2RzHBqDSGP7C3vwPkVk83H7X
Vr3rJqim45PmfsFQQhG85rYBMvTQJRZH3zHCUVv17egXgSJU3YHrugkCBC84+O16SPUQx+NqX2Cr
8wynTCZDQTRkbsgNgPNaBws+geglqmDeevs+KnBwJx2HK9VetmGo9Fuoy3z0RPvOa+M8ZQ++gYEE
QX5UYujufup9Qsd/R+M6DwlDWsssOltRyd3Eawyui+CuooU+2Ct91gopXtb9GUBoLJF1HnRaKN6w
cVrjXZjOM6qeaSKdPJL6tBNafKx+fUtnOanMaSIjJ7gnIq9qPp3sZbZ7TN+hFgnpn+La9jxRba9o
g4ss6jSy4NpRGXqtsup73zvP9bwWEnO2pvoCRq2ph2CTv/w+jKjVlome0nHQBTDNsrkPpGSgNvJa
FuzRc6gn7Bj+1RN5x7+VW9XbtVRWJoV3hPvh5OyLlvu/A0Ns7tX2m3nCgSFwllJAAHAv+IZ3bS8f
FztS9oiFJLyPzVS4BJGuIaU/7UwTLkBi8otBEvrDID8ggcnJ8tjwxSAS+yUWcZgeYSlWe2dvK6/R
pvNiTJ/ak9+ggdbffmea8GL+0vYyeG3GW6LUFGqyUBBrcG63UrfAUxzcIu5X/6zNtKOkjm7cYBoc
ysEsao++zJux5jajE+4l47LTUoFR4iiF5YqqV+9NlHyGmVa09wYGg/E/PZiDeKYFa5bKW9QIEqyM
Q71E2DLykml/wKy79Gcxs3/QYzugsZIrzxPEdd6pDOa1MVgx0ysjZlULiI3dQ7JzPRUPv43z6q6g
muINSNRfOHEdekO2tpJqdwG6NNrpUAGw2jWb6SuMMAwxv9L3sU9h5gshsuNkXWq60jqsolcAMvh3
VpbQjaO5Q0nhJEuWQJuDEu7yDvU52BMeqdthCxknDiPWXDc9obOweA2+2gFQWnl6ho0QPACkgnQb
tFO91HrYseE7TYJRTUVg7jewDib0NAZeA7LejmPgdeiDlA8/gtw9ZQEmRotf7/xHV8K5rv0IGKdz
a02tKWVneb2TBMvVXkA0+ZVyJZqytQ0d1TLK7ke5/pJYevLhOJjhTyO2QrRj9ggWUo3T7MlZ8jpf
hZ39c8FzcFRsVYzXg3xAxy2la/48FF1q/iVrybKO9oqUEBVe7DzU7KgoG6TcyzUDYtpCNGlwHBd0
Hq4otYAvYI6qrzoh9n/Si62ZG0D5uuvFitYSp9yeVRIViKzZUreeX2wPv6fvHps338tI3fSKSwXV
5YRuEzU/Y1rQM4dl/ZhxKeIgeUM+S+7HlGc4EyOswwgMxWUG8r6siW5MaRFGTE6JqYB26+PNYv2l
eRMlstIMRPGM4w44GejGZoDCpunTGmriBBySC4TDThMM6XaUko6YjTYptn4ovlPsrQwhhmDarRJw
opnxuBgLsfRm8sn5ZEcNgxgQPKEYwrsCicIQWojUwzBhL18FeF0rDYoMNydRTZyloHzR21S485/N
S9FVhKBXfU75AhQ0NAxbB7n70HSdmbxvQLnR4zO5ZFVqC+UBNZ9mcKvknrfyMPelxwaRP0rsTtdc
LR98TXncQkeYijF1l/ihyAn0C339VwPgy6ZYrSOflrp5c+NTN5QW33pZIEEx4+6jauGUEbxV9ciX
gO0WhWacIk/4zuCdgAdO5wPbzeiddwuUCmI65vLhgRI5cbZbpoqayQAUP9lpsvof69SrVzYlN6fu
yCcl9t7K6Djnhc1SnRQtQ3GOQtVfwz9SXGjUZB+yZodeKmk5uL0ytxgcTbxViBVp6To/XGLoEv0P
S9DNVA8au6oICeN0BirfT1dpDvShgBWdmlt0oOC9O/ZmX1+D0tIYaP7WF0qx0te+hrzqNF64Vz6D
GNDi3XK4crPVuMzfaVfdcRnCHiLAEXjTofJ6DOMtLJ0pY6spnUi9WH0ZdT+htfCQ6+1HP9jYz1H1
Zap5lFGT3uW3jGxxs6KOmGmPybMc/Pg9Wwx7uKWqCd6uw4p8xFbKKHQqwiGdQn1CWQC17YCZ+zAN
mnnIct0bMUHeeeeU7bhDUBfmdsitTsHKDCYIsdbgURpkISYVbeZvJIdT02WKaCQX+dFj7uAWvkZ1
K18vAAYZfm9dnoAIEsoufLdfilKt3DirS6f0UDImiyAORO2xI83Y93CJTSg/Bg5BZW8lHvlFFFed
hrjx3CHukKF6T45U0r3ksFyzevmB9rFzP0Qa4A3N+fVMoqWcx1V9hH0TV26dRVrjCpZLhnLuOvHw
v+lQr1l4dcKs2P3tsovaTVXcBGGhFCXVUpW2tvJbmRGK+KXoISiaS5Vs7on+JXhiisYpe9QiHREh
G7g8KjdU4AP2XVlQ7Dz3of/szbIZUOmBDX+IEbvoU17NXODHX5YJq8UEPPJsYSu6TPyLrIsPm19b
E0ChOffdIQYREaunMiXhTONvya+q6GcqZcam6TagpW54k0mxDAxz/ldv0rKJ7PZIKW45ICIiULrX
tkV3V+jk/6mxNFkJ0Ew1jwC2F8XYs4cNDOAef6JEUpPAvzGm5vAU3xPdOq1tnnk7g/iz0zMJIu72
JNwjlnsG9Ua6AjOr1+MIVd21eRuICUgfKwRpaBkJFTo04T3KEDTJDptKcFpUdb+j1v1609GmESZm
kzTaGJhnLmlfTBjB0WMpJsT90Z/4WAocLyZm0zK0tplflAsaa/oJ02w2Q7+v+xrFhPGgqlp1vR6t
8q/xhd/sAbSXDtiZytak/7d6Zvovg/AIQjJWE+YL0369qa2VJHJOwuC1j1rUa4STYI7YCVzDUleR
Okvqe7mE2mY8f1lrJeSNDJgaAzGUDIDZdGBeUXyWftcU3RmjghMCh3Oxh8Wt1P/CYVIeZ4RWpYq2
tDAo3QKa8QKxw0NFBH6HJVzsKYm09Ub919iEtrtU/wv2nHrkAFbTu2DAb6qQRdoRTmW6HprNLcjB
uBcuGiqDsye+juViiJQLon0rQ9bIs0qpQ2KMSklr639MnhAc0LtGUjxXCZXmJp3fPia+qrwJd3kB
G26BdiUh0GC8P9+RS+c48QcrF4dZQPyfY/6EptWESyXWNoGHeNz+uEx7f+7Xd6loPiMx6aTEkBeY
KzUblcy2THJla2UwMWDcHaqspkO6PSrsJ6xtOG8in1hZbp9wk88oNtozlyEVgVBLi9+iWJsH4Pid
iDrP0HFhF1KAwI61eGq/OkfMf7EnHvmAOzLuXRNKKWLwSBN8PCewVq8Q+C0ufjw9u3oVhrd/wwGA
xLItTqQIzf+4IuNHZx/8clWyY3n5ib0Lwwfg9GR3OJFhsn0ltf4KxQRDCclOJ8SaW8tRSJcFF/s0
e2FN1swr72am03zftKRfq7jcRWiVo5geoCEx6p0qaxYBmwlqltYgwThftdfWb+KyNNzylcIJQDPF
SJXaKS4til40hixcqKaYPpvWgMYIDdR1vUZzrdC3Ancj7BRUHL8z3zY3KAijoQYNc4M8idApBVx1
dG7ne3FnjfObDJIwa79cl0V+s4FYS7O24Cp17pRYMfOrbAGPWQVU4p1n4rHZX4SyYRpoE7qvbskA
WRS63apMLDMmZztbyhH/cObo6PYINtU8WrdpUd1GOe3Q0l7TFHxY6Bj6WTMZQBjc8GkPyzoJhfht
itWG0gfzjDT9ComsV270/vuYtPWJX3wUo66XSGY0yRQh1Z/AEWqSGpJ6/Dbu9JuCFaA67cAtTU4/
F4vc1mVn551ATGnssv15j4T438Na/yF2SrD2LwwUTFIhVxKh66NgL8l3F+PsPdKPVg4jAfFmy92y
8cqoWj59oenYl8nynNg1EcbJym4qV9MZHqosO4eH2ygOCxdO2/58Ob7us3Z5Y+YF+w/E0VVWsPl3
GdsLJ9IM0F3eoO5bg+34ldkK7qc8hMOpZ7urbt172AA1GtaB6EwiVr7GGr1P4y2JWM0opjUZWpvq
z/qRHBg9mFFED97LIu0mCJLfXNIIyEdVPplyJo+EGczTKdfwExSuRBEWbTIch9559Vxxq0I81TmW
WQCUIIdRYYsKzWTbtRuqzVSGekGYNBvrDGQRSlXQ/pFWSVNlwLLYtAbmpyaCGf7f50GaoIcVxyWQ
e/iVJPnEOuznc0UHo2X87bYPJG/h5PysAl+dzK0HeYWL9aUp55hnDK6VdtwVYs6h6pCU6rm91D0d
8wIzSi3+xJPSrqGgs267bHk/MFGvC314jNUcMttd4ULC/Ht2VldgFCTq3zauo7uyfiML7pHT9F3g
OufO9j02ObX4Lgeuju8/d5ahW69AFIefej6uwp8zIBIR/5ROVrXawrUhxNdxVEmvz7qKB6ewuOm4
3bfeFhtUtDEYsxIGZgbF/UCcjoB3GiBWYWzmH8yukzf7fTBZdGQ8hgheNHn2WbhM65MoDLGIfv8P
yPGldUkrDQoi6afASXpQ2IlZD3IAASMU58npmYlZhAADhzM7UFZvvXRaPjo4Ag9niuXpyhY0pxJF
AJEt9FgR2HZHieLB/BstZGTEb3DCv5w6/QjDi/9lLpej7JWz6CVHgU5Kk9BNuaPtheOrwpkinX00
Zf+fUHhg3bt0+l6iTPx1g+WMRz9rn1UmfXY58RwhSz9PiS6wyFuOKJPg/kV0OiqYzcF52ptrhgvD
VNNf5PY/dZdj8IiUuNoKOd3/v6FOmT/5kPb/2ZgQE8bBb3lKbjrBdVaW9JO3efzOv4kDWMbL6QeG
nGGPk2H983/Xl7syvHR+Ttv/S5d5CKHtfArB7EwzPBPQlYa6uhIYUion62+sE8Cv8f/OZ4i+Pi5d
xlyY/Gl9Dr5MKgZWFH1v65A8G1zT9j9bkRpkaED8P/BCpN8PHWNutEgRjyZh8wfzoYHP0KZpVtJE
qsMmydSSWMquft0zai5xzWxD6dSDNTAEGCoIiQRAVG0ZzaQGq2OuQcKN3aNZgeSvug6mnJj0DYkP
ZLXQanfecj3siraLJFZ6CAqim3z1tm1FqBWYblcS9QUkuwLfDlGMtiOW0gOh+a9DsX9Xv8gf+yT7
wNVe3kNnPNzBKZEb08Fh33WnnKxyt6gc8ICrS5YPorTn/XSJyt3tQeM3KwNFXjnsoNSLXhEfMuXA
0uCcITQ2Q49DVoi6ZNubUKjvPDngHNZDLN5IwH8c6R2q1UaHArj1ypGwwF/c6BC2gDB/SBmU81G/
wNEavNEXvNI87AhoVYx2JluAnN0cG5LgaYkhkmN+PkIjwcwgxdXNpTErKHOJ5TGdefRjXJFltq3R
hbOEi4JBecQftHTWYJgn2wtHFRWRFc2g+f2ilusOdxK2vAPqZfhob2G3sk1FYVlQBtlvkwYF7hnA
mDZefODsqqOEjfBVONUMTGd1kcn7JO3ZMkQbiVrZSqGmmHnFVTkL54+8FLsndvgMdcL28tXxH9hG
v91UuHyQfgx2w87pZpkXbnw2sihT0trgOkGrQdMw28chO5HyIPMLCUf6xQLl4XP6myMrAEEw66Ky
UgcfEdZcx1ysjnEtFvdck+5Kq6AzWfkMOiKyDMmx4aNUXavQCEJkI0zPE5wYhYM/wxuJ40y5X5HK
yfBRxyR5OW4kxIDHW+aArvruGKT5DUiP3s4XjUknOsYGxT8N+TuR8EPFB6ame4z1JprLxEaKbEyE
DBtHhYyDl9eHnCWPsdB3VfEhlyorfaXVwEGg4DLI8F3j5fanOJzcf7f4th/Nth9auv12zXZRV6SL
5700w6TAGjGz34W8271JpSRvpvtfzNRneq6442xmN6/cmhlnG8Vhbjs7VcERhSXg0X07dH/VC3v4
gOeP5kX6h8HQE397vVEneESRZal27V/3gRv2ofJby35lfHyxIrkQz6n/Rwi7VW7254grOkf/ME4w
L8uYsJ9dEffCedPhsSHTRIWJKoMFZRIoRiYif7xAEs7PBo777yYVDmZ6XLBjMyZHD5cq1nhJL7xN
mloA69ViO3CTc06aRrfN8ktCUUJV61DdOMj5MQoH3dF2HRhArCKvvNJTuTAgEzUJgoTaUp83dfW8
qM9Z8jcWPLvuji6wiE7m4ipv893If4GhNAo1f53TyTLCIdM/46vmctE1kRsW0GMR082tAlGw1VWW
coJnuYRyyXJ1kHLOIK9yIjfGyKc2e/ubpG2s7b0QeKerisC5UpgtF+4ItsFdsNa6/BM3MoUtWnU4
qBy/t1DdHxol156q5OxjOlGYHxrtqXi7jmpCybYMPKdM8iHwoVrEqV4lwSTRfEClbhTxX/CSQe/4
QZ5cp85uw+2/ddVr4fM2faONpEhQo5F2VwxuZXpl8tzIo8s5e6Bnn5CIw+MheWZ9Qjw8PmNPmGZK
KZE11tTPS1cgD0Pxx205+uxQj+qxb/RgtPOg/wUhvuQ2CA9p/Ru10C191ui/7ew4MgBNA1e4XA+8
xfK3cnNNn3erQbO3vF1GgH9p+cc8FppgTXP9nk6VLl+dE2EOe4dqca/2JrEN0W+nZx2Y4kpqmQMr
873r4h0g/43nKR9ciTQcMfxnoSAK5LfnRd0oUorQFULgG2Zi9EAedSFxrbcU6CReyoCF70ZXIJnE
8EfGj/FCNcFY8XsOh1tzYObhemKaTfHTMiuOIeQMNVgcoAeXEq2NoUoEa90e7IX3v1Cb3Cir4ywN
3P+nVKBAcMjQBaH9Og2cYmeMuTK38mc7DM2KBdHFidFBwhhFSy+mqK4r9LHcSpFSWb74/sowx+Hl
ZiC9afxZXeTeqEaiaASikKAf5NEUDiamU6wH3Frs33t8hfR9MDReU0+ZoDEQ4NVEPL0mdQmulzpr
vkieCGt7+W98qN+yYPP60KbjNuXOJ25Apu61Qqc+OgtYn4uAvtPSTWZYLbTpV20p3YzB9vIxDxt3
XT2qy+W97kKW8raOdHBWVLrq9S4rAaUQVuadk6AfJL0m8MeLImkFVdA+v/tK/nfMwN6UgCdbbDMt
QAk92NVZxvW0+gdJitk6UdA6f4hphftnd5z+vl3H5R/Za1yJtLgX2WGY+P8q8vsLJMIsKULi/VEL
Kog1+8XIIg+OxacYuWCCxEQ6XIkI974Rm5A1BeXARLxygdKdVTKYluTjN1S9XxrZpJrvrJG7hN5Z
WeA3ueJqTw7ioQDJEl9U/HCJsvDtcaf5Fek6AkEZ0JCTxKifvXdYqhYwOc9QR2ueXPww9S6lAMir
2E64tw7xQZNV27MQDOLTG+o8ZXZXHqJNeRAunakq+1eV7TFGa3AiLUDQ7HWloH8UZmQa+/Jteb0M
GOPRuKKJ2Mqv3Eg+U6TnLT83YKoecvmuIydwEtrleBL32A0xI8S4IR/goRZnRsk6/ynNVPfq4VkN
e/L9JMDjyh5nW08lV1SZQuF7hl0y0wywz6SPQ/O9oZWuHHHbhkPivY0oRLI+B64xHXuaVX1PtEbD
/H96thOhQ3IbWWFqWJqVYb+AFUEwu1LUNl8u153XAUQlg8fQzXcV4IIm42lHNJ3POSfOro+pmqbj
4bLB9zDVtxULnD6LHFDc9v/m+onX50K9qQ+2X0OxJyOFTISmqDHwV4nojIeBLrvD3WzCkmMIfF0l
jbKQv9Fz6SxZrdN/aEKvInNALrzZk4fllnKmR+VH7rlI2LtmUyflhtmdhtSIAGqGIF6c7pDQ9tbf
/7GYKw5sy33pgYRnYDkz2qXoO6Vmx3CpXGJZJ3Qghy69KaTI/+gzkfoPqSi9NwqTQbpuNJO03OS0
BB+emb3txaTWPM2ntzYKxtL60EOT3styqhvJvu5A/2yly3vLzjs9UZoKVaxN6M+HtjiNXb2AWEeG
wmUEvZrtwWShJFEjaVjwRaGsA+3Q5lSU9X5etjTH56E+K+hmuEa3jq3gsjh7KzFXAJDXsIEAdz05
dw+vyTTUjVJ6GvfiZobVVMV6JVQ38zY3T5pDYdXL/4YYl6iZlt0mxJQORLN5NZkOn4HEI/fSQl9O
VaP6vU/QyJRRpEtNDY9j9xO+ckd5j1Byia6Jtvp/Za8MAzXD5kyQ7v+yIV4FaVreonBjbrABJQgG
6RCz9ncc9zyZOhlt2jI+6qSaSS0HfuXqedCkOdronpyXUMq2vGAe1/w5K/bsw1cHheDNd+T7OM4C
p31WFiA03Sh8DfG/qNXfCj49Y/ox0U8mDMXogv/91kHb+8JmpMwQOqu7eXn/dGhlyM+Xu6J+0I67
i+N+qAocxbdefXXw115S0WBzjPq5F2r02xhHPwbYahblml9P1ocRzLc6CxrVUniGWPg7xod9xQpO
+1/b4ZtkvTkYNDu81h/J4ilZ4UFNSgXloEOkhoubWKBuRi68GPMaO8XJl38DjxF5k75ccP92203/
Dp4b3JyPKG5yGOnGkAHs0RIx2M5UL0U9qhF1bCnk+v/EUMgYuPHPsMgUKIOC96p6bNlFhDPcvrte
DveCnhHyraZWMqRF9pVlApxwGdl6emcoOB+FP2SzYmZ8k9iA/r2N9yHbGOg7iSiIWVVFwsau+LMs
Uv9dfE8MOl6v9esF6JY304leFIzcd+n6OV0FIKqR/yPZnm5P2GFxUU749fs13iJ9TVFrpPew5O0e
9nbpx5lMS3RSqFhj/mSuJbvKV2FLFbSNnQRMlh6OmgywmlG4/ibJ/wDmMg5ty8Ygesrt8AVxTUl+
6Kp7BtoO0wwBc47wfS6MJYB5kubl/jUuqk3cXhIya6JqKp2vsYyZfbG497CsSiNi+WhR2smlIohT
QdiQh+IifA5oukCaqqyIW8Yblh0NcUg4b/iTLVW3ECyD+HbdCF3u7xnruEKit3hSfYpYxn3eoE2b
s/TDIuqyV7c7idTA9UUW6bzs+N5gkiAkdC1AHYuA+j6woo7Iy+EidUCCTpRv69VVdp7q60QdMaza
z16uQfmNEd8UZW4pcPUJSnxjEvVBl/iyur4BN42CnxGFcN4sLqTKYrR8dwoDsf9QcNEe+w0eu0WG
OfRmZcFmKfKoj07ASNtCmOt1F3OKy+xCD92yVhLd+woqEvCuzdADQcfQrY79rjL3emyy0AZvk/Qz
0znjWAna9zYahR6q6CFhw9Po/yoCd5FMtrKt13P9ROluoCQk5R78JB9qOKYd+MH1j+HQdxYIMWKW
S+8E4PnddAFUDlHUyaqgtlpjG1ozbqXJcm7A6RjTZ+uTq8yUv99R9FB/Np0ySDWBXFslyHIUA8U2
X51uJ74rI4Qig7cTpwBOaU7yQ3fam7P39RvmsLIf7VkuQAflhhb5YqeMOdTkHyVvONFnw5bS84m+
05Zlu7l9IkRJSXBsW9y80ga5hiMMEInCKDFovDlvI3mFIryyzml/7xQqptG+ZzIRKMpEijo4xIAI
hcAPKwHETGdpdyNI1RRXWXaqVd7iGqYA4F360r13Prs9UrMiXEB8wzvV4jyKMIFzkzHe/4wPNGOl
uW1D5UP82Bt/YU5BZEHCFQJdkByspoY2BO4WZKpSANq/rfZ4T3svdQ4BQS9yQ4oG7nkgk1g9I/Au
oYL3KYXf7VEoPGpWv7r4XX6poE2ADcGSRE/Owkdua5p5k9u2HFQ/V37+7SBukSpay6MM8PQPCpwY
K3fAo2qg/1Wh9r3gfAHFn93ISeFTEvKlimqqqclrNLarL9bDbhMkTVtIpMHYfBZ0NZmtZwzc3Ij9
yJU42xBaf7nTllW5mY6Efw9xbW9orXZNZ9jukCgN8cvh4qNGbAPvUobufdE4wKnWwoQbq5JIwtBB
jRIH9QgXCBoeK+0HClMf4Qor39+Czo+zSQwg04fJAmFCdIzQBgCdXfj4YOedKKpycgsiVMYpiyLK
HNjTtKnhXTVYg+I6M+d//ZTKJX8ixAUNSWhf6Lo9f6+igmIjiXK6cIKp5R+ipd89XvBY8PqdA7hC
ldNyrJzw++WjtGK/ZUMtYjOzqrD4Tg2DAfC3KrTIcva4C86WRv6MtTF4WeF3uXh9suaKsTuB8jMM
RnahtcpPFxdHWL6sUfZ9cub8RpRo7+sQMvI4tw5c5v6s/cDD45hD8C0G567Kgufrm8gqfOaMjLRC
sENQhQY2aQ+Je3QYlsGk07KPLucqLFX+PWe/KvQjkTgR+/Q8l1eafdt45jEz90wNtSkDmAAtUX/Z
B/wuwkPhl6dfURrsyfDzhQG7A/9zhau3VZz9JkMJStE1g3Ocy8xQXHMRRircpe0ReHnPjX5NsTaD
YHpBEDbUV0ry7wYI3ujwwi9DabOcLojA+WRlRz66lZLqG4frxUYKWNlGCmX8B68NLzRQ7+YWNDbm
YR+y6/q7lIXzMmOR+1TNVAQ3JP1Zo/Xlp4vfGtSiD9Q5jOvkK4gC3j9LvlHjL7V+wE0vv0JWDvZC
NB4v/fAINrsbWeAAQTnl4o+ABTH0lPIvEYLXPDkK7JmtGLSAam1eYWTMJahmMc4Q4MtFCPdZjYGm
8eVlFvt+uiq1aVhoHLuX6uxaqvN7z0ADt2dpC5CxofzbYZG2GFcPXAAkPWXqHnILK4mexakA7tZz
JzwIsyUJGJ/dLvrhIhZSBRUPAIyNrp70MmJwi5p6Bd0gc+LNezH9aVZk+bC64tLWaX+nAnT9UYZY
hnn771mPSUU6tklbpsjvj0I0BWienr3x6AUtNKEOL1fknf8Atgr5uYBcIyQYkEYUbasyu9lBDme/
DQyTuJmkHwu0SEaN7o1KWFjXOhS1n4egS8decyY/LfeeMBiPN8xSA/ALC6kq6CgpEQN5oe2gvvXC
NBbIkn8h7YKdaPwVJqga4NGaBrjeQR5B5EGUL2737kbmtp+9pybwvmMKCMa2qJDeMWTELgjHSRA+
0fXe1pYkJjIBvkVnuTVLjtytYk2of0gUPSJKFmRGBnbkhGHEkaCPXBVxTLemflmuVGdXbEsJXdLI
pUQIWrafCZP6ntu2vWK3+T+MsfqXStB9rNQlMBZG+XsgYp9EF3bRs/L+6SxLt9YdM8jBRxxwVu88
66UM0F+NNuonBMeLWQfC5qaH7tNddNWNd+FoYBGmPm66kZVGiKeNO2KN+6iZEieyuR13cAJNNgnV
cavUyrjnfFiSf2du5+eNr8OUsYQVILzkqPKe+fV/Ti61+7IngEOaVJk51emGaYL6flWewQ5JbX4A
1L5THrhgc/3Aw4Am0MNaRTOr8MOnz2jcmANQmb6Wlfe+emJqSArgLdaziud0t8UQdHmguUvLHzbi
6hHLa0lWNilxh6Sawa5l/vyCVODA1FdpCRhYblsyYKYX9NvXu9iSnZZKX+sVsW1Zd6KBtlJJMgVS
cK7zkkAeLCkg9oj1/cPwawjVoBcH/uakr2w4ioSg46i4Q0BRem1DY4/2fqJnAaENM0LM1P3zyNjd
mErtZkGAUsmBQA6IcFNacSO4t3T+VRoDbx6MlryslaF6qYKPchyXZcxlQGbU9n3u7l/uJLmNKnm9
DgqOD8waQkhzvE2ehwLbACQPlLtKBDDVmwnnQ4XdlrGhoAj5LJgZygnxGOaLitDZsU30FS/g29TU
1RmIU/3tYk+YJUeUi+1melARRkQhClRO7U0/TJRwChGYwU9xGCMoJU7oJQ0Xrl/BkH6z6X+iurLi
4V+Oz8dBeXsSiABe/B6lV1mzZKAzjjyvpQcgnOyWRO6fQKfy+hxBjNP5GMEc+Kww8ZxzCfT/kiu7
khe9TtKG1zZBKFZK4p8CwBZxibhVr5xcfcmQUHb2orJmItuVCbDCyTWXcYjCgDSEw2et/QQO2NSc
iXshZH9/EFTeSeJqWsZc+UeRJFiBEVgjVP6DmQJCBsn9SA7AnKIFkiBeWXRAyaUVPsYY7QomIiXE
2CHsYqOPFFkQ4zStVM2/ufV0/MTpx++NzrU8My/5Gm94jiOrWbCqYymxjatQjMdaGmrxaCTBCrlk
WLuLFlfgsyH91+uf286TcQHTvMF3ADcL/4wlR4seaYgMGZgU0N8eOaCwWmhxnS08gQ5LMpFFhXlF
x81LmRhCA1sEba7eKHoO6/SIfETJ2mpq1ygvLlOVuoFxRzP9KE8ulJSyXV5kIIcdw32SMEVFsml9
qrCkDZknl9peQOPTHfD6tIcja1i8bn5tCyEqJMJby5azTYsTcaGtXK2YUzegtx6hrDSH7jSfQ3r3
FCM97nA6pWpSayOyWAv20yfdwSfdyHViJ1+6XXH89m0wy29qNN00G+lyKEW9hDA2VDlUZDLdQ9vx
Ci45uuFZ38iQX04h0nrKRh6eIOS4oPNBcpQG6J5GMtKK3S9ujzxwVz69/wv0OMYDiavrK/Arn0mJ
NbTM0fwjhSAECjMYOc0pM4bGyKDn74DbMenXSEGnHLqrdx5zPmnOkLWumciPgB0B7uhShBq9i6Y/
bx6dUtJSXIXAnaOByccc9ofI79/oscdXZ5t8Z37J135Y6AV7ykB9gE4p1cQJgfovkxPDfe5y/Uby
Dt/0ENqV9605r6yXF9ijSj2u6ZE4ggimMHnBC+D9YgTlobcEi46jVML5xFHtyayqba5hvT+2yge4
maZt0jE2T4umAWAQpfeobUmuevi2dIAz/RdA+iz7tN/bT23KeKF8VT/djTJAGZIQGfXQGvTZsDkm
mqjT4nNMDoRJPyDAvl+B77zU9QKP4+l6KrmPbI+tEbQnxeZV9SWxBKaSMTJpnt44tv6g+RaBAVuY
+j00s3Fu/7OTegm76+5sizLQQQ7atcOwqKZ8S3ws7Tg3E1Q7JyOlOwvBU/jaIS/5pfbe2HdjfOEA
dI7wqOiwtbYE/SD8hF/c0m7vvsv8SLinRTupGUFT2b1UyZG48eXQZU512rCw3FWa4snqHp06JZl+
9L2RSLbmmxIibsSdzPE+2D/JM1rWi9hwsyVQrGIpq8OLz/0A3Bbjwe+jL8pGlVHOpFbYdkwsiG1Z
mWqoHBiG243QWG3xIfcJt8l9rW+wkCakCCI8ggR+oJHqIlCYL0SmepXWnKrgawgeEaz8nByVcNpS
xLxL3QheQLdnHishYASv1DKsbb28oZoRlFeSFmzwotCWgFMTuEYKcWlURLrggd4Niyfr7JnjECxy
dWRFy4eNh1w5FeS5IVZqoAOtEsPIHlX5QVJNySDol9gdDBL2mw2qDKM1Z09y5RFzLOwdBlyb0Ayw
eQ1fgR2QD+4nJpXUYLBDGHuM7gxcxI5UWkRBhP62qmeNOi181vSAYyB02Gvr7Tad+0HsLGCc7yME
/BrDyIjR7z7RNDowcNwESkUVMS7lsfv0kUt/huvWGtzaMXj/m9rLnesuCvAuiNTzHuiyVkrVt7Xr
MHeagKjgrdF2dh83gyUV+Zs7t4Q3VvBAqTaegrr129IPthOV3lx7g1pBP2Ra2GDd1dEgp0hQP3OJ
xyBnOXx1wkxpyGaqu/qUc2qU0v2WUE/6Xg6k0n/4n3tyzABL1cqGqvefDjVCGf4l/n29BAHEMNv9
5T070dfihkKrlP7NY4gEZOQJm9GCY/WQ81+uhyCHCuw/eUauO/WXqu6rp/Wh7fcGhOx+OcF/E7N1
hiCBytZUtnIa4Pa1e7579Y+UYBrcqVnRn2QYgCVQq+c7tYO1/5OyACgXQALmWzudweNooPxXI7K0
Jlp47FBhAdI+3m+rYg2/NPCl6uoF8mUqK+ckKh5+GzM+vtlX8BvnHPRxo7v2HvQ3y1Slh4vya7YZ
qR/ZU+oeqWbTKZDG92ex8XNHUC9BOKy0ipXjsC8IkbhJczY3P+kNEbqsF8sULchSybtur7ufv8l+
bDf3kwO2jb+nAAIhAhfPJHXXUNpDYvr3o4ix4Fs+p8I96GOUUYPDFPalyspjW8/qysFnz5DT5Bpd
0RcgzaxOpn1c42JTzNsodymaSZQ5KB1mFLdYWeib/C8nOnI+upixR/+Ab+qxhPv6dSCexZBSaNgC
VDLykZDWZ3/1LHFz06uoiFlAf7QhldN0JNlF3YodvyfYIe/44He5bT4ISpGW5JQb3CJGOWUc0U/5
I0oVSlWxRWfWeGfJvBAEdLvAVgD1JGw1kcAtD+izPERa85EtiYDLhbSyyqVaCA6V3dYwmwf61Yig
06+sCfBq6jNkuKYWGqTtSTmqOFIlYDu7GnICLW4OnMM4mRtfe7tgEXkEOpK489cAVUx7BKN5zGfZ
GZ5aa9bjZF0wNeCXP5iKUTnivQvGLlf8dYfHboXJsqH2gPyzw/OHhnjsYSYr43oAVXZCkQPJRhfz
4sYeL/PPAA/LgOaBftx2azIcU24hFBY76saiOM5CwrhouHftoZcozpMEFfjNsmSMtKgy9KfxUUZi
tZI9ycDCowqWnghywLXN75lbqCEVpo/BbNf4lJyBSoJjpaI7373d4kNxXK0RX9OtCYzh/VEWtCfy
f15+4GPv03sSNX6zGlJMqPMw/THrarJ8rK3H1i4Nd5Ul8w1hTClFLkilfW+W2yoXHCEy0gcEhVO4
f/rQsF04mFFFeakQszGXUao//zBfi2gFnUsdMAga8dixEcykkBotg1KqWh8dU2hL8TgLs5+miYYg
GCpNnpVqBrsHuPKB8fnj9x0WtHQrhB26cWej0XS1+OtYsFCS9vfcrBAE5adgGkk3J8vG4M9C6PKA
HhoAoCc9wNdV5UjDDFOtw7W8gAKhmKqbFfgo6OEVGsTz5wSiwQTBfbqWovE8QlMAOuWf9nkrN4xH
Oxywpjy6jMVH4r8g/m2JUvUYQK6bYCpUfUt+omFQ8/k71yYSuGdM3eWMS/OtW/Cow5zJjW+KhRnA
sKgfyzdO6g8PrJzcFEjktqZjnJIjSPzKl+l1Lp1EOQWJYkNBMSzGUfbzl7zwQpvBqKHIU+CX5MG5
PMIoXTA+OzvdQrLGSBQaatRSTwIn7T8/CbANBLT9+ZRE3MdQqI/9ar+UMpzEOuvDmph8Q7MEYew+
hKFrQ3KrDd997F6Qff2YfEjTnqTvz/94Y3k8u0nmy6b8G968vzxYRFHcZho8wfkxtoPXUqAeOihK
Bpn+cYp4jtiEayeF6/mZtvYBbWb+xNI9e3VFH14kJV+DkC6UeO1RknSpFtL2Bv46FnKWQ7FxvyHK
i8xsAsn4YeVITvtMhQWrveAgCFgd76ZV8sEUcLFZ7c+xU8EN+14enHUgPWH5tfd+C64js94y1vvG
D0uK3RpI/Pyjb6PdYWgKt6c0k32rMovQQg/zBbggBUJ4ZYaKC/0jw9TSwPgizheFyrZr5OGUXvV1
SDc76NHz5I85g2+o6rYUEbTYgizOtQWH4OVvvDrcGZjHtILOFirT1R8/cwUONHYPXchHACPFiXHd
SplJGaFoDw1lpIOhgfa2OtTNgQtSJ1x5UX4k4qqyPcCqPeH56joRLBBnB4lclz96vfCxSFZLxLVt
pOtrOSXLtvGazKrbjYvQavLWlVphAHRuv+09O+Jn9OICfJ8zAWnGyTGVUFZL9UA4tnjavYH313oE
c7NQimcYdZgSMI157Ti5uKvYWElL/9OgBHuwLHwjVWhu1JImHFnhM4CVp7R0TmKMQjNuIePAUNYb
xgRsSCWU5TRwxnyQqLyF3RNAIrT1lLN564cTYFdb9tMA9XdJ4dEYPeQKGVMoWEC6Qi7VsnqOy2qr
fvZC5auFpils6D3u/akIMR6zPxhE9yMmob948fxUOefuf3izRUT1uRHlwwPSlEFwli53XnP+0qYA
4m+Vo8UMCucmTSaM/zdUJsKsfBPQ5aXlJ4DdtA+twTjr8BszU6DeR9jYNKmGtvoSKfyCzREVs8HL
flNyhEeJYe3KJnlNRNEJEsYi7HDlCBO2VSLx3bpVju6p7a0E2d2RLpMBlixh11UHrKUYdrCpQMCM
RQ62Ue7mCiiVlLdbwXC3aPIUu3xSt3TCp1iKslfxP4conSU4elDW1zOMUXZOWCqqDhu6BVW2TW27
ZhLnMD+HC3THCv9BQOwXMqoJt+H5u31T2/c4t6I+XCJwSxyZQ3nzZGQ/bRCrX9PkGaWsQlkvV74t
/Zmk3hZQ2gPqHbTPAz+Gnsatnl06GvfMqR4OXgVG+JxqLN52NTG7lDgjTwN3fYNnTK1pgh7baqr2
WBGnFrJYGxNFOaGEfNFZImuPv92eyO0LA+OT/d3iEvuTtWt8HaKRyNzBXS8fg/YLp54BtqL/ZQ87
2X7N8SIjllYLNFP7g3V+cywEwkAZxQDDy2TGaq5pxZ5EH8dSaLQA4R/JLiSVsnJdirL4F8hYBNPG
1yxte41sW91EiRGgA03TJuKATr0VF8Cqt2BlTCW91hpnzH246TRoub/Wq76pQBO+M74/ezQDAuKi
Q68YTTgsTXccuJCVoKP1cdVV2NC/UNDV12k8HHrvpzWezQIHtcGyhg5tM5fUa8FZe7gAGxndRlkY
bAopBctIdDUhzjjmhqIU5NA2tPl5Z8eMpmUHJoGMnW25flQN75bdBQvLMPEPOa7kmNve2OkCRniW
iA/vZO21vg+aa7R0hSVkSXYNwAEkQju7z76J9llQzfjQN6fuqk3c/c2CbHxuw8HqF77Q1ML1ei1i
TcVStAqHPDMl6Pcnxp5yjNsTnXwr0FuWsMxnzGMVuZlpjauzj1wMkJHb96i+K84WDM3h1iOur82X
x5CRe66ILIpwBfXtpdE4VxvjC3zTU31xfvY8HIR9H9Y212RRFZjQf4uUIKFkQ7fy+z2j30WWcsnZ
uxWlde3jejHO3BpX2gZnxhOR5wAy9CnA/ddeIbvpi1lzxhTJLKds63WTJvYMjQDsn6PRooLZQgsq
zOA0rrOb9lj6QmZ+usCfbN4YsGhxBt95Cw7c6Jk1WOuDOREiI6GAmNPq9NQUZ0ynjZkKQME9RGpa
onsuAK9JrxAohRNjZFTOmnBJwgl6FxfKU/NWiyzGDIMS/jiBxm7wcTE+wNXKXhr58ZsMC69lg8h3
ppSwgQqaJlo7SD5kReKOduBfqGuM8fPaENmMQUY2o969QFcEbwFWOgEkL8tHM3BNX+PdC2THl2HC
9NaEwcLMMoAuCc2tildnRBVVvQdVEloypGp9L/nocDNga9XKZ9xKXLKdz04gZHtD3oFohel17Yjt
Zqc//kKC6jSJYIwSr5cvlSAwE1upvHQ4XZUUqmNilOKuIuvx3GCsPPStUcKuXH+ld4BQfHlQfFpN
sz8C6Vq3YrVFAqkm+CQTI0cWy0yXnEr3B4Ax55KT3i8VKRWwSKZGWjYURKFFZSJkzXuAwLrpFsmx
/0nv3RFnv/ucBOAjry8+WxRENHeQKXTydqRCCmsW+h8yd77s5WMc2QqCCDtiM419nEiFDU3SiwDC
KvH6DKqUmzVhtIHRz+es6d+vEBUwzr+HbSaCQTwKgfzEnSU3ts8Vww+jiw1gfsvJHjfXgdnPabE8
g7dd+Pc64jni6KX8j39+O4+fotOc4XXCA6rc/vV4pCw9B6rSv/8ynBm/PkSjkHxiBoIclxRHUH+y
D07MlLv/DQlJM7T+gFf3VsugfLkL97pGJq29EmQ/4uKj0Z5rK7IVyXMwCEmyjG24mh5RaAyIdqYt
o3yZhcHfCvlruQ+woZNnUSZ/0xKE/2lSoXbnyJY7rwNl66dVgPFd+D//K6+QOZZGfTNINoyIy58u
40XBTzM6jQa2Y3NnZPR/HbvlYap8PKCxfXsZwku02c/fQciVsJQ+qIcL2c9g0xVq7Rwbird4OrUM
JDcsGKmj4y0X6iCuStLEmgPSgdSh5EvqZgz0aE6ZsYBjwEz83S1GWUw9NL7IKEwDnodKXH7Kmm2n
yWDAwgRZPocE+162WeaJG+zlbqMEpfQkWtglxPAX3yXETrD15tT/qKmfA7sMqCV6KlwADTVmeBIK
nUjxxrOgzxFPtOFKBYX6Orw0e7kxFo78CR90TsZoEiBFFxDJPV4EJHeI5rLvOUvLURncVtlN/N6s
R+lYGQhx8p6oRfAlvibQ8kRzPBU93onOyT4xHovMBvDYgxFtnR1zctK/YaXolcmjB4dmstTElUum
N4ECPX0nWR0xBDlvBkvNTeav+QfEWs25a4idUDbzSGq7IpUGxsOAXMNXtLmkYvUuq77rZrab/5JA
pZCePOkQjuX3KARG9BeIsWvQE1qZ5T5iS1oBYZKd3R2O5ZEJErny42uiUQWohWqL+GY8RzMl7fxl
pdlvETnh87rl125221DHYm3fzII3JScBBs/IBih1BzPF8DTOEohlYm7BkereedEyeAnO4vnoh82C
Jt34zxDsYswb5zJbEnrYvDzwGMZlbzMCdE0cgTux5uA0JpuvArDHYd1nIVGd89K2OmqsoR+nKqKo
wHHMsN+Qk+dzlhs217RPFfqf0uHURTv3Qwfoy9+jgBr0AR5CY5US40OlFWvwLc/h5D1ZDF3o5TEQ
bNCKAeeSF6mRWlzwK+N0FuIjzGwhhljzxXvXtdQ6+xOPdtMsoxH7uUsohRfoALCdEwiuBReNaOte
a/ra9KIqRcOZ02ul1g/WpcDdqq52CarkVLy5FZboUMCSKt9WV+R6h0/h+DqG2meUNbsR1T5kV65r
UFG8mTccn+7kNPo47vgYT2dWwY+B5XJFiG4OSn0p33Lc1vdVb2aZGECvKyPbSE7BEemZi5zMGUEi
Hgu4PZ/4/tKPhLutMCqv7IUYCbfkicjH4uyUl8XOHCiMHUtDApvHCDk2PS8hDHjl/mp9NA9Dcj0h
1hIFqNWrH1Pyen/tN31h7JP/XveXIKdECgQq8OQsY9YFecc+e6anpNK2MaYj5CXL4+CjRvE/JH+N
mMHVbrGc7uY8ADGykMtwnTXGBXfL/+8ktbOwEsVC72mXL7iKBAKPzvykyssNpk+S+AlriZ4yIJzk
WL4CPHSrAdAVQBgD/qBgwHX/sTehZ2A91BPU6qTFPJpKSKvItEwhPxn2iSe1+a1ReNgS+uV9PFvc
Y7RtuxhMD/3yWFaKTWy5dx8IjZrVgvOZ+ryMV/nAcdvF8R+esdx58wShyhs7KpCdh0PlI/ah0TFG
gu9BLZ7uZ+/lUJpOAiPgMJQw9wlNVltm2/l7DARsTSyCN/BGMA/MTzK0mNaOVesxZWHYwYnYsrVa
WmJBFjThbs6wcOfEovO/9szy6OirG5qpNOYEtkIBJjmRQves57UD+/em8nPzH66Sxagg5U1zahim
XPO+ySWi820duubLGSnFxt4Hh9vKBAEIv6USoGrdumZwfVvar3f0WA/Q+mIw3OkPeFvzSc+Ip1xw
DD9J/9HLH325bwcXvKNl0h+2z4FzAu6mqjDtNoySq+OiwR0L3XOf/VqkPr1qdAIrjk4RTLIZMRdV
6TcBipz5JIeOfJoLM4hlVFvO/YvocUCy+58W4mv/xWEs8Ac/BNEyzZCsvr9e89VqON+FFzUweuho
OozoYGNzylnAXKp5+3NfYObGcsy1b3OmM6MIqCzfrisyLzWizE0oi5zSA2M3cMe3+IXYxbbl8RuN
x9HJJEPbHlWISocaZCV2+iB6sbYGQG8pFAOqFob5AGD888NWQ46RxjStZaVYWK11pruPqcMsgmic
hctRJfez0U9PlBuveM9E88HzqSZxs3ubK+1ZZd1pRpnvV5GsRLZv3Ogr9yZB67Ffl9Xi2bSVPp6M
/k2Y5pMEqSdYnpqBQv69dJfwPYgJO5Qh2vyLm6oF5JNX9sJr0eSmFzMNdyADTst2bfl2JrqerZAm
PoXxIHoyRSsJANIALmqwNzpSDPFxaVDB5BT/xEDd8AsXgXjQhV4iF9ljFgJv2147MPQAsEETtp0A
ipwWB1+3VXoKrP3ULJNpeEOj3G9GP677Xj5Vi1JnjVbzEb4NZhp5t1kxrQPPV/3XeQ5Dh8S4dM0T
zg7pdhDu/OgpdThoc4opkoeSLOVtXpnvcVnY2ns7T5VG90OhbCJeGQjum6m5DEVhNjB0V294EgYs
Of1cS6gI/ScqL6i2Rd9Jk0cloRww9imfx8JUfX7XJTkQ4pvhfqBOZeXSnTiLvxhmz9dFbVE2Rk9e
baUCVwfhewiTcxozpeRyuhtp2YgXpvrNZ2tg5sStmuyFH9Z8pa+/NoMr+nn3Aa6oSdS+stzsMjAL
4b3FzuTiqSFDLvh6y/OqRiJ0wy4b+m1rg21TEoTz9Or2kKiEQCTim2L7KBuSqCaLwRVGiA/yc46/
VHDT/hE5ympDUCT2h9534h+rDuxMiScwaJ2ZLx9XyHAcTMB7c4uLeGJVQ9V6NOJtD0pYIK5e8Fpj
rbMyVLghNOmqIE0tyXv45YyLe1+v3v7IY2pXiBa5JqzfhD6SpFLqA4rffJE+ZrrGDyIthPcoAbV7
XUKxXRMk8rC5KZt3nh8lrRCJ8+pcDpwwqW2S75TwgYrXoXug8CJnolRBw0/dhZL3jbxqsczN1xGG
Mb2dGTrlx5lFoI6F57Sl85bpLqdd7gY8PgpBqbTZCrxE1gMKXXVTB8U24Jgnijyz+ROMwKwpaqsT
ku9rUGmZ81ivPp8ve9EOmNUOF6qHaYkEHemeA5hIs+H0a+5mjtCxTtvx5NxBFFyzEqrLjHpOEi50
0dfuYQtx1hvvhwwltp30pcUJA6HkR05mik4Md48Z/57tWLv9YeceVGehSp/x3eallXoWllQPHpic
uwzC0AinAbQfa7cUYej42joxsE2WyKgAtBLv48mgR5cbe9XmH7QPMefKkDZ8asRBmF6kZAEKjbzP
V/KjYJtBw2dC23CMClcuNKAvyl0Kj4WdOJs44e9XyZ7rGH8YjsTCc2nVuUpYxXodo7YllrN4t3UE
ELBsG2mLd+GVkCmebscskciAHMlrwGM6MwbhyNEtUk9DosNVgKJKzFNLxZ6dEoT2otbli5HgilU0
8C4EcjSa9nXD3VvmpFTqgwEh8uSB/tz5oBjZov1gwF1yds5+ctUpuMe53jFDQpgjFrhD7JSiWOv5
GV9UF496stx5c5CVFzTRn1je7Of9azIt29+ZyWYfy8em/sOCgUVY1A+fiT75V24htcZs1+4RoE8e
/CijTqU4Z7smqSXvrz/MtVLQxLU/jQF1tW1x0zYurNswLA33CcKmZkOWdUfPbj+Ld1bO/kVuKwaX
fkaHwhyb+TpK0f/fnaGSPnnqLx8B3hk0vOcRP9X5kuZnA+8mhEZMdVMbYR59fIOmBxrOsb+4V2D6
YYTHuI1GAHl4M8dYHPUUizH3ILvKHJAIZDQ71V3N3zGxpb56TwCkN7zzZsZPuhRfvPYNOGF/IwgB
xOVx+MtFqShA4nO2+Nk6GHtUkiE33xcTEytS1afxQBHdVCRu2Brh1+4ODsVwbn/v4fPsYWnrShLg
qODM9ZcQ5nbaegG/3ck5mAzdAP8VU14jaSsdxu7AaNMWOOf+kZln+aoVW5TS865/qlG4KsPy/odX
mldKnpvK71628hOELuzeNfH55/w3IUFAtJ0hPXPao0IQlURZTohVugI1/jB3NlLmITUgweuzn7Pr
aj1UQjlEHORLRd8U0fhwX5og1udbJUGhZNn7NPo5LK56Nh0rL5MNPYTzMD0FyJbOWjkc3KYsse2l
FsBRKhfMr00E8RIY3EkQP38M+Butu0MyPu/dYJf8LkpmZbohCroqILBWvGapRVgb7nIVBeVtbZtX
IYGpPP3mW3wUyVygIw5NCoSOxvX961JfCz5JNLQfjzgKtxpRPIYmekLTTn5NB4euUh02oT7TBrUC
hZshdOKOChVauHgRxqJgMSA8AoBUWd3JtOTCyHxw+eaMo/CApGcMEvEmZuo+cgQ6kywkTkOR4ua4
4HqQo7wMFYgTkYxOuolnXgdBoNl+JW7wmbml0BZziCjs6r9/d5f0Nh1jW3mIt2Hfj38KqppKjVS2
UDouosPxcqrE+ZxrzdrcOSgME6MP7SB2oZJzNNEx0hI7evWSWqbINoWF01Tw7+y2MIrz5TmmCM6Y
0mkf0wdEz+EVjZIIKZCgdYUs5BC8v7NT9/yNDdzQ7L9d/8cg0kswgk/ynZIv4i/QSjfuVM4mTfD8
twJJhEQslW+CbJLuQ3GcznOPGa9JRUNolv3kxbLGQsltyRaxKw4Uhp7xiC5lnPV9PgFktHzd0Fec
3XkL7pjWM65VWYAWPeJJ6NEW4vwrWbRajC+Pjs/7JIyAA4Qs48j1IFQ4jseuaRdD9ea5WvmOeK7+
vbJRMrh7OVVQ7gH/LzBE5YSQ6Gj5rrm3vUYh2XdyK2O9nRkks3tPT6grLg9mWRXiSGm99LnddGop
yLnN93WM0OTZyN2mBrTOiS2rg4DqwfXOraSZoZVTFRvb1AEQ2v7x+E4dTjxKre0AlcZdZw0Udusf
lrxnM0RkVdRTNL8bF6sMNVp6nl4PJ/IJhqVX5ZUXj9dqvbLt2QJ2N1GSEpfwPgbcSjRkqTNmq1fi
ss9MQB99RmVPZF0uZrcsGa0jopn4jKUYvw3ElMCHwy5DToKUu2s9CYWkqXH0+ddxxS1k3C8alpnD
pwN9KyI8gaA5jWIXAcWbtNzUzKrL5oobi2kZk07YzoQn8WOZdSIBaZIpUI9iofW9TLFLTEu26pQ9
u1yKpqvCG1dtVKso1gRtxDTrHLR8sPr8QYGCGIdMdlChrBZ1cMpCGgcYTU/Wccqyn6qorKa37C/5
38o7XD9Zf77Y/DurpmeyWpv5GU0lRTa7hmVRLXnbRihleXXGdA515JvfiviiAzAIwMURu+sBCMb4
M2h/CNj698BFmYRwjruv48+hO98eT9jhu/WtSQ/KcyMN6x8c48KFJT+Gjh5TmhULshjTsSszd8q3
aMoKeyIsP8GGwvhcUjRsRgNcBEqovSnMi66B2KZKXHSVUsapUrZEKuTYOIeSaoEh9cKsXvBGALaz
ENAeYjcCwxtYYb1u2nvhwWCk4psuJ7q0LsRa3YvWRyNjaESurdfQagRNG5KBqVw1OgMifOls1fik
JNmuM/FbxgA35RZDu/WWDbcpDoJ2NliUJCZZ61Jj7JDvNh3poOa1nglOWOItZOsdUbyoG5WAW24W
bG2i+grifOucGfh5JhCeHCtraqBisF5nHn5RhrnnQiOtFlQjCpFc7SP8hFNkX/lwWLC+9HnjN8hD
AQEIZaCmNTSMObAMLSWECcSyZeDnsz+I08R9nChaV93pAlRPljVXCgeiCnj4LaoqtDqX5AZ0U5gI
aKTcNgkMZzi1i1y91MKrPnbUKaJBqrv2ISvdtUFZpMDYw4fGsve4tOMJbJ7TdUIwoDd9NdzI1GMD
To7NaZHUfoMEWeJhqoTcXu4QM/02NxbnfWHWV5HCB4Sm6iGFctzHFvtkRni/eq7gzmPcIblor8Py
8SwDOh/Elblr8mzLOVQLFBEP1hz6MFirA1T0lF7wi0rX48nLOs7zb8tBRDeE+1jgEX4KbDuk1QCn
Xz/ft8xa10LhPbmIYIp2y9nb8ummRZ5o6g2OBBhvPaq+pNJfxmt8QCdpNPNYm/xA4VcC5/oOR37B
M0yu4c+OhZKyhBtgToJQ7PnV9GpT8Dc1m9p822lML7g19ygvmL/cfGY6W2TquGWIy5tqpWXUGTkO
NfRn9NpdY07EX7cRv09S0BroNVA9lZ5XVpJGIB8J9rOp4Oea02IsqVhMnSbYf1Ti0NrfQ0noaTfk
rbRoy8Bk36kZWKsOmg5UHPbQOCs94fgK2cMOC2vMNAc2hYW7NGk018a4sjoy9YpL6gHwe9oWbOY+
ajEeTC0EWgPHfaVIKSIsFqzUpT3axAjOyHzuXWYT0ZMolMoahjH1ZSuHe/aCQcMdCn82Fho/q0Zg
ajvWZriVlcMA5AL+LD6TX2IV8vRUQ1kV5U69YzTrE9PO/nDNcFYkgez8jlQXiF+P1z6I+TUhSOqH
DuuRUdrH0/oM9AYdpt6q/qlS0XCEA24m/E3mmNAfwc1izxAlsOgMgCGr3dILREv5Vl4Ds0eGfZjU
NeLM8AslRdmuc1J9Vmdzp5X0qijaj81i1SpwIFzQFZlabxt/M/9ky44TANQ+OrCy4VRJBJOgs1Kc
+s3XAlDUAXUIj0Xu+kVTm30hD5Y3ivU5g1RNrl2MrdYh29KoWSV2OX2OVU/ddK8JWolIXVIcX0Ce
9y7w7ZMbbPJ/N+Nprlo3MwUys7J2gjZRlqJqZ88/WmSsCqjWknNPum2qgkRNoHyaOZxiecQa/D+S
qAg4YpMRB8sUYhd+HUZ/HnJTvRy6FBAnlFoIK9xO06sLFlXBfBjK2d+7ITFzU5/inqamuO7Fa7KP
WHPeYNXRzJIcSmz50n96B+sxyzIdGLMRA3uBaDGlw5gu9NLwu8whXglSgzbgG+LEhDpnErhHCuUg
TfcTzWP0awmLfygVbAjD8pdiovBrKy1Ki6ycVNW75AM6U4NFFMYv5oeZ/P3K08hB39u//EoE12NT
U/DaE6sgM0aFUf7D4PXzXZobHunDHbSDt1mZOeDfMM4Wh6EbR3YgQWw1QOY5r2z0uiX3y2FwCY95
yNhXGZS3rpAtTTyatTKGZh6Y0gmyScZkiWw/O41QyN83BItLI+cG5Y5+jSv6Ek/ubvD7s6QVI4cL
xqAyHjADclXxiz+k2YyNmavWr6WiycPiYCz0KAtTauE0DlaYj6Xmv0KcvY5AG+tcEhiprHuvUfH1
MqVZcvEBaltKw4N9jvVe4gnMCg8kITmpDdmXQo/Kmy1/ARaB5FLoy+RUYPcaFUAScu/a5do9dMsI
KIRCAmv/r5gznvsvbJJ7LdIrCrVvvCGDGpNvUmxF8cpAk5lKFLJrRSHdHX8JrwfLr+lcJCcRYi1c
o2tlsILcRDLGg2QiqVCqnY1t3xyxNRzaJweYp5unSueOmYbdq551gaG06uFhNDiEyRyZWufcPQ+f
ncdph0Fd/la0Sn5/eeJwKQp49jE0lF7KDtuyztdx+RqIqbZOjce4pp9flblU2XsX2Mf1QWLicMKn
mbpHwcFcZL6Hf/Sj5K5nLUTxwbbPg4azajfATYENeIvG8vSlMWAEmqMDl3qnA2mfJLU5Y0xpwBFE
maqEUieJ72m7Dq0S2jvhA5qXm1orTlUfvseE0s5jCQBq2gPsiEgRnibnt/dvXCxtiWuQZpMoh6yt
Ijnlw6cbHyUxgSVkDB80BdIf4h/jnraXEBc1EPEtNeh+8FI/D/b+D/Zn1MJd/NGr90UQZHMxLyR8
tOuconJXF3qiSW9uGCjM+YIRhomtMypy0qzqNulxiCJkGxFUMZWxn9gTaeEgw5j0UGtWq1byHS3g
kEIFIeMHWZH6KbftXgyZYYDorouR1dn++xvOGfWgKMMHkov5wP8UFwnlZ/R9MGmWfK0I7fBj2L0A
jgJAFnQoYVonr77ib9nCH+yzli1UcYf7Tv0go/dXBO+ItBm466dYNyfAqm6G8d3oJkgRYCLAiChj
iyCZAKi1QqV3pJYiPMByjlEbbbiyBDeTuIsVQS0cDLj5Dc0VzCZn5ZzY97FsSMTVYU6yyiG4OAG/
ZMURmOObK8BDiFl4wbsJ7eyEXY/KbIEj/qWJfzRHCrJQFuzPZZRF5dPS69hItT/uCu3hBajeDSK6
yKRLcWZYmnyKLG0U/aBB8b+N/ZDa/ef4IxywVkBunu5NMeaXGpkNJn4AT2w9lSJnNJyhx3uwMyun
jDyO/Sb3LV/IIRQnxwwj2JMwMpH2tMrrZMurljq2uknee2Ih5SqjkWh8MxElrdHKOA2DBm+fi2Ys
ktai/m7XYlhbnNxH0Fv/VNy6kBny00iWAt9JI4LKDjjJa+wtXY49OGraIH3gCAILPpx46Pbmv9v+
iwJ8vP+y1DhrZOUn7BvAfaD7dQLh5f6iB5tmXnZnhd/4uAwyYtfKEZRwuxFAzFLSAeY5eJBVMsQw
+yB21p7cEkRckd8D2kThbPGs1k3EMvG+i9uizsS1UFwYx/qyqfOoS2zv7mjr3A4iFZ9GBIczgPXM
1tBgQAd3cXiDLniB2H4QJWS5cfLYLXlMgRtnVtheLjpqHuW9u5cBvxp4Vj8jjkcqIfAzUerfHDff
JzOjbg80U4FN2HNPTf//u69Ws+Cb11ZfsZTkbtfqJJVES2sdIWuhPVH/jOMhxxmg0xBgRbOQkGjB
o0GSQodqfylJDECL9ecyoT70Ql/8WCdJ0DI9Ajsh6RWQlLplQd0dFayK+/hDop10b0wrCj5ZIOpk
fXT0n5K7ReUZ6A6Rds3RUsyOK/gwylrEytReDTrqs02E6i9mKeAmiKwARq9BjNblJQUAnMf/9Z7u
9gzTv+p1O0uB+Z1HA0/RjLuBJgd0u9SihL2FoT+ME/ie+kplFh2tmgIbRWSjX/O/zjB2l1Xrn6rX
7Ar3dADI+UlfD1OKzAG8F7UZ16kcHH0huScD9PXhtl4aNqsOPks5rClQC4sWPLXIWykIgwb+E44X
cGCvdVp2945NWo23qzy1R8Uf93UY1qvBTRfampi4eGa74MT3MTBmLHf0K2R3oTWSsGbOrnhE6cFq
sp7ojL70IZTlNyHp3w+dDMDMIGR2PyjaeqJQmAamHzXxCi0/QKjFG0jagTPyfRTTpRrbcirZcQe8
+tl2/pj8is0GqehWcX0MwkJbksIz0ROt7lZL4aBU69heFL0k5kcc0b9bLCS53ByhrbWMbCSd/xVw
8YWwNypUBZlOo2PIPG3xMIzSVPpFSghsTyJDHTEanjyjqhEqhqzXWbQJzAeCyMqpVBbKDVeKIIQZ
Hcs06NUr4spFsLW5xmXvyc8WTV5phcOYbZ3y0NttifqaYAmpo+BQMLzIGLQGh7BVoLRVqohmKCgD
LGchw74c9VIJYrHkueYyQD1GNOwWedyDHRNbqS/vUqfH8ENf7wgJyNm+YICKHe2okGsnqSuhFKbW
mlLNeF82f9V/5tH0hGjC0CEZtGnvzHKsmYtlpqUfBKQz8XGSLQ0oEQdv2ZL6oJRoPTBv2d9Gw0bu
OZw5JnT5m8BTr5RMpOhRTODlpw5UAmnz5EbNzF+hGa6NrW8DmIVZCMr/YP3xMdE3mXVwaMhS1rKi
paYPf35kzsC6Kqwduph8oRT0RzwLH1ajsDIffGNnwFTHtHlvyZ7pyoxptDWuM6aJw8TZemI2bRg0
Fezi4bhR8BaiYunO5NQwhtL78r7WGcm2351N1xo8shW2KposPifRHIYWe3iBWLrGwFegEEtii3WE
9SEkKccNBg2KaxwiKm2cMXZHA2eIld4PVbbui6ucDIZcdt0YQRN8cclSywIsHLNZH9Md5lqLkLAF
b4gEnOEu8AjNm+8u3MjaVco93upxJDbdp8OPbDtGL/SQazPV1EylWl6PiSSdcOBpCWKNmhUOGDkX
Y+QjH/N5GouQTDUvCbbx0+xoLYVQZwF/MYtemAyQukz9Yku1IxPERHm6Xv+X3ZZxUNcI3CQop5bv
VWmtVwYz7xXxCQCtylEGyehpP3D8rPu95ddrYQTxPX4om8NTLYLAy/pbYd064JoH9pXTNz0i4Uh9
qOc31lJkYLaBSb5YS1p/ujbIQ7pektZIBeTiG2hla6vZNfO1Jg4N5SYx2BCPmilkHQJk70MmN6Xz
gcYXKoXePZXIS+l+iFvQXFwUFKEqn3FUXwJHaC23IUlNkiZnx/PN5LKJ4Nxrm1m4MGRUt4prRF7U
d7lCjKJEqk+8bmxieOe0KO0oCQOX/rb2LPkNZ6/Q+QEv8ZDcfW9khBWVIj9rZj+eoSQaAogCMgxc
16M3f9an6RLWWaOIhMPRq1BCpdjbedOeCqhAs4x42dfCDjteuWVm0ZJV8956ZrC2hdOloXbCriB1
5+CrlvZW96P3ZA9ozN/XD0IxOQ7SVerBK7y+gmqgj+YZe1qfQcmDgZmFFoujr5mojYSlf/+HMvws
EW15/I3vx4Y+/eV4fEIE2gKSNZnebgDAm7BgkAQ6+CIxo7SJjoJl1kQmw8R0sbe+mFP60Eb3Rp0h
6L4mJhgsJADDuHNZPRlSKi2lHnSbwZCfUD/wNwu+iKZ9yVMDv1A6U46qprxegcYyATgvJIKLETai
KRBTR/miwd8tgO8vAQTyN8tK6EdrCo0png1RUD8MXTJ3FlvD8paw/8Tt0vYLSe1o+r7oF/Px6UPw
HZO9WBiTcQ6+deOCECfPoefYmRnBM3NR57hR3e2UrwV9wsmL6VpYkrG9dGOPOjsx51jOHmRlznUF
j9VyFMx9WUlhRqvx5G+BYi8Va/uMxQArv0CmLkO0DGCegjyJMWO93gSt1M+oQ1lS2xCCntyNSUuG
qVNJT9b7bxKoD1oY1SHgKRIEorV9R8BYtImjEoSMOOqIbgY0dmsn0xmmU7wqJFSQo3WR4WNzHt5n
uSyexU7uITKQbz0HxM84LReJyxzsWp5+UqrG6xAwYNqkYfAWH3mdGLVHAvk99ltnp0DHJrRXbWY8
M+l45O8cvJLgsTkWXkGKG/OW53GsDNSmpSf33ycbqN9P38C7I8b4xOr1eAWt5eXZnZNfETqIy0ad
rVTg+XO3/YtJqUARb97bo9f4n24xJE3Ggwn3QMtkIn3kJ6n9hoGF5Qom0uvQgSVwm8hxj6q9AxT7
jDy2GACMXFK2xJyy8B1AbRshqMDkevIXttjKxsmMcqkb4s3bd6gzi3d5M45v63Xx2zdwjEsiAbHN
niS9dDOj4pFbMSzOKKS1lEMBUdp8Z5anW/6f/okFAwc2MlV9XIQ13GV5qsve3gn4y/LZa0IoK/R9
YO5jtyKaqxkGEXGzx22S9PF6tWx3ZkvtR3aHTyNtRiOMV4uLaC2EJ540yByAKDZNZVMmctzc8Flf
KXBjBZYvtqkHi+JjA7WUJvJ4ytXepa9dtWLek6vqXC/yVX4BusWH5Ay9w+h/7aTPAMoIL0Ry3Y5B
BFhdNb1HvedasHjI11JJNOA9CN1N+0O+s94KDaYeWJjCGAjgtpJAKDSCmZzEK8NeN73j5B4BC2Ko
8IdB2YrTLynBBVIul1G1WAE6BVbyjmgYMHKJiYtvEhnJRJ/dIeSR35zNuc4IMNPp95j23HOS8Uw0
2aeME30WvIVpibPHGP4Hy5Ie1em7rR9U7MIPFhb/PE6EipC3+tps76I8vvNw7GStINSTXmnnvuYK
PsYZCl7ehXCea4qPVB0gxylpuxwhr9rZRZmVgGHHVlH91C7wI+JeIBUz5brByI87ilO9o+ThLSOu
KoRZJTJUC3IE/ShyO50YmohrJuPhoDgufHB71epSssl/jZeE/cg26TlbHVTn0biT8CnFIAIuZjla
IFgqrU9apJeBR3QB8ZTZ1cvIBdrLnyQ9ptByE1MS5zCO3FO10/f25n4uDkRDMHTIX4iVjafsLTce
ytQm7qjuahUw9KXJ2GcgE0oWp2CmsWIz92tEO76jcUsQmawug5sMJgwUOoeLPbyG1PrKzEZR8Uk9
SiokWXbI9vFN2JC8rrvGVe5O5EAt0oct1NlIGo3DL6C/6dbRioo0ZCm/YSUzv0ePDJUUzvT5SrWk
CWheRxJWZgiUe6SYRnmO12u56t/ekRbmNNrA8kggj6I0jgBL8tSpyl6Ptxz0NVt74a/VfFt4oAul
tFDmXLzAjoLsDlGbtOgjoefpOvIn1Fh+WxDEMHveXW33IzuRLPeVOTZ0/vVKEphkuTDLTdwIbclz
kmqZmzwAqXWA0FXGtyun6KMbnnFPARA98H3XcI8H7dii2yCS4Hkj2RMELX93DahlHtoaRNapAPPE
HB9Hd4AcuR60G5NsEPawtcnpYPZ99xG9hwb9CQsIfWOdCA0cokKWmkGRwLa52GF8VXyz9nM014Yk
mluHncMG9UP3SjVWAZ3HG4b9ZRIGnhcI1B8aXtAfAIfcs61EYIATI6pQMhuSWiU+6qlZiLqskgok
PI8eBMEMKi7y8LrxXOFdvn633NBuDL8e+7x6nxVmSFRg26+3Z5phZjuizx4Q7LRghwyDRvrsh/Dl
Ay6a7+UydcH1N4bbUiRiLNQLhqXzNzi3RGDWTFTfQoCeqB3f+Epc5KbmVKg815klraHt3Qs1Zl9A
qN2NGkJ8J//wygnd1jOaSvlJbmNvfANGCxv5IwnreQj7wK5uhapBeuLBhD9C6AG3cOtuSN69L40G
YSpECwaK6ihU+tJyz31QixL4NHZSu9p6+GzJGatfsvucwsK6WYVY4E7uunQLuSUL+qbv6GLw1aBa
tpCaAzNX/8gEZjE1DvveYvrnucNPs34cu4VkAVrqiWAc7Exlt81swbRq2mozmxdR6/vZt3fUKCoJ
fK7hhy/XGfdVevtjwxwV34XGSu9w2Jl7E8CmDdZjiHxbJzAkaUlSV8MfsbU33u3xJMYbX1gfQ2xK
8+8C4jzkQRqAqNijnwdU4//EzQ/M0rZIqUiIdVFnDppOhHerapye7zMGP6Al5HZwwmo6kWvbpsod
/pZQXs0rwtHoZJOjdcSwbxma2IN96TPg+uT2rIjr71r9huWCmp4OcfEyiXfYe7SI38BStIAK/heA
bHYZ1H3I9HLLgMk0bHKJtIG64tqxtoQjPbVIz2dgH3aPywNSDcDCP2SuR++eX0+5lsWOOe46f9Cn
Rdj0ypyY6k33Q7Tl3EwhYqSLiA5DNmqRUx9EcVzzZmSPBoQWFSGmIzwx1dBMQ/pucUjPsw4dtZJt
E/fqMHDtDYRP+60lb9qxSV/Ya5mCFFgjFNszbKGRLg3tvs3TWK8XvdOtEZZ47zHGXPQsBZe+vEDZ
rWDFzfLpYu32wa4K+qXx8PdLgP3jQKkCHMYiTYmCzzGmEN6o33xgxmlhX0Yjjz/ksxT0GnvhF9h1
FfD/H3nVSPFSd1MX7UbngCO4crBaL+gMZfsFD/eO1FGd35n76NP9ZfuMI273Ehib+Z95Ot7sCVzL
oKD5LrLYU/ZKOyALeZgjrsTlhedsqjrBp/8jAo9DQvUFfuoijWg7PQCLhmpNlSgW4T0nV4D9/FXT
Cy8kLA/46U9fmXES69kXzJzgTLSIorRAAQLupXdPQv4ST0mI1EJuiVj2DNQLmFtvxtBMxhpDReaP
3qj9BXZmacPJTCnC80xSUxWaHcYZwkyJLI9m0uGGJLT2tlR8xXok1kmus584MP8yFJaxKux1n4Qs
jXs+ooaoMdtrl9MzmFsiQEJf9pAfdMZ1By/18M+BHW1rg08gJie6Bn/IXym4cJTZhO4OkZeyQgng
S6FX94jvf0L92y5t3BqvxF1UkZo+wgXDdTduT9LnF/bNBBa4ae4ipIx8Zt2b1Dwqs04Ky2JEylTJ
NXFBX6/S6Qw9a+25nGaqqh1sydZfapHRaFtbrmD6b3w2L3OPAB3gFTMzQsKRwfovexfKrisUQl1p
lPSzxj0czC8nZsNUs/k1aDiEhsHog5aADhBIO7kXHPVS3R92EsHXGJj54ARYvwmhsipxcJf21wAS
jkL9H58vh0L8Ds2zGZtX27Uo3DGMey024D7bGQNe9aDK2nDxu77oZMiDvE6tgpqgzvIDj5Fp/veV
1kRhw9xwxeBAOp0QqbTQx1uw8OdbFEMEmm09waRvHoNxu/eKF/IZsHUWLANNy6G9M5px1gR1OO0k
vTdzaa9foFHd+WvXQssYg92th5iK7drr+7UDE4Mp+UBXwSOJOYBbZVInXlrUpB/Zo50xRs/vDSxZ
AMIRi88d6VsPAjC+G1ldD6OLZyHQ5N2Fx0+rj0TNrNLTFw6Ok5IeVyPWDTB5jKX8MWpBrKm8iFDI
YokujI9rRUVosASXRdk1bCPTAFScvR7wkMHdnHxEoAfh170BeMFu58azKmlGnpUEHHbR4DW76GCM
5UB/bdUEXvtRgeMURvSeFjQv0t0RpCUrfNT5CcphwrP8oFA0PQfa+L3oYM5NpkurxNo3Tx4ZIUIO
cImPeiUxL+NCiDvFW+a8pX+/sCJ05UbJ04pKpdSg2TnbzEJmpfpRp3CZq2jDNppgKtwngJKJV9Gw
a78X25UsdQ1t541GZHIhdTAMVQo9Kw9jHNJ8e3V32Z8VYHuhfFa8ljKc05jU0V3tC82/V3Fknsuz
Ga3vyZ428ls12KyePxbCKZem5WNgu1kLCX6u8pGXyr4liNlIIlWHakEbp6+JOtcu4dRvASLd+jY1
Dm9AG/HHqST6WCGqmx/MAHy7Y1ynwBBFTTf+TpJeIzvNwcDidcD0/iABD9BD6Nhu0ieT0qt1GCOm
nxKNzzUoEYjvYxuVN3MDTVp8oyj/alGqF2MimIENsaBZcuLEKaySG4mXBmlkY8BDbJfzXSA24Z4c
JYQbd+0MIq9i4jzrPCott73/Mm+XzgNNXWKHvmswW7BeFhbhDb6ujcBZ8YT8u+Ml8Cc7IVitSzJP
yqiRQviZES6J5O043WCgwTHHFOnlNs0mF71YJ+AjDMEcNnizcepVlvpcgvh2NIMd3mfUji+yu96C
NBQ5oykc21U0sRYD2JQTXNVf+PZOXBGRYYOMLaLt95PaKGQ7ALlCaLnkgwzUiczHYK71GisrTHmq
KWcqHzAbOBY+6MBK+9yZDOYZKZKR6bfsopk77XlC1y7k/VROCL7GYm3SLuScKa6St7TNf9gDTqeC
V8rM496QVC4gsnDdXtpLfwR48TQruKKrk15r0/fmAXFlxquGCetjbSrun4Sjvhc9H9T9J8+CoG/G
yBZz9ujL3u7QLTA0CKDGTPlkro0/qZWc7W6iSSDHulvWqqhxYNGN0whjpJ/uRJRw2l8aFTOeq1te
qMUNhpXC7LjaKF8f79ENkjSPPDGOmu6AV3nGR9Iqok8cbmDs/2xcXbqyM7aSm5Sc7IPbMSgmIPxZ
agSdpCTtzd3sQ1ZGQ9Hg3xgsSvWveiQMXAjQHRe07M8mhAFc1igMtwG1bBS8M+HD0yKnZTVgilF0
LeqaEkJrB3gZingm67U4dEcrhViXZtiM0AIayTpaiq0SWxcCjpTuJfHajex+rfnP4VMdJDri8p4f
DC4khhLDsHXWFEiYjXxtEDrjTwTH+8CSQ3Ol38Q9wLVcYp+mfMs3+LjLiKAZEN9tzuOaTZKpeUq6
ZVMaopMMNM8IX+zEo6GFdw11mMxv6Gyc+8NNYk1CLboD/jHHWYit7If5NlvLH/soDIjkdvRQG39p
my/4OonWEX8Eb7NHkhoeobshodqwKkpWfXKrMzO6HXb7PPkcsIvCSNyqFR7w6ZTUU3r91o/ruGuw
jQt38s8nsfnb3Jmf2v6MksY3Cjt/GV2MORx5FkZC8BdOtw+fPRqRpSNjcOysYSelfLwBZ9GMDNxq
VmtSnxz41c6yPUlPx8G1JnmMdfNeJrUEQ8JsBTyR0uQP2jRcwYJGZvRo5jk67WEmgbfixtrqtEmm
vbiiUUADWluI7GQzl1nuZLq2F68GRgYZ65eBreJVBMK0iHyfp/yySNb3WYQOR3zv1kzE8IbC65D2
3cZB+5pvBwjMXIePSuvc0PR6H7DnuGOJrcHRNdbFdGqZ/Xc8oaHV6dQY/WWNsBz1290SCT2oNtH+
wj5MCC3tzlnn2cH3msX2BX+HEHH6fiz/OXD8ORgDl5DCb0PB1onIeFtwO0moloktOqb+zjm/87/o
dRVKPvQaow9BOVWNgbk4h6nIQFmuTybKyNpZ2oLFOwfM06v9w1GVFwaUi+s0o5WPvUzSH9bpv1PF
IXQQf3DFgylI/9RHE9k1BbYmbJ2BgBZd+kD3prFwc5auLJ7JUlfZ1egDfrppM5nx78iB5V4VxF7T
JEkuZz+tZrivOdiRXxWA9eNIajfLPaNxbeHZS4UKMKJaM9syuzqDFtNo6lQslGutdfm6scPGYqhl
95nTMQdAVQaIN8c2Hw8GiCSG8DRGInE2YzR8ooObQvQipaUw4MyfUKDxIGwGy/UBaIvDj6oJyFVU
wwh1KQrqGdKOQrhBut14lhmWuEMmXumKZd66NWAKH+mtImUqP4coshNKszx6EKqGtHfcHbfeHdmR
IeacHf+gDBxs0kwITTcL6/0jNBM8kLNjga+bxjpL+GaPUroqhUl6COim59m+/VUgVvIM/7srmhQV
2eI07nMb9D++foNzurEV1CmUPbgmX90w891vfxq93PI6v+ict1HXzPhS0UT4v8QvFUrsHW2xiMb9
LpuHNzZ6S2MvpXzzPwnXECCNY2zuQ8j39cvu0hW2edFzU8PWIT8JjVZjknWXH+brtZKb8RuEZXKG
BC6aOLX8bwJk5ScFUO4Jb7/J5rCW1qKgXVU+u9iHg4ICH6wfzgO5CRwgAXpScxjXRAtwWVuaXk7P
/nUSTrNViv73HCV7ObUHfRLi7+HYshjM2ZksAZ1G1b5hCwmY8yMYh7ofI3mzgNNNr6plZAHmaXBw
lnV3oN4DyJRDICNNmlRa6vGLSwBQbTadmN1+6/2k7NWYV0bN+nngw7HasblLNr2JjTMO77PW7sh/
yoXmch9NQHNzyWeiP/exckjOQZgCRFznAkA8ZohmH2sdC8JK9WPYoEktGBPhwADM4b7jcVBXXtDt
lEgOwYhGwqdke+uSuiA94WWJbgEznqPGeRC0qV0DVxXaV+XanxpnM6gUhqz6tq4pPbUK1Csd1ZDN
TDhNTe6Lu0PUxTivKYh9USDBZg7BcOilN2U7K+FjJmpSmbONKAPVhKMswsuzurprFH+kZBfBizdU
spJ7gohcikgHcH22Q+Y6K7NUI12xnPTfsiXFmmsS6kD4qyLyhNZcl+E23hs82tgh+L6Prg9oKkKp
tCMEM8r7PUi/vHxHc2OVJwzDCb3hk19eBOhuR09pebPCqry5CcA0PWKQdsQYZCu2U0t3EhOV/GMB
tKYjYrftk68spu8GshU/YSuguwVO0+4Z0SOMNw35bsFjAourLQNly5TCVCyFzpkwENqMYLDFhtc/
raEBWrAsxxPqYrl22GaTyH2ASLurbm5UimRFQW0eMwL0g0H9+79alGYBcGa31+VlbfcUVntKNPa2
f0BxztYTGSUaiVBISzsFVlL8NZfQx4Y85+idpVVNggvTvljH+W2raJfm7gw4thrGpUPX8DIIjyTx
Q3q5Eul8qxMAkq5/nTF2H0WbummTtTGjvOva4huaXSt03tn5vBLbysrD5um5Z0h7QwArl3VWe8CL
G6imF8GIr9XnDphqYAFdGn7gq1Ect9zOWvvlxOejYz9yNiBt3GLZkKMwrrHl8bH0HR78qLe4R+z5
yyiSr0YmC1f6NgA1MccGDMr/xu0qF1E7tgAq9x5xki3aaeQE2x7PZyaADhYKcgwEgjTnXeo03DKM
mjUVBZZXj3XtmyLqzOE/s1loawZsfa81CaZ1cusB6qcMSf1RWEEBWqdZsoLve5s0AwbChAcMXJjM
1yqJcGIOSRnftLw+vweBA01kDbXZ/Ud4SarPPGRpTqY2OEjKiCt74zM+w1Pm/eHEuGjG1kmuJs7g
BH6lCy3gD2q+7Bi6/xZo4K6uPvuTHgR8kAXtggi/cPt5I798D+jL4vL/SLjR8cmhAKCLU+no59QG
EvmVuZwlUHbeJwzW3cq08qrzqyTspPCTHP05WiC3ohPIcsj2nb0oxHLmiGiSDAZYS64B5RQQGa6D
HC7Y0AY2a+XifD1/1Elp8Bt9QcfcqojHwtQ5fnAa0ouH7vhFbERWqi2Edo7TKr1zl0Ulzv3T1t9p
fU4EmyMD6KeB4B6is3IpHv1I85E81yB1LL2MxOnpRRjLo1YAAJcaSenW6LMTHSEMaM7c5PiUgyGB
wh7xhjeoLISbDuhjxUpH8Qz6DgbhVwVSnWEBrcSru6Flvl24vPMVEPIHJq6gOFyZrP9QbnMaNl2h
7UaSkp7MINYFLDQ6IMFa8SPlxwckicyRG8joWjV7FFmtIB6Zdn7mMd6jkSFuFPTUbvpw95fT3vDt
DMeJ7u0746Ch8X8YBQCak9pTMSjUYa7pzxpciavgOcAMpJlvtlJtuSDiCx3n/GNxP9BwHyzyZLDi
yD55Qf25EbPdwZimj6nYEuC9B+0lvIqPx/6tqi0E9CuCp1Xp/CLbbdkjR/lnYAohl2KGk8118FAm
XFXl3ZNNUD8OL70GDplb2KP6m90Zkr4wrQ0p/oP/NxMkMMfzvaNik3Dgnz78UElffNoYqAzpG9YQ
DhcVW9XanaZQ/guFBHrJDcZRZFw+Px4SP2KcHadTEs4AzI6R5pik6qfQITyaF+w6QhSwXp8Gjugt
/wjsVHhyYom0B4rjM7Dy/iee2b586ucVmC3FuXmW4g4aVl4CrdGyby4NmSjltMuFnSuccJDwm/5t
27w0tWBdtaR9dDiXiuV11YrilgjRMLekfROooutsugWqTJwIifF4rC6JIe30PTLf1zPmX9kycaj0
ws8E2P1ejk5dO9BYCB7YZZG8jX6c67CzzgXw5tDgF8P8wn9W6QbkbYKIxcrL4Cnao8qUNIsoxYDj
ZAapgjN7uCeoeBAYpateHbFGha8TbZAZEgLiZbU7CWHbyocxgoz5f6S/51NnMZ9i3ftFfxNMC6Qv
A4zEqMXt4qgdHp5USM1BDzT68vMwmUqJ1MGT3PaC1mgDpXy6zu2FPQblVWKZRqEEA0avZ0UjtfzK
0s/NhqL6bUR67OQWelYkjFoNV2aejtmgcSgjMQMrXra9skWg0v5QhYjJiIZ1Uscsa/CAa/0br27h
HIvoxu9U5zmSQemkRXfhnrYdzHPd3t1JbxpEXckfEBeMM0/YhZ/HVz0UjdeoWqVeDwB8giwNblbW
rxGge1fzm0EgkaVdCXBiV6P7rc8sICwi8YiIJ2we0e3/4UDMZRN0gK4ls3XOjaFFLwGOLAPJc7wE
B2Mol7cRLmVzotm829zPwJ4seGQoRsnOpS3URheoacpLtJ3mT2M3JJkVkoP4h1iq3cYtwVjSocU1
q7/COyt3Lq2FLM91UsIiDhbOctyQCxy2eAyACCsjUQzYhUvU0eD4woWjT80z16BuZ6XLaXWOKmWe
g1QCY3cj7s+cRbAyBpCci/w7Ir/aoFJJ69szo/JxNJVLp8pcKMqJ5XumZfZ+Kpyx5hf1y3ml4eUi
QjkZqfl1zatN/HP7IqEFHM/lbsgFoxbDlF/DXu3CNE20lETcFWPdJWv87PNnNda4/xromoSqFx31
vpeXlpH6Q8ofQ6Quu4H4YBQIS3iCCghBSagWhOTHnpMIcXP9Jdn1WvmT26+to8ZBZAVN/DZ/12zu
g9CdPRKi/1iKGpLhz0pP51P2RwI6hjZEUltLI1oAZESXcZKKDgApOPxf3JlWzOZqlKx+uiVkzJYX
75ngJxjttA60h5Reuy3yVf7w1sCduhSFblEUr5+cblKVJE4vbFJEeJZozhM+WrbGmig3EQ4FW5Np
4UFXWK6CyelskYcQQHC2appnLbQEFtMc11XALUjQBcQn97bL69IF2Xd5CBQGbFQujMSwU7mggrFe
2f6JJJ9nKas+nbLo4WXg9sOTc9ASylN21082EePu1P/oK9Br0ed/4aVlrrdHclravjvaT0e2TUbK
C7djeiO0dWpP1LIZ5Pu34g8XsJfW2CiIZqriVdU5uBTABigIUkQ4R4o2CR17G7qRHmHyk36Z3q64
AEJPc7AhA8+j75ETKnu11tDAv8l7CV43v6NkhwvLj+nCepPGuIiofQQV9RGd775pgPDnWHtlgGm4
C6AGm0qju3fkK7GrTrCFyxyeh47dqWaQRbhu6wTsPA3gfKAhkTvJ3zlS0SQEqw2obHGa6JLfswnv
6q1wHrzPULod2yRIwWx02WEkyvj1bPuLNbVwTjkf0i9ajxfak3WcTwWa4+bgqHkCm9BIMJ6Y+PhW
eiPE+3SUR2k7PcrDfP/HqJQuLNPrNXoc+MLA3VVFEqWF/J17q1Jtlf4zpRRTR0DrJBEH/dvl28Lr
tzCBP1mFBBua6QRCmwCQF760UeJamTI44WHt6NJHBoNAY0F3MfQvECfm2z3mwL6XnpKJTH8GjsJt
4ZkVXhjYIIJJFO1hLbVecjCgTF31gJmxhrwnf0/EadA/NLrFkznYIiknqZ6rjJmqPmjvnvAcEuSj
PW4+P3iT6OTbPZz3Y8tleq0JCAASFPeQ7aYaU9ZeTyNdRS9Rl4nxGjiAmDYiN9Ihi+jfHuiYiQ7z
0EHDQKgwXU1w6xU6PWnEPkadzMyEQ7/JqQO+3nRpBwXpwzDDmjOAEwDDT5nfaOpdR2bDUKe8Iqle
uf9RJKFLb0qbcZSrnJtHp77fkOWycYW3FZG4ZT6b6lJBhmFliGenAwYKeCFEFcyjGWvFBaliusfK
nVt3Gp5qemYHN3HSKfWQ74Qk8eg8DI+utNAlx9upTvok8bXwR5tV7GmP69jEls6OkrxeIWCuXZgQ
0YPIHxq2U7PM6AgyzpcBdvQeWTyrHGj/HKL6yCnaOQUl8i5tWFWid0G7knqZgy9XB02J6topb9CU
ZsE2q4BQ7BBNavddtGO6m4KL3pEiJBHQOH4YmCPw6Phq8TZ14SexDYzOUZobdlz5fNcaYMbOE957
qoOliBvHOV9a+Ab83VNKmOQPHhfugPvYgNZ77RQDeb4GGeOyBw6lHwYwVSt9gtSB9xcn9Sbj0m11
mK7shL5OHECssLpQujP+QApbjnFepFhA52IsLG1oU/9ORrh4M+mbQxbA8SE5sSFYhcnAyMOTlCOz
AMv2YagHo4c6Tbl0Yor9ZuW93Ql9DdR4trKUTocH9/xPsMRqN0fDauNVr/Ly7duYY481lqYFlK35
sR8DkXBwdKLsicCLyg8oWcFSupuOOxZ2x700nIZsikqHE4rA+CjKHofO1hkgXGLYb/viviW9Qoio
3EpS+7wcoEU25pZURwZYkN99nHnZr23ZLBhGocxH+j1B0zrfqT4d7sG2YgFATSU8TWJPiezVi1+M
5fhhkxuC6z2TveLmnr0c7Fj/nju8lxAXBXAmvejPoADs66iV01sDBjKIp0HfLilpLV/WyY+n38kb
t4ArQqg+hm3vkzCg4AKjFYmh3iK/y0H30A6WkMlSdrbTdmk0jXcwloZ9/piUCHPaRWzMeogXKNyL
swXSEJhkbvxEc3DHFd2dwINkwn2o7qC49V7EzkNWz9kVQTD6yjMgB+My+oMBplALR56qorLFOzc0
VRQs0Kk1405D3kV/SLCAy0O0+CtGjyhN4+SRLabkAmkqu9VvRiFaFXrjlWKDztzH/nixwcJ47SkM
l+tLl2R8TEH2HrvukmO9/B5G+wjXwklL5EpGBKsVhb+8rIxDsohh1LZahjXgMZPRQ6W/cxHW4hY6
UbE7v5xDdW2eabouCYuzp3sib7TBhK3AArGjmfKpiDKkWJsgS+4GqSbWzQBrtk+DSv3HQKTo570g
Es69j6hKqzP/ii/nN2/WeOS0SnaPOxJJpcyBLVKubNN7twdoARZNxX4uQWx5/sux/xkVV7LFjnHL
kpGkmewQjIioGKAezvYPLrYoeGSnq+BmpkkSMIDUI92muIOsjrYYWPhL1GvJ1jxFZ9AS0R9DrIWI
sb0AaEUQz2xyQfJQidmItcPpZxphLyqHlNWEg/iCIK+riIaPBpvtoHvbnkRoGDVO3pq16qWQ58/c
burog+QHt8bJu/yRwO70jy5g9JSJdSuiXGKuudCVGSYV07xdbpVHn8Gb4otPLGjY/cvigehj6hiy
3snWTMxHNqbUVlcLRZhWoblHd5Aid5nteUNBWMVRCRhswrNgsvkTxfj5k8KU0eKAAIuGb2Db6ljf
0gV05i0J0t3AJDG6z6pFGzxJ0UsxR+ekAcC+kw48vPSBZUbMP2rzWCC7+Yz3q9eCAS6KfLGPeTl7
Jh0HM9FRXN1ZIE3JSG8YQ/9q8qGPQ7Lu4PLRkjzhPlX3lM/pCmIG8nilosq94SgNaRVgxYm2QOmE
wr95ISUsx4uJUuimO5NTDbbYdzOQLrJSMYx0C9Qgmz6sAPf+I1BesoQFuaj1WAWTzCpp7zZKzKOi
9rLwpZKJF5BDaDYgcJ9eFIwcrEr/9JpfMKFMj/GSRIhtQ3jgyykIF9nycKBwBtJ6RNQsa4jSG6gl
e/jee6qA5HcStpVpktcWMMI2roVkHY5BetJGcH/R3L5EFc/OvhtINhVf45hb0FVXy1DTNUer6qvk
G2MTpST9oVsi7Wp1dsXvZCOPltd+xypHK/f/8cvrv4PL8z7lA8AMIT545HUWlDbE4WMMYnmoJZ0/
0hDdSCFai1EfW8O8Qp5BaZ6OsfdWkhhYWpTzDZeO6JQu/9yaQh9HBUEcGbkGTKm/1I2MAUm0xvI9
MyFAJ9mntYTnm2GX688+t5PvrCQZT/U7K1iw2muu5+OtvErvA+fz2iNTPevkpdk6rmKvHnuC/OoH
ktinXZ7e4Dul9zRlVZ8g0yQJ/3soBmKGewCUuzo9lMsJeKk7YP3uu1IjKMOXYR79HbOWSkWu8rp5
Iy9I06aGJ/pUUGqO9LsuRqcYh3rcT7oZd8mKDwEIh+U9EUk17ngEM932dwWu4xYtKlH9uc7rt9Wd
/9Wwe5/ZXNLfQjvL4lwOrHvqsM37cj3N37AmTqYdAZqv2ZvQH7O25Rg+6tGqYfU0A7GMhum9nGjZ
Lz05F1cyfSN8d4iVKpau4eePy6KG7YCuC8jBaLD3c9xxlQ5M2LlkFuAPDka8bi8nVBIS1MZMp5Rq
SzUcV1Fdkc4BmVgAvj3E15rXNzBjgM164BJIoYvK39Y3vm2F4mZaZabQpXq8nJTBwwRfW1oGL1xn
/gCSoe/lvM0D1uNwaOy/SqquceFlLu8U5//3/lGo+ozZNqqSsrhGciI53wKAcsCBB4z5u/pJHoO9
NpGxHY97nyeCDJUiBmnsHarvIJ+0QGx0m1PJyP6EY+wiY2NHMH6c9PstQC/s/mgJhWFE2zgb//y9
2dEUQ9GXZ29UJ/HMSjm3U4x/QBduH2/0jr0cseHdFNPnlR2UWjGvI2KgFWdgaUTzo1DlxPuUNNQy
Fcby08ejNmjZm1MrahTrs1+aTETKrQWMQ9zIdcEOpLHBQw9m8Z8Tp5ErRl+fmvXfq/ro5WeHpbY2
9tWU4ilRJDO5MADWMdy5zKvHRsIzwGz6/x2YImQ7h5QqLFUAj19YJfXjhh7ebfPxQH1rHycbQq8B
u/IFQWgTbro881aGAnwv2LrgEREgQhaWRzrIO0BNOyERgZEoiasO0uO1NdDtE1frHLI+pJIPYBsP
W+LeWfKGMiB9JAkZUrl+YZZu+ny5Avb5p/e5KGOpuMN7axOgN57kSiLPBCh1S/y+NJRBUC3KVh4F
usXrMU/lo5H4KgT2BFG+fpkNYt6eJacI2lxyhqWILnCK2y4OjdS9IpnQgKK8HsZ6cs3LlMP1K2Ja
Xmx6SUysat66oFtWYOcNQHnTPdJA9DvNBvkvZkCRawK87388t3UX3H1XBh6iW70jQReFEdthyfPX
FYOxkpV40gdSepwH+UOx3L4ZyB7ZQ+FNx9WiGraTDiomJOuTOPZbkDW2pslRguEkdCeq06SaQ81M
C1wp6a7QfQO1294Whw880EW+AqskmNX8/kIIevBK04E9geCBsyL6vAIgLLemjjjeei4QhVNqvF8e
GBO8A7WoeXhpt6FBwi6/U6OMAsikyQLkfixAsAsikqgOAiWjY+E1g9NoqHy9kidFeFGWLCso11Ln
XWf2kdZwxsk52T+9JMFxSpWNnxUg1MNa9hSQjErmEkFH11yWxPL1Hx6BykLZ1kqfGqGUKv7j4g/S
dulFsJuaaR0O/LH23kKXcLVbMNNLqKXsvUIhMyXt8U2efc2sco2sERKWXxargWahGfxGLmSLBuCQ
UAM8a7XS+MHpGcPipfJV7YTBfvzyeZ0CEeJzq9OjTElQtnHqFPjrYNpo5yfLVSP3gbzDMX5EKSgi
DujgeDT05VP7exfGXVUnTC9ZicjaJwdgra9zZSmpbBxdznzFObyqQczlqTSkQ5/ibdRYi/YhD8uJ
WeeTu3e/C+4gst+ki6WoBZaHjaGv0sID7Hhe1v9JeRUbG5Igu1g/rAozblbmTKz3kTk2NT6hXXAz
K/h+zB08BjxXfZxaVI9heUgf0FZ2r1MEfchs+VYGd0rG5FsVekZLHiCF+FTpyJqj0CFDU9jLope6
VAOi0nN14AEpJJwbp0MuStZH8tlUdZplOS2f1aS3cJ3Vc5y/Ld51rg5YMifMz4xai7BIKXQQFi0t
015QeaN8lWG04o0timFOFPVao5LJeAGqy9gob8NOqaNgcuC2tYGrj1J9bfHdRIpCXIsv6GDEpkxa
arko+oM+0wMrIeZhZ4hg1zvCPHTGFx8P4096avtNVG8bg0/5scY9EGkWCsYP650KF0j4OhGD+eZD
Ce67XIkrYuQ6vWvywm0SDsQQ+AqeWAypZibatEL4B7cYYNoJf2cyrGRKCZrMvbgwNpvUNQI6FZfF
940JwFgRGftzdad9sRKSY3Q1mhlWL2ALlQHdNGv5oITdK6bFTOQC5MYI2m/4j2Jwurpwvl2C4Ybk
RgNQ58nArdhrikjEUG3PXoG0NGMxmV2fRSv2Wym3/LrGKPaXFcKo3ZjxMy31oWqdXh6G//PsE8bL
moI40zRUeIJ6FnU0qasx3/Mr4xELC+YsXihr7w+CUd7uVGkc4L60pC5Xvs1DYwxMPGxv3Vh3m2Bp
lvwGg8Di14O1gXnEQ9xeL9WvkToEW+XbjPvL63bjhvPM6/M2R6UB4pHQyiMG/7heqC0JIOfHtZku
53a6nwk4uaA32yMtGHLHvzmqSah3zQyeDcw9CdLTv1d6c14uQbs4i4Rl4v1xPvd2PV/vv20ldkN5
fWoxXRoog8qXLOY3eYX0uasNpjywezAFX1QyUe8LUEFNPDc09t9SXnYFbb0PBKfhSCY6EX/529Nc
JAwu1plLV3ukoJzznoK70ScF1/pI0yfaVrK84wxGrrp8K+1RGP7HNxfFCzzSfAnsvJ+fir3D1yXO
yeQuxivs3LWgAV9+G4dd7KytmVY6vrTFWIoYw+gl6UwDLT/gvAWo6tAJoDwWvYim66xXFNgcHxzg
Cwe9zxVDawdwkGNH0ytcuz49E3eFYqb688DFPsitYpAYKZeNbCsPOdIhltR6x8/KY5Y8WDNxUMYv
xZ66aImeWdu2cvS7c8IISptyKTrU07SW9Qdos0M+BxP0CmoDPPcGX3azoo2cneb44sbuoDcwDgRF
kWiDo6JSJ5go6mzdkw4iiqIDhXG9NDHG4W98kDDJZLC12YHBorje17MJCxIFyOQSLvISyftowQJn
jA+P5RHz9a5VjeF255o7Ud30LKT4tKHC9QBg6S7TelOEUNLa9vE05z6iX8H3LUU5jzNtnyjCW5vV
g/RF7QPQJVczAfwNtescydALHyWcpon55y6FqmKJpk9UNf/AwsK6efH97DrLvIZ9yDwnoszum8Jt
Bpx8hm1ASEoN3T9OEEjYHkzzd/1Bx2fztSMoI74s8azd3Q9DSXYCVKHZ8kpoyRuhpkkphjdHmW58
2glF+Av/hxssOD6aXoqM7G8+X3qow9E2sMk6H5Yq/F8m2YFCEZMZAU0+RGDWvnICkJbLoL8Qvshe
rdtFVg0QKMxJRJy/56+BB+CJgav1d/0cwE0T2EcCEKllL9b5OuVwjwvv89dng9FQLQkaWkA0wfYc
FOTYw5OPzfNpUn9Ghk3EFZqxxHViiWMlCjGDDTZZU8zBOqFXzSAiKo9QLTXikYFTTZbnyIAjKgSb
0cta/mv8Dg66pYeLy81xZsraqVOYAXbRjMv6jRftNGCt9ZHtCD7De6rjD3l66i2wcrOyTDAAKOPI
XZE/OLPVsPtI/dngVf9IMim54TJ5dHKdkr2YJ7gsvh9WWPWf9a+GKUDg9yEC/GFdswmtrlUv0FFV
1Z3UKUOqOIXlK+D4ElBDzUd5FCNYSeL/2vh6Ah3V4Bl0mh3+DgEIgd4EIYqa64bsJTkf0ZSRN4o/
jU1xZeWEOBEKBUsuo5ZvA30ky7txlwt01NPtkQEMx2rX18rglGSg9akkRuJr7vpEU+ANy6OD1Z6R
rECCyBMNM1ILW5aosU5+2bk67oaozSchoGgL3TtXczXdgm0poPJS5SXeDp3N6pdEZxdJ7ltEkduE
5llb1YqhaOKhC9Bnupr0tpHQvjL++9x35gzINS+8R6d43juAeDYorgXlfAmRH3lS5r0zG9vgA0sv
X4kYj4Zh8Gq9AqNnuiW7NRheh77QV5mgc/vN3b/AFT6Q/0SotlnaPn6ydIo8azYbabY6KqiRdeAd
qaRI+ajWDrSfNXOTpPoinGIdlvGWUJy9JD6+fFpN+AFh2kJtrHx2trYECyDNIOAByUfIO8AM2SZs
ppxwxVeUS09KNsQZhvRDz5iBi2SMeXQ23Birgu40YA7DBKWAKQX1zb/AV8uRpfqmsioWDYMjt5CF
+RaAchOPkoz1v2Cr7mwQn8fbscxOz0QuH8UNXoSlKUa8gcNgAd+1SExPttPFKiKx5c3HBihe/Sxa
34lVLuwF0oqFenxCuyBaxsi1utR+5OKcu5DHCm/jyrTS3m5Ta0ODIRLxGftsn6G/I2+8oh995ch2
ZMwAYCdFDPXvx1bMKXbV3XrOLGt89K6WlL3CRB2ESGozXJquIyP/v1Ceo/TZVmxr+d8xk8HtqzfW
vC+l64X7uvXFCeUnWdafKC4t8JZYWS0Nm0XQpu/dV2n5gXGqLTpAZHVOpy8DOvWq1pPX3ybjGKQr
VN2Gm/8B7hUP7zHW4oF8Hlu64l1iL13926C35xSzHkCut2XtwiJSS6vNslOcUt1SK0+oLOxoQ0Mf
Tf0bwlWdZ+hmoCLle2tTYRIIk8P/Yp/72v56wXVlNFoi/hy/tyU+uMHbErC14RfiKMqlvtW3zShB
gaekgmwxtJPO+cH0ZDbNzGaNMhUbBrJl+4crpW8omljaevxj5uEQjs4YYOvb2EMEeWDhbv1dzmWC
v11Tt6Hlrr64DPPYDMTvEUPpgEtzLp7DxWP5uTgW9RI4Q7TzCtstL9VsHFWW/QaqKsV+5xdePwnU
cycH3KxCh9OibJ1N3IK9yBp+EOZPKRuiBTZahZZEok37A4D6z5BBzPtlnDVjqOMXGzFL0tfGaWWy
3cT2D0geP2UtEfWGKv4KpMM7vYf5bN+2dvLqbt6BIznBhQdZ0PepmmYnUcDHaSRLAce6WNDXZaEE
DSY/1THikIqUXwWulGzyQbF2jiMiJLj+8g8FTHaygJj1OOF/5YW5p8aWk3k761E3r/4De73D81GD
TX/RRpdxfbZ6Fe8xJPunVDdMNp4emP8ldKdihx4JJBkwwCfrnvOBpUNMcquILo3nZPAefN5jG0N+
fNdzF1gMHj9TnHn72jWpECNqqt1M6TfVPNabHZ+hNjtnfTbZ3JfeYaJW5jbldtLkWnayZOz6eCqY
e6Km3fCzpyqvrLZqK4PBtZ0BxZpRGRlRa05dkP2E+7/qgqxQGIPiQFE0qrBsDhpKRXZxurH0D0DP
h3wi03WMrtRUkuhAfRiXIB0lsI9zC0ZgVVybuSI/hXfXlif2pUiufECJwr4q8yMU3tsvKzbQ4kkl
uUghivNlwivlYGhij2NVG4lG3UuiNXapO6NVopfKRhjHmo9xPAZdCqXZPJvx1o9sg9xxnnchZ8Lu
mUPqwfDkVEpKABBbPw4eN/+yXXwCNgrd+dKHxL6h2R8mYP65YnKLfPZO35y9YwRXwPAhKOqqNWWF
dVkNxRGNEZomjXzdB7WyiD5D3URScRn82RJTtDxpgT/b5VFIqSeUK5ttY6JwV5aadQB6zy13edNT
sgRl6yOhmiGJ0CsebhDnFoYhdiTi5+xzFNiaAHAk6IKVzcTNh3WJZv3Cb7CCRG9Mw9QDSLr7/F8N
qG6s2UA+LZtDtHF8oPmdx705cOsA6wCLoVt+54nZosB7Ga5bv8UNDjThHUrQ7+gxd7YWQFN4vRQj
aZ991WTmSDHDbTwXCfbLGMahR5abGmcgEDb9PlmVycFlu36HsPPiMjgpWNb7Cy9TyL1RdMbmPmWH
pHBWTLjU2nzjhpqtq9BVe45XxntvZUJaQ2VjcCMIfMrpkNeV9i0pNBlJGhm6AzkMy0y+aOmlEX1z
kHRdUCET7/NPGF9tHGzYjCIloj/YFwK2pU7SlFTL7Lhl6dCwBd0cBm6vs6elDfBhuE3rSwJkP/TQ
6FnLe4Ttwx6S/S6sphovuaO7RDVL70hhF4r1eFcJ/SZsAYs7piRk/8E3ColTv1Wg1Fp/l7LWQTAM
H0dpTLyVvkafuwuTzCFVB/FAfWkBJxD2Tqlm02A8uXfewakwJ3YMiSLv8KzaCMm2U2UvTGKByhSj
xDa9QRJBKAuEknAbaGLC4xItZRe4eKOPMEcKwQPou0tqiODtVlziBX3hKoONTgOfR8vWPODgN4ll
uFTYqHlaDd/e8r/zt9wUfQ6z4c30oPzqffrcHHy16rxRGOWvYoNWTvsJI5aqsqiAoGRZznIvL0aU
w/LvcCK+EFejFIKIFQk71enb8YbPRNGAyoLBX6rtqsTV9jHje+r/Rt1kIkK2alCeB3Il9qOjD8io
oEyKmErY3SakOK/7k22PFLP3ZwfC+y63WGKDAnrZjfjzYr+u9rQT2+58+fB8An3DI+/U0kbp/9uT
zX+BWbal3o+Bj8IGmAHnTXby3aaYbYDG62+xVkLdT9t+KdHvEhTHx1fNVdtEyML7okiOPGykypAm
3T6aXRL11d+1uDW28lEkbVwQR6srNTlW/+6y23Xn97bb4FXmJL3QxhSQkVKqDltqyzZUmWbvY3y9
IokJ/GlAx7qlTUZCyP4d5dQWKjIwpZjyt/Ah6Dn7EZZUzYCUgNUzGkBjMOqa04DudprHZ0sNOwOF
E5Zn/b+hWQ74zvmMfqHHigJEk+4Woxn6XFkTi7pupjxHXAbXlZS3Q8eI9gQyHXYS3SQyJh+zOX0K
ogQhgblzp4zsIwAjZLFld18PjclVIoESKI3SX4KOwTaKMunbLE4C0WSDuNqMzPhvCF0rZ8QzT8CN
E3uF2QnRINk5zDvimE5ACcH1mqKcAV2GZ9rHHUWkD5cx1VOClIgAybWGWVvqqpPdkEwXP5dtX32z
ZRzw/rqco2h39tSmTYCWsZ2WX6eaKAaJhkackizyCnH8mj3pnL1vm1woRDSPzu4vWaXqjYjZfpK/
Nzk6Ru9rzStZDALOXXwycmdZl14QZss2bVjUhC0DFS6ces8ORA+J2V5gVyNAyLrSDKQwKSreXXrC
gukgToemQ7miIHqsNBF4bBhlsaH8EU4bsxU8HMA9j699ZoLoVdz3GkRcqICkDKbbC1bJwrx1arqr
7Ir2YZMvmG/ZA4Xz7wRLTpd8SC1fRc70DFAltqDTfdrsZC2jNvkmOK11o1iokoHEhpxhrU5Jdt1j
A+zlKLSsnyukrhPqpCW354j5sKvqRlplABAu4zOx3OcKKe4N7KBgCYZPpyxK8lKrwXrX95ukSb36
RgAn1Tk8urie44Hh1YrLKmFOZBxqpd/TJwYulRf0SrLQbbIVF2Q8X/XdtDee6A4MtYqR0WV0useC
+GKs9QrQlt/VJg9phCCb4pTq8dUjamIW+aqhDj6l+YQ1bT1ldcO8FEYOQfWZ+Tyd/yqOB/BzDEQp
7ExaRdU4VkqbomApdx1y0e8911SRNju5R8xICc6LoY0Twz8bNw2VibYgZcAdBc3tequKVjER3KQY
dlHspstOabU6Mk8ISM9Hb4aliEwIt3qJ7QRMG5HhIagDsEUoN9K16hgwme4aZJ22M3rNAMDUYXQ+
qpUWUK0vh/aMJOlPGxYBOBdT/y2ebiq8rsk1XBn/C7dtJitgJDdk0CHf6GayUDLjhFpe5Vf54kzH
wg+++esPd3TzFykQOtoItuTrdlB4GBJQvP4/mTJM5EVChFJSHReg4C1qAxrXWRv/RFgz7SEARUrM
8QvMxwQwHbzzPoymtgG8JSb0YZ3H1NkDE7FsV0X/72iw8AhiTWW5q8zgvDYs1WOfszF+217AQ3Wc
4wiE6HpOry+jSkF5zBoTrKcD+yAHv1BpySxGTyS4TF4CMaCwMRIu/0JhQ7NwvfvYI2ij5VKbStNT
UCgKle78z7x1NBFGf6pIbmoo38G667OiNeGLe/qm962qPgYMr0LlqLhcZ9ZcUWaBabL7OBkU14n8
vwrCL0s0bxyZ5gBP2rF/E8DBHW5Vpue5CqoUJMkz4fUoL1AH5qa1ulGisFltVCQwyXcOInL5fhjS
OUTNMCkAmcoqy507HayYi6OLT2t3GpCNyyrfE6Xb7+nh28CnaEQMewbfgE9rZ0F6JUNONOoEQyP5
bYC9YcjzHhR4VFoclZntkECHEh4ues4gympaFfdNGbqOu994x6fT4eNTtDrdsj2W0VsVoDvTkyT3
gwxEopD1viTmLjMXSPoNfvBxJLtomyuOHjJ5VRUDPSDLzg7vhgHNe74PoN6Z4DF53x09gw0Mb9GY
Mb6g91+Cn5JJGztPHxPjZ3XmzAna4FOEBrRc4cj9h3gJUQAEuvM3tbk9ncxTjNHmzC5bHMih5KGx
knZwFHIeyPjU5Avno5L70b8ZnhzhnVyb/a1TDdjQU6/ZGYWExqhcFFRHkoyFdN/VNQaXZB11Dwtn
oOW3pb9Ku1U6v0WoM5JfEVdcK8xAJEzyEIXvcVEWwr324H8F15MZGKag9dHOZfcCE3gQaSKxJRAS
yPsV7jSBUe5Meec7lTcsVKPhHWHlt8Zui6pygkniwBmb3AyD19GCOiqDEoSjEtJM3PFBZoYhrQ9b
YjSq0YnK9EAnuaN50W5C8w0gEZDUDYKUDpiBoj/DYJeQySB0gm8exr/l+W4CKFTTPmH9tHZIsR0r
wS2ovnybgO7fEusbM+SAu0QiJA1acPh5NkdA9vyVte9kCbyedrJKIrkkhrakgMVIt0x4ozhf3igD
rh9A4P1TwBQ4ilIsRhF15q14kKkVhWfRr0as8pzZleIHp0nidjmnvQc6GNU0t0+ZejAaKDlNN4kz
R477+wP27JB5psiOqqH+1QCAeNNmbEDFCVEWNHYhiCazjuq0fh0xoqwxA8V5Ku8zxJGrmUlcC6qr
NTVtxwnZP29pqMLZSDSh/HbJajBo5PSvA8/y8pOO2r0wDCxcZHS4Pixq0ubOLPH6v42O7XV1SaIy
rHwHPKqQHtlogRwXpRwuZwADaN8qrrLwU9FycJlC3DkrlCsvS1hsQKZR12qwbhNC0plRDLLtRY1I
EztYki9tT+/lOs8DqBAKmMERiDruRm9zXy/na3wkBUY8FsNZy9yRELQ3gyHD2w1Hjak4n8k1AROF
WJgBa+K2oGMyIYs1HIWkbuUFgUuxL4jHDL53B4xLp2czg3dcleGhsvoK0NFHaG9X7uNCugVRPx3h
er/4StT1rMIfS3J8h+FjxC4cSlHWFmCgT8A8KSEDbKfqG84Lwua3C0t9qGncXFhsQ+oOSOFZbI0l
TW55oG8ziItG//f3oatQ/R0GkBsfaatYVLN+hO0SGPUuMffGHBccITVr2XT5uUzb7xR/KFZNH5se
/AEwmq7ujpKYw6CPZOTTP0qkbwwENXVrYHtq3APRKegS3jLKhCofxkCvuGEUYigWIK3zwBEtw5Yv
OL61f49+Rzwm5sj8whmkUjjayu3M5kdY/ZtlA3pVaDyPVQqYNqh/UEe1tHwdwhTU+ZvmWte02Y/6
iqmQgvG6q/NIS1GWEPYvvysWV/C7e9tNJdGAThZN7s5BSlRWatGIDtS72VdgNQv7o2uyv+udgsO0
eRW5n9RufPFJx1kj4tggVvBRQ9lecslpwbS+B/jQVvysPYczTTXbI2vB4icBCcj3Rv78wp2ESllw
XLvRPQxj7fcoCXbFgnFy4o4vN2oiodtIHbLO3yWJ/BNP3oNYYJKf2ZQ7/6pD76sdj609ZqFfeNIJ
BeSgdNJioxM2Hnu9HnRcphJgJcpi2hBj146sWrVIzd4X5/r84y/zJN+vEidZzCnxBJBGyoxlg2Hu
siJoHeNzWJMqVMtgn3HwU1180kIQeMpNdOGSXhJY2PDB3zmWH/4m3NkfBE8yIqsSCi4KOOxe8zMu
mVq1+puBRMNvw2ns9irV/lO6wwuQNZQheb2uFZbrEvAiymGl5WJNv4Jkvs/iUv7Fv9CzhiwvDniq
dddmTr/+YPY4gYmQLdeFnws8g7N4hwMx0zYFBUXM1djLzW1JdYQ9IHZan1J3jCBLsVBO0EXMrcPV
UaKDKAPexVFVyHmw7H8AU7K9KfwoTqfnCCh2Ja3r8BbzEyBv+unvhpYxr/v15M6mAKG3p0L1DEr/
IJPxJ6/6sRRxt8gWUjzfwJ9Ei0cu4JK80Eo4lMARt/ATba0Qb4sX5DM6Mti+/UtbVD05uiYtelr6
hXll65qCsb4epJpPaoAU9Awtg9xlLOTRHFBNAtw+HqnO/1Sx9rk+Ha9GTMf2sXBYrTWRw/27ksdD
r27g5ImfpVfaLJ63X4cTof4FUdLts+LkLU2ZwaUIrROkb6TI4Nz0fZakEdLzXRukbtdKqSiM8Fh/
mcMtP1vhiUm1jOBsitlM4ToYTxkqlhg1KqaeNCrSwyo9bA6MMc0IoUXjnyTiq6XYvFx5dJy0/laE
vD3vY05NoLoG+uazRohVNPnJlwPnkYxPeRDEKX/MXD6CilMJ3hcNNjemUBJMTmcOWsXU4qvfz2My
Vzki1/QDBDEq7yWxehrEOGrmwyJ2s8DFVfI0yQWDD0t+MAFXt0m3JNLV1t9x7Cu/dsds4NFemJUk
GrWXnft1LXRZ3u3qJsWprXYSNVbZlLTrPMk/DikcDii+2c91kri9NGKxKLr4KyfgAqPN3rFK9DBy
2g6eBiGfEKJP7lDtvmNL0d1oXfr4EVUgmRWw0o+VTP+6ZVjThe/lCN8ursTFOmIJBu9G9jcFZe5y
G6vokq/lJs0s4KjaNasBfP/w2IH2sG5fNnY4EGmOvSellrMfzKgayAuq7DBTCLhxL7DLSySfYpED
i1EG+NwUv4b/HFMfTcia9NF7m7iq81yRvYqtc1l0UR3tnH9r/vtYd8rOdhEqLTmQNH5Yx3IJd1nr
yVCs65nWAWPfRYFL/GzKbya1eHNBkQFCAMQepPsp1zVSJm1uR2DyD4ycQMQkEcBFv9ajxuRMhL9J
fkrrJvMZoupMEOJmW2gJ+LjZkcMBWAdZ/WdY7FEaI7LVFS31qPC12ZyTek8dWFPlRdmCFdiYNB2O
vcjFPk4BS1weFm4JZ2O7ffQyRZdm7qSmUXA4X/BuNsSS6dA1amK0FjUJRDDHShDLXBAmwbhP2Zgv
ppkURJpKfLn7F3o26CjgfhTZV+iNGgu47HTVRcYpyfvZPX9n8XMKCosilQk/KpI4kQ4QMqVsn6qR
utBCz3e2EMZKsdH5AO0Vb4/r3POBX9/YbQN0uYTtb7cMSiMR5P0E0ESdYiwZoYLHDglHlBzv5FCM
UtcmCGfBTCGhCWSJV4u8kxKIrWTF7BvQLTEEyBrGRJvOTyYnjASIH9e8nitT8mPRg6qmrS60fTwN
HhEHYuXeFnHvRAUDx60o2GNNDYWWOIjdoyszc8XO2tkKsyi6Ipg9rNgGnydMJTwBTmBHRPfJ/fgP
9JlPSGPoO9b/8kVPQkLk8XXLAeexGH+cipaKJJGV/g/MMqC+2UrNXzwY6MHXHBgWWs1fBh19YRmP
u/hxKqprdUHe4OdK4mEN374OQSgrzDg/6IbO2dhkFBVVOJhrBfYN59V4WHRW93yC68bnSUE3DgaN
O2U6Zw7iEs2FYrCH5BOu0UPEZqXtKSzNsbDdNc4qVLilnKyDxGp0o1cBjfYjNX6hsJbNiHRpT3O4
VhnzNJIqOQecGFlnE/YITG2cvEYJfVSYFoRjlJpYCEUwB9q0irAViE1xmEgDpRhBhL/kPqP471hZ
+Jzfx9CkesXFiPNI92NXCJAe+XNut3ICbN9IZBK6hK2j/i18mDaUZ8VBZ09Uu0mxZKHpgJtuCDi0
D/j1RduQJrifskTWv1FDFmX9cE/k0l8GX1hNEuI0un63gc2QodnbAIppEFwGrv8D6D5x98EQQTAf
1NsTavse2fW0MtKUPb/pLkWwcZdeI0pspiBPyiED3AUC3/DsDY7WpqNCHYZTM/913N9DpnXDiIL8
sgZGwgXiO7GvcFGyExcX7/aSsCabq973rilS2gbttzuqtXqpBPTx9XT+ngGxLHHcNpTrdnlK9nHb
FOUfC1n/nZA5pKMRctvbXFbh+wuAx8GKarMHQHrnf5JMqlHmppEohDimLLUl0FPKrwNgXJchbiXU
oXiYQ0skaZNwHdhnfaTtC7b/ZLQsjfhj0Jy5mpdDkc2uv0hFoGzAkv0S6PmptzJILBTHSpID9d20
KQ0Tmb/l00bYmMM+JdeoxZvdL6zf/+SVQVDgS2YY2/TD9d9bYcXqCSKcMWTKWA37cpuYxC3q0Qg8
D7OXOMcn+HPY42mr+RXl/VwOw0C3qk1JZGltPHVevC19qwjVRTnGonmpCz3WeIcPG32KPL3AQ69C
efjC8g8ix+d0OK7BQlz6wJ+e2DTRBxOZtu5GyrPCT7c6z6sy5hD2aUVJe+rveNn08NFcrpvBhGt9
04p2pvJm48P9jVWnqjzdHSEBxy6Zd050hIW6cDShvuHWMP+IfhXYjy3Pi8sco4eCXhVUO/4kS3S+
i42inrBzhMF8TsHCyuW2fzfnqHpZGvk1mdDoOAhVnr6v6j45KM74XHTbTjqcrt0YM7Gu+01DdIeq
eylSUn5Ky73Nlk1MqQCTmB87klm5S0rjeEx2dvZ9bbxeFcPvoQH4C4MIKW0GEfP+aljqog89+Uev
TFV33VRm4D9JPQu9AlME8GRW6XJz4KdSwYi9kQ8F+sLivQL3iFrz1a/8AVODL1MgMgtu4ibkf0N+
2jJzEPS8prFqLzpEPLHKYzaemaTXmnM6wtfdb00NGLMqL8ICaGJvGrsJ4+SmSwiWqOLfWBRmR/3L
2m5cs6wtRa3ncd4OHw+kRafd/JsMYFDjK5JiBMfhM2P5z2qkq4xl82micW8ybR5Uz3lJOvAbnHnf
uT/999qXckU4jOUo3v6h8Ai7odZwO1tvaOq1jK1k3mjHHfI1dZ2VodId7LRwde0+GPiSNKAx773l
JrOjgXuHEEPCDRu4B78enG1Ff5RsMdH0IgLiBmC4fG7oZ6B0mEg7veSIhrnK+H2K+jmRgg33aJ1+
wM0FZY1XZ+cjPMFn+VIrwERgUwQpxsAEZVz72O4gvPV9NYmWS2EuhC7iqhG7avBH+zssREPb4FoK
indviqtvhIaDyLXXyDfX9d+BREUk/0tAobDsnO2ap2uZI7gtd/aGeFIElOz+3hNt+uRlYMQko25U
iCG/1+MT5Cf+Kqrqi25XjyZdqvZhod79tyVXnKeaHAT6I4d64yi/olB8AFjzP+H/al/fRx58uDOm
DcFGbvD42njOBErggvkKyzo/ljwTA5O3ERxNJaqZZc3cQtlJt7xojuzqNnBL2D/GhygLHDQ0dez5
rLIP9bG7p3ESI8l5UJNaw7qy8+9/8p3zfWu475m8rWLF+e1EMhPRMcIS3bnqM9Eyok1X6SBGE2r7
hcr5E9DswdJVOUklItj+L518jCpZkasvfX2WiVpBZq2aMmuP911F/xxA8kyda7R0pDP7OaLjCjvu
y84b2ErDJ3d89McFv1lfZlXEpAR8gNmbq0TEJuP//L17aLvR+t8QIH8ZsNCW6dJXHwPssK6ikaDS
YJGzqxj/0AN4jB70ddqfB8kbNLV94CGTGgtiIryG8deMNRaGLuvhlY3VlrZzuWanpj2XYl8x9S9k
vjlIxFPpKN8RNthKNmNIo1ADlul8iG5CxZYCYvjvIOYhCumI0527tKOxCC7ZnL+b2bQbAja/uCz8
L4+LxhjVdrl9qZx9wzkzBDCFi8zG2Rxz1z/suCM9kFSkiq+GptQ61rTihbJK8qz+562c0OV80dzI
TKwIiOS+LU0iCIxwiq+G9DCMg8IwQ1Spt3qW1Ok94/oASpwDLONw6EA0AZ9IFaEJZPeSPpU98qjj
/FIYkI0j2t+Q498LkI1WCb3FY5CY3i93WbhA1rZ4qTU50oehgAfDKRK7KUUVnmWlGEsX2sESS38t
nHkWUwFZCR9MNzkN2mYZr+yvsb2l9lfyKtr98glBfCj4eOoyPBUh1n8nPxXU//LY261DH4w3BOfo
rZb8ry+DhKH28+0+SJTJkcMo7VWaHvnUKsl0idJSfwEy4idbX57mS81Aex6BIYjtUBQR1KBrONSB
611FA/8bI3w9I90Jl+xpHyCXnE297X64cB1jhqvatJCvqYXDLa9OOMS1yW0WKsd8qeue65fF3Y60
BN2xsjJmKjmYXifsuVjwUxCtbrOU8a22hjE1m1SjAVAabnt8BMB3cZx4BjE0WuTUGLhpOUyn+VnK
SxKkPYftEgIzNmYTWK7mzvacJo9uNGOU2I1tYTg8ACGaf/qNdC6E/KNOc0OOE0h1BQSdzJiJnnwG
dStxL+UEqzC8+XtvORe162XAV7Ef5M4dj2rS2GzrwGIrW+DXnXe/uOWTAEX9vI6mZ0onYLLglNLK
3Q8UB27ccjnDMg5V/33P5gtAZ9Jaf3qhDZi0BuDdn3ttpcTahr7y01HZP+MAWOqmAcdtMzTeeUUc
M+Afurkw2381pAudVUc9l7aiFslNasvom8zGdBxScg5lFvkGZRMWROK7rsxhSlMH1moYK72vH03u
7UPn5sioYAWAXo6MYi8Y51Ffx36tlUNPRV000EDVHaLMX1Vd6bF3g7j7JHBRHLqTeApJNsYUzKes
BYUyBa5nce3MOyb/kC4r7yoHko+fpIJyMfIbr0AjcEtahdtMXPoez7aTrqGDEZIyLVtj0tWku7Nk
PUJ+7ikYhuHWduhkGriMePp1apRx1u+GLCTaJdmgyuCOeO/r4/am07PlEgFkt0mXsEd1aCTvxP0c
v1mKasPRt7qPjn8Co42qcEWYliPW0fPfhv3pPBBDxPsBL2MggCduLVvBckMFi/o9oZ+boOHSz/ST
4PEX+JLrom3ER2ihwVL963i2xFLmrQvIlubvw0aalRw873E62XJGnkYQwuWXll4r5I1RAp23AuAH
ePLU4fmmaYqMfyriDF6KTHvYcpySnSdr+8h3/deesbsEz18/0BDmyW5KMU22LnXjm2nuxEuD3ArF
q1GGUdcECHGRfgMlJP+Hju/3hz4H09mA4yxOnWdcA/kjqtezzApdjnqlGA9xBub9UAUMuyoy/PBA
3puu9oBmPyDVaJOXR/g/b8O77t7bgId9r7TvdeImxaU20U5bYP5RqKeZCm3AvZI3D4YbfsmnXZJq
/5D5EGvZ0qV03Mw+iLmObOgsTHEh9bPQaeyZuoZjHGr2NsUxX3OOaDm/cKxP1eKqv2P5pd+tbUPB
ioKU9P1RexPs4dUkfsXKDXRYDR3WcMHVgfVOc7Btse/RtWZvOdK+0WkY7cbVmyBmaCVUy81Vv6PD
DEuYME6I9xG1GjVon3lIZlmsNtfl//FQf0sO66XCeeORl/3vQUcGgH3LZAsXzYJXOgvESRfj6Z0A
ki7umegCJRoGS6xQLmmvV2aTN6SHihjBXBqHWsD899azfLNFWfm2xFiIZxdK80R2eaMn1M89kx41
mwQ8mhL/MCxUa19NcWcgfJSKugFbgSG2aEG4IbKyD+BlT3ePmCrU26mIF3AxDufwQHud76mKpjVa
YiKHOXx+FRy7f28SRA0aHmJFvEwEm0Aiovh1uZjzpsx3np6MObDtn4Y7HRA+GEtwtwUJR2pLWzRV
krRQNWvbDWIlaE6rpHXeR+lEiKBI5RarcQ2/O4i+mKHFsqmVI/3d9X945nL+kz59MX65YYYufaQX
7BLrHqgyv1EoJk0JSs+WUZ7fMar/G8OWsTwlMGxEtTQvX4jrJJ2sKPgZYf4BOY7MHQwCaFolojsy
8YXMO0efy8iHMu3QcVId4bBdnaI2m5XNpxW95cK56Po+fCjPtUcrarPPj31hLEeh+L8Q4FEBhpeD
TnGXs8wmu6XXxwssvV2+x4NCpy47JkAVkMJSTGX3tFH0jPGBLoe7KknZXmZdw9TFeMTX9Wc79Y0d
SeKfCQqBSc6rhxRpo0mRN2vf1CV+3j7aZLhqd/8pcrHgeO8HZrVEDud43eRhcLBc+72lBM9dODIP
ZYneyhxAsWMC3J+fzJMLJpQgE35gmugUR5d8hsje7N9WwGFtxa6Xdes2LaLrp7jMSLoeRdDpod8c
YA8OGbYKZVlC2Ze/JS9Xp4hVf/kubON973dOEthHW6gM6VJBuPx4C8ISYB9HlC0NAtyEn8bdfpHY
MwrPdvpEwAECKNpxlbrk7QJbV7raBSeDEC+ohTz2mncJ9vW6UZZHbvPGUWZ3qjQfhuM5BC6Qi8aV
9TCX1fwrDzdPTe5iMVJfTgyhUMiSoS9xHx13cS2lfb6uC3QCB+v+MRCTKhq2f84bHUpCJuSzA+Jj
iLrp6P3qexiyFmtH4D4ejy76jqNtOO656f7DuP2jqf76jyNUsnL9YdaaRM+csHUk3LDEJhy9/eeO
w3l05AuNsqa6TOFEl2y1zehZpiWpyyWL/IxijN2Eb1dh39eox0OIRVX+0MMu1GLqOpXyWE6HRSpv
dpBtiM9JQy7/vIUyGrdd7ZUV6V522jSCH9RBDx5O4nd9UZcdJzTw68iXZPwxJOK0MBD9WaO5xMWL
VXuAvEIQJ9GXOQYG9aFLeaL45J8jm9xu/zvh5Bky1Cj2z3wdWl5c+xQYWvMupufa9DBKUBsA7xSs
+SFWxJH/B4hmwF1ABe6G/ZzbhU2ukM/KhWPLMQ4OQoYcEPs94bp/IgKZS0rhoem2o2txo1L+raAP
24rXU6f5zXZga35sL1rIE0gBSDsnDaGNf2xIWF9YrIr2dpgdhFX+O166oM5+J3i4LyUalHFrhzqZ
KRLYLJPsUzoKDw09pf3s0tWFyfFtBWGTdX6ZfHuOauKX6YFmovh600HikqleJgeESk8SUzKNFTK+
LZJzly9D5zjxcvbPHrsz2c15JfuL57Qj49Tw2AOjTqwgbubRfQLlxJDoQMCC9jex5DRH0z37lXKX
3dQDOhYmW8l2gsdVtDmNdRoOaU8qOACILkStT6qqqGopAUDStXbasOyPfwY4unOn/ySG1HebBHYU
u8EsnwsuzQkFrXb/uWaJKBRPyd5bAj0HD1ojs7IgMrryvaBLwMayl8iyGMfNF4gcQQuwfUi3lwQj
5moJL6g1fBtnQxqemCL3T+Y8MPyp5niCfmaACFY/INaGXcTRSA3t0HWMsQ+V4dVYSBLw+KKlDMIi
8q2NJ5C4cQ50frKXvQpHakd8InpfO5O7sYiV+YOZDKs9XMAw7bKvnRersU+Nc/7y4uGaGuEDs1vh
yloRFl8vY7eP/K2Bq/S19VkR3iRkIw+2nCpWFtxKJN9GhHJkPoUS/UWx4sOJbwCnGRzFMqFJNobl
R8eqWotxKNLk0XthwqXvo+rv2jwDjOk9FQoADw7ONj0W0z29F66dD0lTFrRUNMSyf/s/UmacKANx
md/ptILmpsaQZRrd29YlQrEYpGSgPPkChrxxDowVW3Ka2nwBV2SoKUcflncY4xoPCft2PPL/eDmb
AoVAlXJBIUwk+j8bhTcv+W5QKVpwQiK7lTZYl3UVx862T3aRwqmNhPQ3oCsRCGkvVeVbysVoyYyj
fy82mYWxbu8zqrRIdJg5tXoLKsyegHKXpapSg/UqteURAwGrOqPnECi8INw22fyt/NjWjDCaN4ON
lJ3VT19q0+XRfuYWS4j1HSh0dLsLRb9+mXwda2nAV4KOhFe+ulcpr7Pu5I5WzNGod+MlCuH9xAjo
1aB4aPwy59cF0fwLO3rA/vHDwNz5STVOwU2M9ssgCuLaMl2UjRDbEqj37lJvA60znVoTxZZzgv1q
JJnoNT2OpMQRD564kEvg3hv5uI9LIYyWbf+5wydrSFtP8PKH1iLsxw0TSXNbRZyyNZz6j1wVR7VQ
LWg/9pYXZbqwowGwGPCcDMhSBwd5j0nAp1HrPykU8rn4yqdD0EWjvxIGM2CzREaEUcgTpEjefcWk
6IDDfJp7OWh82rHGRkdhxZOlrnDD5CPRcmApN2tCAa7wwYCqb3ile31ScajgOP7YoDyi+GOfrTwt
pQtmBd5J6WqyRsgNApMXdZMGgtkB7LSp+/xb9Wu6gg/QnncYX8QQfTZgBfUoWBppN6FmGfKcpSTH
F1PgOtmFl4n+vmCM/m1nraTC01nJKIDjK+cJfxXCKICAn2O6dyacSInSneztAffYT8QaoffXVJrs
tO3nbiVHo5bhH9LpDJwEPHeccDnux9wwl/1UnkKI2RCgxDyrlQZATxMmGb0d7qyWZmZNgJ2LAR6u
0/8+8wHvx+dLHWWSjyXYhlsSVIF8QQ3or7HRR9ZUxmFcUJUvoLmbU3cXiTS7zDZVG8wzYJG+f1cT
d6YWwxN9DgsrhMCevXSE1gBYkvTUQVmjKzLDpfo6nX9ySRN5LhpXIsB/hfVojjzVSMl+coVmRMo4
YAaarHlxjueQwwSS2u94u8IvZF4cVqDsEYTKEz6YkwGJ8Msjr4eDTPQF20IEl0n24xqSTTZbL84V
ynCTHH3FQfk3osBItS57zBUO4LHiep6mZvY5MZAG5mPfZPDKgPVNJ7sFBRh+w0cGOO4pUA9zflPY
OTKnugw1FCMFk1wDz/s0I9POsr85ljmwE2DaiAEUplUndsmDTuLY7uI6+BUfGIO7SZR90MMQt9Zj
si/gE8T5SQIhhNggLeiH3KjnPG9r/HxJdufr6Q+Y4tW7QWs64GMETu7QiqyBpytEb1HXrmQcH/bn
oxCAfpQyXokz6uL0ep+qATzyn2zCw7ix5B3M3XowmEKtlStyjB6eCWEWEZSe/TfS/CC21aKcfyad
nFjAtsupPRCRkdlnVfHie8ZvWeyMGQfJQMFtJig+sURz69yjkvKCOW5SIHbCI4y0SMiF9GXttFin
uCk3Lw/O8zJeAD8c2YA74RqfevRP2gSUhzboAysIYlrG280lxc4TO6KvafYnrAzn5vhCoOImCw1b
TlVfhGspTWm/W2QSvb4+77ADsmzNE7hggq8/CAVXn/RTK4DUGlc37uaih0qWEp2dqScRcszw58VO
QQn8auYkvE70vS6Sqz/jbju1DdIIpfDKEhNowC3KhSx1ArepzCSk/RQJ+rcryELdPGsToUOdcja8
UC+h/s6zuUEDubFEhDPzK0Unq3PqZ5CekqW7LF6t6uWNsWVaUBOzFiTqjqa4nPYlZJIbT91p0yAn
x/t2pRCDEtzn0zoscNaBH5K111Osq/nsvz8QDCFxheepVCRk5mmfG6KqpcFxxXyCGPbzZ1aGJF41
2XLtdNFiEHr3q9D97gL97/MuXfZkoB4gw4PhX4fU9oSvWl78Of6WbGrDkPRdCMZ7zgPDHoePdtJU
tC675eiOohdIjX1/7io7ix/rPiO23JEEYS3/lELqGDsCxz1Yit3yEtqKx6AjpyrJ+PJgfe0mexTO
OhAVmkedRmXLewYMbAt3KVbwufli5jj41J8EuAo1ehp2IR0unBi8u5RBdDuZbxDSAGqCH01W6im7
4FQVEHRV69SpqGUclg36bVxVvGN9ilaA3MSZoyNEZmIbXkjjr6mO8MgMuhcy2vDItJyZsgV+vrpN
bmIyqI/WTlZLxZeFVgUxkcWSjDq62RWw8yOPQwsoxpySQVUh8qeSxIGpLfEccAkZ1YlnQohjXHXA
4i4q+TjN00UP/oWSUs5EOXO3NBUZYkkF86tuhUVbJBwDGjkyGgZOENx101R4egZoylOq5eNu6Bxu
bmWK3rzK/p/ZCWxErDpgbCyCDw7lomphZerAbKLhjD8ZWpQa01YmaQDBALfrS5F5603EfHiR5FNH
uot/NR7cHg5ZD39z7/zh3tctJiWDrmYqQqoUN2fDOYRjpkTGQ1C2SWqSReUuw+CPkNuUYlJlZHaS
IaVWB7QkwruV11N8ZABmcXUZNcg4j/N9E3XjT49IfY0fbn57phlF6CE3vp0n83z6jyqs9umKlM2z
4yYWVF5nFgZoeVwDkSdpFbiw/xrzj/PZrOspVqwx4bive7VaqGJ6s82Yaaj4nWDQh0wu6weGy/GO
wksSQqd5tomssdJBtDYUTuew+vCrcs+pS5uE97h/Q64+ahszhCu2BN+1N9ExcBf0t1rquAtgydYM
NnpnXkhCKP4ZsZyyUlh8KKW3mfYHp/3R82B9sCoR2mTxuhVBUbxV4we4W/kOtJfeYnyMUiY0MG6W
pFvOacdSq0xZlSRCLzIT6MaKdgTGnPPPRiIS85bPz+sT1j6zNcSP2dDMhvDgskTfQ5qkuKT94Ifh
tDponFnFfYSMG40vJd+IWLfpHBcq+eNjLTphJJivSfLTjO62MXDctpabR2yImbxz/OE2yoJYZR5V
5RVaihQC+0J7LHSvd8qGTsZzKn/y0jZesnmtGnvMtefWbJeMp2gKeNOPjpWBmySVVnqk2086vdKq
Wwk9+o/xV2WpAApwlytF9Gg8CnrDJ9ZIo/L1Y6WzQyzxUGKqnEL5FLpTJty+sQ4KVdpOhxc/EaTy
vcM0MhP0wekhXVSuRtz6QluvcVcu0FxElLs9R/CONq3vjY7uCQKBb1nncz70DujGl5Bnb3HBIjez
pksWA67KbjmXlO3MmS3S2ZE3m7UdjfAJ6nTiqOSpR4Cd4EEJRaRUxBIRxCV3skqBDJtMhWEaE1Yu
C6rvWR/on/AD/PSRB+7vbbv3A9EGO0Kko+6JkG1KsEsQhJXsnPlClQDSYKojN/d8C73RC+mlOfo7
77tPR56QxJ8+6fD+21mDtu6yKOp3JBjUZLR+M8RiyycbrTzpRFmnvhQ7kdvbcOfi73HzXq/6JSFu
J2dzvDKQNMEAuFeHlV7tkztdq0PoPciV0Kknd35yiFtN8w73MeRcQpg0vGU1nebYmXTkN1BgFou8
rOSSnjfET3uP7iP6msXTp07UMxUk8muoSjBIRf/0Cxb336jTTGifd2zwWpnSBhFLpKdwG9bvJSdf
RJ869/uxZg42efJa+iLYtweQOFZf/tYnsdidaLjuQrBYwILGxsTSP5vTSXmeZZvxV7jKVPKiVDXI
7u3iybZPT/Ggx+imnh+94a0CF7dORdSxWc+5HnkChOWneS8ziOQghzPTAjTw79PHXhYYKNh1mghl
5LKqjD5I80opp7vA7x7XYnYxHJXSPrupMIyD+AXoO26Bl7oSERmGsmEQa8ix7ZjaO73Wo6v7+J4y
RRJV1JL4/7Oi4jE7cLj2NXypQJ5lIgdrDMQu/r3uBMgKJAR/ZNIE6AuXgFmFsXKHj/btFGE7XoCl
agpHzPhP7fDVnm597+7Wz9wSEgkR6cWY2nODuEPpxPJZy3+jEe7iAZ0Vtvx/1wFa//1l99AmuvAt
LXLeeOc2YlJPqiccOnTVyNj2T27lYy8dCeW44AVIxNNJqUgTQM0z4yj9bhCWoetglOt4xD0voTpM
ENBb1uHIaH3NO/DEb2QfiD8r6ls5c9bJr5g3sywEI7T49lKk/Rm+8+5fyAuA9oT0nOSgsx4z8x9Y
Xc4sSW9Z7S2V3rRcCSy7/gMS+LcQpN4nxHS+2jAgO/rStelZF8wSnFeP6HfCvV+zwiSvqaFipVGl
568zessTJbqdK3U/pbxNknxZXpp1TxQzBG7tD54J2E4xP5Sstw2bMxRn9OSF1yxwz3Etg9OFaUP6
ms7/natVMiLoFHvtAHPAPNqRkwOTfKEpAoNyF4A9CyPagut2ZEXu3si7SpW9QhxxYhGz7Q3gftkX
Asr6oZfmFDxr9TJx+rESjEYvHV2wrwlJiVo3O0M1QPZQbmVq0xn9MNjG0f60Ep6hdflGQAmgiYhU
BnwzhymjeuWqNaVyFlZ3WKvoBXDy6KmH0wTjwfcQZjnB7YvBMK3MP7uqMild/ZIY3GFAS+dhIc9a
8MRPaowhoaKzU20Z3W+ANxagU+MjSoZzrJAMqzST/+hmRqi7QZ0bnw/kHxIaVVREAAseygjVSyE0
3YOn+33qGMjILq1TuGtcJvsv50Px8WgBXArC6Hhh/ETIe1QMRiD8bB69AMQXehYfIbdM+QV62N31
Xc7QaYjjwXDV7XetvPczhk0NSam6jYF4Df1jCcgqG25L2XPFwjtnbuF2jZBG7x2NrMFf8Yt68VcS
HfQyfDPxqtTDDR93XK3KJR9QXFtfiJ+JDrDNt4+LObWRCRb2VYayy+wujvNNqBeQ1XG5pr6tmza5
Je/9CvXsw6pT42+TX1WH9NFHeoJwg5lJuMzWwI/Q8MURkuhq8NgnQYpJ2olwME79nA08XTLR7FCm
CYHRc1uhyAdxaiqUGe4O52nDDaZenxIhgLM9O8iIJ3/DqvjR+ulEe37iexAJBJ8s7SatnIZ6/XsQ
qua9Z4xf/prHfBlUGFJN2moc7y+6Rn0g8VmKR5JWWQjgT+FsG3Jj5kedgrlJci8nrMpg1msV8kHQ
KTIjFZxOn9C7XiTUwzGJ2kNH5/GLy8k04AFIp13gg05LoaOzqXG+3tHPvhqJdKYtlz7Ifbw+9ILH
CscVHY8zkdPQ/OG8hnQaRVaOafVdG+0b1tNh/PQnrltVObKtGlk+DZV66DYeEkI2g67rSkLH8C2U
Cjb0Ce9d7vsHMCPBtZkA0pmXCFafUMA+fhGUsR8++N/Ilqvz9HEeC0SfwCqS5poCwwLOmaee1oyd
A3TjQTAHw8odztHlSigT6dxGdUp5nmLgcOQxIRrCd+mkRHiJSD66x+GSMwDSAnqY35x5pH44Shtn
7SlGHF10QxWd5bbnPIDa9dk4b5BU+RooYByxUSxIKNPadzgUK9aIXdjqgr8wGy2L1UHBh9jA3L1C
Uk6oNaJRFXqkiqV9Aa+0Ajv/qQoHYnBSUm6SVag9y3a9lqBsvsfIpZ2e65+Z4dPMJyRNfYhu4CBA
+izBOxlXyU+QNy9xPPRb6vsYLHMv6M6OZiilEhvIu/cigAko2I5MSoVO+N0BIVo89/Frqa5hZtuA
bmH2/DMkqglapgyAtgkOJI8kQ27G4TIPLT09XXjo2mYuPX0nIHBinL1OgSucjC5ztyymNGbJkS8/
nWjdiuuPNVL7sgzuq5Jz3tnh8W1CSaqmBmJ0HEuGDjmjIzlDqwkukXOwiokUuumSRS/NhNMy5ugj
WSxJkTxYcXDbmBZdf260imlcTXZlDp1xBUkquqQU1y2Z9uR8jv63GHGU2RoU9AC0pimXAx1lU4v7
DNdYG/J7E0VvbaN8lVvgf+caWR8Gt6uH7qAmL5CusjctkyWSBoePdj6/NEw6ccHxant35gO3Xe9w
PABEGIEyBcFESmmGpbea1jAZBqfX3A/thmG46aOUzCTvADK+GXsFzNDIAzilW7i8EDEak9ii38JA
23hZ/JSM4bliyzand8Ar24BVChxSwrH2m+7SCLGVZMAQiQ3OUXeL3nmfa1EPfB+LNI563hsX+XA4
hkFEYvMIuRQ4eqPkz1Ao36cC4Hn8yw/OIAPAcUDuQ4v7WxPNIrwe5BwNM1u4JrYH5IgYWWyT9uos
4HNzZn3xpApWxSxIaFral7h4jKh2hGKpO1Ptyho/r1VpNvNG6qLhn8U4/R/1J/1arIjZqM07cwaw
GxQvhYL7+ibsp6yY/RuXhHA1L8xV9uhgogwJBucHOR/YymW4TMaLJpZigPkR2tTT6L8X956SnW9j
4t9wHZFGHNaPaoEc/fwjzkM7UDPKlS+dwf7uKRn40faGZMH/Wm9+oOSIwrC5+CBo/KcQH58Ry71d
qkVKigEo5Q/wfMdeFqN5vcw9fAZe4qdMAZCXw00PVPgxOINURaMKl/yOH1tIZbsXYB/YkMpTMy65
YNWIw0R149uNMPTqrCtfeyaLZB/VNRAIzXsrqn8GGukWR3AviF2bhzRvU7uhUzk/zLTyxvi3B7If
2J/p1PKfrRvHGEzvPx4eieGShtOyXE+hMPF2vWeo+Tvz0NHF5cetgvbHxkesYwgRdWfccJwBFGRg
6CWAl3qsrdw3XLGjHec6BIR2rhMVhGZ31Ipm+sDyd8B9yAcCigUj4OrESxJRMvMnCTgRknpEDAXj
vOor7O8b6f0QcSAsSPS1EYTbhBacANiO673cpKVW1sVE7cjNEd3MH0p3SDl1RBllRf+1haP3S/LI
w8mgHKn0OICtKz01HM8LS+hPsMlPmIbo5SlvaoyMMztx7FUaGPQN0L7QJpJrRRLDttmyOgIP30dD
AiZAY/O+dJDepACn3Po8cOnhuB3omesMUD4IITrWB3FmQfy1zg6zvjFTSakwcHzi2+HkyNjwCdPB
nQLC31ySjecBf86sMeg1oH7eyOq7/oQ8UDBo/9TVOEAgY2zWJW54IAaXBGHUBYRwj593A3NPxfFJ
1eZqj+f1kU3VCTpPSpnh0Td8Zu0ylyPKk8nbh6570tQ9q2odCE/gA3l9Gsw2jU5SoURqZRwxiO6S
aq8Hx52A6YrzN8CKB7LbEitxhxjN923GWK9L1ZcKeu0o5t/tMqJ9jXUC+fhykQ1ECxM+z7CoVa/Y
/41IynvzmffBP2Z95TvN/dsihM5U6RRs/oPJfGBNoHi8M+xetqu8fdte/uWFcspcDv+tjb+Tlh9n
oZWSvhec487P8beg73izjeldCCmICXw/nYkgEdDUFLtpU7VrhDYa2w0O/QJOL0MP87mMCaPNcijF
iQpAlqT1/v8s9g2GZ0iJbOHyuoEs4yvT43FadK8Qo2G4milKgUuAMjS8TMyqbbHAdUoEUXMQjOF+
TvFu1rZZCrvs9TMNnNSHv+NlunH8PEP4m0sI/NiCEK9eetJzx8zP0RjyXGNnc1T8fEgxzYK7z2cY
Yzve7PpAO4gSFwfFsHyE3hHLV+EUxrY+wTW4WsMBf90DpL5FJNcBDYK4x/R5XVq3FEzCPJncBuLa
Fi77p5FRR2+YhZJlLwCSZ8SuLvmfGPb04tSqI/4yINhqMerqao2oxoOqzAxQU9CpfnwVj7R260TI
wQffQtKKpIPKWGcFg1gGkHYV1gi3PR6b/ofavJp8vkjgEn6+GcQtieU0yIMQKpmx9KD35KZ7uUs1
ZUM1PKm9Hoyk51U8Ba6ltdUhI9x92kcq+1vn5oAW+DIXFMXNP+4tFyE7Vlk2bE02/RHsUPCRKfTM
COoNWN69tDl5auVsVKwGIycPIyoS+sBzjetjpq/vVi7NMr2Tr7Z817P1b/s4fPvyrak1+OBOTOhX
nTS80ZgEduIbhtqA7XdYrAaGIZ19pZ1w2+KLhQez6xjOgm8DxsARjB865tizIB7Mgm9nQUlz3nQ+
AfoMjApQyUMeyFfwbirjPXwcwiSm4th3zZGwK8nXdDY7x51jL0nkxl99mD6n7TyehFgosgIBQRQF
yMzB1By5MksNfw4hINlXnk6BzeoZgyLfYrlO6bXwmrAyEwD56qrwB/Ox3yv3GnDixof+63J9fXKV
qPi1fyH5t125c4Qxr89QZqOaC3p2Q6pSkxtliQNUJx37OKLIAiVGmkNos6auGjk7PDuSaZ9SIJ5d
zrxt9Z1P+IQwv3liA1xyEzOFTKXWzCQTfKanMLxFnY6M23RcaDvl3mtRBoalV3Cj8ux7LttoQFMH
mnRGeoaqDsu+xga/rDzWCtGk4EnssHA72ccGbPdfUS0PvtFrhpNJFDk+ITxUByf4XhTk8SWdwVz2
TZ3MTGkT9lQJMxUzmpm3vGVPoqyEQglwaZMQr0iYG8oj63OSZcrZMHZHFOzsuhgMOlhLk/ftvw3K
Wc2TL/c7j96D2ssxferx8XfofFftSFAnkEFRyxlfzYJg4OIvstcAS+Gjnz3toIbZ4IQMJJFEnQP7
olc2kvjQLT8uFre+Ib3twvbmkNvhStAVZz44T+5BDLR7bQnsPgLpYTV7nUttOGwU+0r/LPuMsGiS
s+TJpaU/BbKBjy4xDakWSf9mHD7bkOtRRsWRpDw/rkJYW55OQkpjYPLpoBgJIarh6riRcjQ4yr84
cXel9zBPhPejFpmO2cje8mvLSXFjem7IwwY8KNOtFJqlHYQZ2Uf+QCFVDhTgfgu0pPzn/wEr6OJw
KFZyeEz7+ptyR2phN3wy/MRXDwZ33E6Qr15VQlh5Qms7rMx3qWJbit8eWu92ok5RBFYeRHORdlCI
ILYYaaImd6XJH7dDkE5pwKRhpxe0K4nfEaJcSLqrngUDmpZhllONvSuvo5T2it4pYbjQsafAcCY4
BGEblV49exZ1HN8Xt+kulFzcHb0vvQTfMp1aCpwF6dAcen5/r8XO0ic2x3eWZM1BLg0YoDlkcwmS
0hh87HNxzueEMLq+vofbGzFVJwjsHPb6SCKsna8ieBgDCsvhYz265drklGFOfSW9ekSrIe5eEvWH
mfF5qmEtofPLC9XgOhlP2KTCThbeGLt8WIyO3th8tNrYrQjeKI0S8CP0CtDQBfbrRNve+Y+VLYkB
nFwMnrNF3fyBAX6QkOduIi0DnwtzinYfPpuScxT8khla/sJ/fFiy7R8YCMqZQRROjnNrqY+25732
ysToI55oEBLq756vxAtgqKF/WBwesBBnuBjbjuiStbZU/ttPaHzkIeGag4Y4okXHouVdyy7qleQ5
1mvRvEcgOoBEidObqQu8VPXtc9XStBCmGqN8Tf/h7b7aqRjAJ+7EYFfnFn87VkYnwDt7BUnM4mP4
l/T2MiDZ5otzx5CGK6z5KG9hUfTIHbGGP7xbBhUBLbE6RLikQZLcAlySVPHxA78hvGjJb4fJWcQ4
Fd5pPX7jllIZM2mPK8FipxGwyEdRL4dCnr/kSAt6leZFR8vBDMnAUo/VaMXEd7bNAYexqhCxoybX
jOHBOPkB8f6Eujtg4WQPlfevA1GJGR9eXRI4JzAMa0DSGGTDDW8Om2GcEYk/gv4zE/d8I3WdeX5Q
nw1DM1RDwMFxAoYIMLlGTO570KSrqCD+TyctQU51qbdoEUskFrmc5asIEszwSNiNkSLdy8v1EEnW
rS2AU5hxMFuACOJu7z9XKtFj8d+4b13cpLdF/d2jF/yoWnBQ7IoOcKZ0yPyQdnt+FlViP/GqW1Sn
llLW70Xy+vgX/nxaYVkYw13TcI01NxvRIMvLxar/k8OYM0UlUsvOk8g3iCCF1qAz0tRJ4m+3oKGV
phrO/5HkWattxO9UsmNpVvMkM+6QivkFS2C0WUl80fKSlcfVDoMjDCYSOlwwCcfZIv0CNms+eJ4w
orzShRDdRJlgkp/8rz1PmQ9xJRqqxVA9+AIlS4x8/6IQvVLMIiAfmz+4M+eGxW5mgxAKFCRJu98x
vjCyql5vNeFUNkmsVs+pYPP00sNU8hJSuqrfTT94AJVtiPqIZhEV+kxwtF+t/qrYWYIOoPyfbm8s
aKTn4eSzXlP6DX+SVsqSwSnuxum54XqsAqkldDIMloR/3PfKFaCFJJ/qs7Pyl+8/x3CvQ6JnlHbU
CvBRzf8VpL6Oak4K4d8dZDFfJaiH6GlLs7NM9Nk4ieo31i31F+4x73xa52iNyjT2J51p3sW60Gka
q0QfTythO/VHcZkgL7XnktiUNFgRINSbrb63DvovSiboDlE0g0yeXoqvaLWf7qkadZF3pjSOk8pN
Hv8oitZNu8VyFwklV/NNq2AxuHaqsoc8jLhNPpOUsRaLTZ83qfMYPuKUODMRXomLvkirBJ9xgBXD
YgtSkHjIHQEiBdf/ALuSS6k26ee3uyZ080hqK1Dd34b79sZydBAJz+MVqr5qz7I0DQx50RcZ//CU
4G9lx+SiEei4XE+FrE0u7UoACRfg+gfvRQ6HMFBiwPoNZaXSrZK8v5jX5rMh6qwcHvp/JLCnxh34
SufSYjeaey/Gv6iG4UUpKeczQZHD/C5VL5RJTpp5BwR24AOkRaWRjcZFXkzbogwfLEuNQV03vCjz
HTNVk0PzgoJdL1u0CFJum0nvPK7kbwbkAxSMOurODrAAMUyX+9lgwyquBJcTlcF6p4Q/IrdQlk91
hWuqGJBqzWHuV0/hDTDQ5uAv5J+gNuycmAdO73nY7SgY7F52ndjPS/Tx6zOi6lsKzzTzQG7Iqfx2
j4Y07zvPN8pKqTjgid4kK3gRy4TlnizVgC0POfBLu08Z6y+u8O7kOb6La5Vp6HuXu/x/nhNDntnz
Ni3Qbi/GL+902usmlf4r0XwDlnehG4YNo8w+9R8dLkj/zvITKXZYHeQBPZIDIJD55YXR1y4d6lYh
T0T4EmvbApn8o/ldNk7GtlaxSJJuyzEoW/dnQk4hyTE5RAP47wpsnfl7aWbC8h6FADZQ4ygnj/++
Le8BZrC+rUWF39Hc3Iw11YJ++Itc83yGR0mhe4bLhKli8V/Q1XuGdTPgZwPhaaiZXWojcpLGozEx
eIfVrXnVUeI9VMnUbWKYY6lOlPpAoVq4NrLXAttXzjhVxGD9j4BGrEyHb5ue2qIW1XztwNdbAyGt
pkAX0dzdo46VEjuQVzA6YgOk5/V2+NMYtRJso8WDADYbcoPjMRny5yPcK6prgfZMe1AgioS6BPtQ
1/tHH/Rqb6sJq31LifARmmW5+kvsf9CqTo91rr8AMf3wvuIJtFZGFEIl9BZhdp9v+VZSZN3Dk+A8
ZEyyEqz2/OVVWbPLasphePdRjXFfjSV2ym8dIrN5oc9Yv3TfzWn74++4cSk1w6ikX8zD4TTV+0Gy
07Oq6flFChE5PKb/6nHbI1uUEod/i1sdreRVHRSLWkLl7efG/V+MsfZ+cXZHtV254fx5MpK1RGQR
NoEW/CWQclkTMjNQReJL6iEbvCwIhSzjPdVTamIFtJwDhnFUOS8F3L5oOvw7TSsXcw5f1ADD6qLN
T+nqWEmK/rZ6y2FJWMqOa7Ugqg0AvcpHukn3+FaM0Iw+i0N6FtDQ7zu/j7QvtLxejgjEMt5aE6+e
bXFlt6sGdza84Fwltl/gNqzE9m4XbikS5slCX8oTaIirLhySQ3PljUFyObLvN5pxn2ra2T/e5XAo
I3uzrM8pJlh5kI4ZvsDLsGXTUBkGUfnwbYJsloIsgFn3dLheZ7hbJ6cMwvNadYj2JCViQCP08oOu
IMU92P5ZbB/veEB2eB14YEicAmGofC4OY7Evs0A+hEIo99ouTdEN35Hwyirg0PEEppH5CwQqE3QK
IKzHfPu2rv07zEtXYj8xD6QU3pOnFiEdDqYOXgQbl/+AwCBwhYEJs6nihLUkGcFHjD8b+12KvP5H
zAe6fHGXSEPnADTJ9f1S5wzzNeOn010JxyfH2HVmSWW620fpN4BmwkNtuyNBhejB8GId8Tiqdvzq
0g4FQ0ZfIX9RZp7sdoAKBS0LQKHD/0wfe2a9VNjagt0OYZSLIztVw88I+rofR2T66sYvOgxMjHXt
3WO4YsCl/KnDlMOjBN5f6KjED6kLdQ4ddf0DcrIMHbBwM7rK5ln0YzRV5CKais4WVn4TdYKlYrfo
SSzp0m1GDC8fQF3UL0F9ZpSaoBFBf/AqXCnqTEcgRWdO7EuQ2jnUmbvJEL44pEdz6XxlhNxWVjM3
zJd6+Qga7OZZbe1h93nAjTbKGvywjDwBMbRYFeHFCpUF7WXw3o5bZXo+lfvBSNUN4vt/CpsfZc9t
DE5rUlql5zAtC5S5qFb32Kq36gZ0qOjoifHaeN+yzHaE00mKR2N01p6OCq+UfLtX76LK7DYr23VK
cy6a2YcXW7IitVDx1kF2Hpf2OFxWnISmVM4yn9ee2RLOqrjpAQPC5/IjVZ5RWUUXnhbtrNO5p1yO
OL6gsbvIAxLJJrMGAvzMsWg8kkLzxxsV+iatFPCN5CN2624h8mxu+YeB/X8LojJ+1PlxOAofP9yt
yNvDK+SLpRQG4d5kcvz0OwqNCh7CMtmbpiT6eH001BIdECw2Cahk9iJaPFeKwhw4ZudLeWlv7mcr
0bUPNKZlIE0Nnw59A/3NUI22MORCZ7OkVJmNxm0FufMbg6nwjFIHflDAHQD14fmRUtoLdVgolrKI
SGGxwb1Osvhe5uZll0u6TQE8VzQ6Wjsu3q3GhZPW/ltNRQCSNkYr4Lb0YsvH1Q2GXBbJvIaJDIiN
dgard1Nxwzry2TX2Hb6TlpxvY2GkMswm72Ilb7vvF/XVjXtwvwRR8+P1Q24jwka0OWbyQpIrP6CE
eGxtrulcKbn9U5zGL3szkcq24sE92fyppCBqApDWorG/e/pCa6PfV1mxLs9X3uOxPminKyIau82Q
pmgadMBXWuqJJ0SJHdAhH2f1TBO6OY2NKh38ejssl6pkG5kN5/Q3FDoKtNqzhtPMxDOkcfgMm+qn
v4nGKIQ9z+DXL/BVdENAtbBkWx0GOruy0Gp2z60qdLRVunRDC6LgS5wxXAhY6sebvKRY2qIhefSi
mHZkqMx5Fqieo841Ak/4iVuAZ3HUtJ69qIOeQz7APXQBDggXSD9+xXUIk1ObItscPKLPowtcvrM8
dSSZnpqBk6alrvmKLRl9dqVf4QJMKnNIJibnPFUag8IjGtxMnO2MoIVURj5hjz7wSxp/80jRJFWO
JsgrfKYJHSD56Qal8vUobal8VD3SHBho6Su3Rf0GX8ADJsYtL1eKW7ydU3fM9HHEG5QjGso/f+g+
8tMj4VgbmeHvbJqsvKjJSW73LtUgRysr+2XCdwt+1tbipOvdJhKd5he3OLRYE0uaoPibWgGjoywb
5XfrzW3l8d/NwlCBD26ShxHsH3hGrRL89sZ+4FYgksJfjcC5oAbXbOdKHz/QnduhsP5VgpDTeiUm
IUtly5oPNBvCpNPyXv/rQO8J92cXjrZxf/E0JkLZIGrL6dDPz1EKzvrKGs1mr9+PeC3WuJQhXhvl
e9sYfJGj8KextpRn/1JvxQbfoZgAjIyHMz1jD12DZrzbRMc2fp7BnxhSc8PHe3RuYDf232pb2D9/
DBRqMX2Y+TsGDQwJ7/7Z2davLnj1PMjGPaTvXEYnBbpjdWMb4EwVEQ63B6agqksZ8GcJyxzqoTOZ
DSmwS+jyhlygehQHeyWlFzYlCHexd1erk11IJZ2cZbMFExmXkjrAcoUav8qdrUUp2BpX5wkZgvxZ
SFDE6VaTAtCfiMLT2yZMEY2BCz4iwPVAPVMYfEZ4dullTilnTzY7U76v2JOLP2aa8ZRlK3qRqVmA
syil5ccFMIsA2VLnk5nL9vk5BXSuRiBbK/ucNNbyEfEMu+nJUOGN1YJPvBopvKK4uLhN8Y2kWd0e
z/CUuxlh+0do1BBsPNcwS/ClbHM1s7ioWz77OHe321aIWarBXDoLVaN91TnphUS+c/b3BFFwSiXb
drgPzTyp5dkvDQMQ+6m1VTg9pH/+XcDNc4QbRj0Um40HdKO2/s5w/U5KH1YKWWq02bBF3pEBpPRX
uP5HperwP8asC8m/A7fyDWweehSOId2kKfk/CKy0SsC0khOnpQrn+foxDcEbWEelzSDZWIjDKFOy
tBFyhK62hJ+F8yStXPpxhoypcTJmhWOs/1Inc9U2HA+ys/Og/HAI+/laAwY1sJkXl5kPl8NfqiBO
sHBuhIk79K1DXdSTPZkKq8vdcFHQEtPZktvuhNx4NdtRY8ADnn/tUJKHuSiyjT02O0M+rdHiAuiW
PGpWQznpA4omirflXekiSzJqSdt6IFppCI7uBL2BkGvuFw5L2TtZh8v/4C+MfF+p3TsY+8hL6M41
08ypdElioPDI4b9LeXZ19t770BSXf6s2mE3S0Hk9JgTEfguluhLfrP2VorZh6eGugpRGFazoDXGu
azCHMn46BJDZW1s7N/r8Ls5uMmZ3WxJmX3waHqAo3XYVwoUPoV2P4IVvtBSFEFeE77a8k3p64BIh
YdQ1yDr73oymT1amJckl6EDKYwirXMQcVHvKoJrtt7CnmLU6mOG9nc51pfOfrSnZvtYstI7zJWg6
wopx6ynBjQNvShqDjTfhsGr4+MPkjjmu+pz25ovxCJlkWif0vj+7MSrK+jRHSL02rq90NXeay73O
6TuJ+zdV81W4GDLUFRJNGeFsOVR05CTvsF7Irpd3fVQffNrZJYs65bALFtg1vsY3BrR3NfLREmhY
JaBX1MFHc648rOrEi/pwKM9HNK5c62ryIDvroSPDEEsHjUtQkPOEL7jUi5px0dmTVVeIOe311+Xf
DoIePhpWEm5jmWkRr/KN2DwKAAVBwujPRip1zO2virWT4ntySfWT5OYFOmsNOAdPjauNyU4vSwEl
FR1UdHqtLieeAoRdDtDKzwjfNbK3vIOj+xspT9SyLNMJRxC7+eumy7P7mCpy2K5nQxGRllJwYUAC
o7fbM7CcHNIF1BUozQk3caQNhrRMo+d0QvnYETsoAq03NrQoSx42RZ7DsctftuLJIl42OX9hR8D0
N9MwdjM7MWVDuZITbaKqqDdMBLPphvl28rjPkaHXC5XwXFFqvp6WtoT0vtpGGIDMMkF1LBbZyHBn
xg59LxwQTK36MU7VGPFby7Ro5JNXG7kr7ZHCZXb0rj2btfrQ0ogiqHctD/+AqhWXjCDW+GdAQH8d
VcWlnq3jr5uNoU0jQsX/+BgT+6hF17+u4pOA4FGvKEa3Ddd3UjXpkcaODTDoKRS0G13nT4XmvvBo
K4AcN5UC35ioZ+bxWS2iqYBG1WhpgCl5H/oCwd/pT5XAib5YIS+Z479IHMCbpadVkBLbS08+fIf3
+OoXYfUHIJ0vZv0+p9GjrxHKuTivibfXQoM+fXDV/aKnki56PPk6Q6mm0TQ4lZWKO4sP7gNY6BG2
3r8+pXNCvw9kHrLSwDBksFxoCaZdvMPNhC+h3VvXyfciU+kIhynT6qMqUsFHnsfQfHVunuDqKQKr
pbCiioYzYTdlSRDXYmtmPywoDs/jAkJdn7bFLLZyDTRvmjh87cj2WZ9KN0l1kB/5RQ/loO7yriHC
qAG77cU6FmFvp9Yt3j3aiwnm0infvarfv5+7tIdAuxIIXysliU+8mbO6NwYGJDvb4O+DkCrQnwsD
Qj7hIkcfbffa9PEZatdPCMxl6xCT1L7Bh80JVvajCH5z5bdFHFTFmrBoti+5cetumJSw3FRxkerk
5pkJTPau5vn4geIyFPGsGJgBq/3cMzNgI+MGgQ2TjgB7cnMKffkyY0hGe1M1Tiu150olEzRBOjqP
4vrktaNq0mNA35BsumQvNjgUGS7NWrx9xYLaE6Ly5zD/IKEzupBGPXLQjKbyA+r6tOUTEaHfEGdj
0cmlEqadMyZ+P5Jwwv4LJsxTFw1ywv38P3M0so28AO86tvdfLiKfsXo+KIP9lWlfi9r/aiPM7kKe
0HYUQ+ySXZiqJUAi23tal7HxPE84zFeAw9fqb0FoL2IGjQjrlob8W7IiDBOH1zPBv/OyBd0DgS+j
sPJABfFAMbluiUPTYYQmcyhkVNjl9MD2/etoJaWKcqCyRhDoqn+QKgSj2H6OfEFlf3d7FBRyn6bV
2tAqZ+ReVjx4fhMOF0Eq7dxYxgpHQprlMl3kVtTMA8Z9uoVh8zngQXK13nLOcyecutDiI3HNttpz
6uRHkra41m2nD8UqKr3xogomr3sucyMDo+KwFhrTprPTnfbwPSc4UPamt6hMkAmTgs8fmF+Yb4tA
Bt4RBkIlm0m6uH6l0PxSY1rteojAvK2lOuhMtf93K24f7d4XNiu5cWse2YhXbw/oHIyeZQkeJ5fN
N9xqm1qDu2JvxbSlzj4EYKvoW4N1EBWRkI3NOLIvIXSbSSMBeYjxyBkxhVfXrvACVxZsYpUent/a
2PFL0JdhAVkzT/O9P06ppondjPxuTi1a3wo90B9cJfneEWGdwRuWhfFVOgZHDgWVlliShCGZE3BV
vLO0/p2X/Cgf5zmu+zIpIek7Vs7HI9Dk8Wp9SbdzSKZtjTkK3/l/Ht1SZi+Ixzg1ApyvDT5mMOYn
CSXDFRODJbxr95CSsJFVFFwmufvp8BMRVQmdOvyly+bOpd4yK5YY3cC6V6zN+SKwpGzdE8i1gSAM
Ml4kcu4ZpbxE9yBfyiymE5PzKSkBvENo8PD67E7sfH6R/Ny/j7hr0jYlzz/bSi1bQdy15t+o8UU6
j1UbHKxmtfF+GglqtU0j1/hRzufbkWny3Lt+dyMjB2Q60UHshvqt79sSSnTLUAR6DG2Oz07nL4p9
HaZVIagYajbTIB0z6WfHWA1LNaXViP3XsrGLJ2YzcD1Zm1iEfX5VZDj8T9C5h1vtdWZhz5EGdsYR
JRqVkGscV8MaXePJbd985NH13g/9iDD4Vms7qQTrp7HpZ3N37BZTaP5LC38Rhij1hf0oAYg20yxX
2DjQw6st/QUM9AMRjEA99L9zjqQzK47Loa3XQBlx2hj0GQniGDTE5nKUupL8BtoOZ8UOGV0UaFzR
4njchG0unSFTditzbfFOM/dxG58icsqvw51oPcfk58j9B+vJ5UurkjTgB7meb2Kd2W04VJznzfKQ
/Kb7M5hBs+Om1f3W2kjYe41Qvu5kJly+7Z2oTKCBYUdXVYbO4CBlL63xgOqS0+YhY2twvd0+5EBH
4uStmNsisgCkXcYuC/RAZNh8gi0JdssYUw2ctBb3+0G2BAiLe0/DAm8k/WcRKQjbjrzfBfSS/6hS
LgIgJWqR3vjYWM9SscnPTPJKNXvibCJuyFQwYC+PKG9WKWl6ZrLvynsZzcDf1WU6FJqcH/GpDmbO
f8y6wZx+JG/yYKUeQB2QzFbzQH4XmHm6QIGtcI8nh0K6tMT7ErghKvMOeguBBvO+0PxRL35fEhlF
YUF2lHW0nk1pfD1qsbHElUMcLCCGnWRH936qWPdNv5VIWiNVvrSymFl9le5ChlMTpQn2duA0kWcg
O1TkGw0i11bFmPcTfGRQdyS1gCgCuWewuWlTWGhffJhkyElJaWeZagk7jAT6M2dwnddi0ZtKBn9D
rJIeI3kM8pZnzQtGWPxus0b3ahVZJqMGf5PFlWS2qC21GV3VEIlMUgxnRmfLmI3VHiyRudJjkePk
oH5eDDjlUfaSQwR5Ut0w27sU1yjUH0r3AMcVQVk/luhvcW9asvqb1idlQuHXQ+k2VgZVXQU/w+SG
dyJG3IRMA84ULdPAk4ffeiQmanM/2azLHy3T7wtmeFJ1FY7JrjlVOc9fFyuFDWjMv9nQ0iE5CQoY
zXZ+znZyOXIZXd/BAbUe440MFNVfV4n90GfvMJnAFrhtFqmSPYM/WOHhcIz/o2EgSdW1QBNVGstU
UBz72T0hOveN5OzEbJalTvs5SZ0hMu6x8OnM99UjSmgfUom84YIBkp38gl7Gzknbj8fV20RaMkk1
h3Y2h08HTx3oUwT62kyGhB3FZDMEhNf7Ips0WldEISjTh9GoBgbSvv1YREgGPxNJ+1MBOPR1Y7Ad
0iU6EmCiRZDS/IpdSwhSDgxBohIqzU30bxtibOH5JZ0Vh0A/ssGePQZQ/EPpRken7yqQEBgWAoaY
gZGA0dThSLyHw4cIjdrIRij3Em+PuGzVam1r4EgWXKECXF9tbfl1hJOKIiIS7mb9WcNQQDb606Bf
hdfCT2ldhp1ZLQDGOOaOIG0q9V8JpcUmaVsNhszZ4ybucWE4baemrZgXWp11erUptuAMVco0oN3d
YD/RasFg4yJf7Q4fZRMMoecSqs46GTulii34Z2FFGcD4+K93MxxZWj4dpWU74ixwOW6mKOUewx3m
FZ1ZAcl9ppPR79+dx1DdTaYP+sO3nOao4+GfbrZ+9rO2SWqtHlx3t73ZOALytvdV3JWLWPGYaW3f
pxJMHPMPsssqhccIr8WbpLnB6a4+TPQFU+Ti5fZS/REibRA/ZqGhLjtedTSjcHBDTyvhbsPEjP6v
r4OOEAjFZVjyoNd2yMseG4M9p/8lP0Wx8eECn97FvcQGyKjmskdCpyavIAqbYGz212MgzbYIplnb
rIrwB/s5yeuIZuaiWcGFvOrEvk5PEmKBbx8EZvSKn0bu6I3g3iTDtwWU00Azz+rDlgOmQtX4jbD+
NCl7y/L4ZZsvzG+sJM/IwIXPlKnjaP0sF5TufWSqKQucv9NsisdR8XvDx4oPaEOBXZSoRtDSVBzg
02B4G6it754yhBv5oUlJnJu78RsQSSQf18FlNhiKV4lKzrrY3fjClg80FKmb64W5DRYAOLaZ+8Jj
xzCuLBr9V7vyY6la1An4879B5/tELFH1xvk1/ZpczYaP4KTMoglXABrVT1j2rYG70Do79/OUE3IV
B2Dn5jMyhiWjZSS/3MUwdZMPV2mAO+q6/vDV6SladAc/AJYZaYhbT3cr/2+4sXWEL/KqxdIvICPt
Ne8RZ8Y1gP7i2uJ5ZTaL0ZZD9MHcmjRCtqmuNRr/6pAqgjaDMEATcM/u9WDpi3YXBt2kVmGDZXps
A03Etm1m7NpjfJCvatbGzTCtgMzLABoeh6GXO/dT1sSpilPJePxRK/AotYM27Et+E/xKRnALIDFi
1wGuRbhbk6deootw2QYf8keK26/6m7egfZ7fUmNcbM5jr83o3HfxzfsvYTFPPhM3BBiLHLSPxcJK
4irs1T2inDJajJd14UsCpdzKjxd0Z80KdV1vHBa9ztsJoGusOOGuUfVym9+NPLp1JK7C4Snl+IID
9EbeFiSVDTPDE3dScamuluk2a+JfUdiwWRz1sGMd4VD6EPXRrqvs6FwdWfHGuBEcUjeoTmW1voEN
yO0s3gxbJLn9kIyqoIc0FfRqIornVJz4TDGZjn7KzEdjrqxnNiWB4rMLy41H8o/7N69Ma6tArzi8
Vx4qE6+Wtu8mq+UxuGJ0a56MYSrutjMTHAzO5ssMP51XMSLgNDmKcT2XwcInvrWcd++k08Twyisr
1Hcg6AS/P5O+8yeh4KCGebGVOtCBUAgiB4e/QkIXFUUEwAfzgzrI0Ke6vVPSDB7G1+ZxniK3TARf
xqujfxN1RkUotjyY4NA5LEjkZ22ruHuocEIaQBmml5QLGHJEWDsgHvfCcyOkYNkO4LKVvoguPzPu
CQiPo9EqtOJUt0dVg2sg7og7lA7pe8b0gWbWZPxW8dnstFVStEZcla/aovHzZ4b0Bj2rnzqKJksK
h0YajhPDBCcjIykZeKtmZnSUAgUG0VxyYO5IRqUhS+xJjCim6VBazGoGF6Ya4gsljyzBTOrmSHjY
8tVsAtYlbUetP8miY2uLzKnlFTT5K87mVAoCspSpcZjeBmVhbkXgutrUvnlsKq1AbehW3pFWgvE5
jTi8UnVLP4l0VKz78GGeI5xf0cOmQPnSBId4uhC2GcSeW0KcyUOBzKwLeYr859ka2R9l3J51V/3W
gmbs06zeOVP2t0VvWeWjKR8ez010p31FRKIyS3jdTalfgXznVm3b66Gx2PoUGyuDmS+yxGtz1ZnJ
U/3pc833PdKstA/tj7yvJMcYnKzJZQ4gGskgDM+DVEodtEwzp+yCgOKGeY0qYNub7CXrG2rlsaPO
Y49+6k0KV8KEl71z4ExtLEWP3k8wRpA71eBlV1XZnHtut4dCl23TjC1Nuuw2czWQODIdb4vnAA/W
Zotpxo1VJG8fvT/hbsUgTyqj7sryghM+PSHyzCM6hH/IjUrR3aTAkZkK0NKrvfYGfsbHgjnwPi4o
A2zPS6ufKLDYAKlJ2PROClR2neaAnEa0sV3OW3WWdMJyDKMSlqHmDtb634H3pOLUgJ2AMz5dJhcZ
JYcj4g8Dm/e57Q1KWMQGY4vdEvJ3lY4zc4GlhsLIWw0BWJ1GqCPx0FLpqX9jJzkhXAVhtO6tuK94
7Eif/6l9qUwm7dkxX5hD405ChUsMZAIe8aNG6VuJdIO2nRS3M+dMzOyx3ZGslX/CEmwTw7oxmH11
On8ftNIQbg5bZwyt/ET457KicQsEWph/PGGxX29u10kvYZLrcCENyLxDy7qGAJmA2KWhPgi6At63
zQfzIXz6a+kLVZHnRhPc1PpcE4dg9JvUuHD7mPbL3Mt86x0RVxSdvBkzijSmmYjRyaVoJzwVwfjq
gf/DtACXbjp7W+EwVPRFtdSspmK4VXPRYN93owaoci8fXpGhKAP/9tHOloaHPvaKHBCEsIAIxSkN
PZPNMMkPHv5LHp9eBjlFkGVgMnQYtntbD6OOrpEcAtzpbzhdiUuKrI7y1ITYopw/zmfHKBGtDLTj
6NMXu2Qs/lDgvIVZul9ioXZNXojxaxv81ttt5U5x/Rb9mUY7coR1W0UQI3ZaZdYT4pQLpgLo/Z+t
cm+E7Uqz+0kkzm/XsFvc/Nku/SfUOdI38jrC9qSYVqc599wiPXSjZjFF0MeczPuImwXu5gqUKDGz
n3WcOoeH9DGNlwpdAMp4J7WtWIHmezivu1oM/cVN+/wF9IQwwZERweLsBblmq53wLq5G31T3pvQt
DMESso00cdijI02gmTQ3bs+ZsFTBDQQw/yyZfufYKJToLihUfWx03EGvP74KS6zpP6aDzAUuusJr
rksT8QknLai+Lp1klf5HsYxpWtJD5T7JszzCuroR1TSyrT03zaJCVjp/TfbI5jwyYQD9498leNTb
rhqtSKSYPF9u/hafrWpKq8G97MvU6kmqWj3gSkQ+K/6JFiBbpM4dkBsW55f3XS5KyOLuUViR1e25
l2qTM6CxAWWYV1DFsttVx6eH4ui5oM2Hn7ye+PySejMquiIbO6TnrEFCvGTmXRePg+qQffc/EDAP
q7R/us+tqhk8Zu0996vSJD2LOLEgc7yj97d++h25MabW9B5zKo1l+W9w38/HQ6iWYRpNgPqe81uE
F6lNwClXSlDvDI0IH7Hwu2BCUYCaKXnnODyIdC0hB0ncvC2SvxF0qW6J6WAxUEngR15EWNkPMYMw
ynp0HplVv5iQf+d6zoSFw1vbjFYZjN2YbBNtFZl9pLA6M3JZiyYTFPhqvC0ZBFjJw1+BToST1tNg
GOszCT6pMmjqxtTMbsQHuX7twy1atkF+7MkgZ2tjNX/nx6/hGccayeXiTIsGuYX2R69NkE3jIduM
6xDMqzW96v9965XmaLhIYjO1OVlgnyV4bFAiYu+oh5fPcAYg21gv8hWvQh34omsEH2cihIrvDsFb
CGsL8huAjSx7tObxDTrYzfoMi2CnwxbmEcQVvUuCviPtQg+zK95SEh+BLs9jFlIP5IhYlKgs5rMu
Pqoamt+fgEDk3cV0kcVVFYjgFfjaMxH2uH1WeQZFY1+bhyF9yV6QDnQcIF4yZTvp2INemBuHbg/q
GdvivAogfXcXK56hvgvVMKsYd0a1TXOK/r0NW+1HOJrOgbJZWoAsAbId0SlwnDTwT9KC8Q9oD9lx
nQQszcb7iGMBKyPcCe46CLptS3nvCNjAnQyZkHGNWNys/gth0VGD2N7ZQ0aYIrp48jFAwRHIu+Jq
soRwIK/aTKBIGmg0bO9qwWLDZbprwZS7GBvg9mHvHV42jEOsc20Pxf1l1qotgCV5dLbqsnHPTIaS
o64AB6cDKWnp9O3bmU4hZpKSpwT3lPxXN+QSsInJs57O7v4NfeepcGanpqXVJZMnEgwUuSjbkGdo
nHbsjlIqC8w8+Dtamrhf67S7p19nlHN6pLuC9zUkJhuRi1iiy0gCTdcWJRT55gXLSKbWgbUdUx5p
TUC4yzVDkYOugGT12Ix+oXQVow00tBj/wKLSmNX4A8t41j6d6w5jxbIevADQ8U1eRKvPL4GxT9si
rFvon0zs7QR76fWm5hyPcbKEPU0gKN9J+tAAacHLB6q8v4q9W181ZU3M8maPWkzDV7Cx1rzkszGA
2ruTZomz9kltH3O064SLy3RdC12NWpOZEwmr/LhvWx+nLhQkEiJKZ3BCLKqpiEU2EJVZgGj2icZN
O7R9nSm+vK5XzcVpLaJ54fPluI4ugGQd0QbLlB7Qa1CQ+WY/OqTIjl+3jTlfugfUfgea1jSxVcK4
DUkvjCvomV3OD3jUCGKDsihZfP622XnoHmcpcQC3OOvvz1KGGbH/CZFlITr8FG3+QyJNwUZyIMAL
4AKKG4OYCeUUoxnphWwP16hIZonLcjdLqhaEI7hyk21pNsR/xDpv3mtrKCtaueBiqbZMJ8Fk3+X1
B3krZphM6XqwvZSjheEHsgpkmaYXo8QC9wRGfYqXoRXnhX2ma7krPuNAFCrcorYhBci8L5FI4kEW
wAFFmKSDskDA4Lw/utBFNasDrghelzNUVXEKYn2pJ4poT8QxIl4TXwnT6CUL9j20ST5OBBx0eFME
9V3qQb39WUz7ZTPAqE7Ru473X73MgAt7gENQPonDClz+RbQ6DNm+tTT0O+4DcNRSoutU8Fy1eTOH
c4Z0IDr282LO0aAp9VANOw0bX0L81l9/ptmKd0R9R5gtrmjN2690dgmy0xRRHj/y/AwS5xJsg8RA
Bb/mDay/NGNgJrMeFVMFcHkiR20SSnPgtFXJIG3aahF+grZf7gqmRUsjW/wmEsPM9IUhTGHYi28v
piQOzIjupJi+dzMzyrYw6qN9SFxi2u4nsm50jUZy8eaULjKSdD5xGgZzEo8jtPLDq1118iR0fq29
ZsVW9elT0HGXWKIQS4uxH1DKiWYBeDtt/ztkSG7vHuQ9yDahYA/vvx2AGqf0rQzYTi/FOz2QrJsQ
rmbZh4Z18CcOiDhj6oJPvsusDIiaUxDzGWNdcso7xnxhT5n9wSIfTY4LxAWEya+QL0NsJ0or104y
o/YmSydnUWseLL+vBUTAcVpRba5eH962+VN3NPDUB8A2K5TXseNSpb1mDRHxG449bpgLB4atnnsN
UsX5LN0auSMxmwZ305B9Y2sUA/Suzjm9JFPsLwdkEsUtx/uShmorJib0aMPeWPAJsBDv+jYJqGhr
tW50q9URWsqXKcyEMman1itE+QFWAeEn9k01nlmWZYcx90T2uCguKj0wauXGoHNyamRyazLsM0kd
Rf+qhJoHLIz1FabyF1s7DQqQfs3xzHqmxfgd+hYXSW3jZkRu07uDKHOHEeR0p2j1zhC1OiNnLaKK
uWoxZeHa1wOyqx2lUzIILkHyrVwicHDAL0en4B4d45qzp98t+ouI+0kkgXWThbh6A+vDMN+zRsS4
PXKYa/Vvy42nCtUlGJnalqer3R+uwILfD4LelMqGR1LMny+HtKtwKiZd+c+XYZIjkHnRlcBychRA
43j0BpDx7WEZtf9Wmi4SHvI1Ojo4D7qOfqZmdzqqLv9UJ7hyNo1c76c1RoDTUBroVHcHT5v1Y2XM
sAy7MSYNU3eo2xmeoJoAF+egvSZh1solz/Eb35JpwJi2ar8GIQZ1QV6GQj+AAxInQun+Lt2fhT6g
i8M1bd7/7+0cooG6wLEOptWSCBoYMMbDp+ggL9EVhWgpuqo08zt4P4NRKWo8NtR37UATagxb3nIE
LkugTzkTmLAvy9gKLtHBZ8B+shsvPMLZhmCpy6JpbymQyr4L0BNwEAi5sqNIINY2hSU2IhRDOzRK
6uwRSeWol1Cdt/4M9dFwPLkSsbhd4amcm2tm22x3rustN7Ojc/f23PCe2PJAelcIGdUX12ltfK/k
X3MnIvbYbybsJu064ywPbdhNEGIPqNVUTsRwBD7KkCLUDTPYubsoNRrd9F4w01P+y90KB5Qx0box
Et0i9EF1tX+qXRRu9XlNCTTMzWnR+20ABnjjlrY3CNdOiCTlSOY/sd2Xx5R5SlyE6RfZZIggQWEf
rY9BPLn7MxGKw3JZ2k8yD63dHiicZLC1ORcffF3Dfd8DtJcY/K/TUf0rW4B4W8FSjRak8A9fD6qF
YvHJIgak1zDOylRgtMHsU4xZGx6XUqp54SAQgNAXk2quRtu6lM+o88UKwJCTnyGbfUlfdKdFJmJA
trz4Qi8b6p1ipheknKHeTHBUW8SF2J0caBcF3j00trWPJcc89jSaDtIco1Wy0azVxenCxxNCWCon
1Pt599+T8Vz9F3mYRu9qEBxeQkWvhM7InjpVRS0qRKaceuSsRG/dPsXZOr+aAeC6zju8OqLWJ4sI
tVTgyABKMAKNsI1be3Fko+e3KMV9F2rSbqwRACvPBo+dQA8eh591VlvVIs0cYPr5BwGuIBeqX/7Q
pxZievGh89wuAcn6XmXz59Ztewfq7Htu1Y7212fmtaBdkfFSE2jFs5LvQL3ts8dSMHMJoMyrgYbv
IhbpdEG+SE0Fxik1fsHxQuvbTevFIIjSdv7fupjo4mgiw123hy2o+RaBOqXkEZka3tMUwGbPAWtu
/bv0pKnlzw7d2xmpQykCd8G5op+c4GYHhI29+94w1kXZJeCDeY//P4qmHmbyx3WIotozAt8VpRvO
93fRWVFpXD84jaRWCQd3KzAMfSIoNkmqUIAqtkAFupsQDmLFpGfetyCjXX9LgEp7qNt2AvZl4L1h
VnhVU1Pkcz3Z/+eF4xpnocb4dWWgII423KGoNolgZoluNEcUwMuCPHXTDO+Vz8gWMn2Sy5lLng6F
vXhHdcTcXQJH/gGsEBPaMWfgdqnYWtEpz/Wd4mJAZHjjQnm5GCBLu9efhhwIsm2UYhAwbqeC6fCr
cCYPvjebjTHdNbSgkLtMsoaAicT7altC0V61Hc/75ZvFQb2gshgV0Mpsm+jVazDilPvkS6JUemLf
yau/9LunPdzVQ1BPZuD0FckE2qre1ShJn2UfdyZmo2Ktjt8MV3/L1bIXQqBISQzhpruLchLZAojJ
YGhcNy42FUeZVBlB4HQxsLHmcfpYBsWw29l+1EbFcKD8nydUI16WqOLmLi9Zh+LimCNERJLQ93ej
hMVrJTulrJ45Y34idAQo3SWtbsh8mWOio2efXPKLubfPIXkv81+tczidvoAY6Jk0eaLSPUjl1rh+
Xb4yZlmPtVxcV9qXoPaFa7733lEcKmbol4htfIdzUg5HehdJEeVz7jcCu5G1LsCC1V8UFtWdl5TP
0CGaaH8nGv1YPwVby0ZpH4WvyIWmUMt3MTL5r9SbLSXU9OvsusdmoX+MvGgm0/KNLwuig+lpmSr9
q5MNgH/VRJryo4Zf/cC/0SF02VqygFt0dVVm7rFIuCu9xXhh4VW17FAY4tHU75Wf3ftsFmYoyjqD
d5KVlvVlWC0RQIV7RC6xXDOZ3WX2Rk18FyQHFVqsIwDZeesBAk5bWKja1jazEhUyib09iQw6EJfU
POGnZ00fhNF+c7FHG21ROjQNjmutzZMgidBcrvODx0O6MrKrx18nYpwq6Wa/ocxMJLfgDH6tut08
kbivzcU+rxjK6ZZ8n89NM5urEKwxXsZnjL1nFxuKA52pMRfEuy7kLVsAtAlPcZfdwmPHgus8Pb6a
Ask8exoiA4RbQZE/ADA1Jg9K+JDMzV0z3ubE2swxbfzfkllE0lSDRGATFMBBpBXxssKCNI0hl3gN
D3zsZh/v6MVVgQdhAxn28pmAi9nbNHnhK7E7/Hkj6dyxwlT0DsAh07Cr2SgBVRRnlSE5NHiy+7Hz
dFvL1CvKeqpnoDNv0opQ0rfS69JGu/Q7zmQ7NEhjecr3SbyI6qg8Ed8UhPplVH4McQGQ8Fgjs4Bf
VIByhOo1xqLR7u3jhzuDn6Cgl9JbRDoAp6nGxzzeXQfDiuc7pBpFpCU7dZNz5/8QsyT0e/S+OoZD
LjQzVIKxPshkjBdYQPIUhrKJlzBbM4hN7pwPlZh+ek89nIc69WKKvAWD0UU0ATVAkccEj/JIwxKc
pa7DEoJ+dPLLk/m8NYqTwLP2RqaMaJUW9VDTnse6cR9ENHCuFJfZ8oDHEOI6QIlzCZBgYaa+WUV9
bWHeRi6zsZUiQ2EiIjXsPAMitazx/ZuV0e43oPnsWSipIOAm01/xapozp+fGRFyvH7w8wiAu1YHF
g0yDoKk/yDAvJJd+hrb69iC88AK3PmZXb/UidNiXTCI2JGsGSUmCTThzt2ZwS/d2QDgB9tnysZ5c
oeBlyyvXbRrYBuaWDSGdbLXdo7NjMfPt/uErydtirCZ5E9SXfT9MxAlt8BS4bp75L9Z826szc+Q7
B3nIJzbpBwhrl/u0JzwfJ3VSbFOnqdshah8acV+ZSKiWlD/ZQZr/HOe077dsqzQNTVu/93iMTToH
Sq3d6eU4ZibBZklu06Tse34TUjkNOHWYXRoFjKigwVhhRJbXcP9fhMSkW7pUEaKy6e1LYdCyDeRj
r4aPfkTRiZC0lCrLFmizT/cZSMIF1hM8BZDPq/wVxc5zvpvWYANkPBEcia46b54BP38TBJa30HGS
otBnY7ng5uECpLwd/Fddt+wSynbZc4XXQC5JgdLyXmD7dHG7uF2aQNv+AdqxLeVWnD5v1MJA9SKQ
xxCd4Sh5o5VwRF+i/MPcE3Q8D+5uHiNLFQb4plsmCGVnLY2zsdmBwn+AIqzScRmTNMqIfwmKCgE0
/54FFbt5SXzadglrepinGKSQb3nUXCYIO6Y0lOaq0qfE9YNG1TRgFfWUebQ+gsnNmorb6uGRnz0R
waaWgxwsaBPYS5RWOFa9kdLNiHw56AU/Ocm1M6vFgoLPr5p6k5wtCtP29NyAPRckLFEB4AEnEWud
LzKLbKwbF+JF9axHBd3Yw2N0QjJivBWQUycNrnaFkqmBlzqgb2X7KxIlLGec5Qzs/Zg2GOCU9S16
EFwA2L1RGWzwLDaHmfXGh3/OYgEb6K5uPvdlcA5/UgzhHcfsFg4JTf/x0lmC7OXTOxcyu+G/vCFV
a4kwIhc8aHy4V/1praf2f369PZVQ711UL/hO2AtXAIwjAOiXvjjHPQy7T6ay8U4AvhjtT/F46sym
RFhKPUV/cNtZBfzPP/kVsh2vkDbzEN+7q0wf0HOgfuGtHS5CGUfUr+4wKeIJy6Ue3GBfa3u4R7Tw
/o8Brj9xX/Ic7szFp5H2dFssGzO6dyihCrdFXEsqb73ASZedRgxOJYo2JoMFeKXRUI3FtA+OnjV6
sxOF3ISts4R0DPkIhHW+kptF9SbU0bEWyGgJbACktrSwRe3n7TlQKVAyrGd83UMmz1pHfrMTcH1+
Ndy1Mu+Y1J0XWJO/OiTtdALut6WzkzjfDfUAq3YVgBtBNKnSopffTsr7CHBJfex0WFpP+5cu5f6j
c0x1CXBRMzg8otdY4sNQhtekTwhuAqR/nPNIZ3rMGYk5yccN0kMeq2d89L2m4YH4k9SeYrNLAjNX
QHzN6M2EHmlBzREBX/geGh8NbzHLi4V+XD7fjFjE3oj2BecMdxz3KAomk1vbBMdVk8T3CwxIiEvd
pVdlSijd4ZY6UhWAiWDGd0RHM4Iy/hnl+tVJICTN+ODM807F5q3wG/E9+o2jv32vj8HCLNODf/wp
+ucE4Q/iFTIQO0j9/YRs0WmZXlTatOIHBvC8SlPltONZl8Xh5fOne52+Sys1nw0dQFT33ZBzh3u1
/jxfqMzRHV43tRTLxsImdFL9OydXCjKo0tJk/tIuAHD3g7m5Rhl9d5dbKyDkZLsJRz0bcni8RJmb
WyzqS9T7DOeHbjWA7bIy4aqMuu7CGAH7lGDf6vs78zMdFmrxPzucwlipdr44pOnnrj6tPtRNbUCo
1KCJOVM8C8FTGcMQUu5yyrM+fPootxoWhxOjLiwFxAjiHfw9ndAJQzV4gbQK52xibHmhycLGqKSy
9Uj/zmJzwIFdk1ttdE2ryl9Ut+HYSgLxopMHo2WR2jRcuACTVsvPbobjLOFsiTiN2Os5pMx1khmB
tq8rMKC4sWFdVxy3LrtnY2IqKf1Oh24ZXY3lzb0Y3Am+IiSAcauJLWksDmJyuaqt1aEYZSZ7K6YZ
FqmS3mqVZZqOFGnUiF1JqcXT6IMtkfbxwdxysvVX8Yo3dozyKU42wpcaSkVtULzyzJZtXgwLD6NV
ZQCgcWZVGhNDBotrbbclVAGeXo5L3buA9xBt+FhMQLKBMfcmT/L0DaUPyfwXm0HzmEJ2B6z1umfm
+FOgvOVyON4W1pKUYZwX8RL7rh8NlIul/M4m07jmqIoDAYdePxj7grlGQOjrxCwnkzowzhrQEJVu
L5AFYO5LtjYEsVRm90guuzpUvIkujcvXRpFboRJpZSZ12YQVqOGorsEThvn26wOrf4ww2ZG08pjE
bwiA6SFXj+QbmenbQ39CpX9QOZ479BCFEAzsbR3UV0rKi8qCVWlF4Eugqfkpc1D5WFQgOIcU2UDp
C6dg+sScIX/CcEZh59H3P1H+jfC81IpPRTzFTcvavKisM9HgVzHItOntyatErjYySZJ5qIJnx/gT
ApgMayFbRhg0INmzvaXOsJ92XXlMUZrSvEs3LEOIuSx+eiI/iVqe/83SSTMGuj1yvJe/HUR9OqNp
TFLNCQGnb9NJJxa+6dbsCg8GZqNo6EhwJfZYD6kdrr0I+8xWern29Wc4sRzavgXTKDt6RNGVTxqB
JTJKDNt2UwsBC1pF76WNUvbTl0mFvragpWIrm8hxULKsNbq8WS9ymbBW+hbEDmiCviW5rXtJyKfV
fchXK0EXCfVb6RO1OG5Sng0iRIOWf5+pPXEpoVFiDiM4pRqkdQCzOkVh6+2CGoW+6nqabUOjyoO9
chukqTAU71Ukj+QmhLWzx/lXS9wPC5FDHGuslH8cSnQ80W78czqY7TENK+08k1f5yDTljqdxI4zs
GJYZNLdokrk9UfaH7eyDm1D2NR8GR4Q/6XkZ7sHa5OzXYQhMJsjNS6cXXMSZsEL/RWzhJobzHuha
yRIZxK6k5Ht4HlRKKQbfdJi2oOBXv1b5QJx/hHyxAiN3cDS88TOqdKKc5Fc1OrvvyCgcFYgrKdSm
ZgLqWjkMxh3LzZ/B6vUpiLuYsD+bZuLheClYx9bhmRjZCvqCmcZbpM9Gr341512sCJL2x4J1s4iW
kvSsBGxQL77Cfx3jRHoQjKyw+2+ebw4Hgc+0dgana4aVzQSR1gtK69L+/miYNHnSYWwUj8EN6ncO
MtLv+3CiLXfmvpkTuH50cQrhQac/nB4uL7sn9XYDtmhsSe+wTv55NBV8hLMPGwxSLlkeWoQo2qa2
Pvn6cjKCZ+iQZSciWAJsThv+kIZtzuhpWWSaKyJ97A89ok+Y9HS3lX/XsrptWohRTIY+wrsS90co
PZWSjWVTm8WZ6gEXuz3NVya+FrNkE6Bsl6A+m51NlFusAJiC++bNXdRAIGcMdNcyPYkhKsa89nA4
c64VfCvvF8Kmf1/zz+Plr02twdgzlCrJIhOQ/4xhrptGjq6rokvx3w6qlqQDFw1FXIf7i98/8I+0
8r7AWVpfnsZmgdEb4Jxd4hpWPk2ztxuXMEGZbL7ON8RfxLHqC3KfIraUrjTQabN4+FaDenMo1+1T
A/6s8op4+tKtFfnA9VQn4EmZG4zA2e0rrAjUHvUQi3AjLcn1XLYRx/CFL5kqm4HvcL+Hp0/fYGIr
dLqWsP3Sz2oaErrQWRhrM3aHs4sFhD2Gbt7yFpRguGBLPJPB1FxEOLNrtdtrO9ridfKyoRSjWuwm
6qsTsNWebakdSxCi7jekB3AgY0yVsINGqKfwzP4Ca/KbbvzS3wa8UKttWUuEV9YXknfkfqFQbDwk
C1kWxQOj389EvH3CyHyel8YA2kSqC6FjiAB5HZOjPujC9TbGjRQDrT9xBpnU4mSaW8hgTC+H4IDS
ONI+3A3KuWiMZPFUxsK+rRf/MowUITjllLp67mJTOdGuB7cDjP9/1MP/msiMJZgWBLm/UrFSU7D3
oX+w4t1TC6Pcm4HmXkwoU2ujHRwqigsDc2LD9ngdebYtwIq7r6GSajJFrxRftcn8EnNumLisCSQt
u/pTEx6hY9bAF3gyd6MLU/tHA/ZWcQWBkf/wbcou7z0WnHCDUAhflnZhkbCjbzPhk4SQabA1jgBk
Airvevjn3hLxyX9oGe9tyjZXoj56lib92GejF63oRMbIwqrLl20NjwmXENWFgSfUNByoc7syR9Ub
hgvTSVcILl8UDRlzOf/5D8z8d+mUqe3cC1MxxAyg6pVYVfz97ac6d5PIzlWgjPv9fENXcBTTqts6
uBPd8e6dPrmVmxWvNfnegUqI6OefbNiEAMHscMDkna7r/oQc7fzSqDg7IY5emdHHu+hZog3yZr2y
+VSgDfmAoQUNgAW/Z0vwzhT5kwKj6+2VLPrqgvuwgHqj3CP0CKIfMrTIjbn4dp2Wrt9d5jQBAgfi
Q3pK4hV4RRwuRRPCH96PFOn5bZwC/gU2bOHrAiY9lBtJMCUba0ZGpKhzQ9TEyuG2Qq8ngtVNaLWD
BzIx/rLKQlHBh0HrAcDYdLOhrmwr4nNUhrjPqEehhtQ8DEaxX1kcSkLiCTpXbSYlQDNMuxTYMNiC
zmxUllrLdTWwmc6OLtf+Y20PDSXQyrKrHEswuS4bGWFaD9uor4Hd+FQVVu+QqYWsZSc/Fl31pmW8
qjYNfRChaYDMT0j/4D1hWGp7F0o9/XwR7CcveyR65thHE389/ztFwpwMReQYMvOOv+kqz6ugMfb0
DhfzVutEBVGqRHhs1FIiJZPd/LX8bhnAgPmlhys38EQdUmCuJIA+6H/RqMNVrHC0bSQO9xDexRqC
HVJUMdJVytdNrZGXl2IvolvNYr85iZB2fERg2E5WisOyhNi7kpQD+07pCO1s8S2WfMtEcErxYud7
v5Dcng8zNS1GvT6ydE4S4ahSBZNi5v52Rq+Q6Y9AC9QUKpe5pJMnMuMlx0AdYOG3/ZiwX5SE9u9J
fJ3jRG1aSXSKSe8cUSzL8F06Cr/LDdCDCg77y9Nb+kOIvmHVanyFJ8YhhBcCnjSQVee4+UvB4rVH
DInzWVHMt7JCc0FLgmZPwqoRNUzg9mm3iiczXk/02aUoLQ9u5wOqHbW44PhNVxWgmZMdRzjNnB72
enakqK++6OD0vn8Ae1uuD8Pzr/u7tOALjyuAZrUjSYCaNtlQ9jTsvxqSpoAgAf0Tf+sxeNjDGsua
jtTP/a58+YvT3M7PeBvk4RvsWNSDa+snHMtKYrlq4mW5G8x4/wmZDVhL27gCbUepkncEJbBmUmRC
Z3wwEBIbLIGS00hoHa8dF1tPFyB0tlgQLICq3mLDyX/OMn3uN9CD1XpCItlM7AOhbP83P6J+lRHT
W042A1X2rkT33Oo9X7xZ71VNFYL0RNaEUghbMnIJ0fU+Vk2JOpVHUr9i2FnJTXiV9Wo2hx1SUqWR
iKTWMbp3U0rR1HfU3MgViEsZhYrU0jrNLBh3FR/fmpMwvfYqgQiIZer5MtJMT9TlskSMdvvpa/C1
PsQN/0GJ7q6IhMPtSaDkY4ZV7CXHN1nRdJ0rat2vPW9d1dYWfAGDcsOIGkc/voPOxNfq/PVt684I
O3mGVaVKUGEDMX6EhNWyv/WmT+f5v4zTBTt2zbP2/ZQyHAMIGoYAT0yrUlNOENJgrwxze0RzW37A
RK89dMihWh5Gjc4O/ENmaNiK1co6FKIJythPHRNDxzHhcHcpF22BXE+bxpT55PvcHOQGLjKOVjTy
nzmuiDk/X7UupY2qRhJKt6ObgayyvwvSHADUs4KPzYDVaKcItKK2ebLeMVL9E4TK7OQeoF+U8BAz
QWyh5xi1waamyvYcuSum0QKoiVAuGRRw2kTn6F439eqITdMmT/OgB7Ol6yHVzWluOHBSlG7lxIvl
vTVmEow0jsalmmB2GNqHHR6GZ4xpr5jLaEJWoTDr+skOcvypS8IOPNTfkh1nmTqXn6vRfV6i8bNn
15e3wje6Icz02O+eW9WS+20CeZACt7ilQ004/w6yZT48plrBAFQdO2YraaEUnqsh8JQQCe0eVsa/
UIcRK+nnRajCrWZWsQTGCL+W/PPbC9t1PApFALzK8fE6Q29YvbY2tknkZCqxis6wsJE2Jj6K1Yep
1IE61V8+/SPfciUfo3asdkpg/03qrygJ3BHnqBEiIHoDTGT6fAwTW01WAFFhxdqrH4eWZNukOf92
wu83yUJvwVS783Z2jT+2wGbHIHG0I8DUQwI+B8ejNc6mMgAYUDzP3fxg76JWBnayZQU8ngokhHi8
i9VBfRsybvbm5lH32wCLGBDrNn38vpYVrwTMw77oytRpgCiRWuQ6opijubzAARnUX9VkFpNdxgIl
+A5P0QUf2MiloZMjoiSOXKvTKIBjQCs5zQMUhqcbDfTk91oLqdzWL/JWYrxjAewaaJBRQV0BHGW2
+YV4bQJbthEhN5tJddtz+gWzeHbrXAkM17F6qqdZuNO/1eiszYWJQa1mwL3CPi1IcReJcBUQTID/
hc058F6zoaGLUc5iltmn9aowQCne4BMfh4wqloz8IfTrOgLlmjiu8dFi7o4PVaIgif5H1RRobW6K
cW0uGCUf+Fku3rtd5hRahpQD6DZKw21mAQRfU8JyI75YZCp7hP3exXPx6EyOmVWmfSMZHo+pYxU7
bvD+WwdGJcN2Rm380mZyvOX5OMJ8YgtxeosEjM9n+6/xOOmHR+N3VOdWwxghddRq11XXbzqDeN+w
wiiXL1plyDQKVVPBEUbXCKfSn66PVCAloYbfReqH6PAS7NJ6/BOqx6+I+DIR1NSz5lbg7qwN3Vn8
Q90UM17gTMrEFLpo31fi1VUQZW2FnFqVHsVHEJGLd5D+23pRzD60USGTuvwC85n/N4MsyNUgmmHh
FcsGqNfpwqBxZ5IFbNTV2sqg6iH9levVkJ4VhQxJ26jL9DpSXIgxZtnM00w9kY+6wJZ1YdqFPOF1
ezemNJ9faEViT1OKJKwhYoxRs0OQ2cngY8wL8dQ/zQ3I+5NQQiW2T8D2SvULrWJKsOaPGQsNKnAU
JvyC1UfayqoyHIJ/dQ8bPzRAyJRasoEf5TfKhuHlRY4DKXKZ9ec/UKotvGOrVxalJ+mtbYZG//gD
Kb2f6g3AvsYGAyh/ujdIl8AOpkKHvcLKH9XzwynJjyzbfoWlLRXLzLu2QdiZjWcMJ/9GdgWKTCty
9SSChzVLFPTZaHDvtMlBTnQNpEbGZxWnCFX3feNPY1pvdfKd6lioV/i79JnZz7GM/iOTj36aFqXd
UjfoMYC3r3Bfelgm+WbTssuboNleNpxMwJFAYM2CUHxNw+p6FKqaTMOg8NtRXifS3T9n6lVz+CM9
SHg9yk+yIpEdPyRNIxPLU/4Ne3Q5bO9g5mQr3DAn4jmLFyFi2wlh169i+Yr7puBabsLrZbzLTKT5
dHgLuwrBW68wJIodzkJSGnNs2nholvF2wsCGS+HsnceuCo2fVCQlKTUMJd5xh5KMey6dme9jysdb
6CyPFR9K8IdyoiQXb5KN6tRiFXCXA6xMrOCQKnclBv6i+2WqtsQcVTMDYH2THan5bb8nUkmftkIW
Cu58TXfyYfVViQdD+medswAb1wLY0Uvr9N7eA01n+8yjaRW4rUKa8hmcRXo8QO2ts/Cr9PLmofVv
u8Iu6ih4pe7YQ11dV5gGgttdf8vvnCQ65Hd0lm2cXdO3e/o3/j+FxL8pCMguUeqbPXGimkLznN8K
EiiCg3PLPYWCFKMYmxCw/9myoAWZyOaIbDKSVoiXgp8DkuAFYvT8FRMh6s7aGw8eAT0TlV3+Z8Xf
xHhFI9KPlzxFSSraZEbcCdA9gB9eDSywx6Ck1MUr/bpmJjiMj3P0NksojvdI/aAWM/ztTHjFuxBS
DlFbU5WccLo12cPPWET8ql4l3yUFBAYVkdoEAejxlMI2DLiXuxMVxcI628bc5MhozLpDcap4ECuJ
cxd7vRTmDaTdWppknHQa2sxeg8tbXmu+XV8StsE40JjeuCIAFrNoe/tNwHsVZ+bpKbkgKssZ09W4
wK89v9d6CixdlNsU67brYxRwuV863Tg9MNWvjGhLAXsKrpbAJH0gVHOEeypDozfIfXUklNPwj4IZ
XA7mar+j7oTHYO7abIMfN3iRIac8T90/egNQQG9C8jmEnfj04Ait5ueId+dUwnSvDOXttckWvfnB
wZI1fzYflaS+U6NS+gVXjM24mK6UqjdFk+vJqU92rno8tJChS0WUuRsA8MDaLxzm+m8UVqfoAn6+
Ha2e+PjsUO3zVqkI/p77UHHLTfCBPQoxDlpfo+RTNlTY4GiFb70j+ApGyCN6MDJ0J1fXp4L22y0B
TNSvU1rvWUfu1O0fc40DEPrlsUAWTqAZvGaCEhCINf6jtxfv1WU46gHYsKmPuGoPrjGa6b3yxU4t
FhQq2dHVUTzbUJt7gsVk0SBdwb6jGlXkL12549slW7d7pn2Ug8GSjzvgQSTM1EMuRD1VMUK4krWd
BF+3UhmuRtC9IRzh5xi7oLzON85rBPnuISzjLcxux3DuTBa1pRUP98DVkvAb2lmTVk1XkT+V1lRw
LsxzmA4kZqpliOtYAolPVnMnlqZ/JpK1SziEL9EJqXkzKwbSS9J/ixAppwbO82atMFPdv5srpZMJ
2jX4BYfC47trmbsbL+FaX1fK+aN6dJDz8u4PcpJrDDDd8/qy5uvauYoyevZ5aZAlpMZ48TVK0ds6
JJ50hcRnCZfUQnd48bpoZ1y+lJYgMM7+Aettrg8BL9FUNJfAHe/6ucN9onIMscBPZGziiy9C7EBj
YcnWZmnIJnYR5bXCedaTaSrhLqnv+2P4kXUM2Y69T8pVP0imu6ZvB2dIM03CVzb7jFXJq3UdVhTy
nwPMPfK3cHZQwlFL5ilvgcl20Fwix9o3avHg1UKYG6wVIa5/RGg411+fIgkDFNQW5uVrZFTblvS7
t4q/XbFu1wVZ8HX1FGUPWSRaYWJJNIQOsb88vqDyv8L8Ei2GeDoPkU0gM1CL6I1wX/1OFgTHI67i
6/ELjhk37Aw5FZ79TbMS3KKExG+pKZ4Pw6c02wanGRCEmq0eqzsiIRU364eQHtSXwvZbssRw6bX6
yNAUFiZdm1LYg+xPefLYvOzAf7rwhM7E70DOYVQKAv6m/PwEsW+59juQ/FeYJSaGKOiLlvI8ZSIk
Fc17YJBMZknj8gKK9r1f9xoOlQ1A/4CpAhs3RGIMm150gtvXpM6WQYPOGNrRTZ8A8+vD53MZizoC
ewHgSNZaCivljT3qb+aaQjMcwY2LhbIwpDYpJRAhNqnZXMGDDXZlutcA8ctnn5Pmaeff31Y2ABXL
8nFU/fUAEZp11F5Ylxerw6Myez3cDuevt4oR1tmKYdwrTXAqAkkQR0Q/5lquweE0F1FKZ9draFfe
W1LN9apdfS0MQDOaSvylS/1MSgF/WCQxZkdfr563ZvTZ30EpFyFgjx/xHeOgcsXEY60fihpIzEUW
u6MXhAo/k84/fDgC7dEE+S7f6YOUJMbRPr4wS6HFi9OKx/H5cs0r4htEq0VGYhDNBcJH+H8uGC8A
TE161thB4Hqk/rf1usySFOHe8lzY6Saq8oXhBcYbGRuTnuLPS7M62X2nJP8AzvZFMdtbk/X8ILqW
hyKJTxU97gg9c59EOTvwZClx1Kt2bB8SVWGuJplUeijGwND2CgOApjdcxP7qafKUPDIF5AegXKD7
tU1uM6f0TAATA5o0ggq5tVITokWiij3ti0ksz8TDJGVUsWAeRvG8cdagHOuZsfwJUuHxJskiVHZD
N/RJxRHSeGDsl6XkDQSMfONKagAvmNmYTK2/B1UIilJIAdOgX2zYQIgwZ7mwnbHIuUvxiRmhbXrc
r9biRLp1Ym/b0bLLe0FUV03INHAw9nQzp3R/LGyX9u4/i/YXP25sWbirs5WjD7Txj4Q492K7AwGS
vwG9d9puB+aOsU2wl+hmcgRYLUoX+r0AGurPD75VESHCP2c3Yp2EA1TqzgQLd6nb9KeFA5kdbOaC
GEbDuhoRJfGmgBwFsJMY3CJQLgCwFybeOChBC7jSBJZ11zueCfJeTc8Bwoak11k25jXsMjSIS46U
XG073wW8wY/J8/YI2RlSId/D8jpiWOb4z4drIbrEnAjSEnAR5mFRS82c/dWKfufVp45//gh+7YzI
cvNVpZz9M9sNaMyRMAhlQXmsnZYQWGGOra8HWu0TFscGjVZKCXXOzNs1Vowrz4+3RlmjvF3r3AaU
bzD6vHnDesMs4I8gZHZLi3w63umb1psUp/y47tfd0Z2WPHXqlZM8h4iLIqjiTA9DNiA17fNna+nP
SgYJZSxFB/kjU+NXHY7Xqg1K0srcBCsdvjOKOqTXvuxuOJsDCQ+teG+9yCy77pZrqCCrmKkws4wE
PgpOKYalBkAVClTf7JG2+DgYwLc+Kdd4GB02Oh87XvBwrh+CDsg/pmSTSIvQQzRuRhEiNzu7iCU2
wQB3OgdU4OVthN1wCZftfqKaLYbWCRDUQRkIS3UVHGzoTJQtlDKfuFMhd0arr266+hPUPvH1VJZ5
HrclBAqgFuixmFrO7Oz0DAKKHVPXm7USSxccU2E952S+vbzeYxuIi3tphMbnwNjd0oJT6g93hnnr
pCMSjW9QMqMv5fWpO7ulqqzmqb+tVwBEocKUqbk16wycWwNy7DIA0RLMYmATu4AexA3vN1CdcqRL
1Opqe4Oe7uoPZ5bo7GFKEr/WrG9bKGz18fSYa1R/1k9Ml3cIrx+5NdIi/JIq4ial0ukcu/va/vth
7voLKPJmiHC1AZcftIqowErjD5c38aJBWCC7G2HhghrWKQT8+MTKtHF+vqXsw3vcM5rIx9O3xPQt
UlPIM1w++LtfHRsKnnHR6MEj7MU+rIcjvsnOFdNYQVCDSpIwOX9YvhV53Ocb+Yj3arJTYFkJk7K6
7kLTA8PW6Vt9xiGguv2InrU2HazhcbaxfIebqcEt04t9uuGSKMeli2nkODigpsCQyF3UXtgAosYJ
bPyA07WBW8gDKJreNDZTE5JQZIz24oV51WSzOHGEIwB04N7WcHwYkU13kuo9SD0/YGFmCKqRrZGY
T6lGzLkNVpKCy0HyDBF0HAC88AnlWLEJCjcccGNJkouXgZcwbSINQuxXha2DpH+oknevDpImULhM
epOvqARiT8jZwb2dIUiiQ6X519sHfVuNx9BG9KoC3VNDbAFFxuvg2l/JO8shcQo26g4b1617mUrE
+dmmK/CqnstS+8EOzFrTNhH0FoeP3HAp4i4Tv0AH43VTqE9yYn5xtGeh0KgJW/4oiUMExPstimBo
A753XoTDjbCGx3xhilnhdCn8ZXHYUU9YdjzMDpE/kZvgc3/CJ06gBw31QZ7aphKOReN28VBgkseN
WD/u73BlFCrRmbIXgjl472twYkbJUChHp5asGwNaKquPBmw3irc8rY2eBVkZhsJdZq2JKvI4Vttq
BIJdj4pvQ/E5fqV5xNTxrurg9G9Ac3ZQAU8/RW4RRXW2Oj99nTP9AKjf5IXeQx8YIwKN/yLXSnE4
HRwqrGymNT/h+OTE0J6tK2wALD1jiLZlOdQDb4wLy++2JfCWfJ9lstwZJ0Ezs7niEArqUtv0Qy1Q
JfjP/VaO/zThEbnUY7qAxwGTk9+D/uqNyETeLMB+uzDwTjg+Si8dlKSsIakWrQ8HPo5aBTFoqVK8
o1zW3/kb/c6jhjHKPOvqKNp6DlBcBTrsuwF+JfMep7+0PtiHs7fVSbgWR5sLFfaZeAqrP2NO1u54
bds4XALX2SXaTep5etVjvyxU2izMFbPsXXz3zLzUDLP4gDcdQ5AJm2dNDZGBlyVIf5WYOVYq5I7s
40njriaaImDgBT0EesytXImwSuB+lbpkwfyNo41gQeeWmYMRJwcXGCh+6emk/e0LYub+6bT1+8HZ
YpZ0VG8YS/FrRIJHUBbcOQ6K9hFy3Di0P5TMABd8+qRRxGc+kx9PEFQpea2RQGexJwZmrAZy6yUE
8Kq6Z2aIYHjNh2/2rq9V04RGS4ZIXExkVAZN27zkOB2npB9FjwLzHHVq+m/AkJOvNvyfAIbDW1mt
XedPaLUXnAc3Vppn8gamggdoFZhL8VRz8UG739JkPNPMHxbViLr4wX13urHblgBkClW8Ey3ciHt9
hOMlsSlvnpdWn+nWwKDLrnnyEjJ/+DlZboL/+XWrrquxV31I6wXau59xmrPMuMinKU5+7U4BfP19
ACgUJZyqW5wqsViXH88Pr9Y7aRQZ1iG62CRfsBY2LXA+y7Rg/xAOA6Ly9qqze3u9D93K1mo+cxCl
aRCbF1A3t4xrfC47g8BS8kVb2QHNAfvcIkXTvnI2tongZwKc/ZIHFovUvSWT38m2n+U6mIlSf8QM
i/7ZlJH8apVTms2cdoFqWPpGPWgBViYIc4d1gqijsMs2P+lw2lAdB39sl0rHCLCQUhv/fQA3kn5h
5nxIg5tKvCJ7WErcVBloVvrEpuIWhQa1IgBevM07oGYznToHBrilYERMt1Mq1HWri+yq2AXTMayA
gSd8BpsByom+59tWLTe6kGG4MsMJez4p4cqdzg5qcP4EcA9ljOR6VjzGxjiESiNnQy/JEudJHmFz
jBxOCCzyN5dmGAeRFwyOKWRgezk9DLA3SoCdfq1RRlJgJwtPlOscYrMsqVFZe/u/0KgTtA15qzJf
F5d6t0WwTBk8DeCT3uoS0XbZc9tKiyO9WoXcU2zXG31z7hSsQ1yKtdCnGmh52F9wcmxfxYI89aRK
tjwkAUbMILFAYBukiT+xeqy3zBJt5KrJHX6tCWPvPhG85EDvYsuctjn3wHGomSPQRv57S5vOytUF
HBQA0Au2+rcr35nTTUY4Bs6eOUu6dW2DgGFuon+bZ0E0NcYqtyPj/VLRdGeuq8y8hERV3el2x6vw
9zGFFSV+4N2ItzV8cukjGc/7DA1rtZY4lMqGA7Ez8ggrIl2peJwPK9gQZlp6RYl621UP2Cb1mXVR
sMsaqtyVOGNJP6D+suswg/GhwvVnMuqSwgSOHkLxjJjovfBZFfbiIOW4Dn/nTZypQ1I51ICCxiIN
qAUr0lPEahN9QovzHLksO9+ekpEKPCiPcI5DsJ91DRbUFMQiqCoEwjQRjorM1rDXcLwa4UzqqylB
HkVfazSXZTpNcIXsTXfsw1VrCkCrgQVbzaq3OMGnf0D7Yc7SgO6e2aTrSak4+z743KVYtnUA+0lO
2IOZ7tF2AfHfefuPuj9+TOuL752ZfBezZ/5AsOuupyYofg4j7aRsve8xGkWmRhW/BSZk0G9dnO+b
h48woAtiMCYwsFbkT1oXWYSlLtj/X0fBY+P1dSOtVqQ+bupOr+yqWI4dewYD00nSRFsv8QTsaYe4
l9KJ1F8VE5DixWBrZhkYknBd+m7WcjJY/rTWw79Z4P+iobODjb+R3cTb8JkbfavZe71YOyOS3ioB
kiRAFq3ukEm6eE2pFv8nj2AGaQDXI7xkzuuDJ+bLPzE5IWPxg43P5pZfIjkc+bKnfGq7nFHtmzmE
prIgWw76f/Ytet77Wc252aRiF4lblHMHgHNpqHxgi7RJI+qx22xycbQYxFFGGrT8Rp3iRw5d4CpE
+41ED1xEuQjmCDQoTN7UAy8GsmSVlOkK22u9HJ8A4vB/wDnC7J6WttrsZbOtlUfXiEF3gE0Rkc8g
V6C//j/cgUqQ+/+SThDV494AnU2wWFPSSHi++bZQcPpJ/+2KIvr8xpWeEHkxqvrB9M9iNEpzJLdg
jr49rhYCgHdz5szswkNgl2yswQHnRF23ZWcq6JWaMnEHjt8zgvgv4P5EjTH+JoBK/Zf3t+S1VdWL
dx/D/0ym8WBqEvxGzNpArtZsAMV5EiDhZdS/V6/2y4tdX1Olpb+9QYRaxDi6p/CKc+8E92h1tSU9
XLxDZFIkRt0Fmg7Yum1l/MPZDFa4YYWJIkQbSAm4BguLQzFZllsTXc2/bGUM9RaH163639oAyXtB
hV4+Nve9gBSyuOnNagk4zgOLIW7tHIB5V2XfmLc+iASZzPeIdSOr3cXDlos2B5Edj/5FTP5mPkxq
rBguhnApSXv93OEWYYKXYHlsCVetUGLuX1aLhwKiPqUDWEi4KgmAJBYstHZH2Ow+XB2wg2n5btEZ
ShUG1Q8AVcEZdnJFw2aQfAEjJ53l/URd8bmmNF8EsfgyUkTrwW5Vc2/IDWY6rfGqaJGqVUaN96yV
oP36dr0uzREcY659AFZwzhT/mdijaoWwyMuOJtW/ssLDLl6xXkRqZE7CFFcpiOqRMqozU0Gw8Uem
51A9webxl9HGCJZ8xFBhnWpNI8RLyN2+90T+5Fatujw7d/sJlNEiOfle/lNmCJ74a+F9jkE/OaMa
qaUyAEpMdNp+nCnmd6DyXNuthz2dEkjAnJAJkewE7UYU1Rldly/J+L3LmF1tu2vlUvrDWd6THy9C
UCXOdd9vK+82GqxYyu2eI6yGo4NtPAXgVNbPJGyAK8yy4XefhnZWUmqsvaxDRsErMPdsIRYXYrYX
9pLXxoXq2J5IsYxhXU86bGjjZlKrvfoYIN/XY7RzSRoc4ARDCs24A94eW5es45r9aTwNeOsWxptM
8uS2aXml3XBEzmFLhiqNXTZ9FiDcS06k33fphE9b3v1oftbPcPuSQ2f2zaUSyzPjJOPagWqCb4DR
ZGqMp5v8CUPzxkjz2Zvb15ofJBRKhT706eGGjhSXnJ8s03ixBQna7h5LrfscxZQXcHrG30To3ibZ
nYpwj1FEp0PdFHKv3AIRVgR5x6YAY67DRASeoyF/yCgMy/mDhxPhV/3F0FosmkojYDSe/HGvl0ji
I3vCZ4SfRJ0p7MyQS7pcV4K6BpdMSIBSxWr3ZPdVxbeoQvJF4uLI6gx7AJjrobPXn6UwIVaivQ0U
fCT/RvEf2SO8ZIvDvch5h8FJx8IGU4K9j2cHUcAihKIZrKRh5ypTMHu/7p6xuA8IlL3iUF/7rACh
v2F2vW6Wp55cwG3jkWYRa7N93TXFkaO6xhaCewHWguyTwlViaFWHgAdyzRzEj5X2PHKImIMAoL5x
of6/UvFIwb2S7pC0/mnurHcyAKH1HVQm/4Kr3rD70GVAgkH83qBZ/BLr24Oc63ttlJ1AAHGzu5Yb
ZlyrxF2uJ9MQFpevQ6oxIVU/WBhXUj4h5pvY/Y9hIw0YfgvV2Crx44SfBXqlNd9P8D8b9hU6mzxx
50IJs5VOpAHBSEGB33J0o5nnSCOsGOcnXLkBH/JQu/JK96LMPqn4ute9f6rxQsBijqPDUjbDEFJa
Lfd2gW6SFNnX2dTsG05V1++jvp8fseldaMgPTgx1JeO0/bIZ5XotihYhJnFONuZvHvadofsj598B
wAiw3KnYAL5Sylsam2qPM4Pc2rGtDRP/WA29gqxPSt3keDenzwXl8VhvqOz9h9DwiOGQzVLo0Yob
cpVWR9GBsTBywjkzf+0oLag4FInVebLXrXtanSF/IpxazdWqeO0RUKYWFUTFo0sxycxxib8I96Yn
SjZel2w+IV7sC9QhhYAzBG5ErVdjEVlRJrgR2a9TjQnHW6AGH9E0SQ6ZgkXqfIZauB4OT6r81qEr
dWmYVsqlpLwtjAAegnh+AK9PPdY+7v2KoDLyzNoZMZgTM8tWVDqYIe9U0usXfe6aqWIxpF7bCZdB
Lm+pTBT52NlOFMk0fRiCjlYrnqVO9M+Ke/l0hVg9CPg0b5FO7eSiy5tVDnvcrvxLZ3sCtNZGxQWI
/VDHSXQTzl8r3RxwaDKBeEHDhlUKnSEbKOdfYw8nMnY/TumSM9fksjY09ZdL4O/OENrqGV1EQ3Lg
IcyQjjzQ59+zKppfeXmpY3WgQw7pGIolk4x+r91gA7KRT1DVKApfWAca03yPEsCr3l6rK4kw92X0
0bP4kYhYPpq8GArU5rk6/oBd+3XHky38jckbwEbSxS1p9fJ6DVzCa1hNERn90Ypfp8OJF4efqKi7
OhOHf/YfVVUCL9eo6pcwcgDmCWGZ2fjx3zicnOUIp2GcSPPh7661CwdBFAZ6/OdaJ/MkNKzhBnHs
BARZJh8NvhONpvYcMYHx7aFzg4GR7ij6MrslJy2HOKY8dgfNe06ufUQoOHeMmMJdwjLO0YH6cNwm
lmdK+U0InBpVvzjwYr1G+qg+oAZxqmLDWr/1r9qS3kE4ClxzOQ6v9TWprIaiosytHzx/PJIr8PLt
4vor0lffVDJu5NlmbTkpsijCaI7GHUbtXTwQJ0iV8ETSWvaHgA2N6chAZTL9zJluCM5JdGiadRLp
qGEp47NjtILmm5ONkQ/H0GpWU9/UkSOCwgNZJK1oC7HSm10eM9AVSzMfDXZMJR2CBrSl70JPQdRa
p4nkx68hIGol3lF2Yd1/FaaQFVUe2HaqeIYaBhgkA6kAvkYab2EHBqAXQwizy01WuE4z+6onusb7
HJcbc2HbsMNNxUPXl6ttTWMMVRu6YjAMkjxv/5LNq9XSOwTnv1NWo3xP34JvHd3mkEQKxyHNcNep
ZaAEr3zSfxdYuZlU+seb5J8/XU5W0ianpSUy3I0YKjlexImH8G0q4NpFI9olqUCziSnBdkRCRJko
XL6rMnlNnLsXGwdhOFZo6+ZXtDODz/0okX0zmvtu5Y8VVv0/PUNCUmwuhWJ4F7cWyDiqHICMpAO4
7q/YK/yXxkNXxMR/K80qdQoNrsppEsbN4jldiep4Bs5kBaMwCOdRJ3Wbp26KosMnZH5Z06f211v8
q6jqLnaeTcrPhxTK4ztDrbP+Xe5dSlH7MNhCjaL++p+67ecIyFZcmqjyRTPWCPkKGEBr1U6+3B35
vrzuuoSspgDpHPaBCE0qY+jSb7+V/vrMQ0qfnnaL60H+KQtqCMuR8essGsUmDNB+T7nCZebCajQW
GQRBo8MmvNvodGUroxD9PRK6mf03N92XZXNVv4VrzLifg7X5JzqevH7tw+INhYUCFSFcx+zr0L0r
d4PcLRvfjchgF+mrSWa1tQf6RCzzNwPzYvAicZ1gSDF77AZ3eDMhfSlc1g35ZTbRzKZ+0aH9mR5Q
udqu6sCky1yEcKdRJTQk1OJ9zitiMECtpn/QfhLNih10kfnpDWbQEnSHt66FSnF33hLjBXQG6lCb
PX5uPSNDtcr+V5mkEUI7l9xMcDeS6sSowBmZlWJIUZLukNhtXLB/0akCBgyWkQaXBi66L/xtjios
pDevoPc0GBX6x9PPTlPMBimkDEYJ+z8LA9LaShYh+mnPA5UuH29IjDlKYi1Cm7EAf1OK4y5rS5Z+
j/LIJ1p2v6omfT50vnbWENHpeH4aTtWPGDZm9qYbVNT9l1zwHmVrNv/VAXLO+ePZ58VoQlup+up4
RXH5BeasWRz4DWShk7lH6AZBqP1r8PEtWtGIJqP0f4GNZW+fnd698nLBHM2/cQ8lp2AECrO/09Zi
1TQpJ2sIaIVFT0LlLMv9xGguqN6nse2Ffioc5NeHO2kqbK9rYuG2pXT3ZqMsmJntBaEgmdqvNcJy
fbtuKuQtCRq/BGQH01G0DB1q68eG+NCI/uaqLPRWpmpSM3eSAF2aqsK8Xncc4hn3bi+Nbat3/Id1
FUjkj7klkm3iqy9MJF5NK09Y70e0pwtRe4O2V6ZVDBYlNhwMn85gjKjaLbQluCYU4TH4w++g78O7
O9f/J2ZCae3MVoSBtWtP3v0kCp+BML0PR6U6Wnv8ucYVS5zUVGbRqO1QKXqerzpvJYKFGxf7nu51
kzP51W0kGfMIyFbKVmkgF3S/ZHgqVMZeJh0QzaP5Wyrh32Rq8c9cWn5ff7Y4Az7r8+uNsMhMo9Rw
2ULccTajzw0NiF757BKHRG2ho/Jz3LkiYFOY+T1MlUBf8lmbPnoPXkCQ9y46qJxzY3EEWMaQOFUP
Tv5ySLN/G5gEFoQgj/Y7QU0Mcjshma1BFHJFRcqwZCJmb7ib1eVukw/UjNdjQeSF3pafCTZB++mS
kk0Y0xJ/HREpSLHY8ut7NZ4b8yVhYYNTs321qe52dP251NAHWCmh1V0Knz5BAVccfrTjw9MweKQR
d8MVSP2ivQWLw1smpYCuEc41uz4o1UgWiXHf/pHl1u7YIMsFaBEHkgEMsOwHWwnCmWW+/rUO1/ma
rdI8Y7ZkHADgAwXFN87nO9afJrTna7cInnffd/9Z9pLrRWO/SOjlb5dfXGPMBA95vfC9IR1QjTY+
htjw3WfZ10C/w40ZB8cQ/IFVCFZNgrkRdzDszPcJTYa6qMj1c9OTXtteQPvdYmjEno8esNJz8ZeU
fyTQAIr/H4ZrzESA8ncuMpdNSzZHsgo5Uf4nZ94TqR8cnx3G7UvGpxenSk8yU7faxYLm1L2l5LiF
ZMTPscTFOKuVRQ3ZzeQgBqJE5nyYGPK7JQIt4qg9SNR+ULSIL69oZAniNDYq19LWl6y7DxhdZ8Xg
0hoh1EQJVcUlvto/QLJdJCb9/eF1VHl85G43NuN/e9vxD4qANOi+zCcpfllcCZIysw0O+YcQU15j
m+NmJ/CdjTUy49yElkKPT5zsrQLZGH7N78pArjJWt6RWHoCwl0YY3YUchu8/kqmbagvebTtGs67g
RtU049iG3ZfmtIXm0yYfLmPL482UAcfazb8kqhf5mnvKxBDqq3OTwuQfvqkC/Vpo6cqPJRsVeBnu
Pn+1POTOuiGRIYXhT+s7pdZzEv2mR/j9oCrZpzzaypzjawJb2IKC+Ojaryb1BvCQPJTmji/Hdf1j
c0u2pDvQ9pKTKKvm2Cm80YDat28MrdU6RtTjPHpfptT4z0CaSRXAE1ZJtRt8FruH4V4vLwG3Tx9U
2SAarZNlzx34EShtSG/Bo8MV1DTbtMBirOZrbB22oEsrJGK7mxY6WmQl1+KsNNfJnHIsOTCcEEbn
B2lGl4eOnwJke718D74OyhXt26vXSktHuu4c5SUUS7zGbKdxVBkzrvLSlRB0PBLiNQNZ2zTD628Y
wME2LU8IiA32rHz0/4gOVpaJudQtha8/eDkaZj1AV5mN2KNJ0UPFHXyCbzSDJlQOd4+6pwnizlCk
rQVxZcb5ZduZgKapNfXNmP3uMiEv+GiJeWgZ0BkBnCaFl4NjAnGRPtMDLU4s845HBF0J9wfxW5Yp
nWQ8rH0eNnpECezIl0TJpUqc/XJHMwHANNBpqLHugVQFXoOjDotTbDOTUU1JesJvnVt80xiRJ+Cd
TqaH4M2Y9MNWM/392fgi54GsoQDAMvKHQuv7Wh0yXnOFqc/MYaAHx8eAFglNpCcBQJybgTHWLAnq
eYzSSUrMaKZSaEcpuZhtkGnIbkWqvuGqqKNhNMS5Oab1KC4+2Oe3kOa6h8WVlgl7OhMWesWYUceH
6dlvE3+7DE01zRKrWC8soaBUgVSK3yWHqDk9bZDoP4lNxyMT/awjZFveFx4pFwruKShrPiLaTn6d
6iGcfGy+5ND78iZVjhNA7Dln3iP7zBFHCJiZSgPnDoSK9SM+ssTsF7nEWTfJU+850TrHLYb2fsfm
iOJW5aOVnJ+cQJMPLD/FjzBlUqGtfovvAmwdkdlwQRp3WLFzpBSMvGIr65xvt9LziGoaUGHiN6SC
b38DpT+MYLu/V/Imdrp7wI8ZFVbrHcC4eGdQy0UAUiJY4UYlHU/49n+4qbddnGGC/4te65Wh4vnD
KFhWcA8oVXfbnYWg6t8SEppIKM6BwvJyj9IIu8BVAIVJv2btQnnMqoTQjMyO9zXIy6nuRSkun/dF
QQQyXOfHv5e76Tprxhvq5WB0NkkAevb4p3GmLP1oJPHvWkfjM5H2fH3VfuD2AsLipp10cviIWxkO
mUxAuuqZkAz25j2bpvJyVLn6TQVAV0gOrOi9J4mQ3AmkHO+pdGD99xY4J8aNzHj1vhX3bbpMcSqI
StOAdLisrc80++ClxbAvi+ozesdjfTrKOCWmHxyes7O/8UprkcqU1U3Lfh8Yk81zNTaF1Lw3RijL
xsME8t8WPAxNNQFw/otYzgyoSPrX16AQcaKeHHx5OotpUDQrFiZK4XQschy1pWgts/sEx1pJ1Noh
8Jbf3fWGYx+gpSEzQjAfe09TRCvmPywWnjIMWnaXGgaQAnAfBmVoM2KtlV3B38YpbkBgOc5GFkz1
LiRh0RM0IOPrkn5OnDBZQWgabSk+2+1kJIO88tOUorwn+hIiVYJG0PluxsawkX/XZ9bNjICS5oSA
YX1R99YwLZ5Mm3reRn4K7nw7qLhS0rKjLG5LYnXCeVx+NpCwTHHsKpcY7U649jsW388VmaXIeRnK
oaIh086T73NUXva7I1IKtppavCu6es3d/6VH353XJaODvj5Pv9ivI9YpcwkUn+785wndZCaHIX1Q
WpKdCmvHpmZ8D95WEzHLsGtDSrI7OROGmaX/53Ifbfzynd72s4xC0F7PgS+VCVkINsMEidevJJVM
J7rfbaHTdLgp5gy6CEKMTKSo20qZzZlVYQyASVSCa2Z9F1btxMML/J7/pQO5kt7a4ki87seOib0L
5K46GO36etO71bP4Ucomn5rx9tSmQQFyHee2y7VbWEMsaL3w7YP2ptW9buirND5NCEuEL4uj3QXw
Iv5QpT1hQufQdtWkLdEUQS7bguI+yWeh5Rop609Clon4vLLdRzBCJmiD94FI0hM1T3TTPuD/fNGZ
w/jhP2BPfvG1So7GLHGjlaYN8nwlImE59Q3h+0D4ZNiZS/t355vdq7Ir2IJcPE/c3EJNY0Gjos/2
9BB5zUe/woFWV2/Od+9HomTPPcrZw+g5y3KtXwvq9mWNGCK+YQi/yLEp35nFuNLEOpCcpTiKrUlv
uiQ0M+G7oSvsh7Bkp5DKP4fYRLt1dtevqAqjCvfRLeGjycfj2u1KpioIWpulJ/a82LxN4TGLaQg5
UwIjew/2JV0umWkrlmuePwS+FjBy/eldKsySmf7XrbCDi3m1ByShh1mN3GKM4b+W6OwRkOD264Jl
S4kZmioZEIluqOm+cjejPBiCD0lXsdITAhudjLLJysFjhVH2gHl3wyfR/GRVw0Lj9ymr9GPbcyfo
/W6GUgoUmDgyYeEt5kIA4+o30X/lOWa0xQqAY10CMuSEXZxokYBiv1TVgZllBbn+EoDFP29pGN+M
63eaOCyyKQFdnVUWiX/fosdAH5bS6Ju9CNJrRh9xmuZf9w8YXhN76+rXRTc/dqizgDy5sicEFIwK
vvspXq5uiYXvaRNIdZRD15DXo5pXN5ypzEE2NjMRegUXYuYVGbRmrkSDAmH7ZCiK8pt22xONyRfz
yR8KVTPCIpoDLB945kUbL4jWSuMPeQYqu2/zlwyjawDQUbOwniQ5lJxiljqXbNY+32S2XJTcKNhA
JVHdq0/xkJwmXHAY0bF7tCruw+ZjPQ4DY8+tbGGogMqNS9Z+OPsDLyFRcioARq/A8AS04AVlTOor
WCdcEb0VwTl1HEOEzQVAni76f/saXXIiyCMlfBAmzVtFkqm6JBIXXK4rTIcI/8kwQURug3inTYWC
Yb49vx8E101EJ24tW7LtTRXI5gppuz4YRsxhtjLcGZFcm5tzyMKB+VIEUWIRdxqkYpCmhP+K0jgX
/OMeMbQdgK3qu5TfHWBJBHjhjyJN5tnpjHP5s248WP/EufJD9Srj7u27dAnvwFRcZd65pg+kv2gW
z04ZyMi+/QkFDbJFcGI9+XXqZ9DdsRifO0BnyEkYRHI/VlsSsMkRaQJaIaP1yN7xVO0X3lRYkncd
fyTRve+HkeR43t+NmkvneUFLSNTOCX0ozlqj/I6T6OsCsIdhfFClYRQDRKyjSl3I3ac8rhlVAaRu
JRJyjP5A2G48PxuBl/TPY1uT2euLQ4UpkgQnewL6j3PJ/NoT9uI6oIeNP4a8Z/uvdEhQnsd3Ndm4
tIY8oNSswhV0g3EWzIicHzRZRdy74qdFO5i9bv/55WqqMbg9nCaB5IfDYSUG8slBOYVA2CJ+g6DU
ull4dE6Mikod3ZZnE4lKbJyYNc1Rnet1AFRomhvKRQjL09zlBYKZuPyJHDaDvJblazYvhLvwZxHe
ni5zF5/8OQCGegaTSl94UCjCkU/UIjDz6yc5nOb7yIW2sUH07QqrtKrJDDSi4Vj/CsA14wMG4XxA
VY+aZdh4Nsuigv7hhaOaMVLBU5z4WZzB9egzZiQ/Je4n8rl+ksaPEBvFloseL2K3aNTZvEKUjwOc
looYUmyueWx8Tz9CKfsTQP2oA+WNVBdWzXYpWgDy3d2MFBxJnovbkXvf14IHCde11G0LFbnCgcB5
6zSTEYnjFiG/GaTKKNGiY7gg82A32ER/wDJEGiJkjZHR095pHznTZTbeT4XF+5eO5UFjUgTFf3lG
10m5+9Hclwn/xi8AJPIVCB3pU5YoB6pI0rxvhWeM/iqTs0ccTow0u2RmCtJcpgeHvxY+S66BfKni
83npA8fNhicXYGt2Nfk9V8CtSnWZJD6WqjhBRkx/pDeDEkhkX+U4w6mdK21cyRw8gFbX347pHOaT
IXZRTIHghCjSbxgIk/MW4Qe6Q/6b916GrUJjVodiQJeEkd5mZdnPqPvBOwu+Smdsr+XkG09TE8wG
aYY1SyzAosOTnGYzVtlTBPF6ONagDuPF7DKbtZyyyRWorzC/r7rySArsjLyOvfJGEE6IMh0+Ti+4
cKYJheH73/o8hD3N92vFjgjTMx5Prz8irv5oclNeVf5OueqmHtRU+UzkMyyLr9+7GjSvr4BhEhp+
lfjpaELhu4lcuzgv7yoKN46rtlEC16EY/OvXIeKQIhOenGVvCY3E5zmPy9APknR08xilVaGkzXiw
mfyI5egY2W4MWkQrwlpBUNQw6f5m3OD7bOtVy7ZyTtPg3EDAlzn0zIiIiliKBoZDX8Ry//TITCrq
PgxQnMFezxhRgcdY+Do6QMHrVkZED9s6yU+hj9HBMbiX7tyjhmd0D+wnyJs1HUCAt1OU7VWVotQA
YwdJc9xlzglj4QPxY++qHam8pS5lidTyCi93Gs27EH3IMFS7i2izl3XNqAKcnAozGLZRQG8Ey8MF
niHdT6k3qbTvfl/pZm0GzImyI6jxHj5dy+pLkPKL3+DWcESjtaz0mJGRL/cwChuvbv8QEntbN4x5
78v07ngoDY7lq+aSfjJQkaOF2xg7DQAp8aNubcsbLLi4tdWUz2XYcz2TxAYRg579G8Boc7NDDoY9
PnY9x1J7Fp+khklApFzOj6PBNcLHa7wYGyUqRQkyy+uF7fhkfcL1/sBrcD0m6DhUWeYyegUliC7Q
qSdb4RzyjKV67UYqOVf1URlaPs8Gclqjc2AOKvfQKMaRVjl4rJdYjj+hUpj4RIE9X3077zirGni4
bhbIsXJt/T3s304b66gMqeJmAlViLfufoG0Au0vwJmA9tnFETeW75f/TLp2TgSVO5DV0IC+9Chfz
LGjmQwvYv3m8BazEmgkROPK1Loyp/YORvphOZ8OrYrBKc56uiMocnHXgB9RyAykTvTwIUMt+pc1x
Tvufk9q96o0f2zvwKM7dYYhpjLeTSef5XHLxkZDqB0trzw6Bl18f65XzZYHMUDwghxueKNexvUIn
8f1xN/1cXHhGr0bM11SKso7jaiT5Se73ISDBFT80EijsEuAGQVHFY2/5lnQiTTULQSl0ZY15F4Qr
y1zUi4g7vvqqagxiGUVKYYXO6b6FYYaYlcp2Xfu3ddh54lmGXkwgPKDKx/b5QfbXN0ay6Pq0cAav
OOX1Rddr/l8Lh98ylT6D41lI5R2KoYDNd5L82H4HxZbZpYBbJicI5rvaozIFmDdFfXGfap5z3Oth
zVwUm9DzAftjVw2bvHo1VCWJROyWCgVWteW+3pdSDqVNzk7wJmpCLBVzBzPA6JzZbWPJHJzccgqY
mWXIvpCAc+HqGkn/jeyvgv3/tu/gWqtfO3Dh9dL6mdkEtc0kcNnCWqVj1bbLLDfmGuKFWnkShh90
Iwp+iIjQX0Z6qT14OJGo4yiFtZN6b56CQekdzW9h6yTxQxCA+oostJGugb2hc6atErP5g7AG1SPt
rEfmrgLpYK4MvojCtOETZ9/JDeUx9MkUEvI88gZFqmruhtSsU52m9RFEPK/IboknnwGWd6Kg+UZ5
OYzbfHQ1TVctBtLY2DNw6071lvYVoWApPRH+DhF+lqnitIJ5krxZ2pI+YP1wDWJzXPSYhEUcAcdU
byE+/uC8njrIFf0fgZT6SuPTyR4CvR0+KtoKQxYuGRJU2hu3i+ZnvfqQmZCk64cuWPuFtPWpgHST
JmRr8Sy1BevJhJXoicZH8z+46neTGiVT12cSyvpzJhYNdteeMZbhLtYY//QRKAVQEHmifyJYut2/
pLTehxz+wnp81Rta7xpC66C8ooggdQj7j5P4EWZZyiStJcRKDNJoygi1aCYG3Qaj81GeCbK+V4Di
YYlRj2JtFJKPk28D644taj2bz6+bCumapwuoY3z3v05J/OyVRlNT0gR0VejORnYCjXBzpj9Z9v4R
zOJDhqJn5E6eZS2JT1fJjDbKiwkACG3wOTZIJN2rqNnf3pH//FvbSveJIUlpnhuKSfsORnjq8Kve
cWcRdHUrxDQ6hMOJbc9EqAAEHQv2EryD+CPae2Pjb/cQJ2XfUoTikDDmtzDGjwr8sTkaTlNoZz0B
vrsIE9u5i2Vor3Ri2XhBeoilylHQ4LAKqV56DD3WsoIa+HNAUQ2NK6EELn3WVU2MYUYPCUtz2Z9q
GURNw9Vb932zblSFdF5F9Wf8Ulobi8jP4y4v8pg5brqrJJOAB7aCIx18PSDIFABIELOE59Ii3/dk
cZYd+xbdwcZV5uL7UWzJmmeyf+vWWAk8mi2NT39SjcCLXnD4rFJV1KRXXi0EbBpAi9YsV1V273+m
+cKZuxVYvpQz+2ULUj0vfiVwpuimFH6LG7J3nVg8ItUMk5QSLffB75Ca3TLdOiiyqPm+496r7jnP
+2Xcu2PFThSItUky8f7jyllbIITZdS+AVsb3VNpuT33DM8NTXDC8ienB8C+5bLNOteC1Ob2L36TH
TDhoOR8ugqHzpMAVDgC30YxIkbBKlhlv84NoCAWIBUoUap5rDg+vtjXVEgZQwJX6fRfpxkc57jWu
7HZQjEn1OyU8GOT8W34COPgQotQJ0SiXG1nBsqDFQQpxTv+mzwCWXrua/yjjTR07G2NyqM2p/LuY
kSt3x5eKomTPvIIJRjpz95TbtCd5zTeq66W30jAWV9oQNsWDiVU8gUi1feCLoGFqK9KUU3hjAdqX
NS/rtgk0KZoWrvu2UzkLdu3ynkh4stqiTTXFMye3m4NpgayFS87/YteumWngVvsBuqlZ54Hb3f2P
JNM8bN5SZrRBLlNXJVLk7/r7L5AHhRpaxcLbIvn0lXexCHnh6eHrQbCvq0DlFSpgZoi0ZtLFiSbO
4Sa7rwjEvsKLGOjxV2Gw5bkIiCMMMt+DU97q+D0zHBQSVghC6i7Meqq5CTc3nMvP4+4sK4yNyc3X
gwBwyqsC68twkh6tD1RZYu3k/635NAgAow7qP+OH7gWiVvg50wAqMMSzYQZcmBY92hGKTunq43Uk
mBJB5D/1PM8X5zl1EFojI2GQngk+HMcQSwKn9drWP91uGMmSLBLx80f1dNqH9ks2ZR/RCTrN6ZAQ
odfU+Wzns6c1a4qMcNSDkzucRjCqTSkff5/9fyxiTQLv9p0Pc2eZzfnOCJW8ylnZtwYa4geoKqeO
w9+liPR3WLIAGIH0SJjAlqDAy2MQWFwC6cBBYZX8HvqMoUtvF1k/eBqn+8gN/ajtfwHDxF52h2Gb
cUk5vSuNxn+CvJrDn0GEKURlgR0fYXSXb4jAF/JXdH6k4TwLrV0kRq9SdW8AHgEdDTuAmZZGcjBI
41PUzy0mqfmtQB3Vn9OWOm5Z+0xgrWyI0aG09rL4mfvhgfmTTUkY+6W7s58xKMbbC7yf3XGHsX+P
p32SysB9HlXWYXkkG3/kDX1UogwcKuCsXz8cVT3VJpmt7Oa97R4KbnSXPYn1NoRBy7Xe+W5TVJwe
XCYdpSwfCUnooZYkreR4EYqrc/DArqZiUB47x4VFbuejCV538Phx5AejMaFn90j5IYMynZX8q9k0
Ti+1qQs0Ivhb45dX2il8F9NezU962iFAOfUn0D2h1CiG9oPEkq6LtmeI+oOUEScTTro0Eqq4whCq
XlTmYHyktI3wSVtxP+FMqvrefvOuVRLJyaa49xj/d+/QNxZ6T01YuYb8xXHnhrPrp6kTTZ7/F2MK
jtYzRgab0hqmhkoJQjVHQQVAbClbzkb/1FC9sDZlJw3QPQozbHKHbpFqOdk9ue1Qhi7HfMPNmIcu
Y2u8gVsPyIfYh7gK+AYf5Vs9k/Rz+azX8Wno34DmswbwSYExrTqeW+GjzELSECUiKVNlyCUpknmX
gUXh+gVfisAmI+BB/CIPLi8WxMCR6iVyJN+wnFT5ybFusoohN7g1tQJehPUMc0ObSaCsHRFIuKIm
GOXhe3J5NEwAo1nvKy3nIRieOrLxl3cFqBLwG85PTnPPuukTWeQumgaTW7hnJHWLlbYOqR2j6acE
sb9eT6XxomDKZA35ahDNBDYbw4EHtBcFWfD76bS4WPGdircJQVGN8mMti7c+c7d7uD1f/LBBcxaZ
ckJYVg9H1/0rOO08G04P1f1YEGbT3pd9UTvOpM3C2ZwXtvlGf7+qDUNk3cTVEOmRu2NipqcnQNaB
Jb5y59yJuMVPlTsJnNLcEtNK+RulbPYQ0OafvnEMJzokKJfRgdSYG/K7bnDHlQEEmZwe/+/gahRd
b75qpBoMBs44Pvf0WDov/ts9fgZ44h/6LUzjzoU2u+rHwFAJ89SLLq2zbIbh/9Zj6h2czwkgaCHc
3EM6EgLJxuDKYTnrr0zo/1DOl5PD700tVzBnxSHUw6SALIDLWesube6k1aT/3wcyBTpYAgvAENpK
lmB+BplKT+DDbIE2c1lffhYbAR73OKcHZXNqkzE+fa4RiPy+cv9/KsXAax+lakh3l/5g6t778GJm
fv08KTXlEOuYYfXd84cKmaeFH+w14CNBlw6QDl6YqK7Yy3U4F+yCPm8NES1gN5xacUwQbxz2dtjj
wsuLMH2l0QMoIAhH1aG02wLWvz1BmV45r33Th19dC9s9jgYZVSAkdYbeGXgapBWrv8nWBWVxnKBD
PvssPVoRpZcjT57M/ZWZFnn+P7HG403MqJQfoE4HQo1v11u4qwU2qMXdDTYHB9gZ1SEtTtzQXGOf
CZ9uQmUzGr0hxxxFAGxb3xE+0Wy8BO1qr6Z+pFvMYbbQQzu8PE9NkPcjZ2SIBV3H2nlaU4ckyFgp
GZUwTg77Q7/7MAg63VZTIR4nKfu2wBsT1p9u/W4UJTCUiimFyC6vkswzJuPPZOMaVOws6Azhcu/P
GZUUO3N3olphmzn2BgruES2PNFQFT38tyBT8u1ko2Lh09Vt4/qjbl+l3LVgy+DTd/6AR2e+36XE1
oOMzfqbTvymP9vSQgxElevJHpML42GehfCMx3dFLcwin5ErVBzAS/wnKD46Mt0CEiTnfv8kqgn+r
f2/DEEJgBKuCIRQV9/yaPW2i8dOIyy94ZSuQoGy3cllZcDzmksR3ifBGIvpx0+JrQ3e7bMXwRQRd
jlWWkiKvAVD7hMzprxC3QKbUVF1wxOXWNLv7wUBY2zYbd45Ry4B006/3m8flnxffdg3RplXw21Ko
rmsj9qnEqUvOnY23VOtsoco/sgN6X7gm6Btv8dR2KrIaTOqPteDtblj+pnXKuKCI0oO1o5Oo7gcA
tzqq4jtcTajNgTG6JTDZAn8SzwJMKwju6n7XjaHk16d4qiNedd10opzDwVnamjUvtkq2UR0eeb3Z
yyAGwOEio8wD2/sPZwAcHAzknTAv8Whhmn3UfAerACKsVVWOcaWzmWKAn7OUBQHjBFZVczU2y7yp
IpnhvZgDWz8YqQ8ZditJjpFrLFSnfFrKgj66HtoZjp6xzgtJ0J1kGbzkGptFT0bNj8QgkhjkvmZ0
tZv00MAN9nPfUHLzSMAfGlNH3XcbhMeJ0bHMZxjM+BllQSH8drI79I9KpPIq46Ouh+5YQvW1w9wn
8k+Yuz0VKY9UlvJygH30IV9v4bWhHW7LlFPjCZhRjO9aU+8wa+1OMAlxOYZfZt9MaC1/75Ay84rD
H+3Da8KJ6RNTmI+hoXtUlPamBPqmZgAYdST/owv2J4x3jIVB9YUMj+Kh4GjGhG7AXVaIVIKvInaN
XO5gmGX8wQpbTgd4b2x85RxRkV6SMPMUqpBP0xfoEa/icw5fARhE32ts44yMXMyoLH79mmJgh+nW
ehTFjtdDvpm5mlXpBwKn/tzRGtVeQfCqnRS6lGNtLztisyOhozzrFGmA86o90wgZXH02AzfrOJL6
H+6Kb5u7VFzzbiVlt/aYpvAWPsSrjhbkjl1V09awZawtNutXhGFdlbizZn0WtRdDldpXXlGIOT46
N7X+I/Wh4UwBlKCBpG1mn/ymGn9WkWkGboZtbPA1Zs0zCPU35Josdr5tiQ9kAhowAqDb01PsDtKU
dNkB8f+0SdYwjWINMUrFm+/Iisg74QaeLMiNak9u8wOQJ1aabcqAisvxWDhd2mQLLi7qOAJjcMbZ
OmI0vnuUZlYlL//0lvzdT5RX7puNn+2fhKgbdewFs9Phl0g9pGCdGOpAecwwBZ/Mn1aZiVNv2MDr
ERGHkWiDuLeWU3ftqREYX4Ir9JzR6HYh6+n/bI3Mdcsk2NwdwTt4PytXBcYeuHSXCdttIUJI5JXZ
Cbwivhv8z4OisZn+KooScNNekU0PX57nvV4koy53zdyvI5BtHSVkYVAsR/CK+PL1Mv1NEYGa7LWq
uium6fNjnQTE9kGqDoJggX+XEpCkftD81WhMr27/rWyHeT7Sdt3hhVks3obFyISvH/qhN6Lgvp7j
EzrlBQbFopwz3tGUeUaIAzk5bYjLRRHiQa0+yolGPif5zxqmpchl8L5NKz3GwVzpnTVhjaX/5ooT
zcXXCFGGcdlPBZGzgsxbDOfHTk/Hrtw/2N/xWQJz7eOt7YElvGWp3RnUFdk2K+K6nyWJul+7yIOZ
Qar9X+7xymgT+etj9H07gi1zH1JTietjzigiSWWjjWrFQmXYVaG3eYfIz26VvFLhenZpDvTmsmJk
lnkopCR84CFER7q2R7LeCQEXa39dBN5BXqfK7Mqil4PKv11ZDR1Or4GTpPpHlLftGcZmEDTKxKpg
D7ogfarHNcEKIHnPgLahMCN0vtYKFgACkd7NGCJNjZ71tIZUPezW3xtIfSqYspJKby0HPGCyyjzO
v3Q++tU+PipXEmYP1qp7DOfilhvFaLSEt1YB2nZ81yHciZEaySOuAdDmy9nkrwPyi1b6s5JuoMMY
BjcL8VXagQLp0LHDTXbhhrnZOdRir0f7rgv5nXCmA9kCo/o8VQ+fQ5InScTEiAfqf4Yru9M6EMkB
KcO6lPcYDeLVjk+PvL50eyTyx2gC9hGLeRLm5Ii3eprtUs7UXaRtthGZsQArW7TFO9KTqyyHiBEK
QrJeTOWT0mZj2U+cWgtSI1zVvUo+vzKQ5EzCoBK9tFiA+zME02Kv4p9Y02JE9bD54mibfiKThJYl
hhOQJGjHsCHAg2j5r3HnvweVeMV0PWNDHk7qNMPXt5ISu3+nNfoC5O5EmaZVBSQKJ3wcuWddxKpk
6Ty8HNBfncq/NqdF3peYhsJAr5NGlrnpIS3H1pZNe0OD/3et1fvbjSOnWdtriIreX11zRbk+MEKF
5ITs1JUiwi+VS4N5dB4GGu8SNcHkX4XdmJ6OJR9VC9SMdkGdIURq2obd/EPIw93AvK780rXqeM07
aB6DrH++OkZQv63lFpv9f7zm789WAwvSgKLxBcMHLOVSwFmpEv76JBdoT/njoxDn4Ql08zFPQqVQ
SYhy4YYWDjLqMRvG9a/frPAdCxkwGfDeIW+VUrjjU0tyLtJaVVDp1KRgIa50GuPL2vwz7XROuR7w
Y7ZAr/KAL7i1gBG3DVyc1HJ1F4lUym3bAxm2ONnKcqB6WLVP9yxqneepr5XocoIxB23eFxLN9Zmq
KWWdQihRQ+g8tcXqDMAUzFzY1y8L2uFaddAzPxea6sUrmEFwdNp/fMbQmHoi8RfUGbky2cp4DGbf
2tlwAy0RYeYR0NDbHXjxUe6f8bhx24uPSwUpPZavelBR6AQ0wyrYkzbiMg1gpBZDXUowI3phW/fT
JMBkQL/fB4dfDIBR2wWh8CXcbHrR3XDO84VrGYIYq0M/tbJjcehKlTteWb2kqpHjKlW2IEUt1ALi
iRIVE0LcvIG2gXRF3EzJTBGts58qScESDyKlBSr7C65pzckjie7zWocqcerh3HjOmlcoIkpY/6oD
R789BCAN5jcIbwS0B0w4gSlaOASyW4B6B6vItXP9D9rT4KvraQ7yj9y9U9lTyb0cewGYkrGQ05jx
oF6hrAMM5TlYXYubLQfCrRZBKJ12LVrCGuzpo6HOqdqo8K3t8UZAeEfFcqeYDPNs98uY2Ti6e8kd
LztDaidvI1J4oNEqEKIReQPcDwTbNRj2czWXYl9asuc6ZmkfH+hr2IfElc+eDn0zuYHQcpAyU1ex
vCKtnuzNMPk5555aCLZlwBmubz32y0OgD7+zVNsGZ0X4bf9CEUj5vXEcV440VoW7sp7aCNJljWm9
01Jd39cGnvThJMOCpdXK+TycXPJTk7jLHHVc3F6LWpP0GpiPEi6R8nxV0TgRCDBe4RwuXvpR0P1e
3kZW9f15ORbrVPWbQdfdHfs1AMazKwC07Jz5MEAPGQdwa7VXxsdQX0G0irROdi3Lh+23AIcyWbwX
WfUTDhTj/fm8d6TImGz5yDvNlZzsr4pbsL0WUXZjsMK9D8z4/UM+pF+6GO6LoXPTf9dMVDySdLkL
OtvzLmVpTftVoSUnlsRL8xsO+NyqBCD1pa0A/PGnn1kHKFpRkTZufNB2YOnpEjsQCoyEPvVzU83S
bjKH4RRvbBoD+3icVPJfYoqWhJ10lN9Q9HuxU0sqlPuKMIdmZ/4LcHkSqzvtnA9iM3d8eeJ1pwWb
ITZS0V+721TGoF/m7w76QwxCly51rvbFCPAoSkk5H3DjzYO8o4D230kQ4/5tnlTCJGhQsuaM3g5C
gbm8lw9DcCC3n9i7lFL2jo7ZHJZwa1nEkunKGHSy1buuYnoJsoaimWoavOnpFSww1caxMZ4MrRaW
MAdr7DEFS5pN3J6TDeiZU9qcVzphAT7Y3pQ8ygPCZ3mv0AvpR4y+3kgt8cyZ+nMWEBCgBuW/SrRn
oisup+9X2aXM/g4bn0V3ycxSpkuNgTHGkSi1vb6f317UPq6hnrsnikXJSboWYUrfhgtt6YA/Fmm5
N6GAOhfnPwIdL6PArOSbg5BMHE+YdSAu3mr5fGpEGEg2gfkSXmBTdOTgssXwmNcsoLeVOZUDdS5N
9eiZvh2koXUg3CkCz35h9yh/QVkKAUNz+MDZ8WoBQNPzc27GlAvDQ5guQYyuhyFB/CbhSHKo1zSK
EbvZ+FWlFEgLcil706pwhmUathBXMDInsn27Oikj0jmdr/Z8L1sIjihUv93ppN6w7Oar1hqbnhwh
Zg8irZnC/zbvojxXw5rSNuF4OhvUxDS11RUTRfwbVZJUO3NgqE+7msI7PdFgBR/xQcJ57ME2NLGS
UEjr9mHaQJztSj7KYbjVgSrruBMhthXhrH0Wa33MW0kFLcdML+nnJLM3dIXjd5UBNOIAyxWHxvug
76MFwuO1x0aw5HKrYDuQKdIGeaq6h631caXwp216y7tntTdH10hgkKC3lB97HUqHPRvNkIJPCSMD
KPiXFMAuh5IdvmebDpeU9UFD9gPi5lCIp810MLD8VcsT/qHUf5MMgkykX6xt8KONErzQ8DxwDV72
nhLklVpBUc6vNVpGlY/vjjliXLw8NzXuFQOrNKFlud+DJcdhQE/iIjNVuCj33YKUN/9zUR3a+JAQ
smrRwiK6L96fwA/bqEUZLycy9+tj9N9tTfSDXNjsDJfzRB4MJjkOktJh0+gR9H63CrmBED0hVewA
zPFdZYnl4bY9pDBhUuyf1nP014KMn2rEB+qEk+erIhxnwmRj6vSUfikfZx/9xEimINhXNm/k3IMp
t68bgAVWdAJUTtHgjxQCX4qKXqq+8v6HUWxzJ0Y02mFte18AWhSFXe/r8z6jhlEUH0u4geJ2UkBy
OzTHVK1US1s/WKzoTtuywODNW/KTqkPztM/6yc4qDv/46bnd2l6Tbcj7/Y0XMvsle16G+/NruOVM
SsppuINEB/7ifITGsl/1C4yN8BNOxpPg9KTFkR1I8VF8xvb9lGRCYR4b8m79Wcxgyu66EoBPC2iC
3ineTDz7Mu+fPzVPsJg6A0jFOEZyXseFpGA+3RO4huvUxmaUzaCxlKnscKAuSAMp+BkD0PplPz8x
+Bu4jdCA2cod7Stf3q+A24jNty0q981073bod6B+JQhje79eDaRodzmGHCMV226ijv0c5LmpaqAE
uh3YHdf+/xAcuSphXe9MdlmAOfYi5WBVFCxk1AWx2fqmSKr8tGrH+TazY3wgZhm4YJ93xNR3TLo5
QCwYWj7rHJJY+96nMBA++aCmH7r10KDP2Cu38+Kg/VhKCz4xVkOAq6SrZIZMLkFzTr/wrdVP5eMF
6JbkPkiwfoT2BRQpInkBVs5UAQF3hAMyxrzCDK/q6/8sNU8+O0J1of2jSOkyqsMyOzkMCP4CY83p
p2EEsAZnLBrIwRWk6JSELpJ6abXHNAB7QNcjuSegVYLQA0Ehxd7e0TsH7ACSQ5D5Azl3OtAVbR/W
gL5dh9ye7mKT6osRYXmGwZ6j2QU24KqvqtQUh1VP6jiBmNo1XWjqTdZYYgJFoqCv8BLaSnFs3cum
oWAepi4X1aWcZtjzVHHdx9xlJ7aNitUqsZNWa2FopwJoMkkAKwE7Ay676ozQW/CbElOcOxdgR9DV
gIJmo8hg7VSFl8Fh7/vXw0Mrthy5J5VKcv2OxLScB8sATl+F1Kee/rSpk2RXUzn9hxvmaQEhR1qa
llLJN1zOOyFnqZIJOKUJtVFN+tj7hf//T5or0sgeLR0Hq0mPNoElJFk8wPwAcJ3vL9IwhzLQAq3a
nnzORlblSA3EQttIgvXz8gFraS7Hd+RKECKsGqmcbbrOH6jVm63V3qNbeuqCttbr3ZctNdtAQerc
08BKT4p3lAJGzekEjMtSm+1DFIWYM3PsaEARPGQtJEOFk7jEds3rX0xfcxbeVezxzkx5uUhYvA4Z
HjuFO4Zw4IrCthTsXyrf/0rkesqOaI2yCfy5JrX9+weceIyY0m7w01AaUP1lceCvkQYFdEIyl/wr
U2DiCJWQlWloWA6l9Itt5L3H2DRlUXnjhiH6zeAecZikYuTfoJjUqG4DhSvoc71PjR2GMM0JSPcI
ZdEmDAa2FuYGZd4XBKPkNfNzoLsYgnUN/vJ4/4P0vf2ucrE0q+lpeIoedPz8BdHVQlDEdQtxPbpM
lDSDrJY6kUhZAoVUDxioiZiKsnDYdvOENzVGGSAaz1oF4eglQulfjJLJGzaamRGV0llJtUaJ3EXP
31GKpcFwYqoeX/Jiw4XgXstCfi0Uz4EUJryWQxNcRLBRdsQItNkKerr4BVnlhU0eh4jHihvqhn3c
ZxWNuVPzttjfXK944BXSCo0xGHtUEK7r9kgoXXQ1y3R5+fubIkFueAbQbMtkopb5Ei8PIBgPfK+F
IATLw5OWz29v7HpDcqEX9BBudgPr2rVBS+/XQ90IWyX34me678GMq512PvLsuPSSx7x5JlWPHyom
J7TauMgGLzkCNawun9fP4rf/cPxr8y+Hm/vFPG4QXYYqcBcsEZZYi4V1Gf9xfLfqFXKlUI45z74F
KCrPSU4DukCYgG3VaOPdL1xHRAEnOsrJ3G3SoqSJYnHLZcgjf3c8vep7ZMYig1HEAnSSiFDyPcVr
5Y3hop8coorgEZqs/P2NusTO3j9jFWXf6RtowHVQpXSZX0hpEvOOrm++jBjtmRVS/j8tZ6lzouks
tsESuJF1BX6BiHRAd5wvuT1un+nMth2AN5snM+cLs8pK2aR+Xk1YcEFK0kAWVxYyi2QWZRJJzbtB
weabrxo5y+vCQKZpbUP/H9pOGMQZEx45l8kd4VdxrHJg26loPijp8WGrsWwyq0v5xikPoS6tR5Tk
+BlHtB4WiqvbfDiInKa5aOpxDTyGLDJreYqUhGYJJKr9NeN8gu6YmGh116K4nS4EgHVKrhNvRXNr
eRkMKwGg++Jvu1Fvo/Z7CBjTIdPSjeqtqP2ajr2oky3xp2hFzotXmlBk5EHN1pZP5NsMAxm5LAHi
GGtEKc9D2jHKk7EvH6MZ5dyjBfAp3+Rq4tKWDvonWjQxwsQOhXyitSeiCMbE81zyf2Io504u9/4A
F7kP5Tsibyd2G7u5cvnzBL5qMWdfNSQO4vulAiydsujcPXkssJgjfo2Ecogvh+jf2DVkbNbY6OR8
4zjihUju+wEUiFFJ6IsNLkBf5OFp3z2jx9CkstOljL9y4oj7lOjubxMwXljql4zzCSYb1Rt9zNPn
LlywM6ISwYG0VuaH4nWZA0h+yAfiovIgqeyoWsorcNCwsw43EMBk7ByoKHOp/rSzmWha3aL1+x2T
hqILNqq4Pw6ThuiDquXqIqE1dCD+jsjKJSMbSFC+R89Aza1giZTM24cDekU9+U2nCXXcjvvxIAfH
rHU5TaKXHAtSz32jscoFODA0Bo5vLOgcGTpSZtP0tg5PWznfoHWhRO9nd1ZkEjV1fXYFwKnY+lxQ
3faDX0Z9b+EF1p8mDF4yIkyKfhOirTLGn2gVH1rhlLtveaJnRh/jLGcJy9FHvG6I/6kP1KBk5pFs
YEy7K2puJp2GQwNRjjXEe5ZWKsO6wy/t9QAjhm8pKH0ELXBIjNBxEF/b31xhGU31/qkexcRYLfJA
fLkurzA54q7RdydTnKy6VKZCU+TigiE1U0XDmyi5+55vuUZB6eE25W6KbAXnGpjp7eudhbLGXDu1
9W+ykHMV1K+S5egvZuGWgCjxJvqbp/6IYESngZDmPFlYAvBm72sXU16Z4EMPXP6EoggqiW2mnOqW
s9Vvgr6UYlOJPjThzyIaGRrwZ+4OjsoUF8nTgBNL02f5PcJy2Ag/O0p7THu+UzXWxNtnN1s4jWFU
dA8JYkw3WuS4O63wO9Mhexo1f6lmxu2mWQskJpJvfBPAfLVTTFc+vFosCemXN0oVRpqIfRExwBeK
TS1cjVtqL25WLlw/2Laxpvs4KP64YRgW6GfN98l/R9v/0TWnQrv1WvHOS+kyzjVWKamLekXyb1sy
9o7ZNBYOi2cGuxaPnU0icegdu+bO3ytdmNs3HJ7R2avfvDakMr731VvvkQyHeU851AL5xG0kCA5g
QPaqAin+1jfOKiE9rfsSlZG2BV2J8vIMKDGsoDLo6UHmdF3YhJmXClHq/nOPtWgdCFajt7f8FG9Y
xIy0DYHIgIBrglowHY/T3xrUV2o1w0Zq4upioR8bUZRjXx/IAXe8bRb29NnhPkKj8uysNnIipgEn
2g7rjmGVnPwXVuIVoudb3aqF8G8WhzeQaf3uFolr8x56hghiH6WHzHCELUFt8yHJOTwRzpVpUUFM
7VLoQ1zFGueG4jOevy7rQUT+UhuryOcE7x0z1wD/JDhHXYupaNKuflzDx7cWJyTQ/AQErC8HpQVn
RfMaqQd5+Qo4Bf3G30l1OIaCXBf7UjAn5ulRPVAffgRgF4BFj1JVpzYfoLV/vTUKDjPuyITAjcLv
8Kbqq9kNyw8hvW7LglZDhJrPTObnri/45GsA3u9WxkuIKTXtpZ2c7QU3ga3ELGqy62D4P5lCfPlA
YwkL5+ZR1z3s3qC7k1KoYzw9EWAHX8PKodUbZqQRPDP/YiTl+5GUmUCi5sDT4uMerBKbkZ3936/k
k8QTRPT6C+dnP7CPza+yCMKTWOSGjyouZDJ2aQeVzUuwpEvpNvIK9srGXcQ+H0V1HdaxuTsGVKe2
cQvTKw4HTo8jYj4YNoksBzp0u0o3I4ZLfrw91OJEh+Pap1fJQdPr6OjA93pVweCE7nbjf9ab1yn0
8ptNu8fAqzcLc32oVyxhBy00pJcmzEJRgMIDvwZbXt69n7B6jWAuSQNniDHOopXgHSjltYC+sUFi
l1wVoOSv6LhMOevvoJjJhLjBWbQ27ziQksHTnHPD/ZqzvVDb4cxMzWVTKz48Q9SlvyaLjzzbcjqE
FWfbHCwhAw/7XcEWL6V/0vgfDcKEMlMSiIwIgy7EHyoG8qI1K72vxizwFK/zCpEQUSmcZRHpoU0o
eQCSZtQBRPtAEbz2yih7s2M4d1XdamLUyyD0nptsG3afkIh2ERd6UoPsFpyxEJHZjLF5S0lNQMJi
diIpja2rjJc1io4K296bAT7T75mLVuMarn0j2DCZvTDWE5h8M+h9qiv24upu0H84TH8vT7iSQiLm
XuP+W3/wnazBlTlW+3CeAYdrI3haxAAHRmpaxefgmiw2OT/L1hvT9qpYV+RI8CsbnHaBT4hoCEZ7
qqilk2TlFDSGh4GKp+wufimdGl/uqWzeUswA5f/REnEWEE3IZ1/E76opudpLjjpSEeQEpGcgDN3m
46l0QriUU41sohJfckY+GQjI6UE5YUMEeJapxbLEW5fhetbo6Mz0+38erFFhL03ujIcdztKN2zfH
i5Lsq41rvQEcE5GOQbTSuazR4J9r0L08EWGdqmFluoBYpOP8w/jqSgoeD598IIrxwLSl4+LjLivS
eOGxC1kRF/M5/YGXbAQuJHl5gwg+LgZ9iD9EbQ/EEHpjBnKxilIQl4m2IUKXR25wULaHtVcZZ3da
eCD1iDtU8ewzVYShT8DFAuLm/QMYdb8a94wM1BA1KwAzCG4uldAT8KaFMbX0keKIxadgO57wZkAt
7EemmNvkgM6X6LzBHAmquSRPRQ+bkcZV3KqmArgwBg76CbpigoraBrjs6nF5tteA2jy5YAzUZ7BY
T70M3XZHiLmkfVJVgutYK3UuYwV8JrX+ohSx5kLQc0GgBT+zkKRM1s1zAAfGZuxyjQ3WKLMMK0Fm
jw+feCYk8uUpjBMuy4HxzMmNwqnekrE0X79Gd3OMOxDojDhYQChXmZU6UqT7AW+c+U/wyyaggaLk
xZXEq4rjSkWSALh1GjlGNp47sc0RvFQBGBPq0ZtinxtNJqjd+n9PiaArXdDyOkCScGbCD+cCtRIs
qfVm2Nv+eAU46XqQGiVbNG9TNk2YoTHku9ush0rHxM/pbm3K5WdSoC0dUH9slZtxoZnTPY9bUCiH
/WnDOIzg+VI+lSq67tWXsiPHSCLkkjphhL26vNaRv31wewghrnGyQkwTy2KxzZU2KeWUP1RwKJ6f
CObdYBQLTS2P27gCF2mTbuF81SDKnFmmZE/L8wB8HfqhxNETaKFYhZSo9uu4U9Kp/UNxW3O5whV3
EENN8KxKWad07Ek2i0FcHsPDnm2DFzjI9EFdjvopDJuYdnh/cCLq2DxroCAAvRmbiwrtv/pbREqh
3YYzA+x47Y5SXmxymrjHwTUt6zy1/lWS+E5WkjXwaqwWWxcxPwUO+m9jhwMKfOUXT8fRaQYUrbS4
rJ6lpYgSbEadJDS4toUdtJVvMc9sJDP2MXEc0EEDWcE5wFTZk7KLPqKPUxeUJSG4BhUy6hrGwIS4
c1VNT+Vn/pU6hgktdsImOKhbcpykeaWDoLOI1SDhJqh63qyEKQIzjuczrG6BZ/ghMugUFlNM0a/l
Qo7eXlN/v9TXZ2W/0nJsN3PaF/nrnojQfBvLaMUuqiv7og+uZV3p1WOJIA6A1kCjj4GvMoAbVDFv
TRdMZ8EnqwUVir/SMCIDD758zyO2ivpNPWj+NcX7Ezq1cGLSAQO7bX1M9nJIWK6VF5k6sCvloQbO
Jx4oLKtk7od8k/2ljos3YAaQNDW3Z/VkK2mvXO3b46HI4kcYDGgNnk5FRN3lGIZ0M2LweJSKhRUu
XdiDU+xFdVookHGKy1YNO6u74lEKc2nuR720gdxmtmcepI2pJ3Yap0/Sbn+OCxInxzKVuT4sg71F
9PEokr6jINJGe3eROnMbXh3O6F7BAV2i0+f6Y+Fzb7NwpJ0K4TfZIn2ZLrVEdM0IPtUW8s1SmY2U
1IlkNv6VncoeJ7shDbRj+xBqWUusBGhPlExTrkG3ZPVFmbl01OYEZ8Y88A3IXkDYZckSeI/dK96Y
bk99lK8jM70s6fSPLOEluWdvupVVcG5+3YhBtq2mQaCZpaFWItYXT2gzn7DEksGeMtbepOGO3SE9
ClFfh9KaqGQqcqMjiT2nHK0Wk6TXhbh1OS76J/l1k2xL8y1CJJFBTFLC/yIeXDHjUsXNXZNpTcG2
68OC/q6FcK7PMrcNKS3rkH5f17+qBhH9PnXkU6YrQUOVLIMAPQDuqnBOfCOVCDULPTr5zSgZ4z1t
EMM6jp4X/MCw/4b0KW7asyHSQuY7+Gc8tFojOo37eqnfoouM0BaIInHXfBuTh7AAOaYH0UIF6eRC
tE7KzKFKcQ/7EbrctGQ+nw03YUSa2ZTJ2I/VhPlUsPryPxPh4vU/qwEXYER7Nmf6dVmkOj7EKL1C
CkCjrCmTV+qW9LAJgoZcpN0K8JFsvi12GM6ArtmQOmLGTMTgfNgwCK2zABXocdGBD2y1dzgt5w00
8FNPYg243+oACcCxEaUL/fWQELI/E65SfpXe7Q8ZcBgE7LDgHNp+7Al/nudvsFwUa7fT+HtDSEPE
wqcKRK65o1GiJJBGVp708F4WJbYeDP7ENRlZCDL4FMTKkmY6NR8iRUmCU7Qp6C0yTxhO68lpuj7Y
BaRpwXjNMrUQTsKGiGJXyxnZANaddf2yroQq6xXvGhN9efeN5PjXTK/FUv3b6xOGn8TrGWJnvhEF
lTdoOHRmCT9dH8Jb5CKor/EJZErAcsQR+yIgElMN0W2t6havd7MdxwOJo46FDt3+b28JKkW5lq+3
bxIdvGWIECSr0ZGlrFEBl7wBN5B/ZivHEZclZElBIEOMqgLl3fwL6oJW0MAMeGP2j/DrGj7k4COR
1IGTXkizgvjx9OrhYCvjgUms/9NXuDZ2ODLOZbtuY9hl9U3AFMyK9GlCzANlRuH3siqZS1PV2MT1
1Sr94imSVsmeTfhY97EymlJfS5ANrE3+mIGpKlZzO2908Lmg6x/eQMX+Sj0PuoRUTsshSFChQyxj
UKui2SKwv9TvrAiJI4F9Wb602wF/D28KarB75hCWB+rHzmbVTa6tk04wXKfDInMNML0s8FbkRMaK
bYWx3wFCJhw6yBO4f50LmBqSLuVL0K3pLfi1IQInwpiHdOqB5qA8JKWrtgpcK2Ae/JIoTPdqr9t2
VK5gLQzQguyQ/XXdVCUUIMup1J6QwUtx1/LEDQ71P7G0PfyP8qExO2zNOYJENgmLk+IriDlxhqB/
ntSRdS7IYzLaw8eMA7zHXIRI1Zvs1tMe4VJSmU7d2EMjdlp8h1OHBxFlFVauFIx4Xrn6hfOt5RrN
H2VxeyuX437252uXsLMI+NWC2Bjmxpanf4KaRl9Zf9KL3O5TsvVBy/2S7PuUmS6h3m8sCqn37vJl
wKTskd25BXpPcqFW8nfZ1xENmpSbQqrp1XVLS1upMMR7HP6BErzxUwL9VIcMl7jsP0isELIbijRX
rZiiMFo8p2bQeSUKZRgEvacPC9LtggTJVWD7EP8uR6QOqMKm4W4vFzVXWfiRRmAul4/6kng+AJaZ
mUrmEy0VCm485sLJZAuTbeD33H4tF2UeXgmhK7TWHvhV14vVtIEQM/S/m8qBnN71B6VpX9ECMWku
4BvWTOLPzVoYz5CSX85ZUPiwukbeYrlxiyzRqCMsjxp6YrkhllnMy1mbZNcXyohs4qE6Im9yVDWq
sfZnU6zFqE/kyPTRqvHz9TCxgqWjhUDAuOdACLYdtb51z9byveFEPl5kqjdUGvC9YLEitOYii8Es
eB0cISlpfqIJwr8tXdsjgBSecQ7g2Tv2ZzmbNE58zUmm3xLBEZggR5ROg8xA3o/Wcs7oZGpNmCro
M2uw8rpsF/4ijs1YWeFtQlY8xnORVvK3VXr4Tk7cNK5Dc6SYSu6DuxMJGvkcF5tzS+0v4xwmGnEw
DySN0OpDShaxizvTlEvGWs3oozSTFe0hjs3OvUwKcvSdEzyNOs6CZTwE5cnUyh0kZKg29+PSk9UN
yR0qtwlfQbNeb+RlZXOc3F5segJRPih1SX+fZn4apBHGtnomkmN7KU6XGQni4+/hOnJrpO5n7yuk
gu9kFtv0WttPCO1k/f2LsJ0g/jx13iXrIn9Nygw9dUci9g4xgoXL5+kxQb6rbuPOlC8CHepCtcfL
IPFYLansKLjhd+vJfIgigf2biN3QUfNl0waAdeAfNTf0dfKwWDguqE6OL6/JynrOFLs59hIvRNjB
SRrqnHiw16exLLkK7Ukz6prO1L9xT+3zxpfReIOLPDzf0AUJ34+5KLJ/Xe0Yf3pbwMWZ6F0uWGdY
3yIqU8lxelvJ0RNzUfRUdCdjS3ViwSTfnrXiY+7BcmmbdZyRmMMeKbO3tqf+yKuIinUz0PNJDKrD
V3kCICfLJv0QCs0XjzwXeCxE137pP2YMzMPv+n33uM+Vrp2WiEphs3LPGvXQgiZOYtaOdbs78IRc
Sr5oisGRy6f6v68/BSJLP+eAkfFu553RJkVC1zCGlEcaOG906c14JSNaF8KBXhgNTjScK+FmSNpH
fYE2lgiwVPvYMUmFfQNFdYyD5/+r1gZZ8xsxiDO5QNbJKVFYYIkFdrHI3AU5Ngh0Ja96Nfsxl/9v
009mg3iKnXxr8+Er73dqbNIzuVj1ZXavc8OZrW7rswkGo56M/jmFZMMqtRVnaxDz/a8xoBntkJSr
g+TOj/tn+QGVXUovEBFwu7BNVQRnXOmbem4ItuyMuZrCfbD8Fw4htUalkOl5IGoGHuZkeMjifvbS
aI0MxJ/uodFZhVIVhWWdUGcsPbGfqjy1rFFc4WG48bs4OEDj7Vsej1s2fcvWGsN+yKL7SaqaB79J
IMRE8Xko8m3keGATnbfprWLvrnlc6ITV7hZDvxS3TwIaJT8nUsJlrgtfsLoCUlASa4y8DXX6VfP2
DB8EsD8SQ67WuPQX1ZVufpWdJ/+hh2+ePNjDxbAyWLIYwWGKExsQvTYfTj0MH6+A58DSG6PIdvTC
/Ja/nMMNNUkVui4BJE6QiFGPqTd6iwjf/72rp75/QSDAEZMLu/lM9Yc+ogMLZlR/lRcpO6d7bKQH
OaP9RJn23Fg/ggQOdRBHknQFuHae3n7aykdbhO7dez83QFLjAJoV0LxvT3s85elKZxCLwI1Voegb
sd/7hQ+MrckkmqhIrcinZUkpCojYEKTIklK4knURpSlEReVTrktkaq/rENAEOjsf/4qpm4Tw3pBE
s7ismbYsOwAQ5fHhapoz/+PMNH7to12SECylVVgoJXahAWidOiXDDbYnX5DGI5pEQlBkQJKnQVax
j5OrA5gTXdSJ6DqUTgnye0EYhqRavNOSeXha2nAWi6Hh+jgH9CK1R5XvO33NpjCANPKdEGDtiWRI
/cpG6iSvbWAeljwofFXDa5kp5NKpVRAKP2afYAWcYXnMnqmxXY3kr7ExRgaqwxVtFrcUq7gb49+h
d7ZMutPqJjA48CUx6b62eW1sSv9EgW31pG5mkd/Q9GWKPRrPmWkmCfZvLHB+Li4QfnXduUbxCCET
WdvFG99IWBmP9kXBAjaDHViXbQdgTgFt8hD5T5LyVzmWKy2KrBY/JBL5GyuLciQV+jwXH/xi6VQu
DM6ERTk4Wt/8E9gRA5RgIl6x1TxTEJf2dUEndlHQ14e/gZjhtJ6v+zLNt2xq71fh9jM+TJ0GKEuY
Qr11NSXulV5mN+eExIjHe3YYOva1PMj0enmNO4nFpV+neJl0q6u8Qb8W5ZvC1UEV1vmdWQMdeCML
ajApx14NOr/YtMCZrt6A0aSJNcMiOIQWrb8+E8GGYgTLmmjmrKVTDdxBoT9al9+HYXk/ys8zDJL1
YqcFZBoaSh3vZIy9mcITs0XC/e5sLsO6r75oMBBo32MeWxTUoVvGCJFaB4TEsBCN2CGE7qRYKPTz
8BEkySS8yT9umM1816Zp/r2DhheO8K9/hJ2eWVn0ROwkrXlOCbJ8vrVspQ8Gq0NdrbJrWPxuj3og
H+1QBUoS9q1B57LIbUuPMiF3BW2dp+X6FztI4RSVlFB4YsYS/yEpX+57WWAXobVmbEjX+DtSdmaQ
F4QB0Av7kRkjxly3EBrF8QzE+kVNFQumQEfUpBiJAC1h0WFDtnhFLOEz1YQVqqjCqVfCpgtY4NGK
SRHZenvn7mKc2pxeZto/Uk6Wzqu+8wmCtfh7seJ4Nif/LyfFaSRj3A21z39nISC09Iqf02nc3KEW
UfrdtdlJO4C6p2uzPILHS/faWPQb7KI1PsY8ULidiYQXM/mUP5GO0E+qR/5V3Iy05hZtTuKgWM+z
xpH533tsyAWslMeDFJARHgkLBIaYB/VWyVbR2NH1DRHWUssy5+nctvovIhl06/rrlmrbm2ZHzOkW
hLibrwYvdCa01JQbyV9bMHyLQeWloKxm6j2b2ZX4g82eKf7rXazZaLWKcfxnqc/fSHtl96v4CExy
jYyRV381D7pcgbAUsLjCaApY2CMgVCL7sVLGOMOSTu7AVIvfa4M3q3Eym8+g4P3hBNCg0B+8RY7o
Y8/8pxBdE1hsmGh3Y44ZNmgo+4NpeaB78aiDkgTTBod0VGu6rWGcqpD9IT4qURT90BFF5YVGgMf/
XUHtfByf8Sn2Md4wezDbIBJrbxf5qsa59Z7kzqds2yd9E3OKOQ9hYUEg8Ig7o9LVqx9Ley6hukO7
2h6PBPwZ2WPcGa1cWk8q6vjv/kLyusvGwctrXoQDy5JymTgnp20dYAYXOdDDCQ7/49sH8k+VZqjF
FqcnN4y61o0pQ7w3778BJcJJBmLA0X33SyxM5CSManvJ4hX9adY+obFGlY7ltC3O2tC9jjKpkNr/
NTZwHqQllEDJuUfLgRZzi/lWpvIpdJW+UBtptTfv+H6Qi/sbHAiwhDzkDyF/L3TO2AOPSGwYNO5k
ajSuIqtulOHfJBvbDkgjqNo3RIZwYr1PV/lIo/gNYFf+E2ml5WBJoSikDvzwCHrTf8agVWRp34oh
5kqxyxce3RBHilithCI1eu+52cWYCUIkIJoFvZ5lRyn09tpDKODX/qp9mgY7067Gw2lQWR6rxFK9
5hRxuBxNmeIgJHmD7X2hCvOqGBoAICo4Mwx6oDPhZXLL3fquRTPCO1ch9eeAvvCWUutcvJzF/DR0
7lWnInBmg4BaeaB2B/Kxe+JPVtTJYzDB9jgymFTeg2qfvMw8kMndt/EqKrAmGSldbgRpPfmZIFX+
kW/EwKIRR/f3PhRPfWt58vsWbMvw+VRirNAOXo3OYP1mk5fw5ejl+DKjZQzX7GMy7j96s+armxOc
pmGshKP9FN/ygfKqHNO6veeZKqAyiVe20Oh6RRX9bPynrVqER0h0YkZFkegJKgzK2w/bzCXekShG
Q7wOaK3Gb2ZwVfJ0DbCK5Lf38apo3PxaEI+3dkbgVXkOZ4h/GF29F7Q3xbLco5oAYMjqK0f9S9VI
KWdS72MJfcLtlQAd7rnVJUr3TLhrcjcYNiDHYNm3/TxXz08J2s+jQ4ZFajW4zyz3vCAaHQbPmSyr
AOGwk6dyWVI1WWqcgTCJ0FBoA8ayVh5ofLdvd4EYeprQ6IgwAuKekajcsiP604patxFZFPTSZMsa
MyMgkJUvRNnTfYRiFmMapFLqUKq+O2x4P0PBDjfpQNySahI5tIeF6Ri/aV1hu2AP2louGIhE2svE
gHMPxhMsxW0R33EPH6zQSSwKGwaAzux6V5aybdf6pc9Et8Eg5RmMThLDBlAGrF6MhKJMcEJHmovy
itK9jPoSQpNGWTaQxR8vtVC0uTLqUl3/2U2vbhm0sJ4gbiXAnUWa0GlYQJzzmdv5oNwe98DdBjH0
ZBaMucPD0AywVJPoBkZi6QLXKTGIb6qWML9cjEb72OG2euCMszoLHt4f9H+L7UYYBEUO74DFYGZC
GyGlKm5cOrJ6bAoKApv0f5OsWTDOSPmRLmOn+/NcZ+xGGwD3RQ30Tr6BNQ8DVpwOp2e0ITZ15xnT
q4Pr6aRQw422p8Qe+mdGtItyRWvky9uPTQxTqrK17Cs+JPOJ8obsfPZbX9xAjLiciYwqAdd0Ev+X
zl/8GlTwuumOfiEf3WlAm2lSlKKucxzxUqaYXlX/8V0Q69UGkFKcfEryRlITHKx2KkS/5s0fNzb2
7MXr4i+3V5zdsmiIeObIFFckK5C16uAh4lm51xSymFwQZjOktD5PfuG2oslUEEDhCMMA8hXVqfOU
6HQp8YqW42sBC5KfyrC8v6DEIySNF4XMuMJbmXkQLC/7v+3Fo7dVjHeL3+/3WsTXM7wEprf66s3D
PGd9QMqiDZ1GbT5/LQiYcxNx3Go1NaMno7LKhQeLkq9qE9x/G71Yeb8JexPcC2PCcFhWqCEvTueF
DCr8G1UQpd54YO29A++mDS6K9C2kYE9u6l+6nxDisl8VewZCQ1K8Z1GXQTKv1lttzsI47apJOoYO
7l1X/vkdqkkbRRIqQMYTrQXbghsmHtQiNveh+ftxaUEOGFr0WBsYOB5UiCp7zU6xDmfCHevC0E0L
rdb/At3tm5ciaSAHeXY/rZwRHN4YtpeX5qlIVn/GsFvouiPnlMKO0cZRt0KlTY6BTjfv9qFBRXa5
v209RLes7EEcXV1rCezdedP319dJ9atZA2iLAWnHbAHgyA8R/NDkh+cKff3+lDWbskGkYf0SnvWh
InLc4r2Sf2+6nDrnhdEW0VCi5Bd0itb0SG9xRPje9ACd/w+n1SDaleaJLIA59xrBLIVHf1Mh8Ikx
kq2c+1Bmhu8CjiMbzFFKf6iPd//lau1AWUYg84uF7p6lKEUkqpTkd9HDvJ8nkvNfOl559G4gUU7I
nZ8os4qksA4lQjBUv+oRBcl1jU+HDh5Zml27493C/hWnfIvd6A5NdaTsNhfBILwdb1XKv+XRWSsY
0hfC3mtY7U91r23hv73OdZj/Vm3K9jExpKxE0DhNzWv8WDvosF35/ggwgMPG5YNxVcZUrd1yNXXF
9fxQ/UeNBJ3KZMdmiwhtkiLMJZ3sF2LogkJCW2fNIcXMJupZrOL8/VDVF4A1VLVQy67srF0V6SFq
R53XL5qy1url/kzPLjxlzeEEh2Q8Nmz0/KffT9Wp0Tt+FPZkU008cftuJ8Sq+nLg3fRmr8iR0wHi
F0DXroKMvIpkGNMebo8eVs9ox/TnFwMM1nHuIvGT7YgVegupTJbbOUy8fJbCvoj6prE8J0uv2ofQ
Iof7TX+nBVvQbzKMhHS3e8mNqNhtCBxJDFq+0k5NIg6pX2awGNtrZMi1uhwqj2lfVo5NwxfqK05W
tJWPSS5mZC1lgxMaFrZCyJN8BADXva0ZJCxYIPGmP+d2uabLuAPrL4QDzlyVg6/Dk4WRPKKT+fQP
g4y/+lhO30A7q+3khvwnloIl7wHsxzi/gcZTRiK3fo+2AxKfEKXFY/ntM2Qsq+UvRb0mYGRW4rRq
aNKp5fwdWH2PdL3QgoUgoQSqHkEjBTo7xhNRpWM1WDQRpLFnOqN5+X4DVyAgnw4Rg+/NkT+wtCcv
QJDCbiPYpcgK2j3rn8bwci6YpGTdaNUlowT6hsKT30NRNKsNqihPhhqGN9T1mNHZmpa7cS8xYJj4
79z8f8tCrW00uLYGONjvzoRmixGp1MppGXxiToL9PHpPObf1+SGq/gMlz4MUHVJEpPouFHQnBmib
o/J2/+wiIZsw3fXBpF6g+9TMVQ3pxaziNo3uJ6ABYJiJ9q8J11ZyCFjPZHTH5lBr6Nt1T5bjgwCn
kADrJLKIopxwWZPuplW6Xh11UYVrM++lK5Jk0i7diHcPsEMp+qAbUhWoDlZ5csFBy90JYVZayQfX
PdtV1ah1PczJD+7Ljm1tMcwvpfHtr17Hw2UkbFovKgFZOKx/p1EiNheoubjo5MkOIHq190Ft+j16
zhtTN1eYcewwVa7kboypZ7HiPVGiiqZUwiiqtBcMkFtD74YKI1ukFupMW7F7vZjZyqtenmBZ6QlY
UZZCvSyXRXpo6zDsIQz20q7Fpan7ddjJz0wVyxUKgEgqJknKJhPt3mgIDo22CtITFc1WFF8ACWfa
MpeiET2btOh0wWHkn36XTmqv+21+Dw9v30Oa1qmiWLnJRdUdTzVknDSBgehHisRAUnVXVU85+5EX
dqCbHK25qH2+4aMHjojnXZqI4R9erDwJlIoZXwwLs6iZ6YDxIPMw4jXmIPMN5x5/2hcPzPpFwF3j
RMDqsD2UyI3fDsnmAR/CAXU+hor+VDKib6G0SB69Wkc0zMuqqDYCB9j9RkBn7hjzFiHiTnJRjEro
m0bAdYLpKmnDCjhxZvm7yO5ZAI2vFhfPCyzOondeGe0Zlp3kb0SpggvMxUKp8anVsrjJvCEm2oLS
+m4IpRvlhc98vDqyERQemTu5AUnZOXbRoi2r5NbPzsGOy59khpHiXI0T0/MpN0pSgNf4nbuUvtr9
9rFHw2AO+omel5An5tzkE9B/LTWIERTTh77ZZsKX8cO198RpvIPBq7DsGtAXygrpcxOybrPJwD06
oh8VBk1y+WBrjopiAll5F4NGy9SI/4r5/sbTJksY9SuoTsOaedhAqIxih5ihn8C+BW8qV/6n80ns
RI7buCJ4oTXu3l7w2Smx4k040jLdajgiUM4ljeXXKUDFSXpwvMo3g0shIN0FfhKcH56Rms/l0qH1
nS6Mktv92FtV4EKT5QPttiMApB+GMitrbnAFO3U6CVlwiMb1qU3/TF4avlfthcQXHsyd3XSTQENq
u/i0sMBISP+WqbsDH0VvHuwnwlOxDeYtK5DblaVeQHCprdHfVKBc5K1BIoEnGVD0Tmm4uZpOayGd
pUeVtbFbH8d9ZI0Rgah/Iuwi9rbN+Kil+i/Rib7Mzbls6KbIqlFsJ1wI7nHKCgltkKRVcfikDrFz
H8cJzntJCcHBeKCRIseP/Fzvq8KxAIGQWpdjjfrZXvfxN0niUL3815PhNhMwEvGA0Y17OGso2ZAh
fErhEGxJWiHrJ9dgbBanJnPxMPBrzLI45TQi3qemmTG3RES5vFJGI548+i6eo6cCZVgQyvgpiDXQ
b8bMI37EfkKE+/wdYO+xlJyXQeJgrc7JIQxQ3FoDVMXWpsWaQkMVA8J08o2c1Lzqu2jaBhiSA71+
0FXUuSbG4bM6gGzIwmf8vP+NtH1QmfxMhcD2/y3U3ka7vhn73pRVVQFXWvAkj9to6YLxK4U5bFLL
EK5OVJHQhM5QmwcECj30XQXxAH75L792Vnb+Ui/FwHL/hhT5XcQLY+fXpwFBO3CxU5jmVFkeHHbW
R3chNIi1/Dr82RpW1ajcZW820QxPBvIXdpxhOo4LUhOQArbXIXVrDkeep88EiT1Afjx7fWG/mJsm
eu/A4nmFXpP44hCyznTgEuMTgyaDKM9gP1Ltf846hW3gScBHebIItUD5OWxV055QlmpYnFBIjItz
XIMIdRKI61GSb1uYBmPJr1WHB/dn4+1ayXnnqbaXmqzCIK5c1JSay2oU+csiyQfgCUcK26qUH9Cu
rVJ88cNV72Mna/wFVPLxJB9WPWUDtqXpZpKBM541zx2ZKGV6imMcpOJDviUXFyfCng4/R394HhLY
nDq5loJbJEjrnQt4z9EdD3LTD42bsKkfv+mM1d0ZTZ4ktRwZH17/ITjH6gQAggqt/EUGAlHwU64y
Ulr1rbI2HC7jYyC/oaMEnOc1FplloZvg7AweiA2PH5CqGpD7AylQXQekB5tGFBnyjMwvnqGJnsRm
GRTLkzjCRY0hHPMTeRYR1t4fhWuFf7aF3wcg1ATGyJDMC8Suw99Do3Qn1pY6mzzx70Za1gtge286
7y2R0hfobAzP+bwnUWYf8PzhqvHVNpoTes7UVGAU7dBjumaeQ73VI4FrA98fLyIgDexVnecqdwEs
ks+G0PzeDNRC+IURShwBtHxuGA7/1T3XDIA529IL8QoE3BAJ+1LgTWSM/LT2++Af3KDaDEg82OlB
wUh2GJdMM3+L3d25GIT01qVzyZM0Ung6C8WEcWnBvwzbFOodx1LU/kdkqD7sOtaPlmd+yc0PdxZ5
C2uw8HP2cjYbaUHIkFnloBjh4QSYAM7petvomE+TkBtnLNEc1UnGHfdGLqGFCmA5ib91XHQufiKv
8db8B2pKrlbq3bZNTQn4BLu8I03/yWdv+4zyfKHofC+O+WIUv/dlc9TgOUl4CxoxW9JBHjZsjTHk
W6CljhoBkca4qhseLZlGxhBSDabaVIng41wENf2absFQVRAht3FcqEfY4WYc4+u092BetiBNThMf
qkNeYovEFxQXGLkNgctD+1zHbJF+LoFCQWEEz8GoqW8EoKahB6h5YLGT2ewS0C4Bs9AaoKOHCyvB
QbdRBCWcd+ilcPF0EKEQaMZ9P69si6rVjvk5VRl69MbnaWyGVDVbpmKjuSmHbmE56mmJsU6lwQmA
SI2xgCAFaioFwKJ6j+Gwy1Yk5OZCV/U7vTmkgd8sOUDngkvet0FPmF87GR6dP0Se5zwwRqIe78j1
DRC0HXApp8OD3CyHpAeVbrod9NU0mEFCCTG8T7Hn9U/6wu1R+QzCEm0FDIoav0cuTgheR9CuUZ5O
PtgrcOAqFbbxjVpYCvXiLcStpQIFdHSlZpx9qon65OAuYjLIbwilt66IFUj2p9EID6b+Lwm6J512
Xq3d7F6PLICeac86NCSn2l7ZV41yZOJsBGXSlNsj4CLEvbS9WTAQMW+ok7fMQuBFsOLAU1GJSJrh
C/gmrFYo+DGDidR2TayIaefjGL7ga1JpAyPFbwWvNwe5ijjzPrXFSPDQ71/kIHM0z9lyrsQ7lO/u
8DASGnynOsxSd65g/RlUkOU8aaKD5ibFD+m3BZP1zJDVlHfHQwoSl7spax6H1ubUW6OgixQa4GKH
rBbq2m5sewrI1TzaMEu1JzrTbdmtPw+iJdlZRfOtG1Y9gyx2UJkW5MlIk0tlzpG2I0dXL2haGHkd
4ZKE5Mp7tUvDAZTOgzL3ey8sfGIAgRAEVWNDqY/dUy5fmT7m/yws+1PxH+q8upzVv7dTuq3BN0dd
sL/oF9RRPRIzLaUEf2H83XSgGehOiVxutjLLwbemjmDBs/qoUTPFX8GSbC1odoQrgcCdxwZ3m34B
yFIcLnhvMoflJK4VRZJSEgEuiiqjCrH++AXggu9+oNTPBtaS/txeCDBz7KI5SYMFKhJSO1yFuw6W
SWGU7204qFMfCkY/+28pDGX2yZKJF+sVp6BXlqyvUxfSSsoLBlUB6n9jFseDgcTLDp5Te4G8lZML
giB7POLE6S6PcmnExblBii+7M4xgb01ou4arj1Y4Q/adPDP9n1e5B/PQaEOgKcdOqFTpNRMjWQBH
viuZABjpNn3XwZEymXf76/na2sNZyQlrRqdPG6JkT+77X4HNrXX2FcPyGkmIXCjdk/yg9s/dEL17
iNZvEUktEG/Wo0pzj5qWOpPO9/0Tzpqfopk6ydur6KNlHUPQdVQ6OPVgMmFlQNzf7MA2QTaGf7QU
00KKd47BS5J6Lxj0BQ9T1tcvLmO2OinrxVECIxdR8Vopt9hQ2J3EVlxjcmtJmQsn7oSAfYP0Xf36
SSrsQQzS6NWluV2+5T0A+l8ofZe17hTjtr3OQ7NqQdDdvgfkX844XvtWGPz3+jbWXmLjciwGAH4v
b1+IBT8RAwJUpNvaYg2SiA+WLdoU//IGcMoS2x5IYoD6IjR3gFTb2G8MJXmPa8OlrcZRPSrsPRWV
7e1ams5QkfSkbsl+gF/uyd2hzc16W/aSyFTvttZADI7xje3VIVVjnfEUhk5x3IREEkf0KqGHa3wM
8k9s2/b3W0/UBBVqzFtrkGoWBd+ncVNmut28URj7Izu+c7j0lpx8s3SwdcHNkhn3KF+SA+088o+M
GOJHkGrMxRBGCxuHxEyOUnP89BrHszjxTdpRMOcdA5FtwbJDx8fVdew/fbQV+GgAiFw95YK3n13D
mmIZGFvsc3dOyJk1guty4tOwyTUIMow1CGIZ3PZ5GDOXEMNwoovjCEiDCM+fanURP9VltdTqzkuj
1GHrtSVMGzqn6tXxOXvWdrMpMSTcMTV6zcbwAD8Rp8SP50OtjQ6ucuoKBvORDPWVR9AaYGV4WhMg
Zj+b9fxIbRO29KQ7za+VXeuF04CWZlisoow5l4CpXsnX13QcEGrCucNvo37rCydEMn3jKh8j6TKa
EcxTzlZ8kb0ONm/rpMua2XiO01CHAD7PBQT5Toc+003aOQseo/GV0m6Kp6BH2cO98rl8ofcG+DJJ
7xI88OvSiA/9FHnjCI/6gS6c+ExmmkY6rCdPT/ab0ujcrGE9IAMSoGloOng3pnQPWG2dATM4sH+9
8rPKteYe5G3U9R5VMj4ESQr7OCqA42lg/TgtGpxR0fkWlEB/DPHLruVH9M00IwPqCyKob/Q/gS0p
TId3F7SPhGZ/c7p557u0ZSg1Y+g3LAzFiOQx6nLlLCd8pBcOgEK5bti81+B53twcIbXO4we7oeRx
Wjl8RG1BJD6myYtkB8YxP3+MqNNfKKEDSWFFG1rtz7eAhPylpmtOB5iKiX1fM6Jl0TgmA5qlJJnt
+F8NeRixn62NYxi7U7q3TvsiSlipoUYX0w34YDHrX5fz0bIIJRE86qYYLUj/oRHLABoSQPjCpRyv
z7UG8EMZm+7xq3MGzx96dBEp0yk33+AmETtDKPVikCeOEQep9trWZfmroBr0vVNTdes/y7h6Xo+Z
lLE6D5ao76FWR8kU70979Td0xJLnZCNA31WBzjnb8bJ5q4fIEr3UkZ1r0x9E5fUXEqY6lQREmMDE
VsNHsze2mbDh0EcBdMsM30oAJAtt3K2rb9DoNVBpMWLjff77VC0+r4y8S0oqLMVLB1t1gB/Ty9C9
1De3DWur/rDXyQ52RydjT+BmDN0XfNIo0aHiBCigrftbOBuVcTcig4wDXdEJLTRRqSmjjirvlRDv
Gx57Ek5bYg3xfH7kF0nkWqDzE5L4CG3rZQalgjos4jJvKaWsptJ+8nR+H637ueyCQnXJHfOR22VF
o4gV04fbFDI9DB+OGY8gK5pOdoMgGOpNcRZRql0JqISy4xDKBHpcmMvHiIR+kjZRnCg6Yg+1GZCd
5YjF1LqhZi0sCSGtf88WBF2ZU7HmLkEeCL0vBgIrSyBAY28hYcjI0DlJ92OIMKYMtpAI432YFPQ8
BKSlKcuPsoCG1lsla6oQpBIzFK7EL2JTsoi05Rbx2FEHmJurBWlZbyrOTGvm00ObziUeKUiaOEaa
pXiSczv7DAXiT+32NPPOceUX0xzfhvF++t9hz3miULReb87ak9VLsAwxFrrXdFp18UqEATjReW/u
LucZZl9/ykEv75hCfiuCpdHTPw+9JkvMaFsLYvnOpfGqboyapVrWZ0pi0rNJLpuNULOLtGcrXK9u
tcnk/02IiPzvooqBR07L+Hx9bjX/SdvV9Wk/mWxBIQ0CxvBX08G2N6CrBondqvVAdWJXWT+U6fT2
Wff2aWINWreVBR4II044mxf4od+ZypWWIF+jtFtzJlxnG5FRM61vW5iwWwcRRyXtYX38ysUNN+He
x/a5Gwj+3Uok70UzATN3Kd481ahd1/MHQQSYGlOGM7ErkgYx5+rhqmkNCGBCfacfL2rXT5IrSZZM
I5TQbv8Kw3kqIEdm+IEe2+RWrsrRe7nF70nunpIZL1UclKbNMyboqBV8hjgf4SBsuEUlz2Tg8wm8
Yeyelx3c8I9VBwtlWmBb7rXyM8ZpJ98nIG7nBou8QR/tfKz4WZzsdBUis6zmPjN9jwG5jkXehAC+
faJ1x04sXNFxIFZdd02ROvJJzIlLfIHPP46Y7LTAvMMd+1yHkm0ZzGONwRgPhMCqAmZ81jDmpq9z
cjBClGDO7CT2F0dHP6q8/Ntq68sAj3ZF8m8ZVw9VXgtsHKQ5ayMaMJ8+5ZV8KrnmHrGcUau/2jUT
M+df2EnEb4vaEc2NcPBzPVGUuRhdBIgiP2Ux708aRymM77whtQit5K6hy2iDqAFti9ZFJQvN45hq
4GP3+rI4qvA7XPu/5CeZvyP2nNieiowucF0zVH8n0cqM4jpjUdYLrR8XIOn6hiLEI1NMLbawRocO
kWgoKBHPLKFZq8+h/cHyFMo2QMV9cchZS1aY68cy0XGo8Ght1DRvtQve3JaNEw6YYCSFgG+uGXfI
gCq1074JSGzPhK9+Oui6yS0mVGy5wCTYgN1Zs3xuRHKIIwWc8kDSjPGTUW7coBcZzhSDtsVkiJRB
RdgXUSOL02SRpEJTJYftBbC6XaJFDc3sIhFNmQBgF7cHe9SzFjuSik8by9Tpw18XbE2I9ZTB2exp
K06fHb9E+J12vJiZTAjm+SIlPLaLYFYEJtEwSlYgv6VkeXiYUJ+R4ijNOzqrLaqMC0xXPfet5XrO
ajV+JVbxICdemcbQbEC6PAFVh7Dk+PjNlhfqlQ362Yf3wGsLd8T293k16DKdcJrjEsgNc5kB+G/M
ulbNkPieUcsdjF7zTBM7LIEnbp0ZpLBlIDYE8gMGaitpZLOQikqbdmqbUDK8XxEC7Ydfs2Pb3P8U
6J2sW7NuSWuuYMt7bOBLjWxo2RWB9e1FLnh2rN+gqJfJSbt03rscAHP65vWaiIdGwZeRH096rcvk
H5Uh/uAfQdPxuenAPHp2I31RFQe146jHuATttNCdxe7CgwJFOiVisirWddPNhLla03Z9cCY5rIxC
VuaXftgq1VozkH8wtbwCrC8L28ysgoWw2lm9KyjBibFDGGRPKW7OQ6UZTYv7vBi4J26aFkAfoiSb
fzo0iSE0jRNNG7/XWtsMLgVdyro6x2TAO+mYoXmItj8JqxPTFvN7V2+CwJrt1Map5TMlgFyBk+LZ
Oolr1LCdSKVQrFclp0UYQOuZSYLK6DiLNx0/cgVoRIedVlayZY1BniViQGXLi1SNtfIsgPyDSKJF
PNlSnl8s2K+OkJInfm4h5Pyq8P/wSwgKu9x7fDsSx4fr5HYMW2ck18UeK/eoy6SpdfxUW4sGC6H8
RoBM4Tv2HnhZt5I73D35NR4K+qg5j1x6V9IVHWg896n3R8nsyG83U4oWl/6LZvPmemgTo81M3h3B
5c8l1kR8CRhd36R3LQmKbGVUlmHoBV+oFkkz9u7Mwghfmwie23SGtZs4Kknus6K+1hc//UofVxwO
TogB202LA46o6KUAtc6uYqRi54GxA3cT5KWMZptUuD+2KguZY2TFSdYLXTS42/pErtkxpvT1wr1K
TgbKFIqCxla7EvTQWQsi46mCehC/cf6RupBp6EbzYWmSZ8EeVaxHM5y+TVs+Lyv6taCT5am4EY2l
NUyTyDERQDwEctMv0Ubsg7nxVB/XfBcHM/5J7EkFyMZNDKfQuqLNLi81tQAQkfLOJtciNMvJSXA2
cZM41T1kmF/9M8ge5SJGVfUEWOs41yR8VGtZhKy4hOjaYOj0uPcPs4WHYmGcjE8aDTqJpJEBCLyY
Ef7jG31FjZztytfyu1ROuBp5vxHzWJUM+mdCIdJklxcUYbFAuIBsbYUAomO8dZay+OwM5sed+s6E
DM5OMwscaIRg4hP4FyP2TIaiXPfBdEq2nMNEn/kZaJUtG+Crg1TfDA+NtNp+OYWfZx/VYCDVnQfW
jzQ/QXTgdOZZLPp+spCp7ttkkNrvhxw4YrOQLshvKd07T786YmAmCbpHztFc5gTgxMA3CckQbaL2
uy5AX8n1NqSpkvVh6mb2rQj8ftAUilb4GBEovH+ZXtanBr7xB8ljxduOKaGFhy47N2a2FedQSEcB
wJ4xIB6ioDEsvLw/nhnjuBzCgrBJRk+spg6zCvHfKGkl41oKqNzU6GQkqr454WGQKCkHMOAWoBvN
9+P2NOm5eptLF5o/9Ryo+H4iq2Y6oix8TQkgnUAdUw5VZ+jb2KH36Jlr1/IA6g80tOGwJcMqrM/e
RsEcMYI7liTyO9cYRS4nG1OtcisSRmjmDj1wdPbFbtyx1UEY83UGcTEbnW21NpJbnU+sG/MWoB/u
7lLBTRaXAH6aITug0AtrSUxzxRpGrLKtgTOVTWSXA+05SeJcGJSf+91S53vUpq89QmdcpAj3JVNz
pJT9Keut5EADkktMKqtuLltudCHkPtl1gj7tYlL6Y/KCYXyKCC/YVQKIRoHGBV4QGwis79RpY1/q
ZhQFDbmTgCb35wZO1II4E+E3JyA8yaEEE/3SMjvL8DvzmQ5AP+5ZeyqMBrT/RIdaJDoWpxG25OMg
9fUeANVAIi2jdGOhtkLPsMd1yc98+0RTxJSFCePY5ramNbboSKMr+5/8SxEZi21hvhK4vv9r2+nP
8QgIQoElT1AreyhCIEO4Fd8SYy2Es1/bxScDNjjaOXIzKC+iZoXsZ7qETKR0MqYpq0uVL/hDA8TV
kLAMd9o+WQynu9RQpStE6kZg5s2ECChtyCe2ZgEyCYuhkr4u+JWZD54WUVn9EoFAPlL0YrTpji35
X1WcYa9CYlOoryJY+c9XK3b4ruN7GONe/3fxXrzUD7PrsnSU72i+oyNOZ/fB8cT7U3VnnyavmJ2l
YkzM8EWuO2kf7fHhZuQfaL9EVMUw1rWVy+X/dfvaL9N6B9ydlozpxFM6BIGEO3fF9WQNFqui6R57
HjnAK49HTT847Jn3Xx5ZHPXIgQeGC++6swr5GSeHngzEjGThr57Dbs4upcc+UVDkVhuBVfphhhiP
7Be7HB+Q9yt6qQPucLXhEjU9C8sLib6eF/Eel95lBpecs/kHU0LyCa2Xy4g3D3aVSAlS4aXvDCOi
3BtjV6exKA8oe/b5gwuoUb25otwJQ+J9NSSWqlJ7cAJE/sQ9trxZpUlHTXNMeBPkqsdmNkcOKClE
LTU3oAerFFNpdLZANO9F3Heq1x0t4CGmTm4YxyrMApZxPUwCv9iyAFq1KCz52ws7/nJpiVl3TqmL
VXN64FbvJf60719OmdsclLQVwV/GiyXlmAUcml7hgBQyB/cXND22tEbVbhl2TTcR8f9JqraFSUeK
cC+v6yL3vpjDLkDh/QU44tAP1eDtgdLtiorRN4FCt4bkWvJ6hg7oWa9yddLwoG1dOKxTdIFhoSA2
cYwd/EUzWQMFTOJzBwvk5YCatrvNoHY5jzz3oT7J7fKOxRh5WuF5vIhrRKNl8yTVOdkf7+kDcSX6
BzMzHKs0ZqNMGsC4PgfaRKadLgxJ8hhoFI/dMG9AwBS60yVloPMzX1dNZjS8XHLf0tbAWDh6ZVZ2
8bwS7o/3bJDshrLDk/ntfJhZ5nN2MZ2t/G2sLElVmYPtIYQUl5HjBMSM7q71U0QFQ6ulrWH9+AuF
16LKTeLcaNhWBqa71fiOKpKxdn+TdweTGhbq0IdSOScESxFT490jWGh7vdnrcAbTd1v3qEt21JRo
TNAQysxR2flVcUTWz0b64JIli/Indizb5dCTGpsEVtIJzpVj7wVOq8yn64nuTYonMaHKhAuJ2mim
Ei0uJwvJwBsofncOWHK+r3l/qRlNusWeo5Fh6liOS+VvvXJ0ug9FD3uhI2j927/d/eNXosStqJZl
yuLQptxkuaYaHGyPtxOgSMjK1hkLPuyFZRSAnbTGZ0tFQgpmCezGsSY6xAYu0i2yMy40u/9O8R83
JHjWOFqPiSk3gdePaq3HnVFUmVs9NHBNEOB/jwxSAT2yNRO9E+UDOdpv6pKPvCjLsWYN9F2Q0go+
P5DiLMoUgsYAeaTkIdw2FvaSj+DCP1pahELhG/d7OrQoSVCKlpVALUcZwTlO2Q4FPmLc4KmLKSGJ
U2mbo91ZcxcUR+z6HxyU1P0FPLnl7T3MIj1D8Wh1xfDhN8wijMeMviIOtQaYMB1Uu6Fht2jwkWcN
ghPfMPcsS4+SYHpeoZ01q6ROxp4Xex0XcWD2OCB44ocvEN2+F/1aBytXoDAEepMr8DtrlVVu0Vp0
DHJUIORBvHvKxZBO/YAPwsz9diyugWPJ2oNPSikFJ4vlJDcScWiUJnBdpq6D6VLnzXTt4nu+gKbM
W3AcA63YHArAQFTQFlcXSaDVk/lOFxDaIHMdW6R+dirPtTJkUTLfuf/qS+OdOsDSozJ90e/41Dhb
9KYTiNYf6c/C5oWPGsLNl/q5oyFopekfXfVRaYEh2vrMsn24qjpG43VM4Lpf/2dss/NfaiYbbq73
i+m4oYMnzOYryql0kL0l1qVt9ujxDDVoURZLOJVAEzVxmnTxTJsUklezKzq29ZkC6bLydgc3B2aK
mHlcN0RQtt9QrZZk4YGBipKzMZoRYMUBkm6TWrzBH3jPqF4+chF+EgJ7lI6SlMuZlXD6pe6f5fcS
4V/K8iUFEZge78aby6ViRmep59c62rIUIlIJRiow08ym/p7VjSITY5bqFfwABQGI0VJ/Ro2pPGmG
cdGzD0Edkvm5IaZ8663X1/jBJ70pHAdxyn0YOXUOBw9xTbgh9mhCRYozeOpxZ2NPbI3mIme8X+hv
ML3L2TmJTvMJIofu6iDQjpJhcQIWGhfkV0itZgDQSnKFjkGUQHS4WPEix7jRI7rkOCnXxM+jmGDq
8PYZdBwXsZURplX6fjobMp1AC6LhnWAjClFjrT8zVt1MoT5AntZtLDSOudKWQAPLZtgsO2XWzrEY
2Mku3u1WyQHTMwv0oP99KA8kMsdB/xUb5wmoPmm5fOKlQlWTmdzdLOiealxctUKlfHPL4EWZWTed
11FefuSQHzxUyTrZJJGTWaDVEEsB/DmhLt4HH/BrJcAXWQGxIcnCOW+IwAsm5EqkTWAmyToXqbVg
U54EFRwtLkPdwcQuJh3AyOUQfED9xZwinpiQyDdus9AuKfOj0UYsk3MwvruIhdkwxEmtZ2ngAc7S
ep0322Qp9iG/bGISciRAkzvUs3UHiOIuIEwNXQtDPe8U7iZtfGtJKmqvzrtfqVRueTjG8Jl+tSL4
TUda6rfzlb0VaczLYt12ggSwuhdyGmXPKL9ioHC18W/S8JJTtAGG825dVfJwkol6W+kN0qDuXWGC
5Ns8zQBWxQe9OLNDcr8TUyz2KJzjcYN8vUr83eFcScSd06dwO/RBsr0b34ornjXCs4RkQaCQfFUZ
VnxB1xzASLhpvy7zzZKkry4AQLBG8/2Fw8PaSYCf8B6BpL0Qhk6OvxXrCbPpnApQYQjcxb2BVrBI
Xt/NB4yujrStXnuvSEvRGtpzhFL05DhMDgPDP7ChiRm/oXBhKzHJwbbd+3VicHGtNKAD5Dlk/5uS
VHdRrB5UJ6dfykXJo8fbTN++QBK3OTBrup6tiZevPDIIwScESJ5/2DcfI2APbPTokai9vmVNqo3K
c/wSGc8se49a2zUGMG3ePvq7jRCLoYp2BDZWbiaqVw20Be8z2sS9VNQYJmoXOGV5vGWQ+wXyfX5m
nyBWLgi1XJ0Je5wfCoM8a/q7C1Yts58YYOWXfN07KoD/8n2Lzf8FMCuCRfwexDWt2Fh7QY98hms6
bhUsEUJ8q+uZzfposEazCvnNboVEUjNvXpWuswVuX8P2swGmFt/qHY5w/NAFojU2sHQ+J60OK4hm
SZ/iq+Q2K3r3D+JTY2znBjP9/aKPlKP/GwO9h4PywpI60Y3OFGTsp5g9N24S80FaK4PuWPyVUvPv
dJERnMfdwi6O4IsEVMfUbtyhLzsEfn2D6F360WXv2X5UXHMFD2Fk1b+5FiUQ9OiPAMAsz9qVUcFx
hBYgQD76x+MrObjL4DNpbwAncy1z9RwoQgVXjG7ZjedhoiuXZRYLq+DiXUHnJ/Hc9qcut0jEbOWS
A9cchCSdye9LlXvxCwFgkAJS0r0M9jnfb1bv7EdY9/yLa2y3sUOs1VEjQrQanTPrTKMDWjNGQm5f
D1P9+hrFDxjKvQbZ501/JtLEmMpjR7LWeELAPxajkL4BhKlaues0LL/3z9qynA2cuaXO7UwjNEbj
1C4llDVpvBNa+EBVi5qjinRdm37Jt3rC7z/TGKOgm7trwmUX7+7Y36C/LZmYXuIXgTk0NjDw9qJb
od2tTsBbrVFW6gzwYQP88iN6vjSfygVFR+boR6oz6b+UeHh2QYWmdVbc7HeBMUYyd9I0aB1kXoxQ
eFqA1Ljd5jbVTqzdRfIYnKRlceNQpAv1jzEv2Nzju2A1Oob4Fc8oiMLXjrL7CJjCCoY0mD7qeQtD
4qEtUhtgs/Had+uq//jiFTqYSkRQ8zQJVkdYexegkpfxiM2e7a97p6X15hJPCnNGigG4r0qWy7ut
2QWXFrQiMc7Acg/eqorLEl5OnsJDK3Pqg6yS/dRnWsUTWfPsmU5b+QApcnEEhwecozheD13JyS6p
se8yMl4h03Wj2nNhUzNh5FPK+60EPjLDMCuNRBivh4anUNQxPE2q/uwpdCAp6qs9v1ljdkmjvUQM
r/7DeOt8Dr956J7xUh0/repXE9HbG5siLsqVWFvLrWAnhf7jkIMgnBc2Q63Amc0Qavn/SlW8couW
Y91+xsPNn9peJyK9j5ObWO/TAgqeM9Q511WN2ZmiBY4vWkEtlU0LyL1F1j6c8GgFjToiFfyRxgqv
qWaTlWpuAadruS2bs0bbNE/mH764qCYF3Xlp1PtcaRrDGWIEiAAT5e6mg6gXtFE2DvghDbsf4bJB
dAt1FM58ZiPi5WahCFgfgt/S6UL0oZ6CBRyH4wQ3+hOMTrNrlzwPfDiLaZdrzCme3MnxVKJixnhh
bmGnA3Yc8Kg5mB1gMd/RxLs+2zuw8cwUeXiqU2fQRDp8jdwwiGi1pzKB408giWUoTcn6eCen5xBH
GyJFDBHW6T3F+0KfzstXr/Yz0RUtoE4k//pGMQuupN56HBnycP9nTkp2rcioJ0HKLt7ojTvNMxdA
EaeWR1L6yXnBP7MqrOgwY6bF+TZm6EAhz7FnjyUNHlP6YXJ1Y2RGW9XQ22IpaYHVh0Ea6JfGIZBG
uj45VH76RVFEM6mD31k8CJ5urT4G/tHUVim8REXdHsVG9NTttimQr3y+oEmMshjcKTWLBhVB7cHd
av/6BTESRS9t0NmevVZ6QLkIvCQN4JzzFdoFqBqZH7DggexXh8ULsIMGgrkTtzj2jKlriLUOmpTb
7Y58QofIdi7Sl6pRZ/yIrdmOY8D9UZF9ScjblkVHPN/VdEXBfmBIliHHurRWtYb3x+d81tMDDJ8l
9OBzCPo/s61IntD8obl8p758vN8vfFxHdW3YV4yav24rAWcucMgqjBYdl5tsouGrFHHhuyfqiPMy
YUTU/kUA3w4/ZEvqXnGlul7oX3mcmTTQXCY3BhNIszG45f0ADow3EHhz5iYoK5IatkFNqmLKZiCD
+WPqCoi1RHcdILU2MvCByQAyNT43OjWKfPdYLON5vAx2qleWm4TCuvEZZoxLYUOP6eNwzeBOp3jy
Q2Mc5PSTnlmKnGYrXA13Z/wy9FpzgzTD0L2Vom+ofPfLQh99X8Qk/BM+tdFspbDWP3AJhHN7Jp7x
aVLkzMfSWxoxbiXbe9A5etv/QIP0ikD05T5mIuGXHCtT5YaFMYJ6F7s7rxskBbO74hgVloLYx6uG
kDKIq6nuvDhbwz7K9GnQhF4D0j++tX+Sl6UF9tILvWhG3cKBOi+QNA07m1BrUHoJc9WhmddL4gXA
Vjy5jl1q1Ml2FwXHaIHRmEAPg30+BaXVJR97a1HV5gDIWmqYhMmM0J1y+VvcU/6X5Ui6gqEwC2dt
3y6UbvX8fwuYOTRaYLnt5wUxKnV6TsLrJ6ikk6VnrDNN0oZO2RxpUjPvK9tcSG/ujNmO9REEx7ng
A86UXrP40DbTgaxZNzAEgj2DV1r8QhFiGpEUFgynbQEX+/zesfRwqu9fNRP7zRoVYQWdgoqND3VH
6kRkyv59OmbiSmjqYLXKB3n/mQE243QoVLmxnA4i69t+RboBgpCaJbGcdxHmEvvfkGJnnfgklH9y
rXCKL4R6G55jBQv8eHh2WUDFNzB5QEj1vB+LpZZbhtOY7T+joz0Lmd6QAj+n+/iHiAa7Ty6QuhVZ
1cBqGQMuOogzKjJLhd4xuNNDnxTZqRfAKfAQuY5gzFv0IMH89jjS3TU5tIvVsESNU0Wpwiji6JVP
bL1ldoSQWpg7uQU4Ir/m9+AfHTq6xGwp4ii88m2E6C9dxRYwfRzAlvATNUNoc+6GTg56Muogl4pk
C60lwsdPcglwnrOfuDy225bBN0Ihbefs3rnvC/VK9nO+uz1y5WS14W1Ys/xw/ekvXWqDqBoqSc4x
TYQwE9I1RYrrQnt5V0gXizNQYsxZF8dGB4QalTPfmE8uSuEj45zG8VICtKf+tzhwuz4mFUCKzwxF
U8Cq5KdvYfyn5Tu4dvLoJkOg8bafG4UuVuuEmPxDFW1Zhxva902KW0MY1IxR93EVKY2fa3MJ4Ui6
je6plGf/HyOZTZwEx8Dk5P1Dm50qOTkD6t/18TAqZt2dJqR++qtrBujUJKGIANoI8vcQ5jsUD+/n
PpZQH1VYDS8dhGOMMz48Lv1DKeik/B3qJQvPUDQCSUrdJNveKfwTb6ArvfcS+jHwI2uADEapvT5B
JuyZrG+Tw/csX2ndytEIcHYxc5QrQ1UVND1etnCOGFLQ56kdLu3Fd3f7gigNBWXLSXjcBC5HngtC
1UldeMHt8ciiFKQR830zQwP53m5gmrcHEN0v/DKwhfdypSREO0rEhf4FiagGItEjIPoOP+WWMa+n
oLiLzAoxSsrwBJe4l0iogkWwnYpFS2dRdd6OU7fpOWBJpYaEKbtJPIG/jMvc9ng80YQ+Vym3Xypf
pAeBbLrAAaMlUS/PWGhv00aKlZuv7LUafGLZugH7Pll9J57uH0QHI/pu4u+lsktJg1N0euOYADrh
bFwgDjfhF/8KH8S57B/veYZU1TFnKCalicvAEkoN199niMj4BvxwgWIGsz7kWnoqUhIRs7KlDGMU
L3WvVyhnobHoDwON/3RmiyJvqzGqa0n6lyOGyo30PHOnwzCICaRUe4m3HcGheQVFxAnekSfggHSK
SPC3Soa8Rqmob4g1+QHi5knY88/foQgGWboGTHPG1Z7T8WXfiIuutpg2kn46RzNJmB0N8rbE6Ckz
0xeOyaFJnmid0tQ3DNp5Id0mFOxTsAhpLGvQT1nSEueJzxn7GjpT95FL+bngjpkAbgCmBywlbBZc
gBNpyW364H/wB9grWLJLwwUiWWvl7Ax/W/hj/kDclP6uBsNDyEiDcaESRvOrHkl/Lz4tBPpV3qmy
H6LN56C4kJ8IWoVOrs/QHYFL9qfUx8vle41nXX8dYJKfKiTX1d/p/a7n8PxwjqpNFKMlwzNMKjoQ
Hb1W5vgr4XCZ8D8KzaH/zdVCIPYtgWvpuYyPfEonybg95G3Ft7bvfAV2P0uemeRUjyV2Cpi17Ou7
e5QEri+O4NFByYcfi0HrFJyq3jU1tV0CAsZenWUyzHLu0WwFv3BcRgpOiPNO91DJ21R0QzfXrhAb
t7QpAVo493WtAdgmBOTc50ljleHulm1t2mPwEbhXEXLouyUv6V5e3pv1cMwg8jZkYESrHjcMCoto
uZJJKE62B/qu+Kdz2dqCDky1jSCLXPZ9F4gqSRUd34tvptfksVmIMZ2n83bB86OYvM/ORAh9GWyC
F1nnATuBN1GjOuFVR8B8FC4KXNJhauhy7WYitqi3fribE0v+kuF+i2WKKY+qD3JzpJAKn6d/t1Jl
fkej/cJo5Gd+IvS6dgxHG4aRvjsjD/LGpAb5LFoDVXB7gsGrba9ZZ1ufjffmyqYt3DPSDfvnBv+a
82RQVWAjKrQ7ae8GeJQD+Qa/ne+OEutmKlAxqW1VS8cYkG/JcQGZqSOnQ59KGTjJs2BATTPkX6L6
vpcPcXh1ppmNfV1ocpz4g5dTxE/cJyjlDxXz85ZMdo7A4mm+ISGSv9+V/YTyudzFMAj0MMM4GtMN
+tkXUPdYJ/diSm3bIimNhOXbISC3YoASRH0R0OLl2SbHgXH3pJ/HjmICmY9y7k5VoVcVT72ulPyZ
n+CVlUe82gBlLWksosiIhLMuDBuHTftKdGLZxgvBNV4CNcyTwRhyBmLJQCyvR+pjfidj/qJzWvGi
bFdMgr+dIYT5yQolcR96cHk6lk/K+54lhwdNdhRSIRMxEtnYBq6nvXoYER+tHs3/iyYQiNEcS2TK
BR37bbOhQkDvhCikg8YbE2bHIc2M7j/P86rusMJ7TiO8teYv6yYtU71stGilHmFsSG6QoOCXaVce
/DfcAxinTlOjkE1jIvA+8TpSS6pK5whFL0fP3iHaDbZzGc9/HdtW9gPVqHoeCrH9RyAw4Qm2Gjba
rUC/lXYOS9e1VJKIew4xofkfIo6pGNu+tvIWAqGiGYbZCuKksoz/mHIzeWJ29mH+dmoALZzm8SxX
E1TuGh+oHEzNv0k1d7aNAipsQIMRXZxDQFIiieS3kc/7QQxdKoarDeCoTaVxaBdO7A4i96In63bw
cXaXHqmwS3Th+K9Pgvbquyejq9DV/8qHV4FtcCJRUk/TCgemhZYkAB7dKnxTMoVtHauO6mkVAEGq
Jsh+r8Y4GRN9GqKeTahE3ZSBfsEtdjqpB0fbrccHv9z6UgNv2MOfkNuhW+CuT77c3PhddgYwbMfx
vi+6XpmLv0ciXs6reSN/1V6THQHB3UGEKRH5q/aJcyQ6taNbE2gCpaNHpwr+YNb9HrptXZZtvo9g
HsBqQb2BkL/HJS9a+zw3RO0YB/wMWaTFtVZK+L+++eKZFEqf+5o0y9xDTE3qhoCT4soyNHJtr6Uv
QzWWyNGFiYlPE7lIoN/ITqmNmGqA92fAgIwrVsupgwVdLNcs2yLLEE8jJK/CO5CLTuPwmGCVMVwM
OsmzMJDjHFbuTCNz9PCkWoWbgMxr7QKmED+GUBPrSrt+UHF55uAfUTsLGOOlxZMcxZ7nzFdcCLHJ
nT27go90kZaqCndcF6+l+VNPBnge0vQpOlpezDwwIOg9Da1eTuKhr6FKKtKCaX4NYcwnrsAQR13B
xXP04VpyDhfqTrD/vwnRUkk5SmCoVTWMuPO9qebbyM8Ol98NuRlwLM52eCcacoMOwYBZtYGnS5vK
P5TiAtk2/1QDqDc9ftywWePg5P2goWfgTSY7EzJh6SdUF3tlW7toddYdtXrykq4cZkWGiobm1TEC
nsn1IQECioA9vxjHjf9ZNOuglL1rLkxIyuMyNiPs2nFumRZ5jNyzOLqP6dQZVU2SUC5doe4T9b8p
JRlSIY41OqasJn9agYTmN5IYgIDczl2gMVGoytLrhjfQ1ClySPenNh4k/itTNaHu+2dF9fyhHmAi
MKmx2dLYsWG4WRJXRgcNfrifsbRcktMr/8x0lNcejOZQrFShY+Q4Y1zBm6O+OpoUgNiWljmicBOt
T2mfvytA8hN/rPAo9aK6KZH9tJWncr4n7272qFBpV+IIU4TQJEVPua6h0LK9Sg62H5VVhSYAcNWX
a0RVmxEWQR+NgFRdaIDuL707Z1PRijnIs9WFBmPaGLypJrVg3BS7FPNoQXGj34MUZAOu0zcv3esh
Kwpre+HFwlRWoCXAWSVmEVGg4W0ze937yqZVFLWBSMW39iqyRhxxBbnFGAPXVTdJIoXu6LIOEV6/
lu0gWIB5TTo3EHLbEn4Nph2gkR/312Ui5mDkuNJCNOpvJKKTFqVSGTGYxSlltuRhnzdycLZFzBRY
pzgVC4nwrj8T8Q2bJQWcB8IifqPGxHWeNa6bnC0VdZzHbEdwWjPC4AGABRSWYMFqNwO7iTHBCzsl
LRXJ43hDmuR/IqmQfOQtCjeXYSzX58ZsbnBuEAdUG3UaMP+0W0fm2r62B0kr2no8HhNGbPwKg7G9
CfDNJ5Jx0MQqe7UmFw0g5/BGbAE6qTwf0Y0lr6AORyyEqeD/gZJkOjyiOSjgWCG3itHl5UqyWbKS
bVwwqaV23zgWvCxzxCjLoH3uDcZNM99evFo7113qKd0lRAWnXr7Kn/3i6+ACLZTUgk/zfzCcYzVW
eDG4oWV5YRYR6gDIZXGi+o9kuTJKJUT9YqHYoZyLTPnk57DAMdb8+RRsKppUtObgzHcF5nk4RwJ9
XgGfs6LVI3zfuCn/+3BMoBF0qklAm7R1IFGP00qNV6un5c7vio/cf5MuLomCU6z3qPcqyCZTkQnu
fcsO2M0J1nRIKy155tAt3pMZ/JHRRN3RTXGNyTys89JYFoqJ4nhShSzHg+MQSJju2PUIaOy5Wkdk
RLAoqQ5HXOXGVYpzmhSqvwuFRKtWWljNga2hRRw45QhHcnFo8jg2DmqJl3S6kGqxlQ8kc/hkablS
+reQgGwgi78HQke3nVhK54HgboooGcWNmbLqgjLlPfyEmjfhYoWY27epcFCESf47uG+BmQloIlyo
Ql0yFJYyQTr2cqQh0xRYqMKXstwf+ntcX6Ek4gF1dNey/skEQqdmOcBV/HSZPGkzZ8+6LARGkD59
KltS0sgkvnjf+S9iN4Y5gA6mdEK7Q7Zu8LDBf/j+Pq1oL16/5YlaKLw+2fQNje5dDkX4tjCpxRwe
PHMZUAnbu2LAqfY/TlRTobfqo701eqM4dSRNlcg6SxPng7QQKLpE+HvE7S92gGi24u5ar7IlmJt2
aM8dqscdj703ukPtYKG28xgs9/iGceCqmW8hX+f1V9p+RqgYQZd3FGq7qyf7nIY5+IhDnf+20ty+
1jZrE4axQNlK/t6uCbm1uuZCMKr/FsNsBFO8rmmjocHbnak7h/nqnIvvfCO2AmdMVnxJ4S5augk0
+BNR0GzVr0UM4Esg4gl+uii6EeZx2JzpoiyiojKw/h2Geos3eVE5U9P3dnVS/k6+33C9zE+9gI3e
a3Hc1efaYkOp0Xx/UQ/f4Ou4NpKwy1xCEoiPYESW15XFTJsQlTAalfKeellCiIuHtbVDO60W3MgP
chGfVB1MzOolgq3GG1QVOj+Dc2DPNoexkWouermmoyeG+T4kOD3/faK+DSGWuvXiNvNOtVAPKzdi
eaysunIPP819c5K0XRvSAAX7bhduYzd86VJDU8/gymTyqGlY7MiEf76By/wRhx21uzav96Dhav+/
AG1m+RuPOHVNihf6ugLHdWdfKqShIza/9do2M9W9P7QHb2RPTnD/QcYNWUYMBHZMOj1kT3HPBSVn
z/ITRgHnTh1y9uul0LYbQq0FAdCfNUG9J0a9rSE++kohvoR97woYH1iCNingU8dDb8+n7Cohak9d
QKDaPBb9Gcx8pz9x83UnxCzX7sYrPPcIk5jD9btB2RWevIoFyhQCcKfgLfVdzwT50eFDb1C0dZdX
dqr1d37pm1+nKYNMmRwoFEY/qjbf2Kyhgs3iWxDlNBil7+MRGf4wzlU8yftpCvtb/JgOLv4LsX/o
2pDDV+emfDCpzmPqZREWGwHlEvjzLXAKoyOZaYGaEfwhSbKj91LARfr2smKKsGjHo5cYYGIZYPDg
wsd6nPCE6RUCl5a5ki49jPa7OAh01dJRiAO1t2PQCQcD1IfHDN5f6hHPwH+vrN215ZGIJySLTeLn
ocTiMnI+qXK15rk8W1tx1ON0PT42ai6aWWlc8UnmDnZdqxDcABDJLY92jFrLFHTAz2+jsOuth5St
dQqR8vCRRqVzLWD4zDtF+ES04YG9EIDI6y3tIoOKr+sDG5Y/JAMy3t2KQRIQ6huMSC52mOe+tA8j
d8Vn9Qm5W/6Hok3EKOM6BhVXaDtSEgAHDLU4DcKc2sCszq47YPi3TJeLToXplXQrLoyAnmS5F+fe
IXqh9IEn7tBIqF4k7XYDnnsP9M1yy2Q9Si8UuMUbedkCrSS3mnncl43d+rZsqMIAiaMylk5Rnjpe
c1QDjKTwpiAKQNhQFk8ypSQdbthih6t4Kt9fbeeYLzvH2O1kvmYVQnMHGkTqpNV88tfGf3Pwlcc0
tcFC5PwhJfQcQn7dJhcrBRl+yxkcGbdLVMYTxAzhFRDgL05CGC5pQQARmshg6Wh0BN+z92QFAfyX
+T2XaxIm0Nl9SFs7RLG3mznw22K0HtGwfmgIYVM7E6GvGjdvl7B7XOT4ukfz/Cg0guurUZW77pTZ
4nlRhwaR8vRfdK2qdeokvEnpfsJLZg26HSzg1LaObKAoOPdNWa4kmIhnpLDomogTDGPfaPplceKM
7M6cIdffox6n+2Val83AMeUH1U38xIvH37cn+3v3rYB0p3Yz6Ab8CkGOwF12qPAHW8B2axQOU231
DgtlxnYtwqr1H64IyAOAgmtxM8HIXk7gH/SBXsflIMryWT4rpAbaseXtbr7ywTFj5jDd2HF1YOQU
Kvg1nA/2f4scH7eyiS5Km2KzUCo0jJlKyH35dR7eV+vXmS4jtf/5JdKJumSfKhivm4LQ8b50hhS0
U7oHBcxzycykq32fMkS56Mo+qhWw+3CG9fb/c4/e10iiFRMDojPYT3QfjVSN7kdep7Y+/HZ0hai2
8pQfsFnERzynMti9w75H9Jwy1k1HEobVbT/EN3aq0jP1inWS3++UahskM6Ae4Jo+PMEPX9/jHpOq
bG1GPBPaMtTkl218DNCDgcVN2V1erlQillF7tLOCGjXVHH7sJjMvOlVyUinBvGizDJPlQDu4tXsq
UcPEwZEYm1RtQ022fsKortWqEJq/5N6pzo7UjBor6EZVWJeKegrNZEoSKdfYKe1BgGmNw9X0wZa/
b9acZAZnRHppKXPIo37qm/w6x9BhXUqBjqiPvwlnu8zWyTrFNGfX9ru3Tc69FDCJbQev6m+bjhVU
KyP2ogsI1bKkKFWu1bqnB9gXQyrg2wUGNSSwZYiHI8FL+ovO3OPQJ4tejouT7SFQTwmJ1msMPvJA
W9AkgZjBBOFsWZLXEH/moTX5SEVQPLRmomZpcZk574HJ3jVE9oo8eE0hRK/CtK9Z04/Tfl3lMFBs
bbluA3M2dxf9bnKXprePgGpgOGIVQcXTG+EdGd0eGn7wxyG9ocDpcseTBbPSDvmDkChUIwe+XvCR
uf6hIT6VbwwV67/oc2Mn13KWbih4UY8S7xGYuBQ7nTNFNo0/UNh9/Dq6JIz0kBa1N7bZ9xukjPV0
sNBO4CkvNnZ0EfBsdaar14T7X5FwYbqMROxSYPc+G0eQ8p9Bx+rE55GjMWxOPYTdmMmt8bpyqhf+
ccLtnnhfuuMDdKwl58k81viwdkjlfMW9QYls2jdxqXx5q2tYzPop1xj4ju+pZz3zffOKZ3sY2pcI
XrAdItNzgwXRIhvldYyMU8/acAjcUPfdli0pe+Fod8PM6s0OyErsWCZ8OvQ/096Tvm4lwp3zI67u
gtaRwxji6m0dGYN3YQVbPDMvtg3d5q1KcO1NqNLanMX+FmT+ZAa5UMu9K87xoIFi5z1o7kfgw5lf
WoAg4nbcB1czxG2aIzkJ23Y52zxRQ57O2Dz82Bzxc2XT1wwubYtx8AH2hFjUJ/L7RyO6zxWRHbZx
5d3NsXPRspB+WFn14vD+RiWSs7jAGpIQEdPteOzr/pLFld43Jk5DORROHtjg5D3KdITURxiA8aQw
DHLamQM+MyFx8TWHi+WOH1TczEJxorAtWrVWbSoXrh1Vxmz4SZYdDYkUc7z63mPeTuPVr+uqGrhE
AtiECG9vXm5e8dImBjZImuhCnW26ImfwVwWrmvKahhRouvpBixceBYaSlu4sPdlxEtwJ6kOXCByO
1I0z8cS8F5hAs2cC9TSyxZOPcBm7Vw+L0WdhhRT9Zpq0yqhfyaFkm3YzlFI74ZJgdXyJa/ceg1Yn
0I7fmS9Iyn6c+TrO6UEDNASPIpmrg81s2sgc9B2IZKvwvjrklLbsdbOpjTjSSfXLG+j8TSpp5MjE
aBnVmav8SqM2LBYUt0OVANSrCDYaRwuwlI4QdxiOIg8sOn9hFoLkMAufdb9KtzXp87NHKVFS3Pcv
G7cGYg5OZ6hC4c/9UZx7xAO9I/r02knRT1gx6l2uxaEfbYfv4l9tVj8AuspanrGvIbriJP04kjKC
BXCjWqfkW+rheLPPjRg0tAvIPTKAJFw8nUup3oawrek0XFg3CCfXcAHU6g0Ik/S7lLovQmH+N9t8
vaeRGjmyxcUWU22JT6P7YioLufOSNgZnQPXaxWsLfbw+wwdZHKbjSwUvAQaFhLbtWSmD5yxPZBOf
HFE79DExgTA25njzbwuj3DxVb6tw+YZwENps19GFirWgVbUXiJ5MiCn6yYG3uq7xHIokpqxyVFQs
m0dSkOXmGCmxKhQHegGr1P7cRhBwFd3uAaPWyvJZSZTbtXjZzzwb0vMu6s9PguRGEyGFH+5uN1Z2
NJeM5T+zHAN++0cfJk9fgxkwnKtKLh9aaF2EJNyMvo649htxF4DIPr63EF9lW8MA22MZN7aFOAxf
lgvQWX2AUJdT+8kHPaAxneMDlbws9iXCXOMXudlkMMbyz7MYSRt0Ompn5T7PkksuPiHUGKAPhE6K
beyXTYW0Ly6sg5WcN5FOBbnI8tNBy9WuMgvkcTFhtcSGIdggNLucwCa+Htyj82W7wtZrZ4gokClC
9+2l84ShC2sNPyupMRKwmkgmLIsW1OU/0PoiawMN3DL2sCW/AKzlAZKB9kO79dTaXF2g94ikhX4g
0kkXzszPrW5vPCyDdu1uaLXEjc3aa5JL1YgaNmWPDNrhHt/icmPK9y1tyVPRBKSHFDqu6qlUgySj
IQAmJJxYng392LQ9ayCehPWOcwrjxMo9tbCkmfmkCdZ3Q+bOXRTw02M9kgFtokVjw/d69oxUjwzT
a+ERBqW5Vj2K8iF+UCSzvDc0ILbLWonZMRStcJzXoMD+py0lCwIV4CHv5uO9zTzjC90QqCFN7hLq
RB+1axHeLIS3V4jsmyAvwzg4El7lEYr6maKDleWYkAVM9PpqhdK/vHDVzZFjAZOz6E18GbtZjcIQ
FS9dg1cmUr6fL2Dwe9t3J5beAiyXFhzT5hDrZ19dOs2bb/UY9cDYFhNwXbUbtTpkqB4OYZoFuzN5
1wU+bMiakZ5+pargB5yH5oh8rfEoKvhDcxTncbFpmI86aQBVYg5Cjra5d36PPSLUtZx6s73LjHPL
jc9qPu3jeAqtWQCqx97vKdJiYJ6Hb0ICkJqp+KyLxzrQOqCael7c4uM6VtPyK0qE0lEnr960QETB
h2Duet/XSmbZzlF7mcHZOA3UggL+fZjgmcY020FU/1YQOhflf5ELnA4grqCdj4hJoRpmnoCMDmSG
n55InmSQVRisruztBi48dy3TuluHLC0kY/yIWn+vGYERhT3j2pZRNdmJfU6c0F9BX1p8lXWzJn8t
3uhJ6ApceIVkcKJakNfGBLwz7NeZakkTn7mPuj7gm9XGODm+fEVwHGLG87oL6juUzK5qdjTO4wx9
ZMhYXA07BjRsk8zHSlmxpq/mAAPXDmviTR87Zt1pYeMaa88oOJTqqGCZX944EXSkBFTILvh7LtRV
pO5nUvjMd9yTRZDJZgySvDUF+4UfbOGjr9MhoKxE60U5Lmg0qch5ipcxf2FnB06WpHeZynIBoLXg
DY/EnvA/xkVkPuPRiHsZdwcR0lfnOFZTduicYnXTXzHCuzhk4osjJo/tV7Pl/BuveHjyl6dYZ+ug
wULI4402cAWFdDWG5d4IRMGLRXklN+d/sK1U+dVkFz+t4V0w7NKX0kZdUkSU8jBDvxi54gv0foIv
4TQTkY7G7akA1jIVaUpZu3/hEA//VbswMag5TN/52vp+8YsD3KKxSmFmSqcO+JcaSkmvRsah7W84
ppmw5wIBsia77IdQmGr00Eou8ywnzzRY7+gNQH5f6vAPy+/ODHnaJzcYgpImlqxaWOV/MBvx3165
3gyPoBgXEPtti5kqjDeMVlR6IKms9JlT+LSZv1m7rwRONxzTVBDXeWVjN457vfermpctN2AO6cVO
jCxbd/P2uQICWrh+YTSjTrZU3Bb+FaIODrFMggPiVBB+kFyGHi77+eeXnzWkIZuWjj3sGspb59w5
U0tWz8F4UWSw2EaNCZuTk7tUClc4kXv2IF6nBs+6RxtIrg12m4b5C6Urs1Lh4qHOBltvjRr3LVPf
NrFl30KFCDroSR99tCcGGRlWhH7QuyE4GLbrY7Fkw+bn0WyVp4sNmWgOuDYKd+6iWuI1teuqF29Q
D1GejNedozW0SrV56YRHq/zpmydN6xA/qK6GLrbr0qpW7L+iUvrxMXrmkhzpU7p4AHNbcbAosZHF
urqgzlgeRoSxHHkH5RtnOg9KuvmvUykPPdLmVeej7fM1j9KWvz3L/bz+9IW5ZLmBRu9WZYymagX/
8IaPcF5JRa1Lituzx8ETATmbGDs0GQdecOQpVUKJ8tDZaf4g+K4Ytm8ee2SFBa67XXjufEhw63RN
lJDnjY3tmHwgtYAmwmlG8iKhe1KG/bv61Gtb96eHTwvC/UfJyqlH9Mb/oqAfanW2H2p9JbKJ/bkV
UC1zvMZes0TTNPHivXzChyfUjd0IXZWxYtTpIMQ9bgyuGGXZjZnLtN84BdrXt+EXdOBsBkVfwZ0t
kDeBSrxhz/9uo+r0tVv9VMuHKBh+f2UHCiMxoGDboB6BcJPspaAjM6WUe9/xIBT6RRST+VL6h5yt
XmV4Y/dgU5xXYw9Y48upRxYQf1VYFIPsTbAxV871W+hkF3HNcLKfOsp7zy9OgpePAPp9TxIBkATa
072zpzP3eAE2c60Eth4AqGnA2PvN0rg9sVzSwn5jx4PcA3jPqDsCJ1m6BZnzMuOBwxP4Q9arvxmR
Yns2FqaqSrFU/QXdsgD9+QUwQaTH5EJNeJn8gReP769v/BMwklj/CS0qS3cMrUTg7RCAAxoLkh2x
sLVnw6VR71MfIQgpdnPUyAF9Sb/zlHSwmU/BLZ0FNse/itJdO6aA+vOhjNWoKAbBf1EgM8VJeNLY
aDo4sUV1qIZg5PNHfM2kqXYhj/Rf9HKEBjkWIj/cdZ9XLfWG2F6ErEEfb8bVFnxwY8AqwolwN5Fs
4dxfDG/eZvr7BaUWuNvJtzI88srvIf0kWo1KwicjkcE0vM1vMTdCvLAsSY0c2jUC2eNODNShnO8P
uZEUpHJrh9JCmW8iuzEvpMR2yi9fvCOmKOGsSAjkBibVey4hhVmbT01wkmWkD7Y4mNZaMq/F41mG
H/lFPEtXJkK/uzUGAM1FVeNtFMMGc9Pw/iIkC8DukUSKRmjDhnEeZiUfyTSk8d7Xkl3Nvs/ve4D2
BFEztrFo6yUZQ46PEhJBJPvGhfukvliwlr5tMiH/avNWvLWnpV2iHhrfYD2B45LklvKeT98wbTHV
Wqj4VZxKb9kfVPLjOWk0t2JTfL5yNIraS/e7T811BVmlmprfyqOh3M8fKnu5nKwnjk9JW9i1Ck8S
HZGDRz78mRQ1Z5QUYLjZr6acZdv+yjr0J+0S8SNGIS2Dyn+Omz+z2OfDf7ECuMk+Y4FVCyKwEM4c
VjW9mkn98HSr8iTtlHjNdTmb5DKJCTpa3u2TjPQAcyOPtKAjPk9P+hJAe571cXHQpHaYYq713P2f
7D0ZK5ssB11a7woC8zkuz/76Wp61kO0yyh4xymcQfOpbXSpG0opbnFfN6nwFISP1ZFWqpas5t9GN
6CDldDitgPfqOG3/3KrdLJ1NURjUPohc/xFfgdUvf678avHpBdseKVcQKcdoeLo1Y8ZppgcX5NuA
RjDraEBIkqXbQkSgu1iAiKlDfTYarmFsIOu12lsWH9aomEquCSeMFey5Z6YosYvIb5CugKcd81CP
Xq1uwwP0QX7byiCLxglgcHjNUp/krylukkzPtoPLQwHEXSNkKCM3ShQ6qhRn6YvoiHkvY6yBbFoV
Zd8ldBTU+8mAX2G1n95iecc1aNuQNpe+r49La9V7egBbfQT2CndClM9E9iq/1xDsQtItqOM9Kexm
pCGEzYPp6Nn0y6aaoL4WDMG5PfxzWxCztzJ45jDQ39nRv627aFAcenc0kZ/bsGG3LQ5Xu+fWfvpC
Lii7I2YvHFLm0PDXboozx98DkF814vvGQM4bTf3VjD8jNNVnbcXSZldC1ciKH6FV9ZzXd8VoJcSR
oigJbMZ9AW5t3HUoXxfMMh0CnUwn2ivQB9Qi+4uiJJVXG7OZ1FTlxlxDR9lV+Tao9gX4+h+5l5q5
KSnFGK7KyfOWgMeANHUwKUNlKtRxejo4SAX2o+tpL8ITOUJJxE877ZdgMBDhZiKa4FLDNoCZtzm6
3y5GKVMl75d2uhZ7DuQ8c/ThKNqE8qZkuKT+d1K3YNGuSP30/tTBxooAxHjWYRqA7ZQT/VcxK4Ye
ghW8Go27DqYiWfAvNhpV6TmtcCgjcXsFx7oYeZL0IRkfgTt+9L6w1Rz0oz4ZyIMtsTyQlZ/H06pF
/zDQml9ki2AjmZhWYD4hJBJmDHywCS/6WpGmTvKDeCOWbPdHpsxo67gLDihZ1b3fFOMzjWV/hGYU
uY3Gtu7Qs3euqET2x8SmRuhYYUtZu3myLATnYZJ/zTkRp6ex84xzRz9uk7OyQVGM27z2Lq7+Wy87
ppVD0+XypUR/JSsEz+bQM65E+jrpOQAGJ3bkCc4tRL2sSReb2wBzsv4YVAgLn6GOrJdzhG77SZRK
jjYVYBLof/0xG/QEASljBKwYPBv74Vzp8LqtQYbvZwo6yZDwvkq3KyoqHqNd68C3a1hCW9CSUiXt
B9QNf/bHx1P5O8x1ljSvsX9vBbjTxiqR0IsqHTPfVW6tZK/IJ2P5EObCX42l4azyeCQxzUwsVxX+
iUxlLwSMolGeRwOKp3w0Sx4ZK/WiQPfOYcsENTX2XFxEQ5kdKaxhLH0hCMEmDe5Svx+ai+pJOXsh
k+RsTXcz32okfLK3WJLkYPnOW3Wmj7MvQgH52q/8buz7a7xupVzpOKpJuAgha3hthfKIEW5j4IUM
A3M5BJvICI6Ztrk6L924ausU0yVpq1CnYZTRNaTzVCt3zyDadMTgaouWlBQCERdTKty3cCbg4UIL
R3c/dtmwju+2/BFYfSDTAfZpefMB7cSsP68CJwCK+oWfRkdlqdCTHiQyvJx72tYfedYlKxL7XCmK
fiIUzgNMLhY08nnVGO+T3zRcf6DPncg61XaHobNxHwSDy00sxS5AIIf4Q4D0hkyF8Ffh8qsMCJDa
4yTl5D4Q2BnKIITeAwqkG8SD9xg/Oo/5FAMfx+DNhQoXwTSYYDhl136rJNkplomnmP9P1Brx06Mj
mbjnp2tryol2c+qI4noLebYscTn1M7GYtLYCUnViTHoJpHGwt+GqIEvPNX4jnmBtBmRhYht6vj+5
Zv7SIzNfG43QouLxBmEAVOCE+QVHaQx0nkH0IolwGPEsUcQr7IAGZvHWyRGuekZAiklSH6Xcc5cq
Q/tQWbc7yAjBc7ndZ+eJ/VoM5AFr/piwgyT/MZNtGJqoDhYfHtlVy/fubPl46mf6c0LU/filSvk0
LL91io8IApmr7NymyP7qkmj98MJ6+NaT3bVL8XsXwcYLqNKmm+4O+8Xj1s3is+HfyTmiFPtPGihk
8JfTZxyqQJls416DImEAetmSvIKjP/7lmUnL67wiEVFLwlavuCpFO3xkovG4vcR3K1MpdN1jTvnP
ecoDl753xnAyCnn2MWFf1lYlACuG++rmHEb6ruh31m2vCLkr+xDUCYPc3e5oQRYD5LL1ki6SD2Uy
9vavtxibdo08XlZjuErcBbHAX7qViWCyeIurmuF65BuzN0ZMBdubcD6hTzX78jSDHOAQpBlpvAp1
7kB1bzYHQWKPCE5CJJ+lqP5tGx7ObTQMrR+J1YwDnScJi2zuLtjvO15ZnLo2dChLfQtQLQpcAmn0
T7y32obX2tgaJZGSGYJ7/y+ev/23Omi6pcBZA29N0x2x4s2N4CWG+pdddKEBFC/DgF/YTPCzL3vK
nzQbdUT6wAzc896Ke2wi7xvk2aNIeT2+ao6P2byAfODsEqvwZJWWl7wgvumWaSmqALlBwTBBMWKK
GRHiaTlm4bYiHMbBTxHiGZplEcV0OU83ugaMFnntb3SS+wkSQg2v/EnwbOKUX4L66Yo8LoHEYCnY
yZv3qCoEeSXdr5UDr49LjuIQEogbIvr4LT2X2uvV+2iuj4laq22bJM3hPO8ds0ycEyj3C8lZ6cSk
WGWE7XRJ/Ke3Kr+dUzyp0fVAWrin4c3Ak8+/hldoSDl8R7JzbjoTn/XyrmBzWf56YOQO5fxNJJmx
xZUCgkCnjV/ftX6ss0M0l3y//2dCSoDHeFIVe3/ms5leR1desFnDpyJxKkmIJVlL4i0hOFs+yC+5
tOe2smbUBfWJkVLC1UjRgy/a44oZIYRldRphjFS6TK6aIZhffY8P74+c7mNyu0YNzWCvYf7r9UN0
heDzBFD+qCJQ3FHtEUqbUN9/ZRbc6ZQzjie2dN0Hev084eZ20vMzdS1y+nOpfkNmRLNhfzGNJng9
wBjtCj45N3R+pgeqbXkqanJLLen2qETLWVOHzJu+dPOcgz0vA59qfjnlzsdspoit4meARY1GH4G6
7NEDnnd1W5OUacrZAYvvWGM8VI9b7Isn33scj74BrugEkwriUnPgwOFqKYGpFdQ5M+G7C1EMbi4e
RiSdRAtPEzYj+6KqiU2Euw7bpAba2gePadmcET7ozIT0z7JMFcmcY6MkQB+K7LgF+t2fWqb9VAoy
j82mvsE3e7uMG9mmSFjsSlUK1nLZPAyFJUVgGJnynS+zLe/YLr9rE1HtsqN6+F+zAfdbYQKQNIZ6
dp6l/vuLrDZqst3w6c/P7bN05FYdlNwNJHjTX8Mc/iKL8Imd+zylKRMsdP9qG5WPd5EPtRkOwPbj
sBTDtuoh8nQqxx3tiDm+bb7wy4IyqitDBVeqoOEX70wDgD5hY00SBAFqA4QT5fINjLnFk6koH+c4
sSDRROZYlWlrsbiCLb6HzFYqowGo14vQPtODGVsLcn2VlmyQSFTXjRMTfH3k5fVFFW+G+LJiQYLB
dae63lvM2r28cGGd2wy6Pl5AEyxmD/H61jh98k46hEUnkpH/b/1M22vZ8cuhlN3OTFyxUaMZNfc1
ZEZDQXuKlmiau0vIRrnUZNFWLis/+tzMuYKxleWg2XD/6u0N/6J7LOLMhSZLgGNjgRuc9CcLyNyB
TiTKQULXdzTV/iLt8EXCkl0/jZx/xlZaO/pLeiBPVP02LPIBSS/t8/V6bZuKiXBnaGJxP7pf6riR
eKSuqUF+gve61oVwbEab6Xr5dXB4V/8OR4/UMHwGk2sjUjPzuQ106iDnex7QL1wECAG+mT32PXPP
GCJZk8lOZhqNu7ujH3uM6mQKV+gqxLu35L6VUeacDGzB+gYeGIo5z6ycLAVrq+Vd8lpk0/zmkVCo
rsg7Jdx8v9pFcz5mTFe4JFCnS0i2haV+bRgVoP8BfHjtFf/fHnTrt54AVopF+YB6pBIvjiV8uMuy
3aNmbXkkwuHMUT3Q0p555pIrD1gq0d1uIfi2XmDNpFzswfMwzU0yhiTQHK+U4dQFmqd/lL6JOG3Z
a/Vn7Hl9BOyRerNv2umQNBteC/myM2koYqY4p76M8L75KtA0xavdYvCyWHGtT58UHyYVUqZi7tEv
bhuGIeA4i3Fp12jCSF7sLug+1s9js36qwbMRrvk5SprQNef1qxzbZkMNyp3MtbzTUSMTYmVv5NZW
Nio3oYYlC6Yv0tBlRFQV13ZVmG0T0lSc1JswmQaPrMYwhOGw9eeBmJr7m564H7Mw7KYiCnvnyo5q
O0exBQ708AoHxLNVHadiOAhBJoM+Db3yn9203JEFTnC48uzr2nzCX5WwY23nMeDyuIiM2QnycFxK
jcG79qSRabteLLzUnYRFXV53Lj+hWtJ8h/n9M0o8cjf6mbzJ+gyhvSKeaxnaVhQxWWy71/vzCBbO
hFq/8vyvE9+WGOns3pJmyYwaJMXpoetBDegW7KoOYXkHz8z2q9seWpV4R1Vns/KN5263Keu/Da7B
9jwfu0dwyix7QAulMFonseh7NyxZsjQGIaHKNBKIoEyg3yJWkmflJHSDPD5/hRiPHKljP1fWnYp6
h4iRp5Rq3wxWbnO7+FWfurzhHpRJkpuFNeQk7Kbd61vbjCgORdXEh+yKLPH4Ml81GPDPz2j5jhIP
hqlgj1XHeuKibhkdoBjZB2UyIdR1WKkc9BEwm71btpnhvTaCyURTGlCg0aQHx/bBvAsSLkGxXKnC
SnXwc+s0mNxWvKKeHhgAodGcxB3wIibyTiZqbswmpwDbWapQXgWN7oApq7dmxxGYp2aHDKpPmd0o
S7FL96+qgEAhEN/IDnPp1JB+TNj/A0DzhC2MDG18XmmX+zHobjbVnVUY3p45j+aRnGRx1c/CR8Z6
bpbzdcoqjlcsPIMszizsXnlQiYcXFHqrv/rTL2fIw+Y2osWFlv42mFWu4rYTZSD5UiDvbnRH3yWE
imRDgsKdtkXgshSNVu0W7wtYObIoT83ssM/WjVEZFVuMSPtu3bZAMyCILtOoQF2aboJb8zYetJAN
mjjJd5cm9oSvkat2/b1ikdmpqb9VDNqxroYZE7HCyHoj8OEze5tUxGugUuUgNLVv37iiDWddjpVP
pubLLLFNANOICu5twvRji6f1R6c+BIwahfNNeMHaGjAUzLvGuRvgWfP8XZVOLQnMet7t1y4BYZ/o
lmpe8xPTnjP8RvNj3Q5t3/3UUNFCR4ZLLwgSzN7hI78dw191xseerGFn6UwvfbH2ZVW2JTVOm9g6
WubvqRV6J2VHK71fKmnCQ5F6dzz6KJDz8VeN0/530DmKThDaqTxuIPLoVEhhVeas8M0PFFoblKtw
DhkJcus+EejnDGr891IhbQD7C97lbKqz+6RGZEX7sT8rs92aEwisAQRCY374yANF1w78CeKagNlz
LoZ9ueyekGnqWPiReuBErWNIYQHXsCPu09zKypXns72ZexuD/OFImthXU5vyNIu+s4vMsP8sPw1I
VaBc/vh/W0Y+7aoEPcVI3rhef3bVuoF6eFqhjzIXGHvdt3w1+CbCxADobB9D63WGcE+HCKxYLyMI
EcOoquzyAbO5aIFurDUG4EpXZsozKcx61niNbVPZ5idwuJzp38La4p6uDGS1hHtAqRCt7E1Y936M
hpIEflm/h/mEZExgKRGDaI+fgsoN+jEcjb+CqPjdVs+DHoFi5/+TAiEQBhjmkwEvKM1EuNojJ7zO
cYlr2bvxCHFw0cjf/pEBYIMSpWpiAZpdYGETdB/AZpO1ckf02uf3bKfum8AvnZewkuRFsbqHcPH7
Sosm3XM9eMlF+gfG+1UkkLs4G4oJfO0sEG6OFDkHcAFVEGtLw0y5+HF1C8YD66k6TvBd4qdswkxU
GV8zkCaHBICN+zh4CAZX2nF4Ky1mT9KDEbVKCx7BGjWP6K+MOO+6sEJ2oxl6d7d8AmTPdQJAIF8n
ytWMC23IGjViQ1KDLgMZyZq6J++22X/th2JfkIzyWAE8PccJTMuFUq8ouSo30gjympagSZygvgpS
Ze5qTMhNqU3PQjkGiKX65OnTo5LXF+cg3mcojrvSR/9UZjuGJwH88yN2nHACwE2xn9RIqKjxnLpz
/yRYNo7LD0/MNe4WpZG71BmmQL9oMcycxnZT6XrSL2kp9PI40iiSKSwCE5DIkOTA3lC/YWnTZnwi
WYlV0Q5sTEfGMVsn+doaTc/4loWV0NtDYOXt8SdeJSf0qj/VonQhMwqvCgZ8QrqR+4Padrr9KEnn
drFb2QdmARle8NawsSrREj1AP/fgKa7WRd+Ws0WN/mRAS1i5gdt3LBVkLvGPZi963ofyijJEWdlV
+PDsPiMVCpY5go0ha6DtdjTdpEKi+J2nzxQXHpDJq+FJIPvNuRyu8JXwnCAgq59S0AvqTtAcFXmn
w2jMvCvY8UAJxWfAt9bmS5XxNzRFR+xSPKuxczoxq8dKwR/kuPEgv9XDDxEaEOleTWVLlXm2KvQX
BV7ZtKaJ5dcWf7ga4CHihgyrW1nOHuL2yiU44opd1kg+bzmJxKV7BwbTxVq2UqzpetAksUCudIdA
8b0aeP6RvekbR+OdIwd2tvKi902It2cjneniQf+HJy/PPd8waHGDSsS+ZkDTZehWZG9nbXHScY3A
2BfnUZItMzbplR4mtBPDR31pF9JzbycbqVBQrHq7O3H+mmviU+OMe1A3Ut5CqMWyEDZuRl8vJggE
r9fkDYFSvpq6/cxKSFqDJT0ijrB8Vtw5cUisL4pt73Zg/Xyh8bhiDYSEVbUHfEhHezXVK8RiPTsM
UCZN7bwiFNZfQxp4pV1NXQUFO1mtKO7bxd7CRk80nwCEzo4aIrZ5AAtehI/vvnT8obiXWyZ1Tsx3
sTQJSPwwa09TEA5vgY4z3pYLoA5vOL4+Rk3Rz646kp3zLQZoFG6C9QChAmA/MpsospmHrFUbh8sN
9sOFuUvLmV7xCB4GhunxrLEh+HiNx/FriaF6W+Y3HBhzS6HOcCsXm2C99ReLY8JiSw6qpp5V6kQF
kWdk67BYVfJ/HUT3VFFnZDv9NtKYqHjN34D+lo/dnDkCx9VLmEEJFxzdHRn8mCIltFG19OuPmZf5
McplmMdFuQ7Mk6xWB1Nv1N48XR7JEIKd31xx5lix7vwk6gTyMbbxrIbaZQjPCaTxGr2sG/h7frkk
IWSAnk3HSKV7HFJAo+Hjr8iAtAzKGUMjJXTaOgw4kTsSE4Sjf1Wl/9/VjuAhTnZ2HVMkf0xCnM/V
Qg5FDuaYe2jUBkay0S+wYM/AFNTs0iTH1UJp9Wg1Lyz34Wp4kmIYkUGterLR6rYmL+lWLQfEuAdo
SDnAzeZvyUbzCMrSflQu3pD77WcLMErvLwqcvwKmJt/jhnW49qYDmT9V87fi8QcBaTsfvKpkl0n6
YCG6YPMA+3j4jDeAeBPFhc7RyVThqh4WmunANXVj3KuUNu5xd93/HKiRDCvuvXekVWHWe58Cd0sA
+EhNkT8JbCsA8ELMSp+Wo42MnBtPD1502LxsQlzhKg7IprOWjtn48gb04oBwhaCrWgdbQ92Cp7L4
D6z2meKbil7SlO+Wu6pMrGtE7VDnl95HTpOzQe4EnxhjepCsbfDZz+EtFsLfGT5CL5T30caQ7xUd
NWTryJUKKJ0QG54zLwQe410oIkq8kxQfGUBAyyB4s2h52kU7XEoNsaV3VXtN7uZ374X+gwGEmo7J
9CbFDMnLPwNdkVG80w8dhtM+jsUPJkt8x2pgJ7FtL+qsLJEBEgjVvx6n7OYfH/P/ICOWK4eHSPdp
uF75IX0KpNkwiX8fqd4GpfVtZzfkYG+r82QorfjRanJiVD1cUJ2He+FaQsnj+oGwCj2tVDIjNULi
E9cndUiYNogL0EJqyxJHvKkDjbH4HGeadiMNwC9UUZCOj4vnXTshhhe3HKaQdFyRwadA/w7VmVTO
5a7sNeIN0jN+A7TTc1anO7GKR+jxFfoEJ7Qt7uEj8iM0GiWeV2z7lBcKYN1qUtA5AY2ixSd1c/ia
fkghtA450JOmzyRhMt6vHOAWRXUWdPWmQRIl91OcpxlXHLD0byfNTYTqHuTU1WXdJGeMoEvdK8x4
RowLn5GoND7RzEBB5EWjmfEq3wZihdSvK7dqZicIWPQktRc7jHiDECfkd667awPLxZAWefF8xgfV
7YC1CN7fYPpCNbO4gWz8HTLDKAZLqdrZTcKpRmzsN5BIVVuQrbo+gAoYul63Tz0S/W2XhpNutd2j
RdRlrVSpu9CObMMdNlJWzCQlkRGCGvWfjoFA+RsAgIr3V/f9qukqRMA6g6rSJZrpqk0URZAv8P7o
A7SvrDtT1wTHaUykKPmFGRewQnTcpQJ0fLeOjTb2ebItKmXd5rYkIO8HNQCJKzBwX5tcKs3KmkOM
pRjzJf7tO5W7fg3WK6dGl85Y8W/N0WdakZQ4WJLT8t1z+3X65UCxuW2ktjoepB21o7iuMWIk300S
UKZBbZaiauBoSYBlUFYNAWhsZtm0FwfB9EvYe+wvm5cW7bJ0B9mgUC8N0HMHsLvcix1Jr2TgZlbf
rxfpE+39fHhKp6kEvz1buGpUzfQblqoes1JsNBD2ZVD0XQgILUb99+TZGXA/z9uS7cWqUzkRIat7
iN9XPtQKaxVzwSJcWAMe3QkgyS1KQlPHJSeCFgdf6j4E1qSuz3YTQ4Tt97zF571kMeSRvDzTWw6F
1vsp6vW7GBV8KicBQnBgMRXtKp47gHANKlFAxbrAX73NEtjdOaFM5iTnBnqUqW4+vCz9ilzgF6ea
6cGiAWzX1ga0G2sarvDmUm/oAEWXDJfWxi8EwJv2qXURg3+Jxyg7L6JmzdT/+9lQ9+rDrgoteDoM
m+0hTmQuXCQ9Ggls6RAErv2fnCf62QWAkznj+/wIsi4r9NJ2dpFA+5ZkjJxdfEzrySwUh5eiADcz
OqsTlF0/tym3ykhU0LW9hAHu4Pt5r3NbvqbfClZcYSLyPW20nIirxMWXfJL6qhWg/4+iAYy72+53
pYisgK49rsp4yNLSoeXUMhhrJdMdteMUSNsrYIYymKA59GJ9IsC3pIhoTonwliY15RrTQRBmm09y
X7uKthdfgVilEPb9FEy24iUtqll2Xhe33oqeQa6tixiwUi3vpL8HaiR9yOdFFnitbAy6g5n7iokU
yzPyUACR1uHoCNuKhnUtx2gnzvNxsXMRsLnf3C7SbJObExrLJvCX+u05qetIkajazPWtYi/4v2gl
a1h4GCukdB3bYk2pK1AQ4yGIpLpon0pv3rjn7wqMYlkcjoiRNse5y/sbihdV6CQ/wCDAPKhyyYxC
ZiNE4mR1wHVsMIcaGkMGyU5su5PyAcFmSlAxfKpr92CGeYIevCSij6zK56ATpBJFhINWYwSDfP5z
meBt3z7Fdmghe7iXxWuFPRau/tbxiDcfpSoumuk5yFITCYrQGniTAA9qSF5PWhjWs7eQvxxKOQKI
8UylHzkvIEcARDnnRUqk7AVwm40iyPdvTovrUzYcaP/akGAHHE6wteXqrTcyLKBLgHTErlITqR71
0EqO5AhNQhqWD5Nrmh+IscB0FgWvIRrvfXSolbrUtKEXdR6dGzUmM+lb29t3T6k6Ig9+Byk/JDps
RZv4jTzA86XD34z+nYA1V4KbQaa8cZzXKoLFgo8RGLCdoyxZ/vLwxJs6fEOenHbQBEABhWovwLU9
wUvm0RIWM24MKk9eo7h2RBEMkvr1PkVMEC/ziFs3ddBLeW44FV/WThZwyl91ytkN3ZpOYzh1wxj6
M20Pms++6zmz863l3uKMOdc2h+gx1y1frUrx0R6PR50jy61y4bZWbncOifQ0XNcQgVooeRI5kwNn
6Iihf9i+zLuFli+Oy6aFyaJax5RmuJNkGaDtChzY5MLVy2pd+MiZeKGGlZP8YjEflyBMTLmB1sfO
urV7Z4zTS/KSBPD9/S1OaivYQfeZ1tFJICVpLIpdV4Z9gH9lG8yvW+dG9diSihXAwqao7F6jCRLh
nI7QyhotZhYSHQ++0D3upwHljgL+7SW6wBzAd2X1BFTYaR0LH1i0tGgDi2IpWE1WGPombR+FAStv
lLuoNMeBzexgPDS9fH8hoohP59bm1+6f8l8HpgeDlw6NaAGeSOrfxEvSGxP9iUuepVDvYvzPIpWZ
unqzi/VKzH8cj/n4XC7HZZ5oasdlUv+pgG2NvGFw7isQjr8gm8JawI216g35geWLbCfhBRHs8/Wp
/1ygvDVo0ItXiqhBIlxxQ8OYVhuOysvOKOXozshEkk3HMWO8ydP8L06J1rNipWRag4ZOSWX8wx0Z
zzg8/4MrO2AhksUN77Oo3MfctOUiKeTV79RHhx9dSbP5lfciEwoq3WquvIczN2vgm9n9TTDVIs2a
0HtUvvfceVo4JWGSLXnmRwjZAGDeT7+rCsNlz724FT23R3OzZnHEZP19QRPbVYLx2Y8yQRrckuPE
yuz2M9pwzTESbxEOVHqs0I9qpVGnUPkcPMz3rtGL4Ytn9h2Yy0UgBY5F8PcS5ucbQYjR3ur8l4AO
Ej/a18h3dNKvrsrQBIa7nmCryoXfV+G9gwaCrYVLaZRPKbof1+XxxunEbDi2/SI+xxjVYD2DiEN0
gVrckTEOklJukwLiG56uqX2UxcheihUwEis0bmIF2N3zxATwxsQnlt1Ca6fQvvFE1tAKphxn7L3/
adq88D9HuuIuXqWJIkTDSU+8Q999W7xom+PosdXiU7WyOyS5h25BIB4lXomIgIZBkgANQWAwQvmV
2EiM3DDId1nZcTzHcBOT6EA/QyqZq6TLz7fox/EaI+/Rq6FYomVApXqLpgUkgbE+0M6BpEkhHGQd
U6nmzsYQT3rSI7HJDeMsxvey6DYwiHDlbvuz7rwQUzu/FZS1cqFB9gpbypcKalFo4M8ps6uWX8II
RuVq3gfDfnCMoP+BOFotv3Ran/rlphqKUILThqI12xMfsxCgjxez6KASy71L+43U4fAJ6nRH48WP
71Tjx6+zf5+sB7Lbhmm5eb2eMxTU89YCJbp+/eow9SPTcpj8p7ajxfBLiaKvR4WkUkloTYvYEuTJ
WEF+0TuKeeXNGhaKB2Ip6FbXI+H16s9ZdN3D7QabaHwSm8B8xn6sexBWMengqs1EMwlQ+SwOQnWq
abBs3K7grkYenbrLD6tNc1z7hRdNgydf9Dx+N3Mnt1Bs6LmtGcErKjpwt8YcpUt1DxOsM+62sHcd
dIJOTvN2P/ezZ9ZZqnA2N5up4uxK2gj/Dljvv/umII4mIwwkS7fzjgZ8RIOLinr9ArAR1mgBJ6IB
W6+Y1i1cOFRhRIWfeIRf3VBV7Oc80YS0T7lcdIhe/RYyGlvp5o8elkVfusY5qrWXFwagKujZVYw/
aJxzCv4BSmkX2S811Oyq35nEU6FTplb0wBkFyIshMNmg+mE9JLYIW+uZ1xgloQv9A4HRonIUKcT/
Quonft2lXadW9U+d4nYEvt1LIP5MdfKd81/smEr8SF8hw0Esv7QhCmtmh/W+7nqd+DCjaCTZM4jj
/k0WD/0k0r2+wMiNfAR9Ah7QiREX2qaRxXcq3brd2vTN9fAEiOAwPPq0u7Lfi22wRbvTuLJIDeSb
/wtZBcHmYlnGlvOus8yS4W5/3QtHL3OLjRayqA5QKOUX+oOKTIQoL4/kaSArue8BaFvpqN56wqqh
kVfaf0IdykMwZz9+eXK7Zu679m0F8REJaCbkbGLWNnxxeyIuU+TIFCamgp2cQtUNpz+OrkykRAJU
xTDNgK+odJOKrnnb/P1UOW9yaNLSvgppYc+KLDa9PcxPwSSrZgd92BleV+qmrohnFyo++1A3nQev
TwFGBv1CeB9M/P42uB4QBDqnfVH2uE528NqAMU41ZQDIsxWvzJPsNDpSuJLfqOPSMd5fZqT3gtad
6BW6Eu2QgXAChkQ3/mILaQ2i4NRpHwq6IiZ/mCURLvYlWs4TWs5+wgEwyVlpm7biifa2cSsk05+q
VdelOVm3k5ORqGRy/fJS/LmJOqrH0cNZgGhti6EjBX8BJUOv1umw+7fJIUszlZfACFB/cqbUgIFQ
kuj79qUhJjh7zRd50256TIZlEYW9DJdtAZEorwx+MnvAzRYWunJt/+5w8glCX2+pIcU6JJgSnAAI
2TGF3m62DdE5KhBajl8UUIFG6wM1+Goc+gqzgbrpKCa+Cg2kKm3sp2kiz5fCROiw+hQaAnuztC5Z
u5S/bDdDdbWxnTkqiKsYaw/9cg6nqvE/ukcA3Tl/6EBAXsxbOhHefNSmqbP2S9bXHfNw6euVYuT9
7wsKEpzJZqBI63x19p0BLqChV/SQ3sJ6ag5XzDBLMP/WMGEWqKh8WMiEbD0V9D5rluutl/8VeXHK
zhaIB4Hc+XPY0sPUcNUqn527q4u8SGONhRuNpluld1HogbnYmN4usqfV4bQS9RONkhQb1JGLDmoT
bfHOMnpzy1nW4xJ95pLZm/UCYrRbs9hnnNzlX6t1kKIXmkUUCmv6b53pNyszBsfVMV4VeYvjwJYr
jYf0ze+NIXWmiz7JhieH8cjnK9VkvtXjcohRXs48bQAD4SwVjlOlG87GkI/BiQb6T1Aef+OUfTr/
jpEKy6ghMRX9g25z61DTeWJ4OggvvZvEwsyZ0gAi34BLoozBCi+biKJlHdJYmfTzDFnX0SvRQli3
tgPU65rc8Igs8SMR/DnBtDRERcj1vaKK8GXYQXKQrPs1ZpWWuFlFtD50yglggcIvyb6ji2SjbIfD
GobCnZmgIYF4QinR0AH/ivn3cN0Misrs1aGkS3CXgdT9QemlJCqwm6lsFqlJSoq7EyJpPhdJRDBT
wT43eD0H1H5OqRprq4M3PtUEjpJYeamuiVZNUkVYQCzCBMWqWxJgL3P29Tq/6Y/JTAN6nKpa4Rc0
K8Hbbzq9THUSrjnVZP1yr78PgnasKNvT6k/yczabV1Gr5fP2T5JT0H1PC+/s8/XpKOPrT/UOf6ef
/c/O2to13gb6Aij6hDrxnRhVUDoXch7nHhfuBjBgTzWPRrDbCVDUQbPTQ1f9bCizXi2CfPSW8rSW
+SpaU+CDDIK70TTEW8jDxIhu+D6VOQxUdIW+KejWt8riPOKIhHLIoYb7bh0i+UnnKXx6tPd8BTnM
SQ7Q24Cs/FkYWzUJXff8D6sZtPJ0m93/kACIC0m+9Z66JD287KanOvHUhINUcXtY7z206DIuTrj5
65TEsbk69N3XaSQfZEyPkGLGj7lMO0FyqJDPPvuotPtJTTAsff9H/E/doUsd6JT7TMSEyuJW6kDN
aUOjrJ+nOiZmnwA6LCQy2l9O2f/A4VMDRcMYV5YOuAFmuB5/PnOGs52KVM2g7zjCHqEsatZcwYYJ
kXkEfKNcSFWKcmuGtazga1lJu2OJ56k9MyC3gsTzlqmbwyFiN+5bnk0RyjLfgDtbhZXlxffTRvbF
nLVHVjBU0Krhi2y5kvIs7exszlKeK9OEb43IvLo7C+Otx2IZevvrpbyAsAhJWxvHTAkCoLNhnfRd
W6OeygSK9vvCyMrGDC2HMTBnxZTdCA0mjD9i5knj8RTfyzdq6dbfWPlB4c2wsjJn1RflHJAqFdDY
qD4GkyWNKKk5Pomrhj7zvxYhHzicrVlL5XDsPpwglQoO95Ci/MY+nG/PDBowRTA+WMvsc6IOVHdQ
4JWeXy5MOz/2ED/BZUqpQAOA8B3XdQDCA9QUTMY4txz0K8DPaOSiBSQJQWEuv7w3gwjlpyRAUy1Z
M64i5dglCMCOKU5kU5TAo0F9sQFt290Rht3up7s802te7rVpo56jY7KQefiZEI61/UXlRlRa0BBG
4sQdQlbyHSaNGmSffgn34YEgli7gjC3PrzvDPrfzDZRULzXV7sEe2mDC1hgPcrloWRMIhvgKxcIJ
iAYeJabJA+mC0izI7O909HC63wDRQJokDpbxDvZz+FusATjxy4Iw5O3PeEOTAYLE0XUi8NoZh3l5
6pngj+YanLA6bb+pLIosNWZ3bepje8rFTQcqgQ/9LDjqBXeekgf9/g5Q0KBD/dbEGxZM+rFlEI4P
gjvFjmeX4WNj3/eRWI8aVglHMsDCt7IJYKYOWpBJBAu2tt22YXW51X3lKlnhZCoQqXgybF9Ujkig
Gnu3zPDIPcmutIzFn4VxbdwLDbi+cgYfyNmkyhfX1lKCf8RkPUJPNpu+dCcHmnstJyi2DevOABgb
u6wiivtgveGoj24posPAyqjQmRcINksVJELRsgYukTXturdboHlIUPvPPRW4U8l4dRZ9CUSKiKjY
BlZraYTUGtq08Hos4GxA83WTuZCswoZPR9sNvNyPEcm66SFsLgknux2k4o0uzpQfHPQmLBgAEJaP
FuqPgAR86ik1aY+0Z+88k0a44z5nCDGilP/L8XVzofW5F1NhzbDFVVQEa8vbONUx9GF5M6mVvwDe
sNWmxDOA9pc1438hB5d5YZLzJqMTLIQozDY4D9W5Miv+5jZ53f/xA/WBD9TjvNYizKGojoyOIjFg
yHgweHGt67cDwafSO4MltvKzFLQXnP3qsr3Tkw8+jVNSZLDhJoFpTIJOmx9DcUDRPLJjUXk7HNnx
HgOXYFaRMZZmdm2tRjELrwWipZcVdymlfuzLZbS+2qPNgXzQueBU+FNBEq42weHZbLv5b/OJXU3o
0Ru5L/FGNs767Od13l/ocjEIXkAQiPqz3FAxeb0XY2VfgWa3LFT2Co/CZd9SNZYAoqd6YJHy6xuE
K2N0qbkAGhQ1emPDpYcen+zAdPxH+uE6saCd+cEFdc7Y1axQ7W/No+8pDvbQc+c1lViURlbWHBMp
SP1SKxBK7Jve1M4fAZhQaHuKoB6nw5oy98D3kA4hCPGKEDptAznWkR+ZH1KO18voQq9zNrwagh6y
ePFnB2qmtxSvZxJ1Py+UNKaN+i0p72UmZu3ppqlCkX45PI2UkzacLr5Xh/qnw/cdm+M7G+FkqZIW
KZ09kNRwhwz08ETkf+SycHg0H91tnBqCfUXBQBiJYNLye1t8/ncXDUO2zsB3MLknRy9PthzfRyhY
ruomaUFOPkVrNHwlGiZeefzggWafr3WUciCT4SvMhxPA/MFTV2cC6yx4OphA5Ja9oLhPpuJeTZL/
IWqiKtn92Bt55A/S5qi0Ll/Q17knutOkTRhVbY0m9WThmaZhIlGrJvHVuE+yMl2Ln+yw0vHgVZ/T
7QK1JkB8GMAx/p0pExzZ1PL2l5lLaffc/f2gwTn0hd2mwhOAqcUY7/zFv0KiLKb6dA12/i0OgM3L
5JFRKx2o76z7aRzQFlUhABIyO8ht0Na4QOmI1qINQOzHfZtjsbxTBmp6xtmM6n8JPoe1hdJPYNKP
/JNkV0rAgFGnCCHmV2L5tsgYW4XgcHmmhApALS/JgzzWlUQE0o6yMLJ5t3yV0uB1cKN5/HeMhNtY
AudYriJuIEZl9HUjFg1E6dqkVAi5vPg9CTijmZydb6mChwZnGSksBURlp68CYDkIcs3xNnu/tYn9
AcX4OKtILvgM1GmKru6YNX+TyM/e6t4LF97wUL6WBvO7ILI5MopEFYGloehW8ZjP2I1OcRb6JHzP
SLQl+qGB+FOIhIGjd9Mr8bExZY113bMurxWAj3gM/OeegakDLwP0EMIT3rl8VCaKmZEV6+4UNat3
m8SgTrajOfRn36S/RBrvCc+uXrZUQxt9q2pzU30nSO0SbhsoyAfZLEyMVRtzwZegRpPFEtPqrSwk
MB+TXUVsw01iMnYSDU+3B5LCSeEc5X14I+JonJ10m+WcAe23N6pQ41+TRGMArxZOpRCpWB/RXwtr
DZDtO70tVJDPAsnbdLPUGHqyOQ8z9Bx0xlDF3XmZQNFsdtBm81iWSHAe2tDxdcekpE7+tTqk01fd
QRMI1/fsqUM3E9MgkM1KHzjhsxHKPqCSLyMW/qV6VmhTP90EqsfhKC+zmIeRdEK+EwPx3f6XKR8r
i7Qsm4DB9vwES3Qx/MHHUAltUZYuiUqzxzznWD/yCF5Ri3UWzNvMfh4zw8MOkL0twcgzpjqz8VKz
zUVU4/33O5DifZpMXnW2zk5swubtHc/lD9Edz2OaVsuRABw18LD9sQPqaN+J6QGO1XiL+i/ZyRSd
iXVt0UB0J95eGtyq8fuceVMUsGIhcSm+StFO07JWa0ZqbgrmrWL1SDvQBiH9E89AMfikWCPK4t0F
jzeVNIwnHeISGe5bm/pZDZNui0F/4E2c4gnczKgZKImBbYiAEBPDdh68rSFocg4scqiJgS1fnf+O
xjQPOuSRv+/dDvyinrm0RI14L5q+a3vAaUktaF3pyQUk1MOPfIYdtHgB0TUDd2RSmL4hrZs+QmEf
Q4+gTbzMwl1WYtceS6u2mJr9QTf5ghORpGbwP+V9sJpZV3zn7SEqwlrzy4e8nUz33REQecgprT/S
+OJf7SEHSZXIQI0bUDP+qshTmyrVk1Hn7GlKsrv8qr/vESI2ECvSLPEBsK3ZGKj7KDqmdIetS6qv
5gvYn0qH/PDeg2p/TMlYKoZOKPRlJ1ZQmLAj99gMXYhpAJfaLKl+FOj62C3XleOJaPNxH3Oq2Vyd
y/RomFWthzEfdeMDQ/6LFDatMIqsPNITSr4oZ/mSo3fJabB8vnwOAzbj0N9fVvURqjh3cnt8NS+s
1nFSTwbXS8ugdq8fyazzGGWrqyRAo1krF6f2XQgRbu45cfVdBQD3ZEdEOWgTCc/yBQAMqLc4wDx5
z9zYRGZrPC6sgG4LYm1g2G9DD4rZxK2K22t+eWyR2JZO11BoEQldgaZmU2ORp7rgp4it3PfSaSgI
p9hQcfSl7qCvmwnnkqjZnQL4fS2WWLAEYRjZfzgmWMOASs7XDRwhTxHPHd1cic6t5lD89sYms+p7
JLE+j4R2bur2taVL1R09VRdnOinItyMEn6qunS88CMYV3zqvUdph9YN2QuIOL1Ms3G7LIB4jxW7B
maytu18juqCnOeeCvxKw4dnRqcSPSkiPythDwVDTjKB4X+Ce+XqpNkZFbWmOBNAXw9vFcyOxTLZ9
zZWJVDT4AQfQ7xQjGKQ85YH6YWy+2WraHb+UCbtOA/Hmu6hNnMdYIVJ9vqrzBzMrIwrsxton+ykl
js7jzG5gW8ZLlulkru2WSr0Nd1OyDnd/9oswgcW5eXKU1ivDaZLYxG+umYSf8vZfda9qA5VpPgib
uDSFayYAVU2A2DIXN9SvpVOicDBmpgdpqMpi4SflZWnPC4z52Is4gpW68FUFveOg/xPSvMEgbhWg
xiIDKNl+hRX5Oq8/hpueV7Jm9PLPcl2+K5leUvVk6kA7M71z6biwTfyonF5vrk7JzVxCSriczWJR
fnSDUqzBEm1u8C4ducupY9dMTZMq9wtst9W/rrXYCplqKTKsbpZ7t0sNzslN8o/PLrs3ZRlHl3dr
u6njSYTppPjZXAhAXvAG7D45h4HmfLSiW63I+a6pa5vPZNM0v9pceGaRO60muaAK0ZwCItPvOBJg
zqK+SGLKRyR/dPY6V0ao6oIrcNYHLTMWZIukCBescXkF0VpC1SC2ryjwy5cRJyWJ5eToErtkGUKX
zgmnaJnd7Jeh+R+rxrY9A8t/HY0etxve4c9n4C27NmvxdnpBCKwl2ZkrDk8PXIX51g+l8EFyCAwM
YV0SarE59i3mvRiNZ/yYVVFA7ws0kYzWFb8QLdUBOPk0WBTnTsRWgnDE0fV5TdHOeHBNxvHmaUYo
9P/IYRUdpPA4oCKBg+CVZoH0SFyw5ecBotPMyKWC1WDqA75wF+8g55KyBkKbfxT6V3zQuaQmuRI1
XBsuNpDpX9380ZFjE7xHQmkqPXwG6sD1fLv1NTBSZwp3YHZjN6LlNfmvdrJHwUQZ56XU9tI+SLFC
AO52eEyES23HTMqALEfXGllRDjTx+8FBjPoQ9BibRKd2MuEh6O5HQy5n/TKVDuzrRnJetyQxhrYi
UUyTGZUz6tvno8zFgPnlV4M0n6XHwazBKj43tZzEN8XyhXwHv0GfSifRqH1+oJfFmz3LmSwMcrAr
fPoHjemEO3wJ3X9dsxY4CYm3eU4xPkfj8jpIlkuMKKWGL0PH5Q1wtG1WZO61FXWOB3wKWxTi6Gr+
Ux+dnqGvCnJRARzT5zei1Nv5AUgdFoNSVrBuoZ7VRlaqYtmGn2VPJflrASbbzzz3FSQQsDZhvPzt
Ka6LbH92rdhxzfk1mYHg79No5Sg5Ypq17k7/X/xwEkesrtTzPUbhWv3KuY8K040rWo7nHX7iX8w/
V7KaoyEYbpJRAvyDiDvxYaxXNw4P391wkEl9Z5D82Uz3cpTQChziz4MJCxSH+amcc5h+v7hONGQR
TxNlhs8QOwTjG+PU8uDNNdUlnN06jHkQPuiWsh6nH6XFrGsYSzQ8I0I560+FG2AZzllnka+rJ2Mq
rlYxEtt0Bg35sSDBeBrCdpB/ChbTyIytGhSSqEGPKOL7MWr3eF7rFhncICqwegKF33K6BWI+OYa/
lVeriGH9s9J7J6rexkX7OHsPw3vSYsROrU1VeJrmiVzDvKgEMqhDV80MwXInOVA6VhhRt9QsV8lY
C7IENBeE0sHpuaIDdLEWrTMraHI+WXKRUkXUkC4ZQt9BlikvvwZUMu5obY8YF/ZEnmr7U9mlv9aq
xVMyuzzWSu/CoH82DaXh9WCo8cDN5kuvkIt/C2fesMmJEuU6cWSJKsVjHI+q0kc4JrG4d6VeWTYh
Y/tOos72WmcWzbyaoq516Q7RqX0sXbxeCxC13dsS0Av1EtQZskvoUwDoLjNCIzziNU2wfIhRooXO
S5oxIdlgfeS3/NXrrZVpmHH1qUW80Bzs5hWAHG1CzBfzR9STgkt3XpP5n/MomxJCzUTacnQOi5iu
Q8Du4ZsaOkqbJhyARdNlE5/XRSaDk3fF8VtTHysmf5JBWxguhRM9AzsEkre6rWIXJ7h+U++W2wKr
9OFlbs30JkNsS2qDnHh7LGxnW1rGIXs9FwQZ0ZSrkebKCwBRlZZXGeGAZBwIhYbj1Vihc7NxUix2
o/PlebGuD4/T27V3vCmNyclVjearfiCDGaosFXTW+SIDHlQbb2hjReCurBviKimzM07eXvWZtoa6
pk2ROcONM1aI4FZKwNw2TFQPef+prNZVrU29H308miDQ/3dkmOMBp8NmgCVdCScb/MhfWaO3o8wP
T8DdofIG6qtZ+4wCY51au0v+0YW3QUNM0UV/B1ztlFe7f6Ap/cgtc6pgpH/nJPCnOYpZlskfxewb
Kr0e2ejr4oeUA77NDCaz3gQGJznpG8uzD3bPYNvWt/85dFAA5HPaDlKX4jWc8rClyIaRiGhtXUj9
xi8+H5a1u6BLIJSz0BJeQhL1NU3GjqzcDk5xO2+mxiaNkKkTUV1971K3uN04n03mzSRL5r+bum1Z
pACeaI3/Y4KG5zT+Q63a1hVfKfXKGB7DhS8/2p5LnfszbvZTroL5ZRBL/LwjwGQktWURzeeVOadD
kwFeQ92mxku1HERXjHKeC5ACxIikWmAnWfcdMr15YGTbE49n/1AYSn0t6Ql9DEPr0eIMoKkSAgiw
pu0M9Zbl3kXh//Pm8dYb6vR+dQqPpuugpHRhYi5tkD2OTErHoyn/W8Arg0DCmZUgv90qTmXaDoXm
xbMTSw7XqQbo/R9rtKUU9qLRlIC0iWcJBdWc1fLm2ex994xoknqDfOiBmKBLOYZpseV8vYKVUDgT
bf0miD36uVQhNbGVcJOMH2W2qz6LRq2KsTy6raqtSFDIFaZz7Wo2ifKz9a3cnYk169jDbrkhpH7m
YnwKckQ6nL/Jz/znPo6ofHfrk96QBf6T8oV333PjQo3A9+hM0Xt2Cknt2Nm3For1ToWNeHTKaJl6
apU8TdXjId2VOPpJS7ASqGPSRb8mauYVMEfdeb0SAb32LUJC5ciZgEVh+wxgV0sa5nBo22Gi93CG
9wvbZ2fpmJNXLrIYzyKhFKpZR4+uoUd451wIm/cVqs45RK1npCyu28zZSFotSiBOCanK9eJ8ldY3
k/7qYbqiYFtQNr8z4dRBgWBGaWidOLs3K3Oma30GWxgB9fSRVikesQ5v1BDC4r47+9shKitSuQbT
LZeCFhD35JyFeMJxBkEVMzJ+aZiTrKEKjMS5cfd4r5854hGqyJsGIKq1qzhKOt+jVyJb2vnVI+yo
3/9jX9J2wX3A1EohAZLyz0MXEw+iUhAJOlwb05yqi6OLigkXVxPmHTalsuZs1OYvxZHACsPq5+gn
2tWzoRSi1SlSNA5l6bhaaNCnquPtDPxvuQbPK8VnV2aqZIhoHEKd6akM8IraNrP8eShib9AW9Tc6
LBh1re59/DqXUdIrpEVfcy5msZy0GIs24JNe0yVWE1es2fuFhI50Fa2r5DJTsFvS3Y2MzA9NRrT6
tPJesWob75SppZkMEJThD7+CdxnAhq2LMJX2AH4FDYjehPAG5WK1umhqdF277/HUNwd+ufXVblX8
5qf49PSsdGldbYfdBGBJVX1XIz3ExDju8xMRuP6AY0NH4U1aYt0kHabBFtfp+sInIJhAU4JZRxMZ
N1To/xGZfBNBZJiDM+5KKRnOOgxSyp1NxDUIfMocyiDXbLtC+zatjCeV0/HqXd+8wiaAbNITaA5x
dN52E0MU6/TFt4mcLnd2eIHFXBcpgFol9zBoJR/Yp1HRQ5fS2DeBWyeI75UtNf0N81Cb3f+z6aXv
kykF8NQkxZBjH1VHNDg7mHze93R+yyqdTYR6QRLVVD0oPERVWliMmHvt74X5Xd6GEEhPJ+xVSFNz
qDXWgeREyUcE6tXtQiIlTeOY/3/6Dgirvet1C+BFuqcL+A5iotqoYk/52sgfMhiuGsyEZoJxh344
gH+b5dBUYLDQzPDOtCNyWWskWCjtKi6hpnphDyxhPWbBm/DAH8hBcRP7tkwEjNLuAwNBQkutqHEs
ldKyfepk2+cxAuSTUN9wa9crTPCwyVFUodaDJfsxu6AyvtUfnntjaikrbRurwWfPGX+cWDxh9cZL
Xf3j7hhidzKN/F44v7UeFDuTU2SsE8I2tNlchXyzoE7ex6lGMGrY7ZZBJKZQherdoeK77bTOrUsQ
au3LTJWh4YDklBIsJZFN2aL9CahmgN5lhVcFBVPouGXbXjrP86ukWRsA1/DHqVEBvgyEUZ14tZ1w
ETN7+axWDos2eQHiAkTI0hpBMMpEcH/wPbNyNUek0xyDbSM/1vZ4OeTAyBBHT9ul5dS5cm7k7IvD
YPdIn15v2osBXwqnCeLAV1B4HnL+c/8sSm4JWIfdLhJyEMjZnkNdvJIfLNpP3vQxtO214aG4/Hq9
mfJiVUOfnucExpdlCAjDkxUihFwiknGz96QeOY+o7jFSOhgXDdOc7pHL7e1Cdn2wUk5dsRdoeuXs
tZavk+vFQxteBknLnJVElwHiR87Diy056V7zMUvNKQ0v8Dwiug0LXS5rq89Wh/r/6TTvZCLQ+ko4
TCiqnSAR7nC/WPcfFy+pmFilOwDiUVGdrrSoIUqIn3Lw5Nrw6hKkus/XkAMHYHm84QotzQWrJdza
D4k/DdaxZwhVCO10w9sGFc+cbtyWBHwbTiffM5cxZfHBwWMtCTVBQDZ1FoJ/+ucmgXx1AAbO8/QF
Br/EJehX9k5gw+ecvqthWhucGGVJMz3sx/936+eldw3AtY6LdPacxrHX6Q0movLdtxY6YL9zFi8b
/ohrXSHPxJaWHMc1TB97lC5mvt0nioispS6kJSGRhI8HzwPDksgAQXsGP6gnq1KzrVwXuBgKmV64
U8b5wHb7kwAXe2Mz4Pi/6OUsaS5CHf78gnKE/8udxNrUakNxbZhjyaiDitPT8gblTdi8+G76lL01
JdoNksTyg2cwZWSaTR7WRpFqKGjiwlatzKDI14HmbyFkL9kZnyyVL86UtCNJ00nM/QZUc4dkkJAa
YFlMS9ajcRVqvRzTbHcUM4Ti8HcnMrSWm9xM7Pbfcxe4WH2t00XGmB9u4l9BHzXNIK6QhMSyO5Tr
kPPyVtVYeAmh/BPnGv1PMQHeJhLRRmX929d2fIiQ4Dgt6ICDooVmBVkiQxijWFGGkyYv9qmpIWqx
n+Ypw81ZqBpBCkdMOFNe0kF+8cuf0caEfM5D1nY/VHqbsLCbIbYsd5lfgtFMear6j+8BH6aRCpGC
Utr9zn0pxcxpelBLZ027/RsAtf9suVpZYPNIZlv+Kw//R9dZruR0F8DIkG3bj2+YaoHkdxEzCNwZ
h52vfoGCrvz6nNqaaJ8wBLTDgDTzaRpnBnYaj/6uH9TxnGzmosZb8Bxp8Zu2UVW5wCqfHcLmJQgz
nbV6DWop0Br1XCIj6vj6nVT9nkqFHuXq2STJfIktlC1SEuHXrgDC9tYf5ue/6tCMMsDGHUVQfNdt
hHeBZoZATSx3QwiiVJ2p+M2xfEL2cqph9V7+n4otFK4j36GRECjqlCXUgFYf9y2x5QKPMvuF+i3m
bO4+3cwWdchdxnFqp6dv9stKHggSjU8UV2XPZHhUvvQn7QPnwpzc4PwoZQUXPwjjVHJtlve+YxDn
uVa2uxT3QWjmguGYwuiKN89PR+I8t3lMbgTyuiEQf4J0VkDe5FPRIM4fd9Ufnz2P6fy3E7s7MTxy
0Rum3+z25uiSi37a/V2I89frGnwmkBwDS9HQDWv8T23KDGdtSI1+BPGQaln5WAp1TCDjfEbdzrPH
OSt03FY/kgHBIpdmjOAUbIRYozyyfbkCRwrvDnWJbXAjGPwVJSudwAY3l1TffF9ATts5zPSw7rUM
zMEIL53K/LDb5uLpU3/MQ6j1msxXvbvc/oebK4zeIm81ELiCqTNNuYG7L1TIIKzfpq60NZT9rKMu
LUWdXY46g1T3xeuu4fRtnr4SrOvfdGcd1EuzAPgpsjlpXwT8PGwF9TFrrREvbKdzyafxOJ/53T22
Gj9lDbI7n3TR10H1Cc6IgCcYQbexXtCnw5g2nw1+6qh0GAPIH/A/Kz5Fk2R/UnFOm4lLOOWqLkud
7gpd4V0fNtXgJrJibEWGlXY+tDI9ywZcC92Ml5AziDGxHNUfD3thu3XOk/L6IdYLM8DP7I9KgmTF
QbTdyaP8rXajhzaU+fWXpvNL/kvs78Y/2xwRoTWd6pyys8bhDX3hU1MyEHGEN6WLeiab9q1X4x8e
6DgnodEGXiAzJmpl6PxzTWOTy25XvZysD+fu0GH7cjbCpcOjK0ZdhXJykbjDBvB75HRY/86tyMKx
mH74oWZf2BoauYazjS8PjaRt68ibcmWImsk5Um2fKwhWbTb9kjMnkYXirDR7knPcv0JAOOk+CItw
KyFB5u6dhkaIjsh426LtWq9jsKyL8Ic9tCwwM2/UieleGJ0B4Oy00O5nMwq/FItItcC9hkQM16Wj
1rTkFnvTFIEyItGGOtOCdgEzqBplQ6Z8L8YvdmV6uxArzokE30dXSr3/NEEK9gMZV+s9YjuOKd07
UUo2GR3DCkKRH3doBH6xD3Ty8g2mgrCFPCfqThkqeKaoJ9xLhasNN2Mb93HtYIpxfQOS7duhNY/o
IO6F/9PORj69ZLSiewgF05BTJKZPrNHI5nozZY3vnY82ueAeOwW3wOw/J/IjbYZxRvc5D0DokLBS
zcLqOTf7bLrCxtcZYtwHxwIAqAE3VK89cbWemwkhyiXIgd+Ct0TyXno95p/K2TuLOLplcQKD6N0Q
GOU3+IIwtlW4gOGx4hW1ByyOMPzNKIMyOaS1rHXkjjj2QBhrkZb4S9aHDDSMTcBRsC8hQm8V0rxR
jaKQLHCzxA2YiAy3nZCqqxV2ZfCK19uYJkOp45Ynf+lg9YuiE468OG8HXcv87FY2dgTVWMJvzJBJ
wHgOpXyQqkAFfQ+xk166WwOWc6pUApIRzrujC+k2oBQFHIpNsQdusXEiDOxJQGZDO8cmY2rdGs/R
EWHbFy6CRLt9dIWaFVZuR0/b/3AnjL7sF6kctUsAztAUXnns7rZqWy+tV0+l94E6siO1Asm2IDtX
nahAr8znwDzIcwn5cAoU9wY78iyENb51SV5RLSKn16STs5mnJrzwruIVrkiBNJcnu0sT1MCQJ7gn
x4UzMY8CSUX1cOfxdXLNnZvwDykrSVRRYLoy8UBogN5yGgTSCLJbUT090gvOZK08hPDeX5Zqsaxl
8D2SuAK6ue1DiEVa17O+7l782OvIbqHqpghDod0Zys/859ExmBi8KENYtak0p8D/CiHWCQ39+D54
xvZvAkCKp1CQaS6B2SiZ7/U7uwsthBfSM5WwZz6s1171ns72wTTmjeeJbIHKMZJVFWy19S5Hz0IO
0LNVwKZdvm8T4cJ+sZJoaiyk8sVNFXibEC4/enff5h/FQOnBtPUb8HMb3ZErt7DIpTxIcfG3n75R
Uuz+FP2Hf6Me3ummcfnviUlP9Yd2W/lt4dOT+Pky6hKfCy7R7EmOY5vq/t75RlQSyvdbeFZrv13o
pqU1S3AA2RGh+0dXvWpgwOyS1AinaBh/LebZfVtc15QNCs088Mjfmihj+lrNMykyAy+E55Vg0ODj
BHkNChe335d4KbWJ76A3/JRqXUOfZT38qBRloWkAtIJmpgDrmUeIRin/L29z8i1hZSaT55+KI/Ut
XvdjFo7EgdF307ncAm7EDQnM2WNGHMSoNkpSlxQ28cuF6JomJHR6wvWnFjBC0bQE/YHSVDV9aDNF
/urtUwvRNBEXbFFzcrMpMn4AG4kZ1NmVy56hpzDLaD+3LF6st8nT+llQwfUS+5pSl1PoIx/m4NK1
g7rbmzS+zl7msSafvg/HRfYiEkyhr0N83pwpRPmoq8x8eB1fVjUn2lD2GqDPXngC9spm0E3oEcsY
eoJU5F7AKtZUBBCi7I8sK0jr9Cc/JYSz/zPr5d8BRIQ4hEDV5G7vqCQ6kH8zma1fU1pXvfSll25K
1QS+0ulAZKpDn4mXU0l6B+KOIdTTGsaGl/98igEvv9AKHEDb21WeQCjfqLNrg3XLYMdXuBOPHj9R
M3CH9ZBzkrXpUbMtSrBGbQibTGPYdMhWv1iyYAcIzlZj80qrX6wiwmhEf7aTPDqNqzSnuRbJm43R
J8PFQ/ewAB5FbfVv/ToYJs20Nlqj3QTAUAsjhnSltPaL0TQ7Id0avsDX8VqBnlZYkZI2FFBJjsYT
LVWZbNJOH0cTvRZLFN1/OHfkGth2aPnsTDNY8JJMs1FieFn8w+YBP02wMyHLs/GnbnaNHAQbLCfG
HhmIF9FaGxpLVBxTC8VvsshST+4ijnjxfDGEBWckLmnueMYEX5W+zgpwkssd0/IRdA7EZE6bbfb5
ozA4yClE3lgc8ARKkpPInRx8ZhlBfJ3Aa76jBXtiY5TYMApb9m7vA2OkFWVn/b1u7IisX2hd09L6
EaKnWDnKbyPTS49vNAi/5zNFoGea6StbZXWjxcNjedOr2/qBX65XXdf0sPulT22rzh1D8Ay13lcN
1y9Q+WST++N5skXgEF0ygbTXWTBLlq85Bj85UQcdA8TAFeLWkNRzZLN1lOguAoDXiTBIR2hb5uEd
u9XlKwIFlKMr9Z5U3B8O8yAiclIntWzhSIt7sChtFR/Ag6R+QqT07JdP0W565LRF0AYR2ApQkt2u
E8gatiR/i16gXxQOSdLYAq992ul//c6P89Kn1S6ruhKcuKEORl9WbLAcG2jAKc2QXTOikRrGO+/k
25Umu0Bk7r++yUXnE0rxycADUJuMddPFqqmjhUyob0WVU6d+JPtwVMAAkVXh1vlwH2o6w1DCr6uX
n6RdY8MKXtA/ecGkmJa6yfB9YiZ2/+oRmLtpWSh7lcvybisbTXMHJ+fucW8+jrEQQb9zoUuung+D
ZNGqAjXslc8Y0qwaUYUdSb72D6Bzj2iQ5/LlUR2zUJ1TnXtI75IUJprHziY+HxJYobHmDyrlVxLk
19cArBABSto0mLFurXrjvAyT2XOPaXcGrW9UF3mlZI9n2eKcOWzTwxfO+lTUO24njAXU4VVaWl8I
xJaHuDqy0UOdkjVuGuJDum50UnZt+vzOjTt3Ll3rH/eqQk43/L5Og+hbPQUfm7r1AS/UkDP7447N
ajJFLiuEaBvZiHHCfOhzwrc0ppQMG7B8Z/ckkw8/xv/3Hk0IcpHhM1lJJnsm4N7/1VeQv35fuACZ
LAdPdSUQhnmVNL5t1yd62Phy7Yu0uQfGF+KVltzrgj4ZBPOrYeCcWC2WD7wKnS7BVbNAWyqIm91S
ReMx/Bd2XDWymYVCfzAVzx2PuEcKvE7CRYMqZl1l4GHqeNRC0+1eZEqm9CVUaRw3pfQuGEfZnES6
acTH1BbKPgueBCfT/fAakGv0admwBeNL9X/u93o2ayhPCTdmb/2XhNh/zOGAcznsF2At9nq8BdF3
I50y4otRy80QISGng7hWw0PplGCUbhNlccR+mGDd+puzCgxgs8gXB+/wMeyvvW/OElHDjmtWaWNe
iKhqhNBW6cZc+8h4abkWl9e4kwZ6C8G6iXdNpA/t90L6XpGcE20gt2GYKbWNsbX2GBWlEqE8W2Jt
lYLt2cHtXXjSQWOGPdyzC+03HBRPAhw4JheH1LkzH7df6k5kyMEeKCUpjvPAsKh0YIyi/b3M2rTU
1pzrH1T8RqVeve33z+gQlnvckF0ACcD3n2zKf+Vfp7N7L3WA5HgswRk/Adfu2K2h3gXNYjm70WBa
/wRHjnhYnpLKnRocgH8KgBpP7Ey7BHTbirh/6J15ci24CnJcYTXzzDDnn49HQIeWC6C4ClYTXPTV
6smsJf+74CNvk9hp4z0L+iU1UNVf+mHDfFXOyRVl0t4gaPaNREzT4keTX9lRXF2HOpRsCVAlxnGM
/ZYDM5iXJY8gRkl/DLOWGVHUvCgw4cIUvEsusxPme5xnus3tWyHd2JXDcwbR2CAwI1YpjzgtC16y
eg26U1NII3SXA+f7deTBxfDs06glftAw0Qgzxbv6INkVw2y2DOGyV4NHXerPbA9Urr5a/1H2Xhgi
YI2HfI7ACT0q6KdQGM48Jcvy2E4RQ8eZs7/+fzqQevHU6meZrzaTan3AO50ojYuWJ2FvXYjbxoz3
/vJ5vzRqrabAt1aluOHqGE+ETJAgYYvFQWkikrogUkklmSiIo4pbz00F//EkDbeyVALVd7iwcmu5
k//9/e92PfS+RGl1/IXnSUuarOj7/m9kyHBAD+x+EsirK/StP7RhxYXuZWnmmUSSpehamelbBVaD
dvsnZ/svIIp+zmjnF+XClc6BjKv7TIlQ4G8y6D80NCBZUmTTP2UUrXy2h5h+2tq/qw8zA2zpy+SH
VtbDBqGMPyMr6X/mvWXMyMGUDLoZdd/2/ZyTCdKl0MYT40T+yYl84uRwhdSWAOiTcG6wAypel+Et
GCWZM17PKmyaSd0rvEDeorxRqey7eoa1FOa2nuKB9oPF6zdankuEfNjIiRZCfTmQmgiM9cREe6ME
L61XsCKSeBtKT4UenjkQIuKQflhW6HK2tUkywC47twl+jlDA3hl9TE+0Q43lqgPW6KCyf2Pt3DPk
qUymYGmecSEdrdFiJDnLegrdyBK/tYaQYlCwbl7w0lqSJuKPJ9ioimLE2E8FgGbfvj5DJ6ZfSGwu
NfTSMFt0g8vlLttNrMrCcRk7/+GWMfPvKkyCUfLf4El0ja+Q/zQOV4TZDgzoAUSpbB7pQ1wu/o5s
RPod4qpAO9VSld85darx5OVCqloVPS0b+QC7Koh8g0nXgn+tiUjo4NApQlfWag0sn54OwyAFM5ad
EFfYkQKomiEgz6WquetmEA0z6gtmVEGhDzGMxA9GEUPfc14rjQTvMMRHQSGAju2OLhDK0Td6NiyN
GPWxcv6alyHKslfB7fZ/nI41+FR2JafRi3WcPkDcn8tEvdvERzdDy3OkGXoQV4Qzmj2jlCvlR7yH
u7ZvGLGi0VcyGHEH3OQ79suMebiezbmfvehPQ1fqCbqFWhZ1vpGZb//ru/dsZ7J+mzkKvX76A1zf
ZYx5jEG2HoREfbkAZtoGKgNBF7EaUtIPG5Ew144t+L+PeFuhCCZd2UdrA4lqMKInNRRTM/pZST5E
8dnQTzLeD+MsqJw4eS+WoR6CYXfxcL9TsoDQcGuhm6tq/fyr0MhHOY1Va4UnlQXhEtQDece8bhpo
xnCCVfqbW8nUhGbwLgmmM4y5IzuOLS0vbVyhJ363QbS/QY+DIx0ubCdtjYmsmwbqoI6S1MIm8qn8
Di4JixR+k25tCgPbNwm6dM8iyrZXRpp8qVa2GobPY8iRFWSMxmwDRtc6A2WreZ5zqYqY5GjsiC3P
c8qQFfKMA++LErw4S5QAtZ5zmdtigghbQ5MPLs2VaYgxciPrB+qnlnlt4+YtuG9DfSzKZOfGQKGK
89GpSp5HdCA8+klH3XVju9hkAq4SEdAhsVhznqwCctBmiWMx89ft8RkrH4sqs3gBjxFkdJLUZLCY
BP9+UWw3lvXtwa6L9zPViJ39BMkfsrBg5xMPQFyN4uO8Bowl/hbbZdDGJFa52ZL4YXJcxH/GqRMB
YpVvQEQON09Vm3EAR4gctEDSPT9n6lve1eRj5EPJUT1hcSfSv4zuziK/Pb1DHiDQ9+MI5RO5rTjr
IVWWdR7VKr/dN4OVYXqXvDuLOsji8/3oytSzi/4Q4an5kBckJpo9ZXicoJdcFNgIamf0Z+m/sAMu
cIvLZ0nv8C0trEpIb2H5b/7eyCKlHISUrzR/gtMZ3QYpkAPIxhZHQujaRmYo4OTOSxzKw6AulsvU
h9Ob3tauwQnVTQuGj5q27W2c8KcfXiBv1Zqf0Z+wnhjNanRcvANhfvXVO6NMa5okd4S5lItL9gjK
U1PPrRGKBu0ybRyz1DIdxmOzN3g8Pcc696RO1b+AoQVEnwRHUEY7tFlq6mZ139uReg8wf8wXJ6U3
lQ7DLH059eABhU9KUzKAhmDLGP5vUG5z7oJNZLDf5uCsCd6+M4FVA/fDU/qX6A0KRYssOwrFYa7R
qkS0DqXUp0TJO5T8JYrnfL/EplcT1BcZeVbbkgJcbmO7La83qJsBGNyKmVtrm6zlOr75EdSVWdCC
baOOuU5iy6WJLQIIRVWZK7qW0vhmKBBEat7FDXpdGIHEsl6b7rCAf/dFkC3BehNgjFL9FasXwcj6
lHxR8adsWR/XEmggiOfSzl1Zo/gsFjl3E4LojDykk7im17TKJATGdlhu2LMefZixKGWad3gZGsPG
7LVTHKrsNRPUxAn9z6RtQsrKpLblUXjecoh7SBobvFMPpzsof28J5xlKBpK94qE45hg9FlwfK3oI
UVptiM5XhK3LJiEjv4XeIFcp+Ml7ideniUZiQeOFTw8hY4Khlnu3zdVOHjbCCWhe4KB/M2+qE8VY
s2TnQC5wSoc9TgvSrbaCpzTh5KzOdYEdcewCIiOj6FlxrErRw4EZhq/MYqz2cBL1RoWuQXpAzBRj
OLPXFhicBNU+hSRSDD4h804LLyFKcAHNwJMG/xRTy7G+fCW/N6u/QeFIoUYOMGYowLpnNuD0enA7
uPhnbcKvUSAtCESVJfF5tvWQZUxoGR2TLIBBME7UjtMXdO5kM73/dqaprmafS+BiMpRajVd6N9Qb
/WC4z88Oy/QGnTXyWEcikTjUNWHo76JPlXhX1oumlqooc+/V6gRBu0xxD65UQMv84mMy38u0tinw
oulBESroxK6KxgQQvPmKePhy3FhXS2lvQWfGqNhliI+yCrBTZI6JtPGSHOwxV1IJ38kI65gCup3M
N/fDNhplTrhQdC+fhXguzhuKq3rI9L6KFHkK2PAUq5XzMzbZJYbZPZvcN3An8An61/dna//WZN0t
i+I0tLeY3VhemnFzFggdydXpRAyazBNED1QBhZo1hBSmqBKW9kG7R18vvV2GHJderETLjRTNpN4v
jhfXvWUA55F+43qVloiQS1bZRzS0f4KY/AlJQsQkjKoGKxT5pJ6KGMKzO56vPqiMk0vJ0R1c7RJK
1DyuLOhHYQaxsWLXl62pSfEdlUSBLgEOMpZAbZdJq6tRyCiR3Ur2XEeQhnuXE4Hozm1DQrseZz6e
S5S5XTCDbrEsbXQ9ktT1yQ8VWpIRQAwPKd5lpBNzfxmAUtArEx/hDRRy9OxUsvUZYTmCPalEJSfj
MqJ0J5aC/2rwlUP48jyjv34i0fDOfewwyP4icsGoa/HVt3ldsID4aBiYOlBBCTLww3wc4/8R8LLk
HAkDbKzQAwAS+OPvpWlLG8OpeUkUF/4G0f5fz1uGThJesGn6B72xdg+hHW6st7MFh+WkH7j2gGgw
MmyWf8NbWGrXuFtCgU2Pzg9RBbncf8iyP7Epn2rCvx4eYSZTKR7TCSryfrUBJ6qDnFDLfQwwWPXy
bhIp82c28L5cmTn9llf9kMLs9h6kxaLJf9CGa+wqWDhd+meIAfAvqpdrEhse8Y0Q7n999MvoQASq
rmhYGCQkJ6iAXSbIEDfzoNd/tvE1SG3fgrqFF8Rx1yFI3MIdFs+bgeU1URry2rTG2w4KxzhzAbzy
BGesv9eoNifIl3nFtXaj0SrU25aBxrQM3VkdMmqAM+jDSNqbkJDlJ04je5WPnHQ2+RXhxTd5daNI
7ZJNHsKt7nGGP8ITJwjvnEvQn5iIo2BuYQ55gALP58bMuAsxx5hEzsgIsTL8nqQTNuXXfB5IuRt9
DzCTvX2YsrzPISl4XoHKnIgP2WJrI4YyKp1tfgV0zxKpupQxEG/7/87tjEi7PFtQuIY8qD8HqCmI
m1pCrHWoUVxaESboSIJENuQMtTr2yCQBmP+DT4gKY5rZ8HFiaXqwg9tY3fnZB/dFQZlZtiQYw2Rk
mjQN2WKOkGKZdLzRA3Gwr0Qp0Zk8mGxP4+dzjqOMluD2WrRgfnzf6hwvnaH6gU9lphjS35GGHE3N
oQ09dfbbMb18R6zjstZ9hC7pcTRfWFJ+F9Lk/QGSNYReAgp5FjeHhSa1Yw9NM5muSqmvmXXQg4vL
e7rzsp5TIfTOGScS5/2hvVuMUSnBjLkrjzfdk1PHnJr+Cxt9/hJmn1A/vv6vnd1tivOP4f6FBEJ+
aE+p5ywP5OqtyLFtAQJHQO1LkiRkYgt6obcLiH8E7i8N3KG+aCy0lBc3alc1xNDiGaYcw7NkQKjw
QG8ZQSj6LnG4LLcL+uacQqh3Maqtke6jtM3q7pYDbH6QD0grVCvQoLTELEpyeSRlYa8hqJVN6J4B
gRg9SBXaJdVJx5wmr37Tiyoe+SJLf74AstDhgyJNSEs32ClOJiFPq1ARITLjBknM+MJiLIWslUQA
fp8IEtQCTc98Lqt/RSqpJ/2DeX4FS826fb5pvbbpiG0chYnP7VtpoPCCM6+HMnLeiffH/9+SZhIQ
kv222DJ3/FowXFCmrkdMarmi17WQsGlt2qjKXLYp1AhZQewY1EnC/Q6Ut1lYKYrUNlz087cmFSYd
4MyKmEFmGtfJkJQ7jGwDPqGkyZLUG7Nylk4NMgpi59fFJYLPMEYmQ5C3xa1/kiitTrxsTIoJ6HSp
OJMIuwCpWowfKf4UTkNMK/R4QJR1oaGpWHFy6C90lIiC1tXzalr51lruxzRF1h1KXCQTBNtcepQf
5YnGdVSV2ODsxf+PMyPE1qaMSa2oUlIt5UlHUm1mZmh8MFfGV2Epo+T3f1MqzDMX+5c119XVWNwM
EemuPw8Cn3oQ/pitGzqHJ0GsIypcDOfnRsDLaoSFMH2XhQHn2wAwEjCZILZWG722p+hxZpH5RbGQ
vF7Yk8TaEDC0cnBE+zfCbQPvOgNhGi8aWgqTdsIbOTiVKnwP4PdgWTskvtQ5omJ08qm+hi4nYr6B
N4LgopMCFtRhhimtjI9CEwacCnafcUuIQJuIE9fmLz6b+0IKsfTz1kA46GsnQt+Vm9jdtADR3Guo
IQv7v5k3y6iiuCEN/q35h6DkFpgO6zBrUWOnaz9yc4VtisZX+EJKVLgfe96wszW33e53hqP4vM1G
Sy88GExcpkBw/bWF4ZjFWcmrGf2mdWXi1bkTsWBAkwPaRBSGDcy2onwg1mDyyP5kxVWQWqxqUPCP
jj5HW0ros74jz/1hZNJPZ/oLQt3B2Yj+asE5SzQVVMnivna4MbjFybE6qL9nbp+ycOJVjCWjqmuB
6831xyczWW2AtMmF1Zpe2LcnyYd75CjA/btJZOZC4DDwn4Iw9wqTRe1i63y/7dlhcdhXkMkxv0r0
liYUlTxSxzORoH+W5umuDxrn1hWgrU2zha6L9RvZBglWaGi5AURatjDYhtc6HJ+KrtGuZCD7r7Op
Ac6K4gF3riCrcy3u2ENoQM+pRn5FbNCUZeGanxNIoptxWInqc02ryA1kLt1kjiqVl3UVTkPtncP4
tn/0mz08zjcUBuDPU4l5ozznxUwjsfujeL2wU4TQ2Bnu8FSo3kGLViqc+Ng7DS9RswDgOyFbeINQ
kqwNUk6pi73JdQORZf7O50H/fRF7K9I6rCor3ggaYE+GK5c3hHJNI/75Ci4mfvc2+y4hcuwYwxBw
zDBzqc9i//Pjq1/iTY+y3B33IEVgx9Q8lusBTRX0SCxw5h9hgzfQOnnKSA5IEKc0I9UHL1F7qJpq
HUI/DWg2QWpWjYViViO0h240uLaX4MGzSg99G9vGEgtINjbsGSYwUeneWhXNcdp9Hw7zYCzXNjZF
FdIVNXGAHGv9LL9lIy15wID8rwmVtSRqBRb0EygQ+iRE/ww3LD6uzyfRcedSQA3HGch7ndn+kQQx
BlGUo6aRtDq8NPeUAxUMGWnzRszGQjI7R53ChjDSL04wxhenLn7wJQ+xioYHWhh9oIY93gGhJZYf
8kwYEKgpfTh7I34PvEpq+dBsJo9va+kWTjZVZDCyKMGuUpLj0lTwFPJVY8skb6dlTBESoLXBfpB6
H8yoGkuboVjCOp0pJCnKNBReJjZcogRsFL8YOq/Y6aeYllwmXQsxsOPv0tWJxBqgajjcCQzMtcl1
5J3wviMK2zFv9HXgXKiHQUlgIZKq4tNC9+v7N4pmr4RrZ3F867GC7wwFb8Llt1D9Y2ldGKXRv6Nb
tFgDUAgGqSGkdLIxt85DhK3wRJkjv6CX0q3dGV1Lg7c+K7A5zLDej/rCRTt8N7B7J2KuLjq8gjRm
tRnpDZsLOS9biJwuw/EUVtbLHlsEstLGJofM1iSWBTxTnSU17B6At4nHx+yNOSW0IsK8pedjZBCx
odAONsDExvZpiBee9Bz6kG3ZaaTx5D+JfnGzzZqCOe8aEasHpo7Jg+hmyUMd9Wqv5fdgWNPXFxhN
B0nTd0hDOdaGEQAp87fi/7zK4CAXM9/W20B7SCnqVsohdG0eKqHCR5VvVTYG3ELeXUFiHGUeyWEl
3FJxSZ1usVX/mQb0x7dE1IjW7SnKR0jl8/6XvCW6waRgwwQXkd9OnpQpItoinm9BnLFa6f5wx2ff
adIgcNGX8/7iLV1o/v5Hlh6n8KolHeXowOVR/PIS4YUpRpEPLTS6hARGluLrFdXgs+2K4OcB1lab
a1oJghiD3x/WUQTgZdxaY4N+WxKw89Q8im8SwkMUyqG6xCVk9KgOVwHMjyNzESmDGgMd4qR7/Jfy
KueNIWTufAGPmTfwnFE4kJpSg7tNg7lhT3BDAIpfySuNVLyyitSxYNp31KQWv9gzIyr+cPEldwnh
Xi3uswnZTzGVxgnsyCfmvVlvatAX4yOEEaX7/LJfvNp6d2fR0SzWwSOFxYJSkw06dvrT0QsC3/k9
3KNgQNU2GAJRj3xrySPqw2JljMTzRZkTA/6mCNPJCtUAQJKdk6KjzTRi1HG5NB5BWbxUymJeK2tZ
1RYQDn2T02u9WTk6OGsqbtDLsbYUFIWT1ohulFFr+4QHx9+Ab5I1+S21LH7r/n0T6TJ73IIDRr/P
Sk/2HBIcVTAixSp6afGmo6jsuPNV6fNXXNljPCElzP08XhuZVT9JdDc1Cuy3tNzq98IpcZMyZTaf
sdj8bSyKGRxLwLtXnp4yOhm4qvAwxrF6WQFeRjTFvUklWtsk7sZuSMRkEXuLC8/W9o5y3yrGi7E7
uUM7aWHtZtrDs6c6OgFH8s2xW1SoC3YdHVtAJuQGXqzuV8dSokJr9+xXOZhYiiiW/fTj/6ssI6tG
jkj44uFE6xe67CDHPZh3Dp/nx2g19ziUB97GJ+kek3sl6o8OwidfFl0Oow7eVbxbpHhhUmgD7ldJ
oJbXkulwdIn9GrSUyfj+Pu1nBAjb7SdfEV4dpzghkhuZ50B0n59tSSL2YB/U1SQv1LV/Qllo5SPe
X4RiwmZdAf2sNSb1+hvebuyPO1v0AgCJzYyoDhoJ0IaYdwsEahSMgcelro49wVaWh0xORRgIlKSw
siFMszFCoYkJuppoTvjUxOYA935aoqMklKMiVGWekNHyhg+ciUlfdRcW1tiu6upplMRvXURqS2hl
ahPp73yOg+1f6YwOEbg0f3o99g9BnZ7QaFYWAY1fmw45kz54JMtRXRoViDqmxuW2gIlgqmrW5Z/n
R+REwrXj5z3CenxbM5gnry+i3zxkMxR71RhcPZ0uOpf5w4Zv8gTjUYsHDPDEFsItAYlvQlGvcB0b
RqzrF8ybaGR7DKJDSNWa0EYWwF2BMbiTAgzg942kPfAp71GT9aiz/+R3buOMFehRfxpLZ0thNODf
unkSexgfGKQ2d6naPd9eGypitvtY7QCmeGoZte4evnZmHZ8fqyWMnyf6s+7Hzjc6r2R0RWWDBQHw
WfyYaM2n0sfKrARDJcCURNBeYHdWddSwDcXXfui7Yo4tjXwmAIeOoe6IOS3pFpx+NXWsmWLFn6uI
2zCrBqJ0wX0jXwTTRqpsP31pkZkQ2yRnc6bZFJ8cdHcizd++WXj7tXbRu2zB5bpxKMWnEx6FQBsD
Pq/SBg/rWuOCUIPtesLNG5JD3ydjGKkxAvVMxUTvsfuv5pGhAKO37N27iyO//6sieNYsmaDQyar5
YCEuzKPlXQ8xdKuM3CJVQA+6A/Cov/bMHIK8kgBLxlTFe2343LSXgvJzvP6gaCVfkMfs7znecLpq
XBPu5M0Edh0Sjnw00gmdnUVjmYVQxCHfelzja9PWwQX3x/i/yu+M9XA6BgYkDlhEjM+4k6yOdY53
ax3485b6gmQHMiY7O7P5yrGKkCCBHmE3FIazjtRIAXkdTh8Zr0c+Ur6yQy6KkOomSJN77qara0Vi
lOqTWO06b9DHW6CvZsJnmSIB6nUh4bPQ+5rSLdmrcrZRqNYXW/D9eNkEXV58K3obEHvfc7fPGiGI
DExJK0Y1ywU/OTBIyh+m4vWAe+3l9cCroRuxsar129m+z+TcKwNDFQGigGFckT7fKrrZOxaIOhEg
2lQijzN5Nik8Plld8I++0qZt828emX+1TwsFa+biQM99TYzOyldmgSoIBZ7TjqxZ+T5ssv0eWVu/
lKJbScI4j1qmYQTNfpxrk7h/+L3a+i+7385rEwp80CjIHO2Rr7brki5jQzBa8qJfof8huUEEJ8xk
4FWuwzMcvSoTUqWcr5xOopA44i6rFCV1x3qbdv6a8SY/NWToih0x1DJQhz6GRqopZZvTJzQxvIZJ
mhh753f/Ir3vNqcQw9W3ogdvXnnjfq1/rTKAHsNoCiacvQpvISdi26UgHj5BCPaXTQIFQAs1zns1
UPMzO3LuV+lL2ZgTvS9w5k2rlDqVQ0Hx5KppEmgW94NyM+LQUVIi860XIB5VYklYyNpTurkcDxeH
js5dB7C7huvWZwOCil0KbWIKBGndgQl2LajzgOGkeY3BT4pOYyNBaWyTi80bXsWIWxK/eRTkWrpW
M4DSRYkRN1m6flfEBNop9jLYYDxwE4zE5UgvBqntXwyWkhei7nQ9FXsuzVPe7xxXosY4C7ULAm4R
laYUjA+7nmspmd8MKrRcup65TZPliTDz7e43TFZ6VrQAwAwWmHWIfEgOazUTDuJayecJcEKRWGmY
JCyHvNDEXezaxZOtN+zBWkVcyMO72VmDLIj8TzTFzVcIx5ZR9jHfnaMFIOuzvoEQqqLTc7NNmYZk
IBrMQUKT7VfxB3d53ar7QEpUttl7Go5k5+Jne5btnQ7krqjGMQQybtvHGCPA7z4UVuwS9pMM9YUK
98zkohPklM6DElXIMi1Nmf5dJKMFJJ6pxfzbWiDx4V3xecy9tOr5Kx2TdsXVTQJv5/FfnKhF9yO5
mxxzwMz/kDo7xCTnOWzplMhw/gEoAtz5/JzzEcyu09rD/97E6QYvkrh5d5aKlyYzDJjJq+j5fIUQ
v84qJjeGe3b+WwtfpuTnaZk8/0JfGXwg86Y/x3woNlkKnqFMFzSnkDPCwM9XkWJVBoDZee72+/ld
7CFiXQaCAgR63CSl5PxvzgXa70uLQLLgvzffCIgefOS7UUzqv2TRosJrJ+dROqP3ukcITgZySuTd
ayjVK4ZQgJ5LoGsuxw1nmbXph4OWVVAyflY9BcMj8fqmSScHRSuDSsyH3jBjOI0vFCFOje9UoXMB
Nr8u7/ebnKz54/MbxLNnqpORbb00zB9SU143eIhbwtuArWKZlI6vD6AR6q+UvnBO9d/ZzYSRbFZV
8lvNTeh85jzfHyp+WyIwRqFup8qxSsv2RSLUQqU6JH+uNNbrugs7As+JEZ1/tMeMep3yP/mmmp1x
7/vK+AkNSPsYPKMkbv08Apwn1VIYzCB4pRYVOLbBD9jNxq6Z0fUB8Nr+2ZFjkm+yBJQCguh5F9dU
sNlHT4JaIa5t8gjdEY0rgp0gvWa75WqA5DNd4C80t6Of9eHkP6ClDdK8zYSXcVAojcPrRgRENv61
qfB4j0gWlzlh+aSVi0usjxqNaiq8j4keF5QOZS/QOqrOoda+UwmXE1D2/XPXXoUcDKXzRmsRWCf1
98brcQNxMlEolYQiSChpAenFU9q2yDV+256WAbATAchjbiSqIttLFEeLHRu4qGkEIMZfUL4iuoP1
s1qFlYNEAz5ijkBvvx1n2pZq5ZjabL1XyIPPKdGaoFlVxPog9C2/VU3hEtniu6aTK0tlBBG/14Yd
JQy0u5SDgFd0tMnv2JuV76MMgvjQ39W4EUR1U8QGtHhXDqFqDR6erqhIK+tU/8WqlDmoCdat+s7+
jEKCE4SzcwE2s7jx6uf0gIhi0/WJL7DwIe1daydNkb3egyZdnS6GJogsJBQEo5tRY90y5sIDYlFf
EV2BM6msotcMhkz750HUG0Wh445x+HpuEQmYFMhlAFVPQ7azCk/G6J9sDkKj1FM7WSxMYrd4fnM/
lPU5D99uyTGe0luo/RBwsB4I6RzFL9L1MldEWAy/vV9/wOCR16Y+mlN+HpslVITwEEb3yQ8UpRYT
0TaxTAu2QGPvFsQ3Jqe8rmhMNPT/04GSasNdUEs+Bk19DsC3JbH/OUbNkxOlTvFmdAl//F2gEq7K
6E9KnLHdRBE0I+MzWdAqeB/674yKQUS548DCaQoGelg8NRxXh/35iIogCuxf1vdf4gD9p5CFckja
rSvmVI9/kdlPgtQBODP+VeBGEYJ9sTFWoZqxTAnk4VugUstWegB4J4uGR2gGVUorb7MyZEQHp+a6
cnyS1tt4rddFM8/ESaAbTzZ6oaKe3YOAYjXcyN9VKtLQ8vrdJ5IlwYLd+NsUtFOYDKXN/6itLCVH
PsqsmTM2r48/KttkNHRlc2E4fIjYZt9QphgOP4PIndeeOxY39iqmr/jc9YLvyX0ro14vb0iML+gW
8Wc0351nkns8RdNM9Tcyk00jGIsfRDdv4hyEzoA14XvnRYFdx1UoSTUc/P3WL+0AlkEgNez0dSrO
MJFUHfDYMmabrh73FsSOoW+IsLOVylwYY7MYYu96OkFQ75E8pyGiSpNEAHeVYAu6RlcypWhNXl4u
GebTVX23jLWYO+NZY0M8LGI614OH1KOaSVTRfzzoFbaVXYY6TJ2gR8zvFiZlVTlCP1I8jzOqagY2
nxiLrmPDQBKsqgKLkQWjkECA2FPvXIYnDXhyShYPkPbIjiJFpWj1tPbK08d+Lc+YRYtezdcBm09l
j5ArZ3iqbGg4C1zDzOSKyAfL+nTAWx3FcLHR79ABdMYuZSlO76bucS2YU8vKHCu0goQNX2asfIFn
SOB/JaXM9TN0Vqf/f4Y0NleWUtGXA/Ug9MK7dRQNJieg9Z86vyT0DuWYR8tAD8Zpb9fOShPpp86W
yiVeey31IJ3c8K0Gwe+9sVWLmG1UmKq1yHOo82nrqAnyHGUr4uG+L6D3GKqRs+qCcTl39/vCCMC2
w2Hh5nTa0o48iyXbniOPTVoy5wMLAS/EXNcKTJOu1+Vf89wxlvyICsuU4m+Yrlh3DRHfNv1aMNUL
ONNxNDywhcvrOh1oJLmgBnUCbSzJCs6GWJyIdjcZfCNOIyC35AN5KoZ1vqyR5COBf3boA93RhdRr
rjNEJ3jSyiHoVI5FZ5p6N/9lP12qKVbAejdn+uB1+DW3Zo0k2GB3EyK+JqoUz8yAaRkf7Dw2ugc4
hNE5O9s80n8E6mt9jtLjHClKXCXMsj77XwELPXTvTJ0lrip+KjHM/PgJtNtK3doA7vcM5ldWo0rt
2nW9jxuNz+Wp6p6bh9NK4D9FHr83q3xLtOBSbCB90qR/jQqJyxGmYoM7G6AyBzOVtNW+KeCESjPk
aUfw3+QBPbTyTXM7P7ezNylrF6wSCIMm+hgFbEsrkmx1eLF2AJJbd2H7cprhVysfbpmNlTkdnVDf
pKe2Q73lVElVXj8a/KMPYf1TjZIL6c0elMn3Yr0+6rPTlJ4/ynqnErl1dYNS3eUXT1srJrt7S8xN
zmrXrfEJC3YuE7hVEgdUYPaZhHltsowhcKGw/8cHpYZ2lRrWyKI7JdRQO+IHpT0SRO+FOOie68yA
QclRd2xvYtqMfJmc0Gart1zcFTwLmjdPQX5X0IY86Gy1dR3eqtjC/iuahlvqPP5iiR6fj5Lpmm1O
eOE6Ak71zcPZxlOScPYgsH5QKzIAwhqkpCr39Tf2QwUvDC5NLlNRXQmiiC52HXEx4OuHzHJD1nKK
HE0PQ3SkXmLLX0BdqaRbXQK956pjsr87WJ4Ya36rFmPwoQVR/5Do62LIBDdqOmLL7CeO1PPKTfKs
oTwD4Au/lpEEqXkFKPimNr1uFigLpynfDADByp+w52fNS6iq66FSKZ920NTY9cANrGW7CrSEk/BL
yxTa3KAUR/sJfIgcS/tyOLT7PKgVPIWkiFfDCappa7WA3z1eKwStkvkxdW2JU2jFz0qtGwfiTPmF
CeybU7ntWL23od4Ju9ZUWcTnM4HojeUkCRXojLrKnba/+cpvyjkOYP1oymdk45HhMreWu7oURP8d
1CCMm5avHhvNXvixUT0WZgYfhZzfG5xt/sal6nqBWl3be8++HkzhRMq9CIXUc1NpDKwQFNV+Xt/b
VGhQx0B5cdiBJDdhaz6VIkyzQeIdvH6zRN4Ek3M6w2CbrVdGaNihEMqhP4jSBxj1Djd6zmOKydv+
cCz24pz/Fu2u1V//Fs1VIV7pn/pyM3EeDqHVNNED0xWiD8KjyS8F+QLGw80H28Qe4RADB12awgdB
yjA2yGXsp8kWOT/f1W9BIHqGl+Y4wX4E8PDeSq5qW3rofZqukNu7Ex4r2zN4gOwFsUoiUPopLKys
UmEl1R+UbfIHu/+uXlsx2USf09VE3MHIxM5iVHipcHi2hTv1ktSpqMKq+9eb/KjrHUGVN+pVpwUl
ah0m6oOtpj2Ct1/fK8mAKJ+nTsrGBAJN+4BgiVxPBWIyoppCu86Sau3FvsB2IM/f3CC1J8R9oFFL
ufoicDvYnlftH0yC3LUkb4Iy5JSJd1/slIlhxRLQEp9T5uBmAiJdoquJt1a/K7UNOoWFPE86jJ7h
atzYyk5iWTjJ1PQm4UmAqZteqXb2D7ENxZKTl4Kxuh5BDjh2Ate6XLlhyoay1ZXXCVyzB5tMekGn
E1ilO8YCDnhAPY6pVFVwcJywgqiNph6RO8/WU8xlimNYESyc2ggFDgVbsET04s6wvISMOZ+hdbpL
l6YmXsWWF0uj+ov2W2abv8cFeb7EZhO9Zr50mGLdHpOkSKB2AYQqmD4P2+e3Ddfnf+OGS5//+Zs9
u/JRnJsbKH6gns5UFTLAcSuYw4Y3yasItd++Fe7hzUBBiNxNAXdIGHw22ZCzYEZJQarUFwjdubME
0cNBwqFkBN69RES0yuBZhpTrygZSxhC76pcCsCAhZD5ukPUvV6NiWJgVmkSp69P8QTVKekB2j0Re
Lyk4sdIJukoDRfy40t1MRsgZrFWh90GvRr4PttPE3O/fb2j5zuU//9WKWYaejsWtFrC142dEiegG
Q9ydlvFHwvTkRQ7pZUy5c3Sf6IydVqD3oHvNVd7lLUQsM4gg32QhKYXE9ql3EllC9cLtPTyTQvPN
W5qEipAmyHa1dTHRK102ibWmr/CIucryfwlm/bpu8jBcRtkoVmSiHkNpVqhf5N673gXGKIczbNQk
BBWYq1vbja42mYVbkryz7zmVqsAyDQweg9Bz5a49Gnn9b/1UpkkjplyOOFfrfnwjkd8Y8HPyy2iK
+XzNRGKE/3xpRrJ15O/X2nkUE6OPcAUheVkLH7RQoXYjAnAadcYcFgkNFR6bWgazzAC8sPVRAQHO
kiF4HdpfylQaFNnPf21k3WO4pYVzd6roSsqKPrc8zAGf4gTlTc+sDpsp3npPEIyHzVcdr0Sqh2uz
/aWV2/pOGHNGZ+LrpM5Wo/rrJAusHiGUhs0Wlc0aB7N1ytLEnohZ1nBxdiPAjxhQ3gtWch1awT6a
Xy+Nhb6exBidDuiH8LMLvJVoYBxUA+cJnUoMs9vb6t0t12ceTqMeyTvScyu0I7kV3dEDyiMCO8dS
GIfda+l8Us0yvful8nbIjqeO2x8pSAx+WnUjYy9B/RiiNg0F1i7zcF1vMDCxiJVU0rY1RRpF/QHn
XnXcTkdgXMRxh1Ux2KKhALnI9ivs+Pmj/dPSLasDrvC6nkTrBlz8VqIJR7X41R6v4Y5rCxPSWmZY
E236T+bIg3IQv+LI9k7hAqXdwSSTI9bi629yqovyIAktuYduauzfsP8w/3JLhkT2rs/y8i/lhwAU
zjpGhVYTPYkFOzXShFUBvJGZRiDy1z3SyIe3IAYudBRjpXZ4O6tIcaRt/abmEZuUN4Bg1qiWC9Rv
U9vGCwrOcnWkOXdKQRPJvG0NsFyPcw88usaAJabP3oLf00nbb5w6Glp3zdRtb1vAuR6qF+MvDI5S
cEbqKZVzfzDm1uOhv9PraBPCzjh4qB/RflCG6rHLWN9NhOmB+A60h9op0FDSX08FE6gvL1C9y723
5/MK5x8AaTD6Ki/axf8XXVhK2K4WGluQ7lAHmEstnANidAdpOqoR4L1zNpGd1j5bZTGqI/gzZ/NS
4gdcg+8DXFzB1LdK1f/IkiK8SFz8CkLyUeX3bszGTkKT7eindgUXXDi6KV9Lg6Z/y3bNhfeHNi9S
3HXNRrmqXKGiV1G3RAITmDnOCR5ZAkiwlMcXyUqRJnfTjSYLBurVROkGCZJVt+fbWsOF+hb0OXX2
iF1UnaHxPXu3RdiYmG3vBf3C9LwAtVCzUkTeTOl+E17SVPku+PlLNr6t7Jzr9oRnRcUeX0S04ZeW
t+r9QWsipwtOVRjvix181CsscsPMEeSpxqsadd7aUjvcS1husYVnFymmJF+axkxtFp4vkAIMDSLC
BSx6TnaKO2p6wlIJft2Sz2qTZy3uzSSUP+Coj1YfwE0k+E0I+S5q05VTBNTed64bXACW5oHj9dzD
GHGwokiKvXvzC6yjc9FrZipwCwpO1suEc3BJXN60p5w9k0l0jhH1+MQs4h/jsfvVqR79Y/l0NNF1
B+vFQ6baGO7+Kqcz7Rc7RvxRyCTkvk8eKwcEX10ph+bzQqRXuSqxiB50/THsaXIPsGcTI/cYOmNR
RVE4Ux/7TJg/wa5g67M54BHk1qDxobfMfSr+VD72seWNzZSE7lDwN0vB8mV0kmyRrl9lMgNXydl/
PGVpb7L0+qVMtldBriSmamtRvhiWWOblZ0RqFQctnzG0UWA8mN2t7knhrJQND3Lg9S5o5dknyr+q
2wF/ksJplcVBdvkyP9Bstf2EyAIb2eSz5wc5tLX2t7FQTOsBUvvRnpxs4ztmG/kMi1QD2EYBwX1R
dD5HVb0dRTIuy3SkQdZJnPhwvxwRXGqXzE64UXuNwbp/DEGCB9uYe20gEMbLtRO7VCr69rgDotTX
qLy6xUW+KWatyx07KsjIR/0hvH9zyW/BR6tdpKgowRicUnvaVUO9cnPNeDiCy79LUOLdeyhrv/I5
5jzQLj8zCgVq1W3yPqT5KJiq1x33RjnjAiF2oW5dv3Vl9L0Aw5nEJz4u0FLi/+N0ad7+w7GyxWEJ
XtbrtsdROCIePl2x1sED3FMmCbC/7TpmWeXBqOZvtDfUR4ERAlyjq6rXM3weuS3CvYAHM+veXzcP
Jp6yk8+xTo6/5SBVCa2FUOt4v+BRiejEAe2swzZXteaieUu+hG12qs9XeLBz19/mEEaN1fTPAbfG
RUIBENGboRwYseoIKfnpetTpwYMkA2wtfwKNTwP7udAOc4lT/axiC+eM08+YTDh3vNDQhJmsVPqe
ETux1pXTuBvX32XvgTquq4Zm0hzhQlPKmEgf8lcBRUqzx4hb0JmfdygZy9k+P8ul4zTsFmB9klNk
xkSMxEUI8/Tc0Ch6Ox3WaD4M+UIYSFWi3xCpPcd+XmFy2clRehc9HueXJxjGAv1nlPebxb67+bkD
4rz+uyTB/CY45ou/vxeFerxRSZfy0aNVEqKSBZ7Hvth+cV2CY/BuolVefuMSPQdr7j5BBl3UjlTt
O1G45nYZGDmDLSP6Agiz1kCguK5QSDWkb/mBwvXPMAv9cZ/lJvKuZR51QIPmgx6OjY0438PFKB2K
NvpbEA3YouxShr72Mphgl5i2hqaJEJRv5c1+X37wEC0qAHFnmUR79KwUrNb2OVytFKQzuMV3F/T4
FnuQuZbhff3FpcNvnN8U4AsZvVr+S3GMjd0fZwDsZvNkCSTd04rUKUx5355uFwqt+fvlvW2x1G5d
qHdm6nu6f+uFsMrSJ0OhdOBv8xFgG4GeppuqFKPcnmmcBCu8hStorSWd5EI2GcReTh1Q4NR8ESv3
PwgdQioyZVIOFSH2haGXq4QKQOOJ7kGH2NZERl+DvQ+aujiEkMyytCp563H8SjGveMdrUP/dnm9r
8GQStwxQp1GIHVbR4j1FSYX2ow+IpKoBopF4XewrBcL1PMmVXGduSlm9i8tQN+NcYtzJCNb02bik
I0iQt0gUQr7e8hr6w/NbRgkUmcBU/Fcz8/NFnmGpCnjeGeFhmHm4Dyf8xrKT0yQh9GDHI6bZE4lR
1l39nzWpSwytXDhledQT765Jk7Sb7DMj+JjJnIcNpfid5NwtgedwzXWA4h7q0AkiGL6Dyo7mFEHX
BugbVpjGhM1HJqRX2U3fZlBTKHgXAl0rLP/ITtmCYGtW/EmpiM+b5RxmH184z7bsWgEtRQLl7DpV
xMeh8O+E9WwL/QVWWmpt7fJjDHZYU2bg7htCwnKqR/cahgIxw5DUPjvwZjKwUMDxV5nu0ikKY7yn
OxyRQ4h1ILnHx2LhNgLsIzSOmi/VmgPDldDwO6Y0x3TTC73uPyIVtRBLFPOqf4uSndCvozasuLhS
lg4mKEu7LnhOe3fwaNqp9ODp6k46a+7DT/EP7O6OblQcQtxj8oZo6AgU+QQHmGAZfpwmNVfH7FdE
RE9kNJstXBbBoW6F9k6FdHQApG+FfnI/ALFlyMFq4kguyupKHznRMmELxLr6K2awlPlXgiXGxb0m
1Tm2wFsoRc1GBZaivf+pLt2au+QpakkqmynWlG+wvxLL3jE11Uzye7JcignqZ2qbrE8T2KMPDtY3
eJ/mnluJ3YEETRMHdM8kDX9PcZmNAIyULqrbqR3xUf+xyD5BJTyacqLRsxgHnxsZCIEXGP0Jt+xf
aW17ZlKEMm2N27FW/oEHfJYILauIXwGqRbOo8igfmg1RIRD40Na1ODb2EPAXBRwKQLtsLSlNoAyd
ZNueELk5UjiX5J1njgwrunTgad2jt9d+xGn9mVZc/in/hfbeCGmP6vvzSU46buhmQU4HzpV6+N+c
ylWUaDT1OCetlsoZ0FO03aV11Hzu5AbDEqwhZpg0E9pkLSUdzTkodkPYYCchPPklspU1hcwnd2hO
e4LxfnLq9LukschVeFP8z038tGDY+shuS/0U5hj3Z4ewWJ6bsa9ntHbJVlQbOsdRcjXA73D4urfl
d8DcLjpa6/o7qKzTydjSVgkK1zEE5rodpXG4ZE8wvHBL6yhCpYwO44L6g/P8TgbCwSwkKCmOJBuf
+PAZtJ7moiI5oE6qTPiaaIyoms0QP2+ujyRuFVocR7y4Bf02fiRfr8JPVf2DR2vdkGfkcT8DxYof
av3LKNZNi+K4+XNarzGYYSWizFzpnae/fMGUZzhSg+xUH1hFsvu/gThrjvWCA+NgH/kCXIsX4/52
aHYEwaSIRZPVaXq+3bDN1i/qxPu3Ajet05N6PpyOjQMVXpuCw/d7Jsy1vxIhQ+aLa4RotYmBA/21
E0Qi+jkZT2UT58/WjKBDkrKx4Z8eHf0ZxZcSSc/n12Xw/ErziaPcnDQq8wW6cyvUziTS9ZtUyIZE
Tbvt5jdZLobdpe/gtCfTHUrLWLwIdMSVtEOiODTzJVq9huid5q32tLmgXTsxSDSUwzQIcE5kCm34
wpC2dvX1Zi3VZyijvN43JoR0sqxHUyvqNT3Ct2v6+gJFtQ24VPb38/q8KXax4hi30arj90QmaxVd
Zrtde2w3L34Sz8f5Vx932kKjgCznsxZFf6oa2NsYcYCF82Lhq2okJr6XhsuhUf0aHKh3EMTEsDZO
qhgezkxJUXPixycXkumIEIO+KmVO0D2/9HTRyTliaI37rHLYsOHEnP0pd1LxTlnx0tAehWrxBxFh
uW9ZMjlugcGkW6GC2dxG8+PBg4K28Kww62479G+Ljj8a62yTTAENmas9fWgwBk1iN9+S7nJKUkL9
yRVN54krH1tpZsn4rZt8BIRd7k+EBvcPTiwcB/4SF4uf3N1cQQ8Hj9w+7AJ8PkppgBS/4Jc0QjFF
Ptib43sWkDbNPtKwIJW/unV0PciUQyDax/Nh9TFDE+t7nqUFOLNmLRNpwoYHsm/FuO/4N+R0zx9E
Ug+G0CMMn2y8bQpHtT9t9rhE9EylaQ/gsLGfA3wzIs8jtSDJB8l+inrvALZudhrac66abvkVj1yh
H8B+fJKkATDbptR5ZDnycOfs8R3xQEM58Heqo4n1dB8kEOrOTsi/GOpE3x5U6AQkVE7AS1jLbYjk
jYLmC/ek+o1ktcg+32QeXgE+IKJhkfRR1S/pggTAKeodSb7H3QTAO+MvcGa8KmcnpNEP6XX6TOWk
6liGeYlUSNqogOFnG34xL+EB8HsrhuHpOZYKlPcQWAmLid8r8ijhtUY4jZKvyTY47B02P+d3mY3t
fXmRInV9JDvsghbc9duvIFsdUcuVkS5KynhiTe+yN7RFBzXEZeVF0/G5Jd20NAGI1o8OeXkUdAOE
9Dqpg4BBbe1tfb+mkoCXQtap6sb2G/XQwfMsLvXiB5h6ZndrPNKv1SHngbtpTKk0MVlw9HCi9Q4C
gKgrHHsl6EcFt7dmyeYWLEPvSecKz3wTsBiti87UIc+B5NZ9KA7dydWkuBzPs21awORjPRg9kg7u
EntNNVl3zUgdUp5OrDf+WETWj4A6C5gijxWMDDKnfmp5pZKwqg/BjXTyvZkFEqOZo0JRTZrseQXe
MVPTAtVCXCPOkCwpCNnMdDkEr1a7pX8dX2jLK/gTmFXS6DES0zqz5DqRRaGHAQ5inPm/wucNSpgl
76POF7dy3aUhBbdKCklPEhNlzFDWk7XZjO0jYYE6zk5HGCBmWKTtB+ReHj6wm65xTgZOqDT1FuWY
Y7+IWRl2HwUG1v/2mKoOIm+uVgYo8kqCccIhoCdgl8ANU9VjdlwhXeasglvSR3HexPT0g5G65c3w
qm4C/eGQ8Lzi9oySTaXkBYRHw6oZpyroqNkF9NeUk9CVHu6jLDvTrc4zGJ23EV8joHbQ7z9tZV/t
gHf7tuHvMY3lh/iFUGi7XpaxMIBf/Lvj+B9YaB6K5aLGSX48iv9qCegMVJknA1rKzPE/UfExR7Gl
8hMCgQiLtpTu7N+Iizt2EHOBfGPLOiWTvV7eT4rWcBsA60fVsUOCJudGBXP2P/tfspf/VIPOyIdb
YiQnO6oDrUB5L9g5PXjPdFAaVf0f2S2XO2ZWrdVwg766hvQcqit1yht159vrhU9B9k4nvAzpR648
g+ASvauD+P5/x6AGVgunI2GdW/z53ismGQdnsWVgEfmRIIz1pFYMLTbC/eX8L+9Kg+BCfUzrNt0m
rXIRWcgdWyu/eFuoWhzuerbHdHHUsH16Z2M3d+XEzBWRBxNfs7K3TGtJGorZnVdM+YOM8l8DgbQ7
SKyTzlr0Fap5ffaMfkmkd8ITbwEhM0NVBPXOBeG/lkEf3Ak1wEpjjMXw6A6iTvSAqzwZvKS1ycqy
LKSTaLNnzp0VHp5rWTMgw5K7oiagpDhtXHbsC/kXJobDzoADXZ/20o6hzUr6EQB47awyZinmTewr
9OxzleV49ipTpT1tG37SuOP0Iogg44+MwkROVL//lP65tYmAbMxY4sjtg3gc3Xh/qS6tIvfm+5eH
5on/mHcuPhWcHiO7aDUkRIkwQmAURiCy1kSb1jEN0jt83+oW45r/P4AvyjRAHbGruOOfXq1oHby1
f0hdPGiYeXU02baJvMYHAyvfi5eEU6v3fcYIQf5X5qWqfLnlvGN+nz09C+ZKO41Ol9g4N4cYvjNm
PNroq+uI4b+jrGt0FwX/rSDB+2d4vHgcUzljLXPq7Cx4l4miu1+wyYESGj7d/iFDgn61+ibWfnyY
NN8lbET9lp3/bI/WWSSmQ1gr2Y4Gm9hKts5LEXyOhocPUbO2fUGWTjjAw5Az7GOq6UfVzoPhJgL7
Ngkho0sQvTSMHlmB3wo1LtxMw48yWHMwzzInPxKTlQXF5ZSyc1JPXOXPwZMdXU8ZOHksUZZ6zSoJ
2ArTaOSGyE6AfKL06E+GYaNiR2UEEadh35hy3E5f8is+IoZCDwkZGvhwhPnPh8TU3K7PNClWJxCD
ajCKZgbVm6tRmIl0q9Y1Z2ARL9AhnWorUbh8PdeydZOwJQ9YD0Y/G4cBX71/4VDrrmnvawSKNfQm
s4WSKQVIkpI0mIF71Evd0tI2ryt7KJ6qbPBWTp4tb+szYgYX8i40cLSgoKamukGcZesVm846Fi8f
io3c9ncsQQVDvtsBs2oXGzxut8rnqAs9/X2MXkncMOs9c7p8K3j8mJaMDborlYxPRcA6oxDY0OT1
Mcze7uXnOAt2tQHNxiFK+fJmGfFKYzOI2P1hHPyxAK+9TjqWWeDJBLiNeleObR+QQPZuB8F8X5Dn
x5kKbygkDWnhg64BOVC22ModwtyaB0uk5exPHN/tzwBfz075RsmE/EgYrR4W9v+G+d6S0LU/rjJ/
WgWyXJ2kxyi4MtHjFpkwQuQszPjuc4BAMC5+SFqYmiZ6xZT2InDY8qnRW9DnPY1bzi75+iqWo3Fu
oW6E1qf1hFR/9vwVk6TaxKvMljbiY88fHRiZWjSTQeeh1tqR7LKiXxDV2Qii/sgaSbBRpV+5wmux
iDUXB9K95eUCTpulw0dKnInuV0i1B4jJPML/sCtFcuDx/Yy06watxB/EqAGsk2IjZRqtaWac+K7H
i82fYXVVRAb5BgLEWmbzv0bL+zc0sNcl4KuhZUyTlfcqmhUIreWNE3/bCkMbVvCdF/HLsR7drTJ6
+sy7dtJeKWc0J2GCI0u1oA8tX2uZSuz3BO1QgBp+B7ebvu6u06llarRu+7rfpFVGx5aPJMPhOw+O
lmyTZSWO3P7pcaBLrP+JYMBHC3IRgLNT8AsK5nk2/2OgXCTWHHncMCGoyhGGBG+TR5sL5eyzR/4r
nw6JKSa/BN+REmtNO695Fe3BMgbvuW8GYjKCI+QKi5M0AS/zjbsluY3fuzVrKDm5sZ437jNqTPQP
e5kcbCimh4uieE/Y5vnypDHzjZ9JiiHQSIKfuMO0XLS3lPLh+K58NBhRMXfemxAxez8/DcmVUu2H
mk1lLUbbRjrEqPr+13tTJKfO3yUqH1jHADtqQ5UVsF1nCRsyBZLxV6NOxxeOBz8Ar4RpPB1/Xo9U
uwI/40fzrSWbQl/bktjs+cU/ROeHbWAgu0VB6yx+QVsWDEn9/J6zxRYqdgcHWqrP3jPNxODF7Gf8
CyPGsKnkEeLVdQd3a3Fy6vjqFLKCt3Oy/VphUHpI7kuLQTS72+dttUI6Pl0IjqLBdkvpy7fNBx4p
a0ti9IacRg8reGo2fbPl9inbHkGY/YpHLC5Z0+PNRHLFd5tHM+b1Yqr8lYDZxf4zYLYBXQuetI6f
gB1WblWLfAz4OQGh2e3HtqxzaEm4izo37QPftXuUKUQ9GAjdO1b0Z16ANhU+NfuJxtL4xYVU7AmA
BvyHpphRDJC5yxm1vRzT2cAq5YUMDCeeMcGFNTO17kYG7fRWpyIagS/kmXRcFLmTO9hNMfdNz/6w
QZeNjipzj9ROInIx3kbC1yZ/3wS1laEt068cY6XWNEIKFCBsAKRv0wSIK43XoiycK5l++l9pfBOL
/3e9akUuO0raNc6P5zKn/keFMLTadohqIZDBvF5Wj+ZkXch1Qm98cobss3hDJ2KykMXkCSQoFxT5
RuDZq74B6g46tnw8aBnVaIJKhstL6dAaYXJ+P6HAZigGOC/1maZ88qYttGHrp+jmiSndi7OKGnyW
fCTTFNBdhmyvPzvg29V4rDxV/kAuPAtkFBLDrUky3hmNmzvuPnd+ojcZU4j9B5RUQG5OhJZk5pUn
TTEzAogZf5A9jnSG60pfNUJTdtRZkmQnAK4i5kIKU/q6tMPbJCVMvkdr7UN1t4JtnQ1riRicldzc
gVkHNJcfr1420Y39UAOBVj8ct5vqlw1eLU9yEWjELq4sEiV7fVvPqM6K9rKmJ/HYbPr9Vjc6PDGo
QP0wxxkcuVse/+iPhgz7o+qYP48QJxuWJQButP8CM3IHgOPQGx5/vQfnlwL5qHt+S0X6lFlvOYeR
1fVHmBvm8hoZiVJb9jxWz7ZCEmfyWoqR3WLjMOrD7F7gGfV2UJP1FvXrSSgi2PvLUt2HMalNHbYF
eKKfUhSJQ4Csi+YBQt+TagZklPNTCD4QuD640NPS9AcwIWg4jYnG3Zq1WWpocw1yBxzKJFWhHLxW
E8agQZxLKpbojbK0X0Yxhdeh26UObmNurYOhGLR5ksEU2bSdh/cPk9hjEAqurdxLm5xl4vuq92R8
VIBkXPcr9OfH9ApD+53UE7Dot5w8uXuviBy69u4uTuUtI7idwNXo0WpW5r/EAZhd6wPvwUIxkRYx
Ofwm+O+94PHmkcBP8tZKxhGUTZ+s//50aUiXvG3nV/cyStafm5xF8c6f9fAdWXMW7Gv06mTv1rNB
9c8UTxzPxIyDeOmRok46SzvYC2C2II5r2IXs8MQ7j/wp5XAuy+ckDgSL1wExjIt1yP56zHNF03UR
yU/TZXK8SvsAH/1RzfIqzhM3tS3H5nGBp0lasbiI+v+wrYfRBOsy9u2iqZ2dZDiBVtuZwf6h4yu+
EET84kXkvj2RD6mfvzUzzRLb3yY2gsRUosOCegJ9k+7oORH6/fkLDFKYTIckmSa+7ywHctxbtbDS
DJ1NT9KK/IwIxhR3smTy/86MrGJDzamU0U9K/Hn8OwzAk4uenWIZJClyah6TOYoRPQlrTfdEQmR1
kq1T7IUu926TxXUf24CEKbU40FgaEEApjOy870ZijLaXo9YNlsi/3eI2DKOvqsX+HZE8TXnkymOz
PFauWmZWjRfAgejiv2qMfi41cOuhr3PK7Jp8Kc7PiY5/JBJAcnEWXf8ixsPg4LUDM8D/T0WivXmw
xaKpPYHsWNASZaEPFmfPP0DsE1AjnWE2DzR5YH1XZR/wa9vviRXboi4ji3dlB1PcU+nXFTw3jszk
7NDNslMNgVguxc6YGZHGo7Y6IOvctB8ld1MlPQo4qWFVhV1QUk5UmDYBCQE7DybrQpbW0X+HGo43
fGYhINDJWpsX5zU+lZn2P3EEfkTDmkDzg/oFtFICvJvKsQqkH9ojlksmy7+kwtXt+5fN6WyzRd3b
zS9SViOv2a2P6Cl0H47XWfyQaO6J3kqxi89uo+0w5oPsx9jWHOiQQcs69/NEXCobUIYmoTxtU7O5
I8nFa7QPEi1Cvs0P8q1IJz+BZZxB/gJCgQgGxc4jvHv2J/XnFXPK9sIA0rGTAlTtp28Xc7OAtBFw
woj+udJP32v9elocwS5/nlErFLjVBgk/bKea9mEpZrc6gBA/PCobdJnoxS0bej1Oo5TL46gu2IBC
VIr4eaRJgYohbhbj0E5lLqzZx1LFaL0aEaZTZZZUQ6xxoI+wc99UUFNeAXN3Di51wDJRMINFklqv
t+7JLuVEUaqRcuc9AyX9AI5cb2QKBLV+joz/Dl84vXC0mOGMWCJNvFfEpd7f4cWHwf5LDZLSiyk1
3Zln3LWQI7WY3Guu3EVNLMG8uSYO4cPyeBPv/SodYcMZNEAPlBQK1h3de+iHXJjb2tgVJDjea5Sl
joT9ivmgW6H16gw4B4qf1kKc2elNYDsfEr7YXaENfPr4IGnG9znlTSczAKiH/qNauXI+rlxeZSRs
liF3rIL3nOkp8SzDwi8MlPjjtd5IQeCphC0MvPswUS0zHb1AMWJBt+vp+0+Hir0Kk99o0XWXBUIT
w7MRZ32E3OlxWsnPM0w0sTP5V+1ArPFXgCgsS6UhZrexMWV8Ba4ChbUtjvtY+pel8FGHhybxVtEx
tpnbBtk1yL3qAQkf1hCRiNApwSmq4aKzvrRXMX6YWBMIo/4tQDKvyjd3g8h7ZOagZFNSjF1UXTCp
f1LoMXE8pn1mMsfTSI65n25QrtCh/bEVzlQayIOzrhDQmBUrtvLuwquWmz/NvsVCDXh8guz89oog
/oQrmSShuCidAGWedfrurGq5FeyWLlWtsT0lUq2AD0lk96ClkpqHgFISBDAPoAPsfbadhLT2+AEf
GHkx5pC95P1jpRGIJKrr15it9lQsXuEEjhPJBfIFDKIFzLQcOMoweGAQc+XG/CMhZVzKYu1o6DLZ
RhBAlCl96+UxHNpBaHEsUyZzJu/f52CmqHcuC4n/rEqV257G9SCf9wFr9SPUkuGPiRDXBwsbGrFy
PJZJlxzwa52b5vofX+rJN3+mh8pmahr+gjTP56WJDBgvbfvsq+ylqb4zF9uR6ijT8luuN2M6zS5k
NkMAmYHcKkFY7T5i1c45mKQcEIJq/7F5uiDUxHKSJHbYnXzvhZ+4xHpFXtTRFJbPL64rPfATjYgw
s3Qz1c+JZKqOnVrAmbtzYB/prGmqhVIZdqHA0O64NeooyLg03Zgj/P2C38Z5Cou294nBFocKFDor
45sTVMxFjBonwwqyw+pc7mUSw5IXj+IEncnlRWwCXL29w9GKOYFKixja4ihcg5KyjGGhEzq9UTNt
yzNZvm5Z5DgjGmQJIlbLPMSsySoTawP4//u771FdQOWYqNGJOdMIKfWBC9Jpkp5GFH9XeLspGvbB
8CEnJsSj10xgCPKf+mB70EyvgTGxABT7YqX6P0iKOonOkrODqCQQYJ2VJh7EHiJQY60LRTCmkuya
Rk0lC5kQFhZutZQbwapLFmds1vP0EvOxfbx/0u8KsCVFbHJCgX9dTH01TeTwgyGNSBvtq+Qd+tLB
ERcGcIV7D6dUsd+E62F4W3RGf9hDCmLg3lGyMSoZnjevS1jD0lBcANZU1lMi0NNzEeRVgif6eXJi
Kqa50gECYv/NUMSV668P6nJJBIdUF9X+HtIW6QBS7oTEkOKs6cAHBSb9Xcx9VkXxRq2u53swFAow
SlCaC69E8TLCfbvYkK6ciMMlqVSTssrV8lea/QX9I6SbsM1MiPXI8vd/bB7D6qipE/n5i0lPHmMW
JtOqmCnD2FVyUV9YQ5eVSpsVwJ2JhFl081vvsKYTgoKUv+tjvu1OyjvILk60zJvrYnBeuJgTC/Ry
ZAcyap5x+i2NV7WzY7WKTCW22wtFWGG78WKg8YC+La43tjC4rAb5iK8fglW3/z21ZgrwoBL+cUhz
bVv1gEKzNNy9DvaQFSOUr5DHdTySKMPq9CfIKjZVSmp4d5QyCsTOPJC52uPMd3UYLJ6lY+T0dN5Z
iAA7kR15HOs/2hjD3kqmSsuQ02iaW2qcRtXd8ZJkCWT0CrdZcKbSR/hkHgPcQVdtLxEuMdxtiI9m
1VpX0cQOmAsldXKLaG22r5LraeAqhYsxSDKWqyDQIfHcDpo2XUgROuGW30gJzLrjpzHYhUmwq8An
4+3hI0nYQMl0nIxaWuTwZlznKTmUGozLlod//EOEnrhb2va7JYL87aFMVfMkYrRmliMtfQRuLUMh
X810vo8dE5NhOHmnhU/1sI3d5hfrd/I4zu2LPZnBj+wQ3zVzl6sfGv09/CEyhXK5ccKIjj0PWfi9
IGF5ey+HR4DFIOsVdq6cb0FFwKKy4tYdefiXiToET7cztMzTKr7QBxUFO7EZr/uNxfvHtGX5a8o0
amyOJuWv+KwLLK43+uR+L4FxQaq4N1XSh3AkSgBbCs5wnsI2tZvnoTqS//vA/K6b6efK6PtWrNGV
QBPI78qs2kU29QSW2+llJgUv9TdpRbKIpk8PSzeMjFezSN776rEDlgIL2kdtqqwE/OkUON1rpwr4
igsc0AHA/5PFnWjyXE28YCXC4U74vPe9iSwFgdB6Hi3FppKjaxKrhir0NX6FHTNan6D8M9HpkfHN
dsBOUzXrEmzRg2wrWyY1pib1wGFJCa2rXq/MSYk7jNxS00FPpMR/wMlDLbTidgWlg+Vg6G5zZYR+
M/8wLl+uFvCs2esH5tqQxYjXWiM+Psokakm9z3XUmZZWYZO+/vfkOuEoq0Lif0PjL9vKlu232X0O
c9S9UwrnhuhpACRMgfTCzBUEbw5tR8sooqPxvt8/ksCyrBXVg9eJRrfg9NoAOQ5T/ZU11ugEvqAO
RUdAzrPAW2DtGGOyVYGVQxLMKUhm0c5YEC2hKWUqoNknR+HBi1DcHdddC5FMLygQAVw0PcnyJGjQ
sOckl6bXAJmDEyRkzL/8zmynjpj/TchgJKqR0Sdl29oMDepoeBJiG4ufyyoGV9aJZYY2aVpvZUr+
b+nN1pWEiSX9ZokuBtYww1harfJkSVItDM5gDkkaNMHkLYW8s7+c3BopeMieDIjyBptBOhERfflC
nXPB6kqC6Cbu2kuTB8zRT5oBcPtkTEq2lHSRqkt9Woxikp8V/l9fo2QA6ZnVH6scM0tsSNy9n2AW
dgsk8YVuD3XBx9Y0F/zKSzYZ8wqNiB2g6/shzE3HxQja/UEpzllTZB+pPHMtF3m0Bi4NOhJ/jxMt
lBOTEqzO1NlMaCoZ/2G5mPjq2rrJPwGZf+uvKARQtZiOC96KTMUVgM43F/g2SkVahFIuLnN3NczE
6fmCRt7BfIrtaqRuFEKW9HK4Y2d5eGVWKaQLM/T1lLJwFe3lJiQWn2ZoOKpGxdLuNszjBZW2nxa5
6lD79zk7RYD33+BeQ9fo+T8jyO5waga7lnpsVK0HHv8JAyNZQEpf9iKAyDxoOQVOtT7iCq5XyOY8
eXMO6qRpTQMOkqsRzWj2jx1pJzBH2gO8pJR1xoJzKXH8MsBBDky1CSGabYr6CemnhYjyDZbCIN6H
q+SqQJ0krdktx6kBepoOrI444X8AR6g9uU7/qWRatOUC9NYOhdbJiySVIGynOyCl8Im7oMRpWZvi
h1MY/IAVnKLthfarzu7felzzhvUXid1eKvD5qP2BtAkxih0KfxaPVOtJ+NRIoN2M6JcV/TgOz4Vq
4ujHyB3RtSfEi8R+D0INwMpee3SZjEIGFRZe8pYyjj/qL2++qmSbyUKn2/1UhhA3Xu0ccikOsPJL
09uoiPYqF3+1yHAUm6gqOWrOYALp9R0tnN9RqXD3HbYZ1e6hPMV8GetEfxwXOGbpJj0tUhlNn/Uf
DRNLlkuP+1IoU2ap02bAEGOAlAsVQkTv8jafZ7WlEt6s8dZVU5876L2uwAquGocXc0oTJvDbs+Ik
3XLwDi8UsEkrpqpRQ/GbodRnm5aFUvrIH8imjf8AaPrrRh63P1b6fZb8yFgoVg9dNW3+CxABUbBs
Hrc15x+bjXmt7YXlnah86MyzgsUGT65mBPSKOne54Vg9260tKwEP/kRM7FGESiQqRR1GlFEsLexT
02nQBujFH2q8hnBfjKo592aeitPGR/f7Ls1HLWZdF4ByHP+yKYR3frbnx9iCuIpaDbrOGYnzT8hZ
w301i4c8o/HouK72YBgmWjEeX/sZQLIucNMjJqyZV53siekF5Dy3nVfD9KNYswX9SagxD7UpB4Nj
m2zE0zJI7cjTQaW6/EdZmhcXYhoQiqzfWh0WbmdMICDgHzaY4q1AZ4OVm9nZ4i6ICJakkSjRi5Jd
JjrDHO/FlaMBYNMxQ1hKIPLJan0dz3s+hnYVqXcypGH0BILbeKq4cnMExP7cyYvOEc3OirItyrO/
BRKB0uBEuzpL0y3mkI1ASNyMUxNxRmA2t13s38hI6IYqrmTVDJ8h09qvjxuG0TM55qLBXxGE5FLN
oGsSZVVcvEh8NHfNJn3YYZq6JIfRBav3EZ54P1R6qCc4pqP8DrYcuP3/koTWCb12YW7EjT+T9FLE
yVakOlg7q/xTMq1JxvJ/NMKPY11DHPA0c34XERqGjyGY6T/g01+mT+Vm9E5H172MryE8snx7B8WD
Bz5CDWyJnIuu6MbeZ3WcPpgS2ECRxzt6zKRJ5FVc5nJJWHluQG7LLequ4h0jvV5dFBbpwqhr62mP
5tybz7qkFDjn1bzeuR83uYPk0Wy5BHbDt4uOBGZQlhxjjOC7itYtzr2tGTpDputvOwHjIq+dh1XF
nMjK9TRV3oF4aL1hFwLkc7ha1xtDyxQXM1WWL4qZViIM/aQi7Ux0WOHmhx6K98nSvAPZjALTZ/TL
109QSAKL3ShItT/Xg0NOfhCqg1bJZsgT5s0yp94ciRTGSOkmQsRaM2J8732ubspxr3e8PPTQOpyN
kp+hS5OQZ304F/nI6xQ/rbl7wyj0R4gQgvwn1ZMOdlVf8tY9tC7Igto9ubm7D4FF69CxckprNMaw
0QpyMc7QB+0H02+59ptMOsVoV+ect28Ut1W1R8r6OVkwv+nTJPIkH6Ei8X2Bc/cofsuV/wRexAnN
VCDtOg7+COFjh729XQI6SnQN4QxPHe4wRnq2As19Aw9QCPLWvAvGRAWeUsZq6fHOucbJvpygM7M0
jsL0vE3CcUBrWa/uPaWtxphJbvN0DWvsbM0UZHU//aOliSrz0K2f+KrUUbrByrDOjJRsyuFIr/Nc
wK1KNjRIqNtpWOuKXSPPLcGQg5J1hUu9BujqjQWb134Pu86d8JRTIQ/URLQm0vWG05FiBsEbmLiy
4RasjbWh0IJKKjKdU1LsP6upZwvgJpSN2bnvFVEL1ui1LqWnAyGI9BU3rZ7bDqalwWQ9WSsnopXk
/rlyVCCaGqWYBQwdSc96rZZHYnQAh71mMD+iGneEKca90tGs/pCfI4x+c6324yf+tPha1kFpFMR6
ZQ/IGN5riwikXVXffULG+aU9mWdI9Yido/8l48Rolu4saTu+sCFYGse1EyJbre4zg9Sn2A3ythvC
iYrJOmwrmir147HBabSHLuOGq7yWpbwUaXg/nGExiVAJRXVzRpH2YOumM3Zz0qhydPAbWO0qAbtG
N3GNWFaG7fNA71aKrqoQChK0nRCbnpc62NBRZLjiEedHYKrZ/svlwHMfLkDHwu4x8J9oy2bTayJb
S/cAZRcuLRxIYf1goG9aPFBvifN4uSUkH0dyNZdjip13HOTJmuNKzz4TBzIpGK83QQTBO3H2aClz
3qTh1QmhzqqNANEUWrZIVMBQEQKLmQwYUl4d5HhBo5c2IZlQjYF6yn5gi3Wf8Bvoodn1g1J9dC3m
03fBYqGC9YnWgsaSHeceOE/5qIspTCy0Uwwpuf1oT64rS2UDV0u2SMrC0+wwK1mErkiSe8jEfbkV
hfNEOoFna8ukAxVZUGoHQ/uQxrE57XYmGy2RNy1FhhDR9BNaUe7CXCBlLrbtH+S1poyNTuU1prVI
oEZJcVoW0XdDUHgE7FFjbC9k+5L/U46AG2hDKVRW0P1WWLk1LJMHXNsuE/NVOtprAgpBrMRGIl9e
tLQ/SRv0apL0wfmT/r4Fp86QEBY4CqHa150dEKUXECy7v4AF6bfScoRUExA06obLMglR96rsW60b
lRUZ8hMmHClkrjZnoUgsJzdRwXyLsG9zJpBk2NCUyzJGoHniXHv7oZWfoQWHHl77es366Wz4U8rq
gmek0VoCnNRUKpA9jV7Ry/H+gWQDNc6dY8xX5gSfVA6YKu+aMUWJwzJclLb9+/mE4jVWHhn58Mty
qpW0uo/ORO7rrxayJ2Wy/NsPQEHh+esqzQURy4p5VddZzknJLu+3hQhvYeC//GVw2JREfSWvMo2H
XSzCZ0MaIA1LYsis8G5c9ZScMgosDavn5Bk3IncPB28+pGUR949e8FLzAgITcVuFqhO3PK+0Bg5R
gxzmxbVFP+45qrr37SkPgRPMP1FT7YAHUbF0udpP8bIEyNNku8ywQnYQ52OSC0ViLeV7mAndB+VW
EDvKpv4nCX1z3vi/XMLS5XZJ2J1ESP4XuC1RDa6zIWAouKtMVsQbCFTlTxLYgIwbSwWhN57h1fGa
U6W+VsxWI2qT6DjBkb9HMxI9HbflqfDO7Pq47+ocODdXVvFJmOpsR78yeLYGxY2lOxM72DeOOvz/
estUaDH0vgKTYL7UBa7ZJrRWs51uskSknoZ6xAsvJnsUYnNJrvEY7+AheZREnMZ/vLq9bKKidcRy
qzNR11hH1qYN1+ZUVGEZgB8CdM7k+8vGHLgBzvYl1O6Lf8OpHzp3SBTEPrqFRmGlbmcJpCsL/5it
O0j7N/D+uDMCUkYc3JfkdHEa0SKe+3ewhlFkehY+i9+FgV7nUZi4dn58UU2azKxywuxLW46gkhBu
Y/FTxb7+uurtWoW/Mbjhbw445dOxDm16otuLHWMeL9jqFhc+6GylsfiZd7hLQuGJczzNqktHTFOl
iVmgU4qAKaExA2rDhdrZx80UUOwbWRwg/43YchuYhfcxgjRxxkr1tYMuUum1TqCwYYwPD/ceULaz
TA6FveZalvqxDM6vtwlGii/+8NGpkzfzx0EMyZHUX6w9ewTJieRBPwJYY3CkIKSQ8n0bwav9wL58
TnYWtb2qIQwmNp6zdmUVZlPf43muQ4bM4At8gDYUDmiCRUBnE7jHB1UvLvoVz+3Bo6Cqfos3rrvZ
ml7CSSRHQuILbzj/CEZzS/GL5X6nbDwj1Crhyd7Jr/kkb+HLKun7PNcn/hjdDDxZugcpr23grYMl
+r6+6tLNo9zpi8huuCKbRw3VUkx3faUHCdAaiB+cqNIZjYeJhPdhwq9EdIdho89POHvilTLLLHAU
Ll0JiYZCh2zLBVA6yCDeZm2JVja/hzM9KtvMPfVsatOLDr8QnvlwfzYsJQniyXZC0VEV9ZnzhxEp
Fn7EBSyM4p8JAqZNDSTCWsnAwVs0fOkbW84RVoO3iB0ZLzfaf2ZnA3+iItQekTeJX+QH37OZJY3V
4d0mN+9bDdjpaEAprlIiBBjYixBo57PZzbxoVdYJ0frD6UOw09XCNWcq7ITADKaUuAX9b5i/pREQ
Wq9+3WDMJHDs29UZf6Ygx5LevZg3+wtMS553XDs8k+gwY6uUcWKjekTmsI/IAOlc5HF1KpXzuz+J
db7or0kvYihz8Pz7y8O33V4l7L4yG4Wfot+6FZ4f4zsSQkv8THQ3ddcq+udT6Jpb9FNc7bVFJn0d
ljz6/UjlgSbQSXYKwfaLN3PSO7JvjdQUbOkVZZ6WjubqLMkWEooiaPuO27zzB1JUuYe4pSzFYdD9
gaX++0JDh654A5EWrtGf6NbkU9WOKvY4TpfjDxV/j5d6U5SaKv5IDvYKwqkCa0lboDp8y5HNuD3t
S4NE6mB6XRaqN/ePGoqPtlZmRFn4xOUxzK2Y2WJ3X2dc+dmynDxLJUP4ch1W44bBbiI9EyNZas4L
2yLdFR61iQycRDjXgkhetlWup5+grvt/e1lKGCFvHvSmnoX7s7HaqFoAxSJZypnbjcHKGb7dN8xk
mPvp7JyKt7+1QT3iZQkHM7usQ9YcRz5q9Yh8U/k/4pm+RXy1kCvLITCrxCpkDQxb5wgWxYeuWjqF
L6Yjx6sNYvjDtV80yNmMElkGJQOltQrEe1DoqsPc/jMNjafpzuaGIuwh2Yfg7wC95RQ5aa0tt/ID
/HGVX13Rx66cGnod5EHu5cCKFy5OUms7Dn2djXvvcVDrTExvjQmS1y3RUltSsb+ZCIR/x2KBbxEG
6pAwjvb+IlRV/piwFhvhS1PEX2qplDoJtpV2yOllm5CCAlq/5o/j/O0wTsgL4IdYmPjrHulzJ1yr
RYOCFhOy3vY9nXI2qD2T+I6eeU6gJtQg5k6JCzeQWgK7lwPeGbzu75zV4M4J6tkxYkw6GwyddmDE
TjATxTOJ012/9GCLjVex22sLSYIYfO91QHMfUrjM171WfxeZYQYqPNqKICe1UYcRc31AUn0BPRM/
gXCrA8T6RV9800hv/iGfTrlQXjoK/EvBCFPLjQ+XkLVQeCzYU3UI87klqLTWq8JZ7VuyGqKo3Jvd
LFBp9NakqAaxtVjSu1pV2Ed48l3HnWkcZN+0vZiJMdmaTUfQooFM1gJ8t57mzwGtDZtusOavv40R
eEHdvoaDOZmO0IuHqtbQ753+pIaAheH+pTG4y5W5zbeLPGRv2fOjwRmIZiDC7KhmUo9g6WiQNupi
Vd0HJga2XW5B17ohqO+5qhGTYMPO1MxccX/TyqBXXsxVsTtlk4LRRWwtB1jPZGiNbq09db+jcnOf
9r+x0ZPGoC3yzf8KsA5Q4ARHRGWZOnOdpj2GMrSr2d9futCgJ/CZ7JRJel0fBpRhj1Wmw6Jn6Xa+
zO31jDu3JJJpRor82AwFgGjiJpjMhmwaqDToJRgQbXvwlI7TJ9HNCeYhNCP5eWtChNk6Hbep6lOs
rEb2M1ZcmYChdLJwQ3JoV4pQrWpO9xxl6odyMqxz5deaj4LlW/saXEq4f98XNg4xY8Umtw/hziDI
Js06BqZmogqUlTdEh3HhDJg8FQBBPdlCpXLSIfGpAnA4M/zc+LzJRT/Mnbdo95At5cKsBnDzdGWo
QlTAYfE82zzHQwmkfoGqPvj5LlKfGz7uGWlen29Beavtwn0s6/9x4yS6sMFfurwU6e1sekFrbuxm
LoCXPH2jSi/VLTKWMkh4B+7GWMl0pUpSL5+97kWWlADOAxT7uOiNdpwAVpZ92HVimRbZtCweHrv9
zAl5V0WsjSIh468nPOMMlsxmZLwZCwvGOuj3rd1Fh2x+plds9/IUcUJvhp2jiy1Shp7KrZm+d1bd
TjIXJ0Xiz5NjHGTzBKpJMmMwCJPY6uTQqJ+Y578SAQdh5llNjYi3JpUOS6tB/y3+eVBH9fEvy8hM
ph/FiRVocENs6YDPsu4+QPv2MfLsu1oSh6iz9M2gZCdqh7tSKawn9sS7G3JqvhAdSiA/tdFYoMqf
po00QtLDrCcZHcN+xnlK/zcD13ykMxToduL7DWwoTL6qFp2lsDA13ojJmkpbmmctCWVTFGLXTbJM
VeHzqXlUoKtXgj/57zX8LvttFBdcAavzFYLPlTizSp4KbXYdkNbOfPuo9jiErnZ80kwqurhk1d3J
DKJobt5xyHblvke7URD6tHXIpfIbYzCS+P50omZXDd482cfLQ7HEyciJTOICYjbdEg5GSuXVhFN7
HCTu4vLqKYvoAzCUpeam/EvXv67Bp8xxiQO1yKQo3/OqhJovCfT8CRgiJtK5ffr4NHbgAfv+grB2
3Lt1QPCMrzCZygodISRhZW6UKUODA5zSXrBfcJGkc5i8BKHs6id1kr6vv+clgQNhEs1kER5OIdm0
EP5iKYGwZsM1RtR9Uink4FAMFwuKDBJe5a0lyDTecYvImc/UXASrgdlT+HsMUwPJCNloIzjVEpM9
omsRWwXNf7YZ/NszM/29HgEinaPS2eTbDPlxd1g4p3NLf+VO7MG/aWzh2xrG2VnIlCIQwL9+5AWn
SLaSIi7fmPxiLiVTe3840JYEhBv+WR1AW4JS38/xZlXVZtVwkjVtvbfYwHis8pVdsMOO4OMv96VC
Eie9qSg+NcshhsE9X2B85NN829FAPu/8t25hA1QtT4iBgzmRASbOwXZPqW1zmNoNNPwTmk/ykZFH
VNKQ/DwyLxQeZMay6CEt6oFgWNILebLaU5uk46WUNwLV2SfftVF1vpd4mjQpe0zcJFWHvUs1wkUY
twhSUgOHV6jJbKKLKUn8G7oivRZINa/XHlPkU7sRvvGQpP4i4r4+6sXcE+HRU/exo/BfYGyg5yXQ
KV45uNZ2Qp17qqN0/yEDssaMhFECkpW9aOTe122Dv/0InKn3+zjS4uJiI1x46Q9KZC74zuTq6awj
FUEBujXwwr5ictwaBtBVuB5cS9tsug2wsClKOsEaPjPvkGi1KvHvc2QDbfirwuVNmXmLKWYC1aQP
BDjUykV22wHgWlD2ObePxnjyMIOdt1pxkEnPSmv0+MONOXXgcoE/k01zt0w3oZ/NzGNVlrnJRm8I
qpdH/6RFMjVAm8c/c9rzovbe9M2d8oKa3x9cd9etUmHb81XAPvTEOv0/aG1Iu9gKJPRIdFnTUcbX
0OfxwVMNsEkdTo8SXVuHRD84XIOqPurlgoqvm305lTECTLrjCE2dpXqTIShPSDIn/qQdFboJLv0y
Ycdv+v3/RZxpsMeq4oH4y/14V4uIY4RLD3kbzxG2AEssYTM3nhpheyvkOawDJQRAhczjKNERsVi+
ODKnaIkSol0ZGkBrz5SFbYzrkbueXyF/0/d4EclRGmDezdXB2+pgMWb8UzRC2yFMyHbITOD4Noxp
XBPCIARPtZpT2t65wGz7QZVzIthEoVXAt4eO/Q6NcLiCsneSt3WEF5M1/+gEXeZ2ywXA9ET2/0J+
AYT3g9KW/E1xW99Gl2ZExCkYR9o5Zg7KEHRmzeWadERzo9oRmLGOLMhkEowGFddImgDo/rGP012R
UhazBo6GJUk8vF4AmcxSpkO+jFWUbjPxlMiddxmG4tec+2hZpJJieJwLPFe1q9NNS7xwBpJS7gSU
bMHIurvSv204tnZlG94F3v2jIMXb+rdD0uRxaV6vNeLu/JnfEdPCdb75gZxGfW3Yq+RuJZANCKaI
Q24FVeWTc1aSJKKGDGYsMz2zH++7mlwC21PnFhhPDFMtO2batI0SLQWcIj2jkIbKwy5EcgkY980A
jWBGMu54X9Dq1c7GJldnlP1jro2bnhPklKQv08rrlwDEzP2BiqONWcQB4AWxRKS3d0T4PMWzd+uo
2TA9eL3qqM0fhWZdspkGuxrLxLCsupRycbSdyTVm/LYrPfN/5OSUmI8A4lT3KCfV2LjgnYhv7QkS
joThwz80LkggZBw+dDaDSn5Rcm79tVEHLlrmcqgqLobyaar6x0GvDNhRsZ1tOdOic7MV/pTirzPa
p4u32H84wxazYsHyUK5uSaPD+8q855NtxnOfhqwFrk87BYi5bS+IlPj1+/+D9mwPEs8qKMHetpkO
xThZ/Uhr4L2TNIGNdDj4TQdxGyw1VfI2xXaCQftn2qKkNFy0Pef6DKM/GYafBMTu6asBH0vA9HTg
NN8R+X2oPcP5tIn5fZsMzKHSfodIWA1/frH9Jy5d1RO76yPeTIHB+2nG/oVnV4zpa9qmAANXUE8O
XuoLbGtBWLavb6Z6hKNqP2CZ5wno7a5O1zO9iT0MP5H5aBhXrRf7u8VSv8s7sP32EeCvOflNOA8z
lL1jVB7lfWugkJR/2xTaYJoVsbKhs1vkK3b2rK8HFr7grYWzAR5lj+SF2TgP72Q+YDTOMcINmf3o
pJ5heNdMNLrU0q4sEiwzmw/+iD0V4jC03yaYCqgjyzxkR/GMGXL+X2GvSFTgAjd7sEr79mEfGD+8
tm/pDdNY+NQRh2U/rB4svXNjvfLAcsrBvPmgD/XKkk+ebQMJzK0Z1ijkhVvNIYJhp3cIF9DM3wsB
xIlsFhehK89ZPGz7VVCSzICjtxKLProhY6+XqfMzrx+Jf3Y/nEADvzzNy9Inj0Hc2d/2VhFxSK0C
okFiqhqnm4uGFACjre/Arnunk7Atsww3vLp/FnJAiZE7QCg9BgepEYmWc3lihCq0lk1Ua9EUPFRo
Pexk5fTl18mnUWF5D0K2tkxbXprE8x2NA8v4rNuVzlZKn+e1EvmPWdFeq2jKwXXh1A40YGHwJswP
oMBt0vtxaMoQTMGpVvPQ1TYjMRitHE1LGtvi2HFNdxPu756Zmtup72eugdiHz5V8KjgCHpU+PfI6
jzWL73PyZ2doeUIdtg0UbigpYQi4wMx771sAdyf6zYpuPV/rTzE9020s0KrluBYoj+xXkmyFhoye
8D+cJcqyV2dTAithTPCBZx3oj7x2CXbNeNq3E9N6cakkQ/CwtNbL60aVNEHtlm044G0yq/2SllBr
7Z2xkIRLdbnylQ64D0jCPAUuc5BcvsEdLM76fMQ8TaxrwnXwQZjdlErnaKKCK+tyCaEjA02o5pPR
Bn4FKqOwsfoSSmiAl2fo4/M8L1P2LuWXucXArH+eQUa5cbKiRKfELxMntwbfWoSis6slE/MWbaQ6
9JvHYPnCWit/NmI8NNmUoviDh+WjvNvAi/KIIk+JuRTjX814bBx/kJiTCLfDapL25nlKjVRBojbA
+OPtUDEf+w777BuTBx+/QWCE++8RSFvrWfbjaqCxr1Hs3DTtgYPCT0Y982NJvtgOrrM0S50hhRAN
/aD1bmu2qUEUjF/wD0xIGEu5Pqq1LCTKQWhJmLrIGmt6Q378Lmxkt5HzhuCLi4Qu280oWApifp1f
Q9Rqa8NVL2xG8Q4ynzDjanS+iuu7EkzwhqpkbjSPeoCIs44ZK2/QlHXTQZI3y2G6rB9iNJ+WnQVp
XAGUMGwbTenyXvEz5RVz5PaO9Utfhc/ELP76fqWenZFQ+Nq471eCIIoGU3bL/71iCishq3e5hhXZ
2DIoWA1P4mV2qHdGZ0UOZ9j7Pc8aYt0ikTs6eIayH2quOUvP9lFJDrDTImgul90q5resY/XjNofG
d/6N5mduUWpKm1er6stNOooQ5lzc8FgWK/Sj+Ep76VE+/OPzPBa4b9wPkiS8nwTq7W0D/vPPUMwE
YGtqhUj3iq9HtHg8lcq6V7OvICbwoVu7t86kZFVTqQLIR//fdRJhnlCtTp40NLmgmg49F0TXovel
jZP2uJ74/sM2or7Yccy8D1aiSllapiUKf6/kS1q36rNSM0/RhCrDA+mWB92QUPWCGTM8ft0c03GW
bbR03AjgBnuRnoYef8xToiqA5lhsO5TQHyQx137eMJICsWmd/arUcNBACG4fT/TMiazN0U3lWVrP
Fg4wkisIKYui0stecXrKIc6clU87nm2OhbFSh4ErROp2RBMttzRyIQbGgarJdJayqSeX5Aw0tr6s
Zti2dsrnPC6fgjuWh7/TBHTyzbz0L18jlujiFfcYoPEuIpRwfyI1iysp75jyiGRr13chfOna9TJ+
eXaomf/zvnplETWyVv3iLDi2JdQG1Y1VOVTW49Oor6soQGlO11H++n2Y6j4VWZziP+Tt7a8RixHd
xdnyp9i9kQLxv8DTcedFA9IPRLGXCfQlAonDSdlIA9O3GiFEFJ6pP2zmW8W2K/oRSDO1wVIzjYCB
GLnUsNYqYpMwQwMVBx2UsAqh+GX4OiHUqeVYkstmVi4N1ami+Q48b8+NIrwa4UK9d131GUIFtm5f
7JHpnCzOe67EAxpxXOF8HN76attYZxp3YDjdRUssO1UhP4RRce9XvcFm2bcZbD6aYQ+g600CcDGA
06d+BGWULlQQndyS3cOeZOLgXNkQln8QPrE4lsm+Bt3XyIQIzHk2T2cgzJK4jTDAisLuWxHJfFv1
GeqEjhSJfpxIA5SJTi/isGxqZid8TDz836NeH1uMCki2E29YDd8a7tjvhn0LFV29mk5lmsDFSpF7
qT8JKFADjtnqF43VabEThBaur/U0ffyZLs1DiBS45+txLO5MPeMLw4aLiWq+uMivHOdSRL+9xi+y
GlIse/3y/TiddChBSdinR+V24YBe5fO46A5qycuvuVQROHvKLiK5mu9I5mnOh8Esd5K0kfyIdm8g
h7fmZOZfURGvznRwpSC7DG/bkjxAs3PPN+Rvp7NuOD99yTVH2pzxGNYSN/OBoEfVSBa0mNdSXZtj
K5DAs1nQbVDFaaoUbb8enUl+5gkorCbABQ/xdrD5J+7pc3qu10K6NABog3AsM8mDKI4aJdCSBzKc
HkY1kkjSBrNw06pbqmcFOl6ifQracB0vNISuU1d2P3ef0i6XqZa+ul9aDywKOPbgrtuV92ulVIaP
z1ljd53zIfVRMDJgit4ROUfng8gqfQx6X66J4bRhpxvAwCkliT8fcp3rpy4kN8rwp4Zfp4+KumF9
6J6vO8Ju8470MrJ2aeptWzcDYuRiRFSTm2Z/D3Ufmpkk7b7E4GNaGUDAg65FsbtI7qUPJL0cBOKe
p+QMnjAE59ehGvtMxDYa+LIPezyxo40fRtSCXMdTvcERt08NDjh2YglZdSTXWYKZbNZ/ol6/pN43
BL93Ywi+7IXxw4XBeFwGryJTIkAZ1l4S2oj1Z60mdKwCooOGLNz19rVd7OzNZYQlf46th9cbTEXu
1/lRZH6Cb/b5CnRjxLpv1SXDYKp1Ne53bNIX/pjJRTG227dU3Qo5WNrX/yM+Y/1NdmatmvZ4jkpE
vz1wF968SnWCU1N0AO61K68IV/aP7tgAfMK/yJ/7WryU6NfIIRi7CuBqyqqw24wk/NFxCz2jTdkJ
OnMfKsYVNHE5h8iqmTXkvcNbD6RuRKPn+l2ioMoHv9/e3aRlFXBbLhSzeq4R6okuv0Qj+np498UK
lw4h/OhSF23Z8VZdSlgdVBUGGUMZhn1QNOcHzFfYCotXwR2BGUrZBwcZAMbLehBgvuk3xZrU4WYg
rafcEJ62IaO+MX+WG8N1vgvxR2sFGWbNrCTloXjfTWU47mjiOPRWojmrYMa5RXiNphQW/eDRuhRn
MzoskikUo1q6pifO+MrLWhp4UaRYmPC2AhZdxr9Wpcw2FNRmf/+SeIzWiUCoVG3Y1BjH6EPsWq2q
qU5xy9+S55CRu4qKAHXVw9WfV8bCXdKpUW3vY4hjSP269xNwFJ2G12QBECtMZllEJziUnKpf3rVT
HNQTegjCVAMoc9Z3T0TWIZegOKWD6KYhbEmsNU27mRAczrirLfQqmruzjIU3EKwibb624jPWjiv0
m3aa1yZhr40H9buQXYcFUUgiyAhwskuGP+Q89gLgG7832EYr1k/jPrEFkVsYaM4kwp7XVWTJpirC
8Vy7WD87SQmW/8zD+SF0WIfOimL7ib1KeUIYGopdm/zDk9Sm5vSvABaogoxKpEs+p+YUjN3Klmd8
HJUWDHRr7os75iAw+/L9lpuwbGtTPQSxwaOPOBOX0dnlCJTV+oeW42zycC0CaHh2cPVrkPMUKac/
/r2KQlxkz7hmyqb36Us5WPZlJIP0V7i51fWQSkPJNR9skGM+wd/IzedNTZjujFAFoJRS7fux/tlC
P3n4sQZ1HP7m4KiIIj8KijNgvipgjS1GJzfMwoGR0IjbA/gMzDZNKnFLQg1sSKPmgw/q/On9lczR
bUaCYWcBeX1Vgwxj0z/vCAXTybYtO8jZeVvhLfDPMsPh4b88DSmtxpNeG10MaEcGsnayxlKbMfg4
I8F/WTohUgVHvsldb5H1vLzz2l0S8zQnmFJiDhBOCp+2aAyp76pZ5iuJLHZ1Z480xhJHsjQinM6B
K3p9GXHuNdEFj4W/jL3wBHMvxTJvnrVM48P2e/evT2K5JTg5/nFOz0C+OrxoFsdupmizkRy35vZV
lipJcHhWFt98CEIa/qdtP7cFpXdKhsQViy97rFAUqablM7TjjS5U7BynAi9VOEfdT5seBEsyKt3/
MiLdFFlSvMtrdhko5eathJ1jUUuHujlJiOjD/NdzBWSFKzyWZUUG4uJY46cIZuwYSFXK0UYZuKL2
5akgjYCZzlOq/opiZYJQ9cfdg4KLEqKvW/6K1fgydJ4Jk9Fg1YCB3fGChgk4Cr1iAuhn7fmfyZe0
2ep8yxQFw+zHCID7Io8i9oP9h6gkK2gp0Gyz4xPWMh6pjJCJgCopZXK+xeCd66zJa8SjAWk51TsS
WzEb/IutfGW1KIJNO5Km5NPvhE6FHtxuE9pvoc5TJ3I2eKDpuzFsXcayQCQwoEa3WgBaxLaEjqDy
FOk4DevNO5+k6t9Oad+cnbCuyeurjuFDWyPqQ5szNEwliwG2cLZqS0f44OcIZe55iSroTGjolqUE
37kXqb43WHdydjZDI4pTdNgjvBKS6xLEpVaBFZVWhMNdRmXHM9NkCJRrq2UtzmFzB7qhtgps3oIi
DyZmXFrz3yT7iMUkHeBELs+3wnyTlsjvXj0VOMcJC6TlmPN8+QDKDNYxFvnkq98lG/6QzX7mKseA
+fOfvVHRVwIlpsmHG+TYZZMw/tgUv7BUCcb7VoML6tZXFazzVRfR1SYnYAon1o7jOqpnZHj71vv9
EBRHu2zzvRdC0bmydtwA3/molvbPA8Wsv+nhSZUHSJDXf06d00x/S/UESHMDVvOZp9RQBUcT09lv
Kqmbeih7K85m8AaLoQdfUSEzzU55M3meoA6sIOrIxXaaNm0nr79Oh3PzTrysqP/5mvWTrue28WSK
lLyW2qdaNrmn2I78bRXPMIFlOuu67F6K2TR4swt7mb3HHQyZJUg0nUzepMpEOBRIq1PiYYMehkud
jz0XR2aICMq0Ny4T9oF8qB4Ix1OfEOdwBA1wLUynVmj25nOWlU4t+OP9qB4dS+dcN5xv+dij58oV
XCRVSHp2CU6iMUTt7RU3/5Qo3+xejUb2jutmepgUHYrhSdVsfj07wLhvzr0rGx6ZI1L14mKGpek3
x+E7cJe6Dv1Zezs4/zvg8zZvB8Lf7sQeES/y5qO8pH8r/hwws7lC9kZEr8t4Rr2aEIqjklsiMgM7
Pt/BHveMWB4KagcOy0RvU3pG6WauJ8A0sn0B1UjpRQXY95UvEHGSZEdn0brSwMZ8gJxYh4dx+gP3
rNiR/gcPIzoyzqj7o10GzK1Utt8TuTD+BU8NEY8J28Q0U+XB3n17/AczmKbXczwf4kwnN4L/6FEq
6aIoe8iwKGMkVfYPlIkdit+dGVR+MiZM1k8j6IMSziiXuwoI1F0FxMHKs5RjuCeyFLMFvf4h4ERy
yNHdk1ZUyc9yijrq8UROo99/kjYji822MDQXt5U4cqASw4SmU+dlEBOtMGdn5O2exRy28d45jddx
M6eAxaJBbQWd2lAJMWxqAxXDimuRECOmU72CVeBhSnuKainoyY6icU4TmApSfGktLwtzDxqVETNb
3uama6GmJx6orvy6AMRhgW5/Sj8ApUeKktSi3+ch/eHmedl1p7hE5Q0BiGnBaT3+bv5CR1dWit+3
AzrMWA4Za6QdvfjbKsC5U/k8Kyh3cT/4wKejHmdaYMqsnQOMcTalNQzSofnfm0dh1VrEJXwF3VjG
uQRAhXEUlJPKc6d+0MnVK+CvZ/R3+goj0nnlldhx9AjdGI0iGRINL+b6wkEZVcfDrcXsaL3WTPC7
ksFmbSln7oe+RuFA1NqlFmo6SMZYmfsIEsCw8lxzAr0Wvdkrq2qW8W2S2MQlF7F7CxvQnqCWJHiG
PblAir2Clt3YV/VJDo4rAnEdxoJklHen/NUfXondrFmouv2RcV3Sz8TjyRtwWR9SVsnW9sAv40Tt
p2ZMAdTWk+kPqqvXFs8aiMBPNOLeGtYOpbHlrkvqvGgiTEWPfU0yS2BoNZFdHsZJUFFvpXArw7Vg
iv0oQMgwRWttRToAq7rfO36qH9WAc9t5AwVN97nZw93yEDBnfvuqhT2eurc1f1RPGTUH0b8vbMxR
Ovv1p7YPdhYE0FGBefO8iiwF/xZfvNK4I/BDtqjSbcTztI+vBqWH5amjzfCrFK0I39hO+aqWizyh
xsdErlZHtY51VeMygt6o5fivvm5aG4E2je9dhPhcTPX8wxA7kkS+/2eSa6ub/wvZnqcWZCNgDASg
Rm1CTTBSbRI23oquT1lyYxYa8x8ofsF1v7BmI4wjRZ0S7HkuWfS8s0d8nlfrki/iOFtpWTWpryIf
Nl8FpxfJgzkUQUaZvnoK33Gl73FhPnQ+Da81mjvQthSI3SLnwgqeQSim8zjZ1cyzLv/EXOwShow0
KO/JDf1WHw4xupEsDkmV34c8TV6bxnvmimDPr1/UcZl9Yhj60rBhsMqgHeFFPZJQWh3RnHMp4HEd
RWXOFSg4HiHqF5NeowQz8StGDhLxVVeT9gkK0A0yDnOdLtPG/IRvn+9JYKVpisJUgRxacSvpEl+5
XYPbzqw6Sq5Sp7hQVydYQeixbU56lEBM2smylniAhmiHyXPhUXeJTaHPgG82OsIuGw85Kkq+Xaxv
YVSch18AzcFx5dPCSwdfR6uuKYsd1VKaBi+DOXuPEbpmkUsxihzlVcHA5l4Y7xZfgndkUp0VBWcl
j3LR0ZedfDjJ81lj1/0sziBwjuwFaqeSy0GED5AXZtiC3Mchxa3lhArem7KqHuMBZ5rYTimoGUub
fGT3P2YECMgmzH+IK3PIIgJLaQxU/0Vf3Ate663h1mckUoezKELcGtuzNtp+rRHapvxIVAEEWaGR
dlFH7w5ck2v7HFHt08+0tkVHK/Uxq3r0K2Kod26it27IW/V4X8AsfXrHYP+4b9I9XClHid7tf2AD
pyL7OtU38qM/EHk1tEDnpoRXhUkTpyls5F9qwnyeSeJrVUA3tmk1dtxeibAa8HdWtNq1+XkvLzvp
eiU0s/wnqEBhR4DPMsMKKJEHf1ef0TSDmIBuvDxXyug300wZ00s8nVjXjGnGGxSc5XsoNOtrQFvF
F+WThbc/rK9Dtt4ISfNYDg1WGTqZk7Zq0hRAZc/LbRrL22CVYvG9jjifvqt3kJTd1facL5c1tEwp
4Hgs8fztLQDtaszf16dCkG8qzcsxVF9AhMm1lpWorbwBJ7s11xmC9igKvMTAB3bWPuQVmLAk95D+
+e5wAXx2oikR7/lqUup2j6WCHGX0GBBLHKcoYZXymtB7F1Al+M6ptk3ypHwgBO1aqtEexSCIPK88
giidXkkq6ZBHniFDj8aO8TzwOji6soEdE35mHOrfcS211JNuLKCD2I4XZzJ2jMEvZA/MbovoxDam
IossQ+5a9Bl5/d+hXsXkAKkXLWh2cmk3rZDBM3BFsSkKLgls0EWdmCtSTNMxsvgwFOk/TR5LLmB0
JKhodtJt1U/6lDXX6NH2jFnJRJOKdaCtZPJRUwEWKtOseh3Rhxqg69xAo6qIFFt+6QIW4P40tT5a
DjDpjxv/IPtYCCdeWpjgwKAWwsyA/sX6hN0yYkyBCHbp+4nTR49rEmuGh71wp9JGJGixzlUlJ6wX
8vXzNcIYpjZLiSJiLH21NReHoR0a0W/XcamY+y/4bkEbCjzHHbOeOz4GHz1uZ2HtQnWNYJUvRcyb
ijgOU5vrE6QvmFBtt0h1uACDxAEMWDgWsCUxkBwDpmO5O+HQbkaERluzR3LHkXFj8nd/YKHzNdF4
3xBN3PhDmmHMt5s4DPOnIBlwvj1kwWGtu735wdwm+3r663hlcWGFbVPda9jLT4uRjnCBGb8YGYW4
ol101HOatoPIRwuFhUhv4kwPByN9Kxbc7btAz9WpdCll1LLaWWSkW7YHcBBC0+WYG47gu3WHvKxt
fMTDfsyGQdgQnvbGq3fWjGTep2i5Fe2tz0yTvkA95dlq/nOUv5dQ+04zZErGFzcgTDAXzmFhAeBl
fl25UQWuzNK60WoEKRUmMMybFSa31Nzd7tPTpjQrZfncNvlDOhKKaj1hfPusVufYYkbvRuZqHiPv
njc2BK30dlzIS1fRB7uEqq/DX1J5YibTlGyGL5cJqdLJDW9UE+br/UTsvKNotsmkCwDYxmPFkwdL
8zsD2smE2btzB/fwCWCuDMVz2AKIlXpXoWF5cjLhf0tDV4P/RDNTeEzKig/hZrG9eJFwbHX4oD9u
DTxtWMCxAV73rQ4jMsQzLMZWsLH4iOCWhE3SkITlbKHfCS77MVxL+jIdY8BTkOZaa9KZ9xZiA3sz
jL6zHw9dZJ1zAFgGa8mE4WqW6aW2RuoIFTJKjBIG/lGGNh6GjD2u70KINu3Vejeza5u7KQAEST75
d6aCqiOmwU+ELlEm3Qp1PRcLlatgdlbIOeGovcHoPeZHFc4+oqwK3tnc/EZhwP3dXkWtUCAz6dCC
2pG08sJgdWIgCTjBu7KWW62iUgpGGfIzCPBdEW7exc5Knm6b2jB1pRw7aKEV4pphL+XVerrlRzOC
MqdPNuy9KMdXtLQF7zjrfuhEDm9ghdbja0hGiXqN8YXeMvUGzLOmgkIaf4bxdPa1HTlEicQwjLrC
ADZNM5VuuNP+X2/Y/k7OG6fSimnxmG31XcbHIG+0whq1Sboe/opNXXWmRJZZ2hL2UI9TRBQoZ++8
KcSTKG+pm7PkaoL5XYjlzXQeTPViQlI4+E0H/UddN8Ze8CGJhO+4C5xgN05EfmzjytzmM5wCKLeF
jXJ5tK4Cy1OKn/8Zk+28C3qydD2v/K6sjhvf5FkaHyHjQsk+lD0H3RZ6MOyTGGwdF3XG0u92U2ZS
hK3RobjWE0tsQQrDB+as+UygA3gpJ03OGaLB20X2utmy+OUr6VlP5ibUwJEzlVsZVwPPRIT6NRF0
N0ZBQd9VMgWbnZhTwSp73z1ZmL9Fz9qb1FGqohfq9mwZf+0Wo5ZgM8msrAW51quR5JQRRWhPDW0R
V3+jNuVv+FCqf3IucoDKrVbkBvHJg7Yglzvneh9Pu4YBbGSLwGvRvUOFyh+XOGuc/C9thMr6uKd1
G+6HvH2Pne0WUYjM8CHI9F+2KRaw5ipxLSI9PWvmfTVXksep0jsB63f6x8TBg733F1cBC/BFejby
TzhC4ZIhYVoxE0QpEpTPPHN1jwPFiJYuUFfKJ7lILw/SPYhLSa4ukAA4hbWfnkucb16OVA/KnCZe
3SUcYw//5N2+JW25R9kuEjTZ1sT48PtY6WExyZGE8Oyb/FK1GCutbu1ZQ5BByEcbEJgk14yROD8+
odwfMOLdevy2lPgJgWSJ7DROS4+BU2s3GZxZYMTn+8ADt7YSxjkNolrFFmIYUhQdtLiPPVKSs941
6RKf1umBe3+SZPHddEzAYZHynF0/kklsujv/7fxnNOLaBmSmomexaWGyWCMyAzRInsw62DqRrtJz
BvI3t+np0BUd05j+OjpHxkiF0+qcWDKjxNx0QjXClIdQxI6AXleT0fS9iix/YYcwowW8O/inKf3u
bW5YfglMPvf5MBcnbHNdqoYR4645xZoE4t07LYoajiRMaJpWCXNMigko+WvBqNGNxhdupdhnRnZC
R0RTTsGXKZCmWP1fxAJWT595OLiofOi2agxNfx30jFxR+UCLa9NIUugkSw7dBalCNB3pJCfz9Af1
NrfVivO8mYIHHyA3UZVvpKK+jbYF81V/IL/5qdsBXNd1+Wdb4kJcWhQH8ijch2laEsFdlm5Tc4Cu
nphOVLjG8v45Rz1AZB1gBdqNgOPuDTUtLQGHqbtzzjav3ZqN//76jVSOxH6QwoBMaWX68Ama+2VR
e1SboB+C37HC4+j+2LYiXIsh/oFfUn0jWHLEox76QlRQs+htPbbYdXjHEQ0Jw+E7He/sa4gWqp4B
ltNuUYgUVLh1WdjIa+BI/BLD+7mC05sOPlU99Gf//sunoi84IpMOVH3PAe1g3eNB7SsfrihNOknA
aMvbHTqdoESX93C4NE+whHEVkSiqq+yjqq9/aIi5HkKq3/tV1wp3KkX1nj+TFJ4+t/pUqcU/z3CW
AE5L5eH585fytwo0pxnr5/U5IelKnrMdt2Mzwn6Y8+P0I9PTAZqDqctmelf++YB0VHqhVT/pYSLD
EPcnk88FvjjMgcAoWS4BZkWclRJZqZHTF61GNqt7xq0gHqDx/6y6ilGeyA6ycpXsjH/6CRAKTdLV
RtO0qLzXnGCa1aUXfCQxNKdwcxKtn6dwzEFu+FGzA79MSnPh8DyswSAkj1MGo884m0xFOW0WLh2n
ed7c5sz8wgJV3KznYLQJJr9X9ZN58iZ7OuoSAhXvT8QlG0we74vHrTxrcgEXwOO479bqX3l/IUML
kabqLdri+roneaJQV007PdkGVvM5gXD7+xq6l/QMlQg4mrTUL0TGI/x+0g8x3c+g7MdR4+c9u+wA
U+DDqSJu+vIUH0l7b6U3c9y1IsnPNcEJKO4/n29jOdRU9rJ7ZYZHYu1yRvQvsUKecVKFob9U+Pc2
di+GSZUs0NUYmmfD8B4EfM5b07V8kD7kD1klekkc2oH9VNK2Q++T4U2QKRO/NRgStj5spJb2lo9f
6PW2yO+/+cN3u9bvAtpf21IZyeHVSCs/IkSY3X1Nbp6urUAogg+e4aB7Vms6Xz7cF6MsZzq7gBOk
PGpYywBRbzukJBtQodR4EwmKgj1WDlu0M3A6DfleUnqOfFb7gPDdTq0KGzdPb1aAtGpu+BsP1yF6
CDn6CP/Y8Y0Xtx5Ti83uAwmyPCKXJOC6EoQxBZabVZn4Ik3kMYTFgVJ9OCcgPgZxJZeZ+bx2uueo
3nWEhFhOlk9WhWvMAobpFp4Glqaz+Y8Fcjp9ABGacLkf9HuE8ibIXL/tzyFUQklc/c961NMgCXoH
u/F6ZX0WS2XPsP2InLlDXCqg5CkCBS0XUIBGrCz0hOK6J6DUZrxmnwMNFsci7nk5yKhnbtSv69ep
hfVAmWAis+zuH5+mNlFa1P4+rKV+RLKrkkOgT5t51DdmZyLw69ucJxUEJjS7fRe9kX42gMAZ3h9f
J+Soue+ijz9H6Jvon2ug2+4Xto6LR8yrkZ3vQFkmgYeOkmlevwonSK0LPE3Y5IDdxWgZvzpLkRsU
2P4y5xVL1rvDo9q4+LzCdADwrb9JKI8Jx1Cn8nOTyPfVhTsqqDaJXaJJgybD9Dm0cmQ2PKTCocPo
4NMAL54vgRFjcs8088gKG6aty4IqhYfzNXEWWNo+wVUu/y1005WKi10IieJ2h+YjS04jdEfAeYnd
t6NtAzl/tQscjHVU7Pl3BsrYl4tV5RtZztEGwTXAx1MtYrbgK7ENislZvvLu74MAjRiDkeU6UOCZ
GRc4fKnY9o8t9WsAfV75IG6qglNHQE3RJylj7nuir0nY5sWvyTCS9DaxWEJnbddm3fBHcdFfFGT2
p3oJbBBRph7tOFuQpyUpCPqOHv5IXk+RgWjnLYDa3BjmhUMosrQodbqm/wgrruKf9UmGcSxYpgEH
+pPveadaWGBN23+H2KtDDylRKnXiCp9ENx6sB5Xhk1JXKUVWCRHja2DSHu1imCv+yAAoDUQMi+Cu
4twUh/5aIN3hzxccHGdMgalQDCo5zrSz5I14EGMHIE2sYW+NmAphNW43axrkJ1OUk746VaQ2yO/R
gLrRrbj7bDK7Atz4Dvwpc/MERrHX6bwATduwvg2ge3DGomiedSx2ADcatHW73EHp+3I9yi8zBI4S
TGgM1o98dBwx2SpgOY8PiKE7v9UhZ2A/OUaF6zBaXKdV7oQOpXBkRAzmyQnslQQcm58pB8bJMV0U
i/UrBi1uyiYZ3wk2wkTNQ6UDqnJFjXGqqJWt7wmDVrwRGc56r/gCjvJuFI9QMtFBgc1ncpbr3Otd
sJ72z7MWay8TUcTLCDzfpLXzSA8hqivM217tZiBKEeD/yR7oBUdJDNZLdyO7axvvCkNcamrVLa1G
Ecds5bfyh0greBeu5c0gG0s5Qbi68uSlN+1+ExO911QOFMyIEUfPZjOI0PfSVGAhCNbmB8icvh7j
hp54Gfl1AMQHGZJYmt+1TsGuLfOy85X+Tndt6rPH4/9+mFuL+tJRXwl3U0ucDYKNGsY5rCiLguwd
CWH0P+ZBO2gPkfhY2vT2JYapfUYGFS41VwXbDJr8l4XCZ/gzGg1kHa/8YoK6JgILtw61FNmQ74fo
zWt7IbyX8uCtv1tyW7ScIIkH7dVsTCk3hSCHsPqoQvwH4xGn28fWxmSCCX8rHriKre8VCkOU55Oi
KQ0s/lV1P1fY7ZVMqS4if7glNEBGvG95CKjMXY2KNGgV7qwjObkLK8VVoHCsznhmQvK5oJBi9Nm4
h46uAfNX3mgxPKAw6Stc/z2rf0KbxS5iU5ssVdOZhYYEZ5yCSYg3EXYQ8WvKNFGj+tMwQtZeJXdB
QtIBCecgGNBHfUGsppgwHA4rDD5MeiSq2mQsiiJSQisrCszwcJTY7yWZ23cH2lbeWu3K3LRUtTb/
3h9UsOdWtRYUvCyZCVdamNRao0hsLC934Qpk6VQwn134/iPzOvz3VXM2nm8zhbjvy2B9qO/3dpD3
yey1tfx5mFTMpzJCg2+Vrm6B1F93a4jSBL7rldMDdmUEI10k7imF7SMvaq9fFKE1OucUl9jKWmw0
DElUQ2cTSLX8L15PiYC8XqHYm9tJ905vLffpotS5SIW+7JFMkwyMJJIK6SpioNQkfxtALsVky449
+1guvRax/tt393ElUSTc1tkxxhfdBam9cG/RA3HCu5p3VyexH9HDomG5b8XkFh+uOEDJGwDfcCwu
LJbjsd+BHp4FXsigneytycnU21BOSbG70ZK9a4qeIkn73uQhwvu32BrMX4fkDlbvAkoKvvGmMnOQ
34SCWratK+oY8Uail0amHIc2UojFeMM9wZ0QZPkzwD1sGF7xs2JY8pBzLnGbuKn2tNJjkzRLLb3b
GJpnZMSkPZ41PJfcsDb4kKDFAC+AT+NS/fXaSoovL6c+TC+ynrh3VDwq+G7e/ngwBEwcAdzMjqND
0qhnuWgaUM5vJ+DSIHrhiDM+m77FvcxZI1Fp2IZ33dycB57kzVfo+JcOEkGVdyFG9j69vHh6icow
sxCBBC27ZstZOl+wg2BvtrtK+AZXyOJvDcFV9KBgCvX7k4r1+Yia5FdVT+3FY3SxIGdQQXeLqg/1
zzImRJQoVc9f+IAYFvWFh1OBhp787c3KmtfI+fNwmDOwTXEGNPls6aQIkwkF6cppLH19poxWOeSm
30A+RBEheOBAclc74O7H4AomKXy/LCyKdJrn1h/TwiBjHeq4ZHC0AN/JiCKlDaNcGKww26tWMHje
jx1wfyfs+THqNEtbh1syumvRQYLXzY/HboMzJig531QSAG/0/5ZYIc8tGXjZ5VnXfXm4zpI+eR/u
Agt04uQmSJcCVO6UmZ1uKotO9E8787GpJElhmRE1UGsKwwS8j6zranmFljsMjz64OMK4VixauOFF
6LbvU3blrwfhTuNH4THdIsA5eIyGr+3UY2Xx7PisvUYPSsncmAe4VaJG3ZiTzpm73bM8BswucjFi
cib0Jnkfi2la5QsduSDn1uy9XTlI2HsBIO61rGeEo7tYewVtE8n1syrhq8dTP8kgO/a0FORf8j0i
PUow5ItC5TNJJuWBJ2Jhj7p6UFl1T5xFFE1pOcm0/fGAYL8pot7FAi93iR0SkG5TFqCcd4cBD0iU
RmLpQPmE1JAPm4JsisjJ4IjY7PcXW8qbjOyibM5mDTM+2xx8ko7FUBMY6noYX/mN20EN3b0IoVqc
ZoKaXfyXdxrUj72JKHq6+GuO5393+DZQ4SwbLsd/w4zVv4+HfNqrHHTEL3x28MYQBMsHu9rgWX0R
47UefTV1udKqum+f6oTVcrJkbtplPeRnYeudqnH9XO/s/FcC8IQW7h+DLTddvBceLokgGMeI1JzL
w5ztTscb2OVKq33lxrPffe1H4kWJ4e9nYx8xyldFbONMXdBfDuBHHdUL9fqJDiQl6ZFueBd3vU7/
G52Vq0d5aycltLEx3EryIHs2V4DGdlNTIFUG+CLjzBUgU357pWz3b0qETzRW7ubzzXCuHLO/hTgR
0S2appU8AAfe7hXm3hZlsLvvjjv1z6yyiPU1lfXMsXts1sechlrJ8V6DQ+TMQc2uR6O7icfXbNh8
PTGBhbs98zWRHtNgUKbwywkfIIAkCsHBD4Z5FW0hGJDGXaNAYxiIiJvi6wvq7Y2GV0LNQMxxl6i4
bZ60sAz9O55QwmDUHOD6kuKC7h8uW+Tr5eQi3Z/Y2uRmrgzBOUmADxO4Qhhp2J71EytLLyhWVFKF
yY0f6NrpNNfdZIO9PUUSfUljV1GIFc4OgbR4qbXa5fYOycPWPo4weOdMXATLx48YtaYJnPMDQjuN
soaGBzzUvm7UUhI0XOrmq58CfIcsBV9Ny34FarRT244mKSRgiHUhWp7KewdmgE9MOxzGlMsSt7qC
vkS1FWJLBXj9tzPwp28q8P01abXG5U61RuEJsoG1Bo+Ifk5RVdKbe2ZvNjxpWQooEzmNgvhrE2U+
iCClPXVldfLFDWjZ5aVmBOnJtL4lIA3DNwvwPDk6y3VKjUSw8DN1/5zTnIsqOntaLaT3dLVTiWwz
VWD0nzaLth/WqWLUc9JWJV4gtkkJxqtvwDpY1FVFUsXL0GlvwTShwCxbAHT7QLbtrqZ/zrUeEN0c
59wU74tsMwggQntCMmkHDPwF0k6jLJvaml8KtphINEybZxFAW5iJsoGqPpMQ6F6WjXRaIyrtcHKE
QJdse54abm3OaVQwB/s7is24k6roc6i3Y8ev51mlqtV2RcXAIhrmTy5HnB1JInAMacmg2PBILQ9M
zT43N8zekUc3LttT+osW+RbnWP/Z++bgQDUHrccDmZMT2vXxQDBx+ngQxLTPWARBCIRMLMxVbypo
dkv+bguzAGZKn/xQ5Jx9mDB6QLvHq5yE6mxHoe+oPoZDFO60LSz+jcDBBOg0D6jV0F1I/Ua5BMll
hcxxEvb7E+4kaoNJ1I9BWNMlYFy0XP8vEKK4c7TA29Itu0eTZLo34w3yt4jTmqYgv774MeOqdbtX
C8steS2sk6SX0T6yHu3VKZduiWgVq1/Yt/hczAChn66EwIs1bEkv1YhrIPouVpV7eiKZ3PdnxdR0
4FSqMWlgv49rZwm0Xjbh4FdQ/lS3OwrgbUbnntpzka1FvSfayFUXlshLl+6M08BB0GVxVDF94rvx
SRpcs3LjO8Bl/iEzSVSgjVpdS2Qm3e9ImWI4ql0IDwKk+o4eEgyxFf8M+kb+9aaTQ8jWx/yM4skn
b5K8ls/dJDvtsqNn98i9Z7ljyBBSm3E5ZfC9chs8fzCxHZVcPtLMQs9cuwayWzp4yHNhCGeQNwsj
xnYYbVwgaiRbZ/2r1zwnwSp3x90C/h4he8CtG2xDFxL9HpUvv6F4zl6GHaLj1livnUlWWL9ZUcy/
rqq12jUsj3sXfv/u/xKpqpCA9dy13GwXiYQGTBOZF8yS4aJUr8h1gazmUe38DpK9L+MhpL+pVCfL
5fiGyDwm850ZS7xGWIsMLQsqlayllLUraRvUeaEakXU3hnhc7EmcRMNWID9v89Iia4JLVogJ3lpX
iGO26AwbkVsZmi6dO9aTs9FEteDvYqpur9FpAlyKncPH4kZqcdOnQhIOzPVFfcGOZo4PF/dcZ2ns
Jv4iOoFiBwWUxn3I4CRHZnnW3xu6LBx96ViRcRYfzj7/+KjFTVv/sMUOn2/9dCOtROnJAp6PK13B
Sufji/gDS2X183Lcaplf6WpJMoZef4XLgggQEUAD6JfwX+mCHwYJ1bwjSJBFxaw8PYLgKWr8dcOA
djwd+VEDsCJVur0eerQWUSVYDkFuW0rcgCCB1erbz6Fw8F2sTuBbIyoAxKpJ9Pmweev5f/oQollT
XMJvvOGAq4j4l2p5z4HcFg9unDsNRDOdldZZKu5kiErJgsWTlUaCm+vdIQTgUsbsDnslR/hQue/R
7AF/rXQ0D+EdL2RhCZd5VhMpBiCh5q6q2+FIJ+h8D1tYjdzZ+XvtXZBtLrgs1mVHjulfkvfneEUK
kUGr/XHFNbwnEc9nSgvjxBqwbr4FsT4DGKJB7k3VyjyRCLKe/QL4m6J9F+6qHExmIVIetVxdavaD
/aj20mKwVG/w9eZ3bWmKWpth15p2fzvnPnZGyc7v3WQq3VESkyaMeiPns5NvjaIKVeYw2D0x54gV
s+JSRZjTwbvFMcH3Xp3wXUoR/GLKtTS+ryDFqE8FVlgqkee/KfltWtVjxoEzL8PyKdnG/+Em3EIN
Sf/xKMJCJghYfKozXVBb+oG3D7cJqKA3QzqOi6PYWRtI/dQQyzAMOXwnyRaO2XkO8cVjI0co/n14
P5hVOu5VabEzkpiu43RQXuVACwpZpris4MfDRxju7JMMLAWDFR6bnz5Lv5hBpX9erS4FlS+V2srS
DX5Dz4YpBjZs3zN6mZpjMNf1VmGcWPm/Dsp4/QXLC595TdaUWCA8hawEHxDS9nahmaBfQDlBoojy
TtuXWB5aTxpzqGPdnrFf8f8u/WxxJC3rQzZjwMKUva1JYjlHKmJmpptNd1YXHGAiCHFBTVYpRdaB
TBRUL+/SLFxLEkQ0cTxZWO3ZVYTOfXI4rwloDIx8Jcp0/b0GBdBBDPcd+wuQmYqdhYz/b0xwKzms
ijZtdqGR34sL0sPh4U7OayJrKreRZ6TRyBM5IZwYQpB+xaP+9NJARI7PLQ99aE178SGGQZj8vhye
ltqNQEkzY76ze8FFUPZVd1pzFFZ2g+Mxux51acyvAdREkkEyy4UTILrMOMSjNnJ4/PgC7qb8TcyO
v6kma4jKOO8O9z4i4vWNfiWSWFHAaeadxWQfObn9LmVW3ii/6BXgPFjWt4RQ1OIqJ4zNowutjZ0i
BFlR+uOGXF9x6cQb3wKp5vqU2MbOztoRhqv+EGsb2MAge+U+k2/A5Zw2PCGn7ePb3Kzm9CtBzHpe
qHvdAZE4IlxBjNGX7LSf8Lwov/YZVViiX+hy9RHTMBPXXMJTNnt2s49UQGY6U1MP6DVJ8tEC9Lri
mH2VbTs7BIdmnM9cq7RboCVPjcaAnbEkgeA5dnonCYmsFXt9WZz7IU64PTcPNHZ3XYybnTP8bsSC
KFg4Yvm+DHqDD1Nb9P1D+1DoSlvTBucyy4nP836dM+Gncl7bCjAreDjzOo0ZQgeXZUi7bqoLHNEd
/I/u7j5jHT3WTfIj8P6+7OWt+nt22qvzKZciq9AsVBf/zASvmLKxxaHsEbyC6o6i2LI4v+slv7/S
p6xXWdmgakvJPDRMKH9kXmjv+kCq3hdsWlc/5aKfxe+iIWOQqO/UiLK21FuOwda+U+bColqYnS4V
cvcWG4U1V+Zt7su2vcK/Ks66WisQAZVg+45Cm7h4kJI9QBfaRyCa4i1k+3NidL0PBcxqb4IWTX4L
MVEP8PGMzPIysh+TNAIn3+ozKvw8sfHk3/DTQXQL1BuL0g3lVSJrC6rocLoFZvs1HcbFxK7KOgik
2v+yyHuHm+XI+0su490nQtFxr3uaFkFgRXSkOKbXnWOsXnfbKCYLZWKeaLUybpSKH6LW5KtFXTGD
0Qa/DiUKSZHgTrffAahqtI/i2Ft/5xRLd8xEZraF0QbzXC4se4qnG+UTecuTI5ahrLredZbI6bFm
JToCocwVKJc3jYF8X69vL45kYVU4xB6ijESfCz1sytjNVfpAmIrC/SnEqxpBAEN4Yc7tWh7f8QH8
urnOd2vF+7iN2UaFoXFLvWoDfPDddQ9HrHJqEGIiWyyaTsLWeZCIb5rxAs60krPROvDuwV4Ngqwj
sNRU1B2fsfAIyZYrOk4+J2USwHPgR1Oh44jLS3YCE8Eps3MZEx+NlpiWDXugByb6Siq0pOrN4OUP
d6r0n8EikO6SsGfhG7P3KNcYRsu+N1DEWVcGl40p4DPTbo35k168IdaS6R/x97h7pcSUFh3PUMa9
Sxc8a7cP7y/Du4PnqVGQr0LEvZjZlQLu1pL4ZMNS8qjM1084JoSNnVbx69HEuz0LzF9yERw+uD9C
ysFrAxp3G06p4S4kqABbMOzWuG0cr833Ke3Q2RW4XBA6ivtPM7SInio4gtcbX1DmtUWWIJ3eL3oX
PZGzJVlsBjVyHepPpnFLqyx/lyxZAFATT/nSlk9kUpvQzwy7mDHu2dyffneMdyQ+sdqkcOEQWnQJ
Ew0dd+T4sekDjC7iRI/aFNzL2ERl61Rfl3Q09BzJUKy5s/26Rz9IRN9Vw7NhBdLAF6rBKSJs1IO2
9m75CcdwX5fitAFFWtEx4dMrnsjNL3gCPfpc0Lox6w1pYDPZCwRYfncmyEdpQdFI002rVi6TY78E
53ANAoUy6nQebcsZird3oxbdktZ2SbquxhO2ApUlX/k25ow25Ht+5QobFyK7lmDk1LHfbFegHPpl
jyUor4OSgWaHpE2vrjS0ypqB6Rd9AWIEM5ht58r2TxGZIMQTkd+5x0m9tY3VXbzoKFwxgyQsgnBf
agtH1uWFuPgWXvUGc/0PlM4dtjwFOSLve2c5PE93vksEg3fhTuW3zkPtkWb+thzyVkOBOQOgbffB
syypVRJ0FFcnurTcnSMkqzOmA1/GnxcD0lm6IGUbrUjq9js/SLxVQ7lkN576imHWWcaotsmGghYs
YRWr4Z36Y1YrVt1o/FJOAchcsSqONgMV9EQiYWkMAwJQ50yOmxmI9gbobrqfNLKNgln6NUCdYxVi
uMLk5XAHpJAC6a6nLA3BP64IlUB4iIWvTpaxNMmeFGA9M9GYXGe75o7nHAeTm5N6D7qtxdXhb4Vr
OkKU8KFQ0e3al3iSZBnQbDNZdUkqQJ9S67n1f9ZlcxUwUfSbvbt45JUtQMRq4w3XUZ8cYEcZDPzW
nR1V42F6XVP1cy+SsKfwBmnb9UvNtkfsywQVd3hLvPjt8eePvRGypoFNY6SKn32hzDU81g16xSYk
p2to/5gKELbq/LC7j7kDEX9l1g9YQbHmimLKIhEfl/QXXbza18I31HY22+a9ePxigFX6a9u7zUdn
sMFTOgO+des2UnEVwqsrXRm8qhS+/9S/QIq9EJzGv7+kJYbyKnaYyfIaccxOP3QzWM68sxlsOgKX
hZh0kKCQMq3+vQKCQlWAvalg90as42yuBvQYUDDYDVEhY4wz9gTBjQYyGLc1o393scBRXk/IRlt5
Zx9Mz0Da4Ie+JjkbliyX1Ut9bcqbV01FrxsfsppNvLcK5uFywkWjIQ+Z5qmWZBIe4Jz0bTJeBYYj
TUOres9LiJ1dDuRmR6Fz2KRFl6s2/ucFhTAzHDlwmhQdzlUS4jhPTENnIwfvMJMM26R6QAJrG+53
txAE3oO6tfD+1PnhGMfOSdTUta7pVDQAldtK13FaG1MrhjSqLP4B4XQBf45l0YPb1vZXWA9JgayE
qxGgDkncTJDxj00Y3aDNYVhkZBPIEad5AMoVRQPjmfkjCYk9eRsTnDsJCw6k24vrYaA9puLeZIZD
b/A+KtH99Zvl3CTAxE4ti3f+2cOSdfBp7aZqmm+k8g75d2vn5m+MYZGi21n/d2zxjFSiXMh32e67
fp+qtHxj+qyp+Jc9g5zfoa6xh+TDnWpCydsfDuPRmStWm3YOaSqehIDULrRNVDVGEksNETA8Rqdm
ZLhadOmzE/nTawhJdqbOKO+beYU9lmgOlWDDDFnQgX0HoiHuAViAdFawHukYKLv09SM+WPdhhNss
qTE5j2uiUmcX82LX7gP2TdekD1XOocFSqHMXbdJtzHhpP+YN31dsSuXhf7TJn2/rRLnYXRotRIB2
ehnpnEpxaDdbDAfMVnjMiXPCrzTsZtwXdKABerznyFIVJHPqxwQRUheOipqMpRFruYyOmU2p17PP
gnqRbG1lnyeOWSmC+T1pIzh2K9hCH5uHjiHgfFwGZxwyflIazaxgxnzWrHTOK12EVrGWwhnQLSMj
dmBTC0UkGKp6wt8kVRkKF+pMZ79KoLMEoeuRlWiUsz+/B2lHPeadVk4l5GP2F0BptItOuuvvhst0
ZrEMaLuIuWeBB0N0qk5vT0//X9CmNAClHiegRX6tiTvDsuZuLsM6UEf8jg6sYg55uVbsviZ12oDK
9eCHg2GCDx+mCiAanXuW3Hwy5WQDTJ0408tTuchkTt5VraAKZRVwS3TeHAnLooGb5vGByDV8bCnK
t/aOAWovOlBbRe/VUZEI9B0sEXviQ+I5SIkOPHTcGm9zt9m1chhb/hFj7VxFiR5BtO7uoUZr1c6c
9tq2nG7KxjYD5QnDKt0UgLF3lxxSK2Ym6A4Px6SL+fp76DpwwpZk4UqF/5rJDCOrgFp6ChQgSelS
K3xnJerj874vofrTKszfs1UjD6O6qNbgBS/6MPEnrheR327XLrgssQGs+B27lJUyYLtBNWqpbMS7
340tgZ3TFz5W+wJz1WFD6nJDoJbnRmVhrmtf6ibWQpmV9y5D9dKbikvsqCDmdac4S6+4AyDY95gl
BZ/m6qQJiqKQZIzo+7tlVrrq6b38u7byXFZSRfRgooaJMqKBY14VdaBgw0bjy1lj1Iey8mhS89h4
wXT0Z/NwFEoNkz2dFoMy8V+Ol/BUZPKj9ByOUici4Ski8PR8Ot2ZqXWJ0sdVheLXADkBllTzwY6o
uuF61Pj4WUJgIDohPHwX7jSvb4GOakUKCl7femOrBt7bNxHgx8Mnae4Ffe0Zb0Oo8xUEECGGfoHG
8L1EcBaAuPqxrnaCsMJHKkoUPUGoX2aDvQjq7uEH2rj9IU+QSaBTNwEqJGOcrCpmkfBWmjYq2y5z
vk5oZIsqAhitBfMbp0kBLyYq2Cpe6r3+dezhsrwpd38aFOEJKO2/VrPEBmvfy6h7RL08UQiunmfj
PKzA1WaTcu9lWHjjzauXjuhaa/+OIaYx2Ag7QIuwRxtqsuHv1UptO+nSuSmfZ3klIgATp/0+5ezK
LdHJQtIlH6mPsYHtrKj7gDJ0FnvJ7c6jMHF8EWnSd7FQXfVMo9KDf62zdRgtO6Wt/QJnc6LCQTA5
KZAcCw9Iru8vag2MK7vuM8v1HGyf1TQ1gj6jRS8SmOrObyE3vZf91ZMJqoX6rfs6mR0AoxQQxuiI
7ygk9LlSsBDJEUk3VZDxy1uxMhwHdBc2qyrXsvODV63X1nslxLd+k+Li5jbPEsGjdb/11FZSGd8l
kK9yqWSinn0SZsAvFjIHTocUEctCALSdnKPpMfrvzS7piB0BuM4dsJ8o99ZLvHjGo/ObCmAGJ3gf
mo6NFstRKLDQejBX3AZtGwOj9eMe7j137Qbl2VXtEBi2q9eEiiJRHoJMa/zrl2tjLLyGqX6b3flO
6uuPNjx9LX0xjazuZHTJTGgo5yFjHhcQVHyruEaxwq76suaODVNeJAXD/OliqBF+Ags4lKbFiYhm
dYpPGiwDQsC3AYmclFnEVyKxCXOM/0stew8lnR/00WBzsSdL/VXVvFbk7SygkCS0ZNj7bxsw6uOd
/9ltERPSU8B66VgFUAFx3yb+hXk+wuk2nbU02+dEnYq4rl56Q9ylvRzZy5WbOu4xyidRyr8U+6yL
3ClS/8SoMMAbwLy9PtR9kD6k/bnPXgKPykn1PLiP6EawPMH+p02XDmgSC9glZuOyTpQsKOIGQBQ2
LbwgIL7gDmdJvRPBlAWhmiS4QctC2taKrpaaCE1AOdq2Qspfyq6rKBc31XiMGuXFdelwTdjNr9Vl
ECnQzEk4t1iNoKQunoErFWSgvwfJOgU6gm+k5yhPH1EXSWmYXVQoqLhYMeZ4duTUGKLKUAeJJCrP
R/jU74ltkPr2x4PkIs8cgSbPaYpDBF/GZb/WibKm541UwF5pMq9viGmZcdpmZ3B8sKq0M4fFlKKE
uIHTAb3Peg4CzQ1IJBXkFHvhuPQmPqBPVFBHIz75YVVKxJEJ4WUrzwXQHBSsJXg0A/vHWvYSoeHt
oFW/wixiHQtLfDK6O9IZBEgt4QXOJ9+XEKQzcBZPktCzLdRPGq/Z1Cm4jQGxyECjcwjVIKXlVHY0
iQyso2PHS6spOKftjSctpT5mq9dzGjfFwKRljmIgBi7ZIf62jdvZUmhQ7AfU6bZaRz1rte0mvWpr
eX/wk8R60JaPv4o3Z/vmk1XxJPW8tVU3tWj4ms3gvFcq43T45RqhNlZNU6mL9xVcKHRJc+WNGmjN
+gLFvon0K8WTN2x/a+1IpajcgPV3Bww/2EKGHZKViT/4WWGBXSvqVD6wizYkm66enSiK5dEzwCJQ
7xErlnwEPSHPHlWR7oNyhN+ylGmLSTJJ1CUgQ4pKeZ87floKGlSuao48C13MqJGTmdeKZ/02Tw9j
YYjAa9vMGDOeBP7842ExTG17FJVz+L0QJdF93wWHJSsV0ArmvYqRKpCoT7qJQrfV9bBl7q/f1Lug
05/gQztCWzvg7TSiVK58O8w4wDrSdSn7hkWhGTDZmV2RUNAFSqMW0Gt/pn89p2gVRfo2juRjFfx5
P317aarX4t2i5mwcxLe9uIVsDQScSvoq9XIyWV6V10yxJjLbql1CA7Xx5Qt7qjP+rBteJC0LHQ4H
URw6J7Vz1ToHEdM0Cb9CO+s9ghtggXr2xAUWBMarohVQyCQ+MRFyXdXStUUbX3jFwSvBqHzDTdGX
ULzYvVElgjxWYEovOo9sSFgjQu4JIHoynlaUpaJ/9fe0sfJiTkIkhF7B91o/tOqt6g1RZS+HtNbU
QnLpzBJxB/DeGw7lDXqQb6fZg/zYj0ojP8+b7xF1qObrkpxfiOJA+kD/0uRozJe3bamVv4blZB8D
8PRPKM6Z5+HvgD1vOrdwfgmhtMYIN4ZG3kWXnXr+xBfc+Ed0QGSh2rxlxkE+A48fSKvwgUIGe/oJ
n6K+/e3X4Fe2IuwHr0ZKZOcX0daT8yVDpxEnYBvYFeZg+grIdSkkGTnaJM6TN3C07BBJZKlOVfMr
qEFMpmqbanm4x//wukyDbBh3htk01kYTdXIQtDCnQdLbZySHwCbAQny7NxGUYN984b2Ij+KSN44b
8sqspVcQA/vyX4ZYoPPPvPHUHQUTVBAk+8C3w9nhyzC5LUZWCRYoT9l9mVl60JNcQ8yNin3xYTe4
+OT1BwzAWVKp+dBhOU+LTzCYvXrGlm1o0CQ4OYydnQTjbuZ4H+Yyh25hV7ekK0Tw9cBAfGa2/u6C
JezmodjEkXFOxtLEJ99DJzcMpKw9qBhGYIwbknK8Nrb1S+ZDbtfnhc6irI/m496ebwBY5pbx/t1T
mVL09uoTp2TRlkryBV+Mg5n2+cH6q217Sfa2atHG86rvhy6EhSWGSDos/1VIO157GXPIh+XKgSgl
8wvGOBe+uEGNueG4SWPZfhhRfjBpvCs+ExlOz52QKj9QCCs3e9g1FFLo/4tFgjxwJNNP7HXx8hvz
E40EY/dOV0r+X7ZE+7CRi2/aZZ2Xa9kyxV0eKRWAKI66XpewH5caBZIjg57dqYvtPNScXrYeBGzA
quEREWu8q84kImkbTMKSTsAXy/iOuDkJm+v7bFb7VJxjYWvIpIuUmrvc+YZzpNqgEZBH1wu3uMDn
iDkZ0x4ROy4VmBjXOaNhNcLtLaQs3lokdLt6//PD4LzAWAUOi8juPSTlvyPBofieS0wEFRaZ4Xze
/GIBo7KVncLw0Oc11ZB54lpaPQPOgAA7atvQgE3iaQf8BTNdeCjJclDka9ZEQvjLYCc2dUBkBrc8
hJ9LpvC2WN/c/GykUh7bu1SpGpjHY0XW+rDxTDRcq7X013AEo385KNM1eKmfLHLxV2EFC40vG/N+
F6WdroHiQA4OAMZ2t/dV5Yx4f0HVFErC1GXWO1TFSd2a6QxWd6wd0liY6aeo4IT12CJCdwjUB5uc
JIcJARIL5pgv0jfWPKbRTsYwL1D4OASKPrhSGrjN/4jGAgtevfJt5a+1TQ9MsJpimRuLbAZ/tyXd
uNFGPMKdCjYOyYrTGmE2VV4AtSxDuDqCsbkxsQnDX3kk8IO801QXwdasFuSIZM4B3VRwm+Kom0Kk
h5D2dh9QeeHo18bGLeSe0GBqx6BvwOVmHhXADEzRss2P7Dv60xR4+X7aMmlTwVy9kN0H0edzFm3r
WTKpRHPadBO7N2/Kkd7eeRJNWKMT8nzL8Xgu3zV+m78J9iO5f+aCSawb1eLCOhu+n77Lx7dqj8m8
z4hEDxkCAUMFk4KJ+MmzJqdqS6rwPV7XsG+5CmZ97sa65jCfcZ+ecH9Nj2xzhb2GYsyKwTOJ9Lyt
rTFlfqM+lf/lRzvsy9hDSDMkEn12EeIfgSm8O6BkoPXiq2uyTOkttRtCOy/Sb8vkMXvUzPcPIpzF
sr7V3ZDFcAXWpDubfdoNlwwrAfJmuMBSucBXE2O4KPQ8LC3hw1NygwKWdLL2c8MKbjgqUrUft4iB
PeRdzOeDtCd5ssklq8PETvc95wzxZR5KvLVxkelwXVNZItLgNkNWAdwMpd+QJP2edU2jferAYLxr
ewFVjCKbs6ru3DiS/ACp1yDTi6KMNLJdKvt2rD49WOx1irNhujsdw3sugu0iSCdLpQmNGdyMxAm4
CbWOBAbS5A8MNX7keEroO7KVTVAQV5KIKPoMcfDti+0zF56EzWprxw/KvyAbSa7hHst+2ZdaW73a
8FUDVWIb7DTbP3kLfkaPI5X5JMBjQLJE91euDGrvCoDO+Y1U/cDIptRH3Y6/+1f+EjMF3XqAdHBN
fJ4T5pUeAGUrRyPyRKNkakezBYi0yrhpuQcE/lnQECl0t5bCABtVMUveaT+81gTxlOtWQJ1GWY8v
xkHO4QSJ2RZkGtNaabQAGG1bh/ZYni4NTVmZ78VxKXk04kHijQkiFOg9WsCxxQ79JukEe0IxL3Bz
cVGr4i3WLFkKKl+8iV8E7UY3Qp4GJsI9vTt4ApjuMxZeRSqhXwPl9U/XR/QibLavAFriK9q6Vi+1
SWOlSvOvA4dOyX5QVBczY8JERHZUc2wZnchzEVLzt1zIFSrSqG9f20CXaFVY7gGfLxgxErivbj8r
ujZ8UnTWLxFehH9RezT/sGDrR8shz+XG4c+W84skfVmRswfXWFdiJ/gvHRKuv5zveFNfbk/6nLQD
bylsJYs5NNSY++iG9isUd3wxSyOfWXWO/2vxldgUSRoYGXKHOaVRK97kIGb8Ia7hnNc3YQc/tqv4
RMk5w201D9YsNT6sepBBjZH9oAiUqaEAvNtqjKYYysRNnGXp2Z5KV4s1f4Tcy/t8D04iYWnHTZJ/
ly18oKWcutT107ypL0UV3myq6CDN7zTDtCorBk4FyECX7pzAKCF2SmLM/tS7RLrjPyLlT6kqBWcp
sgWzYtdyaXr8SkjxnS1BixhoCJTGviEVOuaSv/lhLy/VT/Z/tvnTqp4/vNcVoaECOAbSaaRbE3nv
N+dHp0UKf/630V1XagLgNsjJEgS/UJH/wvDcGA3F+4RNCE2OjHoPr6oRy/x2oYnHqyJb89PGeZpg
zOAz80eJ+wtPMTvGj/T6UrzGd/oru0NPfKRo+N0xcIEUn6T8Av9YQrL+c0QCHNGbtzth/nb/1YZz
/EKIr0k0pUelYhyipT5b/LQ94KN3oh3wGaN7Jm0bi/IYkYbKrmAfmA4IMmcjn4Mts7A3CA4Vs5aR
W0EEqqHfpwd8LMfKICl8Oyi70/fqrBDoigrRKZutY91MfZs9+W7fqjUKfl6Af4DqwRKVoTmRHqEj
K2S9EwYLlEvvc7MrGXyoyMtc3Fo64zBHQMEVPY9RVP5mTebmwWZcG/U68k+OydhpSeSMOAFyouRE
hPoV1kYyc+23hnzxxhkIdg6HX9fYI6YgNbaGg9ArFvd9ySUDfzWd8TssA1RUiq/vLh5dncwwMODY
CD7W+9QVHyHYepUFpRv44DTooKx77bZAZheuUtPTGsBfNOtMh0qpTtaGgdkJ4rJQBptTbV6sPZ3U
R+i4yXlkKIAy4wOAfBSIXHP7h8t1q5MFEceoMIkOV+O8lahDLiOI8s6G+ZrgPfPXWTkF6E68AalW
PuXdaaZIRdopGrELfbrB9Je6L13SjVTImdTjcAx9WRiygZtVnvkV3+/0urW7CefLcfW/ho1rK1Vk
rijn30jGTHMaLRjRcMODtfHPwqjW2Fqgokmcr8N8CVG3Bf+6uUdgz55Ms1ISvVakdTC4t9h7PBel
iodvSvADSqBPMsKuq5bF9X0jmzLiwYtcALfqkehhXgrGy9K6/eaubpAO1T5vIPy6/1EgUf5bmcnk
zUlgXVn/kojKPmXhPe1xVIbp7PDggVRSKGiETtb057Vj4qUZPVcBIBrTgZIu97s9warMYCHSHStw
JkTwqSsDHSUM5jLs8SUaIYjBYVoX3SxtqGCin759YS98UbbTUSJsDb9fUOT/h567hWUjDZKC/kte
sv/Uotkdc0ZKW9bMjKuUnjgG8ktAnyCdtu3XC7/nJ19Ak1pffYSU4pNNF7lro3uY7G51KE8wMEhl
Rd3pMlftsc8rGwJzMw9sl2Ft2iVinqh50oBnYpn0ZBHl8l+lET+FkzZD7VwblC6QYCmHFv90odNL
0/mVegnNjCJYnFdi0FwfUqWH37A8i8czmC2boOQ2AqXsSGxr+cQAolh1wF3dMOwB8PPzVB1qX6Dj
E2EEOAFSUHnp96HcHYSKecjSndVf4Q5Qs0jcVDHugoMXIhhQt4kAZJB1C2Gvblb8rLFB8KY60Spy
s1OMJMDRomlWmFy9fGh+NRLwrniFYDbQo0kePeSlGeB5mzdBA/fz93cNtoI1qobM072P8BE+b22e
pWxzfUyFevbt9SQeUvNQ2i9osEC2J5ls3zIUsxIJh2hPcPCQPdQhkxUaJKtNroq08cANPbTq0hmG
ZMIh7IGaj4NDOvA1on9GesnyTiEBoA0YYMP5hvWRIohofaiWWfZTQdRPj/bM3Y+2/RV3sTiD0Wq0
WirmAXA0ShPS6sXeNPJ/4g9hHXJaMXV3wX4Hkilhkz4yEDiJfQO/LGaxXd0+qGHsxAh/cU2RxWwN
29m9q5ZhKv62gZKStciAr+9O0+csXlDE9GV4i2O8UBtNhCVIIBxob3BpJ8p3az1+OGbgZB9Nb5uU
B5iIfmSchCDQcq6kuxpJ2xleGgO/uzuljWceEdMRcLFqs5Dm7E9wtRKzwfaDK1bsGQxk29ft7sGQ
jtmyClXzgysVkoiKF+3O2KO1U5TENqYYFyadTLAw9ejjfDQR8gyxUt233MYeRr4GCHhdlWdsmCXx
ooMV0cbA71gVEh0dSHxq2Wh9o2IxeARCCCBZWGfUnYnMW2Vgxvrrfmc8zIFdPLxTHJye7M2i+85o
e9dptX+SajIzW8flkrkQTqbogZngvDxMPVdEtu5bhiPlcEQupRdVLrrez93VHa7wTUgTjJWAulz9
OfG0QArzKxsp3r3FRKFmuwXC3UMV44gnZUtFPPSm6mZbG8xzWBduP67Lm+hBkR9unfJVVEudomUn
tlTkhP+5k7b1X4NT8LsiiurxOuMPpFunkawfhVckZ6SOTCTJDY7BPVqMtK79rTYF1S3kGIX0SH1Z
i9GA4K5PEk2nvscSBHygPmcSviN3v/aBAuMbh4YgBjFwmNifJfmlNXtCXz9j/KVyiQTa2uVVjH9B
FWVLhecS+/K042YvfGiYG0fQSElMo8ae04GoBMpsgfpDT1TV/bHP7bK4y6b3hF9P7Y9Te4N4j9+K
TPzCZOS729+UGoVaYl4k8tUHeVGhhSiwKIk00a9KrU0coNce7OiYRQkYy5zaybwGuEAPurgVtlzD
HYwEUjkaI4NNSmTBjw5z4rvGg+Qc41GTywGe64r1SjOxEMr+aErWDNZZzX+bsOl3tU/KhQDWaD4E
m1yn7AWs13f9fBKe+BCnKFObwBfYWQT3NQ6fE6Qh6vlTo+Ok/TetA+fT1KQiHm4OXcBhrAwraegl
WheQrqZvUOVmXBrqnlwubCFMchOKoC76z63HbPuM9pNJDNfFoKN7y6XWQLeLJnLoSPFWNuwPCppe
UOl9AdlxfDzb4M26VwAygMhjR5tUuEgYpkytVV9gZi6xeMofZ/8TlA5F9H/Hc/koCxULYrqqHOty
LUSCAfP5icTQ5lkvb4eZRA5/ykngFe3CuNmW8ogXOGTl9eHdA11RNBeM7WjEuRvb7PZde7cOIu05
pJbUO7d95UvMF2kQL7FOGHySAtqoNJjVSu2cRBatCrUdf/a0oNqQEveE9mvSHmBbouR6nFj/w9O3
Yl89fCuZ9ePSoQAcRIjBK8cotVXPF017kaEwbKz3Kxk1QQn8yDZGPMacKHZcWL62KrtIr+hKtI/x
y3ZUsRwT3x0u+tEpXIobp0LzkPUkrWahfag+5iQs5JPgEEUGtCK/yWxD0N4TTZ/jfe19CHS94Pky
SL1nRtJD1MisMmcStRxyNbZprsY5UhtHhf7ij7gvoZS3m8JwL8JQ1teshqR7CvqfcPqIpXXet5Yr
6XbGyudhJtew5Y0GGPTZvMzfETQByU56RDh2l+5D/BUDvO0A0J6sLdE1juO/AwlHmLplpLRkH+OG
Bcb5gFeYyxt7844sXH97eQXAKCYWvsZrmFahJ5C+LTdnhVD/Nfjh+q/ZtG8KqQ2RhC+M7J2PZ2dd
S0N1GB1AKKUMRSP6Rg8dIb+mViWYRSLCw1nxFuhKn+bcbrNIs4yWdgHno73OUqODN3paCBr2G9P3
+Zgb6KS+ghHPzq9lmev01VLJZznbjwxZbj99v4gScTQ9CV/GtvTQ7cKw43saWIc/UGMJe5iY9pbf
6O89BnCxB2ht3rtFqgj5R0FcRONVu3LfR42RiWRQYphGqm6VL3H1goEAnmT/vCICNYZZYJkjk6sO
LHFPWGmpBeAcM9tkRyc8JTkynS6B1vsrdQYakQgMEt9HOmkOF+MwESsUd4Np8OZ80+LdhR8Nrlsj
RRg43UNeuscHx6c5rTl9UoKnsYznb5Nwd2EWWfJQjqa+7qbJm1uQlTsnyxd8EVV27D03alWbDAdV
HP2B9c2bAT+MzqZ6NYOTAYqCZc/fitTfWCdTO6MrHzWytg0VUf0yA76X2MsE7C5XcTvFuhuhbhOf
q0izNbKGVzQQFDS3U/ESkpEAtdWMe0uKYfqEAK9Jx6EZsw2AxAGXuaB8WFH6xeZyU4UhaADwRZr/
8Z1bAKteou33UNs2h6CajA0SAPWWOnR5N6aqtahLc+Bqgkitv5tEg9m/JbTSWuI60eJDTIlTUjVA
D3vTAP9M3iYcb/FY4Tv27Gv3atlVnNK36CKC3V9EBytFESovYZMPkDC8QTtMwwvSzYS5LkSzCMMh
ZcOD8hYwr5v9EV8UvoAbVOxnMhMmlizf/4ut8lqPp84TxF17gNTYdQUAHQjuA+HviB75U040gQcA
2ntXG0zorTEqXcflDxf9XuWq+zrxoX946HjHUifDABnswHF+Aau20jPJfB8kAt68ZgtWdfFjt3h6
MfN1AmjPNYVxEtfW1B/KJL2nRW+nTtqq61FSTjETaGosWyn8+kesz8C6hKknllaYshOm6+ZCDbsr
0/lkTgvYpJAT8wTDG5muvHeEiE61oRd/GJTzihraSxVMS6EQJOKT0ZRA83uoMyqQSJb88cns7oxi
HvjBfQlvKN/DzyBWtSS5UNuPetnssZjGhHb+AqNyAc8dkRPrzegKNVMdsqqmN4ysC7EMAjf9ylY2
IctjxGtxn8OeLQF9dN1tJqInGDv8IFgyibWR1tO0qYeC577osMvRduZRotsoZhlU/lOF+6XYM6xJ
JHWPr8zfRSUOIum5aEv2zKTqZzVJ++9vEspXyyGkDdyMR95Vz/uwIptipgUpbPEwmY2HzfZi3Dg1
0OmuspA/AIwypsOlVpvUQ9Csnb5yFaOj/Nm0usfWk3SKqEVp3ch7uVVVMuMvKvhXhz6BG7cPIuaz
3Q7bS+eyvycl3MJv1kBiEil05VMoSZr2UW9aesvXJqkEmOW+KkUB2viD9Yv8BFN1QnQARbMcKQsQ
qaOnP4Ki1R2dUTKAgV8JquucORFuLe0b0yLYUO5M+UtMQ1+U40vusJaBcaHUfYrPY7bGJAURxoFk
chaH+KqLboZNzSmLRIWMO7qe5lxq7Cxr9oN0Ulv+sSj0FFGEJyl214ueNdC7L8FzMtOrIrRi5Qop
HadTq13BFzx6JDdP8aum6lYWrj7qNPoc6Wjd9bKiCsqQDgXjOumV48PI1Ga7zpiVb+7e6nNIdb1T
K0mvvYR47QeoeghZm/+MwfiUCsdJjogXaltMXjDfguwjDGyiTpvcoUZklSBMd+9R3IfRSGzujRy7
5lCuZeuKl1A4kzLeQIy0BffEqGS46W5KWcHcEPLs49Xkgq/G4PXj8ThIhJs9Gkki5Y6opYxWN9wG
YxhOkQ4gkaAI3Bfc70nWT4GhMwoG7blu/hXXd4waxVLntR4xBqPXI4vneJdJz3NytcrpozPcemkL
hvE3nxcWYZndD1YtwGJINJvx7Voav/ZeaZzBue/xtaMp0RKaW0rOliqusPnJOukZBsut5vC8oHm5
/7sG/tZWMWBSW1abLFu9P2tLJwt5zoPeWCxb5AW2/Bke0hvgq93B+wybrbPkKhkKG+cYaiWCOu4C
bcrkD//G6k5OAMSaQf+JCpDqIdWi1EmfNThlxYPcc1eDzxOjdkw/Ah9yAj5lSXsnzeg9moHlgPWS
nP8a2pUfvbQHpd0wg1cuF29F1vPBn5bSgwy5+stRJyGaOhq5AGzJjkOmiO2LkkCWVf4gG0UoIXd+
aSs8cZqYVl9wsdSdENbDC7H7ZO9S+dSCLCrja/bva1/1L6havDvFYBu7ZUZYl48C2cIh6yQzG8r/
cv1EGiYrSAvMeK72UF4mkxlpQK7tXGGMJErF/AjJ9vIm/CAohzn/5Ea3yJg0ZJFYhFluTDlduzSZ
+jf/QfXyvFP4qUNSQor62A0YvftjXwJz
`protect end_protected
