`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
iZLsMvzYxl7UVy1qksvkvq5F+Ify2SXhnMnnJ/du+/+lFNPcpRV85a6SGmwM6fvsxk4pSjCeXNqm
2Ubaqc2mxg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UQbYQdAeJSkAWsX/lPzNC6scSmoXfZDV630edORPPzNEh+jybSRTRuuCaJ9IXoT8iVzvKCKAR1yN
QkGWpPRiEhJ8OXTA25I6IbsZmaXiflvO7MupLibfpUyj+L07fDiYsePPt/BcqO3yBiBVoAFdeYK5
bHnbL/fUnG88jJMY1eU=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jo9ap/fNrLfE+dxA6JJ3KSul8laZvan6VHTnDDxOe3VXOVXVzPItuuJ+HusOSfsZLkUytmA15aSV
gQx0uKf0NY0nTPRNwHWnkZUKsbQV9FajRG4878AVzw5XHuTJkFAvxIPDDwu9jf0nG5nOwwTkzT0V
ClkcaV/NpzSV4a2VqXmiwYfjW9T4ZEoYD2q4rj2VX1UBSEx2MRwzHhNXVqPehN2ru+JQwa20DVXR
91X5ca88BMGlJnX4WBOcILqinT/DJI4N1hOdHWHV1b8mB8ZCFUo0zjughurelEbpSlDcZ4XttFAA
OLd6KUNcfzo0hKl3nKHyMniA3eWaRRwEaJY4hA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Q5qiDOYtq8Tp69As1Qua6kt5SXK/cT5jdULhAEbBlM3hiEyy4+/g8+S0Ob0CDq4WqTPZoHuOD42x
Op41NLGOUOVWsd/2ZDrVnl+EyL5t5ssooOOVoeeENd2/QDT6adpfIuZhe3NsaOSPXog98P6+Qqql
aB4I49m3Bn5DrDo/OgA=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YrqWkZu8lZKf5FNnOeiWG9Fb5eUlWvcESSzA4pHZpVvfz826Teg/X/ss4D0XHwYz3c1ROB/4YzaT
E83zLtZGbVxgSYu9zePNM+vf0omIhlPKdmjPDXw0Em2CeCNjaX8FnbMcYCzBE1YGEQvyIPV94IkM
+lPMnVgXF+JBfJy32LSRLflMPZq7u+Qn+RNb/Ven7G5EwGctMVH9l73DTRnFIzrgMSd8hAGbCv67
N3XNuuL28QrI+hMBvbYU4GrpADMlkJKb5AMFyfwRIZTyF3gT3fKeLJB84NCehjVd9Pd+cdiZ8Mb9
fEXz2PbKgThYgep2dHDkj366YO9rSXHUKg9P3g==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EIDbDab5qqu2YU2pLrvR3jvVJUgPeodJJCXWJka2eBuhFJdVaVun4knhjbB22KTQ8R224R4UgRZ7
oairxCoLr6zBMiZtYQb3TcGEhiWqLweaDqnder7RyMrqY9x1MothAHafdQtczJsyEp9Ut1BFWZjc
wlQxG10iksWTm4BQxcLG1LkX8A2hC5YBh++XA7nEW5aOS5rRU81Ogfq891N5doFKjLywqN6jB3kN
0Gqhu1j3JdYEBObO0mmnC7DxGLRjCEW0oUx5JdMyZbAUHIYUP/71YzFGg+Hk3I5Hw0erCNc8Lypb
JnFE6otWjktlATPfEms+jVIIQvb9NxTvxD3qhg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 288720)
`protect data_block
nILhyQsDtKRKZmw2rzM+0kzJSezy9woi4CyeS53w9KKv8Lde5+SKQJfI6qW0TCtAhs0JcwhiohtJ
hGtVeKD4dWXcJ0l5tuS/0fRMbedEJaQ/hZbDaKvKqy9ngCqvYgWLan2LypmeysPM16a395wgdf8z
ByzvQe+efOyr+5ud2InR9QnlcCF2/NgMzSjHHN3VgYfyr145m6S7VcvZYeDGjuQLKTYx3lmR6v0b
rxIuy32ySGNsXYCoizbQaJVoPnCSNdi+HZIpyEBB/3kSYtMmact0xAlgG96DXxvYkxSA/o453lOq
yfNNCOohcni8hIM2cRXevw2Zy2HlJ0xjJJd7ZvWTcDeibHBz3CLBGLRkik6kbUGnu0+GuoP3vu7E
zhEY+x78kQbWVMUUWUzT7Wa50Rh95R/CbGF1Qk46F2rNMjC3fm/H5oHTjO6TwMq/uwefc88WQbKx
OIKEwHy4A0pu9n/zPgN/E5bsGkdweFsptxUNaoMXkHc8WA1mihunYIdlJ9v7V0hwjI60diSiMsIa
CsDZkzezACE03d2HRxInMR24E9PRPS7xkk9EEVr6flIF5CRcf/4uLUsnLZPdX0UYD8dSQvbnM5a2
8FUjh6xrCPTiy4rfODoc7oObfn2k+OmJI4AYD8FjV+4+I+Vepp3EbQmVAoBO4DL8VXAdL2UVSmuL
PjYDoiJ0Y5GvAcCpEEHnUn2OJrsZdVCWVmjlxC6HihG+KmO55kOnY5FrDiWJ8jUnXcCPVlG/1nFn
nRBX1U0vtCDlVxX2ZPFRAJn+47+bYscQ+eGGWQbT66vJTq0aO/h85vDqElA9HbUsVABT1Mchqc1B
zGfPcxmp8+5f2/btf+actsSmFyyGjEK2F5BQlyclCA3f4HVaGgrYX3TImEbz5T0py/kRoYgApsWu
/9VNXDtPz8Pns8o6ZYzxQ9AxNR0nQR68mdUmwaM8JdzcZ3vxWuIHnkGPEifLHu9+KiAkd+XmW20a
sw8+QH/R1WOFHsz+yD2BrtwgdRHX+JQ0VMz4tkx3HBJV86dz+ReBgfLASFVeiTKAY3eioBA5kABY
Jtn9wJXXM9Hsf6eId236nOADsJJ9AgfsEjEKuAg+bnqXdDWmg6Z1I5fSvsLfSlqqbeFvn3nRYsVp
/Vw3ZOAHhQAigIm2yp/7UFAuz3eKR32Z+7sWovHTeMC2P50yDTHPkVmK6/yyIVtmu7sTIgI0wjt5
kCCTBks4sIHAS8TFi9WLyV3UmKFbLEA6t/dR0ol1ZVDHjNndwrQPs4CIGSq7kbGApuJxIElp5X3H
IK9V8W1xc9eQ1Mvx4RNLVKpJqWyzGU3NXU8bVMHekIChumrmEJohCUFlSgCFGwr1BYNvRruVx4Ym
vK+WGYvVKWNO3CZYBMPIHZRZDnyQCTd65mROm55OcNoeUukuPg2tPwn10hEu2nbj2jrFKvzYtcU4
0hVrSbGQPgm3nx0vY3YOfqJixItGNFQbqqtstpyB2woratzb4eDzVFVcINqxWcR2wWDHu4skpY/7
cnA0u70uX6VsSUlqtJITDNftQJwppg9sLfPxkopDwu66/K56lFfKtANhaZkpel2FgbUdQ2YCrnQL
Ubym3k0SCBgeDC2PGP5G2TkE7Iy9emND+/G/Qo3qf21xPA46FgcShYcaeBOdo8wEpoLViJY4UTE1
7sAap3AFPiVFbuoznfwTO8iwLH8uEhi8QON4wR+Jkr6PaYS61Ui1Uif/QH2Vs3txr9ARdoF9T+ZZ
S9j7M54MkgFLQPyIoaK9kd80Xjhcki9wZaGG6moammqpK6GphWgHqvZfoladaE3FvuFwv1MCI22j
i+5d4Akr1j2kNIIuK4TULTseGrrAcX1T/tI9beAOPKM0V6r7nIWugi/rAlxvycajmnvFUxOQ/rV3
UDNu/Ut+ZoVW9iEOKDgmuAyEMZZQGH4FVkLl8bgIXEe0qKaKPB04YlxEeMv/pR9pPrs2yG1jUYXg
fJOP26OL/8lNm3RJ19KzqGKuGtICjx5G3LTwAyg6/UsckvhGBGLsEysO/Y6dkWuMzjUnsDa8kHSN
rE2kxdJzvQeX4IL5o3C8wmPlZFhL+GBpgwa8LW7IiHrUTmt8js6u5zqD1p9g6tnQTg3VsSfA2kCI
wRTWe/4Wor9ddVUKIn7ykY0jtixHlcKNhMUq6sBPNYuy1my/2aybOMKPtwxNSVPFobupblVSa5LZ
BFHJq0LpHhxk/s4Znw1t8v91PUdGn4UymuzJfJ1lejw/lNDwX153ZnWAjKGQoZ+/4Q7XT5mw3xXN
rvGspc19XbZYUuipwKnNRYr1A/+5D8b21YhFT+fcVqubdNJKuS9g+6xSGAGu/gwNP2rsfY6hptJO
Z1A/E5We7JEXp0oA4d14tbfGra7YJMS0yV8/WqO4A/v/EWrDq6UtXeHzILTyGrGhD8ZZFRCHNPji
+P/ucrTutqhOtjwn5nkDhQ+ZzfTlqz47zwZ3aHI8kRRVS/gtShVeX3vgcDFfLL1DyZhJAhhgelOf
KTBPqBmGyifhkPsJp3Pawx9pxXAp5qbYX4iCQV6or7euE05YXjxh0pJXeMh2Sf2FWRWpOljxKMiC
3jPK4Vr2s+Ib8Djc/0meo+0w6v1DP8PiVT+uG/RTa3qKsJ4SIZmE9xWV1GdED5EtP4zYDsEe3GB6
d6DyAwgu7KngsSFCZn9M1R6OU0/V79g4nJZ0exjQ0rtPPg9IVmhtvx3XQqmcmlU6AH3S40fRHQBe
ymjJhWGbssdxHkYwBefbJacgxIfX1XExrFblr8Q6DSrf8fUGWWFmb2zMip7g6xkwxku1VMbpUedx
lvBYSSqgfW2jpz7kb8xXQSNQxkb3PNtannGKdKB3dEEvDrfjejvFrUbjFW8+VEdCieyx/zaov8rM
UH0/gG0/x5WNpJJn/v3rx/irE3n+VqlB+fVJx0N9KyE0nMzEgzzFSvlB+bXis6iWmH1EldYW94rt
Ib62lfUDb4Q6M3YG0KM0eR2CCJ8dcCsb/87qBR9Z5nLq0grYgttUYUA3lDegiohAh5bj/Jsw7eiz
fjQxquo+HedOhuvvzvJ48JF3meCNaiZAsIlNe6ib+k1rjbEcDNU5FpbQogZ8h9acV+jdojMEcHv4
cL7WYLk1cltbxrsu5CbCCl8s4wT5OQCP6UYiaWQ0G96cl16XG0BLLBp3d4JdLCShcNmYATFpi7gW
s4IjuTV1WiDUkRqXK9woRB/f4oyE83pDRALgcmuu+ZPoNVRgBHQvMNQ2dhhBZ0wk728AfYbU8Y4i
tW5Ht9AXzZMnZrXN+9bbMlp4JNzqhUUikUJu410pgVqRg+/8nhLrJNO8uPKSWGf8wxMhnXyNXIb5
9X6UfuPyVYGOxVW2X0vlYgBk2Bak2MpoBXSk3QicIgVwfDZVJGiTo7UY9qegSGOhyiZBGlh8h5Ys
YnjEFISgyJz/1Fj8UMxaJxQeRR42m7TmQ+1JdB5zL1ZgosVRnXVOjkRf1KGmMrqMgerfho6WIM0a
HmLLiguz/viWzlqSU5unMV6cO4SWiCkk0RGUIhmjxo4ayUNaly4RHI0dPt7zsv/LPzDTKzOv30A/
SAkfsfp99TOeLFQLxLSXD4u5qUUxl4yOT9EZYpK9smysTa66Acybx/BuOF7XGBxAbizc5muIVJTo
quFNeWdzZMnNoiM4iPhCzlK2+UiGMmVZqLLXSRUwBeWxsi/iCfVNtCZawGRIaB7bt9k8YSGDPZRI
FKrFJNoGoZtis1C5cr9AckMIjMoQTWlvPYMnjfn/HXTOmNqH06/1249gFpDNwoyNSr09ngEzfcZ4
E8qE8hwiABgKcKHHZrgFNiUapuKpVPTOOKqD4UhjB3gOKy3pKuVJPwAn6eK0quP7F+GpTje3FEb3
W03bHXSmvkqJOHiUVSa6cVPXije3XOGyul3LwV6ZYeeK9pMs748nRGlDUMf08KefWs33pHn8mKDz
Xcl5uAFlMBFH3BgiR/OW9+BW5+62T9KjpcDrwRUDa7XzyZb3U+zXwLPZ2AwhlZLZimfhxQTAEze/
4hO9+8TbLiJicpGxkKAam7PZ7rb1hDmGGIVBnP/1wBmcMdBFWnOmBiBQuiE1MfFRfYZaKSz3AD4o
OkPpCbCywsD2VLL1QcVyfFXL2THWX4UcCSxHx5EZZyRE5poqHAeYwJUiuI+oVyQXdJeE9cNxY8T+
Jmqa1697kabbLu1mbRfQdvlO1oXVnQRSP6WWc0l+W/1qBWHTQhTgqjSAPCd3Gh6CNCCAbKQFS5Im
7/5s40mpMg8GozHGFILcqv6bi9JwH6xhpstrpiHaNtp66rbrPGvnN6V99VsJnzUPmf8rp+fbtrTq
s1hxLkd8SQiSp49+4EJrp5bUKy4wVITpZ+sz6Z+ow4YgTsBxhSEPxlS1viWrc5oKW5TcFB0Opzfl
v1dSnZZTpHXnbCpwLh7Cra8xdGF5pb/mLnZg3Csf0IhV0mB/2oK4BxQDBagqmDKcd1VJvWJu9EEN
RX9zVU4zp/G5Luww7pXwEgJOlv559jP6ptzU1UXiSPpQBiOVI6VX4Vva4p2oJJNpYM8IPQYpCI7A
JEa84ku7iihfGoaPOZ53pJLRAUkDkdc84I+MRpDewqAjiX4GubWVlL+4WiKcgAUCGOE3WPvZf9ee
dI5Uslo9QeYJluQLTW4HFI3v2YJptNFg14nCfXcsvs6sy81YeGKTy/oUSlIqlVOlRQq8h4ugo6v7
ilHEQ348mNIKQ0Od+49xq9PxV0ALBPkTHF10GTaNlz++Tcbwie4WcxyqKE5qUrxPqyLZIYGTXIl/
1Ou4bGAIQm41CUDQzCwFlYC0GrXCHSM8e4rZS8WRrLcA5SYwybsuvwJLEcm1mQa87DCrbSYrTaxa
cVzU54UOJ7z4FjX+vCT83gcZ6nXQiNWt+ivRSJYjF8j83mZ2bJJHUuDSYi00wiqk7/F4pBDWQJAJ
R7919ji7hL1wP4sw0tcotUTiG/ibrtolbjrEE0+Gpemxu5vm83x4wqcq83NTtpd7i2iHiNT1PCIf
tc8N9u+KpviAYMkXrZ3CyBX7/desVRK6zthpGrIk1ikhyWDqCcme/I3L5e68JG3GuBQLbiGben/j
7oHuX4+lGP3Jo1Kd9PeKONKNF/W5sXhJ/YHDeQ8fPWT89CSxmbLKo5qgGfy6nESyr4CzrnKSBy/p
BdNa2RWadkgZcZRdrzmDhWYCxxEigtu9tUyoXSEO4F4r3jv5OpPRhB9hUjPc3LjjCRCCi98nKnEK
Fo2ohNhr0sOTfV+z377fzcKJCuUZsFtRrAPn0+8Vd2y2DQLpwd/mkm8FwTOdmf2SF17ci39nqTDA
JOOtq6/MNz9GSTWNWp1PysOOzyLMT+k34S4S4CAnbsrP58hzcd99QZ1jqfoUBEtLpCW2pKSOJtVS
RUIFV7uMN80fufPj32Tt4A4131r8yKAbDjO9H3P9p2PnprWwhfn1crc+q1p3y4iu0u99xr0V0YT9
XdDJQbOE7Iu53PnCOoX4wlN3twQWfFhIG9Bxk295AZB7CbYrCdUZLvyZFgTFJB2W/L4FRHbhs4FA
1b6swPDBqUAzJVwE/QjSd9BA9o0jofCcGH+ej+1kXyG/4qDsKhuUvKZ01ck8FtzD3qeX8mmnuB8C
oisFh3KslfG21H3yojP1jXk6wZcXz7WMOVQSNQoTI7FtQvLpt0SiRX/kRkBwb3n6Bx/nukQl/DVZ
pGJhbslMqehddU6+WR1v/ZeZPbtadA+WlOb+zNk7sjR0qn8hsaCvS0e+vN3bAERiB/hkzHbkMe47
wnzXxJvXZ6u8p/KQndL1Z2ePVMd9ordnLE+jhm5xFLbRfcgUxlmnoeW1Tv49ZPZTPjSmoi+aHlVW
gb0teUi9+3FSNVnvZ+qF1X1OP3dcgmoYkFahpYtxZrEvpafZBx2zwftABV/010Wrwm8OJoBYYhzQ
ztNHgFpvVMHazk7ODZaHhgVgHu1JdtTNfCOh2PF9YsWv8VII9SulGnLFYxpDOsMSbe6bwsv9NQkN
kaH1J3oS6amwvnbaZIR5G8jZkihbUxEjvwioIisBKF1Pwsplc3s8NSg5s7YIsHQWa3botShCWHIr
WoPF8KTjOWkDmmaDTrASj17T0LErDWS6PUuHxbU3ffGmKM++e+Mp/xwIGeIUnGzHABJM2m3E+pSS
cYWjILucH74I+ZXewoDHoMIjYe1Pv6uL+oS7Ql0GNviUh4ww/ySRzneT4zPovx7Iyk6DXvgsh8Ua
ioemGRRt065loS1Ur7zh+CupdZqvcdOhM8Ta8SZBToBuFFmuOCm44jLtdg9zBqamAy96F2VBhcw0
dfLOzZePvEWnbKCviqtMx2L+r7elt3aug1kUY5O4cqPSnw0tKQFQEvEQLgBhAkveev8/kr6lB3LF
LX6vu95SJliSppLf7lmU455MRWqNHiBI0GgyJ4zN+CyMh/umGNa3KFU1gIvpeyCD/mPMZQFy0kYy
ZjVS6lFGctJ8BLx7XLdq5kF/ck8shY16QpvC2h8JbxLCY4L7uXR5MwlZONPXqyObk0ecCRN+8Znn
MCbjAloD8UXSmMLFuOuwWEY7CkTyEYhn373rD2bAfuN8pPilLm6Fj0GLr/oGUBblothmwCBwtekx
9pnbaCEGkj3HxqS1QfVZCvVg9QRTA/zrMnCZxOHjR6YHafWNlXelSlk4NjZzyXipf05rfkVvDEt9
AlFuAahvJvXN0d3moIkNU+fO2c1wPGrEcQE5XI3fRtjA+BEJlo8zSm3q55tUaQH6TGscC0VdEvDl
1h3uHp5xnQQkzdGVX2gTe+OM8nfYJjnXrm5SHwsuAr2shuc9LLErZShqWlWXaJqOcmiXuhTCKrbP
XlLvlZMdBDw3oElWVEsC5V0MhSrKvZrH39VZPfISeHIc3i5xz2bWJuotDsi+daYoAdVwxwRSK9d0
HEdiGl4uLOHRX3BEthK2sePbd5zocmf9mN2RIovWolAjtoPDASvVg+NIJfaxAvfq7NO/IZUy2jaD
WR2p8C3/f/qDmO548zWkwDTB6Q+joyYo5XHoGO7Ea8trjVv+iPkVNElV86PgC84frX4bQYlWmFjX
X6pw/d7EAEkktyXgzdPdll4Yk0wl1kohbBdZE8hFa3DZKXzHUw5VRgTuAphwjpL8YXbfTwzL5SQk
m1Lwhg5lZpQQw1R5rSwoNhBvEHf/Ra1SiUFot5nd4F4yBEE0camhMc2rg+zEkHJYjJDF4ruLdOtu
jzronwYRz2VQ3tW5V1DxZAUlQ8iyM8Lb6SRaHBku730mrp9LAnTspZiGYnsNrREvz9mi9eLnDyMF
4wLuOX5siDicZUEuLsqXJBWxFIG+BaijpXADQEp3ZJqp3+N6kgTsagaqKD0XxQzGdplBoeCbUza+
iCS12ewFl3P9CTuCrO8ovTofsYKbCblNiUqjLeBb3s21q12pvCq1gdRBL8sbb16NSSpbwEHBkDPU
7Bghw2vHIMKn20XYvcZGBXqhcIaK8Byo/RakyDXOTXxXMBJ3MdK2suRlSWXIUGuRxAbhnO8YBaKv
ci2O4cajFCroZXdR+Xt12iudOPGVz25V3hmcYov4+whyU9Uxuc9xqDqrJEOLvtTV3/8HNLbBzqfZ
K7sF2JpmbnHl3PhfHkTzg7UNWemoJGoHM8yVmGXkgduD73GhL9J3wzOrYYzLgSXyjbohwzp/XDer
P4i+tdn7cNYKvLmjThNzTwtnh3DrfjVHPiGls7Ew+3SMad6RHwAqMqFkVapz9kcyJxXgqwPOXiK3
M8lpM5uaLDh8iu9Q2MAzpLnsctQDk57A1g6HRe/MGIBJkUVPIg/9o60iCVNAT3tMePAon2DsB9Lt
Pb6seM+QtiLzmKtvdXzdXhjr/l8C3lSFUmHXaTIX5jNV/U3x3SmH2o39iVEeRnS0O1ay4cW4hGGZ
V3Dtcbq19W23A9LNmRbRgSCt7TRaexL9UvOHFNOI/1zQPIL17pQY7arUUrSAg/79ktwnnxDJjJah
78OGlJIkYirsMm9US92Xhv3vqcuttxPRGIPAVJWPXWee/sh4cf4UgBTG4MaKhVqcHgbBvVS4sJZV
bjUhFz9axGewjnUzrMconpIIF4wGMAHO1KymDtO5LK+MLIbEMfSnYQDfCZ2LPVHouWEhEO8UYqTa
6nqwdoMoKRcyzvZ3QJxRdA0mv5CBFKZBq5PLGk1bIgcIBQIyui+0UN2WdG2wPd52ilRtUGbKGQdK
382j/r8bFl/QdFTBzDuz/KeC1YYFvrd5+vzAxN/g49PAsGTMLFou0XVn8acD69n9jkBZDu7EfEQT
zi1NwqBhmgIi+gGvicBAN3wlkSPBC1ZVDHX3cDdkBbZzbVI2awR3hibr4r4QtPSOUm42CH2HdjsT
d6QQwQ13q1Eiwyuo5LSrVmemsSTtyMZHBBnZ1XGYV5Uyi3pxPMNCvxWUrbao7imQCDonsCW72k+z
HkiqYLv3d5zBAg4YlTAJicdfqpJVHefomizzxc9YQ/qo7scA2GYYFDQ7aFmfZiIjUnZH3rrj0CL1
mFy1Y1E6LymsLhWKvMJkl6T/Z5STIp16vLtdxcD3JOVa1I/0iz5coh9VNiyeH8iphGWHpM37MKGm
NfBzIRrURdb5nUSC0bQK9emfIkPGn0YevCrgnoQc4FRQpC7XbCkpsuCLhP5Rmh6QHwFlNB3Ybzwb
iHYA7z4eAvs5wcIpu6pFO/28uCKVRgJxVTz/jNCURfKoyeKSZOOFB0qt3qcwc6Q8md6W4tYme21u
UMIVkO4jcYDPRyCKoG3+KQ+4j1zHsQ03c+Se3DPBusyAtUHKnX45QLZu2B7C7bG1OuGqjLj4Sb6M
lg+ufenj0+kaLeS9EIofY8IBTlSwKJTdza1fkLCz6wO24FyffVHymNR9cdzUuqo3qVAybUHsD/mM
17s84gVVY0PaJFuempCbkvwANfrdXS61o8E06JIfQaR4TPvxWU/jByIKvf/FMX8KQB8w60a3l+1J
FGsWTT3fx6EA0sVUDUur+a+HMfTeNT3K1ShM304bAWqm52372YIyyN0XgwB1mBqRpjrYPEV9BSrS
5Yjvbwek//1iyPy+Prvd8/BSysCVZzDjtG9QpN/ZfSqoORKLn+hgyof6rr0DBXNxEBJCn3b0jGtI
OjXfzxM7cvQe43JQG63jGOezQ+aRjpIOE3QBF6LE2WL5m6FX5vleIiqpWOnVjsBfFNTDKdGN4/XH
+/8ByKednTyG3jTw9dom63tAYBFUuzifFH7J91O50HukDou7Z1n9nfybxQAqGSNS+RaPLswHWWAF
0Pj9bcI3LYfK2OrGZe8CQKMDZDXf/FpTozJVUjzvFrb1q8rSxiNzo57pRfrJuqwZ3MC91KzC3NAa
xuZdulQ8VdJXoOXNBz/zEYsqkI/1zZuoC/7T3CSRaZ4IlJkzZDN4nX4wGb8AD5nHmhAAc0twPk3U
t0mhw697vxe1loUmg6MPS7yC3tWpC9PobzhOhcOHy2bzX4Z6/fCbJ0pUZ5D1vzJYT3Qthg2iTxNR
qf68Bs9UXSD8+GK25kuZ1RC+n568j5MlxaCFaaKXztvtlk3FjgrriB40T1uRcGFQR6KNQ6dc3xIb
odOpQEkOsxD7x6uHZzef1j9MrGyXh4KXumlibTpmjGdTtl61ZKenBg1NIPPD25dKiW51/ohRW1F3
Ms5OhTnLk+gQnSxV5T3ORtH24L3r4XPc3j+LmHyuJug8VmPFAdG11CHlFMPysDdwZhNGnI+IOBdS
gc9+5v0zXl00GE1UATiQ7/Cmedy4qjvku4mkGVV4+wJ/lkyPvshkqb7SOZBaSaVhhRMX+tnpmwxx
6OJf6kwOoA2LevOZ5nWb/6Cx0h4dbkd1KeQ/Mv8hePSXhevgMRRiRyDh2SM0IUbrt5xgnzFxijNL
pJROLacU21g+b4PQYHqahpcKQ4gcX3Y6IZkZ7PfBFBF0E07iG66pxqn2x0prbJS3P+/mJgdzoKjs
KwMZNRPPpAy4Vr2tzwMTlEPbRqtwCcNEIbP15ZsQBm8wilLthvR8UVfwpRtjPpev9glxwPIb3qnl
MvS8m4H67a8vYDcTcUbn0CGTVDZhs3ndstGbe1LBXInv4QBm+bF2N+EYNm9arEleGiY6WwwtvPWf
yC1m2/4oXB2vUUs5HA/McEyvx+amJDu6OZQIr/yWt7uss4GHxk1Fvi/UEv1onrIcJfEDxPKPBQxe
F44T4ovRCB3RTYAutTrfqjmX1KGamdlBOEjP61nqZZHWJxBOryt6e/Kz8f1JJqv4x5bnuYLjL4JM
+EKTAPeuoWokJ+mmtR3veYSnFkvTuYCYzqSloT7XMWkJMaKyuowX2+5u4XwCIFtV5uMjfPJMDp6E
t67HWNAG9p63GT9jewa8B9l+My4W9iqt78YGvOK8VXkEO0S3aex2IAVEDjwQ8xRmaqosNN6MGu5N
2hOvEIh98VaaLilStMVkvJpDMeL6TfVp1n3+jdFedxXlQ3DsxLEJTH02HRgAiDsiChBlD2+ecuFw
v5gPYzWTObgLogY3eLVjv9Rm3YPo9/58FMdZp8DHIzQYukqLUCEtnULJTQqPa4uCV4FCz6HuFPSz
VM2ZeAG1l2O4IPipJEwXigGFIWnDD2iHhq5b8hoaTMmtNGIBCyL5ELXvOaUU9zcjwsIk1bhhcswx
9wFhHWde8TSZYDi8daUxJJ1Uz1sM+mSFGqsiLRNtP1YnJFcFAxvmUnEDHBDLNoiaEd/HFLCZsNNt
54rctuv22yt6+VJANAdyEUo+4QWP96FbwMIiBMWFP0vvcD3yda+CiyMXvxFPIqCoY2mwQR2D7kbn
ni5GY25ICFvncvlfoYUnxCnid6kNVqOBvvMarg4dFVcdWN0TTk0x8Wq0kSaHY9SwLWtZPMeSlkrN
IHlrssn3PXxZkFvpXSi31ZR+fqh1iDmgv2dwryJi5ELIXy1FCt7Yt6Ugw7lIg2LMv6fA1IoT96ho
UMkDmzRAA6MXQkvu9T49ZW4GZgejHa8kT3BGIQ2VZWuktEWe7zEkS498WzHwWVzdkmfBrVWP8OFh
+Vwr7SMAIBxguR/MCQ+SDaFNi3y4qRJBwIeqvGxRboMFnuS6uwAdi8aJHdHGIBmKZvsdmG5gNsl+
Cuq81Y+C2s2Ch5VSzc5/CjROzFa2ftYnml7RA6Dx+Ge3UmoH7GppgTiYl1FbMOwkqQEfyCsauTSJ
yy5IWHeLml6l7Fnk0JX5a1raFg5NH/I7jPvwVlnJyRMK+ruA0c47LArKNu8ubSOVdlgBrW57vYXh
fgkyfnCOU6VjjYadw356XI4HfE7WAHV4HR+oKzE+lwTuqq9ZbbKiCR8Ro9ysCG50X8II6vUWwBOe
gUFBl2L3OA0xSY4+NedSaLtw8Hcbd+3AqNs4WY4WZk02AMSy5Cb57BVTWkbpyZx3aenhfux/Ej6R
1o21F/C+JcMAHzKAsolLInUAasEraMTn5xDR4OzxcHaJhtg5FKcynfKpORKp5h98qpBtwGU/dGLA
eDgsrK/qDUJb8XUOw7Y1CqDFOfbGCCdryPJ9F2JYGCPETCDI8vRQAQugdQCKeYfETZ1cfa9puDdN
6lI2s68o2gHu5XcV0TP4iKFndZSsZL4xjoDNDdEXJ0L2j98Jdp87xBTzaE0j4KjAU1KrrCbKf0Bl
FvuEPlUqNl6DDLbBjcv7re63AuSaP+zf8CBFCTZ6oS/gMEebpkwIxp/Vz+YJ9ngj5Ohe+ttOQGlX
MbZoLH0zwcXnqYjkusoJaK/+fq8h2XMdSSGKTMh2KbE68+NhEEKtp5anPszHHR+K6GEHiOonSf+B
1iRumHjAEG41i9umDfdfQGbRa2Az27FP5eYI/mZNk4LyqvrlNvT6gyIbReQbsThAFIrn2hjIeTb7
umpuC5KUKjuE0N0jK+NuOf7Tlte2GvNACDeDqFFfZLAXJluz+DfA7uPWM67QzCjHKUXHqVQWWu1D
Peoq13UTzfbYqBZp6yYqf7P/eLw5CFKgfyhkI4cTYfjq/yQuXWuKwldVeIZCeFfMaSZqFrdIaci+
8qdGYoColZRxHHigYDwd1suPxNeY+/gNs2IfnywixBrMNiVf1ihql5v+J4sCIQTQiRKOyMqLMDzy
ahe4Ckr4aNkdCaxOg2EVPszo5HJ5sj9VArpEWQo/hjr+uDRcOw6bzV1JpLcK2sxK7TDRzmY/R3si
fpQYSVfLPpkf7QSGD16cAIgw2Nq9c5uSWSoE8zUimoWhfOsOfw4I7F1QB7L9bc3v9PQ++fangcX6
+rSSCkMptQR4rkvSjy8cfVyUy6AJwq0piEP7lCeperTXOqggqa0w2mQqDFkwQnQ9qV7EzpC/B5mW
Ku8nLkuHfNL9U4T8G1mhbq6rde1y8fm2DJhSt8zuGJp0qwoydZmTelKdnoFSkB9bwi83x0WBCeg1
Mr17a3YPsXFxZjnciuw1dKSeO4czwwppepJ2J16LUMJFpnvJ/zu1Nezr9mWjb9Epr9WmRv9806Yy
1+1VftRFfl0Q/0yIvh0LGhy9UDZyqo1stYR5zdqw0jWLEt4fzHz9bu72tCkczk4IOoy6AEYdXyr+
WI3kgmrZFEiaxU0OthmBKdw2N2X1k1wWciz1/0VQsbytXHEPf7Rc7EQE9/3I0b6p7dasQpGAY6kB
aUKNAeyFmowk+PARKf7waj6jdxXcENDXbC5YPSBL4Y/7E/E0mhZ7YuZmv42JTbSz2VDmy/ebOIkU
gp8C4ItrTGNYcXXoEb3pBfQauPSZPWvHdxwwj+vIwasTBf5rpXYE6pq6LvzYX4lpcnNjjLHzo0ps
8/uE0E+x9AhxjoRPyKSpqP69O56PgMHcPqZDUI5P6UckOgtMrPwsD4ZxEtu+3WUb2fi79UWngQ1L
/r6eqIv5t5uovp3FIv1+tGx2LUIqSsOigqtBK4JAFdwuEA6oPCgAonrW1iJDPgMHWRlvCcX5E/86
1lPtYLnHN/A2hnV7uYtqTO4bJACU5As0eAs5P2b8vW+0tBz/yhQiwU47x0L1iXXv6yADsOoj1xs7
jo2uVbGIPKqBkmj+J3hUfg08aDxCDWC4nmUQr3gMYzgmBrfZYaaJR7yr0gkxJF/BMMkd2mk3SRhP
0gHgMJesMCu0FWrgxFJs8efxgSKtVkpB1D5jyuYawkATgbaZ3UwSkgDx+SEyjTrvuNVzro2Pm+ZS
aO/m2xB+sHnO+XCR7MxYfQTlwM6c1tJUYqj4wu0JXYZnj2vueyexWdLVxQE/xgFTQ2FBrAIaVdpS
EZglC+NJOmnQV0qygyYMTaP1W7V53dXL6Ol9hu373IQMRyboY7A0sqZFtPGU/2ROj8eRK/tdF4XK
nFr7OC0vdyi6GmoYRk65sHpjU5mgN9OHyHzCCIeoopEMK77NzMq1bVOJEZPQC5PBJPmnvoBQ8SYI
iTWH3tag33gRVe3bLmOAmqZTrzAsoVDwP3aPhtoNgJFSOe97+CdXquyuHpL7P1/2dJ8OWp5ydKKK
sZ8f/bSK+OUmjA03wQiRGj+tqL1wcQ4ckKbH3aLMm8kyJ3EjmlPatqaTMhSpYKm/idDR64SLRhyd
J3d+h6633mFiDOIUpvm+SjK9Ypy2K/KFVQWJmmBO2sj1CXNHO7HLcu3fBWYZovmZrK9sxd2XiA4e
hBIN3DDaLzYKP8u+7XcTWv7Fio6/fRqhG7MUxSuK3SpxxeR+/yEfoGcDb2Op8qWO9YfwVUo8S72z
OMAQUGHspepvY/61B49SNGVVye1MIslr9wQf6eO1dij2SyVNspqZevW4e+r2ebVkZNaU+2riRpNU
FBhpddFWOKEMKfgDetSCLCMdW8K+o9mC13d0IV7HibcpvufjZozEsg1k1gQc7/ujLapF7kjyFhtO
tT94fWxJ5TdNq/ZE12rSuNBnO4NMszBw6fo0TUdAjVM42w088nGzSjdLTdDln1Vy4xo1iBysmHod
xMO8ZB/WGnjNZBjozPsLjOeUWattufw06kTaTXX1lWWqVcJQvfU0p7sfcVHBmpXKFN3uNb7gbLCT
JJBwDmGuo5VBdNevszzG2XwUdsN+usPmvsiCoCyeXCJNTdCyrllh8F+nOcfqdzSsLtD/fJU4fjlo
k+GA0ZrjljM8YZd/X5Cn1HyG2YNU7+IiYr2yuif2FvtGk94JbHQgu5IT98buVWupdu6Zadj4v4TO
BXAra9JZgFS1FG2PhAADErv3kd55iAUPinNhn0T3I1k50wd7XFmONZmRqv5WRhxerEna9kF7xH6g
tkaUJZDa9Nhs+UfNjwNIypa/5e4WSNQhH14iHp0RDou90aqYd9kmk6y0iGFoFcMCnzgwiQ7VFdty
c5WNDFPXl1LHaa9WA4qwULJ4d/K+XCRO+PXxgpmstliVx99rSurEO1vJye0y8hpJQfVUmEDn4s9+
0xO/yg6JY06FhOx9DafvEYZ3hu5D7UaJkPOaDvnc4POwjrk5JF5To1uherVstz8MpQKXpGpLv0gX
P4Luclv8ysfYaWWnjX8jH9Zm333l7lOFaIEG9s3c1lPFaxWr3dg/tug57gx/KSAnZ8FXfFdCbq3w
zhhxxCgvP543r7tJx+Zx3FZbX0v5mCAyJnutTTM6bdSbjx8FPHI+BASnpErcHxi1R8cUJdx3E3Tv
KmtSRYNYsHybN9raT7xs+3XkIZ9hbInRZf0GjKIlyE9qa32cGgwpdDjR5hIRLEVsXrRBQN9Gpzce
fnpqPYCVMbGXPUfGRXhqTYFC4Pjc+9E6mQRiMnfaV7PvgnhENCKDbmTnUv+VuNlMw8/ZJOFIn21q
raDj/WBKrM9xNBYEaDBg0IqahU6AEQuaTHTujVXgbmga+KP7c7Q72N01Po+Zd0LDwBxUa/Wk36u2
l09HUMVJE203cQxpsr19y8EZXPZU5kdj1JlrXVwIvA7Htnp1rQNMPiCBas76rl8odejOI3lnAA1Q
u7rhVL31c0LlTi5f9WOgIohPeUuqHHNGSri1GB/dF/PmJ3FKBil90ctX7c9xDF1xezibY89CKgzv
5h3cYqVbo+0ujppOz/Mrl89QaTJMmFLByV1A+FSPiZL5+yuxasV9kONMmBDMEes+JmBAV+v4tcee
MD+zM9XGsjkgqllJOjHhsOtodsIIUedXmDvCLn2Oul36zsn6+K2HcEq1wTn4x7PeZyLflcmhxqv8
1sKhUrF4+k1NWGwGTjth1xBFGtpE/imJNrRe+oEK7gbtHYdKmqsCTpeLwbxya4OhifYRx5O6X1id
UBVD0/3uwc+JjeXJvLPjxtXh3RvWd3/djXXisefSLCIHFTNx0TVQmixFbR0EmYNRvsxjUivUu7R0
iISBOKQjzJBzLPPP6otK+vtFuMmNWNvNMUPk5Bt5uOi4Xuqi06BhTC8HZNneoJwN93m6fg3LCSp0
KE1IIpFVPzNnLuLiARZT42QIvhGMChlnRpVDYsMNgCbf8xzyffPlk1awlWTV2fESpXOX4JgH7Bld
6ZoFPfppc0Gug0ZR0RXQpMln1vKD7RXE31yNRDL/QZT2QiWCR9grNTcEoOWI7rAC2c5moWy9fBfr
L4jFTVyJYzFNe3tvyLke72M4u5p+TLhCQejkFxz8j9WX3hmpTmhbey9Iw0RcjzdaXA6BWSFf5OaB
uFUJLJCBce1DFWujljcSavFfMYY5VTBtlmKwNhRnLDF2N74KAB6fjSO7SW3cuZyiiGqbXZK5Rh37
x1vV6fxuLVZGe0dSAbTcPv+HnjrpO4p2M+RAVjVZDncZW7IQiqWD3Y3/5UPmpBVicw29N82izwrH
/5yCDvXDw5Yb6itlPNxPLL8icDwDkPjGJztMEli7rXfMH3WONAgIa+HrA6vnqz8n4Y/hZV3wK/Ez
hyEBs83GNYEKOFQ9czOp/CtvvayHyrqVcIVt0ooxb2a3ae+mSH/2UGy/bjGcuD7FZYIE4aHqTu13
ksbtq2dW0gXlV7XVQntLMQVrFFTZ0R/BNw0GVJ9FYhNLwkNx5hzVkZsjPI+xIlz351FbkC22DHiV
pGn4TIzH+rst9xhX8Zc0KBxihRVVPOlVy4mbocBLaFHJaOnwB1RBk8GjzMVOi/CuEKhLzeVkhAsR
YsfsYCMIFmUxQx9+rvAkY0c3MTXgjh4olGK6rX1sAyzWfwR/q6nkYY7/SKwNMcHai99CtCWHGDii
fZO7XRkfDfsKQMKfC4E/aw6dRb5qiI1z3uwl+0JhRDdvFK96lhdCV7Ir845kONZ4rksELd7286nV
SzyMMeTxyMxzCVhaU25QezazlIIOF6AWDPbpCUrMseZBc0aYlwKy5HdLWiqMis9IZjcWxZyopi9M
s/OeXBn8pi+Bd9474g3g2b3TVMsmE6ArCenc4oO9N74Oq4FB2sOK/UqtDIR0C82xCK6rcUelQGHs
mlkbdNDUFrB6X/dMP+jNEz4Wa/smc1mSQ+RJWpBsG+CYpRIdHkNQ9giFfdFp9x5kPG/OJbG0T0b6
7P2j4I1PFPLZpe2IlFNBFn4mQ2TEBGi1km+zkZUOVlWMfKSaWtd7ZekrkR2EofNHt2LTKHRYYays
oz7hAy2XopvoYy0XEqnspi1ZydvDx6Uad4vl5oKti+/pRK6DCxyf3KqohoFhtZGmJr98eL2WrDKg
QQfKPBKuDFvpyWvbCVz/b8sMInsIbCOri7lH9AFZvPlGPSuUHHWity7q/kikXvBz5AbkHlkDC0so
pz3k6i6V9OtLbfLhq5MJkmGXnY1tdqzvLuyLFZwl2fGILrze0NH+I5knBONj0uKwwdof32AboHYD
1BG/090GvTKH5k5C9NR62DXcQyd4vc9+z2BDclJt4A9sNmoCu6kC84gVf8/984kpP8OQLRrMLMiI
+ZMkCZQR6GvfRPfTIyv9Imbduh6sEQpazhW3fyjvT9R+LaD3xAr76j/1lqjBMKbq1DlcRdUzzmtl
0MpLmIEJKPcakqnYZ4Uc3oeCgVOzuV8KgzYBbnK9UcWE2O3OZvAr/VQAz8r1IXLOR+WkwLnGcU8m
EN0p2MTJKJeVA0D6MhMmtawXEDHlUilnDwrD3I7aUa1u6mv5vzOpViqbrKD5CbWzPh/0ELj4hHhk
7JlYn096hQQYX8JuWV6gE1SxxODLpAYtlGgVFiXeIO8p+1eFmW6Bx4K8gM3aU56zwH0aDKhoR48U
qJrbarGWPgNX3OztiWzZUezd1SA3hbhsu4xcomBV4yqaLM2IMjvzdTuqoo+BjeK/CkDzZ9mR6C+r
qnPgCVSJoNmm+mtEDq8j/ycu0FStA3rdm8+FHvtOEGC+rM89ZWaOXfEyY/F/SQ9tVAO3coprGjl7
UxXOhVjpWFqBdSz/qJSiRT5ltZxYPzB+LqNIm9KwqrIR+s6LzAuhh/wFdAsIxAyj2s10u84ZDwfk
i4oEuKoA+w6kLU+GATwOk/hCOHsbfGjc0JZCwufTR+HQAzTmEp7oczGQ3R/xxplxnnVsDyKA4RNP
ASWifWXl2iFyoEvMN227mqAV8AAaDh6/ML4FaX/vqI8ALGpjZ75rmG4fpT+wPOzTlD8azGMNrTRQ
yL1F9ouVTPqDCRIqjV+V1/ywl+kaLluFIE4zBFYqiFx8iOmBon50fW+BX0KWV8WWFCgkcMXJ15c4
0oeD4zf/wKISHLHPZ0jza8LMeN2aL7LtQ7KWdcVyEYEQm1tr6t8xDKlCWVc+cecoCOF+I6MuuvZb
zDRsJPfhl/4MwtSYuYWz0lMZKGhGqzzSwXXuovn/Mufg66/uzDAAeZK0vuvUCKzUIsKgil+z90TC
/0FFUDWHbcWAKglSdB9b4DAA1XID2plsx0/XN6r4Jy67hYonHZSNh2MC5VFZ9LJfl8O1s/V817ik
70Dbz3TV7AloCiHPKyBijiLBfKkTPt+4haF0ksrVdFooe4JXdokYT/jgHsKb01OfawJvUwPCwUqz
ULpxAhvpNmrJcz1p7iLkLY52r4X6V0agebtdtlhE4cR1MpIS64g8J0qVOmPfgqU0QV5w6SWdFR/o
eFsh8fF36S/wlI6FFR2JSQW56Ic/nyE3gr6hzeVx3iVFZjLUkYq0Yws52n0O0z3Q+TVtRCABrhBw
GkuY91BhW0qNrz9B6HsVgwrsB1K7tMmYfqAVNE10cPugZGJKx16+n17dGL8KKL/4O+qfuuMRCt44
1WBYf7avFpZpdiysMw5cPsS2X94lpGOGRPeECkMVWvwwL5+X46dH7zmJ1OWpREoVe2QrkktDRIin
vXH56SKTy1O6wJAt8qnzD1QgqZ0984CT+JPz/6smeGhdzu7teC8oANOpgPWeZRpLFgeXlpqCrEWG
Fl0dIs6P6yquxqDXR0yj19M+Zhwwd6MK76EBY88cZNO9PhVC6EUqfavkboO2Oi2MOeHC7jlYUcmf
sUAymuJzyXKB2bdGjedZJ6WIDY9hLjyx3sa4/ySRNa/mCllrmevvHDgLh6FGOn8EfZU4wDi3CR8J
b1u5li/+b4ZqBA80Q7Reh0LBJ1A2q7A43UwwfTzI8XhtyROH9v6oDNQUzOKhI+KxLHGnIgeQXjFk
wtrKen6IB3aTDKeJvnwrph+uHt4DzeZogqxZoUhSviM6wdLPf9oX8ulYHtLQADp+S/anscDHyIhz
u0gSiNplYhM/5f70M0BKsX0PkNLODPvcMBQZSRTUcX8t6v/h+Tf8Ahh8t74qqW11V1fpWvVZ97zw
7ohPaI5NiVAAEVIQ63QQpubIuBWJsyxPaDWbkM1zuX4R0nknK5LMDCsqDqCrK49b+WkRz4MFi2Ur
VenCdJcQdhi2EbqYp709cf+kjvYrEGnLsomLbSsmjSo70Q4DNhYZD42c+fKvZezhRuNiCxTncexG
DFM+yL2qpa2Rdtl63M1DeuqiVZzARvTthZigpYbTL6rnkFSG4cUGQreJGsS31Cen5Ei1jkbDtEw4
ZCNuh++N2Gpy+NP0X4mSX8UAVdttRVL9wWXYe/O5vEPDZDTR8zXYiHpPgEqSukB43FdURmMcM2JV
1ok+7BGlKALPgxFvYwglZz5nFufIco3knbNMjxb4i+Lv0Nd2HqGKfCtoTVhktADkn/ByS9bxl8p6
FYdOQAfnapaVm11Qyuq8pXzepw+t9rMGh9qQ9sNGkNU1TaiH4OjdrsBmnwEzHpJHz0Qog2oB63Rx
TRPt17MUZ5/g7yClW7+1/u0g4Aq81oA9vRlvYcqCn8IcumEv7S5gOiesOrkgdYA8YwLGCmsbOVwW
1PwXstytiCXrSD1ugt2VfFIFFRSyrOfDg4kJFsh00A8E+eIIM8ffCovKny6ppGDAqsrcdARO/xGJ
Ydi8xzpwsoduyqH41rd3g55njtYS4+XN3VJPINcze5c8kY443cC6xV825l8lZfL6rgfJQLEsw6co
2CiNm5W1/Pel5SkQHD5CPanosRjCvMps4SPae7iMtqps6LGzGEu2XB5br7kJzI6187qSdXz5/J27
BpYLDUSjnaTjEavBzopMKtTHGJf4LY1XpMQhND7wMpLQgpDJP1WBqATAX1nkAaYiw2Q7tdKpIc6Q
SE326wbyEm/rG4QSo6YIPWDAtcDkMW8+MlGokyJOAJuZYYFxTCsfmrZgECTuGeZof98ZHBnNccnh
1D1ONH8L/0A7c4WLo8g5AfuBYnkhlGFwzwOpThKlpGh0/VqdoV5iNXUbea40sGcHyI5EHRB0IyFM
lnW1XI1qTr+khGNJfWnOjTJzLlF6Qz6kFt7l3xUYTEpAqVgv3/fqvd220LcNbQBod+4DZeWqkAC4
1su6aqRt++x81zWPd/wB/cILcUDzTTPfQqaR49H51fp7vNtZK+Rl5b2oT8BKmEFUfZPJsNmSFMZG
PUNOZYAx4MuNxrNo+XhrKfNox+HEF2NWelZ8HBaJmt99cHDv2G3z6DDh7BCoH4v0IVN7RMGXbyZc
g7uzbxAJ5WOc+1ltzDItFLBlkqtP0EAOEMYDrkncE+VTvaR943AKKCmUmOklW0GyeG+8U6JR1EwS
cf+6zj1xL24o8bY3QrFtLCoIX8q9F549qx+3cfZ3BFK/B9bxtln48p0yHMFB+pjwkW09YgJMn28P
guEMRWDVqmBJ2XBTWF7nUG3U/f/Ne0ys70UYmKfgRRp90RO6JLQrP6XpYNOeJWujh+QVjKwIV3YD
b+r3uU9fxNGYmAGBE9GDKcJhRn6qf4r7KLr3kyiTIM4UaG1/Nnsz7MoudDpvbeUj/KLF4r7SELXV
7wIlvVtyN/ACNYes3paScrhkEon40PN37QpeNl4xmIUuUr0nnhtkaEtcVMJMWCNlkw4pLDfx/yV0
fdal++4JynI91kCWnli5Acib5fu38oAN8vWdHwAlKLEdM5a1U40cB4sLnzuLtP30v9horeRZzs57
5MNFoeWfC6oQgYYm/4yMLS2TPcO8qzrWblGMmuhUKxp3TOgdn8+PAyx3Cjk0C3cDVVJcQP67cBq5
xGlVJKSsVWMj5WdYl5Cbp2gL3JF+n4W0uh0OwEK7KfRZ8DZlvCXo4cAu7mMN8TsuVogCexBA3SpB
haY/R9fcf7ov6WiWhl81q93mYBAuB/e7ABdneroSse93TGdwEgBp1u7lPA7U9/TBZfNCWFa3/M6x
+6WV4oO+Ujtn/JW07krUfcsnJkZ8mq1a7v3MgYKJMrqwAHNSaDBQWeOJgKPsT8gzPO2jbkmG//AD
FycgytjsdWzMKl/z0v4dkSCA2Fuy0wCVJo7x0vxucqdADKfIqHxZH38YymS8inXp1DPmQzZK2/Ag
suOsvcswQmK6mDD5uoNpot5Y1xULxSTWEqFx5ABMzGcIJYJ7mQiN/834T1FikJMwKvmmU1MNwK8a
9nw4oXL4lViMHEtiLLlBc7YDeFdBm9RxNtOVJw6w/A+YmmzZ8M9lqjSsgrxhjbb0z+oSTfhEF33o
TEkHoNSGu1UDlPIrDbNtVAXx4H25VJKoNUqjkItW7P2AprA5/5M9eBgf2TVxtnKneooKXUInWR7T
ZGHiewOJbfTIjcOc4qMMYaUlh/0QM3jxS8SVruLldUahwIW4iuXp6eHVZ1hgIWz6DqKkrA0JkHPl
LE+eqJ3v6WYdIz5+zUNgd1oby+gjSRCRNMxuWKHb8TpXZXeHts38QP0aSdtv8ET/2rjOvfdTOHfD
WSlk3pxPKj7wOgboJ3jTLBbUzQRBGTlq0iSLZXr2q2Kuupf49nD87EOJUtfno7O54IaDLbbk9ObG
SUM2PTk9S8/0J9/zIHix4q4WKWT6VoZmq2U61sfwHAH8eFiIhrUtSu3dX02EwRR9RIcaDiVlLOCr
w/t9X9HyPTjkaTF/jhn2DhUEiizzJy2AmKP7mel5lGOwQWm9E9Z4G/76BvbC6Aaq/7dImAQvsCzc
J3kZl5fyrc0JdeEt6mhwCSlJOpRFqP/BDj32ahcupN6Iq5ne+eQXLY2kRYiOQNibHO2uNM0WIAFS
+tknYDlL4dMbX+nWyqENd/fk1m5cXlkudy/S8zMwvF5OvYDO3eGA40lu4coUxAIkI801hpN9Ez1x
yPSXr0pYuRz040kGgnf9OXnwmeE2nBA43Kc2WIaIU72S257h0JFx3IHly6KH1fGG1/XZ0S82M/IR
EBQlV3ZRYvMawK2sqIjRjuWMpy9uXgoq+mEuXGDm3qxs/f2xjotN77DIm0LaqNnSJOoNTUa45q/0
l3YpZtPlZgv5OQKWm6N8lgwFxNs2aeuH7it+uOh66UyOxuwVJsUUxRru4xq2LhMosXxKEc9+QMJ0
A6P9McjR/KroooJBPD4f+IYui4YmQKEInW8I2Pd84wtbnY5i5IqFZuPeZD9qCejJQEAqr19X6DgR
Z/MbMPDwxE23f4KJtOrzeFHbboNAXQdH8dG/J8nJkjlRWa5F80xVu1D7NlHaPlCAkcFFj367m282
2YQ3aRsm8gJ7h8pZ0MR9Ua2mL9FWpy5gQsK0YlLAzJbMgUQsDnKGEHMqIKmCq85Nmc2G7LzrvMIN
9vmCOwP9njMBRlpWBblar4REWQO0alsQ/jfgJ8LDHWHuzVLZXFPJNMhtlch25jXQFGpZgkg7O6Dr
ehxuJ0Kjrp0Ku5oKVHSy2b2uaFWaEw6zQyFC3pmMvpFF/d64/UysDXgPy0/HYzOFnK056BnwH8iC
AIjiwWgQmxOPmlxU7Xq8biEaRPMOIgWDNJm/SncDGYqazvMNPIhnExVhxq0DXA3Qy3mwvm4odePE
lF3/HTQ5pKpUpVuKxTeeay15digkfeiLR1Njt0ze5uAMrDcvd4AJ7t5FEITokzd5FuqSRhmWNyFN
o32xImgCqeB6gpqspS0EawbTZXf9qnQBmxXzF1mgbH/jayF+57d7sWIGcBojojMNwrcQhF1ci9fJ
2XEmUXDkIc5/HHNCFNwDXUqSzoRf7yJPCzWdiHs0XIRvuotPTMT3ibTumvu7UUPOk2Ivr658Mcj/
NQIiY/27rKgijImpXwe2RGaxvmTkoHY8dphh1EGgIRyDEocaUiPZ87rrKjkpsu/wL7zH7tI8YXd2
sSCafgfj7TShbiYdJ+JAghRA777aVMRusH53ZpWLfxguMlJFSRRCWkLb1LVaLgEJ26jbBWu+h4Rr
O/cyCxCGsDiqkHdJf6thn4/GDwPVneDcb61lbzxqE4qwglHNbBtFw452EBp0fYwj4p2kR6n2ktjZ
L4BP7S8o6chktOGN1VTmWde+nQy+Otke/Fu/t6WB3MnDggsIty6WzOp0UdVvnsFu3wVNlIf//BM7
JlUUpf/hARwXCVQv+ydJlA8F9YyYIMhiP1wl0c+NQ3jhn/nh1N/93kPZAeKC94101hVr/1TfAFLd
WyTO2y6qcbaW85VgW6jcqP+uNVrfb499fcLPzQzEOoUm+yWTCrJlzUIZKndKUQU2mIVUzTT26TVb
2WP/+E3bMtn6mqyMU4Ii1YrOQPzoQ/nDcAmtIB/agVdv9qyMLeWy1N5cJhWP/mqxcyDNEohnlUFY
pL72vLzyfjMAiRl2iWEaMc7pZD3+vFKcyKmwU3C/+m+uOnKuTewbpaxAKjTqCM8rdXHDPmx0q/Au
RReSxHJhyY1jv3f93p676ek3nABPwEelofbTWkpXcR7mzhq5+C4JnlHdu+jbCgveasflmwNXU96+
euan/B6ol70TOF3OMdwr7qy/2BVvkcREVJEJjMYA9LyGYCd5QJ/68HA30WUTlt/kZ6LbiWhzZ7sb
tWRGt5BjBi6DGhnU+Dzw29ZPR6wfjyRIbCX9T2EqKcvoArE3zEj16z0yZA9ZqPRc8RbiWji/m+an
O7C3GF3FKmGhhzpkkJ/hc+toJKG5kZ+jWaKPgRx42zuXs3TR6zzA/GohzQ5sQ5IBNheHllntx0lu
aY1fiJd62pQnI752AwvUuwrqhjOWncrckjcs4lSPf1le+yA+aX39droB70zC0B/FqJlhhHyKD8Hx
dmUKxH3qeOt7SmtkMeZ6i7Oi2UET8XQ9rCKiOrhWGkSw0ao9Mf+NwjwRzg9Fioa38/+R9NUvAKXI
JvDUL9ob5GkekoV/4TfpA+nIXr1CEFn111Em37Esc5EQLx0iy+yVDqvbPu3RTzpCNNoXYlkFixu4
ntSPWTfNRU2l7fHvGKfIcT72Lbr/OQgnVMkiMIVgxYZ5YWGdJq+UyKkGeDA0CFRYs+ZoIhSOzT/7
rO/LYYdGynA1RKoYMKwDNYr3Jv0SM4MK1OEcbfKQIAn3/6r/aU5qdjLniOTFHrEjzmTLm/nWfs5R
pG+vhKqNodLUuFfojMh5LXj/+7L/ZunX+YBqjK72ZhVtJHqOu/pPE4KqbcmhH6rpPF3oi2EcNTJ5
Fz2I9R8tQCLlm9T17SYcRBSY+T8uhHT4qsWTPfJ8v10wJDWrommi5ZDQzF+ZCbbBrfLVDbxapcB/
LbuIKwxwx+a7k9WzKvfAmSU/+CTDfbx3A46QQexfedddkvJqk3dFHF6K3it21PNOe2y97gjFt0zQ
Fiaw7dP0dpCaOxKEk/EudB7NCFLvJdXhDGq8hdFqkR/UZuHoME2z7whs+NQJSH6+POYu3H3SvXCh
yYIrlXt1C7EtCjPodHtrz8PmdEvuiNM+4HzoOkYLK72n5vyJYoUxo6Jwj2OUx7xV5Kv6UIvAzEux
CyAhnwRZPIv+ByNbxBVD58FDCn8LXXLe9QuscYf7pLVFI0gP0FJNIJRP6z5xNIR+3bsVYyaw5dTR
+0N/QB2NrhKd7Aq4h62N6I0K6I8pt2DOixXkyWVKkS85+BpM1d3PDZsFtcZeM/dLUpge3IVq7lI2
o8EMoNeE+hofdBttDrFyBqFcwLg/OvsitRAugihAdIOg8zPx8Ay4SpW0BL2Qnsu+EYWH6jDOch6u
Tjr8Ee0AgDrumBh66qqLVR9lWVgStX8F/wiXw3mChwYAm2J7wIL9/TigyguNRoARSFWgI35txdfc
E0sZc4BLu87o4YKfHHzBTV/Ecc+AGczfwoTseUHVjhqwHo4BLjfxRvIIwIx1q/7+mVyq101eNJLG
5lz8bZUxJa9M5Sn3KgsiVXMnbF8BWZsjcLxbSCGkgTSBKXWhTpNGBc6bLUXMxKveWImS09VNxvz+
bIJvYUXhjc5WpN0Vik69kten1r27W+AONqvsPzB6HJyzDORFawobLooFDAIqMAiX4OefqTVpRdA2
ZHcVP1tLHsqatxp8FSP6VOrnVPu3q3o5uZSeAEhyZMJtZrO0fwqYvp/lsnhdNieMaXamp2z2DVlj
J1R/eFykuQFZnrIvYH1L2uMogW7IZe5p2+4ULHXA4opgZv78hRa3b8Q6u1qlXb7VfIKYTNt77uON
k10tINTF0DhxHZH1QkmXlebUQKMqV/vSncKgraAC/M7cDOOHbCTWpIDg3cUn/UtwvqyIffqNXiva
2/nbIyI/Q8dr14vi/FyqklsWeDv+dYWGTP1JQvgT8NZB8Tdk4T9ngd4FL0fkouxGGawP6FfR2S67
h+YVJcYmotewQXnQtuix36X9x9WJ9PXBjAE+x9HIm7f+RkTZMYlviivcUYPVoxW0i3sQ0vK3CHZ3
AZ1k9eZZs+kbTZmSFtqxcxYSMgIc/T7209OGDesaYH9sZB8SQFtOyOhKlBbWwgjeA4VP1aRfBQwU
Fsih7Ys/1wzbMBFaQOo1Rw3IOLThDfLMKJmVw0W6UsFba7h5MsXFo9lCzUK3eBGd4D/4OCIZ77GL
Xr/rGkyIKtyIERKMXZuQdiBJciguF9OVaUGfsJlwlkxHhHsvRNV9+k2iz95H72rPEWJDXC42zhxM
Y3R+pihMegKBWBMrps3K/2j+cdHMoay4uJASD2Rlmw0UzjnHpMVwrQn4WgfAjJ2xnxS8OczrLAee
PWNOpX5ZrxEFRN8KTocgueM4495s5CKjPhhAtdmsbzhxt+HeBkgaDpnlmhgMh3JfdGmLPIxIWRtI
izUmcYj/YrVFapKtuupr5Uyr93XWgczA2ZTCsly3/00vH9hLwPyPncX69gziK6urAxnuye85IwfU
ywbNaSDOkUlEVIoUwegk/wmy6poaGxG/vNgYFHDxQnzjuWBm49v3ToOkUnrXGVehph5DC9yQhjQL
rT9ZtuMwHiOS5fjWeoe8xKkHOOh40byJWDG9BAsXnG1lJkioYDYQgeE/D35Xm06GsW1qEhnnHXSn
vbTML5nFExY5ccDX9eq13enbMobD/Q4u0zRq0+zU1MpAjVhbA68jyiKyui3rKLsV985jD7Z5+ZK8
Uu+6GXaVyV51vKsK+pVck9g0FOdgKr9PHUV6YckuEK3g9TKFVCVEz/mgoGHzazIEQgNnQZsRrJH4
XNxR4uUS6ObIz3JS+HJyNvFZB6GPltfxdLad9uZqJ0OD+zW7Yf0E0TjIijxo09JGqykPuBFWqxo+
kbjrdq02R9Wyc44Z9lkLP4j73tepXNORTXZ5IzoTkNFjY1tD6wau2nndZe4+H1mO3aIcJL/UjmIZ
JFWEYvIEnYS5iODhFd8ksgmGQiavRPTexcKJgxpXTRcPzVWo/Mi6drst2MOAUIVMvClirjyrPmHL
eSFnPEoBsJ7hzzXTpsC9Wr0lZLDJCORtMVhfrKWMYDDtdXJ81xVGWPjKxsCdczR1/9+tzkplmqGh
iELhhGm8ZVa/OjvC2wXVYiiIRpqMoZ6MbX8q8yKmF9azlHmlg8C9kB/JWO6ZKmKLCeETSqsOP9Tq
jW7LeZABmig1n4VlIUYuO/1QSRybujr5PDTFlGgir7tlytXvYw90lHhCKkmRtyLK0dbPqeaIYs/o
cXmun89j95rVJVRH13jeKgRvmXnwRePJem1uK1X/zMZSDHAfwye4VlWhZ2xD3QjmoAFtXcMw4l4I
VoEKDuI+sHHUD09JoR2uINNoOEDVRmGoXTkc8umQ/Lm9l1kcvCFhntFrPj/PlCp+Vj/CzODU02IE
cvr0AWXb33rBO7WYsdGzb4QbEhX01MBju193TzUOMyCBHUVLKERurQSS45Q2ZxnTRTGfEZXsw/lc
DTEo+sygg6LWi7IaTTHuVfa0xSc7ChKBOAOV/Es3CDvEKx5QNk4MUHkJ6W09HBulMl6jSw8t7k+h
Rmr9hzTxZoSVkr6O1H1hzn85oKsGhHzk5b9bZviqiTBgt7zkrcKxv6S5kZUxknM0ebqAEeD31aCZ
tYsanB2xj7TdLQRu+XhQiWYZ6pROtXBkU+Yh/o88X6kAc2TwDZ4BMTPuVhVcZR1YIsMPr7H5BFeS
lbnjEwgluF3q4p7swOotHEHPbKfF7psRCfZn0W/NhChNZJLgEliwbg3NsObsDzKcvMLiPyAqC29p
ZR+DHAHWYkz3NEIl5xVG07u8KK4GmcDbTxWoQjJtuBog4ZIBDQyiR9nNAzszkcjts9bwM+GJRvrH
WefoV4ywMiXu16ZqFj5+GtqV3e5kqdEZUPJyVo8LywVewbpk3RpbHiCGU4Zj8wFB0Q3utGVGTtxd
5ekxZG6FlJfeGjEPYBDwdKyhuVJyM4ngMDM8Xlgycs7j4e9td64Ba4R2XWnQjV6FwoK3qAQW2G31
zYrD0TAKX5sx+YFT6MedBvy3sbID/uri/mpeOPdnOO/HjkFKPLvamyYwP4uTxMXTkPTO4dKQaUg6
shjUtgcIZC8IT7R7BqXoi7cTlx9MENIW5W4ZYHAA9tHI5mK5bq6OZNFu2UUvqm8t8fZwPzijlTgL
lJxrAtybNNlturVMHL3ANx1DFp0X4/Cht27IjF6SNK486Cy/YQlozz4zvULFMFJIBlnd8kZxdZj6
VOl0k38HnXStT7swFmubh21vmefhP+yi1fnmyJoWco+gcxkgy015u1dxFjcVo3UGqXXmNJYxQA7T
1UTfNM24vVUNo4UfOJdv+aEA7XE/fAJjFwPYP15mRANU33f6/j8+kVLbo32QoKKA9PQmtD+Gw074
VHD/R81C6MrQ2TiVPaxmVWI/QFsdvMSradBIuXYFObJS7foohfaTaryLWOQ1nfogFowkkIn3uCq9
pBnL/ldKHd2+5VdlPoDnWgqH8KMwWwglRLGl8ka7i5ULoocWKWHbH7tMDJm1IYkF6iqCGHlnI4nr
WGfvq6a2iJX0VJtbEcIWiF3+wtxl2u0a6XQbC7ZLIS3JbqlEhfCqBjuqSMASezLTFn0IvALUpx5G
oymVbRQ8tn9YlJaHiY7yfp8iYhU1gLGV0BgQKnC7zIKtUIgpuO0M/Iz8EqMrOzEc22Sy8UHdcNvc
kGFttV12XI85RvRT9cSdgym+6FEutba/BnF94pVptNuxQbKlQJQJe8CCMVILD9AsgcuXLXTb6umZ
vb/WaJXGnyOm7oPVtgv8EaZQL6NCKvHo/fkP4LWgseXzZqa5vxdljwmJPpFD2kIYOJapUPyoMOB3
B7b+X2sMvVRpUB+6kG4IYZChDg3qLSGHA5IHQE8hky57cZ17/bCoFqPAThNSolaO/eQ0NuwMSk3u
CMvEoHdb9McdM++Il4nK7mNATFGZqVRjZgncBrIqSC2iBntNPLK6Crg/Yn7SmGUSD3haUCorTK3D
Cd7oYbh4XO7Hkrnuj1HiPp3BMucrGUmPBNKL4dZ2d6bOkS/uOoz8e1u0castJ7ATjWJ2sX3J4Yv3
O/4t/eDOrfriA3dkcEOJynKDQeDhLBPy5VjQRbR6u5UXRipqcfYMQEShWxu+hybcnbLvaqSFseIz
wVY9+1VNePwDpY2d1nClA3axR+9rLbJxth5w480UDHZUm+O8DGynqNFKmVRpAru3iS7lytxFJ7MG
1UX/HKnM7+7SgMjh4RJZ66FtVZYXSZ5c3PH6OeE4/7hp/P3lbG9jQgCvPinsPsk1YSB1kLRWZRu9
M+BknA6brim4X5m5gDKusC+nv8xKdL2Snw2eHfiNn5PfJeLdex5gYkN+SjFRAeVPcVWpM967T0XU
QZFS2hkNN4iH30oAP9LQaV+/V3eB6MebIreyF+t1Nn3BMlTlasyZOfIVCRweXIHCLJUuDbD1TVEI
Deolb02acSg2s4oCo2reu72PtvHqMbeJ8h5xySg7RjgRVkH3MvSAoxX3wkXcICp6rECusSs16eTx
TpVq6vkydi50+h1wKhIYBE3DQlIdA/2HFyhVBmZ/LYVKcDFxPK/If4TRil+pg8pPhszvogQDMEQ2
lBJUj09wcTvnkMLdNel2Nc5IC7WXNt5bzm7PansV5JbC5cZR2AJBBv/O48dRh0N2N2UNoX2ytOUd
tiaVOk1izVeSAuRGFU/wrQuA66ySsGJb5KyDeOGmgzJmcU7R3qpGTnIkz7Bljwf9ePl10fhU3Yic
v2+SXoKZWINHCgd6eMJunSjqNfmGwVsSNqcQGT7RVqO/W6j1QrxFUvgFkSQWsiJbO55SsZ0m+VX5
xa5BS3FftUfvS0qCwnLHkovxRf5ofiyMBfWTfgQyhmfUc7D8u+7ont4HZmsXV4rf6one5+UOiCcI
YuuawL5hFqJh8+8Gmh1AeSv8kMjHs8EsBrnipTZr1Lp86dbf++S5pr278E0EALOhL1JYqc+5Ij9b
V1gGIs2jUr8d/epmsBlazTiCBHp5Yt1sqPwBdnDX/YpbPcAjsGDhSctHHlNRCUF5bRyrz9yHyeYi
b9IUJNnzygjV6/rQRlYqs8fyqQoAWFtEAuksm+faUNReVBnstRxBv72q8Ad7lE6ehVhxR9eJt5Rv
TiXhMn+zANKThoGWCEbzEHmRaUY4IzscgzAuS0R2cFcSS7DPciwjs/B/QI5IS8KX3xZQJz1vca4k
siATrQSz0Qj/gJdue6drbZH4H2HnqonWIq5YjwBnBVf4xISSiRca44xPhRu/lmvNiNpqWn49PpRT
PSWoP2d0t7bTQN8rqxwzuMQlm9DBGc9RW3u8C7yeEOow/U6N+9J7lYYp4B2nslm0kzGFaLTc9yEt
tfCyDacJm3F6aEedDuPjQ81csz+0zYiEA562yYFcLr11ROwKBo+pKIdWLYi3RdMHOOB7QGUIDItT
/7tDdAmc+iD8U7f9YC7BrMpH5fi+YmuSotyBXofv8GySkrRA6TOUeiXLciSAc5jytiHJniVVaG3W
PyqYDyAbZ/8VE5k3WJlmXyYU05Dmb/Tc/RBrqfbfygfQiU6EmaiYtqP0kVWvNNS3cGXP/U6vO+IZ
/tN6qnTISOmXaDjTPqNusznX8VFdohfDr0osm+30x5imcZnqpaKQJitLLshFsfBsFGcVjBnSI3Bx
u5ZjfN4Xufn6UgGE0kEu0N7JZbFWF/CMYVxgTZz14k0u2yXku1w8Ja1sh8FzSjT/HmfXc4Ng4BnE
W7MxaMdTiFW+5VlwjGBbTLZaH5nGmxlSqE8buHgXhQ5mnLLYn4PoGfl+8X/3KZRHI+fe+LOjKhFK
UUuEfGI5HlMVZe7tEB6Is8VQciYbFT59dJUGlCiUSN4QvnIHTmURJ69kMx3xDqf2bCHtsIIUAXd3
+mfMoeGZU1ZqXP46B1GggKzSdQLLkYI/bRLRPpSI+uyrdR4k5rX4Yl7Aaneux3NmBilMqU97wZb7
bXf/F98X/HcF7JPQnHOU26pB9qJk4wlkZzScSKPCQB1K2ejRHdcoerdcNpWg101W994z4tgHLiKF
SkWz+CJpjb+s3BO8V9bMyI17NCvGWqwd1OTucX45DA9KPzARGT5RYTzwKyQ6ZYOviCJBSSFhsSoy
SEenTGxoVhrRGaYkiazrGqEwr1afBI4XChAK46/VkiazbBEFoqMXXpZNqsWFszKrYFgNwhn8KgNM
x0uXVdMYQfu+2hBJrgncbG4wPaUmEKIBOIxTO7fN5nhT9RST5+HrJIMWYSIxCG8LFFtyjjQuHieC
QVslCu0AJOEXGJijPXTCKpWHMbZkJL3ECfGAEXthkCRNoR3xoFPCRTmPE1s9bZq6UnDUK8i0sJNr
m3I3BC3CUKPAhVE9Q6l9fOTDuuoOtNY5E0R8EVDlyPVjCUju08cSlhM4IJ5GVHi/zKtchg11bHvT
+NsVjPbwmcYr2Nj2mKilLmfvYgzjEzz6NlMYHTXhRIZWrCG3fiTf9ZX0lVH2XSA0p+e6QSIcBaOu
Ez5RC+mnIUR9Spnz1+zVVSbYHVYYclVWXF7J1ZNA2m1Yw3gcug8WsMmn+xxv8j6K37eaH9wZc5JZ
jYQq+xyJXFAtVOIl8u6D5td7mwXohTBUcbB2NA5J+QygHcd8Zuj8CgXXm78NZc01bfqhLrDCtGTC
t0ibGaLOzA5VmQYfkC+fE6SXocS2vilfOJQhOF1fQGSXR0ZpVIGumuzqbtBzLgNs9ewzdB7d8lFl
t/Bq05Y04rqkzhXm/Gg9bRJ42WqD6+QdRq4u/ONhTSL8X/RhdxRplCiJF/qerzU3y4f94TmV7pNT
sQmS8wZD5mXp6DUpVaWgEQxx5HGVQLsEPhp/fI1kMZGHllOtvI3QXG8W32oHNcFLlBiZUkyN3dZd
MI7xAf4cfXAk5cgOgV4pDNQKyPjfReMk4Q5CNsqE1p8oHqZKImwK5q91eEbDqdK0BftPbl0I7CgB
xp5HkWpxqgis47u9Tt3ORNzBbX7dBT2UnZIZ1oweuVbiPHpd0S1CQ8xuOWNGsPUMyMG7NqB893pM
3pI4PJ+PGrR7y948lfIcoC5evmhNGVH4+3GMm65LgjvTHQ/Be6X9XLcM8yVYCIYc8FxaIBPCYlLn
ikCvUuS+ZBj+cmSCl0isBCDL62hPCsf1oHsUNRY6M65ZuRQ04Ts6vdffqjuIbXDHo59ZbBN/tk97
HFalHqHj5KAj5Dy0s1TrK4TLvQpqNvy4o7lgrmoJaxxXEVm+j0PG5yRNovBoy3CjkH+6DYWGEvm6
OfLj6sBGVW9NiYtOZTkbc3k5UM/kZWBbNlYOb5zb+SkVEpMqPuXA0qfVsBeeCy/lmMqAbhXS8Z8I
ifGXxG4ZkFT0J0N4OZV/J7fc6AlW9EtFJZv80kcBoQWKNffQtDxK8O4Pvgg54fe87Bn9IJlko0dc
DXErrkkhTQ5+9QKm3DYP3ZrINOiHnxGAMsS55FCZEqepKdZ5rGKQH6ZBhLAnZJcAChRmmQCgjc3d
Is0PYxvJeR/nbAYuPBx7i+Bf5VKKfFGKHN8FCkppn4+LggB7fUpMTMrh59j5HAyOdswNeyO493BY
3Kpo/zLRanfR2OZ3GzQYn8v/6ne2HuEnuG36t6Krqewy+xpoTVMLxBjTWA4j7eSc3bVjyd/QtYlz
tW8hXbsWna1Wn6c+uKYz3yRTl9ukwMDRbf7FjIwZwBGqL1Xh8zct/7q6V0V6FAjLFWWD1AC54kNl
Sq3fsgfPcqtN2aL8zThkkg4k0TybvQ6QY9yE2ps/9C8xp3o8mNRuIgolGCx9EBfu8JgWdqUoYoPH
QfTJyFW8pe4sNj7ZNi+2EPNWBF8SoNfgn8Wxakd1CMfs4ZQYR+hLDYJQEaUAQWbHaRflliLv3bjp
NVXbJ646KRWBbRxz7a1ff9+bPcfOo1V9em/Vz1Sdm+1OSC/7fykO3j39kqX/b/uP7wNZ8rp3iqHd
KW0PckcjikN4sH7JPA2v4DgSasWDR6RiHalCHP1uCtHVicAt77RqWpef+Glskx/4j4qn59aTXRT1
jD0SWrb772G3GEJU1KPqqI1FIUm4fH0pbz83PCTaabo9ijfymI4nznftvLKbN4YXgvVtBydIQNZa
D+snh+9Z8zjZp18ypIDBXdNpdEEvVIdN+venKtJTXENztVcemAhBNLYXaxJGuloqBFJ1C+ttj6tr
yQXOY73ychVp4UCf7XgWxZrlXQl8zFmnd/2MCYuA+pv4Bqx1Ix6eBw/VB5WKhS7UgG4wK/cEcd3G
8nJ2pVAPRLeVvvAc4CNtOWncMKn4VPcx6KqcIvoWfOj+14A0gtqeCjD5t/S8iBo8kH90gPKalV86
zmSMdfbobQuUY4dGGCQ1PHcU41wc/18yn8t982h3GwubI1uM0Vz0AEjEvJFT2UuWlbb5aUb7oxFb
gP99MeSa5ABTtICsHYh9Ey8lRgzL5ujcSuUyMVIxKaiv0m4c/JxmNIoXsHtGP7QtOfo1Zu1IY3eq
QUW7YkI7bFQSytQIrctlIGCEUBK7yUsP1XpHwd0ZyJB57LJfdWq7Oiy0rPAdX2UXXo1dsP3c+EX0
AnNJ9UURnWkGz/wflLv4a6q71WuvpVSsqe4AgAPKny5UwwHqf8IVFN2m5ZTVIKw8Y11kmMilYDPS
DBi/vlC7frj3eJSDYNs3JPUT/A+S6399fzjBWd1XBXgofXrAgmoriIz1oYSFWwQO/dBVz/AfE/nQ
fHaBTbyu/q6ZLxy+L8cj0CkpgU8PUeDoVlOtp5lmrrYVeSzh+giiKRGJpsiZp/PrGc50B75crVIw
/iLK+vYNg4aKpE+9eMKwYdwMdZ4SmIoyNvKXXXlimKgKuUNGjpDSAy2QS58o15vUyOe9/EBvLG4y
miGJLge4LwIW6FeZ+uSq574d2GuwiVaLomF+yaus+gVkvA5VJKEHiWtDM9coNzTou49bMmtwHUIX
tHdtNklF+ATTw9U+Xyw2wr6IjsbdKopw3gtA3zEWu6hDsFQBxkMrkTJ9s/da5S4SztT1r3K8Usd/
aFpobntJ3mNfA2CPoc90lTsDRMpNlMEC+rp/jlrCIRe+v1KZldKsvVsAzIwetpkBc/kZ70IcY1ic
n4Qu0JK2eQM9rhmBXNkw/ZvPsHh4PbAkk1PW3dAj2gp+R8iTDhvnjeTd8aae36ZfuH7y5/SgP16s
CVo679YhQK09AfwJlCD1V+oaGt8LNf39JoJIexN6wNBZAXs4f2T/wRLueBNusmV9FBBVyXz6pWz2
bJvHEH/1MNUlBLuW6JXYMmuaQLGId0jv1rzeI+pdfGKTVtFGgiuceTs7ULcDPhm6S/YgmS8Ke5iV
fKHXq2RfObsxxW81Eq/cwoezrvH990fVWiE9VHkrYjv3qEUQabT0v+WbY0RznHe/5jP8U893Ami+
rzSJ0aoWxREdopiPPuYvRaCuzr6iWE1VQv2KfWvhJ8ZrlHE/Zxgkn50tMhmmrZqalM1oGeC+vH+s
I+g9ndzTdTyyyQDfJ5khAp1mrXbjdgtk4kknuQ0oj7GfK5f/BwlnCNbPRiyHqpbQP88o1ZGT2qIl
yijjtf690oIdpHYz3cWCMPzfUAb8RnThitTaBT+WmyOg4kCMchctVKneMUCtwhjkDtEQiXB5pQcT
16eA9evMC3tQZEyv6juvOiKvNEWiDUif5DKEkbhFvFpY7bEWZSspL2KXg7Aj9K7GJ6R/lq4H9RDf
X265dcwphZ8dYkTi8DwbIq7Rhnw0yviNGOU0OWMECzWtKm4BZ2lHzDCMRZPNXt2leAViufYY//Dq
GHdK9ZMm5fqAEVWWT4f958Bq04LeTjuu8W3BCXwe7StUPvLShq+F4L/lFm7WL5iCIRXAH7xmlfam
AR2bZ0NY3xN2d/F+yqmGPnk3Un19Vc79bLE9qhw33lqvsXZK0cDjBWdrcvqyay67qiMHQX4uZYG7
3A5wn3DWPnL//xxl+o5xwiYkX51jxiYC81D7Cl3XMH0Hj+dWeX21EIROsR4NO3jMrLi4UsVS0T4M
KLhgIfK7X1ZZgp5NstMUajE7xl6dsC9OtGSzwTw0BpIaI3jJKNbeRNd3VCUADxO7WRboJi9PSSFp
VkCE6raTbf4DzctepAT3PpOtrHlhrNoAp6Q5tRwENeTgwCuGEjJoHLAhL4UHpRcR+JAjz0nPcGxA
KUsnQCCDEyJhRr1aiPhAfkhOSjxHr/bCC2WEMjMCZodCMe75MLl3SWWRb3hS5nQ73GX+UWbh37UT
d+hoAck65Jcp6y8ebUgorssfi+AXHX15qB5SpKooSC9RGs0c7BIfmSQ/HY+ouVjhuW/81mxfOSj2
T0COcDFclPaSuKIEmTBBrTfCG8iDqylftrrIsUTojpM2al/DkqqdIKS4/r6ir2BxngSWuTVs8ZRO
3uGDoX2yhQBMrt0qTFswx33+wZB894Z2BCGuke3pOkL3wLGsEE+61X2Dc7IQ6namgzsWwrKZvE2c
R2BFkts/CeTrYhSdWGGHMkSEothWN7OPrvF/lkRF/4dZetwDeCXCpRwDLpUzXsp+0daWWvYamuV7
lRd+4PH8b5z3IIbIXstYtwVjXelos4XimUsQE2P7XnKb4mcGDrtN7TEcYUV2lT4RShs58wh7sqtU
c54cMkopMRpgjBbFNGL1a0AaaWntWz3ZRKm2CKI7BsmQE8XxfVAMgopo4wiLdkRadjQ1YT4NykM9
RdIfEgpva7YEhzwDZQtBIDFuHgbJPQ1ee66K36lhXUW3+ZAKBCs3l2j294BjQkx5I3AiiXnxzDbv
lXQd5L6GDTP14VtyXlDirhIq7GQkMkxyS8UH3CpAJVxIvErAm+h6sS1qCW2KMZPGgRKHiS76f3G/
UIs5e+UqxsIkQbGznEfwWrWjzjoQqPwze5QkMncENGM2zbyxXBE+FLuSFK7j2WCWlkhNob6qAkL/
Na1GBYCcEYV70XMoHh0L29urHxiXPI7gredr7d+xtcA47yOvc/Y9t/fYUTsw/rZHsa6KRKjAr14c
ETqKQKZKIaglA/TW+5XJrH9TsdzRT1eyCM/YgDUsEK2lb7nXkwptiZDwqpe8KhKmjOOmexR5js+L
cvDnZRCnZW0CLlEcrtX4Kozs/AHOKC0eJLDGOYtvvg1zJl/ZfocNSXgm3c2D2wUAdZnHSrKGvQui
m81+rsOX1cVjv8K94TeNM3+49Xmc8m9KgbOfZAzROrl5BYfugsMurheYujLmhCxrdIsuOWAtfG0T
mzsQocwdTe8es6UsPfzxnEmwBjcoz5CMAsOPyFzEyRmL1aJHJ7mFThE/8QnlmETK1jGVg+pRJC9F
K9FudnfH5Xr5bkiaOBqYq8JDfYtK3dmFwmtwncBeyFT7o4ldZ0a7+Q7Uj7kGVgfqxc82NVIQ+2Ln
rVxqLxFWuL889iHleOYJ6ZBGTJs2Fg08VAiCKHNfnXgwtdasyuw/ohZmSdloAvYPE/UaCoFphYFp
fPZ5lMxsSK4ygu/Le7QNZeBUjZ5fGdKyrWdSeFMGwmME07kC6rBSGh6YMsnBK+LKNEPcA22H0fFZ
503ThdUi80Imy4BkMPPECMeX+yAS8xc1CXVKDNIeuHcIxl5oDAlIlfJyEd/9xeMlLAr1fnzEZAV5
z/AyBJYstaII2J7kc6FoGCi1GBZasqK/yaCDnqp7AER9lx5AOhcZO8suMshgMm80ZEDdqlPcejQp
V4zejzgCuqP2Nc2Iuz9Cb34eGAcz0s+ov+EyEJNKuJqdWUvuCGLTzhMTr2VG1KYx7gOO8AI9IOPh
FIBTx2UhSiwcQ6Vvh47z0APHnVyG+zdJrPQHGk7UCGb/MlGfk0aXd5phEUGuD1Wjb4BG3VMaISSw
3VNeOW4bIZpWvHYWoC84Ui/eDJBgLidnpx+bpdSKZntckZ0ffq38tiX4OUw79ba/+cEQCY41MPFO
u4WVcYgkDQIKq4iQDqbv48cmaNsXtPFeOF8DETqgTTwVYblRXiDY2hYVOeub080+DN9OmGVEqq0z
vKXJeO1t5qagA9N/2n2YU+GAoZXDYhCZ54lNKRfPuxu6wExYErn6NWibvdrBzZCWq7FQbwwJkU+Y
bha/cs8CrDjY4OawUsnC4ZGL1PXstF9+iTuEGh+B8M5EdFZueR2OFvuGeqAwBeMAsN7Xst+ybm0A
+ltZzI6YhuaV5iA0rYaftMhbCB6JrzBvYZcLxkvjvShVdv1+J+QMKGMuudlATSkgZ0rmUZ1cR/uG
KEQ0vQQvC56w4x2yyTsoVUYD5YOwIXOiouYnSuHCSUo3rQsgIi8pG8eH2mqlZVV02ZEguS/UFj9u
c3pJIC5J0F1y6pLfXJIj7sGlYLIWSt2D2zEcSVHJIhE07Ln/bsxY2YPcoCVtVr3pmEE+0xVjZs1D
N3HChr9fe7no9+NR541LRnMx4/XW4L/Ei+T2HqcbjEVJHPiwxTvQix+PGZZZ8PgSBYYoePRYNWRP
EFcOilUEHV26B+UHOLCvBGTCoKdSXzPCtF9qdL4qBMairpikgpP5gudJY2B9R9C6vFLo7c5WrVdG
OVHpCWbnju0E7VVsVDulhhF7xwKbZutUXkdxn0RKUr67bPzPxor0mKiWr+71pw6BNWB+FkmwJUnb
swzjsWAGcyjneomwBW5K5kirvoVNXSxe0JzbmUrWaJKYOMSVmMOCFDSXXVblZl18U69V+Y6cVCk1
+xLRZeDsGGZTFjpanezeBv6dlTAKNPrBTVTJmm7S4RiuuppO6q6goOtwXnNzP3fLuGzUXV69CNwS
OIwGptIbe5saQZDA9TmdG9mXpOgPVSIWXLwY48FPPA8Gmy/9xayrWD7K/GEJjW+SIYnkHrf6s4pY
BwlF5mIih7FQLbPf0LbT+N+WsypBMUyqDT7YNzrsxP4tiRgZL/PZtmi1Ea281qeFldumReGZfWIY
DZRAZvkRrcovKtTmLmtdhfJ1OXjnpm/QPgd/AbtXfImoc6fnC4OP9lBm4QVNezrVm7qjE+Rpobit
pdJ+F7NlO8fm14odqrcoCFH5zORkyNebq1U98BYtkelT9AVN8J+pyBpiT/Ezd31tAd/mKmU6+qOK
zbO3SppRRkUoLhJW/9glVLbLVufQaMAypFOAXIjMCEeaVE5QYkAZ8FmnIq1hv9TLh6iakQnb3HC7
alMJLU8BQ8ZRbJB3J1T0lciodWWb7HsdO6w7qbhonUJZSbnOsvm7a1OCxOtkg0+gYlZPRKlxo6Ya
plDpd16RVZB0Sq1s8wELlc77ny8LD51OfO5ZqnruFeCdBgmU3OHOYAcL6/ZCbeOZRPL1zl0qa3Ni
eJRFExhluaGVHrnM5mf0i91srDkYYKlOrKiVwDLe2sz5PKyiuXIyOWZfGH1olcjZifeDBupRS29L
cZ12hqj42cmd2uNpBc0b6Q9hCtH4N5yNq6ICjz25oXyjNcaB7XPOmeml8rK04u0wiBUwhT3saqpK
PL+Sh5RFSrq5E6dNAkrxSfLVkpg3YbEFnw5c5zi1ubQ6b09ssoPHlMwySZy+Ll7PjoPNtJ3257tA
I0YPPSy3OSM6J7ilwrCEspwREgsC7EB4RqlQCWtApH1b2BbRAtl/c0vrjRGAyQ4EEuDMYuwZ7Ics
QE51KCRgqZe4pj6DZjjFpwQYxPDs6MxB86Oeov1vJ4rdF1iaNjGETOFlfNltiglIboC3s+LuoyL8
gycpittfZh0qctzJ9rYVfsi+mlqEjsYeKw9LZ0OeyoP+e4eXHWvw1HgZLyj/g9reJAK1MSdJHo8F
WiA2I5xlnMdlbD3RtxWVXzBB4JvZyJrGyPwAUjdPVhs15ePTrnOA+jqi7A9wrIRnRpWxSrSJDxIk
91RgafPpvb41t6cz7Oer/ashh17VheQfAYjwaH9rSXk9ls7jxZPgX5dWBKUj05r7D4Lith/DtLCx
6YuaU8eemj4rL8iSTC18CfFhqBgu4FHznzuPlS2wZ73XGcVHaaFcPIgDt0TYKPn01nzGulWBG9dk
eA9h7urKYqYURtjGp3W2keNN5b1m4d+nPO2iBTZREdfMzAUjilMdBDA5IEq62e27zqmoOqw4cfTB
Y0La5r4ZIB9xW++8DmKeMMxUJ1IvTdahUrsOjDLo5wu89Rs7BWKWMibIh/JItdtic3CcdXW8GHoQ
l+/dOqeECHjm1EF9t0Y40P7fA6Hd0unA92uA5uyDfoL1xgdSKbqGiSZYVoCkSH56ABL3ul3D5BI5
hwb8l3k6IAG/GuIidNNX9s4wpSYp3RZR+zIg79wGVCDI3VWdh3BWsaYIroFDqfo08zxUXR6TU7NO
g1/5OFAWRmdSb7miezl9NL4l4ydqx2x+jw5BvCsFazPRLVoqCesP0dspcZNEvpJ7S4KLLpjHtdPC
MKWj/vV+MXW0GS/9P8/xNjRKIfsaYjN28BuCnFs6+jc3V3aVQFbeWB3Y+a+27tywHePosNE4Zth1
EiXDvOPn7WnccIbCSobEGJjrspqzL8oLEh6ACJlfbS/cZOpAkv0XL5fy6JIRhiuymn4daWYuwFNy
TCTUZwzhdWQYKeu6rwrGxtLmZPl/yFkgXi/8LVBpvOl8Q/SSh4I11VmCD2rTvSM+bPtZ2Xx0V9y7
URzOGtBOf5eg3jsbwU65LPwuXnfDImrnhYLQMf1SYOxLBH0Q9Xskdjq8umZYIIqVmhNgrIJ7OWU8
ksttVXzGvQRrlqDIVvO7zhyamutD4tu6jA2YIYi6LqhOI7WDiIwbj39OH5wqlSc8K4EAJP286djt
UVAcixDHSeNsZizgvw40vB0DNNKQqfgdLNaWyLkvOGiYio/UeUtZUPj8Kbqbijl+FXpJx1drY/26
1y3PsURSZPKIyGm7fNPFDKEisiqcOBiO90v+GEwwlS3KKj6qxYs4BMHjYek3P/NmI06555YCh2yL
Vu0DB+EIslCxgRoh9+oPQENIXLN1zT9I12a3mkz80oWM1lZfki/MEIroHa7lE6BNSv5Kbd41ESZv
JCQMwAYWE9B2BhP8BOFmMDoZVCpa2zpndZtTasJ7edoLmg3D/3+NIe7LJaxl7vZ+hQ1VYuOWnIPc
vmWFdeXJuinD14uV+DSMLWaFcj3li1yut2Wp+GyT3bOhkdqVX6Fj6ZMeWmMmcv7FJa/bvNJaVZ2F
0+7PHljc9G4L0Hsuk1ZTCuY4IDVpIYeyPPAtRiczkZaaXe03KnNfw717He4qZYw+p6R+URZ5G7ac
J+RT9ofVN3nFhkBE25ernkh15CsI95a0efbgivkMEpxfXNwpnu375dn60TvJSII5sd7kHbIyDAED
DId7ONyXikfG2mVSJnHYbrIMvrvbRerGJNu37wST+dtyNe/LMY4QDQy25ommWhEwGPID+fPBnGGv
RzMs3nGGZpZoi3Igfnh+6MUxpoqOyeH90x+GAT8hvjfS+WvHGYh9j55RRSELZDVNYhlGTQ2yCCAK
rcIBq2dqp8sUXTIXhpTk+Z52Cxlw9ZnuyDod1vlRpc6sDAdE8rYAD/TPLhQiS2hQILjrG1xmXFkG
7GiUhBpHzPtOGzpryf1a60UY2z1OApt1vCL+X7McUS9Zz+OQjfQoSc+6o8OLMKvG16v9cvTZ/LLE
BFeRUJTDRTaRdk3pu9Mg0eSBEKlPm4YvIy2PD4p4z+XBme33Ixr9+PO8POWJ+UzlPtU8c1sXARME
cUViqlTy2+f+gGjZ+3wyFy5E2Aau8JZAjGP9DxePr6AsDQ9wc/tUrLAEi1RnUrD0yosj7tbRT/Ky
EDIERYLYwaGg6pbnhPEAI117vW4oJkiMeYCxYRYX/wxx34bcpttu+fpDNuZP2m+JVTgo7mEVEppH
TNmm5YjG7znP1gfvQLF/NxzjREJaT0D0MK3mRq9/Tnntu8WhLZ/CwH5/qBMUBjMxIGTqlNRma7vt
KjdE/ZRwhjhjzetS/8FZMQI8jG3U8QJe2qGYAhAHdHi/+AjK13QYbQlLGsJR+Z67wbdhqNinq8yX
M0VAyAr6bz9MtDuYpWAGdWFoRlBdQbebK3EWn2vUeeDEaFrZ1jUFYZVrYNBL4YT7c/zqe32Po25e
8uSuH90b8MYbkFlw2ghnqGFL8XdsNAIFkzib5z2Zm7LztHPuHnSliG2/GyR98K7O+eneY86K2wFj
qT6nhwC++jyCAabBCbv9jIihwA25XHYw1kqDnYYVsojtx9z6xgJbSXRQWS6yKSBP91KolTQBdFVT
MsGIJsx7djL1fTYJwEBDPZ4HG9fur0CjMoQg1IA4qLQnKwjMyJeqGh0WM6a5RW2mGX6tPniVwMEE
Nj8i78MCVzEk1sLgv9SIu7De4lh99hDAokkE+LzkKdNNNinCRhIx06q6YYcJL4GnnLdsaMK32thZ
s9MDVRtUZp6EgbEemBSQ0+FhXiGHqzzWQLsa9nik4r50Xzd1F5wT8XyTxhxDJiWO8chBXg32pbBi
1raPaaphCb0XdJWQ74LftFCZJj5NfaDsKlvtUZ3h/yhgsh1wLA6+naCbPghXeMdm7Ldy9ZzE9xu/
5T9xd2Y7b+5X/QXTaRN+NDCXErfbRAlYKNQqFg3/4b2La2gH7EDFu4F2jrWCec1Tbhkayeaek7SW
NRJbYuSOw5/sBwS/pVzH5w/sM8ufjntruByeG2N93rjGB59+Hk70wZ4X3hAvCkQu4Sj3xjTv74qN
j6aR2XcXu9GCV9BbC5MmTMuVcK0tiaLBVlz5xKEIqlLXvPgQj9+mh076BottDi+HrRpoSpFCcyp+
KTa6FBAaFxbCFVOQbkF1NFsHINuqvMwuxyHDifJpr4dxUcCJEU2yQqsayJs98Ln8WCMrvGHDZ5/L
Ia2ZpKAso+FNnK0PHrBFIgHlqkOvYCCzDgsytUnMcvb88AtDoKyrm6l+8iSh7zGcX9ThweQSlvy2
fpa13X+PKaWe7SeTvblJsiMn/DXXj2Kmn0TL2P9GkYJ44g5Qid8ylI3dTBnVUfyUXpfH18Q9p4kn
QKxK5ywEzirMitsfaHstIHEPUj1C7Lva2u+MG9M3fH4Cf7jneK4i4unbmFtZirqQfPbQHbQPenF/
2mmEfxMQMvr/rm9AuH7Su2AVBDQKYMcvvCoJg1IF2GuvEBLHMHG9pc7h0pRyVcEp3pzGzwSCDwNu
U1eiRs7laidoviZDhemfM82YVfyeTovyhRIIOcnaBXlBNdBX9VGKG0RwkO1syjoXFKYpyy5sR2aW
C5D/1tc26WEcby0WKlTPNqE4ZNyPoPgzZv9BrX0Eh72/B/+WVxz1A5o1/8asjtYN+5w6OFOxyh1g
gb1RGWVAIWbl3YCB4/G4rw59OcBr6h1cfHNqW9CS+WjTj57v9+Gh01Q1P7IU9014MgzQfFvv8Fs/
sfdVqaPCztmUKAEwMjF+FZfyS5HPSqppJsKg3KFr5iK3fi88vJx0EyJlOD/HENI3sCMAwqbAdBub
xi5ajfCfRefgPqQM1WVJU2pBXib8koFA9hqvt2FhKJymPvpYktSjo7jlx0ctxak5FmwLALh7IB/7
CKefCbsRVFtDp2ovFPY2Ihdu4H8Dt4aoiyHTQgojOUdBYinssfMnpHJ8nlXc8vr0v9pdi2F104Nw
9q+DiMz1r6Y8msU7xUqkSfMiSmgdunxmEH82RNfZlqg5NhRIENft97oz25CxQ5fs/AmDyEibMtTr
s8ibCErxJHm104rDiF2G1Zg7C/3VlkqU24mWszyY4ewtacHkIVl3BoE9o/kQ0aMvmT/ulkAXzrDm
HOJco0/FFkLDYMANYoFQU1JvLx6WLNILZBro+PYACDIdPmyk4ezpxVWw/1o2q3rLkQjm2doVzcuE
ydUI8vvYfbaa6FInbrQPfX9XrlnK71MWmGa2uF5KR20HfqAasOURIrgJVF+8bz6ml7slKqYiv2GE
wSrqqdVbLfbXxXr3X3ZM20fQj4iW46G+qYyALY8q94e+kyruK04nHk6t8ofSupYzs0+5ll7QIDnB
p4AECEKX3N9w2xI/fh9uXf7nctON7Hd+JfInbqevuCPi2nr5tICI5L0rB5ufcNlXQs4HVyB6eQeB
n8Dww2VwGkt8AZ6YgeENbDQs9L0b1ix/f4j5JkGBUqaU4nb5vao0IxsckiVMob096MTZJ8U6M0Q3
CBS9HwNa9nbnTF3XqYiNwVknsi+t/9gqLSpD7LeZv6DI4RGr8P/MNuoGJGHlsglmWk3V4ioYN1Rp
0sd567aTud3c2mGqr8pRQd7fRuuRgGOLLlObrDATKJhcKlhYind6JjHunY1I+E+nEnhv7H6iv7wR
8aGtnMowVG5v04B13m/n76W4v14R+sfMg6BsQ36Hhoe2Tt1+crP8jn/Im7bdunEy0xP7UyY8Bojc
Qr361K/9KBvd1Gb/jVa1UyTiL0ucQtiYB/iWOsC1AbdU2BLav0zkTeYGFCKIXFMBch63q2UXqVia
8i8Y+w/oGDy47m5tOiftuM9kdr8C3AV00ieog2y2fS1vO9iVSc7oONSVmtr1zTt+bM2MOOLmtmqo
VJ/Vb0Cd1y69N1K0buO7FLyEdJGRNMdTfHduVRJ+19WWIdpE3aTvzPDYf+V3zAhuMoKdYakuBPQo
uiu5RikvQb8r3UcbIoCQBqcffkABVUEgSRym1GoSE7J3+3bT3ro6mCHseJZEU2YrONAVHljL/h0W
3HkOh0gB5eSDtOCwFEZvG46eTEQVA8KBh7rhL0CY4m7+fxF6R6q+nL5dK9U5d7yZMiFAU47F1wRm
xwyd0WikT3OABlTEprIPTjUSrZ5XdSQkQr4wrKslQyo/t11YA0yeudOjta4Nxf99UULozuXIQYVs
mp2CnnsxkZOSonZDPat6P2SEkzzZ6PFkeYE9arQGMDOXbSE3wIuP++rwEeD050w9sJY321uSRR8w
APNm5CoHi5BupK9VA+HxmZ2+Jdw5ExtdpQgUq6+iYbdCbe40hq1Z27xoMCcV++WfiZaipl63J28W
kMpPXWxvUkJQ8SvRQf2D0cU7q1Qv/mlkho2lBuJWP3lnFydoVpIelpweS0mYk0JVdqCV8ew9KIAZ
KV0FOhxi5Ug+Sq1warbjjHW6PH7ZPeHXWLGSwgj3o0KeSvhnVRvXnYg/HXKRn1eZNHv8NaVETVjn
i1p+BsYjOFaNXurzTbwA1FNcV6hnmWltDm3eq7oSdfkubwzGMzudFLRcfRL4slBhu5Ecqel7ko1t
TAHdPbhxaCP8jVYXnZ0vqBHWam7iSN4yITdEUhUTLbhAL3jiAfNcpdEQJWQ4fXIc6razEJg9qSdo
VA7wruK6lcqaw1paHHEzImXqnCyS4VdrcHhBLaXITmSDtc0XjvdJnIEPLG8n2b9cSR7eBZut2pC5
krcjwTg0HZaGXhx06H/pPzbQIrlrhUltMTU1U6xlKqOrB43f3Mll5yYYVt05YGNmZ+Tmjerz68mt
KB8KVP5pJKAB6+CFC7PIUf5ckqfClUqR1IUzZJOzZxqrhLnfyqz2D7JypfAPWQ8GMpUH+ZaXWVPf
QbwP/T0Hro2Tx5PhNpkGckUQHWorXSNSecDjL6GDCuTk1+LcA/dJ4X2uYEG1oM5xo8tYzfsODe36
RoATLNqjaE7xGY5K8HdqLoOko+XjFXRDxa1NjnYiu/xeYAPmj2oBIyRL7LyzMqitc9QV4jfmH/WJ
ZgpbG69Y3kGb9gHtO4RDHfdCSyX1y0lcuNTxxoVYpH6oIqDlc4jGX542U6UrIBMD1lwNn9oBRwZB
KlCfiEjppxgUTfxL5AVEV0BWBRUVDRMZ4juXb48UrOnbX5tBiRsXuUixNoXxvlrcgrUPBh3+rdWV
q34n5HuzpTplnmYhFOjqiQaxl0KmvKkdUWCCSr5wUT2ypatpkNsjiscAX0Ye1PLHcYSbVMfyyukj
Gyu2iEBCFqYKFEo/Q/53o3qEvv32XGpHGUbzO51Xc7lJXJqnn9CAX8Tkdgq1YHHgpjOwoQmeeqG5
t5VGhTzZTUSomMD00MYXkjFx01hJMwYCV1T6PEGpfoL7lbMIG4EsRBaMMpDycMOwmk1ZmgUtfa2E
MvV9Je96w1Gi6K+i5tlUZ9E3RIlEwz5vEAk++jf+LdqZmvIzcnID0VfvM/V7oGqk6ZBrMYTUYpZk
8HEEhCxadyT09801WLTA9dJVpGQwp+tVaAL47oi58GWwV03qx/EwWZhnjpQBy0DgR+RtOjvMbldl
RDm4urK7Oc6XgU03+JXVU4FHht/u43z1i0tE1Rh9W8a2KGoKbN75f0nztwPtXrh7g8X0vKvDF9mW
kZylZThUyFSm3h4pSupfYahDH5D1KzEZORJxYj5dgxa2I3MdQo1seaOan9PeuT0epWmRC6+ipW42
lKuA4T0U7/sUfhXQ56CbTOq6au9rkesjbfMKieUE52NIXmiYktLUXDxrldqC7hRJ3+zGtAcOBfPr
CZlsAWmRUjlxsePgSNX0Ink4DwypUwHboZ1+NYPyRywKu7DaHk5Le4+j0KBIb6vBICDF/rVSQBfC
uEtDFAmrNJGk1Z/WCO4B6o84E5MM+VVII446leBdFDy3tJEOjNHxpvlpzio/fqjOzJMcIs5Prim9
QtkGmUnC2OpNDstig2GSknR9QnkFkgemkXjQC+1Uxs0NGGJ5b+iLKKJsRessEdmWPh8OKakg7eGY
ZysmzappSkRHCwj+HvRi3ofrasso6BBD8VJCUUiUrqgdzqEo15BlguTjs72HxDZZpo9bkkC2c3s1
/Ejn7wq41uHRNa6snyZcEmRCXbnqXKVDSh7JuiAviSKVpp7P5ANYHBaHpwBTuR02076S2Z2BfDBX
WhKwFL38m93fjmL1ta4Uib/zrJpkLTbIr1cbsJnlUvrnNOXPJd2gXLQjIbexLaSS/GvQU4Se1z7t
osGbxO90WRH7Y2zhRaUD5WxT/Rk1xuuOUwzGj4v6xYsX6mGSvpR8RuW6qiyKlT6y7FBTpkAP5qdL
XrBghlF5OxMvr+cMfbshGKlEl40g+1okElNp3yRrf/lOjWffRQ6+se+FR/TURbu6dXxMUL97FibM
b8z53WEKS5YeT90ordsMp7QkXQApZ6eJ3Lj++tBxc91Z5ivmafwI4Tau9W97yv+SCJuKAZ5hS+7a
pvXNiEe9Bg3/oKw5GKH5l+rcdk/Y9lB7eR9DZi9c4PgUMh0SEtk/qE0dPb9+tCE+hWPwhxx/LGN2
sgSkGm1RAjlI4kW3AfT5TSOBbJjAOoq6wn/msVx4Zzbh8yo3p5PAiAafKaH7nJEG93/YZluf01/Q
RXMXnDRYHthkHa153aUPaPKDAigtWo0TEivNSlefy5QqrCKNE0Vp2O66jM9d6QXD4feTnAu7fBU1
Pg5piHYNSs9RDRKfT6rJcAFjcCgzNIxcuxScYrMHzDVt7P0EWoT7YeLPlTDcRwP9iSuloGe9be9r
/CFtwlLPQQYSdPmPMPWzlcs0gaFdmGWD4zCEvZa3s3eRLpCKB3NpNaeeSHp9jLfdX0TnsuLBpGBO
j3St4JUNJXMn+0HSKg/Pof//OWKUPhuu+BsFo72ys3pJfNx9yjDI2A4aS5yEPR/7dg4yI5QMjzT+
ve7Onidx1YydUlhayTELILhv7guHHUE2HR6jD/BrlWeNgD4L47EpkOlWoNKHb39tJHpdpldqSWYQ
n23JKF3FTxhK6ZZUT50NEJADY+wh16CLpqMrk3BIiQCMO+GgIi6VK24Rg+Gve+nBttz42X6yioop
mOwBHx3QcNTjzj2Lqd37fAAHwB+yjsIGLbowRFkl1T9313KtbPWxcdnvZ2dkvjqWEKR/wOwiv7nX
yuYoI+JdwwQQadye4lEr+Hkf+EuNUKRLJ0gH/+uHGzRWBFo7ycXM3UIlmSqYEuasKb0x3e7SooIC
WRS/BfIfelfH7eQKfKDf/3VfMaLKY3xKAQVqo7SeviQTMVK1D2kJ27kxnuP/TzbM58WKx1idjp1d
YgJKE+ftk6lHRhvl2yuBzjy0jVNaeBRaYvCAw2LQlYWEHUnPVW+TOxsy36dB6LgGZdHUY7eVRDMQ
3N4JPKee0VSrAE288gpOglEHhQ7dKn+XvgPCZfYJX/B9xZcV9u76cl9gZCXiN/8sTcUAVlCmdXiz
1aKfeY77Ll2pDK6pR+kb+hWIy5b8z2x+7LcXSuqbNcnf7WkrJGSg93xRBmugztqAzJl3SxfI0zZd
EEBfwueycjtp9raGIKDwS6XJ6Xn8PhRZrcYW0AJ74oYhlWcbeBxb76wH08uXgr4sJyVy0/5E3PJo
/dYfc7L1OEQ0TpgEyyNFspj9Kji5Ki/1hIjePbLXNV19q5kJmfcs5jcbSKJO+uH+zQistbWsfOIA
V3/2oGz+3qnRXD8D7V4mot+pqZCJG4IxKcsM5I9Xa5Xto8+EcZPc7olN/d+SodtfDQfZNrA+wzo3
zMap+0InRORnAAU4c3CX3qIbjrtBsG9E4Gk1DB6Eg4a/c4plc74gJhi4ogcFM9Ow4yKvH/ENqob8
X7caY+ZQmBDvoFTJOURuX8aBdKxwvAw3MkLUYlNNoH4KG19ufwSIsJOVKaw5gkKO2EJTG25Jp+Kg
+Sc7yQfalokkUDxRW3ToXX9DLPUH35MjsqkMADQg/C9OU1a6NyuoRfV+OKHyk9WX0QfpisRHeC2R
QlRNBVg1H0sqqnBChbj/sY/tt2wutHai4akc7g7mjD+pe6S3EtBymGJ2QQMgMtbWUwU/TJQhgHS4
V70/zf4Ew0mkZlnEAoZ2g0Tq5/yeL+jEk/4WXu+646w4LcnBDTAxA3a+bFWin5Oha24qTqqmKoO0
dd9umjEpSwMbrHY4uUGgybQOLsiwuSXEGmaI32Q0cX9zglS/QWZ/u2TJBqxK+M9JdtFBGXlRSxiB
DeL8PbfSv4nUOeO9Hi1OvRxfyFUDta/myCzHC9fsGFdMTC2TU1ekQ1JOhHgVB1DmL5uzvy8ugdEZ
mM+q/A1O5EBpqzlraeRtgHnyh8rA1vAuQHs7e39Ko423zsTJ3RUFGzRljY8TcR38iRRaMTr9Z4wj
/5mnuIm6YjnNNsDc/eduqFpB+yOFyNZvUABDKrv48oDDjYpQRHSfeuHIZGwTYKc4/4A60c8zQ+Gj
WUaWCl7nz0We230MGdf/AkYiJObDAwE1/XTPtH1kZz4dRGpQqHfELNN3xU2jkEGnHz/tymHBdeS1
beORILdutEAsWATHmfWkucF0IuOP0zAEVDwjPCZhXfNnUntuuDNVXOvB69ok2LxveTHaR/yjuc+R
PI2xAK77KhpBB1TKY/rIS4BndyoW9+K+xU9XoUeq8js69fROoZMmRov2o1nWaYNgyLBElsPDpv7P
XLz5+OsBn3O2NSAuFn+/qmHs2lnPVbMGiyUN06IU+zKsD+4Ef66mEt3i4z43piLEw3E3JTlK08iB
Fv0S12S8nnzAyD3g5io+v/G/EogXpICU2ppm6mXI6Jz8/h6v4eJ2r8SpbhAqgHAr6G9J80IsGeUw
2vwvsGH82vHrCHF5Fbmkg8HCdOMgmt+n8ZXZ8mVoTjZXxQHXhGNHEpXTjBgte/H6UzQOAmOKkNjV
v6fVrRXKXfnIglTycd8u4+NxuqDDxVQYXowXQbngltIlAqfEdv9bgjRXFHW4ZjzakmWycVQkuYYR
taW6aui6v1O7SjIrK7pDdnUpYWyiFOLbvfM+Yqp7FEZIPBccIVW+M6+JbDvTgretuWjRWSNHQt55
XDwnmLqIH5sN6VDceHxQXTETpIxXuy9XghszzDEg8ArLqCftpMW5cJ/zHH/AJ64+4rcfOUDtlp9D
C7hf1kybKVnyQfy3q7JC1ZadlSbV/6YRp0062SVxod2Rbi4F62IHm5wplxzWpm0S71IGttXjVg6y
FZkHHAgq6ilNnBZ4pzbM7hf0cC7+TSFX11wJcbuC5WkrZ0LIUt7im+lwMTQYGJ9HqB5iw2YlmEdX
iZAxnOWe/3vdhpLEUtm+i+a4FwU0t0PV8JbVxM2SJU3qK25L/lLLXg/7zaKQUwpCVuV5rzZLhk1V
rPhHb9GCcv1TB0efpatdjFaLvXJXpB6HqG5p9N2thiG2Hiw+xjX5infYMi8/1Mq43QJZwlFmsgIY
JV94Asoxa53gno8+9PRYOKIHw77F6JC+sfZ36ipgXW+xJqpzgQgJRbc/sY4+Y4NXFp50uexkPni/
bPkodZWlc4YeMvAL66/XIsK4UUxyHbuA28yrSG16qt3M8jTzI6m+3wNZcMKaGQ6a2T4mS5Po8WIv
sBtxjxOz0+oTaqY10XZhcc+GRUgNV7PlX1PYqXm71dhGNVP1o6V9Te2yu/ULg9/0nCdogoXCx23X
SHaCH9vEzFpccuEtkDQ0QJ9OcKe7kVEaUsBWZw94nbjCfULb/cG0tLogedfwTs1Ft4K6Hf7MAU8Z
XChYroTZoDH51ob2rXtNS5p8Uw+lYCh5TM5Mb0xx8aYQtPW73HzpO1n1zmo/6qDiIjl15cJJZXC2
+BjlczqBGh5TWqLfbYT0MqbBQ1txwmrxT/8UZjLhSaVruVHY/30Fn6mS1GDlZBxRlKrmgMrlWjUL
NWV9wUohA4Z7wltSPQhEW1K5rD4MOPwb0qVhhIx/Xh1wqVClKHb9oolN+57xb52jxwWt0d4dl/lk
FCuBwRpIox/XATwnDp2SRnlEvExGAWDHHL7uc9YvRP0T6Pza2cLREUuo1dP+9cTmWUD36Mr4wZLt
L5jMorYY919Sdryx6W2itPpW5NVkZMZXzRpjMzrm0KcF7a8lz22E/iofvD++ZgEwGkSKUqf1xiTK
7NIB7bfsl41aWYshLdp5be5xcKeVdxdEBycWC+cEgJwDkEIjCO4hQFh4niubW5cdsZDsleA6XHdI
bWeLPUQn/3Fbk2wQnqByrO3NU/eb+R5+9XwBwN32pn9FfODam09b8VH2jerKsnoSsNFmGYXPBvmy
Ia2cHaTtAGu1Szyz+5mnLoSrQURAlWKaOxwtTvwlNlC7Ub6Z4HJoEUHexFuJurET+RbBWj+GN60N
hs3Eq62U6WEG2W3yJCuym81b5E1rR3RYpobFPlp6aNnAJohEo3nPzCWF+t0mWiR7a7N9IxY8t0XE
BlZNiz07deu3ZILWt3XjhObtKCuyYvaHA5ov/GhkewI5alRAaYT3UQveNYkHPVcWmYd5T9UKZAd+
NRcwCFEo+OOea/9T1rz4E4VRK/lRha1bGOfpvtkVUl80uH6NDbANKsF/vDP6S9JuJivAuMTuLoL2
Yf0ZtEGus2p3qd5qwag2usyrRtifpKzjMIVlgDVZeuduDcIolQy2tw/Hn+b7FCvm6rXgQn5TUfCe
8Z6HYgLuV0XNJ8Ctz1/wbdXhfpvyh3FkT0DRG0lU4o6LWUkwJZ77rbyVbKDCbhGwrLbpJeALbTYU
ArWCmzEJ2j/Qp8XK0vPeDgTxVdun4S+AdbUv/Jd8pIqZ+LPR2v4xSC0KiQztjJOIhGFeJ7n+cKr/
3umSuC+JWS0qV1ItJTNHNsbcFjNmWfD5qiA5QfSUxLMtB0gATmAjYQnMGXtQ5mbK7lVr8u1vZ/Is
jUNp1v8k3Bd3kv1mC9TSMiiWWvD2acyTjXlpdKpJ8UIT6mlLpKp+scHQygvEuelZofuI9TNHmmVS
Tn6vbv9BM4vkZ4zfmLLOg02xLrczLwqyLdXKcIB5R4w2EbMKtXd9WQtNBnM8ON9LHoS+hyX82Bxl
5FXjIcBZFAueVFs/guR+vil337lrUIyvZ0C7/RyZUrKD8IwtH8xLWJdF8H41TaB2T+XkjS4cHjGo
Z9wTLuJ4e5NPMwQPe+H4IcW34bhb7w39mlnyfUz/Fnn/vjTLHZPYK3qHlcHkAionS41ubc7vmFaA
CUL/qC+Lnw+25YZxSX1Y7EAXliwIUchPWGHiNAfjFD+AOp+WHzLE5iipTOOMT2Ph8r0z2azEDOAG
YFt3z30bpzr534CjsxLQUaSm7sz/C+O4haNciXdEav+oDzOgRRsbJkDjLdX41BSLS632fZ3r+Dvc
2PrExY4c+/nMkL1J3e3HXy6TGtRyk85Ejz2zbOKbqE04Ie7fpT8AS0uzZM5WKD/oMUa7YWMtvOee
foJiRXRic7C6LJaKGec+SXiq6KJKzxUq/0TR3Zc1iZk/YDo0jXcIeG0OLxYF0fJTRPWzGMRQGYP5
agoQ37JyA/rmjvQAAX5biRZtt9XGmdjGaKGPN0EmNeZuKPgVExvXERe7nu2y5wjidrjAYoU/TRXI
SWNwdmxCGiqi0vpvLFpDf4kf7nkxEU48rwWy8sBEQbJQYlbB92F6Eqg8gq76Rp0u8bg02BYhC6oY
JNu0ENXkWmc5lHR0Fgl1xqDbrKxprWAU7cF3AqK4HpMdZEClXwVoH0+9ZRQNNOk0oKukLT14SsHw
4x8zJdq5OkIsJQXDFSkI1B3lK2xfBuWii17RKje6NbHcxZR370vgNS/gS+qZarjAsa3W4zdKmqus
XuK/qXmCumZx3llw+9mwJi0hGvq/riuIihnbkUCk1ZAbdltftMCr85kZf0+JKW90hj7MDdBlPeUX
i5PRea2BDFu2Jcq4h10KSRpUe3rrquhyRHEii0qwqOxPRtf+gRdY3beYPWTD7MbdGKPsVAW63ku8
JyaNxpr7PlVyFjx37Ll1rBKICLA6hX0wnCM1b68OcYwKgw8q6zPfMFJF9aHI/UIbxEC9WH2DMOQV
/Zc+jDFYhzvo2IxrM0VMHbwKhWk4rCuWr7aeXKYDXRDNAvrzV/ncvnVXKL8iSSioD1HAhdmmU2a5
GvSacY9KL5uDdU+e9iYn2tcZIczZRYS1ElsdicPoT7/ilIY7JBXXUBfCQs4q/uhdyDSwbTqpDUTI
d7nduNJm3/43XuIq4zUvGvlwdb3IPDqlKV/p9DUujfLeLIJk56ej88MsotRtDaLS5eQIcTSyiKKi
2MVj/NBJAtGgVpV/ptoe+av4BGtnwTXBqQ7tMyfKNVpfjgvIBoMQVSAzJkEYKSGVPbNmi3bcIh/K
QGHpyuGRN1cNvFZEe+D7U2EzC5IyZe7BM2mKLoZDSAr7jd778lKPK4uAYKM3JYjv6jd/tHHMlHV3
pFBW6tNaBiFhyjVGbgaU+huKdSihvLNpLDeJbMheEvZ7XDcYM1Uew8aJEBh0qjuA0jaiYOH+wOe3
hhqgEXDje7mMqJvNPkGai3OttOp/+mLm+H033ru6TtU8eTIvPDJ6yClCFstxDZWaQNbSiPzl1Cus
OvGBvuXYXZiJDD2kvE6huDyFfyIIncfSBloqs3yIJrSV+1XqXBv7brM6UvT+Z3BrzADVTq7sEsJo
bu7CBalJv1EeKdER5pG3CYsV2ZeYNM4XMz10BCZNhOgIYub6dnz7y9OPrY43nneo+w08L0pmqi1p
LVcCeL300YmhUY9T2bz0h+i/A976Y+SoVrvjPCROAcpHk7rggpncdaXC3TyHZCTgw3EF8bI84FM/
pk3frUuu8QZj8SCDkPg5uZRNbB59ToRPYJeZzKGeMsIy6exMctzdTOakMA51R6iM7UW0fcVItthp
0VwSFa4H2F/AnSgr/S5tUGc1riuN2c+dUS7u+c/DCxTukpZFAYhiD9bxnvsAXJUyrShDGGxDE4Oy
lDu4JLiuhlZMXe5aOxR+R51+vpRPwYRRmPefERJNZBt7XUYRNojYL1OVkLXIDVxNBJF2GwkLtJtf
PvERb2nVWl6yEOBkHHhoMVwI0oVONci6iJe8Fm7cUFFpNbrpqZKGpIrcWqmyObrSwSFyhc20pWVm
qacVzMkQQpQxJpBYdrSO9j8lvxh/09ftV8UF7im4srtwW9eljoIN3dabhJJEkYbNHLu8CXBdvDMz
f3RVzLmKuPYHulWK3aqaPUAF9jcd+lCzkovOUK/7qarrwdxJyfR3kpFUiaLsQg/DloDsQ/gXH3Wf
iFhGcHN4aVi/P1DhT3FsQ9frRKGtSJ70DecbeWzbEI5FdYqR5d3gxuhojio90e04eQnvF5UX4/y/
P2P/fz0Q1O0OGQcvKateczJz0R9P+tMR7IZQDlXbbEGihrsiawGEIcFF1Ghaf+WIBeL8mDVUTMCp
bX5XhwjXssCdejJk9poBRlysP7r3H3Duv2YZPhYK7ISDU9459OIZx5sookja4v4thcBY/NUQvedz
xnYAwkkGWLkWvmO0yIsZy1t9uARIS0Qz/9xq9A/iBMP0E+HYqz7kPPSEVIKLGwnKJIDUYdlzEQRM
RSMMvdNc8fKZlphP0uZTendezsPeT4gGvV5Ivx/XYlvExC8QA/US0anLg9KxMjRoBNnrvPe0zXsR
8oycxPMYwFKqNHbtVxxrBOV9MieQlMyq9kgMmtADL8nLpe2ijJ6fcC8XJtIo8VvdTNKmE4BCCUHl
xeYfEe6rC57hlFTcMttaB3J9QEmMeMekqw3Jhr3UQA8GMVnT2mQvNTF8QBtfIprW4SQ2PosBxVsy
2hdy3+Sqy+UdNxz0+ICCDpsdjXjuVE5Lb54kn85YC0/T2PqTBqD7x/SI6fuQ8G6uWmvChDHw3BK2
o47/ycOMqavpCEmSSznZPl4wM51c1EZ5m5PkggfBLa7sbdKUIMk2aXqPF0MPh2gJLo9ThIAQlaKz
esTHIYBBKYOki4SIqk2c26ocWmOtEmglq6o1CEDMF+RZWP4Xr/EeJhiCWJ2sMGljLZawc5yHXeZ0
+rbl4Q1gOykqDrM01GnSHTDNtM8Bdaa+rvrkUisohyWyJtfGY4TqIOTClGGV51GwLaO7yuz8rVyD
FH5605xTOeJiGrKXQPEMfhUvYrE6/pSuKTGxmaaMPyPOnTxhwTsJDyC3siCP7FKMcW/0gpgw9hGs
r1AUvMIxCirIxHszKrPLId3wRwQaCEOeAbdACOYeG19FYzLIdEHU0a1y6ES3ULdOttQ1r8mogKFQ
gCXQCYgv3iL2k6RqJmnrZ4WjlbyJtfT91+vnNBubMAEP2WemgN5hMFrEG7K53xW7a9IKAdzd1wqL
zQeE3HeBoAP1/NcnwTGUrTF8M3UqP4jdOX4+i57gyoAvkBp28rWksw907s8pNcgdNpRrFq1mtaAW
6x4/ZaxgWmF5btdyzGGgUcagmE3l9+vJuoxdSFnrYgronsTb6PmiOiiw2o5K1JxbqVaEWFoKETeI
reIKogrSyfw4B5z4p/a+7HCD0KXhKos+J1JHiDmYQ9pRylPB0twy13WkjmBCZGHNyLZD/apgqAkz
XIiN3z7Ghw4ut9QGWbkKsXQ93koNjHN1dajYDHqVXOAH2ASsY7hplb99wY6fv2pndkO2XW9aYmgP
k5Q2fplJ45Yt9GIJQLNszMLXA62SUao5ZRGY1HpMiwQoiJkYrBYgWSlYxQbbP6Ewycfp9KLyurNm
jm2+lgdP/EHlr/cMy6wf3+FFHpMZmwllJ6Ky4qtzWx05CdgU68qEe62ColBxd1fk9X4sSu2f9gZ1
OQ4e10fCxRzsvDTGwDnkI84AozIEOMxWLXPQtcCPOIuc839OaYibpdlwiB8nrUh8N3DjoK7mBWfJ
64g2With5k0d2Qk4vXUH5EqecoInirF/rw3KkkvjneUQscjOXpm8Hefwk44yOgDXUI/pT9dbhJ53
z7zWlZ24G5179oqvxVuMmrorqFFgYZdpLUZ7gQqnSqqRQLBspa1EFmzOrr3LdZWtG6tffi3/qNPl
k1E8SSpxa66CYeG7PmPVSYW0wQgp/2nrI5SRp0+7FjE3FOvTUw3bYL9Cq+d/En/8izotnJnrr9fd
FmkOjoyK6oTJ50myeAtMXB+/Yk9eLu3plteePYeGM5QYZTOheK6LSzc+Irqdu3uBVnAmFNsEu/jj
kKOcpqkIAdAJKNu3eNPgRiBLz6UQp1NMRKp2hQgkPdWeWRUJyEgYNJTAKkmX5CIV98CTTBXBQjPA
H3ztIabpuEGKPEDAhfv1keZA+JoPIF4e6Ex/S4uNjSF3ZGI/T/bJKIYyyGTFWFelO7MgA+w6KGVU
DTcpbNZLE/VF1sk5XWB6CYYIrtblOTEGwwlFfNEktyiLREqBm3Pf0hoAddbLZG2+BurMcj/KVVO7
JE9+DIHeMBDzPOJfPnBfopX6Uq6BgckB/RkLzehiUhYPhhGWDKK33mSbkR6ZUkDGN/3XZnZf4M9Z
dT9SuKbYmUBnlTRj060JSdpmyqOV8SaLE6pxK0QbwOq5PlqTbFsTc11pCm4Ku15zYW+zijjbmk1l
hu8aAcNG7wyG9lIUAa+K1iUDhPcgtlh/y6erNskwsEW9gxjq1f+o3Rt1jel8QImhu3Z8h+MUFEVY
fS507Ig5p3ElLC8qhfyGg1yoKCcCO+8/e/VtvCTknh4I1yUsaFtxk1jCP8PRZZJmBVg51b8/TgNb
yQKa+AUXSjBc4qx5ehPeaiQ0wmos6S1oys7FPuEfndDDgYEPorH+0/85C211SzB4L7m/xGpFNsOv
N07PsHsq4Vb5dgkarVm9y2HdZb0LQ5fRcw9DySP0gWk4KKqBttKVxnkLnx1KDKGxvUJjPoWM7RUS
298xS/bUREizGbx72Rkir7tRfE8WuaZpomXDl/I6seQ3KnrPcEwc7I4o8he5jlRoBGYiRDO6H9qs
vaNnpQVfZdUZj4bO/lP7649BjpztSoxV9wkaaxMpTCWhvjqVSBc9u1+SBV7eForcEzR3MSTJQrIp
FrGMelDtl6gRzhXJtYRii6e/pJ1X5EOJmkvS5UOThZGVrz6siXyeEdZfhRPnn6MzJ/p74Ra7PC5F
JM1w9w1cPsUt+P5qKJ7g6jLKbwc28/3Ga067Udq9N/V1fTaJtp/PT5O68FgUPe397otJOWjbsvdI
COL5VqXxXo4E2WdB1TtJbKJFQRc+GNtnvofHwmn2ZIRseRKnh6fl937Fn3cFcpMZ3B01BjTXIgvs
Hah6A8WbpX1fzH3vWsR06aml2dF3gD6wUI6vMFwB1eoD+F/bcpI1aXgfp0FQgY8Cs/i1SZ1105LN
k3n0ffRHRzUE58bufvBIBs4QlAVGJ3FMYWeXpSAJThgXnUY+LVS5DNJtc2qqL6c7h6QRYxELQkty
L/nKhr+SPQcDEvQYfPCSCB2dywSzcDy+D2jKoFJEPsl9HL+q57/y5++fLPAk2GwNE6pUal9/NZO8
5FDDsqofOgBJe9a7tFglYjLTnlEiEFuAoRznlGR4bSBtFfPrxOEuS5MK4T2idDMhQWL7y2yImJSQ
a3zYrx1f/vsTL7ulmg2gPwQ5GarQAARYO/rHbNDq5aJgxJaJhhtzY1Bg30VYK+nxTjbY9t2fCSLf
u/wCMknO0pSfx9JYqGBNL5MFtLV/FEBt+ejp5OJ/VZ7RAv0yDA2QLj69K00swIU4Z9sUseOYsx4x
JFeEFlpDBwDpfKsOMcmihT9z/yw0LHFmWu+iGRiaQjB9jhZ5ODlYY9ww6SwpA+dHrXLB8fwXheaj
3m9mneoDivmp56MfPgxlsfloaBMD12yxOk7kEZ1V3X678rA2ehKiCHRZ4CltRBhHSLvokIc83akZ
ZkpG/EAmXrefIIaRj3XRClSmrl/8saaq7vxjjUwCjJ7qCKRo4n0/6qr7Lm+Ck9yXtP0NpvfYCNh1
rb4VoRmtvWLdH8zSPRXh8iwXK+p3lNQpogWQ4m9Vkig84vlhbgKEfSpcmcVssREJNAWWaD4BTUB+
DopH68ve8h54629McGzd7JiPo51r/DTe7WtEf+j5OQlP/omMkGf7UJne05YZtvANG/t3PmIlEslK
McH+vPDdwBpRf8ZgL062hI+cpWSBcRug5Evcg4ShkFiU62C8NimrzAZUAWQIxEyaDd3QD2UQzoBg
J2YaFYj1sV7Yfgy+uLQqefU6alpNOJKY8upao1bV4QqcRXBf/0gshRRXyxE78Tq1Q1/v0AkZbVHs
K1SA9ETevYTgFyZ6m8t/Rq0xEGq/mUn+I3niArEIefZdHeXz9ztQlQa2NGZNNSRnkrf6srJQn3O2
MPHnX/fbiDVGWnLcQjxbtZkKi4LRw/4NLCml7+BpQpavYF4+zpt13tZfHiLuuX6BWUxHs5jNUsLz
firohJa9ea1DceFqEoDxO8dV3RzoACF7+HARnFXAAvtD9Jv9L/1ge9yKULJBFWPBwteBKc7nll6V
Zo192wCHe8AJ2YMBo6tjpC/oUaMc6IcwEnv2igc7vObzZ3nAhfmNC3/dVIVQNxRp3pT0oHCeOon3
fbEJ8jSto9ZlHfaoCTi4MJWbkYJl6vR5wNFj2Lfn8Ew7riVQ55knG0vs5gCYS6UXils2YyOOdO5q
GsVuGCOFgAjuOvrXOIpbh1RAZ+D7z+2Ex94cpNQP9B5RoJLbLr7HSLrnOmbr/wI0clREwsJJdZzV
HvbpBwR6W313g9eLdsYsQFoDZhWCRC7xzOHeM1A8ksOI2ADfYQqSZOB62SZRTEhCZivoFmtZUClX
o75KBg06c19oPI9mE7OHUEGw9v842m+7c3dQmot+siApF+vtq9MAVhMnWNmxhNnkuDis8uAHXanh
xo2K8fREv1j9dtVg0Cw9V0qTG0mtzjAcu/9g3bMTT+HHJyWX2Zq3xEJAPDtlQ/A8LDrbwZzkfdkN
VVVRhIFan9U9Ls0AEfrZ8LMGh3r/hNWN0ZZEEp3AJ9rPk6T0lwUKEuTKsfKlmcEwGh0xqJDJ6Jjp
raftV04xqkuqzNq0sVuBsQlYuNnoZjpfzmh91F/Gyl5tGfofe34iTZGSeGoerMGKThWdGspzelyJ
RNVK6Z3ILnr5J/Ip1JSIqd9yADR8bPJS2u1Dn+IQeYzdonsH1kznNi9CPZaxIGE/gQAfPlEc8t4h
PiwFIgszyjh077Key5AW2KJQmKPSFlVXLbhvMlKoxGpNBrMyqnpw7VarP4s/qJ0VoO8BsOwRy/Gk
snpf2NaTyqEmF7GaZ81ao4BPgOyhaMqbqiT6FZTeGwfxSrz/dKs/gLr9YaT64piMxK687C8AXCHS
yvfuBcmTRI0jzOUXmUWVyO4tZVA/hRrAePP/7hsRsoIyB4fKQ3LhYB24UMYUa71TwK3jTxRiI70n
2lHjlEG7NgC2ySAJk67/J/Zctxn4K0RnP1UJO0aqWhrdxUPlfj4DMdZ9CXC1T+4UQ+i3mc/7yS/q
cqMynTA4oB3xJ0WYNwJEqwK81w+37g9CqcaZG5ew/qL1G8vxE4vbcB+BkQSK3OCHs6YR7j55WRN+
fdkio08fZGwGHVbqR8Pib9MOMPYMkWU0HjoOJGI8J69qXu1ij0MdjkzOyeuU5Wp0K0fFnrBvpaIr
SGPEFFm3x8JQZZJAoTFenzbBftcdtJrAV4bhGQ6QS0wx08hqk+XLh30ADdc8oqzKh9pHpVhW3GsS
OHVwI+Pgr4zMocZNvf4+FuVywr5JeRYBbdFiinEJ+DdvHfhrnnbfjf6kzQ7bAQKlQ00dc0cE2EHO
yis29D33j1yUOEOG5eSJu8dlqS5DmZ3FXWmcq6peJxNMHbBYfejCg6PSx1nROKctFMniOEIGxHkm
5/3PV3tDus9a9ol/wIhHLwQNIUAYzSf6JFc9UUB/zokYY8UNYBTDUu47XvDmmPG4bDP7t8BM5fA8
6xfq6jpmdXXnP4YSoxUzoW8lVzIoiwq89TJrID1TF6XMws77W6mTmP3jrzTRxqNChByRjWCnVbRc
5CAoyAw0dd0RY992Ovv1EqNyQaq6un/WJoG0AE/48H7ASSWGED37C2DbTg/7ueW0yhnYwyH2qx2P
h7rfwZT3epJ0HoLpx/3EMU0zXEofs1V6vphWIrBL367Pc6zDnaVLNRnG52KtjDv6Q1Oufy2FaYM+
vimhrDhDI9aSk2j7ZUnmUJqJlBgCyn12n7ipvKub1HleT2J1odYW7wqedE5keqp1yqrxOVKS83Pc
BPcdqYDO3AmJxKrag1u+YVNriK1kxCXVLf22G/ob9To/f9USMtMOa9n8SFQPSWIQQ1rbqyvlmIZW
bJs4xizgritCU3dO7I/gsWibsOUR2ZYbMsS3GtwzAjfNMR9LsdVYJrcFR0gFhKn5mw+AMWMqC44o
nL/RzsWlVOgS6/EbQHqsO5bfl1pEKUuX5aXhH8tkpNnUTQqgVY0KBvBZQrnF0EFk34pr8YUc2a5V
nnhatPVOIZCUP81GA7XUaOezgt/6eoDRJcLsUSMUgAJ/MlYj9xC9TfRw/pK/xbUOg4sf7pnBRaCl
ESaMo9BbBF1QfAtsStRCmv5cj1Gz6lrPnvBP8fUf3O/lPcGmKVehAwmL+njsz6YrrHudKOEus3YS
MmdbFF0+mE1BypbCeGS/JVH9zkpk3SF2l0jYS1qBS0FAFSMO3BFsGOkXjzStYYQfpiEuS++kbV/N
uOmGT82kyuiKCVErcaEX5P1sC6yVbyUO6mdaouvns9jlVqkX19Taqd2qmwdS8rcc3P4lvTa2XmAf
7Q3lkck7xAXRprvWr8NGGk7ElLV7WhGr3ILaRPz3I2xesC51YC7tBbjd7tmOQWUnFldUdvmD9f5p
sOFJS2+v1ZqrNsizqNDLBrXz1f4BUJGWo3QAsNzNaPRNvOC0GxgWr0ciPd8Bg7DQcgie2T1N2KD1
hi9vMo7qiecT9zrvtUAYPTmqLyM6sp9it9gEdiib/e4O6N+6J8fWHMJ7NzuBjWnGRdAWRUcJZzqA
6xUHQYTsgHvgAcfA8UvKQOPaor1Dv7zK816HbsJjvE5MI7/sHMNVVshtiiVL61JrvI129Z6u2ypR
70cG7ZER1/6WAtlCkGEMJw27O4nRc5J1sRKjah3u4mItkN66OID2fXj7IH1RPmO1lbpzhom/3EWG
IBPH7TF9CqIv0bXH7CqQVFV2WHAkPJAYiVR5K3i2pnllvV2p2rVDnEVzyNCSTA9SW8AqS0gUi/0z
df+afnAvqA0xOhFyLqrzaWAlfX+/irfm281TesSy3WzGTrImbvaoRTsK4Pkuqxl12phfjFujjqmX
VxOxPXsuFDmZfc0OfnMMjljkkUVXUvZePEmdcHdSty5ApVVfYm52QhrnD7T07DI9uT9TMqzhPSRD
I29GPt1DMlUggwUCIzlZ3w6ztjs3sTcXMIF8ur0llL1oQPlernliiMhR6720sLwum3OUpQnscdbt
eM4HzWr8sahnGCcZAud4no+PxoX68RdbTAvZjZoOGKwRi4ByvsVmZTsdpWHR9nf704zJmLjM3Vfl
5/cIpMK9TEJZRQoT/Urw8CspHOHLYc5YwBlQbbH8J3SbxGGZg99CKFDFxo1i6iVtqjpLUVZ+EsOn
7sHwvXda9BpXOnr7RM1bSFMvyR2HpXfCNn7kA3viF9Znv67yfSgrj6OsLUR1KvJMJUuIk6m06dti
AzQIcyXCc4/ESb1ZaKUOfwM+0Yv+v7JJcy12f9oAkHZC6tu6UD8sdxNQB6Xywep5hJDtbkgGUB31
jz445kWPEqJa7kSz8fOPCy6bO7aaKYztsHKmsWzYO0gGPQ8cQcDzLHN2tHfqT+G18gIv3DhvlnKA
Au5ZYOJEI47y8Zd+XlkNKbewD8w6oK5vGu5Cy6gNimcPxCcIilyEeaJVbew5Sprh4IoYNGP+V9Rd
jQyky9Rvr0fb4bJco0WFgZCOxgbQsMUrpc0De96PD3wYOTwMKLxBCRT2PmMLQeuwJ2/dc8BZJY6K
tJ62BnwWMqSRFRp0aZIDhBK3+bADP7FUux2QTtQyOUchK72E9eAN5BV9MT+WWFdk3T9gnY4j36HS
QVDDIm3DeV1ccHzDmX0QusbBRcGrkEuP4g0sJRDOhQTbIw/g4dGaltTVyvaD9uBU+9bEuXr9/hpC
o9EBuNxmB2geB7ZEytbhD6KpPP7jDDOzjGyRW4wT0fApWcZVG1FFkX5RfT6s+IJ9N1dGXZTv/lVq
+kZcY7Qa7Wox4E7Fv8r/ddPDHS5zK4LwABdtfvgbmapFBzOJZ63RmnWde7UeBgx96c0D0J5P2xWI
bcoVqB2W70PkSs3exWwBux9HaCU1h/DJTqHg/oIY4B2Ra3f1xfY+3gYBOf0qwgWiR7PYf5jSc7AV
C0F+omToM87wrNzMR8UwuEiNXkfg0OhWLd7d/K3B2v9u9vSPgw6uuM7hpg1D4KZF24JgTOtDBBqU
w/0tahs6LNZjEws6x3noH3Ivh6ugh1LboLhtIMSOlggU5yUkWQT25XZSuW4aXxGofp8awkhtUupq
CyQeihjwGbs2Sp+V0U/FlCq+IgbZk8n/dCe9b2sP411M1hfYDclqcVaaBhcheS4zqPxzlqy2Igry
0N70n3Thx534URk5P3WxbRJm2frGiLxbQBLMmi1ws9YjNZWzl1LlkIWa5+s3uujN8s18vXunSrIf
qG5NH5/3YkZTNHli6ASy4BPiVsM9du9YlX7Ok6ezK2C5wJqoMv+2EMTzkdSSOkzJ/MJaUvLpUehW
foBXK8d6sHJPiJ5lrfVtu3ar613YyvvGCXEvIkzy0Il1YHv5wvXe1t4mhZdTLS9jWsSAUTDL48ZA
gRbfQU6Q0l1Ukq1Xb3Hekc66GsrjbmzoJ1FctfCa2ETZhOJCj0usNv/RFmVCfE7Twr2Yy4bJhliq
qRUx3faAxTyIoSWYP6wlB99T5G9SrUUVNQH3zjvRWR/d12z/0Lvuf69r6PfhJ2xxgQFFwFD304Gm
GQQvVgh6q93F0mCIZTWBi16q3BFQ+hkpvcCKD/ayBmGmA2QM/9DPeloFj/Y3NdDo/JqFg2ef87ep
GxPMpllru3Y3vHpavsE7q/XPK2xLRE3ZIRC05aAFS3tJ2amZmw0KSVN8KLuppZGMoPsEnvOgzjEX
obK768z/UAOC7U2t1nUNVU12DxaYHk0dT3B2byBLT8mEhHuTghZqYft6+xX/ko/f1JVtAwc3XCzG
J+4l1aPRCm2NJg+K+YihKJonbg64ro9DmDuxSnPF0WKr9gBBwsOW3ih8LKItN4XL1+UvTz55bA5M
UcFYzl1embggijpu0wy66g6mDOzbw+cSw+fM6IW/+PtwSO7vtoGj7m8a875ySL1UaA/yPGPbskE8
iMtTj/hW96deh39aX2UDACyN5m7rEMxfhJTZoiXFO9K4fYBQVSAv2vNRAeWybajkKiRgEVtzTurT
IS7ZMiwL3T2eYOLbTqrWdfhlVJlXtdFDRB/EhNq6Mu9VDhiZKw1MkFRrTcpKVW0JIPdRc7LyoeFY
m2Vi1u0f5HIVVSPOsF8FHIrr/pRoPi/hUsgsf3raDy+nIKgwV6Tvu0xKpAEMwkjx2Br+sW7UXgtx
Z8BCRPfgUnCRPtlOM5OvyDrX4RxYhHs5xBgDCDRxEyyXDTy483A8xnV4VxgG6U9FVOMN06HPk4v+
6XB63ILuwNyIn43wtQwQoPRdC+HuEEktmvkEVpMefLibuJSjfhuLl8Du4X1WhHDDHKsqWleXjaSY
JtTQPEDcm+cbFOOR++5BCg43T6o31H68KDmcEb4oxNe9gU6uoSh8GH1tC2L3K+aOhil+VcI9wsTb
f+lSyVi4OhC4lF4ENWSVRZYxAIntNKbQGKJlnMcsRfHpj2zqPmqG1uruzeJTNZixQ1ZxFr8Gdb1F
zn7npx/r7P1JrsYYY2EEkZhUbSwg5+Pr/ewCrYf1YE8y522Ncyt3omjfyMQHoaPozwMBMuKm7vuq
o8jYmFS5sn9IgfznJn9mJ6MVOcseCktt1QDzJNLBUQ1BLxX0T84y5FGX7zA0ANNb4hBHh056kEZ6
zr2zJYFBbdwfu7yfgwGOI9r/yzY6L1aPCkri4fx10h25LAwhl5p7WB3JqD2qVoXqTpFFB8tnOXId
nrPrandz74W0LVlcE3HiTXNwEaoZhTtlvypLJpWwH4pxDC+ItvzGyeyv2WODK0rOPJ3wPH6CuAtb
0/25s8e3H4a56Jdrk8Rz1+ZxVcnjcd0Jce43q/PXcW0GUSr5Ytactbbgv9tcA7GGJ/djhtlwimfe
GFMvclIaDkIAB/fdOYP98BngnVQfMeCowGjHjv3a5DhYc2djzhMQYMO3fJgkAw9lmpDaM0ND/MnJ
9in+wD7yTZ3BZEHUBXTeGwpGsub6udxqftCUIaEWuxaFrVK4YmGyDey3a4H9xTbohUs1b2In0tIn
oBvuYNjdzNjtJExeySsEuZ7DG7T9+5anEWjfPGreKtgi/xKr59rjkuKbP2VrYWWlPs7hzIy4l+gQ
4/HIKT+IK3daFrM7D+mCs/SRq6JvQjA6w63RTPZeCxkZbxfN9n7eVb8rVc1z3ZE+P17VxSOVZHMV
qbv3A+1Aj8y2DiubLLx/ZCWqIWSvQWZb1OHYVeBEshXJ5i8bA5bx40sDxkEZxhQFK3RlVe8dIyvn
AstZIWzg9jhPpuDmZlRnWaifWj5DQiTt8N2pktWNprscyX0ztiUDWfEBdmgGfXgJA8Ngvd9OBUUL
51988DcCBTjkUfx+ihWlff1BcOIrg9iDM+okjPfw5cCHY/TVqWRdK8MZotoSAf5R01d98XUI7JuM
D6XGCCmGY0+gtXHVtP7s/z5xRT5VGs9coIMCj/4ZPJ2AKYq/pcNG/cVRgURkoqy9y/acakd0LEq9
1XxWwI9GBK0jJmBzwDD06B2Fi/OBWkqGLnl41E1F963vSrzZ9LC8HA/V8YaqhheT+NYdFGYYR5IR
abeQRHxdi5rpJBio5JVeA7OpIvK4P4InUHnULFYyg0zARmr11C68aTQ2OzW55vzTk4Qt/kZh45NL
RaQCaweJvjWGrmRZFwJBpkvV4tud+twTZSLQivdrkJH9Y/TV3G3wRHOTGufkuYq37RLEj3cHhKFF
cPwyV/LJC3RiACZo5A+wGZIhzof0Yq9DiKnUOI3+SgD5NMgW6WgFunfWFiqOpjm2ZzEXjZPKZypt
rnp9kyCh3CKMzZl8ZzJxOYt5AFp7HdtBQFmG1/N0QBbPUZe7CNtJ7MUMaD/FIF5u9PSPjSnTEHJZ
LdF4BUBZ5LZrNhE57iJ1DB1WAzhSNY5dAkgNYBPlyJ4HM6mt0OMeYTNU6FMg/BPlcP26AVaeR+UE
KXg9JEnzdv57KysCYy0QuV1jiXs9Nypd9kLNVZ+JQLsRpbHiaSRPDaDBGfVZIPFWlrVzZ4qrTKqi
PXTZ98kQXKoi4ENnpFZGtz/pOzsyx9AVKyfZWpOrdNYacqr/KzrNyXF7KCc75mvwrk85clBXCZu8
lM+Js1O1odN9vBQqB82Eo8ZIT9F2vn5p2LqWPARLupcGPu29RNsMm0MhFG3lS2hGOwReAi2BDgjJ
uuGiB8Wi3n+TSUyZfoK+oiWO7Lxxm/V+WjixH+DnDKHip0jz77i6pck71hc0gwbg/+TeG5WsCajS
3270b7mGExQWyO4SaJ5kHIjHHIlCd6hh5Af+JaJR5qKLuwwa4nSKpqzgoPqbxkWUzqgNV2eHZcLU
I3nFCqNHpTY3yQ1yeNIkkSB7v6a4WaQYws6t2deFDmi8muisY3N1CUtaT0xEREPGJYNDC4oYGL1N
r4keV+WEKbXVjosJ1VTpKZC/85YFpOIvYNL3+9cFJ7M34DRITlmz9EGF/4NM/t9rxlnvi8vG7Bwn
WSid3jD0U38a/Jahu/YmDDiNcD9/8pc/IU6zWl0tGfUduIp0G4EJQKfZmdm734hxcfMdKls4iRqD
DhQfdkiAdfkMyylLCwaz3kmuLdhxCorjhmHDfx1LZPVBwkdx4VeoX6AK6QiLvEHnqA8r9PaUAj2J
ZyCt9Ds5AmrjXCyyTxxKrlfS1p098PnTeAvjcgZ+ZoeHFfok8DnpKECTPaj8LsiGh0kCl/JaTFns
n42wCeDRarTWPoL1gJK+pyJTPRLFRWkhIlt4n106/ZRkqs2z5dhpe8vQwO7urWncIXnfIQxeS8+I
LFsZbEz9Yf+eOjmVzu4Tbo3UofN5oxa+Sf50VnZoeo42GmJFJvKgXmCmH01dqVio6nDMBHG2P3C9
8HGdlnaYKEuu2T8T6u2ADwgrvCUERPSZbm1vLYTVm8K1uyWjGdZeDfYMBwXt6E4KnczIqkD0yXUL
5vSbYu5xzIReFrsnoToT6kEOukSWtJv2CNa+Smx9FztKvQ/ZkTdq/cNumAMi97qzs8LqnJD5iDLD
TnWNoHsk+GZkQ1S8J3X/4ahXe6qrLXsrMx8m1o95iFM01vkzfyklfgGMSg+XrVAeFHc57wX4LC1x
K9ZnRhQ9FHpVytXbsX9Rjn7vB43p/a98df14/0823z3NkagREMZfDBmKWVhgwnoLFL2WJgRkcK5q
n56u57iNFUqeC9MNxt59Lgt5Vj38JVzCL3F/Oy4igli4VZCcGNs/hlNmJ98ZQLd5j9TVDaFzjyzj
YkVGIxMTSi8NJ06uAsVVzVS7CwbR1YtygAYMC3ixqSkMKdnf4yihS58k7VrqqUmmpmxlUes8ySYW
1x7zClEhlBfNvjaNe6Ou/0ScImIn3NZWeNF59E1cfMhH83uCdEV7Co6SIyixeB/5KC9luS6GGlxM
ZaWmy208oAhvOBptB7Iz9gxL3FxzJIQ1n0KhJ68cBPMiEUCkqjUS5ViM7gQQ7ap8n6XXiv5ghQF2
yf3aUYzjywfl0jh5lnA60MeR3/nzztTfn5wgo+jZ0KDDerw1NAFvevVesGZuxw+Dual9a2vWTLso
TscgJaAQjlYbbm0wlkmjFg9W0qH0NlCzeKn71rttSwgcsO7yiON3B9LgcS884WwcTwu4/SsBcd55
DT9AcVsgbd2xsoajvXpUvKhG065BdZjtvGeCifOpMbopVu3zFb/d/V5WLiC0eYwWP7yVzNa43NeV
WdyVkWHKpp62BAHsruCNQPjRb3xxqfN57CyGNBT2yWov0i6U6KeVaJRPbG4R0yDd7OqmHD2rWzjo
Qtxo3sFN9eyQVClc8Fd+Elq7rsNsb4Nvk0yemPoSqSBapQb2+i01ER49We2lFqYgbIInVJntuaqk
Kz1dQKugDu/BeqXMonEnjJoMd+niEee9oeXz7yKjB2+QIhdTZgYQ8VtVHoQAE/DIOhR/e+lpY363
CFKKjPoKstqTtf84TL2yZ2vsDhuP7Dm8UCh1OSnhmB/6rVVQH0wOPJWwN/smIC7dGwc6jOG2C3LI
0V9/LBF067Fb5vLINCBDJcqYpvDdCVxPXCqRV+mxjtjRRrBdYg67QOdIQUTampw3osdIbijN1MMf
PCHvXcm71rDYFfGo8J7eT1cn/DD7tavqi/Fl3FOKeSRAi20PaJNEW6CrcOKx45cwG6hZqxBz4ajK
spbwrNMa/5a2BJZ/MAB+V4zBgf5XJ21239RfmBNzPkzVrgYm421/+hWph6FrzwNdCtiaTDAPzVcW
F6Y+ti8Pv0lHTaPIFR3l3R9FCuFSVaN6yW4L9O7M3kN5PrBzULng3tUS9YQ5ysXAm/ogOaDTr+Uz
d0zGF9cKTUqr1SjYdlLBzXP5qSzYRavkZvX3+ulUmGC72uQordk/moB5cbKW23yc/vd02h/vn+br
yYTc8cCmWfNAmwhrFTlUKjt65fFfkf44asgYbGq+Zo62kVfCEK8D6s7QRByQMsdJtPpjEkhHSw7Y
6UaJwndFHN3PRKpyxDFveE/XmB8huUyPR5vCkwQgFMAkVUIP0Y3eZCbB1mRYoo2a7a+ViVbOaYwq
6RUkzHLI0z6pyPCS7k1h1sGEH9YhoPkVxfkVWuLRfh6913Oka1PXOI7/u1TBYYMI8ttVGti3zTj4
PPcl+keIvv73PSC93Jqfxc8kginxPIGEB7NEg64+5NwzcQmXvu9pVbVL+MDh1UiNRVHFKl2TQDBF
7qZxUPXKthQx1IEw+pGWP6LEI5k+fwJDKFl2pYhxcJMPM80RINL/6wAuFu9k37WN5NvwEfP/DREs
wi6JNdV6R36KDus4TgWtWY4glHEtKDlFjMPzwdEjDc/eksUIdRc3sKCQ4uzgGRCG6iz+jsfMbVmv
qzicAU+18fRVcqoruKzWxoot7rWFvCj4bbqRIyekMZGsldD39JXOtnfiHCxnNKq1Ct/zFVb1qEM6
ROt12u0+AHgqzWrKI357J+3/I3rkt7sj7s0UobKji+GJIItjJlluUYfANvqb/+VoNUmdL8cuegxx
1zyysBfqkOI/os8ujcSvvHge1JN6Tw4WPfEgjGjQVnpTGdLA7UsZkv8oZyQj8ayA10QSZYXAOqLb
QarNYVI/eZf8pAUHhkG8Hqsg/lQdEDLUu2D7RKOf212e9bWDNxU47BurJnz8jBIuz7IEUltggXWL
kTUwIpd16V8Cuq5Q3FT7kegox92X5GgZf7z6O1nA/72lWfC/8pgZeEy6byoYBvPwu+DVF+a+FtHq
OE83Za0dd21WxK+Zop65cURlpZOCMXKclIidlAIqFRnDtUy/PCRXFEztb47hSeZZTHouQS82Kwm/
YvdVEHlAyyklxKogWah16bO0fSno6fEIopJdU6jRHbRkNDNAoVy5lOxJvmP8J7s721oW3yFwHXA5
ijkcL/t/QhWxab6aDlqzOnokCVZXjtrvjHhjwiEoj/GuHmVnjVsml7Ph6svXaAk+/ZQNrQyAGW0W
qh7RwnYyjr7/SuV70eZ+dj989RaY1aJGWeFOhgTW/QR2+rABJmxP10/Q1ZNpUjq4iAx8tiZ4xdLp
Jh5He3JjanH3UlIMU7AMc+y2AUnZ+nXOYRgMw/dkWWKV2Lt43PMJ/CWfCr6OQh+Da8t+MYOgqyTf
rB1/jjsfF7Eo/3F9euPd7O4ZVov9mr1urwACgZ89syXPMbYWG2T0ErIbZir/csVEEkwYvQNR82eN
caHVIehzzT9ECi13leWnPwZMSPONyWEUNmyGCfXKQS0g2GxJI5w9Pxv19JmJQb7dFx5L32MSpQGj
7Xg4MAfe/w9wds8XbZx+xgoGRHp4KE+Zf4HSeXlOnZwP7hqJiBm+LjccHD6+G/zBRwhfhLVWVUzN
OSRtqlPJ2zOVuhIaIXWVwLLbbOwVJI8on9wHTVgjWaOUj2L83WEYfcD5X9TD0jw++MKBK1vnrOt2
XvoMY5r40bKomcofSEHC9NM4AFzPlAk9DwA04verYY9Fkc5VR9dVjP88n1WXOhpb/cPLVgatVqFc
/hUhHBRoiuTQx7CstsAtK5DytwIfZGxEEYDPVLu6OFxV7hsvxOTDE8XnbwqZc7WuOZqyVR8MorBp
aMmD0diihexil04SQwfq1BbUSXfwW20TMggUH/2aeXCVpJi/pRIPOrbt5BllIzy1XZnxj3jBGbPQ
JPZ4TZlz0EJv09oi6lHespPH4+CgbAVCMSkGQz4EIMTUJR/eXSGuEWyCu69/w7unoLhuwEl5Fsmt
Ug0pAQncwWr7ic6knuRui1WDmKKMGQ6aWPS4unuknI0xlA4LzZ52k+f4+Vzu3y65cFsJV2aAfSaD
gRWld+0kTxsoURpBD9OIRw0Tjy4BYkDE8JLNB1V8eGqF1bRH8fkRA27s1M8g0WY2IP+QggpH5GSk
oEdBqmpDC7OOz9psl4/KNUruAUATO+oqVNXhiIl1KFDeaFWNrqpijtA2MXs1ABR79jNFPgMKIcYr
CycBWfWWdsRocTBkROImmMnX8m5eqWsRYViulNRjtXQc72rKY6iDGG79AZyM8HtxFN3NbBJ4Cqcr
jOdO+ykN16GAS0SNZKiaAtQTegyzmmsSxTTQ1efe2rlHsYyEB20fBRExBWw1jnJ/jXgqGbxJAJtW
qmrRo5Ve3kTHA6JC4P2kt4gwYogs4J0yj6tZphPvO5nXKr5cpqydTaNxSUnT8MEi/pO0c2Va1S2Q
e/AOGHk9zVbS9GzvaO8WcjBOUIx/5km3uqB7fMOSzeMLYMGHPAcuW4m0dzW2Zo1baaGhXuYEZLVL
pe7utPhcWU3Qu7XvMXts8bz5bQS7tljdKDbhFYFRBfvPkQeuyJVHDRfcb0mlHNzLxjo2Syjz/N40
xHhQNBkBkFASnCY7BQOr27v55hpafIN8/5cqRoOXHqksO13/SYQVnx4E0PwcCL7/BbtCURILwDzK
LLep20ArH0qljRxQwFGDDF+0Ae2yAsm5wkyHu0hcGhx99/r9o6jKi+KHiETBuov9drDEVhHc3sqS
KNY6B0QsHG63Dx5iQlU5+qPuMsw6f0cwjUkPP2B7gFAJlT3wLGyrpQzdvnCSE1u3cSBz1/8U+8kd
6RXGBWIucJusXITPaHebY1ZYYk0TMblh9eXTNF/dXs+wwqDBJ5HlqzaQ4UcTp7eZK3hxI/vrAnQi
jYxowcgAvIjUo2BrBCvQMCrUGOOGm51wAOTt1O4v2CgRGFNCGrjCoWDrnCnA1tA2pwHj2eimwo47
XereD86aenSvOlbQOGt8mk/MuqTZ1j4EMJ86pqKmBx+K4gkFNPmd4JZ5qCD44cC4hhdySVXWlmrq
dvfPs/eXk6b+id11cdsjYhU/OEDpL+coMW8oAQI+aHurMR5yOFW1FgZWSCBKIrOJng5/WPQdeTE2
C5CV71mEONUu3iUPEERUZCmBHtHpMjdcflbpjRmjNUuDdIMxDnBgTxTVUO225lXC2/fNslqKOEVA
TOMWRdrE1ORDOm+wScdUd4UpxzSTyB4DR6rpue8/7bI6xoPu9FuDX+QOPFPz2GF7g40GHpDU8+z1
eNWbaY5amy6W5ol+5diJ+Phf1NshhJuuCqdFZOv0Ux8/6s2t7Ni7Cw8e0MkCKvvbZEYc6YsGwWVw
koidSyB9XFqcw+Gv1t2CAXvr7OXVXnfryewBqSS8SplAMRT9AX9lrZOarCcEOGamn7YbCJSDeUTU
lzlZkRNgHIpGxcLiS9jxhljIdNTs/ttiJwjQW7ESrb5dM5uqPOtZb/Vz+Sca/80v5LAEIFQT0zTG
QHDk4BccKYaWQs7ZTqA2JysF45vySOeFpRBFjU3kEj8IGKBguFH4o9MHVmHLTvqH12aPaD5CoS+E
G8NBXnpKUiyit2EPkiFPUPHsk8CNnWyXCu2lgxfn4IFJIi9gMTi1ZJCq5wQWzt+VXfzlnPDtpVP1
oyyxoGblrVVN9AeV4aRPgpcS+gk6qO0ShNhmGf3T+LCuZsh2q6jwRbcX7rW3gGQKj3l9onAlp+rS
z5pOhNQSq0xqPgwvyVa9o5fK5bAo455ts4DuHLKJSslxBZpWX7xQ4N9FbelVLvwPHB0FGuMbzHxe
7rLEnlHHv9Eo2rS8ka4tGshVCPZfjV8r6RdSp0YLAL/IjAuwkz026ApdmM8NJPB4vr1N7xFQeXIo
x0FELhrBDNSWT0xAItAFzDKsgN/n+gcu9pswTmuWWGXSt/rg5d42Z2Bfr9AH+v1AClEAEyTuCfdA
7fHeWXItZ9slbLC2jqfZ0eFPrICUjLVGeGuVtp0EMggXpPLVf8CBk5FxY4WQUOdDFe+g61cyKJ9D
rV8XPS+L82OvO94TVwMiEC1es3DU4IyH7fQBCMqMbImFEBv/lClnQ08f14mDrxU0Ah6gacvmK+IK
V26Qm7839+tP73q5VmxUTDb0eAq2DDDTPuvfXBW0+NL0WjOIeNdSRxluupo8xxOoP8ot9hjBS7ps
7t5Quf6tp12TxkII8ikUoTXpUmj5XEOHbNbTxAlVMj6zDro+EPquOT927PdMMfvjxN8zBVa5/rTE
50n3TPj4dQFFDoTEU6doUUwM8IsoPS7sGGCfRRXhJwC64RIN/SOe2E+mXJu0XVL9JudcfnZ64jor
k3S1/pErTi2lWSC4j+NjTqGj2qSmN5wGIADUpbos/0YOpTaxHY4Nc20scxVrbc6bWXanq1cWIDV6
0kblo3hAbd7Bua8LQSAc52wQvqJOQ0lAeybFmCiweeKAy/K+uuxSu9m/x6xxL1dbtTI8Ugz4q3/4
DCIawXEdZTKsllM7YQQes9ndx2beStp6+pdAOnRsXhjw17B8gf6ImNt1WjiwvITJOiTV2SWGgJJk
H6JINjlzBXERX6BbwuiEiTjiBzJycvF8jUVqFUj2PdSEK7Gcb0L8vc4AD7q+VNhDPrPcbIKGUZL2
Yu81LjKfLatRLUVn5f75X9FBkD1ADgYRi+PhU+WNGLsfhGDx7sdQ50JKhY/Yl+bLPntvgxW7cK5P
V/yaB7P1tG2ENSHBo5eNa9ZKK2Omda1S3wJ3pTodbG4uPUR1+59BtA1JlJcfyIHyqOmqNH3GlM3w
XxahU3bUvp/EVvXxjcrLzH2RrBN0pu2p/VowNtNMoDcdZUmE/oKyb8csfErKND6yZIDeYqZZU0s7
xIuqJvf45pxb+X6RoMCcnaHe/8rHxM0EGkjEPRFxJFWXkwcialsWxKIf7YBKJdT8xNNOvCj/K7ne
0W0UEKpVAV9GP43RqE7tt32TbU3ZzHrye/OtLMLiSNBTHYh7S6bdm0QpE+241PbgKV6lzVNas/Gb
1HXPnIrEjyfGyX/1QNB2kuNKeCEHVMhwyONxGTYEAurMt0dSW28EzZjJpqhdLTB8cM+HwyMCdUdO
Xe00y6o4pz/FcqEuQfBjaWKMfwBZIx4GN+mUY18jBtgE/BOZfWn7iLreRAk7PDkWLVQjR1Akoa9j
E+V8Fe9aTl5Y2N5S+pWPS4MkJG5T89D+9FiijaI6ycUxgjC4OuSjn+1SSTbNOqDPtM7TkCAcdHBf
l/WTrFz/84HKFpYwLty00qy2G5J7tjKca0K0PzPJGUGN94Zrs+MFqcQtGXxsPlC/cssH+VbblFSI
EAiuqyfmhJFvy7gnyTUG4mjOsFN3XRohsD7tchFa04r4Iye+kYNL+oWjd6l5dpAqHGRFQD5n1JOD
hrhU+TeWznZeONZO331f4KLz++87ExPUJ2W0bUBe7S1FcjyFSwFH734z/CMUbP72pQa7Mxa+JoSX
l3GeKk3ju+H+zphGuf6Jvj5OKoxfEpWIc7BbpQf/Dw0z8hynFXaIL2pfRKO5kgRtvnKjkNQqhQ0z
boQONYQ55d8E3dVpbsKp7lzM9N0HMKZEh159i8z29ib9QFuc/gkbMTyqVS0H+Ki21Pp0CUlhBCda
eqGEbw//r77kIAMxy8vM5u7OdewKR/ONBaMfQx2zyMhnzXV19QgynL6/XLoxPG2+TTW2XrTFY+zo
+cAXbhuMfLWN4Y7PkBG8Kf+ZNAGNmHAZMPgGwTkK0QDJQUWo4eiznBmd6RzEkT/SVTac+aiiAh3k
eHGw0VAeMMsrqLcO7KQmGV4edt9rDHE/84vTvplJhXDLdXiZLvxlVwmf8alVyckMnbcGQFHjEliy
CR2ttiHXvZN5ONGlhFohSk8uR8TfsBafvOhgBwN+DPfDTgi7XyAx0O7JiZbzDGdKmspmcqICrJ5+
QTwhWPuHEJs0zw2OcZI7H0qsn/nNieDjaVYc6fNrXPD9/h6SNG+Uqn/okecwNrUwQOZe+90ou90P
B5xY/H8r6ibpOd4VyITh4eq9fYFx/ZFLCGIxohTAlzBNlSnKG/vt4XDtVKW+QZfxY5zPm4SQAXvN
T2R8k/QdmT+32YDZzDi4lheGbMcNCVjRZRneYcvIVg59xjWRLmq6s5AeKYsv0MqKLYcbpRz7qARs
MjsVNe4OKd8oxYNJ3WRbZxN9x1btLKoHkZdYJQO6QDMY+ER2Uar7M4+Asehb0xF1HgPGHPgqz/LG
Zbv0k7n5bq+PGmrZXdxAzz+VGRME6h7I27RdRmBXgoGo+ks+RXzu7xrkliCbQWo2kASkiBBPi5Tg
lmJaIZnnUszS2eAd/kg08awUH49lo1RpvtU4u7OZW0r/86xe8QyhhNe0yg8w3SDBGQ0L5IEJzULK
T9SyZBtfm6myI00Z9vPaGVUaaKYmRMpdUye0yZRl1CGBEG7l7lluXBO4ESircAKLCAfgicIQ7l82
WuiCGH2rLaQGYcgYjG1NtWnhZfjcx2fzdBKwoo+vHZQH1yX8ZnXZBsCSkMiG8k8fpEvOT86AgKz9
jtc8soJ15aa6ya73aE9DXplTGFknN7D07tU0jrLn1ra8UH6n8LUKCMlKSY/lt5yN+go+k1Tb8Oq2
fm20J7J+FJJ/I49+h2BWbhag8wvgk1Yh/Cgyf9xDh3DYP83FZE2OYRAF5XtcfWGeFIlo4rKIsrBg
2HqkD3BFvW+uUgRA3vb8eLg3pFieSHZJqJrlTnSfLzTu+HlvacjrWyDKCi1q1jj6KrS76Dkaq1HW
5ovGacaCHP0i+DGpJTJQwMYpWCU0wVrZ/5juzdGdAEqSjA1+5kBNeJt9Jz/QeLEDAvjIgXSLP05b
4Bdl7+TyuxRW7hAW5LEAWvyk1RAzndqvh50og45+Gd3qVfEUflWhRCbnOcM3wQP3mCyWql4oSpFk
Ax/Y/25NSwIY8/jAWyzs4a9lFk9vfMOTIqvuTucjXiUlneG6GeWrBsxEIuGTtrlbd5571OatnuF+
mYKclUvHrr9Kb5zHkQqfXse1BZNzcu5QGNxn57OeoxOBb8gXZTJnjHxcujk+394gGrl/PrCp+/ND
XnS3aLmGWJD9ocBKa/RTVRBIm5jnXpLitYwcSEn71bMw0kSjeiBprvOsgIwOkU/a8UvAyGoDSNSe
T+Qt9WyTYuzcuh0H+Vwn0avRkFFmumW0C7ov6sNoqvPyluiWeDp/4JvXCgFuizUnYoatVbITAS1y
GEzd8XBvk60ouZZ5ofGDKkEEywUsyPkEUeAGQDMq+LinZA6BGu5LZxHVADcwCUH1MaGkAYV+uS4l
LRefJ6CEvSMZnMgMS8QwnE0vdH0zeIx6cAVm7BomAHHSrC4SkCrT30bZrUkEJln0aq8aissCM7+I
aa8A0xqM2qTWNAEIn152EGS3qkZMJcPDheSXaC48kKfptgDU2G54PJaDoFN8RJRh812Ocm6hp+iG
0pgMBNuLcSK+GT58qtxi6FaVeOc7yC2JBIlbyL/qQrXU5L1zEdxzEmLeJiIsyF0c5rEsJQv2PbHA
qah+ArqluEg5kxSnEVTho1uR4fCQY+Ka5I3+i93BAu0LhuF8PO8BntSz/XzzS4/vGv1kxxML0K+0
42BA+hqOYuABbLMF/9D9OrIOy148k615KSPTurtdnlCxmA0etZavebhUVKzNcSnVo7p0HZods+2r
ZPtZklpaU873DLEjnPcLOWhm5efUn7nA0iIuTUycRSY09PcTLvHP1sj1U8Lq+dZwcfD6rQplUeLz
3XzqXbdwKaUD3dptZc63JMnb04SMxCt9Jc9pikVfdLZPCQSPVMWfl1EJK0C62llNv3Ujsytccs9x
YcsBFTcMPaHuZyV5bwJwf50UPXG8f3fOh+TaVWETsoEZccAc1mY6gDJ3XHw3kC2/ML9cHYnpJOp2
Rt1bW1J0yHZcV0Dd6D5zs0yR7qDejYvc2tnXt5aIYqCugV2eCVx0owZTl310mY/cSrRUZXDsDS7A
CFbHAbS0reOyiIiP+WXNKx3yTIt8Fq+s8BKs8qI8hC6hv5lOv5Bn5hpRWazhb47ND4Z0w4p020GL
LLyyTZnsu8GVsCx2IUNGNsOPried7gNxWZUAkolvUPQCZee9GweSTjMO/Gj+DmetryMw2qisKn3n
cGu/GrXVBbo+yPoFh/fjz2WGewAcrYK4iEXnVLgw7JqK3CnDxpwRWvzgsc9oQGDY0uqzomUn65HN
uQJZLgMKAnmhXrdH+iTlzL0zDIHq4KnCf1qRr6a7P7pgx/kQa+PBtGk6Ykfz8gqYPmjVRkRwiHQ9
GjI46CUVBygfh74b3kJEs1lIF7KYlbPFaWyxoFxdA4WF8bsw0c+vALT9bYflgKPj/GAJ77gCOVv6
tN6w1szh2YxxYgMJ8X1RHj1WcJE2mzFm3U4siZNkOIxMC0C8uRuMEoPWI2EhV4Yt91jIQKBKopFG
u7yClt8ZCqoivcfdbcuW4Nrh5V1v7siBq7elAiziQ9KnxHXD+EmHiFWDAT0sSVYRmMDBgd+1+LYl
vuBWnlCJoXE+obVMD/U4H2y0FGZJB+BbJ3TEx3V+reNjj3KBiagdC2+AZbR6Z/u51ufczWOdpVH2
njQ49jmp+95vFw7gKzSue0UN3vHHxMnfRwmrj8ZqXmKBsv9SdamQ566KlTgsl390NpRw5uIwiq3C
f73xKD5iHbeLT2QhdTWVaPM2NojwHfC+fxG2JlWfYM8QpoS7lSIjwLyOCCILKH8YUUrOgAZ2DT72
1hPQc/BeETEBKAMOgNoOZWY1ZDyseUJYsQvzWuU6TPBnASvop7+lLUhRd7qT2mQ+aME7D01xEBWN
BTvODV9WS9puP1IDette/xCr3sb1Ca9tTPqEElWkgZ/kI8kj/6YqIH7NF6oyhnel2Zle/8DAS3z9
kARVJUKyRL2tY32HnGZ6i8Di/jGVeMP7BU7rWWdvF+4w9lPcU6+RNd8E9LFih6kk58uL1CPJxV1N
CUvUyLPDBVOa5B7VNJBgZ/p1aka7TZpUipgLPQIrTynXAAQGkwP0xoiApYSDV6HpRUN5c5anpuxN
pnXQxm61sIdMK/OXfKtfaVaqYZ5LOf/1j7YTmqYOJn6V6J6YlumuOtdy0Or9hToda6HWB0yY8zLp
4F7g3PD6buwuaH8HSwWTQpO9vyM4OJLm5VTPq5Wf94MGiz1jWpYdCONzCsnPf0hRn5e9Cpo85mJN
hAFWoCtKGNv3r2zfl2D/emSybBxLMx+fGF1aXJtlrDDvE3gB+oYzy1dASNxSlr0eXFkfo1RaywDW
zhhs/X3Bj+9Hd+qJc/+ZqsnRxGjexsU1kWhJWhtg0w/vuT8TfgV7w9nGSqxKQpizHwoNYMfF3gAz
p8EeVejF6zlFOgFafHjeHWjcEelayygQDtCJv0et/Vksl9SFJjzc0HT4BZfKLiMRqSyJ9sDz2xWL
PXRe4Nv/RZXN4SjRtjAeBYejy85cPYDLVtCoduNaGbYAZ2b7ngad+SnQcCvKEwEdciEqJ34tsv2o
VDNUG56/d3EOpxWOkBqcwlOR5+a+6xu18xr9UTBslJkhKsUYQMwHMgupCrqRSbfZvrYORztLK06Q
+GxJoQj41r9hzzsv05kGYvvMjhAr8n+YQt6bGPprhgEja6TRwHgGDUpavV5g/Trjj6Oq3/DdsPcI
ykkBpGjBxWaRatQlqrdKwOVA0LAQRKvJlQFykO3oe4RyGQyTdIeafW/QmZHRagieIGnDEWIzcWDB
YwExbtORxMi5Te/MkCz5+kPBgzET+SSAyr0kwh6W2buhqwZ2/eSUxkT7/ANFHiAEJY2n9gIK/sML
XQZNpxHxmwhVq3pw+GsNN8vymSq6qmTkv3jnI4HWWrZDgVfFZuoQYwNtRneEq6UA/b3Le3F4BlJa
NnGktpjILnABYAOMkguLaWneF1vn2Hb5QVh6rmRmYPeqZoYDw5sJNs7nSjfirIIIP76+U+tvx9ir
lJf5EF6tDxouHA2pVg3ShYD0JJOfN7mVtVNQGjzTsVjyC5SM1IXqjHuSaMeV9ZdP6nHBPGiVWaCn
LsH+nKEumDZviZrhUHQ0Gl16rIV9wTvA+BJZwSgfE7nq5l/XlH5Qeu0l2w0DRtVGa4zulA7go0u6
BEb71vEKtQE3QpdOVOFSQsPOA0+F2fW2C7E/JZIbu/3SoFYGJzba6/RMY3RiJyUJfqIhkWp0BtaK
juhbnQVCiOYjSo6OXzl/qtSYNl2ue6LBSzL79SuYSwh0QzjVYo/Qzz8JBnBVAPGiRqGra9UQd2mY
ndL5sYRfOiv/zH4d5yR2WD6madPFd42pJZN3RKMslTU6wgmhf56tkg8V9tX3AP6lLJfribYugmfB
gkdyR2aEFurtpn39yID8FRqbVyqtG77SNIgw9ONiH95U5oqShT6t6L5KJ4pjAXinNvkCSafZIEHL
RE29h7IOkv+TtO/IyYA3yGeAHKIQnN8V340d6LufTN9SR69LQolMl0tCGHkhEhL6X6Mhg3N9h1Xf
Ox6fTlGpMm5jYYxGGtyUNnqTozs+BFT7UhPIIdV3a19/Kyi9RlNJNrzA96NxxXA38p+P+NrhpeSS
UiTHO6lY2+jdoEX/UZuXp3zZ3IauBP5ONJf21oBJPhxucAIQO28icy3EMfNCnRKlbzyTMqUolQi+
xTM0URB8MFEWCA9sQ2gx86eN3kXZZ0cnKK8UQeTzjAPD6TrpDCmCIRKTDyE8kk13V8jzkz40KdJj
ZCdRCwidNfpWmAxrgP9NnK7ZxFxMVAKLMKSXhHcDntulHJtwKkxi8m+WCUM9lEi5h5U5EyFeJXuE
rRD/7clNPr33V61ckwfgJx4pW6tFe0wjeTUgtk0lbYsdoZGebfAtWLLHeCY66CGE0b2OYfv9xT9K
pNWaYn/A5q9bQ6I1G0mboIR7AyMvsIDbNT+6X+kQudyhNjmwUNqDzNzTd19jZ55rs1DTO8YP4ZIH
mZXaF9z/krNLy4/kPnf7GGsrms8fkuBVMhCcU1QdF3Thcm0sZ6ltcX6km0DbIZG0pyXPB0TWhucB
LUxNUFoi/1So4IKgmBT8h1GpuMQdSFNiufhGvCG8QLorJprvB4qRq2m0IqdPRfAfCpPg07bnaCEg
i1XBCZHCJ3Hk+fSSosCCYTuodnO5O8gLnYwd4I2nCfGwIr4HCx5MLLqoUpWcIvOv1US+qJpXz9BA
L8amhiga5YvgOcfASv9eiP1Z2tDctAP42gRI+cUWa7ca2sCU3qvub78S6r6rFn2y0YeXrQWVP/yD
ck7MLGWMg91HQRJtiycP4qkazlWkiPjY1ptMIkhWWuD4YzmCvcM2GTpj7yDQ5l8uj7PyEnlwvsW0
lqIDlaiOjWP5xZjoVkzlxV1W9RX/E09xFAUixIsrs4L6tGGOSAXvXrQrWF5jKSYDRB4RHT/2dbzJ
VzaovFhkAmPUUKR0APfQ1Va/hi1IB0CI2CoPIg+XdeVvz9VHLj9PEYZ9l9q9m25D3u9Rb6fYTH1W
7WIiS7yk2mdh6+1hebvqdBDeN21Iumk+Z0r2eyywE4k1D1DS8XhkJM2KtmYVu6R7cMckTFMqNJYr
EVx4XSDUbG7Sd3tkF/YzRPEQAFdFPh98Sd1IkD/tk2xuOnVybnPhYgtVOHlkN408ROwV8/vF3wuC
jus7wFQHJOPGMggW/kUZO+UjHGdUXodhpMa1TxG9V0WXljHMwvvNAqUo1wXMgMYSWdu4UtTvhDq4
U4EGrrqFioEvZgJ3n4aeqeoF39EDHz12A8Qs7a4aFamqfFve3L/1hmfm/UA+CDtPx9/UIpoy3bQv
pYnCAfPDUMmMHlySj2qS5xghp2YnK/+1zQ1r5YYG+c7hrM09oh8yxjF15k3pqWy5oXKuIqdUZbSz
lgjSQnHl3IKtPqK6FRk64O+YKe37cDh3VxrmhPacuUZKcsuJYZ6Av2JCj8PbEa8AcgIH0L8Ob9sT
Q5k1X+0rU9IXbV/+98QEmH09uNe+tZuEIwn1wCE9l9S9BwHS1mzXiQpgkJ+BWPEF39a/PeuU3/Ho
/bMpnZd/DQCbz2nqqb87C2Vrhj0gjIYAokMW/Y64RcOZU+rdv017vKSkwxX1pmTwpHRnGi95Sa8n
JBJTS8YaVhe0zHaCN1aO7NYPGVQX/P8jM1iguWluFMsJYBlM7//9Wzrr/cu6La/M8bhGufYSrJ20
qgssv/nE/6YMqMU7GsnqObbRhinIwVL9ojW861UkWuWPQcxKlZfjD6UH94UQOeQb7qHsRYajYlyo
eNQZgIeINucn/kvTBieI9tmwI2tMsktLH+tiP2aiKihOh2L0g2THtzPdd4wLsKsPnHF8scDwTNtW
qhSOSLmHyfJZ423tPWcOLdBNA6vNDer5KEeB2pmBVGV6bwy0UmJ4LthyEY3xWHSjMyUMDOAN5lBC
s7NWb5yczjfBlj7uS34AUrGvOIYmOyvWi72PPw1uJtfkhE7zhL6jROfuFLEy+L5CDvM47LPsNzZR
NhpzgOFf3J7YLj0wwm2FEnKzKmZNuhza/u2kPF8C98xNlGI5YmaNJEGeItgJXEFWRNiWSrFDSzBr
Uo9PltDTww2CSGXNVDjD/kFC15x625xs3g4XlKXXwMP1tgHy0eFIrM9nJDSr03F5Tr8HoZwbVcUZ
FuMgnW+/GtP9IN3P+//hro1rHf7DE4uCTHAz7llNHkV9nrFS9LGe0MGf0aq1a8hCucuPpX79vHtw
f/pff+kPLAJzmyo2aK+6zhQu4h3cxHyYfELeJsOIOe4+OCl7XJ0NGWuLNvRUswQbpuKbBRWNueAc
edMQmeNMdUROzs9Dh/Lpjw29h0KIG2sPlcsSS7ijidzKQwSjYuRIMxU+5Zbjzk5B6Obtiju7A01c
VeucuxmRtbTex8ChhHaxAnaW9nsxHiwuK/3pgev1rskd7Q/nDT6MvCOV17R+vPWjSHSvLw44Oo/0
mzno4C6ISR+MXGnlaU54ySIZdda5qfg5Z4U2+5XESxup9bHc6eV+6FXj7tkNT9Gpvh8ggeHmW9be
cXbeFar9VW3RW5m59/SqRW56yS3xEd/0Di8i5A9UQjg+tgyZxRvTVygZM4omBGmWz3+nMEb9o9HZ
034YJkKpFXY8K42FNP1grzeHt27zTZiMajLhuRqJL1iMiUhtAuUGi1lfJkMIBh9FhHzMswJ3iJZ9
JTNy8BN7ek5lw3NuCvSL+0CxvalgceWW6HeaZDUWnad9NuCh9dX08tZVvb7aHffCHM3NBHHWtGVB
1CFW70JmRpjdn9NS7OOhRhTwrHAlU7upESe4G9KmKMc0sM466GLgTKAuSpTjFrVEg+ZVqqulvft2
02M0sr6466vriQ7rSkx4IvjnRBrhro0uZCC+41gZtdRPdoZJ7YM1hp3rU0CZxerVrI1guGFOcwsw
1DsLJzcd9e/TeZgA9G0wdExe6tf1I5G4UurMtakQ7g9mUispMo6me1k15Hkf938L/R79qX8Oqh1b
K4GX2bzLrojX/gYXTNXoSjpXFi0BA9dpyHzf/MM3yAlkp98g+uwC/Bd5hDgsf34AWFlm24XJZN8H
J9C3w+apIJGQoR+j5IljmRjuU3WEGIV8zw15dxVZUEz4e2fH5Key+7kNSQeIHA+1l3yDLhazjq5Q
qKsGoJIxPyiiqKbEgzfMpbdDByG0hW0hJHG6hPGlwQAQoCQ/qczDVMdXUcvYjZw4TXHrHxkJMmAZ
tZ0IyyJADSZewmeKDkc2Ujk5ltGlUes9a9gf6D1hhxD8hzf9DP0ThB2rYEwd7qJmveappKWtNbaN
cajm+aMuJ9pUEAYdntz4yuqc3RPA27Xv2UqFm9/F6I56GHb89TXsB/Uu3GyqyVm0vQGPxZ7CZpJP
fZ3Q1w8H1rdHma+hd1cNJif310g7uxj5sjZYsgY6yk8JCj9jzSQQVHSSYPZiLyg7MM/orL6nCm+s
YE0qnzWyMQrBtne8NGwBAKghcWgLgpxzTcYBJoYI8N8pjjZ5Xyt98JRNGHedfv3dSvFCa0hWTzOW
d+qZ1euBQqi6zvU5cjxbl9b7/TLiqXX0FbrI9Lb4oku6VCyF90qnw7JQsumaOfAsMYF0055yXM/T
6m9FyHkt7Rn2dhmT61iYtdd10t6sPsqB9hLg9mEKdjlp+P6peD7z1faGVkrCy+uL3vQugXx78Cwm
kScfWm87T+cjfXrv9PPQkMLaToav3fs2O7vVSHqYFG38gyPDXeNr2ZKNo7X+jEVa9ymHk9o6xnMu
WPyvDw389KftLPWZWhoOoMN29UtXhrAnDuWlgTkwzGSz1UGd3D9DNDk4qXhQUe8V77fnhfp2zvNa
5/gMT+hQRkkE3KpjLLFbAI0Ca7njXzkUty713Dh+HvaDeiYouQ5V24R9tjlErtL8C+TbG+eJ6AeT
xWGbZSFWHBaMPZ8m44wdeQFUn6HU9wGonEPJ8AnK58U/fyC/7XiOe17CvZ5PcIek6vmzDejHK1v5
v2rbiCM2uBMBRy/NiM5O4kzGdckBntyozm48T8aJPGCUWppE663jjhsvFEk9THy52IJYgXF+ctaV
++OgXoZfWXMiCYXHoSU56wEOEkltB1wKjxAHHIWiq6Dwq3nFfakvtIbx1/3S0Oa+MqVTi5Ulu3R3
F/RB4O0vvpR+r3cOgr18zOG5pADdTcedlfhfg9OJXZXgujXJW8oGuBRlukNjdWPKCC4URx93yYjG
LfNPHwOey4pKljCXkWsqQ0catArFVgTm911RNtTv3K9MloC2jEvR5l0QwhbHqM2DTlxv2mbsmDI0
QHnUFlGZXgSHj0oS5bIOtSi9HtqoPSfiirQ2d31vo8QyveYYzAQebLiOcbr88lzVbAE6hGy0QVax
FaCo2VYH8FYkAm3wGgola05Piwy9ZnV7jrsTDFmJnvUV1EKQJmpJqxVe8r/yd1t3yhZw62YxzoHg
IGyJl22zR2bdlbfoNRapcDNGibsU50JyuSvK+Ww2NGNvbXVhSoNk7rtgGn/UNKxfK8Dl/H8Yak2k
AMtDgKFDwBvbQJFD130+hRa6D3TcBBvwS3I+fNtSVYomxMdo08w8uwYpDkeQz5ulAa1fsMuaIj8h
J5w6qyYwRSVe644lP/M2m/J3kM/vV2pdLS5xeFSR3YhYr+PhhnXB6cou2iDVnWPSbblRGBxZpz3C
vnDE8vMmv2aNftnpOIYGunzhPIeORsov4kpTpbdCYaskzqz0PLYgN/8A3TH1Rsu1o5S06iabnpCj
3DwtmfpIVMX+E7osIOTEjAJ17aKPrcSrukgiLFh0P37L+SHFMcnw8a41aANEpbUcUKVh6IoQ/aDe
C5oUUrozuosVe32B649hDfTN7YG/nqktJokuxigi1LhJqQf+DKWHV7pYMh4bd5CfihcW5iBqsTCH
qAVQB/Y8m7QabEu36tqHPNZmzWInJ3rOqTnJdLqCfYGys5GhE0CsxTMYAzE58pXhy6QdEM705GGz
exkn2hp615sUvRZHEAgF52lV2dd52w0BTSdJqrelrPwMdirul8HMFTC7H8gXw4tKwbNwZtkgcoVy
uRwytBOikfC8gVhIrrQjmM2BEttWHvG1PKc2gqRXHns6zohaCStwwTZj7v5Z/tW57Dn5UjL/zp+D
rB5B8Rm0JyMuL8UCASVPwTyEJRI/jHSX1/FuqZPU7RS+sBDVSJuwRrjHHsrZ6ZHdiG0RSUiLDIsR
NDQLT+7H6GMhPtvlgu/+ZBQG7yL5+8r8ogdT00cRVAdd8DHTRP5qDodLU6cx+cXwcr6PwvJGcOQo
pgj92o2oC2DUUW7a7Pw8NYL3Mh4r2F5KdSk/mkbU2Qkrq7UMpeIYK3qv0MlNVox2RXXmLGorGrKY
NQYCyXoNYvxtEgNGpEWexS/42pKyx6t9/zgxaNscxShnJCR2l531ZAnw8JzDqMfresCl2nT5KHDD
NIBzLDkEhVd5bwflt1+fEMGhMUxNUJR35LuY+Rf00wZnQ04prZ7L8IBEnuBodUSdRSUPl8qOzdvv
WufCEDGo3ySDnypVStnqyZzJp2GKBsuj0NP9JBSTXPZ/bHzttRyEQQYFSt9xZhys/yd3ZHSEGeIq
HCfH1exdVAkMcORSO/UzMP2SZjdgBMaiwmKpfA0SW5iMdupRUZ7aEEmy3CjGIMPnaa3yfVHD8ro+
GgIx7n2ba0CqiQ7mha8PK8GqUZ9nPntAc0Ck1B1WAVz3D7JFD3s1zE76og3TRNK/0eB8rdQ5yfgx
9P/7g77BYNceUmmIrycCTk/mjmOb2hxYNe+D7rQHAC0+zvSLthEwnhj3mIcE7BRxZASA7NYpBMTo
klX5SJV+ZXrQO7vAGhu1hWsXb9e+N6c72QSBwcJznnD0poVomLyclsBZEPDu8evFPlQzXbvHC0wQ
YBAvAdN2rLHRix2oTli1pQsg2BAIYPI8FOThweOQ8QJxO6R/ULdAVAvLfUo7tTA2btlA9z2NLa7v
jNyysYOmyWvYJWaqe7735r1Mv9MqlRaJARdH28nCq6oc1eO8j4zDF4liCXmFHTaHMLfZuuNOVCX2
laJ5+5OKitnGO5yjAyWiCbaWuE8rWVx0FkSbvzEEYBoDw8Uv1ptE49OPLRMDUYV6Bqw+8iSmH7lz
9ar0Km0dwUQvO2TiBIGLlLZTyOiESd6OVrnzyNcIUnFfVy639+CDC2o09e4aw8dPWWOWfxrIAPZP
yWNW9d9USSw/e8PFwB334ha01+QATDCuENbooBzHkNeiCvr8tr9CDK5pVgR5OtdqKsrWWbS+oqZo
fvj7A6mG3oJytD8QdslTq922CvvnTPJrxSTBnnyt/tZzlab2TYeN2bQUs6cyKUtR/ThyGguSFIB1
kKPiKnxzloanHrwQp0gxipNsEy1AVP4M5jInuq6m1XoP3VmjhIGlESDDGxnXGyuQ4RIHsrZE2Qbk
jNAMAUaUv3vrH8OYrFBXQ1awzssJLAeyseW86sjfsfd0LSaT35b2/VCBR1nnL94Kdd4/j1hyGeRz
HF0LGXgF6D427i7j37dTzBLC+AZXbJ1d8ShjIW/bnuGFFAZrpG6K4rqxi5GMYdiPtw9lPvyUxwSs
m6HsmYVfF5Ow3+VUv5Ekn805G/5IXywrvrFvkn7AJcFupp8+QiBtQBaIYex6NENr67seeKe39fsB
XR+KFEGydGjAVsX1R7gziATZgCeaIpdRiR9vvUDSUtAcibuE5WLiu+qCv9TRp42koKgJaNxrMq4o
/v6PLgMqjLFcj1ticcb6nlh3u+rDw+XYkMpoRkkk9W+EuUsQFfff48MCn5GvEQLHqvv0QWxqBgOC
jRDSBWIuQR0jDtWpWUHiV7sce0M1RZI7Oa/1B5Qd0rsyH5o4EMxNTzynZ+SfD/bNBvIF5gj/rJ3l
wh7Wkva1VCMNgkK5JAubScluX2AMis5TfNYmUDjqUACfU22DZKzn5ufFff2Bsf3Lx4+XvjiwqQPL
RpGkrRwc10nS/yxh9tZRLxTtzR8Om1yZTQP9sZJ/vImLW+xciLyX8gLXbnXZPtXyU7gGW+5opYVi
w4GEs3pu0Zb23FAugtQ3+uxeAozJQ8G1P7MHm/PJZAw5fFDDMptsKjljI+p51E77B1INB/28eN2T
nRCrXkd6ANSdrp4hE23Zc8MmxYpZepSJkU/iH2IMZG10gPqs4jzyDEsEgBCtto90A5oILrKsSX0G
5Lncr+iqUJAQErRvwujAdflxISMCNrbwKbXmnVjvpjVWmKT4Y80zbWBEZbtSz6IS70PVTM6j+wMQ
ms6UyyWbr6/TpOn4+tziJ6azfqhcX1MIbtqawb/s6pnPbQZ4pUBVYO9SBT45ir1lrm27ua6FvmWs
vuTE8d0CJUpWjKI1aYrzH/MQO19Y2H4oZ8DQCLvMlNTR8mnVSgV5rba1MF2dXUzp82KFIEtnHK0Q
qInSM1yu5iTIOIrT7QJ6asGLUXti7qe0R2oesmyRAAtQnyb/bzBFn+E91Z3ttu82muFC2WAqlfvD
lWnnBgfFhzTWvZlALgztSVQLkGEtcpB+k9tRslhCIwsHKkHady3A+mkgm/teQIi8z7NmIwkXVOh9
vG7ePz9pSgmnw6RZhfKqlUfVBsdf92nETCcJmQx8PqcpTevzFAwsxj85gYna0j+yGzSiYyrO044y
b/DVfPX1qxrJINLG5FoWdfL8XALkJOiaxkEod97Hx8jG9Q2Nbbgl9BSkWl8nmoLdmpK137yg4dlO
BCxMcgEC4desyB1CPGis9gNiYC/Eh6p/HO3sz5xQvcOLUAMOwSeKessXLzhrLdTk8dAmu7XSHZPf
V3PwUs1Rr/Ul0VZk7o+MOH1qqHzZX8ZqVjNrEbEXkqUjt/nN80BwP5zRcqsq15mRmqKS8gooThHw
0rLqUTDiNSji0f4RdfgbQzBKUh10Z61kSZEl/hoie2WBCS8rrRAenS5hpmkSNX7Hs/pA/W9Dz/Sr
dJjee+gtqZMHYR5HN2+PYDFY4KPjc53FL6nqaAjXsCFarE30q5zaC/hHbVMWmctoZhrapd5S639I
xV81sKsViTK05b26ELoi4VR3Bl7oSTiEVu11XMVCBKWVNbUrVztOK5B9CPaYr6agf4uBd6vJie1w
+FEoIcIMeHnCxS27LR8LafBlpcRYlLBZW0ChVPeIZS5P4Ar9XQH0gF+AAA6HAvbS43LzuL5FxXiR
im4D9HSNwcn6WdByc4rpBua8usHsguBtI8giQhA3NUoHEv/Br0KKJz21Rx+NLj6FcUX4ISUZnYLX
D3q/+05a1mIXPGkDyhM5oYVRL4Utcw7peCUu1WpENxsYQBBHWHahUxghY1kgE71MCJIVYCmXq9KQ
frFktyGPyRUmmaspSkwKuLkGTXYSvCCjOjChv+jrcyFh6/0oskSnbeJE4AvDG8nJWw3OC+yFc3RW
cgN8P9z+OF9ZoOVTr0LCdNRK8WLmvBTBz+QFsMgEeRbpi/Ze+mJvYn5etNrKgiQ7qN6tMrGX3gyz
htzPGrn7Pzti/GJObt8AZEWc3wH2UB4o9AYxVVuZXQpncUSyeIlC6PFcB7U7FGQEQdT1pcHtXQPa
aDWPCRJnyeWBaUZ84MEPmQIRzs64tFUV1Bek7Y+YJCqUxOVjRh1nGiNuej6fWsdncqDP+AYleAWl
g6BEU/cd3+ivpPYK+Belv5rbHuba6b+RulS8tAJ+W0fATXqPoHxPIWKRet0XEUgY50DSVFTjxu8o
CngzfIoTMfxVbieVSxWJZxJaDIvdYemR6h4zWUS2GHKOByGaPErAsDhvOmhTK12A9Q7SeR3PTAdd
y7Cf0RRfYClpCt7MXEEomgb2s057JlRCQP05x6jWg4rEsQ901K8S00bqFkTXgCY4aXYO6allra7w
GvWRVOH+4Rewapx75cwQnZpE6p2zgMpoP2A985v4ClIbJjcjl1Zpq/v4i51K7eMN8UoDYL8+p+N2
dGORwKhfeqs/8ntaeCuI+VRqBtcmP8FxaJHMFasMDn9NrKAdjQgY0Jwb1Sjf7rOXMrtR5Lap4mX2
Mc1YEb4v/D+TpGZMKFZhrVEzYpe6JlD13HOGutHHwSm3mzb3c9KkMkOkgtkNlSbowQW6mLd6p8sB
j1eSM3NSgdhb4kqcwegKVE1MhxmKNc3wPyxRXJ/rMeOP4zc+Wjv7aMVVySPJKao73u8PaOcxrkzj
AzcQQhqoejju1mggaTCKYH/3kRwi16bme+htScUH3BWagSWJnn2eaSohon3cLlrkjPLyM6KA8SDd
+FAgflwiYXCv6Wsn2MpZbtpxPSDsadsGaIlITZbEBKF+AmbKBMcHsSHiuxiFf2eRXWCvNuK/qnyo
A72zRIXPxYNL/3eD2EmvURMXeQCwMw4zBdGw6y6LG8LMs4w7zdHiKNakDBjB6r7evOi2jdi9iThC
d7MYOaoXR7U6DiV0tyspKwvfPz+DYAr5+0YdqEKFyiKbZaDCY5/5r9BN359S2h59oV5cyhmJDblg
ka3nshc/GohzLtNkqeCzNOkAN4VyftBWCLXObvLpGw0JtdkTuJNW6VEAx5JnvHDU6m8MympwnUJo
NO/SubgZHQCoRK/wW8tf/NgioM0FzdcohrNwy28us9JZeWrJ6zho2rWpLfxSmHY8nsfjdi/uLK6W
1O5bJzZBFBBjGUv/3W/jZBLwiOHY7clKvACTrZJWU7kP/xeWl91NN6Vnho1BuduHe04iwFvqj/2k
/5UnagHv2NEk6gRfW5y1n+jqgz8JrykW+HnUulw9xFKdOePTQCjgvmtmIbvHWyQN/wDRcWRDjaNL
cc3a3WLJbV+uPVMLj6zQicbV5HSKGB5o4/S0IonDfPqp/O1AilN6+feDxuLcU710HJDns6pCA3pk
Ott9jj/9xuen8pKxs3E96u/lB6nHGyaAnkt00/3JZQzq6/vKiX8f/v7Cp5RUewMc6aPylT+NiZ6G
ohxRX/Yx0YlZlzqc70aEVPtzUJ847zZZMuBwjoyWFv0W+cG847sxQUY6DVXUsQoexNMR1AMh+gAf
9lnRW2ntJhYKVppxGbLij4T6AtDaL0UloK1vKoJV464oUmz3kgFAsUz9i0gSfhyi/zpk+9lbL++7
smUk5Gzo9MGRdB6QFNo0OMz4dFcM2Xqei5vhwExRZ20ujFOydVKA89uLSybtZk28nUIvKB7FNOXr
hIt9DVYHQFCy+EQk3d6shbxiGKagZH8G4C+Aa+Vr+Ohi3p+wq2lgl+1xw262XYpmrvodEfnXupR9
m8lHt18gulymrnCw8FFlxykArofnNJcteyR9Pk6ndhRYPGEEbTBu1DjZqgDNvbKFz5jB1eG/C12v
QJ0mXOXpGcq9H/F0V1oJ2HDpFnGyqD5fghTlDaWHRSyLsc8cN7LkkMJdFb/tblKnwMDkdRyYAPij
GAhhJp25J6wLMDafSLEKrM81Gs8bJXdAy4L5hr/3K9HAE7DxizsvvS65YEXN8TgsF2mi+FXBhONn
1eAdKrNKUrmkMBEQf1utSlpmtQPZWsRPBF7XiJNGmTHSxU7cdta2zvGD/egEDFeoiQQ3e519y2oF
rQ6pCdsLYdMCNz/oN6T6Oe/PYzYrAS7RtJdxm5vEu+HCI4aCIEeuIFPF72zJHo9Bc+X0ZfBbgvZo
yoGN9h5Qk9TCKaiVs5i18YCXbzCKyiEei7dnQMVao9q9ahO0hH4tGeYU0TVuf+WXj6H1mq937Tz+
CEqapLueEryuTpweilpZcZs4HKn63fu8u4gqlBC/u4FnZ4Ja+QBALPqxtVrzTA7jUEDplIwRqhcD
Jz0fC2FWPglxepRx0xwF//5EJvfH+IVVVAN3CWFMJwXL2no6/05TVAfnKYCHGuoI+aswAmRHKLFw
p3jPwvOlE/HMd54gfQd2MrLifcE6SLbDfEMPEz2CW2VCUOnh1PbS5q+DHTnuOx2EC4ZJfcj7XuBl
g3j15nOvMX1gAXSY9LyLlajdtdSthFGtBEOYoGSBCvsDsWJHWwGMw+wPUsh8upafUafDMJJIs48P
5kneglUs5fWyWGseNFeaFobn4Q0ISVRpsu8nA55woZizjsIKwq/dt3AbC/O9AQX432CGcSCgvkHK
T2B7lOWrV0GUAwhAEEvptvS8MXoXFohRfEBGveY26E3c890rzbUF1/LarwDob861r3zSL53YfHAo
pMs4CVre6OKl7hAM2fEsWae5f7p9TVHKtGr0dj0msDsum0UxHQoT9Unw6KTHRe7AGdC82qJnmcTc
yoyF5j58KNcO7K/PjX4KVT+dUB2Mwct67H3HV4c/TulmLoDlikRMOl0sKIQlJ/njlgX9EbOhx2aY
uEkaAfYQqi01onjdJ32SrH6s8Iohk1vrJ3OLaNPW0hjnj20oaDwn0HHirCho39e1x63P7PUUrYBV
vIT2sTuV7u8J1WzyC1QvtpPSxh8yoAX15lK88QEqEJAWujHPd2X8VmfZ3AbLrBEexjx6MWTLSPER
30tJ7uD594dV/6VhxxH/MOo+N+pHOt07XwgPdp16xiURsZFg9Zydf7GQ+xd90uh/eXMXxUTDQXy7
Gt9zdn3LiA+u7nLiVnY+fZb2/YaR+Nm5SfnCFA4iIWE0DUfdnfjyIzmxWfNBy7vlZAHmE2YsWWCQ
FGe5ey6kJiWeK9PfOqEQWsqiRVxzrWWIebL9mLct3rAfPPL3UQGOZtvic9GR20EbZJMjAJnqt6xA
Id+1sz6u9SJaALBX6Gd03cvoyQqkvi1Xx7svlbOQF4Y635AJRVe78LImEEiRvs/ldBqz0pZPeGr7
F0YJQFnl03MhzHiFI3IX1osh+aQjPKtiuW+yJfzfzmu677pP40yR+tMwz4gOLm6AizCa2zx8t80M
SwSFOLxW9DozElxRLEdg7rbiWDmm5qizTeyL+ZmdAym+YjXLKj3E3FUEg+FjQ47m9U2GRxM1Sr2t
wbxVBx2uv2aKel21lfg+fU8T+FDmG9jE+w/lk7fD7lpXVG7Sl0mQp0MTNLiayraWtKoRTrueJyy3
X8XFS7yVcninufrKZny2gKud05K5h4pMoDG2rlBCor5F3YAK3GuvmRC+2Ev/l9HJf7puTMIgG5wA
V/vvdttq7t4CYy9pgRXdKP0jG+5VfvYJXobHPhKk/QxVSV3tC0q/9nVgbRaBOUCd8hPdmpwgu0r+
OARfw6cutdnIuNy3X/jiZoqCsYytPP7M8EB4OlrbtPtT7wNvxSIX9ZiD+T7CVJvvjXhewOmCkVVt
pHnWwWEUPzRLuv7KuPcco3E5gzKUqGvWnVLjPlS9vW+1ArtAA2hk/0cOBMRovZrbmR80KiieG8r/
JWS0WAjSCJhFKzZl5XeFi7tLbLBn+CepgNYpSyMSW56XtDk4hiyu4qgxTUF6EtGuMvaD91i6FJq1
HpJTaPLcpdW/f/73QlIb5m9MF5psV22LL7ZZ5sgPDb8w+nC0u/EriZBw1Yc7kzPopfewV+e8wrzk
n5ml/BqAu/K+PIZ2LmQefaGUA6Wa0Na7bEyTP6a37Td5otoVP9GrZplkuDyp12+FYoV0HD/5omSB
t3NwYdhuZO3+mIHLQzSMWyeAyZ9mvFZA7uC0TOUbs42h1Pn03o0rqluhMJtns7/Mc8DZi+vj5OWN
rntKlF6lMnLuojxqx+vX911/4y4zTYc7Oxvz5dNoA02STMuAlMiI6MBrr3p+pwHWXU5j/XVFQNxi
3zJmU4ZZvQCl3+9U4ef09Qe3DRnPHkNJR6nCsDSE00jbKqNWx4Rck7FWjrnnI+dBjVOVaNVtzB2k
mh5XLDaeUm062tGXRT0vA8fv+mPAVzpOHQeJKVJPorrMLJzInA6y71r78Fj/B+qkx9kcPTJOxcoP
0OaKJr/EuuTJ43GjhYBGaaCELqJB/9u7VDjgOppBP21iYIXbaxD0N+K8kwKQMthti7oHPqhoYzDi
nmrUra3aJ5Qrg+r5agrnPj/f0pdcPpvlBbllU8YOhrPiCDdeAGRXZABSK42smwJT2ZZAQkOL6S4z
NPUfgW5EPfrvwKxY0jhLxJ5g1TNWrfkycGDkIRR0GmWi+3IW1a8wytIkIdJe0Xlbes6ljdlqkPJv
Utz5ns14KMPUHpkPvKigu2J2QSnBao68Hl197tprKWhTrM9PZokI5Gj8EQ6MBSiE+dX8s8w5vUuu
tN+rp11+cscQdT6L2T9o+FEajUFFHk11vBtfs6g51KBvD8U24asBKmzckQnd6Zy1uZOYBPdrHnI5
TUSClB7yn/S9r/nvpndY06L0li/62lJGvBdtyuBt7iai3PGt4EKXuvr///OJQC7Q248W/zTSDfk8
JdRLvaa7VDbm8aJtfYQQ4/s8QhWUm5I9kCybEaFmtp9xq8oKWtRNZXuo9+UOJf0MEgYoA+N0PZOB
D1E7UHbQt9+IT53ne9+FjNlj/Plv+eZjfHnmF2B8Q5FXX/i+5HeTZ7tUlWoFKfbEXQMLxaSklQXD
7cnexqwR4uF/9EVy8lbMQSW3F/2PNCIsBtmSaRjXg18hT9jcrgV+3bwyMLyZqkB7RDE83T89SzdP
hpfyddrJkmxRNilrH4wpK3baszXddeUjb2Dx82GB9JmjOvNAyKFfc8p0c59V0F+jLhghRWiYVWty
peKAxU9zOBg76C2lZdhPJlpRFb/u8pZNRulzN92LAlQehCNSmlXpgH2BftY8onNTjJ1bdKOaXpQL
nEnYlyiN3DoXESRzm0RE1FjiM+b8MwjV9Ty5kX7AXkQqY4zS757xMPcNLRCnP5UCk6EP6s4f5aH8
JCzRgLI3LUAjU3VQyzWywy1HvoMWO5vLg0/q6N7GX4wdXOA7VVv5Lx4q1tx63qENUZRIIkcawLv8
pnfb33ZmyYe2tDAw/fT5/6nOPQ9ALTK7xkS5+W7FAYRipbHq/3DKrPR84lYiL2XG0MHlK80mdftr
JXsEDiHP7Yt+DKpZ6bB1WIGiThyVuRq0sto+O1YjAtdSnq4jPFd58t9F37m5Qa/2Jfx/ahXU5jMs
t7J+cHP+BsLisEMU/0+w6F8UhM1HEhDY/FCo3Jg/pamGsKmAwKe16rCS86TQwM0Gm9yJMxyJb0nh
cDwIWuwibURxcTMqmhQ7l06TjTfouaSVeg9/7iRVS04Ws8sevdjFFlBlHqWnqp0erC3g4PTtj5/p
sractseivdDVVdQkja/uDZQZSY7oSaCkjlAZSJZc1IcSC29W9+cvDJfDuut8ByshEC2Vl9FwnEwj
MTwa76MlhYx53GL73MvdR51EXLEZJcqchX2/mjtcHAh/gsS90WovPkXyw9xDgpck0TiHxb+UNXTQ
XEMzqplgQkPb7t/lsw5Ty5JV1v9R44eb9NZ6A+3QKNDRIsObekiLff98YZzxxA21M7zQzPANBihD
DWvTTi4W0RrpLOklxwGgWdnsZMp6v0B/Hb+lQ4GNFVNAquasTrqbgvekh4e1gXStjSyBfpJtPOGf
bp81GJF5UlYtoHj1Dchgp8nmiIFZkYZBnQL6Te6B15RAoEvLFKuvr5s7iGQi5zU9KeDDqw339V0L
GzwqhWCQU9RN8ll05N2mb/5PCG9/81pz23Ug1AMcF/a6mlHatNS1G4+6nCucg9L4f/l6x9twuf2O
NBNxPI7b0KNj/xiqKUxtxJGxQOHeME1uvGF+tNZNYvUwoHjanLc+4Of9xEtoRMayUviLIvo1XW71
jGYgVIlRNvjZJ9/5H5s1AWyWAV3GtzW8bxq0qFbVt+sD/OiZVIdgA8/kyVh6dKK6upeM1ahNZyhr
7nvv1U25rbUAm1wuaJfZcxyJC0DQRoouX9jnghia655zZw9Tif5BJ5CP5Rqea4yeMNm7R1QQQRsw
/WZTVvjd1GEkZyv5QENqRJJa8ZT+XyC71iiU4e3Kc4UmMGDu5erzG5SYUYp7sA2Q0uJdUp/EVORT
cp/U00+fp37KqPcw5zUaG7GMU8f++KdRPVRQIEsInUwa0BkhghT6rhmGSzMEXiQhINZNBoItNAcB
FONmZPHcQc3jxmx5kmheHl3jAG6vJWbnTRdugirQ7EAtTlejlvfxACzY91LuwIS4pvG07wRBBol6
SqL10cmQ0enIKWGD1jjpXyl+kacKoJqj12QAgrBcsdO+HKxRFsgv9IfpDLUWfIgQhbFq6bb3rucG
+cMbmG+kVJI1HjZTSNow27HD5/2HHGbM9+ruhlZyn1+P83CvBx/GKlhTXgR9qO9yCaWQZrxmJ2aX
7nSQfPcDT6JvJOCuDSP9TtDZzOxkPii4zbBTIFBIxjGIZoEDgQ1CTX+DYumxA0O3d8+SiktWVAc3
dRhD71KW58z/g7S7UAFQDRMZ7YA4UnLIbORGKohpCftiTwi7uyT1XtU0htjEeRD9SjZJ1fLUf7eY
KMiRWNb1YZb7AREhUljHwMuCpNwcsHyg28AVeUVxxqHw+68kXKM7dBLLViGF0+fbAIx8+xjfd0Xf
NWfVKvbAn1/ypvMn3xvtFVs0byWM/N/kDM6AU4fX9v1zDoMTOq9Rj9VMNoxtAs3oIFIcHWPjEUTS
BJyRcm26vhhVoVHQS2bPnS+ZcA4xQkBmZYeL+Sz0ppKorC2J0viSKkiOPnXHg6a626H//DGkY9+G
I+POmUm/WDIalp8cOtmgPPGfWTs/elipiqXp4ghY13kwfvGelpKI82yWn526yoKrR//WjDDVamsd
IiCw41y0huLTZcGaVwMj4Lmxj6VROx+enHopFaqrotijaevW+srmjjL/1l4MmkODkWrXlHI7BIv6
tD2PZkNdQPV212DGD4KHVE5JjXnTgTyMLgmgoQohw19EnMUFe90yVZKdtvGw+iGQHUac9tbqZHAb
RU5oqigyU65PrsW96hmI+CMTjgRnGQFBQ/JweqhszqBcmlr/f2Khvb4PEPSMfYtHkc9dxevfHwOt
pBvEdjABhma5cFy6q/bfXAyDUKG2kmeZRUXJ6s7vmRutMt2B0t32jIIU49H8fK78r7m309vAhTk4
UDD+B/ahL978ot5BqAT7Mp82HiWXH7RXzvX+VGCrIDXTkf3nCSKi8EDRSM2rlL9A6cXGmNladzSB
RmngqAuLQYiYy9a/ToOPX3aeZWOFn3TMSqT1BktVe0FuFqK2BSIsA/13aj/Vq5hgFbnQLjDmE7HC
mn1zJYMQHNBZxu1Y9Wfu9YtHRcoXXNGoutOk/2FclO62gxvYIBIBjj22wOQbfjVht1ZdQ4ktwrM1
yAs3kXCISW1XX7tPDQ4tJ9bcidQZQfaFEykK/lvS24I5qvAw84r2EdTJsnS1rzNMoJKfNLW1xP1W
Qyq1cqH7kqel0OXV2NraFS9jcu+BVigwsYg1YREcH3SDXzNZc/9RpoGF4BiLpPtQOHIQtymNvuui
jQR95v34p6vWGmp4xJmKTJ+o5v/JoJtVWubhBcmEZ4N8oxhVupBasaKFUmSsUxKTwkul0aKQ9FVJ
ilCyfLRri6V9eYxI29K9PStY+pgA0MwEf7GnKvvRqYSM3tkLgV7mwhIqNlFJd1AQY+jTbd5M23Z1
vE7v4PVMTnVMX+nFVyeMp7A4lEmXbHJIa4dRhGbOtGb5ovnYKvM+DEhNzvZ2p/52uzdTWRDWw6/g
hKVbabr9sVqti5CcG2UeBlrSZ8BuEdXokgkrO0Bss6tvV712TcASvck43wgaRGD0FQxz3XShrHg6
bmeHtH/MrO6cgnunFzPPEY1mEacQpnw1hFbjKWS5OR/dNEuChHDBYErR9qzfDTHkGL1EwgdnFXQ+
ImC668v5ygbmW1AGF1bqczl5dKoVN7+C3ivfF8JBD364vrtwahFZ1JOZFDun0vh8nMbIj0sbBsRt
kAb9r3/DFVXpMkPOuRJanrw/gzt+QpIlmT+/v7Iz6NWMrMFfn85wqjLU2psPsgmMMeFLAloI7WSe
b8f3TlkoSmWRm+t0B/HHYBChkqiMtBFr8TtyjXTzGkZD+yUEVNjPf2020kYzAMPVTXxAF9NrthkP
jfHqt1JJ392lwppHUXQPZNyPYJtk/S0orG7uR0WiWj/+wcvrZDpeLEQ7b7rCPbrK6iB7DA9iwWjk
iV89SPK4fxQGIfE0S/BtOyZX6hVOHWHyEihCFACGBLqiq7fDXdqubS+g6cy1+gGHc/friM6wr+uQ
J6ozApQzcwZYyjOPD/GBCSQWldpY5xWrgP9q0nWDuBQ/9JDmXs2i0zBl6pGBETR0JePW4mlTRkSA
wXVSKds75/8MPoHXyOqpeTeAsUqHcNZ7y8f+/AR7ahDuvGEmHehfj9UGo+lgAEt/LPg9RJgk3T5j
BkkClwwzL7IJBN0RMAEATzySyUMDpSUidDgkJ+Gs2Oo0N0Fm+FFip6vh+Nv3937+peH9LP99DSuo
fCIIvZj5vYE7CZZuHLknZuMIsBgrlrokRDge6h0y0gPi1FDryqNqyOoxgTHVdK46azPmQJqaPamf
+ngWGmnai+pLOltKxarfAh0uvPhezDvERpmYOJslN6g4XJ5VuwQuLB6sPJjia1uAaBXhZOs7dUzN
TX7GemnpK8zy4wA/oiwn8ESwai5sBLk6oa6gLy/QPen08AwTOraeUZ34JpEWzLjA1n3CNvn/fllP
4oBbFZNk9RlXD5MxF3AAufbo3/CtotMKUcVzF4yxFNThc/m54xYd5aYXP/lmuRosl/cnJgB7n8Sa
5bJBul8lmXSfbuNZuU5KT0aaR6vLU1oZMGu618ef6b8ji3KS8/t7fo6aPodJE6fNXaZgJtUPOwVP
6pqF7a+cjexYx6GP74qp+hbiI28xvYIc1t8y3jlv9XoB2NxBdvxXrRHVtLeVRsO71wjMj+6z6/+u
k2p6K56RqfSxXeo5vlA72n73hdQCX9foCN0R396GSwHa1WlSm2/fH/TtSSPHrkVaBIwbUjqgsONE
z9ifV0Lx0/tNYxJjvEJQHRThht38oiAKh+tELO0zq7zWDKzB8zhxcSis+nHnidgRgUPd8vSe3fUU
oFVK9o7FyTYGyHOCp7NjM8To1EBBW6Y0NV2LaJwjw3GPQNjpIexTzpwWNXpIy/0Ulbvj9l6vrjap
kvTsM1NqWuQU0x1NLRQuAGQ91vkzo+wPRGo01uCtzOim4R1BFHn4q23/P78scm/OEE+1UrAHhVt7
fapQPLxgt4PGlv4CH75slCGg3laZnWnudEv71/LnM4UIZ+Id1CQBpdKHOu1FqhGcVk/uoVDRMcrd
du/ieS5NOfhEeCiUJ6vyLKUbkPcIu1NpQqUYwU8/CjIMGkJ3GyrxTVnjwZJII59Jcds3GKb+vKa6
5Ni6Jb0Ey9WZ9aX/CvnMik9PU/DIqQ2X+ysdHsxTnQpntLr0Oeo+NeWDb9pskKEknMcfiJ7Qq63L
wSM3fGbsNvzavuV3PfOTQ3bO2sKAviiUKbW0gWdYADhyjIqcM1Ff5Oabspg6/6pPVRa9n4JM7uPE
VXH5Q/Pvc+S0QROi6WPVY8NJwmBqw7KKUtZrIDDSq+z8uhBKJo0IJQrCW0Ny9dCumi7AD0NloOtx
GKi0tvFvS3VlbLm+00QKChB8WGl/k2/x86VCdG/a9HQqZm4DSp0Oa0XPAzG1jElStPKteEWacp0a
wgquSWN8ddNs7mYfBcifKcFxTdnFHHtn8SjhuTZbhjL4h9EPQ14k7CWrE6L4pwXX4DzGA9YBXRTs
dFO6YIppp41fiR3ci2A4yVCtzSm9q/4h4NEOOL0vqaRienW+1QAI3E/8Qe696ZjlTn5GB+IUJysg
Oo3+XgvJzTfkrmRfZiM7fVdCbhCMSwvgfQ1JgQ1KnFkG2+jGoRuHgZjgulXZdjLvFnTF30VdhRHG
20MuN5Jbe+ACQ7qdvSIbnOQToeX0WyZ9zrazrKRcdXukIYbI4gdI5q0LtIki1WvYGs+fQvDNeGN+
hSyYh1tqyzO07QXZPguYCqse28UVxfQ7zAd3NYZO07a0fiNVbt00t8O0BlKdIHquqFGCUSxvUs4K
/C9K9AQGdWUtvQrYi4+ATq0GtOPhoLjtyVSAQIluv8GsqzFAwsL+W81yZS177AvliCtXmf42xM4M
2J7aZbZ2unAk5sa9rwzCt032hJGKrUfVDd4W093S0lc2OcIl45UKOgNtTl1g/ECeBRWfNdw6d0FW
vN6elDvc/bmlwKGiILAuomfxGE4nfnBxUzbTtIm4zOyRF1JIvN9cTm/5pKXAQUxYWS+z7DFIUFml
fESbSxKSzsXPpkYslj/OL38+/hp8iTDk/1jiCnzxxT8kCE/4XhMzoCFjDzHCiwFKpbCOHscIXys1
fZsAuSKGgnjq268p/7oR8rW00oOoZHWSJnD4ewS5FHgrjGcda4hlj5eTrjIPoKv7eSWi1u3sqGbb
uf4EBXjuUriaAHMQNEdtXT+bTcrBHRY//89Aa/qZOnsAOQUmYeB02vdf3YR2f7giAizqt6GkA1DS
h/P5cvmoBxhb0TK6YvZrb+gHhYz63cD01KiPmcVmwMJtXs5D2wvedguq9yyQUF3ED1IhKxVKAwEJ
Dn3lwuCUv+EtKVpmkffvx9uYOWqd2AZN30h9nBoDHpmLbqylx765mNvt6t+ZRCi2pfuNK6ShdZaQ
qRyBZOsG5j5Z0OmmE2pe+4ofYiFhy2QTCSjKZq3vVHlSgVWARIalbiEKIZsuqmeW0KrYB1Yzb6jP
6XyQk7CTHnGX3FtWF4N/bnwxHUeGjk1+B5s7grGNUZpX10g7enf7A2p+wM83u2w4AsFt/+C/oBYu
n8RN0VJg4RzqhyBCEv/c6zrAI1zwupSkY0QOUDQoUkf0kV4BvjJ93QV2zI4ddw7XW2jNUCd+XVX3
/DRQqhqYQQge/VNLcD5+ofSswvDti3CSkp7pRXllGdgsAR2tUJCTLySW1EaGRbHKmEB2uoJAejhD
UN/X3zf80zZf7x3D98I2Jg0nG17i2/Joo135aD35fLNLaemP6y0GIieWmRFBWvveAJHb9YiXVX7O
sLNfmRCN7848ntc51s2p3nWTmtF5ikW6CBjIh8bIP0e8VTswuk97latw+dBZw6kN9hwAXqNirJiD
xro4DsOfQ9FtHiSgQ8rT1hDs6Aavj3tDrWLltQzz+P1RQ/Ka+rSZwOwZt+vhLZpn/XhelN1YVXAd
WJa+EwdO1K1PCfBHSAwdP/1xwh7Q3Jh53wX1CjgAVdRTKQioYs3HX6wSNzJETnSpGGjXbmTVyWkk
oNMpl41owP9LhA1PBtfTAYtFAuOchuNVefEACeh8y43YHPMu1eUEVUhsaPUn3h/NmJg+XU9K5kMm
TOGKKyhf2dVzhlZyCxUSJKoJMHHwr+h12NEMlvnxVZfWfPQOa0TDMwqFu0g9ZvQ32n++7/26674b
Fp+BDTMb3MW+xJ91R14EdgrC/OLY3b1BG+6xVneX59INM2J2bAWAra2q3zDmvL1j461Bpe4IiE/g
jrdZmprChFkZw/jfSun+0w/ptnY1mBJ5IIKegKqzSeEK00AVLqUFfp2LFoxayp32xFs76UVsKMBY
rMwoUb+yhVXbjv4S4GZVSLNp3Ep2xh01LU6+b6UnB1L2Y7Z5tmg2v+pVVySUeA9aA0nuRFMSr6bx
SwlU5g0CgGo9ndaCvheARFG2h6zjhUxSx15TVKJP3sHFJ18ETk114/yThQ0CqQEwR0HJlGH4RgYi
gfZxJHRvw7OfTV4bbP7xAjF9/E9zkWVatMs3kcqk9bQRkikRwRSCR1ExZcflmog0AcBcKe0Ft60Z
msm0U+c3tb/BzTdhv/JVcismC8BjcjYERRH3L4U11CxcVvS1/XJmfHIf0iUxLoE67eFFIrTActPc
v1rUzsU9mYwPRGziJgecP+BpMPFb+1C0HSlLuJu3tVw3VtfQrIB4BUZ5YJMubtnhwt2GZiSOuWIJ
lcs+1lBYSyTjylUYKE9lDEAWihtb6QQ4BQ1P7LMAVwvQ6vr/aR87zQFUwsr7jsHZW6w9J7jSzckf
/GCh9UbYJMzEuI20daQr34PxJ7KHQy38xlUfSjmEiCl1Y1l55fPblIYoZduTqbPGeHsgBJVoYiIX
Fy1b6iyO6iuQ0mbsKcCtCNaefqPa2FxeO63xfoaOIT3Mmzx9BVTUjBK6fwLsj7b8ZWIJRG9F3tQG
zuQedr+8BTSb1O6U8jqheYipeOGQx1boN4FFMStiNVKMhV6+rHw7iTgX6gOo+vTDitoJmgsrUR7M
bq/1p9tzDr4puQg7HwIwCKlIvdCSdlKCD5GegJFvNpyHhCtmdt9UR6Zh6DLY1+1/H7+zYS+CxI1Z
CQYvMLVuEDUKyUuF/kkm2Dv27xdJWRPeQ1xPJbCq3oBIa1LYufGS4o9bvmUhOklm29VyacqP/XT7
Tl4G0BcG4zFZ7xCZ+lgtHTd2Byys8TBTkNjc2YBPz1vFBxCkHNZNp/M7YW7VyeM/l+w7hEjAsij3
t0YycqV1v+2kjN/9resKDkPWYx+u0wUS5UtqGRtNXKct+2cvK7eRUwLhQx/XMEU+k/m+kxeROmb2
r/r5/NIqZW/0TqjU104NMfieiIJiOIWEtB2QJ6DHtGOgJmLP+xF2ZbtVwtOvNbqsAPw7P1x8GUbX
KNRh7hmLKRBPVUFmK83F/hqB5H4/y9jeLxdT+usZ5uaLr99X1BoKkr+vAi5lDNGeEDpd5xEO7l9h
o8mcXunfiX2/5IBe7w4bYO5n4TUufEwNm6erxwVQc/Cd6mzxAD3xNVoZAvk+rffOIv4bFawtNi47
QqGx/nbAx0Z+d9VcsZ2/h7E5C10rUQPy+F5Im1UN5gZYeXagPBmZI57E+vpLyp0Q2HSU+0HtV/gD
TPZ148PblJ+OGruD3ZPwyhv9WclG0qXIXxx+7hAnAiv2LQfhLL1EWzuTsKY3gNexrfSsZU7QWCMA
qGxpnlYiTrZeg662K0rLwJlawcDFa+4GdlA0+vQqzxzvLrUzbsiJ9ta4pOUecouDCHbcdrRv0EhE
7OPP6U1DOLhPxNPPOCZlw+XDoZRPUHDuBlF1vHuouiyS3I2kAWnyhAeUocQaD+RnIrtt1kdzFQpO
9AUrq58TNKfC/dTDWmap35IIfGKhrdASRVDGIYo420MDZr48T+nUFhxnTKIEOoeMaUIZ7tYh/4IQ
5RDb185uVWr0hOx9i+79Rv268D044d8Qbc9k1I4l4zwxYWGUESYY+UG8HCy0KsbvwmBEpb4WsOXz
Y4/fDRgF3NXckNoc6JpBuv0ehiXBugegE9pivyHY10vHbvMRM04KJfA4IiFxey9qdsdiJrjfoUYh
ZraUDVuy+5MXoP5g8r4k9IGzgghkvtDyJi5yf/+lEIcxz1zOlgHGQ12r7UaXdJvBjXUnCfxo9U4P
DEwDFm6OMQroXfIAlH0NOW45EKpOkvotaEda7+cgoNca8/ap0cbstSYPEsExfQFc8FZZ8RWFJO8R
LvJMCU7MQ/zYIIPu/TiopdXoqoNU/cuktivAzhB0Hw/yvokvEojK68qECfKWbpmKz+FKlNr4UzmG
J42roPMXPuxMAm+ZHHrWX3LBiY9gawQM77xjIV1lD4SAvRD2WbWvSo6PbSIc0TvrFmTOHdPQQd92
BBSKk0WQsORJKua7zJ/O6jgRUmtyI27eiueGyoH1Yq+Id+1Ew2KOXiycaYRbRPMaEWTT+o21mrQH
gZ8ZNxtPMNq+BrFSXuC4RCf0RfJ0xphbGTstRjwZTkz93oujHQtl8niX7b71INJJIuwEgR+4IXk9
ooEEulugl+QI1/jbdRrOkpudA7toO4M7Drxzz8Pg4lruQQGaqM+UDNFnAbEbfX/el1Y72lBW6x6+
R6rBtuo3zrXkGgA17kYIZHRcP1iIUhRP31+upRLFNbb+dyG7R/LDgaMAHmpwCbpa77ueGfsn/TeA
2me1TZggVOLFcncoYWI4DegVN1oYu7Cwrxl/9trTwGEWCS6xff28inLWtVkGRJtvhDQ1rqYs1yyx
rRvWaTcBwO7LUfh0phA1+FtG8Ee8jYI28lzQPRRU0MgAxd7gkDZ07ihoYZw+dQeNCBiq6aG8MAYg
yqd588zgzS2iIes+6cO9mUAEvqj1rM4er1fA11nuWXEgAqG6Be/Pfhw+NIjdrlL9rZBhpZmCnyCI
fOtYf0ZDb78tLPsKtNbyf6kkej9q6t6eE3o5STFz7MEMFrbXiX6alqkBYee9slJUrZjZNx9DAmUR
RxbLppO+ZuDR9r9fJ2bokQawMCQqN77dRjDfXDuEDBLvaTwPLof+LyVq6L3otUcb7yKr+8jjsHZb
hetAxmZ66AcFEmVYCw+U+s+478hZKXnHAPcDnrAr1G4ZUdY6bgjuRJ9H8cH0pRiKXdokUdZqeOY2
osegf9XdojDakf245dijZCWPYPfL51gKGVIOxUDTC2G92FqpBhHpYG/YBjnr8bMeYjXyic3R6kMZ
cW7vEVtBOMLGW948HV9cYbDCz6xrRr12VjobLp1vbdPkkS2CRrDFpiuqLJoKVuLDg2EssAkrKUOl
2TBFaOPz4JhT5Y9/+0w227IX5+v1t+nRX6gpKZDPl3dOY0lFKj2coBR7yqKkQ7D9ezDJoAYSKbFm
8DAVX1RXizdLSil8Gm3tAT6eD7ytlAIz/R0g7e4A7skrWt3WTZixRbM50M/hI6P33Q9tT7al5etg
30ARSr3zEPW33AfVAPUl8DcG1hKKyJoLfu2x1/pWrZR9/ZGsrbqv7iUBPo1GeOwBmcoD8Q+Bdi6H
5X13KflF/uW9XJ02zefg0HlJo0UmVXNxeCRNJQHb+/Yu6d4U7IrWFTvElj5HjHVMBTAuT7QW8ZCV
RAH7RrdxzWrrNCNIE1oie9R5zRMA1DNaPng+XqzQ5mUZt2uJiwVwBEgDl5C622+n589ueD5YtzyV
zHU55+YfMNJXenljDyz6M4fK1Zglh2t3md55zJ9Bd3oSdCCzoeuGv3HHS13pg3iKq2ZSsNEWCWkM
C4XHn7bxZRZwDNUcEtUb/ka0yQJjoXCsbLYQF+dlu3iDJHsmIS6DUL8DQzMjiuJVT/BmD9av6LlU
DtkGjyqRy8GW7cek2ngP2Ttvozb2qVnKvudP38OUw5rRkVe9ZklKeD4eFMxleqtrR32t0d4h1E1R
/AQDsIV3LZxxf++Wb9tZIVCAcvBdFPNyknzWJNhEw5fFajgVFcgJCIbaoZnmKCscrOfiXR/6wd9y
txXiavQCbZwIgZ9ACHp38SlX/z70h408LbuEU/7SsTGVt1XjXeW1+6INwOzZhd8W9/a4LtqYDAO1
JZNzhEn8ZZTDNbjZDZVb3nxW5bOs8OwmHS73JRGOh1fBuILiFTwYcNXfEgCZr/kYdSUlv0Jur1Df
895SqT8cFdPtc/X0H6nC7Jv/sr7d3Aq2J9b1cfIxX0ho/2hLU585Rpca20uVYilSxTkxe/HqgkVK
ytIUOK+PBMbLFIvSWj8vQ8GI4RZe7iTT/h9pNy7aUC0bkJIGd+o+JuLw0jwX5emJWFDJjap3whmG
wJLDpWXuL0/B32BeHiI268L2VlzxoLgIe7Wb5SpCF+pZqlXS7n+rCFJ5CbvmCKfdh2FUop0kwbQy
k+NyI0uAQ3mhtty1I6KP/rugKUe3jOdD4xOCqvzu6pYLErmpmm/G1Cm708kPaUgCj5B+4dqLptdj
2eiQixH5tCkg6BW96KOOYdjZ4qH9ITJ+SmM1AZhBP95nZnvpMgQ1THI0MFpquIJPTdBo3E1kGdE8
KSvpEe+IU453rmyIALnyA1AmIHASYMp1D2n9xZkMyHjUO+GU7mMwPC+vRE5l4BvnNUMNFouW6f4F
F+tiDAd2E/rVdGcjXXgeONMmUevcl8p13U1Xb06YJk+WIPW9txMgI10AN29ZGvLHbpkY1o5PQ4Hc
qm0F54ArNsvyqtlsGsttuj+a+Sta90DO9f5SgJeiO7X4x8lLRPvvzcm6vWk8ISl6LPncKhyGTriU
RqyrQlaFx25i5qRHunmwNqeMAe74XCnpyK3++UIbWcA/sZeSXgkKkgUFrkXSKMK0GUlAaB0/d6Td
ekY37LbQCzf3s7pFTxcVnvXwnpH820aCxGhyDRxBlCWdMAf2STPpqcqm1AThGRT4cwzIykHpH0Q2
E2W8UgBfMjQM7+wGigU7iC2sJyLFlqSx3g/qeOuyWd8N5gxKrid7i9aTZ4aokY3LuL01UuGv2f+3
bQomAs+cLIXli7PoLFJY8fpalUZPR+66IWe8cWL7b8T8Ku2uGqstG+zo2NdTVgtBqhBTazL5p5je
VYGG65pzLDqJQSCkA/XVTNfIxqU153zV0p43nrkSCVCk4LE7iFslSGyXNOY7nqLdraVP5pox90IT
fsrXIWblUGmxFOyxhR0K0EgfaB2i6ImlF0fEn9arrI1Eh6QgZhgsaG+ijp00l/7gzBNBE2ECu98R
Mcgle9WsF9XU6ilvB+B06gIO5n+y6YbFQzzJRar/uwtSWgJ/qtQ+pKCEWSx4rYz5CyX3KGGezHCE
Ko1De5Z3KqSLS06UWrk3GBS98z89E0MpSf5SqU7xx047FET7sL8+LSv9ockRHNtF4TqiveAsUJWF
kv0s0vXJIJ9iGe51qfUANg6YaGrd8Jtp11xImpeZ/bEP5fzuJQIrEBifXpoRaHYaFRpKwPPpQYcR
/gLUCUA3S87Wb3gPndEhesa9Gxyc1mMqczrQvg4oq3l3sarBGZpGJ1bBtQU/9L0/f9GYhSUVpphn
k4i38D3f0jzKISj2c024G5thOOJ00gQFiGUgpNvn70/9I/4HLrXCyYXl1wakAN6V05uy5VNQgBD0
7nFQp+e63aAlI5St7IEBHFUOJFf0XmFhI2B3mNiu2+s1haWSLPNcF4cuPl+/E2CEnAJevla8issS
bKWL37yduiI404NtFqWSR+qM8+8F5NkEg8hCInhgAciBhNr3nZ8fbVFgNJ8j8eQ86iHrkfPzPdJW
8/+P0IuVCed29KlGDSPutXxKJ3E/51+n58WOQHomVt/czwKoTnL6U0BRTYExPZUyhIIiw0UUCP+W
MvFTOxmeHziqHha03EM/T6zk5tiwyCyHms9QuIAIRFVjGuHTdiOq3mMrtExo2Ye5S+2jvlpDdvwJ
Y/T3ZP1XLPq5nKyPH0EEVJ+23SBaxreSZZ7tre19iLj+eNaY8cM9uqirhGUfIFc6VvjB6vkB+102
hONCibvptaAfv2QK1xMnF7qgVbpXZWeWIKHSS3TDRGPcrtJXgji1cTYdH0ev38IEaWFViXrSjMq6
xAcjbLpxNqR6oLFzQcH0IRIjyEllwAcLe5oGFQlpsi4KbggIhQteQXiDNThiTdc8S6lRKpRew8uJ
EUnCoQothAIHMoLURJOkSSz0zX/MT+3Alyzq9pu1++4jlnfNDJc5MAkofrOee5wuVLgt+iJtsjlB
HpqIWd8gjLP5EicVotvHwEembeyWZ8WM7d/RokBv4d106ytflOfr0s6ykD8sA6bHsz3bPeuwwfuA
7a8NT/Z2euGQmskOMQ07CsIMmbu08fw6Zv3M2ZAhHAg5NmSca7uGZo9pF2fWNx2/5foCkzgAVh+a
Wnq3bXZksOrBMs/DDgAzvoeAN6DKwtKtbGR2FXMFnVVsdTnYw5hYwfjXTCcyVxsi9o8e8pBLSeES
zJe2qiZ6Hhr1okpREbZhYoIMiurTXBODj/lxctcGBsTIZRfl+cXijdcEJxL/tBNOkkC6j56Avyyw
VaTa4WXokqnzjGKyNwQ+qBvARfnVU141fKrEHa0OWeDvMWY4PHrRZCIZeqC22YEQP3Ekj7rr45Mq
Tf3LVDvmNw1tYsznOBnkqH7teibYU8aOksz0fPfafOInCENSL0Y/Im2crQWVQb7f6cK1pIY7F1g5
xC/KouVUPI1idAaBEPWBS1O22ZBXcjf5TwJgOKI1qQ+D/hnttTS23y1J5Io9DqKv54M2J2MMbgvH
m3N3t5EQGMixsN2ZVvSRNfLju2wwuFcEBxqyKR3Ulz1VcSV12KXiAwDHX7GYkVr3TEHZV1Czo2y6
qpNqGkE++PZzJXZiTHfGWr9uf+3/PNmYgUhvi45Htgd8ntTgdc/2/EAgz5gmCskzGu9VxXnGgHtJ
46vZFH6f0BCqPESBusBOOnb2eGxWQxFSFNnYWX/kQYiPGZsL9fCA4wNb9+Vp2KqMaqN1Epbvc4pr
LcUGg0ahensdxgIDB3KItKgwnW1lnwuZvL2h2+CjpacDVcbj541FTOfJLwh3AkEYvFk1/Q7kv9id
GaMtVcJKTIJgwoDUumcpv38hxBYdyHVIyx8ZL/Oerwfay/Lox6GAE424XuoeH5Ji6ZTIaiS4yAh2
psEogkv09Jk+9AWuK5c9FXF3ocuHVPSK2rwsZtQ6z9IWYrcdLChxzLG6M6dN065Gpp4IR+nALHtF
Dku42eOHjw1pxpay2PATeRpzB3JtFmrfDKFPAc2udP90mUYqzfGFNeuCFz+zB1783RIi8vn4MO07
bdsh3W4uHvVxeYwQ4+jOJpa3tRMGSJuUbRfHXqj1LWXO6AT0Pgp5147N8WwBycWkvcNSA6QB2jVR
UG/mgKVahi9hMEGuLo4BAzAqW93GtuWc9fx83EbYGnEEqWtATd828dH6gz0OtiP+5Xa2/PA9uB+P
gP3ZeSrStNF8rI+Si7RgKAn4A2KkI8wq6vg7ldj5HM+KaHvlu74Jev7kf7almIfQeXorXA/BVttr
KkMQxCIDgW1/WWucLggmhjWI6ulr2tjy9N1k0Kg4zgBHwk9O0OUEb3ae0XcH2+SaMBSPqg8iS/xU
sssmy8uVbfRtQr953DCzjVpLder43Rd9K6s0Uxd4WjLaYsRMTNQalfuPClt84eAB5Z/3n628mlrp
JR9DcjIEcGx4Hv25ojuVaoPb2tGzmwFzMobdLHBCbo2PJwnOFAqRzptd2b5tCa+Wff2edZIafaWa
VDxo7h/1RW6rxFl119UqOMelubidnF/ZZnmdN5uO6zkJZmYZD1QMiI+ikmBdPvD6PGhf4tJ9M2JE
Fn+FHYCBxvNPWNgfo+4WPvAPxsAY1wQ+cFCQP2A4GrHiOBllleUlZWNiFHak/7HKxn+NnAQLTZfY
H4SblqrQPiK286xGTxGF0aFRHODSmhmjaNb2MNmdg6Ms/h+F49GfMm4pNzHSniGoKVlTt2sYMq88
gTQCLCZEAbPKb2++OFf9R2AOhRNgUBQASn8sWsEpiJ1XvHA82JkmqX1SaaQiIfgNLAy0mhTJM8lv
5oU8UReLFSPx0aUTGhhmlSwPWclh4qO9i06RtMX69Ncs05jttKRTr65VdmrQAd7culEbE4jZnOw9
D2/YdSF9GQliUuatwtXedCcpbxxDOHo8gt4r8jbPCOb3aTSGCIXdyg7dn6FI6SLDJ/K4F9VTc80a
7j784mzw9QLTe5V+tI90kr7vK6G8eaDXPpSv2MsWblu7uEDtAQglgUeDLrURKrFB3nWE92RXoL//
Q5zG0iAHf8zUmAsJievjD40O8hzEiYnCGxtiYXFKSb3o8Zcgzax1/yU12alT+hlK65wf9ot46PP/
RnAObZbkCbhWV6Tr0rDtqrRf3kAtNQj4Euz8FE26dOYZ9ggUWtFqaATJRvQi1qgd8Sk0gmH8NEd7
bILfbomMn3VKNshciHP9Ee7TC6A+g3acVLWFwYGm8HRxlSG+BBQOvFTUBU8yMlIRakOWLQe+F2pP
v5R1GTaayRgHYUu9NrvnwVlgDVmjtBLyo3dST8blmt8yzQbex1VOm1ITIEiDeOZZMQaKP8lpc1Ry
f69OelDaiaDBYZP8u9ZWH0oFIeCcBSZFD7oCQXq+A95YVQK5YxzcILOtE0UFL7KvtiCwYi95ekWu
t03AL7Becbd3wOcA/2WUz2O6JpfKjPvvVlB3NqYghBlIq4j91aotaHN38SlHH/kXsWGPp+FUofLL
Wa9UOrMFhaXD0Wss02vtA/mggvDl7luWVEtzXl6+8ae8qv6ZzCbQeVFaZBWpqRwQ1r8C2cVGjOkZ
ztNp2Yfq/OuzsJQXaxsaBGvZthJUk9OP4U3T84YaluGuVa4dSjer+rO+AdUmyDNp8/MTmqR6sz8U
fRBI+pLeKyaFCNYHH8hXaREFei7RGLbmRixCmHF4jqRv+EUWsRR/GeM9/zGHVpQAMdqbemneTmrz
FPwOFh4B9HXa1jEHSF/zh3Ae9Sx3kyUbhL6iIrmO8c5AaeRkG0VtvugIpbDoFrwgOpDXdymCmoMn
UH7rTAOHKMBpGX2Drc92Q/cEX26EjbdEvldvb9sR/v45cW2oISr54eQZLjOhdAZYJ+dMUNFPa/Lq
CxB2XrPEG1R0KH8fDjqFfTTr+hxpCxC6NmoU8R2mjJ3KFTruDVDjpmtnpVt1Pnj3GjHsMr/CIm76
EtNoOdJFrLFL4eL456wvwHR6mxXe3TPlX6kmVwZvAjMLNrV2tiZzIvjbn81wK5IeWYsU3yZOGNn7
iXHC0o1qubH6ahYrlIyvzZYJxZyeim+aXAyfBtzipAz/PYf1hCc50qTp9c1uNeoQ4Dw2PYQy20F4
MoDhMa2zhZM9guWMFhIYIejUqStwCNp8+NvGTfcW7HpbbT/FczH1zCX5EorzjfCo1jvAG992H2Oa
psKe/tDjakVkbXP5JXaXls0bRV7ZM3l98qB8BnCvuQASZ98QF+GgFiNspsEQYtmIjrf0XFNCa2HE
AuKLSdilZWMPBDr+rLAekaw5sCeCibXClbzpQYLPnp1gRQis2iyhI5rV2nNSPIjhwwRQPmYuH2P1
u7YKKCFt98OiyHJ5yyVH393WANYtLMGWPECXxipgvcViGMj5rwOo7JIrruFHCramA6Msir1e8XLz
pyj9aLN0l1sFSdRvODa4XGUfEtlHtUftePbZeNbDJuXFuXvGKpU9koAkd1KQnURcodt9eoL25IKG
TaP93fr+agbyfy77MDSVPOea9HI3YKyEjxyGan2qDg3YcCUw5oz6fTCesutv1lp5mdCcrkL62Gcn
QUy6jlU0PKxZCeDtNEqT6WaeAq1zGuQYCmSu9jrKIJi/E+0rPwMUYIDgxc7LuG5p7S7SSyl7gEWj
AmlBsmnHMh7VHslUepxQIqZieUpJc0MEHVBag/d65tD3P1tWP0FzO65MWXQfpzelTyMiGTkshzUa
ManS5mVqLrW2g6HeFJaOdwCd3fvvF1E/l7rKpUiN+2q4XQTUUGRFonUn4ChwO/uk5Dm6sZ03j/DY
GohGl++VmDz/KwANGW/4+dJXK7wRGVm8q3iRS4NZYrvU0AdIwIsMUAmVuUBFtk8EAchI2gSGR8NL
kzhhWVKKyEMdkNbskFJbZhbshoXHoiuEw5HNeirGUA2guLx6w4ZqaXRAHltEX1bWEaxlp+PSx1hL
CzTABER5YkWlRnDbQjGtCodfxVpSsKK/yVvBg6wr6eEzB0jhczuFb4gMObaWS8U2ihMgStUe0FoK
p50nDYZhcpbdRBjS+JttiCI7mRVoeQJ29jZvu+2LopH4dPhOpAnEe8EIIC0MoVY2ox0y8UDraYYS
gp4kfXKhchgj6er1c6ZWKDq0ItVTU0QYc34Xd1pOFiJ/aj2BbUC9/moQkiKxtB1k/LVA37oNTH4q
8FDxYNhjwdAYM/7/ZMEtXzf6HPMSiIygtvtDkaM1YAEj4AezmhLepMDR5RZ0ErZAZT9M4az5mzbx
Go42bbw3DJebKOAx4NnnN185YCZqfUSn4xk6hP9CrKmrOhTeBO3ABIbyyTJlZViyekhvclpiGh8z
BumrnQvxiQJu8R+8Uog8L+EYaOtJwhj+Htx07OaNnFDY3ut4bS1czQnNRRQqv4Mc/N5ZH/JqcLv5
n6l1HWbTVFHmgqMac73MGFpTL+outod5RcbH+Wj/qosv4WOfcqTQF3CvLoEuvYiWcg9MDEg6pYJF
HhkmTqROkMHLViJf2q+lKKJgrrUVrIRpjeqBEWbBaiQ2ejKVMFITWIOvWQF5hM+MDCNoTvZkZZrD
HWie9PEez5/O3P8RQXUB/OVfbDf2WFTqXSc1RTlv2zVBvVqrXCGESpa+dpxr65tq2EbTVwulATRG
a3bbe4av3OIo8Thnj0jyHu29KOosxClAiyU10Ghl0Mb3G+UV3n6XZk7/OoyMQmQB1QELCQPwb1ko
/98KOjqkVjgTUj+jtRwbLapKGI0XMzLFKw3Yp7twQtXI1I2kOVkGfPHGLMnIv2oinabHlo9DULMS
5vvNGn4gxt5lYzfNXyJ6wYkyvupHLAtCXgacgUgULh97M0LKToU+EwEYY7sVSMB4XSFcMPtWoja3
mz/hdyvLuIcztKPCz78/UPpfYRp/aUjqljVggPtdnVNVqThyHqpcdFOZqPXZTzSdrOQ9PAKZ+z0g
fhKrR0r90qO/WoMGT2ihvUsIot9NGBtdS2nQBOUYBQVSK2Aws4Y1Gyy2uoi7E6PdWRP6S+BISWIM
vfm/hi9iamIOel1zSXcZQlh2/6bfbBCXxpdh3Atd8o+tH9gbsMnhMaMdZGUjjYSxJ+/DWMJSr7ac
sasJeoySNpPfxSwTU9afLRGbSjZIXM5SCZ80VIzfpYB/vOMuA/gCMbWx658twwMvdBciiT0b2NG/
mgzetJJwgVSQmtuHo1L2xSIsn4OpF9JnVtIdAUX37H4wgCAHFDKKI+hdyl9Dxs/JMKct6KckiISu
VaJSElFmGOwF84KsGtfBkuOl7CLfeAB6xEmWQnOToFgGAt9tvy8NoXVi+bWy6I6CReqmYK9wgFNf
g/piQbA3QFbPgM+rKXAkuKh91yhpwaegduoPVdWhWcU1o6XRY1468aSubaIQpO4ujXRz8JXzNpAF
hxiuYqLpqFTVha9LHAwJiNu2z8rdg9QOVqJyBhYOlQa2Twije4o5Xyq1376IqDpp6riI8ucQkosd
E2YpPmllYJPw240547JgCytz2gnD1sLgofYN8PZ1l5xn6xNnidMqhrK4s0GFf2JOD1pk6A7UYDma
azw3a/zmxdw+0RqsQApK/nMmfbffsquzYCMhe0wpRnV5Oj89TOjwnpl9DHOkbzvw/J/Ozm+Sk2vL
k46oOQWyYlW6IbhmPAc/uAhDkeL58/S09HPx9iC3St7ZYxa2gXcP31zDZfg7FOe5p+trD4noXUeC
ilW5jPclrg3yuPoobXU0SKywqtgRp5nRvwi+yoRkYOGtrRuEdkrtztjLZNThq/RFtg/1EGpHBSUO
NRtnVRzJ9cW0Dbm0xfsPc+x+/mXdWamEDX1JKAvaHRh2tFup2RNpU3SbJeLFqyGQlmro3QhuQIfn
hFVru+O79I8/2ub+eKIEGIRO3Hpb8cbB3ukDpbEfK7DOUOgOd2/1qUh9wbJKJuXyFLYsP/0GPnkZ
uW7on58WiWDNS1HNaTfnP/QlRIhfQxFrkelhmu24dAqWXCDCfjYxWjBwQr3X9ZEkh5PHZV2jCxPl
/V1cK867iDFLcX2+yb7h/oSYlhYZAiXj0D5YlDJvZIRrqHG8SYPAAFxZKmEQdPZ5dvkP7S9n8La8
nWiM5P/e+eCsYgM5JSHz4f4fjlPIWaKGroyex7uHEFqTonU6RW67zd51BBqsJEqf8ejEys+CY9MZ
MUZ0Wo6ZUxBJO0RgevUMVw7gN1TPfcFS00Y5EV1owWsnOQHHk5x7VEZHY5Y/Vbv6Bc2WCIXWrSNI
SlT86E97EU/Qf2/RAUVPkby/S3K8vRFlwT0EU9dUuiROdfnfjVWZiOLV7YUiD6pzHAufMe9Bxa60
KhgFvyiOJ8b6J2Mi3asWkR8nu1/gpjPLjnNHNntpyuscBY+zQml9YmIxLoh6SzyPiVfXT/RryJiR
+DcCOYtAW2Q0+D4tIqk0ZThfN2K7WB42VanncSU6udhGkIPSWG0Nyd3S3gTqR6g0VTY0FMLUSezp
vZe+ZUS75qbAvpeSWgXqu98jHNKjCOro5xE7j8CgS/yCRHMdu4d+GbMovq/wsDwIxKZ4KdoaWGQ4
Ysz4id318s9TnnZBBxKGXqNgUKqY5hN/ERzXPM7YYJj9qajyL3LwL+cTyj6/y/4RGNO1iAE8hRSw
QawUdrMlOX+D1MNKEzrfmygrL+0G+kAvn7wwn2yi8V9EypEhtw/f21Zk0xTzVernXXd7COdt47Fr
1uXKRP031YENvz5z3FGrzr9kPSI+Xjc1/vFV5swTf1v72YGPRcr/GZDkiRFODRzfUd7fjfKrl/Wi
UHbybv71Ff2dO8BDqy6GzrC4NLWpLWeOUdn8nsakiwwhqs/adWRKCY6I4uPBSPTrq9msZFHAF0v/
NPzGfzpXm9iWDrbvONKCaLv1r5rqUTgastWWTqmmM7laJckv+bW24VLKitcRtdUVRDWR1cpEFmy6
uE57TZymZzniFcbhzb4gAkVBuMaBNLgdxUOHb+EXGM+fpAyUWHc5N6r/OpGU0Bn/6EQyTZRfAXA9
+GV2Pu30+AKXbv3CsExajnSA6q8bjhQXOEWMYiZgaeuWln53JgrBVK7kXt+RUCV5k2nRL3VxEaxY
MUVbr9ia5gUySnCqC6QnJWtgN4RfHjDXIq3t8yMohvrQDiIU9/g99fQXHM0ZZKyP1bMdbwyI0fCS
Kwqe1/KpyTatqCAVxtEq6hPj6dEgfPCkQO6gHCP3DNNGaDFGCNHhaf4jNRsWGQViD1vOqaKNgJtZ
h5yHU4sk4ZfFdV1QeLvdMnvUWU42WuqBf2F21KZViWGmZrmxVyYi7DqA2AqO6pJZwrohMSN9PFjZ
ZtDOcW6yHa51mTaWE1jl8LqoE4UKJVeWwg1LzqE/otJov1cblfVhbwlfBEw1/I+lM5VVa+RKPl5z
d+/inWuvs0cC/brwNIU8bJLO5qwzy4dROrCn7MwfYxkm+XX6pScmuX1pNm7iqNla8lQFtGeAnWLG
3rUSae4nebCdNoXlXlLA8WZOSJaAQNQXnwxURO8xaERYJBNtHnMOKhnfsIBLbPT/+xjFY10H4ZCX
j5H3qwerCMmmlXJH01MqwRIMqRYBl8DTOvKVkTh6fGylKCxoLk/jluFCRvENAPIxK6u9XjJAuyC1
jPzXBDJQFwY+ZAZeBfmw/fpYKlw4Z2Y5C240MxdcPwprjJDbZaH7j8B8s1VaGGKu+hRkQPCEuPoF
u3bpI746VRtF6HaQXCg6weAEGAXhn3n06PO+7glcj6TmESh6T72tHYKyAlq8rxCBnXfXHcZmHjL3
o2s6R59Y/8BJJ2wC99E3d31mcZG1uMryX47iA7JXSWeJUPGoRojZ9in2LEWORVjOwd7idHSipvre
c/d+eMkfPhT5FYdwNCOLIbq6DPJt9KQfZmMd4L/o5/yE2uzz4/HyTzVx/VU4ccSfw+UAKisLTHNs
i+zZvC0zaWfacwIhnGaINzfI0GIoK97qnhadkik16uqVo+8JI0UwFngjL0k6fZtfKRdo2lZlajEX
Fwn0GJwiXNr521OkXzgOe6Pl8/rX7J+bYBJsVNCrQBE5ui5MIYIg9ZbFgP14osUGQP1owze1s1VX
5LR/A4tmyuVk8HtuKmtuvVzLKTy8+FxhLhlpHlfIUTYyeN8ZDtYlfWAsWFNKmGElH12RkEUSoFJ1
/GpjyYz4fOMOWuhWQC7/+QTErGbGeudLv/jFOODzG8Gl4XOiGLdQARmk4P8RWrNgquqhEA4TPplJ
mEBXQLA6XX31J7l3tnGqOLnLS0ZfeHdz9LU7ErnDcTBZalYQUQ671Dv38mEvSGNSAHT9W7cSy4P1
7SAvgVGO2Vkba1pVBGtpX/7M0yh5AYAlc6DYGArwf4r0yU0kYK9GQqi4GsLnz+plpW9crjUI4zsl
XlexKWlN8NstgImn+mImP2ScTkUvDpnv8pc+WILzp838q+px/kEBjtNIxFkyc9zDh95xSN51jPK+
fbgNDBg9q6e+mRfIpquqPQaRJXlGRHL07YpopIwpamOxxdxS/c3EjXGLbVsG2HwvfWXNwTvijpmh
d8xvRr3GejT9QTtqNC/tx6KNXQbuMG4Yw7rk93MY7C3Ur+jIs69DaswPIAr46caFcCE7M04Dl+GR
XXDtF89c0El1q3nix2crxmtCKJEOkh9qrlyv67plKGMPz/L7DXtx7YK1iBNpfhVHOyjBKXISM64E
LwDAVFQT+VVuopjPvpTCjwM+m5rYLroL+wAQHeSikUXL27usmHUrgCy6CyBm9dIFGL9ccf3IWgec
EQoN6vS5eLQUqLGfSjTzvVwVhhKijbYfAnkhV8KM3A/q1ZVcER3HJjCKTs7FbWCZnjCa7PJwQLD2
5E6KcGVEOU6QebhjlkH8PUtm22gNWfENerq5svKpUYKMObZxp6K6MPNLdFHkTCvyQyRkd2twnTvg
hM251yYEcJnTcWeorZl2FATvG57NY4HCjsaOm7NhfEWuRf1aM+zl/bbv70cDEN0wIA0R8p6EG7CL
/pBpjBJ0vNKJVlYNKvNKppWqs79EpUB9A293GqnIQEoI6Tgfo0xK68aUZQqR6H2YdR3D99MOyAQj
hcPzMbnBoJR0L8q+aPXdb0TUrJ/28dZJUPxmU8FXAC0GnUHE8G3d/GqmtyH0XdV9VWm7mAdHjf86
MSwsKDm4TXAGVDy9k1zg8KPSVmdHGOpKSWSDzXAgU9TicO8tlN2xSxGMyPFeFCkDQUZHpT/S34Wb
e7WXEr2exOCM6lvZtFkWbgYHcfMLb9GR8lBwe4AAk5VjYEGt/Ez5noeA7CIpIFhpLkAOKRiUGWJi
23RA8jAY/EU6pdmpYu7wcpVeouwpgRjVPts4IfSlt9FKvwgw2QuY09c6HKMqSNCkOYA6Dg92Vw5F
6673tR9T1bpoMOqSSCrTukHwAWgwXIqotClxXEErrLxNXFwRO3/z9eML09uTvQgpgo7oDgj17y/b
eVG0hoLBfhTUKPCweONf/YnR63SG2PRf7BIarHcB62jqV1E6TeuuoERYrWfGrrDOQjOt07orkjF8
AhPePN1zMZ/mEPYG3Ks2c3M0ZP94TOJWwk8QhXdkGIqrxLX+7A9/vqLY0uahezfhS7XFDAUzWhCT
CaIaHAxzOKsPCkRFJZmzE6xT4nG2FBdy7VkBel9FpC7TIrhBkcTC6RBPtAn4wG0FY89lzhWaeD3h
E9MCv+5aYvUXSq3UQ8Wd+IkUZYHSPt7XGYSaqTYBbhw536Ir4aGklg8uVRB3X/iUn9SrkaGXmYnh
At90yhYLJRcOGWWQSOagwrUpyzJlcw4p+UtIps9scy4q8M50bEdRegJjGtPlu2bSdk7ON07+iVCI
eF30pSBeZJLp98GUEX/KFrwx02xmGwL+RWsTeYEByjRYgwoG5SVrNORdikD6MRvrYjToiNz4MTBM
Ioj+O7pMZXQRmqwC3tbpouJ6mEJd8mkfubInOqd20nUqeXjTE26PlL486J6yrXOt8YVfzQZJYwbs
hsu2AstGLBfCa+v6APSXa8immViFXL292jx+G+UOTwdLiUYHNQAesQRwIG3CnJNYGoi3TwFAYKgM
7YIEEDbw37YhpVHP+CGXIN2ltCJgStLoGZ7/d2BsG6ddNVAeZR+9vF9nyKjkYqwjB/HGxo4zq/2W
Dox7ewXlAdeSIIl+ZhmnLqnw5sGHEztFZlNh0rIuZDXh62i8JiYIHbtCnolD+iYZfBYt4dSXs2To
yfct04kVmRL4EqVHZIf/u9jInbwoO55ycapCmhjRkaXGOfl6Bo8iKMQRBSO03Ry+62/JPupprcMq
TTtPTE9pHPx383l9mmMEILG87WvKNP/4inTiCG7n4yxV/3ZMw3TRjhthshFgCv2sDZ8R/icI0RUo
AwHnXFF2NNzpggzbImcILyJaCnwM4opktyH+okomxv8Wj3M0Z7OP6MWYy9vfg/oaO0Qr/StwfUvs
/49phZ3FIH7P/wVtr6XO0andUjdsFA1gvbtT53utxBfDXqQIU3g+S0Ub03hB0b7fd3XUsLGN+knb
GvWCrZt6+EzAT29cDpMlDQLS4l2Oh04BKURdLvNOv5nAZsgSt/E/ktgsRZqv82+7DQVPqxpIiLXM
xui5Zjc030RM60jWiYvddZrUlo8OwKhtMfpvRLFi7qRhV6J6gR1qAZU9IPfaj2LjA0AjYy1GEUFD
Xji8AsFF0pouHgI+kZ0BoKQZg+7cOmUz4wSMKJvGeT4KcvUR7DIN6616WGvt+aD4Khcgx3MMTYqP
wJNfIovRc9dI3B9cuClD8io/qaXy/2XluhRI2UeBB6US5Qc3prdwZmbS34iICb6JsWmOhlpjQIFf
W+Fn0lwZt7WKi3NGRgd6nChODVPVSTKs6CddTXcsuxt8Q4G24BzXz9AeNLxmTduQk1sEUCQ115lC
M3e/ajXilEZWpDfsoUe648w7HORca0dhXzs3tytPCVOmU9rPZsj3MlbL++wceGU04Jo5MwSGhm7M
quyPITwhBjxa1L+tu6FPGPeFDCCZOL8GLEUiU1UCKmUeHCgtWhYH+Z9+UFVMX7b4Pf0Bm8ClpR7F
9lq+2A5/eEt1Ip5Fufc9uS5wo18Ob8U5SsjnrdKkm/iHLgcsx62VINDAr+5srxch8njrWoObOuWd
hRSmLmcxFGVnH8XpWWGsoYZBWd1pmcd4HglNghdRREByC3wWQCIBno4Tphe9mP7d2J6NbakMrZPk
lhvArSw01lq3kvEa4aKtKyAynWCQEUHgG7B6DntjwcQR0lXqfVFAXmlEP3+Q+fhinDzhGSIcqB0m
nj+x8hXpeWTkZpn/IZUc5/kOSN0wtwnasxNtNdzaG4JUunWjsIYtiV91xXrFxJ8pw0qjPY48q3B7
uVnBHk64mwwxROQaAfUQfciyRT5Zrxzgs5ETSl+dndsEudcUh/uWKzPHRHgeBHAMzyJffanQZzcd
uRJKbdabjWN6psaJxNK1xjA+STe/jofsTLzk5Bu/pKwxFuW3BxkUHI7XkVCfrvQn4YAJCb+Oevpx
+r+qqSjADtmB/hrpJjEob3VoFX6969/HxfW9YFSV0h4jGScYGx1WmPlMx6W/6MKC9Ii1hZdaOa8m
bg7DXwKAM+Vlm7CtYObj4V7QsoJR6KjynnAxBvhOeCxiuLJp6RdoTKEgWKANe0e9va948IjmcE3G
5DUA1ylv4RY+dXIRgk8dzCGwGZMIYTN2v0W0w7IyWApGKjJ86UPtPaFSi2JYToyKAx/CXUZZlX5x
0gqO0GEXLM+qmF/a/Ew3tH6Gf+TYdQybqn25HbZaaVRUMQ7yA9Mn7n3aR1lIlddURqaUz8gK6Pfh
rjW3Yit1XOeOLXCU47Koc9Cax3Af4xmyc8z1eHNDSCd+aEuFPjYWRNpyO8EkXTxZLdix/Vf3RQJe
lzyYMpaE2H4rsWLGKYu07nGjM2L2xXsSvjj8VOMTQJivr4ia+9ZEvbrLn0aerkLavnpg+TJnBZIp
WAs4foqD1P1OsjbkDmUxtJQ+5wXXy2Dqdz2NmogvqvZBGmUp5IueNJx07nJUXRIqEFGwAu5XD2mq
+7/sRiOwl3W3pw/HMZrUKUybSiZ9/7e6AfQ/y2AMwEA4WwZd5iom3xUE7xY6/FuOyOVDI6+Bytw8
AdVk0AsIHlXx82jg0TP0U0LqexSM7DpnL7I5IzQy1dG3VyRFQ98SaEUBRbJsgc2p5PNpu9gEIe9g
hA6F/oIeOyDFX61SOL+mnJk58JRPk6UnsKTh19D+3LQasMq/shhGNBIb/aMwDTi9Op3l+2fJ7AuE
ntGIyZFrbhrOyEY2ndfbyeG7mVAatAIJ9cqXx/46y+5UtpVNUFPd8gyOIqUwI0aykW0ignsanvTd
ARSOVm7Fe/sOSt0yHon2LQlNgBuoiiY+9BKmyIzSqCnJYuc1XSZgVsKVojThYb/8FEa4iO2kYaAK
MmobFh7sj+vm4Y6UsNg2VgHT/N9GLaDmMNA4LjE3wLrd3PSws2oj0l8fAE800VYpZXPxJtsBzuSZ
J8lBNin8UPvglJDLEmM05dvFBX5meGZ9+/vkpHOHa7vePLYsPG69ffu9zndyn+qWk2SxAwHZTzrd
OZK9hwZW0hrgYHuykeQ7bhN02uBuTHZQxARWCgDaDIS9J9OQC2UurjwqudKWWoRM9APT8KQuSnqh
vdN3kZ7Nh4rLZeHA6HRR23W88MGP8Btq5SwI0SL2Weo2rB5metOJgiiR/m0eNXOe3SW811IhVQgE
yTfsyuJRqOVhDBJY19SJAi+2sMnEjHqiPT5F/Gzh8mYGInk8bSIqw3Z4aFeUAvcSfFQnXHTQBqJw
50oRlG4RIFdL0oeiMd2scln9WLyJVARIknKgy8JuT53ceAsL1cG0r10DDWuWwBQ3b+9Tc/wJaLKJ
qUxmw1iZim4+lmQoQvUMov1eGregmgCkwFvBBa9FLwSpeTh1Kg1GmLfHe/+DW+znB6ZdabmjQzgp
hLnCzNxhL4EuztYmZHD5jvm6Qq07+TPf5x1/CuSut61BCSll9UIOAi7+8nDmGXZRB2O4dB15FrPv
Sv7vkj8hM7BfF3Lkmb3HvRoe5RbluXqa8BZn3nn0OxckEFDDosO3WzUgwe/fLIJsbswPsQpZFoET
D5t2z8hF8ymSg1cHKmSOtik+X6yF0y090uQ+ouTDGHvFMCYiOQPaELyQjAfWCteGgYsJLGlz/Fnw
LCJAysSDWrZIfkrPlQ5MtCBJ3VQs87p++ok+21QKRM6KjT9sdmdPjb8CJqucxoz1Fn2nKainUc1e
nEsY1ueX/YQ/ar2g8zdl9LLIWo8GW6CGVM/NbXxPvRftzB8t3kB57vGVE0BPco3nJXYO/KI2hzml
UxXyJy45Az4+4CeOqaRHssKBgF5dxa1Q/SRolXKmX5X9+8/FlP4LH1tTOgA8OyC19M7+gWHZcOvA
Ahofk8qiJutA7f6qFrNLu8QpIOUBiXeE+sMasJDIe/LB/S2VAY+POMR/kD23eog6WpqpJbSZm7Rn
WDAlzjw0mLTm1/Km8/+s6+yudsGVGyVF1XWnGJ1ExOykO2Woc9BmU3P2zPm18xZqYSVXwzqFFbPF
YmwIsAFzvTWodefgZXElAoBJbjRyODHG/+tCj4I51pkY55+A9Ldh9SsIlDeuvqi6+7+aTtaPQr9R
EjMO3PR2UztdWyn68IDjhE1CJujm4QZMZQHdRiwpMXyIguNiWMs5ZNd1pc5bCVqh1vJvrUoGr2KM
tmKGkNywpskMG0F4mI/zikjCY0FZdAGbW0C1lhLXnwSN+rvarV5tT8OEjuiFf0gfSp8aYC2BhvSZ
+OXHyOlPJenf4yidqtJ90qsOKe7L4BFVbwKkWn1qHo7vO/F0TfUHqo4Pnv7UKyBPQO4CTCGUdTw/
WdBblQESS3GAKfsHDyayg0A0xbbauAy008vb1ZecZ5H93ASzk5zwMS3/pFrMeg/DJzLpOj235S0r
XK2QZfIwVbgXji2LPXjqx8G2a/DhXNdkomCEN+fgqsJxPKpr6ZWhbGzbtpnubxz0ncBRi/eneJKS
4ec+TQ+dr2W/VwSqzZgVyCZKdJBS5wUeLHbQh+JSiOd3GXnD7NXCau2GsB5S/waXOjK6ip9PqNdQ
nfNGawbV+Bwbc+uRvYhKxGdjyWT/V+u7feSdrSK1pxBweDdczDCs/x/jA+hpkPXLBKR0Uu+EVxD+
fDryR2n+m3+QKy06OxTlL/EMsY9yPeUlXOHUDyNPgTj8BoNLoTIHTGRtYfRtpX4chH/icrNZJUvf
XFXQTkq8fW0fa9mqxjztSbaffdMTmTMeMECTwE4h85p9qyw1fnLTDcyJpk8cS5ARMqNMb9y7PbLN
oqSEIo144gEmbrAhWMn8uey2brDBfFPCVBjC8sknrpkoE9LIDXV/M33vkD2c4FdZlXcymcSPLqSQ
sO6s85W+fhS2Oj1A0rPTlp+SF/QLuGSUvi7KbBOKuRUxNJ+mOCw17yLyNechpXkbNL4eRJy6rpqM
Fu70v8Xs6hHfl15vYNzKtmF+9+OSvmwXa1iQ0zazctNUlbDDkjyvljVraKg7z520trLWyaiEXFCE
NPzTmFBXz081dsQnfQ7z/HNm9DWVwxIKXVnHISsSp5DFOCSNxogOH/H3bQeag+P+30Adxg6S8Tr4
F6U2GfWyqCYE2MlZJQKW6W2YrmkUJZTtSoYXVoZuF+6kaCCAjcqIZcMBqXaRFBNxnc4ZcqZbixN5
u/WWvRG3gNV4b3uMq0f4xc1rW46hLQ3cMIc7zgqLaFk0EMx2D8h6vLRXH5asem+9CfLWF6/Kfyy9
XHqtXq8ep6IgdaMfQaYDVVfCfl95VUUgueXA26QODlESYGrS3XNYHU1twD2dXQODseoyFj0jgCkZ
9EOrbBU10YR1JxLTRjxWpxweQcrMZcB9nQ27JVa5GkWFQHDtw/1692CVdUNO1vXd67ZU71FMy8tz
RrfJt8a3xYpL2x3jzIBUhJhE9iyZhs1BROsGikBGA/t5BpzEdfXlH0LHjw9Hl19LVB3vKkXSJzLx
5kHSOd06lzvdFgyuGKQej8RhIc4HQz/n1oZzuMyOcmzE7up1AHEI/qCHdCFQ+qx2IsePRt20nJLJ
ucbDxSMVE88uJN7EmNh0/S6JL3F+cSW1/iPwVjUNpqbT1Me1ofHBMR+4fvO8xQt2htglbYSvnl6d
0Evv3qkZbqRyCzgG0iMV8BNRHlxuAHL9hTHIheFpIa7DIiURt9MZKV+8SM9HTecbcYRIm9WHE6Q/
E+bIdRvMR8cUgquQGk8RkJomoRBA5cZlF0aPGOC1opVtAXMlJO7xijSfHNrXUb5DmSPOJBrbTPi1
O/R3ntU81DopLW4udTbxS84qevPpoWbqRz0/IAkQ0dOi2mbFjFvxXwji5qhjiZ0ujiBECYdKiAsC
da9wcDYZsxujmf5h6DrKY2rhxFzKK5Dnl428a1TD10Tu9+vbINt0+MV4Z7E3FqhkeSQG1DOy7WAv
L8Q5wIRcbZvW4yvuVk/33QGMZ2rLvKoFHVfSTUCLNS542DEfhfc8watz4sh+/5/QioMK2I7Er/Tp
4fR4juOsmEwABW3f011NxNbLT2DEUSmTagapMml4w/TFFx1wiQQkb2Ha+5pxYSYIqICqbg01BfBe
aOnlbTLYaFzpuqwF3iv9azC19gNiPGcCIC0Yk6UO1i64WpVqoksY3l7ECCPAivfeY7Ze/ktOLHty
PEmAO3NyPSN4TU5z0AFL7XsIgSavlR+4a2XJ78MZAlmFE+DuRxxlghnoRyfU0AMjgn7kgXaoeZAW
KoGMaUZwPES3JA+iqU76o80Yhp8xdyMIIUKW6qQAn9aDSzubYvpZCbjH535xY3f94M9TKiEme1Ku
UbdaPddecL0UGL3UCk8FhkenXk6vFZLdc7VIbUOf9i0s1mrdQy9F0tg3ly7jLCWRnZeEOyemVMgt
QIc3crvT+PUqzXELiXtfOWt3UtT+uAyuPv2BB1TnXyJL9lOOkk4h5PWrAlTqG2dsbNp21veRJ55B
/IW5q12FbAcmv1jhPyTOH8qrVNCUDpAk0tde0TADgfPWCA0zv5+uuNdkug4j2xlIT9mnhJtdR8qt
oTtg4BGj0OQFEzjpV7Y0TXU/PjvZyfvKyr0YfTpALtkEfcFUZxDW3E2M9Nu3BWJ/nAv2P6wN0a8m
KOsGojhUdmupgF3t94JKT6Df9RVFIUmVZFLCk01UmZYMJ/jYXp1U9EjVpJ0GD1g77VvFSpLliLbl
U4dxwYo9MmgPerHrFJZr313ARoucJGMezD3S766wF1NRuJt2bVqrL2/MoFGfXT5futOogn8cy0NU
f1I8JPxVUpOC4AYFr27l4dJ6eNjEhQyvS4Zc0Gx0YNuTI7woJA2F670cqWeMqixU4LN0hpyTEifM
/Dp3uuI5qHMWAckgqlcxM+SDacOSJzKgo1lZMsLwYS5K3amFoW682yIJ/RKN4J06UiYD9/QwUie/
e4e9x6zzZVr9Iik9caJOVlaepA3H1KPfDwZ7uoelqddn0JYlOaanHiZ9mBe2kZxOajFTJKLnxbYf
qZLKLb6yD7K4ufKoymOU35VE7aDRWgsFD6lnkV8EvpkbBHh2ydrUu619pwbBnhjdw5d6zp4Yk68M
zT6KReIBZshBwXROEfW/oU7Lq90VYqWThap0L50qkQdQUb4Qfnh1FRMTgD9rNU2Y5VMZ24/Xj/Fv
UM7qRbnLSWEnEs25QdscWEsLEfmEvBCH6IQb8GHpvmI/c9+r9QgSGXpuI1Qu7hKc2XqcHNb1YiIj
8NcSdEjDrQT8e0D93o7bWk1vXlVviSX/AyasG41e03LpZ37i+tWeasKWyXwenvG83dBveI5g24Bx
ch41a4ZlkmB08RZKNVBq3EbExZPxhExm6Hv3CuI+LudZ52N/oLWn/HvswUxO+9ZkXK+nvnQz4Sqt
t1rUHnTex7Z8UHJTzSVtDLz41PHOp7HrdtadAVeuj1fOsHE5CcjUpTnzigveNHKpw2K+NQdbx7ro
MrcIr5K8azPplzifpsWbIzBLm+O8Bkw/v0PWwfNR0xlnq3BSZq5+UnZdUF1BpFgJ+ciCi3xVEMqP
Xo9CXeswPDSUJEtxAfTwn1pSKGEWhdQX5vj+OixJnRC7jQWi4IHwN49Wo3OzYlKG27UVjzjHVWT4
vSenZJwdG/0/NpTd7VXZcfc0nYOhTQxfBibXLM1Tvvd6L4xefh1u3SxAX7FyNYcBUHSO86C6NYTS
q6HUcDMyyU1J2E0emh1xEUGjrHQp/nF/FG/EuL9iSkXM3yedqgZtdTH3/6lO5cbIoABpP4EtExe3
/LHemqLPRNV2RhjNFJxBNyoEkcnxxbcXjyvXXcRWXXpAEkiKhlVfhUtZv249oYeXEDJQuDPnY2CF
BDua8NmzGgY+c0lvicYXI2ZTxkV+EzVPamaA7riFDiBq54DVOnBW7JFa+C4s9SoG+evWFHFJ7ay/
Gs/O6tg74b/eA5XrJ7e22o+bnsaUe1N/T3PO1pWLeuSQV50MXlpa0y1D/5+fGRWv6H9orPD7Bo1Y
1gcznUqv1zFGxIZ6aud6qPkztZ1Ntg9A0gom/3tlsBPmKtOAz7m90X1Lk4CKk+qFUKB+y7YXIMUe
lsETHT2blONDlEgo6vvL0KmA3YfZpL/2DUp+aSBk52AvTz6Xi7s0KYNa9baqVAXHiskvOF2dbQHQ
80VIDFYYp74MMmiqd9lyMWxBbBqD2jXZhXIN9oiibObPxFjrf6oU/wJd0Ac9Pw1sGcJZAVLx6giH
q55i2XEhKIU9baDkAeG6dkQ2SyXxCcF0mmxn2+1Vs408Qz2xiRz0Glazk1R8CQpg5dXSIYB/aDPh
tWuY35gpG1vW50nMw33jwIg0ngF6229fC/TFdx8Djl110NPV5VePS6cPkhWb3nUd5juY3WV57QTc
dr+DlxQajp6VxxbYqUFmtdX2SJCn+BJG+yXUzYrOb19a4nL0TVqGfU+QbkFmBdIxc/hD8M8gn/Df
mkAWAfl1rIUrZRuhIe5YP/+jOGRjXSWBUmEqXu2IdoYedoR7kMf5jtTyg7tIDYtrO2XXbmOULEQj
TgpJx5lxDibBT5a6opUB90/dR/pOuV7XRK1NpVwi2wZfyWvaoc7YUEysNOpBks60BuYpfDwdsd7r
d3XStk4yQqXBtOeicugPKliytb1IUZKF5t4FqE2JxO287uz0T1bp3le4ff1ypfx2SRg+6FK5+UJJ
9MYV0yj2csxKgG2M6g5+QoEL8Sreytltj7sT3CHnrhjznk9b9ZNGk7HIvMOu7ESrjCoL7FlfqsEM
9I1nIgzgzMKFqbck4rA/oWh/yrCh43EjpuDKYMB8jCuPpmKxX63Pq2jtQwVEAMCzN1SWT7EmN0Th
sild+Ftlx4h+CNYe3ANq0coPLIzD661VilM2gT1dwNTayybdkyZNv5WRLE39E8SeUmwU+AMn5HQj
B0UCs8CtQ6ox66KX9zwogE6Ksqf9AFZ1hN5iL+xFbgvPQW+KujYKd7J7EP9FarpnxiI4v0f/yGsT
LxWK7+F275ubqU4pudyUSTIUBHICbidyMZW+ui6gMlQBqiPQ3TeEmNn/MmRDFRgz3Zo8bQeIfav9
prBIII66H2d8Afj/pbT78ni8sEG894Ee8QycJexZF957LSlxknjvHS/ladDL985pnwl1ld8PsucC
VV6dqjAGUO9XBFkAh9QJ4oWZsXhH744WrNHBVqYJl8BYinP+oaEpyqnvwsJb12KzZszXA9PBx0lD
j/IjGp/OWj4QOmdOCWAcNBkFQ9Xu/xxXU+bx0Ec0ctGIgzlrz+GkHsjGNHe08HBAOfDSlEaqYOOD
9VVmZDRWxuyfxRVkjEwqC95FRjytiYrU4HnoKqDxXva9EJL36WTlKud5oSms/2S1+GZJwYwMLEVM
zDsjyQB32gIDTabIyzcCDGMdP/6dKB9O9418uP5eMbmD0/Uw4mfJXNosHX76L9zHtOLTVtcXUefP
+MaYQPH1agvow3+JDDLU5aPPJPnKz/uWzkbmaXqHHtct9JtR3H1A6FaiMuGviVRJxPu6huJZ/VIb
a7voarjAaZx8HzK5eIZ4T5lZ0Xam6fuekznAxKQqepzskW/cebMBl1A7fHi3XFxROUHfZLYRChWv
UAy8ZIOjsm5NFJhNpgYIe4hfqpdo0fbfT1Hq5x64T2EVV49M9/CWV9muRyCW4eo2OjNXDbA9Wkln
v0n+lmcePVDcnwkgkAUYu5dQ1OIOrBiAY9RK2ylEs7ZOS+HHJ6U+wgiAzVuN+buhRo9Z3qoHOJsN
eW9GsX380zArIhwGu5Smg+Hg3oTRv0mzIaTX2Qtsh8hXJnFJ2nkPRCIr2DKcGoteLGUp3iK1CxzN
aFBoZLAeFl7fkbMUmVw3GfU6nvMbZwtNEUc/yH5rmbGM2EVwfWC3SB+hx2x6TL5jQrjjhr+mpHtu
Jx0BHV+BaVEXKuVSMH1/9V2RI0q/4mYNdhOySxdnZd2gQkpQQHdLj0XWtGDBwTi9xK1tLTS4AAWK
v442Qqk2FgE3sV3Ufjbdc0pTpVood7gj2F9qr0gY9eeEt9rioG7qYNxWcKOyORV1Kw/175+3/OvR
w088Fy5cQqojbqsHnKeA8o+TKhDO1fM4e6a7RsoR9r6H3blhQvgm9CDnd7Bn7n7ucNgZELqHsGu+
LzlGmE880eXNAJxTu9eiNgKoLO6L8tRdoIqozKdbToWJ2d6w7IP/KMlFqrfnpuKDU4W+l3KnXnSM
/9DECsg8D09IMs6GkKv2erGXdZkSu4+Ul7G2hrhfg8JvbV+omoBiwasj4JzQot7f3HbamO4f8tlT
FCow3CibjBp9Lowa8+IPnFNkOCJ31LNesUyDvkyiC2Uo7pSWDgqeA4Z2+bY3bP/+OSZzSY19mGDx
hhS1SjBk4P+6Hev/bvpek5GvULkyiTpePnggLdZu8yNr6yeKREVDDQRoxHresG0q/q5zgbenWY9x
5myl6hAWSjQKK15d8HuCW3CSXiJxP6jfww40f4EswFh9OTilP84XDdjGqw2oQBKAIF6z/0XosH15
tsLDjNLIXpqRTuJppXmMh+tW3JtKdtFHDkbNb/5S984n3V7bybmIO68bAFjt+UHiLwTxTpXuNFqn
RU/8IEKUxUCVGzbipiFUkgK8LFTlZPvZkO1fpM8zIXFkECnhk9Qre77KvmdpCAjvIsamStRZnamW
vBVNDgRhlC9TQHWovwl32TqFKrTBNkW5TGLChawzUWSQluX5e41bMfHUd+ILkJj2rmCMI8U6Ctb6
fEddD9P5wquSGjSsZ3iuTGrG4Ts7W9S6JblygH8L7K/wd4Ym4HWkR7mxv/Wr/0v8zXwejYB7bPGn
n6KejJSU3OthemBsOPCyLzszf1q1b6EeNe/xlgAyz5LRwF2X/ALdhP/C8Vvlmfau1Z9LbT4oM9mI
ZKeqJGs8QK9vuiZZCJHXJCIbcyvujkw2MyzgG/V5M8BLbL29/2BFykj6aWPAgaEq1a+OQljLY5Tg
DG0ZDAcsrbucrsORaxZPFzcohHEs598MTKZTKPCs6X4i48hFaZizSljniojNfQGhATHuJ+ywETzu
mT74OuXUF3N5WmubQ7Gm2Hnlz0gOX9MHvUUYXkJ/1T8a/dQ36dKcblfQcjF+DuTxWvucZMM5yXma
qfqmIzIhs+O24z2x16vqaSzGI1lU3oX1qH4n9oQn0TWxfYmC3/+TJY3gsFY7eJs1HNMLTsrT6e6F
QfU+po0vGwX4sBo2h4/WB1qb0h8b1R7J6kOTxZkkaC7aQ+oNkCQjwX7ho9HscEShbmtMrh/3jqMc
pP9gOj7J0ETsQgr9vTNITp0WR8Ldm7UWxuWgf5+8KbLs/JBtHskdhl+NCM5R5DZPufqDo3HBgVM1
fss/eFKjMz2CrJzbcWImMSjy3UseOxi+f9KwFwQeljGznaQ8iGpaDMsYdAC8UF/M8jSR7nV/Bj+A
SNht9km/cxPFPb955HZOdF6+tUwftWi9d7ojzexEhZ/lWIeDdts5rJ5TytQE8mxJEq6yqXnhyMpG
1AxeDj4rXQHz2aZJMcLPBEdHl0u8RdLGKaLGGpk9hoSpMGZaFllyu5wh0o55IE5oiwHR+KIXi/iM
Ce7MhFiPIkFWb5iS1VCKN1OYtyeGofZ90jKwsS3Hdr/oMMKgr8hQoE5Y3cqSldXYbtu1ZUICTTut
SWtviKb7z0G/IyshByX2AKLHtemHPkME9gqij8zf+F9B/TUAq77cggRhv5Dv5NmBCbEY244L3fUo
2ZHGxfLhFYoGGebcrBedJeoV0GUInigVBFYB0Dt/7j3rgqxm7nXLkR0U4sJqowSpU9Bviru3VUL2
V7uqFjxUPjhbTcJCuJmFSeLXPQqGbqEzBdcmT2vOP39R9h+2T/urvaLMntEaE4GEpLBH+GikQcTN
KfYsr2Bz5eP4HQEOUxz/GFsNfcCaagM1HmAoLuBaoHS7s+G/qyXvLta9r+atHiaY290j6mn17/DO
oLOSP5KGxhDiEvtiROvo6qmO8o3z+XrZdBToSQj6qdxVeBDBn/cECMre/7GjN5hHZsgCw+tyIa/r
GboNcPhfrXOLcvsuXci1FHX1+2RvIuJSXYFFjaSfDg1TGc9mANcZZ7HgyIZgoeErva8Npu839fKY
nN1OhUkFPm8bLZKMPdwvnZtwglqjdELwUyZ5S/D2NTd34GXrty0IXgZGDYPbQyM7usquUfFrOX6p
FRAIRMwiMTkXknxmN6bLjFXujHTDvG6y3/XrooqnhOSMxXInlBNNB54IdwQ++VTVYmA8mDwPcI5d
2Yp02qCOmDYbS216GeeKznmMneBXazyBwMGG2XapaM9J29MgoYXeJV9bbriz59KGJW/UElGpDcqD
a6QTKodbKETtTo2XD0NZ/Yxsf14Xj+zD+ixnb4OC5uqHmUtKY1h5y+tqS1j/6DTqCWqoI9+w8FRb
/WW3Pw9kYaUREC79YRH4QyccvLOha6SKQCPumeKI8ZXPB4AqYESu7zzMWaHzhHruhy2vx+5Lreob
x4qlwnJxenlmtxX9HQ+eVgCfy6uLnvgDzuxC7FsQGAAXTPM5s4snJh+NG2YkQVvwtqN8XaEXtM37
qlehHl0G3Qxmqj41vSBg4/RTb6wUQgsBI4neO2QEdW7U/Ji4pU5kNDS6mZukNETj2xrgRLh/KDGS
2oJiXExmpfjUpNJi+L2m6NKRxLMuodRilrrVb//tfvBcJvLC1Dn/Mvda/BgZLNGVWOKn7d8Ai6jm
TJKE9igx4hWqK9I+OqaXZsCEUTp2NjzglQgrfwNBvnDC3b7MOyJ2wpvpfL/tbCtI3JpLBPKe+iG6
fUYma6W63xs69hR4RJ/bjyDy62hhc0kswNxjmv7IY9jcRLnDXX5IIHhmoOfZkEQSS6/7RiOPF6Uf
YbrTxkEgVPHVmB5Je6+s/N85j3kOiyPW86e81DeKQFgW1BvW74Dw8sq3jgQPXwlQwevmgo84uz5h
6OKc4Qj7uiqxY1WRgNESeypomTaiVeI4iXRocH2eZR31A+wO+Ae7qMJ/ZB2ShevywjQEKm9mJvuT
5usQvv9X+G0fl8SozMPBJ9vOcpIuhz6GTsXTBUZ/XSLD/mDb2rrFN2+GoDiNuvoz/Hi/prll4GqI
X6qd+5ewKmRKRTUeKa6+OXwDrJQTILmZQW1sg04Qreezx66pHr7D4Zohmb0tGVZRlx/1t9ObIq/H
pawg00tX24E/3nJ2lT0AVHNSF7dDeu1QtFrfv8I4CjDbWd0kKGm5iISstDDWwI5vXVqrYPcCw+wH
5k2hAPXSLOnI9m9knNuZ+MP/i/P1qHyljfxk+4rI3qXfI0QMtU3n7ecp36vRpUtZ0vaFih/n63W3
h1uH6Piy97i+qHn7NvF/z9NcETFoZDDKevvBF32VIrhTmhBNzZFpsZQKxBRElR2mpwwvvWYlxziV
XqCP/sCB0FD74NrEmnvwi9fsLzF/RPVktq4uzEBv3m64zlouXWBn07mV8J8r+EWqfZkWb5nGq2mE
jNZCBafGf2ij4UOJjS2VwB7ty68zdcKc5VZ8h/v+VuD7xm+vM87j8pb9ntV2LpEqVmzpac5Vi8S0
uu3znKyvBiBD7Lye9qh1kKKDxPjFgF2pxLQmqCKPP2Nio+Gqux9J7/TrKtfMQnyRYghJURnUmRXR
jkjB5tgq2dUh7KD7IAyhmmCkXa2a0c7RbZWk7+BJdkRkLOl90L4hxowjN2wjFeDNUkBx4R/LmwGm
IJJh0s9l9yJBYYJ3BVPqllMe/8Ez0SeZgaGf10Pv5IUj/r/KYfeLTFCsOaIw1DRJknqzbBWO6llv
h6i8GIrhCDk1BLInsa+t0oIJW5jyoeR4ZMKZIso2WytSQo6uBghCqy88M1NDOf48eCeoJLsWdbzP
guRmBK/BGApk0OaPlDTuvV90hF3LXyoLsgjT3f9DbE8BFl2Pmss8YLSil63BItSCW6+BVlcHHrvN
LCIc408RE+YSxd/rDGvA2LeEqQPpLd3/4wxMxHhAcEfXhxHOBR7QWT9u6QE37Fq128PDlIKeQVFM
4JAG71ge7HBQlIE971+GQNfq5NdAoOYm2Qsr6ml7ptWHTr5btuSDBk0iz8mvgeD7E8JjlPCvDyYn
9s1bTSQGn/ndssIjznrfMSxAInOtoFYtxWlupStkPZ3hdA3pvOoxyPbne2RhW0v/qrwnWD0ng9Bc
e2apWlQk6grfMMS0UZRmn5rFb4ux6heV1fv7mNCAWqYoQCkRSgfvyOBn3NQ6gF9ZImx/zL8jQ4Hj
6g5BKvGtjBvp5i1+BiFQVGcFKaMYFRo99dstCmFQ3aeiChAar+5Pofk3gafSQbMx+a1em528GlfO
3OYkTqsCtXvhEgRbhUeFZOkQIfkoAcYttp9lVXz/3sC6GIqf4dUl5u/9MFRCCyqV7JcPhXwQGakX
4At/ZeqRR/IEJe/TDppKXwz+Br+yAj5SvLZusqKp0pNSUS/K262yZ3lGy9S8ftfYDpCwfeQcvC8d
Nt21PU+XoCsZV/EoYRh3VnC65MmuPrbo2b9nE0c0nhpSm1gLEDe8OI/72WeOn8hcNiooqV2qokpZ
2BtyOSS0APWs7XzF3c56pVqKAchcDFIbXCQ0cv+DFm8MUDm5KFOg4dXjdBC6WACusLEx+sd/bpgQ
wIeB04hzxTyoxFvPu7Mla8fHFCi1worzx/ASoQutnaM8M24FQJqkRkddIkWKIn6oNS6/+s50GK8j
e2Hrt7x7FEIdNptpE4StVZRc7P9qKekADxvfBcHIh50/Qc6l7S6wdM2QlPEvC8weF6eTKEEFMq4b
9Lr7IUJG6SH4rz6MwRRksEFWbPraV5PqD3bryGDNvUe/4F7XvenOjcmdUR7VL4BQ+fieZGveUZfn
CyM3UePRrCTG+X6Fdc180c5y9fphJR61Im5mNPeap6Hr25mYEI17gMMGN2OCD2/UJngqlYRQLTRM
8P0amCbM10Y4AflEE2HY5d9p2ABYJuAWlAI7ffIhcyZjnit3TCZHY4SlMoOfBomvpsZ/Fc0H28tK
w/hHB9LaNN8oXxtQBsAMFK/sz5EYjN8dS38pjepcYaRj8l1/NNopH5H7rR8ZDrnk2gHlBzoSaOqb
YUSwYv+FVDN0zQyim50ihdNqK4Ien3V61Yg7Q5goKN/8Bcp/wHUtcZUMdLyyyCMldFc933ZV9Btj
lC3HGKCZwmdO43PxecDY3Bz7KW7r9lx6f31a4tsgnFJWXN169HAj3LCHraXUsFoRxMbGiIgf/QYa
DfB2vQPUYjckjNXNLvvLoXGVdSbrG6bPRATSrYnAMxNgEVuQP3K99EaYJ9rCjdRW8KYzAtlRyULm
x4EdDUMNyZd1GwbgE6AJ2Dzf1/j/TVi0F+GOMlrdqzfaQFadvsoeZuyUeQ7M5QZ1Mjz4BRHO6/v0
qIOUa8uymyXIiMlwFWQ84blywKd1HWaSnXu1JGJsfY/MjTptW3DMnmizhn9RzccdVtenbx1iNddz
piOnwl0HAihy1PQtBBAN3uUtdevWoqAvowlkJlVGxWxR48N3mk20vVTsacD93JMBB1jkIzfcsZKl
acD6m2FQrWdLCP4FPGAwe53vrKGR9FYcCPT6giuGejGHDbDBJg9K7mp9Qr+ub6z5sA/5Pft8q6im
U8yZe8N/dyukiuLKUZFpsRZgO3ILuB/8zsgPxR5eoV/hJRgZdZRgwq2bT+zxTnLwbeBMCrGc72Sz
1TTUS47+oDSJNXnU0lVn1hXMW4Se0iaqTMx3kNPAHNG31zG0X9gofjdzNYgByaRlx+GE19Yg2DP9
+rxBlhLJlDVieOVAA8brxNhgCDqMv4JRL5F8Eit449hGwFm3YxgmjeMd6IbyuGTk1Gc+bjb02yy1
sKkmjZZauf2o9zCWMX7lQCRoyEIsoWlyZQBz/+Sa6c6/ABKRXShypIJPLcJU3Gc5LwXfNDXrdMrk
LS6VS8ksaZNQQRTjeus/VxPTbSMbKiw1u/61sfThDBfxVkDT+jgL1DpzQsen86hiM3Eo35x0wZ2I
f90Y3WXb5G5Wmbm0HSdwsT73U87fC0JjwsEbvXEAyJJs3m4TkmueI6eAEgj8XYH6JJQN8pJxDzJA
pB1fVti9oIOncgEZ/ahF2+PBD/HjDT0aat2UOMEf6p1A+iYqK2SOJC2zTRXk2Z0rIQQGWD/Ii7Hb
qWUZsU7jwGJPY4Fs/DuYJy3PU+uQqserFHy3QfDt+G4C5RSTEuIc/YexNsPqROUbiPLvigaTXbZP
J1tca2kLN7msD4j9ucby9v70p2RMh256RMZZf7mNkLb+1VnNMdCaAkekrVz8uAFBuwm8C6o8nitz
owZRIwpzUwzje9idARUqxJ0cs9+N2tviAlcvEylGF196nhhE1VUuL0/60gIml73MOVUxM1qzgue9
irsS+b5SNRzlxKoDid+w9uw/gC16VbZQUaMDtCAAQMZL+kVJK3pNOdbaZRBVh8kyAiDF2aKcQwI2
Q7AIOA8nQ/pGRYPS8j0sOqSulkT9IVVJ+MexepwV4EnLN5vXoNkiq2lB7TJR8zqCWFhlAVgisVsG
ZkLFpGDfP2QffCkKXiyIROOUHZT1uVP7cwTA9Itti4vCfKhQ66vsnXN/7Yx7X4aowP/u3ntS6TNF
nOafpDt+q4yinWQ9VdPb/6rlfO/fGVQ5t2z55E+xf3cj6SaemlYjJQrVwVws5GUAKW8dV4m0U3a6
aIdeBUvaUoBgFROfSA3JcLHZ9IXguw6n1owK7CQGfOdgFIOqAn2MaP4BgKAFx9CPjubSLlKHg21Y
dy05l5Pn1eaarvnjW+HuXRUp48j9jp74RyoLd8hGaconRBu6/sHugLxH+PE04u7sR9r6N0Xc792e
UVxShTK2JIgB4ZL4lOvRCs4utoUSZ7mnHfCKRIoTfX+p2/6MBPakj3btMeOraBazeN9gR4Qus3lV
ymDvBkTO1KViTZq7wDSQZYpSMaKPGKorMWk1IUDCOpZMvMrhB7RNO2dAHNxlebke8rs3mzeqExpW
OdEYjGGEoZsXhCaw/bGAaNYtAVBB/0u/vaaOaWAvrPqkCrnYARL1vp5w5H6DHAfNMGeozYkDtmSR
ees8WowigQ5Ptg4Z3zTaxIE41dsMevN84gRisbTBWWtn7az+6cc5kaNOXvXJm5vIP6mjP9YW7Kix
NGZZiBQdTyyo1BxOq5mBB+hBg1GNaDugzkhzFSY8n1bKy7DEbuIiHlVdKYp+7LTYS/lgOcO9v1jj
6EtOysoMqjKggLwg7WXRTtWdTh1IycYpa/+jdN1hUAYjt/CMlZ7Z26IdiRXRNu0FTkcCiIAPD/Ss
Cpp+Xhg+kTcVlw+xjXyFtvcHK6/C5j5M7jekqhnMZlp85R08W5AatACeAfwKVd8+jgG12A5F4diQ
0BUUBXRVQg4YY32BQtffVv0GO/H3VjYXarW+sBiaWnhOAKvXJd7QxDvvCiAFIvUc/383FmC8YjbD
aw8N+8TObLpHh68pN5F8nbKXvxIElwPRV27rHJc1OuA//yb9IVdghqSar2YPSp0QeWikzdSjoyBK
7JvqjdGG+4Xe4qQXxvsxr1VZM/UJcsgH1c+wnxzobyU2lgzbRXFaECqLfwOKxwebrVnzJvp3+z0U
WwcnLqivOuo4gUTC4Oi4TBexefI6uBUAaKmHVAlk/jECWx4j0MZhjCK7+4iZFl9fiW+A13VKOySa
6gEBwagmyEkfvKDiMy4hftPFSiDcLJKr5IzjFSeSdeXIMCW2V8MAxplUdd95XsFvHtfh5QiVS+9v
8g8tJhikA1GWb2B/vJ8yBOXlmqmytRINzoNRNaXzdpGK0GlMjoFNgENQaTyYgEJLO4GeSZHAVVdt
7XiTVl30dWign6l/n2LYopcRTGVENc18qiPpFd6H6U5RkJq4ZZYQ2Ek/AsH4qCfD95IseoiJwizz
cZEyCbGF8I4kllhImyoFvPLjGsCEjeA2gZRMEY1tXQ9GVQdTvLFjl1NkuNMcHEKwLJY+fMq7VLWs
blwNBPsXB5QNv6K6Fdn9KDpXof1uvM117RYy6hf5mDXmR3hM2STLbEAtbyZBzdDQae5VtSxnbgsW
1YBb6gsRUM1CMHLpiwuhQ7nWg31q5f1SWYWJ3b8JDWhulY141efgDUaIOqChCjJrqm2XYy4s0ct+
4u4NM+WHFyltMXtsPEwr/tbSgOK1/VWtORJcApaiDimZovqsRRaLPXT/CIe96SNoh8GJCjXL7eZX
V3wjlshMoPRt1ajolu1D+rpxNMBJO9Xvl1SbJ4K4FV4R0ajiC17DVpSGaMBxLXqBEHGDGlsdH+hn
fy20RDNFaebbGxohIvJF5Tuh6lD6+t6/CwX6KbmW6+bHqqE/nzNbh3Y1Da443+vFoXMZy4ZtUwHT
C5oL9nyzoh1ytAqZVxOHcdMHGNmBP5AksH9W0bbntlX/fNHu+NqfQsNVXEOWfaKqhQKWlE7euP5D
/kdDZfDRMw7ZyXNYjzWVCfSQq1hAfiDV2dTojdTb0rF0Hr91dHFLLC4SGPXg/NX+FQCzyeCdK5Q6
UUnyfGXmXbdd1i1+rKJTNje5WoewGVaCFskjyGNi/e6Wb8piE2ZrCwO/AgUQ9uAzndFkTb8Y/84C
D3xDOl4C1mCZ8tYJhkxeveW1rXOxodB5tF2Sj9PcV8zB8So/0RKYblr/WSewEXhJf97X3XaIkpNY
YmQW7D6Dugej8TKWBrUyfgXs/jhHvQb4p1jJnKnXM34WD8GMYLRdjEByW0FB0SNIbHBw7DbMJUoB
aLDkpwzOmN5z+/JfIgeOARFIHXBMZVi0Z0/GZZr+6ovT2FamOkkxIO4vsGhOfP5SI9EEOdLYyMt5
J3gVmIzoghlEGqO9EQzxvPDkvhj6mzGS1uyQ0eAovbKPc+lRWnu2B7FybBI2OYx2Ig+R0KSaI5cu
+3C4FCe3vhD/PeCexOs2NsiqhpRkZpFiFPl7Q1CJMh2Emu6H4n5/jGND0h5N0rE+74yI52yrLLV+
6eyewz7j77tloc+T0yFNam0bHdo1Z94YwHmfPXFIl36MXJ47wG8Yyy4VcrLesNuPHZ/3T7mUCTly
hFF66V89OJlfaOwaYt3Ei+w8AxzhGnYD6T+axcFWdedaTf+7h3XnXnDA7ErLohCGc2xUkXkziDKA
FiA+MsO+26xtpCIoI8ssbMLJi778EK9Ik3R7938OjV23IYCr+IXLd/qbyfDudPXn2lL92SLOI7uQ
9ziYjNjjnFmsuNxLzuUUtg0gAZi9McWqbC6HM/9voMYuR5CdOSZ+MCJHFybsiflEXzqHYJ+OXsKY
nddiynPeIyfL/KOiX2ALjwXR9RQlqq38xUU7HA1rgYXg44hITj4K4droH5Wfug50Y2GFHGQIeScO
dsr4tK527eVCSae513XYBqZpQFSic/NPekXqxWIY4UMSXmyelv49jCCaegbVVaxx7JAofUCZxwa9
3qsgexSsnNT8Or+RO+umGZa8Cg620WdE5DAEAqR92rwSiqTSHJOp/W9W04fwIK6h4R5J95wm2IPi
yH17NdY1xt35wez6dun1TCCbVilXOBgSdAUnArcNSrKgbLcRurfOSzLOWU6/LaHqI+xgaOquueXs
kmj6TnHog6olH+TeSINGk9ZIafkSLNt6VOfEHK8yf2R14qwp+ytoR58BKuIYVdefTjMHWv0dWPWM
zLx90uk9GiU8BOHy5m5sxmfjNND3P33aS2hM8pGzoICc4SzwE/KQ0/iAypbTGS8Npix291YeC//Y
hquYHU0DleibzazFRXFcO0MoI8ORu52gw+Cfq6Eixrd29qlTTcUS5U8qJzbPE9O/vs9U4k1tBTOI
5bwiD29/kBNLAOa1aAKWolYnErbTv/a8u4xNsOHVZ4iEMae8wF4nY5zFS9WHTKkR864Fsa+GBWFc
jaclHphymFU+h4jZQLJlXrGjh3eq4E7DBSEjHYuZudfO4cmgu+m/d01VzZ2OnGICCnthld9zAwki
+WllKZQOX+MqE4M759CkahkrPLIIw0VhAP7SLQAmnV4iv5NSscIpKIpLGVpNHynty1RgXf56hDIP
4bqUSaRjoXtcG5toX7Sy8IWlBMM66nnfgSi3eOmQUQyRGFYJVaV2k74m6jK/cxxZ+SFPWiD/84/G
Bvx5tOBPR7eUZ81nqdAMkSp0hGiaiOQKFf9g0GXtY2HABOru7DDps6tgApmezM31TnBKMpUhOLVx
ysMmWr3oB4+IaY2zX/al1enGhl1Q6mSYhi2mGdfh254f+ijnerZ6aOuRcU1QxS8GHXQKuIHTmj2m
UPh0Hz8EX591J65Kw9YCQDn3NhqvXeFdJpOVevv2ic1KII7cSsF8PzaGQ/jWUNcpOo27yjaKU5E8
xwLBXruSs+exQwDgUIWjsEKXnVrKmXwCCU/1n7485k2aOL773MwUyMUNI4LRucozD8fUoG2bThHb
7reSAw5ERR9ishXBtbuoef72LEZdKMCQ8xAI92zECBaJAEmYMiFjicVBxaz3/FweeccZhcyLRaIG
t9sJ7VYhrhwdEuzMcsezjwsUKSX7pKTXAuvRjG//Mrr6226BFsGHWxTJYdrhMBzMxa/38TnYlZsT
togfkXOkOl1qHJgRe47xTUCfVn9DV/vi4dV9xHN8A9jgj5cjWhv7Aoj+JSnmz6wf1qucyUOakNtl
GxmfQ/T6AlHq/3gwJGknYNoNdaxcFhmF53RXVNKk/nWe9Dq2kxYjPfQBWhqdIe13ZLmmrDVQYXuh
lep1JWmU04rHh5UwIOmnX3tVj8JCK1p4U88zHPGkPekAma1FNSUrhRpNn8VmzuXq7MqZ5c5x8fUz
M3jiCGqg1o6beYnoBbE50sPjea8uG7E66BwxI+RAvFA3o9Ei+NWp5uObQmuvHjXeizUX9PIXu2iN
McJYgg2RaDZlYDGWepibfipXKcNCCYu0J40ULcrcNIAYnYkJsQjsfJpYsgEkqmwDpsCb+n/vqJCu
HPjN2rF8FqRDcaw3q7dx7DBItiDllD8fGBeJ5HnKg0OqGd4ZTJvOQDOluW0aS/JmWPwVS3sQpp2l
BKzExleH6ptvh642iJqxFuYvN2gxmXDkRz2L18gHzWQ5Yv53XTLEZl36oGHMWN8IHtDRGHGC/fUq
HadJsohwt4W3Xwdq8fYVq+wRTmaozItEQWxLvVUalCUwTcRgf626gp1dYyxoVNDKOJfNwEdESnux
DbODoXp5SUvbTIZqTIYdD44nyZAEG5RfnJFMc4USKWVa2udATBSqpsaIpPlwKvBEmLb8U54gqMKn
1hNgjuhzJF76AXBsgqlpMU2xcfD1U90csDC59V4GiYvQIcsS3Ns+kK3uzkmLXfTHwDIsFdGWqkNP
CKBgjPZDzN6HsTNtgT9K68C1jTRpYIyOaqZwOnR40x254As92p9zQL1gx4zfsFoH5SY/DOMkMgTH
PqO3FlnCbX6TVOIi0jBESrfTvDa7ChQNR3JBjMVVjwY4lOlqvzKHSZ+sD/QrUx8xmhhEiEw3+akj
4MdzQB5K4nN+cvXFNR3X8U+uboPsn3chijegkmwb2Xat8xZyZED1cchrzOAJ3f/V4tByWHCA5R4b
NRbyQMOh0yoTqLeOqS7NI7TLH1xAzPaas3WSZtNSnK6ISw5Lrjbi7o3HBMD2xr8qCDBCA8zfszmn
D74U2nI+zpcL4LX8OCwYaeWNgIbx5l842Gw6cpVf+85dltAkRqsMlQKCM55/K0MzXtjtvu5C1N5Z
zsnpVtUtsNgMERx/YpwjVIi2x/qJKlpPkjgSBvlAiAkO8ft9+LaqVwMaK6DOL1eDYgl6YdNnculE
Vd5/g7wCjxdWKi2ZmAt2F6GGZkBWsuRx0eXbNEHzssZkhtt9k6sTVZMvNCoJEEEiZFgIX2Q0cBOc
z9xjft4pguRnYCMAD+jgnX2PYGpSimTYOBWiB6I/VsCXmGHMb70JRsbyW268eM8LkvdFeAEfZcsF
v9TjJIDJaMiZEpddYp9rupk5sdzHoXL5YnCalnKftj3C7dVWe1R7Ef2PZqdk09AccYTl7jo1PffP
NGqd0b61bTasHldw5R1YMisELenkJdZRhFBzf3jZUY+BBz/gd5Z3FZSMw7z5eRWA+WLsBvISR9m/
mnsZqqDWTWMr2uuTFqCG1McDWQVcUKrZvDjhp/IKuhzPfRvqItM7mwx7gKahBmguENacYZ+Vc8Qm
1OCXLONOe4sscHMf4DUHmY3YEerNqGoYa+PHAqDtbYi/xzjAVoQGiHPjmW/OIcywye2CJ8cMu815
2/pqVMsYwRshinTcUMUTkgYdFsVs35M/fmWr8gH2xvHfUfQZxZSVHhs5PHtaEXOuLPEFxJkkeCBc
8evvqpk9gU9eSaTz/1iAaNQH57UJ5eKE6W7GYuNmbCXELIgC/Sk4xLCu2Fj7MAI8EJwC3Xc8Gb7V
FxK38/2sSJjbQLwHhrmmc2XjFXxYOHogd5+mKSNz9bBgBfPopsVbSc+7irriJlB0V7IcPgYYH9K0
5xCQpU7fAJ6Bj7+Iz7SRtSl0837zI8bat5N5wdWtK4IICcRRO1nVh9ZE103HdHwqsIQfM9NS9bzV
4iZZFFqUNHsx8mphwWl4d7M0FLPwC14DdBnx/t9sSFL+ccpPgTvFQdMblCJPPWN8T/5d+AdIHIQ2
uBX0bli0Tl1XGBQXsLWRoxUp2Gkd4F2wsfJlObqr+KKanFf1TToEl5vu67KBHHwuEICTvscxKzM6
kttkGGjBOGmPSIsnBO+K+J9A+b1/nGWLN8828w9sGKjOYBn60nYirVq3t0bFmyHk9sWIkQbxfCoK
Po86wjBGJsFbe/pREek1hwyIJ8qn5ITNAcTdtJhbjRYVdZnlvtwBfQwhLmOmeInfytsQbKYql6qP
k7+CmvRpOTupVUQ0WGDWq2azFVz1Sh0lvJ7WOSE5JMqHHzAw8lZ+NRYwtoSRxwzuBqtgu8RMMsQy
JcH3mrico/iBA9tR/XgseZVqEKmSAQvUOyORgzP7ySHbD0OT2sGlQTplHrWpY4YOwLGBVVXkBMxy
kp8rwahEONK6VDQzjS7B4J/LC/fhcNuRpIzu5HI1I9/cGBlfU5ZcZaXOOOUAqVli8Q3Jwq27/JqF
vvGdZmNbYHDlwlxEpUdQOP/feF/NHMGn64tuzG+hvlbeICIGBqU2LW6lRlRJ5rt3Akq2DjPSs2dT
Tj8jdHjdO37wqMAJxbGBJswdfQlzL50wV4T0ZE9zcKlLHDkHmyEu/EZSCYN/ZyVlC+y6ejKy2C79
vIQY0u2Xl2NnYVo82k5syEnm5S8z2YjYCLziyW1DHw32CU5+SJN/XmM0wbxUF34mIOD6zoaAq9sP
B5bTdM9pObdcVc7pKozaMLInGRWB8fuKc09QqoBw4i1AJ1edkpBCT+oiYe9J/YojS8IzbzTkATDa
7/Xx6LiKoJ8d63FuUcG5yUw34qNas790eoUdn/IiYQrtUb1eV9bISE/5BxhLUlgGjUhY/dGlPDLZ
O5xUDGJc/pNgxMwVN2Q3RSb0YI2vPbhp6CbSiUVGIM7Y/EQe3sClwl2SYPnxbgCNaN+dlemKmbZv
2sYETzNsHa9AFCOZrqEuKop6f+WPVl+vGFPQoeb08MLTK45QcWGp4vMtq418+/dr/EshRo3m7PGo
Mak9lG3urK2oZbWCatNk0QfEjPsAbFqERTnTsRIjpL/v/6XPAHsIWQFDhbstFS6nt+wr4VGOmINv
X2jvsafQMj6zLLtiHI/fMBS1Ia6+kgJHsYGHoDQknHDDy3kwYiQHg9xFhJPPmy3BRTw3/DWeFk/q
vBtvEl7f+KNeG2lQhRDU+JdX521zyjzJi3qySHBvl5+nDgtIL5BeTiUsJMxWh/zVBB9nsOIdmpGP
l399R88LQJlceW8V0JQNMi+4SqKeeMQmEMMvXac2qK+lWtyahwe5Gai490mnNrvM1cj+y/apKqNt
Vk8XqTXmRSykAvcS1IA0Qbjm7SDLGnf2eDIRwbddm/wW48HL/RS/iZhOr9442FhORewgc6AGjXvF
93dqxZcnk81WIJ0pX2cG7PCiynDQQSDphl0LXws9/XCOBEM/U62cCB4oVEv9E3QE00zQnxQ/hxpd
P/EPn16WnETyOKv2mBB8UugXNodLZF++RACjWjU7LPUJXJdEAf6TncgYDw3RITYWYg04G8WKCZoq
qQ4E+fYb075V4Yy+Myim5okjbfvXll1pKP64xHaTHl6fUEowNs8XMl2vW5fZmHQf8PMmAmtyOyQs
h5N/sd7RlDCKLaprJUt6jLadfJlzjxLvzDheN1IBJBdufnEmsFZ6mPWSW7+40KJ8qvMbthLjj1JF
hwPH+/Q8Ju3aiPShG0JUlDqup8oTVd0qZjyiTi89D5qz1pQz/3UIegw++n9TAWQptTA5MBbmmEdA
tcDmxQ+xytWtyIpVxYA3AewWXLQPbYdiTHNXSDLT1JkZDDovNEWVio+N4EXBC/kQQJHa9r7rW5g0
s8iw7yRFuV9saoS0GqsmJZrb1flHfFHM3Q4/0XXfGdiOGH/pi/tyoNpbUJWQ4doX5W2pEfDfHOMU
l5lHtMRLYALaHOB2Be/+woiVYJj2c9wf6MX44leIE9KrxK0BQd2tshppfOFugvyBq+rYzuCyDqGf
d6+oO/0sG/WlzRELWtJCbcc2Rs+J4XJMikKUnjPzK6YS1FDUdpn6vjQUv9i205ziNfVxC6gt98DL
W+9Eyn3fGDshb5y63GhT9iiFxOTs4aeh0okuTdwibP8ES5VkmF7P0WcghSAYzdYcQE8F8c1Cdmd6
XQIPOgCOWXSQLpAkmGMDsSEe1YVlrWepydO3GVnkM+oJ622nq5rMJMjH4TyxWYVOWJA38n9pnHJ4
/XAqTjjpOZjQiK8VRF5flX4ul6c2hQS/VgVbToLj2DeIgWFzSZ/KuEkti1wXX18EC9r5eNYz2nj1
+q1kbLLVKunnXbBHXgeR/zreAuPecDSPQKwtDum7DtF0OjvIas7QFNpIlMl2v/dIS4B1ZYdWu0sX
Dz42HyUKMw5FfF6LWJwgLxrT28mXZg6BKz7uxP2v7pN8dJhYmaTDxE6gFY5Mvhlzh/sIE1rOJnvl
es3ZldM69FWGr9rMBsn/sTvxiD7zpq6medO9B2qbgpw2QICIps8YYExnxU6/G0FgIblIK1HWV/cr
pKsQTRqkKDt2uZ4AkPSTNO4iiKeNk2rcEybvqeWjzxA7/5keAp0pFOZOa0NH9CkhKcetYq6GYrs8
ZfBrTnXOU1Iqt9HmDatRvkavmJ668bd6AExF7tqhHJJ8Sl9826X+atRAJtplN54QJVQAS+RHnu1r
Iaz7azKzUMyvbl2ioESudES/pKNcNsfQqZx/YurphulUqoJamTtXUn9gFA9t1ndqHzyoVvzp2Ndb
0xUjUpz2LqKS3SYKEzhiPtI3zgb666h/tjwELTOQgIZ8Nx0QkGDYyycGURACIGs6DXrf4QVJ9ENj
LbBebm4DYPQYnqsLDbBCxQXIFOVeDcsdb0Qg+DIwwEUAx2gT4b2ibKc1Eh7vIjd88aa+A/qPuHDa
psX11Xi7jsX+nQHfaebi1rGlE20eLBGu1zJ2duXQnUCOGvUNP0t2ax4q6zgPPRmnzXHeeBPtZ4IN
7YNfyOUA+BWNDEUd/u4Ezw+FYqpJNg8t8I4YhEtCWPF17wS9vIVxoZK9KT4SafWr+9nAqZ8XcHat
hbKJxYykasgBJEGJvqaebrVy2pBV+Z5eaez3eSUGeHai1ia18CYfKqKsAHBlEiRFPisvJODKxkU0
T6eg6AMdiRip5Ru9lFmCELJMq/Zh4C7+F8062kIBUyZDU7Pj6+OzzH1h675tXeCebPW+x49NNUR0
fHimyh3oFaxbQe8MVuqODTdGQPQjqKt4VS6dTwQ4Z4OC9NOJy58lMwC7oyNtHn6e+m9xRYiDPyOk
0/WQeLA2+LTGc4tyiEEsSpXDASwzqKOXCsr0+8r/iK/oZr4l08wxuMe4FfOG1JHDD7k9kVL8YTk4
+lt9mLenexW50lcRghA/55cX6tVOGy4G5HlLYt855SvQEDivasrcRINmnhKxrnyjdsTowj3qXJaY
oSwC4wOeAUqM0eJuAfi78IvQvB9GD9hmEryLTiGZzOFORQtuFKjyiyEpJd/CFfObvACRyhrCKqcd
A5TzZ8DVwyeQ318QpyGdYomWN3qwod8NkidkKCesyHLAKJuRDQCOMC3s2AQpUTJUaw4Ky9JUYXCg
Tzt0FmC5kF2swf4i10Qils/pRLI/Lh+wdRS2/8At8VLMnLpBJGG4uX7yAx2SBNk6UJjj3BzMaMvx
QzDbPesxpJtKWEtKL5GhMRcm5n8gXUhnXLNaiZGc+VHA0yBbKnTU8x+SxOodtJF1d7XDZ4ITpSgY
nnnDcmFC32rUOUroep54IpyZgbhqjJX29SYzJDb8DVzn0uf248y8+I3WIartLuG2tjelXT1B6osR
9YOygVK8KkXIgveKAKzJh0pwvOcjw/OUu+30ydDOKx0Nitkv2Rl90Bs0qcVCS64QkEQO6heOAgMw
3nXUfzY6H5BAwOKB3+SIyjVK+eIg5cp5Z3z9eQLQKcKJCXMCLvlqP5PgfO2aNLZk+UC5fkl+P2w6
uOAQVVTDer5B1obbVoNMwZdjuc7oUNVXiHUocUrFAruD1kXeZ5lA33DkHeeU7dFJqh3zqOeS/hYF
w69vyzinErtKPwtXIVVDm8GrS1xQDj605EeT0oPLbDiyIBou2E031wjThorq8t5QLFQ3UWHJu4kE
dfhMvFHjZfzAhlS340TJnA/nfo2y3Sdl9dtoN58+UN5Q9EGZd2LvK5f39Fhkz2fAovYf2lEDONdC
knpc+vgyKFBiH0INOHETf1FnLBNNST4DxnbyprNwnnBkocQzr5T+4kHvSrieZmwhOard83vZ/jrM
I9mis4EVsGAf8DaYGGchrMuAZrg9YcRL+EEZpjPvu+E3aGMrb304eRC1qD+cJ8qKEWBbZdrsJYMU
xip4i7nG1MsjFGWOagck8K2ZnVYBdTybhBmOTejsolwgqpaHTXwNDWIziChbOU9SEpkXi3cNQGcb
2Jy64Rk+zSaFc/1+5+zSZJikIYIiYMud5vbFBe4vGtwGDv8elgOoMTCU66xriNP/htULSbuXqfJd
XLWZ/VkRBZSQewS/DU4/1QQdCLGh1mdK08OutVtcjvwoTDBY8ZXSGCjLEDl3n0lrzP0SBHEUKBgP
89bfLdMn+OyIleUcbnTNRr5jnr0p+VRvOjONJd67fDwfl8YPyNeoDTPqBy3s+btKP6tZoqUrjK/2
n0FyqTKz+wweM7+BQELUp4ephR5go8swjAa2dZvjDXAmQzm7P9sb91eVblDnWNeGsboZnEPWWHVG
QjzEZ0IzxAs7s41T6fmEWhMZ3jgpqv7kjPTO21/xw96E+8Pc3BmFO1YtZPVFLbZWMjIBjNrI3I6f
Lr3FanqT/+bW/n7zYGyVHJKFFrgP3HC59yGqYvRpKxfyDFtj6T9D2jF5AOefH/7mt9j1TH7XFpeH
1xQ2j55wGIP2gQmT7+cHRxr3PWtG5yWEi2SetLr8mPcVnCW/uPsnurDW4kRhht0D7EwpBbAogeVa
BB7R6fhhEA24K/bm5ChLQmEZeb+ofaKimbs7y/C1HmCfnpr09g4Q9d4ve3PuoO34AiS2F+FjY8S7
4jw8QLKlKmBKYlGJlBWTt6wlL68j/JukwL+s6iUMj/x+XwaFtx+lRUjAPdnT23GDig1S/A82Yjai
bDor2F6Z3txkBSLKb2nldWzPecVZPjs9Gvf+ZiqCjTBr/LJOTM00vVT7QbQYzqKkNz2Rt/6Sodit
aApwsQRD/e3PqSWC9JhjdOG/6/Wixg6655ovnJS3ix+M018FnJ2VcoMPAsUvJRz/OBgvtQ2LapJK
aGR+yoAHEGq1yz1cKz8zDa1KrwAh9k1uLGtG2VvK/1UTVJnTFdPRi0kfKfKBQw56+ZydWq6AZUvY
WRdoGnpDxPHKteI7K5GJ4FISHjsFT88SoatXfmn5H83YU78swIOnGg+x3KfHFLMyrKqgyBWJ4T2t
2B+7UIa3BMCw+/zzKDweCfaaP3WWZ+jIqxdWWWNGGriEBlcwAiBHZnjDK9vuvRqknSyCdp1g6rN7
IcJ5xMGSfVlM4qzEgQzOx3G+jBNBw8SO9ZR9to6IqKvPBp7s0XiZ7GyvX2aIjBKOIMof1EaMpWJ2
yYumPUY0xc7u3IitrNg+WJDVImTFIRoXEeCOmjPiZTnLnl9uhxTApko25YmytUYeerbdN+hkqOay
4wZASK2fNuT3wIGxOa5TzabSVdjCGAxbtrgPsDecgrFT8wJHHBB2uEDcD5Ur6KoH2D9N4um1sh3f
UX/OP7NCSd0wY/kohjndU2E3RYjnkqpPfqd6pTmcS1OGp2w97MHK25RbBwyqcHaUBPLokJ+RyYzw
lyRQGT35Xky4zsI26jPoz+kYdUlsdSu4eBnDPfqkkomFXMdT0SnujO4BtSKV5NXkYKpvp1Eq+Xh6
RKBFMITEC/NN960Zm9gDtWZGBaF40RO5O5JdR3gN2K39bAspBpWXjBc3x0wr3WQFNt+5WUXk3CdR
CNIwH+VHKvAuFhkcDxP03vEzSY/P7wt9hqyvvGCB8FepSkJXQvbY7v12ENAylUo1MOFtye+wqptJ
IeHME7TyEY/2833N3jtcB6Nh7o7VilJrMPYT0gthN9LYEz9ZAadENoVdgyMkXqYSavVqUgyPZFhr
2UBhBTq3HOonRI2lVvBFydgIl+E7ZTZp2j72iDI2YIARHzPLFc9KVonLMsGhyNOvYgDPtU9BWZHh
R97mOVuJuqEmtamLLa0ohCvYGW2bwnh4cy6znNYysxhRMZoMKB5yuSO3kf9gKVKZoH837zfae3sU
FD1CH7A5jZFC8e1Duh+0wIS4rj54DB4m8eMynPfy8G6hkmW4Uj6BbApUDGVYmX6jPOM7iZay9ycU
9WgkCILj/Z27KWzueMJeDLPHlLnJrggAv2ri0UOPPzdaDJ47AUPBE6kiX9f5NjLs399faRrAxl1V
SEXlOJ94bGP8XZ5ROLQ1r6+J/fvvUczZQK0hebsSz6vZPF+HHsJhnA4elfdR/sCuYcgKxr4cO/gn
/i8TJGcqb1I9C8y1j0hq1NAa2djZkFgDu/OmPiq+OZUtzEhqyKkAK23WIjNFJqcCUauh+l1ftvtP
oX/bSo/6YlY95cSFmRjYV9+Shm8KpzU9cSGTQ7IiQRTNO1s5mdhJmAa6Gbg5rhGFqhAhz6WJDtu2
95GNKngK2qa2Dwto2k2CzWqZJMpeqAhgdpRgfseFvdKU9/pfZ9idQoXmV2WBINZk3mOPvloBm7PC
jx4ZmWqbT1ywou4NFrUC/QIWfB8xgu8LRlyD4cSrdr5sMFzoxeutXxBnDKBKpYWZKyyqnmxYn45g
yPkB7JsBhvb56hYs6zsYKuIaoCwz42mIQ6OA2jj9XIVh2oy1CWU5nmVljrlpA6vXtbpo/1nKPXAY
6dJK4//hEU9z7ECoAMvozgSPeJ6bAieM8tMR1TWcuzZ+Cr+DmSuoFsOX+MEoewOL1LZnukI6XzOL
3DRWHwEMVWkkEPEQHUuCt1ErnFdYSrYZDK6207fzPANj/V4vc9Prr9oCzkFA8Bo6BErgeLOiGzsC
sMeLu03/6nOVJSNf/N3ehPM3xJZ622yEJ6yeyaSp0znR2fUQ9bj8kK+2FpY8Mw6eAMSpZq6oqTOD
fRfD/zaTNEgxb1SEN27ey5yJCbaqEJTWimOK7Jt870CkuEh0hzuEJp4ljaAYFLnblst2SFqSSN3Y
HmV2GSA5RXqYwNYWLfe0HQnFjLVdOHq4v8+2xVIAcdwSsAYKvZLXJBALIzghhgkwJUh8H4As73MM
nxrnl2f8SvI5mCoDSHydzFyDOO7DxbkYVu+R2SsqmInzNxCTCBsgrS/FFs438hNtXt8yn91dF1HM
7yguKN9CXVl2ZvhFcvB5FkGlFbIiFdaoIhQn1txi6a+JjcgfDaVY+MetgrFa21omoLInubm6ZbUn
5XRmnt1Si8xSZ9dkfkklJhKo6gE2+mC187hkToR82/nlNf88j5uWtuWlYTceOhIREt/XBvpinkrF
xOMrzbws6OVWp7QZqqS3d3bOfvgs4PD68ZxBmgEsK1S+lVVy9nDAH3xWlnnXdas6KlIwliaaD3A2
yblxS+vZKDNUACDZACyhpE3XEqtHRFoqxt3ijqn/hD9u2zX3yBIh1s4/YlQ3ZvgFOYTpjhxp+7nV
ltyLeqKHav27fhYNTdU/D7XUuJYentAJw2XbinCTcegRvD3TR+fi3poLAleR2phJ55vqdixJqV3j
RFKGEZY/Nv2akE6SPZQS485Nz8f9XTt/dxyduQ0lV9eDjzmo7DbA/rLJhUtDrbgzQrF19VJflVbz
QInXPpR0fu+Uda9KMp3bJod/blncKhCKb6WLkOutMWvzQOG152zty+qARrhdbmnrA567ERVcOJcE
J4fSwDsn6GyV01v6srLnSyzq//+g1hupbISnSnoC25xrFinu+kxMo0iaM+/yFv/oEDS8xrUKw/bg
PJ0EURbEqAwSq2ygv3/QxGzAoh7x8srAN9mm8qS6icFDhJynfc+ftiBF0cKhsG8AUO8sL1C2J0l5
fyC6grgs/owJ6u1xr1R73qSgo7Lr/jFvURimOfr1RBi5D1TScTGnQySClNHDXvIQ1lKbr+UzJiWW
ZLpk48jCdlQ2226tn6H+i9/Bpb7NiHWwstp40KyvcTveO4rwiG/rLe1gAavZRuQsMi1/azsVEOdI
Ju+DhTv9xbIqFUz1IFsHEplfYaiS3U+8bVMIZwUvWT/uYzKC5vEC9RDYyv3+tDxRbU06o2X4WAkD
HvoS73WYsyGzMH6yXFXNljyj+x5ZsLe/qMIESjpWjKHuOA/e1Aj/ge4fnuOEak8A/QnnFkqDzo2G
0UNe5ssP1nxot4gl4mZVKHNv3iEPMYo+Iasi3j7Sh0/UkQHMZJfxmHp04hRT90u2uncDqK55C352
UBd7LqfoMss7vkp+7Twq67Des77Lx5/kR1rZw4amLwq72zIoqjgKahxe0TJd7dYi7cyL1aRPCrBm
clsf508wo17oQqDIH+jvb29NGgFzEDABjY2V/DkpLwXdIWJOBj1b/VPsFY67QPeWskTWuNbIn4Tx
/I/IBfJUrNFzOqtjOROWSv/AFblyInX2mqz9Eb8daYKQsRoBWf3NBpN9RszzxXVEmEDRy6iDO1/p
TDIH2aVbCCW+2IyWvGH9Oh9vpyQiErxzaZshGT4oo6GOHlnCTy1FTUdfwgSiW9qJgExdabYai2gE
I1r1p51+CHFhy0I/utmqlk1piNb6eGqMCn+D/4dJfLBTD/i7LbIQAeIlG62c7r89sk7GWbpTM5Eu
AKAblXXPcxux/iqIu01Rm2h2T6ZncgOa7yoqCda1yHQmlWyGTHhPMcN84WOe9PTQzxOCWDyNd7Z/
IVSt5T/StCsHXcLeSDB8SP0kvPBG4oKWL+87qFuhpu+XkgOXAY+rx0w7SiKWkciTg1YtxJ5InXea
SVvYvvCKIsbyn6+1m6ZlzMqEmrNqqOUiD2J2JgYharzQoG0EFRvy2wpj173aNMkGlUCbJK53RnqH
BvxE1HAdZeuhgzY3ZM663f9kfzS2n548//VDOyn77exzS2lEA9tyqO8vHDKADyJNJeA6PB7zafpV
oQ/w1JEb47ThTkk/L6IU8quGRaZSQ2MZiDOVXqd1E8bDtnfr3clj70/oXMO/VJsAhWeGlygFM4cg
siqs//AGA3VXyXobnE/Mm+daNUl0thA2C/aj7mv1bqLEWDopEhuMbzV45PIKuwyBs0fg/5lIRyes
ySAOmrIaAgDBum/DtURiYCTwU5VAlfVCEqjNRAyyg6msU4eInTzk3nVVJnbKsq+akRnY7G0LLsAy
DPz4BvdD/iCnKuDDQM0ep49tMfISsQJ01VmfMskJvKQg8B0qxiIY7aSMbXzAvW+uVZTAXcqBKoma
GOW7lGRSO5iEoQwaeGXpCPmTwG5UrjM5RyZuLFqJTooVWMheyYgucx4+SdjWH2f3fFi0MP300EGo
1w9T9t1/hqVx1i2qjs6cK5brrPZOGunnH5amFdr8g+GNa7vm01ZyXUdHTOFDeni8rEcFPLLPirYh
arhfWW5sVbsXbfqP/RdIdSq8NavWL4t7m8hFGp7z8wRM3JrAwCtDPrVJSHfA/3MwUCRl5cbCBzee
OhC7WRPXoLfU+wWWwuNI7GwPntaDolQFfmJ9zHxcWYAdeCPnSVTSSzw7XLKjoYFk6U/G9TACQ/u6
79CWegvqiDzssJBvyqYkggcNACBCSNATUKG1qefCY+OYReadkhyaJIQnbXM0FIDGNhtl1j+x5n9P
yYkY6EYQFx/381sYoOvBErgHhd3724qUgt/gDk+HKvkxM/bVvuQeIy8KTtfNHzMk8OmsohIViUfE
XJuVLD84b74kNaecvCtvC9qbfRvTWGU3qISov4OyKw3HuSdZRmNSVzwiXvkRUCH+BnCjTqlrgn+Q
EoexgdViW/Lc1G6e26VM0sCFn4kdz+pM6PU2HSI07VxBREGVOUPKelc90U/IPMo0YpdJZksn+DQD
21dXV0k7exp931LxrwfuSr8rd/z+IMRoH33vgXSsCKpA6FI23APitChz7wDurPuU/YJwGP4GoaKO
bPsahxmuvMi+w9mB2puXtOWqhWCZnNOV8ly5kA0322Tro8PGS1MuoC3Tw1mgTNd4PTiV60LWy7au
5IgW7TLI0at7x8j3qPyVxu2M1fD80ouq36x2C+hv4ZuZd092uwWzeHSPZzOcozGYB/sAFC2zT0Ii
niy9qERwsS8whz8GVCgUdaiaERKGAIrWdFbl49U0h5j1f9PcQvEDkvHq4mDzn6R7z/xqgFU8I2fo
iGsvmjG/bG0TBHBAShih70XacxIjPxAd01sb0M9ZhNSroo0Rk4RlFIf+1KYHnYhqBosNFBSYcgcD
ttTEWDnJHayzHTkYArowRbO1g1nayD60aJ90lZ2ImEnmzwHrH2ZLTm5CMIJkNrkYv9P2YXjehkH4
4FeSrxw8IRP8t6q/EqLbshkD0cnXZ2tWClcn1imklQupBPS97SqDS8dNs1Em+aaQ/w/+IS3ezUsU
I9krwscPihq7TqaieiryCepJdYgf+5Bp11D4ld3/Gbz0bbwNJMe5e1xkytnsQ9UABqQKs8kI3X6S
yMPYZtOLf3Glnvj9ITHD0hBVbki+geL+DTYyCVnVicQscNkbfVWPPsuLqfi1IW9+RBAcfYjD2Wuo
Pc0PWvdQ74BDVLRMgx2Md/EpeNbAY/aEbOqnG39J+Qd5kUvMUUgYm2UBEGEQXi0W6K65jZ+wqOBX
PnwmC4acWw7gDVPspJivtFwU0j9mIJri1rLHd/C3V6vNITM3ruzcDKha3kMULf5edam7lMaBfs6Q
1esTs8Vnp4VTqLACwIiCxiKnAJzU0dojfv0a+3jNE1OxsMB3yrzJWGrsHukqZ0aEm4CJzkzx6kdX
8JzlVryDoIdEBx2oU9AMekapoHYQOK55kLVL3zFU92Fr24izm8xwuan9117hUcJWQEid3GFwhZWP
5INeSkjmlCCl14+yjmBYyG5b1g1cNNw5D/WgPHjEQQiU3iKr03Oe4tDvwHaWFBJkGthrsjTtlr1T
nkGKC2HEcyIzxZLm95B8XSVDsjspw0a4cIrgnU7z2cNovtDHZTcE4QpN+yBd6EKE5s2n3RfmhRf9
Fz2lPJehKXjLUlomr4+viiGHzZNr0O4n+yEz3DyLq8RvdGfbMOZA4kJYePgasY+7MYqLQGr/madb
iZd5LXYqP6J7JP/ixk5aR35ILD8V2o8Z8EcqPAShIzRKcXultOuKL2GI9TwSj/B/qt7R2IAx5K71
/a6xgxuAyhKfJMQX3n6zVw35Pqy/SFNuFRynsUQ2qOuPcMS3HI/CCjL56PaeRmjnRFl/sTjhchD8
w7YyMHH4PRll71+DPaTPtaLkuRolYRjYEhOViMLvXihuI5VpejUpUPzkQclYamP/vJ7piLOt5k7A
OfcySbZ2NlBPe+XzFJrN5oL0IWxBp+oRy5VJzfy1RhctPf/iUrry6fxECAZOsLArhIZDAOleJ4A3
tYPWqhWkbyXtBNGxc0DTyu67Ovx4uWKXffHiBDw/n9u3MFJGSKJYEuQGFQt9YVYdXVkbZUs6IdIs
U0Ns9V/YimgPnmIkU7/9AgRSoz3hVkj3pshVC54sjgQ44ymK7ohptOG7eLokuFZwFH54txJmqMc4
4NDkOBRskrdeqHUJ30yUT0GBlhdV2EkdI7eroGcE1qkp3dsNIQHVysI6Jq3XuC1FdRNEvsoqU5nR
aWzyATgu8/vhZRRMLS0mD5Hd8Ljb5u8cAuZ1WrYoZsyyyGSTaskU6ocpxeCitcQHWyypI8AM/xtP
y3pgq1gJWrxuUNfxOg9QaIcx4N6X5aMXntdUUSKmmE7oX03tyj69ndOjoYi++phGNkoeh6QbkKJw
IQbXlA1PxPedE1hVNmfIzfbODPUqXPVq7+3lnl2eCX+cte/pgTJ3uDBe4wD0WIW1gQ0XoUXqLsG3
qWG58eSatzjvrdQPPsmIiEcEy7t/BR5J7xoVu77utxjqMhExi2ECcJm+CFZ7Oq/uUNOR4/TlK5vO
hkGw9aDhem/8ENksGBzvMnxPs38fN9HWokX2DwZ12k4j0s1wY8hd24Xi8yxyDyYUUKXeNGERwHnF
WLlGZ8CJX5SLcjEY6I9cOuKnsbfgtYoA4HRhx44/xosyLxuk8OOwdvxx/KI/qWdYmaBVuDSmSTuo
5mfe86//D/EhraphXEUtDLtBbeosna2FHM66obSbKQ3OjSTizESLoMKGGzqd4owqxoG31BSHH3WF
AiNvzRTpLwT1shdfUdWCM+wDhm4yLjDG6HE+1hNFCRuDueUxc4q0N3kMdvFocPaTv0fkqTPbrjFS
hWWptkI/kIWpWG1TA0OS6bfRMUZwK3YxWpDbunNaVqPHgasdc4mJpc73ErNVi57y9HxEVu35Tghs
j0LMO/7c5Dqd+YEbmO3A/eVnC/f7ANmYIrD9yqGysrpC5jPKh+w0xsrwWJrORix66wDuyVqVql4G
qo3h4M/T37BnJ+gsQ9N4adfrGzsIjZVjAWHNxHZRczNrxJy6ex97Tzutf94bZbNATzqQn76Ib4tG
swfZxJaa7aeN2gN0o4bPK8R1awkyuK3MzXGyD228y4myuCDKZFHg9KRra3KsjrX43MktMwHa9RZ1
0M9S/Z3VYlUVuS7rM695mT19HBYciGd8LB/emNDzrEPwFRZPt8VE7OCiog3xmBCaHmA7OVjvvhkb
yPfMDshzBwNOVGBkwAmTrQJOGpSvORxMOrYlYST9VEXZM0Zv2As9G81/uST8fbubrxSnU2yl4dbd
1bnajj+tpmwzVysMPgjmuc6pD5KVrFxg+pAt6uCqhTjh5uVsi6ajW9Ky3LMKYbM+nS4hhcDrPRM9
b7OMTRjU/kK9MiR54uKrn+JH/lH5u/DthSsOkCF2gtxVbXOx9Cy+HpEuBC6/6nc/G99BtFeiyDE5
8QzfZXM9SLHglmE1NitiZp/20vh/NhqYtoK1Vd0Y/BhZMm54HmE6E+TuzrPROji5G2adGkF2O8d7
9MKN6C6PwdUPV0jaUiNBmMcu0tZqgJ3zODdQa7lZZS2NacVQv4NwcaB8PA3Tx0TWOvtEeGQw5Wle
nNW0D6ipQrFSJYjDbwBkH2YnfK0ps11qDrTE6utgB1n96jFB2y10vYw3AAOdBxxhM+sDe+jwdqHD
1x3XltYWC2mgh/xkgGFnmCPhenJ12F09z5gkOC0ARgo8el2jHtSZCoWsJ08zDi6PnX51kWxfVknI
h4iKTr8LqpkzVksy3NpW0Rn5j9TznkXywyiss3P9+TwmPCGO90pOHrG1hjdvU3LzgXUv3LyztqvS
LFhilGTeBvitHTguqrhJfyLcq+dLbphY4Vm5Mbi6xxFFBQc/vmtFIg86ABpnqFg7c0NDZ9zl3pgq
sKPGY3GFJNivssX850ySue1es3gVjI3rlRTiy1gh6dYTGm/6DFfBqY1bm5b3WwhDhwpECpemaeXJ
klxdQiy6TM5pd/xSlf9NfusHKb/o96xjwna92+COdiHpfj2pDA1S9umsUirwiDxZW9DgxifynMKr
5UstAZRPxvC+6N1H7BV8M0AHldLjJFH7igoOK5H/XJi9St87vl1J58GsITfgUFo3SHx8wBY7IgaJ
Q5Wv5GEBXAyAuldlDU+WYMF1wD3L5U6btxyjKRYgp8RXm1f1KvCQLD/QQe1jI7oXX4TNYPSM7Mh4
Q3XVOD8/iNM1vGAYB6qxOSRdbZToV740CPO9EJRaXa8nQ5k59qNoMGYfx+Zp1lo3F2niiw8RsG98
qwgtLCAmsmyVj9qrG5CD6PnDLVhJCr0k3uVjAw6b0Pl9crDq86sZzFvwmmIbOwJZSEODoTfVm2n1
hqeDDC6PASY/VLvlISq3o1P+HGvIvglGdwKYOLbc4HLVbIgj9mJhWLuUpvMOP4XEtxf8lUJC+eFi
mD+etDtsiKyeNyMOln9Z06M5+dUyDWhJx0t0CnQ7or0RnXBBjElIlgqbi1YC4MBzHYn5TkEtK13M
uR/Ae5bd/vMEZGItUgiA2yig9CL6tVA5qEA0oGnSTazrsTR6pzVGtDa4XcaFIAYdcGszs3ppjCfx
I2XJBbKg3OlTIb+eQJA1Bldvf1aVysXFObQNmdBy6b+NL7Ij6AUqZVrQnucXQSabnpkN5MRVsa4F
ih+tn6Qp4JYIkB3xfS4tRmQT5oa/Q/dEOasrgvE70cMU1g23HCilvLtvCWmDGpDAciemGLFRMy2Y
Yr+Ub5Fh6olSDgxzDzfpVqb1/BljhhJmYIdG1nyIPphiqTnkCOvqGhitutJ33pn47bSDBc+40xql
D3lUxQMzqNS6Oj3cqs3p67H5fOtnYxfUns4/jNiP6RXujboBxWf+hFemsNv/r5/qql1jhVHKAw0/
lW4bOYwq4HRIOOVlo2vyLyGvrNFTgxgIvuYXoKkeGl8AbAlriwQdgAP7NpwpiD/3N2Xd456EmNew
OaC6pKiqFc9/Qah0yYhOElhMjB3eOA1lMrIcCZ5t0QP0+T/TiocWlYJiMHhdAs+b5ZUcJCmisq1b
gV0gBJvXOcXic1EmSFOfjJmkSnzN2nD+QKBJgej3dO0YYKwB/+86Wd1buiNc9yHO20MFEO/EevLi
C6y/mH2O1dvTz0YIGDWAxV9LG+Nyv8XUj6GGEvNlBL4XQ5exNB/ln0XgWFQa5NIqSWHH4rR8j3rh
KzArwRy9Nd/kAWsayMvWbIWmv6FeBEJPySIpH7k+JdQ0gqWSwQNazdicOW/OktCMNgfy8vlwG8TV
OmsEIdvv0U/p8G0VO3dIWRA1lVR/MVprfjhFPd//jze0W7pNmUbPEy5ueHxOZFLa+AUihkvu70q/
z3jEmVeCTiyQrzzDjo8QL3yufxxWGjuLDQ2fhghSBFdBb5Iv+Aq0fL4yeqBVg9BKJtXd7P9Nzy6W
jNsi+dddQIZpv1mK7zSzB2l5gE9uNNsToLHRPutdp7S7ew6skUkV5lKraAVyecABo2rdzH6kqICu
qU+eyOhxiUfnVxxDyvxL4sLlmP3zrivwxOsnvRkFDMyggqS624XrzUDXSQ4p9W4SR/bmkGQpejoY
sP7agTygRR7kst44OxY4QNh/sijSWV5fG16lwbPPjVE6E5b3WcC3CsMBAG60xE78G1QaCYOHi9oZ
fvaSG6zlNI9DGCu319ygsUtTi2y/oc84kelbWOZy495ftKioCNyLCnfGtaG1GmG3x2QgS3ep/F5M
1wQBl/h+T+mE7jLt1MyHNyRVuMOkMYDdMtjfnVcDjjrfk6kqYD1AAfFDLvxIzvSnGBr9w9MpQzKZ
yIr0Ddu3WcVupo4o9pHUiiyKCLOO1zmf109x42OpAACpln/NSxXRBnrDbM1lKBzXGqlaqxngKywc
ph7zY8tp9Ibs3vKXn1pxQbhJmaWtbEOKNwne0mYiCG6i5WpNf6TxyT0xjlOV7zvfP4j7HGXJ9q0k
S5VXnqWjqnPP0bEmHc8Yqp3Vun3evQMtWtDKiOdE3u18DZdLTw/7Pr+O6I4sfh+ehs/85Pywd/y2
+XEs0f2oKAhXAR3r2d7Lz4ZEYcch0jJpYCKjo8zOf1Vid7tgSZqrYUThFfgCrJR9KsBryhC35vIH
wTc+9WN+XMFpvYu4KmxGTOvJE4EyEGvUfoUvHCfFW7H6t8ewnvQPILYHnKgiIGh03oGZivD4WhVV
b+ZcTB4ei8EGjl6yYhym9JtRL/cOIye+xXv9PXg86eLIORk6uAs9DQY2X76nAVeUPXT5JZA0xahK
9XlyDVM+f/g0qAyQzojJsOe8QmMci76XI2UEHWOVYqfakEbgJrFns2U3YHMqRbxWSG0x4b4YJFzu
fmoYFyPr0HYokQGtz0lQmVss7F59niHugkEwAyCvW2Tzd7b7l5edBfjBU12IyU+m/55k8loMl9G4
fT/OiX91Q3158kEcZj6s05+sS4MwbbdR5fTfAENvh1J1/gU+Uih51N497CsW76dii0Z9/e5JgFZZ
BJ3Obuxxqax4pGAfoJL/ETK5kleqCOwcpp10p3q/qOzd3kgkxTD7XhSUhRSGZBqfYJXyNTUb3UOM
VOFxhHvLUQGx5CsaKN6lh25JAcxatc39XAHLUR6W0NjC1szC4F/q6bqFzgfU8EL+YdUMMJNteOEE
yFAUdaFOECAMlMZAg3xEy5ucV7/cYJC3JQzJ3dIAGXusCoEHjZCHuHoSSG/xK+yLYAIUSGXEUy7P
v4iVSacjpJuzYf+NCpLATIVPFvzvyc3Vpf2GCTlXwRmxk28q6kONQswa+s24qWxgBt7nE1Ocm30l
vjp6eywHWpK/MmP7C/T/viVqeTqWf1pWCol/3b/GR47dkgdoZJ5/lkOC/wlnm4IQG6ieU1VgYu6C
quJ5U9QtWTtXgdMX8Ysjr9vpseSiiAcz+ig7Xa7nHnUQKOZKRRuxCjN65NjYb0OWdjCfGfunZWdS
bmadvRrunjCzF/DvgVVdqiIsuI1Kq4ptcJ8xne79IWJJupLW7HGtJOOO/2CJKXw7GnGlehZFyxCf
NBkABii7rppVzE3heF40Uxf5bknGyzc0IMhKfPdAYC0ab0MLgOyFeNenEuw1QfOWuQSpqBi3T5m3
lwAmz2s3i3pVb+XARS0noiv2xpb6yM8HnvRmflXfWrro1tJIUO2uUZ4gBg5tuts93gpwczfjQNWh
SceO/2vzNWbmJhNKeEnF4vpw/B72yD+zA6wttOiTyEH+xUc0As8ZCpMsFu+DZYZYCQakxLav+FMn
n70yBoHrd/f0CeJ0CKQht1fo9gPFj01NIWgb3GiDYzkjZQfKEikYVO8U99xowah4Nu1BKDUnxD/+
BY1LVHOL47saTJ+rjrFLWmB4PLnfuk3dgfNQ2FBS6Te+g32Azr1MEmP207UeNpwQrdrwhkGslNKm
lA7qbKPDwf8YzbEaPB8PMxqe30wUrpoSlbHXOh69NWpyHOZnQd1j4anYsAKo3FzjoUH763+GGnsY
G+/TRctooyQjv/sjmH3UCUIpWITcb2hDD7MPMAxEa9v6j1NZs7fPkOrrUC2/YtpX3w/0YU6pFxZI
1oI/A9j+s2D/GSzsrpxyYqsQlPpH1hkwghVrfPIpWWyGBfhmkqtcX2nm/xXy4hMSn/QjPAZNkj8T
j7w0Jz7fWej1TUaAfHC6JkbGRVWjkOmCJ6rxMx/AHzOmMuI8WCvexl1YeWWvTFdRbI4f1l/zWDwL
IDV9mKl41TR8K1HYS7/7WwVrUlfXvni2gIpn+Y9VIq9aLuAA2tRdyT/hM+gWG4yOZJ2kbFP3TBUG
3eZT3HHgrGrvQfIn+hY5Vqboo1MtsMDlJgsoLRwBpd3KWJY/DomJBoY4sVEVQLLolGOT4dw2QKYk
kwmBsTwbFH+C5Ae/C6raIZdr5VFRAEuzc5orRjiPvjpEwl4DjAzzh6YhSEB8yofiA8yItGKNE2BG
n2FcOQp7uA8x6gnuu3RBA+rIQdjGLYxPvoL9Z/fXUZnhLRhVdddqjj2BMuDN/HAmgO3kDQ0gU77I
T/DLbGLcxJChXNOKYFcrODmwvyCGgziohlNoLsOmwNtmFp8mAjpT1r8u17er7CrZpszTjNKKQCDK
Ul0n4zSG6EO89GbW0j9nl3WfPyWdgaforVaPv8UdaTo8/kr6XJlmDZsRIBT2LOGYRN2/lqf0XtkB
KNUhUvRx7ON9z0ZMDKc3CSq4CU66jpCo78RnT4569VBC/TLEVCs/yG73tO0dbhdZCPU30f0MHka3
YeztWW25sRTg/hCaYfYRo7IAg3CUeP3fBI1K3ZVE+x4KGx6s4Bxz0Qi56t5DBLJVleTnfVQL20nR
YpgakmJnbbe+q+JG9dBNTSIrldqDUedJUFLmrwqAlxYWXaQuL8mcvQxuZkaCK25+Akrrx/xh1Xye
TWWPhPVuCrTm/eiAe+3GK9wEZigeUWP35YTeicpxYAdZW+7UNhPiAE8IrJRzM1ZnP6t4zRHqCJ2x
M3KgsUwIGuyf9bzz/n+PcCfvaho/WOZ7ZzMPy1VOw/7G323CyhmnnKStFqrNcYk3oHm+2yJHBB0K
NDYaFM1z61p9ikK2rRSDq01KVjf5EoGGr+KOQT++mnbzAjWRAgWZWtGiBckMgx/BB96t1cziijiw
qywdlyLZmJgAOxc49qVpThF5HxITR0j7LVJ3z5YRuGA1L9qME6uuFbUAu7Tk/5kQNP972q5ZCIXh
6BOCCeRm1EznBZiIQAaay46+tLnMw/zSxTE5wbxgpBto8nqgdji5ExUtbphieXrZY+u0e9vnZ00r
TyJtJmdxlIgU2OUEl8G+efdq2pm1ZPkzOvisB4suqW0/f0ndJ029KPznVDpHEr6+LqWeKXjbvb+x
bUX+DthTBTEg7rlAaYIz3++0brQCMmLF7p0XePDnfyppQU3GoTrdsm2BPwKO5S/ri0hasAK9TeLB
mu9zSH2dsJWnMfT/m6JwvimVk2jqRxXVpd1oIED0TMFrmH0SUo/3j0Kk9euUZb2Z0WKnsPVsS6k9
4ieh5waWDEHKLoNv8vKpMYzpg9gYWbbvgOgBzjSQgs85ClEvcV1wG1YxYKUdJHs03shmPEKRe3Ij
x9HTRv9ScyO1S/mHSIgSr1pxsqlQ4u/AyyAEY8Y0wIPJi2qHZAhtkZFJZ26IgJAWTIxz4Pld78Zu
ggHO3mUZ6Kc9JakhzA3ELbEaGC57erPVc9d50MokSGBtmrySZIvcR87K/AZdZWtiVrttujgivr+R
8fZ5SSAW8ZPlYt3E6GliDVz6n5InKmaKa7grDYjAFTbkOYvEgB/i1XnEPnXT6NEx8bt3OyIpMcrv
XvEaz8/bv1aeHmo9XfiNujdFAfjdSs0IDbPkgtzWxqTi/M9xJ3XrVsCZ9nO/eAMQhQ7N0bIkmv1F
3PtIj5dyHQoxmlkOWfZfPUw+VM6xvQH9xGk15NmpWGEIQn8m3iMSV0jMroVVqJHBP3J3rsg+/0Av
8VKwm2M7+Bla7VD0syOXLxpj3Fd7rRq/rCM9Mz1mqdBGUmo+X8z2Yi0hsVLo7QxGrzzbW50nyfIO
LDPse9JRNFLQj+HBP2STFmMkGutdED3nHw1mw4InG1N64FLuQ59NzbCMTLJ6Ebig62xnOJRW/c0W
sy+Et53v07nUbrBw+MjiaiKKdHrFY2PmG27rkSB1KAh5Es94Dxqg6w0dHkYIwy5b/lOLg50zHwRB
PC/v77clev8r/X7Xru8UeyEO6x9oSD5QEMzCi3T6zrRuHstHJ8LPyvsmFtcz9yKuuvDbtLn/Ri6w
T22ad9fDXGcbynbOoxbh++JQpbBtxOzMUdK9+Sj8hIWM7xGlu2pPJHaR0e4grDXCjno9UAuZEUOv
TR5tlu/uUZpgXF04BvhfeYVHOi044rCRmPGb0C2ChplSWaLYgXM3KjYxSpRT/XinvxwI3TBKPK+0
/xR8i7Nf1P/RvEA4i0uuHewNzzMvnrPOw0NHFQCMTcOBCNqIDHNlUa4X9opZc0C6Jv78jb6Va0Bu
jM8r+IpjMdLrqAkM83Qi4Wz+DGygO3hh2kV5+hhw8nbqX98suTl2aDBIqXkhGBcvuiEBvnA4rSfi
0opjUNyiTj1I0wTQMs07IGDVdsyuFBP761RuVnjmomOex3/GbKCTW0EQsTucTO8z/fIkpUDDg2jH
M539dKwPAC76l+CPfahCgyHIONCd3SPmSjSVOFqiXIq62KBHwN05wgWcj59Y4nexuQJV08wOfduK
70mbYcqAitFc1m1X8P3QyN5fbsbdux9PB94Ii1qtHwmxjFWYa1gTx1u3+3g/OZjWUYCzLrgoCXOe
QVxLh8ldc1gusBSgJHtiO+qO3YLB90zQw+1wMHNoAvu+Sg4a572CI/9RClT+AGpkCQc7+gwwqmq7
04adrjXCvDuBgLgeD5qHZ2wL+3MLpsGZs04TaHiGYTwRGwA7jTBs8SVLL5A7n5BWGMbESPM6KNtp
ijl//VrhU7QpYAD7iFqRiVWdtd2Nlc2sKlnxK/RBUGwRmzCl1+X8D8zprsnHGEl3SqdSgMAzU+Z3
nb7OOrDR4frKHX61SB5lwRuJkpN2NKJmq4RvjFCn3p/x+EWGo/VTIP87yWceJSHv/TxouU3vgh9o
WUrgQtpwHbfnUESWIIZ/UJzKWiV39YCHrfG/kSOlcktMJu6yCQKw+dRhTwMGmRzUKjS9Op21CEFy
3Ch5rzEXdnc62LdVcuC7cYsWTdobo0dd2m8SqzuQZaVsTjK/E8p/RZkxp7fupLWVoCaoSsseXHZX
+LqbsWE0JyP6kooPgMudEqxLS48oJSqeEEcJjv1fOz0uW+4EnMbfQ7O7pwabriqDIit/5subRXXF
cgPbfqVFa/MXhD0pGvU5C68nI+IKzPiru4ci6Gc/IYdWIpS7tkkwF+guIN9Qk7L7lBFGCInW8akI
63uHTuGKhb8iFuCZwDuDhf9PGNOoXngmCEdLVjha2QfvIebjtRr4Nk0ACaM3/Xu7B3jFOjvb3HFg
hC/9gaqPQao0YK5yq75U6dl7w0QzYJqkhWp8s2Gnd9tL8aBNso7Rn321E7kND3bzaaIe6ixVPU9W
TpPj2E13GD7c7NzFkztQKxNQW/FYEIwTa8NAXb6olM7AOX2Vga7jFv+oNfJri4g41n/aTOm7aJP/
gCpbcsuI0lD44BuutvRQ+f7DWFT1djik8Vl+3wzJxgPeynNh1IliqeolX2nQrmd4Xoig8U7tMWM+
47m1PW45M9qAwLls3szwFa7AnKooEUvoad2evrlbmKZDZz89Kdzs90WMRONVuVjg25x18a/B1HnI
Xkk/bM+t+zD3tB7q4OnlqYem2uiD5+8QqtsiK4ja4iSxDnTwFKp7d0v3IlfoSnhgyCgqKzXWmNDC
OEhqOcAETxDc0ED6KkezfUBAGm1EcHfcbS55esQ1cLHlvhAfvazLlpUUyNcoM8N3sPkpwop/dKEF
Hgkbs98dltJmnnJEFXETGfGLuNzKvi22QacvPHu8wHbqIByZ8cJ4Ih4nMMjXGRrHdy0TZGP+SRd7
ONBskAFBVAJH+ds/vs277FS2ow9wy4dJIEoYp2bgzIr+ekJFomW/N39H2Sim7jR3FugIDhCqwtrI
17khl30uawN15Q4R8+N5wCD01NuINeWYxtsmbWq4QDXkkskr9kDINzqTDazzqMDtYq3R0Wpweinu
kFaAFXy9nHfaFDKrSQLAmOXHvWXFTDQHmuSVqOgCCnDZ55dKsdzR/ZKPkf0rCSyvXVvV3iMVW4uD
peqjRIfKdAVnsUglx3XubhtEnRnOgCnhzL+Pw4ZQuDJN6qi41zJcA8daH4rtItSQR4/FP620aoPh
AaFsBpSoSzZncEXqbe5fDW4XsvQZ/zeKbK7uhRLznmhLF0X83k5/9+p9VVWmZFpDVH5MVK9KjSux
mPyc76Qq9APVIWi+cV0dCGcV4RUphlckFxWzNt2VIyOy2JN1wdM0mALCvtA81e9cfQ92eE9qjNBy
wIRNTkZAEJRvQryUAXnS3DJJMrs6eioVw6zeZVxHs14RQyE98cuPKTE8CJq2KWGco1ABTqVQdtG0
7n78K4RFxW8Uy2mB4F57xH98VAWJoD+G0CQDjCZ1pi4cwhXgvjA3J2uKCmBrpTBl22Yb+cpFh3oJ
qgBiAA/eXm5J88uiHcA48MO0+NC/HLIiUwEL3HZJkO1Uf1qv5p/Kcq3OzRp7g1ovZfU758nXKP5g
4zivotIe84cN9DgXuKzHRlOukezeXa7xcrxwjFvVfxTWi1h0XVtS0JKIoY/+ADHxJHVrrKUM6Kmm
SFijc4Oz4TRY9NbJv/OzqCLx7lrla7XcRqIS/fUkQMs0SwypZ5bd/wBqHS+M43cj76dxa9DbcgX/
0IjbSivW9L5t+Lp0b3Od+H32hSxMYsjzwM6D6D352XCnPXxQCPAnjOqblpv/MAJrGWXjUsXpVZbV
xFKud2ZXDZbBamR1B0AGScyyf/vU4zuksk/oUgSD507+iuYDfjaHkrx6fNF719WJQQExIoccwUxi
qA5oKE3bw0ntWMC3iMFTxaTPGVxjJDlthkpodw2U+AcBrhu8LKyayaNFk70AIai6p/e3U2M7GmNV
GPwI9lmsNkoQlfIb6cuUljRjIHdymb3BKd65QURiV7eRSpqrWi04HErgSQbPPIBsIIRc8e6VqCMW
E4qEMXrOMQlRuHU9hdT6zruSdwE/Lwsv7cproCZkJy5OdNCAwg0jDNcBDGb+NguAiNlTSOmAtUW7
1cViSrSOh72bs4Qo+kkso4W8J73PKBlNVTkZ3nAbUS0N+d1av5oi24irci+USi+k+Dnt2VmDw4yJ
V67gM47cR6IT/yMtrliOVfLeoSGSNbYR56irq/GwqqVW7aPfEA+S/ReP5hfOqzZE2suER2vk8OTc
dqyDJspQ9YBpJjfFpJE9r9JGKk5uE/5LlkbLCVSIjt4Orh9Jc6x4i7jVU/gSgjPRHkpGkvWIH0aB
GbhO2Zitof1u/GkSNEuTwnL+b3c2mEffIUQNU3swJXXOEbMT8/QQcfeWeW5C63ltLVdXSCpa0pZ0
594S97Nk1GENz1f+SvpguRGwapuwgoF4WzkM3QLU9xpuTFFKvt8608Fr0IY7nGBy27xe7C91YPus
nkjOx8Lh/Fs8zPZHGmZ+zQb95vO33hSmtKvUdBlZA82cNcpFPWv2Tv+XusUoVly6UqUQShXY8mpI
nif4nSfI+YSHJxHF8ULFLiS6hq4ici1heFrrReH/MAL4OD/vNq/TkYEkcUk2MznaUpqfS2YQPDOZ
pvesMRuFrq6xwXMPnJDtcDf2xmoocp/F5ExeBeERmK3nsx5PoQMipU/f+emtk/7E2guypP3lUVVB
REnMkUs7hTuL7FZGiX0b/SUbFvXgSS9Gn/1zM1/1/qmJRTduD7Zv3JZfVIjNQgNR5gCVn3UKFjMe
7zQSAnFdpGk1blEaSoCGu9cDxOacdOu/QDBUZoylYnrcPYOj7uxLY4EcRh4gTcjBPSJ8dfb2WDF8
A9oYJLaAgwgC9jkkO3zF/hHgvZsseWCBjbYmqcQEnPpf/emcbCIrquC11hn73uo87VV/98e8dmBp
qXYJ43vMDQ/5euoBHahFs0PGNylycxdU4akYUSvUi4imp00yInTXqCJ9l76nAc4iFYYTx1KTMsxT
2oeXU7mEFRFvvd7F2fw6SU7laTp64pMfdfQWvmZJcgeZjvjvSXQGeOdctkeaaZIP8qwukRU+TCP3
FdoNQUWxlECDAAzsZDsD6dY6+pOKRbZiz8yhPCdi+nUmlKLD/w9cEnFSnio59/57oCVFbtRlrcU4
Lx/stT9hhfdQ8kq2toJ3V74/NxEEn5WhJTSTo5nixzwFzvqvU1eGYXvWaCUBNlZuiwA7O0LALkm2
v4tYx0maHm+uu8RZ3MIIr66oSUSAosrUxh5cEkIXgap+gi9rOkItx7VoAC53wD5DNL8iIhv2Ee5o
CBw127LGmuxQE3cF9+e2NIzLYGWSNJm15nCl5beXONJiqNOPzps1Q0eqwiU6YNBKAU8C3VnMYdgq
62rRlI8CgcYHMv2E76javoN1htahktgsQReiJROcG/qNE/pB2jET3lPTB/uQ/PrigP8XjoCNJX1z
aaohkaoIpkLSRM8kGYI7HAPXCziV9xH7uUrrePKoOT8vWbiNKRkoHJxO68nuDQJ8ArBeCbxOJ0N0
DearT/jZB/3zPc89LYckaNv27JNzTNswXcboD+hdE4+yuyBMnUYaRsgy5IIC4K03JHvCTyvMo6mb
skaM0c0qLbXOIZig0BUOYe/jWdPXjuzZbKvjuCWCP/6rdUPwe5e2NvfC7YgXBNXLdW5fc3dj4UxO
V8FstUxBrEYmG1/PYZixn/InrLlvtBU/6adkze/AfLVfFYIHxK81N43QZnKDCX+RECbUUN3gOXhi
VSXCfk4mpD0lAzrrJbGGM2SZntQGTx4YR7xhDVtwseaYoOlZuwPPEZkuMFpZmQK7Oqw5b08u0RGA
KI5EUwoFAx+5UtcSwLuX7RPGTZZnUi+Ty+9J7jVM7CGj6cUWbFZSFws2iCDlqojNyDh1pSB0A9/m
GMa4IA4dzZKGDvihNct7TT7OoIzOIU4JcHY2Jm4FfSQCdRgiK9w0zCRNSsgqnn4BT7botblrWU6u
VgBkYJqhB9wM+T83+bCUqOr7JhL3hL3lnSo6AHydSyBrGguSENghq4HPHDhWdsADvRbwhN5kUaCe
h31Y5LS5ltHm5hBLRC6Y32g+2apsP7++zOE7rjqCvFLlRr4z17xaErzjHhP9DsAmCz3pRbHiWSuv
QOgR7V8s6+W9YKQ0cTphahVPXJAiG3LZNRD2C5YxtLoBbnpjsVGBjkqtEIWKisRaXIcvKHQS45pi
t78fKIarbAGOUpZhyXcxROjvQwUd/yMkcICcqvv9+Rkn2F7LZIq/yGR0sAKukSVAeGrfNI9ZFIAL
XWUDJ/FdJZUvxU908MiYRMoOApZqNVj59j57JU8Lk0YY4Bxo8AEIq/vLWOD6DI0ZnlLCNWfw0yng
Tp6i6+sk2E4cjfUo3bkzvn99+HX5zK1fh4GUdl0+R6BCYNKgfVUN1EfzAQZAynv/7+ogzyhZlJOA
xCJWQSQ2+8dXqjN8H/M/vHLxR65oI6GtpwRbK+9o904zDYXNsbLJ49EneZpEECN8GSoHdynC4Y4J
4PnHrrcDZJg4htC++Vg1M5FyPwNPFosWToNtGzmqnyU8WwH3xCgmmbd+oIejLcUGb5TrL0CxC47T
d/fih4P+FuSEDiJljBvShvO3g2Y18ltvd7Jgmdft4reOJmDuT7V0wa5tma7/ZkmdfeIc+gO/lQUy
+3iPc36t26equMcoKmkcbmT8HDZpcWUzuT1/rvCSNgGD8rrfVKlS8m52FrIOi5Ve5MTmn5V7Tsgw
9vtXYNyNUTxUxhnnNYNCHwaFlUT8byKBWOHuGhMIXGl0AOLaKLvrXLMXBKU6NZBF09ukNhV7fpaE
z5WafhhvUdD9uQj5tnkdBbLExWNwuvsFOVPwCU761CpNHa894IqCU78Yr9x/e/trjWmrdBvcb870
GFOXHNbro+7xns0yPFgTXWeMJ/3Ry2r8XdhvocyY7CT7K8ML3nJwG7PLqQluZBf/R7YRMxMkImhG
ZWp/LHIHch5Jy5qv9B75p7KAF9pCthOtOyQAYgCeKjtklkGourNXVdFqNjEyOcRE4F6G//TDQWRd
NMfx/3jCHYnLt6EdTuut2cORE3ppXOdYwoW4n3o/gYV7d5uIn+APj9Abkmt+xV2VDFQe8oEckGHI
AbBjHr6k0Xwalz9SThwnZaKZXtD6qlGMbL0Zc0+pd/Vd/MuQA9wRXOG2bma5Z9kbKyH6sNAs7dqw
DqwahH/9NP28cHZ5cT4Zf0Jgf0BvPfj6Z+jKdYcvqrZb/mL4AeAPjCKCaKgsCl1RE5fgSHFFHTyX
vSxAPotquMfxs2pL589Y23Ipr7LFx6IokGa3998ySvgXR9PZzjlxLuqMiKc7UAydSW+idbR8zD9p
eu241eYJ3X8UTyBFyIkt5wGig/tvS+Rv4KJQzDzJiyohU7AoSv1KbHeOC731ky1F1SBuS8ndpte9
H4HcZ/kbGtVcoy0fXzhxehQgaWBIx9Ek6W0B6E2AgMPmDxdcomSwmIjmyDTP/bHSIjjn9r72+lAz
iP8i4vhJEPZB3GMRxlA05zqEhbxZhD3g+3G5o1PtMiEETHe6pdYpQ1yZ+QmyYX/HW35Wu5XtnboV
XfDaiiVDnoZKnc3PEweKMOjU31dRvOweg0GkIz6BL6rW9V5Z05L4h0/LSFIu6mATC7ELHGk83M/P
tZTwg+ZbjVGup1o6gWJB/5IbhDk7DUD7qrN9L2mggtm74yvaGwe7km1Da1upTHule3F/fcrDQFIP
D8gHR/yo41rb3IicFZdt/UFu0LFSb+FlJaJBWCFM3zCAAgbrc6JCL842JbnplB0FGC0iYdM8vc+A
A5Re7QDpe+Hy9Rk+vOFctHyG4LS1XSStjI+k/gJkXFU5yJ80GAaofQFGeOl/qlbkmhsnXleHnDw+
2R5PlIVymX9idrX/eHyW7ufKHcH5ypA/IBQJvHaTbciCDFbUDpQsUs32Bwnyzqn2bEYStvj/Zb6D
5H/pQkvvy3Mu4Qjw4A1ccAvIQ80HPYNzQa47V0e4KAeuX5r1B7N4mLK5mdOJHqESoqjC5KtUpHvZ
5VsHHNNiNqgLLYh0g2qziaH+8jCg8z5HNlKg64tu4J8wEQRIDEmmlY7UdMuUPRfA9b/J6w7SawBB
dLDsdv2efOkE0UEAPMOoSLrHG5nuQOVPKHLkHiLggAUkM03NMocINKdSQnkBRHWYPGqVvbaPXKmn
AW8xwoY16yLiX3blG2PTtzHrGWzbQnypwKpkJAARl12OQRhYvd8UcOy2DjwXrVXy6krjH8E46wdb
s/3C0BPUzVrkuJQbY6AIK7w3g3UmWeFyiQZrF/RFhGVgp1UG+e0yHVhdw3NAD7Lw1pnMhHq8M+Fj
gRGzXk1igmT0Ukqh3Ev2f0RFl5dJTKGM0kDrD92u2dxwCCmB8dJP7h5WWS3RzKFmVfZ/y55IJksI
SydvP8Fs7D5t3feVNIQQ02J4C2RaiCKuTQwRhLzEuLkxWhotO7m/ap5K5XUHQFooqGOI3MIpK26I
GxOxtM2Ejs6l9pK86no2pN31Iyq3/eyEot/XDdDPGYmGHsDs5x0HvFUmvNARMuRUwm05zC2p6eZ5
hjll85SXhChvDoYazmUOpLMYTG6sEKRNH3b7fLMa2UxQiv0qfWrU0/Q5fHvfDeJo5MUhrqjtJzWm
ykfC1Q2WvsuHh7VrN4e+5l6q+SyKMwm0Ubpn/eZb3943/Tb2N4bj7FP7hCRED5UzbSV1vpevRxkS
tIuDmJhcAsF0THONQg5lJQ9BNeVYjioba5yMOp4/tN+r5hUwRt0gPGg10mtyXkY5VdSuoCk8V7Xc
L4uwzyp0796bRaUOiqMsrlAnQ8NqL8tQdvKMuEcHuSHgFeTCFbHVTzxCQqN1PHGrb1EENsyHLjt+
q0r0dilJOSBMU0zh/WKN4Z8s68P2JjKjo0hOv4n1AnhnZLofEiw+s7jtzlt9HOIBLEHBByXLhANt
GVHT2Ml8wgM3gYo4FzdPoCB25OPiNMaZNucnji5nHbvWzaekIqXrfw+QAG238kePBLWN0awaAB8H
QDlOsSkOt+oXdfD1iAnFggOJHuuWIW8Uj9gnspQGHw/jgj5wx0JoqwzHfqBwnqCi8C/Rr1zvvT0t
Cnu65R9Snhot3T45NbOh1voxavFvKohCExsS+HRpu6yLsRPugrkHl3XhDiVHIT2RNFP++c+6mbIk
ZblaEjqKG72MW4XX2Go/gpID14WiwIXuPvyZxjEJz35DsZObWiYxdfPs9EhjlSVAoujILj17lqvb
kRvxyzP44hQClmWPIovAvNhjQYT3E1mHy1Zbwcy1UZIK7bpHU2P3iNzbP3OQoGVmWNMGv1QnBuQp
twgW1qwJdVVPSupdRW3nXhtUpnypAe+nnEbyB8tpBBTuWi42boX079lCPJucKvB1shiQqSqRxbBQ
B18L1nQ7WzHMkIZV/BW1CuMJWp1otcVolX/Er3pRn+h9xDnj/TZyizYGLdmdeErneH74cpj/unCE
D1D2mTIMkz8weqhGQZIQxmJCX3GVs60FRb7rxXrm3cqF9n7/xHdb2Eh5oqnpgfURIpgwaI8O0beM
qn1yVoTIE4fjRU0rHgD4DRpt6psPeG+TX4Emuc9/ASmgkNr65QBCk7IG1haTTvv9/4hn/QH47aoy
VohgA5mX9zx6UWyoIWl9IXjUTssMr1HiaX9jnIWkcVAp+/E9EgpOhLdo7b/aNxppQyssMnzW3Pny
IbUb7D88vH5KFDuhVf2EF1iBwRBRxUNjDGL68E/cbXxPsPu/3/LP3mfgOGIOL5/TPOfYBO8fMxj0
4RufWH/GN54NPLd44c2s09402++Wfvg9zBPiEdjOE5OJMrBalSA2Rqu1XzvvWX7ZOMGMBtxBhAL7
+TFQBpJopZoWBf0oceCS+OtO4LyGRL2bd/Ee4Q8aBpb1g9YVT3r4UeFH9C3ishPouM944k2tyOz8
grt8ORrPcA6PEEI+9MKqfwFTCciNVmVN97kceUWLsbmKfwUbVvuypGQhVRMudfkslBjc4gHi1shw
RJEUsXkLtywSqKy9cWURTBX248Rs332VaZMOFVRcp/74AsoFf6qWX8b5fh9rdtvH4ZQD1C9GeVqT
JHTBiXTXiRvh/ujP0NDc8eHZbbCDNkc2h4VM9rBGdachnxTQPoehXa5AFeqwr7DDvdcEQqAWRrSg
wSI23hGo79UepDcLKfjbEtpXPGQUN8iPp4xSyGMRBLg3NPGUI2ugrocSIYtdltMf/O+Ay0hSX10R
QJeQVp3rGBx3RY/LUx8DwjccmOQJ2jCt1cifCfmnfCNEe3ApJU7fz53VJvbtc/tuauy2XyCwBk3G
pxczuJ98ehgwzjv4jHAjEBU5+baHWY6sMo2qlHxzu0X5Ky899T1YkjNJKdnUCZpHbZ4W7KT0kz4g
zlgo+kIO9jk1a0Y3qI2LMnz0k05V7fOjT2SCjsVz25u2hd0oS14E63BTd8p8sZykClMLUnjpskk5
XS2gh0nTY+aVTimdhX164Sm6RE6wAGOFg8s11o22B5yKPHKovCkuzaBjhJLmtF4+uWKs6vL5FpYI
H/9gUQWVsr74awwH9z8q6BODlePJUBdnw2TQbAc2YWHywT1ojqMQmwZ1xKZwb64LGd8iJ4ML0wm4
D5te1zolhEXBbOYf+rjwsNCXPeC5CYyR49RdOML7YnTFgvkvjg7OBNJfnpJ20WLSVX+99hjyVy9z
OLNbz+Nzif0lU7+NYr2wUgeI1IxFu+ljRoCB2pTqS43lB60Gt7Mbcy0JkCJgjyB7ohtVUcpsyC7i
dwOwRNT6XHBYyLAhDRkofAikPHVo1U3g3syEqiPj15FomxwgOX3RF1D9I7o90hnTv3atA1xm2zej
eoCz1dCSwzN9qgvGIQO8X9swHUxZ2DYbygRxH+kLIU8yCgcdsHeTDwM98kGF+9aLlWcQoXR5JcPH
CMC/x5N6m2RbZQWFKAbJgTAMRyxnL1wXi8x6bLtkDLLUYKa9AETLcLwQamRtEIfFdQ64I/sOZ+8P
BCDrUg9bWzzpIoTl6ze7YkdxGaYT0kbZwf1oHnQOwIvlzBZU+Hfo9tMEYq4CGn36UKlr5qpPcJ6S
3vKX1vYbXFkXR2sBvsh3/1jPcCTmQ1D7RSHzLbj/oaI3b9RMDWS8u6C8MuSpL0LE30IAXJJVKPnl
Y2T3Ela+934ALHXyo/UB+Ib4wm+Np9zB1U6MzfdHEjTBXAKjIdyuyToSpyiEZ0dSFN60baJnOess
gr7mx240xW6DTFYu2kzrR2AJmSgeGgEzPp88nw5MHv3DOeboljR/+U5mVk7UwjZw6PaWjhEjvdFq
vrQSzTCHx1zCwPGr6AV3+ijLihVaSK/jl69Xb6KcXbdS3s1G/VHWnf5K2Q/pb13Phi29pX4uguiL
j7krveZ6ZasHOfjGoxikvcvXgyF7ujatYN8XUUKGalsQsfOpXZ741wopNA7CpfuW2QJir6EcbyFx
kOtNTm6CmcKFIfIDKr2E4mQnlBKMmhIxAm/Rz+z5dykGEJ/EA8QMfySwYoNE3MskhZeJRvk1EvFT
AtOPVc467IfwXGsyZ7lCIh/Sub+XyjHyJ31KcQEyOTIqsFO2xAapkVXd8FqfRfEjGrSd3RyvZJC/
+e4aWqZFH04YIJUxQDbEb2mx+jr8TM8MJKhCYL04dgzt55lvi2yro+MZuDNi4zdE0jjtncs/k/D/
/mrwFlx5tgPwe2RkCg8bliritBNCEK0+9HEQvyGf2YbhCLWNcclrGSsqwadjzH3HaQ4ezo9QYkvh
enZl2L5OB3U7sgUUvF3k9nSO+BaoApkjR1cW3znOW22BOnTY960gUc/wCY3g21uMU2Ca4GjhmeU5
OfMcjbJ37tWtb1s1+sCsNZa52tsWhWXLD8bSTNzcq3Ix/A2t0eyFAXRtLhSI84dC+EpOwapC7FWz
MFZdVTZLq+oytmlJN2HsjEKy9qbeQ8ZSKZ/MIiLYz3r51JMw1774aGNhtfBW6EakLi8aoTsNct6N
EeD7lCiJc1bctzb3NnlDki3l9jq7Z20fw6Gil/uBIlsMNvnxtBTLu2t8RMqJO43trtwI1BxJ9Tvn
ylinq/strGUZqB6R6YX+TW9/iZU8qp96KkKKW7t6mlOE6bQvDYCf6C8QEseX0jsrh3sPoMW0VFyE
mUDJsVYLgv6aQB+3tmQl/eFEw+X40yL5VSmUvK7ANhEFserH/xRE8/GWuNeMWml89mDOiZAKHbE9
fVUsYIR4xKKUivbhWP9tQC5h3Ht3/DRdzj2Q8Rht0MCT/8JzRCGC7KVhWqiHqESR9ViPykm06k+q
DqkfnPLfqx7fN+KIouG1NDyD/OnUDEp7OwCDEGl+iUjySN0vWZOs1maUIJlZp07Ejc1UffuQ6Okx
u4BYQqvv2Xzm0WJ5dM8zg2077UbVj9LOraaPK03IhCx2gt2yqAZN1ot/R7rzy98e3Jv9hS7gTHVE
jt8ulCI9wNSIpKxJkbJqo7hd4faOnk8RAjXNDUzv0H9tvEH4lc/N0VbZNgVdDwD5E+lKBphGaXA6
OdUdAYy5tvUZ194zsSpHeZeRFTHKQAAWRWx4wrX5BnzHxN/STnmMeKhrn/pqOdgvfJElq2MtUfd7
fXcJdkszjQwJoeacJiz0EHDFTliLbImSEyNLF3pVSnedFMcYhUyeUDavB0Kf+ZWQqwsysHHoWZUD
qJpOECgB/Psvm0J+klihxLklFt+hzolwR1U9qCwRq2ayHNNYrwuK0kVJH7tEfogN6mejBqi+6Vh/
Vp/FISFaylldBB7H7zhOfRv3B8Fqm/obye3ee4l07r61BkY/2mBO2E7YqGjlpF3rIf+iQGXMHEqS
epXh32Gv+9SQ9mOk60rSgtSSQ22EDdif5y2lj9UPuSj24VK/U+MexL/QPXS5Hjcl2eVqlj2MxHu9
MPTDl8ggKYr9adsTRnaj7Dj2CZ9pIQzyytZohSL2vONvKB1oXAgP1zCm7UJkFBecjCpK4kkQmV5l
GRAhAQXUrO8ZienB8P4bMylBvqESkYhzDlTq2D9v2usWd5MCYDh5CfuNDosk8eibR1vt/iuIRGRF
K/4Vjbrd6jIeOpfrOb5Gqz/vUgu92PsEgYNZvoVkJ7CXlG8ctp889J68LRBn9XpaP8KRo0oZs+7l
luLtTVuhYaSEEBXKQtsKTMzk6nVYn+GZhZ73SGaATEL7xlykvZR1vx4tWfj0ZChNpTVWC53Lgb3F
DJ/z9lxrf5KMQRWkEOF7tYsQlcOlOp1emFnUvZSwCem5cp02rJYzDKZ/Gm0l0eWvp+Buq3lChVMV
fg/89u5Peak+6GfwlvaCqcsjr4cdIatm5tt3bUHzVho32DYxGeeYe+UCtY82T7cYO/isof4XHYxC
pIC/athkWhcAZbDUlKF/gkPziA36/SvxZHREna8V8fWRG0NLfMcVooOg6N3ZhBROve4i7FJOvtae
HLqz7x0ZX52YXh46XdFfk4X+1J8ga4Gw2NDZq9th6ExkjG4LuxPWzw785sRc04IiWC9ZNnVVN7j7
NZZtC80FLsv8lx9h3h2d1v4wfefcQbyjq9HWLag/mUhQ5FsAVXfcVdSuQ57nYm3zI9GTTdPwwItA
ySfBZc8NfAgyNY6x5/9kUWMKGFc4s0J7Qp9Wn47vuNGEOJA4w0zk3fnhMpSE0RghFkGNOM2LGKup
ffTAU0yLFg9hif/0peGyeaKxed3n6ui0pwDoEotoCacPskIss2CrjDl3ty2nTkdlV7i/a1vGn45b
L32R/XiwA8RgIpV6eucY4IyhbGJAfaguMVuUZQwQGMeHkVdbrUeRGOqLQwb9A3nIofXGB+cSGLBD
oN+AzE3fj1zYKlZBxyD7Xen0YuqWY8q5UCdHSjZ+3oeRT3T5LuBknn8iaBCeq82hUHmOY9WO4gCq
CjB9o9EmPBbmk9Y1y2pvX7oXkiTM9Om5caGb9scIBpKI4pU1EtU6XnrnQs2cXvjsyGB91cO6jkdA
rEsV1NBNUe4gtQC/BoC3IUapwCbSi1CztWs2jCwMTHSwIB5NbaZwTFsE4VN4AdUW7ziiaFEXl+/T
teIEqol81CwX+1BuutIrbJnnagSzBEFn+y1MfHFWFg2iH3Bx4op7ifPCfgDuYfwCXpr+0ES+rb6M
jIquKotP2uovAWvcsWelxISGYrZCVXEH8yfClmYFwO9E+mdQ9RzNNr5d+zPl1p2mchWq6Xr76l0K
ceKv0q9sZItGr0FgqQjyU3mMeNHRrw3Qh0wiV1B5oatSrJkQ11pm5uRPh9IFAfkvyfnZ3JfLYdaB
F+IJ1s4h4iWC/y3kxRTvWGZPFiTEC1n966rfdJozpI5R9lT2BNL3kwDxNgGJ/3PXfQuCdC8qW7tM
h6jvA4NPKrZKrBPfxywLu5PFOOjObj86eUGZqz6Qs7jxkam/xXhL2h9Y05SjSZ254jEgorPYY2dT
MV8mi1DcPgzqDZMybbD28a3Cybq3atH0dDIYW01fjz9vX24ah4IRSyKF49nMTS7ekf+/ONqjbl3y
xCwDG/K4rBgF+ExJbHTT9u8H9My3nhUEiTdL+uJNU30UcAcsOiarTV7zSbrGT7+ysvolXShu2vE7
n9RpLaygVZyCex4dwppBz/yYCHB2Cbb6umGaweBA14QSMZ+bbv1n3PjAHVnHwLo1AJ8W4op1Yu0i
A3NMaooHKzQeYdwqVxdYhVI7sHYurAi6RzKv22V2enZjfTpr/Io+kzYhQVACDB+nFvrKWIT6FtLq
k6Rx527jyYOo6qeKHlqSrmylnallMriz28nf+SGIOKrVeV4Bhjh1dl9FyRRrgG8pjrQkLH4CHYMK
0j8df/r3bWxB17fP+9Vio7E3Xi639hDmWiT272bDzYhE5q3sj02IWBXoI7kLu073hnDxo0+8LLY3
a9l+MZhpbLBrO82pYtZughugFzLtkMIEXGDGIr2/E3qlfWjB90xBIL903woCUOhxWoj0GnC599dQ
UuuYnbkKFL6GydkRyKVVhKjAq9aEL5mjlj58WgQM4l6ReH7K/5BGmrEnShI76shaPuDdl7GQzYTg
EFhnopoXkSiFkC+RcAmx4sCvWV/VDq9MfpGG2a6tgbiD/3bSNNg2sI20e8C7CDAS3zZhZxdXaYNo
YdFwvS56AKY8JElEztcaeexzmA2Jjyz2CWeKLLPa6WrELVqFG/QBwJ7F0uVX1sVxISbDfJu+6Bld
UwLY4Yhny4tHu9ygtxtMefwq6KWjQje0NZKhTbmaZRrZwrthEc6XpHfDMEzQrjRoXt6wPkrpEpBw
06i5Tlqy/PzDk5/5A3B8BK2mrY90MS2Nt33mWdNCQKzUoioHFWJJKmw/uD9ybtMwc4sxv4XSwZfQ
an+wSCmuu1OB6D5x1sO/hJFxMOaWvxArBRXSzbqzW6sdQIwS2kNyMIMkYPM8a6m8U20VfeC0D18o
g+HUFFpLMikKKftv+3k62yM7UuqlIjAVPy3OPTGbAgSxhJQnCJ3ylA8klbLZMZwQSFV6KyI3eo8D
W07TNACh8ja2Ccfeu7YS6jOlUC8I8XOBV13PcED78LCB3gpnUivdsXdQq1BrZE/+9UUHrMVV9bPq
9fCCPUMq14k3oVEejIPoJoEuUZ9Z6LaCBkJp6OqiYhjylfBuFA5huUy5oL/IzhiyjtF5W2HEoAh+
P9IO0iDAaPfmb7cI1LwY6bZ68RxFcTjSGncboinrznKaHiaQ6wsQC5FktkJsFb8iQ7l5Sc3ZVCyL
gUJ0tTB0NIdP6g/daqesa1clyAzE0yKmYgSYLydrUnYY0iP7jHRKzCZYJC38o3RMdlL4ujcgvTp1
AuaIi0eJpZ2RiPjLie0zBcWfeu1/hoECd74ZxhGezTDggVVbUzwOUyzBYNA/LiAh0fTL4XhD7qzi
kXZGtlrm48eihmPvO4hLpZxPg6YeEGeyLq82PvQ17SbqWOjLdgxk02lIBvROszLru2C6Neeg+hNj
WFFeC6JYsfghMrXHtYHxngKjjjtma6Wsv0lqIsLJ19j+dXbghUOsdN5zwqQd32gwGMTBRFAKYj31
aTo/6Ebw+Y457xwyMNO/3+xNGDySLlMeYHh3qQtPUrTKc6EzAjZ8jSKp83h1EIeRi56IKtyEonSw
GS2cKvixDJVtSnfAvdS7IRcJEPPmBBQU/6jEZ2wy+puHBDGBFBHNxOVsze+91BVh0BqMLew4mM/m
9TQss6Lcb2HLjDxwSdTFx2/xwSAun2xl+uy1zh93G0Tmy+EkAzRW9et0bwr1yFZBAQwAKaar/HSX
s47GlRAjZHGwhJjionn1XD+TPw5ROl0MjfrlLt6MT+2olBKutJ7m/YmAmHPQ08ER3zBax1+XtGoR
1/sooNtqeJrdIxv15ewV8hzYNrHinhHxTLivhQD8meF2grSBweFqqTGQs1rRowlMt0evw4GSyx+A
sONsE/3as3zLrMkk1qNEQONCdY97fndmbWi302IflRSB5cdPUgzwqoy9pthMWDUvquRSdtLBFkE8
cpZeoRWkkRyHQjZZnR2Ua9g3g8JL1KHtPBo7Y6pbf2ctDyG6GN7YX7FHyZkwaRZ14w22lHxypZTP
BZlticyv2MiVaEBFHNBQL6mhEPyXfnsCWhkYWesaouy07tw2A0POLV44juCrV1i9mwBf19fPGYbC
9MYJ+eXNfD/d540Ulrmtpi1/jEv117y0AszLyY/OPSQdf9AWnVFAc/wGgsOt9QavyralrWzz47kE
j1ge7DVcHJSXWwjOcb+Gq15ZTz0kjj07wovq4CjLtiFu432ez5jHWLvDxa6B+25SP7q97mLtLE3p
CTb0MImkzkP6Ll1RBRmJem/9pc9Ub42SrZD/C7hejWsDPNR+ysd9r1FN7IKYrNpLJRMppD+UYRCg
EKYfHGmb8wBvrw0yuBnH/dlXqsz/PWSyzDDLYVMy1iYURxtgL+A9xK/spCVJ1O2XE9ifS45t6PMf
IZ1J2CpbDOpetzv5tm8s4xkVkYdUGlyslQ+RVQ6UptsmyWQvpZwgXbHKNJpJ2EzcByVfsCBi+dXl
VqBfTD9XT5qFNh6Ptl0GgUJY/STaQnK/8udyCyQMjzB//t+kP2gyS+QHD65cxsTJtLl+/7vNMSem
1Rvnn8iwcSC9tql0M/E0s04lZXE/HSD22JdcxiGT524dSvwigoNiXXTahviV5KiVNTyOeQr9qvId
wMdGzwm85ra1z0h4QMtxGvCHwQtiC4dWPR3WUaA+XVmNTNwmxsIoSgYdzvsabCWwISrY1Rb0yv0Y
ZsUO+ORk2LdKKmHF4KcRz0CyEu1OGfSlrVo0kNyhMHl09JxOXi5y7hcRhUAYD6Se8hX1di+ebcOd
o5JotdPfotT4peNVuNTnlvLe6TBSKLNkqaLcSPZp13O7e1t+eJO3cjCtAaZoDa9C8/lf+YdabMIk
zLdVSipx9q9/SJ2oxVkxL2+PNLOIWWtMMK+GoEcMmZrsyzIzJALv7fbqVU5gGPp6J+QEjMN04HhS
qUlNk5PfTzmTIQpv50c6Kj5OHsfwnBqV98BgouwhdrYGItc3Plt3an6PR7/WRWJmxF+4BTGM/hd5
yqYgHss0j1ErfObMK/3/8ifKONVHqISljp5/a9KNhmfguxdXVXTy1I9orRvziZ85eiZRR4K+AegY
BnUXpU5mbkFYlDft2ArqTve81MwSl4WXFdJhEKzVscXYJZ01lJHLW8BssLiRElC7twU3mvEiJ9Ho
A9iUd8ZegsbF1uzyHge2tlljRcmGw8R1Ng6M6HhmceHLTYANyz0eNQQkj7SA2v/faa5TVK1V1qfr
snZoenPccrTFquqc0y8o8h1V3jESdiXV/9u8FfNPIGIurVSAvuguKj5A/yisK+iF7Z7SxdAHWfuX
WrjLNojtw9YWkk2xWQdOL7/Jk0tQ4LIo5fXNfeHs5fnhKt0X7DuI51q91ymOtqXTB1NMoThIBOB7
65hrr1cyH3xZnygFsUPkIhfgxLS6xyh/hX3a6txAlCwVSENpCP3dZNFcoIm5whwNTPbidu4FvRCG
IalztyEmfbtz2tj+y9vODzQKaC5c/ihuXtPrjdeKoKy/KFKqMrQAeNWpFi4lf2NU6XcP0XtO3jQO
beShydofCV3SCF115O/RA2FEshvS8TZ9CqbOzShkDuwXFQaGq4o4p1Do4xYZFL9W1yoWStA4sOkD
aEdC7ntunUthZsIc+XobKVobY55BzWDYb4DdoCKkO3d+dvnKbw/lssY1snB5W+RN+6imt2KD9GHE
4jtG1WU/nzoUBeSvS1aBFK9tkwYHaTum7JlRgziaQxtPb1XIecl+H/d6ES7A7hn77igfwAu3f/Re
/LS4zY6rPQ+gkwyil3+ZlMmvNU+sMFuH/UmuC3bOg4tRErDKdUAV6kHDe8wLTqOE33G5XCbKw5/2
co8nvY5UbOSUIKy5TZFCIf4cNCHT8yWy7Jqq6t7eZY5vESjKBtAojUQO0EssdLE+xVPOyjvkDgGy
RsrsH3hK0eZO1rfVoYSSuyLFyUcmNCyvEbzpTobd80HuZUlyr74ELSYDq/8cCh8sTi/yIAf1snlM
e7H/QZfNk1e9H6kfdoDvnf1z28PJSikXJffT2TNIzXUvh5JUKjziE2p8haYOMAGA01nwml3CisZN
ndehSRiWLs9bd05kY+AXGTSNXOSgSi3nm+Xg/qE6yutWcAHZbG3VjCl7TvdI7H1QG0/upP0px8jp
vtcAYXeSAsFnQx9vswPI/+3dtJxar4VAyxmh1Z1zMbjaDfu50hH49D4BeUeoHfGkOD7Wf+3dlwdZ
lih0YTyM9cGF0qDNCklbQpHNlc5Prv23cnkqwDZMk3h1kwYUn6ZSjRqGKEst4msYD3IROyXuaABb
UJD54Zt/Tq0BSdrFFilRvkzScw83IAEga8oPdwDaTkd5IMHn2AB6JItTcSZv/bnMn1kxFfktfDVp
RRqwt1HxDzHS0HJuRzRNc5Y9Kx943RTzAyYZvIfmWN8UvwHM1ofoATOg+JmA47fJfAjFxcqbOoNk
CgddNUA+sEtXNEzfCc/i1zvdJpD1gFR4Ji16m1fhW25biaasa9xlSERSzjF/rSu7j9RtfVrPsYAO
RGTQO3jfkMJzVtbdr06y0VqsTimnLx5zWBzfecBEjMqXlUaBz3HJkvM5NmHuBAP6LKOZ7CXU3ksn
9opiYo1g14u++Mc1n/bEI12hWKtkkcYIezF3yejWWqljT2H5Y/T5LOce8k2gNXB2CS4/jhSvP6lM
pXomqn2A6tVpyf8Prtz8O+Avl5pEYkk0iLNcepQU3M6CxRhYkWjwkR3FOjL26Au3umNVIQ5eLJa0
NroHoLR9GJtFm2j8H0UtN3PaJR3Y0hk8Jjkj9cqSzyFgDiT4Vb0XqciqFEl/7/1/0TcN0747EbQn
cY/K+eHFs9mhtkukxyjWXnow2e8NuovOLp3uK7q7BXhpgfp8vyAQbiCDD28zu6RC4Z7wqCoQJmP8
My7KgK82sJB8thhxIkBGPbrQAM7ZZxfXnWhFIlCb34o7x1eDX4lBwSnWEuSAdCwvTiSaaB9OfO+k
RugaWlzgXO60LZliczK+melUAYSPIOAn25dYdDrS5PPevR1QKyFHhidQ1b7meCTOIH2Rmq3AgoqS
pgeQGp4JmKUp0wjZGK3mdFsqPYsl1nZ1sqLXm2kV7ckF9ONF0IWS5KVZ3nXlridXXN0iqHYic30H
ew9hrHdD5p8ElYA3kcRf2ZYvfYmVAjVObZID7Pu+0wmzFI9vp/n2PdkmHkGoERtDcnHl15C96Xj5
UqUFyMEujj+60R3hNqyPj0tdH/TdQ2AFD8hVCXMrGhJL9fhWeenGo6C5CTRYZxOx6EVuR1OOj+WG
ZNS6OTZJEuAehlp4LEarfyWyyr87jAHW4stOj6dMzO8LTcqekhuU/97prSK//S6kLq9i+PeR0Ei4
a+Rc0AJ8YXQBg6pYLZrXLyJNcKqTLEg4jRUAkQlzr/MDi5RMSNst4dYwU5rgLPkNPPjbEhA/7Fpn
cgIydXMWdi8/xmLC2bAAUNLaKeNcJv3RbHsBYtBrYRF5zTAEbHTbkUt238SvFzqo1/skHk7EfMq0
ucMBKhmPVkoUDzBqkeHsqAdvbNU6U5e4qiPqT1PmIUBZ4UlUjGqh79DmnBCzrGXibHubjkyf+k9U
GOaDsKFmhGg72FiOCMjqHUTfy4Oi2jxdlvgNO7a65u9qUuu3klC0fo+rR/9Rwtx/btHOzOVxblYW
FIRCbL//b4AvL0FPopQkWH/uN404roXqtRLJ1Fsxs/fpAfv7mXjaIMBQd+DPfvgSC9/0Mjsg8Dcg
YTkw4pArP5HR/Xqki/G0ObLzq+OxDGzUNU7qF2MjbUFGQH369xeOi1KKl6iB10vtDTa/XvyB/hAe
McDiEjmMjn2eeTDtdaGY385bn0cl7VK5bjwplBqDPm3g9JRPfeEF3fSVQ72gn+mFsBrjNjmPKbNo
5dYvhBFkHSFRlBkXfRkm8djcpkqJ7hclKsefiRsZx5T4sEb5PydIV1eBT9G1zgof5xqNEr3qLh3j
y0LVmlL1M6m0L2alBTtUzjL0RykiV2EPb4WwOjG505Xc7L9cazzjz8rnHVl6bSP7iZ0xXdApECGa
o3FquA9gK2Wx1ksy8iIuGMiwy/ktOJhmLwJyIU6Gn+DP5LE5ziTPhjapTI0XdM447QSARnm7s1Z6
9K68kl8k36qn3luLztI386Wsbu9fv00NF7N+AW8dsAVpUSxmsuajDipa7CbYN/lQrWp0/QFAfjRB
NSG+hdG/9fIah83qNwGH/FLZOqDRT3o1FYxVAwd7uE3h4iUSzmL+tpCYYz2rBBycg9p+3Pg1MJAI
MM4w+2lN8/6pYQulJMGkunRRj/9AEBeOVaTSlxN0ylfMfvO+rwtkHUmz234qO6DWCfdhrrT283nw
V7MCvFrAuDBnGWUpbZmkNdYMu/bz9RqO9pwqUTuSAsYD1074dD2QYQ/0jZcDFR3xQ7Ju8Nmclmxb
OyRIeoXlWA/gXSWQLpSy6gkcZpdv8HbP1wIZcnaL9VSujnuSPImN9xmoIgcOFwnYo2WsgRrtpB6v
zSr/LlV/a0m6c13qNcAnKkTo5xEyry1Rzkcc+gwcdNcneWAQ9OKdgc2cSxqmhH0D8zcMD3abAAMl
NmB9NJcSaKbnwv5hiKmSRn5eB6iUIvm8FkDV3ocbTST6cZhyhl6NgBr/bOhcDYPZV+iw6YngyaGy
pb7aUDfRhLb56nPZE997XaWSQWp9H3M0/+0yu1VNIwAk0l2jYNnqeZR7aQU4+4j6jlO6XBF1b9sC
eW4BZLeGgC4E99SgMsEcwZYYCrqQBTWS75jFZkYBgVuTdSQYv2CZqwva2XYS7M75tyzQnELcF/ym
umANr2L1ZhV7hNje0FQFhZIzHnbMoxMyRiBpli1YgRQPbAE36Uh3pR+HooSYEEKFcwii+Z5uHNWF
hcJobHawwvfOa7iHwj4pB9ARXk870CpIoO+SyekGtC/w9tZ4+/ZVEktYYBMoakEH8gJqQSAImEIF
NpCubgBJplUuvna/zTUwDPpdSYDlHard9UHcFYs6XX+wrzVFG2VyIbgByp50fnt+7EiiXrvnaqpT
7E29DLvXzI3qTRxIXgp7rhMEBz9qRkS9GX2ndnwotqbCIAkzV4p3oQE3bqFH53p9uAsyEx2p8MCu
RzIay7Ut8zHypEcbbWMHMUbG2nYChNzb67kgivmdxFUQo4d0qLeK8oJ8Kd9Eu19ygr7H/j+kOyi2
9eVWX1rfn1D44KcnqwO/+ofncmWKxVeSwI9gPzQ+J7/YQ7w0zSaKE+C6lQH02KHqWpD4/gDQ77jS
n44XTECrKN6PAAl7macxeOEqw10jKoWDDWuE/Kd+3Cq4plliemr7ULubKhgrIf2AW4Vau6v5ZPzl
L4CQGZNIN09/fAlQwZo+LvyHBXo0UmrPop+fDlFZAtGqOO+0XUArU+6/v1WSFYp/hQb1D7a05uAc
bkmk9qLkrJRTuqkJMvTQ95ln9fX3YvTnyqJ/YYsXeBw2VWtz1d64QgjDfRbyRo5Cw18Nzt7PIgXZ
Og1rHBtxPxf2v2TZmRa29/tW7BP6ZHg9wGwdKnd7C1FuEVRTyKazZaqlpjgdRioapdHX0ZUENif5
+akSwZXZaIE+s8ahHIZRKuwOxSzqDK0RuxK9Y9WktNKDpRtTkxt1T0zedGVwKVZdUGuowXHq+iEO
Iw71qAPynYS+GORl0DXaa2lX5MdFd0JHh1pYvXqyc1dM5BS+CKcJ9vATeAXfM047bPLOBRiU033Y
T0jYIzpj4KxwJwE2MIUImB3aYAUTYnNgW334uHsG44wh/bSLVesCt5Q6b+FUTUbUk5KZ90CXpG92
XeBzioDs6U3LqmcMbBe9RFJfSWbpqI/GWKgQsLisiMzOxs3ppHUs107jiTIiFalihapOl4rJ1BUy
yzRjeNzEM08GwMTUQttMIjlx3/WDt026usxaOwEjLpjVLoeLYioSUGLES8NK6qtqNu46DHE0nAi/
K5Ukqs27s6gV+CkCSOCc7jaGDINjcUfXi3cZLZX5EN0ZgD2IJV3ZjSq+2e744fP78gQlxfE51RYX
5hL5tNI29qV4YihKLaoHX9ypGGC18uVoW86BXpb9MmUD/zyhXN/1uNSpSxk1KIHyCzIQPdWjaODY
A4u8IZfjiu8JdtYl1EWyIcxPOt6M7pHj+PK8gYuOyWPslurDXhX5pfnYEaeEPBZ8dhSCmy6hCwiQ
OBGCtLbuIbQKc9zhdohUrVJs1YocYjm2OEHb7JNCVZhiv/3MGAQ/pPFU05tGx2acyFoGH5SMqV2K
nGs0VL05J7utuNToEEETbmLi1Ct2QEW9XeMBwwWDbgkCZ5WMY0mmQgJtIqvetd/yGmsujSKuQ5aG
1dhZj/8eptGrEIo/y/Xgd+ArQhriXPCJCvwRkDbZpPrMbRhlPO0i+1KnmKhOFLXpdlimpIMJ2nXP
qbLulMXCKZUpyFX1ZZn9oxqgfHW9L/oFlhNTjYETNOltobQ28tFgsg1R0T4oNkrUuEft5/ybihq2
sVLTnSYlVPM6NVvlP1gaLTqRAVq/JXKtm+CIJjMCx4UvHz2ATFcL7+d+hVWyp4Uruik2yjquZkKp
GXOC2bW3q61cgauLGZ934sjHRCqw71as/1dHlxZwyaJjBvqVH3MpUXeI1qvBRr6oBqy78GDX49Q4
Whhjh2f7G+kouxsAVi3fSWrURjAzbGmnhELY46/DBKxWLPKDvcMEmWiIGB4eABKyEuSqe8sZGZbm
te6W4HRfQXTMe6TboGlsaVupEpOrzPq6kAGzayvS/8n7beatQ9gaJANgTDHuOBpmU08iDM6pCukU
SdTrGIyiv0NLFg69j2VQ52LQCSDx6R0AUSnXQ8gfudwdIM12BPayBGIJ242iPpJJ+q2e+1j47WLU
JB0+/7Vo8lBP4/uMgQTP5y7V6h6YH7FWyHxBT+QuQ7VaPQ6nHD6w5HVB8noMghIMKXno6KIklHdx
t7FEcxivraRtNKsEkhv2KEmpTYIyrqi2fYpl57EA3PJIfzDJx4RVR3VyjItQ/wkVTWZAYvByOfTe
t4I8tRiaEKJPKrfpaRMvj/3usIZqKdnqIka+sASbZPrv8Y8RYwMWy+Aoh3XI2Qv4UeTpInKMZPn1
Kje+dHz2PnzWCBp5Ary3oCYnkHW38oUuv1tecRySEpJGXK4/7i/XORr9f60KVdmzpz9MqXRpyb5q
V6GOl9CLs6fTRSjxABKYO2MMptI0Q5zMEKv7Jxd2+pIyJs77NXLi2LKVwY0Rx55kti70GdBVTjG7
Fom4yBSX/k237d/JCitDY88rDKYW8v013QRec2LNY8lw1qTPeu8DLGszXTiiri+f5PQUeENGtb4f
jTMSc4t98Y+BVhtVTP3zHMAeFd7U52TLfV7/A8HVsPm3PooAtGWus51Jv2mVxA0hgCGbNCRoWzjo
2XyEEHEg9Qr9CiKavXteBtmmmX2z16s8015kVNlEz7S8vUZTkizJnqQQoqYp70bRN2vhlLqllrJ1
vzsxqzuVkzRuwZ5JlY7DurLY3d8sgIn7SosNGkGSSXIQBhzxfOXG4S7vOZUNBg87BHv3wmx5N14L
2vkFG4AAJhG2SCQ1ZSWvVMS4aeis1jgywHoom2N6U302BhuuWubEBd+A3Vv2RQvQPAQOaGY/SWad
c+usTUBRIqLERJnRpeV1CLIHDKindnynvyhKqU+pFL1U6wDziOohLiRjcF9fmwA91h0JW6gtRuvo
6NLIIqXlKmLGnrAyKA2BQ783ge0BbSkTI6bbgeQXDILV/bDXjoJ9nuFo84cZvdix1XdLMucb/tao
lqIvowJK58aKhMbjgnd/XXKdMv+s6w9lviPQyikDPVG/Ip7AQrDjBRxQsDFUdEpEoRCbheXSlCsJ
3hQDKdy11xaIbVE72ol5LC1i8WPvfEu7GygIfR5iO6dV7gqpyUeDXnPxHGG+zZMHzLPWllveQoh9
I7Le61qJK9N8RGuANv+digP35U5sPrxpgoyoiC6hXbcUR90rnPW4hIazE08KVcQLmgpDTc+gxUw+
k2WeyADe4B9j1nbBS2TPN9j6lARCDqAWsLzPw1vkI2FZPRUM94+or0Mt9IvzVZOHBhQYMs2NIAhR
0Xe1bqiJRxOetvIMQvl1GBF2u1ktNIe8qg2d5DZY6JGXHdQvULOqrSAqpgitIPCIzbeHklC8dfqz
DcnhE6/1+h/Bs8CKpLgVB2hbNtml8OIUHEumL/ruW6pPX3trlijcoW/jVsC6NsRq2jnHPFnwO7qK
vzR9GBH5k9k2ELlvo2mltLNlSifYHJ9Uo5dBToDgR+XZ7MFBdRiyS4uET7xJdyRhuCuousVD9+WQ
i/I1EL/J4g+8ZPLU1T3+4WfOSy6mqcAUG0x/U2SKXlkdARZkmDVhB8KHtyvT8Qg/frwQqeTtZOeg
u8dy0Gkgi45Yy5WShbZEZYX0PdwJfdY0xCp1LuvdNEhgF2z+AuWCCl9orL+8BMXnHHkG5cLM7c5U
JGe3jTBdGYW5XFLpvzHOER9giH0Cun9EOBsV0/wFn01LaFKCTp8NIf/tIEWxu6x5Qq5nvUwDFSnZ
95DxFe78Fz4LKJp6zE+YCGH9Oh9lBupl1eWdzVIMKEqb8+mLLyLGmqkZlzF4BJIKJHgTpqp1t3EG
Zgh8yaMtwCcyGVJ5cid58FfRev1S8PtpgPfNfL2NmqgpCGAaKHr0mpXT5htfQyMjaH2G2MuibUbE
xKklstB/yp6negy+zzCrvy+a7edt6bbdD/437437AU4caVsi+QQk5dCMVL4lxCA//vuybIydAbxD
RjCIgVlSaC7ehWYlVUNK4ItUNXmoXgr5Iwkt50DObI19GlWdc33Mm+SsJfZ+gG4Qb+as9I5LRbDl
Wuv0wLh1uO+YFN/yUiW0i/vo5zePfFPjVdbiSQgklqWMV41YijlD8r3SrsOesth3Pk6182n613bq
FpiLgjGWyXb+hJ0UwEffsyHHS5SCiOGW5PCV6y2p2WR0OBwtSs5IcK3eRBMw+d21XmyWhrAYwf0f
0BSvgbod88YBCOvH4ifgAXw1vpU42v7W4KVp2vojD/5JaRXxEZe3KuHHOQ2z+cm8DSVFVcggq3Ws
kKtnRjpSpebAFleUT/Kg2X7hvdmP/h0eiX+f273Tw/AKnj0GbFNLHEd0uPNgWp3YFkqVxhdgmNBh
/RkSLt5I+vbwyg50I7feZO2ol7ef/orAmMk+MBdyXQd3p0Fx4oJvnmYtB8zZDwM3AZgcIDAdsjTn
wXCLRc0NsgJcihFvaIePGnKhKkUihGC/z+bByHFEtT9GUItBkdn47rDehBCdtRXDDzd38MeEEQhR
NA9MhudLem5VAT150/59G5CJNq+2Gl1qrglMdwFPFgcIVSTQIPXy+dN2e05Mq68ByVoc8Zd7jrJF
9GHmIB5dgB8nD0ZXXUHtBjsZUJUo4HW9j8M+Jbh5VCsK4SCJi3fBdnok5hmzzfictG8miCAH9w/v
t1LnL6TbvmUZr3AZW5gLqzanvtnELOvzGMhBk1PhYssw8aEHES0NBzUDDeuwruqoaP6N2idNot4q
CX9GuPe5NwLLUKtkxedqNGDTLE2GoBzkognOoVxv33YAk6eliA0L4NvJT8tgjGnjTAeOCWBD/hts
TMNy6/dQAhDss7/NFdt5RH5hRYMUf7SxNInUfO2okiHm4Jn3lfY2l3OAWMh4tUX068r2tTHbninx
jDmO1sgnpEV4e4tfasZ1p/3zHN9iSHU5HFaZFAA6uRU6YC6bseWnF8BcYl66fA32FNQ4XvCYuicL
K7PhfMSOc8niKG2yEg6P22ctqa4xyKlkyF4w9KKiZowMMojjjDan7R14h+pZhUH/E6DdFcPErbEH
zQfZoTFr9DXtdAks60K8sU3O6r2yOcSTc8TIx3UyiXU25V9DQrj0v2jCyRutOepbyMHSyjQWny2F
kEZIbgHX47orgM1gf7kXkWdbGrVOFRkVlDzYrkatsJnbG/QGpGqKFUW4zYiUSbMgSDetw5JR06IB
ErETN1dVmHOf/Ky3DcgZgMDku946dyU75IZzxUYpM3efEnbu1LMznm8sZlroOjUH+2pNGeOAN9JG
BlOodYxb4W+BaP5ScUnjyz91L2nwxvc3rvKfk9U9PB3eMc1HXvJLVD8b440uXZCdUCfEVNg4YRas
7PjH+jeK6bcgsw13mzLEKDnalV9kDAHoop2VKkR8Zib3YU32E5AGuET38HUJcSQNJ9xp1b2xl4vM
+NyMEddxHTWeiODGBZVFNdWm0ONR7m+qKKP3oUVr2XTixlEi8clcpdHidRN8GrbI31slMRx1TZUd
HynsllGXU7gd2gyQ0wDYC4B4dh+SWnBhsHHkL8mgfbmEVjd9AMfFUmBJQxYD/GeoQQ7D8S7i1ed8
4T50dTIq3CzLjVPI6A7EjgGqF5Z3HuolA+Go8OBOQNIRQo32gexwLYnRXIWVIN9awGimuSLSxtHg
Xf0mVGgQxZCMNU6vzjYhwEQ44Ez26kAlGe7Q2Jy0AyW+shj4leec65A0jNeacL3Kno1//yVnN3jm
vVHJJo5rGwhB5xmeMhJ3hG/ZsbFGkP7MZxc+CmWwpUW+rmu2f0gMm1cXheL+pWj1PVttdTlQPWvs
qN0liz7bjovB0Nx5VCO6Bj/t2yMSIpYxPtmDlyn6yjrQybL2z/QPVzFXIcudB+msBY6AHO0sm4Bi
AXmwyRNm4EOaGQNzD7AxCXNB22LdoHHEmOoLROU0sj7n0ky9UzSlHZqpXJQdA+3Gw/tBGK5OTYuw
pnyT0FDZZ8t8rsJnFrmXp+Dz8aWD4kld09iBAXSDfioqYINi4QhorAiobczpm6LkoGPoW9Fd1i+H
drmgpeIgDnLkKlJUcOevhfNeKf+dwQnzbK5SuLEbZdvUVkThbETrqKXn113/XJKQ4o7fxo5vt2QK
9AL3kUkwPWBd1J2FrHoD2ttVOqZWDOLfAeJ1dWJ4ZoBwM7gp5mboxqV7CpIAJmPnqeAJHxo0Gb/K
W3FOToB/KHSlNtri26ljW4aqTze7iRXdVXycOqfKwM598wpJkG0ohfBPFc7nfur1a6VoFtF+rtDv
2I6KNurRNn+zcDxjwQDomGaeDR90tpOzty2bbD4Np//b5NcDQqpGYGjM5vIqLMNc84EAWTEwDM4S
XPHEQJBjEZ00uaTHQGFhX3k0cwTUoWPZLk3Kt20cK2uMYYB3cwnLUbNcetrb4VhvNKVp/uPc6asT
+ksxFtKRC7yunI+9DspR2Gi1WfcyapS+jA08PgBsmqVwqoSiC9EKPWi+e0rxzBr+m9Rv2kUAJHEO
xfqjrIY6Axd9OOUJaYhETi2AjuU6vXW3Gw9gPyj3BLWEbLUXswjTNzHDPbpqMuiLb+2j2Ja3GeuU
pTkhQXbRkj2iHlHHhkIFA+e4a7DrZ8Kj4M+NSB4wtqGjHITqkDnAfqobHK+833q7rwYOaYNQydvg
iAo0ilHU8H/Rwy4PAShUV86yqSfAAQn7hr5mHGCqg6eUHBQQ4jD23ODUSK+q1kZdkcNeeB0Fzk3+
dlSzXD8W+9u/dsiMmW2WGcxmzrDFp5ZFK5b1pRATxXoSYwhf8Hvw1o0FS9grJt4Jy/ooWCIyUeVw
wtDynvkkuiGn4nq3cDQmJ07fX52A6onX05quEviej6kh9Jrut3MF22v9hhOirNJFEb1JzmBIoAcR
sUmPjj55//Fgpc3YJPj4hdX+C9PcpzOf92qSbVh3Piv34BZnhDPWLqREZWB5pgmwr3W6+lp2plKz
S7Ol0zz69ozKM/ldP3GGuit4M+TT1ZnRjhmT7yPWIUfpQHl5abwbEYCzCicJ0EqifIovOernces/
pUoph10Luwq5Q+bkwAj+uCmzLVQ5HG3+pSsE7xLA5yjtjfJhivmnWq8GPPca08tBlcwDC92ZwCev
WFyVVAR5W+NQEhM/h1P5dl+xjDO7ktUGz5SvLcnDkvuGpYXQ+aUXca5lNeIAZ3vtLNJ4aBGAgrHX
UErfifTJx3rRgTQhLim4vMYLjfGEDrXPfBJmGXKDNG3uuCgdGwGlbTzqRpiNe8uPwru6isZLOZr1
fj+0V/Z4AcoQLSYKDcW5T2aMJcAu7A9FhP9Pqwp8vFJadY5nydqYqvGqd4aE+Xk3DoW2pdNhUw5W
1tbTxSE2Fj4v3hQq++Kc+AKV7Fn41v1VK8ugyg1WtjIQQ9J6IvZLMkmSfPTHZXmcHzkBjyY1eUFf
0Yeeuk22RNfFJ1f7vx/Vlrt75IvDQJ5TujYW/49bVsSqiPinUVSZlUkze7oFlkBW49Th4B5dWZfc
0sOc/vqSkM9ykWvIDcfzX4q/3sN7wXiDarbRapkT9So19leAdnZCB0yD0Ma0zeeqZzta6TXnge4t
ofcnxuOITBLQogrZkutESBo+eqoKSsquzcT+QeF6yMBSEU+E2IA3s1mR+oXNLMlkiDuyyK4CVhIN
Y21hZadueldFXhNEVbQl6mnn/wjzKdPZzpb5yVEO+b0kJ8vm/5PEB8M/ASGM/Qod//BOSKqHAJuc
pL7PtREczoLQ04EEWkV0xpntAbaLTZTRXEHFR0il07j3BvNkbIUhQ8RQ4E5x1EimTcYE6CZI+lFQ
501s4xQlfUHnk2hnHU/XqGdYXE+8WMitANIMjvstW+S4tlGcnQOVpRCfUlnVchQ2fzZNVAvcXAyL
fuE/apP1iHRkfrhFB5aCBdCx5EhStPvyIMNyoU0bSSwsjptIeoQZGGIPYaA6vdrvZ3GohqBPwOG3
+e+NhCmHTiXvVLCav0b5s/CxjzgXx5ZqCc5267Gg7HQIaPwT1m+4uM+1bDOminyIS3hONvUaMO6x
iihGdwSz3NY6VLf1bX1lGcKmDvl+JTtyYCC6tHx03+nRIPCu8Rqw8Zp1goC1Z+uv385P6cEBB6rn
PdruRRTG5FiCEHqh+X9LZ6BYUegSH61w5IWFko9xsenEGkPhPMW6UzOkfW/8MvMeautR1INhmFVw
KlX5FBJUeUvvlnwwTyj1fltNXnS575wWwzYesLK3Rr56s4INPL01+zKPih91Av4UMpF958+njm5s
dTQ6msrn7Bu55qA4Z6VDPe9jp5Y6T9jnv/8OEqhR3hBxfnqtHRTfx4uKhuocRNmQiNtYl0n9NlQa
LtWWA8UylRpp+a5hvSfd0f427KTi11RRmPaI6qU4JafFzMlbgQWkTGOb3KQddZF4p65AtwVH9N7d
Qpa0m5flJOdGpfN6MXKVWM2bv50l8hfHfVe9hp965uTzyYWln1S4crE83aMQ5YOE4VASHL2Wwrj6
rplYvTn9Fd3fmgFgiwaPb0NxQ+3F8JzVPKxN4/mVOEY07qPahXXO830IBY/y/PRPWRz48BTjNlpu
Okj2sbAFFW41D5lYaf62U03CpKIOkU/3WUAGfsx3TxU6dpSwuAhm86Su55ACIafIbw1daDoZ8K3t
WuBro4CkrtxKkadp/TY72uh+KQ1arNjjotWkYKxC3n2c5zA/1EzRaY7DzLNIqOPvjvKoVk85w1/u
cMcQozOernJVseqiMyErL1MivYdad/n+47dt0zIUJ0KpzgBd9+P1UqaMHSEnPCxWQm7EplKvaSpV
rPAjsQF+jfeBQiQouTJFNJVjskb2O50rGdgXoUi1sOh6ruHRd7uJjA3pOBtSjywXzb2IQifDlSIC
xatbOzRMChXCQ3ASQLnvVGLZUcBxsfSv9aFxOyI78Q8tL9OMl6aaew8Dftl0Kv23rgRzCya2xMo4
Gu5tI2oG/IuJ7Xl1RK2olOh8LsWH2KcXiUDrjL1IfWa7bRyawkeQR+RsGEh8f1Ozk1Jk+Ngp9ULo
nk6jizp/+9WBB7nxYbIIgE6acHWScVnDROzwlK8lIcT+ylx2DiWKRn3lidSA4PJWGy8lGjLy7Bpa
OFNSESZOgqQ2ya1lObZQlrUxn8ycKbSVdXTv6IL8CC0VUD3zX4om1hU8LU1Xt0DL4W9McftYa7NY
qOYUpoZAtEtCS8FfHqEtO26eaadD2HAE8HzuSkffAGP4IyDm/DztDpW8N7IlvlFerXboExQ+JU/a
oXkrhXDL0ZMBMx/qqpmkIOqIIvztJT322V1McUnnwCeV/6OzV6+TYTRm7/BuvRmjH+5+8AvbVgTU
TyTeAHDTX6i5mUSou+h7AvUy9zwIXo6xPoLuNeAt/BbsXUiLw2OJSbwFZMswPyYJeS8J2ubeD+6m
HvjFVI9utBzVbCN9ZQp9ZI/b8sGRcSNuzwuxWsm48MWXzzh5GxvIHgGZKmJcW/DzUrG3141H5c9p
jQAw90oL5KxfH8qRUJ4tQVogM5b96UfTCXz/5v5Q+b3nJWk1YV8incF/D6rSXPY8yusu0BKcRwD8
2zCmx4hblPdDiR/CHGT0TqQACvmen6gM77YkWzYs5RynrEFESqS9NjsTer5Btl9qj7fz3fmpshg1
IAasW1DS1fsDqrFJRc2LMrK6NlmeJ8i2o6yyK6WuoDBcgnwwugJg/JZyEyennxGy33ZqYuPyrMhZ
SdKox1l2B8JgsphKxONNPYLzISqyF7CfrxkIVl43n37cy+Fv35TLRmAUy7YXQzhm5Pkk4RONldeL
WixJaA7sYpmazKtuK+18m6XUqngpiwqcasnyQ7+lwkNIdQpwyJsjL/a4U3Zuj69zK2BYRhx55pIW
/7rj5beAJrFQjXXPWuC2S0YDrq1g8txN9B1ZZWldb/TFpS4kOzhmMGxWFRWXwbbEQGgD2vPRIsps
SIN1SSmoqmtrGdGAAUP8VevGdnAZ6Xc4vWpOxZKPSxJRPYoSfYOvkoFYUGvcx0JIOISe46FXGj6e
ZX/JJXtPGtScAjP/1JtK5IthQ1gwr2zeaexDArycyLm+AkBP0u36o3IFP7I+jPrsCXWEG0T9gehE
QDnz68n4m5g446oOBQDk9dkjmmxYlnsD7pmn9vlh3Cj2WH0h3jlaerC9lHJCo0gHNGalL0k6F6GK
2uqyVE9l/HVykrR7Y2UxBIV4cf8E0HcsAq1769K8/NKFE/ZYNPVrwexa/Z3P0vGayEBTl1D5If0s
3GOessA2TsDsvoaWAsEqWugmaS8y3h4OZR31nxD470KtUNdEYMDeeDdtPszEHAzzvAIarSE20+5l
KJpo17EjaSW/SvEaQbkoEL23NQFpkgtIzCqWFI0JdCcBi3wL6xCVGesc/ygeZfP5L7VSq8k5BVCa
tFKiPZwWkxSF7BTq5HCTILXgDT7j9i0pyj90TfU3Gk0tk55yKDvBfSOsFAsZ7AM7oswaTnpFqQGG
7EbLVZor+t4OHQyQxZa2zl30Vz1L5DzyhQc9ZK8Eh4m9CJE1ybgsXSbMwmbPwrxcMqhSnVYX7wiE
dKiJLR5bqqnxGdoGu8YQUVz9nns+a8dMWZvIGHZ1aeFpZoqBZkHxMLeBxyumvLu21rW1T0lUFSrO
aDAVpevBVv9VS2NjkRveF1U/IPKFzI16xWmHXf+RvmLn6BoJcUMRsuKG2bGbhXKWDuyYQEqNqcQo
J2aotaVEV0XxiWsTGzo8R1Tf9nPKk+LMxMLX1QS3AuFOzbplPNtEJGtkPtYLIxDNGyLJ113Jl/n5
f9py+mmuwIR/uZCKuNF8OsUuepTCtbfGWptmaQn3eNB7Du2hKE/QAdvMUan2xbeCay188cmc84+E
5WyjIAU14f55HT5z0WJSI8mmqYZ7ydmZabihzsu+RbiDESRdHaWKlaRgHm6V7NNnEdGXmSqgnup1
+6PLZLxk5nPFhN2dlLNdsCYsQCSzN6XVrJrzme7Yy18VwRBc9GzNQNvj/vcZ3XcpVViDlClLvxex
RvdNFG0JbzPrBhFlO0HkWRHhGjkJ/TmrrBoylxip2MHMw1O/ax/IUKYjeImCSED/POx3vv9T+e5e
+jyT/1ILeJaroZanDvfMjoPIOEX82QpScIfuv3+t4CPiXOP4v3uUrHhoXktUGgVL3T9K4vB0thpF
d2sx6sTEZllIiRrPMsQlfylh6mkfpYTZsi5KflAMWms0cyyFhY5oGWe98VPDZvhvZc6Lsnuv+f0V
aMbOQ1i38JOiRuTsXnDvwVntoYJ3QCsLW3QxqfIPrzha34QIOnJvJ2fnkiXZj88ny2OKTIL/d53Q
FvhTkvRO12bzB7wrmR5Tp+lFVtuZi55uJG6P9MIAo/g2xmsZiCvL20Zjtu+kyoo6XSZ9F37JBY3x
fOcHS/vMPyqf4XPV+EPHsOuhV01o6Jfx2lgXsm6Ub0vZ8tyc/t58AGM7FdBzOJYkAXYnDUirBSPD
LJAhckZFarGIurQFFav3HQiUVFLLUrPkV1sjpYYrlOSo/hNDwN0yrlIBJLrgV6UjJ6nfKp+qYNWV
l2XWDQbIbQ1R/cIpW+YjSH0q0LPsoEHC0uThkU+hknoLXQL8irihMCCOfiTXWQBLNBbwokv9EQxb
cWRpEuj38eyAnvGNyXiQDel3xnHvkaLpZlhZ+mouJVNcq8SSrNb2s7VEWwS2fHzxEpP8Xz464w2t
F277l6XEr6fZbTVdERWOVbV93pUVHA4UldfZABkz2F5zj8PcsLYayGKZSF5uwT4klw4aodC+ebzn
vbbou7E2NuJnxuHjYskxb728aLCyVmDid+Nw8il3Mqn6cwmi+ssvbAJtd/UK5WIMUqRsJu34zc10
HsbBUr/3dNK6KSU1rj6MqP9daGVUcarx80sIjjhqAPH1VdVDA4q4bKm83XTSJM93lYPs51mm8/e+
umjrIYT4AQmOo6csUUBewvkR5oa9Fv527ndkyrIqzk3AcXi1C4qTcSjYqnl3HSDSuOufhD6q/n60
kxBcDlVHLe3tnKJ9z3d3mrCyYfvuruy+VAfJDuRNy6e9mi064vQ8YpVCBPefkpj5aTiWIM1q6J6Y
JMPvmF+q5VLbORN2QTdokpBJzwn7Z8R3hIOYorNdgiUBPFtoDHzisgOgBTHNagfBKt9YpY9Shc+G
z2Dnw13cfZ9RbxQ9gn9Mx4XD6RuXRgnXlmcSQTto0qLqmUcUOw5j2LjsMlhVSoEG1NgtwTtSDBtF
uq260SxUtmchaFe922x9wQ4Oe+AlLj/BY7dgO+ealVBYer43XEF8LcV1P+58fUg1wYe4l0CGRsOB
OrLtbPXC5cl7Y9vjrDiTWFfV5xgTu54jLYDATctQuhlW4cgTqLO/kb4XRSHYZXRfaL61CJX5fN56
/AyPG2dsRDoHcGRL6XLMBTI7sCrwm+SGE7HzkUh8Fd163a3dMpAg5CInIiFSpS/xgBGgk/mloSUZ
d6jxwLkoebjD5juRoZ7dv+Pr2kSHnq9mEhe7W5WF5LzCJclKDux/KoPtuyAPQLYh6ts4SOV8TLCB
IROh12JB0EQUHCfsyZSZ72hRn8UoL2yrFhjPRfbWd2zMBOfqf0Awx8jmz4MHW0mJoeVrLOC4TNHA
knI0ZDvteq8JkRYRJOWRC1uAGT7MSqRU3Z5LeHRD8YWTJRGOyFTAICXmOfQhbZ0giSd9UDfVeQr5
IRTQF2AZoLTd/xHhGtaqAAhSqeCZFpSIZKQBSdczTYEPylquskasOodEv85uibWk0y+2RLyKKGpQ
iNvznuvNAeEPi1W0vV0mRpH8VgwjlM1XqXtoCcY6OYd7bFP7pe4AVQiKiKfOCxK/As1YySrEhetr
FgO+Y1wxEm2AtC6aYxHJt8NiZjuMICxynZsCNc6+sG0dx2SiSqHAZCVKlfqDbNfT5i16OKWu8Dza
Fy5e6H/1/dTapo23Q+J8zLTKAQAK0wy6neeOu4rYqlVAbuLtWay0c2MH22+/j2E7DwZ36njRAqSc
laoAMnuE2FZ/dPI3zLaNcp8Gv3CkLoDJJRrAHKtXYlLoTrQDGeMWAEhGaj38sBwXDqjaxaHpIybd
lrm9ycPZG1Juqz/J9GN9XUmsFCGKameaceeRv+Yn49y3RMqsa4KfkqTIh69hjM0p+Ckvc1ElKexI
5i2Yk5Sin3aXk6O6X3M3FIHhz+7Ad1+wk//hvePH/XvZdt6IH+mmET8zJ98TTD0JR/t4XwaIhjCX
EPFP6VO5FocJ928mo+3r0Df3CdVlSEijAcg7glP6zxG93WzJC46+/bAj8fF17Shra9rUX/OGVtJB
B1cZx2HJZOTfTUzA/P2gCGUA8bRYDoa6OuiUUjyqG9TBgdEIN0R925AcP076WWfI6KPKxhIrqJRL
8lpy48vCGG2Vegvb5HSMKmzJr/xPj712FOZuY/ZDe3nU6e9Zhg8zt8IyhFU91CZlkbeCZSXtnk0G
icpbGPZ0piByxK39xMXC1lRTiGRooSRWkHugG7CuXrnSePgE/fXSUpLy50YhbUMrpEHVgoTvbidr
XWoEfZg89nLSp7egSZg+gw1B4yqAfTnTCilntT3HSZyk59xBZuIXFLxnl+ZsYeYF8KM8+11/3N+2
09srePqOw+Y4GIkDK9mlwVn1S7oAmUghYop04Cxm6HnrAEVExlhdCx0TzYPSAI8ghNb5G5InHdh4
C22sIf+LMPpgmWKv9EEC/sa6imyITq9mTmoAysi707kwu8lU/+IfOqhWl68+rHsvQwncjDVo/Lol
OgKw6ebZvEcLYRjf2ZDFpnUEv82MrG8868Oy35AGd74YVN5BBTGJGM3h3itvf1yQ9rTGafxgdmSg
THrd3CAx4foGKySCUbmHJ1PHqT/bNyB4ZvzJNYgB5my4SS2ffwCldG5GHWltFKRHQJ1n29Vg33GM
hc81X/TWERxOLTysrA4F9cY/sQ6H4JbxXjIFSOneYJjJhfmf0+xpPfE47fBz358gL9/srSgChcQG
W7ibYsFNvItOAUfmz4Ej6aYkyq5Le+1/IAhk/xU/eeKaAYzlFSaP46WufFqeCqRqTzUkRjLMSK2K
fnpE1u5l5242PLwsMqwQCaBZbkvlXRF5UAA/2DF4UZnVCYIIDVSUDzTd8KD0vOOXIlyYjSbuaWKD
K/NasT+gqqcybOTq3V2ygNpTobfbXbhQtjyzP95GBVPvriA/LckLfjzFrjOcIEwFhofhyw+r96x1
ks/d6+mQgbvBZR3FFam8Mz1snpKi/FZOS/N9AwhdOeee8M0TlCr4VBPaNcigMMB5/chnZAD06iTS
OuQonfixuu+46BVpMOHiDmh0kLpw1NJqsGOEmRMBYb5Ffmxk1BrZYxP5OcWpAW//H0Tuf6lyO9s1
UxO/cSTZ3rBViw55sYEHrKJFzPA0nUkPHa/3mkgwUoYEmIqudgOSuAQvXn+8hlnXUyZF5lcXKU/P
mhFNuDXzulPaGOng7R+ml9htIvuEdbYtNyhDkqfZKl/y3fC7OdyrMgPvewu0PGHXRhXSV+zxyb7s
p2+CPcA+WgWW11oK39RyKcD4qQat4otC4YicvMO/T55OSB0/39XOkuR8C4G6TJg6CQ2NBWtP+5eE
hu0tZ9itiPLMxBmCE0zbR0Ue5+ZPKFdfO0RpWbXAH47Jo9NuFSdkvj87gjBxQqQV/EAbzvwBYwrm
zJxI9gVS0yELjQykyRVscXgHjhAs5/xaZkUv6ZX6xWj6XWdpN/mdddz27Ky7iSXeKXCJ//7IhVAF
81Gpf0YlQVcv20YRa+HLmk7IVtiW7D4hAKMVTJUrRSPSNp6irQjMH+JX78ph8RBoTnc3z3zjug9e
PbpQPtAv/FVMoxu2BYjgEw9mt2JIGFvjkli+7phgj0BTvHX+hVzKKeywqW695T4qbNwaqJbo68aB
QtKXoYJyI3RKGMfZEY7/XjMiVJXhLgVObrvBXAy2MHTqraGnrZWPCFQvqhvCc77GNS7rFIlwPT1L
jWlWdRNcse27qc9oJyaZfZtnq36DwaEvNcR7Yz7sgnPb8k1mDIj9Edq5MfVlYgWjJKX/cmsh2PGo
pH46evJh4YjBwYbR/gnutl9i+eL+nTjq3LGpqYeFft5DuBqc99E9CxT3ZwPFe6wKmiK6wEqHOwLl
gXp2pYFLK2Ct4cpwIeEC5DVjpD8xSv2EklcW66qqhf8+pAP8oHQz9kwxTYUtNm5auzxOrs5Fweb8
7LVIPrehl1ITBgW0+zxOkDJAHw60Ghi4ssakn9RBEhocQWLAT/AEzw94WshOALWHyK4QBeOtyD8i
in9RGp2VdMz3KKUom4P0afjpJCqXF5JtsAAhRZ6um7gSrBkV0RY9Hn08cLBED+LNNzz3pv27jJP5
Xq5cm0Wds8eeQ1Mc55ehXfTpuGouQhoEOWId91qydskpzFewNJ8+M2OD5lit3jNnTrDTqBgJfuk+
kiubUzyAXiLmBPZqJVjS01A5KXQcSR+Gf83KeqghK8QzNPPyH/QSzPc9B2w3vobudQuXveEUYVIR
LFrwG3FIDUSwgK0U8BHP/Vb5Dxt3s8bHHfrNsMXegcL0tWJpoJcxNG9EEHFRrtcsYg1y+nki8CyA
3U92pmutpV4YH13uWWxL5GP8LhfhvFJB0TyBCDLsPfZhJ57cYB/FZ+rQCGHYaQqzQeiPahsCINNA
1a+ztiyQl9U3xhEYuEkK2uywHF4Sk9NtlaiUJrORSabwuL7/MZR/kwomcqif3z2l6FLeFwypqHVE
RVkQDwD3Sr0bwO2JF3IxiE9KREbY+iwUEkSiV/HYt8w0NLSfnaLuUwVxu5EXut8RJJ2W5AvfQZgE
pP7VaO8+lwLrWDzpyq7SgV2b57RUx20U2TjjiUWW7xyBMmuQrfclmTemm0pH6m2B2g08wr+LBh2c
kBMZEZ7SMQ7C8iY4v1MHwPcpEi4sCz7Mv5d3R1MRjmJfnCmDGm/RthvX9464JADqm+jzB1Q7d0T4
LkAvmHZw2dAHas9FKiYRn7IW2IFuame19nkvWP06XA75OW5cupVHsMXvPTVzkOVwqBdhUgxStT0L
O2QWfjT5+BbGAY+6j/iN+X7LNDYMpvLVLtgGbOVbcXPYsCvh+EBH2lLaVL2IzFwbLGA0OQ4S9qDT
T/ORUGkpeFYyD+tD+men/GW7y8YUE96DdVPIr7pM5o9tvJzkqsedfLK2iDUG8yCGmIhl8y80TFFH
9/gh+0eZzy9aBebn2KiNI56L7iLJnsZQI72wIe/0Oi8wN0hK1Zkg1K22JCBrGJlp2mAaDl7pDJ1r
N6omuA2a+SoQ+qX1YPZmfooMCDWfzUhY5C1mwFxLYwrKdpmksS/35rXHc5m1tpRTwB2mxggazyjx
DNSIxmbG7hCMOrhUibS7CUvAT+oH5u9kPPh3O9IGKdR9FzPv0SoPY62TUHAu9FxTgGx2qDWvzQCg
LCSKf7FYMewjH/Q9Fx2PoAPL6L4CV9sMyl8xWvsXuCxSssR9u03KBgNAENCoEUlewNlRTclFoeu6
SFqaPWALgKQiKJTq5KW2/E8vvOxu6Xh45Stz6vF6gPsVf7rmXAXDnBWJXXvYD/lDI7XO4TGKaWNu
PCr/jo4PFBfzI16e0WuKe+4/8663/rt9a0fICBe34K0hetbznq4/AQGqs5NOFCgqeiEttalpFJOi
2ZEMsSs+MleF3Wc+vsFKW2UurxRykVoquFxj6ru9ZMHjYI5R2ZWHo7IGkgg3r+2gR2/Jc3wwa3lZ
O8a6TdhXX9XnvxVrQlGyq/vQ4T5k59x9SLhb7Nv1Bb0Ie85VyXbRtV8PsT62UKW1VGi+nveEFWEl
OB84gqhpjYdvOw5r4G1rXLSAHYkQjJV7clo65j2djtORzVb+I2xvMTf+V30ztbcxSC9aq/zB6sfd
igxZVHbBbq5bL45b+WpYUWUJU+XLyRIou7/nFWpP7UeZhdMZMpNdrAUxpR1md5rtk5TR3s4vXEUV
cjHEzvE3vOT5NgEunMtvI+QFk9orq7KqnbA85sFBmrYqgV/zVpaXFiMekD4r90It/eb3RSPZ9bpk
znoc3xVX9srJ7m0cuFSqisFyWJ0LwudxplAzx3522nEF4nY8hmi0IHgWOZjy5OOsglj5ZZaa3J92
aVG4YjiLkrD0wahi9jLH+1FwkvfZc/oHeT6fPvxkjNEqbUGQhgDIbcG83sHY9qf7lpmSNJdqG/Wm
bVeF/bAkuS7a5U2X0B+OttUZmIPdS4VTc3Ze1kGx3RBegQztXLggSG99QLm1wAQ7ZVupghLLqSYk
ywHENOCRo01Bco/cb4iQe+KzWMufLAlxuOEtrJjvwXjfsyWxmp+AJddQlNfrr+SYfoExlBvBtetk
YrlUoSQ2iav5jPtQ3amUZMuVfQBz21vyCTdiJCqjWgBOS6Y58/RztKjxiJ6n/312KcSImnaBzYHS
L5l9uhRWOPgoZf6r8e0Hm5WejZ1rnXTRVe53Ug51Tub+nRlcUlQ11m4vKzShWl4jt04bBoyX4f4R
9X9aKU/+30xnrtkPELD3EFIEemR6x6hn1g+X1gqmZKGhJ07IN2FIC2kriLJvovPT6JTzw+bWbR63
WhM6sAD6ebLRVhoDH1EKbXmFy3ZJUgx4ayoWxrLw88fieXiYFhgr4mxPEMYp2AlaZcKq2BfFWh6D
Fx101a4ZO5MEF9fiZeIrUXow2v7P4Ks6EvEJEicELIsL9OCck0yJq8PQaxf8NrAjQGBRsJVdhv3a
eBPK7UNr9BnRqOfVi6GpnRcnJCHJAwDFVf6Ye+jkIua2y5zSF9tgCPiG9kzz4fOjXn38BbyLHn7k
sbbeK2m5xIlskOzB8vPsTi/eBZuYgh+QSedpEx4q4Cn01wtU7lyEFpl8rqKl4fUDDiJa2cd9o12J
s3PUCmvZHZ05ANQMjQOaVxIW1CW8kd3VQQbEsztRG5VIK2mm3lW3iyIGqD66zTKjIp1AplHjrC8p
s7CFdB3lle+ShCaApOU5PsGX4T/HmZKaa9i6ICvUpwZeVCgFNvTfN1MxWfONh0tbmLnEnD5vyg9D
Q1dgFgL6KnMPCnutr5rMTS/bXfZ0u9G0PxujCqv5o73/VjP6p2MYSyfi6NcOIsbTAEQafhqWzue1
eCLNx5br5Cy/LTw8fDbaF9BUr+3D4Xek2Wfb8XNqoGT9thPFqxaH9x1IehWfVPKoZE3/DRH6Hl7J
RRLELoeXwQO7X1tPEPTZ0pHY0Vczx7OHSuJT/OSQ0rBrSg8/6o4xknpF+9Kz6Ei+nNVNbRiJq7qy
MhdtUDiqZGJkJBtpLenaAokYfyoM+VDXEamtX/fErOr0UrcNnSXa5QCPO63OMKQj1P3XzYYsShGa
qExZ9tTUzaoYPPaa+irgHRwAorZnjVoJuOhGXzHpsFbo2+80jc9V3CeRzSqMbEwKXkNaL8KQNw8f
A+lvV3+3u6AfwAnYFEBq2+3cs2sUUSa9Q0/53wiKCnMRaJsiOjjs3+LiVyZu63IOXdGm6KmljxCd
yVQY50CIrFb5kbD+xvpKB3j3XusNP9+DsYVG3t8G/UyMZJyNTxWiC8e76SZeY3NTMd+hmCe7fX6d
kr/+sC5w7v6glHtGfNGKCDk6xdGti+vZPnpE3VNqjlcyxjGIngoOjQP6coNfEKjHxBnKBiZq5Mm5
3snK0490RiOeJ8CJIjCBCdkiKdfpF9vTlyG4zXnTEyu1zX45N6iN64ksbRoCoEF2ZpVX0nZKj8KE
8bNw6Ne3VJ/8RLVIbX4t1QoGhOEydgjE4GG7H+oSn3uLIUStsD+T599Xgi0HNVoHrpa4ZDHlffll
N0VVA3dL/zPELecpzDpLNvjAnzbx9V3R4Y/jDA2NL7IKbKPOgKtx/DLdGkRlibT6kFpojzvkrTTB
s5drK8cGYZ8fMe7aokFJKKd6soGJCdfl7dXFL4P44VCYvHrJd79Ca4JVW/gj6s+58DUCOJEVfxiC
C+uLPs+EBjR1SwaBL/3pUwR7YfQBeijg/A2c8wHDpLh9QSnNLhi5Q9DYaGKIodrOkKB3mbHkbPu6
3i5MOkWAIHlUvjBst7Ls1z4sqre5qkFJey5gAoHpHoo3AGjlEBKcID4iu8l+NMyKnAB235uRTMP6
2c933REmELG+llqZjDf+4lcaK9LV+e4Qs10096djDv1L3yq8vvM3ilGResid7iRf8lWR/glX+eNP
JmW7mj3e2xOGmDOP8ItwVO3VA/w+1SGucKXlqJ7zqm8DoloyNes1E6dxxzVML5xvknWjlQmOmx7W
+H/QzzOrb2+sptnoh/92Y3XNZnPMFNFyiWO388zD8mqU9NiuvXy3c9WSgtOtkK84NXNScLtHPDH7
I5pJ5+i7B5nNFXS5lweR7mzD4wK32/dMvy7YZqcMK2Pr5ta+qJnuWz3ZaNyaiDYHh0Fe6vR8ATjQ
LsoD8dNI5+lQDaoI08F3CJc9HCrw0Qlvln6S1yz+oVgDoFt/3lbCg5lpkeA5wOGN4EfVt2aL1yRO
00EoXuUy7MBptIBQLcCeCBqw5W/ZZF4rtiDcBihqaz2DaAWzWfSU/L3gbh160Rp8YBpVPOVRgiV9
BRYnFnL6Cq2rUVAYPAyoCha/FDrAUxu2+Vceomk+kJkxFxPUo4+hGTO5Eys1PXasfAkDgb2JCxwn
/rl9HW7xBCHl+3Z66vRYu+qDtHP97v6eMY+Nj7a4A1NHcRxhYbE4ZXYxeaqBHwzMniY4JYNX/Xtj
gge1cnns3Cg/f63L8I+Xi4Q96ZDqkMPJoh6GcuoqPlpMN0+kPlUTxP/4UEpZ4IcBUHD3wn2yDdk0
bXwsqG6VBunR9usPsRQ8hp9a0mwxxN5mZTAZNPW+/Ijvg3IpGMh6JYRcyhkOkLbNOxqMpKhrwqL4
VOzaShDP1WFZ3Z/+VWpmh8eB0PtneoVJAvUgs5iCusM4mBlVyH8G5tbawtVIlT70lYEatlZKJRzV
s2cG6bPVJdHcBbFyhoHM87yW/TN3gaf1vK1M7DTs8QL0zGWyJ7v8rfzZifJi2b/24FBd8l7AeOH2
npaHkG0jJqHzdihkN9fqu/R4Db+324J6cxrkya5+oMKEXMpieUbiTWjMhW+O+Yjgt0KcO3zvLflw
YM3yvR2o2tiQqSbcxJ20s4rHzcdYV3qEssgtriRAAi1JGC8R+y1KHiwnC+U+lFqEf5c25e3pkObF
cFV7SVGk+aW3duwDxrhFM5+T40vIU10WjxYTEuu7Wjaz3P3UUONhGTwBr+PRZS9SnsP/STQAmd/w
sLnFcTt4jTX3r3v/xAhNYJHxVhUzoAQ7fE0ICJbPwqMdfys94+dJHFGv34SxhtbijAhsz/I5297m
QcLpp/R4GKyDIvwRrzLNYBkVop1JjBLA3/pJ4hMg+TPzJk88Mj67Jocch9/icd1yOI4cxGDJdaog
JqyH82wZ8UXvxiXD5FxgY+8oiOj1HqE2OutyDyoPei+1Gok/+ybT3kFRnGPtYgW5AM8ByhHDOj2y
SB43VvtNdmyp58cpGguBijywQAkugLQUHXhfsB6YOCdjHc8z9peICAHNTBwJSni1vXB8FVKvQJR4
zx47oA4g5mjJybdmlOxEfYAA4WL14mGWOmi7lVK9uClbWzAzI9gd2UkR9/2Rx2CZxcGJkagsUusV
X16SXlwkWZSrYQS6+JYA0OYcKsF7PovjKNOSONx+JEI4xxCGi2cHgEd+ypkEsuCJoFYCBLKDODJl
UAuy1LuPDkzDgAZhRD+Z3tSUC8r2TonuDYiPizl11Wuze2IEqFMTY8BE0CHzMPXeI6B0iBdNpXbZ
m5LoG8NsRX0QZtT52UHgO7RzSWgXb74c2HEjMfRPnt4AuMmkfs85+H5S6EpclBkW8FkJejkX1QyT
r505TA5NB3PO/e2nIij3AloN+gSagFltchXHtgiBwSvpK/cpe+IV0TssIrGjbfKpLG/0ca4gVadW
uRyqkUkS6iEL/wmBthG2e8coT8luNQgKaAoL2TMwoa69DIZbqltL2XCbCZI0l42F2NqAk+deWorm
41+8mYsd/7kDiGo/b2mIl71DRFVPsITK5XU28xH+P10NT/KhfuCVeuvJ3psg5DTObETC0AmEqsjv
WcZ8x4iuUEUOa4N1N0kxSAZa/Qng2OVZ5ugHDEqs9qlx7rDN3UIDJg7M5Vr6hVk52YCMX0Ey2NGB
/onvImp1kY8E1+Eavnpg895+WNEOsWM64w3dqE9Do+SfFDrbQLizqxRn1LeRtdh55gxzM0YM2gLC
FuKoLh5FkE2V5rtvizwH/wqc0wnY7MbG8KnC32dr+BqW2Rl/DPF/yqF+w5aQbnM/ByW+9RI3T897
0+NnESajHJ03DIsf9YDjNQb6lOJ+bKPfJqkGd/pSYHKxplw9qof70Ia7/H7QZneTzwL/G+NKpKLo
aIP5vij/7az+YPSB6H2Gego7K1VrbYHx86t3DH742wm1veVO1XIeylKAj1Lu5c/yhfs3Aucfl/Dv
xggjYfdSSGBD+YD+x1KsIx5tZO1u9fbWM54MiS6SXGKcx63aflWPfNX2/wOx6WRtK7uoExnEyFG7
GUVqSMO7HBoKPgSfMOXzNEPKS/9z81Ql6GZ6iyFa7FFEJy6NRRHIYeQg6w7dIH8E++U4H3vmnJo4
1uTGUFwJjK7MH3qgFbdLJfXB6MBffS7HCJvzamwIFKXP7kJvoAIzO9661SG89h1B2OvMRLd6xUXB
trjddvceLN5zhFTa4lALV8tcOKhqWIukgT2vlvogrW6Xm4/g4c5syXZePeWUfHVWTmGWICxBgCN5
k34H0wC0foZ+a2a61vk2pb7f1/nrC9vuC43FfqbkTGnLjDTKGVvo53r+ss1OdXvtLX2nHqbox5np
qq02WqnC4xAi3u04dLSFVOGZt0Q4XNM8T4Jy6ZP+VcXOr0j0iyfxky9xaBdFhd5FTq4+hohIKC07
ZEHsvUfZW8Y/pQrNKDv4HZcNN055iy2K4mCSKdG0VwEtO2hQYxukBO7QZsq9/iMnICR+txNulGCz
OtUw6G3gDMbdQACecYk3NpLNeGmHJySn3kXxSOtIH8IzgSeInZ45c2z3kutlLNNR8VFrKDGcTluk
D5g7933uUP7ptqpxuG6MDgGUEpQ9qhioeA9t52XnET66HSl2KzIMqYh8N/uGKrWnBAO9BRL2EPkW
9lyfSrrpwUNc3tpf27+1d8tVRDNthQic4qSDoNn16mv8S1JuYFCRC4+Uk8Vlokq3AMP6FLkeipln
d0Ulr7KQqSvBEyBezcZdMfLpqrhNGFaozhVS+jhDtoovwp4SH2evs3SkIRMkxjOhrHLkwNIUAuKh
6BYId/2oALgIIiRyuXTLg/ePhLcWg9JXVVBqxvKpF5f+eChhd0Fr0y8CB9p7DIDSapLMAEoMEDQD
XVGpHVM+QBE8+hw4q6s3VGRuFTdF8oTuWa8BNnuEQqMOm52O9ac9A4pnvVN8pUhNxiAzvK2pWqZH
cUUdwhULMch+kWl0KHqil+YlZAg0IKFjoeqQFjnZtRuaWB57Leo5Xr/FwsdEfm3qRYFp47WOy3lA
KMzG2oXKyCta7Uiq8Gbir/rTCF73mKz8c9eEwqD/NWPlK/F7UyBbYpcGJfsoLerAjnTx61geYDYB
kx8mQU4Gm3v9XAEhq1kAqaLgpZ7cm7pQfwYKgVXOodutrHUSezunydmlIYcFd+bSWDfWwYLeQuHL
enzyRWKzMUlIL6S/6+sL0gUnN/pc8EL5HxQ5vBJvDIt5CN+xabHjcj/1trmkWoHgBPFFy+t+ksnz
0fxBGshbyyTosgaccbcy8w4KCi6oTg4NyYaNQSaleYw/w66MMev+CBWiczMueCGNDhGSmpZeif28
oXdDCUhEg9HX3T1Y1gDuiEIUC5B3dHAX082gWHkxVx/3u3JkWUaUayJvIgB7isXw+uXu88kil9ku
+Aci4mwukIKVWnlHiBFmNO306zEnXx78dg/g5/pNL7QnlKN4QfZEeumHsutn5a6BMEcGEc2uc2NM
YgsN+ZaHhNwb+kXMo8cUlls25cWhbd96O+BUzMhRsZp8gI2HZEss4BmlgbihMcEc1qGExlS7/Ujn
ydz7ogLa6iub283r1LH2mLgmROvel6KtwYTGj2qVif1GOqYGHmqp5JfN/KYOm395TQ1S5wnwrADJ
Y8WqBRtCJOB6PAth6ow56j0Qfq5PZWeltC4vQXbRa6XRY01oyTGhk5WDTIiFObwNN2zpGq3+Yf9k
bRX8+H13MOLRLnAhy2dEO9FrDCRE1gxwqgM54jm1AHtGEvffbDucQ1URleDKSl9rp5sP8HxLXOL+
3KFsAoWPeiDszbSaSyC3/QLMzO7be4Dwz9wj/gUvo2Du60+0i5H5IEiyzuHC3WYLEjOO2o6tlCBQ
/uP/bqirWFV9E3sdrd48hDqYw8hkMAU2wtEPU/fSABHR3+Rnq8N+rwKVpKwIGHNujV8YPWgU+7r6
wmtLiqddVg4KDRMWNm1IXpxCAhnbLubywJDOzBjKGAnaQPhm9QnwJwOHYrFpO6fV/vS8amg+R1n+
JM+l1aLQnYgsL9lW6PIgglVhyiNAZHay/vpwVF4bfbfzEw5obgQOWeJbKwTTGGksjJfz6BeBWcfB
VDfZBOKPo1fthywGYyjZjHDnkseRVI25K70YNpA6pkFHDLBlSk+iYflz1YHXB4YAGkW17wt4iwPj
RV03TikOjwVNZsgQtIRz9cV07evSKNyzfH80qHcmzCp9AA8Ujx5AuCyyGMkXflXbyLzXH00nykWz
xX6bdlKrDaE1+oGe2Ur7sw6lTi/dFYkhvV3Jh48AfP3goxT04wVIlB4pohkEJnkJ8CxzO3aHChCj
/q208Og5COc4oQKQ0EAzXLfMnMdZCfGIRbqVyQdttk+MEqrl7ASfgHUttathOhEC1PK0fp9CG66F
2JI+TZhNpybxHrJ4pRTmcHUCjS1yDvwf5dUHJl2/BFEqPWoHQfCg08OxJej3d0FPP0r4NxXUChuN
4RS4Sy5qeFsuP3FOzuv8u6l0BDagFVLJ361Qx/Spfs+QzJop4H4DLFbLuBhbl7ARWgKkIfCoj6uI
QQnjHbqUD7B7dtwdDD9NkrwTJqsE9aCERYRyrwkOZWgt3z8E667Ccah9T7dbum3a9XVdhRsr/O4L
mSST05yaF9HEU/f2es4yGhpUfl+aMKOVZUZv/JIqbybJtPYXTcFo1MAR4h5/vwReLS/PreefeFaP
piufDjqFn5OLr3FdyL8MXxHHmI1AMuBph4Ti2PSrrLJr4Cf2NcBXKOMKsifY7XhPLr9XpmHzVqAy
b5IOC8MTtYCF4TwYfrYEbL4JoLsJQT8avRSD1BlN9k4iZFIrS/8Fy6E5pB18kPv+WowRIV8Fbvh9
XtTXyPgVk8gltehlZNfihGCFRAdQ5LYP65NNWv9877DsakGfhg78z9xVzHLytbAbjRgc36Qe+aJH
B1QWRffhCsyaeVaD8OFO7Tklbn4OaX21xEBCISKG/LSCpZfOHkORAwLq41EYpl5+nNk2wraQvrit
Lm+t7Q04oBTAklZfs7qanRQr2wwj2dnGGPr2YGcOgUT7FgiZt95fd3S54LmVXioO3ERhI3m7Dj7P
T1gENoHEYK2cQ7eMlgTvuoBKBa1CB8g7WJj1O7sVAVZmwsqiNuNsvxLB+Dw75XOhw89i8z9OIUMS
t7RMeL91Sb2n39L8uGJOhEX1XGWj8f7lm3HNWLHF0lfxWWbwB7DM8PP5Vxts0ixb6Gf7P4VdyjW6
I3ymabR5s62t9MnoM6A7hszuR+FXo/5GEhLLXGyQ+ajFtEtyNAo2ATKFuFLKezSBz57kKm50FcsL
QirxghRFK1cfQtlwc9W6F4V7tlVhEzpCqpQRwZgcYxmgSGCoMS1ZLOjiHxESSqO/YxweEx0WoLyV
+6z+DvcM1O5CSeN9kJF3CygS47lZq4xDSEbvxvt0qO+cpKzdxlTa+FEtDPcGYtVyDOqq43gietEA
l2ko7aQHNqzglN7Y7aEfgRRY7pdWt3WuotOYogE+VIqrNYUU21wxUtrBDE7hPqK9OnY3ARiFJEei
FlOhocHbfZ/gTH+GDA1WaIOqoErkdwUeHpigHrWSOipYZGXKYo3CE4W2d9w6tPqSyUNFcL/D74fo
W7oni7IywR7QqGIKj4ZTmMCk2w8TjRSrd2/uJkqPD+ZfrkSm7M4x6IOm68hALSpqjgPEZgFxljwW
Br7ncht68RSIPdtIJLqTM/iq7Sco+EmJd1A80llDku/u/cbb1d7hAFF5A3hWQjc4CH440O9/cSWX
l1JMhZWYI0Ci5jjK79XTt7Tk3fu0QvtCwGAKhviehEs4iw5IkwwfKI7THWqm12aaiE/N2bEn639B
RH9EDdM/k5Uc17Niwe6Z5Smwr/R6AzsnyiJpK02ZGO+SlKY60pOkbIlMIu8zU0SBRWMkdLi+FOaC
5ZlyG3R9wkvDmDi0gTafLw2Ipz3WtfwEt8aNVJiM82UGipENou7oH/l+F1fq+o9CWdR4Gwdck4PA
zRi9IRusF/0kpu1TA70zoeYfVyn/cYE4fDhjO2mmMIHe89QQYIQkIeFO92aTVEBT+DqZB2z/8fgT
x3MCo3BeCvt/4BU8R7bSJam0pAhd2yIkF3i/Gy0IKT7bgqoy8CrJxym6V4MC8yqzHDWpxvO1iyoM
p+dMNJHPhfX2QSAL3ZduyAYMeDPL6lB2hHy5f8o0YqJdPA1ME83SYijq4ib55/5Hm8G+BDdsUmX8
iKMPJNOQhQvRnRVwqJLW33o+ztfjb9Hj0Sb6/DRDqYbCrooXpL2tke9T1akUjhwnK9C7yDbfA2b+
N7u+Yy0gAOq+OzcYM6kKKbr46I6O0nnuWjV8+JdDDVSpAHfucBWSXzHt/vrfMs07XcFFSIfuI/1G
2elXdYiOdt34K2/ZzOjHidUlzLTxc3g+6R6mYVjM4Nv8A1jcu30m08ma6t4CXc+Qe0LPAt3jWFyj
VMUNepyBqc+qPe5W0UZyqSu6IrZRl7DoY+uviYFPbltgXDbtv1AAU5zisYJtx6cWElFrg+nEe3z0
iBxJk8xFB+VM+Au8Z1JGdzhfncZyxD6/AQU0u7tjOYq0WlcXxCYE2uOwoh0hh48DbdJszst3yqj6
3rruVaMH3uyVTmzhcw7PJybz358hJyDsSR08AWpmzxf97elmxqRng9sz/7ov9gVZpCsEp1fMCPlq
RWbV2bs14H6CgZCG8xBE5LH+U5AfUCZK4loBv7NTzVVRyKWoUx4b7byFWdUvnnJ9F5Tq8n7oLNAg
zRpiY/M91iEVszALnc2k6lZEpgShpPdZWwnt55uAmAowqEIALP5QNt3r9JTu1jHsHV4Aax5xBxIc
KsHru6Dr6Wg24vu2PhXANZeLkqbcI6XoPuCrLGcl30FiGLTaZyP8ape65d8sQzFp1LJecWVeSUfX
1VJ0Plm0x7dg4cMfMNgTgiHmF69rTxd/gwt29nXpOEOtH5iX7ucSoBqm9zJoKm2dqRTEsPUY38Uu
RTNrTRRcKM0SMn6/XRGyQp/C20LdHQEuzcPhcm7UUVnJDqUy3T9QwACt8zX7/1XNUBCAWV+gULzq
ScW3KuqcbRkylHG8MbpUj79/rFwI+MUCj1qyFP/2x3+ew5yEw3eXEJjmF4meNmelHlMSYIX8bu10
FmW0JUkdWOaE558ItAmN1Je80ouKBz5ruRzQEZ2gCrg8I95w5VMQ9QjWJGKLR7tpEFH+/ZVB2nor
EMt3uDYVZPJFjPRjqCA0H53/TXM2lA0Zx43F356vHA92pUIKvwLsUHv9nymq1Po792nxXIaa698B
Grmuv+bAQia1X6afYFwKaiwBfqB85rxTTpLKOoX/JVm6ptLSHXset9r0cClKvnJRAcMfPaMBUnCP
QAE0mjcDpIKVthA509JKgp+zM/fsJk3rhybcPS5Otsb3NKAdbdTXtvkXuJGUbTDpP879MfLySDA6
iwdgQwiQLEWtLS21DPNLqflRPNIoMtPVus3zNvu8HgA4gvotVF/6pzN3s2ZO5zI6ND5chgwcXDFl
GbUPIj8edWhpx8Y7AaeXnTe4ImeCoTfUIZMYGhRnJhE3pgx7MNP8YrsKKeu4ulrwD9Bbm2Wpfn9P
/l73/rRwNNglEZ932694KmrdLMKTgsVrwmkd71SP4rj1eF1VgRs3Q6CfdoIE0V2xLHTed1AfgQcm
o0oz6agg+ZDAfSunW6MlXUaX1OeKKxJ2AOGOHXdnRsO+5xUkf0e7qsMCIqZklNunhLmyroPbTXzI
T/TJIJ+JQWO0+X9z9k5Mrz4G1HZE4JNAIDW5ALwNpgJ2qF3wJMF605eAbac7YA/Mh5j1TZCr7u+q
VjkV3OhdJSmg9MD8Ft9O/9OlxnGeEV/dvzDMhnTcSApvMYkkeIec0EDdvBWmh6rO8f8MOmHt/cVC
VmD2fw+FT10lH2K/TF2plTMDrl0S5Y7a+DfNDbExYEhMdplauXDQoZV+BsYimCdk59lABvXTnUFs
jZC36UnEa5b2V9L4kJqMMQ7E7sgHftnoP0XaefAJacjuquJHNkcev+elDkzOD4w8or27aXKgRgXm
/CjyJXSZGeGuRtsUFUJkosB26Y9QsL5FHUD5RnuPWWDtToBOQFc/VZkahNY5TJDe3M1FL8f2FAoO
2xQbcMv+fph2m5pUCeyvdmZ+h3oe9YJnQ38m8XfQAZylRZC5e4NZ8c4XmAUxiZ7h/mhw8G/yXFGK
0lMpVau5h3OmJafn3UoR2dDsfp0UcSlHe7gor19UudUYqZopiVaZTtYW1rJn/7PYYQyglp7eH7uH
npqJWca1L+rCsICGCssHckKOvQYVe0E0v80JUoZet2Z1acuvApFIr5+mbZ7IWORtcSTTyCvqC4ST
QC30JJoXSVDzr2paRTA9/M3Vi7K066SJ0h0K9JzsBcU+GvCUp8kED2ozqXV7r7sBntlCEBL/wpd7
LY98atStsYiXSbr1aReB/Xyid2lO+4EHMAMZcexEOF8V7WZ6PLaapQ2vok/1lpJ5pNLr5sFBoYle
q9jwu2ojYIxlC23YvDFh8PPuuUSV3LDPez9tW5Nwstwtvav3K91pLczpEKSOmIadK+q6A32uz2FD
HYFHxPwosiaPJFiyF6VYlPYWxqZMEWUlAk4HAAjpKOUV32EQ+YJ5zOFwUv0F//tMjOxImYJFm85u
q+KXLMSnICshozQ8DzgLZZ4KERo1S28nLqmW9msqMKQyVHOU3LhC3gxULKaKtQr2CLsg0PUh0YVM
GBmoWyfA29nmooeYTe8zFGkAlq8Di+LJ267vyRVU43BU+vH5W7O8o9tgQa5wm1xcy2tRhU8PTJ0K
rC1ScIFuEW4YaYkvcdyDlRQZUYtRIl3N/x0RVQZCEPxP7qH/Z4C9CdHd23HUq+xAerrRV3/3LBVU
eW9X8y7WM/fdZyjDP8lM5UZD88DTBx1KbPas+pbRSjPt3yeV/2XemGepzjpZrBAwENnY9BQSmw9m
EJHfAuThZl1pjm4iK4k9kWx9QdNiBws00jhqPCp9anYfarVkswekhyjRurPHMTWqplq4SRq8WrNM
HFSXoTbBX3z0Qom8/sy40g2goCJt7pS58JtG1sJPJfdVZAtipg/YQEIFiXsTZ1yCj3SttnYugH4E
JB2+kxx/UqsZpxfC7gboT5+MJ17jvOdpX+x0qVgs3MehocxkDNrikaoSk8GtiXi2tSZ1xu+rt1S8
rK/h+UPlbS1zsV9wJRtH6NOu4WzYPERow/LTD+UaJDL/E9chqANMfbr/ZrB40Mew2RB2mlM1cTXf
pR7OJH+H5Z/fvvSb7gSHZnYCp45xiJfTid8AOZ6lDi3G4gsuUtc+xBRDxHAjsJ8x84zGJOdizSbi
IIQraU1hnIraIvE/5geFAx+p44KPOxiywqkK8gDQ5zaxsMwzag8WgYxL9YWr3szI7p/dLFyOPogI
iJYJu12glt7eWeuKM9tOAB+eWmEdWVJKfQBlEDX7eTydroF9atH97zbYWs7aSuuZSzUabTD3rGVH
R0ipi3d4c7tiiTuPTTkJpOeslFcLIp/Yf/VKu4Jf8UnTahew0sN6sXEBAFpCJ3Y78pUsYTXPPe1j
a1XA3xD/9/2aJQTaitMzGUG+uSydrx/bbG180vNVQgLQYm5OMmF+JUOc+4kenbVygbe8NGmjWEH/
jPHhUS8byMEUJqls4MhVu9bWGa9dbWiEAjNq2Cmg2S7QASpVWV72bZB6qhrCe7Gc4n0QF2eF8wpW
1UoM+xJfVysEzJ6f4ZhKhWsESZPIsSuhg8+BEiO0eEQ+R6LRgzoYPgVOtuONxX/jt/o3X1cz/ehT
7xy92yjBBlkp8B5J0XtUz8MHJOhmgTolxFcHqjpokbxYHQ8zZIZoX99RShLwl4z5fbvjag8S7qTh
EiQ0MwkYzgYvL2cYQKNwZvCwpJZsMNy2TJ12JkH2yMkmTxjBZiEl4rWVEq8bBjPzxsxuoS8OuEto
68pZursa3fuVpPTe9ylb6LlBdQQmaG3EcOhCbnBnI1qjGGHSrg1gmtRG6aLwwG72A877WCS7I0SI
cbBgy40jQ+TAQmBwl10JO5hNVCYCwFlzsGqNHKIHng+DtR7uKp1xIVMNAhQ+O9OLyp/nhfhDVwqV
EfK/vFFjKWfqT+VqyuuYksvIwo0VWAR9Yvtry0zxff8PjC4ik5q07UggiHeEaTItflEULOdp6g4r
rTAamtX4BR4iuuHEDJNHYktSQHdssusvFpAIPZgNSlnn2uo3/7j+qvIxhZ3s/EUEaXT7FumoXm41
DEZrRBhadhUTRmVBzDfeMY2Jq/45WX58HnzGh3ANSe9MboI4iznrEh7SHLnaTVjqcIzTiO3uXogv
OrSZatNEjmfUyj9bJT/RfYdvQl0hAigyKDojQ+0M5o/0dk/05loeoDjIdJRf3k5mc2oluXv5pUqX
EXwbdHaveaVWcJ7DO687aLiyrKwcTIEaHdhwDWMn90LCelI1nC8h4sqjuJw8o9AlzyHeffQiLGQW
Knsc0p1SitJpveVs9LxoCbsjs4ZkVokSN6JEoCPYx5bMh/u7vbMpHMejZVFWnKq/R6J5UB0trntZ
OKXOaL8uDqB/1UTX9b0ihmMZXVvsTvoM7TaTV6vUdnvQhNg0HIAkgif44RX6dwi6IRQAiKz5wmQV
bNOqhx0ZLdH+X7fLYWXvqzwDodK+N4yoYPOVcudH9PjgXOAJGMY/J0wTsdlT4Dw5J9ZriRMJUlpX
at/ecO18m901MkEFEIm/qs5sYBYEu1R+WCqAb9Cbue0nO7n8ZD2jjGlgxTHQpsalbUSChW1cbIP2
bFedzScJH+w//G1oGRrEdBmA/c7MPQMOramt213fWS4ovb9OWyTd4emyf83/X3xHjtUcYoTZzjZv
mqtqEtG0VpKKnBKG1kVEwAEwfq29QNg1EO00FFIXiq4j/w8tkRIelxVQvOGhX/nP2whcK2Hi5XO9
mnsEQBVUnDVyNh/MBGkDOy4nJB3gmvDUFsQiET6wxibe3LyesyeyePDj3Ea/LRNmsvZVFYVFQDsY
zyFfvaKZfHT0pPS7OTyAyfIIBvgsz5mGc+DILamPXhzG2a+NZegEZMCXaDjAHcPjvUUiRuUVW+kT
fYwDPJKc7D5kLecfnmQ9PpFsSxFBd0mJ8xtHKia4TAkZp3Qw9fKa5SyEv3o33aO1oCxcGs90VzVZ
kGQ4x9sB9NcRmxoSS4Pq6FJ1GQ1XgeMjyR0+TcY6kYxZzHfVBBm60tEDBF3C8xYpqkGWyp+I3FoW
qKSRXD2rwZTeydAhw8tDuR7evCQfoRaho8iDO42FKvF/8LtmOnJc/2LGKRy53lWXEu44I2PTmf51
C///+4GZekgbT3hiQAmPHW60ZKk5FuRtzSK4gnTxV6m8xJbJGzAl7WRMrRjiPPapLbE6BotavpiN
qfe5XF5K1d7T6nusjX6WyIobctMli8PedbpUHFbtzCKrWM10c80eeyKFkUH/OFYcHC6eLvKv3w8N
wUso7yBiH+nsrZUYjLI31JyLuOXusli3lstCw3S0M355woF03TspoqBRO/Mxm85AVQz1GTv109t3
UgI+KVQ0JprPyuoN1eznAR3B6yQETH2UwuhW4iMus/baNe3c/SJQDorceGGzGWu3FYHiqqn6aauA
0+Hrmf+HrLAeS493r4Sl5rPnwLfPuGm+PLKUwjniyCBP5HXMYsl7OP6GMmubiMeVejdLFzlrfN4s
mkjl4pBRZeANdUJBXI2ysR6RWfrBH40CAV17N6rO8pSz7h7ql3rqJ7LSaWfmAJeAWfJ0l5/LWwE1
O4FxFZ1uM8VPcpdBRXXQw0OOlxQVHNWLAnnzWvkB0ww5zSky2q0mOykJVGMuqs5/N79noxvQ3GvJ
ZM4GLNONQXd+ZEK3DNQgxALyJ3NKg4TubWGrpP5wPaebJU018iCYPgX/nrT0PhAgJAbAQUBQmpY3
c/Uxd6zhHyjUJjsQTrgo8mS/1mpx9m2N3Yt+J76G7lrLZCkK++v5zBLJdj5Y1MrbGYe4SQXRfedw
4iWnXLAj1M7X9SaNaVZbi5Tsws8uA9x9YQ6U2crj9I0ACK+80veHx0KyqlY8bP+AIkmuItsmOw3d
fb6EOxoF89DR/PPsg09mAzKFFbCm5OeQKjfeeL5vV5I7S2KyBWE5XQQqlTBC3H/+8k0FqUhAdOBU
rqHoulWOCR6wefXivbEUA9b0+YJeh2CBpB2jb7s7eOInUQoABD/UqhedjBalLyWSSNyrAE/074+q
bKLOb9pwU8y+8QYw2yiGybUgyfUSrJb6nGMHsPcCvsohuOby2C+50aVV31Z5tLmXHqs1KsInicA+
HW2C1nNDZrOuM9jK6HfHMhiIq7fKbqFZLv4uPhclTsNo8Lv03yvW0tJNR/wscrLvTjlH9vdFkLJM
XJsKM9uyGn9s+N5vuVJi0YXJpmMTrsUnfnuKV2x4Jqn0G4yPxgBLbPzrx87HyEATdr2cDezPLo/1
NmDwk62pHMfb140DbXgLvump5RKcLf+GOBfU3e9cp1iMyJ6EBwQ4SJMVQuxA+K4AF2D3fYCZPkLO
N6Zn2kMjWovdEHBzmhY3tHVyEEiFQIrI58Fk7QT5wm4+4sKaI4FE5PcVJ6JNu7tkKMPz62zaljOw
9SgiRdNuL4JYXyMUFDnbnHt1lYUdp7HLXLKpFjVK9HGfjetjzmW6QfD3PSN5Y8KdIOJGhkO/MmWx
/hTqSfOUIv/KDFEBQ53btAezZ7+bv0j1TempUxxfTac3C4AGt8ws0oEsizobWG6zTko5seYOJ5Bj
JDTyNXH7g8UZwwJ/jkPZpaGxWmoAJiFLCTa9MQcgOF8ylz/zKxM7tthS6aPYoxLeM5FpNsgNPfoI
8fg8Bnd0qU8RNilNFoG9GYKHqWntnqFPPqyZnfHiZFlKMcJ5bAF+nWNjX6jMdMjCn4lzORCf04Vg
Oh5kXUqPiNygVpSv/tnDRfhuhn1RUrbe7EiGrYZD4O48ZfgGh8okMjj6ZBbYGny1Shw9/Fkyp7Z5
qF3lB+ap2sm3d6613Qbms0m4s6Wv1O6RdzpLrJJrP+sQl8GSCya4S+NzYA03Y5l5dniDdyB3Smus
GNZNDmgTZwVrjJoFiuUz7qFtPBqA2sccW4RCuh/PUsNdWiVxrL/NYZojIMRouDsitTT+X7dATrb2
AdbnnLjQzlbNY+nRrQO03xXobH5IXFhOKxvMBipGF2GS8sXxJJ+2n9Ecp8YOx7p20IVfs9vKd3LB
mhAeDS4rVdZ7ymDuBUIk81KIzl9IqH2dN/QlqQXHUXlLj+XlAQrOnhY1a/bTnPdj9Pg40Bf6fuWF
/GufWE6ukIlykb4bPpMjZl1e0M7ECDRD59dpqW2iPoS1KAnw9c3TCb6VeoEo8tDtLBPowoOjxtsr
ZB/XuYsQHxk9PJy26HHSGIrilsd8+gTLhINFRcNelRP3MKqAnsbAWSgHjdnHnzN7XA2QFKv3et/x
2x4rBf808sef0Y3uBML7zekWcWCuoa5wA4iOYT70mlhP7TVjmcLzsggC+GgRFcML7DZTuhCatdhC
+GIXVpsK0a/lDEhJI5CjU9z+t8rqUbGHgGaMJpp9hT9Fdq9bvwXF18u51W0yPP13rJVKjzfXZjlS
NceEdQjfgXa+Iqze4CigjsOE/vXqRZSU6jXOho4Vv2/UoUwhlnY7MluCM7UVLvG+lSCQ6cZoA6Ee
CujwG2jQPVJkDbrOBZFyh7ol8JPLSg00+d6ur1oH5cIdlZ6R6GWSkam7NyfoaEks6VJVdTLEMK2t
joRWI9qN1Sg2MdrilCTH8gaFHP4pnhWgd5at9V0GoV7iI3iGNa61AP1CJUOUU2NlRa6lZGzogLjt
6oYYanP/+3hdVqfpT6hHBwt1Be7Z6Rk0dVQo9jPmZQnDgRd+b3sYSNZmtI8tTExlGiR3WiPT9m2p
/v6SagKeH9XbBk/eXJPCOohjT/M8MXqOe8Xc/Z7xb3Nr218hWyGXQtrq8cTBNZ5sVyRQ8m8H8dgp
SrHV/NGcraIAuzPulqkUA1j8D4NqwueP2pheTid8WftRasuBJZoZgj6WXyTq7TrcB4p8OAHykTP6
5Pe+8PDFpozcVO2i02x8BgbjS8KSOLs/pf8F8HNLJ9vkBiiKqI6PoeFJ8VqTSwwIl5ivVCazAvpH
1r8BVpZ5uUFA5WgB+kI8uOD3fHH8re7F0qY9cGEqaRF/B6QuvH+CH4MVVxTIQ/2beg0Wdi2Nxf/P
XvA4FRpx8UsxjGk5bnHeXG5IsWISrY9iIJle2xK4XFLWPVC3NtPthnkgOCO+rccZSb/XVALRen6i
aZqwiqLsSOpdX8AlAItg6yUOWF0k2NzhD1MZ91Ogsud2LY6qlGoDr11kS6trLF5cZF9RMphtoPSU
2SnCYsjEYBq9AvawiXMMPx+GpYvr6WOPhVR+UE0/1Gd+AlYidb7DQiA7yQbtbsU4Aqf3ttzvLfit
M4dLUy/8BNJJETHEOBC9Criqb9lCNogrDUCOrwPcJeJZE8qkoxoU5tX4d5t2VqMtRo6WfRHROiR6
fvW666O5z2Ao8bZ54x9UZdb5eJXt3wTNfc9Ru/X/3fQ0kOt8pz2NB9X6gclx0MrDWUyWEzvw+u+M
BTkttfNeU2tptJWGcTEKwnZDEMtJAaBAAkoXbINX7caN5vAOi7zojevEwwyHQau2S7aH6vvuXjju
RiTSFZAwvwARPNSaE1WuNB+XMM28kuJE3ALYKgxeoaIdluz0aS9kv3hsBndD8IF/mljRyS8iE8Ts
sP1QePfdVRGsi/qO+bZ2gl4nMaMbuPKdAlcVuG3mE3LUzCOzQ9UY0FVY8bGSJcipxXYuFEq/4s6q
kn/JLl7obvFV73q1RCQDZ7kL+E6M25WgJ7OT1TTrlHekOcZtBBqot0EZ1oIyPFm01tFuHQk8gBC7
7UD+y+R+vI1+ogwOHVOPdOVQ41DXLGR3njd2UkWGaRvdi3Ou+iU1adeLRutAE1l6gjiXv1QVY25K
VztpUHOFdBT4obAo3VX9yS8Bi60tEgeZB9rUTWkoU5Ix9661nCm4YEN0ooRaN1v+NLiKAbRVaw0k
N0IOOtxtZ66nsA4Brl+7sKArBk7rLRLciGrLbPBtdxvkZTpVO+r1op+mY01QL+v6ABL6V5UbLI55
XblrIXnd50T5zGKq9s/rHDmfH1bpCBfNL2fNz0S1K4puzRGTlg45hOaVPXYGhBgQB1zKvEkICoNM
IkxZnIKTyrADYD0JuqwDA9pbsjURO1EKRTPm9nusFKCysb0k5iajKKBT04Ftk/ujSXXd1z7vK9Dh
uJog3IbUy4MoFfnWrfv8i64YYyc9pMfhodC25ZEzXS9zH8xeZUfK5a0BxnE9knWMMBX0Q/Pa1WOk
l6IsjUw6jCxPgrLfP6xhtdj2UjPAcjYD4eecFS75or5OXzCHhTdK9J3K7BB0LZ8t9T6kPbLc/scd
QFS0COtkfU1nOSigjtchLIiECcyE66nKvPUyNXQd3l9XjSe+SMbXwBBNwgFooYYjiJLaJ+NBaYSV
s5us18SIjCGcUPVn7NeyR4zClcSsCkzldkWlHn5LmTaScJNnY7HSAFsDpLUGB1rvKhmxhbbaFbzd
WiQ3y6ScrjPqAE3i6PxzQX407/khynKv87UsF/d2ovrZ461IBl3F650FOhvLoHlzR4hXlZNwecs6
KCTEqQ7ExTheqpRlEtHxkc+HeLZ+uxmNVzRB18ZlhLk4qQc4OxP2LA1SltblrsiHqMFpVEU0txCX
uyW5BQA550uwAa3+kIIr9z1/pC3Frtu/edLTw4hTTiy892e2b8jQOqi5/mmqgSYxp0EASgZ0UzYn
EaWWq4dFPnu2c/xGmjJ7Py5Ku4r9EbDbBDzgqneiRXIWWZjOCKLBAOonakkYup21YdOE0DRdtB63
9MxKsdZvdWscxVGBWnSzRp3/VuXs+XVEp17tyrC38suV6wbcDwqqoF7R5TPYxpPyDjTsEyTZvebD
gsUCMgnzU3dJ8Bx+ltdVNowFinSIOJrehG+V95YC+apQKuBobv8ngUeKR6awPVQFdVHmVU7m4TZK
ZysdvGXeR5a/rSIBh6SItCVD7E65k1j3Ja3nr+VyIjmiRxlxa4Y9LgwnUk/v3DF0bPA1NmHrRoze
Z2LcrkKSXTaxjfJz+sNCQ930QRpgLuKcZkcb/2s/V43/5G+XviRu7Y7Q/L4hC2jrMowOXuj5lYq/
caeZ5/99KS+xfwuV2PxjaJJcnzXfsXsAgi5dnfI+PXb8rFx1s3lOkk5WCfwRA1DwTuRipBu+cGLr
DTSK584O4NbVokKVEe/S7Rtb8bZH08LO0FlBAKqHbufzmW0XBIx6QdPDjfHU12tbu2SYf8gXfzJA
rmnuG0Lg+4ib6A48TOQT/YmhYgwu6QVdSB1QIroUxXeVSH5C0+RTLlaMA0ow/oDN/Up+ILYPncnL
lWNFualefWl15fIziJhR/XTjFG0cKlC545y+U8U9jtoHqFJKvf6AbuWLofjxH67V9bvgg6WS5gIW
YR9QMNskoy+gsJtKLN1N9NwYOk1A1mrCdCOzG9oIHUBFL01/KKsv8EgWZNzCTvgqzkQcQ6a0QZGL
H8B3AobgoTfaM663iCg7bALxLs7tJRz30pTncbk40s0he7ZnpU/wuhTvPuXyTXHjH4q6WICamMC1
HYs76Fsth5rcxQ7WcPz8vJZsRnlwZiI+N9URxipivk/qe/62CBTL7tvLdS/3RBTq1VXOvg1Ci1Dg
N0BD3OX/fBd0owOkcVYPhsLHqAVW9iKk7DSIRIlYRCQVpE4jzwnL37/P2wjuMPIpjke9omKJVEpw
4iO7vzhyEJ3bdDDiwLhbO/EwfjS0ZmPHlvkEgqeeDTddshlJ1KPx5Qp4Y2v5XfBcRqZf9wrQJ5VZ
Idy2rQGctc/9w68pbeQgZD7I/RxMGgDnPLP1mK/+Ptp6yujESQSYL7WvvB9h3AyJ3BI4OB4qdd0J
FHnlz1HypnmflQ78A+LwMSHVUPAJY0tK3PAHjDxwldT7F9EqAgIgeS1dtjJhSnXuoyxD6eMTcMCE
Cd/qB1jZgHjyI/UNzOj/tFcl42EW8Zt21h08kOtkvZ3RyKy52UI60t92MYHl2q3MMQ9IbXE+08XO
SUugy53+da/60FqqdtJ6jcahJzEvY7K4m7wl3//hXgkXKl1wkKOFYa1uLz8lZ0dvWXmn0iJstXJ+
PEYbvwhFxlktUz3DdRR36H1uy9Pv8royt/qbxHe94Fh5YeJrJPMojBTX31uM2FW52M6KLWOFPKwV
cCnnuQuTeuHmSyM9Bau0RzUal5FMIe19t21ZGNq+GfymRIBGuq1x2bEDU0IMVN6fujyZXOhx6qJ4
ESEr/UraPIV9h7OdpcJAw0Rweqlg6X1teF7c9wAEyOuirMWL0+xpQyZ5IxmO3Pylxe48AlWXGY/X
53T19SYUlaqyQGjzPeXN9Wjz70wHFWxl4W0navtrYN+W4CD7r8Ky1ocds+fOxqGm/+2YJ4O0cyYU
pC8t1UoZxAb8kpjElZupXFMF1mcwfXGZwBXOvovQ8mS/e6fs+t5/PWLMsayCqWpuY8ZQzfVAaGCH
AoSgP8Nx0LlECKrEAc1NRETcBS/nBZ/cbO5Y3fP0MqW2D1naMxKs2PzqJoIEpeRHMtaV/sowumAO
NrSIJUaL3hOcP+qcj/B8kdIVy0T9iGeBsb8jBze4iSHsITK8Esvc8xmL2yccn5xRdbfJbooF0S6K
rrFGL+qgVRjeyavBo+VHbazqtg29Y7UtOnHen9R+Fa+BynVewBEyGOevJOocOo8z+KUJSRfs40Au
rIqcltkKjr69u33/jB1Kg0iBcY4BZkOMFFT53rvl+Ju9ZDhGdEZkHtLibHeV8wdX8cTLyTG+tsdi
YjgSr9QhqWgsk0VKQrM+/d9zmgBeWYIQmhqDxijcfGJ0joQONq3rNqP7TW17zsT9DdE3pms8psG3
NyzRcw7BoQkWB0fuddHMRXOL3FaunAQUaCWBBhDxTDLt9xc0VAy0jDXYI8s/MHutD+fHbYm+wnsF
AI76ml6fm9icDD9uXyFu6DAS1TlY1xvd6SS8E3BJ8eJt+pTHyD/+aHugg8p2L+ovKAT+yhprXYAX
vQQDGDnzdVzl3gNLQQN91KDMbPE0ty+dDfVC2k7gnmkhWgnL8Ag6W0Pu9xHPv5RgoluzBOCNjY9b
1BMrcWbkQsPy1cB3MRARCbchGpql+iZGcD4l+6bsaphJJ/sS7xD2jsGnF0kt1sbWDaJnJ0caArEp
x0FfYMJWWBG3ZStAvkK3VXIIEogCWQzMjBUgEBnMSTYFTIvsqcjOV1JgDLszVbrUVsLKUQlp+X6x
K+hB8rKRX0Qo3pwNxC4hFxrSvDzVkkZaAYbAiyHCuukx0ODsdUM5ymPbLbxArPFElXTMFZtw+0NE
V9JWEB/qCLelfAwwq6uod4/Si68FX5xRuIfsIomUHh+OM4PAEx+cQyaJ3K0LSc2pFthvm2Ezmw8e
XPqf/+FRUebPZ2v4FiYT9ocxi5YLfhhDrIYLF6ml6FSU3kbzesr/8KSDBirDPnp49PxnsOUNLswo
95OuJahO/dPnrgQrhps3LmEmcJOk8YxK51/kFgl5/WoTPLspSXcasbJdwjGCA9kJKHqCxVhNRAcZ
ltwhcmwMJFHkFYBhQ1jQQioxt97FBnqlhN00mOyZoQcyu+I7U69ikqAZA0jBRvS671spMwqZucX9
MyYk/eOXUb5BKhTApbDjyKU2eC5Y+wmwRq/hS5Hc3qms8c+SvGFKKG1HcL3jeM94PUbfe6pdfSD9
MWkNq7EH2B0Bea8e+Hgdw/nMmNO9/bRPfSpBs3vA+++T/GjqqkOHqqTV4Ln8jkD6aGd7qvmBcPqd
BuEUUv4Knqbq6peRZfsACX2z7Yk5GL61Rv/QHF0QMYPnuKjChFtbCkjSfe78BAslbtkdYHy3+oW1
nftXX+OPHFTXY9Hv6hmTn1JTHrsGpNjd5yiQTu6Vz9DPBrFWohqfsIFuv64NJ4iI+nRmxt14JbAT
Nd7v8w0qFgBZ2Re8BlwVNK7lHJoEot9GFm4bCzQENvGFHEQ2f13fmoeRx4AIsR5IpTSViIm5lWW1
sS8E9p9Z0+sB925R1OE4JQnCRUzH1Qo5OgSCSnMSLlRY7AXdnfGLAiJnkj/cvArZVb864s0hdy1V
iVVdgu+WVP7lwW/Zyi2c/1r7OCAHqudAwN2hgN5K8jqd1qIKOBfp9LcXGycSyLZThUV5Qs1YOvuT
ug9559g/VGPLB2bx1Cjz+N2ns0bupW7KRpas4A+h5p4EdwfFkQG/k6jGxO8Nc35uhikieyMZNH24
paYpE5GDQVLMSXjmo7Z7Roq3vXbrH419Hg/24rKFZpGfzdfKhIcLWpEgW5EeKzUHMt5fWdV2nP11
TI6eqmwMj4pY+bKMShuHcTEDn1xn+ix9ITRefsrkFf3ASCwTa95gVKywJqa8z0FM/Ox1WHJB7pwv
HZlxzVcIIbYYG15/AVXbDQ4UZXw+CX1R9NdOz8waksYr9HUsIykWi9Xp4qVk+gExHiDOB75Gcldo
F1F6reBoI4zlNYBB5OQLhD3Sq7e0bvCfNAXptKcqrAL91rQRcdZ3hsObb3pJBtM51Q7Q4Y1LDsqv
d0wOD6OVlOaNbudjSiY5iDWxqvPblLZ+DCebVwetp3wAHpxfx6n+vujAeIfA8Zzx1iZmN8ewMpuN
IjIozHgfnE0JU/Tn+0EMQo4r4t/ynm6tLzkg7Gkhx9e1qiMbzQXBwjL6+jQD/7x1oC/5+2IanFNi
nB0n6nZFGFZCOvONNwZEuz4ZVe9SmKa8mM1ASsUmV6pFmXMQ08tIgIH8GiKWciiKoFSWRxvs7PRe
uNaGxhpMsO8dxHe8QGApsfBk9g/LsAKDU9rBm+68XdcxE+VHyGfLnFR+P3lfGhb7S9m+L4Jf4iQ7
+5bNYW46A4GK3e5dlb8Bfk5V+IK5NFcRwyj+ALr/v4vOjVuzUv3+/bslvizouPFmlsWLqP5dM652
8vl6LBEFmoBUol6eBBAv0gDiKdB1u0G5x/FO0Xvxy2ShsCxTXDr48bgyp1HX6/+2TFcoDsxVudYw
hY8LYMuLIy8n8iyQY0xNWxw3kGdjx7d0W2dUSdCPE8odyNwAvq8eLGlXZdcdxxJs6BFux254/v4b
ZNfniAAEraro0KbEEfOb7pKgepnEdFYpG78wwFw/n8TPBt4YXPpc2fUni5EBJK3V7ZB+JYAD9t1l
DSoAUMauX1XA3GMTCNykcejPNDs3VzhjENDaAp+wPvZXUIE8BMkUS+tpQyi3PeD5HAMdOgUZ7DrM
Do8zqo8UJD4dT6CZcihkveLAM0XqFEWFpcactzFAA0mJzuKnhi1ljISshnLVAgYwmbicvS0kUSyO
G4iJc4awUvF2iyIezY3rvrnKv9G2T6ZstjLB8IR31sdfcKyc8xzaIxPHvRzvkA2MUBjuakTGySOd
Y5zqNTOQUNpk0vu1FIF+ZF2E/wI0QTmf0RtYSe/LGAX90O7ub3iRutRQQqtGiZOo+MmYYxKfwBFy
WVPnAAUGZsqG5HU0yB5hNh4keg40PlNKs37GMB3NjE6rXFrpxoANEmHtYQG67Z6r3TeVhuSnNrZi
ZvWABewAg0oUKMj8hpYuwUeoOq5KMWoq7nlULprcntXL4oeJzj8j0T3YNVOBqohMSabrNxLv67Lx
l8+tWW3gdja6w7ruuEVQhSBomhdAtxhIHJeTyBlZherL7iyhfjFQ2m9VMtUtCnmncX0f/v6fgrND
uQIX1HYSVPE3Y/hRDFr/QZsysVXUBc6L2jeYFUa4w+Kh28vdSRVerXsQYEG/+K9xtNNgExkkSnQf
41PEtWcGZiXPiyYPiaujkDwEKu+kbN/JaVjRp4Uf9Bnb+rMroRHjafkbUZhNC5Yz1C3FfARpSjty
MY4PkJO/QWJ3U1nxumpiLrYZVm0/IH6+JT9gIdxBxXUdBJVy1uAkWgl9UjE1NhmymUGZsxP/WTnm
2wrsQObBlGfpDoxtOcputAdc1y5/RMDg6WLfoOGH/SIu5hQ6hLqdnCzLE0VAicpQ5cdLsUbG/UHB
CXJQ31R064rtMpQ8y2ONzfUzhAQxs0RfPLw4ahm7ey3U/goDtC22gcyRFz7G8GMJMOy+APYqx8C2
1A4smOZ8jRW2h/34FvAxNCg6LG7VT8MREGqNPq7vORIRJThkjeaLUmgjXkfljm5D4EsrqrE9BYfi
ZPALmVGBhhtkHfWA0CGkTa82g1wAvGsE25YeIAH9WnFjR4xJ1lQWQmDvQzB2femGkGfRtrQhmdNA
ik5QQZmGTvkx8mdoB67wW8prAyO+VtL7MLy1uxWnw5tGDqFAJbJR7Lqlj7VqdpJtn1JuFAZEHgjM
C6DdaCrzFVQpNPuJkyKj3kBsqGP7pfgrqy+nhYadkpgBApE/Z8xgwgYKc8pqVsSadHuDAFVCXGwn
35jn/OtxdrnwQ3J5W3gSP3qQtrFyVOsqyHBNGANW34aENgipRjsdm0V60pfPZvV1QODYaagu8IEr
hAF4XKm9bQKQLrlzRMT59QWTZx4yL7O3W9fn/wQkreohfplY++3cyy0lG+xpSp4lCsXWT4PkqZ3i
m7TsVA39DAio/PCjM+WUbcv1jgPmKGuEP+R0dJYSvg/4b64KaCWz+dIamTlGzlBGF5ZRJITbU5pu
2SHc+B08CtimBBqkQyCcA96qKBsvoSwEMFG1cMqp0Pa02FwNTC0hueiR/Wgk9T8IxTdSO/O9MqPN
NjuZehaKhcU534DX63/wWgMtbMBvib+v3U8cf4r7VplexNWx1BFsiXAsxUVA3W3s3AYV1XXzK9yr
ztKAmxhOsOZkp7KIaHGyyJ1AoSMoe/fAvZ1ROKz1jbcqspXpa1KjOWbgbhHhxPm2NN4zaevCw0zz
U6QTY1lxfmGgdbvjIVlHkt8uIojTRxYZIOYp7O1aH8rkUpNg7f/rwVhNi/fk6X5JJKrfPSdTiyyX
8udCIVRo/B1VdbhvJEgVFzivuayfoAswFC96s8tF5q8/T3dN3emAAkm5I85UIM8e3gJdHq0+3VRf
VUXTLDJA4Lxh92s5cZu4LLFbZklC9mIaYq8hY7rIE613GzQ1lXEEyy7aClEBm+zZ/pERkQCtSDP3
5uVmhnC9AcO146kb+mPyXpjt1rNFNuhL3xoScN5bJbwxS5OUZt/kHpRr4VvXnuAwCypbZRa689pn
i+jn3Hu00nYUKwymc/GjaWaQoBEetlKTH3NBZPVU8WVAYHEKQ1406nkm/2sOgmm567KGTsL2X09d
Ub7w5gHs6qqjfJLKjeK2mLWXuQGtkWOclrOnz9nlV1u/jU3BIFt7KaUniBdYOLs73Wp27enHo3DM
YTh0Idf0CZeAqfGBFGWrgrTguEWHBUsC1imtNcOJLLj8p7xkuuispnB1ewZ8HOAKBsazWM0FDBPn
Zj9wR6Hcut3cR+bBBjbk1otPxmgG3+FDNI0xb/sa3SO+D0sBMbzQUIsvOjTzSrZKRwgFPfjLoUzt
MSaUz/7PPvPS6Apg/p2VZV9kLl8eVYvZ4FaA4je58gXcYqqP3Xiik0vlLG2cPh/qYuqGUTiwBhRU
PniHFbmQS4MRn1w6MC3U4IRXsCQ2KWSkB5OMDShUS2uGo/AkV62ins4TxI8QE31wAtGZ0mot+Fnh
Xg9ZICSDAnoAyfP6fQj/EZc2gvIGIJBPjWSAGWe/d3onU9zwcvbOT903AtmlWE97Y2F3k1ciTZmp
OJH5w4msQ/gH+1r/FWUz6rU9FqKadyOlF45odj7ZUxXo6TLJsnIoclll1KsWgnqfyVE6mVLT/HZd
9wjR1e5eYLvMf1bFPVpqYEY3fgGVFnv7Yj66V7BPrea6b0bct7zqke5D8bFK3TwCuhcVMo/GDl2/
UXNVCOkHIa3Y36rk+wXyIkxXVVr6DQoZTCfOsZf1GBswypLSOxB8BHDV1Stnv4Yz+uOlUH8oW5pa
CL2+6V71v9ZMjjY1bv1dNJDj1/XSx93WQBBprHa3ohlhrPZp2b9rgLyW8WKG67qOYqaxaGvrBkSP
O/YTxOPZZeyYaze92SrMjLvpTu+G87kn21/T4EiMYbmbV4jZL7VDStEO1IPF7TTviKPdRBIleE5/
fP/01lKi6C1gvLHnaRvNPvv5LmFhJ3RW+ZdIzRA1hwY6StSgOpVYr8Qv9dpGE/sVt94oVUdslgN4
GjbVcrE87y2wPHNe9xF5tEU3YnfZXKwuFzkuCsFFZCu1lh2WRdcOrMV4ns/827n+04hbRtrWD2sK
JD7scG5m1c4cNx4E688jaVwKbUdN2Y+MVXTBRITFtMlc4U/SgX46wPVXs81TI6b17oSrudQDR9LH
Lst/y0U4hDCwt0GFFuOVsPtozkz1JxyR3gCRTNgxcpll9/OLfeUnOyaMDeRl80MvrrXMQSx1PbQl
cZulLCe9BP/Uf6PE1WxfG77SIgTj1K7Eqak+R711t3DsixbrLh+1KDTa1z8sNudGLT1GogtHS+TW
jJF/Fjd72AOKJTUgo3XNEbAeCZv825ojuvBTmNpQtprYMKKZ7Ic1el3rSPwQf7DST632MmNgDcG0
WuuHbdAQP6SflMOVhVAJGx9oanU30b1ZWjee6piSNjsM/DNrRFlD+fOn4AmZ9C/YE0JY8eVBC+PD
54dSLtBi1Ba1JbxI6Bk3r10luW61QflZsWkdhNivyjkmRYJ1BkcUsYYioNib2EcsmU2gdPJFV5J5
dvWsAkPyxHY0Tn9LkLCTsUctwk1C7EMfmn3vpSmVlt4SsbpLoh5xhl1sC+Lf6smjVUaE3C6vz3Up
UYdzExFOoZNygDkJbx77AM/bxlNfRtkL+FyUAjrk5cGmztm2iUbR0qrrRTB+or6X8H5tSNc4Xb/X
NOuW9EIzO0O0NBYdIIsj+rvkGPt9CvPEFFsouIGAQz7JsTg9JDlbEX1s/kNLEFhBlHRCpJA1KdF5
ZQSzRQTCt0eJNFP0rRFmsQjbNNxQtaLtDGvizISRyf5GxgKGWAZ+dzN7bkGbhwCYo+9oQ/NAugCf
2zC2K3HgxyiARe14yJ+UC92MGEtkrzk8+kmSWpIB+9ukS6fDeX+cNXuVXj9f6jso9SWejWSwfklD
CIPn8fsRc6pa/2zdEbloM29V+R6Z5u7hcLQ8HfMxerMMU4yf8U3mT3vZQnhFWep4zLo78boNDDkw
kpUEzY7Aug0Ac75tq7uU6vXrEJm0xhFXTKdS/MKJUYVdQVK0n2Al2GwebUmVezGvyh3za1Uq3NQ2
42tf7Pf9DErfzqiWNgZEAK1qtSJ4un+Rny6mvZ4+MxHyc+Ps6GG6BYyPpjap+F3IVGPoBkl+PyMX
GCTGcWu/cn8oT7ZLdC2Vhmf+Vf5YQIO4hZ7uvQg6I+nG+FjTT5d8i+q9HR04M3v5c/kZJ+K4qorX
FENt/S4YyP0Zk8geKu9cWvgk0l2VN5Mso4r48JjV6dGJEm+PJNg3LZ7Bl0YOnbUfE+dRY47aE313
El7xk5CZMXLi0nBidYn4h9qo/dxp3gSC8kimNGYLe1a07zcF6ZZqGlVw0hth++lowv0kIUWXQAE6
CRSIoVkvheWesPXebq8V92z2ez1wIMrbiiPQPjwzKzcQIbAdttQeHYo8Y0TS764CZzNEfBNYGTZE
lmw/47PRklqPuDrW/qknYHmmmRqjL7222V5h22rliaN9RYvlvUtvdY9xV47TYbLjpT+DQzOae8ow
BKqMNUq8FfGLYe/Ek7qPO06vSSUWLmITTrCHj1/2aGHos9AaJ8UQPd31DFU4HTJNV9wcXzdizkWv
o4sCh1iHJtdCOQMe5wA7lFKY1XUd8tGKnQPDjT3SDGIh5d7c9EkGBQhgk95oVIUW4lj29pPZ1QrL
JK7Hj6L/KC70QM92llRbQNixblvnDNBDcNm2Iqjn6MwIgeM3qwXWRnJJjFmeKGtOOAZzX/MrnNKR
ZlNXvwRYu7k5yzvAeBY3bQgzZMQXWFstyiSkQYKYAWI+dkXlHZLjDdf48Cy67444C3OxziwualZV
WIe/d2Obl+8pCeDVDI+0dJWtynIsDl1/WhyUjJvht4aWr+mEsYSMd+LTTG+9ryvEFvHuSFEIF9Mt
RTfYXnj08iYPGr0XoibQqVP+63/jZ47hlWNIY7X/NTwMXEzVZK6GK8cAKp5RUb6sQ9N88qIblpt/
m2y5E1QcF6zSBlpMT/15+CwFycdFR9uMlEaOfn3FEgJBVNcGytM+g8VlsE9xEqWWbNTPQwC6hwfT
h0p/Kf0r1FnpXQaR3wvN6npwRRM8t1Dece8mCcvUUVCBTZ8yBMle5FrsesdbuFCk4kc+xf90oLRX
M66oHmYvywuknLUolZ5iKrbFxYbaUqxDIA9aKO4oofQl5G6fpckzeRFxtJU5Se/J+mcY8pnjwIbn
C/lRL5m+uvhlreSxdkBEjWzNilFMFt4u5pdirhHPB8QUzkPldpztSj2sagnqSEERpw4jqvrvBhLU
y3oyKmiXyvvjBTAWZjhhMgBZk4rOmyWv0q0dUyHO0O+b8Y7WH9OPhJxOjkIkaqscP2m4vdR2jlOm
hDV9KA/jw+RS80gFtmPx7MioIC2JgY+zt28/ieewmSD8qtespk2lyGdVOe1KH7peBn3RwlGHH5Bb
fWob0JItdNYb/zZKCYAVOFCLZFP09dLmsCVlh8t6dgSEI1yZSjiIKk9JFgy5qheTA6dlnhfa667F
g/TysVaWNN0/Twjf0/XOKW/x6aOqb8hgR+fxYK2ii+UURSGcFcHNMc3euIOK1UkVTWXJ3UIH6N6o
jx91T9vYSOsgvaCznvvbarw65an7jS3Mnj5yTFshcLtkRa/qzfL879dFYf3DIw6vDuQwcY6crCav
mlGAaB0ev3BLaT+JthsFZoF8Xc2a2IFqa2IE8tlJ14XK/1CFT6W9CYA2QR+4kC8zCiDVuq5n11V8
cCL3dDDxJfqgV+/Ekn5ao2W4WuklZMr/xDoPHHRtMZJKVK5ue+k4lwsrUuq16qKE+RCQDkRWO8im
wxdzlQkJwmBsJFvOqy1qSZqx8r7FCnc1CmgxWJ4zU7Mdc5EDvHvHouYzoQUXY+gbXUxQ2fHl7ZAn
1ewumDrHIE1bx8HHMithZdpG09dBH+K+qF+CDPLTyCI77nnJvukjXprlqYPXS1SHcedzqGe5APjW
eayrJYsXL5wPlXxWrxvD+zuIVeByzYRo5hkwpWz0uAKzWoRXC/W2Cj01OWsjv2z8OCt1OSo2ORr7
+VyK29fb9VdjEPPKRqOYGtihbDSpXR1in1IBCSkp4YCZwpCfBKQlwyjBX07Z4PXOhIrJVppTopKb
gTTj/9xwUJOLzBOR016piShfQcSiarwFjXC7ka/z5MUjgcTCH8GDx1vxLCzaKQ5mXCK6/AFkxC1X
xGB5KXFt5xgkXgCQCRwY9xHXQKlaf90FfdEem5iVDWHAzLLWCl6DeRPybEb07HGtZJCmiRFRRvFe
7gUvxOeAUFemBnlQ9fCR4C/+VU/5g3oe/hYQPoK9ZvPXxYfzOaNhWZFZjsO/yO5Gzf0yY4VLwwje
toEqFHINlr0txyGnKh60NYw9yd+JHBIQCBxrgZz7wDxbWtQr1zHSVvm7iP7Bo1362vY3zzWhBxLg
i7jZXK0CynyY5piFXoDveUfHFPsfZj6oFasPY0A9w+vWcTuh37Vd7OLyWc/1Ra8TI/85enncH/cT
bQryAt3s/25K8hJIWR7qAhMqnyfxx/mY1jam0bpvFhJF2R1NsLIXcA2DX36kIYhoeJPzsJNlCwUu
Ch+FaiKnl7fnJCaY30/eLH9Ggv6JAKq66Vzezb5g/RM4uBezLOUdKLH4je7EiBDZaSFwYxYUrAnD
s+rzLN5iXLBoQmGmae+gKXLx5UERklKLbOXgZxSpJM7b0dLyi+h5dgMngB2TQ0ZKiFqlDDT6vQNA
X9Gqh8yqIPsr5LMUKDAFmEUBeR5KR3NdVwSsGwF3twtiff1euCbTDZevs5AzLyo9IZ73OBwjCNaR
7vODULhnK8a1LKfKpORuqYqfrp6JE9GknRsOZaA6QCGOFkT32EErHziPXVK6WfEtrOryrSTgAjs0
iQ2dGks86wU+do7H5PIxPo55C5y3ifQEZXHp27y9hki3eKndwJ1Rwbj4DiZlMPqV2mbGeaQxGPx3
O939LUSTAr3JoYfi48K2Zd5l4DQR1pHQXrvESYBziLyHP8DMF1HWSYRpzCQ/ilIE3Qqnk6ad+YUM
qKWjN+tPA+dNepGvGcsVDEg9yfqIS3paYuflZ2Y4VvvrKWJUYfgrqEcENyxC8fEoqW72b0VQHUXy
YLza0bMThf6HbSjlYYVEMPOgEww2Rto/JpSW6Rb7iz6vKH1b2+B3UOPDnAWGQwgTEQICcXR+LkXb
iHgNtUKuq8FDQqxP0JF5SiJSEE83I+dho8m1WF0+UKh4hzxIC7v8LLMv5toOlKruwFvBQkH24064
UJXR/OvyRD5xbDtrqp0wAwG/JWM22hxTLMeltFmjgYtIhtqlQBl3Sls45ysnChzYrrVKQzskdVYB
Ed97BxwLkzf5JYnsntXeR45hiAICAORKY0Cq4hqh7lBL5p1v1+1EbisI75VgUJEyWFso7oY0f9bt
FT4YFnZEJdPNfjikOOIZhkIvzTM9QNiAwGRtl57vjH2ZBgHuwvyCg0RN1L8ooqgYxFgZ1Svf7x6n
Wuhd34LoReYO978DrRpXHR4NqzDV1bNR102iQfgc8fb3gndUO3Z/iHqVUTVIor4jZ/wEl9D6No2v
WGeHLFF3ueQvDs6Fxhrp6YBr41/rph7Q+1uggcvdeTs7QFPONWu/Z95QNPEM9rlqlsS5w90DAy/x
GxeCy5rqcoJitR41Tb5pasPsd5KtggBcxd9/KjjGxJvmXzsrZ2HWcOvpq9ubSMVIpOmHVO4o/bCp
avXkbYuZekCZAq9Ti6eXb0tabvBHoEX8tvCfIFwa9GKnaRQ0LaDNeYKpPG8Vmdmx479hpR3K374X
DlXzLy7oRCL/tUd8FiI5a4J6IPp5hnwRiS6WfsSkXJVfimwFXXKByjlzOWUTEqg5LfA1Z/p7VmJs
RJx5/N15vigu0x3uEqHz0fiEsqRO1YjYO8rClCAxo6lcazAOOxhpbGQlSZzYUnQtMfkLlPwnnPSq
d04qgVboHClIksc29bgsOMAnZQIuL3cJKkpzSPeH/nWOCN6/Y00kHrSPMgIybDXhV3INiyX03vUy
83mehaUJMbr9s2TKEkWgxOYtIWWFMa0Ea86TXYKY0xlMqYTkiaS15mtXAqY4jTgR3zuz7+ho0uLJ
0ZntrsG92sESid34c5ZBJEfw7di9t7B1bEJhiIXzk/yR/d2bEv6wiOJNXvuTrj8TcJCGGPp5ViyS
3fawWd7Qh+Wmtkk655KGknI4O9g2bV625ZPG9T3AXM9Sq2yIX3LH1lOX7kO+Yy4wfRq8Oufal/8Y
aopxgeDjxWzFp+6mcNV4gbi+mdomnO+sJR8yqi+22HIgeIqJDh0JqZPshak+k4fofnbym6AQxeHA
xIZs29afjmI77Kwn6xl67kkeNuZOyQc+2zYX5foRvC/EuTd2qvjyNWbxuNLnhRJvfdfAaXvve5eX
Wjb30z7GowxcSCS+dlnjJ7LdTAHJBFLkvUeO2bjsVOHPk8mDdrh0XdVOABYObf7k8mT+NhKO1KUO
LiCOQyenN+KMmJi39dOS2UEue8REpIWmFAZ+i1fdRJhZdB31sAjgiNfsjlhLeHifIdAkgDPo+kIM
8yhN9e/jfBUe8tAjNKgx4dRHUIJ8FvhSz4VRGG7vocuZOrJF6BzKgmzbtnulempBvB7CKixfutZQ
RSItqi9xMWKGIh4Wp+s8jBOPBDDiJirjrbuR4bqCP6pYGMBuC5nDLznepNQRzwslinBTZVYF+PYg
xPvcZidIpHni5qJ+z70QclkccuTzmQQSyEyUqa1TkWVb9hPW3+8bpn7SRxw0VEvYPm+7TOhMKI9c
erkbn5DwjIXWIhKT1ZV3fgJHpwhrzN16gWMrEYm4H9vT4lSmM9hN/p6eclHekRs1GaJJsmrQh4UP
hLhZ5YA74deHlAzToZ6VxDeszDhuHESMbTlvgu3OqoscuIl0LPVVUWfGDZKktIobX4crNGoXNtW2
ycTZ1z1PN5E15zZyNNrpFsEe2S5aMGbWTmwJT0GD/7jF28hMnATCz3N3O6sGHC+NQIRDCKhjVnyt
M+JECdWH8yMCqqUT+STMvuYQvrsvOV3M9i781md6UyjO6zyu/Bg0AczcgWBmmuqQTBNgTzg1QPOq
LWrGC/TbptzHa32GB6xOgO1h6iN8q91jNy3YDvyese5S1xLTRZAPdppH+ZgKo4NkPPZ0b5riNOhR
8M+gKNQn+ysNIMhD3h/SKW+6SdhrLlKC4byxi99govVrodm5ReGPQHxzt5DBz87kigUBnNeKQakI
DPMJf4W0l8rnmVQbd0LQRigCrNOH288qrcVFNQQ2krmM82PeR8r284CTQxV1pnxsD7oeJJ9e4eRm
w/4Xr+ErciRhFfiQGD5IPfBBytSvuT9IQ4Dk8E0SJT/4HS1iufym6PMSAE12q95WxYFf4ISwM+vU
bRNovo9gyr8ad4B2E+GB5mI2xCFp1BrALCKKl84eUvyEKQuCMi9oMqNdgFwNL+sskoSCc9BDmG5Z
xXD1Nenv1W6SyP/S3lt+9LIV9Ot73BvUz/iyUvVlFJTQ3UUGmHgLDgvwD1b7Mu1vLDmZN0i/aHpg
n96fQceRIxKMYl3tDW0SKJn97Q5lxSE8R4OeQUrAhLCW8QViKJps0ZQj6u3ol/8W2srcYJKlXdO1
csvHlDctftyeU3X1827ie/hkAUFPCWBFhfjGdlQj334s+cy4audz+1zi1KHTVV4oshyfPxUpGE74
2976RW90C824WiQUB55TrsdjhAm1uek4dmGa1HFCYuCi/Gnq7t6z57hVhddZLe4cEZ4YU0cKJunM
L117Yu7z2iEic17gCozlQNY/5vfPiHB8yRiv60q9YUzS1H+NZKlkqAzmghEr7oMHmw6hXzzpWgJX
/bf4cdorcZQ48aZq7mTRXu09vWXcA/kwEJs48dQzT6d3exDrZkMGVxpefWwhEfv6hAj4jzfslxZ3
7QNf/R3422jubax7IS6zJVBLlKeDyKZ5iFwphllL4ENVhAcQGgmAXO7R4jVsvLO5eu7cA17x+T53
uYRzSFwdUBkNbvGCa4XxA33R5e+plmjaohGGATysRz0JmR2AZVvU+xL52Cv0DrPEIw0Lgzss8cmL
EWdv/c1UmLNS+9b5AycYBeLkcvuqfA0wGiSDlQBwHRpB/LmyG1QGSTGfQcjLZdJwrYRXAa0iQARM
b08HZIOMToQUllNV9xFp9LhUKVfLFViwE6oGWPQZ2HLr97z3JiY1VfRV6Wb8AYOWPSpByQbgH9dA
ev5iFwCJGnu9pjAK2wDR1+tKpV8QQE7P8Uu4Nyng6f642On2lqIbcw3M8k/GqUm3tdUBUlSicI+T
7oABGdMH5iVB4tVDnEZJAVUFTvlw/g7rzeJTxfMAItSZKvWtmpATJgUIMBnWhGA2OPz6bqIFUiYa
pv9Q6CkT8Mi3UfNvyYYSuL+nLL+C2lEdsm1Koinccv4L1LTojY/m8LlqPJ9FgWzSFywroRWtMIIr
ZUCfC7NEF1enNUW4+8LdbMfrzy/VVZFpu+6vfznMBAIBSgQj76buf1f27imcpv7DIfhYEsp/tCSo
oTYb48D/uM+cmkwE7t1O1LPRwoUIoUfzVAZ2GLSy/2L3MBzykHKcm2PHX5dADchX6h16/2AmURt8
OgmMarlXxZZb3ebhLR7x8e0sPJYULwcd8stTOxOaQLpbzo1QK3PUriHTEjtUtWQiwQTZRN51K9/r
XOywj/9WQXTc2bg/Y1a9xZ/HKCKEijTRtgpPP5KuYUjcEflGhw45sJrHnfsKRPxG0JYJJavEEpat
UgYu8WewdraSrnKRdyixRQHLIlxQm3BDVOmQ4M0a+MRyih/d2c+HcXfs6M6S8OfVOpbcEU3FgHvi
lWyMDdinWNQlLfi3LjuDpsuWcMq7xMOUAifdxwQgP9mGQauUM+f31fAT1Ur4RFOKrGYN8pe/ykZH
tfzO1snuWQnGe8/NRCH81DukrIdGBggfYNsDEUL91gLW/jcXekMZUwuF6IXo3eDmA23kjC/Um46D
ZBZMN/yyW6WYrshZawYjt2iMd6/vYfQhbRNrcoxyfff8d0GAwzlBuzkWMiWRSpV8+Rzf8ce9S7GV
Use9MNhiD/ySoxPjDq1+iFJDi+/ANB2e15KBkbiHTkISI/BM/eucK6won3tr4Xba/nUcaF1QXJZc
JpgXRLtZ/eN2NGkNpMcw2MASn77wFKJdrHdXoEZ280jLoiAQ59VLhFnMOC8pObmEOqhiZyPYQq9q
VGh69qUv1hCjGnDmQLF+ILIXcs3oJs7/XGvXUigjF8DOnzJLHeP1/jsy8c+xUA6I5rpokgNJRevD
EeCk402aK3CWNQUp7dkmtqFuGsOjARZJ9PCQy8Uf8zVqS7k2j++I4hU3uYyhUKX2pKDNFqyIx+VB
4hbRkb2DUUOboS97vG39RQKhx1l7LIFkHZDelTVkd2nw5HY/bbRa4xnCzY+ISUCBSaz0ZyGT8paV
J2f4+PNbz0jk/gHFRsTzqxOTKbnJOg4YSxFycCDmZta35n32ouybrfONxJKshSiO++75e1atx7ip
hHatS5/ri7vle08rwyv+ShnmtHd68N1fk+w8WIWLT5ZsWvz2wX2pD1IXKcpsXpIl1QPqtalXEOgg
ck/+70BEdmnqAZay6inlT5qfm3tQPpdkEFHGCga4MewH++I1QP7kY0iJZKAKinE27NJ5OtVqdvsH
SG1p9QulH5Pc27yNaSZvlYE2KaZJmIkpbw7s6LtKPRLqTTx87N4LcQfxlMswCxHAmklODhZXuGDf
Vqey9Zv6AwSAUvlVC/iw6TyoHdKWeu76I25M8AuEE44ypoJeDWYHjtBSGrB1ZYAZL//oe+fbQJx1
tjL561cEOfz6aOhFh/YWpL2YeLVhyhyEpvCh0fkQgxuSXbRVDw9ds0IrUD0R1mnB+EVpo5WRNslY
buoMTZ+ECBcMFMOvV5wJJTkTVUfd0JRZ1we0Tl22En3W938fQ0WhDvSL3UDhfetvDi74o+79vVR6
qqI3eqEuR3tVagi7Qh1Ommbq2t22KAumJwwop/tUcGbiW167nnt7p+uOfgo8cxjOu1Geenyzgfs6
nfuf1uWL4YTzKPCRPVhse1OkmNz6exBbJawUDWwizmnYXbcPWLYjFrIIZCxX9QXCB33QJYn3YoaL
2lw5HOxuCRJrGl5/0s0sYkhEBCz1rfNcpXCghl57V9cpTb42wNc7qzgocu3jqaAJtP/f9sXPxQqo
OXJYQrttRKlsVdjQFlqNARSxpq12tbWTmnr6acn2Nj8E3PKFe0ZvRSzEU1lZ2wiwDnHEnIOMnlaB
VYEfH1L8yO3M6513zhHf3D5gYrgOrTLaJYSuSqMQh+LOuYhyu3IcWV3OXeK4wTe4jKoHjeNL335e
4gvlgVHOdvgWT0gQq15ZX1RntSCiEQlvoZTwT44IxN+wguOQ7fDhwX+OIk7UyvGJ24bYVq0ggpSZ
Fs+dOuHtIO7xBGPBc5dULODSTnNh+Sr52OGyFdedhuB7Bs+5jSDIaOyKRbTzkoFTF+X57r1KSfLI
mR1khavaKYXUr50ecUxsH45g2Qs4zTgGxYG0CLoQPbrl84heJYXPiGxplOTZ5x36/WZnGdjJj1c6
1eRZoADj+0f7hXIlh2rz6rD/nLWSH37Y28QF+akuTpKDc1sUlxEfQ4h5Dqk+zxfxVZBORBT7ojfQ
X80BOLuim8ss466UxsISo5wg9ZYuJ4UnTtro/JOrqIdGCyIzL6lZsIn3H5Jykvy054bjczyrUMdl
bgc22XAdPRWmI9YH7bwRndqPXJx486zwPNmFMX52QPzYM9BvnWsuXfqYeoloA36ZLQgN8T8KO5pK
s5i62w7yQ4fz0ucPqSc+Iog5CmV24GfL1U1XXf3yvx2QF3Oyu5LBo0qMDAXE05CMVkqimDNrD5fs
95mSKLAPH4uQDqpATD29lkrRCSRchtkg9UuoLvFJsL186Y2rH9dqWVFoXTnypqiRIP01qbwZzP7a
rYdl28F5seNvxqvATnlBfK4Ja2zMNgsw8pYiKMwXksRLgpmVKOSEn82iWf885JFjCJLZZ4MN8UyL
IYwEfBJGYD0vRv0cio2PKtDU9T3OzVpuSNEE9IgWfp7vBo0wbV9LIM4yRxHjnmoufLjJXHyMYz6o
ZoorogDDACpZMvaJHNKR4se6mA2knILrzY8LoZw+h9EJwELODl13GF7Tl1kY/D9cwY5maqYLywtU
GDcp7RE4UL7K1n/WfkzidzhjXgtzPrSQBDydZjW5PWNuV17PKnkEhzW2XLfTFEOVMA2VvdFQE5x9
prQ7hMoBkhlmcGtnuasPjfQwhJGvYHMi1s/T7RVzpkkyAxNQsPI+1whhYu2TiJsXYPn+6UNTMgeM
fkSMXLXbocrosgT3CNTfQMy5cAcv63mBAgFoL6vklYLJBg3GiuAEGfm3xWK5I9MsLgfDd3YaAxCs
Xbn2vcoM1XCQ3RJv599Av1VnMakIqC2erNI9ryFwlD3sYUuSjgG/nIW3xOilCtlUFknQiflqH7H4
Igj0JdnByd/NuXBaUORBpI7gEY30Ay6Iip/+l4u3PI2t9UkmNWpQ4YEjiNIor+3rHINa51FoENAJ
ExVbdJyC9SCOsxHEWWH0gdyp/cHofO0CrVeiMnpF7IMifykRnabvXj1G6vT0TFZCWtzielPbhK8T
UUxYLzzbfN8bIhcVmLsQYa8Rg4qknKaJF804jB5USJWyLQIhgiCav1ielcGTqlGs6H7Cq5TnIfQS
3AGXFAfna44nlD8ewRvgLSONGLM8bzgW1CBt5kDJ10m+5nty3E6SObHl23z0/qlwa2A289h2iduZ
5mCy/zrXLRQejmbYWp0DrP86kAwcLUEkOKvb/amKMDx/KXj1CFvi4MAtW9QuTRPgmNLO7pjEyfez
7P31kPo7A/Qg9aKZgpjEMnYrdxrUYuFza0L1U/vKoRfLPB6XsENgqyiwA0W256NX09TXSl5frJSL
7KukKy2Nhc6+YDS9PkF4NBGONl59syX4b1N1sbzYSEkNvTXd1vEkHVEmwcZdtgP3b1DW4uZyLlfP
QpojKCFczNzN6FlV69RrUu+2OQyPAaN1P2+Rzdz/PgtxLXZ2fIwChxCvXcx08STWAxYV8g4ht8ny
LKDec7Pk1xJS/axSZ1ovO3wvf6Af/Z/XEmc4K5ID9v3Id6rQUHBCKUTdOTRPJQRHtjgR9cl78MIQ
OjyC/sHCi2CCikCVVOnb7Ori3XWrUm71iCxUBBP8zamvyK60yUVh50sP51zHKEJwesVzCfV9oRao
D0KpXmr7ZnCkJWYO59qpxj95y5UK6kidW+/3mL4+h7H7xGss39bPwCmu6DW3/chiznOboUwEDfJx
iofIF/qa+hQfx055+r/HrFvKmuj5OHepNs2gtEevss2XRD6uMLWlZE4IMQJNb0k+ZA4p47141D4E
+O/zNpY4YKI9X+QKPuNgOhDRpiV6l1XJ7BNKnN6wqH3b+O54HCxAyLd3w7UnTYWcmMO47A6co6eW
28eOsz1IRSSicIof+p0BgBp1EmANXzcRMSoT6woUCzGQ2meJCyEtX++ZKbjlFrrK3sLM+BselgTZ
e5so+jCc/q3tjDBRDiWepI4OoKFAeKAwu4qUMhfrRDaTA4EKsentQo0oj45hg81YF/h1y8IXuSGV
39Z3FBDik4ATUmHAdkkm49fG5QSIzzTx6tGTkqX2/15+RkjBoS02rpsRlrodJZvTSefWoFPXe+yS
/0GuxiVl62v1R499aNJhyq6kwINNbpSghVzPTkAPPd2OIkzGQvjlfzKdLKzOVf5XsBWhXwRqjZXH
TUxi23kJVN4jeAjDJeWvz2tIsVkBkGnsH2NQbqrw7+vXWZpq4ruVy4oyY5LlPPxIIAV9gEoQJdH0
q0OSDFPdKHvsL/ONHBZN1+NGT2fJXUyh9DcnqJMpuCmVByhwsldjoKWwrnClur5PqjNJnRCQsi0C
wmM9JpnppfIK+9AD4BCi6jx6LHAnPtPwcu6dQw+JEUgpyLGbksaNmiKqfjwxl75rTa12UFkKSfY2
9Hn62Grhd8Izo8ud1XJJIY3JYoA3KkmWaMKHPHsoSAWLbmaFoxrFTRKNJvKx7UaOmyxU2/xLPZDm
JqzNc3LE8SmmC/bVb4SkZ+fDcABUfKTYnZMGxI3ox+57UG7txH10+QvjK3Fpf8RIU3FjFb+oBBx3
1vtfFQbNX1p4CwrvC36J8f3tcDP9CS6ld4qDRsV3sA2NRDZLLKa8q7IiGWpsVnNLmCYziTdFjEg3
/GvTIdT8j4P4nqAziNyWSnF5/9EoKbbDTofu/Rj2V6qbouwpi2Ra1vAhNueiKy5xFt4AQ/GYpWfa
i+zlqVCsBVhRoTy9wzk0GfESR5JL0k6npCwxDDJv/YooyKbeDxVhMsOuBly7PNKDFyPc/BjMlL6A
9hrEp1PNt8aKhMNLi4aZdTli4TYwsKhrXseNoZtEaAtsutADi7/TDsEEs0UG+i0eDqRrP9t+TGdw
Kv20+7BYehYYCvgGuY5ndLW5olLoug8o3CNtFvuBTSRVbMhESQ4ruMR2uZTf96sZNhEjRoPEF51E
qnGkKWZmIH7dPMphJ2NPI4VSZYeBgCGwOtUdjNXvLv4NVBxEaiX9N0/wUFwEX+oipLlhiMju0yCL
4XE6kxfuOsNbmlLKvfT/NHnPdYu5GsdcNHtbDnKnkmQrausQZKAiEqToPX4i1E/K59NDrta7Tz30
5mREgbB4LjMLOtPYII4MA3Iuo1BqmRRkbuayxfGwbHcaFz7Ln2zY2j/Bmxima5P2s2xCfJQmQgVP
3GkN+iqeAr9gf4jx53hjmBcSsQ9YwaqIBZheXJvX2Hq3Bi8bE7t1gS1bVUNPh+OhK53qpIJ+kMsx
3wpT/Ux68K3BZYAwpn8kLOD+w2yYJfQPVxUMtug4q4qWji17EacSZgx3/pcj4W14S8DNG38bUxlE
2g4J2+1Pcw98vPk8XQI+fk/FZt3ShqoXWovTEOSeZYPdfZVjakJiABpe5tllN/1dTrX+40OuE0wj
yD/+rQX63GoLBjkbeziFdOsbeiTRgofsMhho3tFTpTQ8knwn2YiChAOdfaq1L5lo7vq1cHdmZ+vj
jXc7v0qJYjS3/ESzGvwTbYn5gHLhQ+ktYP8M51MyCi0tcB7uIGl6fAqt/FhrJwWU5LN2xWsU83qg
lftrkKyi2O5i612Q6+/+Iy2hPg3tD4wYZSLUotLg+zhZd+7SUjn74S2hradL2oFKMIFro1bAT/Sa
VNEqjaxV3bCYzlKBkxJEN/FnjdssyfyLReXY0pV8z6aJsIoOakoHx/Dg+3uaU9TQiRR+7OEyg081
EzJyK0M2L80ArrNv3zxdCZxW6MuUOiBloW1w3HtBbmqvYeJmWoCYlihOQRvwG/YJ1Jv95rVT0Rmx
0Kc28lB4JOhIUg71XQ+V3MGSctP2xlRPSGjWyMNK13qcNfKiYQEtVwsZkc8ne6ASbriARzpP5Ccp
olXqcrh0Li42LbItPD2MtGymUuKEgQtYoAdfdCyT6LmXFeQjwTPLQ5aEohihYeMSoIyJz35pwWxC
pLiiI9mG/4cdSUH6ue/EiwetMGvYNNTnZl8LrCFkph0vIb7ZC3Qw8NHQRxTr80rvcJYeqNrmZDtx
iDcxE0PwNSys5h1kQSuz9CZhIYqcc8o8CmYxAkOypFvCm7wTWue2skap6EAhJ2YJBZPL3cmD1JAs
zC6bbY3Tm+GUbKNOL4XHbR1lIhhHB2K7qK/FaTpGi9tyt7RT7A0cOo1h/nAj5q5XeMuen0M/VPiB
JduwhFq/QseYoDki6mDwjY1R+A72mLat6ddU82FoVwiGXZ8jeVfRVnRXRk+4y5F4oooNxwAVp+Km
4C84X38+kTd+e8meLvnm8czuYmv65tO6e8+TIlZ2ErHTE4uH2PaIvwbHwAWYm5jmr+VbvNic++Lb
7gUJ/CqW2LEExn9LYCE+OQg7LB3UYeSHN0RIrE0OCMsuY9zHCMKnj+mjS9cPCf9MUTeDOjHIo4BZ
vC+5xIysHTGBhUpyfJB04fHcG1Sq+SKSw0BzwqhnxzAYfQib0DV60O9sWXoDhIsCra2zZenvIYDO
GIs6or+3LU1+sJK99KWx2qwkYgu/CcKle01df1nQ/HRyZ5EdLXTn/bTGiNpXAaXZqF2rAeURay0l
Zjc2tjwPJ24hwWapvu9oQAJ0AwTEX+M33nv0QER/r8ljwh5iwCEN0sKW5zSJw1JRIw23cExvz9LH
scL3BDxFCo3pOks0aCAiyzmx9Y6q/TswngkmQnEuzLZ/abYw+rIPNSfvrq/9+/9yagfjernaAYId
PnHdUekV2CxIwLEA1GIrsc5W3ruiXJ1dKoNGicINkNUCAsu/eH/X78pAF0r79LFKpyqkfJedPyGC
1x3iTbfNkQ0L9OaVEhE50EMIFbJNFemnvqf20fvJHJkr4DUaYZHuH/a37iryg/tp3VXqCtU0WlE9
NxZMk1mOwfLbJhLOWpLXn9wv+mNz3zKHyT9OSd2xumgojYrxOqHov/SarnwWo7Z26ENoyrZIJXTY
rzy/G9ulmLo40xOdYHY1tkU5c/ugC+aLhdzghAQ8H6nVvXuz+Vyhv4oXmQdutBij1GEhR9wuW96U
CvCLNsadK6TFeaLl9JNg+rBGwxMxOz7EPwc/QGpgYMvdovJSwkmNs2UXQlvaLKOp12EImvXBLRNa
XYFfqmZZX71FJeKaLNKkdHUSHHT0/knG8ZMj9Yssg9o9vpkIxU+80UdxHJMskBm+/spz0xbYBTs8
MZhHTgx2SSdF5KlFUIURKoj7xE8U1vl+I++r+IMxxo/y8YgKpiyoBpetrvM4DYFYIdc5Uuvmeu/z
s+HGcR8Wf2rltvsJeM2qUo8JhaPW6HeGfkACUfR3K3Ty0uOllYRb/lzxjP4Dh8PFjrvVUy16HY/D
SyEG9QSDZ+9jzWPBAbtcTK2aobzm96DU6vjIei8nNv4g3rPies17E2RzOqboqMvUIv/50xJBkWXN
p3juvGJaSHT4ZT3WsB60BhFhiy4ulFBJD84PYy+e2R1CMRXbQMmjs85PGX5/fuBB/wPQ+G+Hm7n8
vQdxYXUJDhXGwrXiN6unYR7LVs8GgeA/HBG+uDJrOMXGjYzX1lxm3DeC1t3sdWXSsBVZyOFhILIh
k3ogMf9lL8r1h1fjK0kUrPhgdSVacnsumXwru3F2QP9Lpqzbr0Iwos0l4c3ZoYacbaNcu+KvKSS6
FMNAQv7TVdh3qrHBIdapnleBuUu5IL4Ln1LML7UPdE0XBpEzqp1bc+2p0uI9Xmy3enzNceg81y1I
J/VyLq/75ekFl6lkWEK173M1bOqbFKIzGEYHAsAXsYco31XRd+osuOyB/RWAUVV9l824Ptm4Zt1B
8X0bjI2ypbKYzNDB2IxjmLAdOT7a/KF7XmejBCjGcwDVm3/Wfe9NpsKDK/5p94HxqP5zI4CFHhqp
1eDhbdx5Ey6/Pvic2EhtlfYlPjIBkqWfWs11qsYxBART64Cj6hWTjK2SFu0kQvjtCemJ2kEBauzL
aj5l7pOfIYKVmwhmmBCM94J4hm8Vg8Gnt4dUba6xC5wL74Y+LCdb2JIR/ettc4Xx1BB5Br1aPl6n
BNo/hotWDNtOe1zFAdjH4bWnQ5bKh39L8QF+ACatpwy62Th0OFm8fh74M5ZNKOTb7+6FtsjwxL2y
6Jcg6Pqe3/O+6UGo07fnqsmwus7Z+KC1De2Twy2oYKOj6AZ6t3FEl5P6ulDcrWvfDKy2vaFHrlx7
pr9H9f7rJL0GdK+GujTSCriTx8socsI3AnZyeqzEHaSzoh+csZaavifthO9f5QR/+lHhmnoZQdif
csjqm9BCmAR3IIbOjLQaTeIw5LBZDME0ar/IiKC84tWfNmTP7oCmvMU7Ic+g6jrVBis7CuAXEx3u
mtidzFiYVbphoAu8Zq1CcQdumJzX5Op4gqN7IJxPwdKiocLHFRpNWkKhraAsk+9xvD8K+7a4ghPM
smEEURVDzAJoTXTPyHcwtH1tVPvWYobnc1q1e3PqnfcDC/43gmsQmwPtkB6y14MzHJtUzBJHQ1Eq
Pd7AGmCoFk40TMIKLE/htSFpj9oVAgDk4/WdSImwcaiGk4KRDKjUfctbLBXb0NhJ2y/gmwpxshuO
6EwTB/iPlMW+g5DvWZ6ArxQK120GqwdYYOazYwZOaUdS1N0omZSSTByhOLVnVQ7NnTUbs+VL6SWK
N5mu2uL/z9r7Je9aXraS7HJTNaDCL3zTWRqmWYbJMGu0uPrHGJeINeOBB+58JtaCPgQLZYSUDdbE
d2d6bd/FP3PS0VvpdCd7X5KSe2bhmGfGTiR7XBidsiX4JXQMa54NPrF2gvidu6aHxCeI2JU9mZAo
uHJyhCU2vL5jvGZhq61w4ArQIplW5T/S5ral2yRHjrnBNDD6fjNnrrzWPg+11y6lc302o5NkVqUm
QC+lHUqwNsfxRfMSNaGhANsT6OI/+t5sA5Wq2aga0xYa5dfkXPOhgNt1CZiLdrUaUNlb0N7J221Z
TYTyFfP0o0ARg76d7A7Y7euFVHj0wAv52YQWEML98+b1gSZll9lzpsfqfs6qtBmJF/AcDQRoOQ6a
Yzm0dt960R9tNt7aZTrWzeB/zn0byeV0ufO7HMv/s3X/lvvvsIxBGWHab++r8ZfgtkLUTdzMVyzZ
/pWKd++XCh4oNA/cEBkBSb+PybaaD7kwnq/YdQ7oJS/M2g7M6lG5VBqNqbd9YhD8JLGye8wlSE5Y
aPqR8WPQw93k23QCMOEY2WjoL9qP1SJRWVg2iSez7KVV6dMwllrkFrxR7zoTWOdjq4d16bnyRa3E
I+J8G731aYk6577vzI0wszPXK9U/eQKxz8ivCDfU+xjNGyfDheVR2aJDFXsX4UEXjeDL5NnJwEyb
B7DXVB8ACNlVkmS3NVQCmYLGDw05NxrPb+yoyFiarxnGXbMijKXgJp5P3rjI0Rxgn/MOS/9kjbyD
b9QBpCNwGd6e6UiUbLPHH60SRrnqyrcD5ZLq5CrP1JF8RO0S8uXZD6bwwlERWbeKMbxHGtWu7yhE
qbaF3/cFbzpQFQ2pORaQVytGheIJaKwitxNQkNpu5fjoJb4J/L1p0ghPQ9c2JTC+IwHo3u3r5lXB
GaAkIumUzLrkFoyiyGYLx2pQfPkM8o6BlgTEbwMhKkC0GTUQU7nZASHpxAmWEv6uKVsrPsik/Qsq
AW5xIE6U3tHn9jfH8B+cEU34KWUaJggx7joKOCXnqwyLxJYIZHL6jOX9/yCiT0A0z+qoQvj/lJ+B
O1jCCbNOilp7phrMhy4e5Kqbf19mDveprdOqN8xOMMwDVkKn/8gzwJUyyYKb0zCOd33izmh+hVE7
pjbYCHJEpmjCmYU/qj1mNcFByNsWp7jB/SNMRxUE8/0FcAQjAhXatTWfq6log5n+sAmTS5Zz/t7V
3P3PBEb7nAcsZqhjGLQoTn6qwVado1s5tnCG9F0LeDPg9FBasWu+m+AbO+xaKHTxtJqlFMVGcyvq
EY/nOhfGbZT6eBDPDXEloRHnjgjmGF+xo12OfSMo3Q7/RQmBdsfwp0ZCgC7mICWXwTGLu8XpIqpY
+bMmqGS0bzHfk1yd4TpDCNjs8N90C6Jcye6B5CxrYmD7ibyIy5DhnGRV+bnb0cD34RXuswJJ8DVu
vRUDQpEZ+5T4NNx1MA2QWk8N6Oie0293oDamGscVlW4HfftLTleuimRPCwu6b5beB1k2ZBIyVz/d
2woKV5J4h1FNauU77TLmHBm8UCa+wLFjlJMzVHGd1jehpxAhXlread9i4LBdunUuJ7W96Ps0mst+
jBRar54HgbnaMgyNfSUml9T+jDqbauhziY8RVtzfmOJxdWDYB9A8p6YFlelqrsgMj0k/Rp3RYcQJ
fITrxHEXEKOgTajAzZ8z0SwdGLkdpW3pUu5rhxzSSsUfjE7xWDJo0y3fjE/N4groip8j45ZHhJf7
j1XuwNRDkMHOFi9GyPi6r8fNfqK69y+wutiscJcfj/3cQ7PIG09fng4oMf0MetopB2W5VW6aUWhR
w9MVZHqv6dL/shagVv+6q08duw/WPBD80K9pGesAdFdyThzpBdVXwnUCTqNf/q59AiNJr2yFfEtX
dhAhw8Ogf3Ua+j3II70+b3kK2rxV8QjEOHkMCKCU3cageIcXYzeAAnxh2Qezri8teJARKp5+TNOV
dmA4tX+bmHHNrFFgRZISenWbktRUPExRrAAOGX0bHNKo+jB0l95oqE6hKFShwxQ81fROV++hmbac
NuSs1DncycpuqNUyR9ciDERIy4K3mUptjx1xTOjyBT0CIeChTYt4R9jiCur/uU7VN1jyNkV+AC9E
e3hTTSE6M+xI60CUOPqJ5K1LcYIabGnBIEPN97VZ1Qged+otAHlRs1bRXLocABO1og0plLIKN0cu
4i0sWrymKwkX4WFpf3hTopTkhOP3uSxyayKZrr47pFmzStPgnyrn289p3H6dBwudACvBZZ6AS7Zt
oyRGVDvq+tipczFS+3cM7FShDj3ggNzz0l7oxW/ndabsea/6BfJ5A9fmMKkHvcAPr6BnS9QTMjrZ
lqba2tv58DLc7W1sM3dh+DlZW42ZNJzsjqq+JqENaS6Z1xyN0U4JHqNpqmMh1mRmqx/ZvOT+gyCQ
58Wg3ifLjLwtV1bY56DP1DuDrOOAUO05vgBcQw0F69OV9xn+rdKQuXS27HoysyTvd/s6BzF+NHOI
VTru2tQF+wdwKJllkna+/KXOvaS2D9LYjxj1lWpZycUqIPRXMIlBa6QSbipSD4lpZLXc3Z9uwX2L
kdxFqnLNWdjjeOo4C34dBlo8oVZzH4K8vqT9wRpdioDuqi+IeTYmPxWuM550GXL+qY7ZaF06imNk
rUyd+kgex89/PpJbcP0GBSk5Ob3Anzh4OC1PYGZSo9cNyzuHstV1biKxYJGIOWwHq/wtZrYhPp8g
zc6eCIH4Tbv29+NVOdNcgg+yTvW1mpspIfZSR5Wr7/jOnvTdChesTw7CNnfXNPGPKEzlW72+C0be
sjWMZ3gV9JJgShirM8l07YwkD7XmU5gXCEVzYUjwtvSICKV+/YRdr1TrUcEy6q2NNUrUGY/83VW4
abFBFgMST7U9Yj0faspXe+DnUw0A27QCq5i4rQEDFuiwSGAXX3xbjoysI8p8zwQvVbh3UYsubkNF
4MU6rUHNPriqMWkbudD8SVrN0N5Vm0qT9i/57Wd7LNqpcZ/L8tBuGoJ0JubtA7vgGGKwYJ2KrCeG
7/YYdkFK8naji1H8rVU5mKrHrzJ+2EpDmPPxcPZ06Bq8EN5A6CWGpnG3V68xeKWQdw3phwC6smbD
9yqvARL52R9+Iy0wHwROqkew4lfN4qd6an9V0d9Od3zRJByt5YMl7N/aCAknhvciZbfEfSNVWucZ
G1eyO3bQH5I+ioO+kt6pxN3sAywSjxx2CxxykojQrlxBgl70+WULrYsovO2fm7WRwhfuPFAVVGW4
lpNEu7veW/VPFQbqanqpqzyp3D3hh2KQ9ZpjfuaXEmumdhuXw8yJ/fcy6uAKxF0zUv05WOepUXzl
3EyultOC2Bbg+tvdvD1EyyR4ysFnTnEPiaz2svr8qxGICgxvoeJyoiaD7kurjgXkw5V1Cfuq3+AQ
PGM31CHzg4rR5tDdwuENq13MqjmhwkUqMhRXRbk6QpypPxePLM19HMGbo3yrdgwgkWw2zngaUia9
Vvy1eolCUlx2k9Szlvcb0CtZBHIG0tgi9FshsNh4u6j5p9TBO6zKm8686fJCTczAhhIm48Q4i2Ee
2K+aKaZmVxHax6HEOTd6dq5UA8vp+MIktNpUkSPdvGnze2i35i3TCUcZMQOys10RhabEKjnH1C6f
vB3I84SPame55Nk+dOopzgDzRZw//QQgKgM77k0nY5QUGdJV6C1CN9r1uCyguJEBckMrLjLBDN1x
ciMl3Yi/nXVN4zdU56Wef8d3RYuC40zAW1JMDX9JgxRiEaWv7kImJU7DHas9Dy1Fdi++yfcVYCTs
2xOa0NWXfJZya06CLKOfjIQQRnCD8acnGAQy8345b8xbAQ39LvX2aInlLIhaW5isPyI7UN7Non5+
OF73KVbXE5+qN6emO5repTPTizUom1Qm2TCtixsuHcfgWZ2hvrd5PJ9P0JlirWMh6/gAZC7UVbBg
kfdHyG//yR5tnhxP3QQYDxds2DisK4L4ZHrKhtEkCXeRbps16mXkOaAe5jDKgxM8G9suLNSjdswq
bGbKgAZzaV/aQ6zf01KrHe4OcOv03UtycU2YukZEj8rZ6tG4/vm1PrcH4Hh0HLr6s6zXe1E8+OIW
ebiaPuF1Ok156j2Q822LoxwMld80NEsNFMAKkZ+vOCNliaV4Ygh2GgTzeTAHJRDlEcIdpj1+bkQd
2at4bN/5gJ5HySozA07nTpw1r/5YjREsRfvTdmyJoe0NuCkENfk8l03kJ3nlzaat4gjRvMsS+iB7
ahu6ZZGRl/kp6AEY6riNS6CJiBUUCk4nV+y/+IQqsRrfntoHAc8PgCOjtBJhxq3s/KNyD1RBf3AT
VsyOyF4nJ7xYI0HKoaaaZ0G8vAdNqnn7GZO8MBdlm93w8TtwgXOesUuYHRyl8N4lZ6tzOhMv1pVs
zNW5pFazjx6gUWqgODKxmmy3KomYwkZnb+hTHjRaEkyI/VUhSCqyLxAHM/1z47oesEv3J2Xvn9kU
+KiCqaGs92LbQdbfNl8jeZAQF5rv9WY6lne3BDcwwM6hGKAyQDJ9iTYTONP0rHs8m+q6Hb+VDdGy
QhkEdAb6OBKn3QLeBUGzpsrvvqj587e6lj5DSKEr3fdgwJe/Nb2P58CrfVirK6G6HJCTTq9tcv42
YybF3riTJCfwEanXy6kniPCqK1bxEAgaQ28h7zhob5F4PaWGEURNy5daHj7sqKEovcEEQT2EgB3p
Lb+idi+l/NLet7/pSea3dAHhrG24ZUM+/S58H2KGf+Dkb1VyZ7KmOC6MITki341b6XdFgMNuCova
geZd8oAP4WsmvUcod31XAVzWnPzCL67LeTbn9nrdLqQJEj/jkySdJOpu/S6EwTo77PDAbqMj5fmu
Csgy7gfLgTbKqWmM25hS+/DUBVDGmRxm9yYTGdxBc8TkzJor7XVxD/g105x199enbDiTs1kwBdSp
jKkSpKb++dNhiDeTH4b5mJBxBEuVbNzzAfg5fpKx2aCGrgVweAFpQXssmgNlTO/+eZJ+7qCYh+2j
+uKHXFpbGKGEBZ2k+xxFVeIXtSufOQwjZFWTO5V6fRdU8QQuGj9sQmgyhFu9sTtnIp9Wy4xwsXGn
9VEhT9SVIdCVNCD+5i/S0aDcwh3j++DB9aNpx0WnALwrjhooz/iCxRH0aHVxJAse0/5b8iuOwHUV
2eoIwU9FSfYOVTm3KIS/dBmWQMXgceJRoO/5VZXPHrSVYsXOyNbKhvI2olNp3EIAGmI5omApMAqY
RWqtAZJFOreCxUrdzV7n5zfH92V5aGFcqCXlVfH6gLFxCcef/46obdd7AX6BHR46f3dD823eTmMP
vHtOycsmV4wHCwBodXWlhciBRQswvbCnuqkLcp/0kYCXBdzVgOFjVzY03BYvthsHnMDCdPQDib3W
4FBPCNA5WLKkaQsNNAbjaShatsM09ePyybIUkVtatFfrzhaiXOaTw15ij8Tvli5E8Etzy8Ryzlje
A/SgjJO0/f4LNQmbLVLNrs8XcLw7Vs3wxsCX4e6IIM5vAYvHOm+p6fbMV3IWQeuEhSUV5z+WnWg6
zU4POSk4kmFr7xdzWGGFNLZgA9fwC9b1qrc6bUvlu0nuwWFavSdBuz2hvoEEPCqp+zrxx530vOHO
130j0u9cboXu1bxVkxi4sur3N4rQRJTy0hoAOYogWVSfazUhlCH89MOKSVLcuDHXxbcQmQ9c5VsE
CgInoRkdjvVMbB53dgKyMZrXGHUToK5UXHixmOV7gVbPxp/ECvNZ4kI3s5G3vLlQVkxj3R27MyeW
1u1GrPSTYC+uYEJAy0H0F3cUiYeYMpRLF6+5x8NJIDJgYyfovoieTw16P1ZkNClhEbxvj3JHXVZS
NVkQ2tdw3kNr1X23VRlLgcWqL03EZfSK0PkALBLuH7Bni0S5Td3StBTiLQDXgO8zb6k3jIv+3j64
afkAbE0q9lWnzFhNSgigID9tPu5r878Lm4sBxoCs+R7JPasa4j8KtzgOuBhm7BvUiMYwHzU+pVAD
6OjGCHLwFd453YGYTnkC0NRSCbeRWhxSYwRpRKIvgIM09GTS7/gQVmLZnZODkTkLV5qWemNAP3UJ
BUofBZNF1msl4bdbt6/BAKEfmvmUVQcJJULw7vz6YzWYNVP7gtnFLonSpEw7dXpvMWDyb5UGhRYa
zM7aTpO0F36JGlqKnCPUJ384enx6ezvpW6/+DoXIWNU6RQAPuJpvRcUN3R6b0CIezKzGQgi3/HKl
HeSLw30qhGSvibRITtUvaKAd/GFW9tw2yE6Q5WipCHSocBTiqPd3mPU1AGUTWbiPCMxhoDy3rDPs
DgsHOkHiAW5TchUfyULQzTQV6NptUV/JaKrifB8Wmd6UJd95JmciKtlvHsKz/P6iz3s8ERU51bAx
R3tHH/f5PF9ul52V8wcWrW6lZP+PdkemCXE85bRU1TOWWQN2velegadXLI/NSzJOT0S4wE8Bt9P9
ZGZj8U+ohPz0tyDR7ujIDOReiRD9qCAYkjV5Ci13pCRWaFrl6OsakJhctzxTkiVFVcytN8yD1Xo1
hBrP2B1NY2aBflaB58TgveftjtVbOUikZXKkPG7BGvZXYLF8sN1GfNbHPwBc7b7NU4m2/Ak4i2nA
D37WvwsZYds/dW/8+8pRssO/t6LlJHYx+JdubgJKsIR93/ULw5uQGUM/+PWR478+uChUB8/Fsybp
wGe8dNE8LAtZLgJXKrIyYhNCAtC1axxp8V/Leh1VPpt0h5bzd1XhRAxhwwNxZr+RuLHd4n1TFRk5
udgx+vksayBtamWVcrAvhRHJaxqNDSDu6ry+mam3PrRLPm6fl/1BuMwR8AzNDPtZNObTLffgOpRr
M+Ucxtuujni265QgkakqRD3mQh8pP1+dPyOruU3YqA+lwB+Hd/OyYwM8oSWmrhoNpE3wi9Eo6Vea
9+OMKGnyajFwVmsGoCCv1a+Uixc27HHwPk82vVK0bYgPOWvNWe8cngX1dDQXWcexoTivfp1qwFX2
O8yNNNZJsyMzhyEmrqH78Pj1gtbnwTXPLM274e3TzBYPA945GB9TlxEgKTHQeLxFWy7sXtCWcPpr
ibBK/zjAf5g1b1OZp5a3VFZJDmT+bbuR/hLWE4L5aWckfQADG/tUhcrCaH172k3u/xLkPFWqSCs3
W7jVfsxVD//5weED26giEYB+XvLMx5dLKAvht9p8QHEdWLEw95gxWEfgWGR3zXawOTVrFy8tk/Cx
wQYfrz66YGvCY/g01AbnAcPsLWV85hb4nSBeMjycJO96MMNKyaVyLCpFnbtyuRyMronMhzrlCbj7
l19zpxyI+XBlvpkz/C3EkChOGy6oK7v9BK2YWZ3r6zrM/Q1A8fQvXNl5rDiZfqnzVxcekZHu5JMN
z5HgmShDZDWyaKNWfmWr9ywMirzFKT6n8NgImzIUGWHfSHuRDo6We2kyuMTqTtrjPUESVC7AdlvK
n+v6JuiYWn/VdiEg+ckJiQrhoO5dPTBF6tAdjkbOCfacIZsJnTtANLhgNgjpT++8NQEj31W/9jOw
Gupxi6bie5i6AW8eq0oFOagXde9BV0osXP5v9GsVN6+wIEL4Pfjue39V1/xm6jAqmDzx/8DtI8uh
OD62AwTujwBcm94aNLXw39E2MxlNctZBXTxfoBdTyOmDUXlAO84zo/zohWq5bltviPFYl4D7/bA6
ct0Mh+YsVLESA/E1lZOENWUVlk51M2qsyDmqiFBFSlt1znkSFM/hjrOSmd8zDlHGfaoibDewJghR
jiKobc9Ykd9nLpsnQEYccJiQ3S0m12C1FtPBGVYo2Wov+KjRFJ1vvwP0kGfRjynHNjh/+wBC6UwV
P7K25h5SyOYTacws9p0CVDshwC5cW7064qVOQc8dzY7Tx6IOSl7FLl+E/53UYMmLJoZTNSSlhI5d
CMVE0jaaCwvvDXKhJrWGAc2f7JoDNExIiyH3A/U6DpkN4s6jMIcPlz2M2/tpQDQr9ERlZ+CnCoWf
wvfIszNtmsshIWZIaRc/kDrUET8cBRH8p3dGe6w4u54pCNtx8R14UZUn9ulrW35U9xRHbtoQx+0F
FOgH685NFZhgBDqzwdwcyLu2qNJ0qVwesSCasKKHZ83EZlX+0bWeZj/FMOTzz/Drer4zeghdXNZr
+uULPtHFaB2M2jue2ga2YPBkNwsFq4W1+R5o7Ju5IAsYrzHGp5oqBvR5LWYBLRtazzYEyIn1/8bc
nbds72efaHE2ujxguTIlORXH/cGkeosKCR14P6FkmyIH/zm1tymsUUJN5exrp4g+bM0Q8amazMF6
HTr8PjOSb5qiovaHUhW28z5RyHCm46HwH/fpmqZfZ+I3oAcJA+qx3p4njERIX/1KpRiy02MtMq7p
0DYMvhSgBSDIp9z1RBCxgV180/amzLthFTbAuIJJN4hZTO9lInnqvYaWRKbKGTxLHLvANwG2KCkF
QBlteKyA3s7XUr7qYU26/eF2o9UOxNpl3oZfrafdbpDS5Na2y82qOdMYU0Fz/pE7HWepMFXofAu6
x2xzkVp8GTbJjc6reKHFAFbqzjCd95Ze97+hO3m1/XEv+IeCBNnLWVCYA6Qfq1RVHvFI3feT3vTi
CedYAqgYjlo6aU/ZnbzN0y24jnG2lm6E4jKw7xZqP2Vy5CFTF09bDVRGioPkqZticD9symF+VqN5
3y7/Q/DyXbC8hDDUBsmjNEasfzMai/ZQ3NM1mBnGbYp1QEK6MBi55XtWRaZTxY8gV+23HYG9m5Lb
jg2ggHUbK3I1SOtlNsrnyVdN/FQDoYr686emuRebxkyZDq8IU7t6iqFnAYavZtTNcTuveInBSto4
CeVr5um5WJ+B1Xw2klcCyDVFRQfrAEphEKEMD0dKb8s2VDXWdHs5eHrOL90rKLjFx1nsRElAovWW
G8CPz53edYS1G5LBoAsGDQ8nLkLaKt9ljqba7X3KfQlvSkHoTK2xXn8EcVDhy9UrhySKGQfAipAK
WJlDibc/WeyRXv84PLqT2WS2fakjM2jLss+YWt52rHT485BRFqw2LaR+QmxUH95CiO+DeI0GqHm2
fAQSa9RuUaT9wLsZ4esNag9N7jo1IbPSdF4/ExiWZ0PtW0/9xesX3Out18iZo0bnJggFP9m48nWi
8EI7tecZjeVlAmjiYaCZ3jo2Rmf8T2C0nHvpK5N6V+Iy3Um4yPLGQko5qt9tXjIsYdu1RsN1R+7I
JSbKmSLaeYbmYcRtO5f5KnV9rF35dezKT0nmWPTEUI0aNDHtNym02Iv6iJtk46vSSFuK+L17m9TN
giKSUB4xxScFxVuwBldWHrP0T4YdRITUa17Jc6jHtW2EOqROIkLnpA1aBFVax0UnxMy8pfYQjphV
3XJEZFNut43WRcQGobm3qm3fjl8JtG8sIriv6pHSMoc2kcU7RYH8BJfKqUJgTAzoB0UgNs1RErB8
7/wdko3yQiELABaKYx2AtBs1X4vfIMg3+/Bi15vxRHLWpGKzreUSm3dFAh+svyechCMZFzLeFqYW
2SpLzjp3SAwpbMOWZ75kbWIk7z0ouLHJgGEZK4L54aYAaHnzIJur7t4mRo11s36XLtYJuBoYL5P1
7SWIumiqW5JnrxDG5d+dShVxoaVvaAz0Xs7JWet2HSUvQvRSW4WPW/JppeJ/p7Mi36mm1dW6lV7f
rkGEh3eNzbMLOtEeJ/4zIetLtOSuBIc7xBNdSdeeHZzeryfhYnQijtqYuUYM13b1TOikWhecWyJw
OTzL64ZAfhM0pTcOoJQF4t+epoAS6M3JP7PrPmgY2neop+URF1ScxkBZiQ3Qxz4tIY+aTsFo5On5
Bq3AekemP9A6MEheFo6J4wVLcQSdifn+rp32iiWyc7wASCzh/bao7JDnVg98Tdxy8ZJAszbpv5jK
Qa2OJ4VEqoZ9tcS+ys7u3/GocIsFUtbznL7oD6Rup/i+0El06mUcFnliT+0jU0YHYoABCgsDMBjB
5ddh/RsEZKLufPcP1QUcwki4r2J0GIDWtE9xwu49clxT3f4lT2o36kZ9VlXquX4nHCb6LEGssxFQ
YcLmbFEK+1wmyFAZkmJy56X28f5YiJ5unPFA08vr7H1CqxUrikAKJzMI+OEMnT7LG7nOhRE8+kIN
TdAndP/y6H4s31/jNKCXedKItWWHION9VRlQBZdSPB3oiTA/2UkqX/lGFRmcVtRBSiociHbJ05jS
dpYuyEIG834gLlWhda0mTUQbVsXz4Kow4TmJ+gCICQSriEPhpVKPlxdIU5Nmi3ETc+c7ILQjsMKj
ufzAIJ2LdemOMLkU5MbL341K2Dx2GAca6ersWLu13Bdxdv6T8Y6UR2KS8wOJ3yBk5Hp5LxKCgca2
VDmvQudLYIaHCMFY+3QSYeXJ14djG0iChJ+luFWLT7VDygzgBD4pl/fgfIf14w5FOsauXY1GezZn
092En8Tv2RxMnNCdcrGiBdRFKJcl6oZK4dUC1mlHPCUlZ2IlmpKbTI8ZtmXe3yngTS08X2Mr0ye/
nJ49ls/T55IVTNxLxVn+eYkGVmV1MJF7836bQRRfz+OK8fwIvV6Xftb1i7epixQPiguWj+I0TYOd
yzgXtnuaVmvFsJkzSDh5CA/Pqa1/OuvANhzv5ctgWHmcU1uN77YZqvlWGwV8lS/syhKWtorsEIuu
e16/HNrqt0p+FUnfarbaew7PM2QUdOotgIAVKhiyicyiwgZu4eSBXu4ru0TR0wBLdSedNrqFXWLv
kQFEXqLSo1tdxJh9jnJzgXi4SEgDc+OlriAw0Udefr2zMuO1Dup3yvQ538SXxhsqqZd61wjymtjj
x9AoevTpagcw6XQOStVYuhhy3LcHtvxld/6b4qHpC+x6FInZqnCivboGglVKI7mB/kR5WjqXWOve
Kur3Qgz6d31VhjN/REo0lqS2K6x17peQsKuNj9E6KAyQlcT4qBK2PCeO1ddaMudSWshQzjd06jTW
6xf798egeZisp3Gf5wmOjAFZMmev2pdgxbgGO/oUJSQNKCPnTjmMpndNS2y1wu5Ct0bO2K2LZbmB
q86AtBnKobw1HWuIGnKfJmAy/Ax9os0nUtHBYXSDetlTZtjTBj5EkIuFT49XoGkznbOzLlvh4YOd
RYetgsWTX3zD7+Jnlf3FztsHd3jM9w1tXqWeiYqT+os/NC+JScHarJddCoaTZQQaCciX7stAqoZG
YT+L0wt4RRewlu88iZ+msZyNQjx2YM3l1rurpceMyQ7DBWfdhG8E/NzgabRUBOV0+iY4U73gDRBT
/WexSQWNxVo9Kk9B9ROeUX663Q47xyWnLy/V7XIrq6Wi8vH15gxD20uJ8/Wio+B5hMrJpYor0YS3
BrLgUsgRuN64ibWXyxugxlgg+2VVz9kqDP0YkbRBjpJRyJnaJJXR7yd1rIksDeTA+w+jpjffdQCz
kTTZ5dI2M9mnEYPPbRjzaXg+M/urKBufCUO3Xckg0jSqC2QTyyhae6mYZCjP+mUhKxb7mC6HwEWn
AKlAsjoIgAomdbifJCwjcskK6EbGzzJInhYSgFZ6HfaTPkv+eQgFwIM+KNsYJGDJylRMT9vFp3/q
zKvRotWBODTH3UT0P8BW75N85kdYi5AlMS+41p7UwAasCuY6oKoHPsVcLEopIsXR6bdzYDnknQKZ
JOg8V5Kci9org4C5eVPH4rtUcFaOY8xKk1e5E0F/ICHtUMqvuPH/tuKqlWfRKgCLFWm8IUxPRspO
SZDDGuBtQ2IrOF9A0K9ifJyZFkCyq+JRw4XLy0QB4XX66Rai/ou9Tce6HujXug6dcFj/NGJzYXCP
6BhQxrBVWyhIHJBmBeJFz+JOQoBFWw0NUddi47x8G+fuNIDyNAaYpBKwltBvTZTUByF/pK9yyXk4
Z5R3mgO+qvkCFRmza7qIHwYtJo8+BjMzvhzpNa3F9AsvJ+m6kRuXhf1XvwOOstHfUH7ovNdUp6Hz
Sh5tKpdJ55DHBXcyzyx20t+goJne93gmZ687x4XaDNvaBax6K5kVA9wNmkNyswTTOJvrO14+BJLB
61RFzG6piZWNkz9TSB624qV4hc0LwcfA0zbC6PUYCGbmdQmSRigl7cAHKviPnDqSta/Ooq+LPKeB
7NAb2JSqjllS0Dztds5Oj9lXBSqU+PA6fiGtaUzo2NG/Zql6L3jFg2Rdy27AtIPuqA3+o+qh3NUk
MLJY6z8tkfD5RKhqMmL1a25k+D/3E4IL7SC6XtxKc7Jfp3hZRP9dNvr238RDN7mB0BEsu1kOa3Rx
Z3UkR4PWYXpKeBGf2ws+OIoCJaBJ9H6lZ08cRJg1FkW4LLdPWCybXdKuGNeBK7ipu7bfT2SDnaqO
8dR+B6G0TE3OZ2Qx0/ax8/s8NPo9HZVEA9IfSPLiE4ljqFI7OBFttIPKjUk5an+WWNwQPE7Nd1L7
tkRHaLtQY6l+qxM2tccfHq+Rg8VNlrES2ue6yjbCCIPmRNzVnR9Pbnq4qi1XCT29NkBY1wKBsrUu
euR45oxXpcLZ2trRUS+TLPN4lECAVf3dSlJ4cVZpnBJc6Y/tdBDsNucu9tG+ALcvEiOkTa5P4fwL
SzWRLaxcD60xBEHnTebRXS3LcWcswG3u3P0d2YR/DkL8wuJsaWtWz2p+8/QGSlqDJ5Kb4q72N9Tl
IfDJCadlKqoY4mMoVoAgH3RSX338qhcmQRdTAnE5fEgO7t4nazoLlff3zSDwWHKsTpawFxPmTqE4
8L1uH6VLnKgHemjcw2WBNLrCACrEYauwh2VFHHNM6o15s/9vgVZwmG8gDgDpe0bT/Y9I/sXQ/F8a
tsRcvQjQyEGWZlRQjeZJIWkzlzwLBKx1jJknhSC7cF/PYIQRWe2t1JJgTdmilJOHWwAZviA1qcY3
RW74ca0sQzRzG2yISN8ydfRf0GG6AhjljTSLnsMZIoXtEK6fXGItzcKO79/CvDt9yKd+Nk1RE9DN
87h1hN571MHbFN7TIeVZnAXRRI7kb6MJhuIt58hNzygyr0QMykp8NuE8/RqgmnaSaRWXN7yYVacZ
plkZg7dL3MCpqwdx2qbItyf3gfw1PcZ1Q9U1B7uZVIt/JeRtxfdixHV3I0MfKbXbAhtHLEKb64hB
nYxWle81ZQDlliFA0T64CwjPrXGelYWCDd45csrHD6bNGsKqQ+dQliZwF9xN470kT+OuQLVvZvDa
Hc5kE4Uu3EpLsgyLR/8YDKaBHnTKfeN5K2A67L6olsj7BbiSFk1Iod2MIkO1I/szymBRTPECbY9l
LxPuQCfpJ79gvlf6TQ7d3jy/3EiSDAoOi7j7ZWIijU/ehl6xjJ8lWAFqoTujRsTWMKXlQv7G/MD4
IlhuUIvuuNi2tyr/ub6BgaKjSVY3mcmCIsHy25J0QWhbyg06N0q0Bo/robSaEIP0NB5wDtM4tuky
GWWoI2RiJi4sRY0gdFF/GoLDWO/EW7rwJPN+WL9GaGEIm+rAop/mMgywnD+XlUm3NbyiP4gBzAmb
+SgAEzHeU52oGxFXRQaJNg2KTkGBlKlJgUGpNaepcM2vyJRrVaS6D12aNflFQ1ZC7YjxMXDPRAqw
dVQi8/yO/Wb2svnNl783aAuEz/2Ez/cg+gehbC5OgLqmj2VYiFDJM6WSQ4N2ph75FOypSMLBC7dz
mh2lT6gdNzs3efM2oXGR/fpwoQ5U0IrZBTgjrAIpMCdnDJAtW1z2TMsjZLDkwlTCFKfrqSOt6JZ0
VuLbTGr2xHXTynTCdkS3ktnm/+zG3Ckvx5dVrVbnCCgDhe4FQSFkb4l/eqj77Kf6PfLJF9HCUv3g
MQa1Kv/V6Oslu5JZPUpA5L2NYvtsyd7BZHlS3QT8fObgCvZKpEFgDyO0ovn/Mxn2+iHA0WOvdk6k
e/Dtf0NUZYNaUfdVAs//683N7OvujAiaFzd3VSmDZ57eF6ErXpct63RyJahB2DPe5HSQMgqi+RVy
sI9iT0fQlSIfwZk0rmDlfkNeBJUja7otMu6InzhjMgVUoBmk9L/UKw50Ff8X+lhR3d1F30EvEZo5
TYM1WeuZIdDVwSDa/du4aP50jYlNnUkvHteNF9QAFEaLrrvvi733VLqOrr7C4X0+qWhO9XzHRVbG
fLVp00SNlMt5H8jViy6rt5QEDhXK+gvDWI377ZZzEQkj9Fg2emh02DxAWDb+w/JqUHnbDoO+llzx
L02RI5ugjAfjPzGaYx8wm0stFh92BgK4/fxvYTpLlzFtN2NPjBoUnsGolPWIecq7HYN/IiRjsp9m
6lH3CQcyf/3DNKCkiMdzqZ5koRg6A4tzSF6jyxgAn1YHmYQrIFGfxLx1paM3gzP5DmHiwzRRkSZ8
W1D0iiDdqQ4BmK/q+r0lkx0d3WCj0d7/rn702m0Zlky4Z+2cx8R6H+fgXlFvQ1vRZqybT4pcQng8
wZBGEeriEzjNuJGrGndt5WEb7Oti2u4z7dJ/Q+NsGel2tjTa/msEGkrwk4w7oc/rD/VS/+4roBRJ
OHeBOFOKj2Tzn7678YMAURg0vh33vhrgabBXNMgswKEVVO06gO0k07XaKgSTdg55aE/l8aT+jiML
FLzKyjLsNXc97xrcvY3eqT6gZGD815FBMLS0V8+GdYC/kc4ZJ+coHJOtsW/f/yrHazLW9i935pph
bCEbbhIakY2V4QgaOjFV8bdMPVrf4dXXE9y57NYAtGBHUIt9NzfTrP5vZLbo2Mf31is+rOo9RZrz
ADiavtGC+TWwt34JHFcZiHx9pirjgseAZjy4J+RJ8mpXcrID6PTGVOnmQaLW7PHcd8Cyy2opqLZ2
iQysuppJED9NZXXZv9Z1mV2u2+6K+WvVeVo66XcV2pZe5E9ySmhKqOeAZjpNn9sPUqIgzeKM0n5P
kHbbEGhUChgWPTwijQ/aku7YbklzpC8oCkUrOJ6e2hTlRCQS+IZujYydaC29/NOvt0qnpm0YU9xg
KIOmDoGnPxOzzY/AMcGdN+YTgen5nrIK5cX/A3/OyDUzBpXNQwQJhNxFExjvE+5y3CB6g2mgRBLY
vjU2/Ms7MB2p2qgz0wfREoDC0KqZEfcsIfegVngjTsmBaA0qQgyopkpgmLaP0K/TETAt/KvG7MtP
H/+RQg5V1HCc9FyinYxBQmHbxx6qfsksIOVqHFvd3B0r6ueIdXtrBQ5DxiZSyQuXO+HtAOuLAGUR
4Lcci4LCs2TLydXaXWwhG+rKNIw0C/xZLc0d866xnlqaePYw/ohcPCGFNO2JLhgKqnjDrXeNZSzM
VaJrlCHDhVHNaJF8qeShsiKdDkrKWcVAtgh8FbRN/6nhmWm9vnnu0w9+tUlKwotvj5n9v4cKkvdP
Ky9sUvHLksp5qWyW7MEpHexHSA+HgcC73P8gGUs9der2sEQCWH9N6ck9VKLQq6ZrMCqURuiyO66X
JhjXXLP6HK7RNjWEGDGFpkj8poQbjvh27MhHNFdUhs+/XhzgVS1atmuqYHA5WEvb5Oc35Bf02FH7
ajO1d8oArcbvmf9VxARHouUt0RpSgAgkr/FnIwY+dX1Ahuh+TzUoqaOd6rBUh3xeQiQdq24enRrA
Krov5fPeHplZUWcfkABdtw1JCWnjDp8PF7TS+FMOR9WmpmB58NAbdy8wjhS4l0vEp7K/a+0k4T0H
WpShnmq2/jrHgYXIjUQbbW9BPQTM7i6RSesZDpDvIOptarC2ri37A+cLdtmF9QDQ66Ab1ljXEvBf
vYtNDnv3gVnoIrghYB87ABQHb6SKLIbU0wf8QS0rfKNF/dQmnfWrvJ8HDpAYgpZi+KMFa1h1V8Jl
4dncVJ86GOF74rCij560AHpX0DIf5gAKWiTQBvyjQOwI6jN58mrpCvsTL6B+pNjv/UhxHrgBz5nV
E1to/tyBaqqxKZGw5XNJWLs86TZmej03bH4Jzpab4qLFeVKjWo0vdoY1CZqvtoHHrkhr8l4Si/O7
OQGkdT1LZwifRp03+k+alNQZzbwMZdGR0jVbRN1Ir21XuAuKYowaH38lo7U0Ik5L8FkrrEiynU8W
lj1FONhajol0l4hFXbHe1iV+nIJ78QqWyqPgpmwdX9Xxc7QDMaQs2YHnQ9L53dQt3kyW7w1G/HNQ
SYflhtjHJ3eju2ueLqNTqbJLc5OHqRXqP7QnSeUUkseGJjJpJ/DjlZuWGUIpUHUPNTMKx2urwUBz
SHaQKf1tclhcwmu4Gg0EH2Lwc5EwDA29Pno/zhbJrAtAWyVSvOW5CHhVmS5ykqn3PywuHXtzC3+7
wNrwnqfVPvMEHRluVRyCAsxyEXc5wkYofhZG7UcQQ6MmM9FKOtgfmhyEPIKwRaBBzXKDvlhTEXDc
GgRKW8TWueqVOWxXgOcrJ+5RG1d0sjwUENFa2tDR03d2Wk44U5Cto2XnmAt5LfMipwGJrPo6XEkD
9qcOaBaR/sXzNiGNFatik0tjhbElDCjkbOT2u6eTsWr9PHvl13iY27L3usq0ZO+SE7hbAZ2kCoqg
+vkL/PJGd4p+TztrD7RnDtdKN7ZaiJaKJvCvMr5yNja9gH5wJoK+6toBghpNiM8lioDjjhXg4oEp
lF8XjWFbzsgPr0cf9YGQFo0ShUQYifZoBJFT5JMYqbVZMIw9Rd/dgfiCUstnpgj/weLZ2U5xuBAF
2/rnf/ldAV3tKyhMV6xFqwgNaLfpEyH/x62CcbiO9PdEwkjYDgTEk/DqPv2V3YP2SXwRZ87donVW
47NK+9+yCUVC3UOlB+jPDxQ8JyYU5iD76Ozftz/XOhrVIbqWfxyH4FwpuarpFzjmE2jR1E2NaAXQ
S9AwGHkTLG5YvawQwfaCrLCFiUGWNI/rTgsvlGQxaJAki33sT6ABtSnGxf+z4HYMFCoEPO0yeNGt
oEI0hipOu/WISTWEY5cpv9hIrGb2mOQ+ZVVT9Ey8yNUp4DTv8fFc8UkPh2yMh/jUCSwvnpeS6zrS
HkHUV9H9q1HpS8X43yc6Upb690TRR4FsWFT3KrBQl3ZTCNNHvS3uP59Sv7Z8th7pTz6/CJobEN+E
1u8GKzXzhtg7VtikFoF7GOjaHIRtxypgS7Tn4TmLBxReqEcf9h9xUxyC6HqfYt9P/op4Ef7xF22r
Ng6SnlcDg61lkA2J5shKvqX9nYrGs6xjgder9A4uIcLzskIQJED2tPYASBPRTuPkM7GrfCFLajpo
GiFvPTLJseHnZ2FGU+gw99I7Mmtw609FYquL/mlDd7BqrB4025wub0C+iAbIWVD8GosTwhZ9MJut
E9UkXFIUuIct8a8mIPaCasecVqxOomM1ymOowDLn5dr6fWQrQA5ZQGclKjrr9FkTbTe9FOqwzrTB
I+KvjfsoEE5s0JoDwWgoExukTtYGGTcre7CnT+qzkwVdFb+rRtFQP9O3c2b82XeW0NM0l9kmHJ+m
As993R6AyGag+v527CvPJlyZQ76o/y3yS2Ofyi1M9HL0uJKbcPWGnj3oc7ISgqvi2GSUyOhsz0LC
sp9wVHiCXqzzdX/Bjf2L8trZr5czGXYH/9Art+tz02QL5sa23upHCT8K/hOpQZEusC6M7GC+U/1J
ml9fcMQ/ANkUQ0I/c/9vL1SCioVlfOLIdwdFpniF83LLBO8WXzwfsLqRfCfVyMPkzk7P6D6mmOyy
9qGULxpyAzcEUZ8UdeJX8GH+r1jS1PwE9TP6UsDFmIAojDaJkp9wLtEJFNcxCOnSsCD8jaeBiXzs
hMFuNYyUHYk5Afh0e+Qd64+XtsiyVoVoruhrIzacTU0Q7N9IS5uBq9DsmZXlEOdMth9A02RvaWqW
RGL2gt8bawOL+XuxtEkd+91yj2q4PGFDgJ7ik7rsPqpiEp+Be1PPbYL4Dq7/qal4mIoz918dv09g
csplvOvzBzYrEIreettKFDeesuol17SOtecdzFxwC1J7fEhI6bRdrgXd4AhoadtDwMfbAI2FGWNL
j75ry2aJDErZU4cnnjJYPfXfuzLPEr2kl3NQlQq+Sipon2QtU+XRA0oDcOgKJ+TMSiFJV3VqHvHb
RE5fFipcyDBtw9FDWgnkDuFJU0ZUhvUHOs4G4yMf4/a/A0Td+wc1cKJl6a2ICD9vABelJgBbtL+t
8I8NBvkeZzLyWI2IYiFNJMoMw8xaHImWcSDNn9g/0qWIK0oXsYV3yqVmNyOFYz7yd/DcUGxL1LK9
76+EQZ7owOBTpyxO9QzFxATDqM99236qGVuiczAUyJlFy1+/jORx+c3811nwFKbRRjTx8r9WdtX6
on+DgnnT2oPrsMMnBloORsLmsN7yIX91xuBh2Rc9mDD/3rii7WuW/NHBlVLKW+J7z0vuyedkPshB
7OzazcdPdtv5qCivC970lG0FZiVEe7QwOnJGJoBzgcv62dRSEx39pcYouDJO1IQ0POTRE4rYTVDa
fVCJU9IfoCRVhjbzfjeNwGvdQH8oMzvTxxBv/4fV9ICt2DUU+uIgHVGj1Ex7VWTwpvymcHq6IQ9S
ORJpjC/CHXfOSEMvEZkbXbgmASbziezcfhAf5loEfM1Y4B1aB0Aw6VQl2F6u76g2QkzZ3869NzP5
bpaCFpl3B+cEChB80ZcSemWBEO/KcHKADQat17LqtTC+7vvi6SVn1sD6AeERkb9PWks/8RA8SVFG
oYRp/X8IYa8FyHkeU3zplPuH8hi9ILYs1e+HFH2L2ufgH6HdG0Qud+Xi4Mm4PIU0jinC404bOeiN
ND8PNCJxAEryuD4nmPUuDnLL3koZ4qWApElMvvhU4ej5PLFr6C5TFr3Y5aPuyoo72K7S6PA3gWIe
9GF5pBTH8n27TeNzSClSgdz6Zo4fzpUVq0I/geT9sPXBXMI1fDsWf9fEW3tUXwYmHxpYxpmmABpW
Rk6PLwnytAn9ZEurZN289nw11kQ1zqjbnHRQpdMujwgmXxUjq5pEcdOjfU1vaqAQMYpC9bT1fKrs
ZHI/ITpKivR+HyYNcPPOGHaj1kS8Ncoru+yodX1LCb99VksFlADmMr+WKTZT/WiyWCA1Shtqqsbh
i1c+RjzJRmDlwPVEe/8BvvSCjGewN4BUQBKSkl23Zr5RvSRRoPImB6rd+h8PtKDDhACwGGnBW/Ca
NdwDPLBFY2dJ7N+GbogxRND+Gy6KLIWx5Qq4zx0jq360GxKbYSD19cWPXuZ7lWouKlFz+7gspMOA
qg1jc5Qv6rqRp+grUqnbic5HIckcEhfPwZjy8F6OvJMXDPd0Ya6WwPPeqahaOEdcP6smq3Zsss6g
0kAnv/pPNcXyBht43yraAgMHHjztT+Hip4HVy2KBYQU0nISDiB5a3iKvvQVKkCH30k7AwRgpOgeh
eVTO7fxkqbgZlTuBQyfXYWvvH7aO52YIAM0MxP1LUFBBSVgqNd6A9waZXaB43bfkxh/uHRocxcxg
M7PF9arpYiDp/FD3CGZ5Mf8sIrX4wF0Epzj7Rh0b/Xy1DIp9U6c2WuXwAvNO583O7OFswVvk0iqC
nKW34+BKWCS/sxIOzJAYfg71hiDXBpomI9SorJB3rRzM63vldOf/c4Cpnlg4sn/SdDoOyS8snGYE
Ju3Yve7ryD9dR+3eHXCqUw4ObfqGnuOJxzAql9n/S1DNX+7Ohl23MjOctfP9H+ZZg1mrxTLfqoxN
Ulm5cWCodGyYDIpf4qKxFielFO/kSKcfwyOcUSuQhFjQd0OixdJRDkOx2zbZWB3g+0HK0ECUh5c0
qEYg+HCReEqpBcJCE5+vLejZrrqC/qrc9RHqQaj+Fa2bATdw4H1MQZyeySuxF4JtUMUfLkcWvdcY
FJ0dazapualGWg8p63pe2i/LseQKmQcNxt9Lq76rzuije8RDo34xhHLDbcYq9gd6523xAydz25Gi
V5ZqKgeoBKXjZQEkyEpF8D3im4uzRVBSmWOrmZ99wrgje3xHXeIzgyeNH2gYpnix5Uq5g4ThvTPe
Mo3IW2j7QRAM3b6d+F7964u7WVO6gxkXbAE3HJG9emlLKy1E3qQDy4LjTKWhfUA7/ciBzeheaheF
WzknD5QVVJ9doAcf9aRc1JwbW5wdPCCt9hRDpiuKshM18RT9Tf3Bj/mTc8SutsGCDg1PQTLtWraX
lzVVMUn7FyP5p+zspT8KpOxB6M9Z5qwlivNdGHCle800YL+hTfTq9ExN+Y7HyOKovQYyAfVyIpeh
KEqv6PY8NBtyXclVUqihi9JF+LJxx2MmMbw1NCBKrtM6zoNMLHp6b9QtPOVZUtHM7I7zFT8piXXx
lo3BShQv8iwggMbFHrmP2e0O66R3N/zs8qJ+gHJGb0uZpLawIgzrpUqDia8lkppXiZDsQmEKu+zQ
DacGp5C7zpOeVotoZJfZtrQmzGu/YciTaQfPieSi5Kqk0HEEJglK5meAiH/4b3bC4S03/LiEeZb5
rRoNFVTMRcfzyHY7Ao2j9/APP3IL6gmGu0tPv1Vs9fxOn1yX7t5oR8N2/8frj6DhZauErjVUsgVw
xtBDM5e8e8j1E7Yw3D30xxswl3cjX8rir6cJviw0Lm+4zesLd8ES52SknRb7Bi1puXZFdUCX8VJy
MS5ZM+b46LkoSyQt2wKWZ59swB/BDqV+3n4L4JUwllfG6ForZ7XKeL131FKHUor2Cc4eeC/9tENa
4O/aJah47W/en8l925sGVJXlys5WLy8wchTXFi54FZ/s9tEQvzz8/y9DwgsXOA4mse/IXRF3N1Ar
bsbAPWzgO9uRITYhT4Xe2Xgcatp4tJLw4vyONdVxAmiD9qr69dfWfOT46uKAp+i77xBiyMfuKnSv
xPevkyrmdAtDQ0lnMt8N2gxk6zXI2CS1rLBVyg73mBRMdiWq25uX9RepaaNoPU6WbK6jcC+t1pqG
RcgOPSMhs9hxk8a4gqxgXOJbN11sihptug9zeLUX3BThifNj2oeTYMfJPa1NF9UtYYpGilRXTzfL
Isrht1kDXMgaFpdIT8Pv+lbw2sk3vEuENKlLm64kS3w/2lIctIxUBs2SqvpkYbekLGYFrrPTecip
bplkioj3m2wCDoyHLVqb2+UdADuYX2iRZ3PJGlqImXe40QTiw3GGI/lVob+y76nnRRI8UHCn/aiB
P9utHgP3GMCKNXu3zkoRoWzWrLmx329cNMLzhFLsM1RjMaxtmVtwsMU1JzuYjzkh+t//HuBo6S/H
BmqrrdkzzZwuTkfOkeCB1Sga53abLGVgqE82KxADbI1yf1NMRyIRheLflsIlvipo/DQoOLI+/xMA
5hQvLXbOx8ZmmgCs+3IoynuTGSq5vX+1+rh++uyFjVWNcGrdt5NVeOnCZBGU0KCc1jM0A0R68NzI
E0pFZuUvlonviggrDwgtpnaTmct8D4wEXrK2Ev0XTtdZtKorw1b9MB1cN89i6MJ4oqWEUsAyXJdz
6w0WGdyjQUG5wZTor0HeBx2AsDc+mZEvH5X9UzZwHKd6OKxgCV7JlueOw/Mtu8oTEQ34nXrgQyyy
MJIZG8PkQ+OqA22ywxFQo1rUubU4x5Nmweqec4n5RiYFenRSWRmWXfrtK6XzDA5Hv/2yjsZ7VCXM
HMp0jqCT+dITNQQhSw65E9o1TNz0oM6/5ueJIvXXbS5PNdbWYhoh+T37A4bVu0Y6MGXTK7hN08D0
3Z0cyNHctKfAj//KK53XpefzdPOctfHnbYSbQQcwcNN74CpkKqRTizF695Eo90+jzYGYzwNyH8oi
znI79pqT59v1AY4SmQJ9Iw8DNDJvH1QT5hgsd1pOPz2r7SyvX3HKesk5EB2tS6d9WlMyMaQRvSim
x2e1utB0oC4xXwk1Y7jjBJXLqy2VQuEXzgG8bUx90x4SwBb5Q2oWR26SeyNjVmtDk+c9nz8QjWW2
YAzVh6vnYGcGmJfmNhsgCKll+QzDz1/N3L3+x1nh7MbFxLQMu+Zzf2VbDceRvy/jSYY0Yv23Wfsy
sZR927fXJ33P3AcbXvk5nPbuH5Bc2iiNGebkrUAjJE+N5yPq9MaEVqAJCFLjp45sIf22b0WsBRbn
BG+B1O1luwRFvEAtufMcrWpDe0KwG1kkWm+ZgmfzF9G6QfKelwrqmnmnS0lwy7uY21QX+JwfzN9A
uLqByzggOTdN53UF5SIrfNsFju0vv6xiv6H6+9Ku0cL25o/UAgk2qOiPF+v4WoCrGNZoElQfnPJ1
5Z1Qt66cbxCG+o2KstUxACRoMKhwMslKQ1ZqIXvmDWndmJQqP+lKyGVvnXLUXGRS3xRnMqJUcOed
fFiIZmeJyxLL8+VxYVDuRYrhFqVa0JU57XPBsQem9ab0WyBv5CPHMp/1EBOTMZTXeNtn5o6Yj2cd
XYggYGwb7A2OpVRD3pZIcyE4LouP4rIe9gsAkTzWKgGHn0RLePZoe6f0wtDq/0velgUH4F2imJYy
f0RP9LR7WQdjXnYu+q5MxS+NgkrCO28t+eEXrTCv2YhoJyf3NtWAD9OdDxjj4tXHafJDfk9g05HF
iyHOksN6WhUlnCRYwYIZFTc2It1dU1wdttAFx/+fak+ITxfbxq+OvywNMZDLsUgbrv2Os1Xj3rjb
QnS+q6WI7mT9vQYBe+J68y7puW2gA33OmL/Mnj6S5vMlS/EKVThQo0T0T/I3XJkG+7+I5gozlJOx
jpGC0m/fl1+87DVa3CrOC+pEUDZHOZjp4yNRA0bPciQxmJ+32cGVRBifK8SkRiKxtmeZpj+MLT/q
9wJejPQadBuhpTRLgGPc+lk4amXDPnIAV9FNRkJFZmFGV+NTiq4miCvZDADBZfKEtUj3bT6nQ+F9
TynEfpTXX2lx62nVJtebQnTMblnE2RnEVtoxML8cOG7viks7dDMQsDtMVgZDFjSUP6j78fKcPS30
N6APWnLx7qMV5Mbb6C8h4nXQIjI5Bxap22HYAP0BFQP1jp2IgZul8MYdgkxyLSUeyGsG3dRFomie
qGaAO366FgWzKJxFvvFEyQVg2tN5p5ZeNYEoUiaH8GySlQO4IOtDMNNNDjQXkTP/xXg5g9tCveYF
W4mMjiqC3kdKApEDUdz7wIw8gmpP0dFpcNZHlP6WYIIjfp5k7TBxh61mAY31/nu2i1rZlGkrNgRP
eBcQ1Ft188gpF9RhTeaNHSk8A3JzF7Kq+tMIeKr+EKC4Rz2nJkY0PQZjhn9/spUExmA84YC67hSZ
htYHcEz3cW5SbaeYHjeMfnQiRC9BtGYU3NDP2p4zNhmVpltOroPOUbaJ+gEx8cWq12R7b4j1IhZm
bAUyiJBowXa9VYmgCElVppk6sOwdlFhLB/ulm4uwEZ/p7r83pwn2dIo/nCh0NcHrPT1u+NSV9xo5
GLzgrvibmIDTvL0RVoWheZ/qp+Rl7gl5oFnDUIYTG9Cv/nrAREzfYPBK9kTO3O9o09lQ+Fkd6Zv5
yAzN9qJefwEa9Z6v+jC0f2IWXJDAisE/Pofg01PMkJOQhsnxDqWq3eRoTIFgQmS6ycyKJGnAcHwO
Kaq8KVukW3G1VRy4jd2JIyRUUMwOZDqcCM6r51PYr0gGJz85haD998pHFjGYG6Mw2Z967EllaDTT
txgOEuUUPQ7yDawopYW1+X4UM2BpBxlgTXBJKqZ8an2nZgzwvS7tYIJoCX0aTzm+Mvj4Hc0+B7QW
1Cb6tkhvaTWK2tMVAfz/Kj3DhXhHuf640c3a2L0zzCnshRqyBgTfNWs0gROhd2HC7zW/lRXag601
C5IPc9FKp8pebvciiwmdt/gnFzCgF8f3ToJHuAcjYKbFpalmW4CEOd53OJ0fLNueYQTtT2aU7rgd
LdwSwXNRuUqmZdZJ+3O9ph7BQi4Xk3KczQbd7fzSVLFs084Vhmozus63ko5OnVnOty1udyjFYkdS
NBs/KAduE7K/fVGxonpCGJYxTyFk+NOj6hPLXwjS6mLphs6sybRqSqAT9gJwSJXJ23TDVcIzoZmt
LP8e6lAkslp9N2HpbmWrJvZL9hpKIPm62uXkNIiC16t+9V1NJQvwUuf2XKH+JIVfgO0yBooS/UQJ
OT5VsdjGVopme9b0LINcaE95v8lFSW48csFxhUhm853z6424+45Rh+UHh3exb5nNDsSHYv3cyEKj
sZHWKARGYSDhJcpGOL2hIaOYHyP5gLOZ+wfoehtl9tSAdSat5sNcVaL2dVkQDs344luf2U6ffiyd
nrR4Tw/ArA9sW9zNBbZkD+WWTJWPiGNmHia+iQBZg8YgsMssTyD9n3Od3oqNaRz2ylcSOs3uNUDB
H8BphFJnw3W2LcmKX3YG072ec4piVFhg6vWowZrd1aMDlip3AqOgsRxABjHbwt1egtT1e3AUcLYd
EJhXe45SUcr+YOO5Ovy8/6q7dBxuxhqfc7+qd/cJvrc581WRDrJLw2gFHDcOQRxI7EXdXvMdujHj
WB4EsDjG/LuVqTqvYXMCFPGRjaBSQmmqB1zuPk4BSc1QB3eeJP3YbCFW6Xw3BT8yBV5eYoprr+R2
YmIx/rW2qzSfOXIdwMapg1ypugSL7kmEvb/CG+qFHRorjOwDWoh79JO5GJYIm1bLDytBeckU5Lk7
xSRpGNVSYQ//aCG1tN54kY+3NukIZpR89tt+t8kr9/IU8P70vFsr+4RNst4Qh9RPknK+6SeDiqnB
eP9iA44bhAxKWEClPIIuDAJTrRL2D9ntFU3hW3uYDJ2Jb8S5dwGXKc4mIxHd7/ZOZSbGMbin2Auc
Zn74X1jyA+lB3kAKAoDEqGsjnntvdrXqUy+zqHAGmMeF11Eh9A9WrFAshpQtJ1ILecN66Mrb/8cO
2Wp6wUNSpTvIF1ms8OFHS5rFft4lGHjhtVvvgvAyXPkHMASgUjZWNpAhHAKrDUKuh1QCUDeiRfL7
fVbzkR5/emofntpU07BE4yfv0jN8MV057PF9xTesk5CaGEnXOnkHoTGOPbbHHt+MMEyT9C+fETBK
hVf6iBc4Q17hnEhKY5H+vWrNMiuyDMhNG+BINT+5fGATrhX0U/2T5jPidNpVLbtFMPrBpThb7YBd
Sv1RSqxOwscm0y+U9N37vvpyFHsBVp+tsuKopwcrXx1eBKnGGZW+gmNFS11DvJEwe441ODdXz4Fn
+8ZkoVxlR//0JuMcJ3hn7Dbrfw10PBL9EEIhax0/mV3rMVDtgjRN04zIZxlfd70+HPnosgrzPLef
P1XAyatkKJuWQ/wCJ+8v3MHjHsgxBUzBfMf0FdBzotADKC3rGO5aNX1CTOHMNYFataa7pI+v1ns2
4LKK7gszoMqDj6BGMi45NWnH1pMg7FEqSkCKazWxKy+ilgDxa/ZUhcToohISHQ8H6ls/IQ3t4pM2
sFrrnlAXzANOm7IQbhsS7TlxbQoukEQ3rFKN4sY+6sdYiUaPtKW+YwaO1GD2fVEryFWYyd+UZOh8
0v3+05t/ONrETaSDOKVSmfXOYYOqwkZCLp21xZCDNFEV1vs+wK0DKfPDhkv1uOaZdCSzJIfSJpiP
m1DQMMjyN6YJ1C3COeRlfqBEzk/cKavIYnrFR8uWzt5S4w3w101WEg9oWZczQ0Z8092yLql44dUn
ZNBvqJPysSQG+8tmX5GDNDnFi0C/o5E1h1jWEjjdAJEYmsGnvUOvX19n+j/Q0bCPcyhEUMW2Ypcc
6ASWs4y5Cu63TEhZLYDacOQGHFNHH3/9h6Q+dIp52Q3Fwgn1kcBG71zdJ6fYS6b042Jmv6JIIAaf
yQUknFa7/sAX1kEdSR7x2EYuFNV728aqQMlh4IwPdsyhwYjx61QttSaNtI1OhmhRkxc+Us0ckhca
ElaSnCQ5LTZD93yY2lXSV1pfdGBJDiFG3iZSLsKKEW0+Gsmd9dBHJAKhI5RQECYew6nbrigNCwt1
W99UEKHJfYajCj3/OF1xWRzvSRW5t9zFsNSo7i0Q3hHmpijIj74r6TbQcGXTqUA4/4TKDb1M7vYk
20kR1X+xr2/8wvjSgaEZo0/x/TWFrdiWyW1j8kI6U+GkthpeccGYCs2lsqTTScxFa324tAz70Tj1
B7gKNjXmoPdHAZvdKQJvs1RPjPwT9K6a88bWo4TRhHXSymgqtM/rWHs49lw3k2dquQulWcRg9tX8
B9XlSLKoHBjubrHpBbLXJHuFrlI6cVODXWucNa7iyjzG3svPL29LKckqAnBSw0l52asYFSTBUfLa
087cb2fF8wnTOckCUkoSgDHlkqsnOD8Oz/InLout1KE+F3aqYfjchiE+yNkk3awweLBzAyzQxDhI
v/KBoqOQe6ylL0qD8DMrLuRlZqVyerjrNGNOOyfK/141OPXcIrMP6TAaMRpqSdd8cqTyJ3okgtMR
pFxO8xlmz2LDfZJwWnB1E+WTz19yh6MfxCZ4V/KyYuzv2xtXTFu+sQx6PcE6ZeKNyxyMiPl1w+0Q
aZxo6NVfpfTZWwcKsTtyhm1DhD91ZU9+DIZC55La7I1yzkPQFce37dc0g8yDhyVWs/sp+SYe+r8O
NzpksxjLuPosCHoD/fTdq51UElbA3ZBcjplqdsWwRBpMBloSvCroSc/bkSIt6RB4p6XSD1uS+tlu
xku0ZDbsUMD52e0kN6L1aXbnZ3YFtLCYIMOILSyMDe9MR5uTayy6wSiFA58CjVlQJww43rfKLw+M
6v3LfY5KFhp/MjriQiUQO4PvC4a/AoRsigHGC7vLD3l4Jmu7wbAyWF03HNqVtxJmUPT/eJMHpt/W
9yobg9XAt1nOYddfp34yBZVZbFU9hy9rOjsmGJDrrS5/w9SFlvQ3betRdRbPM9qT3FcFcwSrBP0i
GGiLXgckCJg1uTz8GFXcXBDocKMJa8QDX+dnXxHBDdbjdLFayF7c4ANDLMLV5NXQO5HTQAxCPDoG
+5d2hlUB06J0VnAtg8qQNPxSL5aYAtRySGbxeznRzdoVIqmw6CQ4DuxezckVQTn3LfU6d++4QJMa
/5YSiKhgBSWPt3IcxZP+3mcvs5p+JZXOLZ/zWNo5h/hqNQI7Entyjj4ZOv5BXNzg571O5lsraQ+w
oKaEtTBsfJMjywp/v/9aZWVTlA6gd7D8p8RqwGx4w3j5D8ZrlxCJ/p/pr6O8rqsvpkDOdsEXEAuV
ejz8/JJmP5BaHiof9dPI9AXX1RgJW9G40+VceyeFMcnjvtN7evWBWOvKK1PVyswLkD8+QeYuHdhs
NykfrU2dHAr9v9J6+gF3OHAq7F8aP8J3vtiAbC8KwqU2xTuUxEgUS1C5gf4PGi6XhAv26jfJrN5D
GzZL1UWhIQ4IbdcprafwW6hNcDMNJBJZEi9tDztAvzrANIB7aWYur6WEQKP7KwRMMurFLtjfz126
RbJHR5N9mR+ta61m5PsEy4Z9MUtpOnmdTO9gWupr3F7XBBmz3QNkSnCGbtWPp5ZiNpk7Drd+f/6U
D7UfvuxfNURHoYMKB4IadPOzXxoHyLmN/0jOCSHR6GDjQUf95M4OqjYVK5FzTKxb1VyFPEIe0GSg
RKErji1kBJksfV5F1fkqiB8wfZCNMDB+6cVl3kbXH/9cii4s3vulzlYwNi6n6ulAZGLUnYmrNRwY
EgzUs1F3ujsY4e2fzQ7UmhFNng19Z6+rrUzo4jjfLOpRp3gWtN0Tyc5xtlg8INWHMMzGDfJ5V0wp
U9I+mCtLn1CkieiALom8sAssLWPxibyZ85R32D38hOj9E5wRRQ4+CixlBUNBd5KJUcL28yG4IDtM
IoWLih5awfP8KgHi6mWcoxdDI+KxnZcgAX+rl5SZdp4oUxKxrSu2uoFYetoVS6T1xGW679PyyNyr
L7aprQ0Fv3Kf4nAiJECQMm5gW2/fnH9wxpsSsPww3BtF3DNxb2czDZS2z2npSb1ygWCsml7mGiOr
qQd5NIXYBxzYGcs8qsfvNHGjKpntokXE3OMfgth18COfM7QnQIDtdofO4/4GLTmLYryx7BQzlX4h
pyefoEeMOHA85BntRTN0tO6qXVaQ1VGCu6BL9WMuUWYv0vdcjDMAOeHK8/pDnMJ2pLxaBUrXXsvI
AoW3xglZZaUuf4oZwLClFXYjdKux5G2dYiYtO+rT3T///icdPKegkGlz/Qo86ijm2gTU4EuuXo1h
AyvWN1eeBwODFt0NUer/xZ8PDS8hKreAPaQzj47jvZ4DRUeWCh1VEGuAfM7BDm8pkobbu+yTijAI
Zl4vdCC4OB2zEx84fSZ6bfH6USESg+XfTicN/ggkns/zouH1mx2gQZQVHAK/psm1nqWFrlHAsmun
Nq8jqSOmz9tK92BcVYVaU++UU2WMVKRte52iljM2pGvou8bMsrHlfSBtEy4kGx0ttducLaoW+78a
rIFeU84WzL3HDfYRG/uJ3Rm3xgayQ1NJWqkFdmiYmG0cdiTYw/JnwxZ5X5DBHCiBY2MP8/KnerPe
6Hs8syIlx9TBq7ufvtbguerFVEf091lJ5k0uw1yRGYbOM7597mJ0G9DzrJzYS3FEucaZB0PC+gMJ
+5sn2nTvJij9UifOT/OGummOrBcR/mr6hFVo/9Kxe3ijtGIyJIg0JAf/Sqp9whDvFX3V/w2G/ErR
8SFxdjjfbG5raGVQsPH911OCO3YskdarXRlvWsLaMu/5/ChR33Mu8LLtyk3GkZMwQstcZiKZIZBr
lrSf5pc8dRnxVmpHY6GqzjOLqsI1CiMpTDmYsqXmiP7hqKIrAycXnJ4Wz703sAWKrCSe9jUOoKAX
EIK9Lrl/frxhqFD5kxm+F0N1YsAWUGIGtAQC4gquZSLu4z27pyvsdHqQq0PWMqtY2SMVSxh5+fIs
gtjdJaLHTh7v65jaKo2gOcQOb2iL9Jsa1p1yixKjFLp/Y4o6cSNtLBctpyu+E33srnlD43/aiZeS
R8kXmIcaqJL1S4KsKtSJW3CQQOyWPwANbpu5/jlYSjHMoqvw1ZMr1M4cEUMbUdA1yRbZusBHrVY/
HG3Q8ZBiO4ZGeBTdrSCKgEuKKNII9qqDhPZFxdv+ESXOH9i3H7ndz1QxtQ43t139+u8Sjqdcka4C
lF8ppXwiBzdUg2IBrw4Bi3okz/dN4aCMpH5L8z9qn3ju6K1lZWL3o+oPs4HAkHCryZ38ML+tQF0+
HTpmiA51/Us/LQHHWejRNkaF+i+g6/Dbie6YwfUBUM1frPw5LTgPMzKweN+hqmrjJlAYqUr8gdOy
lgNTkLvEBbbvrtUi+5/iQDx5I6TnD+pG1PgvzAqN6US1uDZsB5/0NJzfzIoVNA6Y+hd6wCDKKPZO
EGHGLXgYiX9bx8dPmMOhL5LELut9REPDVI5PKGxzlvpnviCNGCCaeakx0qJhGyWAUgvG76mK58lm
XpPBk1sdNkDuLZokYpiGITGLXrWjzWKRLUM1/ukkYGZ/9gDHnECZB4KjnyPHhqxzqDRojrdG8xqr
bSuWxDae9hSpNId4c3MKDocdvU4gyIxtl3AOEGLwLGyaOMaKcNBe7x3l0iGLVfsQaKSEdbY2FaNE
DTGeO8OnkIIfl08nHwIhRY4SC1R6qFyl9pRfGjdI5zPZtbtrEeQlcIhM7cXmsxVbeWIwvoCZaHnQ
rpGfc7gTVYDWrALpq1O09moQotFwoDHmqCxcZ562mTUm8t45sEMbOtCm9VBba8j0CeGH/28NZVp2
+y0K9RcaZekQREox6k3v62oS5BGT7kojNQ41hAtr0NP8KUKeFkSM5V8oIYkjEOnYk8ZKJbyE43v1
VabnQ+BTq8Mz1NPdCgNjeXNEd+QTaeG2VP0tVG24EUVcglvIefCLVAK0O03/dQ54kePchgXx0U3G
uhs+cUsSKpgudUvpngeU+NSRNSZ6MttEJV8GPxxcEzA3koEGR9XDCj1ihGka/KXPbvuOpP5Q1wxH
oaIlvRXWGizt+Z5f4UH3XvN/dMoYl2N0qz3njV5iflzWSugI/2PVRE+T3KMjse/uCNURlGSa1653
Fn2HBH9QXe0tSjUmveRNy1PvgYj5pN3XH1QW0o/DeckjN7gQLa4w7ldTemcKdfwVhY1N+scHn7qu
ppQ2+G+c0VjudWwEi3oUZnj/Fjo8vMaEqP2WD5IK35CLXNpv4XjJ/4YKi7Z35TdZI5bUvWuW1CLf
APzGBDzoBraNXzs/aWr+iDnIVnQxUo/OSZ+HPlqpruFXXDKfCb6H2Rt7WuEClJms/0OwDKLymezA
H1w89EMiq7UycDiWzYBmiBI5dfXNHCfNexEsdSsYcQp9jjkNX3lBX/f7V1lDjcalBQYQ/sZio9XJ
4nwoXY1zdQi8IYOylxHOO61TQ0IkT7kKPz3x6U9dw34UfEMWMkY3sF6ZzjbUq2o3JyAEm4WmBLmY
p2rc/Wu194pjfTAondlq+P8tYqcVQOOaQ2UAIMCcd+N8dkiFyzepORfEIeQnwbDLzmJZTifv+hgU
zyQD9pBjiWF09HkSl0ldV9al6dI+rTKRK02MbAWdAQ7DZCqFLiE+O+QcDv4++tYOrAbhwXYQuO8u
wpcX4ReAME2iYjVP647KDmxo/VB0yiE0AZgjRQp4RVqU2C7HE6sCpKPQGG8wS1Uon0iVOh0Szp13
lm4wdSbNJyr1kFGHLY50HqbU3kVRy0/q+uU4QxJiIQqn7WRuqnotkSrjzWp0ApNSWn1KaqGGGzxM
lQVeqvIhO760NSAbP0tGeYW8aq81MxrW/jhNID7xO2sY/2yqxQGlKntlc41x7OFuxeQcdXTydqZ8
j4nIg0r0zc5iEGy0wFu4UPmuxfLZrxgkscrgq9T04mkyjTH6osmmODIAurkxd43JPxOHvMc8FPeJ
fE7QcxVkXBPrzIWEtVhDtWCI2TJzdZPViybSoNPn9V+SfMzM6+VopU2BLGgXfW9KbOry7keOOZDb
ozY/blQcR3jbBgbHrjfm+dr/+bnKQF60uXYjEjibnoCQTXwCGf/Wn/qi73qkMmCg7AX/kk+Kt7lx
FbuzEEP7CUfSiZOmrm29Z7qTHrIrokI4w6jD32aVMD4h+DMQIPpPwMUEwyQkht7PrXjI808PfN05
OsFnjKE6quZ+2a7/dgJspVKPtiUt+qvb5zgOsLALvnV61GcucCM9liDWHJVnKCm4ESD5xR/HpCH6
iQD7cIoGLdMq6kKsbr+j52t5V6UUSU0TAKa8SWcoPTlMX+RCUlnHWUvIeZvfI+rKTWT4nS/Z9L5W
ytmZeR/mzcYA6f1CNcNG2WPtWxe5gggw7Siudd4whGHhB3gnGPkHt9kskNRGi7T1vMEBJSGcU5fv
m6foAt2zvWJg2gfFxJ7Ks7ffq7v9DGH69PDjLyXgcPuj6QKUiEOK/+5xYXe1IFprlquERPJBrwBh
PtPCSGnyrhWzX9wkqCWham02qwel8IDNcSl+aBwe+7Z1mavZAE8FQkBxMPjzJXpVMrzG18Dqy5fN
57XMZaMuJ1IRlW5/ONpqdyKJghBIOzRQ86P96uOLOgAw6nn3gV/ncYdQZhD8VMp6c2t+D/EH1oIr
qURCJtHC2Uc9FFxPBYg0BL1+h4nwBkRqMM/aEB6GgyzAWW2e0ZmI4264qaUphGOxvxuksNMUmNWr
G3Vrzp/vaDhXnxZPuUzREvuwpbi+euk3GwENBdUbfSNCdcR9haIwicUQM0c7BK0qW+sVc/F9nv7a
fGWJ1nzb7MOhPEmjiMUpe26lWcZqk803eBTBPX86+3IJkyj6txYXAXlrEtr86LMNE0PbpQe0fn63
mscRwp8UGV+PXSUX8ojiujxo/0LkVJZwheCd//q/TvHiu4U4Uax7Vkx+HL18mQzMRmavqiYH6hcb
a4LW+rtrUY1QPrdA8GOFqJhQQk4yNkcGj80hsjoeWdfjV4n4+T5X0JjAyvwhifD/xZIPHcKvJvtZ
6z4Hmrovsz9V058MPJOHqvulBRPRsvEXfOhhrptQZ1Fj2ACNoWib704B/XVwoxg88PN1E/U7VP0D
LoSR+EgdpvFU5+EfgftGQdesg2W8OwZrExYKWktokMyHVR1sS3gtLpuo9nFRh+8TJZx/HrUnVdCA
Ve4vPvqcWFn8oY7GT5ZQl7+aSEm+8vcvgrliFtmttSolTEvmMm4GMhZ+8He0duI2oNz1QWfzdBsN
5v+hHsPFUiyMZYk2fBLIypDl9NdOIHxwiA/yHajQ6LZEsjDcBeA+joJw8ycR5oCmtw8R0vdAhabM
eOU6t6z3z/IReQAKjj5hMxR3ucfa5MdXlyYVtBtZ7B3c9QTaidRHDKIsiv0ZKr0nQ//z1kuVX/+0
y4WfhNauFAL5ZyIPQlW5i4FFE5t+LjGj7U8CbkQIN8HOTSzvuxBfcXd5oH20ukFGY82gWpkADauX
bRLsWZEpm27JX4kD5MSoxTDPbqdKXfs1QRVD2enku+OGLtQxeZliR8aM9X8iZpwbVulmoqAObqEh
qAiVxZTmBNFJ6fX+o5vd2fi4vFUUchByHN+0lMu0gyNwtDSrYl3VgwBB1wCRvWoV4CWf3CYmpoSp
pCPXt04NK5s6aEdzwmAZVmBkDG1nfQ4GAmllRtlb6EVsLh1eSuEt/nhYrHypPOVs4OHnrz0VpR1T
f1I8w+XM/b/cqi+bbwIPSGanCOkFhF03DsbFc3oiUEaFxcfs15aFUxSewwDvEhFqsCTr81f2UbXu
ECQ2ki9Laho/zNsFdJVHsNuVSfoAFHlkymIZFpFEYzbDz6zQz5NW1xS6GSmLxgofrMDxO98Ivw41
4Ff1alxzt2QJVplvT1KHcKOLsf9iZhgEfu2iVYZx9rfK7NjLXGUTDiwBVfJS/UL1GguGXrdBi2la
DM6B7Y55TBlzFdSCWNhe3BTR0KxcKp6yyerM4So4Tg/45cky/2iohhClLVNXakkBdXvroe9f8JmN
9Z7rkuF2kP1BUwRsm+raMnupr2aWaNlUr+Las1TUoZUrXjUfAkRZ9sFrAndAZcN5FD8CgBRiH2kS
5H50mjrfe1Ly+wSd4Hs7Y2VHUHbKohDn54/jz7pQpQsyMLSXFrw2dYsCrQ2IDu7Pu7DgwA41oBjT
T26M5aqFEXM5i+8cwiUddVZAyD0VZa1+0wrQjexfJsMQDZp7F9p9WNSEQR0eTQYImI6mtBDdIMSs
UMrfGzI+/FEmmS0ifWE26ew5aOl1l+qoci9NQrJnnwU+UCV63wurzWYAvh9YgaBK8FbZd/yLOmQS
znBhUPxC0UeG5ExsfFd4Qa0o6doqM8Gr+lZ3iBxsFn+yr6oKq3mUpHpWDSvCFt5KHaisGA7iVmfs
ZnDsM5ff4m1gNb3RWGB7LcMvgLcAruZMn9MKXn4GOHRp5jJWu5FJ2/sr0/Fz+IHxGqzpQ+9F+t5e
LAG0Rw/hkiqVpywFK7zmcQlbx3q35wggmA7eI+n6khPUhq5qGa6gZwI8fJiCT5zNMh8LGyW5vvJz
n1JBKs6akag/8onnm7xOXCLIW3x3GaGmREnART24ZfsbO11ktk5XW2jYtU0yuhF5yMzFFrPnV+fc
9VacW7IlTwrm5EJ7mh3lBpmN78Y6cRpaSpYlhkvxfdxjijem+mrHp+2CrFm4T62B2KTQlkpIOqKo
NWHFl3hD/zdyBrxbYpHEUnIe6EF2FbXJPV42ezdn2Vt2hSH2A8O/61lyzEKrfqfl13KcG9T6cQwY
0MHPnFchQ5G5vhDvv5oeegmRTx5n+oqmI1C4vXgImzoS9u9e1aLdSGD5jPoCcR6fhIHJhBvJQQAg
pmLgVXYRBs6mXzwI6pgc29OP9Xg0MWwrvZxo3+JqoSBMuv4vMCymJTGB4a1NG8p6ulC66qlH+WS/
pIjPmymMTj3JtEyJJf0Q8Lmu4lEgN5vKeskElrbYx/ZTWdPOcRWqY0kiPup+T/xeGGgGf/t00gN0
EpQ5NJXy0xNLxkBbAtvgQBzCMG/TLVebAypxGEbfn31qS9raQmO6qnySVNwyQPInWmyYGoL8PkE6
LIbAfS5SSLmxuDv065qHo7l0hk5Gx3xGRuacXJQK2FztvC+D5D5d0E+TRzgHxzaOzkY20OxRITJK
BxglyWSWsV2cElj3bpJaABFKjnUPy1zNvMwO4p88HBWVi0TbgFS5GnvqZxm0cB78omNs8HnctQ6T
lNVDCcrKsf5CEZ17mw+CARVNiEYt4fc/xsMlx/eaohfi+1dGertzF0jjmM41Ky5agmJtXqljWcYs
zaLy3VT4Bxf/NX3QtQlDuQtdWqmDRhaKzm9AtfjJAUrI4aqzf3edb31WZDOYtvLv1vAyoJof0S1J
c6vf0y90UMCIFEBX/hw2HZHL+mssJu+85Vj78Ctdd3t5Z5KVXu+s2VQGBOyV3Z40+aqq8Xd3+9w9
iPB85cFfXyLzN35pCY/wbX4+aWa+ZoFsqqZgsxygNQcdQ+V79nQlf4BGBdt6bA8ztgakspaPnmmj
J3BGssGyqkJNWO96FqDG6a0c7rVfczRnzWu4wvtEiMTNG7TMU6z5XAbTeRJYiAYvuxMoFIeQ+fP+
Xa9FvhNSfHfDmo3zYISGgRHCeuOlYyCNqdnvPEc0dJ0JyMd0+PvNrGNU5wBYXH7VxO9OXXP/nDED
Fe8A6+YK5gX/15xmmG18wd5G4kjutjUFXJ5cZKVV1BDBcu8HbhcSsA5UTjupPESBWDvtSQX4dwBi
50PRkdyz1WPOZq3MIvow35aBf5oi/HB3U8dwlsoG9yTC8JpDjgKQAR89GjCrCH2k7+621xIqwo8B
a7vL7quvHb0eWCHzMperh83b/KBzT/iSOiOPUPVqG4cpuSkxrJUgSc9OkiuRxe8giA2ufLnBczvc
Dni9Ru4bM7ZVJqUKJjw07x162V/ej7w21Ow8L5vrrCjMhKpwV4SbNWrwfcOB1B+23d5K8Z01H4V1
IwxqKPVvOR68nSgp9PJ89oxuNCbqUl8Dn/ABWc5t34vpj6UPsQluE0hG5sfbsGyXMg69IonfUG5S
KmLl/dLiQHh0UNmc9YYoN+neRrHnuWMSGAg6Hf+GuFwjIDijlTBJgp+wnvmSun9V4W7LsghScLOy
Jp+exF9fpDWKIJXzv+pyQagrxXc0zrn62qOoK0nxNjM9WrFex5X9DeiLrmfeVSym/1FAZ5BVqF2y
mRQ25GmZMHZYQZ9+1vKyAFbIgSvH3E0mw+HqDIz6Rg03JWwXOLnCbfnIA0FBR8QKDdVVC3/OZbFs
1NUSt5xKllrZFBYT8O1B5DgnilwM10OKS/KWTDiLsUswuKT4quLp4aK/GPCLr3UqGdBmKsuynCcr
+AZo1rciG0OsVF3iBYQg4RQtJNQMS3dG53af+II4KNULf9xs7iKxscQkzqz1sjoMnYSnnnhiBQI9
0he7j+gZyzoAXNX6jUB7WANShrVyYrSGhRYGsz3zyOc7JtLRVNMSEzONoC9VAkKvjNbGqckPSoxp
KiFN+fbGjymONqIMnI9OOX50rjkEMTUvwAbjBIeOl3UfROFYOwLIh2CkggcN8clR8Kzj98XzYCGw
hm/yCj9RyoWp+7ckxqCspNqWckj+B8BpmJSYyHXvXthXDX/NeJziYdftFDJqbqKLhiQAn5tbIH8C
KRtNDiH3ueOKin1uuGY1pNiYGLpy5q+UE37+Jo6JKysouUmDjtYdvZsUomVU5ekhwWAyC1or5npt
mKtWU2UZ1KgP2m5ETNZlu1+PSGFHC4KeJMr3n8rUJcB+M2XCGpgKw8W7XLMEBxjayeKchx1R0D8G
oyDzKaldnHwWnkWPDZcnpYRz0G8zHSfhUuqAIEEGIzVVJInLSFefHmdM+Dw0d0athw4gXBqQFQbB
v6oktdN7165DGEVhFpWH2HcxRdmV4siZqkw78ASOa0ftbEy4FgueLjeum6uu3G4TK5FJhiUOCLna
7EbZR1yZdFuI3ps8wXEhOb7oXX+ENGAJHXMcKYCsGzCuc5MUjbDzC8ObypLpCjkMm5k7RV85penw
PKGrxEqznVosqiO29gznrFbUMvJmd3Xa2yQ9xg8OrzqTyS903PjsiOKWkz8p1GFRFYqvnFw8ysoL
9Pj7PQlNC32ZFd5ntWX6r0ZYIp7zQjHQJuZoS4rWFMLTyfYI1NOi4bEmoAT2h3J/OL+XUHiFmeei
sKB2W3j5Ex7hp/UYcCzgsTbvgs2tbE3dV4llJLkaFEJaHLKSzOSLDevHiMo0pSJqSqR4HeyEw80A
/FZE7/UkH//e4GDOFXJx8S/EOTRubVSp3jfv0h7EmXfo6ocDv1vHOOvFStJoj74cXuaOGC0NfToK
ebIPIzuEeu7nIWc4XRCu/aRMIT/5JSohWLmgwFN43xZKLAltYGDZKz5d0YgRDD4LdCBv4EPCre4A
EI/XsJbHhYDpdNk/B173a6SDtK/kHEt6GQm7e9tgnlmulbZZ8+lgjFFzd/r3tG9K52Qaj3zn5/Kr
NMNEAg1JgTcuvYUp7NgFMrkq8KpdKdLv7+HnSxxqnjlq23WVE1rogl5JA9qZe6qHVc+CmJGHcd0B
wM5e47ohvj0lcpRree+Gjczg2UZxn4f0ah0Ejk39qIFpRrm81f4bMsC1Kz6QY1vdOtHjAxu5WZO+
TkKbLrTafiWivxPfFbCr101QNxOpAQYGUayTFLXmgoMh48hB9yTCvI2YnV9Y8VdWu/S8wN5yuBFm
VtQi2aqF8CxDPFlfij8ykawo4ZtinBZ4qpCKMZAJ7sEJCQkJ5Ku4mR8EO0wz8PJ2REDuJfrrO3Bd
HBhshNJWRlR3I5boM51tmpYpFvSBKJC/I9EIcHXgp+x289NBa9sYs+oIkxISHjjof24n5G4Ivyt4
2NhwAcwdlgsuNmuTCimsKuFRCiQfeL0TjlG3fe1O3eYRaLYWf9h5EUmuiv6kLi6yu8j7qtJ5b+OR
CuF+1LdIxL7q8tNq8KPsIrIySKMHhI38x9K0SelQKhM7CQtvDOskFBKKrQgKfJqMMtTjSpeK94Zd
42S3pfLVTDsY3891+cT6RwFL07caF622ejYHjn75yAA21cdGWxLnxXcZq/8kUuzZfQvvzh8+GdqJ
3RNZuHViI96Nr+e3Dojam3qi7KLtU8xm+1gkCabQpD9yupcG3P4AYdD/tqn3VgMd5Pes/2vHd6YE
x9oGRp4srjZexziT6UxhRCJP4JtkbrNgqfn0GxPjbroDOLyXZHgWO6GAaYxgBhy8KDlg762JGhtQ
b0LnHTT0qE3CmGQXkLncCtX5bFL+4SgjbP5wW1hfyePpPbf+ixezIsdxMvpx2TbM7UiuMfc/tznj
l/SKYmy6P9mbCYD6k0UBrFXmjAU7Q03dPIfbxz/a9Sa+Ev3iM93B6vx0TEgnOGtiuEFz4Ni5cc4N
jTo4QtFYiDELpP3THRgwwf+OGIajBbpr6Ufs3JAQtFwoNSvbPBGZ7GjgKVZI1i2EOMOyMTnVAanJ
9sDEQj86en7aznca//nI5foquCuk+cnjRBKIkHQEI3/5SsSZsBYpsYYmTmWNIa6eNYxV6uyzyVjP
IiJ6b19nPFWNpXLkfZOvRvxWlbvst1m5nndCkkHNObzi7BuPZb+iUEUO1Bd5qjH9KkaTin10NTyY
hl8faP1cPiXR+hwktUeSbz1azMIq0shxFVdrk02Evuj3HqXRaTu0YXcSYiAGn3dY4dtXF0QulowZ
d3oHpAZXkUL9uUudlKtTlbxOPiUu72bhJgfW6cbFbdajBuZVuiHh89nHSNqK8tIcioHZCx6qWFkL
zMqb8MC0b7wIigukffSJc/KUimC5fzujHuIfZTnAmof9i+v7SXixG2P5I10ByJLlckyPapajKwIS
g/fybOZLI4fWCK7PUHjV6YRkYmyfonM65CtH1HWSNwqL/3jP4SWbhyv7koK174iCzvsZdnlGpuso
CduQtRVLyF4BYInQh8QzdXMVVQueKOY+p0qgh/ELRrnZlFn5GT0qX7GfEJoor1jEbUumgT7f8k6W
YDm3TuE6ueAXUE5+/qJsBTAApN/aps1Ar2TQW3tUuEaQfDtQBwpwSn2a8cM2FKUgozHaqRDYkw74
g9AZ3CIAptSKq84udrEMH6XTYMQqWItGAnaOjlET4fdEK3AQ7YkP8LXMNHAyLaFIo0fJvcQKixqA
IYX/k/9TovVa/e6YiAz95R11XCRUknPQbJuYK9Fjj/3jc6/rhkTamJ/XTkG8+cSFCYvfpKgX+nfy
7ujuK6nytq7ikaTIbzhzBkK/e+IuyYoMhUEaLCLkl+LuH4WHglsnxeOBexRoptt8LDAGR/pca34F
GfUNresGo2CTnVzMGa3WbcT0CpA7Ji5u1Id/55CO48e8rm8wi2T9Qb3eGrYLYpR0f1sJAvHO5jLl
PHMnmvuxNPxP7kVsQlDJH3PNVlEhF1Dx3hwWit6Pk32jAg5mDzsBiqASnG3Iz9M7RLtJ/Uv/AlAH
roGJRL7Avz3nWUXuhPbNgRwWtKQnFnypRj0CuvdtIYTx2DX0N6nogiCSBIq+tZfiqKpMRbTt+pUA
JX+JDHRLwJ7uv/E7pdbjs00aiMrBduo7SK9GB+zB4yRKFhWpuiqondoyWFnSLI0sI9dMr1rz0Iu9
+j3M+1xi5L8xuGkREdfeOBMI/4+BboQfw0+4tUgQ+h01vEds6l9mv1axvV66+2WX0U2PrDjEmmiY
hvteihOT3j/U/vTc4IVqG3f5MU/XnlgdG7exP/rDbDYoYz+qJ3OcI129BW3wq0wfgYkGSvrxT23f
I2OjhUjimOHgH+kYUS0bSf+jKYCShTj5vGn4j0ZdcdSSqXa3ighWNbQnZqrmp+s/Ku+2gIsIyul4
W8OwAXOjJV7i3cJ6HRokAbHMcssVtYW42UxbH4cmudxTplZYv1qMlDv4NqAkQ9bhGfXvpUHA/9mj
jEchHzdhDI5SxnP68sJDgoxA8YiskhfsfmEyDbSRIl85hV2pYP9SQyJ0JbHGPp6NrtpmVRrx5Z98
lPtzCvvdW4ln2stJIS+u55wlrEicV8vL/JvcVCXJSOErXISKmpGfz0y0Z6DRJN11YZIVU9C12ULT
9YXpXC7sGMeEyJvJ+LOeLgbOA+hJFdU7ZF7HaoOSv7ni1peRuLFyJFi2/nRpBQRXUAxKNiK9ot3v
4wZlgW/bnD/YksrlBIE26Ab2mWCEanSpvhoIXtlCIVzhBKb2lEACzXGmbyVx2+z7kt0OFF1dJ5Wo
d23s7lQbwkn/h/p2akLfct4gLl/wdGhbKS3cuZx51j7yNuUYzLfdBBH91t9UCnw80Z8xa6/Z2DLL
KBUn/huIAFo1wpoQaAH1TWrWYEIzpSnblQygf7Zte38w2EziaqFPt+loL4KLpIsekQinDsMrHIe5
ad8Q53tbve9MtE4sOmA+PkErdtelt80warlT4wRTarfIZmDzFM2T305gY3NuXcbSrLXbQZPB3Zg9
xASS1tUQk9cBD+g1P+bD+XO1nYWCQhpaHD/7tw5K3do69z2NsVWCEM6XhvZdWpOm972t3nM6uEoA
Yv2++4GP4K9vwQvcS8RrbD165W3eLpg9qS8ZpT8eqJmwFDUFC+oj3S+yJsBDbJqnctNk8nsVmmeX
OYaYs6S9BQpzSN75V0VOrZIwZlv22im3xmVLGLMUwJMxL89LyKIJuI/vNzwHykKlTLKSKU4pT7WI
x5Bl04tr8LI8vmnmBfSxTClsDCrjJntz9z29BJQSnRJCTmY3F4/74CTh3eVs/NvzYkSwZ43wKAH7
dJgdFmjaiOiE/8Y7DkB1jycOG0Ol6U5YehO49tLXKOwWc9f9lM7q5bRoZFfc/gtmDP17AagP8xBq
dKv632u2PW48rcSlIJJtOYW/WA18nb7zuFSqUsXyy34HwRGMxSg1QJfvc9omjNMF0A1VAtt0niB1
e2wNa4kOjTp1WhOFATs5GNRdC4M3Ov2T6oId3jhbdnJVlT+synhLdvp+wUGIr515EpMu4xvcho2d
aBT3kzVZr0JjuZe+iuEvzHNQEMlSNR67+jTx3J/Z7vXenVgjgMxGpwLIdsXQFGlgxVttQeMkicAg
jecKnT17khXUUIFB1e6zogEVVU99wwYtH41ei+Q/K8f9Qa2Vh9AI4Rt80Rhg1WKa8jWFcsbTMKbq
VYpnq/c1Ch/NW2j/xISpDA7vPcCqSPsCv7EwWHsvt4LT4dIsdyX1f3iO6mV8nYaLcMR+ibIJ227w
3uayp+LUgvniqASzLBStk7yLY1aXB2YtZ/uvr8XC3bd9YwFktb0Dn9UEjghJ7qWQbegTXzKw83lM
bJCeoFzBosi7IFfhefYPQhXncj3YfnN8LhzP56rPuPhW/xmdSsyHKCECU6czZ9DB5Ywm0qMEG4Ap
rhZA1nD9tVyd0ANgQwmShA7m2lnhrdpOFYsR8hJH8Ib8cAPebrTAk0/vCfWppu/L6zUKR/nMjIil
Ufd/aFQMRxOdD/rmu+uo+T6L1glaoT/MSXROYe4rNfuNkIvL+LyzMnEUDP5/250UxU5GqBRwJrng
MN1oawUDgyT6JFWK5fQJ30BO5uZO5A6sa/AaA407MJLTHe3Z3453wFLXgjbzA2NpI+vqcIAQ1ABt
yL/bgsIPkIXEmgncG27WQQzMmEsVOQg2RM41ghd2kY4mjz3Mh5nLAnM8ykY5Dvh+ThwYwgK7e5QB
0r9oHJdHQJai6LO65E6/Sqz+r5yafXwCtVE9y5Owj9vdFh/zFZY/uJfIZhoGZ8lg/lZmW/sOGOKu
iAyps6w+SYWv27sSZOM+LyPzOJxCisz39SGuuhXiEVbknvVosm13J3MB4/t44tW4prNFvScyVDFa
DjMrOO5zmY+Dq2d3frlg4uC1FatpQbG+aXZMQ+CGCJnj7u/VpqIV3jxJ3RXhgufRCeqX4TU1tW12
pK9vpoEPsYCjivYDJ9GF0Fl9wi3LLcFxF1zlPx/+xu0KMTvnIUN95zsJX1m0ueQ4RUsfkvPzhEu3
A7GYUs/xU8isCs71DL7tjZbKTamEU7ShwYUZU3z2lW62BE4CWRcAYSD9eTbfEy3Xpu3USEVodYXh
8hnFayG82XNnmWALO3xK59lxE6wOy88bNVY91AT/2LA2Gh0Yzh5qMgLCVi6LBQX9+EFDVLkioSQV
KbsNGv6r2lBF3h90ZkRe28Nh3XmkE55p1CjkYtUFL3r3SBajpU+02ptWDbZe9QxA1oNeFIV4ZbyV
aFmVWyfC2JHIHmx+kVsu8e48RdbH3clJC/mv1tFCNSY9HknLQvb0kinrdvXRUscvTmS5kbmvL+Lo
IxVrpTR1Lxffhr4shV69IG/juGsJBWqlD5ftkkGHVTV/bHFO52+tLJ06ldH+lkbxG9SKPJkECxAr
rnjFDff4SKnRWPvMcce8yO8dTCrUf3TLGpmDvZ2HLoPk8rAn+nsw3JaCKTEU+ndJdKTyH5Ul5BUo
w6Yd58v5UXgZZaBw4ZPYqFURE6aiNucm7doYdUgQT5mRhLZrNgwXFdE5msvnUUOSok7ZZll5M62K
Spk+1ng2aDKr9L89MMUGjAwf2n1qf0Ub82Iec5Grr0EE4qC6QrOCx341iztwvowNx2Gqyd1EL+7y
tEbXckWo6L2O+Z4+To7ot2Byy87uoGUvZENBIyGHl7E+BhRp00w9TKVGPQOfaJUNOTRieCmdOceX
xtOUgIr1NmlVV8Ce3zPLCEew+Jijb1zXCrh1NfbY2guxhKWbej/9PjPdOZKba4OHOMk0AwIMKgS8
61r/p4WIFMuEzODQNfLFWGtpXt7w+jOWeNiuNI91U2jVGhR6NvbLbir5iW+lJktSbWiOzFxVQrjp
E1ckTBA1BH6WEEBS8KxzQxcL5iy7ySgwzhaOb32zxn2fbtgsjs4aWvnlMaY8sMTBDX4Ws5Xb9++S
nzOeJPqGT7wa8TiF+DZ4LvvjjoMztAVpDOs+FMtvayS20mou3dqXjLGyU7fKctU/fQdJV+6mTlqx
ydd62pNtb1N15mvPS045ojfsVZhF+y8FX0fhjRxInqLmYc5CI0Dm8LMbAmbN1UCiw4jhFa8lNpJ+
RzmZUELTF7zrkbV0uTFmsL2UtKJhe4E6sCQ4Oj/cKvLizeDOnXAtHcY1owmaAfw2TN2LKzinvfXW
Z7RFfrJrDTfGL35aXYBpAAwGfZZhvVaOnUUUw4T0a+Jr9Rzroo0HB7vX0zfo+gIZAbc4Xf1UWHnI
pLcSZDF2C/COc81YESsQoz7N7+uSG4VKrm2c7ZdOM7pOLvHE8/1DUXEQBHqJzbK25R6ItYvhAgdW
Pz3q82j3eH56uC8//Ivbq0cu25Jz7EmRot+9D+VmI9+UP5Vnz8ATdSuVJrS3VEAYdJW6uI0buXoe
MpHYrs0VYcsXA0CgiaFDPjifvxKTw0Wdzi9I6c0wKJuvolOhw4KbgbDdl1lM1H6fiZVBsj3AcxuD
gu1BEwVenCpLQFVXfeYe7gVGEeKkaQkJIDyyG5AveH+MLp8uRFSGLtA72jrg2NeepPPJ8Ad0Lpgh
guG/L18XjhBa1l8W6mvPms75Q6ZP/s/FJiS4RL9+AvSnDMc7RPCcuwfI8ez+w7zAYVKdX0yq2OfV
S4KTm1EMbTcNYL/x4wku+l4EY1IQ7S8VsdLniQAwoulWzT1PcG5XObh0qwCXQctgKR8AwegaAzyU
1pBohMvXuQNtMZjR/o/hplFWmwb1JZ6aGl2xTbsXK8Z8R3Vp5HS63nc0Zp6BfF4h39+4ZKxTq0HG
sS4Vlnt3Lrcx7WSqDNq9Cycjc/gmPU1t9oIpKu/SGYqMioI6kkPMVvJNjhnnYpG/N+BWODXjHz8N
JOeztVy4/eL64fCvKUTQWMwL5Y34ZeSoGUm5C60TlKBt0a1R+h2QJOwGn9vpzu5TDjBj3bsDloQ8
z8Jei1+X3as6u5KsNvDK0CHlHFmE8tk7jfQUXIcYfWUDTrQck1kDoKM0mhmcuhGQm7bdEdPC866K
5ukS6GnngUFXd6fwteov114C1Tx1rGs4o+MzCVb9GIpWvgqd9FS3KHZIso9ukwA1a1Ql9r/nQBi3
0u6LPUYHTlIgR6wi4W1/hfCZBlNJUSpP8EsvTD83vWH1/tUtZdsJUl0EgbST2M1lY0etvzcpJWk3
u/YyTTKQpexBR0BNznDNtu9c1zSR4snQuz+oOcWxqnOtfYnBXePx4OGMnGzuTbbz9r+I79TaSmnw
m/Kqz/bW8XjjdRAC5VV9F+yCPVkpPYjOpyaQ8flY6zj/spxMrg9nJQUQyZPLZ+vxq9c8H5epXTQj
o5+HBn8kgbHvkmKFAe1tiRvblYKnIUsCYVYb9LDYYcxj1I0McBJeV6FWmwNZ9kByrIglf9NlUd0a
osLhvRl8A6zdrpFsMpgMsMCAlr1V9qoN6PzxYOjH5310G2jPmg48lvCjHW3AVym9exseowjvyVaC
LosEC+2AluAL4egMyp0I8O4PbPwuyvbTOtn7pnKJ+PGnk/QT5fYHCpYsYr3VzurXJ1G7wmjT5EtS
Zcqz3s140ikffChp/RNEQmODd5N895w+YkIt/4EinSVr8JnihVUsjFWPNYWovtbpoCpXz+9Vj/CS
+yFY8BL/Y8WizekVLjCrHUZTiqQRQyw2R4SFLZgFGIvdQGV+Nq8Np7WWSDf+LFLPU0cArE0zqorb
v3lJlARAAYBLBa/oB7vrfjUyNWE+ZxlXkIBD33R/WXrUYEDdPnZ+em3ll1WyblBdoKH6HQIxUwpL
ekw5arfs6x+2FhJ37VJC0OUbe6Hf4+IaCyT8M0v2lDaCr9t+iY6B6UV6P9Z1XpyxZ99Ax/LyvDbz
XmqtPhVEJxz715sHAD9Hin0ENa//tETDpkTMEZHbv/qvcs71DsxiZkknesilguxLdUo59vMTDjI3
btA5S65RKg/LwJ+hhHgW1hL5dVtPej37fJEk0RDS5dt9upqmo4gqoulYoxUrMzeHV0CcsYU9/cQ2
2Gc+gXpsImNaI5XHruDRWfnsQrT2pQdKf9ruXdQL85t5srksOjXMDQAh36c5Xi2pK1TKYJirdri6
fkMtpTcPIcIR5NN4lqzsOAOS5bTfm17dMcBR/HMHdR/SoygQIY73DfIECRGdEfaG8tB0TlpaIapk
vl7i2Sxgo6Vk35NZt5M3p/f0i/U4GJwI55q5qTjlEGLaaezXXkUwfu70cEH1vZKGuVeELEPiuf8d
t+XnJtUUlbqQSRan9ERm0zPQ4/2niIB+Amzrm56kggpNwDFGcY7BVesec7WgYab7X/O8/uYrWaWt
ewTiHcWXudNnjtqwgEW/DulfZqdrl49oT5iLPZ2Tb4hJrelqe0TNihkSnwMlQlEIn3oqh0gYbQU4
C5Tfc9HDYjjc1zXA8cQ5R0klZbK/GAS0o9mMxpE2s0Yw0mD9ZgnYQOUr4eGgL8UUkTuHrtPPqas6
EQ5Fn13xGNqLgdBc0UZa/HGi2cb2KFyzCKa0urrIzr91hhGW9Tr2WI50ThpCtCTO+kZ/PtDe2KbL
zepvVgnTNqA26Hno0MN/xNe8nsHRe5BBkHA/NahlbmteN8/2r/4oT7dstVPY37f4wxoMNuWDT4Ji
0y3cMjqPcRdscDkyWQnhFUXT6vtiFrakeKVPVh6s5CYHjoLOiOl2NnT3zpDkZUwRoxt/nKAiLmZG
quCYAp79xFfVtOCPkuRhESxbbXrmud8C6OHCu8hWJtFe6puT8h4va/9VdH0oBUIISc3PGy/psd3F
Yk8MqZt/A9NA58jQER9Sxh9RvIMI4Fxj2G08XqL6Dx9X0hJh2g/YpopBkmkRuWaWfmNkSikaTxwl
NkFykREObW2/pSCiSbxfuEuyi8uq1KfgobNQu3i9rO4YxPbw+URxp4H9wCVoQ0QUqKRsHPrtwdrc
s2WHn5gYLn+FDk0/GqRHFL1pF1kt4541vAI+O7qHqKb3u3HI/mRnPUKdcsQ5JvPA/vx0Ei6EQKZc
IaEc5xhP3t1VoP7V6n2nCL3ElnO9iNmI31GGUZmiaW3P9tsreWjMct6hoqhOow7TbIXKz/0CpaWj
79tWpeMyMEtxQE2RIifZtQDy4ZxXMxGc1k/XfcLV1kFstgdb2p03WHRgwKiGtJ0ltIpipsZK742O
zXWYCOspTbm2tboLt/NJkHErxHJsbmR3ImH10AyJ+jsaywSAo4i9n4Wfab62vhGDf2+xc+ekaenY
d4y8FRtarqCgM8h2VLum7Ax1QQyDLRlgikNoAFGwPwFIJJ+jsAQvWh9t6z2PJIrTK5VK7OiCItYk
k8CFNDXa9XexMUVIzaC+loED9T6gOjnRjDTHJPlbjMklTzUCSvY1m/e84YilQXetNs1wSmlMIkkW
QVS9bnCjLWobeHeK63/zCp21zMnXCDxvGGTOlPjOekMuLhjqwbymFWBKRdIzy49zafxPKmJQGVNi
Di5ed3uJnt59E1OIhEXlXYEfSTi5LTlBo9i3CQfqSJ8uKwsTgbWygTlyFOoPUbmResc/WbY3oBT+
2vu1ijmBnNmL00F3z78L7Otio3MQ+4/cSb6dFuirAM3bI5qlkpDd8wGazvAuf6THM0BwOOOsiBB4
Dw+VGPRMf2vQX8uQ4L+HMv8rc+0wWyuZDyzyvXZ8SRded4qTHczlCpULcmHbMcem+vmJMHr9uv2P
byXSXSt6l4HCbwSSbB5MfYwMWuShptKMa5iql+30Sle+y3o7UOsmiIEOwUoUDDhwSz1fY6r16cfS
J2MT8ZTvqK8LzgzHuobH7SFrP99IcZxkW4d7W0FASzBCc5koCWR+gEMx4GcX7zklF6c/UK2a99dr
lZy5SfpvU7xPTdKvXnjxvZx3hCUiONmoPrJDaBO3bCKmrH92fO5iA6X+DiLJzynWG2SPcxQaPW74
sqatoDtXq13ok2JAfyU8vF+w3tSch4wVo4urI61O+SutiBLkAn6Ve5YlFcDctajil90990l9EiOG
MMz7vVnfuuwLYb7cdxgxb/eiu+ITAEm9dINatILxsRUQ6xGoz5aLhBcO4k42aj+pkMttyzsOVDTZ
J+0ijmHRxQOKlo0h0+Hz/wleFAg9+8x33v6bdDD0ZGdyetRCDQaRmLjqMdPG/Q+ichIN18hgGr4m
9fBGiFGQsueMQXETzKqqRBHlqf+KOw7gYGxaUTc0LtLHLI4zCYdWt6NNHN+nBgkElKJjgSrxKvZO
CQHwxl23UXT/R/2AvUqSPYKfu3Sxpjvh7iCTqSQCf81a2EOP2eP4MQmVMM6rAL209t7MPKnvU2O0
gqKsInMutOA4vUzfinAdzRE4oKepNIWEQDBJCbFtcu4Vi/nItBDMnfbTw3LbE26s+EWQcxqUXJvO
gRakowkvhTbbfsM3yy+b13ENb6t19ObDdYLl6VW13tG0dSz49kTdA0lvwpFm0zLPPPbjqnU1HIBY
4cL8QuxIpIzIP/Jq/MIFnSmI8lyXjD905bvrP/93YP8ECqhWHAw8P7V6VB2lcAw9uv2Fi/5Y7m1d
E3Xtol/3pwLOJJhKhxcq3KryNFUoEuzL13xKjD0Yg1iQXLqU/AvGVQCAwxwHAFp79sW0Aaz4CyHD
I1AbCB5fb8c1dbEiq7538+Y3bVrl6X3Y8Lt8N69vYtK+YsGPVPIPGer9wBiITdeC1VuBmCuqKCWb
JIsvJ2VMqDfUzDD8Cw1JMLrfq1bF+UnQg020ko0T1N4HII4buTH3O6RE8Svg4JwFNsoE9oaL6nVo
/gTNmZoIN6zFTDcq6+L5REonfMeCifAJ3yq3DhV/RnwP4pDGtX6ZIJ8qoSOi5cErUbzEijnzxoIS
WQVSASoAZaUBoAdiiZeKCpnJV8wY6lAMDjq9we1NVcvEwjTucvBh0nHK5nGNhDkSohgync7E9KK3
3iwwVwFA5a2gclqLzXv0tvAznMMepdfLpANxjYRthSfeWKWg7H3ZgfXLHR/SmoX8N7LHR/RBhKPo
zbWgPDLjLghUFD0zRXC4vgTe2y/Xc0p2u8ccwdAxVSnSel03dfU5KAGOOUfO95CV7GMQMkRYgZI/
z9a13W3EG0dGwLqqdSg1PEkXZy8AWIYXgO7MO5p6e4E4sg2QyAkiX042iwyI2R+Qf3F5ildauAog
IcwgMCwnvBLvv639g+hwoh6sd9ER4GWBKb5xulOj5JK+bFJVFqx1lr0yhFZW+9NkiTPlTn4GqrgP
FguHDzwOfbcTkRTzL8tIv5DRH8cTsC5UxIg3vdF7lrwGQ29cZ6suABh9XbH3cRpxIJxE+RHLlsW5
+3Qf0tKNKhfNZhcDH0RDaisYiOv0ZTMYrXa6ClLpoAzHGzMJosL4qnctjFyO1/rYqPcunWDQpjjz
JYpfRaITsI91LL9q9Qs2wUcCddmeQp96x5jjWQLmhccHpOA0GqHoPpt1lRJKjUvq1s2Iiyl+fMnV
SerbSUUPoVFJGlGXzPhTc7kvtHe0lwB6SiZaWl6s6OAWCqcm0v/efXKyf/a6jKxK128FynPaWjEJ
1trlTxh7qNO50zz6yzynj6haEzGGaaoNUIL+YeW1TmTEAIFreeLCmsCm5klEwSwE77LPTc5M6kPv
23IQN7rMVM4+/9MjLAHlBXmR4MVOeQMvOg7bgziQnLsADI7eD/D80oMo7H1i7VHwYjmG6kR8dV8b
ZSDJo+ukH+26t0e3zNf7SmnC/sRxUQSWLQeXPD++LDg7ci+KN6qCj7vNij0YfRVt8fh99VPdQuKU
dQqrUH6uiuepENZP7MlryixWGK5w3li2ujmAn8q+y6+qwksfn3c6vk6SRHy73+Jf0yL1G0XZEB0M
Na+IDZpksCUCqGcmTHkjOFmfpKcTXHjKDNeYewyuP7YHMPTWh+tWjVHRlEoIjKFqhs2ZoWwJKJJk
ZhNMUAUA+pnp2Ykz6ncuCdxiwDpuGWDVKbxtB0db0aSnLUSnofIT/vs2+r6rQdnVIROGpjaQFCGd
eEgOQAZqyL+/W9cRCmTOc/ceOaDTf1v55LRMwxMqrukKUO6vOniloka2N5O4krrq0OVCNwuFpLJ4
T0b04g4tkmgRbshQ4oyAwOD/Rjk+AAg/5vgLQf75C8mRbQQH0S2qyr5/MZ4yNZFmsuElsOylpjOS
Su8cFb9JakWQyW3PFVVN5kkiJw+zfpB7PQ31icQSZVAN+1LWlITG+ovN6zhcyDAHqovI6vbGFR0K
/ccapSIYxovvlcmjv5H7Gm2eXTto9U/HUX6f0Pnjn6JtQ/Wi10yUIwA8SwqapW0YPytdLL6EmiO7
1/Qgid/JJySatzqH2KkgeP+8QH2V6bNaEWMr4QqoG0fewpLUcRQ660L0XEhQZpBMghIcOXmXz9Jm
Y3giY5yC3e7tHUMH2A5hWhR6c88ocn75nOyVDEB9qK2O871l0+FGfe0mIo+Rn4HCcYKmDnYpkCWL
3LL/v7/XyblVlyVl7sVSh/lWNd2KNLDIxGTG3Wmbhorp1AjYelCTKL7D+av9pbI1LuUJOSAtxR6g
++kTSIIbxlltreO/l4E7qN7IRvqvCi9IRDfJp1xSxf/5wYRQC08I4TSME4UJcTk0pixvtv6YOt/p
4/bHLTOGDY9WOCg1+mb5tVwsqXmGaWRG1cQ5k357nMvLodlJqGA7p9rTTgFjPa1pU6oH2IOKVyvv
fxoCBnvccxco0uTcD2w9wVzvbZUILDw1f7YAIF7DBVIifo/UjBhAAI4f6F/PO2GmzSUdq2UBi8FZ
Zx19yeOkWTy6HQY+/53rPjcrKIsKEFQW7APqq6dbFRNHgAVdHn15WQ8R/lJ2ggBiPYDYW+lBRmUK
1H3yv6NfhXTLCAbsnMjeId+6hdz7utMI7o3CzR4nDYUo75quhGS6Eu8vQxZd3E+Qp1ECcCe+6P/4
CO6cNBDkpzFCvrewSrcFvGegYf9voSPZs438Yg5ArrpAYz8WDcqqNzMjTB2fTAx9eFu/U6w1CayR
3AYETQ1p6F+N+vdj5l8CV4co7DVi/4tHOogptonXqGMA48A8dv3vxfafKtaoZJtAopBSQ9wUhgR8
+yk5nDZZTTRsQvYW7iJVGWfXwrfsy1UcS/ngq7a8S8+74rOgTAXcjm7neOb+MvMfxBRPklD9xy9i
K40SRnLFtYNPffLWI+KbgRkDw8JpU4kzmw4dDTHHhsn5lnD+kimKtp8UqTXKPY2CL0nfiWwa90GF
4S5Sf+ntaAf7Nk1zkLDMd13R2t3tkzrcfmaNuYB8lS67O8JRdTfhdGdsAkBbrW1vi6N1uoqTE6+P
wE37RntGdKdGsLhgge0RbM68VCm8wn1vUiPhD7DTzpvSFe9yLdsklcgoR1yQzYysY8XwaGI3IAVi
prAEBSHePzi/oqq/1D0iEmxgTQt/l+4LQZQUX/XyRtNmGgtyxGRsqB8BE1yTAYOG0vOkSM0vkihk
To/9xtAcueoFRbAAYnCKL04HOqrMpG2F93QjwEEU6WvKiAWF368tIVm23WSYJDeFsCFyyKEa6R2c
Qekf3seRxSvCSRyz9N/n/l1KVlq6WBwt/Nc0SWXTe2QYfZi4Aa1EPvY3dRPpoLBj3EBONJK+CLll
8fASofcdUteIOnIzbVusFS9fm0sczzYU0uzkDQYM8nqqRfQ2AEaZ2he+63p+pqxy9Sy5sjHTRV9k
s4vHqdqL7VecERvDH3/ILJWsyt9YhSTJZqL19HVs1CTEgnVuGAEjSENa5LKPNh8z5Z8SpyDWNuBe
nNPgr+R4XvYALJGdIeSrpmXk+Glw6VBpE5M4BUXAvUoZlCF7Zwpx1ffFDfoSjcGkTokGOUS+PBz9
njh/tsozvzikAlkTFZcanXX0CSc/qNT8m+3Ht3qHPue0OXwQHlWXppcc27zlzmQ2phIZFh7kwZZk
NObafJigCw/ZGLhLL71vlnPMCr9ezWIcCU+hx9R1MUSUMEttou5XP/LhBxC0pLOf/AV0Ct0u10hQ
fVOojtzUqGfvVhCazfm4arRH38OaXDbAGM6pU2YOuTFyIohW1d8g9sGcUA/7ieMyHyaSiYBFoE9x
IYDWIra12d0adkcxGD3hr8G7ZEZTM2usrnyNzAJVbazVpJf+j9TXzg3ZDeH79flw+ClbTdGzcGA7
FUl1HRE7d/p+ghytAh8N0XoTYgE2z5P2GnstYL5SYICczeqOss60s3YZST9C9uq94MUkEBn07+0x
kpkZjTGejZyAqLZDjsCJ6Igwb+xo59VVmxDaYE4c7TYJBkKqLQ1GOPj8f/SSKSqNkOfOymR0p376
rmEOgnGJWo5JasuGEyEZGMn9x1g+70vR9vtRYdJ5rzCU/MA/AZ2FZKR+l3bok7PyD9V1y7gPfKTq
QYzbpfslECV+mWlKncpd0CRUAAN0aSNkclmjdeLSsT3MY3A+q146d6gBYBujdbwWJXnaq/Pup9ob
uYfxh8nEdU3MiVAHHZ+7Psdxu2FvMLiw3EKMc9BSq1+PrRJdkvpfwfYT7DxwmuvDdSILPDEI8XXH
hwRrmk+H8Dqq2VKcnYOc/8169ZBYiv6gu5jrQZwv9GH0Y1BqQi18Yd7BYodkz8GNOdsuFZsc+eRz
1Nmq5teOEqqusCFIWdXzFFSlVfaIXWC9CxkZy+vprjYzbDCZoO3cxfShr+feAGnRtZaJ+xwUyVne
CIQ0IFJJ4CjeXvhwuwvFbdQU8qMu5SUZ+76o+7TRuznm/4jTdoDUYNvd4PXmGuNRVmZ2MRTFQFVi
hArJlkeFrrg+oBsbVFnanJHDlR6lVZWBg5MPG51hrUIe0xdMEVeE1joaZDIRT77Q8R5p8zaRX3rN
GMu9A1/mjBAAyba8Yu65geBio4obx/CXHNXwp1Xzp7zcXWZ4AQuZL3ZBcfbn00yEJfwsBFFfi3Jy
egnkHiD3QhdRZMBT9bhDXdHskuP6uThe8e3J6JHJgDqbsxQ47YcjzuNttJ9OWgjOU7jdd9AzFCgh
zaqtt3jsYkf85DAly4BjQwwWD7iNqQ/6AuYB/96z9+cGULfE3QB+S9t1OFkNz71nqvNU2Z/1SQqY
lAKztL+GmqLFC6MBMFo1ZfPAe/EgaiQA4No15rxTb2MUjc6Kbxl7WeoUbK/0yc0wrFUN6WAw+wpj
rNqt3GTDW55FplyV/ZauLW2ZCABshh6Kr5XjplGyM904SH4DvUfcrPW3yjizK9AbkKUE5mMNXDBt
Rr3oBanzU4T99w45ben1imxVP575OgAnABSPJ5VkhJv9T1PfMXJ4leYP3DCNVbmrriFvpAYb6UcQ
eZT4oFiwUalIexuCBfZV1yo8KkjdXOzEI00A3tSda7IA63FFk/Dq512zCo+gDVlSK/lkg6Fyo6Mg
PI01iRzhNzhR7IgT3aJ0xFHJZmmaFygsoIlTAETbdY3aWb82u16rJlQZk4mCLMg1l61n+BwESg4n
AjzDN68RJ93U7mKCavdbZ0ykw/Ln4jpaVyGDLyjYpoItXDw/m00/yr8AAoiB1FqRKthR9rTGylV2
vvy4scFtlrb5+cYi+bVkJWCR9poU6q2KgrMiL1iT5Q8wXPbw8PAEQdWXD+9jduexmusoRmoTwlyb
/o6PWFriBmbtGtU0rtt2il+TUpdMDzNNiw/9v9OiO9OUtfcKqShu9tk4n4xAKqzGcEsrG/JiMKr6
hN9xtwJGFQT6ydZjaMsulWH8tOmc2JUAZ90VrWtowPjgk/Zxvj+ujH/mqO4502XDcURsMkwcUW8M
F05zDa9RTk666p/Bms04EtqDxeE2o4XOvQ+7ahnTLCsUnf+iYWSzs2W4xpHn06mw4uyS0h2BWNxp
ij8K1MNpWf6H2jxBYtsQFVs8gpS8HkclXhUYI8qMEtSv4ONvESKwQtVsiwlUpwwNCAUGVbvMZZBI
lkw3AGmoVQCIuzHy/mdYs/oq8J+HeErifk+qiDfeeuzuz1czdHRFo+PuJgQLyBw4arky2hTzC1Fx
lWkSCrH4hgoUanhKTxKs2G79UfSQqNpVCwnhyId3PRMK2b/tA1cUNS6VcIVVxRYeCdkT+OjNmhNQ
Ezqb1nxSnBsfNGXX1M612ytlZOqUowQkJ+OZq4wkhrqSjEMeRkNR1i/To5FuzOudcSIFk++8U+tM
Mi+LhY/1f+RReKsbLkWK//Kk2e5d0Rf6e5W603X/LsnfoKa+DzHAgNWcIfryMIxo1mm3xP9VJxtg
wNU9w1sHVVI7jYoYDaHqutRZrpDEYEm4Of3OVOl4Ds1dITTFIuvK28CRgCwpfGfhaNMTCQQYMFAz
iyT8qTRJPt4O+jS4CdAlVB+u4h0FwkHy6LFydMJBZyjBv1tR8kxekXUFVSB6oOhOpMq9Jt2HpZPp
gqOw+il/rw6N+VznHlaCSohd3UGP/0Ors/pZih0tT9B5ktDqovhPmvhlUf+7v3GYAAh0NlXHV1v3
YBmZOFreuaUy7H0EvmSOkJoMAI1xKThovyq0+Eps7OHRwuxq3RvYdelLyBOi3dMvQgcHbWfn7hwD
Sf4m6zotWLnsb624s3vIfWTDY5ktZhiUx4dgcrF3EBTQbaYO7GfRxlCY8yUFj8P1m+/pgJHl+VtA
UiiwXncDbtA/Fm0hRXCyjT4HpHyOuai7RNCl+BICVTuF+z7+cdeTda3hNZaLSLsVzcHY6n286mC7
F+nO7MyXsq7BwaLxmkYG+cpfyzL8+XF3pHDkH0Gky7m/KIKDvSLMjYkqE7SWkRiuNDQNX1u6WJ+n
BfJkTQ0p43mQ33d6yNzbITaR7BwxU0l77EWOOnd7+R4APHeQ8cUMZ6wdEfP7NBEFhbMNbu4FrdrI
AqmdoOz2CyKrn2n1a6/knuT3X7uXPVTa4jehul34TKZUfXov5ju2jjSHZypFIL3b2f5WRUr9EZA8
zf4y5xYvtNzHM3es/To59ToyfN4PP4/K7XN8Ay9wtakKEyCJXL2yuhzlteTLXHMphgm+0RwoiGuh
4Hem4my2aUV+6vUDVfwp8rg5y93HpJyucWXcBeTb4H6xlbmkMlFWfjyy/r2rb3KPm3pq5PFicr3T
YwSg71B07eokLQWb1W1Mz4CqPEcsDnAseDwlDZAADPqD5/z4YAhOKA/4dlacw5lPuweqEI3nSbGj
gwAFdMB/0OVW/WwsLVt5AGGNhkkUYf6xzoQ2AQwhu9lu62mE1QOnVcgowf0tS0xvcUukmi5Z1a9k
pWxv1oyvDtm71s1Z0kfJbiezagyLLrCpJvbsEYIMD9I4tIi/r3S/hEMGmNaPZMjkKeHwURtGKNJ4
oRX0v7LL6xK0Gw1ndZdyj64HHz1Y+QzzwESEMTd4UVN7XkEe6DGak4BMnILTx7hx2kN/e9D0vjoz
8MuGABkz/m03T0UjMsWcz0juCIbOGPZaQnEAfOvevlVupQBByB2ElDDaMhZPa8wjbrLfdgPTOGec
aM/wz7IKqUvhQnACPNzzFu/9tXa6MNpFfQ9IADaMnQzdTPsJ8gmxVzAIcgb9k/JPDt7e205fwJQA
TIEkDOEBt/hGwlpLOhFtEQL7u0eC1rcom/pmX+a4UNt5VENDHboPIns359aeR84WAVC87WiOFRjM
LULLeCGZm0s2RrGRiC0IzZHr1G2ht2oG5dHuD7o7e87vzxOFimALqYLUWqCF+E0sCg1brBSnmasI
WiAe3mZHcSTQY98IAxsfYghBL9I/9GnZS8LVfgM4QfKRY7B1cTGR3vD/A44KxwS6Tm1yKPaPcf9t
kAZV1lcriU4/axxfFCdbK3w3441/B+lj+uvXKy/pGujM2dqmvVTmdC08hPm/hDTzJGOh4ey5W5lG
tl/Uf44W8exmW0R9LQRob/+HKqxtcxpHsKGA4Hv7UeyoRMnBnjdP128ChDYHsKOgBlvs3Ce6KAyv
FwmDQNQeHVwxcNJU5QtbshACLyTeIWv3h7a2e4LE6pAg0VBCuzWa774neAyCfjToOPjnKEm6mqNZ
Oa28WIbmSBUdu4DJODL74vAto1TpdMZgXsWD+yNsKAG+sf+u0vsNuXAZl2NP9ankxJdAnNwDohb1
0HKKz/LyedYCG0GVKBFhzrpNTAieAxZKgMOh7VwXXPLuKYVpFIv8qs2/SMa28r/N9QKCaLVHnSJ7
cqjjDt0DTYYRznk0JuJ5Yrg8svVb/OuQ5C/LTlYtungxkRhR8yUkOovaSq6cIUdeDdPDwwZGYAck
19WbiI7f/qKIaf82JjiMc5Xym+Zkbemi+qDdIfN6Ct+ugizzUJfeDNL+sShIRzhbvq6vtwS/AkSp
01Nhm59FbB0ctm4rvucX6xYszrJk9QGBEjMMGj5KtIGxqP3a+wfX8FL9zSBJtmFcK9SfdXBnf4l5
+/xMltA8zNGh0OL3zXW3VNForU9xoUJR++kz6RsAL1UEswBTgHsoUT8CGy02Avlav0qrNp4Dg+qh
S35Lqoct8ASuPHbZqkiu1iXgOHYy0LRwxbbJGQLkNXc4ROaPte+WYeoKWHDJmGLeAZavR56AZeOA
RkIa5U0F4Dp/9/rQS2SEeQ/wWgqvGUjS33gJ0ghOJl0e4w2y7flEggRAlhe0mvJ5inRduA4zBc+y
sJ7VBZ3K3MI5i4xDem0erSUsjWVhu47Nhsd2O0/ILX7Ujdug5WGVfoAPYvoxfE5RJHhK5LI/IDst
wThmcw6JIVBNSQFdCmEfXmOf2st0S/Abt2xm7ttLaGweNoqZJDemEtQTHKNTDBHBnfDuo9sepSLb
YufwH3vUD88JgTDcVbr5kxpk/5QHzX25F32SVr6nBibZLvB/cvWwYgA31/36QSWgTiWB6tZod09p
Byt2oFLS3WXxxr8Ukr1+j2eC5/9iNU83C+xfbTA7VMVGeJN+N7DtPP0knQur2RFcB8wxKU5UV4hJ
wBicecL5SLooc4Tbq/ZbRJHFxwRJ75uWCZUgIQeNIFVp2zTaUxbdPq+Wqn/8Go3KeM9BfrWhikXl
vi7Eb9QW8jYrH4p9L72+790Gyeli2jZEFiTqnoC5sjr9xQRcueMHbTHQB6wuff4YC+ffX5BtbcLb
JAp2VtbnUQzmEbOXtIgsM5h64jIqnFZRXw6luyfmU2U3Wm2yXkYoNDjdgLUXDymdYQEXDcPE7NG/
1AfYxMLvtesPOhmkrjXIskcNBFdOZOHcDUZEFyLRbTHMaG3CwcnsKkObd8N4AHENgPuVw9T+Cs6H
+xN8zKPg2/BA4bEfAnEGlH0M3gD118AZNEvsJuiWi7ptuihhZgdM1gpfgk34qkSWLkKUtJPYzYZ8
S3NkY/DBk4rXNjVGLT0wmeRTsaRNvxxEB85NFXTOltO8wVhRbxxdqBAvTraIPBctpPDzMb4lJMyB
ShEfvgzEY3jD2Fw4OS8CiHiyfGROO3iU/a5d1mkT68n4/ylCc00Bzn7+vGfl3oeX7sPu858LBO1Y
IJP8/aZcgfSmsegNSigs32neODJ8g9rh7OfbkF1pQdg9eOOuRnDJwBiddqUStUUYpVFo5z9GigXJ
x9Lv3oI9ZBlFAiddUIJfXr5Ne0nOq+THriml4gEgC9YKo1LJO+z2x2/64He1kFuyv/3GLwQRleUv
rlXanDjWOrl55a68L0i7JRwjoHmrEKjYVxC6NyfZ9Pc4+Pk7hbdAwIbmTi0v02SwG9UcqO+/KbVy
kJx0KCr6sY+P8pkS+Su8eIynjRalmMJZDYrN/TiXQ687Iqd0ZKCqHS6IPYY7D44fprKuE+/79VMZ
CezHqZyqFhVJa+ELmXXlZYNoMn1wUd5eo+8GIrpw1WuZShZfo5yWneh6RqKyF58wOW3a9JrIqcLW
EoQUKON1mQK3Sn+ZpJczU5cYyWM3XYQ001UlUPvhkaoBpLtdWJ7ciXB/FSZwm6PcsPe69DxG6T5P
Xx89JT4ts0Hk2HxyXD1YRWv2EujyneQoDItrccQHUowb0pdRbFutudixkhNwCgqJ2jb569tPZl/c
QiJ/hzqzD9OPa0coR/B/yiTIhyPAUScJO2lrs4xecXR0Fkx75px9XEMIaWyrisLtoskxeXYEcdJm
7HoU6njCcxTHYF/hGQsoE9b8pE23F9TzvnCWiHhhVSv/Rn2PWuWP9cnLWLFvpV+t9SPG/Uw8x+Qy
vlO7wrFmV0cn3oB73sAd0jscIdkQUF4gD6Vg3zquNPoELKyl1D9vdSNVelWiDGjnjDMXgLSqcnSa
RjCVCHXxw2765GnGMqnrLUf4y6GuyJ+MU9pzW+h0LRfqh2eRpkiTg0gAl/rr97G1Fq/LKzoymojX
py+vrBUQrzXdQKYdr5H0we2TkU0gWdHy/6Y9d3U+3QtcqUPS/g0/j8WLySjLmaAbYtnpwUhkfUY9
BtyO2DsnRhNBC5W1bTFEh+sbmWG4TB9ug7+9GgGfcjF0HbnZ0hSzIO+SDrsRkhqiCcWkE8BY5Dk9
mR49gm5tcOOicqJM3evehiI/S9XEdNExXdpByBTIA4L/PoKKADnFBIxiTNWjzpySwMnbGaeaxASB
1gXxxu4LconBqOZ6KtbNn3a2AZWpWrv5aUPUXfN0L7WQkP247tHocQbVbrG2mOGNy5M0qEa0vh/5
jZn5bzGhjZHhB7vjSZxjkL9ErT03JgPDQq/VnBoVRS7BtpGk6DBkDs7zwnr4veXd5m3oN7w1SmtH
nROsxJWN90y03DmwFmb/Dm806iBr7uavD0s4jM10a2ejIV4vWNNDxlY7Tei2dG7I1kbqx1PkBz9b
vZyaDKoJ7eGDVm5riCwc82h1QIUEQ+Kdcp6p8T+VycpUQTFhxg4wu+cWUYB7IYh3K0NxkRfEsCo3
YRj498bQnPPSmYSfdDMqgUXFvj7FHNKtTSucyeASnIdQM/UCLCK5kYv+QMx659TacnNWNP7jZIy/
jmBo5SdQD3PS/whWRPXozWqESkQU4S6zt2+jVeFSmiCSx+O2VNMTeZmn0Oye7Y8MpRHvT9ceUuA6
chgPg73IvWKyEmGUI8/mnSS8cceAP6KuiQkfjdZgBBlnjBkgZLgdAQeAi26tu/4Ugd6Fp1fZyA67
5bMMwA1iBgELgA/1gJULo0sdEE151aLxt51md2D5bIJ1AIXZ/ut5wwDwb6JR608wS2flXQxp/rI/
9SfAl0pjpDUr9TbbrR5F0DeREdvTRx0bsp/2IEAPlpruIBcvX7a2kokMOWIfqPAX/TWFHdR90bOC
INp+vSRzCsYkHvUvQXfMN8dS50G3s2jHX0Hp64CbdZPfJ6g3uZ+7oAyZ4DNQQQrDOFQBpUHFh4vI
PC4ztnNB6ot0z6VexkwKFoytGrJgVCZiMpvJFUfo2O1b408NDlRo92xiK1Ju4kIA/RDTV+eJyNjl
YqsGsXyH1/na6nwrCU0NqoWiw51SXlnL0yVOoAcvkkn+IYJ6YBzPQnVF39ULBR3F7aQelAbDmLew
E6KZvP3muD2vp5p4ksBwgmr6BVd2PHUKXRKoRW9YTGcr3qsQRvzTS+Dl7lhlAaEobgXPQ4UuqqfJ
CwPQyQrVYLNhaX4dDhL5f5BythET8706BiIMkgbvZ6dv+GYDahZuHFhP0/bP41r3BZSvEm/CE0vs
bJop0HUozfduDmx1AP9o9gWvvPKIKaL1c9nsUCakclvjxfoYT4QaFp//f0ZKhH//AEBo6bytgMy8
HMQnR1lepe70ARtnk/U9bpGq/u6ruETYvm6qUEXS18Vl9yTpyZhoAE/1E6MiEdbRGwPi+cQzdIny
9xSFYrJi+hMygM+Hk2mw5oGoD3VnPrO1r9KVYQOdr/wWRDT3ozjJwDNv9Td7WEdfmstmxy527JjN
Z7v/BHIMhPaZMHUqXnbfb2FQWmzcndnswao/CdfPR8pCiQwVX3me3qlDvWY6nP/0Mvwp4UHgKDgl
oiD0e6czFG6FSvWr4VLoyiBRRjk21tUFIkZLeRpKotWh95OhqSbkofsTjaWkhE1umCRi12uhcM0U
R9QqKBvwTffV3NjaVPhFTBQ+ATClEVgH+CZ03ffwMiXNZ950PCEzIVt610HbtIODqdTKkuy8V4Gx
gHtMz/GbwFBsEFrXjr0ziJDUohHZ46LpNO/wccE8cuvVkc7MvUQZYKkdOfXOoC6S8JXAQ8sPToh/
d3eU5iHCuLwG6zXgLJUxXUWDe0TWnwEQz+fJJR5ZYw6ZmXSRjTwPsm6t+XuSnUAUwfPFCabSCwJx
eYllSILvKhM668bOhSnVVM35LBjcu9Zp/D7J6cDCXxQWgmo/NHNH2NRNBzQDEvhakIPDfjPiRj57
7aFD1xSX8Y28iRjMVqAWqmeb+P1E3cfgUcGE6rS1mnTLtlf7tRSC5frhi/9U9ZEIETES1yd02a3V
Soeg7uL+GRLfz7k+grQEFkbe1NLbEVX9sUldsFBylJp/lqa2rb1C+0bZbVNsjYVMXNT0Fx8rMTMF
6343Iv1UAHnLDrJhBoAE0VtLsOiPtdA4iE5LUJQReBNnrbZeT9btOsOLaNMqtD0Y33fkNtbgYNsw
Mog7icw7/vqzw4siY7hMJlwaOU/yx9nuJrvScMzQSvaHZhbVcZEJBEla5Q25n8MZ+lFPjoXgXFVh
MeIV2NccIn1zID/JTTiZW0V/IKoyGyaPNBfVX7DHK1nAthnYaaGk099U6anQwCw399WZe/lHV3HV
kqZ0e7p3E5ZRi6B31W1eVOEB1lwbXBiJ/KTMiiJ4V49GR+bhe/s26z7i/Y4AtohlvCvYRjHyJusr
9wSm/+KhA0g/M98L55m82/92LD9a3EoEVJ6EhI6MvXP9x7553Yr7EEj+Cqwku1G/ou2+b0hTnBHK
kMLf9y0dcLZqXge1GlFd5PqSNUYZLLNmyGAXKrJ8huZA7w51UUenA+DAW+UPpYwRGs3EbcDIJt+2
nKmNg5D2ktVkRiCcNghqiiOMJ/e5gLX0gC5SLIWqsSEjkupk79MN3+KfZW/RvPT+q8ykbYOJ6q+9
zIbUvOpE0+94chycvdXD5dXbazX3nNqu/Lx11XaHWDmQN2SsXJk2wIQnSF3p3NUyhjQC4qzNN8oS
uGxi7KW4QlyiAiB1FJLPizmALCmZSvJsz81tftvQnmwDgfMLPtzsgk7AfTGk3hQ3cbkc7M7SSvI5
Ro6EwS/T6BRvMWhS+MytASATFOWPDPSESTXCahv9hu/jbBzaXCkJZRSy+E6TYQQdy+Y6f+3WVEh0
OXDOcYXXOHhGDBJJ//id21WIZ9hYJFyrhWElcVEtgzAcWbL2ufXbf9Y8pl+3Mky8k0Wv87F7xPiq
7KEnzxdrFVGfILolXvoOH+9ZmQdJLlkOCUj/AeDT8xrrKOA0D3C2icVR1WTS+5XwSKVy1qsLhY9r
xoJYpTT9tDvDROGowZecBARyGtKP1Mk6qg27lybADWdNKcI8o+Ig2OpOVlO8CAmEB1J9tJpzZkYd
Qzieev/OWQMH8EJNx5nuocnZ0AojJcrlRBorlnVI6XxuT8GJCmsGvy2+gsBHI+Gd8Tbe87kXRl4e
lZkQyWL++Afx6//VnagHRwOb0mIeCRyegX8pZAdWtFt+P4qteSvh/2qKLNouTij0++xMQoYiprOh
jnBqqBhoGS8M+cN9RWETcOWDcy56GCDQ52mELmKQHtYYCXifsGXfwg++kSFZ+XpaSt8EkadBd2cM
w7bdYN6QzYoINOH166VlO3dKNB7ggf0LeVP48oVS5ri2dDC9bo8MAZ98dS5GMB289d2Kf8W07OLh
oUBZaF6vO1bJMqkH7kOZT1cgNd9OBLQceYWGnhRn3TxIMP5HpeM+e0nxWxF7v1lwAYmjrD2twiag
gCgWwRqdq2m+M/jlbi30X43ANBpWX4tCKjUNtQqhNgPOIv8BiipT56XqEv/0bcmpGOpUbs866pxl
U0CVQgEoNIXFe7SxDIplHFSIKw7zF62pCiv4EvvpMgLkeUiDAmZ+8poqFI19PkvAjKytHYknHYx7
HXMI7ql+m27aNKWr1UK4DbtTQ3W5+6mRqTsIGVF74ZFq7SL5eawNT33scbqACI4KX0YIqmXrzRk8
9ox3jEQ+T0O8VFIl21RWP+cR71C6LCWzUuQyIYb0NYvaIdeBQria8usyRo4wkVptPIFRCzACkWt6
9uEs+/mcd7jEM84qMvblPL2ODmv2G87wAte/CpwrkrXvuPOxiqhV/SG0/w0XEP87xk3L1DXuv9TG
65A+UsSSQytzYlwiCOpl/8mPvTGJBfnJ1ua83wWA2Hoh/g4eakYbUBo99nnuHDrt0aPBwYzMzSso
SINCDtKOkWK0yJb8pONigB1EcwS0PamCCdnA7ZW7zPgBnSy+UaEe0YkXu7JSznFlTBv8jBPpW1dn
qv5b1RzaC31OFEnJZeGHTa9xfyd9rl6hh0YMLsYxaVosgHsVuDaGO7uZmgdLDWRJjhVmoPTQJYcs
uu+WrMeznodsVMVBTiN5dplRLdIQXIB4AV4IOjJOapr+dZAqb2urqBO8EGn5qvrBoQBULvRY1q8o
ksqhD7Tmux/38J84R4DwkBqjhjEsQvGeQCgrzeIbY1dl5z3T9q3eegvVU8VoNPhxKfnKie8P9Wrc
BiZ5/Msv1ywewTnszJiBvGj4QURm9ZnEyF2zWLff4TjFgfQqczvh+CRfYzJcNTJkM/OxLL8Cdt7Q
wGGCeU17JeDZTg77ApJveitOvYA1h7cO47v5uJHE/UWzOSI7C/tBvU+wIbOLrX3spXiyu8HjTefy
jIRUkt5dWez+n4xmPPWobXovP61eoI2FLEMO0zaJQfdi7GPtMA1kbOSu1Oel5MMtW6ezjQAx2ugU
A1RZdRWJKPumCnQR7/uIx1ICtLNrONBVLdpG3xOeVR2gbddup5JQYLD2WS1AwAwgtAy9+8t+jLlj
0JkJd2UrsOszLNTicyYEnSASDNuZDDGzeqI/dx64wxT2w5a0XB0F0OVv9TXW4s81Jlg71bnBompD
Xd/vpOJZDZqyaSAQVMj92Xf1247Z5ilXV9AiHldA+FhL3YEfM8IX7lv4rPITmDBMzXjuKDzU54uU
0R9Le/zygosAoOlPQmQr60wHzvLQjOqvep2JaQqTJQ0LRdDMwtvREG6sxAqRDf/QMgQWkEq2xvcl
YWrI7kPmvblet7fBleLOiKiboejmcy8q6KFOUF2eixpZCpoSYuuccoQTjUjqPYeQ2QbmRkoVBBVi
x4FvOAS69pulz5YRRZU/fahWQJiWlEg/Wh+lt8cT6tprsDeLRl+Ch62LAm8SQwGRT5zUY21dXZBh
ZG2TPoUA/ZuClE0cJ0X0bUcI31ybkxQnku4ahx/enN9z099y5nN8JUQc6SRG+toUXcog8/y/GzD1
tH45F8KWOa+MAzJXeELJMrF12L7upjWreCJHTTpraxfzfjpeFTEU6W4dhvz0f32FjFOZHCBDllFe
cRxofzVA+4Ykd/R2YFCGWrhUjiVxAkQ+/i03yIp/bIwdrNgc75EkdQ6sfGwUbhCDI9NGvjSb8FFZ
typdScesDnJ5r6Q0sXRx7EHieRfC+who4NFvJIUPlsteiHuOd2cbr9ihmk8QGlCV1DEzoPBEJHpM
WR5o+d3FlWSCAhEZSN2hD+pOkzh+tQAdmos7t1HfqvqfjnUrkEw3wlzNAUrrnRFfpbUJzDH3TezU
etlzHkJb+Vy7P5oGVRFJg/cNg0GkjkPhio9O5K7vaaPYddHGKrywRNbIZhLSrXUs7w1NSkEGtP3n
W7j6UnIYOrDP9gzYM4LXqvctE2ZLuK3vcBKn1Lw3S/4yqR5Kp4nPqcPCT89O580HYgNUsirLOBpF
aF/V7eaxRANqb3g8s7KbJFBW2xIvDNEFME13QH8pVZGZ+o9LKsugokvCdp18rz8mGlcCXjdWX6Ac
QoMhYYr59/3ehcxtAegw2HbKdFOOh24XxUgm28kITGNMLrxDR+KcSt22C6dkoJPw0I/wlWLsJ6VT
V/jdBEvSG36qa/IhqI+q9m3C1lnKSAVKA3rldDAil7FBCcS8xaDh/cOiGlhXK1uZnIuq6eGH2f5I
OXY4Md/hFUtjw6BTSLulsMAyapEgg+1cX6TPJZaORZOi32fc4aqs1E7bXPxuDXhDh3FBpIlDStgj
HuYtERpK+gEudqrxcrju9QjpUfiGU1vRLhJUvtIH5ZzIX+VFhFQ9eHZgKv9YQlx62Y7B4qUz4Yex
rulRWSZsdxROrJggLSp2b2SXS+7y1A6OAR7kGmj6QZEycntPq35yw61UwFYQq2AA4HuE4r492Baa
xPqjxKrzHxgehwu0z4jStmbCbougqJOlS9LUEbioRKQj8pjUFGAJg/Ri5/4jHEFOBmWhMOG28YEA
beTn0KcMBAIJgRwJqeeK5mLPZXlMUEpStS9AQAX3AUvOmM9Poi7BpiFr/JGQWxj70RxPnswD6L29
N5hq4vYCvJzxDZGOwn92O9YRDXmTg+z81sxXMRctD1BFGLaXJtvQs7SfekpZ9b7+SOMcLEf5iXxY
k6EqaK6ylyjPWk7CMpxgT4x3tRD7hddn0PhvFRBRjYHtbMk1Os0V1v+ye1zNdD3rL6JQOlb6Eyd1
n+thATk04afGXoVYWyAZzqV7IqPsU977cMnVlJeYBN0tl3TP7P77K6TeVivNpPOUU+bYoiHjrUJT
WJZ8biUkkMz+nHmPq4ZF8YYZ7p/M7kuT/cnLp5Sq2JKPe8dpImASCoZTxbTMl5SwBxEW4z4wGSNh
fY5a7wwjpk+ak0CLFyKZOuVYCoHw5LcrrCO1zHSGGPvLxlpdPliiqcM9AY6xvZSlsMzHSRPFsNJu
2GDR+5M99iQGiDgAJ3zZrkWqOCeiyYZ4jGq7QBSb0sr/tpm7w9DT2bGIXpDLAyL8+mFTLPSSnV30
hecuE2tqgYOUK2CM6eXXS7BmThzjI1aFFzQx/W5bjSbF/8ONAbMyb+W3yIkx0T0eeYMLWdytmUcX
mUz6PG0YasF9o05m6bLH3KpwOGmP5ONhj+e9dB351NvS7Xfw8WAwhgNhGu/l9Vd7lq3DrWB/XXoA
bulm1x43tjVz+aKPqp5yTv79+0Cw/QZdFHSobY4kld2ZIEX4IOLLcvTxvzAB/sMj6h6wkZuWFOLv
Q07JkptvBQ/UNpyGPSBiG49f3Qlw6PpdCuM5jSZK4+LloZDcZFKirW8QNdQzluX0V3K2VJ3k5CIi
9r7UgG42qSysVp8r8LMSGRit/YjwdiRIavs9ltPXXIC0IdWiWmF7XKIox+NzMyKzjUFOL99yBtsc
pfAdiiI3bFNls63cmuCl6ZC5G0A3R1sos2TVIman2aaNza8Wm1zwKdXuHCF2rvtrcH4JhBxlidUr
/2H00zFdM8PgJQiVKSBFrelgpehqeE4IAn3mh7urenx/n/zI9JO9vUtliPTNw+ATbZV3hER7bynd
AiBtVDCv/Laxe2QwG+MiVlG9uya+X1PAu09TRO+E+tWe0O1frl68e+CvcpBxe3LWFi7iLIE4Vs6m
jK330SGCTfa9U1PkCjjP1F/pWO/lsfMl9kLr62Rv6J/LA9JRmY3LvY207uL0zboiJz+JTSYVv1fJ
XJw2jKLy/XWioLqZP15FXmWJHkUPOW3yboJ3PFxDu2rGn2Pufu3cwRkZ/xHhI6LwoU+uTGG6dBd8
+LPDdoE01r1mw2WKQKRpDrqsK0u1ravl1X53acp9FpiKWhJZ8ISfXWd6pqGFY1oXBE0uSgOa5z4u
nsiCNJ0q6hDae20qMoJJdyfhVe8coiDRFDCfIWmD985pDBIdHvKlrwBU7WD+m7J1W6wAdWCpF1NO
20idHo2jx64V4PR0/VYeBlszLSOOX60k1N/0DXH5cAYkCw9mmw1np51M/o7tot6/d+t+3GBhr6KM
EcdC9Q+4Mp51KRYsh7gV64yzYeEff3yrvtnXJapScUfHwoiWZoeQ3bKo2Q/sDIKHB9GLjG/zJPph
irH3rxad/tUHq6rufRyEAIhL0V/LGQcaUcu9R7BpFsLBikn1E/4HVx9eC2pcMqBgy4/DH2IcGZyr
jOJ3YEmYqTWlfsO6jdUos3MX1a0rQPoifncwCvdtKx4nWMG22M9GjBvufcdxMu36gljlH1qJ7kaZ
PWWpjp/KBf28ABOD1QhrgGAwmQ9Gh/jy2YBJrPYa5cEVhPryrUNCrW+cvBHcZtx14/j0YC9K6Mz5
BGzibN7iCjf6d9N1bpc8GaCPgVVjSmQ0X+qVn7GMHE9RfG5tvFyyHOg81Y26xJHPaX8vidqnP0aO
yoDy8cVzrrXRiEC/j5cCTh9X+xcftrcWV1X5G2h76us2qrC/5OfHRRAqZkYWop7UKXdeW72vOHn7
nAJiHiLeeinUPur08fW2utkXNYY3IqIBEJOdgmbayMRc+hTO42gDfrxiMd00asI7LH+XoycywHIE
zB1/2+oK1VCqg/ykyhRmxPD8Ibc5a3TiIsnMTeDDwDzKv6iH91uss2huSWxy3XfE0rqARJ2FH7za
EVVcLtLp0mvaSlEUha1lB9xDxhaKnOYBKr2uM6p9x0ok7JhgKv50f2bmQUWl1a0Yix7g03nDFcI4
+zSyRDfiyM48GJXGqJ24jp3NH7rmsgGLtFbEANHCy5aP+feN9bXzM17LTj/lqyLAYaLY1uf1gnhU
QcWoYpEevmu3d2ec49x8IoI3PzQunNYK+qF5OF3Cdwgn9vgqVd+2wPrQW7lmMOzWoEuXrtT8ApcQ
IO8enMA+79O8wdRHz+E32JL7qHpg1xlBhkxDR5ocWYCLuC9JaPA2llBvIf7/atDswvenYUeWVMPi
SBtQ3ibFhUKRDHvLXIsgwPmSVEp7k2oBSUXB+kkciQ9oMGNxrmix1DtboKuSpnMBhF3oK84V9Uk8
IbwuaazhDgg0M2sUZwgHpGm4l2Mqtjum/q0oJNMtfNmAC2nMHToAOXH66TfBGYaYzue2R0HN9fem
W0nsaKeh1VQPmWVMFu8rhEL6gm0/SncANbV433aedTdiCocRTu50WEMoCOEnOj9YOozlpWmB+QWn
IatZvD0cjNnXah+y19MuVM33mWUekXzry9YixpzW/FPu3Z6DUHKPU905u5qYlxK79o8VO26o5Vmi
0av4idOLioCLgONjOYZ8q/uML7ou8hC1veENFctMqESLrxZPviIZBxDxYFdWVg5/i6zheqblTiKH
t0IP7z5/wmuj3rwTgU2af63ZfwPbg4P+i4shET4Ya47YmRp16lu6+dKHpuDPTFdiR+oUvYXEZuZN
dWpJgGOoU/xh5WTynKnyK139hx/n/ef8I3XR34NrPd4DjWCApC3T3DeBed1I546dTJR8tsxO7SRb
bA8AwTn+d8DKV6m6qz2rRVPmwyfZ1ZNv1v8cjEXd7EDjfnKPfmzG9FDFKS/PafvTVS8aA6JOnygh
3N1rT+VQuqEd2fdpFgjFGW0IRTu8spTbOBeyNyydFVKyixDJXxSjytARWNe3xbVhtn5VEt1sNsX2
98TLJuCx6CqPFp4cAa5Yimq7BN332qKRylOy934ARzHMnlVkqhptqrV+uUSF1NrvWHuOPZT7uz1z
b1BwFlcBn0Yqj2XezhTqu9g3Ng+mKdARA4Zgp7lBrtC8/4ZHWRzMa4jAhLPV1gtwpurDAGif4Xsi
C7wtnjkiBLeW6TUdwdYuu+KVNUBVQdpwe4lFrsWOW5t89ybdNRYxmioObabeS8xK7Em1qVWhNfLM
No81WtRLHw/6lg/JfVquICKwA5rQCuoj51SjdIqPj5TDGPLllzaRjPxSMiDOmpif1lm+X5HEjIRv
yKJrbyAOwMfZvLv6wegrkk9AEMyNxX9DhVASjOl/oWTmia9QLHvmoNmVqzGXPzcDi9xqxD9pFEyZ
qXMFEvALqSsWaNZxNuFPTXxP56RpeHjpoSHUmBOrKx/lbl8hP+Dn0SOE2Mdg3FvyWUdGKJeC2Obh
6JG2T5QhkS8LYbOFt++rDomHrLnz65WltUmcJ4hV/RZdlRFU6Qk140TH1a8+gRWoEWB4scVmDzkA
rm/nPZgtdDd680NTB2e0k9bN7aNxLNWbTDx6aLBteZQErWAru7IrD75SnNjvIBmFdwQ/Viwgynxw
+7ro5iQpp9U1oGMKnkzb1aSXBYBR/UKUdzpPnqeGun1Di0DgYP0F/mV9Ltl2E66uqHCKnD8mFto/
IVOKMguuckRfFtPGjiJCKUHKGvdmwoW5Gcx/TbYiljfMP/EBqr8ntm395WCIu52HCDLrLbsQslk0
869JYnQQv3eMMZNgNitqzBrHCVXRexkKySas2vvmRW/jE14dZzmTq5dQSQZLuE8k7y7WMgtQV+ZS
+LXl6ANHd3/Cz8CAI2JZLt5+seK6uXbmGzci0XZ5zZD25jWpFJFVW9PaOSve9udCw8RQX7kn7c/r
4Ckz1EnkJRrDeiDbiZxMlnuVePXgddZ9aDZiiLtfT5rnu+WJWIWkRygMxNSQp3e9nS8nJt6LLh0W
S5k+WOCTL6KCWtqMTHzF0uZkc2sE7L9G+h2SfmpOY+aWjXOeed+cjMQNt1zGZBk6LAXRAS07V4uk
TJITHJhSacotTtplf204HWXqPgcohFtyNuXFMz/fEIhIwXQvb5UiZgZKkYqWoI9OcZNhppK8xFkW
TwfF/fpB3kdjTvgRKcsR+D/mmaDwrd+ZRvY+adaSgMs1Oc0yfMTTwvuXkoaenghX82nOX0Z+1wl9
UcuKwMw+UcL7QozBb4Tguoz8lJtcuGlQV0Y2Ns54EFwVnjf7u80ttQHZt6Cktt8hOkawAuiEQD73
v0RVsmDhwouaXcglbP0PVexaE0B5qwt/yoI9fqzwO6N996e7kgUpyJfVEPLhW4Jro3IxVc5eB1eA
sb2Y6x9HvEijubwyGJYdgTzHQWToesPigt1DjRrA6AwduHxL9S3MpQL6phKJdUSycWbBdn7JqQVU
VSZkwzqHb2lv0E/miOiZwvP8mn3AoKACS9Z2Ri38lCqk/5BtEmeyk/u+09qmBCa1vQ2ZCBJPh0Jr
FMumYfR9fdNMw/m3CkJO7OjP8bu+0b8zslzj1wTjTo8KyeOLqLVrCz/l8KOAgmo2Yh9gqWVMvoJ/
XUMFSkhAXIiyXuokRkGWiaAT+6OOkJoqbnapoiU8Y1arBYLn2RSDkvxzNa/oKmKALSdndd6HuhMJ
15yQrCXILk/yVFjXr4A003L07P6WiOJey7xxVxdMcR60rgProVtL3l3GrlQbLOpbhyK+X9hSX4po
6ONqMc/ZFVc2l4ihuA8rsA7fi60UD9ZtMD+pDvDpgVZ/Dw2u1xuDy0pg7BldqqMySqR4d8xgqDDn
wcDM+NI0i8zlXsEirmKCu3ULd03MaeERnugNcV5n4yYZMG3j5ayHup37vpJ2HC7tWkv6eENKeGws
B0tN+KH/GTd4NBSKRlDdipG113DHJONpDe6JnipteZWF6teShLegZU2bondmWp8rQfKCsfGXpJOw
2+/TibBcn7bgSkpJiWZBNaAEgmRK7h12ibwp28b51f0emqgCRafNJTfueygBzpQ9H4njbj2OLs0P
WfE6ZClGf3XTjUCMcWAbvtIWlZWA97MIBnC+ps+VV4oLt6ov+v0+k2vTrQtuC+Z6A+Z0qU0W10+Q
TtWP8kyChY6g/w03/A3TbD9ZemMoBKYMOM+zqtsHVy32puEG73kzChBRJdQD+FMIcJpFaBinKjb7
9uwXzbGJjeQUJ/KH1RDeCSsXPFAPUlYSV8K7HlkGDMRjHn4b4C+bbOSyLy1hQEQTMxqlTvBAZIRz
0uUVnR19VISLkwgm+FfhbOk/wAo5od7503/YvEAq84COVopyopFobZVwhd/OVD2KemCmUj8eniZF
F6gN2AYx/YxjlU3Tr8l7xGTlMJtrWYk9sPntSrD3WZbMvGx47srMKd8IXh77uqHYpB+V8HOg4gMz
EkFawX8LIC9hTpV5t8gUgyEyh9pcWY0ii9o6C/TGGJxcQomtrec8It2gGMJDcGoPdxaFFBdLYwLN
fIWtRu3tTU4PkJSPBBJFhXlmsssTXgx7HiYHDRCKxKN4lk/fzhTM/0tYB3aRxUVTiDN3sVj9HKOe
UcUjUt9JTsfw3myn80SZXEeoGhsTL6B2+qfkgQh3+ENJs+oLH6u7qk+Z0/HYf9VcK4O/lOLOkgN0
l1P81VnQyKt1YbVYWu+Q2shBdFTpbbntOs/DoWpIqe2g1ahtlsjSRDaMgbjbZg+sSlhKELjEH7cP
m0KKwN3mI2Wbx4wxKeolqzPgG4Wly+LiUk6gvTuKkT+rwgIoHRb3rIDIUBAcKptF+8j44Li74Nfj
AAp45KLx3Oo6RMSEGMd1Gbb+nozewFDnTi2oX9F5AwjA65hXxkvq2xw/zmxDDnmrw5IKiGWdfaLQ
6aQu96F7OHPIsFFm0m+fZ+GnGYtJQ/20V/cP+RvTzJVXfpxNUPn6bXj24U/8bmnannoyNp21Z+eh
p1jMleA0O0bKjF88Jd0DmQ7TBhQ3smdH7Qyk7isMKsZhyPMfmBRW8P8+JtnT0nD5rRC/spPEfAi4
/szI2AlsrA28LKxoRiKgJW5zgjNRYD69lnGGu6CED/le6tJZWqMLZoEB7B6EtLdpmMUIdIrsOH0I
jY2M5L6DgcFvevTTf2AVC6p/2qKvz010vk4aXUHj+o16/+TKauSIpLT/+Gs3AXYuXeFl7C6mQkFT
4kH9SyXRSYRRTtYswSDx39srMgaO6eqXaTNd0OsLR6LXFx/kW2uOMZWTXStQURfKiWlxxU028ZcG
Ic8yPT05xvIDwdGSWX4RX39xNhcrKiw9kQbRvsDJ4LpnSuIKImRCkj2aKyv372DmLiDlPiUDlmbv
ZMpFo3jD6bLgLDxp31zl/L4TECC5WBJidqFg6DDw1OD+Lck4v3BDXlrVVlYqHG+lJnohANCBjBl8
4fSeXelPmQCVViFgynTZ8L2feFJf02Z+QXixM8K2hMgNF6xRQ66sPAz/lrnN5CbKxhPhEL0zuYdQ
sR0skus1mD4Emc9V1DJFkQRBGqD763ULRhoBYJPsgX/X8mQzOi3RgzxI/EbTrNn2XwKnc+eNsL7Z
Lt2danMCasdBFCP9C8AqBh99rCgNOSw9o1jU8j5dLjHsHZHCsKjcmTMn6iDAlVgnf5TkamObjFUO
2TCCexSLbPnVMj5yhIdoUtmbTMIL/MrowetriNKDMaTuaQT2vVFxvP/R0vzBc7CfwpLhn9hJnADH
QR0LlMshnkv+8WYn19oh3mP/DoF/1JB3LDqFoTPpRmkHBRiaeust7+1LIOLDIKFM0ynBOSxllreF
FDCagHDqcKwXYLyTiN/A6tfu9mY/mSDjqfk6SdFG4ck4tjl+h2kvZAf1mCVPGMzDMtgOihNqhCNz
najj+SPBCcY851rRJHOD4CGDTJsv2yn/EnDExTSMPWVdlEQ8/Uz6szxJblakIvsqyO4T04rZAafc
nI3UQ3krf3bGb+SV7pJ7wS3bS4goV2NybnS8jDYSUnuK3QppJEEQrpkTxB9D7nChAPC4zf3TMFXM
n456xMGS8l4iOpDq84gP65UNSfZne2a8e2oVpdJxKBiwaTrlVO/4bSnE71FSyPvWAEb5EKJnyP9m
FExTdYOn0MsPRObj8t5ynbLJLofzCdqthNCeW52BctgrYshnJP2UWZcX78HsqUkylPx4nGcpxHMu
SZYX6POmOCX9WXsRYplgCgYceL7a5w0j050vH55XYX5rujPngRmPo23AF83soMR060GO67z7GdL7
kW+kDN+WUJBfLtQp9jBGZ5qVSleZQsM2qYKbBKjYWosQfj10uz6/CJPciyvsCSIbXzC8SgAfL3Nt
88ZR0NHO2uYps141Xbib9lXqILVlzADS4TaBI9kPJoeBO0C1ezNivqSOHtR77PTiG17tMivg2mpS
2Xwvf56hrb8FlSI5CC5cb+ihaumpCnhzGRUt+ITBu86uWjc8d7tym6v5eW19iaGmsFsmU2ldWljA
WBJwt6Zz5RxfPzCLG/Sruzn0KKMAH7lyrUflwUvDdOlCopNXyPOflIjKwCvWqrn01vVWE/TGpjmM
EJZqngMpxyejZ659ZgiR5jR8J5V1pw/fvJG4t1LgjzeEdT9Yu3lqjVALRudNmW24zwAFofR5nR6k
Gp6JblWu/fCL+AqnATU/SnqBTVf6aj2yM9wHsfzPqzAz3sUAmcZFtyD6TWN8nq3EveE+Zbr7F12r
Md+skQ1lWh5cDSzJEgAi0zz5GE9LBOVLuyOb73kwIQ0dsFVtLCsHeoT0YCFcE+4pTsAAESam7SME
VZGxTOuC1UeKuBSvUZr6e6FlwAncVAyhyC82yGY/IzBdGlXytXUX9JQ0HwtcJGF5ZmqRxgOsvxWC
1yz1MicHN7rLH1bKn0E4poxMdITwYkw0OFqmd1LdTGvz0tQ272c/z3FHIl+WC4UDr8EbHGIdCQsh
/BSCkcsXmD/p1XdCf6/9JAVNK9PFYnabz+b1Gj6vOED2I/JFnZSC5JK7KBJwlaapFgdDSlP6Ypjt
BicGGjDDzFNapTKR08QmoFzDsV2LCmYL5ByNp4lf7wjGnbBmSJT6WQmfypbsVhI6j4pbqeonnJO3
rsIMZXUNdrwnSNrh4ejcHY9L7CN0uM2Wf9kJ/wGsv+aHn007vZjCOUO5kpC+KtsD0SN43Lp1wr9g
EeKq1DY58DbTGtDhCZFKzgnkCxt9KSuXKZXXbirLj8pv0+Uosfy+ic+8rTCLJJRYDieFvvAA4Ptx
yzZB/b+nZmAfk7wMGYkKUCw4hZc6v3lSRs1AWc+HcCv+m8GcHV71m+Ezx1PxjlFH95LPmla/BkrH
/uYk3BoAPdrPR3v+9RjD2M2NR55Q0qzZajqs3P/1vlRLZNfVb6VcZn6ifZd0VbALLOs+/i18VtZr
A1hHxEqgb8I7MTfSAS99jG04IAv0I+2WvUQe0zI2LukUc3f78Ot87IDZjAssroQA3ejQnF49ZF91
vF6+M2de7axryGSS8kt0lLq3V0I4JSDsm16ajuAjxqRznUXNg/AfiKm6fqvFvlbyPzlaMJ2eBOKw
Sjlcx5Br1KJRZH4zbpa85pgLiq/tUIOHyG7SJMhGxDBCUynWunhITS9lw/in2ZG/2pcFSR9oTYI2
c9rRT7W18MO2MKXdd0MZ3Xe0R/xcQ/GmtRl98vyfHTtKDb3E4vCfdSgr9gUVbtMHyf+eR3+UTgVw
BNLnRgwMSBcoFHliXIfoC9SukbNO46yTl4hq+iMIZVWSq6qCXUFtAjsarjj31HgCslOJOxzHbQOy
iDgwz1fQ95k/+sRKlhLdzISphvUlkuu8/ajQaAUPriUSm6rTyvw/k1jy/KEVSG0MJDvYpxqw256C
QUg05sfNFYZB9VNG6s4n1+RYJouxDukFgepFeOQFIwZXvThd/F67tb133bMValfbFxA9/G8c1tP9
+Wn2nTF6wyks7KS0NuT/JSZZTvQRZ9a3YnP5C1mL16DhDduckZ7ADIPFM9BtLGjEF45gz8kn6vvx
GIZ3/SQ7MKX/v0upyaFFjO1rKSQSPMLizQraKK34YdghwVKJAraY++2YgaDpJL7U/Pui68UkKbHi
PByu7oK4CyFw4iwyxU5aD4l+6v37W9dS56njoLmADm//guqKYEY00MOsdnMJqhb8v7ik0FbRGr+s
D4uLf+LYfx23HlHBx1oORkpZU8d+cXxasg/AEJH7diQIiz9LeuPt8G6yYFWWjGo92ZYPrlRh2Pqj
qcorTY8RDD42h+7Ri4Qg+Nxhf/+EZi4V/x/jZAU70zTWRzDoAp8kEgY82gXkkzmp+r+dCjMQrlpv
bePs0C6aaGLXuNbASgoJl2vfzA/XwgyH1KERl+FRdt3zmqXbfj1a3ybBwfKAgmYdRFB30sZXdshj
TVZEnmnDmEed2RE4dmqZVrGILUgNm+MhBGFgWIjmeTq6wq3mnsGTkoHo4HltSyob3evftSB2wEJh
U/mUKB/waje5bRJb/Pr2hfiOYvTkv6YZCOr32u13dfvNsRbNNnX7syDxbtEBiAGANvoLhKNlCpc6
IHdBvuVgMmKRaCqrenzhu+aanzH8tszba3ejqJ+vDD7mAIRbIIzDtZD6LZt/3pd8MP754goiFbXx
OhcVN0cEL8KZ8xwHRhMkSXecZrJTYNGzuO0sqsvovjnImLqRePhUmFGgyk9yMAF8/WTzexOYS4If
+RBHfgtJfg2E7cCT5znvrKBIO/zSR4NAl8nk+veYH1xtuPlgLyKgOjaheAN0E20wFgaQ3umb5B6Y
OBGnUrj4YaOaCpGAb0gMgG4vVeAib8e3lJCRxl9O/ROoDiVtJad9f//uU5x2E5yJ4qzYuSglIHEQ
4t29rQ2MBP0a0fOqEqgWSD02PJvab+t7d+CdY+dILYnhKNfMUS6bMVQpA7XM3yF5aEUQ0Ewl+mwZ
uOtWs+leMyNeHQ9vtxutT6Kk4NehhDXdwTFX9KmpKrWs0Yo3dhVRgyDr83aJtHRtCc9NNDqHnL3U
V1XGRGRvi5FvVRJkJNg9sm6urrjj7x57Fd8WGD3EpBl6j87d++GdGoCqUqZm3eYCdQHTrI8pQWXH
8hBOol3Q4pIJ7O03O8XPt/2utUFukjOB+iaNd0M3un2v6FHr38qPD3hLoewUcZ8mjHXtMg2xzrlz
zby+92KwNz6XCtMVEtLph/dhK+uzHZ8eNdMHrNkP+W32QsKcwu4Cj1PUoxIAHPoKP6s//Ur0RqpU
r365SpiWaaC4Au4RlcLkE9k9b7cx31n3jAeLkq/NDC8/QX+NnJemcjPwcFbhwG+3jye9tVXBUeso
zKskByr/rIgu/fY3jbzoDMgE7EaJo/ocnrNSh4zTDxwMFEKnyUHhhv1C/dK1X2daJMBBruZfAkdr
lcTyu7BC8Eole4/IoI92I7fDf8od8IhXgVMAuajn491V8XP6vWv+5dcL6y94GmA4ugvt63T5K2/U
lzLRvWgsyYM8Sahw63HpQswudIME11Lf6o5sJIq/fJ+NyqBzxYEQ2JzdcVB9SRHhEwltYVICyZw0
jHDkfWCuBn4eHvBUhsMKA1XSdR9w1ya4BQFdp9RwbNEFJsY9+OamDeh3wNllyk5fv2H+V4xUlQ4v
fxlonpLjr8QADWEI04c0gN7g3fsPMOza4qaBomcfG6leqSUKS4ZpPY4tUAJghKqRnqhIv2vtoacb
OWGn4DmM3MGIjMth44pja2IWaDnbHOGkXdOM+54/69H0wqWaJ7/iwPQNE3jZhLhBAva/JNY9jbr2
ThauFS45PfN8ZkohIzqR3LRMRA2nj4G78U8YVUlkOdAXM0eVYoKsrdDLbG9/i3y6vNctnNe7XfhJ
8yxUOg3R7J+bs4ETchYxm3X7CPMQ4av2iRuiHC+iZ6KyR2Y7rD85WPZ2YBEtN+3ksFb9qwkFYg9S
B6jPvR59aoGTIRb6NBcQ9mOtog2S+zayMa6d4cwdn4QWmW6QU9jszaXEkJSoMWXgPkbqpTUqpBvg
BOGsAVkGgGeWEdchmzf4ttVYzVcxt2sTrydx/UKlqg3AOvHfc+3gU4HolM4TnqKsVL09CeQdl/MC
LVY5qQt9YNY0wROfIyX/GAIr1y+v2gfQ0MF9b8+ZAF+ZoWIXpi8d/rPU6vDgDEy/DbmlnxKLPq7P
RhQOXWVDSObyy/SRBNbNfW77+SLXr0tiID5ZZ4XrTwBSYzOTxWZKoWv/QP5Y3xI17AYX8bmd/5m0
qr+OB0rfb8baA7YRAaF3EHkqa9yFmjx27hUC5FDxh2CugUvmMzh2j/nxBC+ED7xkr7ULZFlMwYwp
6a+RjO9TxiqU386LnAC6s6Zw49gNSyfgZOSYqzBYwe3u9CjTV+siORX4FU30HoehfMzuP9wrQUxg
Z4YSuoAI4UwqjskT7QqU4Y1fyN+GLAPDLWVW+92Mpw0V48VttjOt41CSOGPc+SFySg0wnIE8N0Nl
u0e/ITg9QOrAho+7WY5at8t5dUzaffbmFa35I3lJMgqUmLsdVtbQn9Wp+zdU9lGgu5Itgj3wUVSg
XoSNkJFC7OFHS4BTJTTXTeklcwi9/3WkIm7LCKqvutFJthCx7tA+6RUDYresuVwU8m1xZO4+ubvP
vqPkbZoNUKcZ3e6byPkVHoGO1BFKYscTygkCoIIj/dGpvdYqF1ZwkFY6BaFqdWT444NQ5+GgTEv+
dnIgG9UmSYGUSwerQTsyWQq5Cg9Zm3Qo8T13nroqqYJVqO1Dn40II/31UDFH5rRclCXWsEshXFOR
KVnvxwy7xpGw79JF+aahbWYiptNEnEgc1r5/4oK9tJ63rzDv+yLSCU3O67pKqiE21PGGAh8KE6rU
c8DNYp1GhkrxrX9Q+I9iS7DJP9P6X92fNi7xi+zkT9njxDp/vyW7fPF3LN1q7ht7DpimEyw9kznz
N/cxUwRAx5aoZ3+v9Wr8ZK61JE1db6rTzU8o3jSt7W+O+MxPZS7T+lRMbUc4hT7qgN61+vnoPzBQ
vVPXUeFUOynusdMssMRWvKzjdybANjXKk1iA0dWFnV71c5P4jJ9+GGFnQ43a+JKLbTMEMNEKDVt1
XZB3iSYyvnbefLPBcqRb2mf4fNWP96TWL4XKMzjB2NLhYhWdJoo65B811WkABrJp0BWz674qplXA
X087G2NoZpsN0XuqM/B7jQbX3Iqc0cBjLsDKI7NyyZqOhu5cMUzvtwFG2v4xFkbzPn/wyxa4Wpzp
llANmOrr6ebmFXHAHkkTUo8mtrZPBuIBFTzO/MifPADyXuOls0LdVdU90Wcq7HcDU6wqwEfvLdLr
o8sMfEnXePBzgJXIAojmvYUNFlN/Slh/yKcuUWuRxVZVDQHIrigaC21Kj7Za9YXMEE256TauHcWv
MJn+2++qB51it7DXFvh/+4qijt6PFnMByv4xfVCYTDy7zSci8T9d+8anWFpfODcK1xERN9lKcDQX
SirefGpndrllWHn8VttOHLfzEzic9EsdiWW8en9ExWzijKjJOmf1K0IX4dDJymrEhrfyohH4wCmP
NcoqV9uMzMx2JteaVcxquMty+KnL7skOtjGzdXp7DzcstJOfS///1awmtF/rozSqdoFUbEROL3q7
3dM0T2xLLCW2f73yWytEPpJ65Dm8iFbErZP8xtQzoirf5bRikdzCfoJ9WZACgxrTkKd0kmx9oD4A
Bh05AARZRvVSLLY9NqNJno8pWNZJdteFpbjLDqPK4jm98E5Av5iuH3vmmgH0yPeN/h65tyKrdpE5
m+gZSuBKJaxIz6UGPC/iy0y90uoLb/7vYEzTXo24N61zNoS7VhHGL55E2WjI8YPgH+OdG2vG0T6b
1rWJoI3l3hbdy7yiePiTmbB/xUy0jCWLcwD9vPSdHbTLKBAn2lkc96gtnTCw1Dtz61D/LGf6383S
e8faEFKlR7WCEYDSAor1IhKUZ8jw1W/L9a0XjyLmDJZ5A/L5PKKBWOTKZ2SBYNbNNn4STbQTcR+Z
KyxNNYs7HIqQ5WkO5/b3jR80TbzH0PN0JPQOWqlnoKfHOaGga5vAQbXSuI5pNPstSfK+yYdNc0H1
MgdnlJ6tAl8ddht/cbZGNU/Fvii5+OHY7mrculku2zMMQAmHU/s0jPWRdRC+qrWf0o65Y30iJhlI
Tmz7lwKYeb3vCBbqJ69cb+GEAtpVKpUKZMQDwtQrFXrhe6KM3sXZtMUJWvnUXWur5J8ILp20DnKx
lZwyTwNzsvWC4VNwxzRKwPsngcd3vdN1e8YGiKPYERy/ASPhqCeuUd4pMqV+P15RpkSG+/EETfVK
ObKU0t2qL0ZNv5nvWk7VqDezMGyEHK3sZYYEdbqgbH6KloMoK0Awt7VzGg3RZ1WrclzqtbcZoMJe
x0Cx1nX/69prxj8oKh4MKCIiDvMRUlUaCSO3pp1y6U1iHvUDo7WLI8egCRvZ2uCMd+1qskI5OrcA
iYC8mdXAeB7zyQUr8zhA4UGuSZX2J/CzWEnT+CE9fMYfCtEvXfyxTV4suVB6mOfMOoY9Ngx32mFr
y4AOmGOfbyqpBBAFu/Yq9n2fWVWv2bVe2e3Zqfc2u21DZdbN6QLL0z3E3cN5vK9NYDQaQcZ3m2Un
J7jbkrkNpJFuIsFinO64cTHd0cLeftbxkcJQIb+eZFcz2/THkPmozMRjDDAMVOHgzjeosBuNVSAd
8+hQW9lTrZ1qaBJ1311aXi3wMqPtScbudJWk4++g6q4QwjYlERvZHSnjUKpuaY9sLKI56+qrx3CK
6/fYxsJq9ChO+Ypkhgx/0kjX9wDhn3SqMq+Sd9rmeqAVOHMvnS7MasTSo546Ny1cIyAUWU9d3Dk/
aOVOp3XWMWC66xzKbp/G7t0PnLT7CduknCyferPJJqO2pdX7i0tjsDlKx0q7hHB026NXln2UFJ0X
r3lyGcbC+qTjD2I8064gM+QXe2OhUpYZkEuOmci3Wq9VBT9/ZyaU0wwuj2jV6G4Em4pyP8Rr5Y8E
Lk1Sj8Y0oSg0ZRjqg1IH12IcSGYhi3lXd0eeU5B2RLQXbyQWmh3VorspVSHwYmMUB86sJZvd1uXw
YLUuhUdp1iVMFtj1XRz3utdsGkf8AVJ7iSER1Azg8D1JL8w9DXb8seApXkZ6wNq7ab/tevkOc+gm
42VTStJnnc5yufYx2Q73l7vW61Bnf2Oy3gVPGUGbpbBV1fhpB8EmATIjY0yBxlndPUuscAIFX9Rl
hAq/0udcLfgabIWCxtex0nXKS4We3Cx9YFi2f7M4SudiXqsX0JMH1uTNoOCPgfEa3VQbKZeO1ZLd
zzrAG/cUCtphPy2l8DfJiWYt8V7kJGZDecehzlTGm8F4EN1fiLdY4+xNai865WFiOnHrzLfvcElF
sglxjMWrEwvkUE+uNJFd7Q+mKhoSpJGb1Ghc4uZoGZVm59xDazK/ibaJensq+uWydEDo4PIkq/iD
y1Tem3v+9zGeyuVgLVfcC/inZ2/OigL9F2lUQLu381tGKRXG/l7VkGKpeLf7GD2eg6YxBpdKk9Yt
WFyAvyY+XDhtffdHfjvDBXom7eTDYkIqZzT9VStEF//1fdlDqPLADkvVS6EsjAn2taXYvOJRl57P
ErIQE4QDaMNHfhZ1QeD5rQT49fwUz9J3EI5LHzgeWfOT3Tqt74YhciK/R5jvkD/ByW7+VAn6Hvg8
q57/eBmT8zZ3tr5AdAYbZmsy2O88eadL0BweQLcWjEUcckiZNxJhLE7x963uq5jKUkQcQE2ga68Z
ivfO8lX3T9cGccPsesm7dKQB41Ea/JcBf+cMH4/yL4iGK8RJ7tZA0XhC/rEwyqKe9CSmEtgp/pOt
ocPzeB1yj0QsqtsRmPAJFTtP82D1OEZgaWgFE9Fnxbz57FLfVR0Srl+ateT2kb+aymTgjlkONT5t
KXD5VajcE7Nzmv2VLAA0rPDwjkbzkS4t3R2RaT0IGc8VvmVxRbuxs2C1GgF6XYhk78GViXQS75PY
RunXrieyON8qapmb3ikDRiqSa8nNtPg71ajxn0h6OAgbDyjgScwhi5BJtwzhiLP52DFWyuQPw+yc
nKipxf7BkmUT0XSIbZup2ZgRV1USouTSrwgKVxutrnchbSfSi3jEKnvPI5yKKK0UPTaLT7g+b+GJ
nyciD7fs7zPyNEdxNltnid32fdIPhEBPFP89xZFm1ynJ/r5a6PjYkeZ4KHB4OfgD2PoCOnD3WJQz
uobn10mJOJwniEoju09mdFuSsFBkZd/QkF4GY33YUPQNiacSwyT7kywzmfqvJB6uXoGyE2D69d5k
HiD4RP42auw5LO1q8ib5dWR29Bj1l990nAIwgorxB40qnLLC+XCedsy+MqoSRCqgXoi5YS9P1BXb
Tq8gweoXfw8a/UCDIi3zovsM27X4axR21kOh2dp+DmN3JqyXcT1Q4eIN19vvAU95pvigBaj4VWxu
4AOV9Pwgf7udgAZZ89l0o7XF2TiBbLeEhDAXpzM70c656myx5tw53LDShMcxEI2/Rgmcka0UK57i
4o+FMjky1qvZnZnci/tLpEQ3WKOfEjKoqnrW9jAS9zEcxpq+Dn9KiuJYaP8hcfpB/G935DuibdWy
oOZ4YylEitB0d2mpK2ZvbazhET6pEPz21ITvW5ntiSRnIAOLKYmoVyF901RMrqf2XksbvpJG/Vt2
kTJa5cpSfSTB5/ZemiaBX7sABtczIsAN6lnbovC1JZxwvY3WryRl9MSGN8QzYrKpx4fuv0HyZxd2
ogajirwIgKQY8Euf9hKfJ/E+s/Ie6T7fFPLUF3Av9Qej/zpNUbUVpP/lwk7s6ntIfD4eFkxYe5Fc
+Fav//YdNLseRFa1WzwqgIQhp6hQgwJHBrnJINyup6MoOgHDxSZ4BYEs+1Zvh3j8h3CgosrYa2d6
az92bZ/V9+SWK7E8T/uxVrvgNgV2OeyGV4YR+PKZnxK0BI3ts6dMa4jJziEWqvJw9GX9EDKnpTsp
yDkkimRShVQ3zmvovQ9COKLSKENEtGrDg5WgIlt8A5gukphGmQQ/sPd7l6GxrSo2INUNwRgsXioc
dGyOrFE14a5H5Y4YSiXuX+nYgtBHZkdp6rSqeRxIaHa0SDM6q7FIgLtw5TD956RqpHCoPCc6IFw2
sggt8ZwZkN+2TMPa7v8mfDIztUIKGXbO0J0I0fGHrRxlPScZdBrecs1Je1ir9+LNvsFO5A032WBx
PUZid/40lptCLgh3gv+Pz0GUkghsXBcBAEx4xbCBHcWUPurRMT+lETEshQQdOd/enZ6PqFv3H/HW
AgJNx0xXCQL3XBlrSnnGHm+spK6xbjmPpWED1aZhf1LgyDMbDiRtFEAsa/yn7MAxVjvKPnecRhcD
QeyC9H2hadmDd19wqfrfl74/xkXNF8qjzu3f583VJ9iZpwDTYpbnyOquhV1LyaOlNcfUm97141nr
awUIgoldrbRs6HA+91ugu4qX8mYz+W/Li8tKSSbGW2Hv+LHfIW6w4IS1T39ibbV8yXKZ2ixKHV0v
7KSwvXTIJ3Uph1e6qE4F83Emuc9+UL97dqygYpZte16vrjridil+xedvva+l+8EwEnXwJlFNE5P1
3AAs/LdDEkTdiPRJBOWdh0kgDHNQcV51P58kb+P49/hWaCHEx0/5oSBV2xWWiaOvWeGoPKMG32AI
Z+UqCRAgeEibtWH44hOBCxTOT7y2xChwDvDs4pqyYuL/ha3mygy3XfiqoQDKNuyW35PbHtC8SNgE
klhgaslFbhJyv23xHnYuW6FncNGiY0u4u1Nc9I94ZyzWCM18n41R0c1+TXOUANQAbyZHTaV2f7h5
jVOrMxWERg23qb7GHbE1XUxQyp5ZgGRnhT0cfMdeH5MM32sfRIwRlXR+9ylGb3RPMYeX8WppJEyD
hS5AfoM4ULS8vKtdQbSsK0fm3nxvSQ/kecf36iabYRtBzK3MJlZi/x1satunbyVrYJyCJt6du3uw
oKzZWXAIKYnHrTf23/V9WgdvboM/TW/lMnrGWp62h3A+eF7SCtmrx8Y7KMrSEQbhXjXJFCykeimI
VGQF/29rOuqTAlFKhmUTpDmiQ2TU+EN3cDnEigm6mw+4YkgxJm+kqrFYhF1+QEA/WUrLBWzBMAwU
vtALclTmkH0hhcnFktxJ3yZvzRTVBCpgZSAieaXSnQOgjqhjyUaWcTBKCzO2NuM+5eMfMag4oM76
HkBy4w0jGCvU3rPLW8p4pBXmT8SBdqw9jLGVdV2qiiP5oz3sqAR8I4xhWLwCNroLfCByPRQMKJtl
g7TFjLh+rCXYnpC++R6zDzdKZ/zCst0O68tVqbvgoJIEU8kUq5qHTeJCyGFM6EOYkC2XDBoJXokN
MOj4gb9RlUg9bdnCVWSLpfHe4tA5K0rLGXxszte7Bzmsl0nFuVY8w8GQvSTPBD7oCWjJyDBbCJct
JeDDk4D97v3Kk0hKyUmCN7KNiAMmDfz2Uj1apXoqVGgl0YoviF0EIFrFfo2Rhm3G9ogMDZqMylPY
PWusPjilRdtd5wAfB6AMPbeYM6rJUqTIL1Cgq6BecpJojHxqkFVUN/1be4ApNaY1jZKoT/A1orzl
3nvNiiuqLAYbHgcwhLjDWVyqRYJ4ib7h3VhSapd60FrQCeiU91yKw3WyEqPEUhAl7wjpnnc/UE20
MwWkA8OUE8/rlgXmqtYkmN0OYoR0hpXnIVqxUbYrJQRfpSjRLa8ZfNjcselSOEC/a02baWwE5bek
+j41KskYCc+NDekbstCmDYkOhWc25UOTw55GugEykZYAew1Ru2LjDVRxG2XzgP3v2kWYoM/35pzh
7zoERyViHjunUv9R5OI999jHEXQA7QUwoHMburaq5BhrHY5UdiFwD2Au9/ivxWut5uLu2nIFX6/A
1ynJVZYF2CuFctwTKvnmwlgPRQjUe5EZndhObo3YUSvaXKZe7MbXJC0dHU6FcuOTbqmFFbWv6mzE
eFA1dm2OwaWaE6qfjwl8/9iqO14oE5sOeLALQizga7bfJOxBWk2E6QzXdFYZPfQBU4OkQJTGGQlL
jGWq2l+/Li7CPnW9VmXxtu6O7YNgxJyjtLvo2n3JhJ3/9pO2jGSjFcKZF39BTuya0zUFAgeTDQsi
vQHIdSBL9HmvOD0QFbzNmbMhiWoTeO7eCBIfLL8fh+OmqxL/jmpOXx4yn67ovlC4VoF8lAk+DbjV
77MRI3xmNoGDlXOHQdSyGqL5ltpuyH4tqZSZWCM7tlVunT/KVMJWK3V6fxxfbRmy/1Te58vd0rmq
mMXYnfjok0o3gy2hvjyrAj8CdqUfc9cK1wfOUJ0s5R55wEMgRdz7NAI8EEhe6+vHQkVoxJf0BO6P
ba93h6eFDEblpf/BatWDj3IVnrOL5P+Bzby7lyxNyhNX3UheNiN5s6EQuXua/JRhgbxZorJgCUNn
DrAM2x5jOpgHzUFjB4sFHsy7lf5a0wqqEiAgQFGSCY8FlMyZ6/rfW3WUxf/aaBfviRYc2/krXcOv
5yeK0V4IqNnzO5P5Oo6O5y6rOv/PW2aUwgjSjbGWJlcemA3QMNrPoDWvkialIoKW8yoiddUrKNV7
JXgzknULqCTG+KXNiLptqgDWlp4rW5HJ8aodxStbfMgta63Obvr63IMPxo5Th1d3ermdpLfW/bJa
Ka0XWEuQQUKeICXST2gfZ+pv9DbgrBahd9W9eouxFaUs6IVoRATshrFe64bbvHfw0B6vC7wUwtS8
ptavCsvCXxne2Y+beucvIWMzUqVp+zI9z89uRWbnMJ45z5ai+stLgP1ngYuF07DLEny2DZRFERF/
LuBFNsEI+xwNd6kvWUcIbiQKHM5pEvXKZG0WJXvGwjKNiY2DCtnnXwEM3xg4A6sV5xfb9T4InIRK
kp18Lay7/YDE4BzlcWcYGytktlrfyO+zSB594Rx9EUnNnvZZXAlXB154X3UPkBK3xYrQYBgMoh3r
xP866HwoQQdjeKth6oXUj9VujvQpceMRQj80+eX6odiUzgHGMVVUWqPOviqgkvkI+1tyQ0pgRQi7
WgDXgo1KPHZmbFlrtWD4vaNAxioVDclw/3uQ973j8ZvfhHlirF6yKNi/04iQKw9axlAjiGDDAgvU
+Q7a/EVWwRc+AGLSLeZXOAoO5ZzVURAR6nos7S1jp/fUI09INB9whA6BC2FC95D11ethJ6PEtefL
/AKiDI4EKc4ONvoJJteHGikkCR6F7x+epxYxaDTIupsCn0UTmqa2YJ8l2nga5OsA8pH+M9DszIKk
XwqwVTkXhqu5pu8cJms7EueZ7GZZWdMlQmvwrW1OAc/lWs2aT6LSmZMbMZfTGiPPBIrJ0fN84RyS
ABN8FhVOJ3O8kBB+AwtAwhTOLFYm8qMhGnjn+kJCuV1aEkXi/lB33P/A0pqlit3zyY2mAcyKSatj
iIzQ33DdPinJsY3LplydLKNoGZMI1O7WFnCh0LPXaPDFEL6V5C1zeCuGcVppPw0Azym5Bz75ULAL
OATcI5cT3z27QDAPehbbHZw+Uy+ZYuUmsghGF2IN0V5mBTJlwtPTEdJuHNmXSw/u328eIPRgyj9X
Vmx5PRTtlof+Rd9xjcZMXE9AtOIxE5YoNhbjEe9aXL+092UgauOdC4C9P1ZiLXLcFHZEds2RB169
tfW4bUvNMYJrSbdo8ABX7TYu2XW+O5GDQhf7PeGCoiXU/MMb1ftv3AGQ6s1pRi4YhYaaKSHti46M
QZ+80xLEgNVVT+sdM0O/ObE3Af5/DMsLJc3yNp4CHmL2C3W6ri+KBYLSC0RDCkuvOTJkPX9DBZ08
2oUuWeTgrPTpHk3rOE/jH+Z7MIbimBJ3+1rRQLelJMhq733T7IMO4ISp5FGDxpjxuoi/1hySIR7z
p2eOH0FUyibNUsk8o5NfzYI+CnE8eXKfnovagKEdo55NgKscG6I9uKJJI+2qXfxlRSqJ6Q2epJWp
wZZh/+3OCMfTVRYokFMU/69ymqHobJUIgfg7jL9H1ut1XQq0BDUvW+RPXDhZhu95y2GPsHsI3Oql
/LcENyktVx/oXhNPHpe2k9vvOz01kUV8sV05/aTJW374jNIxyYDRgL/7FNdvIjLLvQP7Q4/iSNnv
m59Y0pTv2+b8v0JU8Ge63/tFTKlnQh81ocdzpWjWAzA69sLXFL1EHzkKyTfO6chxGj+6f4pOh1Pq
hkzfgLw7cuMw88qy4GFJlprgpNXlzEmZZAegZaVmoZWeIjdLihfjuUOzYxOwHYBZDVf7dZUs0Oi9
EyejIUun040fPqbfugKOxmQ6kLWcaS/4lPiJXoipuABD+wQHkpXHhBMiJuCN+TE1zSSz1Egc0pmV
j4USYOgzjlNY2DvhTHuTgO67Q8gErOIKMW9u/odyqwW23WaYYg6KB5sFqnnvAVy4yc4pp7iVy1K3
xDq6R4bGESyaiacN+jMzkO20fEY+020enlZDT+STJWlefBjAfS8R4EYTGoJmcwn6k4CPMPMBpjBK
NuMG+NaluB/UsRzQfYVABRuY+sb2ZVOqQr160yCrg611lSWMbdGbUF30MehmgecX1qUIDmKx+gF3
K+RO/A0IwFUXaCg/257NyjeWkafQTRsY67QIk1Ac7qb8yfJSQZKZmmme3h2OuUEfvpz68z8b3vbk
+vK8A47QGPk1JewTt3PoUQTHev2d+uOegBSuyFqc/sN6RTx7mNmCj31ufRyfCr1NcMyI2ImYENl3
uOUhFHWqw10emDJZmM/GtShviltKpuhuTsG4jrg3BpDhQWso5EQXZRDqT3z3j/PLYPAeDQsw4mCk
UtHQVUJ+G/A/wWH404R3JWHM286yn8kgGdBFsOPm4pNhpymo2ssYeHRQmhjtqlYQDCPyAtECFvuL
XYZCdjxxA3Dm1rJeHYxpe/VZBCnYFDmZOI0HlD7z/28iAyVB1LnTfqxRiVG51MopUnZHX4+mihGF
QLBe3dmV1PYXwkahnI6Sd8QXy/SplNTrV1oPsrxe+jRs1KUOje1bGDtTtFR6PTPq2ekojTPirOll
E4TlfpwPw8rz8Aj2k9as1E053FHh2HE0kt5csMHOfBjnu807ojTFtBB0Xrbu6xp7DjrKdfpEyh4E
bduY6vD6ll3tSUTREI4VdPADOO3IIjz+gb3T2zRORlXcmH6XxLkngb77ZRcI6H3lGgfCB86W0P86
yJO3AKLUzBnL3A9Cktgne3U8vny1q+ahTLHse44cxn6d5HtY780FqA02h4q7RUM5MHOVXAf2J3Xx
15sCPMdN3h+2J7gCO1NouEn0adJ2aSKcewGHV196nuHF13PcCZT4eByqVT4KVFD2wqwquxK1rvZW
25aOQCjYBx4ikcBbNnkqGLSZV+iNI5umngPDDH+YRHu0prqHQFTPylwxAsT7FS5gqon0N+OUFm88
SeR+kRed2q4vJ4ULFep72OkoXI9cbxyykAkYAU7+wKDG2A846xrUkbtaDF1hvGh1cZ5V9hAbsoJW
HpG/es1sI0f19/D23adcfWNBDBKvkBz9XOR3Gd4aJpW01rQXetiUHhxAe0Q10lHyGtJPo/8UDs1b
TT/z+FvFZtIMyXGfOM7wj5bSTOo01YxNyPM3tr5G5kwDlBjxOPk8pzjycDMp+VYr7ox5hx2N0QZL
Rp4MH65jBrWnxTgkZZPvSgPwCoMCI6SaqKlseUpVq0SM2OUraJL/KAzd6CoivDclQWY8dF+yKDiw
A3AHpVpqDtohy0AuDpmLKEbilYdE0vj4TrzWkN8nNcfqMuoVEmhdJoGHni1t1pBMSFy5JRArVKe/
J1/0wONNAn0B4sI8PWPBXPgtqwHQevw0y9mgqe9OQLFhtQ5F9+fn9FQEaQz+pIVq+Y1b86ZP5AgY
sIZzs4DBe1cRFhT7lumXxsq7nzi+tjx5IfI1Zw4LjkBTFET0QCH6W7pymseRlyEQYsqioxcRVHsd
oAHd+KFOrnegeBYt6u+eUL7qnfMPNwnD0NbF/ZTBC9lpodwOXMXqkcjEPHua7KtWP/P9zPOQWkSG
HQ4LUVHouxjQ1Yqu9uK60FZuVR/UJrHrm1Q1tuCp3V4oDJ4rm52cFzfdJdPWVIdbQId9WkAZQjBA
u8m5CFdlsE2RqjZ+xC2ky62OzuchixxWY/zQb8mlwsWxjGUZ6dsb68RYSOnZ5zNZUPJ4FNPqckdo
guSxeWABgMWU9IhKiVuLWk1sG2U6lEv3S/rKbfVslv4B9Rf6KEi5ucuNZuSBExBnCvq8UHZePZTN
svcXWSYeNHqJSyvA28VRzvSotw+9TOZb/QpHj/PugsXfmhZy0CSgPReyob4wLkixvKH9e++SeYTu
QzrzWCWitOsD9FetvtFVUqcP96dX7P0BvCVSmiHSwW+0unPCYqNRqbBBSF6QQ0DFQUVUbQxQv2LJ
AFgmV13pk6dVWlBLeELcAayNrt5DKK4OldWLg9dqHksqfBWjjifMC93PdjyBTHio4IxTQywkBaRY
AxS5p0Uo4vGx7BG09FJRbQaYrTt9a0D0tlmMOB2Bf9jSYdUttEGPIjGeUDYJHcUf32KUnwzfgcgP
vpdXOBvL+YVXZnQ1K65mG5CgKbWI485V8usGuyFWwohE9hrOMS15M9YDYC+Bvs9/Pql4QMmvYx0O
GQoa1df8CjmJxCcfQpzvTzVuGABNuHRvlQnUB7snFkp9lAH/IG4eQxc7/P3ozdbA/QzA6St+wcpf
6kBWNRny4/RLEHmM5NNLHarDT8eh9QF8F2Y81lknwsxVH4y/VRgfjtbZLQ6txJBx/2WxAJXaquI/
sbJaFWDAyo7bViEUHm2MW/HfjvEgXPdYjRbbmcvt3/V0zwfKkcpgN4pee5vuVv84HrvfOOB3CF9Y
F8k7NxzqJ5AFQB0yd4XZt8CktBy8/tH7rG3jw1cIMNgVnYvt1Uo2Z9IQC6EDDBGEk6jlygM32/wp
7SeRqf+jGrubyJgAY+SOvn5q00GXxCZGufS7gDSyJCoL8lH3GONryebNWfRmfwLT12YFjOf0t9yk
uXBKDU1zScmkO9uX2FoOydYIMtkjjqJkWiXPDp81/lFXVXpL/lCoXond7123b/cJOcjWzygqmZRP
g+7KE1XKeH9KVoXiN75WqT64WP33SMMRDsmqYySB/GguQveCsTkLyrBYyjzo+TUGntQI7HYlGWCm
2ePRU6JcBuViRHi5wDdU0FI2Wi2DicoEWtJv6jhnpSlEufiMYLIh6iRyZ2TjVBpI+ZCUe2xOmgxO
ldXHjT43YnCB3yBaY4djp5vHBPFIF+R9+Ffq6K0jpULiimajyUc06AdyNJOxW8TZe8WkiOaO5px2
poMr49+alLnO96WT/PMHNWZYmQeJFqhJGL+8TGcWtmZapA12fbgaGgKAjsZ2lfDulYMuHSTtLg90
YGoEYGF2YH+FAtc5hKLpOG56EzaDxmzqAMorJKFonSx6aU2coFhiLSMmOiSI312iPqEgdzLtHd40
b80I6LHcBe7kVL9U8GZ8SkAsphUjYap8SccQgYnMpxeGEmBzTCyCctUT5kxmha56X4aWU1DuE2HN
la05FE9NqXnLstQcswUOEmQWznaSQzUroEcrFILp0wKCz5vnVjS2jBt0R/TKrZG4Xtv6aaNh3XFa
kMwDYFMVk7I/cFhnUsZud5CFDvXlYITvYHtFTr7v/WovITEiuILUwb0xvvjmb/Oc1C9V8yQFqKvQ
CJ45H3G4I/Dhw8taWciC79Jqt2FZoxWXt4b/yrzYcycDI6NOdVCOb1n3FqUOduTGpuM4OZS61PN0
l+lcmQWmLvSbbSWdID4XA+KogN8X/XTfpU9az4Cm83n/oDGHrl6vUiSsD6z/oeaDqhc9lx9z9NB0
6x5a08Qaz+1J9Kqw+hpvPrS+AvB4ZhhGiCrVlvML02k5zBKdRt1e04ivPpuYG+YQPjs0OGBdPWzK
3Ou9jSdJUa4uDdcdpmW79p9QOJF1/pTQwWWJNx7j63iJb4yXt51Wm8TTBoYv7hhj7/VVUwtgMS3h
jfB+Jz/b3IQs2aMZ1UM+Pf2QpBO1/rXz/InaShGoag02Y3o8Vazhfd6efLR8+aRGGFvxvyWalrAO
Vyox8OsJSptpCLS+vgP4lscG6pvJOEpEA2QK1u5QaIc21lND2lfiE7zj2FE6ozSoZbSdlULBEyru
/4BSgOPbgGW6JD9go7fkn+oQsbe7diOKILO5FpqqjWylhZcC+GU7+mDbaXNroH2bAE26m1JRMrqM
Sl9rykCMiNyiWXC+g/ivttvOheXcH+qjlrqebfO/MgMNbGF0cM7G3gnSmDpScP4kmyt7oLPEo6n3
juLSO3mER/yNoYpJlnQfSyVZQJOSHtMTZl0em3bZA2uRLyjRlEo8+45e931NLXWSmVpty4tRYq/s
g59AaUVDkF8qlRJ+F2m8Z38CiXucgjuHd89uSn3OwELhO4qzZqJ/cQXmGRsRG+AFuD4h5ox8e9zy
hA6S6fCqe0dx7Deaap8+4Qk7N0IMya2/0iQp+OFY3BQRI4mKLXZ35jUDpyGDNQ169pnPdoAWJd1G
m/oNlH7t5y3BbWQooJ76UpunHhGqSV9aS4P7ycmJkioXH5SyYRYdZa0JCowpcvDOrC5B455zT+Zz
Y9qrDRkk8pPClbdxrilJbv1sLvs7+cpJ6c1ux4LmIKpEXlC/M5DA5oHJtO1IBKsF8bSTGiGtvcXE
OAiUVnxOw7bOro70uwCEvtMSYbSOR2Z+6lfiLZZuKfKN85AQ9nu6oIdSKdV2vPXf9MsalVbPbUPY
qO9ci6K3Rt+u6GecaZf+3eK2xmKEB8LjOpePbnuleGUjpRL6UOPG0Wk0NjkhA1daJG2hm+MGJdyS
JWhGZVbSrCAkG0SqRASzR60e39sZNVjXu+R5nxm3nlWcjQGw2V+uXIfSShlzRUy7CIVYONDa8wbQ
A6F0HD6fEZfYM0MwcxuHNVrjSbB3EFPms+clrr5jl0gbFFbVJfijE8KQe7XqjWMS8bwUVJGh0mW9
3uipsyC8TqaJAEJCJVnsqqo5vN2/cmU4IA9/2/rrIjb/OSyc8ntOyDgXgbWJlvCsK+yPAvEBr8uU
rBgGo69RaSV9ksptg/l8V21yrqE0mDlC4MbGd9op347l6eMCU7ZA7zkVNSiuVRUAduylBmhtyT77
tzbeqJ8/ctN01rwbS4/AgHLtqqIfdRPDUcyFZCl9MnZaYkRSNxLmCUev6/xEIJgEDb8wr0IBmYmI
oWaG455onZlryCmcaFlpdrkl32u3RXlRHifldmqd/bQGHP+dxkcC7cBygENs9n4FiTFcEDtC6TxO
en8DSk3BRnIbXJmTrZKvIniZslts+9pmTUHponG6PiYnfkG230rHp3GvBb/QWjG/2u7AVT7cghcb
Nhp99OLrRpyQ2Qj+KCd39M9JPTbopWWJS3JrYJKpHsUUX7xI4xWOlERvcfJ7iG7pxFD+ypEfNIyS
QRwIjMUI9J3CJCNZErBgBAHcft7Huq8UR3bNraZ/ROsj9wp7EhOHEATZeOncV3n33MNwZptAxarI
muteBoDch0PCNEVjIlDSWMMgfeVWFs+RJ43Ti1uUwRL1SaqXsj72qPW/licBBZYcdS0r8nbDaN1X
9JfGB9dCXx1NfHoSYF3HesBWyDlE6zNp5gy3oMz91gOTEZRUbW+rgNWHnd8HoeRwKch4bl/WqJJ+
sbmoKDHWmb5mJ3IgpScVRWx0vfoF98NZpeQHEhu52GWqLuxv4hx6/0l/ZIZn8Fu2nHDAq9ldIDAn
xR9AJ/xd+P7jle5jhUCpe4ST+rckIHuJ4BNXgHI/7rHAbH53ZmR3GZNoykk+XZNNgH6m+WHgCklV
7qx+ILPQ/lPtWKX8c778FOWluVPFhtEsnNmV0Y+YziT7v0cuTMRcAsDARKKrSwWej1/t9fCRRNAm
qVITTx5TP+Cs/MNUB0nVPwcFftiOVHtW+wy0BK5nSjjTPq5S6TiTwXAxxf6q59Shw8Y5Ho92YgUM
BLKn6YPf1OCtb+3YRHCZ3yiSjfv+g+KzUD0hpI1HN/LF/VCgV11SVW0oPk4w6cziD1b3CRgTTWxc
8fIgl9Fax/XE+fC6sL3EUU9FYh/YSNpININ9bkT7RgoG5HwEGkE+LC0SyNII619AOZgkSZ7stl86
+9Jn+i0OYjuU4iyOfRt2PzBVrFUWwiTwQv1F7k0WRc8TtsYtjrSSuLkPcOYVfUJd2zwwaDYT7/mW
uzAyY8/FjOxn5oswYppAgPOZnoQbfQt/HYaIQnksQ9fDJKOD8HYifbkQAal+ghqgtyX37yL8h/yN
/aaaOU66xLIPvmZaLq1+ldDMU1dz69MXXJ4lNbRaPju9Pun0S8nWcIDpe8OmrOV9p4j9y6GlEmSO
cZzeubWX3j0ooBt5rOgNXvh3An/8P9v99iyElQBMAZg/pv7Z2ycGMmo1Y/BFdx8yVrqkIjpb446T
LDida0/hDbTYtzYJFvBuKZv69Tjg2Uk0hULh8RKxojeQrNPIV6802sGW/MPx8OTWjn+0NvT1mWbD
mr0JnjQRAFS12SvcuRlcTl3YIsbm8b0jAJN9ftcC6UaYXPZjP0vHNJ9ayAoX9U3UoaUG7ChC0RFV
7oyoNXcaNSRIyeJRaQOIn/H/gJRpeEd0jqkNiSDaVVk7xs99lfqtKjLY84Ew5+e8uoJtt61SlThZ
BmMlXv5kzhpUc1cf87oOdCnzpCQ3cHCI8MDQjKU9lye9B0udSLP6kpVsTqMx3VRBlk7hXBoqhVOf
iSM+jw7o5OeF+ZMho7/dfNdhYaIuo/lyKpiWIEHvA7VmytSZzVhThxEhxY9avLByY+D0OJv9tQ7i
EaiYJT0LZx5aypSaSHaHFvtI0bkvUvp2kmF9Xn2M6q9ThzLCP+8PduQ65SWf0sJKJ6mTZFy+5I5y
BukpzPuZL/gqBo0pBxbNGJzi6zsgykIzCYFNSjwaiMUizhwPJTvXb8QW+YDDR9Jwf1u/UCzbb/VL
ESWM5V+65a16BuSnSSh3s/mCEfuAx8SwEUl1BAppJVaYHq3WqC8Mq5caxEI3o74LvNyMrJOw2Uzg
cfHKCdU8AWrUK6M4QCFqsgrHOJpmnzvqT7Fm74y/CsMHUdxI8TVEw+SDcl9UynSLAgQXEJULcXXD
ur/8FwpOY0AFwzgG5qY+6gK4cHM95dF4r2UFHfeu8TbqztJQP0T5Q4l19CR0xqBtULl+GGw6oFoQ
N1ZIXvrjrqyY4IoWVrV40rF8fbiJVKs+91XIeBat9Q5FP/eayeXls+cbbRASpmFhGiTWiTrWkfMP
QffGx+VNhKRWN61Ge3531MTMugkIsjCUizU06ERZDzrXxQq3fKQkl1wpdwwKGDmbxyfY3Iw8CeaL
GxOtWZHbmh+lFQyxFZ6kEdgXapqdhO59dDKGmltjpga2s82LdW45DH/a0wPeNIQW6bKhNozNUAED
0Ow8e0XrmdPRiXo0R91omxdLWbdoaW0AnBXcgwftg8n4BLvMGLX+xPHWdfOapWDv/v+05WI8haPQ
mrx6rJcQd7RZ2n011u0NZf4C1+FKOiYYpSWJJ21YM3IcvFHVwAk65//ZHRo7rmmoeSOm1GcWl/jN
PmOdvedfWpI82TF8gEpwEvylbCSw9cwnQ+KFvQgVVCvUEDQFOzBqpZItfvdbXwossqIjEFJmUxC2
Zh9N3mr1FhnLJKOMYqPM++iG7GFnSm2VhKlDhgXV0rgLnS/96aKFBH5YI+4xE2gOH8fouytzoumW
/oED3Zg6uuk4cHgGbhOKF3gg3YnUJ7h/9DtPbXx6wziQnqLfrTdoM5C6PUG7GEU6BaE7Ng2rgKUe
hjKlM+f26HDspkdZrbUM/YecP6IH5V7Q6gUf9kYMXEnjtL27ibWgW4/hImHTcd+eDv7n7CKS6zy2
nnDWlW4Us+iJ017FOP9Pi9MnZG3POlzx1XbzsNrnCOEipaI64ulLMSzKTV5Y7Shwf23fVTjA75+H
36FDUBTCtjDgPyKob2XvYV8gGVa6n5ys7hqGDfu2e02Ety64jGGJo+dd/YxurIXPmHOiWejZFVYS
Z1bEq7JWJQvJiHkHpzoGu5uOGwAx07X9oB/9OAcJKL/wlIyK+k9lY5eY0Fe8onKnOgBYmqyB0v96
VEHwg1RAXRHKgUn9I6XCmBpRG8gD9eD+vNIr6pdsE9mYq2LHlFOjZRTAyyCiTTeDctcIjioVF4Cc
FVEYU7whfi/wIEr6cZ0kYne3YgAp7xOiB8juQ710QM1ZqQagmB/i1fRcwyYTAiKuDYHEh/0n9T4u
mOGU5S1jdjCBkX3OY41cF6MT9/edem7/eIE77FyEQBMZhCeykEzZ7o22ki+bBWEpS7Ebw+YAvesC
JDIug7IbqJg7BzGvevdg6HJl553txiBDaImqsSitFiO469WIqFj4ObWaaHGt6dsA7ZVRqbDMRta+
NuZzUthWAOgCmGvHswg95EfNb52koTH/cdPTeyFeG5m1YZiBYrg0B+VAW5eLrODKIkfXt0cfND/D
T7pQLpJXPPceJbzVASVRpLFjFTvyUnt+5B2EBh/nk5vSpV8lUmQDhQZgiDJ0Dzdu3w6eQu/FsM8S
kwI0QcJc7e30jaXbyE0AXD/J2TqfJ9K3V/4/RW8zdXQRAC+o5ApOvZYo2h9CSQNMKPTTULeMd41P
LpRtSi2taLIS9uthAfVZvDtaPihO9w3D497olHD6RHApo45vdPBpDjxsw+mVM2hW+KZc73MMmTg+
meQamnWP3h0EOgOIhZ+MsYGSor7/t95CYxn8Psd2yu96YimTK4/XPoJXVSRToZdcOA10sdqgrE6v
qJsJMxoQ772NHjkj1A4JBUVLhzL0KxZXaHQiZabRfqZseT2CCznmIa/NyPLm3eYwnFNTdN6sD4mI
+3OihPg75gNla9+WNg8G4TpptLLSaqWCXFubiTIBJ8hZyTocWRXjO4V1bpVt+pqHSMziVtnLJEfX
zEWE6TodHD537+f+5bGRSJWGrHXyY4f5MF3AV3WXtA3htdkPB2xLgCF3A9ouX4cvVqokRNGgyLmt
fLDYx30v2+qcIw1bMw4n2tpOMg1lcY+b+AVHIFE9qSS4X1GHtZUSlCNX8Js+v1P0+dYVk6v99ys6
wdT6zmJsfI88hFtiXOFA/TxCGPDCCOylhlUBjB7P+v9nZ9ohhWPm2cVJQF8tAHWbULLD5pTyplOM
INr2D8eMw3q3hY5OAlbsFvShPTsSBjZr42HlW8wy6OSeoKERHePuStlonuQrXi/E1sDO7GtHZo7z
/ZsxtmRcSNyizanZMzCmnM0rG1S9mEpYLW2WVCbG97PDTf0pPCAzGuT8Kn/90Au+W2BZll3qpSTg
7DhQeE3AXn1xzPHkVzFEoyjr+marZ1zR+f+5pss/QfGRUSAlcvzykvCjzDPRJIoDGN8Cd/ANptWG
auij/rm3Ld/9QHNI7/5knpVt+ZlROnmCiKyCDwqNn9KUllmvOAiuGHPZDAk8sl5grOhRIBd1n+5M
APt2g1AHdvYdDdbWcyt2NhFV6orY3AGxUaihzvL8hZH+TIXCRVld1LCxOaXTXt+00EH9RxYuEC9g
Ikxfo+XCClGt1rfPIDpg8bTS9IwvHGBizwWZg+Al7T8DR0tpxyRUqv36GvU3SXAh7EzbGpaXK2L3
dOrX4w8nD0Cv2ZmW5dafh6L05+DkzUM+ra9WvnlhSwvHAT/zv7ren9o7tBQG3QGMvJbocoWeSiQz
ofUV3Lv6e37TiK61ue+vvC4nMiNrgNSu7Rxs+haMwlTt3bwxX6M+zSXbLKSPR5GblNoBfvBaBpy5
wRCCPUJnmwxC/fCiirb/+9vqvKU4qN0AI2zPB+t4sTmiPeMuuDHx9BwnaJuOmHn8swdjrD5ToqYO
K8f9CL+83X6BAGhagEMpORbsVl1M9cutUl0oxS4beAFof4dAPVWoWX9IISHXacYOaa+NBuEjgSO7
J8P5aU18aRV+WOlAZEULx5k05QzqWJBVBEnge/Al1zOsYIYwOaXGJAjvhTyxIFFhPl2Z0ExKiL3Y
ji1aNGeF9TcxpbtrY2KUaoI1oWX/4cx+FCe7fXT6gyGYAkw8cMDiaL7MGUP+UC39qcPz9Eepq9+K
a+1n1nyrF7sDE2G3C4F1jvQFSEiXdcCTZayEzjbbJP9QtOKW+LPfa8OyW+5mXKaqVkeJ/TY5YK57
959yI7RiwzSmMwykN4VJ1spXsl/H1kpUB39HIfKbt+ibva5H8yj8sP/O06rRqI3O2w64l2mGaJ2V
t6dmaCs4idbBHXA3nXYXJlZfS0CMkQ+x9BdsrL3otk2rjF+h4Hyl4bnsjVXK1IRk1zzexa6x2X0F
0QGTu58kliqZPPAaJ7mfJMkdUC6tkQD1iLijlZYd1FJqsOaPXvFlqevYkzArVgRKpnRE1R8A/MPs
+HZSC4L4t6n2dyXZw3THbMRyC6a5fbNkSArMwEMLKH3fptXC2KZUx/U8g9igxHNSHyPa3rwlLh35
77y/juptHCzy6ZRzewK0Ih7udRymLEIBP/9Zzl52evRU22cWaFOKuSJ8WssU3rf+VqIq3LErrh0h
+Q/0KqNTmxIKLU5Oy3PQf02iCu33uKb2ABqhAggGevqSu5AvjQa7GGC4FkSIffB0LOR378zMZJZx
uetQ1OuQJbmJE4YIZLVMkFlq/gowGmJppL0+LXR7jhE7UbCDDKWvC+PQLFgtY10xdmNUh2I9Ny+5
D+NEw8tpRKPuZIuwgRVjk1KE+1u6RRrgDP8frwOCzRfvgkWOYf4yojoJM275PtpdUHb1lraD3nzA
MDy8YYP1dQp0WcaGtp7zPAUZROY/Budqr0JeJ1osv+30N9UO76muRSiIJhT75cuhcOVyA4+sAz4t
LRgbuIUxSywUXarrHCZaBdthpXhr3VqRJWC0dDSo3+Pgd91NaUPib5XI+pxhqwDtfqqrNnUa1tmd
804r8sYhPKapD/9LKGb/CGNEPEMnnrXEsJajQ11ANVvL5pLUWInOwVaxf5Yvk9degue9QtmEAr7y
5NXvmhxViEoiMmjAaXceAVBs8F5hSIeUUypn9XDRLZan8CBVOp4BR/RpdJPp7j00xA4T8jtP3LA4
3RmhO25ZCv0sjr3cWHx4j3BzOqg2SmU0qmFES+7cd/4beWh0X2aZCy0bZ9dxUEEtszt8mDlu7HEi
Ipdvk4pSsIwzg1b9Q+p9hit1S/szbJRXaNWowAKEsnWd9/tCYqtkd9sFUPW8sIBl+yIOhK0TyXF9
+Kk9eZk3o8cGGUXteTn6D/iN0BbI1rc8cn3yMScp2Kya3kTacSKz1L6a2TLSPnbx55WPbRIeZ485
BHUeiFFLyCTNZe2bVcDATRafmTPq1u1kT50GDvIwuBibCrAYwSY91rXVU8gnozByBukX3/uNx0iH
3XldNgRUSYS35660muxTK72yWJW679zuJw5QkM+eMTQ9a607K6za9WJ7Wy2Z6UQ0ek6SXHFXrGvz
thMd1UrFw39we0BrCRPz3tpJekEEXfFahed3/PpcChEHqJ4erVGmQoMtJyToeOaONcxIdx3l/W+1
QYNwwns3PYkljWs6I2kBKRucP5WWRwt/jGVbDL+P3n07Tx/vayHJdWrlwQMODacNQ9NsHw4L/KA7
lMn+k7hd51hlrVVf9KkG1/qbJmQxx23iQvfCNuxww+fbUK9JuMLDu7oCUsLvd2pQyiIz8TbGQSmO
8Uiuyfw1nnSbP0t9uAXVBFzdWu4HUIPAZwxy4WseUKZC0g4DHLD+ROe929N0wpc7ERHC/A7c6Lsu
nkQoTZi/yq91wtIZJNIGqNy4/dgAHmhe7VJQEPbSWZoysKtA5ICsRHHi9KnkOceahCNsknR23Pk4
jZW1KZAZ/clpNjkxq2KyLMys8mHKh7hE4Xzf/rKKTuQwFSNHxIdLT8F0PaaWxl6MspfK+uL40PGW
6PkCo+MLUDbGxk+nSLYZDjzmAPqIQSGOeTH5dmwfGpiJI8/1lQ9Mc8/dS/NqdCDMVBGeagcZassh
LhTgGsCT7lJSyU9DLLEcFtMCitOyShoYbc6nmxpGGZ8sNKjXGimxYimwVLVsi9IZGvrRGHlbfS7v
saV4CJt5Kl9jWDn2Z5GPsS8498/yAvoL8XxzbnPf12mTbVmeZd5m77hN/GlXl0rcf9IzX4Ow9ZgJ
A0jKz4t0U2q/5Ufp9sgGahmCAF3ZhF+eVRfUspW22QtuB4WN7HatAaIX1g7zRen4FAVA6EhcgyQ4
zKBz780QG9GSboMFiXmfS1NoEK9RD/TEgL4NGaSs9+au+hqiGOoDWnOjaSO7FdRblhXsIZl6ACBl
uaj1RKKeZEPp0OSOX9SalD1kjcSEzDsmO5Oigx5jk0s2z6nhFlOTAMF08z6agmrloylxpKkD+PHB
RDKE9ws97GWMgwpkyHZHIllwx+HGSDxbqrzYUNTS8uoNmz2vjc32/IXinsjc9HLDRnGZ+FW6lABQ
nfLRxCJK3iPyvuXiHYzriDcC7uxloXDwmzIMB+fBHz+FEsaWeetXqG7U4i6VghbMhxcLS4ZaN0+b
6bJlZoUnW1ugwwDoP5S02LHvc4PNIMNjnSZJ85PNOpm0NGIu23+dDWdYPIoi5scUC0lubye1VFAn
pMGzckX3zMFJINZ8R+RqmS+vdtqcYlupW4mStRVGp2aeRA+lZLv1Y4W514A94DvAFG1wCn51LGBb
byV5jY45ptBBcaS9nEu7FqU0O4PmEzTM5fQVBIGlO71qlcETCqTatkdCW3P+SeEFD/3pPJ7+dxdx
xQhgmkK1/8aNE3pdV72le3XTGaXVwO5Q+Lk+8DRgYBOquwZ6NTP6i+ml4C9svITUTYddii+3e61Q
BCz2KNYgH4eil1QQDkLHGsCutGi23KwxQjVvxXXb2zwccBznibEbF68K6jvLPbS+SWfXaTMyysEp
Bfl2LA9BAhUtf/DwMdCrOMmzfQecHrqYeOuQkzV3SxPosu7zLvw21hEeSpbIxELX3dTwT6lxRXIY
NXjCx25WEP5xLSH9A/B7ketq+3/2t/01isnwahf3RCqrIXxpuee8drYdAzJlZDljy0nS4id+FDRr
gtcfledEvHuP0jirExmCAOsu81ouz4dm4NqSSW6IaOfa0pwi6cddU00dUsT3dtx3SNZeAEaB+jDc
AzwMbnhH0sfr08aIrqShKAWYkAU4R/ksujB0tazFzfNvrOGwcqPu4jmqtvuYp+uQQxlinnbbYFYN
e2oTH5ufFje76z2kyM3nVTol368fkViG5NDKsSNp877l5OG0SFP0ygUvFcziypJflgL58zKxQx6+
/wwYxnGciM2lPmJtANeJ7Yn8Clvjkh6Q0it3qd1wI6UzLBfcXfiZaciS6tzHtybOFHKsyDTv7aeb
ipxGWRXBchnUHptfhQ15AXjIC5kBW32cTzF/9zS2Jcy17p0/a5In/74DNbNXFixeasNYIzNUzfTD
8PnmlHy2+M3aIHx6HEVtF375w9ujJSxqCDPHflETErhbRw9+UBdEtNgcUjYMB4a+o6DggkgKzioh
Ixla5cnrZesmSI2gzkaEeMURPAReyc4P4kMsJAlh4vBrpWTr5biyU1vt/4/DpMTJfCnHvnjW/t6T
dXoeo8svnwvnHl3iJ/7ru6PhkGsgr2nHAfEEcA2eDYAFp/NnvLlcVUOKf9zogdD0rHgUGE1J3kPk
ahteP0w7z/p25V1Zurzq9icwnMdtjtqNaTzKZSEWP0G8/pdG/QcmqH9jrAc4mutPOgon0qxuRhIo
1nvqvkkfMP6cbWans7Iv2mV3Y5yHtDffuF44WbNAlAhAsTkhztiP/Fh7j6LVg2uQ2xgkjtJXLK40
7XZIHWiETouZ7PcatIHOjC+vcOtWjrwzCa+7gZlfUxpHLN78eNnBEB2K7r4JMbCvjjjuepnK/cfm
bqGPmlY3wt3081kf32P+LLOcS3m73iAztDAde4KcWGk4v1zcK1VZFxm08nNCQRGG5kEJcbu03GKP
LYrdUgVp51Xi/jYYQv3yXlVVF2TyEot9/rm8XpvVSLxjqMaQ+IRjjeZIj2MhI5BJND60EQRMc0eW
56fZMd5oYXCjNPvLElklk6KeK/IDX4E3iCo7/q+X6QjrEf4vtcLpDyZtKakji7XD67jBR7RcotnS
MWpJJTCWyVMGE1tETkrQNEL36Aehjxlf8Qav35uGhbOTyZd1/XxaOFKGUtAzrM09SNYfuh2q/FtO
firPsoos5Z0wEWeFzK198L05/Kpi1iayEslvIBUWUmxk35XUg4+Z+Gnu5Dn84K+xgdzeKAmRF6Wq
ZckRjEQ6wQLwJET0DD0XLLlbKzw8s9bLfv/LbYH82U/CD5vZB1FBYU8j+fP99I+ielcOcwJhtJK0
xVBCAPLyEFq/ZwQD0FfZIFO/kVkpAPKHLbZMWoRwfwuYQIqoGNDMOQna3ZCTrfxcgCTGvc4iVZZg
3unciMzC07o9hQJNetQJuf3UkxvesIZSPbvD1zLFKB1Ab/eCqP53PvcPWCe8/ALnmp8IKaAYOgWT
Zx42+eMbM4sZngbjjSN88LSJU/MzI+ZoFmOZW4nYCi4DqcTqEOZx+8ul9Fo/eWU/7+6NzIIKXe2u
uQCZa7RcjC8eY6Yb8HZZ2fRQ3r/SwkGYZiKH5PQSyrrXDm8icSSbXUsqPNKRtWXM8qgmgvAqaiWU
b8mKFtoo05lnWXcpwsprFxTH1DXKR45cXuarp4AReZZvgVeeo/EQI9wKEYGzNeG6n284oKaBp2fv
FcuWt67eej2I+ZmUJ0wf1pmucv9C82Af0/UeDOX7/ORosTsmyzuhi5NN3njSSAJ4vI0JdXoz8Mq/
iqsVhdcan3OBok6C6GbH/iQhoI0JRX9cFDj3pMbPGNwAS5PzS5/RvVYNl3cafLXSjCgkR5qzM21T
KvtgUW8Xl5/ilDNfU+1XBELVKDnEHfmZAXzTnzor26pUyCU+Dga9iqqwybiPwaAgcJJOK7JJQ0pg
HkbFrZH9mCZRZi1XQgRS4YkRlcIZZ/HxLcLMDwehD1zrgqXCfEWSI4IBk27WKVlOwxmf1MK9Pz8w
zuEWGxDukZLrJwE5YOe2ZOMagbPsQpsKliY8DpBftVsym1erWwgUVKfa3T6NEarop2DWS/t/kDF5
mGGGh+6eUjr9FIfjnn64xQTsklK0WkWS6XsbmY5TGuvA4IqFuYiCn7hfRMik8/RLfW+5RfwIQ7X/
edIpV7S1sTgKwVP4O7eRHn93MRS9LlZG2U2qYTLEl+f4vN9sbDBw25gwhD6/aWLEXfNHATaLy0hl
Nzs5dbKqtI7jEzMriv9Jj/9JK/CwwLGJhf1fH6zQICZaF27882whlOy0APkkIdn+c3j0oHUUHUqv
5kFQOQjCm92F5+Eh29P/56c+xvrg0vKzZf98zmC4KK8V72MJGmA7uNG/M+U10BTn7FultbLISEKa
hj2iCMhBP6CZqv9vdapUYJGL+tB2/gZ5eGI4qm2r0338lqfGTlQHgkgOuvWKrIe8nTiEpOsLiabF
VRFsryds46rDCnjv3olp4q0WRw2vHUi9ca1gVqeqZQLYdyb+XWu7WD3Y7nNZwzJUkeTwL+Xa7RtK
vuLjHgAgL+SnLfSpDnWY1EBCardYkTARYAnqR3uk9f975KDgqGeLQnor/XbxbWhjsz6eHub+Mk35
UR6Jh+i3jHnnkxax+O6v2cyEIfVw+p7inHS0S+EoTkGEyytnhsVkSQyJkc6C04EPiL0GVe4I01QR
NoJ3CEigL/Z/xmbm/hmjvLzjcVmv0+IzzBNUKvJ+84ChG0uFP1h9LhWUx7BF7AqRqGhaDYugMLcc
TatZKu+E19f2UAAJNX6Vm2Ivd5WonTzt/ls0uzwqzZi4jYDLSbp4yfKr5EqjY2wGjm0Yp/P/Y06F
vvT56reS1Fs+10rIkLLIJBedqHZbmkYNbuR8yNPI/Sjst9dW6uOAgIePY8ZlSoD4tJWjLQMJLt6b
pFgRqc7/10tDcYvjahWu++rGhf6mjeg4D6ssq1bFrYuKTK1ry2kQhjcpB+Jc4qYTla6WLlfCvIPi
VSjw7cI8vWiDk8v0UP+wClq7PSK8WDGVvhtcN+aKDc1hB/LUQriYUqqImIfcEfozndgYTaKbxKi0
FdJ1tOQSz51mE2PhEXUgoNsyEzGVlVS1QcUUeizw30BQmxf02TR9sP6MENRtFlalPH2WE4rjurdI
Kl3MeLoYxzyCGU/esizRbRWpkOHiugpCijNduKeBosiow/2H0kPrCCn7PxqXI+5RjA84obyBMrzm
7xzY00N+ejQ3a7chFrNBb18qZNfX1/cLTquEARUdzjemYoyuF1fb/vpOzxt23V7IJmRru/QOmfBT
rv8FSdMLOh9nI5Lzt6ImjJ+ppUmLIWnretM3Du1iTcxBEbZPepbPnnXhuXtsIy37jwwX2Ti7QX9V
5eDvYVydtnPN+dWZnuxOwXuahfda0o545XUhe9QvD2e2zPgEHYH+yFPIlPff+30xh2DjuheyiK2F
Cr8xTtfrJeVNxFNSdd1F/28H93LK6v7K8d5A7+t8eIcAOayOLVvqZ1qo8IaJSq8UHhatpHPTar1g
0lrT1bMQcWTMFDu+FpLQ4Ou7EWNdUEE1dIx/wjmxvsjJeR5DXfWpT1gDsK4sBF2ZKnMk9qm3lhnQ
/f1+vOMUZc7KDD+noC9qX1bgCvbGDvJkCP8gW/H3gGepxoxBVp1eouNI0hQ0peHTAoKoFlqvxAtx
TSi7IlXtmzQDXMzGxRAbOu/K27dtLHoLQrgasrcN6vzQ8lStDrlt9BrZ4g8p+QScbefgnz8D/qvs
rAcaEss8jCNsQ3pdVNjz2LjcdRMmlPf1Need45iMl85FhKggH5cgCK3XzIrXPD2k5qF3QwQc4ta6
CLRG5a7zaVeqN7O6B3NfBja9MBje5o7zRmFL786w4MtAbw903m9kO+HO3ybc7pNlUHYn55h5ArUU
MpHlq80Zm/z/KGAC/7a1tsgV+SXk4LT2pbGKJ7cCJq1kKyJi+CGCiEObGXLihkThm1PNZNRXKF0B
Fr8t8h5iTuzulCEb0t4cRNHEeev++MAfQ1w5qbTmCK5WtwYArbQFEeWm02rUH5wuqOzRSu+pNlYW
Tlq6i3MxPlygmtf326kB+uH5d5qzfOwd6NDX5k6H2FuDkYZ5LNo2EDU6grgFcv8LfWeTfe2ftiiO
jVx7lRBo5dPi7APRLUSQaCgFi7YRNjkQdrX2f700tBFuPsHS1JbSY6yop5p409xbghlHLzHCnXeV
q1NScMlc+s5fc7/dC1dY26YYt7K6leSoJ8ZbJI88chjf2nxv/ivTYb9afm740xk5rRzVGtRFaVEI
s0+Es/Q7skThAZF3f1O+ipnI7almrvXqhoJNMIVuxfQOFZqZM/cVTLyWB3/DGg++NPXSY18BBCVJ
3uxwlY/dMQ5+ESS2SI3OlqefnhH4S5YpGH6Ih4CmxsKYbys0HnWEwvzBrixF4VBYM/HjIW7wj69a
7xknmE0FJNFh4usg6r9AAHKmZT5rNhentzDd00AT5xA3nQ27UoJJL9mPqHryqbdS06nV3nbi7JkA
DvaFOu4LubFw0Qfrs0+5t0vOQo5m4M1hTFhJq/NzStZN6l23RCqqJOw+EwlPVclYAI6Rf9qDi3nO
Ju+c6/INd7fEU63iJxjHMiQ3vDReJFobn7awC0JOK8+NnGxaLfD/GKMgLWslfBSwp0tGq3NUdZ0b
i5eZ4nsr5GQwEHuQWXV06waUAfiTs1N48e0eYJ4wqVR9qlTWGr7dCQBKpK1MjYL+DTeO6Nc5fljq
/jMkbqTixo8wbi1WNzkT/pc4SQYHs0WymWnR1Xcfqroo1Ht5QXzXqYCcsEwVyVMyIFUnPvsJ9pdA
dqzS+kZUdSO1JsCB1Op1j99+rebgEIgw/vPx9v+9dsKPfMgr3czjXrzjnkbjwv8fIKNBvjndVL6X
2t9Gn9vWX/Pa4TSzIoD87lqaqovNYHqOMsXwvM80MPORKtVh7S8RLgmCsGECoSKrBwRmdLHeO2pL
w4z6XRftA/0QGY15klpDkPdlZLDVw2csB5RgOytQx1LVCqsQU154LLKDKdITZQJ94DUnV0arAqAj
v67qtBtRj/X8dVcQHf9Vmwz04zBp+LcButZVT6ix9Gkn61a+2Zi5en91FAv+06Cmya1Gpa4H8K2h
P/5jot1HgUcNFVy7l1vb9PgCQNZ6kVMISX55M6gcqvvwx0TH0djZ45tkfW84wKuxLUIdKtHzbu3d
KucvVh7LNWrL5WHE8M7G3w6r1WQwL0etl6fdWuHzcAgqjm8jAbWbJrJRr70zWW8Z24UWyyqCUnNu
sxHQpOJmLLHCY+g/xQudGOt8+npZCQ/wmzPaU0T/iP2aY1vM8WCBRl6jRRAB8yCEdmQ2mcsfRas9
86bjxmE+wG4AzE/jP6nadSrUgV7HtxGXg5M+uRwqh/Zy10owBZ64rkp4xIAINyM0VFajZRtLRK5C
avgkHAm+pfAtp8YdWZxLiGrwANg43iqANNbYBEZ+STzH1cztAkE7TFgJwvK5wQTJOKEYkoMLpBJz
4vtjS1T4SMrTtPHHsrImzLse79hfcUH3MKMSjumeYXFkhEjiAFo9OwqyH/VlMXqEgJBzmUDp5/j/
5pol0WAwgp34BFGyOKKoUCFZGIArGX3VaUVT7JMlntEHUCegrlDFgGQEVnyt+VRPcAcFnFXenmzQ
9StXTny2DkQR9+Ve4Ij7lVm2UxRwNK93rYq/386BX66vAZnaKIvD4ry2WY2Z6+r0QUAf/u48Xo7i
MQcwK1SB5XPbSrlaa00XIOiqvrD6uChgJ842+arPHtsrsN2jYWIy1ZOn9WlTr+94M0u5K4SYho9M
Dqu/9eT0Wa55fIv27AY/5qaGkpd1ZxbmF6Ob/VVmV/fkTde4W3iIkf990yHjMVkhqs/ePUJ22sfN
QcxkK7QVh+sbXk6hAFpxKeTvSjEDHMHPPhlaGG07nIkSHLg8W0R6RuQ1ctvi8c3NkdDs+4anELXm
24htH2ZMGdDI5QFyvEjnOzI32YrXgRFvb6ySNnqWX063Lv/YjXyW7DLWuPj0XgwIKtnVCk3VZ/QE
pXHVXjDBReEvR4AuSIonFDr6MqN1iNUvcJtC59Y6vTrt4/29I57qiVfbS6126qSc1WS+E/4F7lLP
+3WCJi8qKmwgTgJXtHrqgbdIwT/CwP70QN9iAHvNcAEL+juHy+9uM6NA0WcJfNmdEVbVYj1BsDP5
1/upYgXO4M044UO3zhKwYM/i7FSEkIFV+vaOCihrkS+x/vadfwpIaH4HRmuMGTa99gmjZvrOan9D
kYV8SsCf8hq1IBcCmyrBupvo5e47R4UU1EGflNMFKbAJHp57WgwZt3Co0DEa+l82yxd/WMoIUcbc
Us58SvDsLnnQPuhI4W72kbBgU1o3HKe7yUS/hSoD8EZ+h/M4z9uTpUiw65GscB6zxD4PcKnOsz1x
ZEHSgqhEDMq1Eo7HW+Z0+ZdG78HUqsCNO1eA0YU2p69yw8pKJ9q/kLfsMm4qdH0DJQdLOzjtZsEN
uOqWLE8pyJhmJQnehHFupJ0+MmuKcUQHAjXdC7egQXQYJdD3ffQmirqa0Pj0xDgY+j+cuRX/CE82
XFbKiDa/81bqu5YC3JNTckvmXbqQ138BE5rnng2sUZfAVlFdITUXN6gNqxlwV33hErL3E+c61emV
Dq9R/TcX64/pKaaGC237jAaIc6SqJzpfkmS47+HOfTcUj1k4auQgHfO8CAugLVpEzHdu7Pg6z5lA
1kSk4NvTqZWNWipGBFDmrRdDabq6Qu165q5P14FUVvYnm7ggLUrU2lt0gwn1IyvE/otBBUB6ARO+
btqIIlUp+pE5DM74W/AtzYxz68xJWZ/Msrdx1yTjF+WMaubXu6VkdGLqIklmv7RieS11BvFbkR8u
Bss0xL4efTLC+CbyIKVie4LbGRajgwy9crUPLMOiEf8sXyEGH3AdiWGtHuK8fPtgEqRUtSJWjrrs
mBL6xR7NPTgqbB1xMlseZ/ucTVmA8H/TTecSaXH4nq47SWBrqffDmso5OW7r1j0QuLaI9dycAl1I
8iX675DjXZANYjasx9xoxkkWJ381527pJCIRfv/JzWlPjfu4dQQmAXEv9HaeTMf7RA57fhMbDNpD
s80Oi+zSVDZH9ayDtr0D1M4GmM9nTdjpE6R8NAl0ANeKE4fMqUDAz4QrjLNYUkeFaHeKZb6szobO
mDl0X4YO5oS0ANfmTALhIfmP4M/V1ToCIwsgWXF00VDTK65lyMvNkaU0id8e6ouR/lseXShMgs0T
gQFyXxZlhKhuINY/e7a3THLIx4DsDB5ZfB/5iSad4bqf8sv5JwYn3KhART+eEr5isCSztfewcQP6
yZksbCcg+uQP1NTYawjcpoKtsWbusw/LSiD3B/fh9r+QXlmsoM8FjOS6K3vXOpLOj5W1TCFJ2N+K
kFC3GTWzV6MjfKeSecdpgbQtBXUpGTcJntfVI4ZsvmJH/ohnnqsFsodV4Y8WZ/+DiLYYlxrb+TAQ
vybOZP/Fhtntz4f9HF79mRZ2SMwCK3C6vc88KlfAjF2r0k5ST8AJyuCGyMDgPaq5TeqKCYnlADYK
OPrmC+cqZSzs1B10SIpayHnAyZhWba38PZg/PebsrsJfwcnQzK9Zj81PXJSkt66c28VW6du5Z++6
bX+Y1rPZwTM35Ho29KHxF9ODEBpFF3jNKmaduX42J5nVXqW7tz6vjvJq2h3pnGnvnQZcIhc7uEDy
6u29CTHTnOF5ZiVFdtBqzjLBXrF/SYRtTtF7h4PC7/VEOdB6i5azR7TAXxMItOk92m8WYNa8ncje
bOGFr2/7m2NS8xm4O40j89lJW5BmWs8J+FsFoxamNrfMwHijQJRlb1SM1eASFiCroTKT2pp6JTRa
GKH7vAZC2/pfeoARQfxHquu1U+VQUVHHbJqq1V55vwB1zu5YF4xxSA8DBuqcxpSQsG22fUf9Lqk1
utwFcpzo7BZsKgBhgwfVVSKwGOZsiV64KaaP6TKnOo6VhVG3XHlcJPygP0MtdlN6ijUM0jfz4MD/
bO37y+rjWOIPvpSjsCPUBWk1X3VNPyZA0PMvTqBzsBMWRpHyyn7fUgZ19PozXXrwW47WZgNe0I6/
wdqwo3Ws+jAR5nDrszCZBFFyy0BsuVrBdKrc+NCXEJbglueu+GTlg9OgqjEUIT1zENfmzx5gg/gJ
PcRC7YF8kEXxpQ6hjfMglJwUrFWeNFwxyx+NHYqCJkYfJ4hhWcDEx8twaYWjwRT9IpeERpMlblY/
IxU7zxchREuq6EQIKWMDUuTAs7SrCPJETKeMMp9qqNMIql7ykNQWr2mIXcSGvTJMtx6y4nYHGFyR
WT4okNwYL+S9gSDuqc8fHr3XdWozYMFujcSoPzhpIAmDg8DFJrfTODSKdc6DyXzysY/aHEbtyMkP
19gy5ET7vjHP/Zo8JojuuZRAR3UkEzhReKlxfCx/p4Aug/kA4m9yRzJ7DlJeDVr5//mdUPEL6LxD
TOGG+mltpU/rduzRRKxx9MHWgcUyMoatNQbX8w1QtoI1zMGkbLeE7kg1rnqACRSSYqpE9PD0Ersh
C4JGmtV4clIK+HAI1v6/bS+fMr/1qy6u7jHbSq3AmzQnj9EWmEHUYTgPvHRior2j8crEBusNMEUm
zSODyfsh6FryUGWmgKMBuU4wPtYwR91aYPoMy8WGaiExAOuEERs82sQK8k4OtLZYMPrKni+abeUz
UxfJLSmGCWMeg77Q0Yh1U9J/OfcGXGFR+i9TsmzjV4ztPOwnQBkJ1ycHUzL8O6s1isyT0rwFueDo
5hurOl15pJnzMyS861oeIQ5aShNdCaRqkUv3C90Hybrld9fpUlXMVt3cEufxTo0BTVNkgBdpGudL
fW10hkdJGPXTCmArIXAEO3m/7pl3c7MS6RH869A5c3GCqvTa7TRr6ITl+10KSuLm7Xb63066nMmZ
mdIEIuP/tvOxMzbRNLv8JzlBZCcTx2HWHFqd9cRtleIm4yjBI0Phus1PKRGrmz1ir97UFqMNC8Om
CoLv+14Gq3wNRgJiwJRI0nuF+dy6svKmPgbvaOl9KEIaLzwYLAsgKuGHMiSfFlM3TSz+WEF/HGja
YiJlA1odUcmC+Ce7RCPk0TaEg6cOz1YgG5xG7PCtmwqvYUzzNCVN+rRHzfHurQ9Z8KDquiK7ww5m
jeHMX4DTpq9rzHL0V31UWFp7jmDe+XTMVe6rzVLgvHGzYSTJqEY76VS2HU3f+MK/0dj3bBlObUrh
MonnK2aBlVvcRfKBz10ZSvevA8oqpGocnVShtP7xqhbU8pm9juPWgDuUL/6SPVNN2L1Pln4C56F9
uh2e/ZMHFxe54+C3qWlPHyfbm0oyzJy3VzsxQ9wGrfy1Y7eSbnN8hlDTEbR78AlggWF5wp4YiZD2
MjG9M0PKlXADiY/nigf9Nb77OtK6xbitqraiCrFotRkGgRZvMGGdXCNw4QKAWV9J0QLT1Iu0w1+Z
lEaV4hTkllxtqImOjcvX6Zvu7+FKxhMJRF3vBz69Dk85scl1xAuJq7E2ePqFcUS43b386hFip1zH
p7J+EguimpY2bSk2EUvXfELLh4XoNQR0Gk9qrGKNG5gZLFVH98R5DjZudMB7kxREe+NIUXpK7g4W
Lmc44pA8jD9co63IYcmXzc06mIqeXfZu7nbT1rHS+D2ajavONbNkYYc2wHif+BT+UG4pGUBuFDqR
pUiCJ8m4RNzXPGcS3V02PcwTBeksxLd2pkHzzNRLcOmDgX3NCbXNX1QEm4N3O5DjP9iBFqieTl1P
/cB/SHl184rAbQJTpbV+1srnLaG1AHzGyY66dhYJH8p7/ibO4S2Th8YuKHsYnuujZzgLc461IKIp
gOHbcePT7d9HPirIFamzFKgToIPukdMarsYcJFOhyxsSWrV+VW+hWt3W/TkuncSTf453IxwlQKho
j8TBwkaG89x3a3mLmnqtpHyOROR/4YZx1Mr7SgApfvXRJYz7sUP+RfHFGOMmi/wCkOoZp1ff7p0u
Q9NBz9kR5cblJADWTqSkvTHlsBMOk0l3vTLEGwfOpFBZFej1NGvlKGRkAYZWz5V//gKKeelQMH7J
S1RhCicjGfgeeEy3eW1QEY1vqPUnNAbLUrTtY9hgEMEN3vwe7vGKZ7rO5lgUlV5OjtR1NjqyHoR9
fgeKj8AWi7grvUxUS/ggws2CjpEAAgBAbl6xUKlrvRQJ2SXKOHnXnt8ZAC+2VkCFGpYYe+YAlYzK
zZuEw0/6fPkumuCHnNouQt5bu7Hy8VNYsWTHb/2WPT/iOtta2cjFrnIAodSfJYsuYbhvK2w2iztx
DQAHa7QvcgCYB/yD8/qK4GAZwyy3EsV7uZjI7+x8f7voiJOolK30crluKWMX0UhUcSsL/Q1dAclZ
eBOemnQykYe2TAAiV9y8C7L9eDcHiPyqTeKIxb11p6qivmLrGoCJdIsBw/ZhVurDjLoO7e9wJYQz
2ekPmtdZgtbNDyxtrkBDG26PuS1qB7/P39yFcp9Or8hiRF2lSt+VA2jycdBcNsPU7fynITrgLYcc
6ZRjQ6Alo8gOv0YwwLNZf1xNZAUbhK5Ph1ed7MZfGVHN2MJzokDqDt6tT7rA5etWhGOEjNhEp3Hq
1M+lapWEfiIU9KIrkVO578LmB6iqsBMGfXNwQO4GOJwIkYVCzjUSQl2ki4ao7mTZAy7Jc/1DGUdx
fjD506Bs/kU3gAn+xvhO82hsn7i8ZNKO4nH7vmuRWwz1g9Mc7OWeLtgQENG6DeEH9zjTmHDU3XaK
L727Ym6TTC9lz0RUoUAi2VOFNpMVd4vIHGZ7J7QKs7eWZdy5ZKAyVai+oXjH7+rILaW0AZ7Yb1BO
KOLV6LXoh7K/SCPCR7jddMSXNqycT2QdalBA9LPt5MT8UEyoiRD84tcZ87G3ALq43DXlQ9/aM0lF
/k+7TJoW4ZVR+X/aViiQt0QGeUZ9pJ7t8+D0zxM71MqwQXrUu6EzCpt5mHIhKXF32ZHxliQ7ijTc
EnK9usJHmmykVbyPmhejKrHfjVpr0kK45gbwAfA1/7TmpZ8fuAbnng9VYYdYbVUYD+kIb/nkNwXl
BMSfF8Lt+uPmgNTmueboyUVeV/5wZ62c1aiwJcPFfSuGXsrLDNte6XLpBb3VQ+0ORQude3M5rhBE
Q/kwXz3/l8wtU6e9mfYqYAsAfNeOAFX5RMD1DURKr4ukHRi2FslBa6hkxHj2+09Uen8UJb8HxBOZ
/ondQjUexeEdQh17sD02acGb+VmCjBLY5anCnW3VRxJ91zAuey2ZDPI0/1N/HcG+xlvZXIr9TwH8
pgBzbzN18ApO6BgYp4UdrjCYyu8PoEE1ZsOXs59+Bn0d15Y1Y7MFDl3mKBOVZAtDH7AYFSQigJJz
gQAT44hLZcVgfwwyybNQK37ADwejEQ6fGUgd2sBPavKagx3ebGkhWxnyOjMX+0BAP2q8Qq5sQne+
7tIzGxhxqLuNfQsN75PiziBhD3aYFdHvljXtJi3gvxmhg917hT4LRucBcr3V3fInPYmkl0dDp8yY
uwAkJISoWKGMf4rJpqsO7zoUmz+cnKDXKKPsOGrE3X+Ga4hWMUxG4z1b6Zu0WdEOpSRLcCXDMF/K
1Iqgc/2sMy6/2dmHqRfRCkhSkt0NSk0Tu+4T5KZ4yhfPggOHEQYIsKsci+djghHL3fTiwTvGWxD1
Oris8SxxTPJQxEp0wx70PZuZsH6G44LcrQb8zZtz6qwViL9fWitRp4jz/H5mY6R2PhNR6QQP3WVu
9+asVMpvMGhtvpTgHEmODu0u7jvQmw936MGYsKbfthU0VCyml8RPev6Spc2TfY8EH1nEuOyRPILP
vk9EyJMTe3cH68rQx7GVP2H4R43Pm3/QVp//9wqIDszFjb+YwBvpglEj7iSOEnXcLMzoCVF/knOI
j5HicYl3PG01/G2kUWpB2kPea+fSU3Zx8BXfLn+MrxEU96mHRxEgRGV3twInt5P8j1wSeAT666LM
0r0srLzUtkk0MhZ8m3p7TidxsUPxuSCP5KqOnokq7CqOw+LdtEG6RDCohHjtaPk8WldQXUNAX6tL
EIKyG8D0KrXGKgW+AOpHMzoLz4h+XxCGiwu1X1zeDT0ZdvmS6ulP7OrC6mcrchjxDNVvPKlvbsfB
SOvfMm10W+cEn+nuIUmckq8VTSpqExD1xHLhMj8aFxJOjIug0D7C8im84cItF9krFHk8SWV0aoVe
eZ71E+Bhm9a/g8j4l1eg3T4xyXm3PlylNKk/DJBSN8Oqw4t+TWL6mBdvolRD0UbP/c6zGm0/u8X8
OT46PoJByy0lg1mxfgzK4AzYT+XKFaCHU2px9N0BQFdwhflH+7kEWWvsSC+kWHmEu5TkNc90VY0J
A7Q9Ak+XKiYvfYLChM8Tm4yN3hSPLkQGE+WRARKLyOEHWtbk++HzdAEJaCAYJo1JfEgyZAsm1ub3
jubdZ0ggLg1ATOKfxUbVNoH8SzQ91n8tp3m4QtpefHXG7Nt0HKx1YyE8R81gM3vaM95SwyIZw2Xw
rV0RvK+sBYGmMWYFMfjxVfofi95O17UEgLmV3iU9faWF2g27f2BVTodP+g/2xP6G2bfcgNjstSO6
rF2SrqkMGg6fnJ7EAdW9bvBe/1EnOfH8sTzZXl6vK02dQq7MX4hQi04EGyqHlKAMF6/D6rPWHinI
BPoebwNYIVgX5/vpkEALcq7gFwYF05/df580MxTQjDt4KP4O1D9lleUiYbvxTFAPgehqyBEaWYBg
9BYTwvROE8/1yaHD09Yf25Pue6XefKSZSzOvOeliXJ6HiOWsQizIkMKjJCYagD9OEh7cPJPpXjp2
w8Fv/AGP7IJoRTka82a5EZHgF6C3mo0uEgkhZJHjPKUAo+T8yYqRD/C6xIkfwpFBxVciSbFeGW7Y
cyQrzzyxgXBhvrjkOPV8mrDsigWKVx8prv+ry2tNoNh+cbNqOd5s4zYsxg+bu5SFqsTspZEfD9UZ
JEFGry+ngfdps3yZfOR3mwIMMSbXMsCAwZ7zOpNOfEUvzikk2ziE/yZOdJm/P/zrASrtI59YjJxr
J1Vxz3FcKMke7YSrmWIDx2pzh0IXFmZaDCPfW2uCVic9m9xjOekPQwhxJ7HrhLzz88G1cnxxbqMd
cqX0A/OEYPrPG5GbtsX4XCnOlQKVYGECGI4FLWdT2m3eoJaEejy8qDY4tOqGsod8EbAh6dENQudP
PcQjL/QyhgylmnzXazP71Iu8O7CA7d+1G11FvvI233j4UjqIbMcBVNXofBJ7E+iIVuNZ6ocjAB56
z+kQ6qogxbyy4ftjHo0Zt9217bB7UinISIQ/O0QHZH/HVCxKo09gUrDiMthixKkpshxZtrkI1mom
3s0hT3VUX6MKovnXlpsY9bFBU4BCiNWrVoCiisIHARye8sgQy/9E507rlf29+dsVAdPOpIXw8Ydi
qsEnVUuQsu4KztnHWotU8OMrnH0X8Do5+Eb9sM4RlrY6inbGMBX5MdRbuW9ZYIyXZN+x7hTR7Xc2
a8z++tpViA34CDbbvIyEZ72Kd0tgJFFTSEZ9t3nGKHRalG57AqCU/ijblocHxYVmYDVobgtgp5+I
HRd5/FIaZTKUQ9i29GvzSCWvfSOn0M8AxL+zMstfaR6bwk3vHXgw/dwV2tbjziZ3OSAY9cKO8MDB
yDTDh+h+tT+h9AxWQCtfvbX9PZlb6eo1FiQrb5uJgbDP3zh3uyuSRE2jd0D88Eix2LonW7Ge14AP
ai901WP3v/rk/HpbnQZLYroQbqSSMDeHnXc9PH4UoWmpTK+blV+3wsL/u7IU1ECcX1wZCIhJ4fyc
NlK679jhxdnrEm1mvUhksT+BBgadhSjA6YwwpjmNkqhYdWWahF4IhGVQSzKGc3XV4K8FNlrHF8I6
mun5ZJLw+l9E7r8uQwsc8/JPh1QO8x2OojfPbSuD7esxggr9SR1HNv3247+HwtAWVSFF1zzDQuln
HZbzMDGNikdrMBwri3jZbv57UfOeggHwvhP3rI5GatSAWbK+EaNlUpUQmGlY6ZDcrnLtICNWO5X3
vRVB5NuGqoOv6mJPXDgkO5dMiOchxtDtGvUrgpXvGyOwBYM3+xUTjByrCdUl4UYZ64964FFvYkMt
i7qaeE7gnwQIWIhHZfydA5Xh8ehv1Mc9O1gOu2lRv4zMzO5QKHXRDfEjFxfQcfLzOgBmj/1SAb8Q
NpWE+JP5d3Hd+K04V1QDiGMU1DSL81nPEK5FZYWfUAPJo/qKGm3txDismEUt5C3NUQGgsbRt/x0v
0KguYwSAUbmugnDQz8p6buJG9dDegry++19ceeSTwml8L/En4Ku17ejIgtUMKRM2CKd2J6yxV19d
x8J9MzhOy9RUjPYG7hYZ2qUGZC7QMXwGyLPJCeg9AWVKfvZm+urjT8m0qr2Yiq9Nbq36TNqiRy/J
+cHZEEvD0u+QNUFausR5nck0noP8ym/HVw86agdp/78Y1Wm/5pVt0jatFM6TvLY7F5K717WVOfNZ
0jFDb/s3+iYozb107Cq88315CgKFu5/c3f/c7VToX3ejaAnV1j/z5GrHsR/4l5kWeKV4qr7cc3bJ
yNSTCtEhl/JM6s6e8zcjeYi3cdsH7MX0RY6pKL5AMpy7E7FYCg7/UHr7QYEZkpAncOapPZ0VhrkY
8E5bzmptQvNj5Q0soQJJXm8sjqRtUIhQH/We0i2hY4jJnTU4fSiwOR+WYEDLHx2RBlnEcig4UAyr
CoeVNiqEZiqU0FIU3FFCGHCgZ3WoI87PX3MyUxRukqg7Evu5qrH7CuzLM0u0d3KHE1GbOGb56IYP
GYjFksbRGA9T9SZPoer10JU6YTBw5Skirh1yvSBgylwOC5qDmpfR0Z/LEETHArLMHB8DhswKsHm3
Xk2Rf6acsvy9tUnO3jwl1zgr/XWOyBT6umCAQurBfx9HAB5R52TojmG8MBVns/bDzG7pVp8aQWlm
HKCmDVCdhwzrZ8/b1hAzlWwro2FlhVYI5W8bEc3GW8kz0rHrrIuTlI8a0SDKgd5CjklDT+yz80wW
4N/BC56qZ/YYjblhPxcxD+EYbzQNQHsTZexgxHj885nI60O2h7XR18Yv8bagIjzdLRkpR5EG+3RM
68yStSQLaSo7yK6HFq4EIRGMkse4S0F+6hrYOIbHS4JhhelMUJ7bV52pOKtuNeKuO79+CGe+G0PO
gz9qsEx6JhlSy06qRe7rzUVlAz+sspGkPbQaH04sUTqd58Fb94I92N1eKS+o3XYPP0eejCPcUPDm
rO2ZjJ6ImfbBn2T5jLJFOmfoCO0+kudnuhr5quWKU/wMZywcnc8ogVo8zVqXe9903iuB/OrAQpb8
bBwnC1A9B59xx5LDiGnctPV0qpYUsAnxXHJupUnknkpF5LGkOfHRWeFGNi7elWlxxRvyOqfWgrQ1
dFpLIUMndZmMWmsneHbpb8RpF1XucC0UCaUlOXMHKtGnsTKa32gkkw0Y2pWDAN5SUphPgpaer/ny
4DZn8eeFwd/uty/kBsPWDLyCF+d4zdC6UOvokvjIMz3IGbGEl3M8TminMTwOKXvEcPZi5mJ+8Og5
ArPOCeuqEw5Ko55OrxaCGFvjSSKjbPKAN90nKdULG7OC8B5wTtAMgYGxE2UQJASocYw9CNWK2DII
krX3l+7kVMqE8LYUOcRWkaRnKN2KmEXNfQSVR6UXmM3cLpXM70VLqcc874UgOMoq3p2g7ceZA4SP
Quz3/fESk3YyKj48RVLYvD6vMYaJfTXoW/o0uymZnwzb9gW3L+YOJ0r1scSUIgzT+cHHsZ2+Zm1D
ee25kfoiv7kuIgooOXADUNA/W/mk0bG+1G3glPvf4xepoAW7qw/KdZu84Dqyyb1sHPPoS+sZDEkv
wdZGOCe2kMnCIudE/r3za0A3qesyjZqCWRjINIFe77YsL1J3pTKJ5wxTzCiYzoMzynLp9QGmpHWn
RJXuYihYVtPF3W2fdRRrB2diFOS3o584eTQSDhPNnel1T6ZJ6zbJKthzi/tYQeu9CmjJSfF9ZC6J
Oo+FW4AC4wlmsbQ53F2EX3Y1K4F5w60B3CNxCpTxzs3ZVmyxMkjDiVYvRmGWYElureI+qlSlE69m
KRKh65OwkJgzZn2fvS7cqs5IonvoYHXucy10p16ZyFXap/lyjmeE0cufE8CC1LGbU0QdiRuYV+Tt
6n6+P3muBFpfpg0kbiyp4czrB/s1p0dxOM0tNMw42XSIlMnA8cVb/NJrUQpKYTwm3mGAyv52ARmZ
gV8ZA+rYwOGHFINn6ljnQGGZ2BuLwiB1x9QAebpOoU8905MUFn3oXhI9omXbBaU7xSHtxr4Zgx3F
NJ8csEXFFdh/ghzRa9T5yby//3dD2jxPEpI1mZ8jxno8gn4mC/Ct1lkCJLJqM7Z5UnqOfpvheNjo
dmrxHBTaJMdEZMjlWS1z4Za9cwV2PnKJZum6BMutbIh+R/GGmFqABL5cNhJq3OlKqrwYC89idNoq
+PgCQDWEGwLVQTC9wEWrRK7KI6xdHEtrWqHsyrdD9i8TH0BOmd/nJgiAyhtD5+LzMlSZgcmMLKvl
hNQh5kvRGG64oHtDmzVLfaCsUwDGc2lkpSH39v0nA9h6nCjqEwM/zAC42wLR25J5gMyPOu0YErN8
krvr1XpbIdSvSyQF5sM91IYYvhQflT6tz82DTArgaxMuVGhFIVZpc1oeLOlRou2K8qEmRANXT36y
HElCsJXGr+mVGQ1AiyOP68JiUwx0qCaxadFC5x4rjfi9jaLSUkt6phm6YOpsbznNEfN08nXnXcue
9pXv4DJ+Em7PAuYv7/gy7WqXpM0qwkqf/gaR0/v3Dmo7saTzkTFiHmFGRNLJKMPK3fd+QfJ9unyI
WqAZ4VoQXoCcTmNea9B/AQVFU7cqIZg+hL1qvgU4Et1eas0k5YqUlVB7UHpUqRdigg9QJfRjKdAp
WpnMF4GfKCKW973ZvpU96IWR70h1k6mM3iAlBT+9LpIald4lkFFf7zII/VoBnpa+9Nsxq0dko8Iq
2a5I7HIjH+YVd9bk21eC+l3rTpU3kT1ZUWyG6+f3VX/lyog06IutpGfD/Ndn1yE14gSse3RE4s/x
bD3KB5z69+6yz3mIXDB0sKp1qh5FXeJAqzcdPAZri1NCdtscFrCXOoak6+6/XSlTnFDnPu0BygqQ
bEEmIJZPdxz6z8TySil39T9YFHFN09jIZoZh3OcwNXdqrYLWeZJSGo9vrQ7BFNcYSIch4iJ76E/8
zisrVVujf1bL8DdH4zX5doaDPJlp1MgmsgAJraokag9ncnKAvYeH55/Rbt2A2nccICLeyaJqR3qx
pIKpg20nbJjR3ZlNGeHFg05IcL0t53lebYLMmtn3Od6MF1unP7K+fZ9CrVwpIxeghJRhHb0JN8Xa
khh433+0Gskn9gSUTXaTLMakkmUry53mywbOLZpZ4H0egD4Qz5BFCP6RRH0qltBkjsTraOB0wXmh
rEAm1BVSceMa5KsCZb8F5913OAMyF/adFkau7th/6i92LViHiv3hS2uhlAwn2giShkuSbpxb9y+z
MZAaDpNiD9YgAYFenHsAHPkCQzolY0G4BzeaUSJFycwU2V1z8ku28RtyIwJHOP3O1DP6ovyDA9+a
WCR+OeamcFQIsPTBLjT/i9GPWSj6n3PRndkCsWcKGA585Kf3ES2rH7WGkdytus65fUUUPa9+2ok6
eKWJI+Y1d2/LPlhlIxmqXlYZ26YZOd8puDwF7x8HAiTgEN40IRiSROqrcSZ8NDMDQxuPxX4KCSbk
GiReobxSJ9I+CeWIBd+4HvW+T4iOVUJoyfLPecqhYiMj/sGamW8bhNs+RveQEPzXjHr3hF/d/dio
y4qlEd0b3ixbCjqMiycLn47y8snU+bFRidXm/NMvVcnT8wi5OAqfK3Q5HPLAHj0xfvbVkrn911ld
PmzYm6HqQ9aW39HRK1jjZ9Us9M7PObgL7R7BAhOBw+nh+N4SHznLPE5/ZAhjByCffi5/kG1kW8Ek
TADkxzdm4epRaR5T9/hnccYVmmqefcogToDIowmCGcDrfComnUgk+gtc+nZMdBrjGa9G4u5Wwn2q
YxMkjwhs6S1kt8CYLPkV0YuBWK8/0erRoJJFmTn7KtZaPQgeHzkVLsrBO8WsoFntjvP/IsxGqGHd
ColVU9YLLH3Pf4qVRcnW/adXsobCzlswTw/bl/qxy09w0K1OxxhwGCZ5kDerUN54gQ390n95wgzp
WLQJondDd7GX6QsWs9jfRbcwRW+Ii6rEcs0KjmEsV3luUp2a6Z8fvHwy5omjqKJoeslqc58cT5DW
IphRvZ96l3HawcGr/TAYSzxjYOTLay3tfbKzOZAS5bP6DArSXSC9gJK1A9yod6ALlr/RvXgifbh4
KNEGjM3vgr132VyApvDt/I+SpDpoMor3CN9FMHG1EoY5AfBpUUFdIFAkiYK4CKd2IfnyY2jclNnp
ltSX/1u10c058uKn6a74Gu9UruEO/P9kIoKmbnpNdjkKZWrRV9jPbtSDzcLzO4Qjvja1qOqvPBpj
F/t/reppIYcoBCD+xXf1C5c/6+P9XxcZm20t0eE24q8xREnc5NHLvQssl53GrkJ81vvUrLtzMDPq
FHYqFApagQM7iLwrvCzSoT0XHeAsYZG34V7Bsx7nsRetMBslxHFBwcCEjbKazU0EK4fh4s6UpPDy
dKMZ/FAOzyDnYk9oLOk/OAO5RSMvzjUpngdKv2nFtMTJ503ui6F9hOMtjPZn4badmoobRqJWGGfD
DiSLQofGaLF/8GiYWEYlsG/yx5iCmmM4BH9xdaK1MqfQ5h9rpOr+/6S4/1IextjHCxeyviO71U9t
DXT6yz9p9ALYGADDWSDLRzwzhn4GTcS0/TqxqB8OlmxjMhw5Dv9UI142BJXNo0NGjx2bBNUhs16y
y0+cMi3NFA8tuaZbTUwqktu5HBeJa1usKQyIB3a9pLHrb/MYJS0a+7Bq9XE4qvUXQEyIL0At8O7A
+NnLvSbRbaPdQ8wRMH5xGWo/Z8lySFCHnP1dLpI2aIBr2lo5wIZQIO8LyMEYg/TWbgzmcmjBjs+W
8JxBWnd8qzDOkj977LqGOwbuDuRttwBfC/OXhfA5BoxRfaVXhGu9/J4yyGO7EVsRcqG8bZ9bWTSX
okZHVMt4+6YWmrHM/CnZMQWjWoWjPrMu6XeSDoDDpwzHXklfXeqfngvR9ZZ0SQFNr5+yxdtNHc42
BAUsAAwjfNR15qHlh7TSjc2LHQSn2SLnn4qzNxleH2JAGl+er7F4Vp7PeAtr6TWUvK8pXSsIE207
TTVetV2TfAhYBzxVbguPeHVXu+XsR77NW3HeB5iVsWOexmfDAbeAYjLZkjtiDpHhgVddj+Vsbgb6
R/J0TZ2K20Pk/1+Hi/amTPOcnKl4E3C5KAsMuz7qrUdw2ccaU8reTKFjA5R5x4u6PPgvzFTYQ7BD
GDaw31oiYmrNA+39Q1SgqXMJ4Ii2kD9wk9crgXe2RYPdAfNAk+cF4matsSDETFlCm1m/styZMuaf
WkXVfLT4gwnFnop0K952N8t4OXLaQRDhOAdF+xubp/PLYbBvfNnNSoKCVssdyU4OMcCDdzPUugVw
KrngOfpoh6j+vriblIsWKeEQWofymu/7jjb8NnJUH3WQ7uFrRhS4GQY1P7wVWJSKxxoIGobY7/qU
BkwoYPcLE/o2jKADXrnpUubCc9Vf9fbUbbB/bMOa11jrFq2i2v3LKIR5Jqtx7u0Dypq3RRevi0y2
wJFtG4BhkqpaZp6Qaj97RZn3mnMqfUT6Eh9jsu4kCX3wwLbOMnMLDJZOjKZGY9Gy5FZPt2Wn84bl
sfZWI87iQ8cstQmT/w69Jwcx22BPT7QXp3H7a0zt/E9G+1vcLyNl9aQvt2LFZIb8ZzmO608JgotT
wwMBnaT5VnOoALBE9sojnY0fc4cg2br5jcKM/VAxgat60e/1FJKJAHDTpX+yO21CCmWAAUTzNugj
BGlbyQo+4viYII2Gbdy6fxtgGh4a41z8pd6z313lBVhc3zrqACB+El8pyfcRW9n7okwPoMmPNbYu
nbVkuDUD0HNTHDIQM2vh/m5VNF5vEYlBqsl86xrwN+8pgrmQVajja3t5+2J2OCqJGG1LCfYVMtJI
qnEuolyliCrvY+/RQ4fzKTj5rDkhvznDoRb0eHmX/pzFLOkRX1NzAfgWGV/jx1Gfw0KTIO8C3OFW
WBgI87F2r9AVUaeXMoPAP0HsxI1OXGfOXC+L4loVg5vtco/jxOK54EJWer1VZ9rsIAakDPF+kOI8
tmUqMWI0EHI/OAzqA0jZG6Tgt4Sa6Q/Xooz3/T1APoOWOe0A2MxqoE8kMtFfai5zLg+ohYjXQGjg
xiumkuujuRkccb1izuJWpqS0sR2QwLIb0lI5Yg7IgXhnTt8hAfiY2UBO+AjqMcDDCZEwG2RDLOCg
fs3wqN87yzZ1bMtub4p/lsT8anPtUT5GemSYs88OAK762uKS3SvF5Zi+O4+eFjBHpr0S3CJTZsof
NKgpasqk2MxGbjNaXJHXYGEapvSACBTPEkyaURMgEVgb/k6oTMGU8yDVJ4AMRaUiQobnkE5YrV4G
PTr/CkUJ7JE2LajuE6YU5854Iptt72h0KJeJKVf4wsfkrLaj8dPgLSTOantpFZUUMCkvgB0Sv3am
YZIb3S0p8MB8fIwyOFrII2XltoJDBheiElUA/Hybful4gZ3UFRghnrDuZvXcmrOXLTO0mXYxatkZ
jER9ruztyy9+T7Zd5ntOFHMLdJMqiwmbqn4eSeQZtTmIty/QhogNshxmY9vLziyvD3UAa7GmXWaU
1KkA542raDdetHdB5Bb+BfHxsFdtfIEx9/b5WPrAE3TgAwIDVgTyC+v8hY/b1sDrj3OD0qLW+QR7
wAxviPq9ZwxN+1GYVNnRduaFvhe1AhE18MbcYYKCjF0DEkQPh3b+L2ANQLZ/Cb3yyG+jMwVx3slK
Tu0el16kzaYJNtAVSghMlaKl8IOeTGAqtRVJCAKs8xUjTIajFBQ83j69YXmFAJmyt91RzyOCcSSw
f+ZBXHy7UjcET/rO7/MPfntkaKlG5OVnk1WvKZOCH9A2+N7wihZ1JjVhapd1wYMaFvPSD0d4y3yn
wuu2VKOMRockyCb2Gob/bq6dEYD6A/V+OhGjDhquSOXswwVBdHVpRgbOIBZ+AY5lcix4HruAGQXO
KYmCV2ia2QhEXI9CZpLETytuJA8GsSFgudgQfsJG4Lkuo4xnminz13aKAKL7V7kWZUJp6b15z93B
41khA+TQBrnfbB7ancapOBLqbhvYDzP86qOwcVN2OOu54dblmrwZX4NiKRJpJJ/TMOE+D6CLyzAZ
IZ69TLuKij40N4J1bN8GtjAnjKR/uJdLBIkx3JVM5bjqA6N6NaHtwFQAFlE6vrB4L7fUHLcw1i0m
4sW+JQYzmgDumM/bEmdEPjfIW111TGleVW5tYzrKL89nBlKPjRJ6ehPnShpOY69WnNjsbGCWGgIX
zjKMZ9yLk/vtvVpro5ihFHYIulhpETpQk5kYcGcocmNoz9Egba0P43rcw6vmiAQNfCo81AXJpA/F
BZ6/UiAjROzwqKXblElQ7uQBcvww4531cnIUg+2yfD0mjzCSU4VyBhTBQhrMloOgnzopMsayUr8p
zvsybO1mspmO1uKxkuA01/CGR1yNSHgpl8IM6c9tpOmn3Os/IE6g8EUv9TQBymfVw7DqbvEL5DFH
iYX5JIY+OsmKe87v3TCqptBJXUYJLV2JfMjw/PspIlTrJJ5KLTFAMzFx90tse6EypJpFA6cxeYT/
YhVcQAJ57zQmO7Sc2Zgkw9ZPCBB4VH026Q5HW6G8dTLoLAyL/6y1CRQ5dRPLy6KnO3CC+WZU6qbp
PLWbOgfBYGzNWTbt839RwBm7BxYMqibkmO46jKpvZQyPB6UHsIuCbJWGsx50yfF0QeuHAejcPalo
68xY8iOSKjbmI9lPBS2oETFniKDlF04N9q6u1PNWL2kuc/IM5GI5nM4QWoRPnuq2TEFNt/aN56qX
XOtjfHsu0AtX53VWF18g199saN1LLOoBk5QIc3m81cPaIztQz8QosbPVZiiEGwRo+y2IynRWVWiF
Rk6fLp/jts7QZl/rHt5aXrQjg5peQMSZVpn15bkgVqNl4PgDP2r4XjOc4uK+k68excd/kwZ6oLNO
bC7iT9yJ9NwOpptrjhxSQJW5YoqX8m9sameLTbLlOmAdUaWd2ySsR2KvG3iutcXW0tI8YmFgxq4z
t1nqw2/bnSZt8Ox+/p1HTTk6wI1Ds1w4EidqnUoT0fA9qDJFSQFSwnHY6htgtQm/yYf1bCdLdlHL
NgBndUDVCYfHZW/3t/d/eWPwOvVhHE3XASanvtEfR5lkuRQoLHmMSqrTA/eAAoow3/q7HqjH2Csm
6v7VsBPn2sonrS9NEdjZGkYdeUKryovgCrCy3MN9YdfKdJtjfWQMh7P8JOCQg19Tvtmr6J9awVDp
aDhRoUZPQowNPF6Fig+0f/352P45DKGXx0sl++NU1HRA+Ve28YkNzB31gSUNnpx7eGWHH/pA97x4
/APd4kkcyjsoqhKPy88fRqLaw/i8C5e42ghrNKEjBKn51WJzT8UwsV1mDKbJ1MgL2oj8eIxgsd4H
U5W82jJIlzUnJSRfotvPhPUi3WwnLnjroRf0ssScyorzJLpIn7mkDxpuVVdxnGa7S+fO1zD7oAnO
TKBFJngGUhzDNs/3abuZWwmysikd2RZhf91WX4tITsQQWiDfsK+UGJzq7xEfe67SLCnQ1zQieoD5
ITGHhCr5jqVmRSy/vyglmyQqFMAX2fqRWv/oVLbEjTXDWHtq4Zl3xn1vlCZnZZbyR841DR5HP7Oq
KwLzv22A+BYuDpLBYJ2JxYNGV3cE5cUPwiMZBx2/enNS52MfSwB/IzdLkhmCusLJkqdalOipwIPp
Vm0c3AwPYReEjcvABePgMyRUkAr+pVfoAAgGC0YG1fjnANeo3gzzbutKv28TXiDcCNt5z55BYrLn
aG5LaPGGhaJdeNog1j0S5kwZ1NFfLSQ0ZLI9Sw/PnZ8T1M5rt7P1ttvGbZG5B7tV79s7drnxOxzh
FUGnnvTsmNACTBme/3loVbADy2v1EsTzfTWZuBgrka6yB+HD4wXJNdyy7HwDvjxp14DtCvrV2mMT
C7gPS7ntHQ6lfy2nyc7tGCegsaSARzhLR8eQKunoU0+N3KjTKXipWtmesvCRbdzfRRcQD+6a1FUJ
4SqMwsDLFWjtIF3ZMB+F6AfcTGCrfoNRqdS24g1llFGPUz+vFWDZEpIBSmzv+MWcfSdjUZisaqDm
5kRLn1vmeCqJZ+PuWVcHTP7JhqAM71RpAW9cXG7zxfsbaRqJRPo0ovH5i2vRj1645t2WBWoUzA9I
UrIANGi20HTyWg0NloKpnLCG2wkmRFzK07y7uFXgjkbGKYdBVX9+zGcDqXH3UNBk+WlDBN2yQLI6
udNmbyDopZZyX0wvPvRIVbNSd3AvzN1U3WR/r6HkHWOr25mDwa6hw95iiXX/uz4nPMv1aTFQZDZq
BfNtg48KTNz8x2b/UH9BmShK1aZbiHvlB3el7bzGTEdlxwzsD4YM53OSgSryAdKvvxiplBds3gBY
O6i05Qb87Dg+dhh8FlMHXAeZDd4RV7UHACjIEPY0/89mYO8H7u1GBuqF2TOtOAyyZCa21KRpslO0
9FlMz7FPrZiOAS1RzD7RLUlTNFuLDtrGFH77QShYi94qInwu+odkwYKu3l4iic/xHEiyBOT2hCNH
fMqr97AHabzNUR/MjMpv4m/+tn9SbXWb6nkyJsox5xnUQBEvrA0ZCldS9uor4jLyv0jxf9pZ4ySW
vZ9Z82KICmWVNmWRNkLz1+z3Krvo9DxqzIe/p8DhQRqvMKNODYVzbpg3OEVWaWxXlxSiZjWd9cfO
p/qQO3EmCijBxTFA9ejxumEEXbii0IkA4U5UKCiM4wPEHCTwxvZuvtDocaUaCIYAQkeKdd63PGcn
IC08fQFqU92eb+0bv+NYX23TsFiJvOP4QiBpTZGID50P+1oOQh8RgfCqLABOKhPChM+/jhaNSjNL
dZvb0Omzdr7d0oBS0POzU3tmOPhOj3UPoZsnpg+DL5R6dPPYO9K69dU18pitlXt/2RBn8D0TofIx
3me3l34sdsyhp/x2xklY7EloSHbdFQYY8Jxm+cnGrJYO4Zlzg4X3Iw/oB5hE4ebQbDGDm1tayOVn
3zz/FGw5/QFgs5CooKj/jpcDxYB0/hBbAVQCuO5Id6bQ5XiPnffKqsRInUUTiy56eMRJJBk5/vP3
6n6C2zDFPTW8JLcCg03c02I3zUc2e1FOZy6D4J9absKIXPuvDvI6ADJsVMKFr8RM3dqFs0Q4J/RE
MpwAECb8t/p+MmvQ6RPktGxBob8TjLTxzWtCHJz3fMyF8AwM9IGWsKtKq24O8PueOiSxIU5e+oTo
sGEAZfKAsYnwAbO8ncKN3+bBJfGRJyL+v5EYsgTfL+Ausy0Jy7j6qiC+74Ui4+MhDlsuxsS7+/dX
joiWWobJQ37iq2zETnb78gyx7J0p3YdhHaw/frsNR7pdI7qOrTG6OEFz03IlZtPZ2hwrLgYkbT6t
i/2jUB55Wa19xnK6QolFRHNIqHsAa4mDwMEknj7h/9UHW4B+ciPQq8Sve77PdB1+yBHCT2cCJFJO
RZlm6DWT/cw1AZIVWvwdqV2VuX4wQ6C2joHT1Jm2BI35PC5LD4gnVOEDSDzp81Zfr6huLWUG2SG/
KnCaPdxKKoqUzLe1rVDHFX/YJUHFC+/07dk3i6FmLTEFwseQMt41OLzkIrqefGuuBcWPv09tjMMl
CT4Uzj0y4TAcQT6GzvbZxxD2RkE/xMTyLOKcBoMc8n+SToQO36m41UjGXGS6Lpmp/9tMjgz/jz02
plm2qo1zHJFc376lscrf2v3Xweu5mUPbxEaeblXlFP1Vf3HFPkn0bQ1t4uHD8MZcHkw4Mup5NQyR
xDgddpwFB+E6p4mF8vH9A0KzjlkB87BRum9c3i+ess8EKWFTsQJErmBciOoETljprlVRF+qcRfrP
3yZyA3AdrbbIodpmnjqJACgAbM+jxgj2Y3fIUDFvEbLudJf+flrlAz5tDAh51aCpCmRfVAHDPLz3
Nt7dvLgzH65Cs/7upD39ESXAuk/UfrcHy9lDY+EW62AbSHYQthxQGxu8uBMvqFDkrhbTwMpgBNw4
DfN0zrO5AqnNxFVb2Y9LpajidqRizilYHAaDKAxwzF6aPXokeHCUrtlFCnR2sfKwLTi0R0VxYval
n1/NRqInPYGQx8/Ptcp0tWKpCC62BYKvmsSmGonoEbGiDc81isUw8H7AieIdpi3Y0IRyuunQnALO
uX2nOScdxx+lNZzPi4sGVaRY1+od3A9q0d/WeOudtqTx+6UoGFBmraPeWiaXaPlHCM7bBbPdczfR
4cHZ3IDO+d7FxWpClHdA+TTTa016YkQUdNpLDj/Ge9GaUXHDxQh6GVnad1lvqsx+a/64vkGO4xkA
H0lQ3XnKchYeC/8hIF5XJZuJ2wSkl4Tb832dBN6ei8VyHSC4AlsvWX7hf5MD69yRrkolHz6M+5fR
EHEgJFTPc92lptUh9hkBG+yqUNXy+h2PQKe8FlPMoD5SOohcEOjuY3FEZovvXflCUJl+l1SFGvyM
YsmO3Ybo00UIrz8UPM+mV0Zg+tO3ui7bgz4WQ7XAbNXLlQPsGqtDCVgfc+B6ehihYYQxRJuGAHmR
sr7Ki7YLF1VMvmdvBc3kMaFu1ukuC1aJtonau7ewZX4KNptQ8pMJTxD5M8WPqLqEmjmg//rJm1Dh
EEC7I4NBJNS0y66QH2FxVlFCySq+jWopYb6NK5vgwEW3vrAbtwDsDrbpYcTvDg+uLoG4y+mZCC/m
kZ7D9llEeYJ6u3YUnHviIuN1nIkkXxz9pto476bHmD449pyyMsE8ZtMgqwko8e89Xy3dlDJm33x/
iYV23D+RfyTTu6wdFSpvuhXPbWAt7oW7YH+bDfs59T+DkEl9erVC8AszYiQWDwm+7qeJ8GIg0gnX
kccFGOLi3toShMthApkIGSQfGOliSFxp92PinMjXo8mBB92EHsY1CvISK8b+oeqpMYFsk8T0TXPW
0hQh5usRE09of2771nVe4NRodJs/7KnnmTQE3jsEnKvCxhP6jrlTyeytZhv0r49g2BkalpM1P47R
Mto5mQKEwIF40MImF9+r+QeZ+KS+bFj/JgVqtjEERSh+fD0lgUQe3BVtAtmS9XiMAh5Bx4XcywUh
dmfkWRQgPvUG12SZhTYO+SsW2G40Qqzc1+XCz534W+Av4HHqVTN6v41FJxqeCJ02AHmM1ajuihpp
Eoz6qIAVnuSNZ+X1iXLWJTDnKXczJrRQkJqAbq6ib59qQy5bVIyelO4/WQGHMgIaUpXfmSDlGpVa
0vV7AflPoGNK6A7NU9Fkt4ACSuM4ByhC3KYt0q0zxk5m/vD2huTMdOWiFU3I7feATDjlMp+cSGuz
Wziuk5X2Faze4CbN9penUh5awCPnq7OmJQb0gmzAOpVZ+VHkVaYFFBA7JWevjT7yq8JMtF27eFwY
/CIkANIwamn7mEgJ8Ed4wHftfJAIE5H02uNuba73qsOchHaNPqo2sQluc3jm4sicsywIejh8Y4Wm
hM9hk0tIcez44fmxIb34ZG041Lju1n5AD92dP49ZZoOboIJ/65UckK3x9s/uQuOVlwjHNjKGXiAr
W4zzootWN7rK8w018RuXyifucuSEMRdvtqgd8s7BOKEc+GRmv/xLnWU77h00meVEl7xIpV7wwU3C
Gd0odkA145LBKi4AuRYoXYRMVQXyqcuSN/iTiianCxcyoy0U8FYLHEEeeCVxIwRYsQhtc9oY9w7r
hse1hEoVv/9fPzaFGXg3EFQ94IhB1phfa7iwJrSrm0weA9wNeTVdUC9FbAW48/0UgKf9XnW7UcfN
JN9E6M3xHV5YXLonE8RXTg1mC/EpsX7M1KmiXPHj6T1AEIsj/jyfzz0bJp9nCx3grtNqJ3wvKNPY
/8atquhwI+3rGsJdvZZLXWHqCR0maR8nTvJr2WIHGJq1rvpHDNgU9v0IdRqAKBF0NTTw38RDHT4E
RK55EcSBmlWcOVnaS/7Yr+sHiPt7wGCDChlIZpDBQnB2B1Zx1BEg1mS53zut7/uclUg5VUIJVi7n
BBm++WFov2Fqx81wLBvgYk2r8KdOTKrRnAGLL208EHDuOTZqESiBfhIFpGZU0jQWkTATbRSFJ3vh
IknggTljmxZjW3klcKyhBZcPDqv+s9Mui3KPybqUj1itJXoZKk57Ty+aJgYn/5hg6ndphbbCX5tE
wOVFE+T07gTh/jfVGTqak3MRCy6FTZvGb6g5B2SvyAwk9se0qeWgay46wTdXpyRwUP/oeFp/srXW
Fnm6cVG5jErcWET6QKzt4gP1PMN38BwQOC/1fvL+8UtNXKIBqL9d6lndL4q9z/ii+8pUIbmHy1sL
F8sniwHWGIeFQ5lK86JaCVhTCWjDknGXEaCdaMxLJ/IphYQF2e02JipHWeeTqHHZ0PeVelOOj89l
pNVimkatuIOJQX50lEHia85DFFq08Bu4w82hScKxaUa5ODmDnYi+fusqffHF3onFKzpbRbA5sdc5
hfhTrR9395LABSUi12iQx/WWj3tR7zyP5qA1leuiwl8EPY0dMP7iU3X4DsCWACq353cdLvXEG/W1
a2zSnCQlvPv/Idz87szjxKMtN15pswXgs/kr6rZNmXMHDOp0uePJ+a1tLGtIy2q0hBQJ4JixYguT
87q80gySqZyRj4Oi4WTPJQmtiVtZrcqNwn0/emqJA3W5ijtqI16xh3rZTnYowhm7qXP9rXcAW6Fb
4Yd80ZD7Adm1nJzMEUR9Ij3aV/yR/09Xza1s3k6U6S+4xRtL2nFr7Cs8zJ1U/6PLNwq4VJsp5pBc
kUXPSENRfrbTR4YUrjy+9bQiXzENLoNgO/5JArBMbJ/qLdydE1H0QdSjB0yj/RhlqUiECXbhMF4x
46YQ0ZgWG3ru8TLnV2VqoeyrdkuvYE2TpWvtjU5Pjg5mPHHrTLBetFGuPE1wlDgz4iSQaBuZ6Zie
i/zSMpbRcSjG95Dgzdi0qCzGtkBYAjGiHRW0cAInq9JHmHk5tvyYEUL230WVSBIdJV++JRXvdbkI
ZPhuHqTLkpl80hZnFSl5ZMw1x8x6qVkzYoWj0WNBq8DwhSa/GhBPqBY7Sy7ptt+KWR85uHvV5uXE
So9rn6JXAqu1Cg1pyNWwIxymIqvCghPCmxllgqxu2OlB5as5LW61gMnGujwU/NnSq6tSQdPCo8KQ
4j5mY/01/diTKef8I6tRFP/s2wIeWXysqpujAb1gLvBBWZgJ6+SpBgE4xhx+wyGTySTvO0YyxtEZ
TIFmV3rB+FW1ET0zpSUjBd83P6e9lwEgPe59r+8o8o8Hn8sZgtcX6WmKy+ls+oICBYqeXfV63fD1
kDEzQ0UI9fzkRniHDA9EaUWaep0nynVddjlTFnJmYpFH/2P7dwe5o7F2HCNhB3PBMfOW3g+YfFHe
8bZToBBaOZrqZhhZtZixkNPtZGUELJx9S4ghSVPtQwE1HukolT83oX2BMkJ6Vqre4xmn8NZRLNQM
XvkwjCi7ufKW77XHrPqiwnie25h0O28aVnF7nkOCf7dgNINKpH2yanelFWQppCzPQRyKSrLutwS3
72QfItstc8xOLiYWDsEsJAwOj5F2KKPTqIEN2N2fLMSXTUnLwFrjQOteAIN7aDYUu7scchyZHSD3
AERpeSx8T2HY60tcPd+fr2Y5co4rkTlmet8Zm4uEyQxzWMbfhnh37k8jJZwkd5cqKlyavbtb8s14
oR/WndkPA2SQ5avqzLIfgBIj2Wchu45v+GxoFuB5I4yHmcT7wPB8bcg8N0rZO//SoshoYlGrLJpb
oKFIzPA6Q1LenF4TguOxhamte3U3hcxUtJSU3vodL/NhIor6i0SGsAV7lA7qoD5FGJ6ZNDNc90Q5
qgRPJwvqcpj2v5wjFf+tasIn6dR2Z2+MFz9/s2DU1f8tv27tm6r51IK9CWE7tBb4LADQVLqUvvxp
JaQQs/ONgcV7S0XKh2//5CVf6XF260mkmT7SPIxq9M5EHOD/8MW+++NIUIEahz+k8mYUYWOnZaQi
F5lqrElVOzOlG3Rxkry2pYWZMilVWqKIO8WCZ+ypwxhYTrVNkGNaka5quTpJjelBRcwVbUHS4sra
1EoNqQEJ1iu8WE7OK0NEMkX4QrubzOroBTCIr0t/OMbU9aQphCJMQwecEi7Dq9MjEO5JyQTIU1Va
mK6Dy4O+Ws36P6apxNwxZzBigEa1YyMQ9Ssxa28XLB+WtXBgdMSLuZQvzmDtVxjzhff/blaf39Uz
NfVZZm/oNFoKXXRaApU3OyBfPZ+G8IeYp/n4sExkCpveHn+EPGjkwLJLg/txK5OGVJ8TCqN9/axZ
KQHUfRtiHEpyaBxrUiNoaRm7p9n+jyQ9v7DpnyKDWJFyRPAww2OgUFeOnJIe4U6oVACgVrLTEFs4
G0eZL4bLJRx8fAP8l31xzHALnnQltGa6GxaTVHdPSsUO3m0QPwAu7hL7u1PbNnauC4b0KnXjlHYs
JVkvZSy8+mCoYw3wWTM7ONjwkSFMWMB3VZjun9vGPx6VuxI/3nbAifHsMcbb2CcOu6OoKME8JjNP
pUew6a5/IiQeZ6bMWyjy1n/XBIor60FAO1pIEzS0v2Z8Aq12vzkFBHihycqB0pJOYrA/4qhGx8ux
c5Ox+1c36iE56Z72+Tp3Ag4ittgm+ubSiZ0z04pwo4IQ5QEZmhXW47mQersuo59PJwPsMulCPLz5
VDW6xGBEp2X7BLVgES1FxyAY/lbrtlvKMHR6wVWsx+LuNt4avFhVRbzCnEwqxFfDtwB7xaFo55bM
rd5tjO8Nq6Ju3HlxmZFRd8QjThiMJb0+1YykBUdSiKjIrvjBtmzgVNL8YzEhCnUI6ioi1MfZXnW+
vRqTK3JxkK+HlMFuAXZ9wig+MH+jML8EC8A0fLLQu93I0eBtzM5qXeILBC3pdd3XxstbFX6vmXGL
RuhevnbnIHRDFaKwD219pDJfOwgSZo/x2QBl+8G4pmMpzi+OYjE8SLjBpiXko5vxfPTTCGispD6L
8HKRTdFVnv4l/LypLkIL7V6mh+1OgypDxNnNU+TpXy2XWR+KG0/G26DHXZh2F8fSYrUqCUPHXlg/
qvSU09hAWb8YWIUuEocdKcTNwJm4tWeuFn9kSVwiJ1sE8d5t+oQuvWJujrOO51ywtX+PDp3bKA6D
HJ6Ihyy+HufhNHHFVoiEIos8HROefV4tWUeieg9fgYprtgCqBnYnTZKD8aDV2gcVXPNPx2M/y7dI
eKnUQ6JfK52I0SwsrCIKbhhHs+zfwKMbDypB1f04j0Q9HQWBzsVZD0TbeqpPzhIvbpOrnPjq/von
rxdvgcju2IqQ9Y0zh3XGKUw21ci6K9vhkBgLGmf6IGmRzrcDBAD2rgU986NLmDIjc59HULKvjC/R
zksoW+mxwOREGG1lV4A2Yj3u9GJ9rooVvAIDQ1Mortj00YfFR2CFGJ8KQAqNCXAPc9j1kK7xG1Gl
1nI2yJ/Pepu3bxXGr8WjZ20wrEfAwQOe2HY9QLV+Yzgs0SMoerT8QPdEyY6c0aE3FfsF80Fh79xk
zdgy79cR9rwAkBxeNMkE4HoU26eHZ7JlKOjwW0Klh9lMu7G+2IqlbhE0lBQm5ycW41dDKsbbnazF
ciaqXJRMR7PrIBMKSFDRjQ99JRPQzXfzhIUBo2dSFIK7Zali8xXpmDXwmC3wDo1sdoZU+7Dsurpq
M59LXMf4PCQHaWHgbPnIovg7b9y5wTB8YLvxO9hBNb3sii78tvfWmVDcPyt+N6Xmm0ugnh4+uZFJ
5yYKR1wbp9oKjKIxMA3xEWpEVQnr/coTDwmWRvEf1aWyHfXHOJnFa/i2E4jaQCsL5ooO0Zqzs3bN
bVPHSJ4Cj4lOCo7GxjIc38sNN4OePpnFcaGanwkd5vo12wMGSYYXQmqJqvxEHb17Yl5SDH/wtA/T
+yIqOH9gtpBT+j14BhLIOjZDNFHKtZP3MyUxrbN6HWxMtBGaMMmVx+9livXooHWJW6C5706DEsZ5
cc8CwUPC0Ye2ZSmuB7oy5rXDLesx5VFEpchYVQhDgX1SWpoQIHydOZq/CDS3Ij5NNgCjF2CG3bmi
4rIiimbWFMAezYvTv8F4xSq4PWo13Zta4sx/zx563oOwgUaU59mOLxPr7N10HcKyC4QIzO/KrwG5
Ub1k3hJfoFh3Cysh1JdbyMkWCFMhu8zjdkjg8KcDxQA6ON5SKzFFb0z+GJ2af/KDPm9GW56FYOaB
5D7DgeWOl448Pm8Ft0gBNGkgHSzQCQtPmDciBt8SbJyhdGBQPtFDtq0WdgvmIv3zNxu71jlDuwyG
c72VfYkuWTK+yHIx5xeitauwdqTEmM6xklUbG46kVYdXLsKrdu8XYCq9DRu95SkS9k5FDNE3afmO
O8c0aCKK+VVOXB4Zdlr92bNR6NXhQmL6OqCC96xN5li25vnJnf8fDgOvIG4rtvNpchI9M6ujLQnS
XaEHl4iE2hgfer91cT6WvFDRzFAptDWWaiBDnUpt3gq4pc11z1NCtZK/6fCHqqBwPc84/WLd+VIk
zqCTNClYVAV8ZdOp5qjnwQW6WLjOixcS9du5w+3HcNJeDNINnyGIWF2DY6AGg0mgK62eKXT574tA
qTxBe/tYVGP7t/2VuXoAjmli3uCP2fiNrWjWMxtRWiND3qppChP2HSF3lD65sRiWcqYOEMIJAkBz
Wb7Yrq+10XygUDo3cIJE/+z7MwyIU+otK6zQ3OTLy7si5qdDfFYBPICxQI8v8I1EYAARvgOaH603
IrhJ0TnU6DTth2/OS77r60qxNtr1EQQHcoOebi5Df/Jb8a7Ch3QcFWpn9WJFOhe5byk4ZDz1R44+
IjfvUuF39L28gVrZB0lJdUYbdOvdj6UsUbCLir+15ZkI4JDvBnIk61xsz7oBToeDwHT4scieMm2t
Q8JXvSgvDPcc6k9zwGDAi00so/GCDSBF2POtzUofo/fY7xkbq+/atcPBkWcy2DZIpk7v9Hx2TrJz
Np8G/sZQZ06HTL/QLF+UouVPvKOdYt1xS3r64DInbGN7MzQV5+VvxU2jtbSR/TsnsqhjCPmgDhTg
4AiqsT0QorsjBv5XMYFxT78EXqX/bvmh8Em0sZ448RnyOfkwTaP9zzHfLUFQACNjsoNIs7PthpVu
R7dcN972l32hBY7JiPUzAwg4z7VDe+QwqnmArMHxwSjdAI7yS5AECQPP8uzHs2gmyn34zDfbQ6/1
SvFQxYRzMUJmItSH1ETh5CkiQd16YfntM6CAO99DsbEehbCI68iwCK6wsMdJmi1+kG3FaEjifPS3
a0LOcOC59sq69Tcvd6a7YsjeZ9xtLxcjK0dS9GiIAQ9Nn7x0vMN4W1xlKIgzt1yKcDEJhKCts0Ku
4ocEgxIlHCuCtm+/E4PYkxjGf6H8SycHrV9nOKvOFqJly82IcAlWXnZz0EZGtzyGKB29M3R40PTC
5oDU/23ab/RpoLXoU8nkqT5Wtkk3yg4cK8V21UA2FI6yh951D1pUQ5xIbk8PlsiudrLqttiI4a4n
bxlnvm3Cas7cJa07NrOhzglsE6yLjWZw4jbTXH2URw0HTcz0Ab+BEX8AsLj9XaApEZvPeJ92JcS3
Ea/9Xcb6GTxRzODwbWmjpMRavV8/U16oASW9X37+jMGGkwcxbWry8vDI/YXHHZx/M8NPUKHsulUC
1M7DowdkdFhi22Dv1654AM70UNDZLZijjOt8ivlc2IA24ODcRdNje+e7wdJqsIyDNzqs0t1HaC61
dxJEN1CrtdNCOGoZiEDMGiPmI1dnCRVHJn3p6USDYIplDTalOZPSAwHogMn0sA9eViwth5xcU3PI
zNsuMIydoXKoP3aNs4LYg3jRU83wSSFe6NUc8cem1DqhNFVtKtGvzE2VKovxdDaZBlegC5xa3pe6
RBRw0H8oLbRF9M2TLq9MeAIcbPPjdyrSaYSp8fO0FH5qAhFEeHQ6wxRvkkPUntwiZQIt9FMqFqxD
UK9dmX9+4gCYuA2YQvVfgtGXcQPDrhDqsbgMOvowfhFWW2RICgQDM7YDcqN+A8Xrb6JV+iQMUf1E
T1lfsjfF9HTdcHNBbkEYTEuKLL7njJMA9zN2171muHPTC20Zp0SQdf3/EOWWuGKlTCtx3j2jraDK
p9FJiohhvkdBUwK1tlQeZPnWuDUskZa/O+oWYUj70MZ6P60dFwbW9/vBLRzVM3ZY07VhnT1l4G9g
Uc4gGE2uW2Y3JLQNjyTyBcNtGZSucP4plQ1JW06mXRVpGyvi3+bDIbueIPbmLKXtfV4Y7g+qGsLs
ogmicGHNGmKK3dm34wtH1L2y/g1qtfY9ICRLis81Bakq9qNyOYbdxVTtEO0oW8tVEBEAxKfsTjNO
KNmy8yl+A1tfwxwAOLwq1+hvRNhrGF+mNyg1Fzv/3CJragiHegSfoyzV9iMA84EzR8EyDzKubIoy
Zbzz5udd4eJBs0mdDiY3dn2UOVrT2vudB8k5i4ds0+1o+GmLvPRTA3RX8lRk3oFq5dS8JecVGA+g
DbDylEIO6HO8CkhcirwPFTvCHxG8Ij7Vs9rr6jRjGUJEV5U9DFLVLz/ylMBVzQKul06xd3zctF89
enzDxb6CCpPfohs/X0b6fOlAg1HOoh1m/k2jWly0XXL5Y9tA96nJrlb6eHF+YHLbLh/U/8wiJ1ET
P72Fj8OPaQ8/mkl1XcOltnKXsbSsG9rQwSdN+bQ+Wq84E1dtsonGuoQmsknoQ4f0M/oG5r9XI7go
Rsu4Tqod/ioeQQ3gmcKiRi1aERRCVL38qm3TvH6UpHFioF4CMnLGhy+pTqJA6rjBmKfR+vszFsTq
CzvepX+utxXhkeyW/LTQO1Fp6EJjXkeFSXFGlrX6PfoQoI2KmbMGD/x0k4BzRjuxjf8ZUBq93+gu
7RE7C/Z2bR3Pb+1JUj+idrWQfuf7L4xyAY4DVeDKYhaM+BtJLLSN+lbihWC7VtR1pT07JbGyTmH+
2BlTKCmoucd5BaPfPhyPiod8LH35IEdXAukSNydKF5Hm1GxRQ/Ev7JRGkODT9Rs5htkv89q61wCT
IiKxqZrL789FFnc8ri0//ymTZ+2OTvLQJKxGfEAerDe3oSO5LWrt7ho3nY028mQtHOnQ9ltFpDRN
ZvrKKrPG+Gu6AiJFrN8eqspB4kMOA1YiAr9NPKPq/k4wGkgXWVpRJZJXyvhruGTKQlSLHAgAf9Bc
7QucEbTWng3jO+Gm1w1BKZf+bPwC99GPpYH8KJ6N3vDo0FzQsN6RTVoWkngpQb1OuRdpoaR3Z1d9
CnVu8ik6tKqpzibT5owjmDBptGVlRd4vXLoo8G9KGfBtEpFnRIm2Xkmr86gPV9fL7QRKMQbNM1+x
2UeM7zEmDGMibPy5dd1VUpCCe0KYsN/Txh/3V/fQkUcPqlrhdE3/dzOLIo5USvYPeQ6fARVcbq3N
skczpSO0FMG8Vb9cna6TrewlvCH2ZskJ9g5MJcCuYLvXWG5fhvyCfYSHoT17DnYR2auDT4mNEuhw
T4iPUPFsuIbysiPfPIZSfIpq/4MUu5eIwY7WDQda5bOlHl4YEDe1QpFpNylH/0uJF5dksEvJiGZ2
bwrt9ZTavFE2hx6CiAYrMW62+cDHvWLYXCQeGQCuQJA31aIaWDpgFcmrKwD4T3jRqLRFMNdpur2X
NzgQvq+DTopaT76WFHDMykih5PzgmLQE/32DiQ62mM+/XXsfwQy0NP7YwVBRggB60m3h3a9Qnr1Y
kmdGdp8aqoO+mZiDMaxWxIETn0P2eMNPbBULwKtchsyr/z1o/+IPtukeh9jGco8YccITouoTNY9N
szUduyt8v88T52CzOH+VHDVqTV8X0jhBVPVBPPygPwYaiEWDF7uwHFFqu4jlXvQ0K8wrdt4e3wMX
tpYqi8nlkOf52akQ++WemsPHG6YDjPdCSAc96WDocnelYtU4aDz20yIyfeFf/LLd2k69FajlDz3n
OVcs4tvpcY37x/+JMJjgSeY4iIUukkoFdF+z14hOmUfSjHen2YyKw5lcvYSpWm9zSj1Vo/LDC8Uj
YUIHZevPU+26d+QpRNviAIveyJeyhvvfF9FSGm3wdK457a5zrG+OUZSOzGOzySluN38fMCGOc/Zx
4NDtimOSnrfjvxIoB8iK5wJurmnT6UGIsRGoXWLdN3xtLQdiIq6vI+XmGFOivvi2vpG5C3gsU8dO
B89Z2N+v4aQgAdqcY1pJSzwYwTQnqzlY3+MHhDYQQSi7RVfuXb3XPZ8BN6vnwrRfo1tzTBoz2IEi
a+0CR5CfczfsAEAfC6L/oLVxF/ZytUhdvYW2ooP3ek6TwB2RBCh2AJHBbsBHFtQRE6y3V2/zD6Ze
Q0kPqQ6IdiprR7P40yGkjatQx+lQjuwdtnWZx8F85MFM9VyrOILIr0UIL67o8Vcpx8xmkl1otCJw
U9cwOYLoE8dMKSpuAE8sQzCe1K1NnpwTytVo3EN3YR1ROEJ+YCwD9O5DWjNXsHZf+EJ2JZ96I1Sh
DQ68OjNvRfmF8qEqtDn7BQR79Af8cqpBDwBl/OVm/NvWqfNRh/EW2tPo/lGRz4QizEoyZw0J5yOq
IjlE7kF8pxezMWTJKb7ERurzgdSfqsZ7BS1hZf43PPramHfMewzxBqRXsxGpUBdecpV+AHaf0AsJ
QXnFRnyPhH7PK5mo038JW3ERODXCBvHE3a78lIPMguKPB0cp4+m1wGPXoZLL3dRXMwR5rPIMZ6RT
65/pIvRGvzbIQOMBiTqQ4mzxl2b33R6Uk/iy8HBhqPTIMbDjUyJvsu7elpUG3bzddGSUqeextP/c
yTY/Pzcr2ulaGfcQO1gNy5Wk9FQZHiEiPoi1ZwmBLAsjNHpvb5eLMh+YGenHEk18dnLZvkCZ1+vV
jqwnXP6MdYU171YWhsLYQrUZfLGYBREbra2lf4SdH7AWyUyjpFMHHtU+QA05FEiKjHRTH5c/liFc
4QdO8dQnttMOBu7EVIivklCujeyO5yKRwzuF+/4bAVdTDLRyRnZtfURsUadrSIbEJIsCzaIzKY+f
heH8por4yi15uMgugryRjyXSMnamKNDXJ5kn80W36OLPZQN+8E/43KFHrjMaBLSXm0jow7UdZRhB
PARinbKICmyhfQGcPsg0t09w10grK2RyAJ28BcAteUY/y3TUIs7g3n+bAsIYpojGOFavfj4OkMU7
EXCPmlCwS7hc/GjrUs31ij3+tNuIP93ZANsMePBsn5H8+frxzDAs5l898SCPsZVAq1no7HBTjRYs
1zQMqvbSuTbdgF9n1fGp7LtRThaHN6A3ZXtxtS5O90xxh5f+aDwbWG0sDdZNBVhMv0Egj2B1rCW3
nc1dDi+UIzy2OOJrrf6RiNv0jh1myCKaxFIUcmZjznuYBS42UG/J7STLN8KGO48w8ra6bXAjzW9i
aoe400Lrrl0ptOzS81w/OqIMXTO3ezGzL5I0SccWZS0lk+dCqHx9lNqOezNYfUwVhGa2uhxn/X4u
nq12Qu4Gq2pgySyjo7bVfigiRfEt+leUf5tJEETnayap0U0daIo4sJfL/loKX4ofpzDb3qRS2SWE
onDNDglzms/RMEz1+JUfaAhL63b2rE8SSqjjuI/QpNTTG3aKbLsqvDCRF6e10Zko2SWHYBKpq+o0
xetP5HXPvkFQmYrInKFHtDVFyLL/JvOyLZoGkgVffsUP4JBbOKUGsoPJvJaGBOfpddJ5ns9VEwhU
IGR9m+r27maYsHZ0DlPOy4RYJMnscV1/ldmoUNqJigMBGPZ05fLDxd77MO5BDQRhvWVB7ZXLYIGg
1O6RhstSOJDHRnrBeX7Eg8DR477ybM5esoC5KNmwjIXnC9U8DUyNKsFbux9wQUy87Vu3GSxAwHqh
ISDG/Lge7mqGRcxgSJpN9rgSWiB2sjVAez9DfFEHH3jOZYaIrXJAFcHoJoqvSDnlJZ0D0uKbF04C
jNNZUmflNvHPlfPSg0s0KGgCiU07p8zgpyBgGVUssiWdilBjFTu68nPUkaMZ7r3+gD2vnidD0nb3
ry5eio/lXUPlS/gKZPm7JBtp6BB01a5vevvvRjLn6uPGk9EyyQ0qr83A57LMpM01wr4ZJ4FrfKQ0
q5gdnW/piPQqqP6eiSfYurT3oNub+6UtmpsdriXCwMel6TSSfftWXaXvvelz4qynDNyHedOGB24T
YP6uNsKEy1RXG1YgxZPApgRr8oFqbloUQj73Igm+JfsCGiB6bQuhbDuvymKYk6Y2IMUgqelGDM53
aiz05Wn+A7FZrqdklmrYFDKGocHd3UtFYY+/WOORHNVZ7T+3Vw1zJ/yD+LEKejhvm1m1+t7nirg1
+iyatPGyKj/ISGQiF3m6F36Ww5Iv4+65QOnKHYYfJRrh24TKjG42C7468qOMPV6xb3Ce0zTf3e5m
t4dvXQZ3cMNGvEuLR9gU7oa01W2aCNQKSCp1Fe533JyP3Cl1moOftz+7gZa6wTZEJ6PFZJi+retG
q+nePGdQlZhB/eo85/gnqv9UQca+2UMTjI86TFyeyO7fH7rlf74Eat4dvyJUtAHnEA/EvSxcOCVg
gfgk0b+D0CnmkhhPWT1rWPj20eIzOzsCeTfQnTGDDUOvK/xLMH1QZznuBIDOU+N2a2QOf3lfJvcw
Ai4QzueRWqxK8llmfQsa3jAQECVgPHp1Tk+y7ctbu3hlx0z+LRYyiG3xOsgGJZrXuBahSu6HqtbQ
HgQWfCH0AgChEWgma9uRhMlCPzGxZXGo/Pg1QXH+OFjJt2/f/gTTiw/nkTr8iQi6sXoWtAivE4VJ
LRfooBH9j8W2ngdr9hVIbixpHEmR/+TjaCjqjiWQLi7TiOSZBfJxQD21dmkNG6ApRmhUkwj0dQYz
6BYTmONXzyNvGQjeIjc5nEb0SaXhxyI4SM1BR9Zz6iuUQRKEXKuKZzi+Epf0JPciuOZ91no6Y6o8
X19ONK172fZgIX9dxUiP7Ezf1mtXXV3Iy1TfaCaO7BbsCs9aPSVL3DTpLY/8H8B5bDim9nV16S3w
hseOJpypXmWB/8UX8UmY8raLXcggKGd/pVrePav3VBvkf45twx4dEbld6QEjJIGIhJrcFMho1HJB
QQ48jTyWPe60qytmVMOSWlAuYP8itUzVAZunGBOjI71J2/tZslpjrhAlO4ukjVp9ykQWiER2nYUP
Lr2I53d9USAq3jfSdQQezW4qo4ohPBSFMJJLMueKQPLo97J7t8zr0uqsCupLStkFrCCWm4b8OuQs
+J9ekovCeIVnUie6UveJ97pCZxaZ2BcCgQNuh9wFgoaLsXCz7Lwowtk2Yk8wI6PshGwnRXxx43Ux
2XolFhSqNR0fbmjUSBkwiyVJRJS6eMyfKpvXMIXBWuRtnEyMZ7Dn/dk8w/x43dlBk1WIngCfqrXe
pQkiJLuLYutUX2Yu975LuiHggEdpL93DFLxXNidnoraSbgntuvpgEToX2vuXNcG0TgztpE0m7I+F
igc6lARPWvGOOVeSxWZUwjd49EB8Vf1MYs+JiQJB3UbiGnlcUwTo6dmJ5OjgeWUQIvIMTX749MGO
On+QII3rM7ISdplFdUt/8XxdyCmYz7eR3h0pqPfjwf/tPO7z8xhQtGys4FKO7abFqZ8bZSu53WRK
UfjvV9gSew6AYsnP68drohVvEi+ejk0tQ1JGWfsaoZBcLnX3coTMihRG39hvvS0pSfmqmP9ZIdl8
hQnEHBvBJqRxuvs7cbiyF91cQPBElmvFzcY6zS4n2CSb/aQiE3IzFhU/Ee23z4SMS3aKmYw1lGM/
nCGqNJnwubg9vMrGlq4o5MmBcvQXayqEBnG6VEjESVAXSgBUCSWNFRZR5QaJ3O+fGJB48V6zVp6e
c0m5wFnhG4vK13/Vk1rp6H4PTvnzypyw3TzWJv5GZHBCJE/iQYhaW3137kLaE7sykdoRRIfMtz9N
4KW7q3R28JpKn64Mqp1vBgSf9Kgq2DcvFm4J44IbxldVbhYvjn+RtHPMm7i5jsajM661jEY2D3i0
XLLQQsqYvT2QDTaqfNFo/xMDXvMM8t8EaLlBmdsLKhvPhxPuWih7ZV5DwYYyu290ybifs8Avgary
KeXK4Uihp7lJUKdvTbY5x5WJPMxXyRh5sCIatmxt73AxlWrFW76nPpSn6wwmLOKY2o61IbOKyS1M
s1W/juqHZsDKcYOPDNBnB10PXSA+UCiAHUYKPDBwfmAGRw8OwIkliMUyzUou4+O3nKArnphR65yN
HjhvJ6C/R+ROCA5ovdHsyrYMiSInc1NrZSm9R9PKWbbWuGkFI6ZRfOEai7lJMkGNQJt4KZ52Jhbp
RscXp7RWpLKaltzdT/j/TCT4OuyUiHhuzIEyQMTP2qsvqywsctJJsH0DzDm4x/bdYVjfEzBAOe/r
7AGXOiSPMbNfRkqZ4PDE0293UvWip7lKWTz8vYSW0ImBb558kkBVzb72uVb6r2E7GEud8nuKt6L8
oDTRHgJojYSULh9YtamsZBYeN6MLiBIpW/hWV0USaMnPHqnWrM7/azBvUIov4X4VAI58QAkrySnx
T5yTMaYvfnPUyTofcpUYbTAIyr9WJ9C/BvC7QF1a+yAYobbtnXgJTFTBEZiLx4d8eh4fchIYU9do
If5vSlG26WLasanHV6s3zhMGzITaIcl//nMk8F68wdpRyYo+m39xcLyHjmK4D+E0GblmTkZkV8AK
8vvcShDotZBFlbZU52GNhGO4AwobLxBIWC3hltxweLN5Rdk6jk34IjZyeu2M0jJlBrT1FGy8mr5u
x61q5UVsl3+88RIvWSpeoxdmJ01yB0eIY45kDrmqJtMIQXLBKkEhyJmlXAPgMwX3waHJ3Uc2b/XQ
aMotuOTzTpzuA+OizSe9MCGlXRoIHkdkzmCB0ooNsoxIuTIIoIQzeGz5OxglbbJAKO4JufhaMzsV
AMihNOPHs+grObiFQu2i+LrDlcYcaaVI8D93E2d27xW+O/zsfkIQ0+HmrnwQBf9EJaxk8Fwr/GKL
32EkrfmFYE2cKcleK2kqaS5fJY7Mc614XOTRWG3wOz/Hi/vpOFxUlK8wPCbT3WZqe0gwfFOM7li7
2rNyJvmxkEDUwVpkdFROHb1yHbQPKWaqCdtXeTGRYE1nQG3/BqRLOvdzEhtznggyL14DsQmI/TiC
P6VJ2PKnCseQkkmUOwXZ2yDExIz8n1QCmHT4DUNxVlpV0jZYsQ6EQM9k/2GTab+Syi0qhZoWSvHS
PdwF/QZWvYmc2YLQyuCoj72IX0EOsgG6lPAAoAUvW4b77Sca20ujDQrlKHhpIyPuRXTzUg9ZkDXl
ic78cXnsHW7H0PPyAshHpIjQeNnghGD53w6BEh7ccJbdn1N0d6vbMdHTh1OlI2T/ay1GyL0vpqbn
QWFa+IKCWzIPnbUyCdc2rnBUX6VXX5rMFGZ/SRbVmCMYiYGifTZdDwo8N01GhSBCqZ9dvyW0ybTH
6kjw4o5BoXs2pYi3SCroB1+m2nGIc0VXcKBouBMRz2Rkl5+N9shVwHcXTQgsTy7cPLlzrh9DOYfW
ziQH1zxdyM2aq9inAVUaFx5Xmkpq7U76WdRYS5Hj+uVlZZLIQY5a0eFJdPhVKewg+Vdpt6f6v0Pm
ON2fNKCi32j1CDFHLSqthXowsW7fgR6ZKe+WOmZnH3/KByT5r2tRCFlZGJLIQHODzzxTTkQ1xfsd
Juska+LlsQ6jtKNJQcfO9GL0uKJ6bIPU3kyvY+8PXYOvNHMzeoQXIE/YTozQY4tbueXPLImQ9JDO
KbGmjGE1g9LK57vFzRnMiqGwidYSZRMTYXYcBYafSDOiKh62xB71ZxdP/XiEwwhnyvURhstozb+w
AOMAhj+V/3+wCqho+2CTaVgkVPl8x2l0fUx1g0/8sUugF8g/Hp+u6GAMn3y0nUUIvGm7TeSTN7sc
T1yMzFIPESwou3mVrj1788kN3LySgqtIc+Do4Z3AVYFchLsKIwKJ11qTaAvk79mfrIWBHwe8lGkA
0vlRTZb/VfqWIee/uMq+JX5RG/kQi5/GfX/6JPfJH/iamC69leMW0A9aW6jKsTHaxczniPH7O+x6
J3AdrC5m/W4n2x8vE0/7+9hgRnvFhXm73g3OwGx8JMt4yh8325qsPMPM2npJaloAXzsa26UkCyud
7QWyNc0M54sBcf08eo3pwYtAInoaUM0Ucg4zea2C+WLvldNLpJoPD7VmQ/1BwJWp9VUiHsPduP8B
LGK+PHBeZeK6h+r/Fq1kzWA0DcN8OGfAKSLk65BYqjfJGVMsCe9hls/1C9Sa+e+GPyuIDhbgTg8/
VUSYfC07QrTgA5POMjQw88UGRKtM9I4wEjZ9mCcScVcwEkhmqPmtwxYY4Bz8HkX442XTIw8m7zlY
Q6iEoWusq8CqUIpz+K/ynrHGFB98NCA7Z4xZ/R//pagH8F5vh7FtLfVOTu7yDrvCbfYcFGUB9MLE
pnCdnyJXm35JZWxqqNmbVq5dZtqVIGByQA2kwv6pCpxulhqDYBsTH7pmcEdVXs/beInguP/wmHOD
N5DH6qyX7m+jPLTQAk1JhJ00FjFzAD0+lblJi805bRMt/u9U8ISUEhQdQ3KaKsCOCTOstFDD2sRa
Z2+p6WFtYFtgANcz4+JQwAb7LuT2bUwUYKGzf9loMXUfCgQ7lAYy4zuxSkUBmYD5uyXywWWExtsE
G44X1zarHvNOjjz7dZXBLSn7xIcakdXshk9bmNPykioYs/Wir10cvpQ5NFIxAzzt5nVLXq6P6Zw5
fY34UhUgMCqn2+g6wI++jb/bjvqmi9KTFTl+Vxh0McdJoSU5Zd/Y6oepW8VK8EqOiWuHVkt17Dvj
/tLkIxMRGECOjGYv8e7a4XXlZlei3OJ8MKfljDHrjsWFIvFw/98+1N0WoSdxPtsmvn5QlIpepcml
sN6lNkqEhObdHtA5DAibLwBzkICjHbGLJfZsqEEVdKDFzscEgYVbZFtYvj0Yqx739fj4eV4VxBbb
63R8txNPY0fKd/CYozFPBGNZYpHgGJmuxTJyt1kZNiIWM81zTO/y6FgpsB7HqN6WQynlryCxwbCz
vrhaY0MyZwoPxLte3CT/14KQpS1K/529hR+0wSuLmzUIOVVRwH1e6QRUd+uJmECm9ESc9iZk6pj3
HGmG6UNm71QfEyQ0nCiwKNLHhZTxPsicu5FThCniRdBLfX5oyNwz77igQ6LpLoeGUBuu3Md4yHSL
nlmn5ZXgojTwHM6PznC3xzhgY+fONPsvCRW0SgW70V/SbG955xlcZC3llMXQbuRsO2cGXWCfIeRU
wb3xqjiBciluUkDfgx11dk0EpNtfHywfe61tem/JDzVCvx+1Ky2+nrMmoE4Rbo/Vq0R9CNIJMypJ
MdZlRATzOI0lTIbeD3lAW2E+P461UblLLVUfHyF6FpHaJpV+zah4kw+C5Z9c9mzBajNdLzvwt4JT
kDQCy01tbCcJiuqfO3AB6P2EYuerTFbl6i4GvZdtFY5Mg+ayxMw+WazSdFg59vg9kEB1kjWXZhpS
NqFJ8ONEZL2ljqrkkH8cc+uIN1AjcRFU2KNYPLLMFvkfGDnVfAfXs1qL/Gp+cY1tolyZreoxrk1J
Ced2BlzdGYaic8ofX05OL8DfjZ9LOJZ2TCkmUbpS9rn5VDw0zhu/RoJo1F+iEiU/OZSb9zjV4fJO
CWYduPwPyrfvzIwtW7M10EQ9RMTTMVTQbRizRwPMQ72iN6lCwARabU7Ys2V81SPtXTpYe/txiNPE
Ga9N4ku3Uq3/Bx5NaUR0bWTvXOK6vVG5Ox9qUNEiFYvqii1G5Lf2hoLcdTo/msRqpzhlWkJExEDx
ztTNNbB45APXPZ0a/C1FZVwaCgiV40Y2CaBnXlJEMmuHYwDzRknKKyRI0js/4tz3/HArsJ/0nvXn
Zh0cUy/dbaF887g0uBaofGFjS9C4ouJFaan5ble+CV2mjYtPYzbhvgp390W5KXlqBMlocBLm/dz7
VtVng2N3EJ06RJ32actU3YdSundfYDn9EHrvmcWpyWLCD5pa8ciNizDrbnY4C1Fmk6LeuIrLfdTj
v4PXjKyEBoltWELF3tQpvS8xHDWT9+mxXZmpwGc1kpkT7LOJQkq9KmDsjoG+rVb3/ZQrcQS4INBl
dFdpmuMSeUyq0qGQXUgwDd7fLlPbm6asL61MgEq2RFDmbCgYGhiCEr9yck4Djwt35mnu8LckSCD/
ywn+o8Q7bYGVD6QZYRFUO/e50DECVPWHc8EGngha6+7g0cFO8RHVL6wK2Bu1McDHA62rAeHztMPX
b9DsKmpJQIjwg7QdH/jxYJ8Ohqt6PNwo3OAwM6NVz8tadE9Rn/GnVUTvEV27zhAd6gyWB6f+gnB6
5fbhIFam7UbKYNqSUQbz8o46lUo8HsokcLJN3+3uRr2qY8FgTr66kK+1x5iftiZBXPA46d4v/ah6
9gpdZGi+2/XjpPyiHBXfXsxtGwkIqwYifStx72X+nGRXXTTiAm6ajAPcMf9qiVA37jkKx/7mXL9p
78xJHHHVbQih7sHwVhsDxktkyvmLosqrwtjE7JVCZks4ETuXy9hsu40g+iGmuLPvODBc19VjpWdl
NkiV77KNQkD07zUrqCO2Fd1Ss8H/cnMgl9JgwknGstPVMJD4ezfCbZX1r6WPb5Zm+OrkkOGbcX+k
uSbM6G9UXWMikkbkjrdk/Rb17bvRnO1eSGfESk7YFIagwf/DnDp4zht9M5mnN1EzIN7btGwzmDbP
WPLBrbHLmtLZWYnpTY6YBcIk6ug4XZtD1/EVaa5jQgWhcBImFzSyMUflEibwMeJlbvSm4blG6jXs
Wsk2EQSgjQrk2kra8K0p6qUcMSKTCIR34mCSJ3Bn5mTYlsNAbqhvDj8rQ3oKSpNXG4rCFvyF1Xta
g4vuX/zleTLgPLB/7IuJn/+8tGKp1Avy0LOA20dnio9AvMr+eAcAG+4AbcvXQjOZmh668nMTf9Mt
astexXFp33KQPCNTxgynKU2kb4aBziFCfu+dBFivGZf5RtP5PRj2wXZy2V/FHb1tvufjdWszCx6I
gg/rJoeG4ENloz6yxTQ13KTa+9bZQCYNzYyYXXNeUX5MkzJczb3GLnOPKdmc8COmPRZ3BJX7sWT5
w04P9LhOk48uPHuW1LbuEgJ5jYpjk+9DvLmm5TUXn9BrWfIHshQUpuP7GRJNX36RlfnsScfgDbHo
QraNtBACdlag3JNyGNzakqd/EeNOLT1zFW4Ms4KmGR4faFSwi23lBdeLJDGaDpSNl2guZGmAs+IA
qNRlwJ9f5F/GnfgBNVXDajb+W0+Aoiqmju/h/PWyQNoKQm0cgdxkav76tuugdBO20pJMVR+JXoZk
nYdmYlkngh90Vv3nJ7qjpMK8+upoFdusLZZsigh7gX6/hbUhhr2Rf1HAK8a6AquPQWC7T9NfWrKv
ib6d1qwNFgEFwQFT2biIeGegA4/Ch3efp2BzWzKqcuusYWsRCINwEubn7/SmCSNDmB4ZvAKL0jYG
sT/s7ecqcz+gA2fuv0kX2mq54hFOr8ZQSSH1hhkhNKyE02ofWFXJu7G9E99di5CWOl1YX/i2lt/g
G3aAOUBJXpCAR7OhkJA6xEaePn+xYmUhBsxab+HoF3ifDoVwlW7/MN7X4Jneqv2HAgNyLkelp9lL
51wswd2DKavY3wovnn0EgRdlPkcro8Ec7aoZFK5V14TwJDeblZQagDkLtZ03+kMVkHICKge8pA2s
gUyLuF4LbByDwQ/k3p5ebi5wH7xrjwm5kIR0cPLBzFBeh8FUT9NBdFWyC/xFvlxcu0Ao9Tcp0Be8
OusCDGdiMsVKOL+j3CzmGiKROvXJLLK47XpcJYI5mVtrvuEqDZQkytIxtzqDmKUmm3++Tm+tzk/t
u8ynwyOPJDJg8HEiWV4P3hBbow7V4fQpXex9rmxUb3J1xB9D8B48MX/IP5cem55YrFe4dxPTtH+G
S3T/J2PHtgypR7pJ4imS35U1FRYIC3Jt+qglhFL4Hcblr5qJtylMRR6Yvp6oepfNasCD+OL8dZKb
y1k6Z/UX438sKkRIZvVXEaQTeXeusmREURogHaIYbuatAhS09wOZMyGVps2EcpF1LZia3vLxf3Dz
TUq7TDvBiIMO9ctUVAhzHwZrMnXx4fTDMjBNEduu4mShBdQB7iLzyKEQXdICA3pfzhlWGiUaTU8+
EXgSEUhYriFNEoOMCAWNmaLSqsb90ULfk3SvK//KoENdwc3KkjicTYv6nvgGRx9IbBP2Wu8Xbr5b
4ClZ2jZJnvkqErCRI0TjZ27UyedJfCx9jEuMcbUbwCggpg63QUdPWAJK55V3iiCf+L9POar9YZv/
/Evun2QqfjXWFeCEH17rxDC1VwTzuStPYKXR+wcd6xs+kjDhmMkAXLYVG4gzlKVSPdSUWQme8mbO
AKZKrMwa7Ew0IHssswuxexE4rtOtdDgMyFYS+h9IyFf8mXbtxt/V6VMiW0Kj/O32RZ/T7QvUMyen
7z6oSkJiiHB/+v6PZv0fGcgFZdefkEScjOpBRMbU+D4CgiC2NPXX6WgJOO+P2wsW8uFsbqh2cFi8
qyt3E2KVzOPad4lALjEsZ8T96dk2IuEqyy+0bol67AQLJv388jtsrSB0qwxKHEzTbdvyE61i7Zh3
IfAukdGdJB230mEQwFVFv62EULZg9CQ/gJOXeegdTqEp/YJ0kOgcI4rcOoXTLLTNpiBvd6BYgw+I
eviwosbbm4AzGmg6SsjYeTxo0DDZPaVyEWtuV5fOzL49gs1Q+mhasiz93T8wdkYFOwys5evtUyFP
ofnfr2BYhUjC8dFr1yFHPLVsXDkMgRXRIV3QPZlDlbMv8l7eHtcI2ZCVOLJuHn45N0dpmbT2mSHW
fvBxYNhPoDltT2m4JUGPFcG+gVh1O9K+CBAql8HfSzU4saPwkVTSqeNr2CCd+BCRix1ck4v7v5+U
rR8kBfM9H/PZb9xjJcwiBYCwuEdnNHEh4ooD6AsBiMdRi2Susmu/sbTaVj3urK5MSQn5iu6LNO1l
Vmq3svOaaC/TRwVjqjH+g4vmRv+IbklOcchZXV2hPsTd6ePG4JdobBnHQ04WC6WgWTfJoF4k/H/e
HzyMHYZjEqGR51dtWBZgx01kriOE6D6wqUEHl4fTqAPw3rwxIqqQehzKpIEyqB7Lo2PEs6Wafc3H
uG2HrVKWMX3EKC2dH5JHPm05NMdD6B7urGLi91iNlCkJeZ8A5GYDoOr6lMJFHs1zu/CuYzpv8Fyb
RcWUj4u9IqOCCM5j2x+ZIY/Jvx8SGmR0GeGyrN2TRB8Whrxn9gztEFH9ezv5vwmrkc5CpPG4LYYO
DDWDzOyskd2mF7hGqj1R+KaWXvn31jglzzjo44nfvs0k8yvFMlc/iYFKobVcEpdshFO9iKEyOrrR
8nc4OnLjWT4osYYDWB4O3FELryhS0T5txCefwoco4b+lmsGmLTb1XtEs8TN+Mb2RF/FcNDhL4yyz
mX8kRfDWacyG/vf1XmIEMuw5wterivn56bxZJbgzFVbqJctjEjdA/QwXiVJbLg6ofepxquvZqPMY
PFC933E7ZWJb6ACvweELiBlP2WbZ5TJzIUTLVfs98Sq8JwtpqIYOK+tFZq9ig+mICJZgFnTLkVn3
vGGo+xoFkYWCVkbuFblWDk/Skg/BVN7Q+5Kqj8d7UMnkFgX0Eo69t4tk6oPh9X25z2GrQ4Ad1eCj
QO5t8H5BimIt2S9mpK2Fy8BsRt6Zin1G/BOsvEv+WNF0lDCD4KO1FW2AV/mpBovFKNLPDl9Uq2sl
RJbaoH96EVZJz7yo9tTOOW4oTR+PO4g9VQFeFsIUCEBXpTexYTLmhcF7VnRZbMgC2AAD2UYIMl2w
sd3yBrLwy/sr7MjgauZfC8V1koYqmmJG936xSOEXzwZhTNHPZ5ZPl2R13+Jq/ylt2SmjeVPe2sB+
/qsmX7F3ErlmN3m3HyLXhCNES9Q12cdbI38rpIuiwYLOnOSg8VmQI+mlnwzcCkfp86jLvQbCz05r
cHpXHA+wGWwXav2xUDlhtLJWKYYu7HrqzXyP0gd5KL+7wI7qt/cHWu9M+QFTcj2ZqHRva7CS/xyB
BclKzq16E9UuA9dwN/XksdlFmU4MfFdvOp6v3K6YQ4pqIXTWLFF8YTTNMlCsg2+ZUFiSeBwOS0EY
vGGj6qP+3ZzXIEBGQigJwj0+0yHnW+eLg0gFWd3wzVE1N0cqZI20+Ta2nNUtftP1zpyjWQtc1g2H
pLzc8YBWtvCQZI0jiKapQCZwdGchXGUHqSDBRPeVAdrJBmvGNhIvjiRirEmMD37KPh4n8dgG7+Rz
Wns5jzY4kdmUfN47u1V7RtW7r/kGE6bTdb4Q70JB4Y8O7WU0m/MDisvzHuPC4UbSiAn8Mb8H04ib
RL2WABQYhDD/tvEGJK76hQaNuvjbMS09Caajp+92Hdv1tvv+a5a2KQDJMB2Uz+52EgRDtdBQKzPE
KJsgusZqJopT9ur0Vl5B9uAwIsdaiVUi3s2UDtDZsC2aufCVNHLCvbPjFzZdQWHVZZlyUduzQTGO
TPLo/3HbRw6E/lr3X/cumXM6yitS+aqBllsSMVAGVgwjXD0mbkyC4je9hWJ72zuMKKSUjXG7Sqa9
JGhZUShvAuO/8gdAZPt3alQcSU2rmQSW1aBN6B7uwZ89xfi2vhaqPyDPIYDgJ23opUvQTI8BpeiE
H56qhtXI2yZWZRrE5BKsKA1Nqsl6sQc6VomkO3eqcmnZFDJmmV2Kg98Gu2tQ6aE2PEJ+BiPM1utp
GO4xty8DXcWxfr5uHtzyqZRFzJisVaZwBnxw12vGRCI+teRMTMcLZwkZnBVSB9CLCksbhd4V7+uN
Ln+SI+N3e6KiGcPLPh4ZpAidpjMih6SezQmcxwP2/Uao/rWvdFfhIGVKa+z3EIe2rPfexg31Ze9A
j0bwHlV3NADuDrkolB8M5b4QjuFKyfgy57YjYWgKXnl0oXvi3YT46l+P8ZS7VmzQHhdvgM5FL27g
1aqWbL+eh0aCXIY0IKT1Ozh4ppqRhGRKyMt2FQz3C2EbfDVYMkXVGqJeVtVzDeKt1jgHt+/7WUUu
6zaL/Vcry8tfphFa7otxx+83+G7PaN1BmgQ4hSsoDLxOotavYOzhxKL+/0QfUr8VJHXROEFxJQwd
dLZUHOl73CMrUmV7TJIYW9EUPJdjZy3LI5eLcrZsohKlgJaEXNNCY1yTESVupuwZ9xcrv62rMiZJ
rDIQ4HIUqJ+Esdzkzrt+J6uiAsCm3OfCuzUvSYxyxscEy/uT+iZ6qtQ53F+XDH1v+OSQaAHZIAyw
iniIN3pud0dwpL5OK+5KwJSc39mchibCJpnMFqjK0eKWfpKf3JLqdrYDXjO9v5nxP5+HMubUdFMn
mxa8PFcbJM0/QuH21pRagYTHcuictr0dVQeisOIEyNQ1wwpEe4trIUuZsmvyBLPV3IVKBW2M37FN
tCTkfrj06cNPH/qS1Aa9lZNzRHc1L69KDZPxW6opx7z6CQeWqGsxRlKBiLWDa1wzPddVoaTD13UN
defyVRTIafQzsrX78W/Hj9MNKlX+Ny6KdfwaCgAp0aHhmf2cvlCg35Dd9WJXzXmfQ6ykiA7KOj6o
BzTHOS3jHQXXY/ML+rZVHFN2QVj6nlIIDIknK6QaBerXRrr581qaZE8ttR8/ESkgIJcsHZi/v+5F
5nyEol+QIXtvs5FFt8JVc9+hSIOAHOVnRTra7WCselhvziwz82mXiEJmzk7oUx8SvH26/ai5nOW7
GW53C9id+ym/386Vs4ByALBpM5qrMEE8Q+w/XAjzt8uAYSuTpL6LFWhsfYKF8UqRSS/Af1KtDj9Q
sK6ISrjnOMRfcQCWzZ5TuVQheUx5MwXUYhjwAfxRtWbtN641zGHlol7SGzxgg+1+gOmT3JBRc5Dq
QIMShtl3GkUxor77pSYbVak/WI8XvcdZ1XY241H/QYY83xF51AvHbZuDTo0aELjKhj4y2AuSU+tA
Uhm/0b7fjqEOKEw5VJAzB6MNKmVrbeNv+1vboDhdj3XB7sYihZhK+bp/u2N05NOuXs4gHhM4HEDM
4M31SoQJu3Ks/kBHbIsJDeKTaZ1J57dcQpVltKWTzg8Y6GUscpfIkkRDbGpjsNpEljwlwITyILvN
r66BnNYAkWBbkfmpxSxntX1Zda8AoJi+OBMo7zBXAjHZtChoQ99QkzMXBIyCACOuX/k7qFYD8yzK
edUXwAnnCtTBB1Pm7pEu1mQkjapcG4MpWFin9MYPuydfNfJ/5010dlLdcAdQO6J2o4VwzF1EpmFJ
HT7C1SB1Kl/52yw31/uCmMRPNf8s7jYLXdaloCEIZn9c2VenJuysVgbfrgnElOfx+N481Cgm0eL9
W30E+7cAheZiRrgHItzu8WewH3YseWnaynnonhCNNCuf930T4KFcHX1VBRV71L//l55YRHCCbCF/
3wmerWjayI2Cnp/aHVOblPyZikMIrplu9zgfcJ49N9slL3GacjlCfohND4ROTW/ykQtwViSyzTdw
mkOuewDZJlJorNvQPm+wanjZyH+5EJUA7NsnDjHyZhpbfK4BNpssh0RWcyIFqJC0EmfBGdsZo4Ne
8ixACCJGjHfqH7V7tCceF73+W++Qgw4VP+PVdHQU3buFtDEcAm6vw/SCaclhOM/ueLb3iqOvRZjH
7xKyc+MVkFQJUrRkwXgmnisvECDvFTVFlMeyUQL34jghpBlJJDWzoPDG0YTtnr8szaJ0b+4eLQjP
ge4kPN/c3srr0+69gmbu66pC1IfEKqPi4AQd/PrdMBefBHcLY221vVw2jFE59DjlNSqfqhs8QJCN
483phRr/J0T2tnWaVJdP/MeioZWAemXu6R9ymp3r8+g5Xe8RWTKOvrjBh5GEQa5WWgapCITD7fQ5
cJZvXJbcdqBtxJ+6cEuuNXw/ZIsDhqmWmIbuRUpoPyusIb+ZPEfnGtvUF/7k9U+ng1yD92hvkwnm
nGXjqAoyRWlECa2q1PtLcKIAuwdrHpNy0UfGsS9F/0TSYYfp4nm3dXtbfAMZk2jml7n6g30qdK7k
14osDjr9K3EKPP6PLEWjDZcTkkS6pJBCJNAe4w1REs9TUqrjkEF45KFwS/o5YMxaotZRIyMKeh4b
Ar+e4jImUW92FjpPQndlvtKLRPdmJPhHb9WAtxmz4wzGFZC45fhXsnQVYaVQ2IR0doSiFFWuJXcQ
nK0+GSZqtC5J5jq1EOh0mBpOHK12xDEeESOK6g7XcRAOSzdTFEV0VI1PjVNFvYmVLW6KHFP6Dpbw
9BVS+7mDtVop6ignxLsUv00vR75b5ZcksPPNot9FUSey2B1RXJQyfEkSotY/32AeId8bd+3Jeqvn
0c8EwSr2HnHsj5nde9Pf1TjQQHvjt6OGe5Ff/A4ojlSmZvyBHUQHcbecT3+GJ+cxWri4KIePryox
0pihufNeyq/O88toYcvrAT/VuvCIS5GR4Y3T3ukdouzWCTgvy1DODKWVxrMlS6ApY7thpFHmCFzh
Z1fBjJulBlmSOI9VHEtUzz7/Ru1jqIuZqpp8VbkB++h0QHFWs8TUTWjjGVVE10zIzfp5gZigRiTe
mDaeVTTVemoOsdVrCBrInwPd99YjfXT789HUPRcnbLUv7/QczXRw7ujqfR/aA5Dq79oDhulyeVnK
3AZWb55xsNq84P1SYtIdVcWCz95zV2m9XG0FeR11Re4Q3UEtDL8BhSoqfvEMMsfOOLmx3z+0n/us
9Srz8Z1xAWN2mjzi//XEEv+l+whhdppuArai3CTxofwY1l9Vd1kfLjGWmw5C6KJMvTHR6BNBWEuN
KeGdFDYd2qhXkMHl7mZ2UFFjHfftWnRwO0xNkIPXj+APpRtZsG9rHDZdC8G2a8zxNAXyA7lvZrr+
/W/o9vgRViyVv4v3HnBhLjT4JxENL0woljMCYylKkJz2Z7AzIDq90OXnZa0q8b3FOVZWfIzvf4ox
5EwCAxw6Gl03VYyhSB9KoGrvLqSQmWCxdrcx2bjDbeQbh1QvahpxM5o4O5Ng3Pgz1CLyz8zjDso6
UbaVim5sskQqqyZyccEGRxMtO3nNR5zxYGU1bLDJZbXexcgyA7vjPR9FF8TnyztvM4cE8akWYplC
oELeZDwogG7URv/bXBwmXUAFTE5bSyD8eAKBEhE4Q7KuAb+CZnQZoMffnUZ3gL3J1UHWN0vbJIhf
lZvDL2l490jFFlaRodUXK3k33noaZTVRtgu/bOXF0lYsdfXXgbS0csnyVHzML1OhiiX94fcWXJYJ
bqPAxDCUsAk3sMllC2pwb8VC82LSQuxsGgLtuh4xQ7vjMO7gSPBBtG2f9bGLmU+bYsR7/ecDTwW7
+FzTeE+R+sc749yOPIN9zO8OYPnpDRvx2sFgsMJbKOch1MBXOzmBsjcizNvScfRng4hJAHpYSB5r
01mDQ+ifB2MemkevXxSOY4Szr1DhV/gE9MhIroDzEAgWOQ0YPNY3yH30iD9r1lH2t4tRIs/9fhPx
kcpzEevZp274x7qIpcaUbfcXQsAe7GLhlae3f34Skr5ify9oCy4dDLv83Nn6+W6QbGyHDUiQ+f9i
E0WJOh67LzJ8bvvggHNHHacJCN5WiMVDpfdHrwm6nxOY+JZmI6p7Iqn82z5Bq+Xsz+BxF+4aJHB/
nrbK0pvP6EresBZdUim8zVFVqL7dkSDFFW4Z7+oTaKakxzJhfCq6F4PxXmoVZV4D8OiPDWkUTDY9
rIE30u8AnWBrHFj0TlnOdIlqJzVk+//IAEE+FdZf4qalf2VmN57UODXX1ENTJfyQP3nRZPQASWuY
KOaXe6a2qx8ej5tjcPGPowMtieaW2xLTK+vYTmnmdU/OyB/sAmRKKbce2Fws2giDbICiA2ErqINP
XmSAJ97UASZWK03/GzChsgAJZAWdFcKyu9iTKmzTfIBhMKJdMhp2x4PvurjuATqGMyDyqVF4ZeRS
eXS4tcG9ZnXCvoNM+tOYfnSMwNsaCmQWqpfyrXBJ7Hg+8KdBbrKpK/z+YkCZAifAHiMZuOdrEXt9
kULFo3cqlW63QeykNuOkmCV0G477wC5EFi/F1VVmk180m7wHP062EopR7EMiJ8+QQ+O2PoSSfG+H
j3k4pUhs+IQUXAP5/iKKt+wmLaWl79rBDRnwoAonoYOQZb5YlauWOM+ftBNCRSlx50jRYDsaGWNL
zfqaRuc5SvC/vJjjqgSsVwn4/htIlCrHh/XeAwuT1SIgTVFR5oqEpwHfHZt3NorKYb407MhNrrA0
/6k+H3QAGPdPIVSjxJhaE2C/5bntev1qNaBeAaOR27qUcXDgyAXv3KPqait+ByLyTZ6IoMpG1DFQ
q5nbr89O3CNfWn13W19qhDacyafGCGAkQF/9f5eHLD6RHj6KbqRNqlSIBeOO+6ABYbP1haefkdrb
+mpAg0oy1rqgWd2g9P5aVizpZHnCzuApeoUEtuXM3q6GlVKiWJWlTO7p6OsEwJ0ZGshz7pqpOOi1
C5MQi8aB/m8qOX/FvlGupBicvsCtFxlhD+ogxcWz5kIW/Qm5eDYNs6xJEx9vPXJcqbT/z1s7K1tH
8ioXEIAqGdVFqgVV4E9TPM7FBVmvjd7KEHM04F4WEG4mV9bPKnSscrU4J0r3ueZeo7gMRYY0/AbV
rk/KGUWRx97WMgqncXJweTVvanA9qnj5w0rDvs43deRtPFX8AA9NwyQKlS6F/4/ZfzNp8JgycfBI
HK8z0m9zlLp2ZtcSQIZ2K+xWilX0+w3mDDixZuDeTBoXwO3o5hc60v5Z+OT3jIfbA05cnLS9weu5
G2DVRWO3Oa0DYb4uJTK4RW+ofLBXRiWpqOpdIhyORWI2PlWl0jOW8rd4zabF28lXahjcFY973CII
FXGjaesfeKvpiALkxF88ynefd+A0bS9sCljfkYpgR3xkVOppheSvFZ5ZwYq9W9usMKeWCMy243Lu
j123ZhmuoOd8St+SjHy+1i92y3P1miSeBvJaiIPBgJj3uNtOuTcWliiRbLgCZuT5aZfLMH9HmtPC
NE6u+XLq/Kln+KVqDXou6Wi8/KVAgpOd8BzWXPEU+ExBFWV4oXh4Fz8SlayEOT7Q2/TsgcGiApqe
mXszyUvOMYe7g8cQK9IpksugSO0VT0D+ZEAH+DwZVuTkHaPRywVs2+e9RuEQLt8H2geEDaMrQSX0
lWs6Kqfk81lrHbrWQl45GzaDRO9V+4kGOjGViSGu8AQ/2UJ+/RA6tlJ8RyokH8NXxOLQVG+KFxuf
XVNiwBx0g/6JGtSqap8uEXgQmL9Xp3UoczaBvmoH7A1rwQ8qefhT2mIXdJy5QIUPemh/XJS3Zheo
SxM3f68lwpE1fnZ1AEV8pYNFQ0v1ygK/3UKbm1bDr6c0lm/ZqbjsKXdQ2Ecg2TfIb8XiqWrmOFdl
un/13nNFlii5frZFI/ow+MxOCfojTFLM2er0nunJN2OqDKOO8Wntpl53nvelN5W6G6P4MKSYtlNj
zZaK0iIhI2a/TnZN9ojavCO9FU4IFGTaP9/5ZxHGZUCKpKh6OJrXJocjSFrNgVS+027FBNTjsGOc
rZ0Hn0Z3s5RsOUm7n6JpxFNlMRW8kSm0pc0JtSmF5B8QdLQ4Jn97jhRUw2NAyrr3PmkuD+5CjpoS
J30XXNo3xDTk8k7PXUU6K8SOOOY38hIhtRAvOCtmwlg0tRioE/CM7QId26YxyZebpBHv+AhFKKXE
dz+gdiFkRFW/kUPKcJXSgALiPqAY9E0/7gx53JBNbFLf1GztomG1sDFL1s0jrBsg/piIyZVTGAjC
kFAkWskjTENuMyV0yP4TevcRy9hbFnd/sGjnw98iI9ZQMa84uchTGG2W0FLtHdx8bX5cBo3oJZjU
tB+8r/BayVk7CiTKxtsJdFRHjwRlqNU5E9DObZmIeUUCwrBliMtUFlyiS/HPf0hYJWi+Y6lX3uGZ
zcka9fhCN8EFK4R5JXfBOB+qEuNArS+dVTDn/CbWIzRrMkoMgyqh4yKbnGXEoSHYDygiwZVrkk/n
FtNnDVITMTzlSqKoB98O3q6IyZG+0Xap++VT+rgrxoKHYvUVYMp58C9i2ZJLjcPX7r5aEcI0FXl9
hnNzsKRXLT2+e89zuz7mwEV2qd/yxgkM0wxS8WmhsQvb+sQdIXARUSwj8TN5T24m9vGVLqhtMUhv
CsDtPcTbaRdiWPa6rkvcb9agQ/yI50WZUm/G+KtvrNEacQDWYqkXoE7FAGs5ZrS3OSM7cCMSqoje
GeerkpjgnBHE4phs5+rE7KGRVVqUPZSe0c3ieUgwliqeacefbGslkBs4hRQYVKxUxBBf29qqvRa1
dMoxjYpYtFEfqQK7C7skEtxzmjwybILHYCsFJFSif0d8clxu4uqOhQE81jTalhIYobe5cGIbTHNG
AgXwEeBz+h25bodIOhwHN/ni4BPhdeuU/Xb5Q/wIg0zB9r+y/SmJtnlo6SmTE50eLgtkh2b75X8M
Ir5wkliIni8nNla/0IKE+1VsGsTXAxm0Q5qCr3/j/FXm3Olnj31LxCF1MNhX0qLHGHRjVpXs/H0k
a5oCBUax+eyCETqGFHG8c6z94I5nJ9pXH+IHyG+YBlMUNY7Cszf86exY+4nHVKq1GvTZ7pBHFvqU
Uaa1G/nGGY3HkZrbNXRxsxj7rD3fBVVzWj3R9INnibklC8XNKgJjV6yDOGavzMwHF0Q7tORCKlx5
RHnoL+dPxDT0FLR1dUR+YpsLxPdpm8vnmNTit/73tVEQ9CeJ7vcXKhgObQcaB7WX4C4GwcwVmmlg
COAr1stnSlmpIlfXiAlHSocEU/Pc9eiYSRAwOyzcy3D5HKrBh9Q43hcElB2SqzFRgaSOPy2Ttlv4
nRGOI4YxidVynGPZuYb8VmhSWhTRpNhX4Mf/TM+e9uHaJO/BWPe6hWiTSocm77Q8E3hxuzY/7nIl
jmPh9ChwdQ7CXwrdBK2nLX1za+WqrfCfYsVFyrNt98IKVVnvA1Q/xGPP+MjoSHxeb+nXdnqSgjGp
FpAbOnhe91XaffS+rB9mhtg3Za8xx1qKsu5sLtvogo3k9US7VwdUqXQJu1OCVSvyxK+aDtJlK7d6
pK1Hwn5l6CmIzfb9kytpkylNqgXAjMJmMWDWtOCPlDCgoQyBP/Ghpj/4Tg5wWbhTI5uqHDJurKST
GoNYJ99sUsOT+ynY11CxjfjrYoyKI411iVjqlHXErTDU1GcXCJZrVlqdTlhLu31cmSb2hAjZb9uX
RygyqGTvyObLPBCkVBW+X+hQ/za7tGsIjm8jSgAWpvmcaZtrCNBD5ozfhHuloKW8SmOZrgoLIgDq
Jjq3GGlt1oVx+b2wBxOsknnIaWGaATHcfyMk+7S8+/7tsRSo3NR8kHulCTrRqbE+vcydmVmG9LiH
kAx8m73fFNqUqmjtPT9+ZLqEXDLeWsCjSxdC+UudwlmJhdbhaquAO8OILg89OJvbc1AEiTYv2hkc
aQyyo66xMbnn1z9QkSPpB63iKW6iMS1uzD0hZiQc5j7cJ2n8Lt6fg6cg5yPSJgTWRncLf9lyNdoz
why69wYoK9zojG6NigxNbTUjNBVJ3HP1VfSmDsmGaiIyBDtnA8BvItW4QO+nUQLck+Ck/cLwhkoC
yKj7fwTSeI7JCIzYiDnNpY1S6tdzFS9vey0yEWBpkw7+gtgfnAmEmYW79X6Zf3vsE6BwfJIMq2wm
invodVFMe/HF1YDqNco7LclByquXaVpvnC2UEYzheBOV5N0rNVEd/qb2WjaqSBlqQmr6+PCO2NRi
l0mDTeQaykoDeXr4PULvKEXeXvaR1l3px7aoGFZoVX/X9Gli06zLe2iUe0pEVQbi0XmlMVnuPeXa
TePyvasKVG9b2SXNvYXQQnumsJxCYkNaZbBNJkmptDQCRvrfFTGkgwOvBIFIQFpgqq0r6B/Fic2U
ac0I/hKc8bW16DKn9ynuB8Y5xVqww7azuHutY5pvaVT0TRc7Cr6T3D8qnjOS21mLffvkPGSWuDqu
ZK1NPVw+wmJksndPTZUyeZa747i8BnP/7VmUGtyYPHbvlOEhAhs41xe1fiXWECDl/oCI/mk8/iVb
eYgBC6ERU4K3135euMtbwozMLFt8kWo1PmGG6/p21LAMr4KAZSn7f9dso3N/TkYrXSvgt6T0EhBU
XQ42l+czJCAkqdpp1OIvJpya88d50FUS5PdrirwFPX74RpxyGN2b/W82LfhIcnsQH6kLPsQE/TIJ
lcTqkHs8zcyNiUz5mUeT9ce209+VY6zYCu1mFWU1A1lF9nWNshO0f+wkqd9tM2D+xoCn+s+p4EVk
k/aSkBYJp+RNaXdBhsjf3XMHZ+VUq1DFpBymioWE+ecb+50zX5Qnl7Tspoc2A7vF468NCTXgL/xs
dgBlIX1nU8qS7Bf/fQd+hSD1TAGY9yqJ6jz9CCKv8FcI6MA/1PmmeAvJSrD5a4NNIfystHWijdnB
ZKW3L+x0OpgIdhXr2NgQJ1MA80iZ1qP2dWu52ozaz0XBC3CN6hNRGh6X57AKqogHiocLTMuCGEgQ
aGzMXpVrIyLc8fl+ttWsKxlxLaoISGMMCYh34UzkkncIocJDY+6o2/gBCxWlTOejC43eLFEh4YeR
FtnB6Cdfzb0EhFlyjmN+wGid9lxmn8k0TLgXMq82q08G/Ry4AcK5BUlVaqYpsC+BH1Fw+PYw739i
q70JU1raqFFaswZAxd1yHdQM1vDD3It9Ev814hy13B4H756/iItz2wloWu5JErCd6cfxApPxUzJd
KgXQsGt1IAPz9Lej4+pYTTSOL2mrgIa2KdRTdu/ovItKiPOEpja/OTDcBcqJLQTZOSi8tyNBYJpY
vqpxV5esP8LI1xjYCc1VevY8m/nVEGBIsgxBsRYKepjyqBEk3yXaouk8ZV6poUv6/+3RGgYaG7qY
3V8KcEciWWFMDNehBFEnBmxiuNL+vgmckjHqeUOZqfh2JKlKFPuPExjWCKRqainFymS5tcbU/7BR
S/SUOXcvtk+4nielkNcO74FCGeBcCqA7tWRuRZARkfxveGM4djPvTEPeuAQHvggmPVU8ieLfDzDD
C4AZZMCewghfsJV84fM8kDxwxuR+GakOMS4H4TcRlFK5MelpMsnwPTAnsj1Z7eiLOBuV9cS9ep9p
a10Qv9QgnGKd02Y5sjsCUA3T/Q8JRRuGfFVk8H0XMwxz4p0A9gEl3cgkEoMaTewsxGT2ycO3RLOA
+cK5bIZvRKzHF51HpkkCJcbh44X7ynwnJIayRfNL/IKM+UKVbe/Cxh/WK/8dLusXZRroLT2HXBXq
oYwvk20KD6N4zqaKY4Q8G933DiPmPdVj3h+DDhNmPAvkHqReDM/25itaxG7CjiPKDjZfm7rWuttv
c3dy/MBOw9c7uyAFF3JMEA9w/WwGufi/fgvBXwMbDKzFkcuGfb8yMeAVtlt8weOA4j8+bdqIDGle
eQZPUCZNIiG+c2Ez4y8hf0cIcExL6JGuiJ1vWkc2qjQVAW5wpiyoznhSs/HWtGDrfoHHnkBIIXTc
pRVuGAkUjPitiXkwgdYdhenM5uREjcp1G3xCQlPhByAMGsoRHY7d6A9Eu5SXrxNgFplZnFush5NP
lAQSUbw4wkLqStZ7yqCpoVRfRMyRg8TT1MkjVqxtVPjEhdPMRkatk3+J5Z+85pCXM/GPBE7bJ0ZW
sRBdxXShMtBCHE1QHvN35cSnOr6y4ZQENTgRM/BCuYSnt6kkXqf2MlBRRVa/CaC61ChMik30nGuK
aQTQBpmwzh6kiVExusMb30mphcWoDEun31TH8bw5l/9r+NpUBO0P8GWfhY1zQQZWdzdzfYTcqkPb
0p7JD99fgTCP6jmoHvA9eE1d0A837dr5OjnBysqci51sZT+XrLDtFvmexlOMrybxgofZ04bY5zdV
+sLw0AH+/f6C8pad0RXW5/1OWwjqU4XNS23mdTgQ1Gl93HzX4cMug3VIR48JuPCV1a6oZ66Mqckj
WwubmQmjF8pPGs4X9jZIUXFQwc9dqfEw4BBUq6SaIRvgqntQMYuz77hU3+ONJn3jJnLwkrroFqT9
GiNnxhfZAYfxN8o8/zmyBC1LGSyUBPrw+WcpfhbTVEILvtxTeIZDfC/lbNB9nUtbLZrAyE0VyWLO
Q2hqr33I3IfcK+3mfbZ4fZnPpojGYHhtwx8s6qKc0AYJT0u15JkGHR41byjM0r4AGb2QYQKzDMKF
5XY75EyDbjQkEIZjUTof
`protect end_protected
