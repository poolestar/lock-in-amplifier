`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
iZLsMvzYxl7UVy1qksvkvq5F+Ify2SXhnMnnJ/du+/+lFNPcpRV85a6SGmwM6fvsxk4pSjCeXNqm
2Ubaqc2mxg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UQbYQdAeJSkAWsX/lPzNC6scSmoXfZDV630edORPPzNEh+jybSRTRuuCaJ9IXoT8iVzvKCKAR1yN
QkGWpPRiEhJ8OXTA25I6IbsZmaXiflvO7MupLibfpUyj+L07fDiYsePPt/BcqO3yBiBVoAFdeYK5
bHnbL/fUnG88jJMY1eU=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jo9ap/fNrLfE+dxA6JJ3KSul8laZvan6VHTnDDxOe3VXOVXVzPItuuJ+HusOSfsZLkUytmA15aSV
gQx0uKf0NY0nTPRNwHWnkZUKsbQV9FajRG4878AVzw5XHuTJkFAvxIPDDwu9jf0nG5nOwwTkzT0V
ClkcaV/NpzSV4a2VqXmiwYfjW9T4ZEoYD2q4rj2VX1UBSEx2MRwzHhNXVqPehN2ru+JQwa20DVXR
91X5ca88BMGlJnX4WBOcILqinT/DJI4N1hOdHWHV1b8mB8ZCFUo0zjughurelEbpSlDcZ4XttFAA
OLd6KUNcfzo0hKl3nKHyMniA3eWaRRwEaJY4hA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Q5qiDOYtq8Tp69As1Qua6kt5SXK/cT5jdULhAEbBlM3hiEyy4+/g8+S0Ob0CDq4WqTPZoHuOD42x
Op41NLGOUOVWsd/2ZDrVnl+EyL5t5ssooOOVoeeENd2/QDT6adpfIuZhe3NsaOSPXog98P6+Qqql
aB4I49m3Bn5DrDo/OgA=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YrqWkZu8lZKf5FNnOeiWG9Fb5eUlWvcESSzA4pHZpVvfz826Teg/X/ss4D0XHwYz3c1ROB/4YzaT
E83zLtZGbVxgSYu9zePNM+vf0omIhlPKdmjPDXw0Em2CeCNjaX8FnbMcYCzBE1YGEQvyIPV94IkM
+lPMnVgXF+JBfJy32LSRLflMPZq7u+Qn+RNb/Ven7G5EwGctMVH9l73DTRnFIzrgMSd8hAGbCv67
N3XNuuL28QrI+hMBvbYU4GrpADMlkJKb5AMFyfwRIZTyF3gT3fKeLJB84NCehjVd9Pd+cdiZ8Mb9
fEXz2PbKgThYgep2dHDkj366YO9rSXHUKg9P3g==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EIDbDab5qqu2YU2pLrvR3jvVJUgPeodJJCXWJka2eBuhFJdVaVun4knhjbB22KTQ8R224R4UgRZ7
oairxCoLr6zBMiZtYQb3TcGEhiWqLweaDqnder7RyMrqY9x1MothAHafdQtczJsyEp9Ut1BFWZjc
wlQxG10iksWTm4BQxcLG1LkX8A2hC5YBh++XA7nEW5aOS5rRU81Ogfq891N5doFKjLywqN6jB3kN
0Gqhu1j3JdYEBObO0mmnC7DxGLRjCEW0oUx5JdMyZbAUHIYUP/71YzFGg+Hk3I5Hw0erCNc8Lypb
JnFE6otWjktlATPfEms+jVIIQvb9NxTvxD3qhg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7184)
`protect data_block
nILhyQsDtKRKZmw2rzM+0qdh5RwyA3oBAsYg1TRq9DYsKCPZ4RcyBvQz3IB709dbZZQKika+HUk5
CGFoi20jvgd9OgVqMWPN7qti3S3uzAIYA2uE1HNhNo8SDcLsSZPRkkXXr+I9X9vw2rhMzY4ky4yJ
OqpvTHEexi/OsacIp1f38o8Zm+nAmqlELJxzuVxjXPFFiox4UNXMgWNs2Cok0EUFzGqgtyzVYtiL
iN5XyEs+cwz4aQp53FO6jEElezfcrcK4vtZjKeep8EgJjKjmIuOxGZeee27zJA9N1NJM9mmEJIxP
JmSY6eQurx1H3oGLNGLlzBjmE1fS6n1dFB2mZnL85scR4xOYtL0/IVcmoIIiBjtUwT/Ewd5b5sXe
wqZ8mvbhXJpvi98HE5bvLXQWyxL8F9rhEYHRsLGBCsHNomPdpI7b/SFRiJ5SvF+l8kREi9trpCXJ
8Hzv7bmw1ECEaNOHNQCZxmcw0BmTW0vK7cnOTVp4ugmVesr1Ib/0/pM37xcPAej/BGvP2QtKhsob
+d1lNinP994emv26G+m+7MIJYgO31Mnuj5tAoi3rMiI3pw5fPWdJzUf13LnyX1Tz6tz9Dhnw9yLc
TOkM7aNlj75styBYPENvOIF82bAg9G0MURLrcFNRLKBlmW++dl6Mv/Z0RSZSL3c13HPjnwPxRW6g
M9uV82+f+DW2J2DxJm7XsDQeHFzrqz38ylIS3YCAuKynGtyVbOcXrk06xqPvFFfxc1RTCzzxvopN
o56J3CUqNycpv3YCvEBxBT2eTE5iqfhbNcG+0AMgvrQy/bkz+cr4bwkaO7mYrxHn2YqKubLyph/D
LTUgqS1/bAcOOG73XBlHrJf3GZhfrJcQjfZLWq56t0QlulPtWP8mt1hq+J/SNu3lOz99x1TLegVh
A9Y7stb78w5qwXscXj9c11XS6+nxXJ0IhsXq95hEQIWm2xlLnl+cUkgen0QiTJfnT7ROXeNKIKrD
I0uI5/Mr9ixHv0NEPlQvUeLOUyzCb9S2/hWtohvsIgiPfdYF+fzJF3Vf3CRTKQ5IvmBdZx8eLOxE
V2xHJsNp7s/7eG+dn75x3neeAfRCJLECWVepM+znw8VLtANvR0PckmZTsIOrXFAXDQupOwRB04Xi
Nya4mUxwlaOQdFiXb6i+/3MzIG3t/wSn9u5H5Og3ygad+bFBAojBjE+Bwovt6wPDTa2ltoqshC1Y
XLub8Du2K98LfsoOuso2SG8jWiafavrYob0ZTUSmJveL/qsW1ukUzicBL8vufAiHeS60c3iTDAXN
o+onuBXSj7vJGEwitTTBmUwxyxk2kbJhi7+F5FSj7JwY1dmHeW+jMOBxtU2qSd6RxiyP3SJTUq8+
xCpieS9inkrp3miYCbbZIkUTRaLdzztUwWHmSQ3/kjBIO963sXshcZL8LoN8yIyUl4A5DwPnHUF4
Ay/hhpfgxBxTLoYrQco29ozlF8+TfeX/zBIOz8kRgbEkIMB/vwZ3f1S5qB2k0OxHVfbGhZdCTWX8
ytN2w9/SUJuD0KA3jeOH/VfBkIDH/ezFUPbv5kb6oR3G6V3tdIh5mlSvl8vsG5ZtDOhMS9s+8Cpi
BFv7VuNg4v+YLFBUudFgEtFAfpeGU/CC5/K5uac5AovOPCrCxBzVj1g0rl2ST8hy2t9U3WuoeFtD
U8ycb8kC4gVzEtWUZ5okK+o4ObcrgY6GmeBDGBEe1vqs+ONZNwROJVpjrntklbHBr03OaLTfG2LM
/0oP/SH850CpdErHbkY8P2r26RF08LUQNklup9XVzXRbK8l/XAf/wMBkvWVRKrc2Gqhea3yB/C+5
pqXDbu6+QITP6Pm3sTxXRMsxYWKWbI2MGvHo+UkbNN5ujewBXaNLgD6LzgIrbrwoDg5HEuZBDhAf
NXofdbHOapliDsrS56BiukvKp+lal56JA3I43kzGYL9WThZNr5JbQ5H7Lzwi4+Hv+PfxjVeD79yd
75tYatDR+VPPDpIdJGmaUsqT5iDGhnZQn6LkxFkTf15ADVDr2tkYkGpwoupx/08h1+yO6j9yab7Q
emwwtsms7cEam/Xa2QayHY6auZR7UjdAF0K9VeRodHXglP7dSHxeFAYq6qhJHytpFYyK6QQbY4MD
bL4Xx17rR8Q1yZAkur+Rgp1fBsvaPyyBgPivAHFeDTHZXJ6f1D3FE5xlDO3UBAXNFjHOxcowNz6+
vyEffrj7P3Y625aHF44vGUFsZNxnn9k4jc7ivIZAo2fTBsf+pRIDVMhds9aA2DG8tC7bTBVFHwwo
qwRYFZra3YHbGJPsw/7J9gYIl9v1AcYuSRDdopJwwWrTni8vbEcuFkH+226PjS45mJ9uHvNL6iL6
rXb77Xsdn4ebkT3ySsq3eAc+BTs0BWHS5QjCgOvsX70OWKg7hBxTJLZC+FBRJwjOrQJLmVr3gMLo
t0xQuyJUjsYzNYZbjWYWyJdMD+Ywf+MarSSHasfLEomEASh207AYZubBdIthgQTAcQaNx4t6jZL1
6QRGONXpr7YJqBgOOSEgX8EN7YEXvxN6lR+ZCmlUpKm996eqsuqAvHNtVKYfAVY9KOLzLnHb2tnH
trymo1puzBJw/qsbpxt+RMdnWnmMkur8zE7xoC/nvdEBY935ZsY5dO1SLxU/yPoOFWm3m+2DX3bB
ZbFspCpRs4zFhp+90kaobyVQxG83/Qs+VPUBjbNgrUGXhdGDn90U3n2grjaWT19TCm1EAJ+z6WPe
TzSgwsBV/TmVYYlmxkuLds1lBwEbQdnJtLwkbEe5iFBQFG2NZbPzE34sz+MKXxPO/Gf4w8ka6k0N
SvUmFkdl9oMMA6+oysA/0cjk4RhqzxLOpl62ixY+cF0/3wH+uVdP+ddhKNjabu4RBDbdiZ2L7Z1o
rm+ky9O11SvfOiaMfjmW97vk5N6gpC00vFH5oBtt/ScfX3BzhoPxmGYUXjky+eSk660XDf0sJxo0
1sewT1Ib/FIe6h2cHj27DQzWFljOPLZaRQeH5FrXSZqnMmg2jNlx9oEDTP2yzsfzTRmMXwI+SAce
dhpvX+Ln1w35bcEzi0OcIap/KGlUZ2KHf8UwZRlnkdJkKiR0+OtZDS0U9pxvC08/hfbjNJxFstY0
GYYq9nNAyrknZt0vwmwG4I4/6JIwcxtGEVJJ76d2Kgimgld3FLxqbzAgqdjMXstn8MpfsMzxdeyn
xtlxXsLZI3nEH6+U24xDOvtrNhyPo9C9DO640rYyJwdeKrMWPtLu+6YwMNmkTwaPwX+uCC0QAViF
p3dNwR/sfWk4OH+ECkq2jzX55Ug/VW0kjK7gLRnIjzAJNbfj3I3epr2ykkhZOHP1e6pfJVMpZkrQ
a6k8Hwe3myzhAzwoF8oA6YYW2M1EE/qQA4Ohsp/JTU0f+3BFmUknkkcwbBnWSnFTGc7nsPwSXh4Q
HQFeI22YxpCxngHwCS6+zpL2oCX2KXTtULdyG0Uv3X2GPiZg4a/W4TZAq9eP/qKY7paCml1bn4hs
2XRDQGKlxCjKwTuhCeNZszNRu3rA/j2/xxZ9z931CjjNumqkOZa5hNOgIIxlvGRqKt/imgZlaLBr
0O15R2bCIGH+bwSrICfOPfbuUnTOYRGGBF0fFHhSs6+e/cmNGo7rEs1+1u7HpzpEXeWruPkuW01r
FvSYdVW6F2UfD6slx5ppfH6lye0VZZc+k8ywsvxus42n0GS7cuK5D3TGF6yrDUYYrZrt2wJWWsQe
+AiqO37L4RLF3nlFMwWT6dfHv5JyKXntE63R4YEJZu6oFdsBnai94TYBOxY6BiroR0h7s1kYJCxl
9w8pIlxTuFVRSGLsEsnyJ76JjeJYKL+dINl69DxnyOQ9TUKOmX1TMmfBpIpFHJgL+cQF+TIZLeGt
0XaEtyrIczLn/ScTsRwJWXQK810UAkIN3F+fRbW9TSsiIYnexRFy+/6Fc25s9A9W1SMRYoRej9/g
UKgCcfnD0CRGu6QmwtrbWDmaddhSrhwNj7k4hGoxxiP+PZXPrbwvzJ75A22PFFHJIfu3B2uPnElU
/EFLWzHVhGcrKNs05YL8pS2fZCNGoMUxhiMm1ixsyFkjw5IPl5nK3aBsFvopo3gxrOqmXVlcvP8J
BsdUiuK3+oXebK0r9dQPHZCHwefuL2ogT+RnhIqgQSDLTbmoslHPPW8k8JOm8pzPQkIppHCPY8p1
BTlsDNFDWorR2GfXO3iDhOercOaoSEgIonKJyzobNDHP1V9oXRnRULX36Teo+10k7em12Ha7Qvgk
Mi5O+tFAj8vCD25jbLhA/iTUyOLyuh4aaONtuBWmDU1R+pPusGE9Py0n8BFwGzZ0TX89T6iD0ulB
D6SJ3IjjdmBTrbBCGeBb918n/msa8F5s0KgDnC0BVTVGBG2wbtJpPQTlKpM2UDaWV+SBAbyKz0/z
7bXI3T0Ss03ZIPzPc+VhcG0rfpix/xTCCnYEMRBQuUXt0KTLM/xqzpnv2IB9LmS7FuUZido1dSpf
t33aq2xg3hTOiLuMKfv5h16l6IdNUVB0bOG9VNWFJ484dZO4T7ESIsXME51JaB1wrItX3V7bjgui
9+tKCHYrKig62RQWXD0nreEl9Kqpi5KJ9D7ij8qm4/2ize3UK5yroYbRCSPe70ZxN3U8pc78n3YS
ZXYfM3GLpD7qQgC533yrvWg9XyYn0eesv7d5HRVzdASqHppHnUtVM0o937G6dcT1N3bu5tp4nvVy
68p/oarWLcPbTNRkb84xOZ+mLONqGPP5K5sMYxpIQuFA7NIogbowe7mTRzP9yPzjCs+51tPrr6XS
+JlMLpbshKOlm5BUIi1W533ggWVTt1cEk29utAM0yolZqyrjgbq6UhGeoZKkgm5WSWzBGyvYfcdP
bLhgsy4zaufUVlwb9mfMi23lhBJuATQf+q9brFUXQRIzjxabe5f+9g1GYrN4FiG4BSJ2EHxggLV5
fWwWJjIqWPPClyh/JUSWYejSZspynIBjrt73Ml/7If9c3Y0fimyoQp+mCdueCvDxmU5qYy+O2Pbk
I/bRYzlL3l7SdkvupOAhGQXFVFm+ycr5olkhRDrTJtBeMnkYyr0BqqM3qvakv8lby3DQ1VZrQyQH
LoYELO27BELUGulkT58bLm/hdyCU5EROPyAlXx4+3DbqZF74doe+EOCEQ/2TNM60aF+hd3oVe5WN
nGsNgNbDHcBv5wyh8v2iJLOR1HCsf9tzgWacFfwyHe3eNbUFMpvmlhoeLhlel/nm9WPKhe6Ne6w/
g+1PWqFQuDHAEPswH6/lCiNqnjz+ZeT4CrUt7rp9sDHgNBkRTVL5IxVRFxSlXmNK/ekaIKjNMqJx
r7SzGcTn6Sw05Fl4jIaHzD7Ms88ZaZD+QJ4nWs7XoBFXdoYTtXWGOLvlm+EWQfwDiV33rpaoslug
lo/FfXyTlfW2Gt8lZrKv+9z4WyRP+HKwlvYCs6yoUwCn6uTkGl7rtZ96SqtpYIKZ/uXnhP/urly2
8XYALaHruv0+mogXdGV6evpzqPN0TYZ9flXiRBTfn2bTp/2cg5eUTDJbiYVHDgV9kxdbrifarTuS
Vw+Nd1aTYWN5gdggCezc4w2v4LTQTNi6Z/yPafGvscsKHbd5qBC9gkiO1gsJXICcP33jzs2zLL+H
E+6o5iyDtXTA/ZoXKAURhk3wrNt9e5cHwUnnn/2dwIe/j5PuMYZirmiYESbYGKjXH0LUNphfIb45
YpyX0JdF9YdJbm073dljvbkb5pEMa1LO2EE1lHrVI0lNJ8dQ9tD1KSc844yrIa9yX22fhPwxsmFH
jYNOppA42xrvoSR+4HPUUMRH7NXFF73U6rjqEWPU7mWcDLHTrvnuezIaqwRq+kP5O+agJcVMijmN
pgz4Mh78KoeSydg9xAib9MfZ/id0mib0h78xXu5DYQ83uax4bGe+j2ciksbIYzjUeLFVLd+c0Wq8
Z2DKd9I9uNUmoF3VYy1sY7002wiI0EALTjvF4hJ/8PmkL+wNthxbBv/Bf/yHk1Ppik3stEN07S1g
wF9fVMpR1PaMwNuUZSu7QzXX3V0ibwd5dPT24HHGNhb6jvpin0AnACoe81UmUfpmWund+3ts1EeO
NdleIbG4IW8JAyZG4jdL6g4VaxRfuKIEn6WfsgfUGaaoJ4QvmhZ8XL+7Kb3JT9QC+/KPYVToZLyG
bAjUEpjlAaDgV2/8OXfG5CXtLU8afbjAbeXnZzFXDvOAJVopYJ+AsOoDKJgD+lNaoYcKcCV1i2zy
JPoD2EwrnYZE56krVM1bHbPqmFGtY0cWBMrKYKOrIeN26ldhqlFwWy+bhITxEWRYsDvHo9nMc2ur
ykJVo3OcCh1o/TpwU55vVn6453wORqMuvZ3McDP7piZOMkH/1gsu+QuIQc2LkLXARaId2aIr9aAY
siSA+sthRkyfcNWvilTzD4vDk3OIUqA3j7UWHZzmjn81qOv6IFb4UmH1RuwF6NGeitKuMe6N1uQU
lt7jW2dD0vNBpnV15Ic/v9RyMHfG82RSYupdBqovAGyivDDgdGjedEs557hFq71j7yeSUE71V1jC
Mb+Xoa5RDuEiMWhkrzJx1i2xfpe/P7u/5xeVtikwnJyGP0YIOfHMONIMO7m3TeLWcVc0GIOi2O8r
koUQ9np7djHvWGvDqjKIs82+J9v/Sr9XDaNWNGIacNb/iOLbemGig7Zu0LWj3ieVhm7SKomhA0hD
ft9yEOmG8lo2wzb7f1dd1MndHmj+hZxlf5muoW0X1mqPAg3Qt27icWK5gwVK3nnczeJK2VGlb91z
M2lwd+/8+QF0klsIa/f4ZRbJd0AdvukmKNFDYzi6jdE3swKpfAVdZgZvsru9S/4LpHAR9AGcroG/
uBSCYxqVJGCkTqmJQAQPrg8nCMh49pL4+bhE66fSQFpzOSF6Q9ekDMkpYxmLxbO0EccF/HAfcny+
IIdg939cBBToJ83hDA/4q7bprBRExBDbFZ6GUtPn9z0eUP/53aT6ErJ+k7eCx2L+fIrLd+Hen6Zu
bhkSy4HXMR5aCXAg3pfcIJJlYQ2ew3XMVZTSBAUfIMDqn2KgcsBwB5ngQWPrtCxQiDu3Eqo1MSxY
mxXfnr8YxsWfyvyPjp2FoMtCGgNOpZIHMY5HIWSZWkj+wjedcXRcviFJiGcTNN3OSuniYvaP3ZSF
v0MHr7kStz+L8ODinvGb1rAvPrpKq2/ncepNnUMhDgeK0bEzOO2GS9ipRRJg2b3G+Q/FfA4lbyss
uOug5JynRgnBVAX/iWsQ98peI7Xy9ipyUffr3XmDoAMQEy3fLvSeP6bIsvHIjSJJskQgiHd8+3m2
G9SoT6whDnr4hEcFq1UFLQkpuOz1f/7X8w355rYeyAVBoidZWKypy+C8rqHKam1N4Ab+L8/dg6XI
TPx27w6UVcHEEskgy2z+HgDqNPYYTfV4GkCkhbb5RWmIxCAlfEkMMj21I3tJUyOMhxxaIP1ySqGu
fpaWY4TUPaOnA5ozcNKHNHgm4HT9h35wIdmw5nuigAT4uW5bGIRWEidjzJ6lGHcvgZuAQBhvB2Th
7Oy9rNcovbSjgwQqz7mP0jtqawzjEaREvKZv4LX8Splc0Eyl/ZQuQc1awXwIjtnMhw0R5nMYB4OE
wr0Kh9JzXOkXBS/fOVOs8wN9t6kNQhrWeUEaZ+SmIhhUYRJ6+SXrZ2WdWLBwfwgGfiDm5VnsKysO
67g8TPImAPFEMOvS7qsbaJ/XBrS7NApduacufZiRKytG669t/MFI82rlwknYoHXXFpyEdwx5SmXS
n1BslaJNipsMZ9nS7nX7FhQqBloqDRxt4AXxvrKtNIQXf+06NV7nsXEA2CMXcbpmqNfy8FxzP8gl
KEcXo0bvhIqvQb/r7DI2V6usr3/pxgjPpUMhreAm0bwPprsTMlirmv4CMpj01w5bz0zdMnJQNXhi
sGbGjpzs8EFXsMkbItzoBPYtuNsP9aGo1zErpVdrUJ3yyPZJaXInlgvMjTwz6y3721TFndPup0fY
bez4d1UnN2NQ2TfxIWyRR4CJKfCaKNjSQgp2Nx06yr3XIfkacKfOGOXwrOFGq8VpFCn+uCXOUb+h
6Vh8DcZkLhjzEdzBjz4h7HAmilQLo2YaLQSVpYqv1uue2BMu3W011247JkcNvIajHLt9NwdJsjYs
lxsVT5AocjU3XLCQ7kEtm6ftwPqM8Fd4TMkTYw7NCgSCs2IE1DtLv28HkgQ+IvzwIDEgVijjIX2x
hT9QY2VAEZYTWL8Us8Vi46gZlEjvL1dcb8AaRgPvGeuNtnbdSN8IgGoFB702QHTfGigbD3+/GD0r
0ITcjR/GIzoWLcxc0A2ojS56TzChk/916rH+uVIgEDcxkGcxgC68rWr141LYCHkibqpP5W/gRFjL
/TBcCToI2lUwbM9Stg9dFBhv1JiMTH/mTlH+BZ7of3+33Wu6/u5t4ER8wD4Y6AaIA5WFZW3w+4xZ
Th4j/jrkhVkqQm58FdV7B2DO1nPGQL1Cc6JMbK+ZLBWWJQpavmx10EcRGSZ94nf40ZlpRsLuwtHj
6LMKt8QtMLARkykJ/4W4LezMSCJFpOjgonhLq83YBySnAek76aLdvBxgwO41TPODasXQ6vNR/gV/
k3kTvaZa5DXMj3c261U7um4OZyLa7txtAyNNe8SayznKX37/4DJPjiJRynQT+oau/20d34/1tja/
EtwtOqYJoO/MQvo1nz3HV33U3f5uvOAEzjtYbLy42mMWqPP72GEsLlpgPg1x89CQvWnstJBIlQ5u
XRRj9HkXEMO0rQ9FvyJLgG+mOH3EiYCjzeeX27NVW5UJ67wwaqROC9yROq+oa/1tudROsnV/399p
qXQqhzuvXgiStaqAXNO+WYWYcSq62cHGFwTehEAhiv9J4TymuVIIvPud7mlWW04TsAwP6Npi576c
8cWaSarAPtwNCDWbqRCz3Ups2I9vcDG00OzCOmPl3NTQfVn1mjWJlWc6cYTYZnsVtEn86f/jL+Ea
2s0G2abGki6WOC9hemUfHuS+Zb1xgDyWwg52p2S033srCqILYNS7lavgyDqLVGDn1TmQkrZLz0XK
K3GpIwMJCJYhVQ+325HuxjOipH827pztpc0ol/9G1uOmwaKbXmXP3h1Bx96MoKuEIFnsDPU57WoB
iCT+pkiLzF0neCDTYKGF4VTTPxbn6OST01FN30N336rhTHNU0IXPlnYQnRNKvH7qID+fnAHvf50x
fAkUGofCZ6aYsXP7cdJPqTTI6PjNFditfXtKDvQXtnAyoVgFoq1RfdnqmqniWRlHwIdd3ye8mknU
YC2tJLPdCQTXgvLUpqeAFh4zMXaTGlEiOPwNC+UkioBJEw0Eem937ZMqrKLJdH98OTG/HdYD7oRs
SGfrL0j/jB8tnEquIGElS9Ofv/tp1gCoC8aQiGYsBwj4DV2s/9iLSbh2G1BJAp0KlA00LNUiqF00
aDYm5Sfedrrb5N7Ds+QDv6uPPKNFu8b9Nbdh60GXs6P+mXH5oruS2kgZ67UOQTkbCvz/wv7pg9C4
1mWLoYq4/fd4U8s+/pgE1FVA6ffvDgMOdq4Oryvol6ejY6RisBOSjSF67bEMWK+6i7RZ+CuBBgyl
p30=
`protect end_protected
