`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
PeqAACiKacdbMOWs2XqEaCOpUVm6letI2uGLDiD9lX0yoyBIWN0n2TcEOh3r3UNckwNHImxwRo1k
8kO4TiYYhA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
auZzPkb3r2HppBydOd/o3UXtK6rJTIS7GYUl6UfoNc2fuxKNxuaX5fuwuO2C/xW9Dwhj6txvdXSl
6P18m7eILIWtScQY/zFG6rhvGQKvakLwLjdAKDz9A862+2PgGCnRM2oAlF5f2cOeaoejq4NzIssM
trMP8apt39JggmVZdB8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
e3IEv7/wkdd2X+qJoUq7FlGbH6ss4+2Kprvx1c80iL0+RtyfFn7gRQ7KRscg+b2pSX30CAA3rZvD
CipsqO/c9bZqj5VfXOrjBqJgQUrqinfK3Gj8SXPHczpmxpnKjMxM1XpBs1v+GuafN4/8KAQ6I/7A
Jq/CcecuA7nqnwT4KVIDPnkeewZOWMG0knXp28/+fOLVIYeEjEvtOerZiTizJTtPwmRPVBH+5Hql
/CtHgmxLmpitZvSNmWW9DqPhkuyODcInEJrl4b4SGqksRts8kQ0XcHH3B397/Q+FarsF7xsdta1b
9usdtMMhglSriQUPZrBPHJXV5L05ik/uuXMlTQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
LnIK6f68C0hy0aeBngl05Oyvlp8vnvOvN38tYskLxxJBl7ej0TpYYaSJOAL2lQ6FLR326CCaFbhs
xgb+zjGCGs+DNfMLn0hgRkl0RBaX89Xm/iK5zeBuUNRjw6QgyyQJYYPDbwCrfTi3xoJkSoIOaHFd
3wNNZCBA2WEnHKz6aJY=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CeNA35IAS+fDRdKelCkD/EK+Ucq+I3G7pjPDlBGYhFEdN5nbyHo1Tmux9xdwRIy9QvlICCoBH21L
SGTVHtQEB/e0aTmfNHUbwSEwnHaM661voBhLiRTU5qQpjAS9zNbKrA5T251UZIbuV7LOoXyp6Wn7
yLcqDCJ7nNnXP5/aFaTEPJV72kevkZNB26SVxFU+ysrxXeK21y6rHIU8tS9pfwjRqFWl32wBNBZy
c+7uxdI/r4KVmipuD4kHmdb7eWXM6MKrMSjlgWvKiolj6goWmzi7SRLQT+U66YMNp8BfQ4XlcT0c
X8Dx9zPFetvak2ROciLf902FNilYtf+vhnmdWw==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
c7btEZIH+CfFksJLkG9oOMqjkJg8WlX8pEmrfA41RU/4n9cvzFdASG+OulihbL7e8ZGDk9ye8tF6
4FRVQH4GOMia26DiobkTbtlNCIbQNYQQA0gZqATjTqU8oSo3ORD13OWR8ak0X8/ikYV2tHfqKP3v
AM5v8u0JTb92RJ73Tu8S4JX7VYwvRstor6o2UOK2t5I0EVDSm0q3pIekgq0RtSAfpZcEmIQbR+vD
Qi/qtGGFSRYICGWxK647oJL+o2/OS29tL4cj06NQV6MlPIUUyt0sgT2hr6dPjCig4QSycBLh5w9J
KvMskGHNUDvoszKAr2v49s694p/o0Vt/btsOkg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 600640)
`protect data_block
EflAiSgk5UuDa3iO87+I4LD3g9WT+RD6XpTZ9NTGD4cT2AjUw1o1U8B5vsB+VEEPo15MtlyZD9Qu
OfIa7LXZZYSeua4ze+zILXKqxwZ/jMhcbSUdWL20tpdt7xoiV/0sf2Yuc3jSv/1vkfBmrimQigRI
yo0nCSVsHkbr4MvMAAlpjiGHgSK+JrlCSoiaf/flolKYFqlwEoJ2bUbWal8dNWOZ19rfzQ3wrND2
vgegBA0Yj2JHmEB6Zi4JFtDw2oPCYCTP/ZvJW3KmGDMh0S9LUqkNvp77VROPNEb3NFmNhOb6UG1N
0eQ67QelEazL1PwrMsS8mTtQELyERRKqx0W1vgdGSwEAWQc+GL0hBv5mZWLNUQUN2/VWIs62Mgqv
WogOFEclaRwMyLa3vh330yoGPRe/T2cH6Bo/unSM4jkQsSk487sBVNPKretXR0iUMrZUTBZHtmuy
f7kugNnKRfdPqE5XXqiXqZWldzAmZ0gl6HpdIQVdJeQJz2Ht37Nv/6aUObeqiBZxUq793qrcZVb5
VEObSBo3xcy9JBesJLqahYj5kqM1rPTjRx+12LzObn9NiXrxJ27lG/GCT0Wnyh0mfl8OzDAkH/O1
BkczZGYnOBM1OVx5XsLxPaEig8NNcdM11pM5w/iYV+/OjqNYUMKT566kXUsfA0Oz06dgLc8LqofI
8BSalLXDf6Ho51UpJhMCPtDpmlDeoXeKVo5h1CrwjOM/4u6L4FEcsWk02yN51Re5n7qKRb0Qw9pc
LeDZ7ibjyQAOyWiaeG0c/taRG6JE6UT006btPmsdy5S2P/2nhyzrz2lR8FLEQuoKnkguBlXorurH
0gnEp313ucuphkV7IJsYUqi8OTQvOKtFQmtWsZO9kxj7HQXxFHfe/RDq0XODjfU3jUxyF36HqzdR
ulOc65zLcrxTgyUd0kZd7P6rniZPSB2H0U1yh+8UNrZhqgreF7bViig0SVroNnarjzIGOEqbxFQn
vI7PB4v102PJeZlDlDkoZH/LziTpGjiKOnmeb1cbQuErtAFaw0t0rT1a5pS4sJ1d/zc1e3fZT28V
oai0uy1H+eTUZAn1KX4zyjJJSIhQCEJVDUM8YjSiluzvtp9gwkOtVYy3cSbty3UazJndMuLoYhyN
U3Sf3Ww4p6BCCd8zeLVoqjX3Xg+bHUHHVjLW5MuSI/ldWFbAvAl72fCFv0oTT+U12KXG6OAjcCZ9
wmmpcir9bdHIt/w6SeDseTCRrLe7TzI+WFMjEqWcXVOVBPbRwmP/iOdMLIC6CVc+RQwJIbynKhZA
9VGFi8a9jFpnlHwJpSTqnKGdgaFqMRxBO4cnkONBglpymZZUrrPJraxNH8+KaIPYyPFWrhYZ84h8
XLl7F6j0GTP/GrMMFGaUYaF/WmAla4cNMyfyznpYbcoliaFLa5zOv8vFkS2pokVoborXsbOy1PYR
YBiD6DA17GYyK7hLHYYxT+SPtIfXS6pX8XM6j7pqs8uH3o0l8pHCMvVzgUII9mKu4XiQnLQpC3FL
YR0yRIoePR4zWP7zTlwgrLQdTeL+i3/eGmtvShA/+FtXcnqVX6S7JtJGAkiyFKJ1Z/MNEGp92Q8H
/IhNdn2rlK5UAXOxA01XJdMMDVpIf8ooxlMR0e+Ku0BKmu6MfApsvi6fzIgvgiC3FD6kXrUcuUIC
UQ2TfyovqPO8Rzm31RBfIVBKbpLSQYhvOd9VR6vyTACRXKW4PhMfrJKv5ywKwsMYDe8nBKjWUsV8
lxSsSBmPTGLjPeDT5EoJ7smpwkZpHpethf2//tEkTpPXHZxkDDlmIRv/r+3Y0KA+70H7yZsCw2eU
4We3DNX+0ashcGSOAVHaAnZrZcbEi5MZlgHIqfGB8fh5940OxFREwCqxpzYE9xHRxURWDuOyV4sz
gx+AHvaKSyQ1QwStQMTF36nFEVquhjU59b+XreYu7n7kGfWmG0nRK0Ej6ZPuykWFI5dAhjtGUUrz
F/ox6sB3n+JF4qLc+MWoki9uoWt76AfgGYIQE1Yt2LrGoAj/9kijLUmUjoT0bacSWc+UCadA+MVl
hcZw5Ws6tMR5klVPn2AlUJFAXU++4yy7A2frfxcqENDqWLIUmLZIhRmzmYQnoknVqTxTUCLIuqgB
kLXaCA+gjsm5ycn5xv6xOvFkImZSmfQF4xkw5Lq+rCQ4H97uJpo2vFWJi2QpvePYlBKU6GHEcYjR
sEDcetcolwPiNL4xmLkZa6YkT4W3sRiiL/VneUDOJ+FCzNX2F1o0R3+F3dFlJ/LpwSePQoLIOs05
sOpYOn169C833t9Jwa8yOX0jrn5IxVrhX8MP93WlPDBWbF9bHt/TTLX/4VlE9zpXwPFQyVcTWOoX
L9Gya1XoX2g+h22A2ke3ScSEz1L/wRiRU2CCzGtGg2YT/57MpyPdeE8cXqvD8OSeHKe9h/F5Em9D
wuEht5VnwmPAVJTgVZWE5szXju6bsPF5Pa8yzJNgqAqJNuJgSwrPZL61AIy1/y+Tisc6AW22B4ya
6xeuIahqObD8k3ohUgmWG7Q5QGy6TEYaUGbqPX4aEwA6H+yHYr5ERrQU+S+p5Y6lB6Uo9BEqSmcV
eN7G9cBn0DFeQ9UN/kJkpi4t1+Ad2tTpDQOLxNprNYue8lDB3aUmDgCUTwJFsRnLZshp5lokUDdV
UYVXGX+VpmoXg8T6pCKfTJmZvZs0bRCdJSBoVgOSAvyXVfA0jqXcGqfvpyI1UoAuANbSkGqOu/rR
+RG09/vjF4QSJt2Z3/mvw7AfaXc99sCwqG8ZxUaSpa2Bi9jb+csWk9wYzgnBiDflishxQSH0BLwj
rZnV6WP3CJoftCt34F0HwYvmE9S/uxCyG/PP8jqKmfiUERxExkl7yVLjmiCxzRr+AGbRyK6P2oJX
YHuw36mwxnzIjXZFfonr6Kb3W6NwMaEn7OVEJMr+b3RXahcFNdEsrSdCAlb/kEp/anQTxOCQLki5
rRWrZn5mCMpNwLJO0+wAHKTcinrCXji49v2O73DwKvGmKejJh2wJH0//DvkSXD3nnOX202vPHOUw
ouVDkPqzNVetoulstdTrF0AsYl/m+S8tA81KBAlomC20CQvXEIhW4pkR1MFLlXc2tx3XJVUuMya5
uYKYyacQum4FU4aAeXDT6sejhaI02G2YXSgWb5cmOBQ09I2WJqtamc7Y1CdhRHyakYnrNvNWs3iB
yo44lbft5SHVzUrZY0i63e4gptJRMMk+r50rxY/urfnjochfG/jQ0f1Om/r1IqwSiWYk1vSDZDr7
k+uRETfZenbmRfqKWaqAqtUlWNhBHxoyfzoq8Ug4z8MPH0jx02LNkddUtBPSewyvQDi7fZe/pELP
N5op+CWxBwn2kyDOnQYUwqgVxEZIZbxG7J/fxlibd3jxIuiIRzK+kq6BeEmZ7vFwIGdjdXWWrNIz
qYXjkEUJMJFDBkY1y9oRHjZDPl5YdnR18tEp/gg09x7JH4oQY+AW8ZzOx+QXTq0hgGAsq7M+YZJm
Z2H3/6vmhdnYGGVQ71zuXTrD1A+kaq6K2XW/UN3TsrNrG95vag3eyJbsidnaMHwlHF8x0CzkTD6S
/nXsu9ujnBKljd8QBC4vG069kcOhKAKDyci6lUohSZUXso/5yt1S/YHDENOf/Hpp9tuFz3Lskwdw
HvQqVeugz5lkLZRIABhn8lE1tMMVG/U4Zs265a/DDUK0oQJ6uh3T6HOwj0BWsgesO+Lc1LrnPWmJ
/6KW2lPKC77OEbLolI/P4fUjcpXulx3KN32kESDbQXHmR/PmLfYx7SnDoay8I7pzbgPCOnCIO/9u
duWmoXCdAOvoMmAShGKS1WcEIvgI27AdCbFXRp8Gg6iKSumRYIavexmmPfHU8iVRLrexzgo8cdGf
MdPrjj4JvoOcljv3ciB35JvuH5xGJs6YuPSk2MPAXq+SVKbqQp8zDqCCJUiRevKBeuzO/TJ/ZBtO
zE7Neb0RNB0n4pY5gScRrRRYq3I4TYYne6hRRTqN7ivgIGIV7d8Mp+hxHDsbwaUqwwCM5ceIzJy9
QgBxJXnmyHFSoyMqIf+iUCY5tkCbUQ/qd+85cr8Mrf3lG+0d5IhzHvlA/BKg8iNgcE0r/X4XBb2c
BJqok0IQdzFhV0GFOlzD3d+5gj72WuIKkdSSWicf90mhMK4WuUqhs8sMlbv3QCoDx+JaSOGQ+HH2
1dtRyZY1ZO9KUAEu3vtkrzNNeURJvW4N7tP3XPUXU0bv82Vr2e/3DeO2FlLWVv2wTTHbXnvEz1ID
//UD9njAgETNTFqQPMhMaXwzfPH7sbkd3ioG7/0rQ7edjGeJ/Kz57xGSGKoJPBIXxK1wAllXCUjv
/zU6XPXBETjXj1e06zxmdJ8jB7mgkFE2Tv7fbFJzxAMaDhkAwI1PwuZSw3RKp2B1dDCAkiQl114w
NvQZKq+HwXtdHJZjPXOJ1gLQ9sqpY95mDdM0vCbP1NFppWCCEpWVS0DeUBGRdXCpyna1lP1CN8AA
V+xwH03ROU7NqA7EHnKePV90Gk2hyuW4B/akV4KMIPKIdQuKKw3PTVtK8DpN0JOL6Eyc1ziN6122
66CwWG0LgCPVDi/0jKak6SIPrzh7akoOm+otJd4iSaqg3aUWeHxxh4B+4sIeu++WZD/RMulz3VTM
XB/N4ao0+gf1aOS4Lvcg3NKPNYj/fxocoxMdb/RTWIrWTdw6CXNALMY+HQ6si5TUqkrVyRqt5QGS
lMEkHkaqHEpgRVKLQ3M3Jh4tHwcCxKTeA+ttI4Sl7NqY3UfJLuoT1YIl3LtrFJ5zBUGAm5OZvxHy
pjt/8FiUUkzI76WEd7UwvfO9Q7e+pnjIvr6/z1CUXFlAuPxIx3iNyGxDHN4tq1wpKnLcu8I5sWzO
ZXhpS4rwxJRyVCGwql9ubFc80iY6S1N/TyphXghV9+/injrCcojW6doIgyf8h1CX2ff0MAFy9CG/
UCV7X0wUvnbqYql4r7Cr14NEiAiWdXwG9uJoOkeSFFwzR57gd32+eA8cGQ7lNBED+SjClilXlSyn
l4K/eM0lNpFZR+Xftf+weo9B416ZQBc0jKkLkzrXAEqdSbIlp3XfnELPvzKy296yZUDT11SaFwjW
eShOBVNXl6owQUOGHaiFU6KvBctShokpGrNYOAIjuNRB+p9zCkQZrvJ9280Ty24ZwGIQE6qNySdT
dGgaTVRCTmMTaEGiMX/KTx4SW2+bi4SM2t6HF8emzpRH+OArfHMcT9IufYoA00/0RFXmzl/ETj4R
24q5b2f4b0T3QZt6Z7VuFNFlYPddQlzar63P1jtV6LIgi6xYFA6kCf9/Fup4W9ZpVs7+0bOmsPl0
zvKzuyCSDWrZzsHTHoCrTOIPHRj5HULR/fAgXyoMO2H7+AU4RpuTjOwI/mQWu/+HmbqwL/rn49PE
uSfi+dT3NSDbiZZ4rzTOK4VbeOUCjEA5ZRhPdfru+UX4rnpwbjSxkmtv6vSHS10jbiWbkN+N4sFl
0LiNI8xVe/CtYS2cV8hDdCBAPHsfRlaD2Vi5/4cpnzOGdn9W4UoXOWMBfAENS10cQkp1m9nhDEt2
8TKwswaWDDDLFYcOD55vQu5TMbqYsKHK7ZqMjbRJdkKUIFoGdDqrAq5dPcvo0BbQISlvjTQC0D7b
XS3/f9ytUisUiFtceaXeLzAo8tDfLmOnHZEHFAeBkQNnazrByuc/i0puwMupBlo/8UXU36gP/CJn
8y9Vx3XwocGWHlBR2Pkj2Cf44OdmfsvD63sI/wlQp/CgxCBK/AP12L2b0J8dwsfTRFvJLS9CNd76
rILSuK3olztYiQoWtatgE5IqBkDh/ZuoosnaSDfXmh7c6EmEtB0sB3Tp3sv1ZPTEjS+8AYr/fcLT
H5ivFPSLDX3o0qElosF9U/vFijEVajnmg3VR2RImwhSNJ4cgVwQ6IuSSkwYasVJD9c5ePytKv96B
mdHH4uxKrSqM+r58Ko1TIdTXdpUbzmv8PCe4mmZ0pvFOhbeXB9Ud+QEuWQxl4JDCeUBOxRgDmayc
aKYSneXzHTDtPnufnq5GPhs/DxWhS/s8ssNgrDciHrkZ6YKFd2mLnaHheHaaSwQWUqA6uWPnhAWr
pnOPQ4+fAhCpB1cBcTLa3sbDB+A2XJru0gwNCi4rFRUOuA0JYejBGZanAacWYaZOpZHRMbv/BOMI
Etufix5p7d5FSLKxF+wz1dyVImF90d4qO9CSJN6OC8GSbqvJtbB3D+SAZGnPQKnLPePNww1AiCsZ
1l2mgR8eVkCCA5WLa8nhvZ1h6X2hYHdgu5BBR20M2+sF49ovq5a9haWp7ZM6EDDxcSwll8Uljhby
FejQpxVhophtm81OsU+2fg/mYzmXOHr1n5qmJaWk+yF36I5RSIBF478yv7Kw0FFczYdJKaah178Z
lWro3vcb0eOr4yAgcbkA4AnumY4Gc7Ar6CDEGRSMNYj85R1ZLTWwKtplHkIza/SkevvGvzZPE9UW
QpiJ/qyKAFXwYchLOK3tgCqC5GVDNCXpP90c5l/FmAwvg94lt4W+DaURNXA2/3KLhw/saG+BAkGm
iABRl2hlLsNk8HtaQk9AfJlQoQJKkEx2Xz/z3bFvor688ISE1C9SLB0FiUq/JVqym+eWRjTLwIrk
kUL5c438C8nmlOyZrY+rzYQwjdeG54be9tPDsZufT0aGkbAHhn+6UTHUL4H0Ji6suuWoHKmh2Lbj
fdSRZ2VPZqF/xwDnYLrLXYKE6oM5FMeThzcwbpfItCJ4gdNNiANeusWKySjdjdZxJaOn35CG8u5Y
whdfOLREnSRhCRMdmRD4BquNkBtfkvzXbX+3U9Q6vtP//EnqwzTfKG8AlzULO5GVVHgKOKiuGqgB
IfGbcDXZdYIGYoe1hSUNHXSzSdDicW1uZON9OYu+z5ynMK2efdwRAyHt4Fc5OMOlmUnTQLpKTF+/
JDgXK4iakdM7Y9JX7AGGrMAjLwZSPEd+kIcR1fIse/xJwTbg088rVOEnTITXhHdAiOSX7V99aTma
c3/QjYOIJx1URGIMFb2zDwzpelwER2IQ1dvbb9bvLSFtEsbmw6nS2/AlFmvQZi4SFwg2v5lPr87Y
8RDvsGMx85kKUCLbCTmVwwKFlVW6ziCMvLV654sXAFZ7lV2WI/1zfgW8PdTqhIX35zddWQFWJP8x
9a2YY1iklHWT+UZmhqJY6M8jzAjN8nArCtt9LGTaKZ9mZrjqY6um69s+PzogGc5mmwXXBWO4H3Pp
rs70i3o5OEwMTYvKs80badRQIEHoe7PUdEmSgEelZY+FqXG5seUz8FPvE6WZj3zwYcZXJAZRhAzi
HkKj2zKh0Tf1F9W1eDS9K7lmWKKL+nq380hMIGjzOYIH/qm9FFBCBRVOqi0m2T9MJD7xd+EigvrH
xRcPJ2CJ9kJ/LTusGjjoNsb5Tf4/dzlHAR8dGjFFOjbXGW4CJE84VoceT1NGpGW6KAA0jJXgq76V
Ko0q/WyddHMtqsdQr3bs2pr0ARiUmvEWbfzHxwVoLBahetDZl9ikZsdWOpAxw4ib+1XftBz2VbFL
yN0IIV3m0uwgbZhMBZkXsnYTEIWhQ6ayffShDvukhuwgnwlLDaFOSzMqHZ4kCSdPP7dHtbS22ixW
qv0K+wdV2BovUrS7pfDyU4nd9XzpTf0q8YJcrlhWQMjw0CaTEKNFkmJ49rXTR8kA5g6ZCYmIG0Ff
+fUm1+QFE6U21MHXtUzIHHkyjxDrTnZKvNL6fOUQkPCvQ2L/v+l7Z20MQNtlKe3mQBWjeW1JYIap
Sp4sWanvd+k3RIzFTB0RyNVNJDuKEFaCOgKzBng6e4R8EyxuK1dFmB02PQwhuNgeBNAVJTPY8VuO
AsJlaICu8OXXyQX1Nc9hU9vScpmddPQgD82sK1a3RHM5ViUD6a050imzBdN+sFozoqeQZiqZsOOY
nW6nwwnGq93Sm3qYo35MCuilAG9u769qqOVFtAYyRVik+7ztiaK7sJUN2xHrgQnYG6sKeFfsaULd
0kAMGzhOIF+kA2CrhG9uDbpwTkuJZJhj4jlo6NwpLoJXpRFOlFEviBDpOPcx9FSt6HHis6Iqh+lC
7fn8cerNyQ+eofzt0E86D3Mp6+fYa+9OxQcVg4C80Db0q5VhikGYdiJan6x5+bg1guAh2PU0Ircs
PRbP2eMbQ7LzMaBzV/U9hu5AaKyNA3xPmWPno9fILeZDe8iL2sUysC5ikSSdNRYKWK+GXwnseg5x
Ny/14/cPhJLNVMgaJ5ek/6z9b5pw45oKbskFGH3WwFFHSUMOpxGy60NGopBmVQAZzZuWiDsDifBG
osiF6giN4AcPfNeG20HTHQnx2y0LpY/mvwvpHaAm19V+NKSTPq8VOBcn5m5Fr6SaReBF7TRIVhDT
qc+bKc45WlaDxKaRStFkm6D+jfZVoagxvEb7EBCEHqkIGqa0D7uz6emU0GbM75De27zSswrukkYM
MsPv6cCRUrWZlu3CW2ZTpCClr1zn649UcaNTNib/wjI/VZi7am1wFxiKDX6Cn/Qpe475IeMEL5LM
hxIuKGMAsW7U4Melcz7adw/5j8BzwkBpmyItLZ3XxRUwDQD3+vrz9EzSJv+FWVTNdpt3JZN2Z/Eu
++HTAkWyqMTE9RgbmIcjKiZH8fLoZakL0ZULczikA7sNf71qwDvQSaFjJBJNbjphZpoAV/TuK3G5
cusDSgSCECWpWBnBgkOum5r823XP2DNzQmnnjgIbHuP7TUSD2FkTZIdgd75AUb32ctfWswOZ/E9S
oT95iPPY2PbNb7Q37ChQSO9wA1DuwpSykigLmn0H4r3WlSsdHyr7UMokgDQ+y/MWSZ1cXQOiTkOj
bwds6jx9tRmalXtkR2dzDvAEH5Jv/4iIAmm8CyLCQQjmVfwsKrbQOsEv3kWsucks4BOjnLXwJVaw
20KN12RH61erTfei5+nkmvenOAcCv2IbajmLXpsYnTjlOcA6u31ojMNefqAAQv1u+h1nKOzV3bDM
ZRtKut81ITkAyUjj90M5pGGRMmUd2PCPiu7b9/P1XOtQ3647tbUzI9G2tq2iAFmpECsStQvUPdDt
uMEhVWRM5Ayy3YISCoZpRBT83WeOdS7vTaBF8UnQfDH2zjUUZGrHy3ZaqxZSENuQpe3M1dl9mxg2
IaiJ/ZoaxywEC+/ojF/ZLVbaNC92iQO1P8o3d0v7FEq5e94mx4cF1CI2AqahpSazJ4w2LJjVoqgc
UiJ59cXsVlpC5em7Uw4wRCLxlvZu2O4bgHuZZzETBiLj6lijMbe8FeSs31ez+PRkcN2X2qAPvFwa
HihtpdVTvRaBgiK4kaPLaAyXGzWGLtuIU7hLyJNsp5YrLgYSs1LZLixBtzFRjQyNexmfjlTHfaxb
maJi2XVqUi8oXWI772z+WHCQkudRQL+Ujj6JUc1Ktpm39Oof8Kua+qeiS259UEyMKqpOwaAp2Y5A
7SaN/zL1ekaYyxf7Um+wy689heUxEkOa3MrT9cCPt9ai6Cd8rGs1HviJY9jlC7QDMQ0C0PcmYsGF
dDNSVbBajXEQhra4WsUDZ6Xhs/8U01fF4fwBXx+zCqONEhmA7Py6CAE/3mDKUQIQJ1OU39blkkN7
YyIIk8We71UPxhjmvGLxhpOueHyVGWgdEmF90rrJgGi/zUuhHUrbv5zFWOz0lBgMGdQi4AakJwvW
ATkubO2v/PfyWvkwFYcNM8hX6Y8kVjeBZc6xPeU4JS9NFShsJ5SjObFTzn4XVF4jqsKgOru9bMcY
h6ERnD1txRicsSetsXyeT8viVX4W6XKU5ZFOu0FUcrMd/7cT2heqrKRVrLGSmVPIdzXMWsLBgyLM
r9FyrAeEK2lhdnNKI7fwjKfsfPGd8Qu4y6BZcUS4XUnf8MMFoAStez6sNgqsIQjskjhZiylrfVVt
jSM6ntKolp1mS9ErIqnY1BEYkxX3st+lVnAwyTly2jx31Ruwi0rs+koeVvyCUtY2cP2GiKQtINO4
yjfCZsu3wGBCcPD/Wr/gndSl25f4xkgYBjgyAjiQ5uWXShQeDL+Ffm8+YJOeTcYpQdYwwVFIQlpl
cC6yuTHdXC82t3bmVRnBTFN8PXru/GNBzKAcfg7/7MtlKXlskCll8LIl4BETQbsKMAtjjAEx8Nxb
VUOqhguTzLxgwT4w+GgJc5uX+1NNkSfrUiTtIMxS3jKDEcK9QnNPvpAuPKQ157+tQvVyQ2Q+y2gU
B1gxKR4sAebU2jWuJtk6MnFTPxl4Y+BM8KFErNp1IylxQfw5sRf3652sg5P8WJDUhIcPZwd9Q1AY
n6W/UKCDlU11wPcb9mVx9Dnv0Ati3Ak6j8X0PwvdtCjChx1nbdm1QcajN9w9mkWmAJNBeYWW2pF4
S0f6/6ByEsErKAAGkiBO+upl1CueqSlbkZe4CbfGbjGfoH1PS1qClXV/fH4oL6wd+VG8zISG+Gp1
q2G3JrnKKgk76hCMcHP3LWmQFi2wMANqhwyMQgb5AZ+DM3fN13Umr7l9guoJHm6Uf32u6UWdI1sk
W5jaQ0We0AYGGBJpRLj8lkOL+dvNVe9YRfH7UH4GSzz3+tA/88Ze8Y1FZ6flt5bDgZYh1j9HrJQB
3JygkIVAwOYm9LzoS7ZcYgDbnv0uePisilyllp4ByQdbqIGrFXQrXn7gybdSJtfaBtBuQmuxWNV5
vyVYkMkfrgX1mto4BkvjIquKQLM2VGkz4XseG9wsPgPHHXtZ08VBqwM1ReraDwxByPVHlFo5xQGK
h8ZMn8JAEs6DZM3wQpR7Lb08FZy5zjKHPTWaQxn5yHugRWRIIdCZzU2U3GjYnTB3zrCtm3r4LtMI
qwsu31dgvy3Ge8F7PU/U5sKQAQEeSUcoayQlZqhQB0oWAvEni7WjRe2JfXXao6srr9KVhyphMlAi
rfr2HmhZeOxvPBBi9LWWTfBPG3gb56e5/r2PIqJbjj93/uPA8oMClaLyc5rpWklTRwKZAVKLoYhl
iNVRv4TW2RLx5SXn9C2FhTSgO1fvHOcFgXHDNfr7n+yFetVCcwbdNQYcmP5AbQNQUB9klLCtGEBI
xnh3/yU7mGONtsM/+dA7VDS+aXsg2+hsQXWVtNEhm5kokM70hwbPUYCrSHTPoxFRriyuGWfKaPyZ
M+TEB+u+IAn4Lr2LCjGcqkt0DyvrR3S2krbVHeBssfUjhFgwOL3HSRVMenEjVRoQeEgIu9Jd+mtX
2eQPkErtAPYnt+CMmKML76n6Ai+mo0dwTR8Q0qtC3aR075bom6+JaCrVi6OL82r2+mYf4Y62RL3/
hH9NQX4Pj6PywsM6oRbrK67HSFU9QGwSRkxa1OZe5QvOwe5QCG6Dk7OzRbrbQQC5BlqGJr4PuGwF
OGEAj6bDYfhEQfb2mE/DKfQplVVSWXVsZWDI7PYpikFoQ37T3nbt2r3b0PrkrvVb+13tw2jG2bFJ
JZ59fGfDnOqz6421eVJxVaauqBdxCE0wlMAMEhONyVWnq0ZNwk7ldZPuzeXW+4/1WC6Rqsf+pjbH
4KPqewIG4wmj4E7dYRl/kDDx0RCaYp/QEzii/c/UoDrM8VlJlbooXS6zwElxOq1pDkRT308kkXq/
4ROkeWUOEeoZokuWiAxuDOhs5q0+kg00Gf/npVHbbkh2HRlpyQGh/h6fXTVI1uq/AypOaoq23h44
9qvEGtbYFYIF6p5vV6SjGaTbuqcGv0yT+TGIOEeQR4sSQjDoVN1z2x+DR9HTy9bXPTk8N7HH70q4
5EujCv7CnsDV05U7y5VYo9suDQGLM6GxFZwb2traJ3qTSWrbcm6iSwNFOkNDLhrvhm2mNdsQY6+Y
+R5vvvYxiF2/J3DDKggHxhv7JKSsuR9dR8yJ9kHmVc5S63EwdQgxIZ8lLbDA7UR6go+kIJ5uOoNT
vjmIGcE0Kb+1Dh84wTf6MNfviA36ddWxYf2OyaK82hKBG9sg8hoi00O8dbSmsCONUZvpRUWLrBWH
ltFGuabpcbspfN4Qrf7+Qes+Fk7jsOqcHjGSX88Djr/gbx5Qspi75P5ALazss2zConsNN1YosQA/
9K9E1CM6L5v9xY1mfjVpx/oP5wczTORlwnX1pEJEG9K4RdR0BQPO0kCRSqfB7vHoblLUdtjaUSuA
ZOaVjGsDf9+76ZGmOTVMhIRLqRiruOWL3xLLD3KAcYlMDXoUf2PCGyPufmgctgPHJ4e1Nud4V1ZV
Ll9yiZebOT2VXlKkoGAHRcS0gtDEaC+ysg0Sjbq1NmxKFBCWTWKjDttcqoT7bCK2lOy9FA31JPaS
wuBldkE/HOZgV8965RPTPVrntmMPtKnBPTljF7jiYQF5/q3AJxFIKj+C5OFFo9uad/wGXNYZWCE8
N+OnEulWGnSic0IICMeuPqvlOJMvsKvUfOyRgq6hzvoH4eZPnnQI6NdtYI1RpX/Ffr0+RlRYkw8O
GIzXZ0y03Xi7CN+6uzF3W4t5hNgiDk3Dpp+fgYoQnK0ZSwbzoxqVhghoqn00XQEuUsOut3zDrBqV
VI03OECT6Ap4EQ72DidBuEBPAikPPnmIFlmkIjLbRBEOdbBmq+ByPRCAfbDOi8QAb1tIG0pWZAgH
+Dj2tL32aS5jNOB4JcWHpIx7PdbQIi4GuihIt7/7ZrRaKDLP3PQWXDHJClxf+l4QrHW27My+Iw3z
XYORzy0Uul00yFzNu1w6R/tYV23hNE5OuVR1pPnMhDl/8vfZOCzFPINfGX+GPXEhflEenLa5nYWd
l+moKFcl/ZThSYn5RPnmF7AyPz0pDXOrlT0wQKUdi9002ndNkEscUQp2AKEawYZ9NTpnonFtgy6v
H3W+nvBrF4kyuDFQRGUZjAN3eHse86S7fGpfDqZMIGMRu//zEvczic4pVdYMVsqJWD3rZzJBFbia
ZkmiOfQuvatCdQCzBUtBoFfU0FZEaD6QqGEUMubm1PBXs1B/8h646P30Swvp/2e50Jek+ZcAciii
89I3cKiqfW9HtPpNpTi739i/UCGw2z77cxncr8qWLW4FOldnKODqU3DDOoAYi7QZjtPN4ix6jEqp
Qui/KBiFSMqwswLnLfwDlfwEEGVKwze2VGuDW4wx+UefvyE8JHG74HYmv2Eewn8aMdUc0VntPgLu
XG3gQr4mh10RzRcLwx1Lx2B50GUWBANC6zPZUYvzYRuRc/Vy1MqVnCkOEe17Le3C6cRiXhU3pWd3
qXo6iHEetwHq8fqBbLzwLgUWPohqgbgKRx5qZeRdtY/1q7g77dZkKsg7i7X7nP6bs4vru2cDtDGw
oHk89vPsquz8cMsSLPIqIruZ5DaWWl8fWu/TiFz5X78KWMnFHQznhX5T6ZGvrZ+G/BIqMqCFI6nH
iWoTgJjvd9B479CpAhYkdNhD2UaytYzQTwg5lMoHTvNoa2UO5PVwST2EZFAKyHVq24Km/kz7DO3b
AzLgEP2/KAM3yDyfBIdVASRD/d640X5rG+Wcy+2gPClyd1ZambKGcjaMGubXE8JnLYZTnzgu2wbI
fYZMnQubYljCvWa0Kgv3brvVXPWLetv7tHptQMZh0x1v+a5AVz4ZylZlPNHO+v3zxw0bpPi1nx/+
B+i1H2wB3lYwmop54rbi1JG4MTyYTgB0QpBCUnX0GxOhJfXVtXExgxmHAbHceNqaJp3xpXKXC8Ba
s5SgjPBTOytWHVH6ULRRDYzA45dvSqmX5inRWn8gBQTuD2IPQ2pm2acpIEzvjo+2ZxgJuRl/29R1
8fmCP0/tLkmz0DEo8hQ/QAheZzOL33kw+aLrZucFw1G0nkn+/fL9JtXht6oiBiAs2CLs1kHa4LnM
3xdHIWarq8yI14vjkf9XZer6lYkbH+BkhHPWdZKfRsxRGOlgcVdWcNDAeH3AHW1ncoNyIhJfXsUQ
JfIwXrpOHV7qmsPs+muXHvCTWNjxDWp3AyUMu3Wo1of9ZYNzm4RZrEZzKjegJ2upM9x52IVdXcRa
Y61bmVz8hgIv68oEv/IOMT+C4QbaWuSUdeVxR+tPCFdecCdOVkPml1mLdGygwlHoRN8S2zf9bcUh
pXrO6hlLSHtGtbL5a2aZKxAfCTPKXSdVvJLRb0QnhfIH5BSa6BiMfCYztDCZ7ZE7ZSvbXmFXYeJD
YI7o1Oxbv5DOkZG8KWInl2NZ0vQ49lkfdK1ZIThQI0GCX25fvUlp/GJVj0834G2r535dWTqoQ2mT
Bw7uHKPmPnJH/Gpr1WKQ1wQJTDqF2ndCxuQ2TVyS6JtaVOJsWzsfokHwUtx3sdxwZVbzoQzoCczR
/W5WM4+Ny1flzLMAU3tiem1MYsIAzC79JX5mNqv5eLy8uC0wU1WOe/kHip0S+F4v7BJVtEjDFqB+
Y0B1Fry04KSs7hKueyPkfK74OC5uCLgZd1LBrH8JyuG0icHzOblJBx6+QKGyw3DBp3QfKTFigIC5
kr/b7moIIMFE7PJ4N3iayV8k/MJTzIT0CK6wZ+AkbyXYzmwzh8VgdvY3bU0Y+8+/xC2hOP9Vy0RG
acfx8V5wxPcaZQxWK4IxLk1n8GBt9AAhOKG6B16cYvf59Xa86Mwemy36+1HqOND7DPlEkMWPjgLS
i+CfVBqhgshBprFEUfiHuq40J5Tn7QjRoE7a1Zso6o8fC2MqPTaqO2GKUP2G6z7nyM8bt/DHYF3t
lAD9oLelR8HHzaMTd1w8UFEjQyzIGoRwSpQHxMtgw5L7IxXtSXPjWZ+OpnpDewYOUBbfL7Wi5lxf
qQCKECf9MZrQHa/9ovkz6BZyGoJLWX+lgbdnN/nk01ATMuCYP+ObprbksywayMQby1Ugyce1ksd9
VvFKdCFWCIk8F3tnEuC0d9gHwQg0q05PRew4cZvULPfk9gmzIwPNh4H2w3XuGznRFTRbobQ4JGDz
LM5VE/0pwpqBAuTF/or/ybnJsCsdeEnl/bdZbZ+xlaa079+ltvW0B0Un3UK5VmEQ3HtsnNkIckmu
gHadhOb3Fj4PqzH9n2Ywgn8v2mEqaUsEhWVQx6XxOpsHchzB0OFvroECV0jWpgK5uxISZNs97e5u
r0aVETd1QNUudWdqAksH9U4BbX+mUxITM+R5T9w1P3/+oxDVF2SiZFZ5CK5lVi39EoxD40A1rcQT
sFKv+mnwheaNFLMjOUjlsjS/g8/WEAC+4NoOeMqcQ7cFQSnPIxNq7Z4UOWYL3CZnPD+2BruUoBUb
Bfu0inb7FMvCqhxv9cAy9VBw/XPp0Ru+p8Ttz9bU8g9dmH2jBkLvYtn9Hhi/r+lkqelz8nN4HqN4
cd3lq/O9+LcUrEEnZh8uoKrtm1C2dpLeh5FhGz6KA3rurnVc7T6h5DHd81u2M2FQKKpzc6RdF6JQ
tG8g6i78YpivCUthNv9ziOZoD1z4qPFfbBvRoOWtj8zkfebZKc9oJ3Oj8RxsFF/bjciVEXEIy2aO
aH7WdkLqoWWHWZnBC1KKpZ6DgVWXwM2x8nRgs9/ok1eyuBsVbknqnqS/+qzDAZixkPu4qHpUhRon
WBc9yY14U7QiL0XFKtNjbre0AWMO89JhoWNfnknXp+uKqxUNLoVMTHvf7hdO5emcLSlJ/CwOXAjd
gEi2I79ybQPXf5sBTrcbBEO41c6/9esiL8IIehddTHCn/uTxRYBP5XvthW2028B4rvpQ9U3sVzta
u4DOzfWSl25ZHxMgd+cgxWq6tsP1LPGAjiR0IkAcAh/WMT1urBfBPZ4+4cHPMTlSZYxhLzHjcU4X
5qAtopJ0GbjC3HofkCFfjUPzAXZwuCzeZjNz9+1OVbolJu9ToP4Ec9r7TK/8QmKVgMtfVKrnNk6e
qAhRL5p5tEalMt543j/S8Yiw1r2WiHTrcK7qw5fmBMw021/SCYLrm1aEPqJWecmuo28VzOH/OApG
h9ztnFAyvw53Jxw5PXHhy9T/N5KlIKYyXvOZj7hCkBwCX7r6cUk/SJ2jOUyRcASyGtjxT6QC1bnz
dcCvmiEsr9qBqLtiSIAPuuS2rstlxolimi8FETQBNtmqvkuABCtcIvfxIthunVc9kQuBjT4m3DcL
Gcalggvlmp/3RvtjHm4Q8NDjvWiq1DYcahOReCECmgGpzd6O9g2msZvJ+tsSAdvvpUMbqqtQfpF2
47WD+CpPzT47kLL9xA+BKDaapp7tGZUoXHBgrJU7TBhL2J2Hq3+AAs+4Dqd/IoxTP1uFDum2J/JX
WB8LCAIW4/Khzb4OPgH03vLDDxh1OyCXVE6Dp08/nWf0pdFm87RorOuGRIXkyhUd8LnwMRQwkTPa
EkK+5RTRg6vHftqBY+BLV/5308C+CaGYkY3ESabn7hGqKlF8V4FmjbuYWp2RhvXgXwJzTgfPmi7Q
DruuO10pIcP2TP9Ek+JyZsy+U7gYRvisB1kA1JCB7rrGQJIbCw6C8DZzVjNHJFVlvMypKqbSGPOq
S6cQiAr5GEOO7e3+Bs3wY742yAnwHa1b+9VK6ARwjvVUOde0i8yG4M92U92DWxo2XdGt4j+Ts9ID
CYqdUi6p7QqX3zm84KKhcBVBM4k2xnTpkbQqMM4OrMHIu1iWM35DpOL3aPQdspmKrGFXq+Pcd7+R
XaFEs/fgr0zsFwsm2QOZg5nxvo4KSfjbVX+cgoPB11JsdRTdM2Oi/xYAqfbjKlJf/mReP/VXaRwJ
/ciC7j7xnBg9GRyQBWpPRTpa9vFG2RiQjnI1ux8alotP1VkPQAQgLzSidu74t/9wjT23iSH0h+Iy
uhz40p+FAyhFkGXiiEAC56/QSywbNNz0E4tKzbFfOef9kLhfAekO38FaPUfSu9EEN2MyDKAcCsG1
Vq6EG3YqQo2xt9/jho/62WzkDYB1Xc5kAtQtG2fIWxEfjnlhWanhPjfjlDjsnJoCCvEVZmZ/Xyzq
/xCkth0EUhcWpeh2NpaZ6ouuoImWDyAGU8g34eJBWC3H+v9xIwGQE0ILrGCgYRM3inY33MH00Nrh
RuwcBX/BG5NzUdux+TSrOX+V27/fWCKi46K0pSwpOI9RwKdd9fudTh7ltsuP2+pStjh9dNOoKCLj
oewNrudRoHyg+sU8nCjPT322N0R/dThtZHzucauhjG537K0DbRoQWMI4TcD2vWt/1uV7e+scl/K3
bWs4JqRDMFhGt5RWDY3agAwhf0JZjxAqFstGeUDRJVbsU3U0e1jJsErKFiwpFIoeqKHrw5nIzk0Z
u3Hdih+k2Ra1XljFcD32IXZdrj5EHIGbDZRVILcT54BNHCxCtkrMGFJYAJPdwziMk7D0GykNPMvX
6sp2sBMlKoLYVliAjReiv45H9vWhnD3xhx+uvu8y83FAYuGMcDv6zY/znttWKnxQGNMlTP7Ijdni
cGN+spjMfxMTVR4+InTjklBCme3fqgZgqLWGmczR7L8RD+XFZUShaBqKI7KdrvVCyToNaN0Z51uE
qFfBg1FT9mkGsoVhvGh21djKXl3fLB5W5lBzaI0nzjYlJswE673xJ9s3RogeD+ilfRNj1dj5RzzM
JpXC+URGtRc75rFBtoWiB30fRigERBzVUZ2SMibZheKE/oE/QJ6mQCPiYA04/3q0ocLTOCLw8UxR
95oZr9mKI66iLcyTutO8MruUSWGxgZj/vNR3k3QOH/Bn8hzcLa6Znkh0v/1JSgE0wtEjisk6F70j
gsRz5uEs/4h7HsFezWh3ZAUicjYkywXIYdOpr1Z6hJl7P+vKWeYa8e8m7i3oUUudhmSf+XvyZJRH
qAxmM0hyxhsh+zK2fGKiQSLve9mnILEARmNxSgoIMcWuAhbhq8wSrWtl5TFw8Vgs2qrhBVBujQV6
///D/fVjwAFi5O2RwBjRJ74HbWxfM8wjLVyjkCuyv8fVlIc+Bd3gIKQNPsOlOy9RmaBItisknKAG
mTyKTNm8I2RsWQm0sa+ELFKGWoxbl5WacBBcUmBMNRFIFl7fxqrq68OrVsgIVM3X1vE053bKJebx
EVTaAgpsNDaGMHpftIpK7dhJVtGypUedpiFAnCt/vX/i8CpC55AM3fbkxXI6sXtrJG1K4Ivp8y0I
ZYQn+eOb4xPo0qrvb8aS7n8A3Ln2nOy/5+Vfv9Lr0UhQ3IK/C2EX1QL/DluDBmO5lZUAvSl5+omJ
kh1cqj0fWCwV+Mxpd8sv/ebuLHx6hBno/WHqqMv+u2y8b57Srfg6EWyr5gOUtrkHvkQKL819PTH2
usT7ZUjSB4LLAAxrKjXV32YKHcVSPW9d/RFH7uYb5xGyKnJriq7Z4NTctym4RfGxxDW3ahK6HN7+
Cc3mhLn/HXaoMd7fX1hEA8ctOWnHYuFzNvyoPcD7QEFh0ssa3bRWKP6MYWC/JlRZs3UqWl3wKRvb
FPhQOcK2cb9WKeIAQk2CJbHCZS+zppGHHVbhmr+n1p5nhzOTLnm+vQFLQ5weGi0gKoXvDbR2sImY
WG2iiROBql/0GM+eUxi2dw91d8xbuRkkWdxWi33gg7E/gKygzDHBy47X/qCF/ZLFkTBVfNl8dTTR
wyZqYRGT0Kwp0U3laLcNjhfBBHzh2hQCpP75tQJEbFRQVqXztIknQT1u16G+402UakyByGCkLCgU
cfsmSPtI9+6PnjL0GFk04MFboEgy4Fw82CR95wUyTIalEmsgz1bLW4N/dt6naRHHuOUx8Cmn1/Xc
y3IK6KsfFUgVs0k/LZk44YFnDbNu/6+/t4sa4nvuC31LalijWZ3XXh/mBWvGQweIAkt7DefSHoSS
QXVSy7vZ5vHRzC5XOy8It2NtO860VcRZk9lr3Y7RII19r6O7SaFkz7d0BYwZYSpgdCGx9rhH6Eiw
ymQMx4VAspwPSWxQzXRO5RndW+4zxuU3RzZfCPVtIulKJUBYOhO5GDfggBVObohEfboM0/LUTO3a
yE74bV32OkZJ6QyFhl9MDXmhxI6GWeuYhKG149wxW6FrAulzGaSAzQ7v44vq1iRLCNVc6UM66jNL
7OPMRKbIMcTF8gvuTaio9t4avA7rRuRwsy6qKtPKvuQ5wMML9S2Bp5NR7/6/IHcz7tJVTHnFtjyJ
A+AazE3ODq7P6wwunnskLUVrQpvL09Ep9KJPxSxx+YSoO6UxiiFBYxTlO/C6BAlcQMDUj9uYVAZa
aatAiMXA0fgsy4k85dGg2gGtiynfkRD1nAf4dzKRwvYs55rTbhwXCMSML7ztsf8+98DrLXu3Adm3
hamOoGNoyzcZSR5e7sRAS7I3j9hb+ABJnL0s8sy24qj1geKauhpD/sxkPqXsbIid9AEPnEKQVWXA
xmfcK+2CJivI1kNND9Gfbm3sRwFc9hZbaoaZJEgGp0djkHzhJhmuAVMFrYN+HuEJlzbgms9SxYRC
6ZKsQoOUJriA54dtB2tD17ONGrQP8MwkroC9hesjT97cwBVXvNBCOxrmHqoPHmKCw3mvUuCbqWQ9
OLvQUBhBEP+AebhtFv6KoMWtTzY+wlVTuYPBwijLrOoDp6+sJOCVqPS9BNGtX5t06ufqoyXDJiPP
x4JsPVb6rZb4Zzscxu8sxaS/e6OVCPVjnn2olojwx3rKkIrRZEgBRijWXY2VIVHe9o4fvgWQhjiZ
5VivFvdmmd/tIprCFI6LLpBmK0OMeuFy+RhLpqlpDDmAb5q3MUhksX3awMoDJyEOaGlvceFaOW7Z
C0KmNQu0TIq+6I7kiN0R3d8ymqIuKdEXV/qME/pc8P9zQnes4sSr4Ll4T8HnlnT3KYsgebEDiYbK
sQP/0xG4sdHBad8cP3HjnImBdEk8wtfou5UFhNNXV9SybcNBuxExNdF8RXcDt3Nw/AV1gaTHIjkz
NK8DVzZH0ed9YZTwmyTTgR07p7Q3fWxMQIYmDc4ZCiaQ/UjEYOmxwwopE7l8N09rDcyxrzZKKbcz
TYjmxCvRrHqPa3gNfXwAIBYmFedr5/Xbr02gkefY5RgBr92c3it84vl1wCGk9FTMcXHTPdO5xX60
xg7wCk44INvV93eONNDqKfbeceTBKjhE16mBhUx/fRYCls+wbjfugDCTjvVC7ER65TqEyDrLuTBx
KDcoF+vGII4e50MXPu/64IEsiQ8pEtyOrwDSemIkQxWBJ6F2lefPDZNxZAmcFmedFS0hnkWRLhj0
Y7pkvpFY3qN5+FAA08UYsItprGnvA2a5abv0LrAqtf2gAKr9JaaGJXJym/sVJvGh0Nau6yqBW/RA
9EnxsS4QUDzhQrF/guZZ5O1iJyCy8aevTCxUhqacXTXfSyljVBkCIvKziBSCLvQEqNFNIYRZxQ8g
aMS1XpISHNf7mGxoT2RoPpIkMmc1bdBhsIU97VhaWBxVofMYJlgMRsj8WbwyIkoMq/ewbYaZtqFA
fZzqd1sKVGWr9IlxamLCa1oR9GQ6wIg14evFiejXZzZpWklys709Qe7NtX3Av2YWMvuHRLwMmazj
i1R/rQOxMmXqx1HrKPpJt7P+V8j2BlCJW30dMuOiCm5HydWpIWnVx6ETsmDPJpdbc7B48ZsJ94OA
72q1V5jqM6FKgno13T+l6Y7HlkW3JGB8UdNYivUBTiTUdGFyEQNqrPS2rBNrajQurPs2hV/FrwQx
4GnlDu/78MjHUgK+8QHN4Q1S6Mo7rm54aEd15xye1iS/at0xXCRJ9IUf/2tyRzgAQzlWPrCTcSzR
W3JDDBt4nejciB5lRsVw7W8P75fi9TBrAAX7Zgf8WYh+KEBeQoPMqHmVrN7zBoFABvWX74Rq8pBO
xQw5uxaBI5T+DVAlnT1fGr4o4Yp87DQaQBatwIUa9Ckbdt7KsQyrKm81GlV3zuKN3bcBzCVTst57
7io83znPiCJd8hudxTc1ezDTaegDE2wiN8LJL80iH5mZ0JTVOGZ0F+9pTYXT8rOErDDSCX6H5Nvy
qeTTXyiMJVE6Zvz2cKjJIQrSYkhvu3/qrxv8d+I6mazMD/bRdehLQwwuNp0/cPjq69jIxHpydd/B
+qIdEhYARnqP2X1UheYzD59t7EaXua9L4Uf2W8udrK4MRY3udzqZDOe9A//hkaz59mTzjmL1wRMi
MJEuzU5J+MBgu4Ky53Cv1dTy0Ir8OekxPZldC198mGPkb/fTleh0PqQRdoY81KQOTXXDHNlelylK
B4GcWeKio5C0vYm+G09bL5OQnviES7czBufZ04Kx0XYqiXE5jNLCaEZDJklkTANuX4pxC5+Vfjuv
e1YPKVGgZMuLU9W1uzddCX7W+F0z7NPj4l9wjJordlvO486s6LKGg3cID5FwmDF1VUSPpWMBqizt
RDrGIFL83fFdjhjGRPEcf/qXK1fnG7tx0ovwd7VIdqzAAUr4LOgKOtSNczXnlACm6V6LeEP2RBm0
CWE/EyTrmqIRcdNMJEGJx1xv6V0IDCJrIDdBYhwHYNHEiSJQQrPZKMRf0zrF5NmGLl1X5++INfSM
dhNIWLvnwEBolCJsKC+32mA2FHQISEJedfICjOX8OT1bf0+rCfrhNs7ISrKgu0E9lrmHDZCvX7GF
a1HVgGFmm7WfJC2qLA1H/8TSpARcL+O7BpsCGltpaPN+WmN9ggZz+3s1o/SadCuhhxj7BvuX4HGE
x/WebmEXFERHhcIDRfFDjlcyaR19/7Y6zPbiu2NB1r6Y6qXikCRWujbEC3yp8LWNNsSz/TYcISx/
rgOj7hBZ+hRljnP2aoy2yx6zP+ZZvKlKNYIZUavwIBv1aE4p/Y3zHCRHCDbUQqc6AhWawvj5ndQg
fwbtUE8uiK59RpirALBJrkrBrWpsWkjk2fB+sc4UVytxtuZobHMfWJSxmuznuAQVYIpIaOOeoJYs
CdKsRX6GTA8gEp7BRsm3DqYBwnJ90PXOeuluG6bfoFBjyJzprEC9SlECpV/FwI8NpLwIZIKIraOe
wTOZQI9J09+YLj/h1n2g36cVhNlfwl58tOKuZuquABRxYsYqqCz76XQXrEPDzRZ4bZ9lqWQveg9N
emUMdvBGEyBGYpSY5M2ZfFaPzpYSVrEXmukRzUE/fzaZIB7D+z1tZrv7QAJP65q+Klvgtn056uJ8
4LP69yRvDTA8P6nDZiqSOO9vK2Ap5ulQ2F9yo/kDXgu3G9Ih2SqdEz7dKwj0svRNa/Gdwo/XesZ4
YbRDfbr9KYmriTCncGuRfEyrlzJXCgaH4Z3O/DGzBqx7/OrpxJlfPjpABRQB8GgvMyTUtWvJTrWz
eTBtX0C+KB2FSGLuBkD7OvlKMZ2A5mbVBYLx0dbuEV1Dd67HaQOAsk9zVYC2gCXUyz+9cR/UmTkQ
i8pi9LFZ/PwGcMjExiHhPtn6d38G/+B5jus/ZFDPiHJf/pgqMyhiuP+0O6ndpGmXzah7Y1l2Zhmi
I9vt5hNukeNCJPgI9Yo9q746KCI+xUJwkCvI0QfVk4ZBUPMNEXM1S1HnUF4nMKv2waxqRXqBRqUf
tMHKqdEoRQhOHc57OV1sjhFL24d7L+QlggZOSwvpxSMhOPuf28t53yHpajskUBwPoZPgwJxFET/0
8VSLrBwWUmNafUxd2YQH5yZHHtl5iz+ILwyCtsn6/1HuV8mD+45nYQRGgHLxeHkDKeR/tlj7vfgs
ixgWdtgfsAY6DgvSWZmhl+ReFlQIqh5o032tEejSz43xOc9nAhW0Bcv0UobJIZekC1obDaY62/OX
4VVyE1HTU2x1J+zKCRhIPUUn9ec1t/3fQQomdVWxWUH6QYOUPnRnQmNuvhC/FW4/nkwQbM1hB4Vm
/L7OSKtcCkLdpNQl44jM5PkP4vPmYTKX7KKypbm2nktBX04kTed5mjsBKdLZxSaKrvJQY73poyxW
ZaVi9oNK2JHFtcCPQD5wfQWjxR0u6MROt8HkNs8TQu+6jDTGPsmgQ4il7F2ewELP82n5VvHEpvca
IRBaxUANiAD0g9NDlO4jBrcY+VjtmiooNca1lYBO89EvaOpyIbz4CTqneeJUX5osOn725SAogwO0
jaDZdfXwJkXHLl44wNxsnAWFDiPmWQJetPa4cBFBqeSIQAXuCAkwfuvgG0hEXKLI3/fbYO3xtIFb
xSmu/EJMpoYvMH2f2IwFJuNcxaMY7BUD8hlm6asaq8n/7ZOY8Y6A0D1Vh2L0J18bLNrdvujmpytk
HcXuRo8XR68uQz+Hxt22UeOp/LWEwWiaCR0hj2OQEsxEsJy186jx+lelGZRkfJbnegrOfXatMphe
AJDCkEzdo41/P49ghaqfwyOCP4onJXY8OvJwjaGGPDIwe2F94mzb9ym5aT0Igy2cOpf18pKzoZGL
Cip3gQzmqO+X4o1X9n1dc9OY5UAgLGketPm14goKI+7bgSCrONULItgcVHOB4PLfdS6A3TDmg8aX
298C6k90bmO2RCsXWr89dWWfr+r9I6EOydtUodtT3ZrIn6lqFnBuUmhtkBoRpMXF/TcU74jY1h68
wzYDE4B4lduX2SoUi9ZgELRDsofz+LD0Z24j5m2bV4Z0dGChe42ykpJcQDSvGkSeABgP/fJQBQij
vfZX2zEqLH6IFb7ffGJOH1/ZikySjj/8Lv29RTfEBmd7ztzJSNJaiqqPewvtXYCiQDeu8NXQBL2+
0x6BAkjr05CkejbrrD4bV0N4a/JU0yK4A3dY6td+k7249ql/Bw3yhAYFlb2wsn1Ba/Qy1Lsdrd7e
+t+6knhWc0mozPe3oO+ali0I/AHalq0RYI50pGQXKCxlalnQUiNX9925Iz0GbP6D8rvlxo46IcKT
neS3X8CfDTDfxAbnFpFz+5ImsjUq/JPfDLI0g4Hn5JqoAtYdIQ2nR9HPjATgL7a/09Ln2iwSM0LB
9TJZDDmBaQGgBwj4/zE7wf9fsrAy4NZ9VbT86Qx42VGnb8hmNS7UZnMwoSQMcFmFqI7W4+ylfnyn
cFTnYDaPTk7CMmxOAg/ArB7v7PeUKQt1OJS10WPY8ln2FzJBF0413DxyVOoeO661w81mDKEy1pNC
nyhlvP/x1L6YMuE8gScOKRRV9luFJplafB1rC1rAewylaRMyYrT3UbSnhPOBfDLEtzIXqz4QO1jS
GKyylcqQx/Bt676nXj/MtE3TDJ69yBG9vblxA/LhiMgF5nUxJng6v2S884xcmi+o3LUXXEcje3dJ
u+IO9rttWRrIqVIH6NmuWxJuqp187AdyUWlOHmTdZi5PBQc+DaqGXDWD6l+TQWWQkXqSUokO7u34
wFeRRnZiXPiEGxWEf5a5g8iZ+gjdpCbtycUdA7gnEXYjpq8OdXEz6imvBINKnJgpFGQGI7NPAKQn
7CXitW1bTJvi0sVfMYDu90XKHdU5/LcCpqcP8ORjfiWWnUP0Nn3dl0MZLg81HjHE8qj1XB2zrboM
eufnwy5STUZUb7RRuib09+KwXQ5EHctPAlmSvF75Wmz02xO+OXYai3nYYa0OB8F0AjKjp+F/TPqq
TG+Y2fbzSBH0rLE0rlG6cOM3PmKi2p0tv7bEloCI63c+bcdCJTD6qK97KVQ1SFgVinewpv5hVy1n
sixZjHg8wSUxq/fKb9QmQyA/naREwORJWN0Rx0O3jfk0+n25B2xwNcxwNbXiQVC32jzGp4go15Lc
kl5AHl7c02M37JoG0eB62rortAT0OcHLUseIsaRgI8tM+BBocfe+kUsoNjCzYYKIQMfbokUC2QFi
dITbwePINjlk68Y61rLftuh75202KgBkK1KD/piluFqFJLwTU2hMYl36W75IUdbX0284F1DIt3aZ
iK7mqGVjyR0FtZqK4Fq3zixHAQ8TOGsiYjFUPkI2jFk8iCVufktCr2UrZIXeOGGtgp+XiO3cTYI2
7oYoze6f6Eb4YZnuN88rw9XwgWHXOczETzBlZYWLqLHKmDWQxJ/mOJu3eWoGSVCFIwPQcYKrZPCV
PmXgLdRVm2JxEr3CEDr4poLFiGjMihRBSdDEr2UB24O3YXvBETwrPc2ERTwOQ6TVFhYeEtzUuSHx
4PcnXxxRvMU8j9eeIW5MkHzdP/uz73lprAioxFYtdy6osGbxF/CwvYmgwol5nz2vxRGcYp/Bn50W
SJkDfolgDo67LYFWsg0b9zh8ff/T+0HWOPBoyIC7GLKV1PuI8tslab9B4FYW7QcmhWWpN2bHwQPe
PxTowERoEPIQ1OIKnwZoCw4KLkW8nkW0WOLQtFqJ/mU8E5Tc4bhfD3dloANasaTob5MCH4iqeLpX
c98wPoNV9Tr8ZPDa2qlDkx57EB6X0T6sST8Cw8lndCFltIKcAgzibLCtQSUHAXfGR//mtAvo9kYm
ixhiy0hudWvXbM8jntre6ak0JGrImVbHsG55wWNXMup8DzVsB6NBpT2QxwVDUe8oxajG9vmqv0+L
6LphPfsyx2OxX30oiogNxm//fCPVDOGRmz8gXVvilXGHt8LiV4vxkqsiAbkcQH/yvpP/GI5hEXHO
0YtC/oyTbJA4Jckn5AD9Sx6vvKLZoPddLjR6VJCsXZVNOSBqC0VikRhiMEsE2ZEPKRYjuwq6/9bq
hfDkBB+jYGnWGPbHVsj/MVCybqO6wJ/B7V4vA2NRx7n0ef1n2vL1/AWUo6VvZjKHHKVO9YGiQ+5k
2LjspYMTNrN6ybLB2d3fHogRfEPZaDWP40uwiSsI5kGOUVnrIaFe9eNPSfRdE03gUIe3MRVcdPeQ
a079/bs8JwyoMpuXAY0lWV7I8G6MM4lxMXXRzs/FhdVL6k7XRyalmZELxaLCJmZ9iHC1O3QBN4jL
j+D0YEDRb4lft29+8a7aPsmQZdOiuw5mq8KN6e7rLIUWSnm+U3Rnmxq6EE/eeoFztDxpPf/0lhnP
9qMAl25N3mssPTfU2g3OmdI7EveRhGtaW4F9atWeH8cXTSOoy4SgrveVJ4UESdJj2+QkhRjbiAnf
z8cMKjlzeQ9Et6WqyFWoMRr6YjeIO13wWBWeN3kSr0ea82gobE/Kc/nv1ciHFiHh/hc0CfSY+vBa
3c17woAf++b2F6+XAjgAxd67wvoDjKZgDUYE1+GmsaP88xDgyDx64lVN8ktzpLfJecet3RWs4KYi
W/gW/MjH9qrHEgDoRPGrOjfMuyMGiLGPxhnpBwf9SfdRNGy2KbMmaoeZO2MPfJcUNASU6vtBzU+j
mOsCiwwD/QuS6h4L+Ll4j6xXuhQxvjVQEHuzQMKxGqya2yoJSSIZAwRSQsycSibiHzUy0yuWgfgm
Qu3E+k8NZTanJHyUtphu3roIBRJkwZUx3gLTk+rRXjqhRZJkwvXkc4Y7bDcGMW4tUxva8m85vIIk
fmu9HilxsbBdYaACIzrdqlMpDE2pnnajkEY1u2ORaahgi1Mn0nxdQU50rAsMEY18ReeUYu4iesG+
p5EYw7BTxSu7a/MLg/CmrTa4bdG4f//tH4ZIf4giIVIZup5nNST7qb3ltkeJXKM1BLF38a3i2Mlm
DM+pOHb2Hmc9hS7wwJdOFWWzN7XZTVkncSXm6tjiADDtcuUwS1W7DeGoI8dIxwWuAFOYppX0COqi
KUDaFbCLx2rOwGDcDy27Dmjy45FGiRo4XE32lytK/Kd6tkr5cWgiJ1s7OtHFd/AB6rfB5lgoiaqR
kOIa4EljsKsZzxDYhXblDO0sJLQFxm3DoduP2feHlko9sULtS/pU1KzcZDY8lGnT30YGV3nHxkIP
Qvse7U6lziMDiCyVv5jzl97nOHBJWu0pTsLsba5McYhu+9TeDkJ0GniEov96DYNQTAjp/vkpVS4L
dtXnPgX/SG1zpO3hXQ019Ak59eUBL1FaO9o+1KSZamjMEZr8hVBRotytrQRmlcT/rQqLQI5LMAdl
az7ItT5AwiXEw9Kvf4H9TFHgEwGxX4hnvIxe2cH9xLUrTxTW69UV1JASSnJ0fY8L8V6doobBWkJc
zAAn8am/GKi9GSCpat8DlMIpQ/470h7ac99++eYeCxrVVO8ESTcpw/BWerRcIw7XAX7UYeoWgZpE
nUipYuu+pco40910jBBLofRk9c6nB7r2jrgKKkoN2cEJbpV3ZPj2/S3ZewZpMjUnj+xthvFd5ODi
pHzEgWC1YVbbVcMqeWlgvrlqfBwjESWitSeT2Bwnu11j5C2QFODTgNkBvPFM0GZ3jwrGTuyWHoJN
8jvX6HgWgw1a0YBpZ3RkpFquHFgTtANg2NRJzZsMG9HAt3zL93bmvUBWGE9nm9RFs9TzsixgRu+c
nHBPe6RVKVllIzXN087e3u2NttLFeJ4aJ1jY64nbq2+3z70aekBXLx7mQyz501+zjXllOK5+VFp4
F1Pd6hvwbKiDLbA9JyLfAvZ271E1Z8wW6y42swy3ikJpJ6AxDK2uCilBueQBt57nvKSravzF60lo
OvU36ALNMO2KXgjRTbGDDBG0uxAETRtksh4iRyBBEBluGd4F1xKIv/Mq3z7fbVk8SILB0lC2r0L+
vBskKjx8p8m4s9W+s04UsYRUV+4PDzaez1O4lXsAaD9J/f/YGz8tBmpRiE7mQET1NzzdYsNmBgvv
gt74+bVk505LRi+Joh26VEpOK8AIwtihKC+GAYhdmVuIGg4a2h64piBFmWAgapKYHcttWadOn8aE
pEwnua8genrgzOz52mz2uhO5O3ADQCi1NvTl4acrAzeVG+KNBynrI/fv8qgnRnEA8+FX+UYl17t4
XnvaKI4YRvUkkw/VaA4MV0kWMHL5EhQzKJkGPo+9snLmT45YDZbnYtqkkNLuk8NTBrQLcY6JD2wU
IO731iUXnkPQwfJaVHGCfvddgIe3l4JGJ+I/K+lQ0VreMK1SpZptnFRvITlx/wPWPLdZr8G79rhq
qQkJkfh2qYbacOyyyvBxCOSvvCX+WfzRzLzNaR1o3TSn2Q67nks3nEw2MAbDa25Yh99PIamLr+DF
QgI/0xiOJuQLJUUeUpg/P6rD4s0bFUq1EaAk1ObGe0cGHZHaWh5Wd203cslxD5I2n8UOAh4rXvUG
9psHPNwZJdqVulRXRhGhCkNHHRP7QSuES4Yzmx1Qk2Q+jVfm6akfgXlNQ63pmVA3ptpLE5EQdsT3
MLbS8Ae52Ionun/or9Wm3Q/ZndJ0zTaQx+pT/106Ygcsw4qoiLSXn6/kaPzoG7GRxeZ+Weo4wrUk
mfCmOQ0+rmemnJWTULTmXcTCSS8mj0lC/JaRmJMNZi+ZZpkj6RIrue4D+9w2kH871+wtYK+/zAXl
+t0lZCZxrkU8CXFHgcb47w6DKPensvCPaNTmR84R6VXkTeppmTBfRTTdACZEHG6bO/OU/IVHHDjr
MLBU2s3VmGbispj+K1A8FAcWcetFuXP7rE5S3a9yhsjgJdZ3oDWGKgxy0S5WRKlfb/0QLeksSFXh
9nfUz6dAzF0DQjEruGk8Ugg+vJsl/7EAtJfCk1oR+6hszbF5p4Tzw3x6wV5X5v+xnDuQANZCs07S
bnvwdcJ1xn+Y0WhfkEPkNFsFNjvx7T0qJsgS8aXH2Oe5+hfWWU9HhpFUzigNcjNrjpBIx6E9CDgG
lxIvGMTMTCLqJ69A5BkZLxXiLrZGBA+gWAvRmYpX3h/sfphMjYKZPPV8kHY4+Gbxn9lNTsQgQC/4
rXP1N/gRBqrYUTrOHoCsFnIJHjWvTiJcBpNXqcCW6u3Mwp7JpWwOhxnBxKbm7a8mpS+pnVyMF1jx
RF+zaMeSrAjuZ18xK06jQ+HGvQWmPERUqmnCTWpYrUwZStnVeo0DI1ErQAGm18Y7ijOaDV+xPRNn
8td0snEOnERn8TRxjrrxKg1Dnzkfs6KE3eqIiST61JC8sHx4hlZaQ6KrXfRwkqNNcU+fI8n/DWa3
tz/a7eS8xUBfmNEWRJhzYwITRHJhNGn7NmAuH4SduPx/3UWj5XEMyLGEZ0oiX7YExY2S5O+xOuyA
ROzT9AzQrU1XQzkQREXVJTzysksZtJ78qAO4Sv351IvVg568kh9Wh6eFhHvQ+1BhJPf4oiD0wv4N
lEfLY10RUj/afB5em9GLYyMge4QZ0IHyr1btlLU4KzAkqAla9UkD0/9vu3IBtVXPx6xBC/EcPJCN
V3ru/sNoZ4pmSjTx6zh89bRuujle7nby0eplAtDI1O+BPVWP4EYSFDBbAij19MMNWGYTcXWXbyZ0
C7XlmZxMfCcdR1bg1hQKihHyKOi54gj64Ahpw07Rt5bRN+H3knxXPnlEyl+niJitltKs04y8lrx3
c/QgvUndIZeY93wpfeJ3Z+aZT4Hy9L+2itRrSMtARP2b6/sjYtBS9WK3J7A4YHqE0HFWxzmuS1lP
n6aqDdFOqvZoI23sci3nD3R/1TDJdPJxX+UxQ7jJWYYwngJa7o5C1066/BimX/df8HFlBRKRHrXJ
da/aCylQcsD2w6iMzxK1tmo2V9su7c4Ls0zOsd75sU+6rzjUbD8G/f4+BAM/e5LDONzlIKfdlLgz
sw4/BsINIJ4rjdmTUKWvsElDUBxl45GhzagPDLiMB9iKy+i40x9epVzJnfZI3/+YDId9G+seOe4i
/gamTWtWYZxQHC1vKRaPt7dWlUUD4BIQRW6/4+x8CQHUzhRm8OPRPWdkOvv+ba31cM0HuB/dGY/g
SgLbZ3whzeGtkWbEWSliHfHCup+/LLu4VoyprLR4tAH2ysfPI5VXJ5HiPyTPLol2VcRp/A4h8Ed7
RIxeuw4b7jW2pwz/xl7lt/enGLhqhKgUOEG7IjBQU/gAEBlD/TxDT/cB4lTdHpXtx6S/uCaK887e
xehC0VXXUf+koWhEJBFqMz4/APk+EgSRe5xyFew5p4lcoYM2bNDsulyQfgGvUcQhI3+2LN5OfqV8
EWGa+hShfeaU5uNdSe0azt/CuwCpX9Q5Ug89hTflqdActnZ5awotYiWVjHQklVgcuZDwrOM2oDF1
mL64W28oq5dSuVOermP/pouEJwukEdKVfUnbkNAGrcWsL0hFZuAhiVOr6zzxND4QdLzK/541PxB1
vLR4SEQwvf3NGFehzApJgI7RR6GBAtxEhIkvnoTF9NlNAgiAwnmw0koClIJtbXmmF3u5v91HOynm
dRgyFkBsOYpHkNHcs9sHDTDe2ZmvBxQSw2tjo+luzlirR+vO24+K83+RRKZ0l0pL4WxJFa6GT7Of
3QFvAQA5U2nHuedvqTtYDIgpNiJTjXvrbuOth/ckWol6nxJ6y2in5nLxRJrBZFFPrVBWbnL9A9Lt
mbQ8acHKUYZFBol+FG6Q+OinCWg48hTthOkm/blQEnohcruvVXJgMcmVxbP1Ihsojk4dUtWT8K8C
eb5ynUHabWb7XMaV593yM2Cd9/Ha8CZbf081ZSHO92WDP9LQDiFnjqGwrLZR1enQqdktzZTpJCHK
/CxRwhCfhnhDqJFW+HYsC7aLAAQLM5UklUB/m1l7DtVlMwK4gBcovuzAggIxkZiHxkxKIUuO9N/8
n83a42UziOG/PV0R4OvCgWYfd8xaM8XDEechIO210YWa1bN2vNGZEM11rLilSb9ckd4XmdMDPaCe
6rn2HdQ4ZdMrIBtp0TsYyrTANxx06khI9f2VBz21m0CaQcoWfM05cLs0zfGWL7RfJaLA39k7Mizs
5GIq5E5Jm3lQ2tvGCua2hS2JLp1g6aOCFEiYEj++5tqRec1mXQDw3DdEb9B8W2juP7ktnfo1UR6g
T1DsCO/usGre4yVMbjbAnTLDPcrDDqtW/aLXQ3Y74e6r4vPpG3AOeM9/vr8kzbxj1bG9w8JsiKQm
q9/uh+kUiQ50BXprTHVkPVlMTgQtGZBiuTZP0+cT9eeIERchKMoIopEbcrYQtrzwOUh0UOwOyPxy
ouumnl59QB/gAMs1Sc+W36oIvGMYuCv+uLOmerigIBh9txWVM0I4W7XW4adO8hH3fiPER/Megc73
I/xDkmSNplP0PvW18dSJ0oHtHFpiMAyn10SLLL0YKZ4dSF4sfpK2HPEWOPzARCV7Zu/78NA1Rzjo
GusJlBWXbP8qNs0oRb1BWO/dX9LzHLQcvw90FqlGdWMrlNSITXDbVW9v9FUr2Y0lOdPvT7Hnrx6G
CFsLLfBvps1Z/8H61uFiAibaLpG/YhbCe5GRD2Srm2q/6gGvHpxIo7K8PQr1M3lL8Il5XAmBmS+r
/q8Rw+xP3Zl1N+Jb9bWnYX3AaUUpm9wQ+F7JZ8Gv8EcnQFYgGmgTexRuQWojWvV2+0hfn5nMZ8Q1
oERfsY/36nQKe2iTBA+fXOT8DLmnhGha/7TNwjLafeSUwHcUhFt8uyHUWwc8GxV4/q8pfltlxivE
UE9PQNWLUIfBnf1UCz/P854bpVp/uNmeSMryXwUt7YDCaMbO7uNaD4verg4h2beAoeHwgvM7cyAp
is3DjrgLy74SFsBz/oUomtgFFE+XNdZYqdNqB6xpIvNnCBZgeSZFKDCrf2DtZBgQ1rhR74brrsO6
Rurl4G2j4mlYGCxXx+Lw/56/lRSYQef+v5XqDPturJO2vDXq/lrTJbaOkREorQgz1drBuqhQQGwv
5uChmpU56uTbfe14J5w5N94WlPdue+Xqdkpoq/YTsLVw2QSX8+uXDs70v1VDA/hDG1Nqinfd6/4j
e0n9cZ8Z9gZbC0eQLIVQxJO2jHfk5CcfcISn9alB8m0jORFG79MtLtaAOSvgZ6baV1cDwf2VmQ/8
FYkM08j0Z73PncWBPzqzY9a4AzIrwBsXeOSaC15Y7nuo3qOxfgQC7EYHThZTD2uLc7SMZNYWcqJ8
d6asZL9AtnwxTf6Y8NAi03AsOdA+INRD0ai9Yz1iyKWmpBa60JnB370ts0O3OmO36Zjyh+wQABZf
IrLe6Dq3ysnk1iDeXRbO0Nb+YOQFAQkAqpRbsmdOBq0E2ePApEBDQvGxLIBDTJnDUXIzmpiw3gih
broaZ+eBUEgRI5U/oZnj0IqJK75hKCampUD2bieiHa+M1KPi6ImhW4OZJl+iRZG/aN6Pb9EKRxXp
7yRYyIWCjjG30MDO4ufHl4GL3DKeTZ7WiIOKfi9krqYpY8Exzx/dpLcDErNqhLlFx7IRXLSdDFUq
TjE4bsU4jG2sE74DuRZEE+SIsz21EsCTx7IKHeES93X0didS6EhjlX10yfAFx/Hyt7L6+iCTFJKY
KcmDeFMjG/TJcQjflTJmdaNQgnFbtLyP8W89AGag2PDJo/Hzey8H+Hgxsp5AvN0b+qAFL08jXzMr
GwvUuwgJBBJminiczeKP+mTfmRe4h3up1DS1f4/5nV+7FWThniuPr3PGj8jKniS5s+YmVXNaEXyq
cFH3ExIGjNBVXFOy7IrzPs86J2Pnr9FcSQfJGxifCaMxaen7w/9yJsjqapPOIWLDPDaTRryXyshn
wF2CwY7f8TWfhzVeTze93PekJcQZakMx/9APRKcdQtW6WTJfAYL3AA/4bt26iNd9x7yrqKRBcuuU
/eG4uLKqOHJDdyVrjLzshzBRr7C1HSOiwRQQSHbC5ZRcQHoAgeVze04/E02ogqrjFiknCPnhQ94z
GAya27UO9imFgat6e9PiUcyMatCg20eHwThgNfZXd2vVV0e37hxz98JI/dys5UYtJZcfLOkpeqQb
prAjd1KGdJRguE2ztgqzND6oGgQtf7t/NWM+X6PXv/oIJN8nRD1tiblICl1iQw77SbDOg6ajeU0c
pwvjUN22iGadRhvHGqGJmzj5RnQYLZr4j5nmfhtXLRXUKdCcw/2vweEzOaN/gewFGKRbg4ApyKXW
pr++HgHvRiNABl1KaX66QuEGWGAhtaawIBoomPt5DClXfNmxbKgEayKqSdIJ5TO5STzmivutKXw2
LfkOXo2Ts8pz4or1BrxRXpb5Y3bjUQ0J5B/2bingJRurLjjSmOzcLjD5dS0tD0weMRIIcPVuVtzv
st+zWPNA9thaEVEP3RQziWOYoA92NVF5nmuyyPcvnOrEMXqYHk35zZyifgwCUjd6CHspDUXNhaAc
+MG+z+YW68jglPNKCyCimOoPq9BL1im4QYXnpBpIAmeV0r+N7hH6QnJWBzbSSnVWpbDsVPjJV0KW
Gqm43kbQ6mah3EeB711ezVa9InwTGYqnoH4E3L0K8lV0kwIo9AGMdhJFnywiiHRwGLXLgPBn4luF
cFq6UVP/0uGkrY/GZ85Ms2UPRvxucOzkzpyqGOckYK2C91b+FOoN0pel2Ngqq4++NqVTTGhlO+Jt
ywwSKRuxCHE5kyR3pjnT1DFzBNdgu1YvHdTS/JY7+eKcjFw6hKQIs/MSkSANqtr/EhNb9j1runA4
NdNx1LQG+ebYYpV231lGXluwcxH/0BGDiRS6ixaJz50islUWmJf74kI9xtnV42kO8Jfo0bOIOqEj
BPht7USBrFr/bTJkiS27goK7VDyyEDguGlFBWwm4SHSzdDOnbvTH3pK83UgUipqMeaHNSwIaMySj
xhrH2oCopyV8AdIHax0Bpims1KuQmfFjVtklazm/LtvkB+BTphFZYcGlki/QjHpKiL/tsAsdmWeI
avnj27ckH7yXE42Y9cgop2Tr9D1qQ5mPRn7cNDwIWZ9B8K6J4Ta8/S7jDO3Ajezu4FNdQDkGgSiC
VpcO08Y3WM8M1IxgSYSv+oHw46MOdzZDhciuRt9hL0K/XJ4Ivlki1063cq1ozEVRpzy5iUTLuYU4
iIwv0KabWkrZ53SaUcA3vifzRxCRIVXhqEmTJa0hEzTPntdsjMirSWbWkv/Yqw+5TUIkiP8VxYTa
uwppgERelnGcikYlGfJWHLns4TTmhJ9biU85Lcw/L4dnXo+GUAduHdNLDTIIQFec0SYVvK7yCSbx
6Vouo6CkHQLC1zsyxaVOpwLRE/xtqx5Pt/4w1MFFZ+ieQ8r78yK5tYDDUKaRhbHlU8BBoHaROS//
YQoUG3XhlebEx6VKqETsMAZyqOrMT55C2/HfY3zT8JLNZp2f815IEtAA63p2ChxOZkj4RQMAjPW2
EqBSRCw4P5zUcZoq6GmfiUvwYMNMgYI9YKammizGQmvqRgv7ExI24gs7onyA95uGwhdCIDojHDkr
QGN64m1szeTy6pUCN3TvYCVu0Ec3lc7tD3xLPvK8/l1GbWRgBU/dQqE8A8+RY+cpMcH2NHoE2m06
QYBQMHBmmZcbPFDialw76ZKMfYph/M6Ef5JnDjgnCBGJornoItRUGBdOT0qwQ7JyYBl9VzVGWc+p
57B2D7JSA2+S5ZyongVDhOqo+iQ+5nypl2c//E0FIXG8hbav7uS+JVsLKGVEH+w1fGdKd56mSs97
pYfBrmvIIGeoonbnA6RyZG/MjTegIxE06wWZzHxAXHiJ9SzW52UKGYuVB/HZS0k9p7k3JdzUR4u2
lg93Xzjz3ecd0z9mQiUStILCNXivIrBBDs8JdfD/4+lf5VDDyEyBnqEdkL0NyxbWj1P3lcPvlCbx
fS7j1TZnYaVcSnkZS6qWOuhvnWpO8t/miblZVOCsxWhAuarrcxQ4blBy+4/ODud6vQ6CfWC4ILgs
BCCfYS4qp4hvC7xD/STUAcE1yEsSEIspbx95+UXZfBt59YjKzw50YE6XMcFxeOTezFy8XZ7WqJaG
L6BgAelnr7ftWy7GwkENms7hIwy+iLsS310k/el/UaRHJlQCsxj1ANj8691hJKtOo+DyFvMQlDa1
TYXGkYe+A5gE2KoB8VCjXK4Z2TkKRwKXVxdw6F59CYtFmbtsVdGeXdG4lbpqDUdZgblvw9HPfUhD
VS8K7bFB+UyBWOJ+1folOEYYmSXsEqSTQG+YTQVh70Gw7SzAxYpbpkO8W9eRo0GzzKi7dzaTpFFi
Quj7xDRYYpwhUQ90whBFFbz/xzn61/1drthUK0tkcR3K+1dUBroScjbDv9pUvDh3j9aIsFu6MxIV
fj3SSIo4zi/I8uxePICA0Gn5CLznMtnO8mKvlu1MmFaW0bX6PrWgvxeDeGwvOMrEOCjaq8WhUFHA
7esiNUvLb0cKN0RYLKQWMTvJSHKkPgbckgyrulyPNx6YO5S3kEDwIVyhf2fu8RzR+M54wse4OFmv
uTrDBPjZ7vRHYaaZDP7mq2Yn75bAh70ZxggfiEtKuc9sz0/OsLs9wrc0+aV5cIRUq3xIhyRQrx/Y
0gBsX9DVPwBpgfBAGjYGpoBfoaBDgqJjir431f7GqMmxPd9WjuX8CRmSJTy1lHYR3bBWU2d/p/qa
Qo38VZLkaYy4uE7cBM7JAYvkSZC4Gm84R1imgTLyeoApcdd3tLVNHwx3NIOk5LtjGZotMXg7ZzMh
fe2PBFc6IXpQMKFag273JcHcGpYAd2BRrY+IS9EJLoiF++FXdi3dF+bK+1dKMot11iAFNIju5svc
5ttUL1trBAJeeG9AXW/1G8wdo3c/MkEPDoceyJ4Ddai5lrHGAZLSuu0MpCxcATPyxxxfBbxEahDc
UJxSUtKWeQ9JSTuKhmC0TWpnnu+B7SyTS7Neh3u7z7gYtIEDbEUZ7P5W6gaRr38v5p4z79miqwTQ
Z7oUJfsSwTmXzYg6Czfbnw9ITYnr9AIJqHCgsFulFQthAG6MFfZ0Nd53SYZuT1eaWIHjfP2MXx4h
FPbAIRsGfDEGvJQIBRj1bAOGkRJ80ERSGDMEi7U9heXTlPWszISTjW1PgfWfY/yxhdZuyUDN3pyF
8ehehhiBufLZS+4cbGF0GNUibeaqR7TmZYo6TlRzRWo8HkosWX3dFWzDSP2khAcV/IGIuRgIstvR
xC3uNBQeqWXUT6fjSrKJ4rhHPVsJTydUiznH6ALCdCKEWcoV8xdbO+DypHIZ4OJLJrbqjn8fvnxB
jCEU4a6VlHa7ItH5bCDiWhxZUOVr9GIWK02TdosHYgzYQjlyZzfNlYtuW4RSwdlMcpb9PIXwgdyI
ELUbehKeaLLnVonCVDbKapdLKo/1Dx+MPnlNOeJGnH5c5ySvBkTfXJpBb+7j/QOb1N4CH64x114v
jR51IKHi7McTYXR3luBCHmIkVrw0Buu2M7SAmISTFpVPpCPK5mEDGs+r/2mKyxmgGxicdVso+r6J
4GsVTd4cHEDZRkSfxowZERACF2YnPloLx/qXgGqbvNaDAcWPcKx43T+rEIwfdpPq2nSInFep+gkl
WNgDpT4zQFk9nNl5nQqQKYSU96YWLObaHbHFiKaR+m8UNawmxCSPOodHx+OjWfjV0cBI5L49Q0Py
S9ghnNntVeNo45Nka23hIEVbppr6DGXamx232RXpmENqdtFgYf2gKGsVCnYkwfzPXZ3zAtDM9Jt5
pkvtOFLm/gNeC+ixR+bLy50222HaxeGogZKc5uvyk8u/YI1Ejy9tmF5YlWRZktUN8noxQ7qOnB3B
OY4OzmxH5CFcrY2uiXvez4xojeyQXkDenttkUwMfEwJDgKtvq5k2iH2huz1PXIBKVPahKYfm35Gx
xXluyUVyntIwyacV8uiU7m5LTLY42VvAUSvg4LT24erJ4e9vn11hwc7Ztt4NCGb8nrhX4fF/H2je
lMN5WpxUOKhvEYjsXjwklZ6Xc/vHtY4oU935TGdnigOjW4O9V7acVtrP13yL05/vvkJpnYNsJJTE
KgaEP481odC+zPLl8TTQdsDMMetkf5t7p8dQN6+7nhc8US6XwHZixtD1ZeaVHWqLtGnfiW2fa4pa
i1uFmHhZVVhGMUJ/D+0bTaDY4OxHaofK8eZTEjhPOa7609lm3EBlDcjM4M6DH3tuib7uBC6ffZXb
NG7FY0Vb9ei0ETVXRtjRo2gmmmkGdcZNRAfdAsRjbiUY2GB0srxBRqlTqk6dwcWfYCh6rPchN2FM
EShXRijKoVbFl/y2ud9h7ShoYCSgjrW6mTdobkRDZZOCcG4ih9CfeV/R7wH8HqxipDsZ0kQJ58Da
iOirQTkTCpg8UPH4mcYZNEv7tdV2IgqTgilocbn6204/UOrJD7bJrrVESTlNXRmBg/DjydWL0pyJ
y0o1wy6dTIgg0gq0y9W82BEhguKisPPvEka1zdNWbapWMC1WFKTn2eujefjWMuCxhvfmk10C2x3M
04IFbh2NzKswyofx37/3M2lHCYtOseX0ApdvanN+j0ZhWTrCTwINw6medioP5TukJSrV2XUURY+O
fvs+xVCNvYN5n6rvlpoL9iwZhN9NxwMEl+36zpjYH8jlN28afSK8oSkuVfrPc1ByWWU33zVD4L7c
qqjpm9uoUvrw4eANLanyjqOt+OfWNM6fA4CQiaWDnECfL27064MYRZ9Fky7JhMkaFanWqcofqJND
ubYalC/9rD0MANngBHh0v1aUsqwJ3SfVW3jUBA9MvSCKHLverh3+rzXmb9VgvuCcgI/3BLQLJZ4J
GsBP5xovW4xJZI2pbyohQ0eh/Cw74LHsnmN0A/WdBZLvzqyq75QAuRYv2dfHdfgDpiwDz5wXsJca
lJu1E3JlKsYDLfckMBQYrJ0baeAhCzhzcEZt461Dy9QYpdzLXRq2AgsrtkpmZHqpPQ+VPbMHkki9
FQ/+0IXky3Us9zDEGMy5rAVmgvV+eZxPshagTvJq4VL7XdRMHS/wFaBPYCHDsv/UTsMnPtniava8
tauGVkcsa2jmY5wDtjWigggjoSgweJ6DxYavTuyRC1zdJ8Kf73y51lPmri9SInS4FKVmMz2pVtLm
UDNGY5IMRhskeZNbB2rwuhrYqqqmq6Y95EdRASMMV983N9vfx0tjNM6HhytArEnxdTIa71RGfkWq
2L2B/9jatvWtYgNNOdn4rjjgAgdAVeUt//DBMDLeqt/GI5d1T7SQI90VpUsxtAaGgVHKVHBdN9GL
j42A5pG1lwKuoxBWxAXlYLQ2LARmcOh9ommA187EKhXX2bKHVPLhiMRLfV5yuAPcwaOJ0V0K+ydN
+a6XJbYWcK+jrOlueVVa1mJ7MXiO4AS2/VQ+4p1xNVYWDFOCa3xGQEWQxZDVjqz8/0jyBz6KlmLD
rAxJ2gplkZ+XcHhFOI6U8wOL+t/2NuM/ZrPFyGITfNQydpUgh26ImQHSQdhPvxmHT8bTeD64Ae+L
YcbZc1LgQp0ju1/K1+8U9htyzKUJI6MiSE4zH84PtsPHJAUXARkvojTUbaAPcAliUCH2WtNuiyqw
3a7BML7ykQKqEP8//uYIQBHGcnqA6JXDKlP7zt1YSpiO6GG7hbCpMMQMF9idmF47MHGPZnuc70h2
pqm97sx3YDQvwGZSZjhBJEVMAP7J14E3peHq6Vx+4Qx/JXErIeA49QCB2IDAl8pOzE1Q24Zon+Gh
iD1zwPwwOFOfTAsJNBzQn8KUfn3eySOviYfJQoQgkdDb9lwzLT9hHZlLUZQOoTE74nCEq9/DjEfw
DxGiXSfAYZl/Z61vkTYJOkGhF2d4fidj5RUkxER81LDTzCHhOE9d6YNBf8LERa/fB1vTxO0Du+BS
8WY2MnsQL1YwFUVsvJhsGbh39RkfVDMrCu0MrMC0C8nj9xcfKNdXKZbDmJ6+pYl0no7sBEBjY04V
NS8z/jBhA+ygVCgzasUk66BBX3q08+yfM1gH69pQjV2q1HtrSvTEE58lhoQvsG+7Tq9zlu9dQPv/
z5/33+cJ0w0HlXJlqsqls7FknF0AUhnlY0VcaNiNqGASkXvmEw4NmEj2oVqH/9vwEbqGQfk/KL+6
l2MV9spD+v96KVv/iQOWDdK0NU9oUozn98IyQd0MXWMUs3+7W5IkwZIbU2EXxFVmvSSg4NAQ1xby
Tf5eQWFNqZX4kQA7VYOJhuxtrwpM6p0xxgndgu+qOCmhblPOu+ZJMncFGRlGQH5W8X9DuvojAIcu
b0AT6kDsHg9PBs0PjZiZEVl+VYjB4y89RBFL0Ppc0aceiYYGWzwUt/umqXridfpukEuWFm7m6TcZ
W7fwlMtBDqGf85t77eV9uz0tH61Bu8P3iivmayvXfc3uyqvzJ9n9akc2H7W5kLXjXeQqOQ7YIFVz
C2GnnVeix6OtmICw6FJ4ikHsXGOc4CnzxjwpKnb+tb9QXLwzvh0TTUuDuze79PecImRXll++5lPp
dmfvmKmIwzN10A2Z8Icgil44oObg0oQHMBdw7MYChDvFuuzvb076m6yM7oo8wAZaFRr6ZXxdgF/k
N/jdOK6Y68u8K6TON0/BLWKD40snJLrIGDBbMouN2GWdd220vzL3/otU3r1TRgXMgFVzglFLhX0T
NsbhtM6pdaHHpktdAMoA2O3/rqGgBaGdLfB9oA5sE6vRn+iUDAPA4qHObDE+bWVuY0/Fn15ktmHR
VddMpLuHIE+uoj9Qr1e9df+1Wwrck7yvypREJvxLwJi+7PUiU0Nl1MC3hRBV1g3XBAgR5KMDxkEW
hP0Xc7YZl87JIxxBmxyfjEAbzhEAxAJ944MhpPIFOCPHTbPQ5U/coGY40+NJCACPKXYe/4WTDe9h
3raln7i/wPboFpIa0XPWQajL7mYIEIJNngZCKnZ1zTf7Yb4DmOsE69NO8va+xcDD8s3K1L56fCGR
7wx4YJPyeLF349dzAG77zZZslQkTFuhmYf5egzWNFVolNyG6vHqDbE3LncHwSlD4cKaHzoNsKney
UCopvJp69MGdX1yceyMWwYTDGdBIpsJ4lnhPr45dZyVYRG8uNAxOi9cbWJobjfcfsJrt49CjEI7w
4SuYQ5EeWtFdlxemV8unbPIqYS2T29SshQaKm5rDcUYopYb0qYl6/ulpCnBxUm9FzUKYnXTGqnVR
lc5VrqcGoLNYCbdIVa1G3eItgjIikDSDvyAIB70fTXrwwYE4pn5usPFntyzEl2nXfOs1uiQwfCio
cWzfjIzqgRDevf1Uz/y2jkGYWjVtysoAsQ16/Jm/9sqM20XZ1e8g8uNDJk+9WR5uvUfTDMLibo5Q
dJr88WcEVtYKj0sdL1qwCK+DI//DvXjsvvM7uuptYrl+QacuHP2UgtQC58lLLfam9yc7s4ky4r7u
/q+1AVeQ0CFAXbUYNyGORjFsFYreypKje44uUiidHGRA24Ypw1gWCcuMqi8DkwnOt73yulCwihix
wdCrHA8U3N4U4I2BWoaFx4/THYY/PJXOJJBlSIQUiYE+rdO/FlCUAFQ6A/SsACnp5EQSeffoEDiM
hjxLTaHsEJs3kW8U32B/4o9QTm2f01l2BIWWZdpc+PdCeY5M1cKZc8hSW8A6olDIN8/h6G8j1OdS
+/cNTbYkmsMMEfZ6YjIe9boyEPt+r+HxGi/oBXfg3KHplrfvB5mLP6lOH8ELyQNns5LiEJHX8KmA
yRVN0up2wt8TydyHTpd13UNMtcMi76TrqWuys04i2v0l+lIeYvn9SUgCZG8xXwUultoAg4bQJy09
5E923D2BUdRcUjvDHmE2l0SGMRQa8o9ZX3xuyDPZ1ZgRj4R38DydqWrm2jtwnugAomhYMlNZDoJJ
yR/9YDZ6oECTfZVMeIH3uhdmIhzmqH1xnutepIWb3+DlG8I6ii33qSgkduQpm2KTL5Oa7uicu9Zh
k4dIhQ81KOc84XrfIyxihe/nwO7La/xia9wl4Bz3iwbrLyWyE93bTEa2MvbvkLV9uaQDe//Wis1P
qEhhNQ9f0OInL5qasKr1FphPTAdIR3JlD6YuObYS8pMGTcsZp3EltgnxfeM/+gMmNJvlkH84t+8E
fhd5bIusJfXZpktz6o1nWqJzS07ZWvdVYMqZsV75dWlfbPcqqefuJH8BNCGkZoyi47VOSYP93wGI
uyugn/XTEELUjvorsH2+vgVRqaD8Nifu0Pyj6XMNjLdMC2JFeAd9ag5jSt2SFLT1LY+EZ2hZHYf6
UJcufcvEt+pmocPvCv3H9a/t63ItS9CAYCp3cJHMv9AwFOFheoZ6XECMEbbjPFqFblxm/sZqyTcv
QOVIC9pLrjFbUL0iLBaabQFSwkKUaKG6sk3M0Cz722Ox2qQduo+sOdj1KQZG2V/BpNQo2RYhAYuD
4QsTAEodNWjV5wKbZpTgIyHixJ8Vi1MdHeGZGCd3vfts34APa13EMmjx97j809z3e2LMFpaS6hpp
1ypZnj3gYhlSqzpKcTbt3MMB6sexhcBwq66gsemXPusR+jg+3hJx0ws8D7/0RbwqlglJPWdHscG2
4p4gZHEN+xZGS/48urwPDZIDuon4QEzl6SQTSfKXq4K7FjoiTDija5+1CFtoQ/9WL5SnIGPUZvO3
05UgG0FTPa70XwhneMIy+of6rLlLNY5x2VXXtAO2RkqrEAJBetKe+pxYPLYBQ1aipCF1iLHjlZpd
4dvCsj6mNYj2/jmViFZj9JjGFi2aCje50GUbn0pyG+e8WRgeN42AGPO7Yn31GQfJNypDjYLFHk0L
wDv0otm/MEMPHlbSW+OJoH+RTGdTWtykTpjyqXJ/E+oYNLBQ7eU/d7Sgf2/M59Vve9I9pflJADLk
vjNdKGXO7bbOiKG9/jmyG2sFipqB9Z+WPfIyzcbNB4/jlXSzGXUi+egEWoAaOz+8Oy2MjEw3jL5r
PNU8JHLCk5cY+E8A5KAPhVfZ4HOWaceD5UBZNL6z0WAt2gTtCjWpC9teSkDGwUgVDAuNe8zM+SJA
S+ghrEvRMBzINyZRnp/g7J8+WBsYJ5wvUqZNA4mZs+smywyHeT9orDnNCGeo72C1n69FvAHDIs6e
bzxv1C6gabBjVoamb62UhgZwG1nb25pUa6HU4utO2n313/QqcJhLWsSW8KkGjXJIe3TMJMBeM7oW
Kbwq2ilUC4Ryyj+yXKpyWC+/2rS1vyONIh/iZ6RtKxZF3104H0vcWe4CafYrdxFL6lRWzml4lqTG
VsWPkq7JPTsDD0JQquYKHPw8zGm0ACs/oQA+17r6IdklfaJG6iWQK/VcOkSareZ56sfE1DpBmLfJ
PED5zwghz3KalArbGPvY58ajEv53CGlUm4AElA45CzA55RmWL2plXV+n5oezhCWJ88jDbIo3f33t
Ik0c/8LhI2G8kJz9Pk1z3u3UIR+vgp4bEzaLQMgwCn5PfX3KssmtTp7lOCpIDhWxmCenQnWsW/DU
kGK6rmVsZt42xxxNDSfFpCdyxzLQPmt6C8SNhKU/vsczj600aW901OAvZqmQhcZRbYuKNGhNkCZE
yJlRL9eZ9lEQNaMQSAoxwHTRszlp1Sp+fnkYirFHoiQSU3LgAFy51PIO58hxRM4SsMsTIbL7GvlZ
tDwMayqtnirqZ5lmhvgC6qcTpvS63FCDTAacRHTL/DdImNBQr5WjGKNjIxV8zaJRjzl4Ha1lxilF
euUbwq007Hn/XdFgWuwCD53JZoEwFfQvn3La0jhGztBud7UCxXzrXlthCUa98KdseRNv2oiRBz40
q54lZU9wYBKukZpzM6ErPLJ9EduwYE31giRf+s/LkDIjuaV5F980aXSPAb6Ku0QSX30buTiYW9Wb
1M3zc9EhH60KZleO2wQEpYF7V70IK34tLbCB72G5ixowWG05Eeoy3zvxZhEarPUNab+GpDcS11OC
U9pcItflqdSRQ999GNS0lZkAtyktGIFIqBxdzIBD1MKo7HFRwxKtbmGD/6RVuNHkrHDYJX+Gy65Q
lRsyL5FwMS6jrr2G3lCyFy1QvXRoOZuruj3+1CgxSGVl3MfF2+WGCIsp0PmFP5ovvX7Jp+SOZ7iU
UNsA+QMdccpbhmskuxJ7mlbC0I9eHDMiatdaQa86K9MjOYIAEj/4mYAWi7Cmsxr5GllEgIGmy9Nz
KguK55YWQ5fyvnnln+PTkpvQb5v6DdYKyLsgtqnR5V1TQBjasz/8/m5IF1odhPMKrG/p3GWsC6wM
l/gkYWcEZi9bXTLwYgboqfwfZ8QflkbTnj/Sr8TkY6UCLVWFO78jDnMHwrw8Gyjc6ns66qHHcTxl
RZbXT/jtU5uS8fehqxEci1JYpcz6ZaionEkzzuMfSPKgnKZlo8xlQX/hepQ/lhXvlIzfUQ2WQ1R6
pO63+Fq/dYi84Yz/n4FAnwLvNcrqLdQGQH7+Q8+0DjucjdwMOOevvyjuM+v0BXhx7BCAVqiPf217
2bLNpOF9Xne4dyeCIYm8yAIsm+9y8l8mqFNLCRWnbIjJCL3kOCgkC3vAbbevbiHRknEfPShK40eP
0z1Fqz74DoB31Nslmwh9Yd7zZHkn3koWgTDJoEG4r1ylhaQ5qNmFzaSVdumLmOFRa27vEZSNF5oG
05+rvLINdd+GhnCycUL6VbxwWt+bTMWRpj5SzJHrsgrPZqZjoysrWaADr+pYN4stfAdn7Nf5mr2h
EoQSO2dZEP++0mgYubvSaGlCZsQYbvL3e35fKOGbbMz1f3Fx45p4mkAdE+XN4ZrkJyFptcQTApRO
ckPDYJSuoqOg57xVkpHk8t5aNQ2M360ARk4Ku0jHuxiH08l5hHDJeLcFb5w6d4kxqqfAN7VvDT61
V2tFYGdpO3blCrQswmVBa9OkO0krHPB/BlVjQz5M9SQSg+O6MNSvrZwggc/MG5oSgV+cEFopL7iF
e5tdV2FdL+6aPUZlisybx2rRuBCuMMJF3GUSTzygPRhZFkbxY01JRG6xf7oSNkUDAERYhWnOWrjD
nCBkUCG33fgmNfJMjhVcd4fHpwtfgBRhD3od35SRQAeHIVI88/kqK3L6+ok3rBDmSsFSxgFGyprc
yIykpUnci5wLdPXKuy90ygNsJDz3fFy5JZ3kZqpHmI2XSPMOd1bl6dNUtFJpus8bKrZgiwXZK5LN
2fTdkLjMrInK4fvRvX8eROPNOnW0hvxQIrWeV0CtUAW9yOb32/0353kAlkVicsubqwrgvNX8ISH/
KMASS/4mmzWnEYahHXR4VJUuaq7WbRsWZ63UImyjoI9LLemINBdKV6NVktFCTvKfgZuJxkQwFYGI
9d14y+8BlSnfoEJakwlgQSPWSHLs7e53QKNIULGePtd/2wcacyhi3L0dgAfmXs6Ew7v8x6zJBNts
rb9YA+9HHMGKhc3XOxr2S3dcSrj6P5GS58bBn7y+aLdVQPNRpa4RiLoUsp4ao7377tsHDce8PeVO
fLTBEHMzTHjo9sE8OnJRjZyY8pStRd9oZZrz7ecrP/YtQzkg1xhnz6NBLANC8WXsNR0cw4jxpI9Z
vi+jJTX/+GIEddyj+Ytpo9dgd4Q7PVsXkY1PvkIam6XMXmDLTs0bJWv10ppxjwVq/MkUx9dd4//K
SqGQLhlgzlfpjmW9CLCuIt0Cm62DAPUHjYCDCmubkr/7LW4KSye/CK9/7LcbrUBmwPT9Y/xICqzD
/pdTbx2ZH2dzJ5O94Bylzm3eC8qTG3X1MtNyGDlJ6e2a08FEEuIw0LbD0tarueuhSOM/BXQrCbv6
sctlgiDX0A/ruWREZwXzMWC4Dl1qxQuq4VRCZ+5gWfKPjttgtwpDnGzk/UNctdfOUSsDq2mMwN5s
gigZ8oTrCP0zYo6OhXPoQVjobyrCrr0SBwc1fCJUcEJaHv7fCQbBhyeGoRaHCpKOmTh4hByWrRh4
spxplgeOpkmRIvaT38sQc4Mxx2onme6gunBHqZ94dOr/PtgKwBAvkpLI9oFL0+tjn/QeuzfChvrf
urmxCK8V4lKW5fDPGIKz/qVL3alMT4r2fhZCMnFiE8+fYbfUa1WMsF/G4BbYkuaSDvH71eZG0kom
ZExI5RK0d/a+WoLC3mZunCBuP1znsYKIS+hvbPaAbt6mgW5ww9ZiXS2M5yPe4ZZIFlEqTir9Ken5
miOOHvWRt1MwLsxGXVotHT3ntjmMgPvfTzNSROiZ7QcaJeSdhkAMu3a5MuPk4FzYiD9XtUju6gCX
urmSYxDpgcNwpKMzuIHmxT4xg53ieS7QuC68iQF34LHSmkol6JsA2NnQWFkBZYOj/tbD2Bl/OYtW
kjBIU2a1r40GVwoPvYb+gL1SX2m0DbiZOcM2beNsgTPyIYrdgb7Lt8Vgqxw36dSlknIqf3kuVWw6
v4ZuuvKSlkcAPx7ti5ybuOnceC8TAqzFTu8ftWsJH5ChvKd7TmNOPdrK/S0z38yBgiV0Lkk0Hn77
anei97xFbmtxo05KlT8EuFPmjBemDTCAxbvGEGAJLXMA99DTUkCn0w4FPEw2JG/N4WhVEQu/8bvI
VAIsvVnUVgTFZu8/nCp6OCmCHXvDNElwl7tq0ajA4Dr4EAsxhV+RZ0ZVT0Vj4dcjZyh7/19UnhAR
TikUetxWqxOnW059y7XPbt/RwUyciRnKFp3IUcIJvNoeoEVbLDnxuuI7/sGDEgNNPGykAIl+Rv8t
B9YWock0Oy8buGNZN9w24JlLAcS9wsJiM9vK+d5jpX5SOr2Qrs5Az23owuIKzu43+7TE46/YrWFd
1kWl1538vr90MmTMD7QPePLA+bOSqK/8MED9HFt0dCdE8R6E60HlDRg0ZJ4TYvpxn3IKzG275wOg
6IxOPat5HY60TdJzlbPtJNAnQ0TaDssRZLFSpsBEjV+raSJE8FXLUqpilCXaDfr/281Q+r2aS5jH
Kg/199xR0k8rQWl/Ewx5aLXeLnN+c8hiucAStPwa7xJ7XCkARY7FGrimP14uBH16X1FqaGG4rKe/
jXQeCRdoTDlSjL/8FYf+b2QEC/30Q5rTvshrrUuEzKBFHT3Takp2T6+tWU3GpkVDDnNRGXhaK2AY
prhXQnFnQ8vaae2Z26c0nsP6lp0SuqliC6FtpI1wvhdXL+1uIH2AhIl/0hkn3iDT9f9P56p1Vrec
wZOmtwk/fiK0w3v+VpBSx8yWTTd/UCO4aKA6zysgzxEh0Sy1pjhf0MgH3WweFQp/S1RW+jfjxvZM
IbMA+jOdOdsq7DKfiDCCAdwe3g/VGGdc6AaFsNufPvWehIOHfxDeYIRduu4FfVIKI9tcHTlTyrf6
tRKdC+oCK8jTrGlJrGD0z0629a+sx9de2S3EhoD+iaGvm0QZzPYrHmvLUQ5/Ca4rybfcFvAdpWWf
KiXx1u+YBdKfvFp3WZURuLoIJsIfiTB8wYoAf2ixkzs7I2ukzE/kOmonTYTEw/pIhvHGI+0qxnXa
FTPAedUtIBPZ+5HV2HTLtdO8RIUzIJb4RfYTKXofIJdlaFZPedR+KkO0dfOV9Mfk7fHBXsHTvUur
y3EDl6GB1gLsUeDfjFCn3yR2GFredKBLlUsg3zmsqB44+pJHvy3ooKNovhtKZ8mphV4xGsEzUeU5
FqJtYqnuCfZtAbAGzp1gNVcw6vpVBKL4iuzdq/TrO69ACISixmRx2Xcp8urAxud5erbEhH+iFIPe
jzRt+rNnijvbLwt5Dpr69km2UImBV1ET0E51FMXEvJATqYCGHlcwTcPVvbk1qKRpp36CdajNv1qt
1hbGV2VMI7QAgAN68E0CzvD5rd2Ixi7smFe1vsy3v1P1MSHKB/i+YOWscUwJsXQLsyT6pr4bEQdE
xOxMqMAjTb3iPKC7tO9K+cSp8bzwMc5Un22zfcGhw3DLXAVFtJzQgZd9RNYyJrBLKHFUC1mypoJJ
1TVVe271EFbUTJNlnsF5PQrvrJU5NfzwXsUEk8WcEaOkufAsb/KIg6qJOR/u6FpoXxIgGwpKrsKJ
elG3vcHADx7jirKtbK3KaO3BOD27XiwcZF9EODFse3Oreue4ZTUbmnNuChutH6MAYakJ87UoPwp1
y0Ag89u0rOMq/kOB5OY3HeEgdjN1SDg2q0HoeaFBz7glC3s46Y106yB0afH+tbktmeRzNfpfF8G2
NEpD5HtjrYC3093p1+D5kzkpQYGUjeHf2g7wiIMiQTQCtaYVeIavtK5Gffn16MOWj4rHKCfO3KZw
m8QluT/XfJAhSU5ICiNp19JsvZa6C51gIEO4q2pzRAqE6PZZv9NTW1DgSyuZiSOzSNK7XKFTTPYn
l+VK3Wod4QcAq4yd7wPCGLcjWDzp2e5KMiQRvlkOYEi94GPpGhu9xmXXtuTOE02270xGlzPj2AtD
eS3fMkYUfKt0br9tjMVC5O9gL9kadLz6K1yIJ9UH9pzKYBy8Zp0OsGxytOHHr9EtTggL+WPJ77Ch
kwSokgba1DT0xt7X/1u4oieM6gkeAmE8SZ4M5D+zVfBxKGSWbLxfYzGl+GopoDSXLk9+Jh1ZQq7G
Ss8vCV1Mxf+JktrXARnn45D66lslRAIwUhuD9t2hz8nxAHCAJVni1g1L1I3xl8xqSpw8Z6h+Jmbh
bvpl1UX/JHF3srsRr/cd/rrGiIvhnVRdN5/ch9kPdT4gcaQ5ZAI8voK/sP2QoZp4Bti324X09p5y
1sp2t45Wput8hyWppB+Bpq5UsMbJjpymAgYBfmdN3Uk4paoKFD4CJ6tuCZb+7gsKBSozTaUDjVZk
ULxTgQZ0aoX/FHR8fq3JqHN1H9R4h/9RLZqRZQDTaJRI7aoDQchEvtTOQ2hugmfoTog/il03aJ9t
DTc81MKYAJlKm7Vj5nYfLGYKzi+qlKK7kPpxJDW18CKP/zom2NkG381A3m9JdTLvNwbOllpfLD4s
pZY9ZoF/2jbN84gnrR/HM2XtqQst2MU9h36DGxqDMwXvHWV9i8bCRD2XoOQghy603DMrePhqDEJn
6IRNMliEjCvfCNW7IPpKONhRJKsryqIm3H5qGmMHs8JI7GZVjk7P96gtvOaYOaOWg1R4L/bGJb8q
h9aTa9+NWiS5WpNhbX/LlJbrANJ6ASR36WdLPsglCATXTTFfFpKlTFf8fFp0vbEiRi/tNr9hsBav
0/D5x+mxkl5NNIrjaHS4P8U+tHTLrS7AmxnWOS0n2FZsSl7albcTZxiHDEQeWWgRQvmfIC0tg5rf
9IkeOj0bizKA4Bujca56aVZjNVXXVc2uawr+9i0qGT+6/7azotaXzILZ1qlnYO1Yw88IzKJHW31M
94EpzhXHPt1VQNQ6JwxycCGXP3BfJtNRaRjhb7PHx7tTUOuMKvofcoI04kM87epaKxav978kjjV7
i6lpoFgoEIaODAsdOyDEuaw+iglr7OajgsV58mllyIfa2zdhMuL21hWaRQZ8we6SSbqTTPa7RkU+
3zp9cvIUK0tsCryYEpBff5WZ8qbFYBJHwrv6RpF7SPa438PUsZTLkIC5TXS0ztI8Ap7HNCDUO1vO
BFaZSVc9OUAPyWRZBrlWpIxEClfo0sra4LbW+7XURKI2JLExj2aJd4+w7Kd+DvLiUmbkwEMfV5hA
FG4vS7TekZ8Krhxw8QPjzYe0uvfOtA1BoPbx+nj+X8GfxIT/WdkyOHSQHPwmtD1XOwuMJrG61fsy
Mho9MVZb/PDqFuHEDl0kDT2euNGQtWqfrMbQc/lIIc9NRFoE/C1iqhU+FSkb/HWJy+lVOqzv3gAP
Sp8rfu6QzV4t+CY5rSnQoDYvf2c+Y9a1rXRP2Z0KtdTX14T4ZtT0cXdHg7ihk9Yv4H48uDQbLLtT
K9r7Kr20EYyV8QJVJ5JLO/gjfiziy5xYeITRpi/ouWyxBwR+iTz5K+5K7MoJEOqyl12d10MkkYWr
2f5PDjaW+IJHfPqvNTtIJe4czFKyirBEADA3GWxBi+l6t1zo62bx2Z3dI+D/UniZ6WZKqQ3xBB2n
UrdqKUwLz/gW2U74ZaTMunCcz2rf5gRnVsLeRby1iBHJyqtqpoDB6eMZJa5Qdyx6EJrnZyhVuUY5
7Ochcr9eCEDdP+dGPPr1ebp4nzjzjC8qGyk1C/ibPQkoZaHO3F3yrTnDe61zgJ2QdiOHSXxE5iHt
nkuEioSxMhp07QOfWW3uRObXJyk7Hs2+fLEFyGqid7PwkKAz/LOHwSXy/TNBmoOOeFRzsUvVkoB1
7OghvXqLEnS/RwX0EvmYi4G9N+5Y4A3IEKqGdJL9xk0gfyu2W4oFk99DCV+HicMdjX3DgViewrln
JB2PUBpEH7ozmLMNJHw9zw1y9kkKteP8enEaftdpi5ZiTEaM32mvdSfeY8wOxPUbYZquaDBQM+c7
oRRhrMSTXy2WaWVNy+oPjbrP4Efif+52G+eh4mr5Rp6dkEk/EFDMp1gXb1Xci1ZJ9t4YzF6/gms6
buwzR5YTSIyk8syBwNcNWMRUya3ryQvOySmTqQ/lVG+JWyeb4TE4wDU8D8KXWjlGd0kgnkXZ127j
Ww7GvEHYNzvCF3SRCk4NAzho7bTWOkQGaQ8xnxh+GsnicETlbBzBymCfpqYedy/0ibDPx5q8PNot
LeUoHLCIc5gd7ITqGxVYmOqAr41j4opzVrYsADeNvNEzITrWXPtPk8AKnL+B3RH2fZAE74STVAN5
v9n8g4OWZIPE4SrGLsEZlqxZ9NT/jEH8RPyts9BEP3nF2OmeIvR8KHB7uVE6bUa2QUx/wIiqe6lw
rzEhYaLjbr/qRsX2SylDV6LjKbgSR+sTDjFoiAgsgYzWio6Vd83te7AWAqeiDzdgFJmK3FoB9pF/
AcbeXq0xsCG/IwZ8DSmQfgJL4yfXIZW5oFTy1uXC4a6AlVt/sMEdJlY/3k264gmSzoI6ahYWYLYC
GntxH7nIHnZmVdc+0ZSjrgvZ82W+Ge2QVqrGvNYkYkiF98Z293lQqfW2sIJ0rKzT2S/8pzwZO1RN
R2lRQVDFdk+l6qroJgrc2sektcwg70TJam7CRW5rMWNJAnEAOqtORDAj2/zl5EH2v5MGatUrDO2c
85f2FmViUbGaiLiQnYVXj4n5TRCwtKCbCjNttw5BHfoDGGPL8t6qTBVyrYdAXRJ7lpDXsN421laz
5jREX/JcVBts9Ao4g2sauf7mkBv2vQF9eF95GuBRSh0cD0JVJ4964p2GFJbM889yw2jxeJKkTg5H
PNDDSyqm2rDrKsFV24KbPXRZcvRUtNZRRbEDbZ8fU6Tr6vlFjFKX18omaSyPhdz4HGO4/xofcbzP
ZEUczomxG9s4zrBH4801msWDl3n/t5XMNR9gch+nJCCbgkPdsGgndSWpoaipx5gJyFoyIcz/hONv
JshMkP47il2h2ARSZrW7J8TdkIW54ASVmB1RIe2XdpH8jX05XBWQ2Ij3e6/wU2+YDa0u7TMtYpvV
5DVghYWrcTmgpz3jvXVuI9QgpuTJ8Q029p1IJHYgwFJqIU+KoXeanYxIUV9Xu57O6uP5dkH52UlP
F3wbDYfBUSY/WIiY2BAbsgtNyjxAxbRI9SUe3CXB5V0eoPAC0GXiwQhLNf8Kx9vEqfM7eLlKmUEZ
h0SzcwddMTmEwqE0WmKIlxURoFxo+T2beQGPvJrdTunrHSqxmLE85bOWCcj2ErJSkVY0VWprj+U4
jBE7uAcFOZvQTVCcN52O2ffm+GJYIbQyLaZ5GoDoZrUjUxp3h09YU/lpfBp4R7p6UP3Hwld4cTqA
XW1QbVxFuvdwIEb20DKZuG6JnegMECOSBfxpQY/nGZwWzgYs/nwf46mZnz5KvX90qGFhzzJNp2Hu
JogaVZFajsGwvtBn7zpG7J34W9ZsXjJQgS5+xChQtwrL5nm/nSvGmfg5QRiWvhS7lYeR1N7gQQt3
7pipcMRVePe8LeafqR+x1jFDCWg0PTlEPWJBLnAD2Bv6iRbPQeFzGsfBrhDsZcp8pFwr7CTx2eYT
xSYhasIxAVIbI5umy/i90EWMZJ2ZoG3aWVbX++E3kCT00xeTqUwZCoQ/wCbI3cHDLEIfhpf28qoX
k8POblqoag88jQCXVnnVFkUSVW5KKu0DO8GEpxDcesyLb3glRmDRglidalh7ES7rpagWlm5sPZ9X
dHlVOpLLZYw5F9wE5BS2vLi4z7Prp5+ttxHStgwJ/VNVumelZIG3rz0asFiS9Y2rR4dulKc1M1RB
vOWWZNFWGSEfSOomzEhJ5u4Q1b9r5qyfwkH/9GCZlCSuFAq8IyHSuuP/P0Tty3w61Ugfp4E/gD3f
kQ+p+jHNDzYXk1IOiU6o2QrhH93KMGbhFIcSi3ZgBoqo+Xv5ckRhjEPU9bX6DwS4nG6e7rseZZa3
sGdyndtjQaehrYte5yCUccE0SOLWZBa88pl6rNaIdM96suAsL0nRwb+Smy79igBl85iNC1tRjztE
DgRBWsl/bnynb7bQ5oGCm+MwgCwmBrZ6qXUnfgVpZJOekSv45j8LYft1eMwY1JiPNjodHvf7TJhK
GmLLgphDs23Ikv9mfKh7YVrcOFJaXuA62NWmvkFkdYZCyeOGmoFLGY3z+NUqI5rJI5+6zFpPSJfA
3OhZAHdt8jLM72yxYgFV4plbRJGLji6lRsWzXpKMwjVAK/aJAQp+juY/Jb3SI0M7XKfJRFYP7Ms5
05ELdKeK0sfthXgTOcRn8gZiGzwagSE7RNBmOa/iD2bOxbFqQZv+JrJtfzHs7f7zT0yvjkUTSeL4
W014G3tjaoc7QRwu2fajV81eDiMMVAdHi/qMsDgH3FcE3BmfnqhunoLU+HdxS/hFxf1+fE+mj24Z
YrZK7ce8x23jHzRF+YPW7NHzyOBQ2PDoX7z0BCFjq1/XSBZfF8lWX0hQali5y7RwGT9xYIwojpwN
Uw5rbq61Iji9Tv5/2oZ5ocfDd56UGFTvmQesN9lbz+mBogpk4bth+0DuYDHPUcwM8xqroYWt1Ady
DwMfNEOECVmloiLvaNj/iS/7y14ZdvlnEJgldM3q7mPP7BqlKGYRp/iOZwYafBKqU+YYj/N4lauC
VWN8aYqRNgufOXVfurr46pIXeRMCAiXsKTH27eRbhkSX4YiV7999APCzoZ+btqR2Uvdggp8GjUnD
lX+hieA6u1N+H39NBF5sdQRFJ83fFlFyl4VE94Z1+JbE+ZTlXHf4Eb8dAaw1PhMItYB9CBU8fvOS
rGeL96Vb9twD9zpBwx+pLD/VoW3+qTvQhUl8enTlU97qxBkaICbJomi6oCWAK2WQdK8k425KvQ9F
fw9qUJCCxf1zZlw7yzE0bxljhnbE3Aj/at5sut4kxMLbEbYy7yOaWsCUnDR1pNhiq7msQHDSg9iX
El0mdcCPk+nWeKsHRTGc7H3gUuNBif9kKWc4lodwkg7CTa2uj/5X+YyGlSxJmmDr4PiF3xDDq5Xu
7PtLTQhYM50PQ4aQ9rjKc/C82ch7yRPHNoJLYFmYGtuwkuCXsXGsFiZCGzokxNrG4hUyHB83Ai5D
ffv99xEIIEXF2lbb7CDV2h+ePYqLs5tjH7rHxZzOPCZtPdHPHMT03tiko3LtYElwKbw8lMseTmon
PZ0O0FLnGHGmd3/+XNmqwWw6mG7A3Y7DSMZLR5K1BQv6DF0HefcwlJFJWadCvClIMacQQ48Q9fyg
x9sn7vftxHJWO40fpiM0WfsgzhiF6Ueh6WnURQb0o1TBkkfZ1/jPP+Vrm9cEZ0J6tRXxjMIhEs3F
KlH6lgyNzRRn2PIIvJKwXWVqowgMIjnU0ud00ujO4Xb1m6td7iDcjefa6BsZkjZNEpoPa3rEfbdA
VNj7a49+25ROhn7pIrBdtFwfp77TlCG0XG+/0HUiQsBj5WIw3VI0KWHVO56NOk9e394MMqO4t3re
EPe6e6cJ/m3nbwqwbZ3bWu7TtcrfFt2LboH5i6RV7gYtzdRd1xXYDv79nWHc2cviwbz/DAF5SiFF
AR1JcbKp8PC0bQIM9UY2HI4Ur8KvkcjNH2d5a7r71Y+j2KoREiCW4CGQM5sfFDyU60z4SHhRr/yA
IvPYRI5Roh/YOU1lCS/1WMAW0kPChyCNfZMKEeiQ6qrpyQcYxtXKEGfj+S72bJSir4mfxnEPzn7J
7ZdIEZ2NWrl3THCGvu5uVaa98M5E7QGpGDksX7DMkBpYRbY016D95dKAsXhEoBoTBlHS5HxYo9zN
GpM9ae/DqW4Vz8+aWiWtVlqfb1BOfYFDGRQGaZHB2cKwZ0fjD+5jeu5f2K14UTbcGl7IWnTCuRtm
tPYqpcnB183CZVOmWmhuhHIOGC6rMLJ/fgpUiyh30WEdz0lOaUiF6SxyCmUmr3680c5Sis1j3lHt
04KxB71PrlkdzcvMYNIzuSa/AZ1MT4wZL6rHC0GhZgv9r6zqxP5Q4RVsSfpU7LB6j+7XFU8y1S0K
to1TtpgK97qc4uQ+Okea1dIAdtEvP0D9S/3hs8ITHJoUwTXjYk4eLlB8KK6i/be2VJendfBw3YTV
cOl4ccX6BfTFAmXUU0poqNUKjhNxD1Rkf5B25B61aLNm/IXmpzPrV7Su29wSBwzD9k8zmpLs2ySq
a9eeir9yYiEB6mwUeq+j9UQHs0gI3Te0MNU2xY62BAM+mSYOM69+QMjkoMtD5qAuXSQWisvRt5Jh
3RnKeFrY5p+/K+QTj7he+zNvi5apFTnFg80fqWg/ybyUAplniyQCdHFDt3aS1uyrLtI+eQ7J66hL
LBnrwVfxTar8T2yG9Af7CXfyLILYDjudrmj9obvVcCdMt0H9p8QHySJQsRz9NFkfJMpDZM3kbYrb
85raBVZDBvEulD2XHFRhaJAvYzV6B5EY+qCltw7rC064khkcQhIK8R+mBz/YR6uL/uQ6uTWsw5DP
k+O6iZ7AY/uWWSwjA++KntdB2ciSCvYpZ3co/CbAMgPdA6Ty72p0YApSUzmGe7rqdv0IRggegmeV
rt5a05QZAiok/sZq+/cvnfVsSL2jWx8iWilUSQOwdXgdaToaHXO5sn7ZgUKrl5a411g/TGjEmUVX
8TZdyy792ZNCKpgjR/GraUcJRq1JoySfdZlBwMVHJAdCts7v21kadDvHv6F+iENfGdHQXfLLyvjJ
lRASSrQVfwGTCfedFBXBsGL7MtXa9S7SJntcrsYN7MXizmUXBFYXbpxlH5Tk2YHV+xJpxJTvFciU
KVL/T1otke3vLp367wMoSlmVYQBWPyTtIoao2c5gfNO4dYAodPRKBSXWvIHCwYhUCIbwi/jdDzUT
XBVtHxTND/K+7o2iJOf4Mcn0OVxK1xeQJcZ0fw+dKBDrOEiQRI8WQNjhDsrEOE2ni52Kxox/XTwr
qTFa88wawD0LGIqXIoalSwsp8us/3iBi7gxatvc5kdt0lYaM2UckPsEhSRkbsJBIxYg7U1EdBbQG
bAHUXjiP5/LU2bVse+DcbLrVVCZewnhsAhmPvnUin6/aKpSuNEuu1sRuYVP0ZILE9yfFh1RZkZsH
IkOvbJpk2Pt44sN0qcJzvAQnIaFQDyy9rR6vX0PuwhJrepvcIqc750MtbJiCAmSSl259YjyEIjT6
Ob+7gk5oCzdElMOJ5ff8VtIbJ3mqoE6Wtu6hX4ZAQ83j8//II9BLdgyIV2/eGYtOhVgCpVRTS0Ih
aYX0CbGiUh4bCEThSGFGVwTvZIyQLHMF8LLg7o7Vhci7odYeYwPYyQXEfo6ro+dei+HayY0intGj
ODtiEMNj2D6bcdmu+OkBVD86evr4JnE/Hbdet0xHsHPB1s34bRvILGCKc9U1dmHaQXhxTeJeeQq+
DO+QzebHKw7VbMHFTCSDFdiPL0alPL+78F+lrQwxajdHEV7dnPwXgKjFKBfjfxCyukSU7hPsyESM
WBs1ZW1eOp6lv8/UshyGBwqC+7JyO7G44l5tjrqM6SGDgrNIO+QdwJ6lo1th7O4g+TxFT8IxHZSa
u2hQ0bjZ/OxXarOfi82TBmiKgaUoeVLpCqo1nkxWhccxUZzGiZfkxdvtoRnYlvQLCvIYbnLYtssb
PgG4S+RYEJKvFl/TJLzh6GsrcD29m8FF/oQXT7iFBwUio24JSyk2SfBbEbFOWfAuuNYzcJfRA1/J
fhIdhR3rvAoIgSxtrdz9vH87bPnQs/Lb5u0H/ia+3eW8+GEt1+CN4DJtoBHtsXALw87gLpJPkko3
hZenK6ua4kRk8ZLankO/0ZDguONvnV6tXPVdWvt9zKSGxIX2am/IUllAf/AnfnM2UpokzgQaAX1l
m+2rET8bwy505BHqjSA1nYC8nrkHwNqKo5q4y9BGzrQWVqxGAKBIaAxJon4048E1oAhYPAhQFi3F
YWXRn8B2ckxd5NCHiWLdmuckYz/ujzs9jByQPxedikkFc6us3Jh03q5UI5SpF0QePWVlFjVhr+jr
94iktfy4IAs/68FfhX4Blg0CstV1qIVNw5CZX95YaiBxhnla2JFGQO34HaktL8eLKesQxHChIVaD
gZienPivn5ZKVA2Q6xYnC7VDlc+WLSA6A7kgjaH7JLnWAeFQlFH/qr0v8S5ADfx39dv0BlHKIKBO
4xjbqhQk8IH53i4yCByQL6o5vddz7dxkmHt3l3lopoTdDqQXCxWcAKNMr+OEipFanAD6CUMnUj2D
bau6TDCZ5GX0CD4PucZk0YfK7z0/c3xlm+CIwotH0FymL93OYNj8BYomWTsHO0cbquwGj9AkPg6x
Ebm/c9dgsg103PDA/IxhBOosQB0yEBE7mq9Xmk8IJ9TfHA8l1Xwqc6olNWrRFe4C2EGozok8d3M+
MM82wm86RbtV0QoYrAqpuoqVJb3RFD/twOd+U5MPdtw7gPFBqxbvHynRhETHIL90KsVHTljeo+q9
MImUol0SlCWD4gL6FgoM7O/En5WIdUQPN9P2hmB+ZkO/1IHaI1IA/3VYFtJLXqulFv3mqX8wadJZ
XK95cqCC12aF4QofwvS/UuL2wr/Ctn5MGESfYD14n2LGqaa8JaUXzjND7sq6pByTUl/1B/C+EOea
VOtiCV9JkUhZ17aeRDu+BxhcHpnH3xn12In4L5wFF/hG6w0QfwNt+8ViZ4VEZY/FqIGnduYeB5vE
psYr1vSsrqbto7RrmblZ47m9mBk+MEmEYLcNJ8ja1v7MX2N5zjp8BHfMhR/erXCliNdGh2rzOYMy
7CSwcEQ5nbksm3KTYJn1cqQdgQWV4iTadwruHnDm0HEZR6Bs9arnshyRshqw3aRffhgTBY7ZarTs
3yZGdl61P5pY1cpEe7lt62Uz+FAjoPS5Y5sgODXcJv0VPEEUnQnj27NLjSMCCptjom24gt1LTi3b
s7QRSfmMlZk70AlM9JYmeBSxPji7VwPaiOYAuKA84NyKB6VxJvYWuV19LJqiK3JexI5y72dt1MdH
sf7fUN1bZEUrccilAw1VtW6htPP1B/4bvaemhIFNZtw67TGPlSmBNddhV4Wbp/qDVULtHtuq1x9I
2Cro2wqIPhC2L0kuB4J6jC8swr4LkXAIIXJTBEgtWGtpgMN39AyochAcK6Sy1iev4MVNwuqnYHnC
sOL2rbyF5GwqHj8fajDyGAP6FVP/Nrz9E/g535EMR4nUAXrTP9nPNx7PITDqgl4XukbMr2d6xNek
pX+Flf5DYyFHgZEFqOqfpNJ3Fxi+7AlbU0ZqmgBnb1sQBA63GyCjf9uyJzfW+Q3G4c4KUQnophA+
ktzl7PBCwNqUJGpSGtpGPAuRI4+0Y/B656RDYeOJlTPnZQfPICylsM5TqxyZr+csp2DFP6UuyWhZ
9HYSzd2aGBq7tmH94zRj2mqz7I7IyCppMSraVP55entXXe+2d0zZyx5Bp7+KEBrDEDqqMfLJJ9bI
FUiY8TJsjiWKu+b6TxEgsUZWS8/GZDm9eKJmLj2aOyMRW/MdGPUwEwdRVB2PHczmzRMEmgTxVtQI
/gBgMD5lHkKMUpBQvnOS7nyhM6XENXZX+FiQzfzLMI3LqT3hvFv21HzB1GtCbkKNv+YjnPIXDsf2
RpbgsQbbM7zCZqeH33B5bTb3uUYwobn/D2HG0W+I7SZUiv3F0Mr7kD8xr5IdZHzIQ7LjGxaNWuCC
J9PNk4yXXLshiCNWFem9Ey9wYcNTjCR/COl3+Fcf0rGc6VwYBwAKWgYxxE0zrDS1J+W2fHDANAci
KgLlJG+LstlLbIg9TBdqehTfWQdDH8V5fl6dp2/pVjJzKB9jCtMz0XIqw7NPaeYKTy0TzhbJFatC
kp9cRkD9Q0V/Am0TiLJJHJgq+ToD0/7I3RRWySSKI6+b5gWBh2b27nqoZ7yilzOLR9HkdrkpDjrJ
Dl/8HO5EmEzBMrsDQT/fd3gMfhC1Uo50lF0dq+p72IHhMBtBgyeOPyRiKIJWm1NFGtY+RVNmbzMv
/eLfcG4XmGB5A+fun+3ohSMqy//TjKqHsl+8jddGWfZVsSQnj7Wt8b63FSREqLWUXI9AHqzRcN7u
SdNSY5xCPNB4btYppUecTzo5p/A+tBut0K8MKQBdmAcunSPTmANXIl+NKvAY7Y7y20mVpk0sZqfp
UYF98Hbw6yVkCf14XiFjAbxhLXnRpk6sWfbsrvEJvCk9+0cp6ICxImpdhGoe8p6LFNRUbVbz4g6l
7BTvOG+lhkocW1lqq5Xt6WG53BrZVQtIMsDN5hj2mG5OCr3q/7wfpEn4BByC4z71qFenqwv59p26
awVAo6efgYc/i9rxy+kL/wzra4JiEm6AaaJNw7bMeaVlcNDeRbd0p4itFbtX68xqC3WnOkA0EVru
05Wo50pijJTeyw+Ugpm5mz4021cVsbTGhmDxAPHl6MO+pvMZkC+5dIC6t80kyblFnWQlEBaDkjR5
VJNNiTLsd0l80UpCh45SGVJYHznYCqVw2XciOe+RYCbziu5u6HL6dDyCJsaefxQfWxemBXfriBAE
Rtp1EpGaRL1Ol2HmY3ZW+yDFPoDQuW/SbqWijwMS6rpOrhwuPJupGGEAeJwfFaewA3DM8UAxtzGX
AGzBVYzru87DVclR/JqhgVo4pw94Ei3E/Hr5LW3zm0ztx2bAg8asC5x8nDpyLN0BbTxx9zOnpAay
CqBjhIKeBLlvM/ZRm2St0z7LmJ8tvERGgOhLcnKpCOpv0kggFgAzmfQfPI0C0yIjBm0L5VDnBeBk
BLTY9Ro9W1n1qVaVtmoTPc1URXeK+fxt4Dlx+jbov/XFUxG/zlgiIrubbCrAJUN0B+LLqQIAJpwX
qYWPPNguZBxd1Cj63RhfWLxp4SrfQYDRaNV4PQyW4VHu6cJ7QzOKvYQ3u9DlMX6zTkBgEu++qAlK
+pblvB5kGscGR2UruG95IG5ckDLvNV9xn2ebAujiiFfht+/cblq8r5RPhWpRLhNaZ35okqtMluui
AEixT76iGq9FESz5aivRLJgOc01DyG+iM/iCcRH+rN1JPNjng80G2AZFPKmlejwEuSGl/T7jABd5
CEEFw4cyT7eeWRBQOvDN0GwlgOHlcyX1GgbPZ3bn3tDCVGauj+OqEaQwHz0VBme0+iOfQ8qk8c5S
Nj8O1G7E8T17XMgEc3oYyBqtKuVxeM/UzE/kHGNb0UZvi6Gu6j+XIXBkf4AldQcqEz41qfW2X4Af
wzFskqt1RJSS0D4COliKsQ3ZgWXOIAVcsWMcq8f2n7fQD23JT5FGvu4rCmEG3ft+QyWx51r8qsjO
HK7A6A3lyBAr/6imenWTZL9y2/ML5pg9GAu6FoJdgD1Pi2ZVwTa4r8z5LM4GeSPp8S6F4k64YaAM
y4XCVxPdYT3w2k+eU7AjMLF2MzjYhu2He51E79bM040FoEP23dyQ3O9SEL9DSzFBdDWThQnbJ6sf
sLQUqib5XASH15RvNPQUKxEsSg+dLIpu+qUOVfrEZFVumlm2Res8S/mlSzxYeo8HtoaDFRoIDL2V
8fkinqPW4LnruwNgvZ6o5vTlxjLr1fAVEi34E2holghI1uhptCJeutH1gddwr9OTYQWfWMREJPzB
VboIExeXaOM9C4gyRha4wKJj7yBj3WJ+Snon1tXM9tG83K/M9vVnyvE3zWYqeF9Qt6wxqaJjH5KD
wNn+wgAn0xg/cRbt3WHzrYu9ZMsKLv7d6NZEkn9zLKcUF1FYCdktf5qzBQrKYo8EqDgwRpr7lHLm
DJNol6PaxjmiA4BYHDlqeIJ4tPMvM2gD0v3TFSOqxvUlZtVXxT+WQxv8LHlg92i0ro4OpaCIpnQK
Da1/DAbgGAwRfNPACTS7YAec2tO8xUdgeV1fQ7V/NzKy04O924sZDC2n7yh168OrGAlDLYyldXkU
omgnuCvKSi1NDIBig9bu69JvnTPjN1zGEq/Evzvx2gexZY++Lavwtj2sEYqUeibvAoxI06/Hp8dX
v1rSPsjGYXX5VuA8xOSmn2pynOr5aMQdvxCAAP7ReILSpxZ4yE+PwyRqCq5a+8kDBnkDNha/f7HH
takzaJuatJb/tipqVaCFJFuJBvgNJI3m6tVYiFQfTMry7GYizM8iwlscJZ0SFwU1jAOFbL5F/irx
9vwQu+RsEPBr3djexb7CBwoCnZnCsYUN8Sea0tMnIpMxMhILpBDFvW+WEfjzbc+mgKnotpHDU4fB
GAHDcd9Xi+YOEOOOVlLAjvgmGU7pnUgSTMe3cWs4sZuk0l5gLJ6C2pm9TAR+Gf7e6vmQh1b6YtSX
lPx3dLGElBCFRq01klqaPr5wBhdJSObv81fM2yZWBKqR1yAYzWza6RC3huF9ZPXicOOpIlIsgUER
XuVo2j6IMShBpJxnutS9MYwq6RgY1MJHsdJNCr/4KaEwgTC+iTuj2+MhZYVs2EeqP6qccLHIZDJ8
wSl/l42ET+N4i1GyXv7NxQVDY5AwIFbC47bagVVy9/6GXSJHYrNTbYwBELmkXblUxXypj4tWhIvn
/isZ4LJeKsWRQdyAQl3hcre4tQ4P3vq9yyi+MzMKVWONFUbZYlFYWZ/hI9AMkxRpXP3+WS4iKVxA
klFpvttkMd0bkeIjhKVCUl7iybMdqZkpLVOMjB1waj10U93B3EnQ1qWLqQngoHpd7OTcdHh4c8PS
2N8Pu2yFi2Ju6VKqpF2+AeBeQlKswTqiVVEc4kWGd10m7x0iF46pLUyMBLqBdQ1XcSmomGTrfAMu
IHcBLTmxalUhJfKt7GOmEYsp1czmVllh6+O/uplkUIbBtE1V3RJ8DYNA4NSsdS2Gk773vRCBQMz+
WNquszIU760V81snsePLOSKWo2DU4LTajLejZ61EnU6nRgSzD9pW1YBNeGb8NjU82o8aMUX/ZVj/
MyaFgLsIgilzWTHwX8o7g+bA+Fl5auKWrJowOXDQd1Ysb1xP2QB/qn4Xj/pTlW7vmobMhpqw3ay9
PCL7fXOnKNkHkchGcj/i1t0fCJ0OLUEc5gJFcJ4lc39iL9DJa8EQ0xZEtc9KgsHBhbqZoKrODDgd
R7MV5/hb3fIBg5ZQop5sV1tnEBpi0MZsS0NdOwPwh6F0MxYiRtFAEqY29MPlKvHtQoz90ych34SO
uNQbejZyRh3+cS6MyR1R+4KYQSpVeMqtYWRqbwrPbABvOYgnuboZXim5nvjeMFYpioRBcGYZvBp5
iphhYVjDjp2boL7LwOWuO2ofutH1sVkfsk0QqhqYkTprEf8ntCAbdFrzGVMGa2VCvStPQ+IZzl8f
MHLnfGPioVQLtafY8pGrtBmqDq7p6grQl0G18VgwBGkyE0iAu/XbUlXkFqYZC4F5/MeUmY5xPvXm
tYqa1HQ9+i/JcIWiwyBC9AjvJu4yJknpjSjc3Z1EXXXkPUM4kuGqAWd5lgJ4POs3All/SKgoDaJ+
T8vezUtcM9FYVvHcgwVvDzWI5AKG9vnD0JMDEZBU79+rQrEUEZXnOkKe1qnp8NaMBNBOJMHhkmBN
dO79EQfHgOETBO633TtqSeFjP1TUa95I8ZHx4cYWi3znBlOr60t0HviUehiqvtwXSSqrCwEFBUK9
7orGreRXk/SM5RljxUHQqr4IVOkFJjOpqh1ynL2MlWatRK6JBPzI3iHg6tuLoPoiFNb3CEsRjDMY
CkEDlBR7gQlEo4vn59rrZXLrAVZbBRaMEAMJMCSzPiTT87vvlCTETQ3jeHC8juTd4iODPVGbg6to
vX9VGdyspfvkII6wJElOkMu8xwRRg/WaHggAQMkqnEvAGGIZ+yUzOZuPX54uPaOtsUzsjldQxAbl
V97niYc5yxcHB3mSEP5os5fHCMkJVKacETBQZ4RNRXGybnzim8iHl6yB19DUAl4QmpZJld217Klp
YVOQOEbe/RJyF5n/el1yFoUny46QHaFVDRyeLWLmr6U2fI3WhewAvlKYYQPHE3KA23IEcc0um/Gx
vI4DdABNxafZiM2pR3lhjCehMU7/nLh36bzg1haGsa5s1IV3lVdf7/p2kmyWoWsPFS0yAt9U5ik3
5GSbCDWGnnfbG6GrMlXbtk2cZFZbZOCs3bYwjUNIIUoJcPibwTp3l8qu4aDQwAoloNybZlO6ajWe
yR9odjpn6y5b0fDESYCnYl4NdYCcc0jOTEtsj0K5q4r2E0+qUYjFBAN9uMSRNsBg/SMW22MPLiky
1br3/8usz929DO6dpr7sTJ46cqk8BvyIcd4gPskYJbNZxDT7b0gf+BfgEWagCuU1bTBxwUTt9ynw
1AM3o7O8TA8HB7XRGQopa0b4GITFBLbVTjkR1YeweoG9/iRWnfNVL5Gm8sxHt8OOqQ4lZQUEoBIT
eQDlfWNHv/RzYL1gAgJIW0+Nn7XfNKwH29O13FNnsxU4BJnkTJ+b/3kElQTdDr4heWWA+NP4lo2i
eg9HQoCid0kHJeJ1KK9Ja6DF48n8PLkgBc1H08TcTobMZGHE3tEchBtjwTcFWWJ2zMrBZIRBivvE
8p9PPnO78gXfdWRMGeItlCfiK2TbexcGLg/VaKQrvtn7kO+BcvUI61f+Qc+yGI0tKjvJvj6nwrn5
LkG+Y9LtyCkeNVOyyxyfJCjvnqWDKJYrs4iOmgHXQ7mGzHG3yfdmuHuG5e3hOSu3TKy58wFv+VZY
A0+msWzMXLJ3Tjpol5N1N4bAVLfGEDUJpKk39pyV8eZX1SwTE/uF+DHratvr/UYH9uIQGEtDiyqF
CXo0uWdTAPXFo/VAB7cTrH3IzPpzlJr6xFvd2N43c8NM702WxztabxYkP1LY08S4a3hCHxrGFZBf
jsF+d/rhmPiGQSEH3C+BKkrCcs6zqds3XQE7Ug2U2qfB0Sg3rIqi3KHRU8RfobsEQRkFcrfGN7+P
AwDHC23CdJ990hhPJ1JvkCIcFrNSfTQE+ZD9Dx9fQcFrM819ITORmknUPM2keH3i5jXhJZ7mW2GO
skhqP7A5FlMQW/BOLlQ33eIYwkoCTdjM/aAWWYtMDwzbduxzi3dCYonCMyV1guZbIOFfBqTgA6Xz
9HgdTeW3g3QSWRDHRJ/3sPOjPnop5SRa6MPxkc14rZkCXn67gHc6z6SMHTBR/sQ8HwcMkJpWA2/T
B+sRRERr0k+hXJ8iYFZbZfeqjZ7bWhjVezTLj6uvIRBq1UkooLjZbvVmt05/IB7dt0zDH/rR2Rg9
HuvuJWpYdSv7+xtFDH46YXXvkf/K5hnEmOdvW5uA+GXRBhRS9x8KrrHqUKSYdH5zDPPit/EBF+Yo
y99ZbkXA0poa9bY6TBLdUyd+U1spuqoBOA4Th+nKtwVnaBMwVoxlKlJXkrsv9kwApabxioXAkRXA
wyt7EL2nOAmXocl4r1iZ4xA/FBGXP8Q7hTFGihdrxGyZpWf2fxJjIJE7sSxv2QzF7xfZcEtLeH6Z
D6CjeVfXujKgtOI2r5RHc4/AaUtppcPIbN4SF+pAhSlJKrQmJgmiw8w2cl/1wbzOHgtxgx8h28fn
MeqscdrbYcA8ykc9n9b3M+AbzijdMyuscZID5EqXdRRbmBYR10hZNkoX6yhEUexCZgSuHzq9vRTn
3wTOw46KCadsxoaL3mvKo4B4zOW7csAZWTGE1k7VUBMGnX93bMmPbsKi92qQOSEg6vYELT5rh9f1
ir6Wca35fYFTCFYbxY3C6L5M2zjyFPRWOOT8Fh2YCrfRc/due9FN/i3nCxhUmPbxDWZCBfHBTX1h
s0W9nsk+sqHea/QNAEOxDwei3rUPhQCOPmcbSb2osbLhusDQk9NcahDf5JRZW1Vvqcj19hX+3XY9
PqVz9Hca7qsMX9/XCgDcybGEiuIrGbfvYSdnls4IQW6HX28ju9gNDL88/JoV08QC17GD8jeBdy9+
kNA0Ze5IJ3e59MK02UNKBza9/8o6esf+TpSZEiop6Amemf4jtSkvYl2D5/L97R14f2eYPMOE0m4d
V4OFfWiy1R0zB3wQUc1ApnIv7BuiUQWZHuI4uVt+APsTcVWPCFESURI7z1TCWn3/avrQlImvjHZI
F64pqoipvfojjIPi9vPmg9e2jQJ6mrKDXDCdJrIy6oLWYpZ6gzajnzepZO55okPLgtswTTf3/TUe
A43qA4fWIkIKgLzDLhJ/9y9E/Qm0M8kksA7SvTeWwD3jWHyYDDqRoGGwIDS+i8C547zF0Mry4ZgC
/VpzwEESW+2Xqvu/7a1vXR1fB96Sf2sGasvT+ShyoESBi0yo/2dwt3VXHO4FjQNXUoVm2UiV10ox
W2eN0czraW7lJ/Hx+/V15zlK17J3d28fqG+jIjAD8KnoJIcc1r7ljVmkTaX1Ahc6euhmmkDkxb7e
j6G5P7qwlu52vGlyvercyLk1Y8xE9K2cwWiJn9iTCFl4aroKtAPzSwArc2IJHIFVZt9eNZbtxH8c
1HVi1Q1jCU78HS9ZWT5Qy56vmc2zid4tJZ36uazw+cDYV2REm8nGxFC4AGffHHjwqD/92K9GG4OK
VWlvkDXm5TAaKFrVkqv9VKegLyPqpvjWn16kpkwUi/Jc54X4G6LWc5x8+yAPjT2LFaFMfaVM8fMA
57RFh0WI+Vasc6AjdVIM0GDBgVSmPsujXqmZgMuDoMVBkWnsPvQ0AqAN6pkAP6/Aa8/VCEQhw5Ax
8QjhMd5uGNsZdI46qPO0VrKwgRqzxkBww2vH1XBhMAoDDwIQGUQ14YwyO3Wf6YUfgFwTVjX0FlC4
KLE6OwlGrQ4FS4XDDKRXOvNyuo9wERRqMNANIGO+sVxxcGCCWfTYAFRd74YQ+e/EG03mc24KOKAd
vrZlLwmniEqu6Q4LVRDYZHvGTlf2cHeq3Y7Hp/OxnWlIcXmg8j/6NYmN21p+xAvDqHRMLcViLQPV
kyrME3gwMpLGzF4auiLBE5CwlKPPiaLc68T6Zt16nekOi3g0XA0W2yJYq3Bf+YwkZaBZ7xp5rdTc
Tqs5r2y1shUME1AV0osO/9FqVQzqm5lzkK3Aeq0soWyFBb7y63ZDNu0U/zY5P9bD0DSfKVHWtjZ4
HWzBJ8FMPUCZiIu8m6ww0Nxa2B5kc9vD4Dc+32IJa3qTXNruOZmovJRZ2IcjJt14hLqaKAek+2J8
MM9yZnfP/2dzXAr6GB0mA9MHTuYWvNp9KZHl4kiJ0WQTcZsJgnnUhSAWOggqyzBAuhbC9IkaGxUw
+B8o8s7cbfdt3F9ZUpL0sQli6/BnstYa/+BR8c/iMqJWR/zDyxi5TksSafliBWTEpHj7QNw7mUNX
1lR7h0HI9/L808SkcCiInL36JN3ejkPWNH9mDidoHGBvvyQIXKk1k6Igi643TYYETek6tdc0GKIk
jZqIL/knd3XQo/MgYy0oan0oq0geul3T1xBbxmA53OShoIh2sTZxlf9003NajV5aBmTAU1N7/CCA
YPB+oO1KVIGgjeSAfaXKqrqmnwfrzCLfXshzDuMJrQJHfZKGd2qqp3/9zauzHWSbTZxd6zDd+W4h
Z33WIdMUlHa5ci3uJT7dLlKxyKgZ7g0kiMj74fBCS9S35pm70ljXYxLMAPLFcjsMR//2ZBqrIjfA
nBiTQISWK8UqYNgCzqSor5wfNAm9SDkROx5i5iEfM/P2aVbJnZxItrCVmbaxW++DBsWsED8yyjYf
VE3dZKivyUVsphjI9ctkwMqB5QC0XPvkCci9ouk5i2yLwlhAUe01rGCFmHoZ1SB2UZ+mzTijwPiN
hbYF33f/h6ixkfN0xEbK9BxebgCHiUDjaNaUrSefzqjUSGSXjiaGrsaC4On6oB6jT6+oJyc27s/f
OlwVlu7l0qqECcgkMiIl5rAvURIxKKLOlalsQ41ozHf5NiTKWXmeDgeILzc0BUbkTkK+opVv99Pj
ySTtivk+7XXpiSoN8PHQTReb/u199E6aaN6Wi6tpIxIv4QsBdjCtx4ikQECatcKEnoTljT6+lwf8
YklEIvkMliSfhilRTLH3L6A4f4uhN3HiGgfjB6eyo3ZmD52LC+76BTlAwJ90LU4ihWzpHHMXSwsB
7eU5Ug/TLpNDkcWzJc7P6LPFde7pqUsnagxgK6uh1Y/2IZr4qD30eG1HEz+qumzfVZukRL4/SQ1s
6sZH3QaBoYrVxD6DFRpzZ6eBr0tsV9M6ztPaxcv8TxYOv8Aexs02ydji1+G3ycokbQFphIzP8FVr
w23Y2SzNyH9R7qH4YdJCZsfTI9eo8WbdZ34o0abxfuL5XNVM9POov4p4Szdr4YuFp4uXq2hxAU+j
ExcaZu1kzwnre4+QdBv01exywvtG1/3RfJzSUzOQTjd8wwgKozj1zmkPgZSsTskZB7hfKwR+ZHHP
wc1JsbfBucJ5QEooybR+qDUOuJ9kslS02kKtJpJdXqc4jfjPot9MNbbYBNOaeXBoKDKeytQefsWh
g6M9rKF+lk3w1+Y9Wwon5CCIhuFXccoqD+aoaf1L1Fb0nEZYSVa0XTN4lFNFoQQM7H5K4Efo6Ij1
E2a46eDE3UR6hR8bzpL7sJPjNyxSmYx//5Li1duIquPAS6zC6tJVNLqHx2+SICdPcgoza9XOG5Zs
TxtIhPYFS+H1tmXiUHMK/SaR+zW2W6E6WYEdw9POrBEYiijj1YeZkHYuGMMwaDveL2Z9yd9L6RoK
ysY6TCzfDvcaC/o0c61ydCPUGh97bZ0gEaLsPry2dzuVRKSuEoRFb3B+JEgqwE5R5pkTNv7XiQeg
yI1KhPepJl5UB8IjDstTqIJOJADcdI7TyFVKHsQ/VEVEE3HTU/LegxvU7BdD06cvwzvMajPhulmS
3JIWtNgsyjzh2jbjdYs9ZLXDkNyHH7jEBD8Fahgydc9GBiM0Xu6W8TGSk2g4pZi/JRGfPulVEOeQ
gJfNnkJl8TWVcPgILjDXNuVzHmAX61bxbKthwbWbhP6+VC2TkWERx/ZWUoRcm7bVrWjrft7mYXrd
4s3SOxMvtgtMknSfn7poXgKf7EJQ2kDdQpNTYRNLHaRVi1joHZMF2zSgUaBr7DrxNywUl8iguBrn
z+UJi+MVOIfxuaOvGK/wdI/a2DtQfev7iPu6XwOmrmzCWOtIXm2jsd4oVRF5fBG6tqvhggcVQALL
+rh4IS8zilEIUaECDUXtE0nDchWxdcixmdSd2G6uRCZ5Ki51almKV9Wyq8jkOgo6uY6XD96wBrsr
YT4TfpRzYyWjMSsMvb0DM68Epgkdfw5QGfwPdsM6JqpbL/I49FYIXDicgjPVxqPjvuyboPL2pWxW
IxSrxFXV8iOfR6WOAVsG2H/+93vWH6KJ3xiGAnGzyG7iSWK40+e0ddeovcwGECDn30LhFiyQNlxy
IdDsBGBx/Y2UW8lSWYwMZz1r8IvaSsGw83lMbMggNBr/T5sCSVP2I3Y1RLJoucCUz5MNPGGD76yg
tXU22xKcu9yhKXjHTHSPtbv/K9EibhcoYVmrW60JxBoFvs0PrlAwYpTQeXCddr6UHHeECIcC2cfl
rouM91JhXVt20JsnYhJd5E70JLY1fdTYYKJR45KqMAtsN5nmwdgHO15Wm7YLJAMeG1xHmt+QXO3O
zn6xe5Fnbg82rK79ocjdrJXHF6SKa8ZZjaQ6t5ySGUkUUi60q+cr+Pbw/0d7Aq7TlPJpwGollGdy
UjnZYKR1GWr0MypGbPJaKEUZr+wms+peay29L5AEIwcxfRfJ2OvWfRFI5zttP6e78OngoBMUd+W0
+t2I7Z/HSA9OnOIWsTesgr8N78G8xmL4D3aKJn2DeHj11QRlwV+iZHQnRksGS7lgiogCLsclGSwM
6HiUtAiCVKQggsfv8GKSD4hw1+ubNFX2Ch1bRw0/Faa89/5RW1ljFulwNteuSMgNFbgCuvEMwU7Q
n5Xus/3XNJXw83X5dU+cAHE6GxJNR9pfbWn4f0t7Hy2rWD4/GzLoM1fbEqq2m95SkG0xbHlyUirU
/hVyr3LT49as1Hk8dcnTL1+Y9C2E+5ALPA3NW8UIoss7JkWAkOi0IvgY6iAZ2agrkBcqr6AkjEdB
wU2fVQGfYVpN0RUSIPy3iwO3rJKiI1vXNcBTHowGNNcyuH9E2m92nfL+1itxWe4hOSGd7m5xdf1J
BMoOGxiae4ivgkuqH/viHA6JWjNF01p88A3FJJ/T+jL0+OHGZPmW1fKetbGOuzxV1HRR3QrA6aAB
/apBdzMIGEhVmVe4zfJcHLeSOFrnW05DD8Us4e2teaAV3+TKaqe62YYcnlVTWCMXV9G7G1+tb8AO
eZT4kBoo1WiMWshxxRSYvhk5gzHMVJHbvb8kqkad6Cj7O1x9L8A/mF+gbB1aFs5lOCIDjCIQPqO9
CFlIZ4HY+2ubo7sgLwpFlbP9Q2yoNu6CzfnRKnpDJtwz9JnDwkWi/MY+QzY/xzyTPMZniuiTMVtS
L84cO4Bv3aU5sQ3WHLdC5J8qJQntQUjWngAvyS4r29di2SrOTs8bWjLTwoRrHcMatQkfiLkAsiVI
YM307PGDE4wB7k/G1b9MqyPMfBkz3taD6OYjAvJQpUqVtEOWov0qka9Sxiebd6mPnVlouemAh/AN
DSerk2wK5htV7KDvDCnp1EDNM6U1aOzci27PSN/jnbqxycwtV3ewa5molhozJVVmIhxO1YfR3PEY
55Mqlt/nRSjNdvRnxZgV2DVKDwoS5tYcDtFb2b5wg3wTVCMnr11VyA5ylnhy4AMLlsvxKeRJJboA
1DiIaO5/deR8ROCfnkLilNr2yLhSQfbxoOfsbBAz56Txs7AxACKLgVcgJ38+qNO0FdgEEgWDPj0u
f72u0PeDhdBuV6YjYmA2iTCmctRuYT2AEnuNYtS2S2UuDm3oIHBnyrtRwldYDigpV7aKPkYPOVnm
AeK27bQZ1e0vn+eRKZkCSAEF2lo86TiRb3wUkTze9mW6W53Lqi8Cw2GEtdcfRjhNbWyE5pSIeMv9
/wGSNNLcozcW5YubFfmZpF8sY2o4YNe9eUbfi1DuQX/S6m8xRt2CD8UhMDt4/p91dvdk1cx5xpkg
zcpS69oYJ34aYPSF0ZHxbasMhdU8SuGnCAynWQioqK2rE4y7KQK83Vy8hGqLLcCrrmuDxJlMGd+b
39X34kqVyPd49B96fPLJE2/cBjPNNP1JQ4wNexRQhrDnNOTISJDD4/HWDFaZ97aXmLFR2kBN+X5P
Wl00SmeV65yqhheuwfktVgy+NbM8EertTN+icUnlV905MKA0y3RqZt8q76Jz5j/NuT637s/NUpkb
ZMfHpbuyC9txrmoyybVdjtJPB03jkpgDsZi3A2sLlv7tCV+KRdZAB4OCfsahkVzv7ZEy11/Et2gs
vFyWENbrpbDHXn92PlcvpI2yEWCwQSG/D/Ny2F/aMed2zJFgFqGSE20asvmMm2HpzYo/Rpe8JKe9
lCxvPtTf2dHGww71NskiscC9fr2EknRLPW5g2jB22Q/i9JLxanl3cmQls11yihQO5G9+mIEGKnjQ
HpVpL3fx6y56zI8vCeScN37GpLMxBIPsQWBgy7bld+2zNaUeQUrPYiNlIm3aqKBvyDJl8b0VkGCb
mR0asgVwr3lIYGrFeqGzTY/m+tCkWaJ13qWAurqb9a/s1qmHVLTsipCK5mosjFzXIRWoIJt4prAk
46qF1LSOMgEe+1ByRz9J6j8FSpmXV0/2CXO42jOlpNInHxOzZhIdIwNewyC2jW0nTh2eArS6gHg2
J4GPPOozdn2XjwPOMnwta8+gMzJjUCJ8mcB+FWVoP/CO06hRab0rp7UxD1UQ4lHiyFfwNUD376Wk
NSi37iQIutbNFyJkgSMzHMhnhGkFFIQdHJ+3zKRvpdR6g042BPKmZ0ykfxVYyOxyw45RJD6O+2t1
dJ4DUxeVJWpjtXBr07iLBYOgov3S9bjs+44j5BvskPTk80+glQXItUa5JjoynGjmwTBVbtOAoC93
refmzow+L1Ftp6YBVPtMkAYfHWMPgWir6pS/wpoYaJaUYKTHSST+G/NNKgPtDE3uyCS7dH+b+FQp
ZHNoAFQD7zv11teg2FiBFDRhLfD0y+fZElADoZ4s/hdJuHPdaybfEmyhNU4oU0YWcYx3XYTxpR/Y
M4dbfdOXZeqPVwPquSlVded2xC6xHI7E7NAfM9o+WEUVF9YQnnYtL4v7tKYtvVFniHEEoCwKLKxk
ebkYSU+hPjsH6peFnS5VwfLFidGxqA3Av8VbsGtGq0DtVfBpWryTR80ToaqD+HpOGygSNK3E1yRz
+49fq9xruLAQ7K2H7FnpZ8jSVgoJXAm5HMWJJ/RXHwh/eISRNj0vpwBmA2BlMu2jHk6yfHVhJDuq
pgePuHloSPgKeyfaxvclZHajHlGEvjWlrmG662fyoPXH3eRwBpfIOaAKGwA1N9rQvcoSVONNFFFE
4yBmlOHsKOEFeK4TxYn6gsHGFwTyzDv/9yne54rdprC2uTll0m5G59T+2GKLWgpa6XQnIZiHSEyL
CJRpaSY0sKHHLlU1UWnQPw2Tk5XVL1Q2eefMDVl+Fncs6K5i8xUpqYCOb/JVXNPyFm+5r6RLYPMl
geINuZD0KIXZQOtFhhTB0yxKpPya3TLB4E6TdOYOHirQxIiMUZAAIuFdW156+pOKBtEyMk7B+HH6
k5JA3oQc9uzTVYumORU8Hvabwl4hsF32i9nRx5OYUIQYqZ9dvVQeL/8WaLpH0ECE5x6QZbHAwLWO
0RgZH2NURVTK0y4aExSph2xyxfZgViSY7/zS5A/BE+wKKOW75F/zqUxC8713tFGxxZvjek9B9WQ6
e7/spMevnssceeWB41l/KgoRFXDV2SeXpjKMtsWFCLztkfZpe+jviIxR0f6kHSs1n64xBZk+MUUQ
i0VPEe6OfE3jxYbrS0vt5pdF0IP7dn6Zfcw8dHSrXjs9hXBfpjA6957LICevHgXpAjmg2rBuFZoL
LStzpiBf1AzFyfGiJkhCHL5mwz/3uPN5G1m+0nobm8sMlkxNtYVino46VfmqiLmQLTUaxkRF/LvA
ghC5jtzM3TTTz/Zm0A6ah7iMMMNygTSQTOVliK6VsTBbcKAWl54KhDhQkTKyHCOFqM/RvXAVBZtn
4ITEVARrAChnJYCMxvA8dxDgqSuarX3CkIHEedS2zEAl0hjKpgzPpZMSSZcZbkkzT+L85HprH4DH
n2pCk1j60298hekCFP7N4F/fvkkYFts+S8c+aptlTuY4zbmxzOo/QAoNreo9DXUP4YB9ABjsrF6l
2+AYMEj/zUoA8tvKQHGKwaBjiqQWQrvu2cicyNRcKXQfcM8Iu4losHGoxJOaUAURJsflVeDOhR+I
6FrWmq+vBVo843Yyf4eFLtC7Oi7YW4JCOWPZUVaWJIdC/sPc+TbfGJLMZZqgOJaniQlDbAbm1hr0
iUs1SJVbXtGN3i3+7kfzYUhvR0KDyE3PvADQpKqUCAEWluQDV7PkcZg6tQgjp1X+8/DOYnnzBFZM
ZEuvqgACFsrRRRnGID/LY8dz/K61xnijOtx22HA/fE+JdsT91eFmYYDmvPL1Sw8niwE9IaNsIjMX
uuo+A/1GkcH1C+eAQFuRxzk0xqSZ1v3MTwKx6kQsnB87MtOc7Ek2QOz2K5sJmFgRCFXOLuKPfve4
+9iCSIHebUEiC8yTBc0YnFzsEieB/gDNzZ0eQOBlatNS+tn6ITuecm6Hi3/GcKU/Gj1d4TLMMca8
ISTRpBfrLWWkV57SzkqyXBUNGhMZ1fG8MpbRjTbNfp0MN8NaQ8TvLc6d9y+kqLy7EHyvQn8aqUY7
m1Yv35+EiQUlpx+hzgydF90/YxQjF0x2X52dageXQkbvyeg2/pfzrKf3YLWdLVXJPTpddSl5VAn+
5V2aRut5FFNdEJOvf5+zKrCjFIWLW2MkYLGJYhh2k35n3MxwH5Fj0itz1gv8+q80pXp+/9Pg97di
RiqDCDlmCqV8wL8y+y08acqIiZO+SofCbLCO+lQniLBDKvtVUkgUIwiXVtq22hqcZiQotU45g9Q+
tQh2Ul4mIgRh8nE5jDfPK+bix2bK0yWAzdZkolsZmmsYBAIv1yQ8Lyu/UiYkvQCdxz2PnaTvayZ0
dflAqUd5ZExStXlxZAyjUNUwiJ+ul19uCPM7daGHTCTlMdPq3s2uu0hYxICUDAFecJZKDYWDH/GH
Nh8+nsWQJ7bXKsrijQArc+OXHiFyy6ZPchVlDiBFMfEgJGRhwUcYLFjltuvEaXtAqhcnbZdCGyp0
NjSjWwR4vYYLkWg/f3rUnPfDwILZAGABzO16+Sl8xmH9TyGCRmbcqtXuWSfXPHV6RysmDNcdcW6e
aiMiV0qKofiW59kjO0SIK6AQv4IK93/KTpBheBg+adXdnj8jDP9BMtn8ZjbA/3p6K1smMwm5sccn
nBKXpvK7CYyJI953vo4CeSZYAAPS8ix0eSqjEKadbklTMwcYX0AZ4uYLXnPkZ7ff2EYSqnuvAIXR
Ni3+KcB98LB+vDi0dPGqKuw4PEN/oid9rljW0xJqeHS8z0GGHYn42n9ixpeVMUAHpQPapZPDpL7R
4VzlJHejUyHHr7sI4ZJDQhnNsRVwVI+1MpbHEFByuidb3Q5kBikfPk7BFqx1vJuIxaN11B4lBP8h
Lm8IPH5+3BExYKIs2UTGtSe9t/Eq7HVwxUK/nDXLfnC1inoTnARZ223tTo5b+DD9vqpHsAyCqcEY
lz1EN7zLtutgAnM7ylxDTra4AuVgk5ds72UP2ttbU5G21yDY/EbMOxA454nP7mMUA+sB9QV85hn3
NnytbmBAUaJ0yo0LEXQqWpwlVq6123pd10vGPjrwNrzBtv3MbzbbkvbQyXnG6quP1Ek7FY8imm9f
o9BFfsp4TUdxM/A6wNyZ4b8ICc6nTCGlZka8Y53WumYOvqzrs16rFHAfD+Tj6s256yi394scDfiA
cDx1bEqgHGxcK7CwaeGEvNTxH3LCBD/24oON90+ANeQbWFwHvBOkJ2RjU9k8nxSApzscEarSsPcZ
QKN7cHimZmSjpGMkPneYaKB9QuFmsmzU5s1gHIzJkFBqPYx9BSGRxjY3ristpjZmzwCe1WeCOn9i
9oEDXSx5gVFDkTFjNMpTJ5yMPMSROwXCogk9SN3laFypUMdWV1imzwgpIl5jxnUS+m1x4hdSEkvr
3zU8xGMRAntfW9iA+BYTVKrmkBA49+5q92buNvOGDp6njvfFUTlTDeyECftLRqeVWvQFNPbUQK2g
0B6z9UUnVAJrS/qUnhcyB6Hdb626krulej6mz4THolSWYUClknY69del3KWkCv+13yFkkZ8HUMVs
WZuMJ/RPJEbUV9uEgcYTlhFUy5hp8kA4MrApE1r2lmfkIyh+OrWZQwYliNxAHwGLKf1cgO3vP75e
aqhstyU/j/mWwGVirgmdj8+oN/i3MVN6qD+x8d5TOz0jCBq2XQv50Wx/yx4mMseeIu4aRna2vOKr
73wXV2li4WJ5UradPuj3/+5gFu4PwHsTN5UKjgmQChCJRIbo1xYLSNYjfq09Sp/K9kWJYG7d4D1u
lAPE73IhvBJy0F9KZKnHwWCyCWx9AIM+7sTh/VF1poR61QRVbuPoYCeWDybRklUVsZ6cRxthv32R
vQAAWOu+wMo0K55blQ2uwXGOhuEuLoiUu62Z1Lk4oz+GPt3LD+oxE2ihqNSY3/d1mqSdTobHe53Z
KVW1F2GI691GmobZfDvxwQar4cxhv81LUHdfSI56RvtU48NzhddmYCp0jbEaZR+djv5ZFcA9AnD9
ANSCwverrHaS7o6QSwsf16/1T1mDpMY7P/tG2NHVRJ6cZe4cSWX4e2SvdReHfdQy4CDitoN9a0q2
A3sAZSZj+XC42ZrI9JcePTrfq4TNhoo6zZgUAgBLGGF4m1EkOTtsEJdazyAB4M+hFlCBtOgZgnss
5M5vMj9fEAoDNG9jfVRvxUzOUCNP+Bpm4VKxfkZQis3I1uRFl1KM55r+r38TfWh9TbKOaWVfjS96
O7/2G1KCr9XF3bEhH0Se7IAEGXvR/bOfwXwpe+ffvkiAljGd29ojr+UuxMUNpDP5Btq9lrLxho/L
r2WHclFYBYUr1cneL+Ltj5VbwoeDL9BN6hf/rixEW7oTEniT63bI4ZJzlEv0KkXNBJXgCyFwYNyX
RWRW6UZsmBSY1/P2+ny6bjUqC9W2cpLkjuEI0LPVXmWz/CEFBOSEd0D54yzCC3TH5iETvR3bE6ps
hvnQvNqSY1R2fe51MLPs7mmD0vQVF4HnhHEQDHotlmRLjVz7k/yszOUMIfcMJ4dKImvu5D3KgCmX
gqrOfDpkFPS61DdlaqoXd8S2UKLshUcx8RpVPAMbrotpdOCqQMzTNQqH/Q5xhTFiLlyb6XSFdjxy
4IOgRi6CBBVjfoN7tCtrADfnZh1pxKf/C76p3wcHMd8oSmXeqFVKk67oenPk3jVdXjtJtk6hbvgv
2DKDsWBZzYiFRRMDmDUhdT53u/oIl1D4QTzQeHMacoghe02YdwpvFmJsm0ZyfddBnoD9EPpi+Jmh
zivBYGV5/y8hmpEjuO46wSqUoi9/7yjy7Bgfp6QPfYnQg3ViCDxZeoUDxmilmowLqjEOcP2EIlKu
Sk5+bx2PmeKv6nm3C1V4a+bhlUUmfB68uJKB5LXwDTkDu4FbSw3KNdz2kTucf3S2Jui0RrsPPqe+
pOYG/ojJMxRIiQRj7FvUlDHehGFvQ1N1ZWs7VoS/w68roIP5ziOznJ7Jsl0YrTDiAHOEi9426Icg
n7ah/rFaXXYtxmQMNIJvlehKXJ0rO9RQRKeOwl84rth0gSebx4MJfWZz+hUkUbKU8iMQ27xoZ4pO
2VXctZhzmKiT8TdFxr+txRfLutDru6NX3JsCoruDK8kNiGnBKUpDFe29LGzjNL9ovUwOt589Kwgl
n48w20ZQeIDN6GqrYZZgN77+04n1L422pI2wcfZ3YfMm5FdUhnONHAz3yCrjcBKQNV+0xgzKkHKe
hS+XvFsjx39HwUnQP4uHG3sS4ptKLOISOPEuolD+/sh9j846qvCPV7JQEGrZWKAMXAKIRNDJsVQF
nKY5iuZ4+ZFfiCpR9ODQse0TC8vzwySUlFy5+E3SYYGH1u0n9Xdri4N+JZTpKq44pg/T/QTe0tU+
zud1h3vZqLEUl7EaP1j3JtowNTJK+M5t/dt1vBkshqf43hpBiV8IKv+dlRu2Mk2j147wq56x7/CS
lEmWFK0LvYLw5HVHfyPeD+7RtJhop3VgRbNI3u0yxQmpbYtGqpKH6A0fU+3whXmzu1WucnHV1I2V
FZMQYk4zqk452HLFX2jXPKoWJ7f6gNGodvGTPxZNKuFITa+43ObQEyLYmZhaV9aQWbIZpKLbWYhG
G3evNs+sEZWaav0OJ992zQkq4JF31BYt7V2uUjq8GQV/ZGxJEQ6tbDJws5VyyLrXDgR4UVDcS0QD
AwC2FHi6XxHEMvabhukKP9wEnKhxdyNrEhkGpNGb1yxgXo4tooyii1H9CEWnWsgFhDgRqozTSq6b
FuHyurv63Yq56rwdBav/R3bO/DZjpQfnL314Cas+WT2C+lPYcT9T9iQ5HQvPGtvLDcySLTNK+yaT
h/dxQ+OdZG+bWveHebrZb4u1IgbPt84Z/BjJdGySxqlOUtNZsi7VOwnKA2bUOK6OlUNuNy9LuzKy
XuW1ynPiMMVsgF+ayD21NgZjNkV87nJua6VyiKTO5HPHGl1aM7Ft+b8z6nCY9CGXc2dl6dfibMYV
Ws/Z3oztgXSRAeYuckMbbvf01BA/5unZybJAj4QiKzG44QV3jYfo6eUI/aiuEY6lzkYKn9haeVK3
3rqQ6oXzB+vvhVd5xhEpemFbWy4hOKkvS722TPlhLPX66r4LfkHHPKaJAdbEOiYGUdg8yXlNQ9i6
TyfAFjfBKD6/qYsCljDTl2t0KMSgYRVoptdLGGIfjr1BRN8rnMlIyl20utzfiELFfx6dUK1pEhFe
Q4bqyFOxtO44QfFF0o0vUYytsvyF2PwiUFfQGKQ2USCjxvsL9m+MNw2g0MyfS78Lrp4fmoE0kzVf
epsMw/kMQ6FkPyafZKrb9W4/0v6icYxDEukXpL6sbvsFLXbDHGG2yf6K9fe5gHqOcIL8cXDUdRzB
DenEPGXgrexcx63WJFsUX4dBMXjMCVOzrAzGhoLBELNUrDO76aR6r2Jrd3pLRwnktJh7rL0RwU62
ncNk/vzRgSD6m7MV3q8DXBAoafQGi1rFg503knrOq4jcku4WyG/APcrsorzqjcJh9ygyvu5rK6OE
PjJWUxhtSaiLvy+uer0aZsDg4USquCoSEWvX4I1SpJG8T9dv4aUkHvgjtGIG/QdIWCs/ABperwCk
oQqyMvEhycPn8yH4xvpgu67an8qowUMHyVI6QZzV/kEIiJbtVTGRFstZQlRxWkqPptpHjI2KdLXC
OxAl+kEujeB/K5NGkXe4gF773vz8LL0S5vtjdgrfT29VDnIuTXPtLHiFf8/OhGZYzhGyXwOQCEp9
9HgM9vDWy7hJL5vAZL403EVJHYJwxGKx2/kXdYGPvKZ18Z5ePRz4BQTiuVZXDbFBHwyEfuJk9SqG
m1LXnX3ps6SObKIlmKL09ghskFspQrDQVuzORvRX3xm4+pvYcaNL3i3XqEp5wtJP+eIfDNpVjyze
/Jcqz3o4MXAwR29xuekpSi4G5LZXaG0U8CBRmcpwfZVmVuPPb697yQxXnpF8wi72nbLdDyqPS8P6
kD26IBsR5UaEnsN2RS15GcSVsT1yznbUDa7USC53cBUgec03ruTlzAm44tR/E6FJamGbZrpzaSCu
LGFXOn1o+/P1Cs0E1YdVW3fndhr4zifoAp89NkyEfl3qNr3dVyOKYyFV1RV4Wa6/9FldM8WAzCZA
w5wjC1+FBYyWcFJBmn3y6Q7kJDPxt8pXM5nI8SYVzJmYX17VaOHAbdbWTGlPI/ii7MQubYCh+TcS
xOnpya/viAXRSTwP5zLt8Eh6UurLSExV7fgXVVY+tJQt7FBhIuscF4IGYF3Wxp8FCmWT9gWIurdD
gsz0pLI+mc/sUswj7Y8Jg0ZMMzjrmx48UTyHa/ZhNq2lk6cDobSFTgdtaHzK8N75x7WgfZlyfn3L
jtFfesGcgT4R1iiWwktCvu74dG/Jr1EX+IEBe7xTouuAvNvPKaiMnJu6qafxKEZ74f0LumJJAFfw
dacl3lbzGaZraiIMXnOQZUeHvbvk7811DbgPiygaES8qxkkdpeaB54DukO5s2rq2QzbqljozG3db
kXVE3ijngR5InzQ98WBOMjhn6XWh9JlSksQvtRLuM7HXS6tHKy4j8/Xp32cFrrnUeyC84tBix6h+
z5n0X4SDIfIGgrgDBziotpKfUq7mzjD9Aiy3vxE9Msd0EzgkKJh1yBhWN76tKa0vZsuibhVHBCsG
FR/WYKfJvJ4PhOHcec6dOHc7KF4TdYvoN9Q+OQ0o4VIi0umj+kFfJONUSet1mgtxrdZKBH8E1FZh
mcoSYFAvAuu2NDbbnX+7tp1dObDYXzlxLklzqiQYHg25k4FLGUro2xdrfKZ8uifjN4Jzgy9wdTJG
k8Dzz67A0g6BJPQcOickgHrDyONHvF0n2yiZWyRJ5yCVaYP21nSX223re0NQjpruq1KDEYufNdEE
fnTc8BMcz+d1yRO/nI+DzKWTzP0/cZHg5Lm2daYhr3T3QlBo1QLNzzpqr/sxGBHAJkoxe6oKtgeg
pIjbuVdk0asxaI+dYQwcXyFwTQ2NqX0iBN6ZtwvuY8pZTcXdGpOTOq1uSl6vO77G3gNNh7xoCqL8
VFGhpK8QpHRhttqs0qyYu0MB6T3lUIrjux5xadQIiPp7wN7vTP8jY7xO15sne32y57S60QYzQaR2
5JDlr24pLGpDGfMRUAUJ8W0ONlKIMY3efpfYFBsuj58wMU9jGGlNsZHJRDjVptU+3pbz+IWWMGjd
zLL3Fl2qR+XQV3NKkU7dhhPEx3R7DS+NGIl5+R+RsDwOxrbK+PRxnuyrDqCM9c6Bv6gdCnIDkt9h
3e4LfNKv/CTK3pidDH2AQdSsM3UEyg2tHh+zzGo0kwCw/jbna6RfBhygeUDXaz8q0sji/mM59OLg
J+nAlSB2dMqxqQ+RKKh2nZ/KZBY8a57fETpexpEoSrgW9OIEvN77UvPbT/NWOhV1KJo9Qb36LrJ3
W44woYwoUOEpPrkSj3nLFaPbKGt0AzPcHLT1ejZNrqs0fqUxKYIhHKyIaSkW3ntNZU354ftYSJl0
FWD+BhAXQEupAw2VSsa/B1ZB0CLqE2QmVX3EnYEBRUkKz2NtS28AU76dUyWHavc2uX77y0vTg/dg
EYQAgvDT6z6k18Y6DJEDWUivVeOLGVzhmR2DTkCN7ZR/tuSpBFtz4JRRYlPeNwzaWZ1D1KXKpEVR
fnB1IlXgFjiSZkKOT4dtTiOWwYCK2GOe1Q8WRWQVt5t96//XV+6inRUh1e6TISXYoVKV10eGDRbn
6uUKN2N+yBNGtbMBtbQhJfb52oKT6jMV5mCLhhiJaTmezPYrCrzkju+yCB6XGKHsGaWk3gd6Z1Me
o2oSCyFyfKcpvkZWMj43lDtyeYLWtEd+qIF/vXHP3XpUA2IarkKThq1QGvjwYSHWqHAcUlX/ao8B
W4VkyPXitx686k0GqhQ1ma6czwc7Z0dfRX3Ck3Dn57shCX0232jvft5IqFJfMAm06GGGM3gTdVG5
Gz0A18WQgPz5O5sLm5EE470YBuCTZgJZ57x/+pPfdNHVHN+KAR9irzLYPpvKtK7WLUtK5ghDnCdr
V5AbuLX+H2s3oLNiBG/ifkrM0xxQmq4VGJEkulnsXPAMLcwCrY+P57OK8CtdTQX9yHPWqYo8AcPF
wmVh3+tZfrJgvGpJCub0vLhAwZWHZTBS6ujE8RdPLk13bp9Nk0jO7g6bPS1STQnvXQaU+ldPNjZJ
YdEDScSsDso7wWX0H93d7EOevSmx9+2jJdEyN2JgbV66aVRzMP0L3hiJ8aAJ7Z1n9/NHoVyxf7w3
t15AyHQKYOS2MXng6FrQFMaVZPLXTzX8hX4BtulbZiFjea/52on1PEUCP44oaIf61X9mwTu7lKop
BllCdUOnjjCjTKSCbG+P8QKvuiKFud0Wpxt+PovWScLNFEnfskaERhWApMd2jYNkVTvSDG1zphgU
ZMZoegJ5UQNPT/1AxYSX/wICnsuP9q4HN/sIc9QXyFRILDoXeZeNx0kw9WZLZshaJsq97NWIJDPC
VJtb47onUP9hTIK+5qBNImkkTWmYxFH2B/dcZFry4sO5LYs83yjw5XCD6wvaxDY6CXtQM3dnYM8m
Acbg70h3CZ3FbFop0tq8FXZ8epspQTfEugoYmNJLZI3Ae3+ZoHXNdBBMQVvnYJs4cbHaMNNCRziq
QIrHR0lMP7tSTZ9JHgYjnTpRCgltUUIChj4u/X8yz2zl09eKocSDnwZs44AQQqxNuGAnWqnluUKi
DzNkcH1K8eiIbuyDfDkJn1UM8SnWMrquL//1tGPU7Vfu5F3aVNXb17qKMxjwiSbkFf7dHxbHQB2R
p50xcQPdyMu+QzpcdvhwZSCnGBWU5YU2h/bnphQd4mgV2Cigb1iVA6Y73pzSYKWLiX7uAHdXDOob
SnAad+u5bqEwj+aR0v9DoFEHJbSV9MtJk2BMv6eVg0GXp7d7PQbBjQYRHQIyIBlouS/2JIx9KEkF
slie+2BRilRLY9OJ5+RcI067s2VPdm/scBvoHyBhPlTVhVb/WN2zxSLh+VvZ07HtiYq5KOIJ7hJZ
kLwk4XbWQwcJl6qE7MixO9wzoOMlP4DjMJFYipC+CsyISwL017vjd4FtFPEqWbTEN1PsSWFoPNrd
LaJz8IKPuE3QHtl1wdgimVEq91+YePEoK1wqrKBmjsCLOvUU0bsJuDhFUTtfeD0yFSWqQw0BLJWV
1SW+XPVtNiw/0pk3Y43PrC0BIUppD3RfJdhZZulBwh5ceRn7dQ0hzLxeyXmDz8uWpOf39LWjlRN3
gjXvWGv2XO+qSmyvk39YMDdFeMbBJtDj6fcQuy8fPEwdjomTyVczm8hlnp6kDCMh2Bw2cPCrpIzW
oo20f5t9lffBqiQHFrquJklHKY+0yeQRUUKlvXcn1JPuj65DRM5R6rpOqjKc94QbQ3e9Rc1E1AQN
NgHMoGT8t9ZRbBwtMzurneasyuO7Db/Jj4ByxT+wvDlyQuufF//D631ZkfPAh6VNf2kqPKyfyN/E
nKapHLMvrMHGVND8IpvcoTcHn0Caq5/m/BPVBpznErjRKMZiwRBpWrox9YcSbK0vV38tRkS1oSco
M+9TT4T1XFTjmi0rdkWzvEM3pplFzVCquE4HnC2yNwfF8YKVqHWT0OwR+ZI2Gn2k1Mzh6mSJTMbi
Z79pL2N71PFXwDSkbsBtbDezFguJxk66391vW8rVrXtktAuXMrVHSxs+7amN9tGnLN/nrK/dqllM
2dEibzB14MUULMk4RcQF7bN7utVoAQr4G36OOMrmEb1kuoa0weQFptB6mwbpzbu5kMWyCE9Okh7H
sKW1DUbwtryzha3JNorBRfCfNkZx7RtuvKVt1UAz8B1y7Lpoib4fsUoiK4PP/XCfKqKL1Ek+417c
PGtSL4PY3cnDpB4v5TcE4f4YRvWxBcJq8kfWfO2x4GT9QhVhU/Gw7MS0Xe2LCQxhQCc4XtNyoOaW
tVCmjMa0o5KwALwo1W92hyLl9lKKQbksVA0kRVNvi8T1BUytm5CjtoElnhumFN3kVFtKhgsioasU
DaKQGyBtEvRhd4bpF/ZuQs+vDXTxkTOCLGvJjAaKw3+/JmYrs55EGElcHPvfg3LAn6EnfCvE/a5/
0B9xpJA0E6NTE3fCa4RPgm2o08XpLtYWPs9DB/+InvJfEYHeWuxoRitxgpVqh5qz/S4w0IaFDaaY
X9eTg0e6hh7TuuTjRPdYGSWqq0TyJHEoykYGRQEW0wuT1f7ywrZpApcK0e4pzMW6RzGBbTGDIW9I
A2QFym5qmwTeGWwZfjM7tb0RyY8m+EkamkLBtd2qQTM/vGjeIfCMyZQwiVtKRy1sINJ+aiNeCQTC
94g7zHSLy7N8qIzoa2KMsnZICnPjOWn1mnxPIBepe4EiNTs0/Z83MJ+aP1Nyybr03saBdcFurCtH
CJiFp6mPdKjB/UihtYvBB9XW25hEDhTZYiObPYtSjcFKgOEyjejmOIhSqZADAcpBalu1bKahXFxI
c0EBRsXUzxwQoYeCkkLe7kyBBP+suCQZy1y6eUAbGJ4PgHADylRg/AwdJ9nXaOICViWZhBU/AKAr
0FPJkfb65kLdqgaKuuCHu3892UYJQm9k6AWFqALK9hNznp/ulipb5FpxHc/AMaE2x5JxdYakhDPL
f3ditpKMh4ArlHsYh4BrDLdl9Qc0txNTbjKW+bgFjtLVX+6ytpFnWQmj8QieBF6QQSJ3btqHOrNU
pXnhNu/yztd8kfRf899xRodjb4sLKbQV8RHMUiPWoav3KbxzmOaRLuUUg55tJ2mZBBHkKrGbxFNB
JyRpTTr2gfver/3am8riQfgsm2R1GfqSi/G+SiSF9oy/fqV7JSAj2gJe+dxRtUYIb6zcLv7EPVQ3
tvUhz3J9RcM1pgZnlBXf6srb1e/aXASLuhx60K6gJSba258c6WlcsNLp+JQXj4MQi2HqEUN1iJQ9
eIsqE/G0L+iaS80hGzmU+Xg2aWERKIBz2rIjaQabxNPEvvoa4/NWPdQF09SNXSMvftNKKAAhRznu
N6W6hhN5MAT98KLLja709gKxMWAXOD7v1aNUP28StbRsZxPFiR4f3HtSfayvYT9WpGRZg8u3KOCq
EiEwI3h+ptapffaDOQ8k8rLTQP4QuwA4QVzoq4XcVcQO701IC2pWN2R9a0dCkcKjKUFhS4mZPqrh
g7/UmOM+XgM3IBavsbpSfsqyfODj6YR0WCkrG/+xs4H8I266FD/NXqEVqkNgJ1B8mcFs7mKuWJhy
DaxZrfium8lonld2079Lei1INGAEAGf8A7ljVLY/35tRwa/w72nPf1S9pO2WXpcb9DLyZtXQ5P18
6cYsM4VQYrjaPf0O2uwYWzhi81liSBU7EeGQU1grvxdNsQnSktoGd2MwQ9VVIJDfoM3gxrvu5JOu
deRqfmKjglxffWTH6MY+jS6XtUdcbFtga0tdw69H9/TfEWCl/FNI+gFzfKwml2y+kx7l9th0eJ9p
UDl751JYAgI3GVdQjuhCRRcXCnoRnMczP5zguXt7NfyIGrbEsp1+dEszC8kAFTFX9qz7uRQPo8IT
XvXhRznIRaAKMBYSJIaEiFAXPnxWt+FamQGBWzI+N6m3mPhjUqKFxxdW4edbsqHLwd9DNrQVnCpA
Ox0j2e0YT2ptTuVLva3Ct7HY4lMuBu1jfjWFXC1MWPfNPMjLzNgC3Ljv2pn/5zHRvYk7l7a5wMVY
w0F9G6GCCtPUIHd8y7msytO/lXDzzdfkDH8jtcYnylreQAflxRuF+Rqoe8dh3gmMOnXu4VGsEevz
/9aB8bo2jue/z0+HoxF7HswRZE12Y9HPOx1qDtFmhjRCkXPouosaooNrmtdIxfIgu1nl78HkakhB
rcIeLfjx9fz+3oEUfAbGH7HgjNfss7TBgJoH3T2OCcgMamdiZagVzCXWgbxJ9SGJl0jg5rNJXBvX
iZqnKGp3e3W/Ds60yrbu97ILfMFRhBAc3uip2EHtCIH6oBM1MddtUjOHSZdzp6K9uQASdAan6BP2
ewxmhod9tas+i57Zb1FeuppgBqbdXlaDLsKHfTluTIs7btbUGG0ie6ssACuRpa13kyGm9OVjrguJ
Zz8tj07y0bv+ino54Q3rnvB6KvwX9GOO0WK0jyGcEWdyYc9kOG//2a8AXj4XCiBqXJxH8dbRW7rn
9fGSn7KlpOiuYN4bqHaZZoRWbGaD45FuVl586PS42pU5n8ilPlUUFbQ/vEwsGMA7gHEDjHgA5IkY
9gjv++RvZTq9MWE1u/bZWzr47ssCxoOpWBQO4sZzRYQ8yepQWbK9lXTlZf5hENrpnOGIoEdPvVDp
s8ZberGwpNrhky6MW0dgOmajzJbTHHUdGyO3YGHaL1tufo6++5WywcsGZiWWVjBbfMamZBxIl8yI
4NytY201JVc2W18kywWys9yYVZwkmMerPnSwaqcaIY9DzhsATsisMOvlxW5C4T9I8sOgK7knUf4K
LoT8vkqogTn8HCYvoysTiPZzatlC4pAM7e8s2Gw0L1iGmQivYlcfWsy9FMn6W6GZYFIGZ8OzmRIX
RL5E7zRB1zytu+Tdbxyb2dGPujJdamp7CY6350QtuQ8k7Th3LniGt+9+09+H3LvTond3u+akXQE6
ihLHkZIWYtFPfGSNacTjM+WsbiHnC8aGR5csYn/hj8b1ZgZcCMZ3ZPa/Q3mSYUMclNCzLksPKz7z
2xhTA9/6Zk9y2biASOyoxMPC5smNDAwg5UyTe+FpGMF4EumNKmasjH3+Lpdz7noYN+a2NWPxzE9/
nJJXO6o3Tbzri17OxHnKUKOT2264amqqKxZS++fs/1s9eLbthkEQrIFqnYyzQh7VCJS8LsR+9LXW
EsMgO6t0M5ubTmx1ot44HZl7UFpo546V3Aa5aiC88RgSzCADgEcu2eA9Lviq6NJp96E8yYFNO28H
nx4cZjcc1vOK4g13zStBlXI62CMzOs4pWoYNVf5rmbvUEzjZLFLRr9MFh0zx9ZC1Wn+fedtBkQ92
WaamNUntSBXojlOvfFmqOxdxpeSMtBTCChRCh3anOPkfYK0m5wJMTvbjToL0Q1RgPv4igsMgwKVr
MMM67uk0KOhykK8NylZxNl39SJGAxgYN+R15XTZBdm1i1ztA9PJT+r+p/vT+gH320PZCOc3TwbSY
zJMbUt40exRrgmm8zf8bG56KUxwQ7CFGPUrQ/H5hJbkdMtoBZ7XuzZyplbkXKPSWXNe1w/DfpS6G
drB3S+G6FbPbk9P8jI9EABpwVyBNwik7vYfbEZhX3mpQx+Weiq/iHFiJpOHbVuytyoWgvV6lR6j3
SzC4FFdWZXRuoQno7krmlKwHpCe5RV1fOir8n4RjOt84L5oOpsEwNN+NRNgveSZB9kRgL1MnN5Rl
VFZS6pEL2sDCN+GP7J9O4S/YQjytz+U3EZ3wxetqLC3CyFtliTXHM4KHwo4Smhwmdd2kMV4oZI5f
OaZ7ALMQnKxedCP8HlEhCUjyKiuhiX2A4pZYaY7Ha10UJEZp+x6dLbIAjCgIeuouh++zAGDdHAaq
EXI174Tq+2foNi6Gmaao/ve2h7qQCY326pixLAdWl7HyXF/tPXiUeH/7GpVbrV4WjXdJ276Rzw3N
6z20Dl9YsynPqh6018NMYN8lUZzb2dT/5IaO7O/VhG35Nf4YdmYF7Ne4gkLKPFr0BrPLrEMzCAW9
lLuxiBK7jAnVS8W47/JQ4tTEw8wdf9mavv58hlOk1xirE8t72JM38XIC1QBjGpJib3b3bbRLkrgP
jc+dMJIGU+LNk+28/U5n2lbk61T30156htluRWaXqARuzFNL8fbJW2hqwsMavCsFi3mw0rlIx8Dl
OU8HhoQ05qS5aCR/dgShibwW152c9NupknuRgpMCP7baeaR+bxegzwVmplTFmGqt191Gfo+j5hRL
Q8975eK5WeTMlqc2BvcdMToqfYwmH4tN/EYQjIzBQty/PRB5NT9Zs/YNfOrU3ylazKYxLwQRRcqo
eV5BUyY3WTlUXYkusrqZMK8sqTCvDPEgduiAkPuxJ+HUevkrrgl4KJViSEP6saqUaB+Cs0sit6IK
B2/1EAYjCkJm/4ywKEqQVmD2/MT1r20sLk8Cyuu+l6kfUY1eUEdZhSsAWECeUu4GXgaLt+Uhg4xb
hIbm+3Ip90k/kdrTUJEgErWHjfDA0dtYBvWqAoFRlE73fgdYSz5j3Mo0OEf8HNh0rMSAcac6gsIW
BLFUZfLLbLy5cTCUW9Or8X/Zy6bplLLtCT79nFhTUhCfZAmwU8BgfyozgRNyjn5BIeKOg+Qx7APv
p0NJVF/0PbEgJFOPm4IL09onzL/IrzQttaTkt17F9pZvdTDBDG5iHSk3pPAR+kJgFa+UKDi65fBD
PSi1DYxkZ82Xzf2JapjLOzYDZphKYPrTK2FQ1684SVwgOkyKJl6ufIe2dt5sbmKeedlTxgjDvCfY
483CF9ARaL145dST7SgUVLVeOSWdEJJYveGbDFgOTvoAUElGvlzUMm7gecGIy/jy056Oacx5xM7H
D98ZhpG57WCuwz07vjaqwY2azYQt0UPM3IGZYPeHSiva+JLKWMBQDOfi5x8EjueiSjRKBJ484rDc
yVOyeZ7+h366CQdpj37KhASQMJ+mfmvhGA/2mRo3lK+2a2Arc66WtW18j8APqlkB/ENASGBkBIcn
OwHH4Sc8DJ27p0wGmMyzZ5cC3T8d0JfNsEnoS0UeQsC5E3JdZX4L/VyEUi+3+rauciZVu+XW/qhF
rpIKMmtx16379M1YnanvcQDrqzNU2ofhMu4BnGKshaQ5HH09i9womBf0OmwunCFc1Hiz1Fb/pO0a
j9iZdeJoavSIr+7a17SeZmrkvPLjnhAwnyn62xdDg6J9W5VmleR+PvX22lrea8lUkXEkJqjgPA/1
QqGL9G6euuQlSstY8PmFQTYcDS6947/igimBlmTNPTDVeCrGtueptvIz09ckB4/UvusG2Knk/LT/
6dia6yOgSKfJG1pUtzhWp6LfHCzC24P6GG1uJzgHbDTrIZTMI/MfNr/2sDbn6owsfEES1z+7d2D2
rbqIm+x5gzOxTatfJI+gqjFswF/HhJoPNDURhIwqA+L6Npwx44nlZYIYbsBLWnTomNlqgltrKOyL
buDZLp8iqSzQXVWviGBxDhhKyjKuZeTuWab9SIKrj3s6jRvUgj7UoIysww6c96iOVDbhNvzDu0SO
1yhRQwosgkhRsv4QzhiUp08wbUTDx2jqxN9JeP2vxMLO4Wj9i2GZXPfKs3cbfVj96WMLBGllR6Yu
4ar6b0UQziVJAs8yhLEFch/u/nvnk6NA2I0euG5j9vxcZkArMnT8TXYHqKpSafsWikCVJ0qNCLSk
MFKInAZTp6SCbPOJB3xkQzRPDM1hM3WeEifUmvs/Uhad9mKdlSUEyWvu7MrmpcWT5exeOKZlfSaf
duzFse7dLFC1ioYjpZX2Vh83qJMv3Op2brRwYOLsLJH1wSkITR0KtzBUloT5rVmexF3WmGznrJS5
4spIjvWVg6WiTXESe96/r+2Cxi3WrD75ZAnD0IRIuMv4C6qDZlrGtfNQvdDQTPFLxiKn3zSzvma2
8XDYohuWiUohL54EBYP2Zko4QlzyueGQQsTUfDovnlaAAqzGA2ut1aSXbJ7PrHrU5IT3gnQkrcLX
sohLlN7pT/BydQ/ZlWe+oZXk7pMMQsiEq9SBYLvaIrl9ME6r+3bhiQwuWyDiKALRQVbqnt3ffjtj
OLPNZjzshlSZlkztKjSPmue1epHb8RuNjcA94LPdgmsVmSucp0ATammDpzGXz5yg2tbHyPLh+hUg
pglvBhNL8aNUFlBqiiEtMB8QUsaH38g1M+2ucMpggR3tlLRrARuvfjW7grz2WbmcpkjYGvB6HRYA
PsZOqbqaGjoy2QA7EDIZjlmFKnes9IJ8HBC/Y82fqwNjq7JU6s42tFJEHeFmDV0x7abFiv2EZmLy
IvB1FtFPjgk0XZedj1sjhVstRXc9tCnRmJF4a2DXjQ3Qu4tDzEMhEXkITz4Y93Rec9yrtDPYdd4S
chsfXHJZf3p48BN9F83rq1zRTf6WFXHIOm68uCvWsT+kfOX0HGcvX0BIhg1SI2w7TU6ihp2vx41Q
4gYILeBXcWcUKIPv5DgQBaqR+1JHEr1DR4nW3bAcBqyNDeJVymKfGUaF7ejH0/mz8964keim5yk2
CSro9YoAmQDxCQFTNucG4P+IXRhWl2HKml0czUf0aDabCnaLjZUH3dmRJLS7T9mQiEeJAPoRy0w4
yJLhwN3fsVRj6CeIG8EYPJ5tc1IWYQzJhLWbaZ9eYSVWU4KPQHMPB350ly22VKYsFZ2JiI+6JQP5
D8OGh5Ilo680aY7Z1U//a6LKhuXxthzwxQUqrxUiOqSseBO5x+eP505OjJieGlWMn1BEHk+GTMsM
YyFFzm69u1h2dIx4wu2nXzrYiinaHF0VTZky8sb7P4vgsnItlk00sCcIvCyUAz37Vbunv2evQhV0
Wp+gONIqj/fFEr6Z4HPnjPBCnf6sSL/x7o5DuVlNyEOUH0M720NRGDAZs7q9X82RQgWHT6TJAIPX
QJXvw/JGU3hiT6u1wUnIdnU6ZgYv9xB07xuhUVjVqsOET7gqHcl+5bsHyjEuC9hXkkqeqrdmnFsa
c8Bfcf0BCujGI08O0e3q9bMfUX8q6p3F+iuS1eZmrudgJdMGKIJcvbJ6enFF8VXVqZhazp+YZDcj
xy33P7c65v9uz+n8ZGiGIRP1IyoTWXeUYGVA0oYeQnkFt7jv8yXSqaXHjvCw9651loWY6h3ZAYCD
rWjMZnNFBP9CuYIcq0GjQuBOAWSRrAu2jOOhF1F8jnaeQPEVYpjGHWQDNfbOITvZXFOoH42jU06K
g68SvEQy+BIl0PxFG/s2ZCoGStC1AZGgnpJgRMIGuRXmcRgXl54ZR07WWOFt4afQnagyzZbU+4Wx
upCpdGmG0tuP2G2OrJNmOHeZMriztf2uzFnibkDZy7/zRiC0Ed4WgvXxREgjFYXg9hYY/LvOVT4A
QwTzjjtT6JorEipR/GDmVdqVNFGMoRJfMu0P1TaumuAtLuHsDWpJnq7PP090t5t+UAuY+ZSiM5Mq
u+J30cHsI9GlHLOPqoCVmmAjuE/56yiVsI6Wj7GIbe4iZrIbbwRf9S9iBvz1V4RFxn5Eh/g/2LVg
zm4P9w8AUfAplZcpLD3oCmk2aqvbteemmzulGdEionlKzKFOfzXbDrSGo6aK40bi5Cqfm+6EfVXU
l4o/YUsOmRm7s2yJZmnXnhh5L93lmP83TCup5rG9GWsdaGCZEvZxNYfpjLF8PVLWj1VdXNZRnHh1
kpxp/Nlln66X33pXQTOpa/wMhdQBtNtMgjsH7n/0DYRDU82ut1t+Io7jCzQCXz/IE4m/SbZgfVps
1ZOJrdkq486a0PWFQC0+cYyQB9oXd+b7yOg0CJUwLEJXEhlJ5uSf0UE9z/9eiDDK80lHCoCxquCB
IunGuYAMsdtRuqHYpCVqXATxihNef358zCV499q/uWoTssIuwZAzVu5UuSfV8yhLTorPhlvx4RW0
dlZUAfLrwQqS2xTrzlpqtfgKoeI3+Hq3OlhuZXvXyqDODJfB79M9M5tk+z/UaYJ+sFHbKtw6oHMV
wRiHaGY02DryOtaYKcpPp7dZGPMqqBZimefB40l3WnhV8qoo+Z6pgVgZJM+fVpj5pF/Wx5jtlrWe
T4M1aEJMQLtWLDMrxsi5Kj1sPHdNKuNIVLu1smmNNkbStJ+RV/mXs1EAII+2W83mudNWD+sQ+7H5
5/y305rwAritSncvxeFsS4FqYyEMes5I8gx6CV9O9teUF0hh78enOUWQKuDDtb5IMeYqxcKNJ7Hr
y84tqRsJvu7edQK2Kuuz7woUHcV4bpbS/7ImHwUyjeNb4eTmZWn3EHYnUypk7xckYohGENNkoQhK
UIqIq/xy9CgtFqiBzv18kDFe7AF7aQiTxVuCQX1rGD7WwbDZs60ptisqem5OKMTvXQTaPiOcN3PA
c3MmPn514xUG9wgxtkfBlGMEOJ+47WpshGiW/531s6PZSY+qK/PcxVhBY1Svy75oXk4uEKtAfIQA
Uld3NqM787gP1E+o/EvaJSdcGb7CeUlWjrpQoymnOJwFtdofTtLW6rUVBkjpBX9xjnWkJKrn6gDi
ablOa56nyZEcQuooqzUAEAXbKE5gsTT8P5aqIGv9QpxRMRHI9l4izJ1tzoy8d3rr7dT6uHzlqdAd
R4kRRPOvsgAexwzZdOMzn6cEN9ciV1IHTjmiZjop8RB4170J4Loro221AEntyAolTGCdoooQq6JO
YUEzSv7P9R1t20SiI2RvfUH5tk0WEvKeMHxCAdyZhOIrhhii/v5dTikGzf8+7kVxw48fAdW1lEuS
jE/Y5Ho0KNeta9acCXgp6WXDv7OhN7ciA2viYvOzSFLQTq4QXvSottu4b0ikKhvuBvfh14u2RU1B
OX54JfT7V/BHZ/aUOAlcW5Lf3EU6buF2CD8MooiVNKq2UCdSM2nKQOf14D+wYz/cTDBRezhYUGiX
FhJ26FLTt6LHW417zuNTTm9jQRujT/CB84E3fZDVvVEiiLvnNOMwlINJSsklb64Npv8xt3Ox+w/e
9al0ZerU0y1OMBxRWObN8n6v2TbFc9/HRYwEm9+jnVvxtTQ3Kb80GnS/v/+buVsIO27ISx0N3xSz
0k0EuMyRbxBSozQV8W/GPaX0TiS9ROzxJKoI5PONMD30oEtPf8ql2Lv3zePeigw5qSaRW+FlDDr2
Di4hsJXo/qnoYqH2PN9AtC31Os3nQxPPKqz05uZsgyB/aMdzsSSTZvXqfwzfgESNd75Hr1n3G4gC
y97foeCXZBSsfYFeUlxpThCwW2V8Ldd+cQWzNZw92XjVjKLubpAlT901ZmY7RWAHixRJb+z4yZa2
eHjYtblqnInmvxAuL2XE2pd9V10nl0OIOhPVhqniV2n7Dat7Ukm0jQr+IgardBbcP7ibY8oTn2ms
GSBdcBF6+u7wnFvTCb7vXAMntJaPaOU0WvBkMyyf7yo9IFo5NU9rHR1jESchXkehvyqVDyjCdm0u
Zu5ZfVlYni+/o8OZ+QWTlcLis07oRjD1wBvbchi29rzZDfsEiJjnDw4fI5X8fAPXbjC0VPAawZDg
+BAna7gdq0n5rNcLoHRm8Gs9RVh74XSKpIG/EvcGeQFGst+wpNfTEQUzHPuZ/MVMsUwloacVjz33
n2/Ck0UEDlwBqinP6QOrO7pMgHgEPAZhQHV0zVE94GTlbufYCY+lBKHGIBiaZgrOv9EpOSg+dBiP
s5iFqd/Acj7tDP73esTA9uD3BfsZzXovR6O505htOK2QpGVODlAECEykZySjmBujqBgaRK6TqN2L
ksD8NLVxFU68NofKKZB2q6ZEW/Tye903cIpF9uXgUpeGWWmMEOktenKTICnRUopHiobqI1htW+eL
9KYYrKzKkpc5MwlUkZ1YV7YVjvZMgASYKn5ZQAxS8/o9fEPxMN4MCZa99jY0r2NmBiFX6EdlMyYd
Kwz4wsX7fXZEWEqfRYELkmiyfYoGZNl5ScsHZzsCh5axAwBUK1ck4N/p+4MPRcoPXyi8XzN741wO
C3FX5EKHawO6g2gYLwxvKsfQJqjOWykz52UlF7JYWJn400iw1+oUxW8itACE5zNmvX5lWgAczGsK
WenPhO9qkvDzHFof5nwR3s26DlY4JAVuNHaZZhznSXw1BPYu2awK7HaL30I/sfYjaCkbcmoOM+ig
3jJpZ59uNxpsmFCXeOPnI9TqhHuDYDnwKGJCG1KvXBsKvNcI1VBkXBFGC/MFDktWp88clyUzZnra
VcExx2wB8nbL9DV2fbWx+9V8xUIDq04LlYWEl9pYtypYf4f4+EeYDni4m+ZdVnMma9oAlmyc5ULd
ZwOS5MHFkovzWymIJ6Uu7AThgtR9fRh1KXRNM9+pAp85qCIy0AV95FVBXiKLsNq0RjQjc+hqzmyT
vCSwLKEeiWlreEXVTpHZMrBE2/u8DdAcESSWn0jdeAlkEIuk9EEzobcttV1ZziS3KX1bHx3T9jkH
OZimKhqfcnDPqLafR4dUOVtcfu6ps+43/qGH4BmgGv/Chvo1LRZqFldMKhR0rDjRgifyPItvzLtR
5E6aZmxcfUfOx2/EXGGOFItTaDfMoqhMraNzNMRrkAr/UalnueOc9Pek9+3P0OwE2k5PDusplwoA
k6uNp7VK+ESLKFR5rNyy7cAFrMMzF/OPp4aWFCLXZIpiL+YM17pZbPjGLYWm+zvq65voy4j3oIs5
FaVb/kqGg6lF6b0Te8CswNIu6EYBQBrMzCMSX8APAEN85LARR/ISrIvT7UDZZyOVGEUx6hQ74IQc
rM+6Xoq6qch3ZDnGKLgrOs5PVzMwpK2/NwjkUOysbO0CVmd5icuTcR/+3DcfUDIRlyoK4FCFmYvA
+6TKC/DBHPyGMyCBNMCLjsFCI0Jmlxtp4sICVGrKzgHNg79v7/wCj4bl6IB9TaaIHwGXYVeBZ9Hf
kqitrmqtYvNhd2GM2JxLQZQhwzRemMMMNHLyqwQSLkvan/HtJxBwOuEOmdHn1roBHSAghoj+hixv
wDOqpLz8IrpS08vvyH8mmeE9ECi5fHs6DGOviAnqIKAIvBdo+9AfpwOf60gDUIi8JJBL7X2KFYQO
6GnzZumtPTJeJ8sf7VqHvru+sZYsIImzpfigjqJF6xwpobO+VjDTMETntWIlk3G/HKuGEYIlP945
iR182eHzO2iDDeBvg49l35/4jOpF0Qr8CbriY8XJEurSFp6rLfqj6p5cAgpBDtdgWBifW1Sxufe3
uajCOOYu3qUqwFQkM29fWoOD/fZ6/5NuW2kjEbyMom6M8snQWAVogf+8r67E0q6Zy84b844+dptH
IPxeA6PW6yGjkayTOaVBO8lBrlsBIkoq7xFxOhiMbZLyNteJpAvVWqdT1jZM4UY9J4wCYNcjB2v7
q+6dwQb+W1VXiUfIC3Tkr8VueABNHit/3m7FzrrelYbf1YNERfp1ez2PtkZxLuYLynDvi1n9R8xH
CbQAxJ1kQikLT27+vMiS23xrOC6RJy2qovUe0H1kYF8678G5qW4vhHCjByp+tto/NxIyqHoqdObE
9ULHXVVwPJGKfOdrJ8Ot9pDJY/lGJkuJJS75S8ps4fW0KsqRxOlTi/pwWpkDf9Y+MLfEwJ/QNYQ2
ih8LtqwKNytkYb8ywRS++ijV9Rd4j8PQ/F/hY7+GND0UK6rmob3c3nSdEIcL7gW2fv9TO79WvqGQ
HcijJxmXXUtpXB1zZvxCsMedHHbbL/tm1Pxactu7KeXzHEen/Ehk5u71/5WobY5Z/ntLByHlZkpm
Wc3eqF1qlwpN6JtF26/8BNiZ2bhlh2xlIgHmdZmO6w6X0Lcx4L64FHGaHGnY+YNcGnUWV1Er0eD+
s4jUrPurs8lNSoSepRMUbVf2IthtOJf1u3tMjdmsSLfwH0d7PolZgxBgSgeB/ZUQBbyy4o9lUWfG
9cHzTDW4HZQutaSI+Hbv+JbaKLxGr1zEractnbXjQsiTFmSUk6WuLeSmACl0mR7aAVFFSoRl0XU/
TsvsE+0qh51WsWnwZ+a19x5CcBdC1/xRnJQ17FpAvOXTuVwZcepLSN+upRQIy0+ikYp3m+yoGLo9
vYEogv5j9taEqiHi1hvaY3Fcb74oPaPFv2qAbrL8vC7NGV+tvj0jwzR0JvErnRFrWRJE/NaSBXWk
KMk3A9tGLNLIXX9MTfVW/xZ4W3gvEpkrMyWAo4BUEhKBVyDhVg9nk0as+iNcZ4YZ6nqEn2Ly4UWS
qcsxE53z+G84snNLgFCzogkal/KfbSoYLxx+bf1/Shl6pvFxOxQ9N3Ipm6YE63X2fc7UV7BdJX9w
acIHwmXfxqsdz+UiRS7kANyVA3Qbz7t0yC88pyXaeCEBdKAh7GjfW+Oak5OIhuUciAGYAG29e4L4
o3kpAo8wVcbm24dW8sPrH/kyJSKMX9QYQS4ad1vqcAn+Z8gvwX5KCqW0VbIm1vG7ltiElKM+ZDna
EM1JLUehJsOQWByFBNoocWsxibnTybSyxH5K5h5IcsIYwKsomxkrb0HTCfQCkcZeFFvx8tQ3ar29
qsEapckjSgSqAhI7Y/Wm3PDkLg1rlb+WJg17s9u5j2nqewMyPjirRDfz2TQLYfAU54xWwTLLvpjq
BgxEic7Crz1VXG4zaIyqSO0AQwgG4mntefgrTNz6WopRq7Pg/JYmB6XPxzWQFJMc/LI+/zv6v4Ei
mnsx510crXU0ht8O3WrvRB+AFEL2/QtcmctE+t2nAm3rMn/t9ipNJmkHyPr+zz7LL7ucVtQL5ko3
39XJfVoJao6i8dMmSYKO2SsP5Jvthe1bndWOpoHCP+MFDgCd/cBPENoPmh5kNjAuVj3zucqPXRYj
GrNEQfBtT6/SUxFkoUe1i0vlNJ5vDXRbbIcXGDk4B48pod96C3PbX1v4DtlT3D0P20ozqaTHTv8J
6BficVjXzYjXBGLTS7O5F0KkLXZZz6gwtp88PYVM1YjJAeIAVxMzRytpXEUgh4bhFXbOJ/uaxXvf
5nwTbQ6CxG57Mz4GzcGF0e0yZs7yzixcXz7uFn5RJP+pocbCMeNsbb83IEvM5bdwE73ITUj2BG8Z
pugFG+yZ+YJLGrZkPbRsmeuB/RMb2CdAiB+wqceEy4cQPuFZB8WDSRLGuGGgpj0lPGxwd0TCydDc
qhPK7zJcyKhldR22Dd0CJLZAcDi1GM+gTRpqNLOLQ/cN/A0LYkoxENlfqHnNmE21QShiuzCIqTl0
V5qrLRgMpAnMfX08/H5o+xaOhhh3TISHV6p3djbJow2lekH9NHYnB/vDeyGsMl/pJQaBOdjDxiGL
DARhjqS6htpB5lBwRwTrZqDCHioFKdvcFqVLizU80GwkYbVWY7Bz3EZuN4ZGc82m49nao+S9jDNj
/MKKD+PnpRQDP5Zq1bQfS/ZNKvyeITfdClEds7lG2/Ai9Xdvza3g1NZ/2Hf6Jq/48A59YtqhjnSk
k6T1wy43heMlXlRC9G82TVHqvK410NMO5IxkBGiMrFELaUGu2Gkn8wxlvR5hmVClZ62UXKt6Pwv3
AeSQxG0aRdwh7cw6nv/bC+iGjNIWWEVtSWYZYfpgJUvtEsd8AkBrcEBzOI7ZFbYbuj6qwrluJzyP
frGvO/k8e+MSpoSDpSBIN7VRN4LvFYApYgBVc5BAsQD21c0cJRmUrFZFqM4DEjguYC7+uF0O47Rn
XP0xgtqh7Z3uBTdFI2LJ6NHhQrIn9g+x0KuQdTPzNHh0qW9H1yS/oMoz8PcZlD1FtgpfP32423M+
SJgOBWAAb77FnEM5i+DrTghu+Q6ydNMW6b40yMFZUvv4VT2WwDbi05/oATzgg2jGxTC2sux8z/tt
ThMChJz42XP1Va4RgDg81yWfqqTW4Q4K6Yts2boZtdOXoFDkakcTvjYyKP84Om2GW+/AZYwxtZt8
pSZezuXqrVq1NMamOfFYLRLWAJ9+K6YMhE76DoL1wEt0XqtkyXiuNQoxjuLQjitEl4d/LT5b0ELG
gvtjbOJ1uQgdyC19WuzXM2QKkeEnFa6aek3MhwbhE1yP5DchlcY8Lp5I0lUeyIG2eyypRoVyLFZQ
YVxvPS/RYMUD+DRJO+Gd5GzrMAU6pnm+zREP8IlqcMEpRoJVqkrpdCx6geC/giitZ7MJTijR5ovo
tD9A62TMnJ5VMkZ/yYVju3rL6ISV7pdzS3Dq1UghvMVpNC4Jl8sRgQoLg28MUG63CUOg5QDDJT1L
nFjhlmpwPXeHMmHnbmJRSHXKc84IcUsJUYdEEJ+QFm2mEHibQ0qIjz75tbtA1x7tDaWh5Ea9TWzj
jjg72AiogdykcAnnbNxVSamdJcm2DTmPMQt25GRW2mpTyl4Lezhxgk8iaiXJfykbKNSNCMbnBapk
yrH4D3LmKzq9HEuG+quv9kcbxaFqEfb8hZLXIYiUpuHhIKTWqWdKnUTb7P0WwHu0/2RIs4EgaDKr
IiFBqzV6R+GRZRGziD7JTMJpp4wWlCrKlpTKDp+rGD0L20ju9gBkeccF5sqD7DzCJEyzSLV0Mv+p
LFZHZtBFlzYFoZ1PMD6ELq/GNwJhAkRdUGG42fDIdgd68691QXTYMGPhM8z7Et9w2+DttOxFaiEV
fkj6gRya1F4wUG6WYxYAE7bOdaZLKihd4NHOh3f3Wsk9vPHcyvT6T7cmuFkED0Q3tyEdY97FViCW
c1x2YT1bf7Dslx/ipvk+0tUcUy+s0Iy5GaOb76MzS8aDpSnA74QryxrodoiGgTu9kNf3OKBYYjpj
kuXuaDmqiBrjP93F/FgLpjXp7+qZFS13/hW1Ljhy/X/FdWLDBEP/ed6FVoPox2v5HQ2NGJZAcBI6
gsMAZ1SHP8xgR0ECI8qVGJKF8gAK3z7VTZdTUL/C5js3E69We70mw5aJDYgXER6Yy3vkMHA08v16
0S4A6WcBFDGx3nVrSCG8fSZ3+BcqZ9JvruYp7H5P0UyzTZfCKXr3WDLyEAtB3UTd89ncIUcviCB3
XCKtqo0p6SAHW7BmwlpUEdaXa6EalGJl5KLF5Svem9SRO//UPrX9GjA/Cc/9ykAf465tG0g7EEaI
MnbYo/fKr2Z80DJCVwVLf/cvbaAlsy/mLe5uG9XSEhREy9z1dyabqaddG0IY0mK+bD8bTkuhU66D
ND1VZnSYrkArcKTAqHkaBxLbKZym0eXbYxmmZErKQhJsJys7JlH9OmfSGloVa3q8147V1tTeDpAb
NoEij4b3cl8bGm33OlesoQhM1OGk18jvnOy/PmNUWQPdPu0DXV6yxm2psjQPtizUyupHQ9Cb2AtM
9jPR2WdvOB6TMI6A2LFNecJLzhRJajEVNLG6qvUIzpUZp9KTDx5DxR7BhvmpJqNkQZCMYd4HTFIs
sPXW9ntYXNWZzUiXw4uvc0HZl+lYKYJQdJGtEsxV2wDHmzvOZn1bS3u9wGYb+hpEsa9wsPo7ioux
8yzwLDX7H6dGl1BX3iIHhkjVcniPhXzcZYkbAFtemK5810e6ITIk1XICabd11w09nIoDEK4r8ffT
ddhWLzOufbjpkjtHVQDj8paeJbs7lEndn81jwlUhPhXF/+gpwHt9/E/gNPk1lQyy3F9+CIWpaRFC
k6WDlt5VXDsReYAXgHGkekXKBU5vQ/cLJpsIjXvofZV6iFMdpgkQRhpu2GckvTZ09lwOS8ss/Npb
2hKf4whEhl884SXbxYqFZiXZFCb1kuBfXJTZD4vCeZmco8CnG5nl8e57o0svZo2hbVNfpB8+6N0F
RtEtDeFoS2Oyv4z7KavlqWK9TA5hxi9NBn5QjX6MBEeoD/AZacTFbRNls7JoU8Gw7adohEUM4qtb
Y7jtUta4l3jv6UGB0ZfkQpCQrREpRqjtSPPIoCicLb+1JusDy65cyWjhZNlaz4e1aNNKsEJe2Iuu
fDpfMMIeAyZPwlugViGqIC56Jy8IAa5HP7yLTmIsC5Xqzej9Vj3WdNmgBHig4z7Gr+9KfycEDlBD
kzjxVUp9eQf+uoQCQQhU0IFJ3L6N5i5hP/gdJSr12+7kuWcAFCQftT5l2Al80LlCV2l9d9jK57Ct
0g0m/01qWJNZuOFoz2gxpM4Ih5ZPeP+cUOrUGe9rccKQ8TuJB4OXyVRuFvTxhoL9mcTGjnF6/+JB
Ah66Q2vMU4g2DKENz4PYqrukjm5ImiF70dQmLIEwx7J3WAWcZAzUvYViIOaOjkhj8NIKGWLxqNB1
yxwZqJ7RZ7xu8iIeSUd0FskHcNyuABqc0I3/wTMsG2hC7i3Pa4Jupbo1xsyGVEG37pYV/tDacxjl
otTt3YoM7ocn2FGEi2VWYQ9oneFVBmOFIAlFu6M0OpgbvGfu8y16ldYgzcmrM6JP7DGIEgclv+Em
Hz6P2cedMDnoGMPbO6lmDSMZ5XuSgOTkQoag864lg1/4iFWHjSj2mCUaAfs/TNyhioo8b6Jtt19M
/EjJfG4B2DIj6m6+1/QPPKlJke8F41PAf3je8oyxOiD8sDJnsB60em6JGw19m6uCDZEwZ3QEjTE6
6jqpKzZiCVc/j3lSwBAiRLHbdnOrbNU7e1E8MUSowTqfyTs6aRm0wIhS+CHz7u4A9a0Mw7Os/B0v
kv45AhYrZNMENCeOLt42VRQU+UV8/BByrDBq7vAE41lKoJK3t+6KcMVLRDYr7cpta3bMuQoQrTs8
gl+yVKHXIyjU9yi/prsSJu52dNA1u8NxpJs0IoHYPAHf053l5nsHPho9eLyzLxCLMhhbFewfHcf8
7RmdSIBpGYgjHG1968++IjdiYcfPgv5ZACgBHTdF5Tcy5CN9J7l9eia4vozqDXpgi/PNfqGRQRyw
0ZwnzoVg03RwctpkAjcIqEMG7AM1gboxgioKJwyQkvT06OoZoe6RK9rZAo8MKv39p4pDQG9LwB6T
OKC9RU3GZ98Fj6wv108AQDlHx7xE+c6RDzTHaCLCNu7q2E5BoaCPheRNntnORMT6GYWEkw8ycMc/
w7roO7zuMGA7tIurBaYiyRBRQ1betWvAl+AafFtAJuDTJ3vso6Zp6zREwG+GjzSTJ6i4dbaelpjD
0okxQat4YXmiiKviCh2MB4whqy/7wKn6MsMf5EudosPFLIdx1Yi25I7oQXl1/iEkxXJ1nwkQvEEb
9MJm12tnFNKAV+4LJferOVbejkrqrLTSmQO3kTPNL28lcE066Q7bN+KOmOOArQ3dIfmbTFiflrpk
e6THSo22pzktfYHZtetNMxgi6zI5hw/eIQYBywmTXx+FKjWp9yQSFHP8bWqJR55PtXb8piRO8uiK
igALAn2KNMXp8m2tC21/HnN4qIgZciAMMjTjn/8iiM4/fwHWPxpyndXykv592U1tWPG7jQKyVOK2
CbX6tX5mxyxCennpm9OcMyUTiUjpL5ghQTUHijnF8gi9thBb88eZ9P7H/QzyuzXiQrV6S0NAV6TI
uwjyX157NMCDqBdNFUs7VuAYi5GBWJmn0hciaieTkf2TeMmXtFhjifSsOKA6ULzsP5MEvNPtqjqq
E1Rvih53M3DIEFgamP1+/UruX2l9WMvsf9ZLvUN0gdjlhnAYxh2sKRee/+FcvPRXxiDqHN4t8mRa
rChqsSRb36ceOfqScOClGKbmeH88/SxZEOdLCGaOxOfpVB4F0w//ZKYHAyB7GTrjdjU3qYjRSlF+
wvWw0S6W6L/oIPUqoAsRdI5u3Ca1VKalL1yiUkLDc9oi2Nmw5b6+cMnkLlpzjN/MMNx4n4iIEqwo
CRg1+sHyDT9WIVDYcIWXIsjIDRVI9CGvOOKEKltV/bJRY5A/uhShWAExpVjRRLwHIO14iCAi52tC
ZEfgvYar8Fj0MwtC85j44vAd38bKMUCNQUg4SXUpXcQfe1igdgoYUPcdpEh1RQcp+H9C+R1M5eNh
z9Z7xQCYHJfFtqmeTExkjS9Pj/US5Hqkj8lRtDiKHYr6k+nn3sR/UfZGOtf6o6+7i42t29shGVYv
nAqJigyWiFbpDszzBcmp3YS6YdKZ+sBLMkgGqBVaN7f5ecr8hJeegmj8WW+kTaqEjAuJOLRC1M3C
9GSp9wW3GsgGu7gKVzzk7L/lYzNp6+vZoPI5h7+/O1rJ5wSp4VMBXJSvbvORkH0ZP/kA5qll+EGK
m6DdZ9mdaKdCmvwuNLL+r2jCmwEx3OR3bWtkW79QjuKXcZkR84fLAY+8PV1LAzyM5x0J0xx6qrJj
vZIvP8z8ErDVrCMtj8UpPG/7mFLYqqV+kKGZFEHIBh53AcXaXgzbY1EV1XxRLexM387ZPbNOIRN6
QwlZxhSDlv6PE7Cr+9JjID8OS7G/aXxKXBMmKVrLg68mtblXVti7ZvDOA03TR/pxzrS/ApwDEZpm
t+oxfz6BzeKvC9YBw36Y56gzN6HMVylUzIgBgcbjIVjz+3t9SuFNm3IMSn2Ccp8bxKQAih1dYmol
2MZqoRkM+Es/XDdoS5ZAPEWdv2VlqnJRV1TiY9jkrWhZqbJajfKAi7qgPQAyrHZt8c3redAOMHqK
l7A+xWfVlLMVB+cGnjkp63ksin+N1a03WovGEodb2jM5hmcx7rMDf5A/vPP3ggTdXTX96rJZNThS
X4Wr6fT4MShvYiZhOk8kG2uMm3mltpV8fdm2Hj6XtigvRCSTmHlQw6Xf2UAciABCztlNNLk36Vmf
J0foBhxK/H65TrhvBXj579YfTbf1mzwVJf26iWoczMcn14Xo3WHKYToNwj5+VePJwMQKy6Jx0OES
8aR2CA1IqgUxG/QkZ2HLMA9rzPwqLixHYeb54gaZ4aBwTDxkoBqxRwun+geQj6jErhfCnJxzQYss
gO3EJSPmj9quatA/H09XpGNFnHSn7ml+16b3Xby6wrhYxEce14A0TCs7p5NVWO8yjQJxXrY669JG
1/51LN2GEwwQyrn6AAhcoTmg5OP63A6pkqyJxgFg5Qwq2lRRm3P+EyOsGRp3aAYh3TNed9RkUiTs
SJqbtW1jG9dt2wY0hyH8RojiYy7z4gIsNCnKze6kSBFscKKgeeVPbRtSEukt/ZmxV6jH0rPZsH6g
oYF/fMQT2nDRG97uHJnBUuJY9/yiaO7LUXsbKp2eNkJCDWESR+yYyLag++Io7l8/21Yi+K1G1VdI
70JKog++/ZtruMa6z5pi9+blBw8v/ZRRK+VNrfazPW4pCC4VR7yxSh4BmWCYSy8aLGn5ZDoXpUEC
P+0FPln/OmJyCP6F9crQ32dh3gtty/ysCdjpnG+47nHNAF5QIG2jHhk/RXbzIGzPsXpdfCh3tjEu
l348ocpKJq49wUaKhlZRCioi+UVqsg+aHcfb1srO7Fo1Nyw8IdUjkiLVtvd+the8lvVvjc8gxAbV
vVu7iiniOLlyU9M16dbcpJ5cVECLjE5LVrvTnZUacOf4oKDQT+qGSEJ5qanHKYXyuvboAno5SmLc
i3JEP68WvkXVHNA9+7DF41Y8oNiJB1WiQsPhgO3XbjCnT/vGScRfMNZQVhqwoRCcP8Lx4W6IYCUX
jQwuSPSVkuGGKR3eqovu7K2KDfxWtfq6iHnB/tTSd+jZTC0XwHAw3JC8eo1M3yk4lRwsM2lE0M8k
DyoiGn4gCJu1lMJUFsgiIvs8oFlaHK3grK7XM0l+izKNhY3+nKD7p1BQQ8rLZkdgqUOq+2ZqRNkL
MtZhrPMi8kbo5JZQbMjiV8TBut8eKYG6jbw9rXFUpPkJty6IIJyX3bHkZ9piaWnjt3u1s/dAiz4a
ft5iaQbPm6SFMEJ4v1VAeeMJNtsbcuhHmKHNTT8b+isSlQjkAijrLACug4XhXhSbQvSpDQ65WMCr
D+ky9jXIZq3RPIM+Nr80hWS7T8ucpMRUWrasv9WbF2DLkNZxG17Nqp5oZVXTgV0C+uLnDk/vaQ08
hAq7oCQ+QjJqUPHXRoFW4rCTuGGabsQBat/ax/PEUiz6CZ+/IVCHNQIJ8QkQe1x2OaP2qLtFpj8G
Lq2R6AlrhD+Uhqz/rn70liO3QmpQQ5PBSFxm3yarIW6k+gtB5nJvI66oIeKqr/MHxH+4YSuuFPB1
1U4O/SmeT+4N2+z+VJxqSVXIdvKX5sbSPKvXaMVYCsghhWI9pSs1+hTp2gL10NlesOLKemlt6sk6
n++GdNdHBZrqvsLulozVgwTWAIrG09T3a8OnLsuw2delO63uo9ObmMTwXBwx5NXbw17aAfLBwM+s
ylXU0LGES4cOSGLfimPhJ0KHVcpgFEKORwpONlWKSr/4UE64fHk3SrkW2FGX3a/7mrHc/gD8/OQ7
rIcje068AQWapnt44B3CBZ15LbC/im/9fI42U6xtrKDeB23rY+W1cWGeFkI7vmGaRdKPZCtN0wap
WVcentU3isTVqoKgDt7oZ2Q9aUeuujIi30jJ1I7fGvamqvG8jnGloRq90RrrzYbGR4lCTtU85GQc
GSeSiuETT6rXb0socu61ozZyI7IN26OGiSHc8Cs7UrdMqWZrSqji3xyy5mCJwBtHvkb5sdT3yk8/
SrbcwcsfsAxEJT3/PVavomccCfUhHMAap92EjXHlf6mKg1ER0BuadfdQBOvTze/HQ/I5ESxeKwok
64NmJ0j0WcMr+bQTxdF4BXzoDzIpP3dypzQvZICN0e8X2vjgrI9I0xbOuLn9EXUg4HKiymnkuxk3
PwM0WZOFyIcb/wDEx1Lf2lsYStaWKaMc700Hfr987teBvru8BQVT2MN6CiOiCCnAPGWUGmfCtEix
M5oaHNsYKisWv6CCyXz435zOHKI8qfph/LNxojZJ42JJzVWruCDiO3u03p6kAc7rzRUD0fVqLYGn
xFtZ4YrbyDTrsDDLR84KXQ0183gbooc8LYcH5l/FO75P22GPLjN7dC7m/Ao4O8nfcZty+g3S8hwN
Tx1ThbNwYAPs/0sP15+UHm+TdtUl/nh2B2dpGYpP2HmZBiqYawKC6jskitxFvCQNaLfz0PQPaXCL
P8ezMSZUwPRyXrWJ6pOC/YidGXKL+VArUJEqK2Ejgkcqad55j0GJdtIOpFpg5o36qwJFx3mrlhrq
bTFCrSJtdWFUgtwuQXTe++ov9MejgJBTipJDRpxOGyLS1P6EzJ+Fn/g67kf8Lw2BG2bc7FFTqBv5
s/DaAcedVrad9knKpOytFGizae7KOuF912geYSul6+oewxyS8YUHuiWVnDnETYIVPIAbhC6itLzc
OxlNU/CKSP4Vy/9b0BX2uopqd7e1VAeq23NPv7hKRXDGMkY1LVMekKXHzicVoaUOe1YDXtAndO3X
OumfeapJVVpUAru61bIpqCkwdoM0sQnaSvxGgItoj375BWub3dmW1iKusM4aRfIvW3FuV0ZZEUqS
zKGpnjDZrK0GmH/DisMNMtBPiN5sSjwScCXmCv4BmxgqNeatobWOSrP6cvWBRwEmsB+C0NEVB47K
D5o2WAIHKNJm4RvehXHrYoeDMJFPtee05HpEOcACHZRgYWFijcUXvb96bD9h22LlR0/XqPZZnupR
sGvrNy3hbDKOqL7Ld29E7N/ulZM1rJ7hAr6aAf6Bmezl7HcYg3/R5E3BkqPSfedMIxNRklDHCeMR
cEx9me1zASjdxgCMw59XtW+W3IC1hcc5aVRzKNs5FMT+R8bSS3AxE/nyoEJjK3NuyzAxNDiVt3BE
lyKsKy5xnN7WlcajtX/wP/6VYVvfYyCcJE7kHPGhcFvgInCCwVjaFBVeQ5J48Lbl99mFRlzdYZFN
X2Rvk8JTenVDpNs2slcNA/LGvZAxsndQNrEzHalHknmCffnrRn0biylaXvkfQdoqmOO1ldgKc8Wk
NksVlDT5pAGKPJo1ucVz4PK1a+pHGMPjN/WYdFh0Q6IIL6adEV3aB7u+oK5JskXTcOmRSQN6379H
c2gi5LfeJ9QAqhRZix4RU1w5DQr9nMQJzCcftfxEgRlIzmIto51YGn7v+NiwMIXHormQWb6yAXPG
KSDgRtZP2V/IQ8CLX9ZQGS6eCK1lwW5P63b9mNLVFcVe2ihS7Luh6b4UwR//24dQDYhu4mMrOwEQ
Nu2/vr+IZbPl6gfCXAKbQKnYamdapcxV9oGMyrzIyIsZFT5eTtw+l3pHUbZZSmOOYjyhgD31T/8p
lomuMtqEBxvvGvSaAknhH4r1TbwTakfq61GUw+mi9xZUYJwlDxL/Qp5vPbU4RdllBU/OpL8Ge0g2
DZjlPn9GkJm+pM+K2pfK34wvDF0gfJFkmFgdeLXegrRSbQlZ5llskIqWOg4jUJxhsZIaplPAiMPj
4D5WnY1j07Ay6ODVHK6wJrnVxnjfRneaYp4ZX6IA1jSxQowCsaD09Mxk0LiXILVsWBxC1eOSFzrM
EHfn0i/vBV7ZVLxgUhievZQVCz5hAPikrLC2wig0H/xaMNZJHRDX3s0FOjF9eo6VlRdVYzniHvwm
CSCskk27XPqP1ZnfzjXwvmC6veylW4q2vgPxILdrWh3qYOEvsE6ijeHkuHpMtsvB1M7CLHHglT5K
QmEXMq0IhJHyONCySGuXpwTRtwuvsOpa94pbxX7dBzzZUGOdlia3PSuxgQRatZcPOEPUWIrordGr
xMwaX+mvH2qN4aKtlBP74DKei4zeezFmz7nNR1ObOLHwS61thVonScz2zJsNE/kj+huas2j0GnEh
uPc3kuv3edn9ZVrlgtK9Paqm4sxw8UEnMA9FWmqKkH1TCgidBDV//y2YtPOCVO0fkl65ww4upUqn
dr/Nw0ZPR/tz7+N5nw5K1hFJp/Spg1AeBA8NvSjByxoakiS88L3RUanV2uekaQD1z/lm7OZhAjeg
kIiAh3zZ1UukJdJhaiIiEIzDbBZRb8pmV6fYuvVEWjW7el0xYex3xygFT2jW1h1YKXzt8dhLWI7s
1qIK1FV2bmFnOjk3ZWeUmVU3OM35wPtPbS33CwD8TK2zuCgKL1o2fPu1vdxIM+NmLTL8/cv67/E1
wcs5U9ueEdH17eIyBvalUOpEpZ85qkp1FiCELFAJNMTAv50lKtgJGJL7VUK8BNcHcWPHaaAEgQLA
ESaAZFSDuXT/vjFFYf/TijmtSYIMxkXrrdUUNZRStq/Y7HBDRU8g7/ln/uuwaNsuKYTtEM5XZkCA
cPjWi5asRP9x6HdgsilQs9YAemMxhsfftG730LuxRVbX8BT7pErr3Id2sAe8nOTYx9c8xAKfYlET
o5/Vg501NH/hckiitVv/8aQ3PAn8BCcYlrmKjlCxpi4bPDLn/NbIfYpm8xZqCnPcUTxYA8+0pRhG
c1k1syUD4XGkv7U4NGUQJiSi1uiNjtbszISs78w85aGiU/OpD8J0pCOryPHTTCs0bP9lfCPQbgsD
ws5WTOmTgI3NCVZARTqvALx/lX2jEuB24ZFJ2+Qs4AsXOzAx5gU3yJ2/8+/ZJWJRESiIqxRn755R
esLFQLgPJWlnLqufUwiXXI11H5CsOBqNnd3dNJEFMRplAz0d7sktEnVmIlorjT/xhv548He4tXuR
zr9WCCaXXq9vb28Gn0bKXmFP5NhDKs9FJGPU0s0VIVn5iGhu7YVb4uiXG0pKsuF+cS51QWu00iqP
AmTRWexmwNbGZo0NREAwkiyj0cfDrr4iMJi700uZcBGiT12jU2xeoutd1+zAhJyrjKUqtN2ch/8c
95qVJxe2ruFuElVtJzSA8uv908939XQ53tb2l8KOoVrT4fVEKEZXykqLiZVIVWJ+LuLSKZw7kg1A
doFnsp1QlB7le+86Y1Rc/nxYcGm8+uUiHX950ssjxayb1e4nWBthywAyqeDPoH1GShonhYnATvVV
XjyGcbqQ1HmaA+iVMjPEeT6m0+o+m1BD74wFKsnD93ZsqiAUYCteItB2GnynjSZJg+1jvRho7H6U
ptAlgSj/sB0ZMSwhF65fdsMnNJRtnGDovWYZP7cAsNEGJiikCabyYKhjKhPx+Tb96tRnFqZFO/r6
tBLvw2UMDAjdW64I9w7ed4moIAqI1lOm254F01ZpnKyzhYnnb80YbwrQ7stWle6flB8rtqNWmKzo
2LD3vHhEaXrorX/hQOqOGevOeRPBToHhUY4qudsvsz6KbsJdLEQqcpn6vTFMN2a72O2i3lgjocOB
UYYQdmcYOvTPrUHLdcZYj/Y+8b6fBtvuYwQ6VkK4iWBqfuEorquTu1zL2oGGVX3GtFINKWjJW9FW
KUINbw7wO2ihc8CA3qDgX6cLmOeXsGldkvOD/y03OJJ+NrYZY10BaHJTtBajY7L3LJsolrfkQzQG
KxmbaWqiqV5Hm4s9c4lVPZ6Tj1xm+rFw86ZENmSIH2xjpPtcLMAjTvQlkIY7OKiYyH749B2tS1nl
45lKqORwx8P4sWOJZjnu+UVgcHMCXBxq80n8DxpXjB7zLmjzEZd8pMZT7OA9WQazauGZLf+FqrQ/
WoS0AxWw+HWqfL2NfOclTs6FiM8uvd0kaB5ikp99GR+9z12DU0qG7d3sErRinuyCfsdimTQ6BG0N
A1LdyQRWqoDMGAKmCXGOiJHJFD65adkrenlXvrnk9qwFlPBspu60nZeTmdMyr2fqmnkXSICJ01qW
fV2JqbYevvliVt02/Er43lqeCjRxUz8e9rZi8LGcNXIaJtH3PdaqhzoJ2xnJG7EV70msO5g7MCCO
XhN1oAZC8q9R7OEAGB+A5wJ3dsnKX5Kh9YyaaxyyV5kXAtdj5hj2MPbInSS9xvy4W+w6xanf02CA
7nB8tWKEojcCGy32igu1YJ14jiX8EtiABXJ/+S8WutMLYXdUBzZbkrWVl5AyFVHVN6zTmWZ4wsA1
hGmsqh4lfP7aLcPFn1JKfJHUOEnrJ4738D52k1AhVOME1CYn097vr+t7B8algDpEl+pqJcWRzTW5
829M6eBNvPAOcxnMhcW+DX5dlxTMZewV1Ur8c8RtZGeN5PknnMRdKO5t3nHNfs1A+xtzoCh4ZRtG
8nHCezq5kVcXnuSBv6EEpmLh7UDik3YnAfyWGHUPYwwcFfN2MSGieVCc89vJ6XlU7c5v5D4yGxc9
Fk5qcE8EL722H/2cQIsdr7nm2E/8DP+8Yp2UoG8SxDif8vtkXQA55TnTQuZBllGWUH0CNfMnjaNN
X2/dsmGF70B/p5m1fuV/Imxm1AouBN2p6Fuw2iGFxXtQQoibEquUlAMDHy6wATA1ujL7dmxFM2qS
Nb7fm47f3Vf78xYlQ8Ma+PlLqA6qjEg+ZjHWC5qkyiUUmBR/PrXNeuSWNkJdREji/cTI1TTiS6+i
TBtN4duvR6nCuf5n/L7S814mhNxIWCAGkGATm36Natp52oEku8TqxyNZ2FVSlZwjOeM25PkRH/NQ
6OO9KYTNMsmvWzfMinc/APvRjQA447EzS+DrMKc6XPXeSQcqFcibb0BnYKTaPt4mWWfoIuZhDgjM
fBVBcX0o48bMw82HOsCI4/fCKrq82J7dU9M5Xxmz+EPPDKFfo+D42MGxpfoJGpDkEkH9M8XuUyI/
b4AuYmgaaK7XLn2wnQlHkSWLEo+DpRW+2waVNZ44LD+/yAtgGFPoHFwBgoKNHqDqWFQT/OdHrpLE
lxGsQAL6scwjcrU6buJrmh7Qk3lj6q/fuyROGwXLVfDkawzuSMDQROXCYy2B/SS2QE3tbz0nS9B7
nepGL9wImf6ZBVyki/sQ2QmucRz5uuUJ6p+WAoc+ZAGctK9xk/Nt1dcxXEUewZQ30ZQibeGqY9kR
+tXAdaduWvLCTM9oB/9TZhsy73pEg0CFnR2n2Gw9KOkXNnCqkK5u22bh6P9XAuROc2LZgORkFN/5
ChOYhceG/avr8LCbC+BtM4HWENZlkR+x9v6DaKa3Ewxeyo9RSx5CunLNEHMyuWychj8n3RHTkAXj
48fzU57sKsYjRkO0pvNZHWJzClmpTBtT7hoKan2RCbMQKwGY6D2uIkLH/klokmpyM43PoTj/jeqJ
EI+L92nUkIlcUxnelvlVKQJDv/iE2hhinlZaBjEUy5yWDKnU5cCXgZrhU4II6F4CLYKqHd2mx48m
+6CF+o3Y2u6kj/sA14Y+mAo0+XqadtJ33lP/wF84ytNWnXpEzgch/3bBH3jEKpPlSpWakVtGBhJL
L4E6h7v6ofbfgSzrtSDPLlOkTL2rtw1RH3wjXj9oif3dKV1aqnQO5ng148U9yuGwxY84BRt/TTTG
7963nu7HSqECuTWRkeGctnelZURrYWXyWeY/xm3D/7U8GvNnVCZQUZ/vjoFAi/puA5d+FLwIWnl/
7Kpk/skx1X0TA6HXtmYRcmDkX0MmV/8uPl+xcAcEolHiLQZ6J5cC3JjMW1ztvX4Fz6KS1e2+9dlx
Vx8JGrNUjS7idNGsH12I+IxD8b/Gks3vMR61eQZ7l3pvcxeuS+BhzRZWqx6ek9r1bCYuDDSn2NL1
k37uHWZTPr65tsPovw9fKs+XMAb1vz0kD63ORZb3kfBY5w4N41bWuYAkWCxRW+N2rBcS8jbi48Mi
KHKulIvZT+0TdWt5ejeImfxvAr7e27HOqnGE1wW1LrCm5LjzSQFKQNAasVtNCgWt+L7V7eV5sUyp
LPYT2fMqvCYxA7GRv7Qf/W4N7nDkowfsy2CrtXCmOIhMpD18Oh2bgS6/Bi8QfMOuuCEKa6tqIR7g
S3og4A92lLQfntVtYhndVnT43g0G+88x98YjjgGSdl+p4SgjMQX96cX9y5W5ZE8tHmXZdVUfJBUw
2DDkPoPgZsfflmI71qF2XppxCIWH5IujiI7jB5A2FVVcTgEKut5bVLnLkANWthITBhiY/5IvHmXY
BfRlA6QxwaLQa/0TJHUTfxLXwS+5H9s0HumMQElFuvt2rlnwlbYgr88SLH1vT48fCaW71Bz+2c28
78a+yAzr8kIlRKURwWBRi9klCeIFqMq5fm8ACR5IBzUEkl87oEKZrphHjADlpoHUUDXDlQ7yYE0k
n+hZwMMSzzwVR2r8cWwViakb4QZ1GmoP281Ly6s1HttcgtVUnog5IAGbdbPtTPZm5k2WQ2ojean1
KXshmmaFzNF9ZOEahcOpB6E6xiJthIVMaJa284z9FL1fHCydkY7vHEbwb8p0NUlglieCHh0DkfVu
CQRSP/P3nERgOLb1WuXNhoQyZb/JX1Zt7VxiDzJLCF6OIbehdInZ/vvXypJsuYiz1zIW4rreAhbK
PTIxK9UDGIyI4ysrymrOxWTNs7YZYse10hrQYOm299i8xOdQYIWfARTIvDstWpSldqEa2emQJyFA
Wf4IKu8fHj/RBqPjwxKbcd/u/MgFy/MJ/l8v/wGQr/xY5MPmSa++HTiXDg4l/qgAy7N8E3TCRRav
ryf/rlVQhxRHV9p7RbASd1ObyrJRGIHYLGfzUXHm7S1zukwEsgYtuiKEAMl/yD2oLyFHbj3zODzC
7BVhiC8g2hBYEakH0EEmFwGlPUXtGnn5OZ9fmQiX4WbBhutPW9ubxQ1g2BEBBi8Bd14agQt6m0Cy
wfb51UzQv7Jrk0PloeNRZH/tpHxtMoPO3lvMkY09S9oPDXlp8n7QOO92tEjpKF0SeV3N4Mtot2PR
cTsCRLAUixo0uqX27iIiBcMuqhdaC3KJCgrRyxXtKU347xG9cT+/bXDOoaLQZcmpxVkAyRpEdMFm
bkk6Jm6PEx3akm891tetQJJoNpM8MdIFGg6MGuzN6U5HH6HfT+LJo2Sr2kcuO4Efm5MiHZGLZdUT
mMPlGeD8D9ZMKraEPZjr8X8hozNOmZvbNkPOFUBI8BqqR3Cs9gcVJ12OLqgz7JAZJekX4b4id8fD
sfrA+I4NoInSsM8Md6HuAzmD5fOERKZEzCSOMc+vraKXDNDI8US0wYrRs3nd+9YAoVNfzI0T/bbO
7Ev/k6giALZ1APDPw2kVWCw0kVmcaSw68/1+MU5x9qWX/W41xILXYCz5Fy36o0EHs7QlYAudz9Ox
vOgJ1ocb9UdBHh22VfGE9z7/VnBlgU96voJlZ7jyE0oy3q1mxaTJGbE+HeY9OHRpWazYZOPABjJ1
sesThaz15ig9tivMGMl+gyEyS/A1olMxNI9n5fyqL0WvQ4CJomuzeSBmvlOo3aL3jmrg68qyk0Ag
B+hj3dPi0646CCjMGKObQIrkhx9HX4QstEVtrb/dH4hg51FHpEBfICey+QU6TgZR3EYCFi7KZkBk
bxvD8612Cz+BVrg8VUiCFIgIp3D5IWWHOEGr4J76uVmdA/hH7aTG8VVRtgyo13gOH9qXBxOOfyX9
1HpVbDq4de3BOfHgn9xV8NKHmaNnupDqj6RWVi1oYw+cAr12BFULXcLM7CAuNCrq+sWsFKUPyVYG
Mp7o43FH4lSu9urD8jeQNpsobsDwgEJaBX4i+pxqDZ2QYjsglKBJTOECDcQys8Uyq2b9YIeYF85P
quS1fI994kJVnrZd2LEmEtnTv5slqPxBC2CpZXNgkaWFMHrwtjYeBBVhrSCR4+LYG1oPV8+LDRUm
EmrNQIQxPOOlOhhidqZUr1aRvhu32/btx+dEGXnEq4BYo/kfgQdYhySYjkrctL3F0kmwFPsjFjZv
z1WItNSi8XVACVsy5jQeqXLFE5NPFlfTuEPnZ186I1VmBBhyhqG4yAyeJBhnnueNbXCRQrEYwIWW
5SjUtDfaYAdVoNPLgtM8rbeN/KxEqzB0H7JE4uCieXfMWWK1B+5cPGvHnviWDFQEQI+WMzB/LSNJ
fsLMCvdZAfWpki3JmEtRijH/l6hIdqnNdJIHTsb54WUGllNtLsCjZPGgdFd4LdKRN3ehZjtFEUxO
7ckLl8fkRpe15GeFcGTRkWPENRVQyP7fhb4q8Q2gD44SGSk2RFdqTgosLzxmcieXC2Z8R95XVgiP
ypjEoM3yUQ0qV+U7TanztymQ4XhdIBEox2GU8jkjiYzaf5xTihxO5flFUzkcLohtv8TIxdSIyLgv
/7K7moSWgQUkHcImkwPDX5GyYk0U4aEj5tj4tavpNTfUDoorO7vpb/6svs/3Fb0ucrelmcGdtx7l
BJ/WUr6HPZv+U7ptFKaY4vepyG3ME/VY95ojxojS31ynPg7FnR2Y6FlFhQVKTppUst5C8UI/9+uC
8fZQW6iLsETUO6B9h+GUr7XAzFf7a1I1Bj37H8IqGYs/A/UpL3NUm/TxnaejgrkvF8FQoI7Krio3
Wt7ffZr/yhNIq3YP2553HGJMDNlsGJo3vOyeQxIhpiwMirXp3/ynIjl2o/tdVpEOlM41OtZBxNQ1
lqtRhrp9W9b6ThulMMpbAf8TzreBo7ZCBoBW15DjHhp0uYBsYpy1HvNz1mi3/rqMvZOVoepEhyoQ
7tjwdUjgNWXJCj80n+/xRB9KKGgBdoiQrT0fcpaJj8tgPItr7bECr6ZNHn7onbaRVUXtzgd2aIAg
mM/FM6wX2hK6dPq9bASTXdxMGdvkBu3d+WPjqxWTogHIDpR30notuwW5HrLDIDvmBfYWG0UcXOhg
7/0UlvI+25pfulqkWbzzDDOKsz/Wo2LVcDyr2w34aqGpV5VHoyw0ApTFMn0dznoxOt1GLRBH85EL
jjFSt+45Pu3rtX+boC5cBm+c9h79sJikXbnu5FSNscoHmKO5WYW4RmqFbBmH4KdCpSpoJQUI2PIK
9mMpyhi5OiDRsJWlK88RPoHuyidN7cc3k3pKAasZUlqpRZ6bFuUsRS8HGhcmOFPPLfu0EyV0Nouj
ML2BI1vVutDjZdXJ91rdcJkQa5iph96eyuYZJAppJ2LbCeZYSPEtVdTQSL3WW+xAMZSKYYeWlZRl
QV9awIR6SbN7mDRdG+nnhvPIOPKdaFfZ5XjXEFbsLS/23Ay2RAq9ieB+6D/oQijmD97g+Z+0R67Z
tuJX/b/2MkSxAxQHw8+1W6qzdPeIYQN5+wbudJHwe3zhReKQmJaJJUP3NTRZfA2WBpM+htBsoY/a
lFESk1Fxu0TYoveXIf3Eh4N3YoI3XfZAkyeZx5dDRcrl6NWR4OGtyWX0ZuqFPnPXYTitpni/SpFE
6HKXmlo32PQ2JrGcjcbz1aJMU/6Or+gyBV9vwjM/mznlnWdRoZX4SNAuhXn+wY2149+dF3KV/w7M
dhGQFraBALvEy5FEm52WENk1xKtxW2tGhTJiMMhlNqpVWkumi2TwV/zhfJqLLKhWl3Khe/WBwt2m
jqcI99cAjXPUfJVlNbeAmvJ0eYkl1m2v4EVKuuCzYirnNaywqporI875nAE5CaCsgD7I76PylL1e
ZQADBHlqcmNQIcUU8V6VMUev1y+4SsSaKG/s2nAOoNT4VujFHaKkOfv3jjW6qnY+4qrSKoGBFyE+
1HhFJJM44O/7pZJ4rDvDrkMhAD9wFuI3xiFM/DqXMTVF9EEwfn4hYOIpd3CR7O4/AqJ3h7KVkjKa
ulXMTCWKfeLSW1LWZ8U/fKe9YOxff+Wqmzj3V9H1E8Ipp1T+rKQktkQ8mDxbDRkc6ifPpNVB5UJr
QOuOjRIfsRcs3D2aUByOyAMBpQyQOPL7O/7VEytWAig5R4Xb84RDJPC+2LK6H/b/kHcYWfhe9pGP
hMZb5RDhU6qSEOV89aQ1Og4PQBnSeh+iZjye9JzcHbKtAY4fAikNdc/yc+UeHAP+0tM/1DbsafYg
5W2jiKQ4h3a6ROU6u07KnMbondTXNPlvxsYC8J9n9xJK4n1EZNPEmCh+c3/luMmy7kKzQ34Dc2O7
Fky977xrmsuz78gn1VngyYM1HLek5PG6SWcJ5SPhvFttU55b6kGZxtxWndD7kMjQuOV8MVhZybRI
H8UpNFCGjRAQ41qhLjE5Y6VjG8fnx830nEN4b+z33Rc1zJAgbNcta6svIca/DALuJa3Po4/iew1s
xehrixz0c8JAt9lXEL0M4+sbYJflT0q1gJ1hzyicOFHtdLDurVDg076RCYXkUrDv7QMpUHb7YjAT
uU9bCaGqi3UI9u0C9SJk+FJJIoQ0HvltIPc8oZ0lOAfuyki8NQmrlJpPr1U/7bBM9BEnRFxaB/bd
Ocw/ppYqyKZL6yn1MnLAlRHOI5EIud0XpG0q74nrYy/rWruQPNTjZ0K4rEQs36fgelxg0EcBnOjE
HLNQsxXKYbRQ5eIwT5I6vzRjgt6A35mn1q0Ll2swLR/8+sQamPlQdJt4acLwpib4gQc0kThzkDEI
j956PDPUOjtKR54QpeJZexS90sKC2uXa2uqzuIqTynjK3KVolsD3dnspMLfiI1FTZBg9sezlstW7
X1IafGMEzW6hOnxr7RJWSd4tsoWlXzHy/NX/RjrRsHUebhxGDJKwrmi/eEGv2r6g411G+zNIvaHH
qlVRqWcAiIcEWO8LpDil4MKCgjdFQDZ3+dLhaad08KsW4A0jD2U6cl9+8TlsdEhHjdsexRyfXXJe
bjIPpP8YCKn+n0DNAXwAedxdZye0OzVYrpFPIwINGVqiBcfSzGgQpWrZauGsyfNdr+5t11fgqDo0
yGAxEggsKTfyRoiBLohTylk8SE9WAJABMEhq1qhJZ6IrR/+CootDXzGoFhYPyo9dQAN0O0our9eY
qbIW5eAuv8fexBoNYHIT9nV//iQYTOeStLD9VK2V3ro101hGTGUAs3rT6knAZt6HXfY/lBNOayTn
ZIjSAWryxeCkis/KGsOKDBmB36+VBT1zIhn9lU/O79iIM7FMaMaGZFVio4nzBtB6x+BU9q9H72f5
5DjLLuTFyzbs2pOAIK+Fm5ztgUS9UI8aV/8kaUjz8YS1LpBOlI4NMhHOlKvK1xknKgwFWOj/NRJ8
vgBiBykPv+4aDEUZO7iu137dSjkmvVwHqnOMoXY43rUfAoavVLcRpSB0T5sQLxzqXKyCjAzK9Mm7
+AbDnBKV1PWF8kSjyTrnEw52sBZYP0EZ7a6mNTd5UkWjiltL1owjTQaxNQVyroEN54yDzK5gtkhJ
MdVMvrQKN6DOe5Gb9ghGlckXfl/kIdubt5NS+vVnwk/FebSYvXTh0trv3cWQLVsjmKr+mvnKcEOc
01JeSMuAJgQoC6Z8GIH8YyFwlU/PzHefj0CRS2v0iJHAVIY50UswLD2IhO6u2MeCqxZqVxbQcOsx
GwUPsS3xj7VmSqBEd6So0Cd49cX5I5tryBFAQ40LTs2HZ147EGXOeiOelCiaWe9IxpEW+MXw07if
fKKD8wbNCeCpgN8OYZEynfZlO54wAZerBHU9wfsUyRHpkIVT38o51MrNweN4fPHK/mUL/xiHwHTf
WsvRMeeZJDKqOldUWbv5wswpP0uBVHe22J7womkzNDZdWQtiYhqSSZJxrM8s1+QM/x2+czP+2ANu
IIEgvqSVZEjaIro2NCpt+NuH9XPwXGhmRyO0DJuKJXrYiinUkd/QpOK5Qb9lkfccWLhlkHwwGm2L
4knx6uM7E8xmzc2w70/pAYQlZRMvgANHK0EjGmCJVbcy2A6/rYS2J/J81Dg9L2r96+mtXk/9tiKX
tyGgUNOzA5ecuVERHAT8nAi48g9rvveQkeL0Pg1ACEWRripXMQaFFJ/rBAqTGGgXAbMynxs/eH1L
ugigsOxDQnFQjz4y4tdjHoNBjY+x+huU4EDr0mmy6ZpeBTd54YSoJXSa/3E7JfcJFqHDySZq/1vT
NXiNDKau82JKrbu76ckkrR2PkptclXJai4xap4b34tKHeAx5V2bWBcaxe5xIQe3VVdE7HBTCYKmE
nHzdNXMK9kBb+nRdZZq7nU2IHqZrgi791gIIfEuWHTIv0AzlBD00DAin51Cr86uYkMC2RgrYdjPA
bj/6RUty20KiW1Y/LYwW0W6wIO4ObkmISk9fHjn906+x0BYyr+rvPys61RUzHjesFFurspkJmFJJ
dfJZbKdhbriJcby/5hxYweQIkKq/ZVQDTQKmjnSgW802Rd/Lfxx+qcAkV54hw5+g0aECSxW0DDYM
DU/n1oqjj/M70qUSmIwYB5EdTRcnRFmVbVJQB8MVpZWJh4iGGkoFwkOLZZp+vG2dNSVwjd6iZN9P
i/0YmiQG/PgPOXLto3yUtUNd0BSsgHccw3o3CpQNOLmE5ZERTR/cw70SQPHFbX8FGhANiI5QzZlW
3wq978LURWleYik6sIb2NR7AChjF76K9xk2u8EpUutDO4u68OuZTe4jdLmPNLG6120S7xAvyJmiU
rhD8q1JSnYwyGxt7R0GKDur95tzwt0Pez/lRh7x7NpyFxxJKCT+gxJT+ehSo3UTO940Wk3M5DAH7
jcUx9YSo/5SLr//6eYAf8timt1rTbtKvIhp3pkC99LGoxEguILiiK75Q/89aiJOxNfzW7HOpeaHT
GOWcXAY4V2N8CC4ULFIq4nQsEbOr1+Ww0C7PGyluXgPAKsvPlRwcGecSp2tSSXscs5zOudl4J15K
aAcy/5kj8CgdxfKav6H9OC64xyIfuLkOd3kk08Fwnd/vfq0sgFV3QX+NKCZcSzuo4gNhRIAUv6hO
wcfT4PUK0wxTg93UZiDHamzC7goiQgmqcVBcYh5y3tlukihEZzuNgrVaumsiSg83zT2PYZvaEIvI
ZlqfR1OfpMJjcTVNgxUrtkkXFzvj/HeaPVtVzJr81yFArB8EQpBTo9HzBCxbbCcoWqz1UjByGsAP
eGYIsmcy9HZxbi77MAg4d5HwlLB/JTz0rkI6awOvFbr7+0XRRhc2Ad+xP1e7hpfec6FdpdGRhFVj
Os8jDxG9UPCv0LgCmSdGuNlw6lPalfTOOQdog4JE4x5DKoiVMpLNKMNNRM0FBX5KgahQGnsDnFHX
NsKzlmZuPxkJC/pi1n9kyRJdsROwIFS4e1mYUBIuOLuxbso1BYrsPwlzVL4i8dH7kQ/nbpNj2Bx+
JTEcGMMW0t8HvVw5Afm+NRyr/fa3c0aeHxL4IF+WZerQxoeCfQ+XrHvb7L2Ko6xoaDLtPviRlTtC
RvNyXRmv9tP4x68+q9pHiquyFc96k2WcegT0n+HHLmDkXNISByus0QgDcOBKrHbnsdqsJ2YYd6mb
wqPKgYdKk1u3zfFC3HQOQBiLUZwvSeHuh9C9sF6sFYaSOTuFgZJ6gH/WoFZUIQsqingp0ch2W2ng
ZdUHNp/ibAwGxtFXl7KlYARSC4Y7jf0v5F7kw02vTiPthNKD1DFo4I18bxVcMfdv9q7VXTHkIrdD
iJ7bhgwh0EtyItfzzPdqAl1bm2b7g3kFDXadLscZDx68sli1b84oLq+Tikvm0R6w0QcQoGw2O+df
Byjl2/40/Yb7QE2c7r5/s+YzNG+6OwmNnYzje/mnwZN2rKef3Bcx1nsWeFmAQsvJsl1REuC6OOfk
FMPNVX7/lLByGIA3eW2jpf9pab6ft64QXlw4wPCXr0OyZrMCLq6hmYVRRYV+rlSjyliccacR7CHT
2CTDzOvlxxjhWaU7+PXbVvEHF6gFn3ImoB+Tb90LYMm6uNGa69inepWT2BG8l+z+fwSIS2UHDKQt
BrAkOzGD95ecscIzYn2WcEdSN0TLtOC7tlG2oE37QXJCz17Bwe9TgZfs+6RmhlGTEOu7o1D2S7Z+
8gIwxBEImnS4ghvLOACZvsD/ky/OofkXqZ0PNFIvj4Xiu5SEFugeYhp0iTD6dRbDCgJ01Jya1PX6
q/2RCrcgvjWUNFTkDYW8eVt5JpyL++RbydW11zgma1qAvlkqiw1Ivc+GvyldC1oXzIPz9BuBS+Yx
LiGx0SD6hrcONPsqMM3N1JpG2PdcLTStYHVYwJ5csx505g1EtcCyMPznp5rValgN6cUPqUSMz3m3
mC4g3i+FUOEkJ8j6w5saJF9Bhx2Jx2FrpZqX1u66ZtPuRe0huY3JOmxToC8MQMzeKFHIjVkVKLI/
N0SLHK20N9k+Bej6Vvau++ZzXU7hMPMERT7xqJ1xPGVdHRP+cQcbuxSftvFHR8XY4h+sHT/XRH8i
yExWqo4QyHVCEBZYzwVHtrRp9La5Kptt4VS+fpYrba9iQpfyLH3y+VY5qmRBOLpRDkEieR7DI4uM
6vzbehWABIhjWbiK89ftD2/VUMQWejBB37Y2eO5YEW9UH+0OUwL5Y6GnMSuwVC3ZuZ2p184H00dt
kogKi56Y3Bc92y10zXfbTJiyVgSe1GjQMz9rk7ndsgCoXHZDeB7TsWVjwV9O2yqao6MW9hHJ5+qs
KG3bARvATb8qMcjMLpL0vqjAjX7uE6YPrkHohpDoYqwLM8kJBydzTX/0E+8WVi29GuGgv4WI2zeC
MBaKCGLdV8l2LQ0dGv+G3zfDfPlkYqKkIq1bxoUe7iYcTTEi8KGCWHY2qI+F4wTGAyfPfIdML864
QDvDpSM9gHX63toIk7uIk9L4ErEoMj6Pd4BJK41Hrs5j+gl/TAqLOiL3e+dYom6xhAkt3wngdnzF
+4Oneke/vryWKpfaYxpd0Klmjj6lY5d15jPCxc3lV7KY5/aXtkGaakW1XKBqA3MKY+rnxEka7OW0
esIk7UuDRs6hz5EX0qiuy27t65ndb128aDhh/61Jh+krn9u0y0qIn0MYqO39xt6ZAtR3mZMPwBwe
9EjspC8DsN6ZDKMTQFngCb450CUkXVK2MhHKftSuWnkz583+Nj30MVllETP16s1hNbJC+B3wVtcV
dDtDwWF0e4PhTX9OhBI5868OjwUrnnR6KBNz4uKpdDRKciT25Z4VGiM3XXuxqTsMFNAR1bjqPQL5
zTEGFAKHY5ZK7JCzFgv3/FKGqIXQr22UxE14wvkxIUEUiLun1EfLIEv1oWi/ovK07EIrZm+eT7sZ
ceCdDGGxLXnImcJb/rBmMe4x9s1oOU4zwRCSTqtncHQBA7oAIPp636SNe0MGRB4OEa1MzZMVvItu
y4FLkJJkfWPvizRGjApEUOUQmX2VnUVcS7A7badRwz3Fu/sPMd7a9yj7J0pycbkP+BNigB0hYmfk
fwQK1nWBWvfrW10+AAu0+WE13rm0VTubuuYoGBEeH5oBYzhiMRnBU53ypqRWEtTBY8u3SefjNraA
Cw4SzCCm0KWtGvOAVhbIw4rzgV7m7iefhSnZZyjE/ICXyODbVzS8wC8u49GYCyw33vjyUUESfhxt
TJnPEr0lSyveRJibf/ohCHZyMLTA5kPyeRpaNvcqZMSy3yJU3/kKLMcb5M4ikueQx4IXlQVDHt+W
GjaRczVIbNkY8XY/C9DEoxoi6Nx07QcZDpXP1pcVqBJjcW8NZN3UJLtKPB/7hRjA16kppbApVgsj
q+2DMRK87wkBL0lJHG0jLww+VN9wfAZd1qH9LxwbL9l11ZLNlYCxbbhXG+7ImQ5Rk/9WiaHrwZif
eZgENgeUZ570Xvz6hcvNpWSuDOYSQ9lnPgI4MPyBQfoMZnk+3ya8Sabju0zFM0xKMCEZvLAtMrry
EmYVMvCWNZZL4p5b7IPdnmaD12HOdxnYKJnG+14G75VaV5JtvjHYmfFCQ3J09bC3GvjqoDBNZT6f
J9XnxqYeZywa1pYr06Up7tlxVyTtbixpHgSpwvaSl/RhVq+EG8JqMyl4AP/QY5zl7BRAXMEqtIxQ
dzTjGdGdbsoeFURMKWRbySvIhFH5f2R8gPKSr10J+THXje+7pyQbG1x123uNVpntcSG259aFW8Xh
Je8BQOrS20zjlYviyuvvOoMJq+7smDc+PLvH2Rts7iJt3RRGyqm7MnA+nqh8DDdULwyp8D519azv
/fWE+LQlmojdc3PNa7i371q22BIvDLajTeJ0epgC0t1R+iQKwyGucouei7OEU/oDK+idQ/xxuDmA
/LBZT8yxoltAAtkzVsceU7qOwXWe7ABWAWCL5NzX30K+TaLJ9wzPaaxwPAQzXa1s5F4ZP8d5fq4c
Ou1yqEloQdKF1d62mQ7AH065UzbSqPM1Ss0JBIgCe3NqQf3JsbDYO/oZ7TOKdklidm9fTjJXNZzR
VBl+vjmFNjVboBYaOsw3wqm0rY0jkDh9MBv04dnidfGHoOhGYvVaQShJI8guDNYo5ENYOrAj83SO
V4ZVruBa/gT3wX+/OjuETq9t2sXtSlb/prUddFur3oyJsfb6jHDARHmc1quPLDGig1KXUqXypnEZ
TC+0TYOnjfOozbCtI4ms5sQ/xAFZPw5A19b/05gQgVKYmID/jmjwiEA/vJZDLSBsw+qc43k788xM
XiEv+86SLeW9I8uVMuoyZDvWeV8PpGrGNShA+1OLze4LfVg2BWrIuw8X318xBCQDFtksCFkRhTPR
m8LMn72KGKLmh5EyIwGmEx7Tw0Ry/nhY2mzy8WBk//IJ8ugh6C2t3NRxhecLxqtUQaDoPOLljofV
uSNjYQjYlTkoRTJIF3M/A3Gl4ANptpiSq6X3U2JBdjjslYLrUhliBXHQAjDQoqx4cz7boV2u70ty
SOH9E0Egl8QujiSMPdSFBtwtjtTOxRO2uyNg7ztlsIPoiJ3s5PDz13HNG5EIwAlRcL1zp5A8V0r5
EP/522lW3RG/IOlwvTcbfQAQU38YY7d2UixpMqIedwK3W0wuFMjmj6UtuzLsABMeIqBODCEdgKwf
94ht2svmuxmx4ugXiwgwy1u4/YhMdkcqRQ6nyMjKkOJC6qqAERZSmJ608p95PpQmbgv5dYia9bB0
8lJxBmtV8boRNAoEve4p1Up5/7rjRY0FIzTllkT4t37/GUPY/VTnPST3P+TNByC0Mwnunue5htiL
8efg8jLBnD5SyYENzVqNESENzAjKNyZ37c3riSCxNzgGBW5pwxuGhceVkqSsKCNl5F3OzjKTWTkP
53KHY8MwLaP4viJ61ErdVhqu7Q7fGoRs1IJ0Y9oSVpTqelk5dOso3LScsU9VY2yyraSGSJXaVqkB
9o0Yk0Vulw7ky8GTXkzh95UZ9SOeXBSBLSg9gF8hJBksR8UyAjQ/IKG2YoPj1jl7P+yORAQlGZWR
L9LX7TDN0I0atLfaaGf/NkiCicolP5CNS39tonxuDEgvYkKh6/2eGHPOczUVFZp2MWlQnNYbDU3/
uxqRRRSbZz014MgljXrTKmGN3WW+bfP0SxgQDW/C8PWz2Fjsy07OV6uQ5ko9tNDRYwEv+PgtnY9R
Ar2Ue5T9mjXkIzi9PKi5eIi5uoQloDu0uFOcRJBbOtNCG8pIz0aToQ9d328OTDk25UlP6JwwDrh5
P3xRajMOoRJQUGDahBZdP5s0U/GfREWzYj0FnVemZqj+ZCZogUKCvVpHigzpfZyIK/KugGbFhwJc
GURNiQaIc15wZLj6/VKaijdpx/Ca9EpQJqwVlbhwqSjvaX0P87pO59M5ypLv69nmOtDDojeKlbt2
A6YyJifff80IvFLUiSOpS7Mx67NfptCtfdJ36wvIa0rueJU5i2O8R20+zr9ZjQuvv8dhcD0jBYRT
LLAOmeJQJlvvWrJF3RH9rSjmENd4KSvsKJ08+yxiF6fgTg5TJI6bQMCz1ITzawGTdsZ1yqQQ+2cP
FbmDkxUksxnd1Zf+UcakaJFXDT7i2KLJqViw6MycSr8Y2PD4rdX5xZC5fX2e0lsTvcuyCTWUSsQ1
DoKb9H24FNG4dEXFx1pQNws1JKAMz9N5reFgKytm5hVF4pdm8T9OKDQtF5wFlAXjFSP1Onu8XHG4
IspNCmarL5BtpncYXGegKhUdKS/U8mPt+Xz82jiT6h2WUyW3OdjyXcdzzm/X/jCfFLkOdrodmEty
+U8q90HsiKlQUp7pq1c/kMmHSfkq1/CQRpHqfV1R5HTRjRllNlRKGhlMmtr5SvP6r6D9sMXdwYcp
kDxyxCdvLerhVrLwmGMrAhKtJOjD3vDbMR0qHNkH4jCBcCkwvTjdXxug0YAT9joSUiFvLc7gQa4u
roSSXh3N5IC88Rl1GHB0YxbTWmZH+xjqqs+e2AXAtyqQNjpq4d/Ngy3cx74Me/rUivyOahTcTp7h
HgPkD60zm2ZnIxMcYR22ZS6Fmi3I1hLzpE9IoT/Q6GRLpYz6oSkDviv4h2oJNVQazQLMLlFBh5ZE
CeNO0nIyTWkxuYgb+DTJW6iwhZmrbUuWDahSBH399FnlYW+S7b/5LRiMqEw//+yvFW7pX3Up8bB+
RNdqERjbCaDDzzM8q55AeNyw5wI66BVmbodkVWWOftbtvVLujQoEg0IE3OokBpTFvpoQp4gV7Jz9
O6AGpDlDf9qFMjQfzfqMjghxgdINHKIsHYP/VzXswQJIIAuCSFZEXcjcW+0sCZaoJ124GLbEU+Ma
EGRvFzUy28Uff03CgMD9RsLXgZfJ/SyuwU99PEtZKTElaTopMBDSLYEomf9r+V1U64LlUrMqKdxs
lKpM0ToexTcU0AwU3Jtis96QN4JTrlK+lXCUkHoS+2XeFM1xkpmG9wopPj7g7jU+ROTnsihVVIgs
nZbHn3V2R4XL646HwjEHx2xNE7fwXW0nXiIYkGNrixIe1wo6bJ0ZieHDGSGStdi8nuAVOAzQtFgo
lxzRDqPlrYX7m21R+7rwn/PoMC0lCBcrhKb4FIboNboahZlS5TukIGWIJqol9pHwQH4A3Ti9xKHN
WGYO42oPtENPseVXyXtsuFXXkvZ4qGz76CZJaaGejpTWsZMskCNvL68gs3Bc/UsstO41FdRC41FW
B+0dUg9qbUnlppCetSqRZnhpGakc/NUcz8b63cvTBxpUz5zQbBgFoDrdspvi0cVuH37crEbSsGia
CR0Era1qh2GEqL3FTCnsJw1jeCri1dTUhhOkCABsE9u63muOAsqCbNyLebe+5yedFLXWA+RztxiI
3/dcrtCj1fCoKFToU6APuCh+nXhBwb44I0jIJeoXQG5+RyfcaMxlzC0jJevPg6XOnREeel7IarjO
sPIQUTKZDaVjUZLiI73nFvq7CYFLHAZhqV8Jf8NcoiFHCsABIeAd36JlWbOxNX5It/mw64rVtKAh
kH4jfQ4Fszy5MvcTxIJFjQ7oN4Dw+aa1REKPNpayXRQo5dLSIBXwWRqxMdlzwj9E2bVa2wug144h
C6KDyZNnQq2cOjxH3FfQF3W+cUXCODVmhgr0P4kQk9ZTy6/bRHUZFh9joqwyk3L4ySeAiXh4gp6Z
pUfxT7u5DyxsFg+LrC9anmFz9d6wOXNJfdHeC4QKel0Bvf1KC6OWA3I3alUGR+CTvVPPOhLG1Hsw
6qdieNXmjkEX+pJ4B4M2oX2IUi8S0jEmw+gp25QapJnMg71kv9JYgS9V+nKWasK3seTKDt/Rl6NQ
QHPjXD2FJaZvlV2MNPplJBnO8N8J5m+UGZ0a4esExBYZB1jxdwNmu9Zgp7lfFhVzShhagyQnCROa
Wt3wsOmA8wZqvANdhbAy1GNQpi+SqoXbVjCX33BZ7DzAGPT5egokNc/uBSTKCrMll9Ft1Km/0IKZ
Dqn1MD5Z5h9yfE2V6aRgyiQqQbGVvk5QF0jqL+VXsrNhHPF3Xl3G0t2G5pz2hyqZUCWt2MMdSymW
VNEDrGNan9HvoeMBOpkCyFp/MWvEdgDJWnSjcxxLa1p3Rue/SOtAiGzeZnCV/Y3liiahZElzDCsO
wxAo21ZkhTKTlpAnELQZfRECdE5vDQfes85kJziSjpJ6y/CyZeiC5wV3aCNWRrkgT3W+wegopAkW
OEAO3VhhFwp/zzxsePUtqE/Fq+0Ooce8X0ezr3kVLL+Tia33h12EG4l2jXpbvI39R4mBExld/IVI
0UkeupUUto2C7epcVi+FJHq77iIdcG7Ofexi/TChsNrpc4csGNCs8MesDYru6FU8Ty6pKjItI6WI
aNmCiypl65KvwViZjzCcKgwPaDFeYnWEQ2A6Lr+jfjhVPpmHD2QXMJqbHeDqKcf0u0T9aKFWKA6z
bEDh0QAYmaFDyCXl+5iyh3llib5YiMEi+ulq+qAoE67L6fo+1f/0Lmq+4IjVLz3u1crIhId7xzJC
+r2PR6NG47bqUJDFhZnKhrWTKWXjAKlz4ueufhI9CL0MRugvEBYBRKkef7fCFDHl8CCjEr5cNK1h
9zBpNzconCn5vEfR/c1C+NZTxJHooc6qGCwzOLx4Y3eZJSJ5tyfyS9mCfnIRvYeDckEvldilOOcv
tzjgicJ/R6TlWpj01lWPzbgW4dwf/lBg1FxaILxLFFIl+2/4Z9GmQNV/kSK4Im6qgHVtV4FvBQhm
BJsetXcKfatK7popg4Vg8JBItlV9kXmscFvQsO6/Ok6Vun253AGdpqCFBj3cMPVYdSwLliVAdlEo
22TfcfvUEk+B2TmEigdundT67tWIH5IZzpdLNeINoCS7rOA9M97ehItbUluwjyLzfzXNXNJFAmNF
gVTNbAwE7hqdHwPb+q4M3uX+tHwXM6Gv0PYiSP4eS8raHCRp3r0GiqY3gAmynXPCezXQFRcGNac2
LXytf324v1RlBuByBvjfJdJ4m0Q086+UL3nXcVApinwTifQEk+uLZmOdZDzapA+9F2Am+cWJTD0C
NMSkWZpSo6z0S0l3AvoI8YqQQ+ymrATwdVlGlmgSw4GrPkKEU0dG9bX5HzEjn+3970M0jrYcqfyW
dTDxTHFgyeEpfdOBNOdHso1pm31WmL0PvnBqUBB3f0pUp0TxKnsrxfFMNg6jhuJwFfUz24hiiG5w
NwoEjW+/wdv9tp71WSyIOG2TWuzGgAHPNctGg4mwR+YfTbt1Ja9xBlsAhz3XlD3zEd6diBICxXjH
78vsAmbOzMpD1VaeRnpn3SHKdD3COhvN2kX3dsBLnFTZhrdeIRo5rlLS+e8Yy/kmZGvTzHyqUjCD
qlYKNSxt1GwvREXd4rCbc52G+T+VS6fVERoROPyzIndhStmW5N2la5Ejsrb5kPzShOHK4WVAsD7w
73biTrRf8X7IFowHUIc+1otN4h2Um6pl7rE4m0P8o3FK2EX490zoQSlJ2grLFJB0y+rkeS2uwE4G
Hwe56g0TLC0wi6Cze7TJqsampRNHsG7rDVbUSwgkEQ3zFneCfeZaWDSHWBotzjL9+eUtVR8MSc28
3lPhJfq2jYetKq6NrRc2nHuKPjd+m5seKGq5n2N9RNoFWparJ0KwguPotFhEzoZQbt3DVwat7Vxv
3AmMjhHziGvGsTFQ8aGqLvUaWeJyhJac+fbgYiPMUUJLDbsJHBQp3e8OXOll1lFewwLf5YKpo+Xw
Yy7/9UME0WYex1ZSWtAae75aF8foZ1omBYg4oiQFA8/+5on2r1Rp9T9OLjo5S0rBwacSYQL7999w
ZGx3mDyJTEAfFAKUtBRZktxGfpLuHPsnD0mOMAL6OnQOFf8a7kfBVqA04cscsnCLd89BzgEq55qN
WSTng9NLEgoxZlTqR7fQH8WZQUfjgF4r3MxHJtxutMknjoyJFRZ4FU3Q16sLhsXmf5CeF10wQ1Lt
qvhODgvzhCsWSX8oBlgNT+9MdAIBhE4HNflsuHHVju8+Vj6Hf4bqoH37O9rOALpkCpAxX8O9Q043
Rand2B38z+9aXu28LfyY2myxvrFpgymg1muF6GcrtDu66jpS+zOgDr6Dcw4PD5jxttBEFiDOreH9
h9NbzXDDthEo0CH+1xwbJ8FtVolVBRQU2sJ7UPl3QsC9qgMiE+3do3gyiBRS/0JFX0TpKDXJwjHs
L/Wrhofia5m7tX+RAYOEU5uqEt4IWgiuegk0Al0gePO1EVij2i5yQ5hh6ZaemAV1fVVJnAYYqOhW
mQhtd7MV6UYGinUpm1rYWPWmRjJFGlHw90AF1C5wVDsltdM8qKA90OU+KOnTgCVM3XEQoKQVuJfi
c9BY0zvW1/9E/tvhaW10HKEcvibnnx+D9HgcqJHRpDM0F/28LjNuZojeB+zAoMJ5zJrvTe0hoYuj
fYiUe9YkEedHQ/JRJ5val0hJbukqb/plLGM/UYW9J7nkoXwALlEgD32ia/ALsmthWV3OKCC0mhhH
2eDbp8XL3ojnel5S6se3fFHAhWIG5QY6ll12T+xeZFlFebG1MKxP9utbxwLRF+U/tLkKeucZEVbC
7pDDf0rfVytQqPLV5DLL1TIZR04IQJjr5j8rhqkLhp3PZtYrgcpqUiDVS9xwJy+IXmqxWXaREZto
OoKbI+LMQL8ebaW+PHZIZTGs8xR6YOryrmPXoFjDNzKaU1wk19d5MK8lNt5fo2X1fDrzYCWIrM12
+Bg+mdtzR7gGZVj2FExuaYHyEW3ULTOIorT4Yrpb9xyeRBV0826tel1uOFhZWBLVUYALbwhLS2l4
iQ8A5xeTcSie89kRkbnHHnutwjx8eOoHKH4x7f6HdiPW29mCgbpejSVodQZXZilizWB7y5dzxUft
Ee96/7HwsZuqjaNgN5v2WKFgHlEVKJkQrUASzKWM0PBmxEKlaI2k18rZVJvS9hV3DUqcK7CA7gUe
uy7Y7S289dwRAbOWGy2q+gPv71Vcdx4tL6GvF0kuqH+T9HsdYe7JivymDS4HQhrnDIhnlwGH7C58
+WjA+a/BIrqFojlB7CujdRHKyJ2KVWj4phtrRlZZWbt23ElCrQcYX8GqPVyx+VhMuJKzv/wqKLax
jAX26pvkbRlaij2CwCDYt/HtuYoMdMzdqOrR5y9nkx1jbiT2E5P3d0z++avo723JAT1wKIzb/rFH
homEOdLo7dH5aHkkymPX+McXJOi3ytkMq20XCeQyTjupcd7HldutNtZgPRjohERRU21ZJNlCBFcU
IlovhQxSnvzkwuGDgqXOncJ8fCqrKDbhNG5b+f/li7gPICxotLSkhJJNgwi4jyjlB1sTKJOivMco
N88+qESX1m2lEIEYc9TNm0tqo90kvyFEBehTl1viR0qeAUzuTTI5MTovqP0GRiCoYQh8IuTD4m1r
jDoYzxivECHWgDRELhZID5qeo2wMI8lxEDNGemop0QdhZSR6YgZ492x9J6qUcAF3eANXeQ0JSM7A
WQRIGOaKbjwAzJOjObj/R+F/mq+Qg9uaDSsHgoh+pE/c35CnZIBDb6HsycOA99kQOsDzqui8tyuA
G5/uz9uFuEFYSMpYcbVX3T/pSQOUGPpsOcrg4399XBL321eWbOqAm1UXgEfVEnzSaC9uhb/WBs8L
IhulYUMSDqI5wltS3x32lDQY1TbS+6iyINDzyUOs0qGTjZKrWfrrbHXWUCn30jLTud06LOWkaAJE
oJPznIchEKObJCbWJMnoHk/2HC1Drl+gnIWXBkYtnndi993tt1Aki+iGW0PmYOjGXYxvqcrWyxYD
IBV8eaIY2sRV1Noyo1FJPv5heGsfy2kHyxdAmL5Mx3rgeQG2XJYRjvx1/1UCl+QfZm91nMKTlBAe
Lnq90x5uFGwXOtVK0eLqrjpENVrxE4Ds56ODtPbbE+mDjWQ1zRU/iuEloQEAHqDFLY3ZP+HjOhYv
TapXQpX5MFga9GtlgarkFjVT/cgdlm/EnVR/YTVmfzq6AwWJopLE4FTgWpwNQBR46XocGcGuHzrp
XWgL8/oOjX9wbu6BFu84GYKOc4glYQeUN0aplVi0sYSufXNhXjrBZ6HHcrtrWKLxs2YgLeynma//
5H90bqkRLJj67ZWbhxd4Qz18N6VxTWq0eUIsf6JhoFNU6bdDDBUpuMscG+oTdtADAIQ3G6FbHLv3
Vrzb2dpAg532GonRXChQ7nHJDhS1QzyfiF7GTEktg6xPiOotYbfXF3E/MWLD+7JB4edpTphe7YBY
mx91jAHJFIj0vg/UCj6YwgkhRlnyw5BIHGtE05E+E4jnh32vw5899N3J2ILH7y9uShOkfURBSwkc
Q74PW5Lepx7K3OBP0h/eohZlV3o6EC4i7r7il0LWSmeWP3seFbZIxBZtLIBbhEgKMuiThMZsEgXq
4xFFAgG8hUFdF6YdMGm7qk3a0UcbiSGQqre6AiXlVlzNThO8Cpn0XptpQcRy4mAoxHQjLQebTUtl
FUfhHTqsxnj2zGC4s1xHvNlTycYhLMsglbTExCOMFMho1Xah4E4eBV9IkfVKz/g6+KxqA+yssfhu
KRlcjJt7aFG1qVDj6prFUriXeSb2n+nBOpFDHD66Iu2lb05jNxl9oP7XNagkK0nlrOfHW3fuT3qW
7ApE6V4wgaTqvXi3HQ5c4CNhVx0kBPyoXw5zU2xtUnWZYR6kEHcgEa8AlHffZHMefHkZRb8J3Gkb
PqrXMM1TzJPAliKe82xzXK1nnWouEhVetIhQJRWOLd8oqfvaY28C0C1738/A+kTUHT6vqNI0Thcu
sbcH6VmTUHSBmqBCCuojG79vuPSBpcrMj7BvT5VeGfD3uu0o3I9Ay3uWWjnknT0cvPiyfxZ180Q4
5dB9ZMGacN9lKsumFKczKytLn/HCOrpPztGOFSQxxpbbgX+TYlFfG5AC/IEi7s6mgxkW6FWZfMJ4
qBS3Eh7zxMOxmFNTQ1n1NxDNqX6LPzj8gao/9CKCECPSbnE2xqz5c73a8kHpJ8RYwexG6G5/ScBV
umZWBYsKSc1JeiMXHKEBi6118BoBnBnM4W4KiHMkxKanu2clph9WaIssZmBms1v7qjWAsx9c9E7Q
UbSEJ6WbQrhm+NrMR/A0gd+sTvj5FXfM+1+8Gn79uX/PdBBn8nfiKABZLuVRH1T/pfXMbacQpx8k
peuR5n8CQ/uEhbfKwrzFrFJgxHk+IH7X9D8eX/LaicC6D6E/JIc6TDHLBfyy6jMmNUIN6D7smLkQ
ZG9ZJ5Lc6nB8RA+VMhflqoLsxhqf+22aq4gxNAm/BuVDIZQJeMdhwoWZCF+QC9yc6MZiiNojPQYC
RNPhJgDW24wr6KRUa12pbFIsEoNRfrOC0sEcse/FPZQxOqw48glmLSELGXXQjpPFYCw3H9qfy1Wv
/iR36eKjiQz/Ad7zN3Ds6A3oMIkW69lVKdpZ1E1EZ0JKEcpv5ZnhXiKUY7LB/YXgmpOdfjzQReaM
rGAhS82uLc2JeLtkSL30OnHmx/SEmcti/FsuUU7+50i/9B5gvmSlBMb6VRKlnxVrOhbXE2fFZOtj
kl0aNiuUVBCei40yT2ntuZ74kjbFIl/vvL5cfLNJZlYpqWAmrl/dyA+9zebwDs0M7cXA2ndVYFOR
bEDAeX4QzYHEceGTmk5mRI8prf7Amwkm2/O5kCbI44sK9fAfVWYbOaMSZ29KgoO3COCXmL88nRm5
2TZjuYHi/sgvX6cbyk34Buj1IAvKJ+r7lEss5gafZyNxTicOiHqv9Cm6JeouUG2XFISLrxJ/w7qY
K7YBcuDQldKNql6lCFwaOEn60ntVXh2tDDHEAdVw7Sl7un3p+yBLoMytzUY+Lb+alu9upbPW7bBH
xp2RflZin3QOBifj4CaWjoCn63pgsyyFVl+7Oz3iR+KzAsMmH70z2NOP1NOqM9ce/V8Br/JgOoAp
mVG3mtMGozKI1oMEdOAHnEoZZCXbBVKlSzusvIJdMPEU+sXLMGp9Ada9x2yRzR5NO6kltLciFiVH
z7B/XPWBLyVW6S1SONJ1KBp0vQdohFBGbbHxiz4hqyIk2KMxOU8thjAYhfliTSwErgDuh1BFsOZG
UAo58bekBoz380OgPWlgLpSOO7O4BVTx0aQkL9B+hBGjvM5NWkYMafwqIlby74s9x9D4gXsg3+7Z
dojef7CGkNK0RU1IlLK+lRBvKhL7YQbDLCVD28wn3Cqnqa9dt5M726G2Xi2DWnY6C7GG4D8EYrVe
SPTMajBCdUmQGu8rd8MFJaW7yPPO16fuEeKS9PSd3YC4Pko2uBaNuq4DuPD4dhKMZCnd9VYkH4zA
Q87R7gcSL0QiksnhftWCw0jDYNhW7E+I3WQ++96Lb2tYMs6lP0dbo68tWoR0rkKZpIaiQg4q2Wl7
c1JcVu1UCjyUxMOnGfxn3b8tW0rkB46WPVjKzbuBYRVypkqPm0I4WbFCdTn9IbXjEphBpLolxGXI
Ce75YxlKEvXDh/JR04iwMtS1x7fCe8Dd4TXlEr4ObMsKHDetVunMO9afLGVLfuak1fXn1EAZngdJ
e6dWy90kbpIKa4peoxDUf/lw177okW+ItOl7C1dRgFpf8bi8hGAod7i/4G+MsdvqWv52eFuG1fG3
xyOsF0suvZ6KMkN0LBEnj1oNMWXYXmrUMB2Ypy+pDfgt6DCxnayUVbvdAGfX6NgDIIBb0PxXx32g
OebYO2+IwgzRd5s0p7mS6XRzKgvO1gGbLtB0ua6/+0dTYFdWHDHoiHdVdUcNblsJn8x9eLqCXO3p
vOFFtecsElzh7URZF4AHbemjaeIU9cUmTlF1wP+egf4CVRlHHuV5Y5FeZJfucFCyneHhHAbO4Pr5
iGbE7Sd1mrwp+mfyMvYouLAXt8E2TrUjlGuRTp59tYAG+469+NVXP8VQJxIDg3YR/Vzlorl0piGF
pURh1Kpfk0oMvoAVdo/TmbQDHbuA74hghOQKwUhMOPO/wg9bE6oWRTLYWtuHH9ihmh8GLhc7O1cB
inf68gXUuTWuPpwv0cnE+xvwkBEMN1jB2KxKuSpPIxbBqs2JMuoTWyQj+yDVSyz9ah6SLG/vITZE
YuQKpZH1v30RKNOXWb8JZP2PcS7t5bMZMw6I0gvIyyEwK2WmK6DZK+2boeYwKo/Mg2ez4LPaj7wx
3EtuHpUljckoHUxQyllaPcJAOPVWyCcKG9IYjsHMh6c15X4YK+QgRMnDSu0eF7Sa0oXMQrM/tXxH
HSQcaD33vAaOoZytcbzl3z3gA8NWy+11NGBPwdcznnHPQBNYnpCGPvN59QE8Ys/lOP09XyMFIm2i
6re2EoRFEC4KiNGFeno7Q5ROGGmXOLt2iqkP5iswCVzJl1KBREVz/HDKxTrtDMnY+En5I/huJDDQ
3MpYfoWGR+ufd6GS5XSYzkIrtQM98dRyn8/+57a9nlgr25eC3adN6Ap4ht4bkGkxn9QXsYXKnMm/
n5hHs0CqmXC/5k1RqwvzjwhuCF7/P3bh/7iqM3+rCtZywq74ud8wbwgsisqM1Mu9mRavnZoDSrWc
R7cmHSMXGP6R48ZGPqEasmXCPQJuOMQ23hUyU702+GN1KdblEkrpcNQDfZ23cRhCf5GB0uCl4gMv
bAP9UYeBsY7Jrfr34qQ5IxM1Hl7OHGfJej0zsIn5CiHB82o26kWbYcMxdgljeaRV59027UM4YNgs
9dX4rt5ujW26Qcotzu6axphMKlqPsvUNDRrvSvye6j6zt2D/tq/S2EGCXtgG3/m4k5AnKg8I2X9O
LGHuzbhZQ8cwolhGwnvgEzfhQPpbBJwNTGylJ3ys5XEsK2dWfMqmbtGIByIQ98V7uSsKOEjgpOHk
DXPlKqsSb/bYYRfz9NclGE9xXAnmhUtM9AiABOm4l56S3O/lJ5Z06pbigtR3bv9AhljU5SUrBt0Z
nBpDDICAWfQ9pR+gJbFg0thwL6hhQzgbiQYc88BUM4Ootwc6DRvyNTOSWuX6TfmJmsG6ar+N/n60
914ei5oG8oydWOXQx0L8nWVrkQNC1J4eVfv17FbieyPyioPAmzkjP1HyIB2/z5D31LIebSK5GouT
A5ipUWSPL1S8kCEEZUtNQpncFwv9X0kdCMmeBLEAgGLzZDb3EaOH9JCMCuW8CoFlTW6tZEVoh6j8
NDKrRgM9N774gnHi4FrMnPufNuz/raqtbf/BzJwiCxR5EPqFAza9x957TrpUAHQtZmTKUbP5/q8n
BGSVXzKyn6J2geCwCp24qzA4kyJKEwNnMUVA9LVYs0FElP1SKywaIuGtmnfyl9WgDPI5Gp2IGHrQ
vzEHc9KTRfK0uHEi4/Wse2V//Mjix7oZP4FTzJZPcb9oVjEoBLTLBI8ebW/4MvYRpGvjKitO0TGC
shbAOodeGIqEv0ol/2QvaznWG133FjikgT9sxXVn51kPgVCnQQKxUfXD6C+kOhnAxBmB/OrrV5rZ
J/L6WWcc4EVfxIX9q+eIl4KWaJBKqb8IzYHiUo6+xNcA5qQDl2hQ3l6/fmaLUzRUlzUQTkbakk41
4ayiV9ADhYQbyrHJvHD10c6o5ka0Ike5HI6tVjRHAoBWH31FDrEehQQHgl8BJeKMLG9PwZBkphPz
V2lxeVpv4YUtVd/lE1DmLDHsqndfcqnQcYUIROS8cQhmzmWKgUZwp5vxM5l3ZSk44s46HztYEHBy
o8ln2VHlvHF9kURN77bnG64onjxvCVzwQZ/VH4vThHdCQQraIBYj7YHB8asdkWSt2eoap6odGOKM
hLzBuiGVqEFz8WmsnI+AZnCXYvmye9V51dIvEa/kyqFA+oPVsxiEDhsQPimNHR259Mp5KDlsrKQY
zI3gUaO+UxBgvYaAVxTOQf7kjHZR1/fHo7F0/mXTbipzgax0hNko6tQonDPal8L4LzcO7Z/CLy6Q
aUzSVOnogoAapDb9bRKnSUPm7uslbMdAV3iQd8Ii8CHlj4BxnDzRUXUcC6QJIKSCbuKs7OKLF+an
wUC6OlvlAfZYcCIc9eftcO4hAMbP+jykh36Ap3R/sV9ShpWhUrCWEf1dfM1LQXsRv6GnvAksMbRH
w3JRDilTS7ri4mrHS9vgvTJOtgru2M4L+2tMBY7xoV8d5RTwLofPc1XjVF8m1uCjr57EewVpiNGX
KmtM+u5uXQxUYEXMIrNIhqHrZhwFaYGP/gy+6xR2iYv7QlcwMhZTYnYc2mvAGY8QJbV+2Z35WN8p
pKpbCYsPnjiKrig+vOe2JPk3EJh1tFM5qn2BjZjxZv5PjiS9BAWJ1fuwyzbHGc5FU45dZKFvWlhC
FiBmjFTczu1K7NkZ+83R3RBAfwaZf4iwo1kn5wHGYcApydTy9keWAmwevWR520DSdQitRpRIfIGQ
cfMBQXcX/7SPCmyPYVUqVYu2YM+eutUZ22DIOrwTDpKYX8sAm8qehsEBFVG1QN7Zo4NWkDkhuPnR
hbdDsHLQ4BWxWQG/oUEXYrBBTi3Iwgf4RK+J7Gw3wcs6wQOhARIr1//7NIzJfT1hpLZsFH47kRbx
+qQNdvh8Em4MVUNBRo2dYhXY7n8yfUPUv5tdoxgsJn3LjQVg106n/okNn6sXrkWzr+uliC3gtWnM
RHC2o5u9w5/yhNzpC5PX88DkT8oDZulxPznr7QmM0TGdhCiP8O97byjCfKFgjGHSqeVPFJKJVj/2
STM5VstHgmeE1cHTK6CXSinlt5nYbV9TuAJbGAgeBvOXFAXupmc3kqCv/YZYmKHO4rm0jheh6smi
vTuJrxNHMCy6ReRmeD8rCU3eI2aNGL1gh9gNBTDidMBc1nTU8FNF80JKb9l3d+NzMc9EWBoXvU+E
2VL1WJy5iOd6oqaDZGSvxJ/ktUzkbzo668SPWbmWAv0WFPqyH704WLRurkRlinJOUZMYZYTrnoZP
uKezWS+08HVYKFUt1oyawnm8Q5SlWtFcvT2b0xhqYro+AOlJHrGyn3TvguHiqTT7DaWPB/7Udi0r
HIfDNN+zdFC1AEFBC60B/buX0n/bduHT07b+Qc2vGIxbkY8BYue2FPNpnOuLtiu8F8B0zPSpzQWX
FtLAffTa8J4bTIVHy66/bFIwB4x11AoaK6/dOZAR1dULkQK7UpaxZIaDMNxb+URnqAIGQmYF2TMW
4vQrGPFlaLm/yYlP/W12vtky7sIA3xQyrkff+87bwHli66dDKy52bp/cMAAZ49a+DZ/ozAooSZLh
pYsxfi9Cb1iSOIKaNWu92MuzGSJ+9uBwVBc4srAmaqB1x0dgQkhdjREppl1Sm9Q/X92SV1S8h7Pr
iRU76lHdjvh8CTR8J4lnapSCyrid3ENIK316xcmmAo/o2jLsqXR0NnKgcHg1Xx/GDFwDAV756R2z
sByvKKlt6vvpUWS8V2EbhgzMx1mkXcKQztAXQNDH5qKfvg7NTkS8JJrJoCmrtTjQuthBssvhF7hv
CX9MxlPEHdz38/+TnKb4a3W6vtbkyMGRRF80L1P53dDzOX0yynjegaOm5GJUKQvQOFuQkRn/4IZP
rOgmj1kGgZlGXo4tbAb89omXY041uMNndDerW7kYUPhlgXe/6NMRjBGIR96pAmqncZREp623eejJ
vxuEpNxhgoQZ1uNlAOaqJd5euMiaxfj+f7fC3NXf3+6BtnZ07a0TR5qX/UUCLJBaPxe9Khx4fKDW
/1NhqvvX/VHRZVodukJe04znQDMNig7Jko1pC1is8rHBoayJqm06XXuoha1tQ8DQowGazqRbfsrX
hqL+gb82xddbbFNjXbAreIfaU3XIENK7j08NqCQfnuuLy81Q/vQrcgdua3qbpZ7WZg01ISYRviov
HcXJZZ6fGDeSPeaTsjtFFnQeRPMxY85FQQnb1l5KurS5RI/dD3faBDz+2pzBT6QV4HfgqWfp+fkn
JjZEQ4tEIxjyHhNKToeXojLS0KDsPDNJOe1rz1fz+xBBlMQoQvtaz3dbqipUpArL6fA/jTigXQ80
d+ZGrxLK4v8uBkP41Q3nk1nsb+zRhGYrr+S6khrdcY0Tq2k4F1M+NkewgOFcT6cmnzGjnlvIA44D
6BMNi/xzfgzhdJL9zVSX+/YF3EHEmiPyV/miMqTrDbf4FUKgDj7g/Deuze0UdWy8sKOWAhT1mx2I
ERr/aEWZjVsoJ1zmIy5en8hI+Sube9yQ9AxqWDHuYMA+sSsx+n0xem1hNfbCc+iWx8DOpk8ZkcJN
x1T35W9DyaWBaQPgY916WhQLXE3nTsAWuZ2NQU+U/kSHJlveLtALFzUrj8p0mDUObLciVWdPZZEM
BkyH5NKF/g3UbybwGbD8U0izPsewG5nZlIXSgr+Ux7ZwpnJAFjWxkJAsaaan7FH4Lke3r9S07xyU
3iFuwdgwk5YwkNdSi4htBzwSaLG4xbaV3q33tZwiumXQCTU7QE95yzlZwDZRoMuBrsmg7q3XqPti
1tpuIJrKVNdg/hDQO7XYRkVqKL+X1UqJqad4XisTPP70YBF0YdvricxXCvY4gBF8bzmBITcY977p
rKuIOPsk8iYN1T1sGLcUj0le54h8yoSqaSxHlWgECDx596M7oA6IXAfpqcizzUtFWjt8vOryoDDq
DJUj22c4Jk0Aqwj+XwRi75fly3u6ZmrrsvsKkEsqiBMn9P0khp5C0SDfnSgx18U16xY3xY+7P3L5
VyzKXYBHdmhgnRk43dDImnQvBJb60770t5SPrAB1m1Cc6RHyFeKoFU2+TxHnBDyoc6NR9fAIoa/b
Gx+MaPPeDzrtOVv9+S4OQ5oh2eb4j4FtR8RNt6B4u51S2tjWjjqbwCrFF/QP1ctLsiFqC6T70B89
LLg2fLqrhbYHzOAdNBpQETgzeNi5z/i8sUXux0JscFzH8KctZ31DujlMW4KNdFQWG+G9PLZuSR+j
9y/tR0xe/Q/IpVZm0E/cl8W7ndKvqx3u6cxoU5uUmEo9G87DBygn80NM1VlWBCXIAL0Un6j1pA9h
5Dm5YkGNOv6yPaQDxcB6q/sBTEVmcext7Ft7BNLQ+k5sO/tw2WbIifLLKxIC793DUNqU5rPp0DEt
AujbznY++CSo7aL6LXSuC0zP155Fd5JJiuu7JJ7MLj3hc9l3TPYFtqMe7rICuHABZcqM9krH3Y09
EM+U5m1gTnAhYuX913KMTEp1tosXpF2NhYwlNKHghX1ad7DedJNS3jZggrbDYMKAjGxTALLgatP/
eIAyLJhb+1etOJ8vLRdva833doHw2xsqUl4t349algyVDwV7cGj9zV1QeV6+uI//46ij+RuxoXuF
tPAokfIaqDLMoMe1sOB6a59ONqFPfyLN02R71JVFgrwkSrVNLrmOS8VgVN6K1flvlNMW2Cyla+Z6
B2RAAxE4iGVuASfrVhWY1FibIUH7k43g+cvw7vcD+rhu1kL/K6BJeSLFshbBdI4gTBO/agKNYdh7
9lHXKr+QMh4mvdWjip/AyC9+pGq+eVOP14WfYAbUi0EuLtnPxdQ5s3qPxLzbITHNAGex6N86112E
YtvNEi8/yanHtmXScMD5GEkbY92sT2e3VqaVpp+NB4i6w9b08x9aOl696wUI42rytmNcXCkrm6E1
DU5lz4189N5svsQKUV0PfQbKsxXFLTLYrnflDtplMFrsu5H1JoCb5SewsJkOh2rn3p9NMyuPTY4h
uCvvvA9ceIo/ylRBz+s0qS6/mOqmM9plOd+RrbSZcw0RDY9PcJr9fP8hGWoRlwTaOSGukYey5GLa
408e5Ma8lqSRjsIAQ5Dt7tt7VKl8/VA/6NgK8Lg3YbUJbJCM5FsJiZ64PbM7Uy2zw5ZhodF9lmdZ
5KTcYfBqhDRmf3+HpsUenqA74NEI7GWUtV8IOMH8oRJ5sJrL3TBO4gBNXLYYOpRrQCbo1cn36NwM
77UZTBP9DloHb8xZmdQC8yvCLa5NYAxrV0xAY4ZLN4AY2Ch7Auu143SL3zuzOu/KX/39XGkuf2Ks
zGezQZo7QHqujJuXW+kPdefsDyoHuXtapbk356y+PmX8+lclPo7upaBIBfOcTWtv9wq1pj3E368z
LWaUhaoayiOYPKTejSBaC+RiSu+VxR+8lYYW3IQUxA6mw/TQ2rc8NifUAB7XO4liKCNK0Tke3RZk
1AH1sWfLzzPVU5aaFQY66/nrD6A8mCqM/5VnUbtfQx2WUhum0OVefsuvl4tf+j5/nsNx/tv0eSXG
uovufaoA5Jt4MOt5WognU7PB+2BhlSa0NBGSzz93mQttSSoHpH4XtYpxzswbcddV0ePlDjwMPEPF
dd1LE7lSzSlMm++qOxWsZOaC2QyHxux9hFSzGUuQQei+yCMlYr4MSH2z8nu9I+IGFuMVmGY1/za9
dBvXGIqFsyrTs42NJ+I3xjBjvkIn0UTjPhAzbLTnQXcEaIh8Er1zd2DNXNd/8p9JkebfkA3Y62pw
vkwkLuegdpTWTWkVPcjCKpd4SwJhaLEoo0C+5z3QuqV8MGg+dyZEle/58sVn90emqaF7wUbdJ86b
P6MeYi1pLZsC4CD0+XBj4+abh65L5bEp+apayYK+6SBJSxpQUibKA2r4TJMaUFh5G/8KIr51r+0l
mXnq0VnaEca4TsBNfLnJF3aXiwsEmKrVyiWYLnlPTaR/SqVROSMKV65T2qleCN60UVQJZGWvbe5n
DuAwkwUbQOy4udgxoeEBKtZ/l5qulsyxthE4viRaDJMU5iFYhMiF13VYLrHqSCmC1jQPn1FhJVnm
Q0q4STIqth00W1WYhGbuGz9wKJwSolhcQzjXXmPFpl9OdGaSXSx01Kbi45Yva+VR81gkb3YHeR/X
QzhmNAd2iX6qHNO8EFsLrNfgfQ9YEDwQVIGodnEljYnybuzue8MNadk0gHVOVCk/A75ipkF8NYMa
z0RFCLXJjQLR5pT2sPZN+JwxxhzHe6U2dQOcMPTedJOgY6MISZ/uVV8+Pi+IRQuySFnbbZJ12S68
E3KUxXcGvZMRUVB9Wh+/p40uLwKFCfJwpV+zYSjEZcLedB5LPLd/2kt5lN+VfUNHSlbcQroRcGoy
Ih6W1lvmaE5fiQWQQzkX+/pXE8la8l9/VfGSagvsIZr66Euf8CgSf33qSbkpo/yTCrC4+iQ+EEhM
qO3qYFVA8e6cBvCKgbz0ZTDN4Eipreix/VI20qki2qJbpoVdC1SHpXH9c5WUsuf6tt3BjEnfJMFh
hjvgTen46GXH0DPvtWh+1sgStDZTaOYR8GH4nXRwr6t13UeoJeBrPZRx12ZCiR4RJM0ju9VR/Ht0
jjqkg1Q211IR2UV2s2xzK1ZDnQfApNHUH0dkmepzBegs5G/h09FyVtCpkQGffgdUKzPKv+Jn4/4c
H7rfEdCxAvBt6msdrebPbkjNN1azfabxurtf6Y8N+8So0PhlAuOdilAeXRz8kLY75LznjDhKBfn8
4Ooqr5Sdmne5k4HwYbiKg8x1cZDQcddby+QXelCo8Mn4nm80eeeST7VzakVoUaA4kFiBRwve4FQ/
5gALOzTLEtoWqbeDjdCa5Jfhm6KKmMD0xiD9DJ8O0+WrXRwumEWUC8JAfSVwV8YU6VgXsFadpgf0
0/N0BJSla/2J2EtajE1k/gdKspBmQUdf6njD+q/wAMHR5CXz38R71YWPJn0dueeA0sSLA/Dy3ITU
oba+wBvmScJj17+9UkhjUL5SHfgRTWhLyajz8PHigh+P+NgoWIy+zJSa1CTpMRFnpt4MqtdeL5aN
/OK3R3nQMAsTyHALKgVRHySn6E3mQ9ubFj4VTuQUj852ibOgsuCHCEIValzGKSf8hRiK5oZiHtwC
R4cxGg6YQbF4zMnFOaai0ovZVJSNeE6KHOT2tsfJ1qcutWz2ut3LVBM3J7OKZG6ovKRfSLcCcGsq
zZHIfmbU8EQQYR8hDGUniz5mhs+qY181AVb8vy0w2Juqe0p9juHDsMN1Yt39AwiC2fhp0fk4g0eJ
TYd27ihnxXu5wfDnbbBfqnlxPRZMqHA8W+d2AtChrAZUu7RK1smjVUgvoKn3KtbPuywraL4n5pHv
PpnNRHOFpXh7zY64DPG01UxxvJjsM7tyeCIjwKotSghG08FW4dvQQh2dpGhhcW/uttndMGV6IDtb
huQRdeMbViLycDnHZbR3hahbb+F0KuSuqMC+9LqX/iVNgfxWDWORkqllQqvUfbXvuXsqEVglVelx
YpxBgB5jpR0M91sdYSaNwqJLds+3gDHhDC6/jkFBAmoPN1D0p8cyYSlM9n8SHWKYcKZZw43Ibsxk
UTg0w0NO2Zrmqi5yOL0stPAoVzKpuUpU/WinfAbTYknUzFhD5+o4eg3/t/P00FP23jjNbhn4hNo7
4pVWuntv9G3QmzMDYJXb/px4rbdprtDoRL6KRjkBghVBHNgtsCLbfP2QE3JYE9fh7YZMpE9wPrxl
NalwtO+K61otp1NW0VSXzxRIBLUvpZFPU1FahzSAldJ1tq0UQHoejq+ctWKzDAjI7nBQHEoMRtml
WZChN+/huQ5q3lFDrtNOkZqwZOxA0MpkGWfZ65JWaNJOB79a1VKxg/cW63pL8aVjidngbpLNk7yz
UH7Xw2Qd8vzBDSTUXrEahxBRtUC6/k7VGqb6mi+gBSiA5mBb5ZVVIN1nYEuokZeng/qJD2PA3yen
YrakBuxMDTJmZpiLUdN2FqIyDXUTeQeqRAmT5ol3bLNxgPp0hMZPK+Dtf2Q8mv31Ot97Z9x4nR8p
QoqP+kR27j/V95UZu3UKL539eyiJxoI3x71A5uFUVd3lwm8rRclkDChgraN7T7AAv5DM66WkkTRP
7xzJcRH+waAS2yJsdSmpMAXqySuFu/ZndVqKMteWJn1pmH+HLgGkQlJ5vOQPsy16zfyDIZcxivR6
oxX6MsZFv1PILZ6Tne13N5s4pTNxECNRomqBLxSiemxuToJEtoEjumLUbmPlx9y2YWFLCEdTE9KZ
puj0MxL3g30jMOTuBIG3aTmXehzo4t4zR96xyPPu+cn0jxWNrJvz07gfDl8RMstjgPfFEZs9vg24
jaK8Yh5gMgKF8IZ8pO9mb3jCuoEqhfwREObFIefUaLmOIpgEOJLFfnsOUGkDDD5BfPGtHTG/gqtr
H6TeI9RRsthfw/gr5nXtVOid7by++ZENkDt74i/9TU2h6lhK4iXod7F+FsxsaED7usb7QR8k64sE
85pNVqb1k05/XnI+nx9QQcA3mrRCcpA6vBaGmPd0m3fZexNMqDRTb5GOUEFB7rJLmcq4ggNDSsZG
KQ2Bv1TVE4MaRv9piagqyM498wVNn5YcC3zF6gUkFY4LBduzqEamIFDxwUajZr/hLph4ch5s6bo+
apHxElpkav1btfWh60vfnkHjSpKkkxaRtj7F6sbUDsSHA9VRL0oLHzwYJFeJQ4GTiQBD/Jy+lNOb
t02SHbd0zezZDwx0g9XK5QFqlhfm1dQhFOvEzZcASlLREHSAk0XP5lT0i9mlmnZX2w+NFx72nF2o
BSH/r4M6gCsh0Er27LWsWU7kzwP+LIaS6oyfeW9rRQpA36hAPXGNOcsYgWcWw6DeSZsC5XxAJ9nC
od3EVOJvssIVVY9pxbBdi59ow99VbaokG59uoLWOPTvlrYVI3ex9dQksb2kAmvmWoxdH4gNjT8Bi
V9vArDyFFdpN2rnNxPsmvjOfVkR9m2ftRYLTdHClvOoFfKYD6NaNOIPr/eiX1LIVYOoXxkBBzbf5
UEgXinpEa8sd582acMbP/wCxtpVeujOCvMCrSMXFUD18Ot9AcB1p6tdrWOHOIbkJM1PyZrw0TjAH
wsK4yA99c+QzxvACOdwClRvQgvRDIJBq0UJ6EGy6G8BmHjWD3Mhvb5cA/JTA0fXYYplgVL5ZT3c+
Ex7mmrVlWikBxezwUHk5EvWheCpm3MiSWVCx+jAYxQ7zeOZPlvYBM3JIvWikik6yFhjN0c2/+h5+
4QQdmTJAmKdEoMu3fUZSLJGaoiiW1q0bR61n+r9KwtKbzIR5Cptl1shlUd8hd65D40PXyaRBsQkL
Lquj1w9UmJkggnv67TVmioLYsDlT5syJArnTOBM8hx3TnEwmGDY5dXSgTPnR/PLP2Jk8ihiI3vDn
b/cZ2fWR8/shr8LclS8zs2YMTCV14bU2J4DiyUXJE4NBfzY4GcgI0KDpJ0HfXRmKVCGzbemQ6wJ1
1YVi/OCB+3HNLtRqlEVxCP1ModQGG+qj/+LB58xFf1J+o1loVabuobfVqM/NO1+xe4VQDGtespnu
lzmyj41tjNthK/2YAHS+NhpquxFYq/H2iO5tDG2wqqbDTlz34LMXUot9OfB7+bxzg6G0GeYSrtKH
nwfhW4D4QCpiACk66v30fygrfsSEfweGf9+DO3NY3akAFtktnl4avfnR2YEkr6XXb58kx8oUW4h/
rYGY0Cn3IYbWCHqA90mAbgsvvLJU7msuoQXMnkjbpB2/6k24+9LifxrJnFTl6FZwtZNr3YLew1oq
HCctRpgBA6vS+pkhGIp6YbsdjZe3HLXVWVJ+2FRr1SavbaCp0Us90WqCVjTxZIddOR5Qga/Dfw+T
c8mTP19WqyJkrHMn+RUel+9oGj+B+k6VCCpBT1QGY2f/GoDPBL8YOrD7E0/mY91wlVr6Cg0u6vB5
65m9LImvKwyAd2zVhj7sHfRj4BwOjgVobRMrl0Zd7EK4yNkCJuXAkgR1qCk5ykCDuasYbHvhYpfe
Gl0oWOtjZlBs7h/RpMNxeu4N3KdpufJdcKlhoUoq/PqrSg9zRvRas5hd50JlBtv/g8cO9qgGBkAz
z1x1kuQ5WQQyRoErrrK+S0SWJ08Tfp4CIlv5sVxqPNcLkSIcTr9mUN2XUAnHmB6Ek3Jh2d7tKeqK
Kg10GewDUFbn460ZICvk7VFkqCc8T3U+dTUOhUO9XikGEb4sbY+gs1M7BM8f+gcy4FGqrMRNA5Pj
IY61KIMf8fs3MEpJFhuMMjJHHLxHnlCweb+2KuiVepmjjOfEBp7y1yz9WLblSmTRAPRzvf0lxp2t
NzODvT0QIuYypcvjEggvx05Q9A1aq47RhxEbMqo+TYoFDr9z3UflD+QbAAJ8hcDeQko6PEQj+hdK
Fy1ntkcSmJL7joyY4o2dOeLUGr95OoEq7d1d110gBytkKB4mrOSyhBsyqxDvuNkvkZIvDP85P8X0
koFQ92suzMdGpTQiupCcah80ux2+/HrS5ElZe2e2Gv+M+U+GQRqFqptZybJvyYPcCIS7MJdMvmlg
wD0cpH4mrJdfeTyYCxRlg/cTJ+HekAgh8KqY8FxRfIxERpDPXeYEs7HRZ7CIwzjscPq+UohGdamC
uQfoFuT+mJ1TV0+mYwJEXoejXogmZqm4c/RLhCOQEfHsE9f5vXnImGBOJi+Om69qf7eIoBCdI6hw
q2VRRSlWQ9Src2oDsNCYcG3Dh8FjBdwZqBIFvX0PFJGB2FZM83idmcVoN2C+18StCJGmh2crxXdO
I/xwCtsIMLW9Siw11fhrE0HkOSvp7HJa9NhYR517QrMrbmi4xbwUDjluTCcEULo4CSoQph4tK258
wlgTNUPDgKryP422laXUTD9OYlpnt0GKBajn+lTTcYy+LT6QHz2AB4O3KRn93cKlgffgpIm/0zd1
1u9etu+MmTfJRTl9bf9fOo9eBLsNfwxuPb+LbS1sePTaaldWSk50itnvDC1p1pcaOfAc0jTlBi3v
k0rusghxJV3r87VqQbEKSNuYt1SCtbNHPYf88h8tjY1HwEtfh22PbZS6kURKqNn55Zl8lIHiY800
9sGtonZkpXdGkllZjBBpNw310SW3bIrPW0G97naOMKMH1YmW2Vb+W0FXxT2JlloqAM7XHokGW5DO
uz6+GRwlzrhTpZ04liCUAzYs0oUYnTvyaLtP5AKr8hO1oLW+wIuC6faye2Yez4lH01CDlD56yTOS
joKKIhmidEImK4tmsd94mjxKnKMw78tjp1EKHjExMSLJZ4pRlJjRdcoWm4DSlBHcWcpKEEuyv94x
nTbKiE6xPwPdspsJ7GKY1byyUEGlj5K6YBSjv5kUYzXiUHjq1eb+pxgphIuVnONSKaA8413FQuHV
5cVSW4XoiGGqQ80n/HyS/ewU+53REHjcP1p043lCUhwEk6jSSe2q9kA4tbFaUIhu51gLRF23lWdj
ShL4nY01yHtjForK+Yf8qWJzk9rpx+VTgcXGU1XtU+nayrH4J0o5fVZfEHLexA0MvYfjMRmPzgkD
M3CrZ8XDo0o3tvK3yOaa/tvSY1zCxc39iwRT+CWYl0rlTPFjr/WqiwDL0e8AVHqwfnQuaY5/vVHv
X+zMds3RYk7d/80WlJyx+iZH4Jjj9n/dsbj5Wy18o2R7ZFMi62iTyRLFvWywbnYuooYfOJ9x9ws6
Ct7DsB72vAJKhKouqHoY53HXlLbzFIs7Q97G9+1hgXnVzP2W0rkG7qKs3zxd9PlzoQ8rv8B9g+Ra
nDa/WxmR66/3N4g+fOUgMzfpgBJHUOcbkPeaXY5DSoqeYgSI6AjgZP9d5FfxLS8zpZ03cZkPyOFm
AWnfzC+iTHqu4uBlsQvIax6dCzUhOCfl4vYO0pNC1//eRy693A/vf5wwfi4oatwIN/a7WbJPuOeI
gJOI/ZOWNlCBYgn57MaoHgHBkQQrqfUFgNMRPajG7/4npuoE64gyoIETz8p564n9J6TloFIbt7H5
tBJpT+C24yUGXpKeH8ydBkHmxcC5e74+HOCaMQ2en8zegEAzogwQfeSXwAed9uaxGIeKty9GvArX
8BNbfeVKWsrBIxM0DLmr4RwJHFic08+ucxkDUUX1yCV3+sUNXp9g1DkYAxLXtdZEQfHwBvNgJXjx
Q8Rq5EOL8Auh8lBBbPKDCAeVEqvTN8G3ofQYYlLd2rifblzvDgc0NGxWr5zpEOCxgYH6FCgr3JqM
pZ8JBJODcdb1+DBAoKP7QxepNfzhPvcnfUghn68PIFIPI8Hkg80ahRz0KfP9DAvvZy6XZaxG0wnI
usA3gnS+lqQpNB02t4z1MMGObM5Cq0w0/iB4d1KV40AjAydQ/AkpGLK1xw29OVK5qDdYbwBK7w5o
Q3CfYOlPbihlAWSC+5/8IKwvh4cUviKSq4SiswlSwE1sUR7NbXHRlieMyxqCOhws0Rtw+gLS0Q8X
rLz0JETYtarHOpfME4r2p5nJ6jwhDr7xo3OO07Nj86S3ciFveVD9L8xh0IRCp+gLES04m53XewS+
/K9zbXh96Xtyyx69FuNqRqFgWDN8FARPE7Vbj44PWSjWlsuj0V3qcVcaQyhMKO2ZE08dGa8gmeZH
xdFXlmqGREYKI+SiRvm0CZ3nezwpww3PiNXVwd/tceWVb5xQTCppH0CKVYWnqxZAby2zIgax446t
MqiWxD8F4lvs82Zb+kJRRrdLwmPVdN9XmY+V9PY3Kc5wW9BN1NJi6Er8diRhHDxoeMxDFHesXv0Y
0VqEckW/te+9omXJjJXo5jeFc+DQLhAMc3yOjwCrtnpVj2BDAyn7WYwxhWzjuRtO+L1s1i4vwBpv
NkymIzwwCHzdQHsEAUgWlJecjEf8jR4wEm3lgz5n28kMZc0rLyu3ovVu/1HsSmPA4mYZd3UQ9LbJ
QPVaB043VjdaaxrJVNoC2nJO5HaTmeZOq62D9Mtj79bTI47hdJlzXu0hPYp38k7+g7jgF/hTqPDx
T29WVoIcOqmbvinTd8fvbBcBIFTy2027RzvwJy49wEiA1DvlgHbAxXwFBlhLQ9p3XMA5S2JG42w2
Db1Fav4HM/ZmrTUPDyoM74CFQOpF5aPF4bw9GwhjumBtG4QU0VRkP1rEn62hvZ3VGZRi1q2EybZv
R3WTF9KPwP2tCIV32TFOUwBMTkxX9PPobCOJca25WjjTQL4zmj9l0ogYX5OlJc6uJbJn0ft1gCu7
XceTR9pghJnHBc8fg+L+rSDuny4sWs11RgPDdQ8xkB1p3N/bq/aizct8MuTgX3HFI4WIE3t6cZJ+
Gw8NkyI8sPBqx1+HOQk9hoblIVQGahkPEos40gnnlUKwX6Yi/clvj5U7lWNmMRIpm05FjoJRxUxt
byJBcsaW0OiRsw25OCkB80ccT5PTYD6e69i93Xcpej4n2W29AxN8IarNafHi3TTcBFP2iWcvbGgf
1ondKppOi/oEy70X1M7phTN3VndUkt1SFcG1yeomqmHteoxCHbOELqMIKi30IBVAhudtovOW3lpp
U1G00yAvpT4AwMOMqh8p+QZ/gJY1xXr4I/xWiTbAwOLlGNONnL2sZKWrdnYR5ysoDs2cRSijL1To
lAmUAFyHwMHjTLbJN0sZKzm/FCBKPGmzYK8Mi/XVGAkH2bAMCrVKtZWDa/HSLcZpNBdbcZCetTze
fxndwSnj57gqVIbZxkJSjiVpoAL+OzdhUIBQRrxnjA/FqP6u9x7HiNznBxlSb+imLE69f+i/BKzV
M1K5em8LLWthHpOLkx8dwtN7NA5myHt891T6bT4A8wjjKS0tZEwFggq3CoqQExV9q1PawhCBFHca
+Dm30nNmf++05XtaFV9XmSmpX03JokShc/1soRKXRBe+dBxmmW0CmKu/OrDsrpNHr/oLg+BM+LEu
TZHDGHEQ3u9stVH3F5psN4KgIiTF2CidmJgbqun1uYlgqekTid6GYdLj9uDbarZnAIK3GRSE2BuV
HCRzqtctfg42JwtcYRfEOyL1xB2l4J1dAocZugKqzy2CLGZQ0ng8ZZvlxpSEDmy4D/o+LyMZD1m0
2tdHUEYXZG7Fo3pre0SBpO9BNygaT83FMcR+oWUJ4WCSRkmKXdgeU2Z+X+8uT48e8fQopykeuR84
zb1kDRJFbIk38h+IcaPu4O0q/PJegc+gHeDSDGaPRHQl8FpULXcXGaShXAHDTF/BJQjhPyBZtgW/
0skF69FVWUaM4nVkCpQZ6nsSHaSpotwYB5HqP1cLnDNrWjJwibIvlovdEjCSKndEYWj4d5r38WiC
PXl0Gb5UXFzXI/tw6fYmfbd+zX5k/a4IKQqGtNUhKkH0Y1eLVAi9IkxAUo9BQOmjdQ7rOa2nsgom
/O6bqmlOT3R+g51Sb6somVDHMDpFHsFIYGuLALLihDUrIB2wubS8f3whojBfTfyARSDjAPUK9erX
eHNth5hVKCWDRzPtmO5bSh6J3IJcElJeLb0IDqCJn2zrinMGfSsdtoQPHS75H/oV4ePLCkOWpbFz
MFiVqnUdb6Cs9Xq8fHUow1xfLwvIx1xHagizC0sOOiJpWtUF84L7pbFOZoqM44G/+xf9wRIRnUJx
LB9D9dNGhn8hdJSeHBGp/iHkYWwgwp0nc0N0qiuXjITnUMNr2BHYaw+Fv2NDC2p6I8uy87/FH6bs
y1+BE2g3RFChfFQLdAZjtc2xAFMt8Yr6HECWGJe/drNypfEzWvOJMHuutcZDRWUWnGbNeOVJIjsZ
rlFdGNdNrfmYljwAfxRs9a4rQVemCuRHNUfhl+IGsUb4UecA+FmAg1GqYcBoruqdkjeO2wkgQmsX
aeBv/futRghmQWJE+VHxFFpOgWMhgruy7IMtO186IN9Qxuxd/LD9mWv76QRgRtfwyUPDch/VPKH0
4Y20OW1SfO059GUDzz/HgSjDbJbp1n0tjLf7o3d7c9xD3Yg93dlSvMt9f7jgP2rpVLKVjCIN1oxg
OXOsyGqTri11Ek7F/Xr+9hzlKfPFt5drqeIfqvsqpl2cznHq5Tw8dXTJVKEyPsM9cj8b2iIcLNIW
6OjWIDETiJkXYHOoogtrem93AHz3w2pow9qiJpWYObmW2NjHiqG5xMIrDE9wUM3rD0wtTRKKKEB/
OdGBSz8eWeeRHDenCPBMWZkz8f1dPOcrX3JXjtyACoRukVqUmrC6sleQxq+s1vcHVbghIlONFqn7
cYUgO3IzhnCIpAkfCn6W+fXpzTPh7KIyDYn3DDju7rGdfvz9AFWfwUQGa3gYEfgFIANG7t70/czq
4Xl8LjmOHJpnGu8U2j+b4s0W+zU/O1w5wy0ZPEn50p1ctER6+0f4ZtWxCuPfaUxu6JZdIdLF6r6M
731hnsSNkkWFi2Um9jvtoJO+wIVLj4LHO6KYzVejVU7q1UJ1IC4BGeax4Ua1XwIF+E5cK5dOA384
qx3zZENxN6f9YQMc2muwn0Lzw8ztOAMK9zHZjzD2b/Af4QY4HzhW9IQEcpD85hujEH+8vF3Wjh0i
FdIJlNdNM4PI/YD2/CNlf+onerA+xuGr8HuJz9IG7Jk6ftK7HftEXnqcaW6nDFftIeTfW7vrW8ks
a2rNA3k6BpzaO0ZgO+9EN06xMePqR4z+vQEHaheJkKIDyDH0RPH+uyg6Zx5ZUCLkFQ1iNr+k5sOs
3UhTtMSNL1dRbIIDRLexhroBupVoHLqCmNRd5WJnItxeOsjHNILb836+bDOjHVwefNVw0YKB8GcG
Qjyol2ItyvmJuTybU+TWxwZj6+o/24OW4xj5rO4uoqgrlZxMDv3rw2Rngbbak/RfgLYuy6jRXDVk
vU4FqTV/CfSoQUFaoDldp25dLS7YO8MYXk0N+RU1DCQLi5jDRmUBCa1R8QYZ/7P3F2eGM+P9Ci2B
7hiAe40SA96fAhbYnqaoQr5XQ/zZuQ2xtyvczssSozKC6hHV4dIBK183CtY7DaaQjDrd+5nHFBRD
v/BZHSsa+wvNKRqZI7b++SapKJALaMNn0OC7SdplwnIZDudaOBfUCv/q1QP6Cd/TBQHYSQQN+xzS
yATAA5BYH0NVentP8TcsHAL4SHDIJDhaloNbERynhWzVSvNruERKZ8ZqI/eAxDHikIPlaDQUpyua
KY/KkIqpVsPnh8CQEStaZ1cuzowN6ckfL3ydqlx7/dBKwdfcTF5J4+nmARKiGTX6dLlz4kYxBwbZ
nfxFu5PKAw9fKdVl65ma5woxpQSqiXDlqQl/NXNtzF5aFo0Fuo+bScbdTTwkF+ItfXJwkG5r1a9+
8IrMNiu+hOmsEOVOu8wjfWCxxZsz8T3sYRxN0XgJIuUZuv9XvAoMJZfQfTjxrD2Dz9JGHc+cTuFx
5wrVDlZhv5MsDsUlMgWAi1tLUYuWrq8GxuBg07wJ48OwoN4mhT9rx+2nNv6efArcfTZHefWlXK8A
uAzNUcn1x8FjBfNxQXVkBfMCJkFemdO9Ur18cdZhxBFKctL+Yon6GD80HfuanaXKvGNcimDz/Cur
xq3bV3RabG1ydMbuG017qgXoOwgtp9odGDx2UdPMczjoqLv8qkuac0lWTf8KP7mlDaPyKbMkGeLh
EVHKNo+0KUx0u+QbGm8g2tHjfdQYZvKbrJdfZQgPCAloahCsyNF4mLM/e5DRgbGGantEp+ca00Sh
ypkcgZoBbiz0zw+1N15eEa2x6aUhsR+LW2M+ZGRse9jKHbkrDgHAf6U9lLrn+49spYw6XyeOoLxw
zvGOK93sPhZ9hbiUbQFwleyqwDdNsHHg7ekBAF43a5fyPRcJNyQPC5NBGISELqRoWE3X9uajFmmM
er6RDcm970H9Ai9DKEpngiSYJZXeJtywBAQnTDwc86xFORo0kdPyvqhtUu2F3fau3jK2A+mAMeyw
Ez12pYV2jq9BQLGb0luiYe9JrIdB61c3jqt22EfxMqQM6vckDKzKaEi/PfTXApqf291R9FqEFe6s
V+rIc/k9WERqPU9IqZHbLjjcznQehGX4yWH7+SsHYlUGTQRNqcG7zz6bB4SmBTGOEbULsHpAKT5e
fLmWK+jnaIpR1A0N3fyvTwo035/wJG479pwFAU+lnC15hmNch5qKBG0mxE/exbSCV7i0EtE0AXJc
GH2KBk0SxAcvTOilV5K20MPnbr25skDpyt0Z9z0/CqGR07EQU9pO9/cpKQrwHsc5YdO7hkoTu+So
tMlQLskdvgVVYT4U1s53jf9IVODM97A1l678h5jw+9qw+Gs1SC39MpciCjhg/3iNteYvDi3EiZot
cdrMdk63mtP4YBFHEGWavpp9JU2fFVT5kyonEOeIZFwij7EgFhYuDbEVBLzf8J42s1jecw4Ny7It
MIipIBzasz340kswmmGU5LhzWth4V0TMkPvO4XAcrFJZUehcOnzmTRiBcySwVgsvKJQcbC7LNU1g
6kZSq/WSUNn4TQnX6h+2mxm77oOmj64tapCbwEY/K4acRgZBcaSFgScwUHoDKlP/CmvpYS9Fy/Sj
/XB8C5VSa8hFE/8yx1ljZ+VM7U1wKQ7WvN+QcvTSI3foCusn9OrFZSfRXCiyek1Tjib07Ir1ZyhY
MO5bfvb8TMwLpmRnpAgsfLq0ux+hRumwxJPdTvxZiPxhDa88UmqNvSuCry2hzdcy7Xr4h5F+xa5m
Nw81Rj0vlso9MeBfx+PwKtoixWgH72hzpMnbgm7qapKRUZSy9LUlDV8NwDT6PlbPVvf0fAzkot4r
eaZM11i/4xO5L3w9LWFYdmU8soNYpaqO9QLhW7unp7GwrzfrJWn0r8QPZaCRVbsZNH3tO0t0zmuV
dhA37bWghcc5GpaEeg5jt/I0htJr+VV6zgk6a+zAIB/8mvHBeWMPu8tYbxrQ110FVuSPoHZ6IIMt
8sfK0ABjI8dJbc0l0NrwpnfzlWD6NkBd4rHE3mKmPVC9mRZwgqR4rkSINO1K4dUKf9CA5DLB6v11
FilQfOALKF0CZLHTuyQakroX0Wtwrj8x136/1HxU7K5G3/pJUiIMi3rES0Hd89HNkIMkLXIz0sDJ
JvEJiSEF+Ge+XSDA7OhaRUWd0Lt1YzUtu9051wiLptK+YK0xU+MzauH98BUSnQN9huICcgCGJMDg
43MCUUulqXE6OOhtJZvuBjyfmi3CM9JHmnQ5t5tsYFO0G6pvn7xdSGLUcWSaAdHb5eo4xY5XOcAL
WIJPqz9659hX03ayw9Zy7FAckfns65vqA7FpggexQID+iH8k1TC6JZgml1FXsL0S9To81yLuRVuv
4If1icegLWHTefHjy9uStDJFxyIInV5G+SDpv/ZA3XtXU4lB7ucvDdlI0BNznsvdNpYRPaYh3WkW
EmJ/hj2n/n2S8y4ywz8HrGhdgD7l0YGsV74o4tSNaWqNviMgPEuTOFyXz5tIUHptDkhHX653XBh4
J7ryVMFhB6je4u3OkyjUfGomu27VmuSmV/WVP6nNIW+9sXx82f870+md5TSXwjziZkeB17u/pmxP
xg3/6MHvjCsE7vV13M9ZAsRQSTZrhcZiOQZvgNZZaK6aGYK5Naik9ruzZ7lQGObf1JCgbl5tP3Xx
D/1FswdGJ5utoXMBSUmeXjcA5vI0O8MzBrkD7Jns8GCl+F3fX4yRTB5c7RSUqvbDosC8JiS3dgGF
IJReDtYFQXJmrxYdzM609Y6dXMOgKW9pB88Sy0ucrrymJp74MjazlbIEeHNyWHtvLSqkXGx3AziL
hbBpeGFcgUk7TqhGJdiaBqtpLF6dKaGRvyJitM5JBZWq2N/aqa11uFAUQRpdNS6DOrIZgM3MBHud
0XExksuJx3VYEiKYeKkw6o4OM+XtgEFhus5HC61G611gDonNjZx0lBbRbQx8HVNmrYKx7drDpDr+
FxLkepnEOHYV6/PN0LW/QrwhZjVY5dqxpRK4jpDLN03QrVBH0yEr7gDALHUm7G1Cx26N4PXLpQB8
q+wFqzXcB9Ctx1f6cttVKOPvZavsk860les5/6z31BQZYQSQMmK4AaUDpo2Phf0qsvJYLYeZiEF/
WhYO5xH9uVv4BjUXqzcOxXkwSTPfBpYgS9F/YrESTg8jP6FWrVfVAsLn2wnI2KQFTSSwhmqY6TWU
HZmZtxzHix1kKV79jqDX5L3AidHLaW/2O1vpdqj2BPk5qxw7OQuOpWwkVaPDmcLOYFCR5LYKrrgW
HqpPHLuaXNW38s6APo5f+POwkwgGH8clsG2YRYT7h/Bzbta/YMc8ATC1jyrtqAQT42uUQEYMsGT6
C/qXJZ5tDTcjNFcjEPHy3yfYQwTzOAGjMY7aBUQk1aQrkqnIyryIG5SnQTCsJryVLKzN2pmpbQDO
6xN409blKSZ/8A0IGoEzsBXiP2TaK3TpLhwtTZ1Bh6cgiS0DnD8vjkifGDumCoTRyzbLyPLU/oFL
DMp8McKTR3NnE08lHJZi5P7kYVbzNke9NLkC9f0sE1kQLwg2PpnT1qqvbKUT2QR2YcK8dbTXXAQD
fEHx/kICUfvncy3UMK/M5MkLp6WGog79fv5CeYPwjykkkfJGVu/nueVpY6NAi6znecaCWoZB/29f
RmfhSnmbU8hnsQnhDW3MYJxpS4HHROu+Nz1RAdubnhVMZ0mXfDlt/O/xMMTJ1MmwmSKYn83Fom3d
Yb004ZyBQvjiugt4it5904X+u23ksRZQqdMlnPXvHuBsReJDoJbxt8mQgHLEInV7B99olFCEPE2t
WI4tuH2KVnYii2VZL2KRuyFtn8Uir9sw1UZyznIlatbn0zq1V00oHBbyWsuvGQS4Aj51skdAVkdY
QUS+cHm69cD1mXTuzS9VGuBTu/KWBk6a1YY+7CctywC8RlVW45mjhce83kYvjYfS4H7/9j+ptzj/
74/5K/hm/BUTXlMeh0ECQT7zOHtaNqOLaWGTcCeCtMD7ZLpyPCWKGKrWyYXyfG5T3atqk1htalNE
ST8zI+VA22MZurL+QSRq/69Dy4qj/KMhXdVhEGd0STZmewwiZkTDnhcLRZHfvvBhV5ZMyU45xs0I
rVgjP2zM/OWiQ/leE5mVRjcoTj7Sl7B85xGgNK76dK8Ou/77ey4E29FN6MqqbQJnL5S/XIHMaMLd
ZLgHDtB2DZdILU+8GRdnw7sqYFD0eGWLt5Xgo16v7OrRfprYF/HzVTMno/LsWE/bFZs7A7cXJZjp
Dh5b6seKNtLYST5sQWvbEVOwwcnFxc0YJI4S4kt3bldDKsSGwkw37PaHLuuuG+clNxGU8NwffVe8
wqGgH25BqP7z1bWm3KIRp0bLYzKo9vGh97BuybLFefwyax/jeGU8864KaluZjwOt7uhel/WwOKII
rqIQZh53aHxgD6T8KF0qbEQbKzgOjOv57H8Nf+HFd2c+abAA+t+bxlJltnwWMdeKbnysYlRHwBY9
muNCqRds6Yu+c8dWAyABfAq/04VBv1tEPe0jLSExQH/hevo5jMZkiesjfpkZwht8NJSZSQmzWdrw
thjRLc7pTqJAzGcwyK5i3nDKZEebSl/QS8ebnzxpYnoOpFYaq/b8k0bWZSoPulDK/sF4cWDE+jIN
jTo10fylPvVtS4zC4m4QAgIQ8W048JYfaymqMAkFJyqVLAP5obpKSh28jWzImCTMSRUASBLwaJLO
70w+DZHLls+T5iT4mEm0QFN6LwqRgLPEQGsd/F2q5NBGrbk5EbE0XJ9vhTLxTQzMvd7bVo+Se1Vd
bSuguijPJ9ud6w3m9V0cPlekGFMEXSruZ1O+vAg8ah5Tmqs7oyFMzrVZTx82HQQ+o2qobUPZNlKy
zmT9UPcFtH4nQgAUXCvFt1aU2iZjad+9ZD8otYQ172y39eB8zuw9YXR55usSdRxb35cnJfyUGbB6
b9JQS80CgRdwNh5Q+91bhQe9zmGVONrxlqp8EhfmksyggoA8HiwumPdZVueyfd8qx5F4n46FdWoC
JJ24dCTiFn1asJ+ge83rgiew5BRvzSy0ClKiLb1JtXfB+U1/KmT3Oa4tQl+RFTnws9rrHS9dJwLe
sbxJf5LNIjuIuJIoateeLoE5oBJoAo9K/2wuBY4cKAbo9Dh/QmwGtAfmi73gUoiOSERo7WM1c6AH
hVGtsl82BYPBDy8kWGJSvj5LMJl6Pmr7ieZJUTiweW2Nrp/1pDJuTQyh38AocGHqi2gtrvZBfLoj
eq+ndSYRFsv6c904AaV4p7vf07JfYsNuIdIJgqTDKV/cU+hLrpILmgOYF9eqiagHW0TaQCb7JYOz
uQhHMQE3f/ZoVDRE4irxhPmpA1M15OholZyeG+uSDo36lcJlfvZsoB0VZ+ydfOBJm8Mw9QXE6CuN
4T1BgUM8trX74pKf82HubvD/RH9LRlcc/qyNTTEK6+6Ju3Kbc69AFAhdBKAz5kCOoxy8Rv06lRAk
54m3LQiVKKzAClXN9uLs00g3Du16wvZu7DSEtHoZLlj1Sy7o4Cdf0D1cTp2kfpwfz48kVOOY6fcH
XKLovEkk6shyP9pNiYZ5u7izm0+hG3bxw1n3QUGHduumQw5fWFEcs/sONS6zDZy3qtctLXzqgL9h
XlTy0ypZdR/ZATF5rY/dWurhlzZbwpHUZNGFT8tDAKa+Ystp2Zw9fEF48fMkS0z10LD+4XduDeGN
sBPV0nD81oUbvXk6Z69eGu+vGc590zRRerdYu5XGuWyqVTO7so3TGB38RES1vVzq0yDVKcmmfZ7C
MVlfiIZ+m3QV4C6K3dc6aSTAShjf3z74P+ASLHDpYz1yrSLyBFexjfHvxqiKNh7/OMDvaMxl6x2r
70sZal55zVNStT8j71Bei7QSetTFXtZ8Fak8Mf84cgoGIfTEE9ryD6L/ZMesCsG5UF7Ser37A1sn
ep3Sw8Kko3iYjacOsryD0mjMybM50CDU4WXr0YvVr704JmJGhlHQrwkefYnAnugu23lF/XOnV6+P
iWjcsmMB6p11vgL2BfZman/EsAlmkeqlWR3tFNd+fx0lUVpOKFiqexrv9Tl0B2P8jLQs2XBeCkSw
8lgqpGm95fbPILi5YAdoRyBySvB6+V8bs/ekG8Q2YaX75z4K2qhMcQ6NsZWygx4Z4PdSyRbp6ojI
w7FcIPXKzDIdrKjStxdw/OUlRlN41ObbBiqqDkhhMnhz/RKh4ruJwbjqk6BPuvpUmA//sK4cLxvp
+w/XIvVE0TISZnIpPD3B3KnQXkyejaM0Nrl0gwgkoHK2vJbDcr7es/Wuooiv8UZRzeYYb8vR/VII
kyLbgNLOHwpbhsQdd9GXsaqPBrS96lJ6p+/P2iP27uAGw1eSZTD2o2FIBa2dimRnVWUyI8NhJUzm
wKydXsNyOmngnHwUFkKqTG8IJmSISMFsdmC+MIzSQJJ1hzCo1jvPvoUev1GSQojgHfE1UpPkvPL/
uFNSVl3BHEO/shSfP8P899L8vtMmPo062t/cUitveKG8prP8dxDjdG51uDU31nSeax/2vbI3nPTs
/Ka+rcyY+e0VjvJA5tsuAamlOVKUW3hVlkNMqCxyX4v1lOhioIoVpWHUoXGRDu9dJizIGFtGu4d1
c2EA8vQK2v1+ncsfFoti7s1F9jPd8ov2fKaZK6GpVlnIyAeHXPsYywQe3QOB4LNCZqs179gQ/TJS
DB5ksQjoNGNcK3n4ai5hvlCQiVF2w5s+cbE+KJhf+PqJnNWcjDZwDtX6/yOHhUIZXbDfO2AMaHug
WLPEnkUAOlS0k4WfmIoSShXpr4429FgaPcLSF0lhqwIQohelG+XZQmyVuWIEBdXenxahEpMxE+5R
WF5MDOquotPZyYEM1ULF7JKg2kziaZYB4eumslfBT+vg4G8PXwXhjORjtjz9XK5R/LPbOzRPegpv
sg8QrANawTbkq4yJXUzHza+rKzbdFDZEUYa2EesMjknMdcXgdM/zHbRSQwb82Bkp+uwc8DPsmF8f
GPoa6a7wMwJdjeWjbYQXKoC32EQSa4bfEhqK4Eu1vir7AgcRIk8Nx/87NhuxketnqYrEQ0pzJyw+
12VYlpouTB+bjcY7CaPRRJe1ikWanEZc3Nwby0DWJKh1TnvE0XW6WsBMcd7/C2KlLbBUoO50NIpJ
HfqPr6wvFN2k32ci+QhRAmchpz90w7xyvUSIJuYyPRyCANT9Cri8Rdt93XTOqPmiC8KltQJhIR5I
rQvW3WuIrinnm6yyZop4PjPFlUTlKXF3iG4idqWlmvZpCSON2gi/L8qCZhzMKb+1vRvHUYEiP0Ny
HnXvUDfKOzv9LD2lcYP/wI7mq4EroYj1frRd3ZWFOSGzZhLcOS0GlRcU9sBNuwlR8awZzigomAKX
O4s8gRPqSipQMb6lXK5UtdmqXXISj//U1qQllHqgUbADnc+OA+m6Wi7XqYfOwFYSR0Nb+loilOnp
8IzdbiFXNONlgn0UkOQf1TxbgDWD6ottACRIyMssx0OVQISEVGctAa8RqRrQJfyRrm+5bMODccUR
t28KA5/FRgTzl4U5RSyqQ2YgRjVA6cHSzVNh+bTob/IQm436UO7vJEdWbXe9NShSFxAcgQS1mrwK
+4+YGpbJN8YKhRDxoNnq5OEi0okYJK1jevnAhPJQAYL0oHRKwZn6C/0jHKvtmuCB6w+sZnAX8xMQ
GDQP6Jx2dKEt+3SqP3LR3+UvFIr1O7NEw+VYcZdTUYZi0UdbMLRVp39/56x+knQzt0uXgQYOZfER
Err+hkTgmPp81pSKv+nGpFQkHvv+TE7Kdx5ZT085t9jwl6ORBIezgA/y1zcvXG9NruwH4mtjyszs
8Ramfb8btPcIusmKW/e4Bl/3yCmYYS0u9+F3T8hpPbB4uI96InuK1VhUkjfsBt5pCR4zCK5tkuup
r+60AtqPGm6jp1tG/DygCShlvzWI6SkRsTuWFUVKIlBj3CoprJt8XrtvkGv7U2xs+Eu256kBOAiP
PbcLye94y/Fl0B35hQUWxkITN5qTY6rtbQwVz40OaMpl5rb6V4i+F2pC04LCv2zQwhfDPJD5MgK8
pIFb3hkzkGNkzxNLA4kwTChNJ2bZEfe1v7ZgU3pcdBRNdDIA+tetqKi/ZhostLg5OnoWpsuLvgt4
RNOfJT765/LyLbWogSu4mKPF+SZb1p656+bLPwtapI78r5jY4uUBJ7gUtlB2evoQ4LE+Kf6ECMZL
JHSPfB77O9pBVk/Y3FSalZMgJ2FnQub+OJForLHsxQHzYjPVJdVrHSBFSWSqkgwL4Mv7ug8JwTmC
Nf/zBPQZNJy5PJawhDUfmIjHBvgnMn9R3YqwskHM0Mr74X69f1wuh8Mh9g4Pa19jDMtP96et9nT8
3dCD2JwVr0Q3IEaL3/14Ugg7MDeoccnHdekm2PVXxhaJNhznRkycqAaTPWpOPZ07srINfsE08ftp
U4DvnIcLIpzXK8s8hK9LZWy8rKB0BtHVeJKDVeqy/4trpdwNdrx/wbxuA2Z5CDCjFyySjBARrm1z
4Cz0gVRHVuFLfX+flkahzeOrm4fA5y2L9iP62IeJ7ulJ+JK+FZhHhBDUzoLwvGfsRnCcX+gS4BPz
tmOFOpED9HO2oh3n3lcFEtXEnBXMBMjOxLpU0NWf4dIk9jsaiuIAG71jjTZOXI+agMOrJSWokFBP
CEGHGrEcTmFCc0hbOQKu6oUF55NsUDsAY4i/swP/3u4cVc2XnterQcNY2WqCSYAFzIZttaZ6S2Os
FUdpRZqO2+PhFPh1ZMa/c8BVCAf8V7lkbcG8qslMnQGJ6IruLwCR34UxyxpdhKgoljaGRshmhurp
K3ebyjnq1cXFItuVxG7iC7laNuwzkqvdw/RoRJI4CI2m+ojpG6vWl5PGDy/pNXptDty5f9LgolGX
Omb4mcskMwcWzEBdzo398gvXJu+BCkcY4tKb3u2iRfYxmR4SN4P5G9Jxw1os2tG4mXB2EGQHgvC8
/RYtuFuWzLIG/I9Ul9mI2GE4bH8w+BagkCdtUUzqhhjiAcMHc8fd9DPUwnUzZIiA61Dw2o8iXevs
agUktWn9jQDsGcc6bcIxoyls4BKdw1b1nQW8nte37+oSmTki0FU5iS9H0mzkUx5UZ/K1GHg8hFRw
l+xrjII446yFXhTSSkHMExMXh0+IwkllpOSIVXfmuGWrl01jijl4bO5mK8en0vgJ8P4VYUrn8l6+
8E82PATyOYd+VamWltsy5VPNy7shOPzET5VPPLwAoEf/y5tVQujb4vy5Ak1IgK0SDJRkA0a++7T4
JmwaW/LFC8WjIr+T/XUovLeH4Kj5+20gxxkvAO9vks9ni8ONJv/pxqFCBi42o3KJWLWL4a/pyhjo
4qrJQliZQ71PBySL/22c9mbKiNned4GFsGbL0xh9RVWd/mCvRwy5rdqD+cQWulY2k0BkqinaOjOk
pOhAAIcclCFx3N8UeseT/jXQi9VuMXxys2MHVsAOiYrejz3Zr44VM402drZdhHzxa8PgsRJTL+lV
0q20DmLseiiukcAnLXn3IqrZJWfkakZN/7CaCM9GQAPVkSeeSqvscK+rWTNlli4U0daKYjI4UJCx
JAbQGkeaFMjMM+t0Z6syxzY5Cd95Uo2x0r6jReqg09xmgHm48TKt12324SqsFktESq5TD1VQILa4
ueOxiFGBSgSWRxBb5yS7j5SI3NZhqO2PLfUsfyEpO2kJGl3SA4dUcWn0i7PizcLpczVvPz5NV48t
Ol6wWbvBcpIJ98PxN4aZkbPJkDAV3FlEnl20UQsGirb9dH5kCgbe9CV+UjhvmH9DEnoXlHUHYRHY
AzSkUTVOoYDdOi3dwQpT+gQl/C+b+7tFiYOW/fYtBvBFhBJ0IhZcPkSI2CtczYct50PO/3KNSMPX
2JE2LUfKFvmSvVXQaghONpPugj134Glm+XX2z2reUGdT8EgMZxga8UlBkoP4so9eSYrrsfeGYxz+
SkGRbaNxPw4Dbw4ldz6eZAQFCtUnkgU+yljFSc7J2Z7Y2KrEKLktLj6wAu1H0VmG9up/fm6BFyLL
q4lMs9ZLQvX4lS66dISvlz9kNVaaC1UmxRNHezqDegB0DqTMg+XJlL2nmCIlI//IcpaJdbEHLdGC
HVCBrpafIo0hljbsdpP/kGzUvAB5Ne093SsRkPQATG/Inq8XvyerCnjSxUzV3DwMALV6imfUwwh8
RwhLmx5ES9OhM405UMfIh7NHONlOstFA/VMNPIJpc/FemM8ZpQbfWzXH0Lg/P+C5ZUQKjO9xt0Xt
hpCqi175ajRRcbFNV0L83cUYKv4BeCy0XEbXOGp9P/0GHfKoxIQvGpKa2189WlB6DkS/Cv4P/DgX
GNDz/ci5NczEvbb/SqMobJFUsplrnqSffBuVthWL7EwL0LKc/lK+sRbc6uubkxaLzBKfiyseMRG0
221u8nU8llApWwQtPgfP5AUde2P3RLG/VPXnc6IhHjGIrb6m7HaIASmCsYUDQROO/2MDePk0ZgWY
ONRmlOWrIrqx+Sq7imdyYg/tdoHrrJHm2+kGH0HNw3L8Utu9DDdX4eIh2uVLDAl8LRjMl67v/oUV
BaPJN4p9bwGMwtKx7HcCyv/H0rdBEvwSJVhB8s06UnaOV/L87IFPcXc0N0/eeswtSQNbvMgYgchW
lJi1BV/eBMgVbt/BC/7ZSP3w59Ow8qE9KBUMgHbDZjwLpN8hJxZi2jf1qRoJOrOF9S9kmfYDAHoQ
xFFoktos9itBebuZbv98wAEKCUbCCkJyT6QjTZm1o/AMnr6HSUjNEJTKFTMY89/4DJw9n30HLRU2
L8UH+XlX6t1epC9FqhSD5ylJLO93yEFYPukd+h8XRpwGtWqs+EXs6Vq/PnNcvGd/uTd86qZfFU4O
HNKCaIYfU5CZXt1ORP8jiHPu5SV/XXfhLwP0o/pbyN0eo2I5w1EMxBLTKt5MR300HXLuwyqd8f6m
2oGa0e6EouHcoH0NCxdOrBKKmBbbbf4IawryGd6ezTTknbxLg4F/FWx6mIq8iMl+KEtDDyyJFv01
q3IhCps9Wxc4kjr+EwHpBlVmRQCfTdeSN2LzQ/53LrgjXfQatF/0q/MU6zt3nhiWEXBAM8dBkB7P
wAQTV4FsInsuQL05LZlfsRVy6ZJmQUwIqjm60tBDJmjiKDMG5PxAQEf/ZB2xEffSfRmcjjEfGn6o
/JWYDW7l5CegNOBCx8Hazo4MN5cJZqej0CukZmYfR1zBLWLtd2gRqVhu/SjPVSwgJI8aPpa5lErZ
kDIvi4ag3eBbw/2qv9qwHzKBnOwEpussrEWps+sfh4nekeDcbBxkr8AgKq/cAQXTzT+Hj5wgbXVU
UDwQ8ZIPNSDc/TJqfmvyjgYpTDc4kHc+fWSJPanxcbD4tSeRIMO4iv3NQQ3kApvkv+vl4F5hQgr7
C1to+Wmt5KBnpLVBsAqVtsmmra5PfPoL5yMKljdsk/cTxYTf1rvxZwVIXPoVoBqlOSDvNVQbmpP4
i6k7Ki4mt3YllrrkI/hQWZaPUVvbeceUn5J2hBg2kzNg+5MfV4gTut0Bti3HCpHZTU3h9t/ZgOrI
UjCqxOdbrRbHZ7OyGNoWh8v+vv4vfwVPPQxVV8vnZ+IWKnDIgqXybeNlNTKB1iITqPhCq4w95+yG
+SUhXUlY4HYqqUaKnkw/ciymlMV++MVORYTyaUPWV8ovEH8/buiFnpERQv3w/rA0Cy1907+col7T
NQ6TCLkk8EcjsYJXJZrZhWi4N1icM9ttCzNXStgOS4txE3R4X1IILfmZO6DibCill162PjwVUvmP
WX3uStZcedBZ8cju1Y3Hn0UYN4mcN9/OY7QyIzD/vLI2mFLie5K0Tr4QFcEIX7LoGAo2Pf/jUoUs
CJ6X+iKnc/4MiGCIuT0oZefljWaEAQb3aWaVH2hscIIDVPjxz8ILKryMdIWKwnQRMse7uQ/i1fzD
ligU3MCDTDH8JuT421n40k/XoJFmeLzN0Q6G0VRYRfdzqlxYJrXWGR5Z31eSx9j9I1KbqxAdZI2g
wDSeAZ42Z576yTlvbYAKsLusqDVgw7tHCEBKzbckzaYltSeE3+/ohhFLCNGYFJNy0AKkQyWQJ5q3
vsT8ldeux8i7V6wPOhKzp98CBQILxRKTsybQfX9fBF07aX0mPdvWxtxyr9wGXiUJ0m/YbW+X+yRz
JLmeK/HDgBa7rf3O1Es3fvhpd64ojWccK9K6AUnWRF/JBJiw7uJizkozZqatlbouPbD1BjbWIkz5
WARWBrS/Ee+8pKc4xkicL8A9c0tmArAwL2FrXFV+tJusniQmbSxlyGKo0eetF6hh4+bvRv2K6kC7
af4dI+N6k5b7uu4GX99LeNdRxwZUCgK5M4jrIXkcUuu/tAFwc6FN/PDuJ0xDFzUGVOrCksUubm9T
dFVfMOOY90cnQdxDBDKR0HMKB+WgiPty4T74D4109hAdd1lrto7PGJLpeqM+bLsBKD/rEODijTbA
afnD6VRV6PPc8XE/ByCHd4juhjnjeqRHocqDfw61WuBbHyMAJ/pFAshzro+RdKaEtHekTqYusVQR
CTpTOkFi0BRjWI3olFYxvaEM8SYwaiExtIiXlJqT3jQ8xVXZdl9N7qPGi5+43dGlaJRt9X9UMh8D
n2N+Iik8oGDnXuujTcPeFGK2/TY9AiuIEe8Ji9kovPcQrYVaAjXmkwSXFffX0qC7V+deXGaFugwk
jV7p+YkmDPolKyF4+h9YWUcTLAxpGIssj+UdFq6yRlEmOSoGVjxfgzZc5jahOpnq1bvAO2VMxzzd
LHB58G9ATicR+pYfJLTjeRw+DLwerFu6zHQ8/vh8jekVGBxyfs8fd6ZSBPhUDgzlwZ7rqxLBj5GK
yHVSFEC6KEY3dZeu34LO2miIKH+pP4k6uw9YY8mWO5Um/8V498NXgkCYp1iBtg2z1GmT8qLDZZLm
uRLFX0TbFhFDb/BQaUW22OyheXn33vRXQRC6q/6lXxjYnJCblp14NwHaspeNJUEReD8PCYjykA1L
0pWdLJTJ+pWRQHWh0F4rXhKX7oKz/LRBx/9AACFiKuEJJsdfm0RCY8u7vcUBp5my52ysFaq2BB88
dozBeOwU9oLXpa7pZ/qlWPz+i65mleCT3udrNbih3t0B7dbQTLQQOcRehCRloQQiC2AmQmaGCHnh
S0rwJzgiaE2HwXYZB21UzpA8iq+weABbadBA2d9FLI/nB3MntGJRJ+nGJ0vQ/3BgCtPKp3c59xX4
NI0xb3xqqQ7yxRsIVsjw9IMwhYAwEjB2ahsISgK+mMl1e63MUATEPi8QMwnaJjwszlvQj5uVX588
kktMjjP8RwTZ5KG8g0okKfsDZ06McJZAmcHPdKKq4m4FUfmBCf6Nv7IoqEhBrpnNufks3ELe4Qho
efiC6ZHrWaZ4oXv4A+M7IvehX7179XyOX6xkQLJEK/bo9+hzGREP+rGqLwW205dGim7kcJ1f3Ix/
gf27r1tSzWNO+i/TLpeALSi75YC6FX+auO55fa3o3eBKSssqTahmvVYEAli+zpJ2gZT53HpCDZOk
1233CRnCqjWC1zRQ04ACpE1FKfTiTIj2ibEpEeJpF8lgfiYkQV3BxNr9GFaxdQlsK0Yh327g9VK0
FoCChqWg/vmKAY/ZXKxgS6fug5b9XEluEievypeVrnihJ4kBlTj+xUrbVJEBHljkSyquaaEpRFwX
0zgpNy5Na6M6bSCbl6wcb2by2svEZooApBhBAIrcDRmIa9MHIAs/uYTpikpECQSxtmTl33RezgyR
VBoBDarLDe7OeXmYLP3S8mY3TMebWrHlDGNpkdnqLOtayItvElrL4j5yqi/sc/uUiw1gpyH9qdjx
Fgq9TiMpIxxdyHwR/WeCXjKtEAEb1md9uA6xQIddTqmAeFflTmbB7EdLY99LFLDlEnHP0JN/Tv4a
GHPTzQE9vbNusyXXjok7xxpjQ1x3kieQ/6wQBIyhaw2rHJhyDm2+7t4XMuPCt9FFlWDKb//jr5JH
t4s+LB8zGXaVaMD678RFscQ5o9o5VwoYxmHomyjUMxaq5Au501V742aXAO8iGkTG/AW1a/P2LguI
biMG72A5/BBV4x5lS6H68V5c8ZuDUQf5I3JtXk2BobjPYVIf61waBRcH0yffGx03RyvHdFpK7XLC
IkQmN2yOR03O8AqV+SMFEL9NhvBmixPlPeY8v7Pq7KguVSj/esTW6WxcDhYX938RS14dmK8QroLs
6zPfpZqV/A/VIF+6tL9AggdcBRhDeW+rzo1C0FomnQniPyy7itTDAhtanO1AvpByz32aO1kUJi8A
Xv5FdoViiXCbkJRuRuV90/NvCFgXNGSQmUaEyQ9S3kOHxjnC9mLYDbuYo3TsPWo2+JCBsOuGsoOC
AEK24cj9IiGA1hMP7ESgWx8tKbEu56yxmNBBueLgEV3IpNPL2cD5b8G2NaKqkXpAlC+fOZ6CTxjI
MDsQse/LLTnbe63svDp+VYJOl0DPulQAIYK7hD1tkPK0oOCdzzbbqFHQBBX0pNY8HAt1o+GLNdgt
tEsqRUfWXpy1yPxAPEcUse3h5iaOy4OJOvAqITnCIN63/DKNwg9h13hdXh+tTajneyeQMi5SHwiq
bLENfomBW2EdFVdczVqGrqhch8jhw12hfugZadP8Iiqb/LbxB7O4S7kV+1wqRF81xAyMQpBq22GB
4VTNuXJ4B1cCND00kfxGEuAWNNwG3rNlixni5cMw1F5VOrAbFl9eO6rPzaeDUlKXKUG0EYlwjBKx
i2wYDsWItdFX0rMlnrHmAG103bQiKS9DgFrq6dGb/Lv+Ijqxiyg6p7Pi8E7tGfR5Zw7VP4IfJdP0
DW4k6oIai9HqZiHKFmBKFmaeAreocBRz0a8DKI/xdRfCk99kexc8ejUXRPO5L5tJSFAsKEUB9f2c
146TWatq3Mie5PVnuUEP/CpMqHJG7hRxU6ghka++EjHENE4tVMINdP1S9aAdFzgnTy9dEygJowVF
Yo4N+vHPA117/zyaDOHooM1uaotGHFhdzxEN/RUue+pYhnvlCvDOfmf/vOzNhEGg2US2WWbGOgmC
OxipIqho1VkmoTy/D5+PEKuyxVF284Tqvg/gL2LDbEuGHObHPHmoINMQMfFeEh/qJYdbCAU8lQyk
uqQiQ30ZwSdZyhLuQkUkndiOOb1G5QQGCUZleaWgVCdwtjj8ehNgoID9ZlWwG47OGQgrTbH5RYpy
oL4+wcJKL5Mxy/DgxSvWgeIv5M5i2GVRv1u7EviXfHLFS6ccuiuWr5PGO+4xzjTc+VcvXe2Umo9h
deaGsa/WZ+XUkAMji+o3B1oH2gri7lF2h1BYsdhiWmxWHl0UMXqUg4miP8Dhm3eEwQU/y/AIaU5B
VefBfhMwPU2X8BWSGK+7A7cm6syodqO60MJU5Xh8rhwsROVl+9mYH/NE3oqWZFbUbJTzeXzwUAmn
2mqGNBsUkd+8eSxagKFdq+m13AdBjzs6lpVfe3MuRxSy4a6BkpxAhDU8NbYsOdbawSlMJV2aiAkr
hhxgPYbOo3zJ9k/4C9IzWAMKu3y1fSnneOToJ85bFGCmumBbCM2ppJyL+30ax5MU1WPtnkHDwJ2u
yF5pgodCBbeFLplSTc+rK2+opHOginGlFB4Fg1kcSkPbhAGG0ofZpQy48NUEJboBrLUqRX9g3LxZ
jbvtyK9t0G+hqlMfP+pqQIJ1T7c4UK7yezWPUmE8QPWtqt2Off4vBinCNVWTec3ZLbkWI0pAOKlm
rBq5bF7ocifsOZ+SIhRt4Y/msl9JHGbkxUAx1SkEGPoYEGGSLrHGWhfiMLzFrkhyRJz0E0RxU/1q
FBTa1pgrRTukrRad9qqWHyUu8lQjjZ9XktLsWIKJliNDap+yCbwQ0mlnI/FIVaQmwyM8TCxnL/5c
Z0a+AWD1aVT3EfzSFKAB05H5GMgh+kcUnCB7KeB6aOiZfp6ODG9NHjGJN1XvKBkvp5DiyPlE2Abr
Q3uRnb0nUqEPGq/fxNV/Y2ajfPF4jLEoyE4qxwdeSFyYSXF0SqWH6AL53BoGaUmLMary7ubm15oU
gaSSpyaZJE6oZVT8+UgiuQGaFSZn53/mt2hXmTuZ+fg9D8SLOw/cSdb0JL5AQolAuFvlIe+Aodwk
nbm7YbJ/Px8XuUfrGkMN4cDpwlVCVAbVFcYO4jEbqq95hDasDuwGzbvImXJEBfkvSR0geNtH0nyi
q8TFuId14Hzg7kyurLyjzr3p1iODs9P4fvplxrgPxFcT5kUsNioJhAb5pgRMOAiqpVkLIEa/nmT3
D6XXhGONKiALuFW4w+OjPTq0L5ao8PPxCl6mkJrMavSkc71m3P4EMJymI5b9z9oYovW69bBdyQZU
sglhaxK/bgNp+JzQ78AUsa7WM0rtyR8O6QmrEJYvcSOWfips4ZzQHiVUQwrPar0+FGhfCCZC1e8e
lO+ryb1tyhQabYFemPTOMcPWn2c1A6fzgqernU0fYpziVtOHfKy1V9eC3oXE7CyFNOO69siTL8mE
/3bm4Ns94+qRMjxo6QeHVv4XGKaLzSu7pv/dFhUKsyi+EPllWWpu8B+YS+MmW7Atmlp3hIFLQ9lG
5c/8xa8CbOb17+CLVGKDIl6elKl5fuy5wdM24X8RZPVxW4HOsk5aN/XA7jA+0QUrqxcupFqoZdIY
axZKJzs8Bx5eZZFv0vnRSrMQTdqllDE1eowEDJiydVoNd0JW+3pRk7Hl7Hnny33tHGaV0osOtlE5
8p8jZNt2Azao3NAm+9skxEZvNAmaFjbP1gtJCUsmsVI9Uv5eD3S8XJwGdqtXNakhyq2NukYaeXq+
HxAMD2G61MvNT1CCIC7pKddMK8YQL5KTH7K6liae5Flb+afpw1L3L9tzCp7+jxAAZVtnN912B9xB
UhwVl11yOiW2cCduCdS1xJJakxSw+pA+B2WNjpeeljwBIES2nPuY1PSoyJlL9ZocbvhxWFz0a2fL
2qb2MqzmP2PN4oDOTuCMud4v2ndWgcqUWEWDgbYRVNwhMJ2Bl3JIax7CmkSmEnCWOqOAV5gVNoNn
YxYfJSziuBZCh/7TjK0TIyhYf3ne8p9W1nhwsMoEwapy+z5IPNw60YQRZ1doNnCOIsR87m57o5Ec
TAQerVyo/0J1BsUfx2QS8vGhNJ/n25zNLT9rS0iHqlklG0b1IkLRjrvZaiSneeP9dUcEalEcY4OC
jhn+2ojGg5IerI+DKhJiPLTBemjbNlESRSl1nl38Y9EM3np6Wv/W4F4MWfzvTTKDbIarSJqN2Ux5
pUsh9y+ciXpCiwk/juV/XW91ryhfYf/oqHn6Vjk7mAWeHiEWrSRVMSBwyjDyKTMWLuOjY1GLDKOj
5ewiWT78al4XSq+ZH0jra4C1e+JhCNNgB0CWMNWLBuYAMhHqeS5lJKbPUn0+itHdvzvXq/wQqE4w
z4D8UsSRK+6bNIIPrLXzNlstz5DzkPxVKrxRfRY+nOVEWQjczLyiBKD9qto6SKjPLTeHlKhL/oe1
1IEorhSi4W9aVa0o1ad7NFPXrRZLF+BkwM8frd15euOBeHL0DdO3eXtwxvoAJzmZj3v1K6XsgAVx
1wCE2BAE/4W3AdOfUMpE1S1s4dBXHDcoYgn49BINITSCeITd0g3eH7gWNbxu23OiJpijJffLu5Sz
kcZ+/pMscRlTLIbGeDyBGpS042sEOTwsfAtbMobGnrWlYoXRO4bXvqHh1jfCgfN4ihxkPFOBFtIw
Kdxzrum3tF6DmMJheZIy1qr6v0UoioE/HRmGF/mkkRry5+4vwHhduCDI3EQpu0nJRAFkgFgBuJ76
3vQz5DE2HCn4fQEscH3P5Bs9Mr6ORBqVxffnE3sH2tzRo1pMu7IR7h345P906+1g9ug/jHF2I/ID
K2HqZczYk/eyiln4e0m/noP/1UR7hLnk4nB8mXSm3mJdTHPsQJ1NJw6YHzDCeXihszo+wrAGJ033
/jgtwvcOMqk0GyLzAYfvW9qUHBlEjjicn28ON0SBjNHT+BYYfCeqIEvguGVExW5sk7R2k9caS+xW
1QoDGDZmQPt+qM/Z+TRMewNcqkiyBhrqLsUq5eiMhfotG3mvjAUh0JeFL6Q7Q3fj+bABkoyT+4Lq
MPhdvDt0nhpgGHocvI3jPlhkkdgQSfXeBTwcBaRsI149PCj3c04O9dvDj9x2D5TCZGHzvc8ZowrM
Wu1cE0qmVr5fbpaRmQeweQp9+1d2mnOaxB7h92VJByTJL4SaYAaI4WCkZNNp1jqpJGQPRN85YXlj
x65r8c9Y/+R/Lch63Hb0KC0pcWFosRjvrxEg5gVpsTNkd62QYj4K8ze2MWS2jb4qTUzauD1JsrBE
kWWHJhjM40WqPt6QQ0AfbMJPk/kmT4mN5kDrvgMnbrRZv3l+obyGuKNkMUjI3f7bSo1UDoVviI6S
aR4BnUE0mJt5sy5Ogb6gYOyI535nQp+S1uMdxSr62zjoFxcF/S6/W2iNSTSu1j3qAtgdmZ5kHGhp
mWrRaH4k7L3s2+bk5XDl2QkeRV2Is8KaOX8LG9B9/kAVotY5AvUG9Cy48iI1lPOjrxa6MceQ64wV
IzI/epk3zEN/ML+VBoTPMuSwLb0NiB9LbOO8dF48WgKOLUJOHuwMAmaP9VfEeVWMP3yzkIRI5ses
wP9XdsI6nJY6XTbWM6Jpa++Oheh/QLRhi+45VBZ+LqRtV+S1Jg8J/v5gDRWaFWM4twGqO83YhOFk
F4olpdDxe3ePbmuPwqPsSenki1hELL20JDY0XrJhcmaIY8yvetZa/T7uhIywhCbpO9xEGkEqVTDK
fjRSKoFgJzj/03OtPxKjQDb43PJF+K1jv5Th/6YqTpF5n8lWlVGKwosTeRWZ9oauWr9sc3c72jme
poZ3A7neB1YOUWeajhbnuwUt9zNeXl9WFXEu0IocSycakDnKIthY4K7qO9FColehGjma4uo/0boq
GNtByUzsWuS9sRB3qYzDh2FiTT6itPGi/yqWLsKY0CqtRKiZCmvlHDlOx7GhOtp1ao3guK0cQGo/
29WGSMtOAPVVNaR5y2pzeRcWdcabG8ikoHXhQ4CWDtURCRjGmqHwsSA6+vfFBSQF6kN8+PRsHu0z
Zm4pQk8Wd3lskBQ2OsNYEA2CzENkb/vq01Q2RnXJMqt3KMaZ6V5avJr9DDbkiolyLMVBSEkfTyTC
M63jvZxVejCUR0XARqUmS209gNTUtt5QxXRDAEiNm6mUNC5808rKSBJLzh+oMtNRC87Gm6IRLfiD
YcLV9HZ27d9mYVkvex7D3qG3oOxuYdOOioBH6/WbKzOEbPnt3F1RYHQ2OM7vDybeqGC2SsrakBTA
acck61PEcILAr+yQ/x8/Ph6VJs15M2JsX64eEQQ/IhZp013Mvjq+2/DWlQhxqLywosIE74GwhG/9
WyLwGT/Md9d55FAM0xHgDUUrKg5potifEVlQRtCKbrjcgza1kS0OwxZF7TEtc5lBVO0yLTUBNMo2
DvCCjWzaxINHVwecrHC7qS8pGkAmdO8xLmW8kny2YkTHft1kPZnGyphMbNIHtVBOHFxJrVlSipcq
pzs71DednN5qPE78g57I24k9czXKvthF+Efs+yyecymJWz9EQJ9ny0mV1DiBaIBrPPouHxj8sBhO
BA0UF0/uhO8DUGwo85Lb2mWZHN62A+YuK1DGvf/5zSZgLOWoWfjRnrl54Obdqrg43wBJ59HJ3E3L
kWCpx1dENNYdfpSVK+EUr/AZNU1tlp00W6luRzSeAVVbX8EmyKyzs2KzHYsTjL5vXsdUJtpJV73/
v82whzPdtq0RenBQy2I4lY6CKp3hXl0wsyk86Jc63bqwm2jt2rq1RdB+LMN6YOG5TRr9GPW5Sin3
bZrzlmRrCLLlYsY2m1jHOMbMpe34q5rgqhKmQYqTUl5iHCpg7MH+hHd/cWLXlwpI0N9+QmkygBP9
C+uCJcz/hfl9t1Vaq0uGyRKoh3IHmHzargXGh317YRmjcqRjlAVXMU+RRqrXCRY5j70R6cilDOUR
mftLg3p5XIyqP6MT5j/A7/6xylfbTgVOcBmgOp+hUf98tJdGjZEP5LYNRSE+OURPuEY+zQ5aYI2x
NnCpSyjLvr4lZCr7+07cVixZ1l2oW3IqkH6P/c2MTQg+CItJtgNfI4KBL80y6jUd4/yYG1an9Dgv
d3RI2Y74GahwCq3cRE5IdaWoVgeCGQduXyUhYfy/WHPxuaEGlNgedhWo52UDVy8Dm1ZpH4Kx3pPx
ta7jPmo53EfoHhnDrK5XAFz4zPQH30jaQ1RIDBpT45YA4fD1JZyYvcZIV87xICxC0D7ugpa8yevW
RgSOLXRUiXyXt7gebYvWXvvxQ220D5C9VwOru0Q/wWpzavhwYlgiate95jZ/AAtWVeYWUhZJP/Xh
ALx/M4og04LmBYFTo9UJ0mXYMWHKrDCCBBgDazQUmawxTgdzqYI28jOn4+5Df7/qx0AouTkURIDA
RIHePd6DsReCG+x6WWI4HvyeVngrLAPYVwykZB/lP+h1fS7IFHmbg5xmpFnELWSRxzxOcZecHvA7
PB6YHxtqvhy/9wqlR4UySYqjEVoAQxfRNgXATyO2VA0LWtDobt0DORxbz97R8aNx2Rqtun2enmty
w74Jb6YYxuxqI9URyqRek76vZJhvY7kckun4rbK0F6E/WJSbqh41GuF3eeo4pCLdLF1RuD2p0yQ2
hfucwgQWfQ+RGkYPWo7Ncvvityb9lUD4If7ohbYG+6z+qhG16A6O2IxKv8TNIN0cTXmH27fbwe5M
qQQ3zChmA2nImsfqx5E+RHX6hunj/JwGJoRvoyGVlvrNWGQPOVlHSPQDR3Oog1lSyNe580/dS5ff
By5Loui/E5gCpZtKuJ6NFwnLH/mNpav5sCBtV7JvPsA7sg7fjceXGWz/F3BpIPOZD1FulZTfpMRA
fsE32aUoXRpALdtAfLTcY2rPSEc/16pSlC5lvwBDSEGYipZJLxtTNxPzcHOxPVv61SR1h2xqYI0Q
UgrWs90bXNBFmZmwUX40iueRamTFG8bLcqw9tgV/HLU1CrkcM69QJVPpKoXWzl2xmIImf61gygKC
Dw54d5W+n7gq+ed7u1RRdn507h5LHxEz4VXJRq5EKotcQKo9192uzDJdK8lXyOBEFUhWxaPMKhC2
AZjvexGRXcTidmU5b43eM+7EjzSGwFYrnn65Oh7j5lkboUkudrdVYSGLP5tMyZnP9MGcrvmQsQo0
2z0IPjalvZhWfQx6RfW+SE6wkNWgSav4TZBudzi+5HeZo9FDYh9DWGHJdj3ZYTPwYVS2NIFqr+M7
plaKy/pFT8pNfn+mNmCTom7I4YNh13mCfWRkcxwCkVM3Y5dUhPrYjxYUtfg11r9rToEXS39lQrfq
8h9niNsaMkYbMya0Gl9BpGpSmgSGzzHD1iCc+Y/0i4FaJoGZew6SdCsrP9I+vHxWc9wgbu5NVSbP
o+2hwvyGsPDV1Nt1rh8ueOOIk1xwbORSDrKl2qcBJmGIHBpZ12vrOALt/lyC7kOMM7eqRY4/i4hH
j/X/R58i5/m0cSNRcmyxuDiwudDhwj8mPqzgu1vfafDPgyQCjNZsOMO8ejmCwfm+HepE41tR9Rt4
aaEDy/yhDiYnRI37c9Kt7GQZoTw/WGPshOwUqMUr2tpdNefB2fOaTxG/AftV5FZ5xwuQUBRCnwG0
RWNSlgUYep/RuQCjVLDXlJkZoxj7Z8a/RddVR/DhcFaMHhK5173HXz55U2e/I0F5tFDhEgC9tUMr
39ziqOBKw69ynTkxe0jdizVkNow3rO8AZZRZEvfDbXXAmGFJ52v3M0EzQc6Hk3iZMbOBbuT0SGi8
fezIsnhlN4/Sh9TR05OsL695pMmT1FSTCxXe86Jx7xTEqsWKHFcO7LyizPKQhiym4kgkoF7023f2
DaVjZUwJWIO4bJyrVEmpHjj7g/2f+oCW5tq/biHQcHe13y9v2PTUoL0Ju8bnfKrGwyo4tUy/jjJp
p/G3sNe1IBeSkl9T0QkePGWboxijOQJ9JCtcnpw6QS4GSseHx8/pJXO2SDhMBs05cHUN+RiMqeeO
QxY0wKBEGCOLbECK1kiSq6DwAuaaPL1Pl4Oo3Oii18gQwhQbKO85cnWCdf2IDLeshhRwygh7I6zX
I0bLl/hq1X/+U61mZBACNszh/mVc1ZdRSjdPMAgC3nvb0SfbeUtafC9uOmwFxbOgJBXs74AlGHkX
kKZuSna+0miCWpwjFziAw/E984G85utEg1BZlSar0vVdGZFXDDbBD3Yb1lsSNSBtqOYhyAN71MfD
jQaUXqbEN6d/GdFiboAb5nXy2dIePk9k326jQNRuHXXAqmZmJmPQhjq7C5XGM1kEpzxU2EuLR4ha
h2nWxwEpemDnmdsull3honhqwQ+oOp92wI99iWILPvbhSldJYWvAsnuu3hIVZ75RZCz5UrG5Amz7
JtssKQ+HrSOiBRvuU+VY2eGrjywg6zyVlU7IBt42md8EPmFudnau4+8Nm1AqgzkVIjI7oe67eOxm
CLzTkRlQsA6kFHTRTYLG2TI0cnC4n6p0Crb1AndePJexZa0Y/EfDuhx/IT6EORRY3743DFZQoWj+
9EHM+zRqZaQC+UF5YgG4cKnJ3eL1DhhswbzS9Wf7U1mxxWEkDo8EZDqeezFSU+tit29MOjz2sDaM
JOxaDb7W/KEem1zdS7UvZJ2238M1bFK3WEo0Eb2ojY4qKq5uffPi6GXmNnaPS27Revb79H3TDITn
8WgDr0d0WfrM6mPJJzOC49tjPVFVxeLl+jGnSo+C8xs9HfZIgTPVv04T4+QuvpngyPJqN8Ucm+7R
gMvRYVXAmTGjzl/OUx7IgmeAfZxHI2OFMaHzp+3KnHfLj73+PAVyNH7YQlBp/JyialaG0sTLa5V+
JB4R+2SWRrbCeEXVqiDMzyDkvFNGiaode72F+bcRvWeNhFDW8Np7GtgHakUMLWnTKSSsue+G+bTU
jnKZkfgBL1Oohm8rFUT3db1v8k9b02rJeGlGMVfx0ndDTa7Axv4ScqX9MpP+AqhbFtKQCAJz+crj
IPG6uBLK1HrwuvQU4tueYh5JTaI2IHwT2mRk15xt7Mis1qfJYsGZIRCziE9B3o5KTHwum4HFEJCI
E+3FJgpvyh4cQD//Lje+6hkXmYRbS9IKZCjFvrXFoBtZYkVwsZ0BCHQ3B7qxZ7WxLvwRBYiVCrWS
eRh+K1GDPnuDvO/YukRL0dpEIs5OcYM5yIuhO0U8fxkHFA1vvFlRuH8W9cR978pfaFAAcrx6chXe
LINqiJ5XmzrHMuMt+6R5ELiMljAghy8hA6S2pjp8X1/7S8GkVzQe0BK/StStXX73bZKh1rp+qohV
YJFZN5HJfjFz630cId2Y4HNJJQKzNNT/61DP1Z1fQ/fwVYNtulAxTZh/LD22oKe7jHK0d327co6Y
xzfN2YgPyZ5V+NPP5Y2UmaPoy+fL7V78tYqHrMFfOlGKZEyHNdZDuj/YtShmRZeIwPChjEJy3DQU
iNLIsp6hlOlgJajYGJ3jY0Ey1Doxk/MBkKD0ZmeRpAdcefxsGNB/XhELSYoTDW5rgg5u3uHdncMU
FnKLkaseSCgHpEziGMxYaJ6zswpngnzVoDo6MnSvSAAye6cmPoGmZtua/J0b87mzDxfTwLpdHTWC
LTfbyLOP/xEI3fwDdgkkS9mAxUs+AyeddKfeKVoyMhEb3yW7i3nco1LhKICZmEGKiMK5lkZtIPJo
QAgxUITNUMuFc4+wGXQkIcoVOUV/v8OQjrWhslj/vaCK2Z4O+1AmYJ7/J4Qn9zleOLhAInPsL6eI
eFaw0Ec8gNeosBQrGuh/xC/p7erYmFaQRQQfSsARlnTtljo72/rSPHdmM2rDvxOVR9jo/WnUHWmh
yA4B156sHKtjko6LOiX6YoT+tGRDfpD6wns9Ct5oX8QZMofgVuhMwC1r5PKZDJMO30QiX3pCqA9u
owMq0UgmTOXWAghJuHW2XSBBSq1X4iWm1klQyPmcFyq1OO4LcdFZmY6HO6OWiPgmwJv91M9Hcc9A
8IEDxwsI1iyqdfRMM4KZOGgviaO0P/E5glEH1J7fapV/sjoXVbDWHhVY5ypNL1BEyLwNvI/n26pC
7fciTHNC8ZlyqF7kO4fD2/TqOwWZG9rDctWQLiwnHIgW028sQsHHUaAr6mfENzsZDwRol/oVP9T0
HjKwESTKO/LBiTrntzRUcTJJJs+3kbCl6kxnSqUBp9AVcpuSQBd2LZHX56OgBYtu0slNNuDbKZHC
taVXFRc/U0tYY+8igFGSMA6g/347KNqG/glVpnEbcJO9/zJs204tpAEJZlriio6iFqa5z/ygTcKN
JELJU1U4WLIs8AodHGvGjN2FFtXrYFsQhIYQYaC5GrCcdoAGj9FKY06cGIqcapG1DqmFisrmy0gl
bqfXISY65RPU/whppSqKXw/Bm949CeSMM4lJeJrEKhOsS2v9LWBCbFHSRoYErhzHfPtVgZySAkBn
OgsiB8stuNyKNNEryXEtIYrrv8/tVKieJWiIHLOEOLsDxCgcQIpObh8DnaPqxe/wmdCl8pDO0lg1
I8B78n9DnWAfZZ0ynIB8nlhwpXEf5c4Y40HiBGXM6qWK1ACMWDw4K4v5LqAjLsp8I48G8hTw+Yhs
Ub6fIMsQcwEUvHr32bx92u7SqmGv9dVAW4kR5+xK7SxyIdcVdeHsTVrIxo1u2LMtQgI1Rg5TdZpq
xwSEonqV/M8l/UKP0WARZoNqx5fXbEDdvjABdy3XD7pvspP++BJormBstW7/jC4mFsjsjwcBKqnD
HJYTQjEeF4W3eWJxYTwx62D3/DQ5v2DhrL3IWOsZrnPJXLfwkgGZ7rNOshKIJsEzb8dySk9Pg8x7
dBwYOTLP+zYotbkrihuZ93N98sMIL3/QJrum/x83IxdsqX3vjIt4WyDn17yk7XiILvauVvYqxE88
2Qop6bbapo0r5SxLBWj8X8h9oI1ylKmog6CZRt4hop8cUnxDki9fVnwQ6aQEriVf2ErhAkaDYwuC
p9ElcZVLHafLaYwJ+7wXKVcNjbAtL+RyumMv5jJX1a23a52K40vL5M4sGV86j1TqloAU/8zK7AGE
GA8NBeypB7an5EVy296Rf/3bhhp+qoNmuojKoQ+E8Qt08LA3PJaOlgWqUe+SvwQ5TDKKmLeiVviQ
eZiOrswCuOgKuBMU+Yf0EIB5QBEDzQvr/ROrv8dB7OVTMK6B67UYgk+7gidXwXZq/9GL2jGcuyn7
Jry8K9yzIc3nGLJUU7/j9rileec38ulQvQaWZ2p+1lmm6dwkQShpTD5nUXl9h+hKbI7DvedFQrgI
sPWKy27il7SPo5ShNo0trjlRpLKLEPmOu+jImiUFMVYq5U1JiiEHbLjfDoevQwMtcdXjBL7+GKre
ChLGL/0MddyTDAY4jsMC++ZOcXCmImSsx71Zs7vsXcu5i0iLQ+LClViEz78ZC25W7sBaTTR/BqDc
e5xEOSkBb4yz3UgnbqON5ukG/AqFePlsIIhTignnsXsOGrdhQGvYXtwp+gtmT30R6ebN7th4tJjV
/BYdOt1pbGtAI6E9CwnkKZlJNTvGx/thB46N7FI8n69L/5YVX9+dLLeJkglCVldCEmSifeHeJUM/
9IdrjaKGjvo4xFAAXGWEquvLZOG3Z6SX017ku3E/kjHo/3t6ENC0VScJJy6oywCLMArIIuUAZ1xS
LYguERR7uNH0wZvvh5uzcNC1hyOQHbGA3BIqOwUNBZo1+oFBb92Hf0nxU1sHnZNMzShcV0rKdPto
dqDkc5qqAQ8g1zTHArIUYTYSoxGHSsWz/lAMllrDAUva77iR+HUkC/iRKqtnlcY72x5vndSe9seC
CMyFAtecgmTFYsBPM97t4EwlhXjIRsvlig406ZuxJmkGY/k3FMyp4QpcmtDLq9zpKoXMb0Sq5jNb
nzWve8V1BLrltWgP+b6DZGMrhGEJLCRjOH605/22g9k4jtGErnofNwIRxysgSoi8KFNJrk3MoQCh
axXA1jDAs+ajMIzNEVHMQesLnhQs+cOuqOKyMxCjI4G3qnpTBJF2uTBLMrPzIajGL7etmdAVf9nR
42qgqQfzFW69aVHcekiEh/pUQwj4XoTlvO+5/4uvkuS8OTnt1T+2Zhn0oBr4kXsYr2yOVAtffk6Q
ZqyIHev3vWkE46u2UiiPaHEQLFAsWlr9X5lC5RHSpMgGadwSKdlIL3fGFda3NV61KoHiSf3WtuJV
bFZcPK65bMj20SMo/IKRe6JwutO5R5znmW2oLar1h/PJ4AMrbsFT6bj8Ehflo89u4zLN24G3fRaG
Zc7cWa/tOnrj1dmUyIi/GcG4SBUiFMW+n7trsXnHwHtkZ+ETnP2Z6Gj79yBCloqQKoOF5eCnca/x
ARzl+GVYEVXSPEiMZ4YpYJsGjQQhVykr6X/JonhNarsiWU6Fi/jevw44rO4qnqTbWvhLZg2f3/01
mMVjr6Yx3vttJAMOIOC+0EHStcL0dF3ZEfvHdoO4n0J3TwZDTJ/hXQ3Ybqxiq9GOZoNe52Mv7YHq
9or8YCZrRAOWXSN0EApICIQoms2unvepkA4gPGuHRc9KO8JEMp3LP4lH4LYB13/GuEKD+RdY0PXi
MGT1Ck7lPSsFpsNFBWjrtY2vaKjZWhUSxZyNiy9VAbhtCYrt/4h5UK1dvNv4u+R6/LD9O1PvF4iV
Su1+SfgqJwPgFwwkGu/a+K1vVeHxaSaSEUgRC0mOos4VooJtCcBPsYYKGcRBhyC/i8tg9EpxZvpp
VXj7Z+ZtnpK6gK4IWdPjHXC9EeD8KLJrkBBc+weVmNA3FHzDdgcYc0xhlFAL/lOKUzHx/XOpnxL4
AIX3aqZSXJC4Vk4CiKMeodkWxDoCBzyCU5EexevCxkpH/fRrLBcMdZl0dXS1I8Vg5HQhLKNbIhIe
h57459LLs5wUsQZpwb5j4CRo2tzoeSjf23JPyzTzz6mTGUA2sZB3SG1N7V5uzdUTqk0zgZLUDb0g
jgoUbHcOSUvC+LFTZZr8UPrNxBLesof3jonPXSf35sTGiU50r/2f+dhiF7a/6cqnw+EWcHz6umU5
y7BjeO2atGxXWjsEl0k6GXdtfUM4niL1HZZ0dGytK10OpzNfEhnIbwfDAcEIpAjfBIELs6917APZ
DTFTwX1DWMksGJQ2pd0Rm8cLpco018pEO0Q+y2PWX7wO2w2tH0nArL/iaJMkbZ3rwpH4mHguPNA6
a0K9RTe7gCrn4VQhJJvDkhQlPyqK/W/U8TPifGYUQe84YLCS3/WRkL2cXUGNjmGH7KIVCmq2CCeu
xNkIs1UaLor4qRev5SEyi63emDyQIRICjSOn1ixsVaY1RGryZe8nfYCBBRAIhkOo9xaFBR6CWeOn
+DAoVxVsqkm7xVBAzB098E1iEr8oCNPrqBAaskWiXYpoUE4UtHJMdSvGfft8vUpi4Hs9vK1d6pjK
Q9cl3horUzJI3hT68HYdDpb3tyY0D+ShKFg3NHendMWL3mh+o/FcFCPj96Mkz2P+9LH02XNnBNvN
pri0TR3UUHY6E0AyT0r+HpzPEzNy2Tankzc55m9mc2WMX34rRx2eUjcMtPIkrY0qUrR4uSJCkxNC
uiqchat1KLsdPDsoHF7ecVjzvaKUfci720VbLq9mzJHZnZcdFVH+di+oCHcwjaFBAA2Ms3kRaosS
qoPx7r9eBoqqTwL6lfF+ji3ITkTbz2LUzzesapitK3qSTS0/wRSHYaUXBxA/FPMnoznWv/yszkil
/tIPo6WpU5Z8pffYXnbABz4iNdrOflZh8/HUIRpWSuF7F38fbWpjMpdqdy2C9O6hJ4m+81f/CHJh
XkvV2rYFsBwoZqvbEiPabOXHCVwgHDdVGyKvkeE+/nmpXQWoWo1Z3kWz4oal5MUdPeGQ5H1ggQ57
b02dWZdvHtj/B13q4iJscWS1f4mVg2vk+5a/PUcJWyBJ+iQIlPWm37P+RL0Tqz6tNz1zr1OlTCdm
TkKfLaimhHZlIB/9IOtssTMCZ4ZGBrMO3HphrVH5m/7ll5zsc0ID4yMip89l4UFH01+QuG0q31w9
w5HIIEqSudRed4YF9RjMBnm/2Z4x6uX9lN37EzzCJQesmGvY588vwNugax9n8mDxEqbM4UWWKQTX
Gu3zlbDdicKmq8DzG8QLKfNk74K1DsOWnJNQ38oGlZXUJKqHkHBIQRtf+ommMvU/vm7K6mYzWC1r
6fFfsync0JYunt3QbeK1QOan1OVl/sjxss8k6byDscZBd9Ew3HwxOvJb1WjhQMIO22DHhqqNzpHH
uytLHyRSE26rLr8ZFIu+0ggJHCu5cBEU7EN+WoeX+pPFXQZMI4/7n6l4SnoHu2Nd5h+ZbQhBCmsI
ZfqtCg6AYI2LqsaXY+Iax1TW/5pBA+06RkmsB51nZb2ykvZyU3LJ9ZHs4qDrPUzirc1+6NmXkaqb
TQ18DbDfVgk86+TiPP3AsHvHY+Vdx98CqJHViArcOZ1BoIzukBQe87FghbXrH+uxRKJF4vsE28tW
CwCA/2dsXxsh93Hd9oMk9EevH4oREF4EcErfZ/J3xQR5gfBO8OzKNK4BuAcCNpymvVSBtFJEeUe4
qdkouJXJtgP4XCKLhloRb66SJiTT/OT8JF8ZFDSQL5b4a58OZD686glkUov1qZ0gMuZegLxA5lfC
BICWXcbBOTr5UzUIRIXlwCGA0H6iMObMERV6Nuy+CYdYceNUmulksum/W+AyRzll6tqpmG8cWLp2
9Y0/X0gpW3Famd5JFzmprh2X9ShS0csuAFPOPmGvA6652s5u65hoKCE0yBTYFMpiEhupKOprJTKx
qw7/3SNrw3YRCUG+uW50sbBGFilxOvpdn/fDzUr672FSmbEvhHGaF2pkQEjO6rSaKwwq3vF2YmoB
79PgSv+8nbknaLtntfZlIqRTXdQTZwEPOcbUfIzVcF9ZiPmuiQ09k44Z8M+JZaGveiFRaqSwffAG
2DjKrxyABUsiMc6fPPsqHotjYGwf/Q7lgqXLii7mHiMYkLTCTkdwqmM7zyqYlhszPSCwcEa2FAxc
8V/GnL2dbtoTJ2TfjoNE5QXvRtGZsDNO4ePgcR3BPuNxMMyNE78FCwo/M2VGzqKO1oP3dNYQ8M0f
NxUthlO4nOiDz0+AZFR9KUjvaBcLX+0w0w3BbtKMREC224CjPTKGusPrkW/jSC6LaE6lXOoXNJxj
OJ4xC4sD5jThSGwp+Rc+DZKF3cmq45Hvx34dYJNoV1HO4bdY/B110a8yb/jX633R6j6D7+oHnCeE
5FVoqwB52bf9Lkom+OtWVfCsyYHLFiXlEes7RlPXKiOochWuyqeCUPP/oKuO3pK76xO6GaJ6eF3G
w2mm5VGF2ldRo22+H7Qlki/GMSCo1f31lU90oEjDa5QDkbJ1J9IM4aS8Ita6lJB7ib0403w5xI9s
cyI1pulDx6++e0d1vQafCl323vRaAoNCuP+6elALQF1MuPJ2PFqG0TlSmINIa0wg95GBdSpeA1EL
LXL57yKsbfnOGF1p0kqHMjMkS8T2gP7VdQMAwtnLZAUvNp98uzYrry4GPqV/H8WKMthxtfzKkLjp
c9ZqV3+8mzHZdZ77iSFeOidnkM1Xm+P+A6WQvP+NQ1d1x/peGw4Pu2Y6dEomdEFxYDc4zImnKo8M
Ux9lQ8Cq//iG5tZOZ9e1FhW+pZd0/FIHz30+fYR5dxMcBQEw6yy8nM+aNFbV6QRh/juapVMt+9qn
yyrg4APNDODn5FIU1/WHWIfseZBByWX1cGbMtdRkakOIiAfKhnABJbo82FUDUpsEGAfWC1kOwMCN
zmlxQcGmEcWjQG1UAviiZgIjHQuGOqZdo6L0XzUvUve1GV9oWQrS680Msu4yG0W4vs5XVVLoHyl6
uYhoi98hsNxygN0E21Tr9cueOtiPPnn4OzmdGk4BJAXNshGCEjR5J2RzxLaRO6zhuReA2m3cyYQQ
hmmRfyU4fLE40i/oVLyC2wwV/ccxDLovsWHstG1JxyiK5IbvM+EXZR2LyaFjR9PqPwe3kh18IKgK
VXUf8uSore9FafYcsirlUGCcz4WWgHeaceGQ1OQGF1lagLzbNmisdh4HmpTRrwKMiyEA7bAI4+Ro
k49/u9HlONFTY8BRsyfyWm5Zf8fD4PJIXo9IGCFAgwwhFoWpSzvFBt8O5xVYP3MMDfWWNaSrOFhc
NS8WY1f/RM1FMICFvYgsPuBYvFaD6679Gk/FfB1ZSPDLmj8Xnl6qgR9k+Dwpat3mphcENHZ26jdR
uKgIp8IbFoQXHBmfLgLlJL0DByHmfrdfsZB61UKnhwlhUPhCqAm1AyJfXIPImfTi5xGxsPiEi0bf
BCyNQOUK+ipbmQAKHwLiyTjBNKqrpCfu5Itvj2ewB8Dr+J+SatjePiuuWlIEAoUAzsDDDGHSuvcP
USJmXERNEODv3JjWs2h5k+gEpUGTL/3vkWYT40JzLfkiW1zNL5lDSyoaogk1TS1sFaSBMAtKiwiH
aslQb1hPDJGO94DYhSFLRO9cAdRUgfar0u8fhnb8mEbBTAEhhC9Q3Dt/kQq6s7sZWE4z5WIUn1V9
hihgEiqfaDicKIxpNHd2o88mCaQD2lJDAXgiO6J9nPe0rEKpSpO+eN4F/rjL5VZcxW7MVhIi4on4
mYqC5Xr2VZDX+qE6k/rRp1yhrmE75ZM46sdLT2o3QlNQfPQfp6tu3otaJwY1y4BgpVgeMbdoFSdj
dH46H54B2SxvJ0n6FGOnZ/HnEXEPC9+h0bhaH+o3RLdxhF+8PP/hBfv4unoSJ1g5gKRN/nzlPq2q
334ktZanWpHeLWyEJ3WbDY4IuKpt8tyDBW7qvhI+pjeX4D6kfwZjmDQApbblQrPDonSkDotMNACl
tBHZX9ASc+y+03PF5X75T2iliVduY+++cFgAAKoG2BQPXhXVKWM597tu3GueclCnUUMUNZI7+LTv
RdrTWbF/yT0RQ/hCJg6a122YdFxAeQRMKUjLcR/cInEUvYk3y5ZDcn3EqG4Du68YqnW1fXr69Dcd
LAwL95/4hSKEwcZjtV24ZjXuq5AuFkXqYWI1oWdB/QO0E+UN+Ph86FKLLjD9eVIcc2Pbe/hLeNg7
s7icFdAtjMSuU+EmZrSZPxWGpNROA2lEmONcuG4mtWMlPhGRy2HhSxKcIVUml1LD6MT7xY8Nw8uM
s/6iZb1KmUks7yELgNe0bAik2nX6wprjxc3vC+RC3GkurnddrrBbK3qxvvc1eCa+TXh9wnTCsMZf
9/9hHC7FfuvaYr9OoD5o6JV6XLhHGEYje9Eb9PFOKnwnEn3QYmnLnqw6nbojj6xoDGpxdfhkmjsr
nb28l7fRiTg45Qrkcu12C4fSKxmEule1Elql6sl44IIESNzC1MMs/batoyo+8E83yGWwCzdlPWH3
f4Fu/LuXgXtt82bzqR1D3FXj3RxGsJp6SOTDuRlDKjfJ0nmVYWH8avdCgaupr4/yy+9kdbHBl5qA
hVOtVPox3U7BJKMjiCyGEInrfT5ZqbOVD17E657ViwN2hGhf2x9vdYbm5i6rjqp8MYnyPqAnjVuD
BFuHKoFt9lnI7/h5JhP0ifc90mIfI2X/OKkO8A60Ve7jtXBoTmW0wmEmVus5p7eIJ6DCwP/2ruyP
20jfX4BQPJEpoHJ11Jt6ekEL782FzVkP0obfSnysRT0AQaxRhQBHT/Ckz/qB1q4tA6d3ahWO92Z1
14B4OpWLmmugZpHYCeUxJxZY4tf9qMpK05MuJcskpCnU46AjulmQ2beQVs6TWlbi1XE38CuiFAjl
a0WUbba8w3+pUWu6EYIeYFEupBRDmNxiJFxkGaOXAbO+HYZ7XBy9EckF/G6JBbUPRXl6p8jfswH/
ehxt6wC2XX1snwMpdY4VdkdEEVh3TqnA+ofye3+DQH8e9GOQgX4FGX7nHmwar3QCbsE8hurGsytS
1TAyfyHvFxpX2HTLz/SwmS567BGcemxFGGU4+Cl62oBA+WmwUkgxMB/SVc7aIqXyYa3acCsuJpOj
dA21bbhoBT5u/OBSW0a9dS9Mheqy4BuJNUpFxHIXZmGdzyMbU8QtmWjP/2GNfBdzPDj2q+P3bE64
YweesksjWyOSzLrR9jH5J9Sf+RmRfGXxcEjuY5I5iTDyzszKgraF9/qIkAs4IffV1LmILPT7EP+y
CZuXCHNQayxTGK3TlaaXHiVXVZZTWovbhXpbniiSJBh2KBWxVBTaFQw1JBCsZ9lYQel0GT/8X63b
LB5PIIqfxW0dv9Xo/xkzOQtbyDRcvL1idOr8ue5YAZcs6ZlCAr/bVRNajwgOYPCdP6xI3VFP2XLq
d4w0u5scJNDiUUz3BSTpjRCtqt9wsLvsTirp9bIdmCtKmiuYsxHE1Objojfamx8dpL6KpV6evKeu
FpfVrLjeJ4nO5Dynohjh3a7FMmFCQTbHxpymYcvQklMayH6SD+r4yAX4vcRPuKn8kmBNsnYNKZPp
ef9p1utripTZAL7mBoZIhhYe1wFBSVU6+/GQBKhcxpuz/U5WQCYPZdv+Sduq4fZQlAHAIWZ5e3G/
roLXSXkmAhqiBGmkJQkjLOXg70YpdJiq4buk9wpOG2NF/2DSG3TmiqDWBPtunH3fDlmeJzpz54I8
NFUJErVHy//WNOFM2UNxVayrQif7OP51n5imWNfQYpDH+4fZxuROtv5gjABi575DkoX8ivxxmG9K
pdo9bbPN1npmh7mBs56CFwJhe4gfluiZZFrbLCBFGQNdiqmA5w2JvNK7Ckhps6nwoN+B078LpH7x
EHsC49T9BogkOYp0qJdOntgW8LYHtOhQ3ScYvTdOdLmsCE6U1LglRJ7v5DejJxCC547f4+TODcy+
ymH+FFHuEOwZqtqvHn1SNtJ1286AZ4fyGjEPKXfoNhWN1sof9uAXBvCoZjUSpyE421wa6QeuXUvG
Z53I+spXD61Hjws37OGLiJ1mRpE00ODCXUJHe/07HrHLQhMqQ6vgDOvLb0lsy5QLZrdzzfF7gZWk
4ZCf7tfKc8OiYTUe2fLjxrJd09pCpgN4LzM+ft75fW8lBT1PkruSa5eAIs9PP3As/nONA2SBoINz
RKR4rEzVAd4vY/W4qG6ULg5Pd0wOG0A3jpY1EJqU82c6e1adBuS+sxIXs0ucw3QEerr7QD84fScl
8Ur4pveka60LGuNlO5QUql/WPsY4xSI+E3la1hiegXxbtdbgwVLIXOy3YJwj9Uz70pMmJyL4v1mB
HZF0dP0Re1m3BdFqamv2pkHIK2TijS9IWJgLYzdHMhYpokZcyvZ7vFsz2WFszGAgCt1uCGui1KdU
JUKkfnBiVsrgG4jyg10wA5kEhIGEQsNBx7nXVoqpegatID4HV46xiVCtGB3KUDrTg+FaKw8bB/H2
YAm+1A+pj03e6KuIkBF03mtoFfCY2obpnWvpppcf8GekwV3H0nFJ7qWkgV1UyaPZG+Z98vrHp2qo
7WbKJcgxJhoOPGUHvf2GiN9xc7W+ZZF8F3tP8LZ4TMubAMam17RQt9QMI2qPsL/FYG5/jDzDKawJ
HTiH0jQyyRWbL22oC7vaINO+FqO15s5LO4NBcC+n4VyA8vaN7igE3HZImJIbWfQCR+JM3eeb7qcg
mzVqv2JVr6nfQpgDhYnmC5Xp554xRhqV/2vvV+5HQVsRhCmyL5t1TtzkU/HtU6f6Gnbdj2VHhR5A
7FfQ0ymEyiafGgL+pXURFI7ufurRJe4T//GgcZZTCJMUtX5F6muWS2RRkof6/NTd2nw2UBfmuARb
bl+aAmUbWt1Mw2Y8KXXh1yOvzIQgVppNrIIN1J0ncGBgH7pXz4enXDNnNzXDwE4KhaKjPmW0buj2
BoS5dnDVHBpgCzXkCi9A//CkRUsfT8F6Li1k8I59pTZ2p3xmdrWnzwxw+o/9UsUjV4fPDSsdt3AK
Cg7jbGQbh5ZjPPp+Oku8jo24TM2SM7NSeyMUN6QBah5ZwWKvwXFUxL4oBLxosChN6P1KwoyfmrPn
Js6e/1B6W6eCVQ2FX7ByWptis/N21kxdysaI3UeZa2HIVXLksrHMScEj3SUZj8D3vNC/pG0lAhsL
Kv40zxvHMzAjC16Szlp58RBnb6u82uSIYHUP4KA2ukxh7GaameURECJ++F5sUs7W6ZII48W0GGVd
vDBhwlkSiPCwdeFeM8oy+VoYsWNHod0yCm7h1XTgsh+WW+tYXjzGs+mF4HsNsCsnnBtS297WzAR4
HPzTDxbRUqOWD1HLIkz3bfP02ZThr0V9Y0K5fXEqkY1qFA/gw+gNXGnymjeF8ObMrQ6iJoUz1yKD
OZTTIssFfmVwU6NHdMSrwXJvM7VpyOWC+NjXientXWybd8U/0HvwmAnAq29FRNXt18acP0DIwlWd
DqXy6NjtBjF+zTiuReLEcm8BSLJbcnjrzFqy+5pbWa+2zwMI28Jsgi/qqjP7QAVvsxrJfojB3RZv
yf6xDqHhcAur6CXk1nXA9uieSHPkamcmZsNSN68o/6/Et4K0TH+dbdFYcSYFK0h4bKz1F3ebmSs4
FMK2P5gbVPtLBcy7DYm/8rZ51KsnZYIXlNJu1C48aqx/IhmtcrHI+Nyb1z6hh1/0iWON+PUn5FGa
jIMkLBy9kXEijcpQCL5OqqKL7DlJcGJFxfYkt+NmzEjZigDgLEPmfZoalN1ES0ttmw1oaQf0HZY6
ik5VO3MK/kOTmrqf/xZYiK3S4DYHiYzhbgYJvi4unE8GFVSi1hBD/iLIRgJ07eh7wy4n3/N1C9ii
ECHayC2MIZz4U+K0v1H/Vi6Yuvhp5kgskbCQdmu7Gtw6q9Cr/fY6xOvScV6MXA4f8mp8pSWvgGb9
gTPb+2yJlWhmzNa07iSX5nyyuEx2Bdjr5PYaO87uBtvNePLjGIEvHPN3sCKMol5xofYyO1OWSNhs
cM18BC6B+6cGvIwHuA3uMuxWunGDZnyIqKCRfgbpOA+wR6bW5RlcgxeVZz0MgVusk4Vm687CapdS
4MA9X/cI50NQfpJt2UhPfmbE6r4HgNx7z/m1sJln4kQipOdQaxuIZiNTPpo069B3im6rwiR4SnhJ
5B7NVxKMQsX00FhuR4QHRTtCCYtsYV1ZJCu7qDs4qLf2xtuhBzIgFceOfgIn2hl7Wi+EPvVqOSob
ho3OLHNAW5W0aEy6WRaY7F9dUFl8lHIFBeREghtTZZOUKvi3pDiAFAar3Mk0F4gIVL7u5p0lxrkA
Tc4EJbXtAla05RrYJGB9itV3iyISbIVLZjrGnLTs2YpsAOvvSnVQxI29T7/hTo3G1J/kicZj2zl9
WlVoC9NsJGAoTd9tp5QZtTJ9ameLlmH92cYxBrGJh1ZgVtDJccRvbxk2zcEx8O/Ztrb2tpftGCgl
HSsacaa1rjhZ7Y/G0wIebiL3Z+fiaqFvv/gxMx0aGjDu1qtVdOJDCI3bC1vPF8J5/9tJjMCrYI1s
VnM/Jzu36zT0gihjYW5Vt6RMZM6Sycs/40zIEPUUmKuZfzFDEzmibsG33BvU7qzTc7LYOd1o59wY
n3PyGWGXk9U1ejemCqDVyIt69lifnF79jU8LS24k1ZIqRTiWApSZBvynsH5bYKcM/UKYcy1r3GoP
XI2awptlUBktdmNYzqQUKC3u9FoFrnyNG1rguqhrK45ZeGvHUQgacJEEV8HNnBhTf2VqB72FLVRt
VrTT0Y70Y8UNKN6w2pbrfQGKpdrDodBF5oVUS5rCovmbJWvEvzrhkblsv1N9yP0EGMFTw7v6M2e8
nZmXMqAbnoD4ic2Qj53SQLWIazPUZup42Xf4WsY+ZA3GeVKpKMUjqoosIseqkP8OdsS/R8HLFx4F
ZNuFk4l6FFPsO+Fbp/kugv5QsdzxYIl8d84giQ43vVyOIK4DtITyBWM/No0dv4C2qpQxK++SdmPC
tDIVkuQGuXHtZ676M8zyC1HNHNKr5YGJOWAvqI2gmhpnjy3XICNOAes7Gl9U9k84dajL8zUfwfbc
72u5LuoqpGbxmns9G1ga19aohNttp8ctxmjMSw3zrq4BeFhVwea34fcmFPvBoY3qlTKFhyGC+wK8
twqYamJ7hQ26BINSSPvQoaaDQwC9s1eRoV35LYEZxaVZ6sM87awfaiSa7GipNbfjA6aUWYPsOSyK
xUGxtEb5E+LUYT1qS0cfOEbwlhX0Kyy/vC4x7RQzjLxJP1CHWZjldumrSudwPREM+g/1KO0HDwjH
bbN/8BB3QeJh5LrBpMCVa6EsxTvUxDAdnYY8ZqVDHdgziGY/Lk79JSzTVp39+P/SY6//Ap8q9UTE
Wxbm6we21G8l+kLISSlkws4lKi3UdTYUIqvOS3ezOR3IyWluh0yq+FpVfSNzpAZYnU461l/B/JjJ
UE38FqT3klZDZcEv3FcQdmqn4zW0cZHQir4x1oLaZO1+abvx0/y+G0nhuCVCiPmEFV1b1Dx/yVyb
2SMxv8XULAxLz1/XVG3YY42Q6aNJOBN5SUF1dXCIXrqgeUL9aPVc3QP9iz1mhAi+Y4U55Gvl9jjR
hVNZ+EuF0X02GTG/p2QfhCVlWlSiL8WTMYjSUEe/E/CrHUi3WueDBj7v/Q8tHvMDKH5vfPK3KDEe
pewfqDeMMK4N+WQfhtO8aREGblenljmwpIX0nEcnCZSoVkNY3LcROoVXVveOyFvy3Z4hw/SbkDjT
+1NxrU/xJLepFYsJm3TcEWkFprhf/90z1vxII6u7RxPGHwN7ProS93NUc9lKDHh45V6XF7jYBuzB
eaVA0Erc/jYDploEipP0u3YtXjY9GFYKzQR9KteFb6HRD4ae4dSg4ZxJZb89nUZ3ixHEreVHnHbl
4AZhqLEeBf61C/RNnQ1elubDKcLAOY3B6ASg+rq8/cBqI44mkPx4AK2gdahXly5Lc68vgQfDbPc5
/n3uMrHG1n8FP1H8bC5u1JS+00D+r4KTqCJxFMxUH9tWWQJEFqCEWjV6P9wJ5noVhS+7F5QsoGbD
pUtkZFkt5LaP+7YwSVWfKcTVzQk0JnO++DhQZ3Ya2FwSH/W9cYtOIfVUtO4WJDMfVt7XluIlTzZw
4BkEfh/lTCSREarMK8/HQW6VNir9ubNjg/e5i2unD1YAidtDaTnAcn5puozNozdUYd0PSDjZdi7n
uRuw8Z+eEkUbN5GCivp2uAl09+EjanFQctOkp5+ANrrWxU+zYTRbc+LhjlN6p/hlxmqmw77flt3U
elal4OZc3zI0aJMOHHWqef70EQZvpuNlRs7oZCWJB3Px8uKnfBfEhShljXEAnEU1W65TXVf0y3BD
le3es29r7/WZ6BLi7R8zBw72BFoIE4MVZT5RqbRwK9apKjbv8wC3Cax/R3ZPVOl2nsI1qga4strT
Lp8NTKySBslhsnWX8ctGr4Pd8OEyVhQFCidgT8JAkavr1vrT5jr50lHxPlygz7pVsaKkl3NypLjQ
1mSjv94EBQZPJix9P1KVXTs9zWHsCRayrdt0SZQFnNQUrHmueMBRC+zr6qw3UFpjxXr226RXr/cg
O74Jjh+Yx7fxdxjYF0nc8OQmrM7BjRwwPz0ksGqcYagEUtMTgE7PnD78fVu6M7LjKd+uT8NxYoxn
u+KK0YFqFqegZnaPMH3oTqU/NU8UCftuA69cuUoyJtc77Rb/QlA1YRB5hxV/b4o17u2hltoHW9qc
finLKlAQI0ne7hFwnqhlqGl+uwV57MiFZOPmHL+Kln6oLJy8Mw08oi8xn1JEO4J+yFk8OJqo4rQP
OPQZk/w9N2TB1LlyqHGd0uN9aF/Y8WWR92O1EZMl+bCm9+YgVkyBsgToBvWLHAIS1t6Psm5THc3s
kNH8n5XOK7ax6whO6Dqtxop0UgBeHKmfGhJX/BdnlElQRqhje/asd+49UzvYTo5iFjA5olESvkOl
DaykKmMA46O2KeYSoYSoo0LWlxdNQao4ekRfcK2juAiGhBdz+7m5tphrHu0N28Ivy395g4m5fEpm
xA1iLu7sTQbbkLY/2MK2xgXsQ8KZIG3qzFWcCe3HW1Th5f1Qd7Huf54373XrSfwMiOOqBWGZBYWe
LgqePccGGH6gzmuEUbEXzbh/6uVo/Hi9lzNLgx6KCa0mMjzP9ieDVQO9Kx1275Yo1o6Cv64u4tr9
qncMggtN684T/mLiQZYopH8AvPCfqU6vZB0CbPnCOJauVQsMJfDzT4B8VIT+vdvdMxwTmbq2IHfz
hkzI/X7GfDkRZIvO1UU8qAM2podIO0Wf7Vj6gZ2Z7l1BrXdFGQDdgZsX+/RtLOsyOHJkK8j8z9Qn
6QNjnf8vt40V1eriJ9Qxs7lRe7fGV0eX7RE1f6LkGRrJFvGR66nx/fJi4fRueZn8nOotCflTnba3
HBETWbHdJXrNv9PbV7eA90dyIFC0IUbEiGxOMkGl7TGSeVV+xdmdpKsA9QYhI1DKsVVB4NDzbs/v
w7wgbC8JNq681RwfdpA/NzdCSm6yTREwOYMBdbN6ChfuU/YYVsXhBgdcIRuPYD+pydjpu1FaAmGE
svDm/z3dCap1MN89ZWHhfv55YTGpdgcRfKMuxuTlpw/yN0hXSqmrGgeaaIBBqKxk/FbK+h77Xs70
svDp0OFncGaTpf2a8rvllz2PxCqAGWf2Wl5Rqh2gK3zFEzknKeaFZ8fmA9OKg8O7c1ITM91aSMxS
QwdiEg9XCDlD+XjmP1X1CcFGyfR9oKUCr3hw+q2Cr/tKA2nsbcjF/Cbtu0wcIcnrHhSdSY6g00lz
da9lhhGTHJeyEb5ACqjsX7QqHKkEyjeFUetkW9vxjKg+hMO9g2S4OSJbIgbX8O6ZgQ9wJos8i9y6
h98JRiyTEIrOCDObjzPgQPB+PuhZBwOA2VEkLgsIM9TbXM+02r5RwCCaWMNJhuscDlcguZ7HFQ1Q
4ef1paz8RXrKNoNEWQw8UJ4eatWgmtWQcRTo9RQLd6pp9LLVuPrYX0SWumIjldfk23QI4BjTAami
OjUFW4zJdPsb9rHvSXyHtw7chXrpUDdkUmRBzkk20H/tKzbhzSt5NWNuQ/ECAZZI4Lfz9cTsov+s
udwcEXekWSUmhhPKPEWzgIx9taMfji1uARvGS4ZZUYkdRSghpmXsHBm+gGFURJUzb6tQ569zZEOO
KuDzeD+v73/+k5bJaKcQZU4e7KND6KACCn0LlSiJ5k+bg+gYi5dZk9EmqJ1ZkC5GksQx1tMwbB1l
evA6opr+kHadQWJjdiDWWU45falA4XWHnXNKdNMteSlWJy/PRP3d/iGjQvvr2VtvhGDJRaJXq5OZ
Kgffa6o6lCHBtGrrVtTE027ru3jcduKD/xjTPXykipB2K+dvZnn8S21hS5Kfq1Ma958GQUBdqK/K
YUkd1TghklfYrNy1RXF3fUsInLTIcZTU0YEMta9dCxcAWJWMBanzmWhlNTkSZcp33Yw52/Z/IdIh
ZnxBHeam5hZn+3RAxINpxSZqXHrZy2nyb4vvfyzUqtmVrlIWEq38TFvIoPJIYsRsOvFnJiT4N5zk
Prwj3j1OyGS4TEgqmlThneBPMJJkJv80vkQlEW+H/5OCEMGBVba0BVQfPdRNPpu4Sb1E9Z5PK3od
kn97UIB6v1K/oS3Pw9mn4J5kue0u6VOIO9MeFBtTUVvZz/15coSmps+sB0G7GQTDajmBwNpf8KNS
dx2nMvSq/yurCqSWIjLtwNOLkHxFu9HF+4roJbweUkgtPV1wOyqvxysDzEwQh+qIuXd8PGjWB04e
dLiOtKspn41xg+F4C63hd2GNgPWxQCLuWufOi6H6fVihKTUtU8W25F7gk9LT/9ps5FWaipURLVsE
LMwlxuhgqmvOcQpHYhDqeI8g1e6OQb5RhxLTQHgVHxWkFwT1xlBwrujBnhvBkP/2Yv3Qbt19Wgcs
9Y2P+cpDMyegYQi44HhvdrtiOmuFLUtkbXnpka8GYYv/4M317rGYpyA3yn9thYBlZaztu/1zl0Sv
2wK5n/QFjov6668obs6zGpjDufXJTSNtZEcQmUlbgjKl6t4eXDtW2LOePWZOsE2O8Fnf58dti/5m
HTRQXbOpFdHx9VXqUcjANPOv18EpK2H4f3iezEtmC7vY2jxrOGLYE7+H+5Ywuqbb+C0j2zIdzDGO
mw/f6WFRGWpE3IA6KA1Z0s7SgGEsTFKJ+Uw36SBwb/Um+nd/Hhd9q3Nyso+gU0Ovw9J+2a2cHDhE
ZHglNAhJU6x/9Nzgw0J7NaHk7Bu/KPzOPORLS3hNX9slqhVwnvQAP7Ghmv7dqsevATInXn95qXVZ
Z+czZ+M3Yc2ky4r8psQcbJYkdfBbEWG6PJIsefO8KctkhzMsIVtBQBSzAbbSY8k1vCCB85Ck3CLE
Wjqer5UgJmz2WuibT34c7MsbGjPkVxmf+IwEIxhKbc+gjVWirw33vU1B8w6FfkBqzr3Q3dPSgGBK
785UhS7wRAjQioob2iY3O/GKznQ3IY+gyKYgS3a92UP/0vNt4sRUM+XbKrgOa4xSDN+zFWI54nZN
l6Mfam/H9nRL8mE2AaiuFNZJNZnHqXejM5tIq4pImodZDX2TQKYIjamFfbjhU6j7xGCj3YDrvckS
9ZgT1K0vbkvfYxdnRUXu+U3D/UKC142KbHDrZOrnxbGdps7aO/smk2qpGp1Tkm2j4eM+SgskfQ3h
kiRFaxxP33lxeXt4VkZVu6KYHvFtHaPM+i6V0R51UB9GyYPRFkUPB0MokOqC36jL3l+IqsrOEXcb
eKb/zJnwu+DmNvu/tQ9idJy4izsaKS4sQnbD/mc9AxVo6ApWfXZiu9BBJn37KQI1l0L3uydRKX9f
xWcsRUgNBogkP22HndaCfk8pBN1bJuz4TGMeNfM83CoD9xWW6Vu/+2t4U13aP9iEgofd/GzEBgoN
+qMNl7oAmQUVvNusSskF4ryUHkZMM5IyLDPEMPLExgXr8A35ZFEPr0wm3Xf1oE6j8hSLNbZHBfKR
CONwZO5gvZeTB8nuXJ5e8wnz7xEUX3Y93dyD8A5lO8QBmQLnMZ0xS79+DTvoWZ3eezERgJ8tc9Lp
l0hwBOEzr++Yy3LzdnkCEcK8WCQ1aKqE0yfrefC+R2GKq9JCK/akaQ1xXLtZXV3tMVdunM8U3vis
1+0pOoyY+3YIDbNraDkysZRKT4qBaU3pWtvMR0h4r462s0KFEO4TAdJzKR84mnDwH5QvYp9t9sDN
+hPPw2wj8RZlu4g/nxjYVs/pCBk9L9WElzRRF2RBUIg/yl3fyTKEUp0L2+3V5W96i5lHa9r+d180
ZqUTpHMWYn9TLesIu9J4s4TzKk4H7fWCznwjp572fx6GOPWS9v4d+nQql1xOXUzsrrAviRxo9T9N
W3zgGeBIXrAGTXu/1pcG8Qmpqh/N95eIm/v0TaRuZ8qX9XgKZWL1MkB3PUvKHp9l9F/Bfyn2I/F1
g2eGkxZtonh4kdJxuEgmOH2godfWBrE437EfQ+C9s3SO9/3puDjZCDnNxwSJBlWZHY43JjDn/n9E
645IhXpUzAsxDz1TUcFf5d95wbklqv5ZgM0YUeBNtC6gqbLFSvtCqj9tGOR8MMf7bb8k9lFyxMhX
jXhbQKHLR20cqT3CKB7Z7M+a0U80EeO7DDlbgO/ZBQCjBsGjzy6nthBCE+S+TB16nKiSnQYBpeC1
Q91yvx1PB0S98ivHy3b0CDe9TivfQTcT1urUQpseylxFrbIdxE5LQt6D0zS1kyKxecY0kDu6Cgta
QqzHL6Wn28HXDLHCwZwzjfY+1GvOYmgi8w9KZd66AGmvbWSSJgc52v3g/jvdmxjpT4tDmHr1/WwJ
LyYh35+ZN612NdX3PZacdm3ddu5pI9UOEDLu56UyLxC5Uiqn5b1qipO5jVjkN+WtP9kgf2svmUfq
LZdRJZMsblKZIm2HPhfO26mf6DzedddFva/qBzh7w3DzHUI+4HSsjbBe80QcZ3z/runXcLtd2Ibz
IkW/SwaUC6GV0WZzZAztZDIB8s8BxhIW41Ma0Lcq9XyKIh4CbbsuxznFxnDXTTSGqo7FSTFv+Qiy
ArBwdnX/9W6v8PXvK2cfw6VDVRqKt3FBr9itCbFFah8qnmuOG6wY38jc0SRfIdAIJ+iV95ppKYMP
a0c76XSpIi5IVFHTVMXlXot75EgqigcDhPWgEYO/UirKglV7DZwY8zy02iZOODDLNWq58N6TDgsF
ycn4C+n69uwvOujDZcvHXQYJ+0JcXu5eQZKkN95M+Ch3E8OQ6u8xVjqV4HdaS19OFfnSD6R6wy21
1kzTfwrXstwR2dNmWW1w9ipVgQFRg7or6eD0Zh8UyzO8GxHPfJNbzXH6lPwLcLGsYkpTpzxAGask
ExCK5ILpNzi610eVn8pT2qXbaZR+74YlfoSnXiIj0hmXPVQeXnT+o1Sm2vQErgJPeG8UaEd+udc0
2k+u404KxcWmRI6bwnr8lgQ5lihCglVbPSo2zT9nEOofPLhBevAtdfDwUZX3sYjAkCxt8irzhbou
fGO5fiwMOXvGr5BfT1+xHp5nMkCywNIrzk86RDRZKyoxs5VTnAokJ8x40A3DIuRExsVBG0PldIrh
YI1Wg0eT8jnDSCfuzx1/figmL/oWfYbF8A2drhWmWbLWAsxfDeWduT4Uq6v4pqg6Hv8Uxk26JOMg
psvqYBdDcP2aB6jGwwNUChpfPRrr0L5TkVH5UPxHIF2n7yD2DIJ57Cd/CswZ8JesKB/O56T0uyZ+
R1UVI4z3hVattdzV2g2hQ0qOU6wLMpVLuwQMZjkF8haOLokAM/cKXrhze6+ELqjKSOtjD+vIZ1K2
nQ6ciW55lfP70X00eEWoRnFArGGM8JvweCmPx6LxEYGYUTO9A+uYs1PFliVurADuvimtZf9EPJrR
WmO3YyMO8IS/dCoRkhCLKBvrIGAn3gPq4zbmd92gjjeRBEVHyf/PyTW96a4NgD57tZntKUw/V3e+
iKNvA9JP0TddaSPEKCP/mtPX6id9tjn3pWl1eYWaUeLwhhCSel8H99pXlgVeXOYCuo+IQZ2nIWXj
4K9R77UBtQUPXsVig6RABSDudmUUtjODGkJHszpF3nam08TX4HFLqAwVhT0+jTs29XZbtLEwRCwO
G4qU/cvu0nrkppIxHcCMYszQ0I5wiTudXdAQ3xME8o+RHsesMKs96nxz9deM2bxApq0HDgcU3wLr
t9vkElZUD6QfAnIpncL8Yrn3fJnGTLdqob7k2hwB4xPm23koN28JlZ6LbbhKSJk+9Hao80fT0oYH
qpeZCFM05wsuYaBBSxZuXXR5q98yt1RmMa6czorkZavg1T7/Lc/yZt2ZeFnzndt9u4Eo7ff6NImJ
j9gd8c/BxNV8C+x0WO1MAYGvaLStQ3W+r43SzGks5Nf+PYf4Pk01TrKBw8EXsHqBJsQKEBDxUyDt
9Dlt3UTLZXANvigdbktv3cry3C5kX6l6ctjOypXVT32V6ySnM8hJVFXJ5prbnCCF13BTiCAXBwiG
DRYL5fq3cwOPRXksPGZKYPNATmn/zzJy1a80JU4y2/ihHNycfHqjSiCAmphj/rKWTmLQB12Hm0Nv
lf0rELGSFdpsTyQ4HE+rWRTcnvmvQ+8F4CgGRkiq8sy2eeki4PQaEtKGY+AgCiDx464cv/TV2SqT
iUQ5WbGehPcmBt0A5+P/DF+PpEHP1q/0sdhIGFMbyREU6ahbmCy+xNx17CvWgSMIPdVMyKYfogMQ
r18GCF6lUoLQSTbTgeSfqufXJWoS9hCIEDX5hqUPBXVlxfm4kj2FPhvOcyS6Gc+TAKIl3ThtYepz
v2332tVrhzzRADodBVRmwU0FIKLYHDYXSwPTttiKtDcOGtb7mzRzz1szKQxMqxYw/sXe4qGipLK4
aSuysMX3EWi2+Frnhr9yO3B1emcLEn6fQZmIiYgyhma114ncsPGAnmSm831VFtPdNLXIWRod/j8D
LRhoKEiZLN09OvZwxFTvzq8aavOmEHKc33ZCbxSVP1yOxp6l8yYEgGrdrknz1S3lHTA1XnSgkEJI
YHthq4bSRdFg0mbTg/kNgDKUc6BLiCPk2JsjQd/8qNcjeZUmRAZl8IbJnBkxN22NxsmdR7ybPhBS
KBfnkKN8c3ZWzxv06+ml4MmouqT9FYYh96duLQwVqPcnsRzx+JptWO+pnBk/GtZQ+Ed99vnUnoCF
iANCwi4Ce5+fBBSdgBky/UV3aF+frTLIuybbSt3138kM3V21tindtFxjYyLOMItnbH9A8s5IwaOm
1Z9fB32g2ncg1Wrdtbq3fBKPvLAhaDFOGUMb7KF5WhKv5wEBa1DVWH/5yp2NxMmfVZ6FxoiTN6nR
XsdE0I1yfi94nca7p/7v62A7+E9/sJ2SvS/KZAeUAJinhnJJyxkqJPGewy46w316dZaPKc67YaIu
0cwAJiklIfcr5PHnFk5BbHGuRc4OohXTPmnm1nnavpZeYUjI246XOYuNYnUEVuX387B3Q07A1unr
HvhfzkEEqtiT8FDzyN9eSjPKbMtlMGG91ZgPMlztkN5DJavrJDTAh5a65LhPnxdUjKyWaFxJ9grQ
oePNrwsacAlFOBBkfiCgdWsKR3xji9F1JgY7XHYeGaq+KZ+FcDi0jgTolKD9dwHnk2fPcMiA5Aig
jgH6khGNfUOLiUdUnyDeAnqnusg4ydreSuXaMggDDiVsyvcY0XmcbM/d8njd4Fk3OuFBbRmfp0lg
AotklPaeLO5fZTa2ze2po7mBiH2pYCsvaSIaQ3Nauqwz65PSMlH1OjaubgU3o5GFrd4bAxAt3IDu
0IM9DLyDPnisYflNkgvp1s6u3eXbYrLpGQ6iyumM5pJauY9uEO9DFKBBzWudrZLacStMjpKvzxw+
IK2YqJ3F4U2ZdmQskBzhsudwnmJELUcLSGmYq7qRWE6y49dhLBqs0b56DUZldSfGv13LqjlCrbZk
NT8CqSWVqUoatU9Gnf+J0ynZ4LijoFGou7ig0sAcG7/jVgi9g/SjsO2ey8UbXg8FMAzVTEDGW+WO
xOOZRADdqe1inAfPi/eJ1i44XKr93LR0iS9Ix9WZPHJzx8N/pb1BjrGnumaQRh/J2mR9ip2IncCg
lOdE6IIH1CXZMMBsiiA/tNdySaSgwxN3NQ3tz+YULNg//SNvljND5jrJ+rRBKTSD1Hf4qR2xBNHC
pRCBhcFVXKNC34baIZSBPu3+7dsw9hHYkWLkjUqsP0/ZLrogD97UJ94+spI1VJMmLKM4+p53FNvY
KRucW9ChCI1rHMDg2oLgH8NsoUhgMFgOhCbykh9RAS4EAcfELfjmQvCwffBNcoEF0JCu4+0QZIjT
g7QB3bMSMaVpfDgbJJseybiLkJQcS1ajjbhZiMBlqavJ1eEhsXqpvEU2lLnFNF/EYcKKgcQ4T2YQ
YdMdOjmoY6qTr2OyfACSazaQbfofeF4zRf/GcW5HFZkX7gUMjftglcn8PtTkPybyGiKDx6WXIImY
cm11E057rg0I44IPTnPmsn+/SXp1ZPLC9ETwte2HYUg+l2Z2Q5pIaAbBcJFpg5QyY97OUeybutt6
HxAxtNvk75nuhkhGoCxjtIVcTCzkF+E5cfp1gdXMpIopFZI0Gauv3+QgOeZJzP1AkE5vqA9Kdhdq
apJ8GQuLUwPoC7Abcz05vWl8vtLjtET7fe305d3mF0F2roQxAqMeb2sMSGIg16hBoGFoIutqR3lP
OyGe0Uqaa8OwIYeK8UUt3UpR78leTN1nzM9Hig9n5zjphQgjgLlWplYvru4WPDOtTbNeQoAR2PSK
o0t0RlOI+CJw8t5BDKUbe9CS1dvilNf8R4YWaqsktFoI5kBjud5bk8Qu/Dg2+rDNwZwgU3P6QeAx
pnHjrGMzb/Pa8qYruhZ558IGDUgCsIPVC+OWYMT20uPOiXSM5gTUEf/F2gt2GYvvR3sBbQU4dQI6
cYqqGYKpkL3IO+/DTBVZGMlTLg+tCTa78bZB5QVrdp+yfY6EzjaSkFAV4spUD56pSZKFRzKHQeAp
bJuEJlbYPWkVe8EKZC8EZxaqKbTIcid+AVMfxZE9JuQvBWZvceSfg0xIZjLR9gtTdYy2XaqAdm82
dig3SI4OXB3eH98lfcbAjOB9lAXf6l7cEZJ8MWyiAsmxVG+Uas0J0rZnPGMk/65egQs3j5RxLLDI
CCkfn6HBDtkHBFRWRMPuqBSqXKNhH11rP15h6GV2cEZN9+59lMZThGqz1puFiB/eS76zKpF356Eh
4EgRQ/kQyZ/kyLAw1lXGhF6bBQyPbUNtBNMsbG7M8ZzL2VXWF7DY0pPCHWNT73guHFoZ8Q5TUuEs
QELXYRnutjNZ/GQpLchWLyeL2FiVzDBJUC//CkqVSYa3c80XQ32Whh9jpkjvHY1HQRZy4YWnF/m7
Q2QbOofIL6HM02jF98qyOAYcmNswJrJ0JcMg+qa9RPTCgQRormPV3b2tR3KbNYpfGRcsnz6KrfOu
4MthRA+HLRograKV8BCPO92MZ0uXgAkV4Yr95Y0t0m4Drxx+tIjFO/a3ciXCM1PcPeYsgXZldN9S
8cq9jbhkgcUCkOBlR0t2v+D7ydLVoMTsh4ANqPlRlppvTwAeoFUagrxgTgqNUiNIx5pW7WVY6ppb
94kX2ffX7ud4OLnnamAphegGqPYIJNuJ1tDtIVH4yoxy8Ku+fPUE0PZTTvF18XVLAyd+4LeOi1fQ
r3NqeiKWTTO367pYpGRlvWwE2axESYEMsNOk9c3H9+bbLy/KWqZSuXfwnEjjERwuHXxD4LJFpPSm
FCIJc4ZOMcAgwFhUHW7qssJa8UPl1mmwJ9dNnrbYqaJv/HYYrEkG+h1lh3LWLtIMVA+BIvDxwNLq
T1lbGjVWDuYfbpS57UsmQ6HM7Zz9OZIgceysoYLcqTMWwlMHrj5Q/ukzCCy7ssqET1V9WxvtauD3
hOTXe8Ih45/0lKQph8TXAD7M4rRJBoWL/oD/4vUHFJjmsHDdjiCABSwPbke1oQFq4Y2bBjRlZIRd
UKFY+xFJr3cOc6Dn7Y0jX5qoeG2MbK214Q91sKjEn1OTsXEHcPQWRe7Kdny+wFIZeQI/clhFIm/f
2LeHTw+wZaG0NbBauCNqsh9NeD9TRNnxwXGHNMYafGtsMjCezTthgNdt31lWYiECVm1yng3lf7Vg
tbvuV6IJeRcykh2DZ5YIOG+vWGUZmiuiO1wV9iWt8uvntnLUqJl5vDptHImhWZiA3RKyvTynDs9W
CPCNw5jXyfcSY4H/5wiatFeDcX4E/5G+NJn0R1kCig6NUNtsVk79UXsZ7ndCa3/kp+r5QSFruXsu
NoDAfQtQ9JFYFng4LTGhOaYMROzAGZMymf4rLRvVrHsUNGslOFvn+Vkew0TavGfv2kMf7M3bbvDL
u0Wdamub1V2Yu63czQGp+r8nKNY+h5m6qr70et35Av+1z87h7fHbKjItKCJuZPtzd+XHjbK5LEW0
ynd+alFdbYlYn2vA8FxD48bYRC2N6TPfEf52tLYBNhSJlqv5egfbXoeNVjjROz46ntfBLnOocpHi
glVqWmj5QMXllKIHQqstIt/D9kP3Gl6F4fPXOKtrQsnAZdyoqsi9pcz5NiRDRqbOI3DXQupJBjam
OhxcUzSIdALyJeaIIrtf/b5hej2uhlj25hCC8Hdi7MmdXHt+Xxhf72OTU/+F9+kJI+rQUl++xP0M
40Csf7NjkzZfzAuMtoVkUUv8SBwrwQiBRukQUVn3g8vEDu86Ik7aAH2iAR1FjYGa3G7ILb56i+sB
i3pPEde6AopxWgHQ98qfJeigL8oPYfm1iJpi9Gp114711nIqJK9PfEfrZilmGWjC9FCcS7oFFsRX
5mLM3m8ZwrowR6irnBIwF65lD2v9ISnxCTwge0kafenvYubyD0/suJHr+Nh1AlKpvnYF9H98ygXH
gRw6dQE07Q4neo0Xv18SnagYWK/pNH9SCTqW4z+94dd8Vu+SeLeyNkmfZW/rWFaPK1oeAFaPhG+E
Ex/4/rejB5Jsi0mJaN0Ivo0N+1n66kOd7O1QIWcMFi2dmDxa8pjGr0vDGGPpI7crqKh+dyo26TWd
0UdZ24tsDJtAR1rNa74mCMAR5/cMZxmq4AY7AYMLPZbSqWR0Ts2XYNLE83/EPWUq7lDEzeuRAOS9
3BOELsNB67zeXPXnylJGyDxVwmdc2WL2aJPsaxJKMHsg1vTo7rFdX5hBmwt7UEFvxHfixez5+k2C
EQ4G5SKb8d+opHvWeUjHo8Tvc0CEEVxI5ESu9GZD0QP9pP8zeRa4xpzEYXLP5tufbbF4b28wARD3
H7c6M37dYkZoxyZzvjAOOzDxC6iVaXjknWc2ysnqB/FqKMNSIkpX42FRf4hhPBs1Hr5ZfQMSXEw/
JpBQg+WIdNKNdyKRycMmgGi1C2n5W9ryvhqNWkrUaganHVDQrO75sXK1eSwoUX6lbi5xwHu0KibZ
LFIvVKYPqtQoDQVgTEmEpRakpo6krht50MI6VAeOVFaYCm2xWmf/atFPZhFfkbhA+PqiqEaRZtH7
g1Wp5I+Ix+4h3xeyvfBBiMumeWMMxMSiKyMqCMB9Sjw3Zn5Y31Rp0RUb62w/GqnSaToUWaQck5z7
FuEG1FQ2f5RyvBexot0WpnDesHvDPMRy+BmKSZ6m4jG0jo7bPTZH5svH+cQj4sqpupSRgLou9i0q
s4gO4LA9VZcN96exuUuD5kRxX46Hk5hkRZkekT4f4xKI+wo51zK/PY6lcrY9E2rbyulc6RjrIlMb
3wvylX5WA7e4LthkVXEv3mewg7ixMERmesCX8wkHqkSK3RsjERS/gAlY+iqK+yoO98oTgDJUKwC9
l1KuPzmUIfDi+C87xSX+yDI5y/ZicEQ7PabpqjHTkyhvhkcVFHYsN1+2VLhQi1/e1UjrTxTVkGtW
D2LL1zm/1IFnTT3iEoyQq0ubjQqHqob6hV4AWK35Wsg5UxlFIAr1IXPPVJw2p7MsnStYdpoSyu2c
uyZruBNRaAf687odgxLy76enXFffqIzA+mviqG60r1C5qfkr6l3h5w4sc4OqetxxO+eDj1NsXnWe
GYC8YS8MJSmJHwiP2mnzILpg1JoEgz3slBE3nP0Me7p1FJ/DhMf28WCBANssQ8pATH5K3QgGJODO
VEFq1mRgvth/dJnL2GN8pzzbY2B8Lzv9H2lzfacP55jH0eesF8eFiqz8jK+Oa05Np7m33j049wwW
4UqI4PPvfWhMD5PNqhr2V3g4PJ5cOYXpKtagVT6wfUVwywFx4eqgRYwG8A2KPixvQCuW8nI7OLBM
EUbY0CcUYtHFjfJBblDI/C0iFbKih/IWOUQhP857iFQWsMYXzSouMzp2ZJimxenDpvcod14dxmkM
CLgqJciJXJsnezEmjaq13wZeR3g86MJfCHo2ahMWr3B5HUyHNM9l/9k2IYXU3QgF8K7zCrsV58ik
sTKLTbduog2gqhATmfn9KR1UneWLucC2SSi2DfBr6AuzdLaTieRyOScva/xnqndD63ZI25KFLnTm
/iYUQhOQ8jUvrwDnf41SDtQgVMrAzSk5SwQB7QZm796n1QkImPwP2pTQF/zgBakq+DECOmzUKNOS
iIxeL0OQLjXpeCoaqorNHkytf3bcyfQ1VJDVajtegWME+FKKOlt1oWNYc7aOGUNEyMIdF1kH416y
vFg1pvyMadmAJJbZ9fp0MRyWVzX1R5H+20HCJgVRu8QxtCDRJa+Zsmr4yPYPVsj5eIjZ+Z4IIiP2
fLVjoU8M7vgmJt8gLxJ2B+38cGrsH5n8lS8TWTeqK2civu9GQjvIbDP5utZjYFVrlpXA9BPs8Fhi
el7/SYYVhPP3kVVAzYXWQYbQ1/SLbD93s5IcSuLdJkx7tVq8GNZLmUR/Pv9AleKUf0+wbg7chLE0
7yD5Xh3+eu4PKIRcFpUp14Z1CCRZbnbmwZSKdL8pQgG9YOCmbrorltGlCpaAQZp4vuMOVTkT0HKy
VdUYE3rvJpeq8ATea5cSJh9Mz/wWtCwUQdYJTneVTUI8EzW8vVqCMQb6dPnv3SBViFcqrb4/f5nX
GKj+Hm2fPWuGzASoQlZ6O1cWj/Yt9FFGUvoIgu8OFRvmXlNevhIpCclsSRsajvVGLhoFeqvBhw/L
5z2UES/rA+KvtywrzaoxcPgFQKzhRxe3zd8IUqlgD2AaQrjtz2LWrfzSwQ5vAWsPH2tVI1jsC2OF
BmlCPbzL4Bw3CcXLUf6GZuqW4sK7raqOkhXOufnDrRSCIEH3JTak3kR8wgGA528mny/5WC5UztF6
u/rxM+tiqUoRYk0OKI8YSazWENnkXklznmcCvC35c07GdvRgDwuV/7f6LVu/4VR8EUN/GjuRHnyM
y6hk8W1dmaFEHWIlMf5EwvQWKJ3K169LA3JRXmfwl5ma0NXwQvxydX+bWMWoub6p/2LQfW5cRbZ7
IwApNoWkw798YznZVssp4hAlcii6iEWnCOJYSLs5Z1n0OrVTpXTJeQwOXB4yWj+gb9SH86wyoRSW
XVWvdVkRs1bPelQf7lx/esd4YKkqMmff32W98jX3PDILc2Jzz+wWVGlqfoqxpqtH4q7GCUcRFIea
pEgziXl6XLzYoMh4kOsLBL+Zs7zJ2QNod6xqN3RMCWiNDHlSQ9YiAP6a+iPbUoJNSRApOZ12y5tz
AtUJTBUIFX8LukDG+PrxY0C3dvc/5VLw346wl9wuwQfEM6gtb+Zlst4wdTdv4pP15OzzemK3YU9c
PEgWInw7PKjj9w5MtOpGLv4v0aLfeqojMCKZm5ZgAKDN+XbGiX7q2++elpl4eR5A1v+PVqMB+an9
NDcIFJ5/W0HmtIduHcu5+tOm0tktXLrr8ysyGbpTJ69hGEMZAsc9beW0f4Y9okAbHRisTkz341kI
CzA+jzuC75kQ9lBKkvjBvOWtehGqzhAD3zp22wmvYiGVXlbdQCbsbcglHU37+mQfdat8jSBJA5W1
5iZ/ZjQL3++1xxv7Q5Oo54d6hAVgGEovMTPidQqhdGcA4QuRcdR6wOswlR/HjJ1qf2rgh6ncwUOn
gQauJk1xmR64yQpWt70NQqYVfzWVIqrLK0ycogH1NrKIDgR5g49XYNTUPfems61Ib6Ma8F7vlfCq
VrnUfLV6PJ6+ogQTKgHBZym8cHAKNskgUJFqh+mymffixhrwPs2/IQpcTIXWaCcXKYC92oRowh6w
lsJlvGZxG2/DnmARugVA6Tw1of7OUR3RVQ15fNPagosto5hbFLlKNPprtyuwursoE6L4Cfz7hcd0
LQoXlwQH04Xp5h59fm5JTXhL4cLd721SFksEFR1ktYKarASsRwndJFckHkXpVIsuYxP9z9LA+UOP
fv6GQ1nsITQyZfHv8Wv9aenALqrbCNgPc69UGvPKyCWaa6kVsmB0GLC6KBWu8SbnL83g4VU24OXM
UmVJrxHKdjJaPQSYAw2qjQSDWhRk0kSy5ynTgec+HN9C0Zz6mwZ/goHxv87zt9zVApw6uMQ2R2uf
mJmgj3t7we47lsxf3maLMRf73Npef39lAOSizRCv1VN7JdNE5w49x1C5wnLoFRtNfcjq3UhE27V3
qhNof/CcCOoce2m+LKAlWRT8QPMFSR9whWUY5jUXeJ1huOpgoGiyalhNEIykv0Bs2PYNSC7HuYdf
RHxBifquvLXSriHr6bOq4hq7ruSB7s5A48RAblh4lrRAE5phh/eHnzb08j+ZWZWQg/OW4vIHnW75
zVZZdDZBP+KETXU6mEuMfu2tQDjpExWd/Ug2TWbq3dGmnF3NGjSQgqCfB7OhBixW81TcFwk7y3EG
qhQyDmDhwMMkI2ZwbiF0kgfZpovSkCLVwzigzGmq5h70iu4CUStljhQ+fruBfEONRPQ5gjZUsaO9
jbE5sRrJqjc5lOvaTy/i2ViakMy2qBrkKQIpinFSe1Cr2CIEAVkg6fMJ1p+5FESQWLGA8e6CVhyK
4Uo+rqVM1z6CFVhuH+G6PetCA18KPGwh7Ush02zSxnl/2g2ueeRkOnMxoVvvM5GxUovH9mz++fB/
bOYB/WyfTBgv4MJiDMz0hMpESlGAoQSxrrJFPtWZ1g0yzksCOwsYe3opyR+BL+4H7Oxtst7ZJoP8
IoW5lZ2xGh0VvRjJ6I73I83C/YIAYio8jwOQMnb6JPAK2JV8DyTFbKnmPAw5L4oxcuSq+KdCboEC
0Ww7VNwi0xh0xu8FfI6Xeq/K2Ze/oSQjwWcpFdL1a3P5L4MVRnI0N43GHk65Jrd0Gr5IxxqzPttQ
exQAmKzeqDrlVRFlmgl0Bq2ILyXqOD3EuKPZVoyVonLCsJz85S1qfcTHY3GuT6LoZeX8iSJLuvJf
kpOgzKN+Dc5YcKUEM2+4oKTsQ/IMOtYinh+4JwmfwjWdvfs8cYMDymU/+/3Q4yh6hZuuVQjrolxv
85Q2BRnpPR2RXuBmlFkoMDBznSdISIAVQOUePkTlxWU+ji9yGJuGFqqTzjYICX8AK+etuKjmO94L
4j3TkRyhqBfnHpiCy+aQIJF/VEsZClqzabng+evxihyBjhNIIq6oDE+xy7+go/IfbNKxvi075zZw
Qn5T7AYFvjIGMwgevfe/3MW6BugqQukQwkOUJgArGMchLbxUR5BjT0Kbg7Y7zUIFO657/lgku6J4
wYMMHbMqQzD2SdamVRFsLWeH0gjQVm89lDzDjBXmVqpOxQLFto1bf6V4DLwVUktbc86abhwSimWu
7OUH9wLzFmdttVPHsYWyIYmIBLz079sKw86O3jIXxawEHprvgIAEQOFtKA3L5FZk+4fGkPbjqZxD
+4wfyRtVtcqhAyxIzcEZuzJ80TUD8ELS+BIdZw244VpT9igv1gk20Rfuan+0e6gpqzC99Ko1wazq
L1UdePPcbSSk85b8sYy7QGPucHkfGgIf7AXwbdvTfYuKItQG0c7/QsZAm0Ra8q2RbsQKWkAiZmdG
G3GMJL6e367Ok8GZkqdVVxM9D/m1GWAyp3gmMP1IytGarYN142qQbEhuln5ic9GC5u8tUBzj8FWY
8Alw5X5Bv+3pCqf/4L9P8i0ECq30s9LHr6d8XJIj6O8XXDA04KJeGLr1gqbntjDcljFY8qJromAA
QBAjjfRooYoAm7FD6Keyn4jIedFLMLioO/vkCbWBVcp+USZdxkMuU1W+zV3NAgVCeZVBZu5SR0t8
/Gwy+wGeDtJyZwuC4Bn5+Ll8ja4Y8yu4ZX1mrHPc3IhLn0UWSmgCO/MstZmhzHVhRYVrO8kR1nEv
8z934oJ78wfi+PEQ3PFj2uMbxK8zxZV9T7JhioQdwZNrwi8E6CDIT5vYBUr9mCn4FtjsRAEiM+CR
L85phjspbGhpSyvCgSUkmYqJf/elKD4dZX42TSA5Bxc3TiY2ofqiXJLPPilxtZ+bzbifnRnEKI73
TNQcnIySiDEFXpQNOyHPge69E+EpcP6I7OsnAT3lQKXMrB07tR6rIaQZCieCyckFnkx7pJeEEky0
/cV6AGD//iuh5A6zGqRlTwNEe4xJtPMDgyp5N9DrVG1+Dm0PqJl77ZIA6gn7WvEQRq7CsJWiNpYz
qwILtcUPx64hfa5MOO/Ig0T54duGn2NvfmO0Nt0gHhm/YQgd3aN3ozR7R7DoCpisXHWAF7v09RT6
IivrZdZurK0OkdOMOXThPSzJ319K1935vzdnUHEx0TFrszwH/q2nqhese1MH0ULaqB6GkHHn6tbV
IUFfhGpEDs2khvtO85kYQffMocGL1KjdlJyMbngoNxnDHDxaCK2pvXPdSVyr3VBLR1B3YCm7iWdx
zwJ3gTjMvFGhvbetpwWxd9wLP+gd+2EfL8y2Ws3+l4mEvRo7aOevFN3/uVozk2pwbKFL8M/tCz83
75a5+SwMBR9pHLvg0sj5IxlwcyfwVLafHbWX8cT3SzOxZ+1ex0gwLuMa40Tf6RcMaNXitqRscc6E
15NLpeJHnfNkpTxOY4up/trzOCzjeNkaD2wwkGKAdxs4Zf7WmP+J4e8rp2e8QlRMnyNKvHO297MQ
AGRwQpGvvbN+U8JA5o101D7P+5vJNcGet4y8L92t+tpTL9D8l1qqjaL0pMyMqa7siTlInsYHB6+Z
1joOMt1CRQjGWBeveGW9MSixQe9+wQW2PF8AC8mjD+yNkzh3nbUA2jyLsB8Jh/Ib8g34Hj/hGNuz
qEmO86xjdEwMmArSYok/9jC53soJJ3fpUkouKBd39fCq9oyafXNHXxypEBANG28UxlskAOiKzmLp
Co0Jalx0j271UoFxLnSxOSyPalO7WNp8weudT1wtI46OyTk7qfIphOAk+H9DlHPcMyRNp+bFzm84
xs1Bzq8EMidXB1qZ9Xel7qlm5ESFQqaBjH0TYBn5HtBCFlRDZucTsn/Lfv9b//d0UxDq4ip5D1+U
QDh38Hw+9cYDUyxg/FPkNgV0FOilx2qCEcIbMQKh/8D+fOTX/obgTxae7w03txdIyt1bHgeLcnMR
RtiVzmlEXvNbdpJU1Nb9WHD8jPJcmvusltKqC3vpnDVojFFgM407/Q9NzMw7WH5rzxYc99CxgMMU
O8bMvMyCXCPt+Smf0AI/qmRaR/atlN9VCJAulV16NGk5s5AziWK7skiyBE2t2zlxfwYdOibsJz02
aAa0jq0zeyBCQcCyx4P6yGGSkrvTqnTemo06d5fzVZiSFBPbvzSqww/MEcE9u17/3TjnW43SOBYA
yLam9j/v4fWCcvAEJVVV/1ZMh6HFE8QyMzxwjhR3A+zb1T+bq0yjeejAB7ghM8rt7zIZEJJjm5/W
oilkYuNarOiV4ycnEmvK8xKxQ8AbAEIawo0KOJnIKlGzDSBiij1jkLfYpb5ggZL1WG/N13p50/zk
0JpSawmb6AXP5A2v9ZXALGJxaNrSzoHrkUIYMbwKyzZOjpVTgjimQLDjrZAxRM9AYRplNcow+wlQ
tBiCkF0nNEmlQNpTMmR1VpHoy9U1VEgfc37MoM7vvF8aMfI5y2BEdfVyAA5OIrJe44F1MGBjn+oW
zpXXHFI0KWQRkJf8HRCY+wxhhAvYSQsIXCUC0u2XtUIGyXhtxtxXV7jpmJGufsB52uFz+JZiRhKk
Q8KQKioNF6ojU4d2KHZv56pqQ95cloroYZbW33OirzEdFLDOVd6byjC1znk3DdPUZZ3b4IHBVT9D
rDfV8jQijkQsBKph9A5SuCBvfKJiy/ziDcap4F+9Jgb80JkwQsqwDdMYdJGsCxRRmT8KwkOezZ3P
hy/OS+JCXMe96U7EqQtgE80Q4UBLSaRFPGZwrlfhsrK3Rq8Lsl1PG1KTj0hzD4+7LEQlMfh3eROo
TTjJcTDGnkLhqyrfvnBOoKouByPrIem854tIiyEPdfz2ipMEywrfRYRh6g2xg/H2KV8Jt8o7Gnaz
RXiRB9sVOzih+uH+RyT/F8QRx9YP1vJDS8q2sL7+fNkndzjHBzI+dKwMJmrxSKgXTkIO4IePh10k
yMfa2Kwkg46FC35f03CUreSTP6KQGgF0ptc3B++gxDCh1Dr24FS0QQ9Q+bEJuav4ejv+NBEPMADo
s+4sxnRuauCSW99MAFOYITWGM+1X7zUkKT3NJWhncWq9/QZN+LKXAJRWt8I6/5fDN99pmIlTd3uw
fYG9AEJwQ7QhaVTvcgpKf1hmElKjCQ/lAWTqUim/r91Z73ogdCGr09S5HIEe7gRqFxNV3y68PoZm
SOQZrKzADp/ZAKbRdlb4NUX8cDxB72TZkKEunyn375sQiXN+evFxTfdu+YalGykevmJGn1yN6QgN
uxSOP9eHx6tLxJFgK3D8iw9h8YNonPtuqIBSCIIF+hQ3trXtdJVzCcbLC1o2tMPydV3+dmNgfuA8
NZfbQ72/LD0hNwuG0NB0fi8xi113JeiUM1fVGaN3lsrZPyZPDcjURaXSefHufjNqWY0KGJYGUy14
jgZCrKDTuQ8QeNafyptvz+Lo/urM4JmDkhvqQf5HDX6c7Geg0mYNgAgjqOfyrg8u4wLi1F0sHpHM
dForRGYdgYaHW7SYOYuQwbn0lC2bYONHTnMpcQMq7PCkOYXGO1emJ0lpe1Nc7F6XruWYbvvqVk07
60Z9YbMmSJHmnKPfTsZBzDqEoPwrdD0W6H5kTdSbRkaqXPD8urKofeBZdmxeQVpSnqFJDEd599nt
p9nC1fKRe/7gsGEbn6wGhOdfoRTcDa41mwC6mPZG/gHxFmgNhyabaF6VftQSOIx9RLrzMgWZcner
FGBtG/dlGYM8hIc4G8Gowa06oJkbyPKKyEDjxUi2aD4xY5pB+S+Wps8W7CbYFG5kayGax7XPqzYO
7y1pzABHX2tdYU8zFyV8wsqFZSA+GN1gTYAmz12udMAh8FaqfLVCDFe750wr6hWTBaEzPrGPsHru
0XWwQZ46owYJ+GpvmksQRelo0jFwVBIp0VYQl4M7Wnld0gQENG+DQQAQ9jZOCV4dV1BLg24W8nFr
m8eQMIFiljODuhgrq12usnogRWHXCg3ZIq1aypnHKfSadLLJLwdigcKm4oOkx4VHAgqjIvFbd4v+
BtonqHRjUizhQQkaf2+M0V4QNfYX31nmdyPyNMeFEi2CBS7Ius1phmfJgRY2yTE23zGY870ElMNG
vVzcyYVyVenRat8QGhquQF+Q4w8MGZp2zZcyiLSrOvO/EWHmqi6dJx2MCPD+RPdFD8/1T0OTNlWU
vtZVpfiQYxBsWzr0b4FQBmAHSzEhTXtGjoBWBI2rkxaGjBD1CmNEzihWLEeY4W12xpblg3nowxfq
Xbrj8nvhDusiTS9snfHPNB/f/v7X+CiKkkRYc4voa4eHpNumgXQQPxaqg8wwSOPN7S+qKdcjbvvK
dBDLGUZXvOOKEVpfXfIeF5b/7R/3E+i4kezJ1PFN9zLz/8D1qX2HNk3p8Qxm090ENfm7k4wnM+kw
B6BBUSsmbQQaw0nFdmBu9DKW1jzrQCeD33IDD0Jt6Zteo/rL8DZcrmLTu24jI13fMfUpnsM8o7hd
KoKXsmLRTjvLLyXawhv/mtp8rUD38fJqZt1td7nPW66iyBkiVhZKYvnerz2zRp7GBkhFBmZlLPSx
GIcX8tdnnfc1NsgZzU2U2r4plwoL2SJxkr1gReprEacizX7mmYlRUcfKdfdW9zvJqbG2s0NJ1ygh
pqIweOuouhsSY+7bhRisNzgwGhwQOJp941gTKNE7cnccX7VwEVfuoMIK79ac6zrCSW+ST7E2oGuT
vyNABA2jSkTxIR01zunPvw6w2Dx9No3xUT3hoCf1jYQNkMxt3GJWKUkPvkY8+ppfgSHCQJlEs2C9
ItI/7/i74tf6eoVFVbEEQ09+2Z8xrJ3J5Kik1Uqw8ZlnbFoKnXYaT/0Llxdb3M4PcOK6NGeq+jn1
NMxLzA3RCn4enN3lJBmPDcMd0nVt1MrlGR4deUqqIO6v5RALiyphEWYZQe7ySi18cqkRKbAbKVoh
Hk99+BGSsCUno/loKz1V4UXlVX8P8UTqpk3kmeLbkSfJMlyBKVCg+qDrMn2eGG1uTZLP+yvYmDBD
chA9jhKmTk8GVIkLc/c3V7GTaThnA7dfEb+JXjbYmY4IumkOPLXgwowFSDxhT8jvo8USMxRbJPqW
8RvzusfuqAoKbjjR2ckHy4O8oOxaE82IQ9da49mTAJMW5yV7SfBkXGXnDhHZX7E7uPfVRhb2yChx
VHtHTaonMeqs+7J96PqI92KGXP8Y6VqX3g8CxwYUMw+9VEBbB3DXBflFTE4ms+xf/6ngVDF61JuR
Ee4FKkEdW/8hG1ZyJqE8kv6NIPPQ5KEWXms1LTAIIDqJBPN+1AgL6IghZ+Lv6gV1yeEW70wjUFjk
dCeNuWA6jItw601HJo//ALVZoBvdieCm6kWk4Qy1LfV+qJEJxUUis2F9Jfd3pZsQ4rEHhJA0Q/b3
UK3yEcCkvyIwkcBvQ8TuQed5N8EGuzpdSWF7hO6wMJrCrTrSMSMhmrL417iLvX2RRiZOzD6olIvc
DHIx3ftsmfc9FBQPyzgpwnqAXDQgkfz3jfIUlurASWM7uRNzlfYOldqKfBYF3+YU8q12VqMdx4wm
EfvxwicLbetYhAQHLs0nbl0zPesnaHmhW3dMfA5nr8Eu8dXvJdikR8MLv0ETywYFagXM0PhTRFxr
xKTGj4wpXcnAv/+UF18Agg0Ol4gIRm2FBTrO3hGEwedpUTqLwKikQFBYO9tHYMu6n38f6+Lgvc0R
22yxdBYUwpNepGKB9aRVWNgWwcCDJQSk+/wwp+xsZrndZmlYyJRTpCHA53lRYAmTKl5bQrrBjCAw
8AZZ6QgS4xfZYJmdhdaOPPqt2iR0eJ+qJfqvwYGmEZCAQEaDKTV1AjaxHkU6iA2CwN0haLcwJF8t
CkoToWZCAiJPGnd9r0KU/cSqtSCDXDd00olh02U8xWms7EaEjw897cEEpX4OulsoaTzWnQkHgka9
erCQDNbzBFTzrg3MGQAVr8QIWEOvBa55RA9GzoQH1BkQm+I3yLE/06jEjwdm4r8HobKycY4KkSOf
pxzZVmD608SxlVLdkjkyOfxrVq/3yiWtZ+o+43Jqd4UmOlUIVxhOR1tKb8pCIMAqS/dWaZzzi8aV
Neb/65cd7zShoLw2zYOlHpwayRPDXGsyS4LWYiSl5vh4nT0z7ofllgGV7PIycc74T/XdmrTGvaQL
aK31LJzB4TABibMITpUZxSAoLgbp2rqsqr2MZWa/V5Hy/4RGpkqcv82258fOUmqcCebF/3iivCBb
dt5vd5zS4shP9+ECzt00xgUYXDS5LceqbK2DvUl4M1Beb24fImANPXDEke5VG8s0XJGNYN29txgM
vdUctxRQUS2E5zyzkf1IvZe2tpM8m4MzNRVOUpYzKU751bq5wYqikTXu0NprwisgIXDhoUKuIJq+
T2IFpqm6aOgVk9OUnPDlbf1keW+ajVC9iJfeBvjOhJrWMP2+/MiZTPSlE4Me+wBc+aksqu3NBQwF
nKmCwhYulGOg9Aq2Uvkk1diaGD13JLjjrVuz8LtIUpEsZoP7kAycw8+f67jMdWS69x4AnQCiW7+Q
+tbiiCDuZRDlbYBhfXu55vPOCBZ5EuB6qFgzq+/mqy9M9cD3SGDkkjQZjmtbffkrbICfqsVN6ykh
MZyYEQ8drUG9NYwiGGEP25OG8dB+fBlgrBwk9tLTTTzqD2bh0aM3gyegUwJ9aC45DmuQSME2ZhaP
tbAB6VdQoTQ8Iw1PUFCN4LeSsdiImNl4dWEgNzkz2eoh4D6YrImJmIfItNKT61RAWhMv4nq7D6Hv
LCSZJm2SmyL6skGXpTWIQpwFZvuauXWKKv+m2RL7nv9BY8juSQHJ0QZGriBZdVw5/rsQDqHeoAHQ
PiNi2zMTnWyt4HBPEXVO5oF2XXo9dvv1dG0IChQhFPAGHvx4T3oIbDyFYr8hsOdoVOaeqe3zZmZ7
/D4/q8XGT00OM3GfWJkVOk++2RI4uTROeGwU8o9fe+1zQWGVWspL5tRjJ+YZPCOjCzKqj1jI7gbl
OWfvw4b5zHVvv6bOiUnbLj/3VJhY8f+oDmw+w8xxtAFm+eAgvaZsXLriaD7HlxQhdPUKxOojZn63
TcnACdOdj6nbrYWlHVEDbKTr1hUE7IzhwrqgXGp1ICYh+ClATgQB8VyCSAwj+k6URcD1IqJr5ox3
CZt+kgLLOwe2XAbxeI7ofotrxNEMr1MC5mpKBjDJ3Ovx4ZEV9VHdjOnZpq+ezaB+Sujjd4DJrwba
ApEbThKdE+HkM7vVgVAB6wAWk5LlkM71I2Qwki275pRorKtRTEeq1XY//ZW/VG2Hgbn6Dwj4g0Ms
rE1QMrhmuCbUZSEaZkrPiqjlsGIBuWNEHHE9lyA7DecZZe2XPdryOTBKBNQ+hVO8zwuoEcZG+lHy
zznww6knJg0/2u959WEr82LIXYnUBnM5GE2G1j4ePKj9ckVDkYh051L2XbiG5bpFl4skQNTmidIj
D98729GAhOh9Vl/ZJYdyo09cxNmxe8yl8FWQX33jktOyC89PDxcOzQGS02/ATSsGidw/WkP8nOKG
cp0OjE5MCKqUhJDK3qhQtujx4W6N/qPKuZzcADh1cihbhNavYE9KkycDbqSuOQmZleA4b9bOZi+y
nCoTQXIDJikOyezoDMTqrB7y3D9g7xPrz/+zasDcmUc42NDBnoqGdBY3miFZOA2ltwWTsBv1AQgN
S9idHYRPzotnkViBEApBv5Fk35jrWN2pOfRZNW5fwWYo08gr/Pog30j6agSwcrgVzbHbF6P7MTLb
oqY02cMWK2D37Ra9AX6miUL7z4SEtgrAq3f06gHa36zizb8BE6cQyE58iQPHWXPA9XZLmso0BkxK
mpEC71DmC9uYozYPOyENBCgT9S8psNpBQEat5wHVc5t0UuU2J0Gea5a1dag6U7JkvMF3ZM5T+ie4
4wNTJAwQ6LZtoqbbVIe+PHZa9dVgKr5pwbVCItLOKrO6d9MiPcqbRE+3IgaCbNyc0+l72Gz4QWdv
EfGgLvcUSA4WuvJZ97kC8fjdk4z5iNSzotUluQpL4/ujUKE7umNxzOc6erre3iWuX2eyzpbydhxo
0bfY6M5kyIenbkh+9Lp8ipA0e8+SsmSmijq+KTfluC+lQWPJlqruTwMfpVT+yiiiqQ1JcJAgpIGe
trjsqaRlAZg/1idipm9DoIK9GM3DeBKVCOyxR62j/rwhlc+6B+JV58fnKlse1ihiblsSyc9edggo
ucpzxz6eh2/PKop2tjqpQMOQX+E1Miwi8eLxU5r1bBFGqwfcPt2N/bQKV8G6ErKLbeY1He+juXPf
XlmXO/P7qdqU9B7DoMtDg1MbE47qrhdFMq9jhivRpFj6SZ0UAXWV4B+j4fnU6Zk/uNnLYo/oAhLe
UqCbrmQYxJ5HjJFrFLCq/jmKs7BaWh9O5HhFcKLpmMpCcR7qRMt/lzac+NCVhRkBntwQsQs2LjM1
3R28+BFMJccb34+iCD1hRvFp4RzPWWG5ANKjAxt+BHmc4M6MHXBGyGFKuCNGTkPUkXSdbO3DcoOj
xIgGVTf1DFL+BxcMfMhHXq7WIyVjGeUYBu2DsbGOatJwdbGdusjf51n+0QmgDe44z5QnbRxQvpd+
dtEw5sa1TIY0MLYkArGlrPKv+nyGDFcRp6VMoqn6plt2Dq3Ir9tlXQRLefDJeYQJp9+3bJbRR4wx
2aCCAJzUaDzkqBM2CLTLiSEv+v3vqG0+bNRszlRd5Phbet9hNIvMtMnytXVw1HR8bxbHabbl8Ph9
Rm6U24vkqsdRjJXVTs+Vf0IpFe9ZFcdvcnwC/VnfIde52bgSV+go22MSR9taoNS4br7Y2a2HZ3qr
k3tbO8zzPjixLYFUnPo+ifpK+rKE2BFcVDu8NEylMjWHg78L1r7QBj0GVyExBw8xjjXooi1z2a8S
T7FDSW4hu/zBGCp/fJqLVAoiykyy6gpD4BreoBzQsmDzz2pvVoUkwWVVcX9u4D0ydPlPoRpVxzwV
YCz8ogpbS11rO5/9Fdrf+OveiiyFJ1ZpSeIz1I9RbZFdeEO1HAHx+O4Qbt+CK52fWPXWFgw8gul4
G0gF5ktQuWobziW6FoP1zFKN03LDqCYf/mygEZjJ6xpy1cUBfwVU/VdnF1CcT5LwG31FbWxqUc7e
ubBKvfb+HsPR2cH06as16VFKCpMbpFzKowQKNUtJWu5d1Zoi38zc8wDqFi6F2OI3rqhHdVZFk1VQ
ptp5ojDF4kmi7ctYrKQHyOD+ONSKZc3j0QUnPMJ69hn8ZF/g/fCgZcKXb7m7S315Q6znDFGWHaXa
Z5dbEU7JGSGhK1H8q7KGRJrmIoTApc3385OTUfAS/uY+88z+jOfjN3Xyry8sR1jlPAD/F7rO03xT
slU9nWc16Ei/MNMKjkrN/aeErPtepteOzgasrxQQq8g5A1XKQBwvQkAwLHohWlBaBDX4fHkXOWau
7lJYD/3Bh7XnceSzNiAP81BKI5ov27VWjylJCPgM94npUHc/2ieTKiAgYDfMFpxrUt4jHxxUc/Du
+lKYo+qoVWYcfQD3RIWCOKst1WNetrGSXchBfx9DM3qaFOVpq+0643VArE+rZiBcwDUiALiHL8nQ
U6yUT1B4cp2YdkrB+YSMt1WorvRJ7AIZ3slnCVALUz+uEZ5wclLBDKemsnVoohAA3fhPE+Nlq5nD
79a6ZJRrAgUrKBSjGstDBTntUycMMZEExhcRSVlDAy2mUpAvQ4mE4iqZPm2Hs7acVEe7Azbpy/Bd
wfQxmlvKJHotiojeDyxWi5Lhs1P28Rq2B4R0zimU7HRiMxe008NecZfKC9htwUKQVUyXswZ/feU1
qYCi7ebxaTfp2LcgV9qF+fg0vopUrCXeGIUXIREyjQ4ZrdQWJcGFBxeip/nwpv3AWlGYQhbvqtYn
pvi2lJmdju7cL0Qhx8agvxFKcaQ3DbH3JKqBVEqBQtUe5MDZ/FhdxOHS2ZqssQNnFu8Al0mR/sQt
Beg4AZiAnCiHE5jOCyNLS1W8UABvAl2TKPaxcYs3YPS15cJzUMTsh68k6q8Ugkx77tN8KWer8uU2
9iaCzIJh7w/2XIg0KH9XIrzmPZtzwC4Vf3liIsw0VBngmkZ7FH6npIumrL/PqtkYZFgJgnYlmz7i
eMl/GkcKsi8IYUDTJRYmkhrIE8oObaLoYs+ANMqrllUjV/oGj2RA9i0G2EJT83xBZqHmWKvrp6R4
0AN3cKOSV+lGqm9SoWOY7Q2V7ScOlzm3KNl9A7IGo6XwIElskxxYXyTR0kG7fiR+/viXd8t4qDWd
34/FYVP5ndpT1i+nZYg3P6KEJtxppHtapK0PGrs3ZilOEiXO7HTPktjN3voaXLZngjrdnjZCnm//
csK3BPzufDpCWxUrH12Icih67JDu4eCRogfV9i3Bp28D8BJCFVFKkQHNXvl3+zjDWFmDMUaOfrTN
6RQmgsF4t9HhKqwKvYEhCblYBmXgwhm2ZVfQTJ17TXnecN58lVYm7aCZkolgs4ItxRxLwOSIrlm1
wdJAOrEM3O7diwxgVlpd5yzdYENiBc2TsiKO8Ihx9KeNmqHfia0LZOAS+wuu1/s3TgaEPhQlRkel
8HalT6JVqgYbH3VlB5zdAwKV11H93GN1kMAAMAhRyqpOTzxMfFjCO4SHwJy2tOEJ4gLYcnFfma8m
EhazM8zYhHQBiHLMNF4U4QMUaorJhFVTumMmkRPI3HZpUB9yB3uvzttZNtkXWQRdJAJupohUbN+G
xmUlZRGBSh1hYt4OKT7EepoAyBSXHxwZ3RjqJND3eeH7l+AHek5UWYm6dhaUk7rbmqLBzh4fRbNi
no5Wrlx1pFajE8jVx43zS3OPD/oFtfO+zwPw0JwAry6hZcswIQDdKyeR0Pjks4eyyMSgNl3rHpCK
bv1P9rupoDGfYoE5mm+nvOjc8MFVjQ5shEZfQSKcP889+TwTQF7L4DKeWMHA0AHFAn+34vvKZadP
lJ1jK3W9fyhQil5CPhCQD7tYRLktge1ZZL/4EepxUul4gPl+EDTWzzfUsSxPShs3m9C5GVVb/BkJ
hov0bF1BeAgjmF7UnQ8DP7WE8d0RFZxoXvyjyJCtmHwwmDL7tGKsCkVPO3oQ104LERZjVyM91SjV
AtuknQY4hTI1CmfVVYxvw7GIdqxGfydfjUAt8E3s7r7lJl5jkLzGfe5m4YgwpiqyHJrM/6txjACg
xBA3tEf2zXo/3TfStsRWk3UJbMqan2LN5aFXbZMoyYHyc5pPpmR0Gq4r60ks6HdGLkWr/z4IA4zQ
kUNpon5oB6j8sUKa7xly8xSZRc+l+nlLnMLJYKLrHr6cKw5KN1a4vcR9hxXbMWVvzRP4451m2rXd
do7iKvz8Gd5VvxcIjhAjq9Ne+jDBE86YLyxXIACIjsJ+FuL5BkomxESGKyGORKpTqg4+zO2LRE12
aoatALmKeyFrBXCj8RnDRHYS+I2YxQzqgoev0YvFMABVc/fqBtb8/nImu2qYp4wopRtmcHn4e0FX
b4KF+ElhTIXtsIfF56gJWD10O8EM95zhRR97Zatm+q3qE7IpM3yuyG8ND7OBjzemXusjeEn5ZVNs
8VhRVLZOM/mEL1n5v5dth2RlQHR2S2MIwF12o86NUejtJi8fHZK957EJWgAlq9NAOihEv461Bcu2
enPUVKzSBEa23lHq1Xv8XYhsQLbFN5W37ixuqGrr/od9cRm5lwo4s1+EbCEkU6c7Obu585D6gdps
mcbGJ7u7SF8mraFoZAcriAEnVQnJAlgBfz3KMYulRgTzU/QMLQh0aVYJHaHPddxXA7sRKAFxC11n
V7mm4WPA/juIMnX/hkoCxhgoks7f6PQdQdeeXpH/S7F4EmRIJMmkQeK0TNsY2tFjKzUT+CwDxE3N
AYOhSXZbVUrZQBXfLGkXBMjPrigMSlCA1L4581dTVR4Iau5jD6CJUVTUSn9pnS0NkJfEve12elAJ
KDbTtcOW6niHyy9324jef3vyXuQA4mNV3jW8XLYb/KpN74WMpWFWWKPAxeCbE0OZ67cXZq7KGxF0
mkj2wUSinp4yEgxWE8akIK9kdCC524mrJyoDe3awpTe7R2lL3IcGXJNzWTRT0hfXqHcCfhdrGhTt
ctXH4J3RRWM++PBTMJWt8FiBeXJv+bmM8YNKs5TljMdBuN69gLRPkqG0DddtJGcaKKjNbc+oqcOk
M21tmJuJ1nHJLJztUw7xmicJyoQxtFBg4ZtfzLikbBeV2uasR0eyO236KfaYzRzTWlRN3o7T1cjB
P/tuxz9I9FM6sOsI4JkFFxNDCbSHqSDhdjcWgfFvzXRgSGBz8Vuy1UVJjSRz+ISEbXRsjABElIxO
hvrUseYUS+d/0tkT4WonTz82+Kfvdm9FGGo6W9fQ8G6MQiOJvSKIpGuWnZYl5o7hbfaXtPC3woL/
JPScD7fjuxRb/opmm/SjYcKghe8QEvyA6pvaNQQ7wdag0+PcK2uWuxls++UZzSCJNYRTUYhgqCc2
/XM+4gpgFxQJw+AKBlryujrTm6jKvfaTHINMlJUJoRU1S0mI6+1LgS6c2+3tudpBiKa9gw9SMuvc
HFdHaXlj+PpYWcryY5634XTCkcAiX0eME5QEIBMLMxCh25WlcUoWPLgFPOH2HtCK+XfVjKa2Utk5
w4Aae77uJXjkHGaS/+YbZQM0r12CMmIZP7xNNxaBZOcKR3eYfl76rMZM6SCSRSKAnxpKERNWHFZR
lYHiTdM66pvfCUEgVrTI7A6ykNqxf3sIAqUnVHlSMKfJer6aASaBPvlN+Kc0Ggeg4av/VuSFyfzz
ptKC3WYEJ3Hvs4/SFCT/wltZwKNOGMGFg+/sBqSckx0TRB3KOvgKB5uiSPNgn8JVvNWJJGS7OnDz
FbzqRXVMR2mleNcu7m29gl7hO3RUqUUZ6beZHEfc70LFy+692OuTNS7eqkZknOrJkMJtrmHLoIh/
c/vnnGCVdLB0lJdnZ96bawecDnaHG2HrBGgZPdXDTVf4pNk3RVRxE4QXc3qePNKN4bMDfvPkJb/b
iNfI5IQZ7hXMnl0ciqGV6M1BmU3w5WTh7jlxqglXDXI1Dtltu0C7js74Xbd8xyDs/z+TqgA41ZJi
RwjvYQLRc7Q4RWGkW5F26/SNJKKWacdewPSh/GPv6Vmscu5nuGrsJsmNR4V1oY8UzCoqpM1PYrik
Hyg9KvQaiJxKPiYUHC+WGJwRTh0M7zWNGagxKUIgyocNPs/Mb6D15q59tN2kz38PzyNKF44eA0Y8
kNEp+hKDqIYgGu54B6pwmRpqfiZTpCYv3SX2J8sCnwqp25jW+3ukbFl58MIBYXIYf1jHBapqP6r1
/XAr7Hlsp9sklw/2U+/0qjyw5C67F7/44RgbwIfO2c3b++FqeD1DBX96eRLywODlipCXO03M7yaM
1m8XrqrqoUhSd8XFRU+0P1hpOAIEvXTbvm/PxAHwcNB3HPVltYmNG7SyVbqTtE7IlI1KcNDpCgsR
GZUMxN7WEX53ewf0P2yr0dGA+8661b82Mc/0ePVDW/oJhMZeNRby7SpRQnpqorb80s0cLVGyysre
/9oDcFZauXRiLWJsvMwuxo83FLw52pDs9/A4iiNzJqA6FtvNWacOTbaX6MIWpdc3kCUxb/bxB7B/
VUqxV/B3GLQ9IUiiYBGdXrIeOCvIda33hDHbCMfk7WxyHlywnayh580fiBk8FjpivloinMeG90yR
Ovc6rCHdQACASQ47OliY0VcoZ7eDT5ItLOixHvbAdI1URM8dBC9pIJ0eGqyyjS7CZQyMqlGfJDbl
u9/JXG/U6n1hgkeYovczmuFPLEtLwAOD8ucFMLTaxHnpszdUQEFT9vbtOoV55ka+r0UIkLYiU7Gn
C/QUcbqg8grX0NQLjYrtPqoAjJgX+MdKEKf2lvaFIfhV6CAqbqLcf7a55eBhHN/8XDCO/8P02tkg
+xDRqnmuDylkkG6o9Th90PzhoiRWZssO0DyXcNpnIdo73ZligFgt7yRN1GDoxRZIL922Vlb+uOCA
qsVlRcU3dshCeSQ1S0XFoBYiqspJKPtANUHrlkTQRayj/YvBMAJJclNTB9df/3Nceu9o5glEhsUL
rH8HDKRW8YxkEhetd9xu58cOxqH4f8LiYuSDiVKlmWtJ/zC9HA0itvU6RIt0H7bo04NQ1Co2Yb9i
NRg3xVFo9wMBb6D6u28IfyxAjiAf77VUFwnb0qHWu/1HUaCVLGwM4+HQZx+EYlX3M+/2V42jMPqk
45ls99/dvH6Cy69UoLxxX+D942QqbnHAdpHrzXNUkiQz/sodemsUJVIBlTV5I7xZP6s/5emcmBQR
Rq5Hr2VHpKqzvLkRwcva4MomSVnyI6ON/FuVqNxOySvIIWB9s4mTHa796Bm2zt9jHTtVR+x1F+zb
taaXx+J/rzv8CqDz1VAs9cVnhzfWXlmrm+v7sSVzReTZY+QfVFlyGamn9BsvrJ3GmfB36U4JETYe
UbKEqSvlGRsFm7b5yNzi2GUwJPfJ3AiUn0PDPwJshx6NNrNpARWr4uLmtM4rOYAqV6UQzdNhd0yB
MPj8uf/pCUcCnALO3f2pinsqqwL4qGI7bXjJ63E5LVqeyShu/daH624/+NfivxIwsqYn/6osLcTr
+HCWI+I9t1wfiT8251O3o/dzCsJBI3fu2PUI6QjYKgVm5Z0X8kk2rxuLAClVxLXiIbtVtO5PDhhz
rmmTi0UntPH8l15ZknIt39iXuwaeLTFsWjQy5Uy00SNlDdk2Fzk9CQ3AC2CA4yNXxYekM3ciOl0i
80np990Rxv7yf3Y+0zeRuhohUqsIru03yT/RTEOtzsJx3Zeuk+xAedwDa8O6ABV8Oi7QYGKwDeCF
zGNb+s0Qngq22dcrFd3NE0VuFGWDwSlLikxd4Afje18kZLMOjne7seg0Ryp78j7U5+HpUtZ4bsne
SJ05XVysi+83hk3YxzUhWOfP8qEIWLnETNso017LPLJjCwGHGp6grsASPd61M9YJVlMMBgKyzMI1
dPbvQDVlj6uTp9Csd35Ivqrg/peIrmbjbf27ousYxlH52kKFMfL6KDi6MbGAaFT07oB8FfvUbvAS
ayR0tk0Pp2c61e+Hwm44gwBgRePiKE7u5hZY1aIaJVc3vOhzCVqXK1ojGyziYdSEdmR8cjGskwM1
mRnB4FMih7jFLqHqe90rF+9zkNjBT8PM80XLw1o0mIxaN8uI0d/h/UbweDQpXWeEiRMTYgRfUMk6
VZvcC+seZIPSovca44wHbH4L/ZnggyZR/34A5ToWcOvDgSpJ6oxn4c2/K9t48Xc1CJIWbir1Es4y
7anUJj8HRTrzsklP+0xe1wHx642QCH4HVlc2rDDirpVET7Ndm2DF+jeOBJ6Kl0GiqyT64LuBcUiJ
FtptmdGY/jHAbnY1UISvS6GkytQXey1Do/W9OMgCOw17Fuq8PE5pR+FSxGfFcX+FqrjgwrOvfiIV
hcBhiQrGqSMgHTgEgTgoQuP7biraYSLZ1bxNfDFsK9NWdKki63qDg30wnJB6j5xA8fYdqJWviDEA
1ZNZisgpwYlC7PsNvbxZBuHEMYVIno8BdhHv/w/3CsGkC79PrA4tIK3UPvhUibbUfKwbpWuwulnI
UfGqc6U6S8CM+W8w34td3GWwsEoUX0+0FwJz5UfJStPkm9X5TFK8cWs3Sci79NddZR2aNsvXusND
HVfEx4MfLoO8cGAhULUmjFyR5UuRti1uO9aYSKxzNoB/r7XYYKVB6eXRiXMwYqgX35XIxW96UE3F
vTEr5stz99RFFI6FS0rFmNyrVrXJkn0A/NsymN0TRz50KYu9IPxsafl5SJfmiD3hTbld2SjWNlQS
2byS6rh/5gBOI8pB7fW/RAruuRIQx/eZBnOZWjhydEJTTsgyZz71dG+0cQ79ZnW2/gCg1r4nKpRE
t1rF/XYLaweMwaZqU7czbApQxGQ5AY9z+3iRNF80Gj1t562dv9D+mH650gabMyVt/DofiJpB2Df6
p/JIGpC94m4SFDX3WvhkB9InE4UonY8qt13Ib2wnCjIxeb0+mOvGMH/QQbIkrE7moTqVAG0ozqVV
+RXb5a5aMppZdrLoxrK7q+KKRUcjlR8FgtB2YYbtr0uAbdCFzZK/ldG0cerU5PdXBapcgYxHioEi
d/TZfo3pGxjWJr7BGiHz6EusvS7kdTy77xdRIi0cUKzQjXq+Uj+xrhqfF1R4DWBDpYP81LlalNNy
Nm+s/eR3+ReLUCYl65c9Td1GMUlBErauv9V+D7bfR5mbAeSeDQv6avtAy1jOijpctHeU4uZktZLS
X+s0oHOtMeXKIG8acoU7VumSxR/Z9JLDOVZlkhdUhrrv0i+uJ8AlP2aRJd1hM2pe7/9xXSQzb6Us
aqqHDc2aqXPUE8CGC72Iqo+U4vpCDNt0Vw0n0d/AZyHcWSQi8z6oBjmP6EHcTLXPwzOXmyK5SAJK
3pfdPWEAwTxwm/GAKLRsHzbye+i4+NpNjvLtoXynwpuyPN7LtU0RhOI0jj/OlNHfWxe5WXhiwULs
DXrWIrb7BntlJkhEBRl3IEkLzrC3Im/alXPrQE23W24Y0IxT53lGwuGztRGp4AlyUaphRIrq3Fsx
5nFmvm7ZJ8uag0GWcvBm1H/EZvMHjVAuNn4WKKmjGwU/ftXAo0K0f4DIVJ0h3AWlTP5z5V5XNqY4
QuRzRI5LGsJ1netmTPypkyDQ3PfWmlGTEMCfj5xPmqOMHVzb57taOqJfPUpUBRe3XbvXHFMpg47N
KSVRJWFXUfJ0esfyPajn7dvAOhVxjB0J8HMHWRMfZ1O7ql7EQB+lZPuY1ed7Zdy8nKfq40TmAAH9
/2OcO8ijACeqabKLf7HV4olsiVig4oCjQKUbn/slKUhQcitB4/gecnT/0zfcJN1ex1mJ/MlBShHQ
VSEvAvxZkSoOty1X6G/O2DYpmrUw8nDWepc9GSKVLVNzeYdK74SsxlM1gozBFNJedap94XuDajN6
vKSs6Q4DJl1LEDIIR38tVb7FXG0EPuqhtvgNZM376rNW2bupSs6dp9BDx2cVge4LaAtCxjOJiHgt
v6JhXm58zb+l4zqLnLgexlWr7dq3y3t3DTwW4g4F2Obn0tYI4z1vlGKAKkp3V2L2cfRffotao/fb
EAKG55s8elHcEQqLwYzA+YAZ0GwButZOWkilBWhDwxL8cOw1YbPbrs7aVNayoi9E18dnXQ29n/9e
g0QryoRuManSoRraSd502Je4sYVxw+bkBvzrgWl9snaSrzo4qJ5uPWpQVMxb0tk6Frxr6qDw56Rh
A6EJGXYDOWSX94eIgvoTgcTnUE56TZB82LR1A/p0qRnqTv6PEABKQgWwQnprHhrIUszct/6C1umD
tLgBviA9O7Anv/YQ91fIkzrKZOWDf6goECcrZv3DrRCcWp+TknmhLfZXTlT8m46/EOGNoQ8fU+XI
qleEwNXUKmIbK87+qizHw/GwwJ4rMLtenS2yEHkUgEpExr1N5n12i1PLkvcsz2iHD/WuLGqcfRzq
AddAOD44rhmLAk2ZRY9sBYD+x/vD4PdFcBD9Q2SBpFqVxk5gcODfAhsvfNjVJWhJ0PNu5FDsWfZW
7vmV1DbzN1dvaxHaCweOHbq54OSEHc6mso/I9aXOLtH3f5SZQGx4P7dVRzEcQZ6E7vOl6Woab7Pd
5OOLJPBMFRf7e9m4VdeX+O+jQgMwSs2mvsgNWFS2QZ4YgsGdFR9K4coH4V27pKhcaLF4dxDxFt1M
XTg8SuSHLonWI/DnbkY5AVyBbLMMX+DyGALcHZvafSL4/yt/IUa3tUu1yXvg25axiAmMQYo/+/Tm
ivEX64FUiAWL/ClL86R9pm/5t313USAF2tNauY8xYrwQsJnYcxY1BJdXtSaR6olZXTAdSMsnbP59
IjXdySYurlp15ygmqIICP+T+4yY5DAbJqB3bWNZAXTy3faTy7QQSSL6HCQ+sVk5FI6FsEicG3Nsb
VLqOQPVmd/rOinTHdqO92b3oOlsLTq73o23WKTuRQRZQqzYrzUQ+EtQ4Q9bd3HQVlL1zOFRmbokk
AmINTxplt5NYp83w0mqdy38euaGguB1aLCR1pqLNoOATY41ID3eFJwaxsIYiBxAjOB4tlK8ACf9n
gofldv+goXecFiT+uw/w7dnFdT6xzGN3pYTodJcyln4DaibROT6efKno+n04YGKA+lOLvsy7Fiqo
WWkf48nwdUZ1w/+BOXJTzRBeyad82huzThi7jSt9hnNa5LPPu1tvRsksyzXLrpGXDF7Zluek70RE
hI2s+TY7EDS/XiBGwEt7Bc/4lZCtbxLDQs0TsQ8GKoZI9tj5N512UgS35iLADLbxM2F0fzySHk1B
EeKniivYgG2GOGTECHBGBa9oTxTAriOWQ6wMNw0MT8y7r1xeXz2SCPKGeKgKLjfN434AjhzEz9sU
l2twWsIUF3RsawUol07KMRhddUHeiSnJSo0TYue4oSpOyo161C7GXeP1y7NkU+r0hjwBDA+EXF0Y
Na7NA0GHyNQVxx+z8EFG5GJrdStpbrpUHA4o8BUhe7YWQhTV0jwF8Q3V0T04UCrdkEvEJbEudU7o
fFM8It8avOxaZYWpZDdf/9XiXzxJuylxcxNiaIWlSRqtKrP0fPKn6XkFIHbREWj3yPgjS1dvbktb
hrD1aK5LPSM9DsJcUymL8mL9YW0C3YzuJy3lae0D2S/yHIsDC394ik+hillazRPHKBU1nCpQUI0q
RHnHJtW1XuYPUeHhLUMNmBT+Lcm3Hwkpt03HgwBKMqe+TuRtKYnwGUiiaiHFPv1pf1/Xl9p8xWex
frKE8R2vcRrueT26lXY2ovg9o2X535KyNhRRC+QwL3POoUl/uDsKAtVhLtB+p9I9+04BdaDJW89q
piKcKYfvSGHUFGSbDB3FZQI3TQL+EYEi5GfOUO8ATonRD634eUyWQorcE/nRNRhSRhaHZ3Vzgh8K
QcM8Ui/EF2P/bgA+KeiZjyjg85mgOZ0yNVilTunxYIRxp5bq74bHfQHLt9qq9awfOPZF6cQqpGz3
HAKCQoOLUGn+0HzYlHivAyHawnC2yNBTg0WcDr8iPK9V7xG9+xC3cnRYX+5mcURCjO2ItPfsbliU
t7OMbX/FE+IFc36atP8u2BBcw86nSQox0ZwUBYgUTBNVlh9KsAnz3XvxLR5kDIx8vTKHE3jTM1hK
YQSr3jWRjczjd6693iuCym/9dcZw+rAF/7funzTGy9JaLGu02KCgsbMttYg48+dfragWTUheGHhy
KQmngmSwSTM6OXUVCXUWi7+6McNP1cO1jnPVZbvw7STq7UZjH6gYzdhF7Mx9dQRT5cwH+qoAh7bR
TJ2q6KyAVjhJtLy7fXMrRSysQqxyflJRe//wRfhxXBPNgxx9Acl5sqAH1vuCXcfXUgJQgn+i0HS8
tcxZ/29DXcmzQ0U+xsYZxAY48sPQsJNPG7vEqGqWRfyT2i1/8uijzPwfbHLUyjsvYDyHjv3/rd5G
D0Y7HSzMm7b6aKq4ImlyMKBKqGZ9qnlM6mrmIJwEgVIP0t/L2fGFFM5kV5fZJcF0RD40FT8irBnB
kuJiFqDCCYxXtybC/N+UwmdetH12MhXJyzH+nHKhrSheZqtSkynSR5Q83UkLEVZCUm6HFixvQhTG
LyNj5HrqXuf4KKeVCEUmdRnNMFG4QvYPIHumqjRzzHki29qOO+hwtQAxwqzqwc81VeZ7HjZ8nWRQ
5Lg9v+dF4s8VArKNMOsbw+j8arxQNQ52D5lIZXmEwlFtUgDnDW/g2qoaIZ/CFcfp8YApeD4OtEUY
3dSEz7urQDKKVdwcGMQ665xj5sd7O+dPrEf5+9leb659j7SIaq6ZD3H3R7rnmB+54JiBIwiE67UB
l0IC9QJD35XIoAdt5QWNGHk9azUQagj7ZnmMq5bITqWkOcgLjZC+W/xZeWvLuo38gerxVUheu4Yw
3k0AEJrg8OsbN9FmbKhfqkvUYkTxd1IRY3vfyjI1zNiE2qXJ8t0dZAty8fggmlgy/bpJ9dnjn7zX
QlUbC7Z7oBr+M1PlpMSNwkYJTHuEw2V/syRypdatiCTBKvOf9sKJnOUIhae628oCYbEUzimaauvw
o8nNC6+xLURZ/djTma9KWj+ToqSFgZzfkU8sgoZtuUED1gGGTl9SGBGxf8LHqlp+w1HvXKFWz4c6
nCEDSaUbz8jW6JJQhQ13UyGBdL6EDqiC/FDipmXehw6ofswo55nVOEBIfJebiJ+QVD/JlMIrP8XO
WPOWC9B2/9p7Q8iXD2eBLeKzdwr1IjE6tPvNGvRPyTIL8rF+KzT6aF5Y6L7JQCrWL/83qNztxUit
Rkspp7DlroT9X8syLoc20nORL4Agsi0m+/jj5ZgJFHKIpJo/J8HTe0J0J5LKl0NBggWseKvJ1Jbl
ZfJMz2hcqYzyEY0HJnpt8UZYc56Y1bWbJ+57MnKKkoA5pgwQ8vOzPe3FGry2MYR4QdORuG6szrXv
KLD24MPBiOdMquYiw8p4tgtnpUN0RpGL3EV6koOEsVoIXc3svR5SrxmY//hMBHsAEx0Q2zILnohY
EDBR2bVSj0mWDr9OHxjFtWO5r8yfXxqRtVK9ueByjZEiKvAlS0EScxK4YyDRp3rPWwFa4TbVGx3P
yLZhF53kf3U2ACOVBmXXU9uBvJ7WRzH0Qlfhakfn9JIByuesPLidD2hsjyHQtFB35hJy0v8S2L+I
wn2I5o+0AffQqMe0V+piSQYw15hhNLm2Vb59ClMvx4/1KAqSe3OsQPpBqgTj0Tr+rOQCbCEZ7Dnc
/J0vzvfZR1XnEwYmbJUjJ1KO12MijloKte8autUJ/SHR+cOrpsXWuU2mdRgyX2qyslHfG1Y6Jb9s
Y9AqfWnRrec73sG7fQ9gS24FtL+MmgH/1434BV417O+kHh0C8cNiIMV6ghamfqPAU1z+/95Anci0
ChEtgs6Ha/7kn8sl4pxYLus+xcfPSMPT4l+AmQM8pYXsOOL0fJQY/nAtp6P08++LtZXa9UzHvhRK
i5kcwLAu6+UZpiZTJSwo2BT8Dc/y0oCu/C0HLWE1e1uaQKNFyFbdwTATB3VEnX0kP39qkJ8QqJKo
rwFs7HJFPGRU37HFAQ8UKpzD5P/YLToGbkwXuhPa+ztMY/H6UjEEc71t66TxVfODjK+ujluhScmU
ivqaUocQ8th4ITcidLkfw77BLEn14+EPBhCONEVt4nVsZi9jX5yXCBkuWZeyTf6helIKNndPosvC
oC4PqOIgvc6D8YD0DMFd3snsv5wxZpQLQNk3BCgY3hGj06E+wYmFPabIcIHEi8Upp/9P9/L6/0I9
Afm3pVWuxJBhlkoCrIwdt9PAgcsCV9TMFVOd3JZskzOTJ0ZAIoh2g2DGg91d306e0CDlytoJwS+4
Og6xP1ZGcKC0Akgk489O88V+RA2J1RK8F3uyvDQKE1YpOnwlbRN/zFdQP099BypBUktJQFsW2TRP
laz2xTb0fHKhgCE9cEpmUCySyeBXTMYo1+DTaGJUghBGv12hsMrbDhwzKhe8L760Q5EtSeYAqku+
RMw93mxn6jmPEvMgvLBKRlIpa/D8idN9za6e6dpzVjQSNZP7FI7g6cmpDo+3cYwa4n2EcJwCpEJ2
GlErh1m1OqkfPSvdfOuhDiY+BxS3VJHWb1NqdaClfNLu6Bft1BTK5nJsHLUsjGlZi3zmLBbFij05
zlgCrg5Yn0FfSIVPq17ArhxwxLe0MYUBcOn+xu0lg/L9iwG0UgFRbsL3nboB+8ebcuXZh0VF+hFJ
W5+jZCf4Vasl1u0OfL6QTIOISyybwibMml23BQUsPJgdGoRN/vAyUkH5xPpXKLhF1vnJHw1k6oB2
SEAgO6gINjYBqrA5UqHtosfjQJBuUbo1GdA0ksiYns74g9ivzlOGgCndC5sTVM8s/LSye+1Q9PRd
2xLA2vMOlnnHbs7k8x8yBUt2WcRClfhCtx6V4rKN7w/kS6OmQdlH2XDSvDuPVjQmylF2sQ2CrUbr
CvetxqOshyyStyv8wbXzcEbXDJjWm2w3+bacPXsB223HXfDCWzUDV3oFqRyLB6eWCqQcUJL4fWpX
8jAWnopVBPXCPsyhtTSqM0GgS8WncYr9Ad7FSKG8odHI4MeY/T6VGix36kyz2gf4WE+g4lqe1DzO
9/nH26HSoUe1FCxCbcW8jj62epF0B/L8icSMWrBMfLJ78jVd5qxpgCng7BURgEoPamaURXFV7KI3
UMfKLeTBcKE0Y4+FS4RNKNqCRlnTC3tNBcfQmhb1YzpbmyVR0VpQ4pTcgOicj0FNkPqK1pnW8S3g
fUluRuSUvg43iArb2DI+Ce3ybEK9kcrs/V2YQ8wEVdJIGN7EXo9PEVIYYO6xBzWDX/akfuxA2c5a
GVqTjaXvTJZAeQmqdaWftsMHMMmMfDStcWKVbBi0gJ7pANfkjMZyVYvmN70cg6znus5K0jYobbzs
kynjmjAw/z5/5PVJCOhNL0vgBXWqh9O7NnbWNPkM13KTCQWIMHl/+YuAtcPPqpbzKHEzfJ8Jzn7V
V2KQRXj37MOI3IiAOlNo9Rk06YspYMA8xgZzmFn9AVBGE2/9dfd3/fuFF5dIdVAsrN8L0e3K0tZS
PYOFTCrRb0Z67mwcy2o8Gc1YhRPBSE20gL3C1tccSoD4zoqoFtsLT05OvLYf83gVli6o22jIBYBV
E+ro9X32rhCsWEdkEoF4lJTDbxDYrygsSc+M2MQx3386iCHoUxOX/WCJ3Fs7aFWiX7TDE1c8VA2Y
Q4wYxbaAGu1nf+eh9Gm81aVI1Tt8oz4ERW0ia1ibKe8Ezk5ezQG7pEUDLgDm8DQrhqq71MO3zaiD
NEEICZggTUjP+/aJiU3u/IGm6fdbniI/QFLZRpdalbLvlC2JCOi49/BXbKutxV8Tm31/T9Nc45X4
kJaoODQg0w3zGNy6la9iAhqfhZ4f+2jc02xK5j4ULfPMr+jpwTI3SAxlxnY7HK5/AyzklZNVh8CV
IFsFsddtw2O5wRTSxum2M/jnmeCIYh1c0C7p2uEmlYeEPifsaP2am0PvaGaA+bGjyu1gWtX+Dg6q
mEEEsehG+ZKLk/3AB1LtY+HYJinqreLbNaFYXAKRVO5WOD+8UHHthiRUPJohZXRC9cBWCtdbDzn/
VarpeUa5UzJ4cry/rZP8H90OGrcjkU9YOY04FqUWfhXAlBBxfZ46Cy8HFOrb83ti9CzJi4YemVs3
unqUGZYI0Y/HFATVbxP+L9B446d3EeMUwZHVUws4iW6ep3jt8zhEEX1OEGMnLgWXS29by2qwrTr2
arDYVHOCz9ggUJ3s+VytRYuvFYRZnEKF1UUQsFB8OEJ6RgJA6LbKByxACP7ViFr9z2VXqTpOXO/g
C434jaDgmzW1jGLvirfjMxyViZ7fiGVEQ2f5IO1Z5RweLMjsqd+z5Z01riLXOPQR1RBnBp6GxCpw
QQZ690jieyOFKoKAtqThuLqA++qK4KPXkHdKsoQV9eG0P4dV6XiGcw7iakIWLZ1dWwLBCaeYUZsp
3xLAqvOy6GbdiIOYOHih3Rjuh/zAgKBNaRltxb3l46IEXz/5bpW4WcpiLKMFYtifjLsopiMS9625
vVvBs80rCPMANVCIRrvxmI4pgRrRYIg1ReJVyR0p3OUqaXWMyClO9+e8XdZYSt/v4UFHUJz0Pvv8
iKYhZhydj5fkQsKnTMH1+uACnp7G0rEqwiCAX4228RemiQJW01bXTg7W5kJE/iTUVkJ9lpNC8A5K
RICyGDqamN37N77dxk4H/5RK1BNl4PPgDxcCmSFYph9t9FqsYmPBy1axQIMOj0C8oAsmK6T0M3MV
qm2D5TUYSorMPkchDUNV8hyZnWcghAB+ot70Um1eoNJEnji5iaLQE6FqYpuEv+rCRsoe7Q6O69Hj
Kwl6J/5saJgIj0zgFSADKpABZlgOqkJ9lkbppv2cMm1DOKSjr3NUSehmrAchkSH2y2ZAUrFt9WPE
E+TuD4AAM3l6H8HuwN999I0nciqMs19nKfp9pR8BrI90+hZxwYXTCt1BSufSyQ5hXg7qjZ+jA5G5
QgQsB44/42VZE6qBmY+l+CMQJ676D58JqPkr/1uec+wqTZMI7UKs8DtUQXFSknDRi82W1T0c6FPW
EB0Kws6482Ob95G8C5E853wCTioH9yicDmlMKxdljkdOBXkjBWgfbpPl/Pmcfr7R8B1QcBNz7P29
VVEtCVb38+sHpOiPRQrhOjNmavmVRtlvR0aRejpOXsr/0hc1ZzPblITG/HmYua2urcJ6QpPIsV41
FfIGTw6XckrdYSaYWxEjqiJJ33f2VDm4qaC7ah7No84xls9O+vRy2F2RqxUCcOmc5FT5RPSESEMi
nfpqPqRKCWIVccgwWkZa2PdNoRKcpY547lPLllmsr1yx/YPzS9XZ+osRMKPNxtczxcdd/CTnKCOc
EzctwrHEIAAT6EzmGsa8Llk2a+tLyrwJQ43dq+UGURAh+n6SGJlB7JTrF2Bu/XMtLybQzdfQfcOT
Y9eeeTPob5RgAT3fE9qpwJ+egEFHZ8GuCwVUa6AqxhwVrtjDFp/cVjkFpLijWai/gPaqlQqWVaJV
HohfmOcGACCV7EV3jL02rkVBJn+T8FVfDWDJ94+x2oRZWNQVx+Bc0HukDE0PPQPLpRLszAY7X5x0
ldqE7PHdlCcOqfjAaf4ZaAF742e3BrNAxdNmWWzzmi7S2PvOwBoxUcQ1sr2z6acKEBA+MmwDxjVS
IcFJ6GaQi1P9U+Mf4FzqSVvKa5xJyWapC/C9udMNW2YbwmENBw6C0ZyrGbOx99HRbCC447tpuOuH
9giSYRUgSR5n17oZ23vilBzLZgLyShclf5hEthdebmuGtLaYPHGxmtgLm/z2bGTbpAKqEAr9IPp0
HDrXwrLC7uxKgBKrmj6XX7L069AqT0UKlXv80a7ITHOLRJB+7r5F+RpYxLFjcT6s0QWe/zn6HHlQ
nbqiBZ5EwiTp5ke2Dj2XOkv10dgo8m6+HRJdMUl/Nk4g2ML2+FDBi+c46DElsdj03K8fPrXNQZUv
iRqkI3ro15ttJVDSlerDxOB36CgwH8ckxo0GpFE3/2EN+Z54fmYGbHjatp7xJniR331Q+sTjB7rs
1DCJtpEaRCxHE1eCa8QtLJGjR9RRXLv/ggaGgfFqGWOTvgoaPbAjSI5VtdKVu2Zf0z6Bbq1a7BwD
A6jGmd376iWqvq9y2Bac0aclGUH5cknCKGJU8xdOmJvcHVtUtAO1+mOawp10ULhqpn62Lh8FMPzU
/PNU0CwfGWWgWCCMDeBFRjpeUBpRwI7KjHWhORQBkuv/QHqoFbfoyLFiUtoOCxiJrhCZ92UGsoBT
O/zVY4FiEWqtkvZXML4jtJ/0ulroVY+VhobqytS3LJwcto+02hIF+Ed2sHdNgiNJd85ROLJCSOxR
cuvHz5IxG16xMay5Vpl5u5Rmwddc6VOQbRTaagQZZ+6YmiNF8qSVpTE12BIXOsF1VixintH59n/t
UTdvwGZ9XCIlEk88E/ZrCcyh6QzfTMBxQcGOn5pVirlvzu1qz2tRCO0UiJTvIIZqP7Ql8685Sw9y
wK1cmrZ7VnH3ab9e9WN4pn3fwVoJAQ6uJW9WQN6ZRxXpgMk0bSxDGnfTzCZ2+13BV37SWe2mg7PV
4OiArB14VqfrJ08aTzFNr7LHaTfpYS1m6c0G+on+lWNI1M9H5DzTWB2QP4vP7wRYsaxD19fH8JyQ
Ogs6WYleRitsPmzfF0LMCLDL7SQmMWawzHu22Uk2VWZFX49AEsQqKAqYzHfUbN0tWwDRXm98YCHF
3z858Xs+4Vgl8vqkOj+umzAxk/JBqAWt23q0rhEfiuXVTNBLHNMl9Yy0YCitJ9/Tul2+VQyC2aTs
weU6WC9/K7/AGSPGrksADX+K+6wqUf24L7XqUiRNtat7dm1blXLsNrVOSLw3tURZ4x6/eJByPUA6
PNP42yI0eJhOcv1ivaX1f4yRfQ1yyON5VQTRqlq0aoIdtvYKhh0que3NA27f8MOZjA8gnle2/Nbh
gAH+93FJqFMqUS0Eggg6D6DLxuhZfpXt0mzonR9uqXlQOBVhcX901WLCq1Bsb4O+eFy+10yxfzRA
yysRaYq8xVflpoziG2nS3DcA/XqE4izxGVPqPWwqDKrmRsvmytgFjLjqjP1pbUX+moLzaarzQ73L
AZvDFKhnrXrdjHclJJltAgxoqDAuixckBE8sUhl7V5ZQ0/lMCVAhTpMZyekxXZz2vFwD4qRZjnZI
5YEoSP7pYClqhzhL8JDMrBK8jKXIPLPg2W/Leh+u/w/Oq0kWr2zwr63d4EH3UEySt14YuXrsZXVI
3C9IyhKxeKnMWHWLr8FzaxV0bIXhkHo+6+Kd8bShffTerkySikgEBthJUblG4+DX3LqNesMZUqca
BApektHmpkOjBzDw3pteDc0iDCD3PaWQKOn+Bl9ZQf1W3YgMgalMbDqVTzz0wxls9XE8OTYbhzCb
rEdf5TW6NXwLYC7Nk0AQb+joYxmgTk53XeecRQcKy3plDRy9l898IIMxiRdUFDlGTNVxuZYsHKCu
RYR/bJzvZRgdeZK8WGjh5f1aYdW0JcTK6VT3OKIpAPNNTz9hrdQEGS7vQWmfkyZeJ9gzNvT2sqDT
4QfG35mRefLeQTNEXLsq8MM6xqxWzZeb99JO6Iv8QQD1FIlI82UCvp8WxxSPoKhl5X/5oXUrV3xy
XnLvI6YJSDv3Rxl5ltEprBSmHic+jSLg/CUGzGzMlvcm1qLheiQL3IGzloo3a8N8V5bkC7P18lx9
8UoLmMEHDjckBGdgkH/qsh7/WGnqWp+8oAtQSgnxAGbc494kHI1l9a7X5SpmJ08SKq6QcQrHptMx
ys4sZR697WAPpUcsPIuFVKI28rX5gWWRkM1POLMwE50mC41XrzcPgR76VxR5oxf2M4R2+JemnZj9
Y2i5NwO+BmMKUZhjqn4q6hfQC2C8MLFPqUyMsCD1ccLRuZFo4mf9PC2EQwXEDvrc7ucmBInvaiOD
8EnCQ1yBmIRkhX9Rs57JK5nHjX4LNCfzQvgKlzaGijQvea/SjqJz47LWiTQWDcgEOU8wLzxY2CZY
XrgRcOdvQP33+aUSdXQzZXWLAzNyneGWNDSYBmBfo9Qi7MjgYOEuG5b+mwFEeSZ/KDlqr2wOR6lx
sYA7z/LgLdKp9rYmesUYRjjSI+L12FUH3ah2SIOBxyTOlnJobCpBf1X8F45vQqqeWvHQE7omt4OV
w/r6IzdTu9TfH7Q3bKPTB+s6CW8rgLgPvzDNc/Sec85piWClefqzEK5H/U31g5km7LxxWNzGA/t3
MK7IH/8E0ecBaIFDPx2U+8lUASSjwVHunXmzl4CWvaV2lkPyeqDJAtsCiaWTxqVLdXS6M8hHVTwG
bNTrNvl4o9EVTMYJFRztR5bN0IQAsw4wjV4T20ePUAxAwl0h7T4zZJyWpaV0fN6nNCA8U1MBIHLk
tElqoaLms8bComlrouFA2VHI2k+GHBx5kEk5493/8zvjFRVbrv4fXocyL2TgumaNyLCiwvx4FmIm
jPBxx60hOf7kBgLpwAxUCh5ktWlx4I9kUSctcw3Tq9Z3zB/dL71apfxUwkKnWyI+f02J0NOvtl0E
7n2D8hUc0ncCfdS88lLRpw5WLtZLFqhQburAbh9ONRHEs9rgjucz7nIwIVUSnev7Xc36kxFsAAz/
zzdEmNnLXoTDWdkCviJOGi2cT1X2P2/0e2I3zQRFHmba4PxrKUJ69KzEqpYAmXYjndobNAZm3lhi
wxjtDkbkyC38bVda4OPmswTqqJK/ykH8AZKsFIdT1C5dM6BjKjXFHmQlp1W94BpfVTThI06Oo6Cv
/HKTfntd5OpY9OmO36vDZGJWiH4khsG9exG1zuo91A95ub9Va4kwSiq0F6S1TjxXxAD0KyV9QHZf
442X3hBzk8VJqaV9OOeqWTPZAtuO4j92pTtdMB314QHG/vSfdo61tkli+n4wE5GOSgJFXP5v7Htb
GnTwQEyZ7FKhwhivboGKoD8auqBLPJoO/SKsFGOjT7V0iBFbhSw0lsNr6n/Bnddcjho1pintZ0Wv
egJG080WD/sUQjEPW9jtFVMI2y6uCtsveCCKDNt3goYkBB0+StaM1ZF/95MLUA9cg17AtYBf25Sg
hmhqKTY4LDbx8dc/lzNpTA2mSjM8/FQqVhIupRwnAD+3SqIkYjU3oHV/r/KoL8dPIHjTBsa2avZd
EFIp7Vd0T05NvgQ3Q6dL/A4IXf/P6XisY8xUZKOH/IHGWk73whWTHw7pGooqwTnNIsqo2ShC0qlm
vVh3TsEoDqdrT+IK4D8rWt/3inncGdYz8NoHeconMsQi1F7ghOD3zwLy2EhbEVW09GCx344k+3Gt
zXNMGQdSkuYbv4iR689Mi8UArskuGNeaSmAY2Nf9ptAveQT7P4qrPBWwpFujfqDkOuM/XJGVltHM
K3F0NhO2DMJ/1a2Y90SmRd1J1orb+GvhYN2kNSvGQQdyqo1i9TZYQUYT+T5oEl06+FpAynve4IuM
kMQ3ku0nClGY2YhF9yceICb/WF+yl3i1fWnVejJHtfQsKJiBcOlmT0+91umwt/dLQJE9rwApuOHg
CcvPFuGZmr+zAMfWkPGFs/ImuMelAQeQCcTYJVkS/H4v6aXElISH9F1h9jtcK79crpnwsgXSCGiM
H6WauCnEU//7EUXnezFkBR65sWXoqG5tYBMM+SHwCZBBpN1iyueb5vTMGyHoalLHuyPpL3qYjvxu
9axrNnIQHRsdKYo3yXhuoGBfYmGV/W/HvYTQ5lnrcru2mUMT0G7n2P/RHpwq1Yk7sPu9fKiGzj5A
EoFFQV2Z4jKZFxV/Fn3sPt+6ipejU/H1jUPSD9rqlAGHb/PTkp0Eh5gn8lURYXXhYI3u26CPadhu
gx1nnD+QvYJaE447NCSTpccDrmrX0B7eWzy9SVuZKaTqufTkODQVXmIKNLpkAyj48pLqx8RSGeeB
MtjA8tnOKrFRjtjdJNVy3nEJ4ujwV+3Xm0rQGZR/VZ5R7xie7l42A56MWUcrA9bUA3HC3QCGQTf+
5tlpmUL0IicXUrR9z0yh7VE/B+PmTzbmiGk9EiO0luqB3B9ohwylRddc4wdFIM7xOBHvWL2UcdCx
2LD1jLFz2mifSPL7sKNDDbFX/J29KLzYgI9HCz7bMlWJV0uz/iVsqH60nEnLupBqD3FCiSTxAajN
VWji3m5pFiUH2IwwYBaJgsIlONFEfp5xmhNTds47hq2tz7wuBCCG+qqapMp2pQ/331Eu5OlqfLTa
OehWEQ5RDaXI1jDzvMrPyIyK5ZJm+yYrGcrsBwiunb4kIzZ11a9k3X2j562h2czdBbD+pGd+EKPl
OIXMmZDATiYDwwAw1E5gLSLhmA4ePje3qigk0TQUSSfNy1KOaoUb8vI2cP4MJObibKF+pyZD+7px
IniKRGtk4WgILw7A0HRZLeWBQAAM63cnpypu34Bx/0DvthlOsJdkuFjAHYlPANzEoPGKOx9TnlR8
fKBxfEUjoMm1GyLajR5H9SGj7vcH1uJ7GYRfuT/XkAV/75afOEXpi0HUsOEN+HIerfG/wMB4y1Oc
hg+BI1HLVfTFMsybcnngKWJJ890oUwKk6rJ+64qoomRLj1rOcs8mKJVUystyp46OEVhNVfiesOQ6
QfzGjC9F9B7uu523qrPsxqDiUAYW4NjNhAnwd/WV4Y4O+uv1nsMJY8HOS2cEN0aWSXqOFrhkrIMi
Op5vc2G+nqvh/CvfchrDY/skEFsKVbuZWZXCPVGf/QRktQCv4eEPFScSr4bu2J1O8mLfrqWoBcp5
baJv1+nG1XGZ+hRlZN/3IbKsB0+59IzeCbT/i2faPd9BUiI/wwTYM9tqNZO9jVA3xekor3zvk2PA
royaCxGXbn0UEuTqAcQZq3ewCxVF/3E/aTukhTDpY4ZUPYufZ2yqJYu2fb5U/qaUy5RF5mz53lzP
twD7uxewekP3B8LXaRlUGc3TbE/XddOcQQcAVdd0y6QiD8Y/9hEWyyoHQwLAVfLzNZSXLJolpuOI
Kvv6Io+uPqxbArtgT/79EibRrLiOcmm8juRsA6qxudKh3m01ELPMU1DuCWs+lyzdhFLa55YCWnFX
zKyLPmecqMWvpPwzB4wXUqlEBKYNgR+arMOBfZctCvqaml5IZRyiAtY2MiDjqSNWTiG+U90UcmRV
AdntLJVBKBbAtgRSMuGO4EyjKGF7Pl3YfWwY3cKduyoE8bVmwoPOe884dPHRX6cSgweom5SGxeSS
x5JnNJK+fvRPtwDP+eCpdUz8PJ31gCxQEJEc/qJeQfa3mzmf25o6oi/MFVn4glbA7Os6rjxD6TfC
fLgKHgMocTSpVBvRPKvqZSIDI87npWGb2jlnT3Nul+cqRyAmFLunnskVFwOVHAB7robvrbQYWkFI
BbmXm3vP2wWs60p/Dvm4/PbUYrwClWOr7XQrxZeZxkD6FT6Xtn84gOyEw9LNcHaL+suJDp8c202r
D3kFmdHhVyh4U6HXi8iKSbNrULgJmy7RlJBuQeRW3uLjyYmiH+nLp4GppO5XOjkYZd0T9WTg2azf
4qxxN1qnYDE6Dhp1JwRVcnYn3iKHuAm08xNczQHYoyiR8ZKl/ATU0sXdT5CX639C9MrO0MzAjGFs
FbF/Z/p9z2Muq4SJbe5ULcuLL10QNKOvR58G8ILkLBOOecoz8/krgbQZ3yZgeGgAVqNuvqv4Ujnn
ZU3v/OK+uSlXUz7SqCbCBzT68LAU2z1hm54WeqFdUomK7KNHim8oNGUOHDoDR/38nT6gxWN8kEYx
lrjARKuSIclm8CJBvIBrxAiEOZ+Ca2T3PIOrm7K7OZZb/2nOBYGkY0iEUuxZu4m3tRsQDLrtf+jJ
Nw8RM68ANUF99EDOw6EwpsNAtHlbfTnXALLFfb6ff6yzXVJOTA7zTXtn/Gmm136YQgeRkzZz3S9Y
YKbAUJrRBWmQke4u2B0K14FvQfbzqoqYvuepVWJO51G7wQk2XVHQQz/QowHSs90qW1XmHGu68Ao4
WByLZGdQVywKaTRMboWZ7lV0HPXXAV/NJqorzONH41h7+d3+53uV/hHI+iUAsvw844h2CseweJTo
kHwEzz43l7nfk4AZJ8miL6nNI+AbG/VAxSHG2GpFyFs6G3Dm0dht6epf6ammEaqSx+i2Ba6MLA8V
YdujsaFDu8m4bcuhHy2THsw/O7PuXdw5juFmzBFWZ4QPAy8spet5SCZ92G1X6ogEhNnE6p09Wf7P
W61LtdAUcTYA572er7yZEeAhlktoGlkfJuO6BcKBdTE6Dy4FwzybUHf30lVWs7C+uPWcd20VuMpe
7BA4vdOhbhRPu6WKIvPvy5PF3Z8KDtq1/syh4dy0UMVSmiGYUEqeJ47XiA1/CeDvqH8Qt18TNxlg
oZDuoePom88xxSKlqmz2wirFz2Cikv+i4hJJLUS3OorqAgqxyHhtfkvHeiWFrIIM8E7HaRHv2OPh
j4oknKdxYpa3hxGfC3bEwT6zcuvKDBpocEsdivysOvn27Jx18ICxK/mr68hHkjZfCVnhI3x/8vcO
IBPeNvLYHRsWKnqDZs6XK1UKdsUghqx6zJsBljZ8uX5gws2kASTCzE2tpbYBt2UndjAK82Zh8Utf
MqDqtonEj/7FaQnlgB6NdwiYtQVFVqZNPQoqJq1ZdfoqZkAHUubabxVK1PHI4jLLt8S2kX3e3Sq6
pSPhGGRKWTkkX29nrbNpv71SpHiscfwYJX/Ufs3x7OqFBLfAfuVAg1bPkffNyxW4lzSj2Stfu7iG
3lzbKtHvAmFzBqbF+okc5SxJoaB3pPkH8rqgeh+JvsJxo5xVotR3w7OP3+UepJPwjvdkr1XCdHP5
R9cDnhpsNo1YseUN0ypkbXsVuxlq9tTsOmkJQMExgQHtnjigUpF+gUcQGSKILeFgAjKYJS9iRnie
sckScf5G7onT908NJ59H+Slqm74e2H428IOwZtdu7itwovHIOYH7o9X/7w1qcVihg2OGKcvh2G4z
coR/pOXEaXnPdBNde4V2mK9SM41C5j3CzSVXrembr2Ty5grmCy2F5+mUMej9sCbjRT8TYmuNNa3q
8ZX11YtxNdZBX71fMjwmh7QCgboPoF9JclO6IybWEP6qyIFNmVEWUh39r5OfoJgn1hnNb01wgyL3
Ih+v1i4ovCmBex7ngfs+Xwj3ryr+JNEFaNuRxLJ8FLIzl3D8f6P6q1CXf8+I6Mhf4s5ECvlGln8x
+iWdzFk1H/XYpRfR7EJd0puqDRRoqh9BKJrhsAkKXNtcx0jEajW+7/l3VNpxU1uaG5ehanWGCK2C
llg2AYPfBAc8A74RztfvLMfS76Xx877jVA1XzDYKnZlwMNuHn3brg1Q3YCM1lAgGtt3GOhKWCXA4
WK7KB1OpWgOyyKP2OB6wAKZqypxHtdzda7G/DgWX5IdnPxabK6C+CqvC/GZ0Jc/K8p4eOIgup0U/
DXMo5dzQrUuya8u/M666K4bWz2ZpebKDNnVgn+N2SnWR5TAl7CE2cmz+mKffXMlAeZbLSb4KJZoG
Z/Mf/3lf7h9mLjzQ19HMAWAAL1wZHmGKvEBXfBMVMvqi+yPe4mQfeTJdi1Uflizu5DAvI+DIx1o7
GdQYrKwy2vvt5OjM2psgDMfKUIt0chLxRS/Zt1QXx95r+Qc928PzTmG3krxAfCzutuM5S+szNWzj
FbHwmKOYw6Z+cJjLvEZ17QIePt25zE2WxnsjfqMfoxoRsyplOHuVxVOyNvf1+IVCJMGMIMXzXgS0
KqSFIESV4qJ+OgLqFmSIJIjULb5gWWgneqzSQdEMMsHNI5UCexdE4BTksEw4Nw4VJIuahUNmXORM
PTPa2AqjivAZyGa8nqaPyNBzmL9/siBW6IqtQ1WdgPyv8m3Pkms5y5KWg7q6jS6UAtFXVuEh9XUS
r7X4Mam4pFU1qR+qxj5rv0j8ncVVBsnTnbUq6aoIs/OvFZIURrnHtty6KSzmkQbWxO+h8eioFlRo
CTjd+FS3LZ+uOcOvzX3dtZcIu/ejRZt2JfCuPEm0/y9gl4iJuzk6KecB7rRmCQOO/vIni7fwtFku
qFhqHn6o72T91sR4Em7uUk/2gXqKvOkiGj7R5UguP7JmBrYzQch6g1XASnVyYAcIYscbR7OT8ldp
1cU7D1vlvCrDXzletTMomTTVRN/S7JTtbUGh1V0rUkwZ3K3osnX6mG12nVgaYCNKNUT+98jv4IZI
5Oq/CSKgH5shYeQECCzFiiWxvZJ/65NO5XCJG12ncruzuzoh1PGQJ8tG8PrTVxvN4l4SitLifQ9c
unkpNZIXNiQm0u2y/ul6d1yE42d25FXvwig9u2jUvpQ4ImviJY9jik046vXTG9LAzk3jBHjbsDgG
JRemgO1v/h3Funfma4IjeEd/uNgKuYo8SiXGHcVuDyV0plHoSRUe3YzGuhruk6+ysY0Ac9olDkTI
LBRY67n1dHaytDFakyvCfGpmXT2AzkMSjfDWWSuNVT61kjmsoLunEPa4naPNpjOkPrEnDS+WBqgA
xrNS5MS+NOjT90C7Ps+T8jq+hO3cyNercK9aTDix+KtDXrVQPg3zpDtPx0R65VzdsvYbYFf307Mp
yMee532FElNTZ7F71Qu5PmSwk2FqWBid0dyD4hToZSsyvklXVOwRqDVnGvrJ/kh9MnVo2EXg93kc
oGN3dfaCD82uyMCFlOiq3kyqmAjc0PLH36GvTpH0xLk9+D34IA8tbCADU9/liTZlD3pwE1k37VqP
cHMhbof5Vfy+CoCM0JLzBiHGLCAfV7bacrKt6i5i9Ie4uCTG8jHKe2lybJOnK5jticekSlfb+gx3
HH2/eHTlNEWfAfzOLEKsAp98Z1LPe+2oboeCQVYr2zekTfl7RPjVIGyh9N4bFn/Lqt0IHJ6lqGSR
2pEAdvTCHzyK0KNcASxlxIBIYwUJrIzthVKaG3oyEDDQSCKFbe7ldeGqtMsWKKNYV745YEfoG7m5
vPZ3C8jIIKe/dzQ7WFwmIDSs52xhXeOnpWk3AdBvlnyef5b7Dsr9h7XlMytWn1pvWBYh/5NcJJa9
ntiMT90gs+IHitKXfhkM/ISOqMIfYVlQUQiZOe1+MvWpAxUhHu6mkIYOS4adWAplFUsIhyaqLPmb
wqqrPaytfjfWEUiaiUEcrd4gdHnuOaTsPKOP3hnV6kGeHHY4sPZdT5Z+EvarRVeFkehJZWbdPdeU
gY8oHEw0Q5r6SqjkZg14QffaBFZZ8tr385MfZLaPQQ/OuapyUbZUt8XbJ+xwnnMNMEKO0+F85U4g
/JGrNhmeCX8Qk5ZS/JaxRC30lGMGYlt5El84Mv3Vp2ytjC5Z+ym3yowTnGaZPq2VScQcKLXDaDuS
ApXThWULxWxac9em/SH2ad27QqM8IcGewfhnQOYDPjmkG1luXf456nqT2HIVVagFenEeIVVpMSBX
J96LQDBW07+1saYkjxicpw6ytVFyVL+C9i57hczPoKflsf5cSqAPNnQLdPnOE5tbh+/G5Lt5d3eg
VGA9lB5gpI6MeTGidsuuKEjDnYD6tLAY0H99Vji1Lvt2dvwOgzeOdhhUhqNeZPENxJpnRfAwKxX6
O+lRpiq3pZTvnneyMjbxSsX5eCqPVzgCC/HHSWKiKVojHL4gqSUX47fwQhxS3nDodALxSZVufDG3
rKLM189REpIj11ZAvMB/rK2pw7M7/Lz4YayNA+nAlL31Mxr5Pdv1OboTvX5iv0kawR0kNUceAP9Z
fuQ6rZU2cJBZn+N5FGbeF4FXMp3z0cNpr3W4PlZPyBDJVNqAxrh79jfqoUafHJGmm2HwPyiGL1c+
y8ECHHlKi4MU5As5GGmEtOACF2/rJB3RozCELHlORhGaZRkvYFfLLctdLMy+1TKCcq7eBtei/yT4
uyVo9ylVt6XQsOB2sjWNHH8IRo/6z9G/6eqaFVGYJ8cFoEgeTlkfQ867EihG0QUv3oIdOz+CeY5z
6sBqoN7r7VQ1pMbzuxWmN4cfweSe/b42U50P9s68Opd65QOU64LXJLjg4Y6bbNLqubjVwFLEsxC+
nB7/JOMQFu0ZwYx/MTt1G5dOAN0cZN0uQQiNhQMo8GHEoOT9L7i6FjIyMIv6HQ3pvtagZJlUTHdv
8QtVO1K6RcypH0Khv5CTzKqUShv4fywD/btNR8I0Lj7D1Y4n1+EnJDvz6GnHN0aTzyb9u97QX/TO
vGWHA3CLVBgLn1Gpm8v/45DDjSp/+2PPjUHuYSELvD5cDUvPV/MvBj+kOWSwK6FD3Uh4fV9vwgjy
CONOVgxCN1PQLKQ2u52Moxl/ULQRGRRLHWedk/TANcQQOq5BnUlP4o34SLL8X5OZCgV+Flyo0CcI
ZLapejZAQ7YPurIRPhrSKz60bEXzYDyrvSwIkCwuI3BHTmVPgcgwO/kUTEP1aeSnrvdeR+6xmoGz
OlhiZp2KuWr3M8kjxWy4Z90t8jiYwVrkQGrIym2SktZ0NhmzspyU5lGhY+NDKlId9IXeisocf0Ar
7ONJJ6dQO+qAKhaQY9DmChs8U69HdDb4iEYkFe9/FFr5ASwSizNz1NpOgTJg5a+lPDHY1tULK8Mf
CwtXMFEpLkilPAa8aAl8/EqPROMzZU2YPrS9+6Mm7Vsz6QPC/NLGfJGqPhx7bgy6K/DRSFMBy/hs
r1QsfkqThy/w2eQUNd9slFPAjzH24ReKEHJDqS5RZXZpe86I7OB/mbexa10EqcXs1v2LfkhCCOhm
1sPhpH0GpjfmPYXsEbtm3nDXi0pIL/5wQK+VTP6nrhQPCR9K4dUC9MV8r2rUbKi9uF3YVoBWNX+U
fl/y8Sq7j3DTptaH3seFsZHgLpNDBL6PfSn+wpjc+Z7AaDdA44g/+O+HhlLhl/yrBvjn9PDvWv7h
swlk1Gcoa1m3qwOxWHxl3FYumgaISV+4gSxvRcrihJlxYJsiOEjKCb39DvRYTYSQhx7IBUkRbYMx
2eDOzDfUZLJCxaPCIKtTR2WTFuOCE7DZATK7Pi2pVMDB8Xk2fXYL5tU3AVwnMDIswtRR2FEaufyK
035NZvJnf9tQxhr9L/nyTELJlZh6edgoHGzDIqNEk/TkB93k7o8G4jeDsyKs1cU0N8ZgFefj0x/D
QybMif9Z8Sm3MhhADcStkdTYwn853dFRvRYOu9sia/suolxbPbQZxOoM+9JSaxvK5Lpy9EdLBI4U
khA6kcZYbMVEuGsO2VriCghaG+fh4iQDo4iBrMW0tcf9QV6azEbcQd0zQjSFZ53pnM+oijR7RXQq
bXDNYQBKhBmctbBEtO8KVW6g+mFB+tmQdmXYoXn8ndKeXumUNXvagFetM4pWTzDkHG6CKDW8P4vJ
pLQsB2cMVOgFe+9uD9e/dbewZ15H1hTalGguq3EgVDtb/PO1XFpiXFFgb8V/Sqim1O3WsaCxdJz6
A28V+ALr6ZOmCOcMGT4XKfHFGPo5dg7Imlmq2/2JS9EaHaNZjPPHNHHYHKA9Oo1AHsWJGm1LIXz+
/r60NgMIb5ZlD48Su8MrmDSIDwAcS0YkMap7tyf4dXksUkbrKu/awJc/aitBE+egFdKOys68Yz6E
GcewXuyRrCZloW9CpQ3RTu4Wywb8SE9R/L3S30v9lbWEyO5sR+BE72WKUMo1i8YOj07jZJ64DgZH
kZuMl2VbP1AXlePOzSXWu6WAn05/OsLphV6xKTUacdX/VaQd8e2kngRwo1HrTluljpZ9i3dkv8Zr
rnG3fPxXT63y6dSpdm3LbsKPwDP+HN3/Cz4kT2qY+sa3huxqhr+9Sd/Kg7PC18jm23K4R7ISNZ24
Ng8wf4P9ajsbvalrZS8kslgrpSEmCtEbWSvDGUyu2q8bNOYTZRv39LnkqBS0gNPBapwN11fKVMfR
Qeu8Kw/zZwPzGEJGxAPUMmimo7qYm/MJL7KGE7M6h9fud653E1dfNPraqKKfJzu/T9/erRziZeJd
5YnfA+GOjOhoQjwnJNGQ+KdQL8ClRfDqxcQGA2lfcWWYAbALf7P3p0ZZdgbneVk1HZFviz/7pSDW
QKxd96INxaSkFBgCN2bjsHvhAVWG0GPWAoLJJNlVQgyK0KKj6I3EsQz5yinDYnPJrwMsdFxjPt2S
BFQ/7P0t9ejxwLkU+UxA0sxcgwso8Q9ml9fSpWyBb1lB70+LLcd8kqo3jp7uxGYLtFgvxIVWPZpC
iEt/xZGSFJF0fYXa/pnVVc6ic3588YexQHrN8fTXTJp46u0B84CATfdMz7/INQNNs63GCGku33wc
tBcvYpjfzJdpuv4BDjYgS/R+bpP1IvG9r+b8ig+DEu2RapTflM3v1ZYARM9CBJKAg8zAFgRuSJyy
8B9fPMTRCuiqqYT2+jKtjAQI4NeZAjlC4MYaWvdZ+HlYQIBbDZsfiSyc7juDfS8pV7he8d2XclZ2
7DTMVXDNXdcZinH7m9c32aeGYaoE4QhBr50zULKdY0HONXuxjBgmIvl/QDhl0KqJYeiVtiCStHdT
GFubksA+hW434BuFYhducsRIfasTRgO6jITYoOuxN0/eWGNvXK7pIyDG8EtBmW1BOyvl9m+boiIp
IJaw84gXpoQa3I53bxv7jt/5EVHfUD12KzOH16aYWqQyRSAcmIQ1JKeOzSsa2nFinOGE0XBGahIQ
F651LbrTr+o5pM+AGnVTBqFbuPyIpkXhDCaJKy9dNFwHAzUNwutF5ymZJxzpOusZSlZ7k25SarBJ
jgjb1znwQzyr2Jz+WnD4ksRV1uB84HT6YSSDVbBChK6pJkcHOneQs/qDey/VtTsxhO+kU0Hy3ArP
oB0VW0zSPrzDK3wkaHnl4e6B2WjfYpdGDMyqMUWnJAJj8FG7o772hiyPkL/iDltVx1HUufpy3zsd
8+Vt25xv9+18LGS/lOXCyQ98fgr7z6+ZOd3P1Dk05LiFZTuYboQV3G8EzYHX2Pc/Q4uMtm+eA+nV
68ufPs7k06LnXDcljuadCEwZq7B+XZApsICm5Z0Q7O+bmHkpWmVYXSqBTSQghFHUFzt+8KcUhSgU
CeHegAmmClpzfA3KYW3Iwj/X/oZ8mwneTFdYXRfWjv3JvvklEIG1WoPfNhrLBIQV/r70yjL2Mufa
J2QrddQ6ahCW5RBPWLyZkxfdhGQgOhOko59nAxqLnd6alnY5xSiAH9LhFDZQF22aFblXCYCv2teA
4R2O+3e8RJdzPlRWTSplSzvgSyEc5KFHwQBjlTVrWcIuZ8wrXIcfZP3GEVGUUVnOZ/7+7OSF2+dH
ktpSr1Wu/ADNjaX7mPmNgVC2XVZSGHoaq3oKg1FTiIhxk3KsV6MPfaRz/VffSV462E8mGtMEjhJ2
FEiX6Pt33GOKOB6XdELCozuMYuRNtqm9MX/igc072W34V4vWVtb7i3cidEYD5Uear+/4GJ+1zIO6
AIgXchXpnKJQ0u11KXHl7wRliF75T00sJMLItevzpDjWRXYSTqSC77XaXQmedOEmhmDh6bpgg4XH
cycUBGIMMoHo4Q7o1RYSedLdIBHxjgJxPBf0y411BSrEZW0oiRoDaW94dHTcl/kvre8WKfteS2JE
Tc0B/dq0ti/iIbp9/BYHIHtroW/+3cM3gzWU6ivV34A2g8EvGeDuyRaNPeSFfZ6KFYPxC5dHYNxD
U25HJiZZW/arz9gR8bHtBJLpk5Cb54HweQaswTSB3KocnEoAL9o/MAOv+RkpzKOh0c0OTZCR38lb
damDmh9vd/Ldc0NWHSFTSJdLbgpkMJ/Dwef8r8XT4QgatAYG0wQN7NrWItq861lxuMn9om2xFnpa
E8DUYU0RwjowSBOSWYAkRzkoIHT0DTeWHTNZsXQtd/lazmMAAaJAVRmUZ83DBEZusDWv+RBvc0KZ
jekznXVcgKjIqvRKZ065CQViF78XaloRZIJyexkvXIgdXEV4LhmEuYvZ2pa+8aocqLatG4ETJ3Gs
F5NpVce9jnYjP2jiu4GJP6G8ngoeIZOFsnLUYnpHrxtqeMSvZn3IQZuTCSNMRVDKB689RXbu5NCb
esqsUmNThB4Ji9zD6AZVEWWwFhFo5sZunYhHVwvOr9XFgtvyBdNl32ntNXH/OTEK8KHunvhzejQt
DFbbOBH8F13cdJNgYQa41PwG9xGp2EnBA7oAD5QGQRJY3FXGMai9Ufwngqjd2acqYRRqNOg3YBlG
z7CxBbLxChGFv7fZaLYsxyR8taY3pCcNu+HBVIhTrZ8+vIP4sJlEkzj3KpCEEr/ErRdUugxHyxb1
U2gAFdgkG85fp9HAth5cBg4gqspbNTmq9zeQ2ZoyTR5H5aXTPQmH/+MUEz7DSan8KeXPVlUGw41P
Y7VetVi3qA6cL4saGa+nt0hMS4QCjww0KFNuH/YvhIq+3g8kB1jLq08yDChT83a9ToFj1c392OS9
eA6/hkEIUq+ZNx6/sY0t3NGknXZ5DuDXCUPcVECRRK8x3PeEQ8YpWNNIU30u288Dd6sNYFxtTd2/
tO7zNA6w6cloa0ksz9KUxVDAj/RTJueueugLw06SBBLACoqUyOK8ecrUgM6Rr12CzHICBS3J0I4Y
UEZaW47oVLO1L+fCTIs/IpeT0DWz768B3WboVTPEu27s5sC60nJL8HDQF9cT1PhU6Y9gpgy/RNNj
NIQR0EWJ81Rk7c3YgdTHH3I6noNbfLwgmIxWn9akEGDH3K4h8/fHbwvGE6cpo2RXUaW7XCClp3N9
tCFbGesxmC31jKlDLBCJMUiUuiUyuOwxiLyT5IN8Uwc4niddJthMXKW4GFPOUerl+qlfUF7RbR6m
/33MBuoJNiavKZLqua/mrWwHXe5ZwwRhEQUN6sKPmv1dC9z81b10nWVmfAeWYMhycsMfGPV+Ec3Z
JLFWxOX9kjxl+kUqnvsc80GnG4mfHoXfNvX8kbhG8NkZPFablpzB5ncL2BZydL9jDIbQye7DOgHI
OV5Q9ftDYY88x9za1zFK2LpkSgJUDgIwgzLe9ViGg3yq9aNCMahb+T549lJurG/e5/noYgsPPiSb
1lknkRMGWG5nT/CzjsxAqyE31XtSZDxbcT/SBwGTOiw0UWegWeTDx2Z2vOIxzb9wHOo3yxgWh2Fy
WI1BlHzdy2EYeseRYoC+ZuZvXTjVGz5j2B4JjHSBGN9Bur/SouFas5/Bp9BrKWV9RjacWgE40eOP
jkf1iCnrGedHvDPjWzj6DQZNDcsVTnRVT277DGj0L26Cc/IS04u7msGxEb2nEhiMibyDzlKaBOK1
G5cbWHp1K225xdBCKXCB72/FTUhTTzIrNreqgTjAsfMsx00jDWrP8CpstW654oa/teaLsEH6L9xR
JQTwg7LhUGc3wV21xvuH+vyYSEzkmddFWobWJrSKxD+XFVOzHKaKBdM5zKSDz5R1AuyrtN4WOGCx
BbkTuXcG7nxRFSb4blx3zprpaZP/7JnSkOQ/YZX2f6vB8YxecM332aubSfn/pRSrbygqHOniOVyX
WaseijlRhRo7J6w3ZO7M3X+ZjF/nK0TSOPQ6dKkUIUgG5ufRNKqzMj2/Er/WY9bZX77X4+dTjtx4
glzfTyTFnd018dy9kdVRtauChVDbwtND0FmZfyTkP7YowspS5bbuuBn3JpEz8HDaINi7ovrGt9nk
/T99rYCRzO/J04YPnFAtWfs5zyTSy76YwWes4NBbbw5CKbfK04bJC/LE1TDCSmKcU+k+NMCchpkl
1JK1vknDJFpvDB7Vntvox3G7cOHkABf8fmew8okeMMFqrTlRfoEEmcKBHK0NVe89wioRoQMSHqWw
UAc2KRxpG+UORkBHLUDaLP4lEPJGI9NNQNPR0e7MxCqr6+0eSC9sfGmo9kdfiBWK2BZhkyWRdgiq
XmToUGCmLRFeHTC4F2IOfYa5Q8BpNwT8BFcxZPBMz4j9fWOQ7U5ViPJZJRni4C4AxeaAF1qjMT2c
kbxWIr5WM7H4HfUWgJq9fh+Y4zp5wQKeDl5alGYPQfzqKlBpe6fcbAeZ9HMvbpE4MDS5RVF94EFY
4MU0kgZqZ0spnJPeFFxSabKjAMsx9mEeeNwe9arA8LzuMt13Cuha02rxuL3zV/h/vq2lO8gyuHGb
8gh7NqsUkFLcIfEVNrNNWLfFGPys3tzsDdvn9kGI0KZl8EF1k3vpM/kkuS1jqF4Zm1dG+fc77FQa
enKVMkRnazXHfiRa/O+DYusY2cI8ffz9XswNaN5diyX7Hx3+VriOS7lWKQY1xIpVDg33cWzM+Nd0
BRo5jAj4gcls0MRheyhkjg1NgvUKYZuGjsIvKRkATy4Vdj722yFKDDGzdFi1S051b1sPtf/GCCEf
2UBm6zEtW7ZH1BBqNrN17PQvpHemNcts5j2stE5vc0eQ5lx85bVlvzczRp8yAiezvpp3fJe9wDPp
UgV65rRkFX4EY87qozH3Hnw7zhNnhG7of6JhrazeNeuMvMdOi3dgEUNIx/numCh7xZEd8hayeEfo
DRylFOSrYZqGyO0zCm/Y3ACvhSuOPwJb9L1A9FooK3/NoZhjwRlc+Q3nVMXbMivG6Z3iUaUsx5XF
DFba4VYz55Lz28+4yr5lI/gvd7L0EwYPDp7NOcyDycSkl4OklDl923F1x6P+NUxwMz/e+ksZY7k4
zSuR/TyiJK4l5CRm+eJqRgWatTO72ERoGI5zZBOl6EkoFdkQm7wJrHpJY+WE//milAJhXPwl5qov
7SMgHGZaP+mIxGBQNQWmPodJBTYUwJAvGpjm1LegmgHoHhk0QgDJc0vWszth+1z662ip2Sof+0TU
MVm4Nse/0R5ilzjshDYzioKI3J7yihNCwp/yKJ4mR17IDJn98k+LA4L/skOS+tDrChvX/i3rKt5S
nTt2r5+q2nCGQseFwuKq9eDuas/j+D/bUG9wQ8oAfCK4rkXeN+BvclGu1ac4WJgaSmnIKBsg/bQ4
ORz5IOSbMElJJX80VIJnn5Fhtbkuy/21LumOwaw5Mk54WRpoVACCGSmVP1iFlHWoVr6cRN7M0e7o
jQK5SVd45cNkEirKKJQnTf6FVDZud61CGMq2LUylLAo+Xg4dAZK9WB54l8H+nIKZm8ACfrNYqkRB
lDIsNcr6Idk50SZUAAhVCzW+yWPtolWpcP+i49JKR4Avuk/PIHuRxPWlKkMjee9HxwL+5Yjip1IQ
kmVLNMSnXWxYLZ8vKw9ZHvh/PQrkmBQbzwScGISOKi/SMMfd333dBbigxLUirhraPd6Ye6ByIf4f
LLDClXno5YNgeGUABjTeno2pkXJpWXw0Qtp92jQ4qzswWrb8y8xt4x9xGYoHAVxdfddNfJ6UpDre
PMV+IvgA/JdtYXyl6/7gypvYrqf5v1N7iq0kCEwcjC5cYT2Xh2JFkBGS/rc07TI7AzB5o/B0ndD/
1WywgcMjZh/6UUm4BVe93jtZkXHbTymqy+OsstcfVgyiETc2pFXP6RWudM0T2LCAbVFOyQdqwQCL
mUjXhO0KWuNz6e97n+iolO/+OMFE/RdfukJCKzfA1mQlP1zIYPtkKSeziBBWr8gk/CQTfz0Ilpco
b9zp3C+0W+V148Flv8SO+qiyNS4HgNL9iNnYVJPkllQ2R3US4iL451sm2GJTCt5SfnYH37YYS4sz
PLfNnxuYYEQ6JK34FgKMyi52ilErjME0Db0NyGKaRJV9zG6vXzEJfZLeUiHQ32RQu1/T7Pm7hRWB
gL5UXK6r0Z/yHfun2e/FWfukdIlhQ/QtpNLBo2RlQ/FEqjjtD+mDUQgUDFOH5s9jh5iI+ijiHLxQ
h9LLiXk5bnJo/5wxJOMt2p8l2Jf9WUgKGOS5oOteGDHORgp6It6Q8u9rMskMR6geQTuO2zZT7pLd
tocW/z4xd4yCrmcBQTbCIfY/VfvCFMcIBQHBPIBYLcisowyuuk+lD48SvgDBzzqK7ICpkemFhtmS
TxB4nxNQ7HF9o+YaDeE2IaoG4+ySB2Sd5iwUJH2tuUoYnZs7C6XMUwLHyv2QUwZRGa9GQ70DXExz
74BN8qPUT7W1GNEyH0M89F2sNIL3l1V4SrIM+GmEO6ONxazJ/ChwI525UC5V7ejT74G4tLLbMgxQ
trnrRx/RtfWg0uJK9jfp3NYyKgBkrxZ+712lR8ORAEg94b//78aEez0veOnTb4vTEWEagvIzcm5G
Ip5GqD++uD8OmZbFILrOTuAQtnTt+vhTWptziHIE4V/GkB27tjzPRSErUmJW9T0Vie/7T95mc+9t
LH+3yqpUY5nSNKp4opN0gKRb+/IABjMWWOWnQXFlT2TOPhkfkdq47aHzZHPyrSDKFGS1UUGGlkhb
pPAwAWZsmWViitfy9b+1hO4t0uoAzd7uGNrJgtbLerNXZpB42ReKWYiOHgW3NdTvMURT9oGIrxNU
8MtK8sn6eaZKEGG88AKWp2pd/wpyi4SjoEbESylfhtrA78TyISZmNr0/oQX0Wpm2iqSdvO5J7QyM
U7gkWTS/lhHiJZJlQ1HPabdx33Xc2yhTFB6Nhv+hlUbwamooLwcgVV9wz2dc5wueEVzufMcE1j8q
ZIGP1uFgTT/l/eLMhKfzA6CoBq3tqHOvfcm2BWP/JKy3JZdzub2uYWpxqhp07nKeeZ6KYLAtaqLN
XSc1offEftoCwmcSK3XoG7Y6taVRd0WvdpnjqWr0+MGBp6Nixx6UBRSIh4j/fQDJu3TAc7bcJtIw
07zOg6oICjvibD3U1fUyWiyow9hxvcNsSE/bNh5fYrBlfGW3xqpCwE3dP0peHNGrnHinMbW6+Q3B
vIZbItX0GWHVsxmRzmAXc4By9P74gsNcYNm6Qw5QYblcG/aptDceIA9gINfn/ZD2wMRWR3mQ5ZWU
101+l2mCqh2T4BEf/VxZNEnooiHA/wgkQLiwhmeK7r/keOHst83PY+teHr3I4u1ZrhdAmjtzc0Gb
Ruj/iFLSRiRo+qGNyiH1Ae/Gv1EUdFCfhQerxHkq9KBYYSLdaNosInMSar9RDkmLnBW31XNBDEHZ
SOm+XImfCRpf/NadewrB0UAH0kjsuhhTFyxGEM7tP2Sjk+2avgOT/ceIEJuqkt5Q5/GksggredDW
ma+UkONgTVYz9nPlcZPvj9mL/7mYSPlsxs0G/4aonshhvFIE1DuMtMxZO/9BNDPLZQhOs40Cwb9e
h8rf3IXjurGBSL0HXpDJBZFksCXIlqVUR1bzr/KeLB571/lxPWKopa2lmhZp2kRzSw+HOzvL8mTZ
XjgS6pukqmw2YBUsU29nRmFvy8Pnqn7O1wIJZO6jjgcDBO3qQp/C0me8ncCE9ZT7t3Tv8/kYA2dD
zad8QX5b1ktmQE6wvlrfbYapLNmEKA1EhPs9c/A4+VU2rLMMAwHfTNHrSJqqCv1++b678+YS5MpI
m9ro7VqPq4xVH129iA4pMFn6x+JpmqxofH6VSvFp/OyA7iJZao1rlEhBpzDjFLpE+dr6SmC9yCtZ
gnq43MVmod2CGn6FoCYBrlSpla4Y+L7HnKjrH5OG1IsKknTZ7Mu1DN6WCR+7GB28ZhtqljAoVbHH
okzCLK40ba/4/jl7LFzdp9W6NMRCsFSLoTvjexg/H1zJV6kktyAhKjSi2ebuABOSh7n9mukXL4vn
eyxmi0t/DVDD7unIr+UatB/R4bk9jNbgs7gAgfFlSulDLooN6gkmB4J130H92OiuET/aj+/f/nxA
zxoaGg4btmhoKcBs6lphNRzyPn1ASVWRGKG8DyWb1Tr98SxkePnhqxCYVJX9M9HGW46jYAid+mH1
Zxdep/oIfl1aIxocZ/7bbXtrt9jP3JutfQEGXqBIiFA+Rxr2YCLvRkPyAI8e+OZ/iOMXtCJ9+bHD
0rbAqmmqWqjz/ZcOGthVB6iOK8M0Q9tOceVsxItOSq1nakodWA4WZ2fSqNlmm/JftgVKDKQXiGMf
STvdhf8ounM/gv/oyoTiSJcHGH952IQS018YyKgm1f2yZR/aaJ9KHFGlTpAh2IxJ4qlxgUBVxWwy
jRZWXLmj8xDfLY96VBoj5Rr+RJQSW1ydssBGCPyUlrU81szbRBJd6kaIwW2YQ5vjj4s/CaJxAVZM
i1N0d62UQ11/8tYIsbWnymIsIw0K4HpyPEaiIFAv1ZM39S9r84oZxWd155cv/QGUCh8K+Rhx/cT7
dxbehulCNOfN/4mBeGMI2NP1gDRTOP0IQj+1aXwh04Mwc5AbOCn8jqTE03K1zmfIynjkuWEnmzAP
Wp7se3p04CQkemGtl5jdSofFBfi3e4XzA22fqKdetHpdndbhMhzqNni8iuZ9nrhOKQiTkXUg0OW+
dIQ57u93LpWiFXtwjJZoL10DXN6l5pfEkC2jgjB9It5I+pxXBvSwgvHfGpFWQWyMjaj3eh9kRRau
uRhHngHAIaRfKAljGeOHU3gAEORssAhQRStaoVe/IYECqaWpUakV6SrOi0wiVuzKAqgZVd8k7ecs
iVHE35u33AW24luqvdj0VqNMVbifPGvtVqal80fp+eGtjzLUI7oK5iCeJL9895tDrzNvr6vi1uGi
SYglBiTVOxb6UeQhq7dZ88owasZ7/lCiiH5/A3HQck3+C71+FNvSWF8T8dt0ZAEME3ylYWkFCmKz
dSghuQgCdaRG7AXY0M89Y5RkjlHPwdNh2NgIeUi3O+SN9ZoGfIriSU5YN07rUqr6vl5wuXVEXg2W
JTgSBuYMvfwEZelFFNIIje0gCFTc4rCRk+EdeephZpBGT/Rf5o6kSNNVa4oOvkema3HoMiYQSEOs
AO0tRCZqcbSXta1RRS6oZJPBn1pB+7C+giv8jse8z3A1Ag/IYbNWv9z5BZNDMNjD3r+g/1+y6IAg
4xUmCLj1F7Tf9Du+Gio1fhxYzp0MDF0mYnqhPY3B3dPuGyzQt1Nstu5uSMdWMg8rdeniL/uGGYtC
2E9CI4b6vHI21Kb+aS7TBt6XbTcFzpL8FWRWTnN68fSOy89CUiV2p8kQD7oM38i1v4a80uef2psN
dSoxg1VKU7jMO08DqQHLMNWRV4BDQJB+Hgl7eo53NX1oX0sVkQCQoHwvXi9bomaR4zPYN4+hjC6m
fYTrpLyfynQF3bBxwZGIjoauWch+vKjqeBwEPfkFaVAGO/P7Cq075yX5+n3jOu9WKijJ051PEj8D
u4CmN4KcjctctU5d49bmKmjeA6wdg/UN4dmIQpAr2SR2hJYzzKxz8PdN4XiPyuKomFmxmmDuZGrm
PlVuauxtYjXg9O15v+ZvAJ1CXS3/Z3NN40YtJ8oURi/yJe0qYHmEv+a94QrjDljV5vC9Eq7rT5ti
rdSVXGm6I3bSbdHxBTj4Rg77Srnx43C5a1yDjyK/Pn1nOdcbgsia84SlSqqQYu5+1V2JzAqrSGWL
z6oHxb2HdaGo8FLRBPDYtiTWSXcFt/G3EQ2vN+nhmS22jwhvGVzvJ2QIXCdvWX65/ksClrDkNeZY
/fo4uvg3VZ8wg8A1sV+OR5T6d5sZRBApeGpq6E/dEIAYKQ5pWiWtFQYaGkYfn5TxOF881OmRv1fq
U3fL558mYuCgBwB27Yo/nidXz1XM3yZDXVyQDrABLinbsUciqtzvlTwo9nZApwKeurWGu/+gr+wr
vDu4rRR+TYlfIJrQwp2FmykdylwPXnK1NTT6oWJTWDXcOqHHYyVFQZjgsBZIh3ISCPq2c2SLNM3X
84zu+o/67WHI6bsqqrTdEjkAPgP4AguCUsA6iZDadtZd75WGfrxC8H5YIFE4kXH3DxTuhTxqg+G8
jGVcXYtMZdpyE5JyfPGf/H1nupXBs0I4XCF9IpisiQNlQSTbE/4zTaigViwsUTb2dzx36isCEYvo
AnSLlxvyf59GiNqS1JGrHl32ZK89AaMIt6L/ifVnl5l/DdWzGLhZAPRfhQzvkWlWi3UDAyIy7UWq
2pSAFAKDbSJZecM4aUGHtY9aG3xMCVlP2U0W7oRPnx+PKyZXGNoxksmBlEOJJaaXTcuIO8wmzPmE
k0yAfLHryXgtHoBgOZ9LPfgI7d1c7o014N4hOfBpkhcO4tZe6F2u2lAziqh77/+8Up+kTgKDBZu4
xS0Ocm5whL7VKodjE4BkdWsf4Jh9Ynu7cVNyU6Qn0X9/y6HqTQ95mu4RTHS36Nzu7PbaXpNEB6KV
6KjWgqkaybOCOM46XNrZ2ecbYBWdCjHalSuCiDRpxk/KF8R41JDavsHk2t3gnpdsHL5kRLdHfryt
UyYVoRmY48KIOSyFcRI8ppM1wKqb/520s4fr+P2R+mCLXsmphDa8OktSVYiz8EKdo/0YJLzF8SWU
/VTonM6huJAIqyn7wpO76/5NZLTcLaEISx84lwUI7jcr3unV5DYXC4w9RKgaTiN5zr61W+8sH8K8
DVHBlN3wif8yYoLheFuOaBnI6Ynd7VIf5lrTSStIhnigM3Eeghif+wf9rp+zQDBWqYH6P2H3PwW7
3hdvVD5DSAzf9H4+cq5TG+Ekw034avetsQYzeJAv05H1euFzPYlwG/C8ahCPv8pG2rA6e4OZS6uz
pCA50jAfVHsPa+QQo6t8S5hLUB4345jjmuLuU0H3z9IEOwF8O5X4cJaCHpCSsnjDITfZn6AXt5L8
6IGhFdXfVhzB/cwvVsU6Zh2P63aHe5mPgppmU4j3OBmCRAnITJmdUl70vBUVYF2L8T1iohByrAps
yELFWKIGfRcjDWzSP2xZDuV0ubUim/w7okI5QmrmZZLpcR8iPZtFSLVsxGMdwcyjjjKn5CswhHxo
zdcikFJKViOEO+xYtA+5HcmfdZQlsvmedgEXNbKUm1VDA5XrqcopxyOCMy28vMkqhDntpCIe/wG/
lyKQG8mSx3Zl6OC2Hs9TLsJW6ih2b8Bx5dA1no/9K+7x4WwV7aQeh5haIT4ixXOOJqrRdJu57/jD
EnO8R83v0/hhhsxs2iGHQ92gEPxaHTvaT8yk8saB33pQaIM66QexppidJhq5t6K9B/HlhSxC33my
RjSl/suDM5nH9lQlApB8XZ2rlYdyieTD+MVYJ0+vSwtFo/IJwFFNH16IxmfKF634JYoyh0cYkLOW
z9f8RvZgI073zqssIdY8QZDSyR/Xz+KOKyew3r0eMquyV9x4SEnl499MlYZ5jryuLSjjnDzuOTwx
eV6ayDoizAcyXZvALHjdwCxSxF8cw8oWiZkDfFvfpGrwot+FT8eFJj4P/4kh2ZbTMIYnS/qhPVZ5
WU9TNsTf73Gy8Igje9qOiNL528ea+I1BUgvzjK24xaTrW0klslA+CzSPNp8a/kRfFwt9a5+J3N4d
b12Wvu7R0JsErMlY/UKh344v421Slp6V1dZIjU9sNqILj0HItoFT/BJq5DdkvMZkyxLJyfNKGZ8l
JYNUW+hL28Vx7BiJqJULYU01fTKe9cIw7BYIjCBgBxa5YR81k4FBjs+bQOBqOdv3J3dX5Hy5lchq
flnWBYQmH3n33lfGM08MgLPQiMD4I9zG2e2zwbI0ZhPgUufbhI8rMRD22wqeSpaYQnkk+YdPAh7O
MzsYhheQBtUmXrx/+lFjsKCrWMJVsb49bI6dqdhC3eQFNLfRNgeMI3gbm1WuZn8uFZ32UPjZ+1+6
S5uxAfBxbVY/pIoaqE7hQXFnUiruWIWTCxjLCSSuFjnMNCr9R703Yy6MG7wHJK4Ag6HyasBhFnPD
otqPxJU2BDEbtzZAXP4DE+z6KgGG2yvqJH8LXG9hLA1fKK8mRat9Zf85L2cf0WIL5wXdhuW8FN4Y
i2BuWHN8OHV2Pk7PdA6OrxjA4w7LOWCbyKy5QJBJ7UAZTSKli+6nPDKkzPlgR+HOJAqu+c+Ay0qB
HyG/KRtKLzgdjJDqcIW8KYiDtiK00HmB3cIjQ96Nmx6d/LRhX/Dyrnn954VZqb7m38kNdMswbHel
/GXd3+NhULSVxUIGXx6JpVYclIWQxowHKagG3JzPGyXH2Kb0LGQypHxNx5NHJU+AZUGYcPL8pKTg
EdEu6Xait+WMl16UHhltEBANaqvQUmjLHjoJMdJWeeoH6tjo60LoVTkLERQPoOuhfm15grwP72Uk
3TvWQykLJudyhX88KcsW4ESTtKvI90/ub7fFohzUzGd8FUGrvo5KyQ0jWrmpU7GaNF4+n0zxgqSm
SMEv6go9ALh7kqxnMpr9y0+oMBIDDkfXQSJwBSSNIeosL0wKUwpJa+GpjOASCfLKcxctKET5Xykt
yzbskgiHCGYNphmUC2sdJJn9JKCghhDtTdZB1keTPsFwdA1Li43jN0ndNlvjpdVXSKpI9Z1bVSR/
wzPRqoG6ssE5wteD9UlzlCtx4NEzOZk1iTOscvbR+uOsH5VOYCqSUGpSRqWJe/+Y8N8nz4CI4bca
vKbqx3OuTH3Kd86kEqR85ooGehAWYMdSwdEV2JNN0PO8qXkD62nB3mz/S5fvWzTyvrV3RcCJgJcs
sVGRIHhWRSFRmpEOqzNQFu+vGQzI291+Uw9tmIJ7eofRS55/QRIul+/J6McHUCiff9GALR+zq+5W
MigPzkQGth+MahKFCgBTIuYAX1x5IMd2q8anX0Fd91ncJaprcRy0ThYdbMWF/dZRuRFjyHoySr92
fR7xCMxixrMPxXgdDzBYcj2TEJ1GsuNVLCD93k0zN8z9rxPUZowORlQU5q20elChEQr4dbWKb9mQ
D4nEZoCA63yRO18ZTvM8wIsssRvzH59rUo/0I0ilwK+h1eSn6v7JuVH+TwCFfilV3aiBj0HVSuHH
pYlPxIGhB4l+8/0WxcxvIMmp76rd/wfHSNp4IRP60KLLev7o90kf6N3sRWFoCO6n0mJfZFSGBKjS
QnOMFcYVRcbXAta69FP7iJEj6YjL5IOnxvCeTtYK9R+DgK5so1bwOyT3mXF0TYzP3kUUVXOoW8fl
45N8znpVbDCWAhIgER+WqztP7yEwAYo2+R0fCNS3t6YuyfYWLRQ5o1xZybRxCBHFXjMzbxP9W2Cv
Cr6lH3Qb/pdFKOTW4aoLQXsndNkfoiMtPMFOQRgUC77aG7utErNIE7843KvbFyiJPgwsx2H7Kbc0
/4hIJS49sIXThcTR+ZPRf6KNIn7XWcXWIMVJvB8Mf0Ds+FMYI9Te5Hojw9Q397KdTrEt/nRkw+nF
CpBc3aMETFBFqPnOeRJDIvS0c/kpLe38YZHY/LarS1fWscen9QIGxaGk0xpuNMGJPOwkUF4C9zd6
ziyBYzJ9izMup13pUaL7GRdHBxe3sdISc6sR9CN0zRVZdfI+dY182b4acto/o3k5Jb6EA2Geki/f
ORKHCwkMSY6YNidbvsK+ZfDJiq7YmB0/uG/zY4USumKRHEA5Kbwq16Dbx3ArZ0yRt2hqfLPGFmQo
b69h3pqnbjqzrlrutgjTFEYRYUQjIBjcoIJxTTCaN8RtWkxuNg3ux0pw2KVwa/PKJj/WdA3vkj3/
hx4Yguf+uL6cLkJ9hBUn3kgPlPCsJNhcJdoqaB1uR0uWBDBU6ziTsVIEsJcDZRjsP8EMrO3gupDY
3xfZv/+YScarM+Dd3fOfXvSpxC+2qEnbzowscSSsBGKy0IS9N657DdbyXs9rQ9EqFmm1S28473m9
z0PF98+4hAegS6lXL8MNo5sGF8Ir8QfCVVjZFU3Rp2ddO4Hxki4WuIcVLAzHRFAKrB+25SjLtlko
LLnfi0JzJjTwWDuzlogR6Bvfp7HdQMV7lAZwa0ljSm4EI1TS2SQ4KNVAy7lhUcOtCqTsEmVNbHjT
S96KOE5xvWDi07DlncF6rL64itvDHY2JRnIJInw3gBQs6S3UCxSW8Eb1guKyVwpI9q202nYk36VW
tV07CmxbIO/zlrQuS+zfEe7ji/2lqlmbgz4Id+A8008FUPDz194KLxxMsbNuOTNsI/o1hI7Pde4E
CtJKt3XYi5HnnId6BRI8gOIpyTPRo6Ww/k2eRR4iQOu9ZJrjMmrB6gKrrW7dpO+yagpUpw4JRGPn
RTRJ7uiYd+ZUpfCeWKXTgFQ0EFeg/I/MHere3WbM0ijXOtB3EcsBh8xVqOHzrn5F7uZO8GKSNGmo
wDSGYRjokt8HI8J8IO3OkjT4h3/Nvdvw+85A1tLoDVnyq+tNbR2lqwjL6CVtAgLkEpfQZz/bmrcn
73miyXno/Y4+9jordP18+0JQbhv7NFrzkoLrU38ggx37Q+QMm2nDYylPJRVVIk+X3+bKHROj7jVk
ExjOOWsO1YB16FyaFmLc9m9J4rX6zitf41dG88K0k8PYwIOBUHPVMqbV7MJ4SmGwBBfDjcNIyT3P
11BZC78NUdXMuBQqIqoTnHclaSRDpKfvBnRXSCZVOzzUDB0ZRWh6ZqYzBl5ogpQspgtFUiHxYmC2
UffvJIzoFQEkOSE4ZwU+h4wUQ4Ptv7AGfVNfYN4kvnjOJPFQnrhkpTjcGsAA882j7TcIAM1TbWKV
k68l3OuekDZ47rNUH66t4ol48WFYCajhzpE3kmsoxsCCS4Mu/o6SYZFyrxpXHbb4zFu8G96DPYNz
YcHIHgwlzzG1m35D3IlSR8tZLohRfW3GuUYC0ni44VZ2W70JmWBdQC1Sc6MYTpdrwLUvB5blDXal
dCgitxhotGOTTzrbZCVJlKH6HIyOsVbGpmS40dge3n/5It4dOna+Ukk1JY6YXDvPek64m8Xs5BfK
LGN/SaLX1tzvmcGBa/9vZhOvYqUxjUesBpgClbfJE2X2FxQE9JlSTZ53n7QRuvD1ydh573js7QJq
eKpJcMVCfZYJfjFq1EyWZEnB75J3q2D1tnxawob7LrftW74MIPK78GdkRRoIIz44U4/GwyX+mhBc
aQ+F+Erh+1o0RVA8hb4OWLzyYaG3e3WGttrMw27SV+YPLDgExansmDy204lBfoefsrbLbYX7saFu
nHuWjIIpiwVI79POyqMVzghZM4hVuDA5RAgdlbeteFZA4TGRzONRaXs78krQszC+BpKAiER//rg5
gwtqMCFVWyESipA8qCAbL4TYLPF9q/oDaXG9Y35iN9G29ndiKzctSlSM3+N7UCLogI2t9z7nalty
n9ulyefMgBUrt6KCnNCg702+Ax+oam7ejsLiLeOCcG2VE3TUMCzY0SZIUGjey+GYoQby0wKWgxcm
ZDL269IHkl6ABuoGlZDZoXnXhPSljx5KytNUXigTnlwC5r6ukIynhVo6Ck2VVo0Py4L55cin089g
QsjKbpo0yC7hRBJAyZ8G7lZXl6ySNSN0QnTgk/NbryfH9N4rH2LWaU1n8sBQWKJ8r3/wUIBEzsav
k5u6Fm3e2JOHhIQVFNQxVBEg8IhP504Qu3x/rjlaPBfqrSuqi45jz34pdZRNff9MRCsZH4dwaZyc
olQv0Ig06HAA2L6062nqn7Vnk7MZxnShTlIznS8RKCwVTso+nwqrFjeppN4aYSlX7oCKNJjUSuEJ
OTv8seKoj8ee4/q0NYYDr0emBzxVhpV7NZIglf2Oz6ot8Lxm0/aiR8XgrZZsso1s9mQ2IvT+Qy8v
k/EaG6NeAO8Xjn088xJ3dZw0CriRumT1ZyA1AIgKggaGd0Ck1MUP/lbqweSj1/J00DsAXHwoStRN
vFCC16sVtuE7nv7b/t8hkfVBGbif/D1ejp+8i6zxTAo+wnMmlu8bqAEHlTSloiLD6tJzU115xbNa
56Qy5bpR8UIk6eP+QLUEGwmGHia0xBcAcVYie4fBoUABg5aEbTdJbtSLKiIXoUTEn9QuLj0c+Xrf
i1hF/8rPxm4cTgD2xDlA0WfjqgWF9yxu2V3Hftwk7E9I4azEe3hNMeBYMwPL2sNDLcmwdK/Yx1tr
Y7trQX4NAC7c3YFNuHNXTxHaggVBOpL0W1D2cdhY9Qi4KMuSVG8VWcJql8xdK4XJkyrqFxaHxnYj
b1npKtae3dsFCQj1LLJDVycbbDzVYvxgaFmvoMrNkEtOdXJ0SL4MazHJfvcQf7hjEQUmDt3cPG6I
zHnoDwYiQvufb/WNjLXMKI7+F7lc39eIDm+SOmgx+5zXU5jN4pNIc2Y9bl50/Z0ePOSLiWJ6cVOS
DWJQjxDEV80oicoVbNwJ0eNyTStRyCaFTv67tKbxeKHzxktf5fyojx2eRU6X7iDijc59hwJUScyQ
5juqVS5UQHuOnRrtrxcp+bFyWrIkQYhJT+N+swShyAz7jKA4l1I5lGu4SoAGGCxhwUlQCycbQGeu
a7yjAQ8yQi7y8+HShZ+HTyzeBWXDKN9qdK2AA9ssIeOPqHFVB+QMKQwktR2fB70eIYBuqXoSQSd1
9Qjj0slvKLs3DDxH3lJSUsEUDnqNWcgOHk+cHi386ZwY0WovOhjt61yHFyF+M5Ug86FDUCiNzYSo
nYtWnkN0IgLBn17q0jdCPO2HXrx2A01DgZvzzWziqV2oYQKaqbNjmsUnUknOEIo167xI8PixtPLC
wxsVjYXdhoXmR1qsJmwYsknvjq9sR47FmcnvW8QEKOqgZEM7YzTRmUKBcWm3FOdkSnttata6Q4Yk
61NL3NkzOVKYOT2+pYzmEEik2TMeO1IorKZuLtzkxeCsurdoN0rWycziEsRDN7cZMOrDAruJlE/3
kU1NL+GxMatl8GNjOafLKydMg8L3HKJNCnqe7HWx8Dlps/Nb+axORS2tezzu42AlV/cU+KqznfCs
cbEK7bvEb2OauOyyNc5pHjwSjTzEHvnvZZxzmK28mEckVfm6ZuJ8moMgaHiip6bMd8bu6pcPCTnl
CYa151fhSW7ty3gRh7vLauK0YG/PUiLLjB3pxQUKH2YKB0ZaCVYmeA41kwPFer+RWYMLqk85Wg55
gEEp82ONNDGIpNHElBErUPIVjbVGEHXBa9S4QzYp2u11DnBTbpUcmdvWnOkNO09+BC/D1YmedksA
8+rmBluyXRcjq4mnD368VsVJ7V2/yz6PJE+ll2Tk8q3X+nyzQkqk1NLLYcK4S02fNPWW0RjYQ3lj
TqcVb+s1FDD4dYTezYWudoiPag1NS8mHfoEiW4rBuNX44+5OPmDc5EllLqWDs0TPdRuN7vZGCoL2
whq9pXbWuHbGfCYKyqd/hza5lLWTUrk0enGuGCXxxfvenjJyitxYkzM7VeBxG67k1jhJ50wv//2d
+ibcQvZBaPLN7GOXamuuz3wanRMqTR2Q8rP1NvQTPFM7PFo2rHry6bYO3Rs0uDnykpvaen+G4dHB
NDwKWcczVahjRUwdH0Y69RLHP48lebMQhBi687awa7p1Ev9htRpvXqFCZD+6mSGjIEKAgxQqCq35
2yzWqKGMTpvvTXkWTxdKc0mrWUO2kTe+iEm2OT1R24xXlNPM2yW6qlxigQknu5JpnKF6+EDlaKnu
gpm0zoryGXPJqk8dF54gz8QGkIfws7D7U3B2v90anC4yIXlWljkUHUV57lvpHe5Ud61kFZJ6SSxG
Z+WEuFjD0V0laiHuFdlz9riDvR1clZP4BCuYn5Bjo3yPxmQXEq9dfjtNuTM91HgP2zlgJLBmfFqD
Ms8KLwGB+G9dfAlYbGo8E6UFr0ltiArKHW1tto9h3qdQzTJC36gVpJfWZAoTKb0qzy+3t2QlYqkp
C8SFW0TUbM6ZpevueyHXi4Sdogejlz2YphDV0n0luh9jNiJp7DUae9r4fH3fsZucunAv9GGmThc1
SjcfYdIiHHsfOLZfx4pdhJOxTW3eJ09slx1/b1geCkVomA2CmIGZqZCCI305DMx5rEsh0Wefqrob
ITvYGKTjc3yxTmEZKsP3Q0fO+ZyLcyPAZ+Ij1FoTlXb3xPrN9WAyE/6TjtlBWAC3J5Jx6lGueHGq
wBy+Ybw3v1L+ARjMYn7Qa521kRa0j2i1z+hFrMatWSQH6AQmBrWr+4+s2AJyR84ZqODgNLBnPL37
3koT7Q42c/xQydtUt+mpk4xpbFVuepmFdyVrYQpppcv3oF9M0x9KiYrvk1zMmdRJWyEAV6xLAC2Y
ZSMULXYtUfU42RwZ8udAvK3ZSqLjygSk+DfgRrO6kuH7aONebNFtf0/U3N650BbInGT6llx5vh4/
Q9/DccCFBYlChQTQ1q/sGW99axP7zaQn6LlPHy5spMul23ujQwLuOAzVsSR6rYl39GCdom6VFgjT
qnVrCTVpGZiu3sQRjZZSyGduQYKM+WrSE99AaCS+2OGpgEqRiawKJ13NL+9dXg7FiOOa5TW2luwM
9sw6sIPWP1ZocLJpBhVv98lU2KySNgJqRHj0Rp+M/GdMi7TCCY/K951qq9dpAhY19brPYGF/t00X
60WjvhZphga4vkXqTF1NqMiFih0ZX4+5s+/N7lL8dUP1ZkwEPVJoPrYcA30efuWf+Z40SXJYF2mw
3TucWvAIL7QqOXX8UuQdfnBIk0rUhxpnHPmHenRs4YTNhCflDof0/c+C+LnAfrMBwmoabFidYTua
Q6G6AwGids26vEQjI8MNjNeqss5HDR54OyfUDFLMMmRZc6Y/y048zqBu4o9XtOJ5nZ1XqhcHs7t2
gwKBDJHlDSEsdlNzFjVv7JFdPnF2v79ECtGZ/6BV4DhsHv/VvEjLiS/yzyYX2yEmHvToguVHkncV
Gw6hHgqGZ0YkuX1q6h9TL6SVODV9wcjtWQUka8Y0gU40HcQfdHi/DfOClgN7VdR4Dg1hVkVRI3MF
RkZptmAC05PIh1sEi9GmZe7/6U+Y7zm4bekcouh1qcBE5RGRQHYRaOqqyTRh9QrJpF7k163wleTb
7+O9q6kWK3ZezU5oMEnoW68aBGVXrOEstsSbPU7zM7ZW6tdB5Fai3RikfbRQmSvbBtIJy6m8TCDn
dpPMLMcFVbslL1mA5QhiUYA9kKnKmU5zvxwfJFIgggWmkSczByjgU7XcGQhLxULMu27/317ow45F
5NkBSy4SUvqtCPJBAHtWTeNp6EU2VlrtxqII/k+nFJ2qUfwKzlNVrGt7eJlvgQNUJj9jfiKLjwWS
aSGWp49F5u3tnEO7DcnE7Z/a9u/kFxdYO5NYxyBMFtO5JZmAFkj93jMp4w6Gy7/g8jo4WLydbcuL
tbJfWIpeqVHxpYonW9eRXvSk5kaPmM5QLYbVc077HTadlPfF5Lqw5BDndTO4WfMSiopXUDdXdff8
CZpPdbhfnB74aQQfa6K0vofGUxqkuib0HrRErQryxMI0yBoMA6+FyPRBv1Fz22BnmQqOV9pBR9qd
PwM7sI3w5GG7xNsUgedTULW7SmCJX9Kx38e1e6fCSxLSSwpTNeI7rjATz3b3GiRLtWZMM3tRVXGq
OaxA3b9xy8Xh1w8M9lF9SFp8oYFdkAtwWVsrW0NnW++mbY7WvHk8fYPNbP92YQuxk0mML07uFmyr
L3MbAiyzTr5LLjdJljKCH+STEMrexHdHhYOXF53SNr06Mce3n1dzny6+miS3hTukYu9nHLxFC7G8
dLW0nBm6fFQ56y0EBeohfwWMMdulhFRVichfkwtHfy3s+FtVG5ORGSTDgH2Ukqxj7A0fIkFsh3bZ
KLIaXvjFSqtP2vGJCSau0kP4Wnpf0tL5reD6I6zi1PyqshcO7pVEJ9hlUUMCgnafQBlWVTFOjqHu
CfGYI/aYWb75FUN5zrWVyOkqfWuAM97eZgyU+HSVyKWODO0zj6JVccF93CikzP4w2V2od3jvvKou
DT9JFxVdcPh65ALWYlZBx3n5eTq3SKQakFLNGejy3GLXpmi9ZnSa8rpJIdbU3uai4DjoKxfQzGcq
5hnmOrhoqJE2vGG3HdQBeMb+9OzmqNcf9vyOXh7yXEcuB75KbGGpTC0oFctQY1smvJI7TahhIPfu
aFxNtEgXyFJexTqfGu7xP1wy4DQDOkwNxk1IQJdMpfhgO7vxpPcGlubVvK6/T6eihxDn9OiKpuFx
EaUPLskJ/0KC72n80xzFd5pdICZc1lgsY9widrYW+LCxRNacd9yOfBK2CunQpp5WUkXiDQpSn5qK
+KXLgfqG/zvVyX/ONnWg14tnhojP6H+HKD1R0vO/HWkAxZ2yR9nHXff6tKOu4mTviJh1yhXRNFsQ
Wa4o4THA3gqGv6j84G6iQYmuDSxB3bQzeo+cQYvyPGj9DNiXS/jBjuOwBrro/4DtNeeeqnA83jHP
u/JbQ7p8m2zJvvJtI5/kachaO1lqej2+voft9I8VbV2gmZ/4uQyGweiVkWkOLXxrvU+RYAD0n7C0
Tm9FKtHD4YaQU2ErQlH1RmgKy2fZwjAzVAq4KAzL/9lEsDN3R9vb+T5xswS+qTbuqU1QMVQIFeT6
zVFYhsoPg0zZGIlbneEuDoW5iD/wJjTIDpc3fWQYVJuSFtFckk/h12Qx4tu3iByMG2RncFTmxfr+
SmbVE1ycePhdj0Us32HTIyiLgtp5UGyilSOaKqq4recA4AZW2xqXPhoxK/V8+p9Dsu9ED1CzCcNO
JNkCgl9JhYduacrHExWfmw2TgI3nOUULQpK/efVDf4x1LgxB8L/lXU6co/o3wFpBaptrZR1zFFVU
G8nvceK80zoFWqOWhbdJEKqqdFRpw7X+wiBFSTn10zOUeFPg4oj8LNyIxAMD2wTn+fbfW5Z60d//
TCMQKyFt4cxJTQe7B4bBq6HGi6fszHeobUnqcbbIk/slUKB4EOzInsmmVfHWgrTJC3t+5K2iJ3KK
TUAu5Vs3X7k/WxlkwgYyl65QY9AzC4bV0UgBlr/bOwkrBJJmdjB9PD6eHZibKT9PPAWzFE8oayF6
sZreuQNKUeH3dbCkr4QiMZgOvTouWLUfk/vT5spLATToDeTcsEg68b92lqxLBVaNGGvARVhm3xoI
kdLA8Miq9+aXWVIg2EwPdD1qtqEa1Wak4gGZ/qzo3HfvuwpLOm25ytKJ8VmOqKkNXLC/BBGB0giI
wN/s2c8yhc+oVp9IWUKNV17nsuTESXrA6Yvr+Zoz4ZDXQQM2s1idOTCaTjQE9+DhWhrQMlgOfuvL
d+EQQNKUf3AoFxlW4xhe26GhnFLYhL8yr45nTgN4ljMYODilQ2k+qKO4JDLfaGtFoaKzZhhH7P6Y
So7MdHMl0BEtwspv7OupgWnCM8Lte4FowqSGavLFetIVpyMh7V/V7CrhGgHEq5rklbEdlWKylV42
92eB0amYmHTCMFi/RN3EyZhQfb8+7Zb0MewyFKF7xsSTRl7grMA5fUTtstfBKNqX/zAL9Ht4jxvH
Mc4EEOn3xbJPHTHM1WQcSInPDVN+3umSbEPziM4suSdKfqADTLwLWK1WY7SVg/D7GIwgkiGhDvMo
G11/9/y7mPU6T0BYwfz52uGjMvk5iH2JGiCKiqT5KSiR3yQwgw0jve2GyKLOzUYXm9r8JnO2odb/
XiUiEaLQZKuPsMqK33c9u99osegtEO3uU0bXV/K6sWTSFGSAdIYn7pI0zfEEKqfzy/CoClpARPsn
1wh7SOmdUKzGhLOuqBTBtfQcBodfNbvfhmomjUwXhnNIAo9GaTbEFKZ3sTWiXv0BRxHXj3cdftTd
EicEXp7Jgq/33xjXMu63fmBDAAzaNZrwqUxzO3P+P6vv8BvzNu98OWLQlAaCRCULBlnA1ikJOg03
dkOcOhO8+I0JOTyoeDYhsWYJVPPAiUm/LB9j9FfPv4QShO41yNZVoZuPiy+SPiVh6P4V6/bQiF1A
84NoqWxEJxdEihU3FbCbmz4jFp+7727xAvqmUSMD7e1OKCPCUsmn6T7LFlGmvf/e0RX1EcFUxHj4
GH8EnjGlSm1Uu3evdiUytNiXWTXXjvicNt/f1nuhNTz1p0lqtXtt+kx8nwO1crZP2YflNIJBtC8Y
xvBEOghJssAc89AkC67eeqGxLkUYB3SYFrqoHi9FlQqvtDp24skPP57t9JLhY9hwcKeZPJ12yRUy
mnqX/raBVDVFa+o2pJT6djRRJoZTKeb+f3scCtN5IrIyUcj4cnAAaGTziAsMMqspFyGPDavpT7H6
K64gJoax3Sgh4z6zQARAaIezBH5Deog3qozD+6al0Bv788CLU3lZ4CuVFeOqa0bV6UdjDEeceHz6
r6dUqQjhQpIqPby46YPNYlXzvO8TpP0V5jQBA50pG/c5TyFcoZCqSZXvsPQ5j81fCS8FWSEGx+lW
a1Rfw6Ev5yyymZXbtkfbpPi9qYQcbg5B9h9FJDT+tb+QqyCNMow00GNkNI+kQOl3d1tuCAAcfd7q
4/IIeUWwZujV3xCWYM+uOVfnHjVrSxXHqi0XmQDpczkYIHWB5xDSciGw7UorNDbE5P4uhjz2DcOG
7d5MEMEOlTe1EmVz/N4I5Y66mVxNh4j6lpSKMGrIOuyhZrq/BkVRY5zJWg/P62H18X2TP1ob3ADB
5hj5lvSX3Za2Ds4c7OWsrxEYjqkGNEGJWBALZ4nmpAraebE1QciczEJeCWuHb7Z3kzAEy3uEpaVG
sl2cFYZRCNZivwXICwm84v99SnG3JRldM9gUFIhtQdXn/bJKn+ov+uH9rWuaKDLX6EB7WPva8cfi
c81wGyBU91blGMjqIom70b5QyHa3L+Ru3JEX4qQoWVWYUWsXnZQa8Ni63ByLAVqLNEeyOSJ4kKRT
hTXhkog/hnEAwmkCcb4ytg1LNezqkZXjSm6onjQC1WcwoepnrFOqGN2uBKIl76nTmGrCqYJPvgeq
BxLL1KquacDSNd2EivXpCAcdZIZX7xL29qsRkdJWAJwct/vVc/WAZDMOoQuEKauzNrVUVceI1wFY
M1UuFLJcaQPaDQYs8hrNN7gM88CTQPF5kM2PE1Y3FboFhwGrxGckiltk+BonYEB3vgmJVxbJNWad
GJAtTVwjQurAZPFhKGq7UsUtuF+HIfyzBgp46uDZpo9KC0P1+Jda0PrVHyL6cv2Qj5jfq1EeDp2f
5yBjK1TxvKCyKR1BvMfJGp76F9gwyagE3hEe4XxRVhfUgz7aigDjuGdPQmZTG2R1aXL+3V/21ddV
gcJ1EwJJY30FO0qLBHdzkYzmJ8vDLdfamZ59ypYLolkQiF8wLsTo2SSZOSkjNIpBpc8Ap1WtGwQw
ClY6CoNHRC5xEDc8d672dRlyOhi00e5NhSagUtDgqD+p8a2T6PJq5d0jVa1PajRDTXrirB3XKYxM
jKxkGx7MSdk4JxcuMFAuC8aETkWDLpJHmKj+7SOSK5Bx+mdt2hWoP87RpIZroQGN+KsRhR4DCOiG
b8N+XFYS3A4aL2LHK4LHif5aIRcgAWEHUD5rZXVe0mug/Vz9wpix82JxIh3PXdA0glAHN1ttg09e
EkVPof3f36G+kDngtrzTYoHV+GT596V80bcPExLZfJljvSmiqYKy/RkSaK22HcoQZCyomkqlN16y
B6nd+K83wh3uaK5Dn+OwIfm8wCmzNj/UExnoffuleatALvBHcyc4sqmgadIV4qRnkOATHpUdvWLg
lsVfX+nAcdsMFoxmzyJjvvMq4YXAo0EbLkWXu6cc+JXfbFK8noORlhPdo5fgNn3Lu/LH14FwrpxQ
W2ez1J2X4SYPB2KCT0w7t15a2lqaT7LmJLVLAu6ieI4orK1xz2FtlQQKdOjy79nnwR6Tk7Wj6IEY
7B8HnCotzPnTbtQy36sOIvQ3E4C9o/wJNyMLlCv0uBW9SUnTcJAeHdc0tt9bSAI7MibR+L/xCJuR
YnqW3tzUM1BF1Za600DB10AJKeYqPittHN7nHA3TCz0lroJxVFlD1BcDX+xP1QrhMb8dEn+rQX+/
niNO1o5yRUz9oEv2rucrYveQ/4QT5AZN9OjFVolUPxw4mfPD+2DtSFkMsy7w7gzwv0aKsqPtQelJ
OAA/8GCZF+hXdb+MK4rkGpjybDoLNakekjK8Fq6RkTbPd4fKb6qduLl2IjLNIFno6vh1Lzl05SVF
kXgI6/A8E4CRX2GUWjL3FvvWkoDXFY31CCCkxd5mwCauU32fSTjNYmPckZ//OFOPn6my7S8mR0ct
/TUv841DaJKcJeaCFDx91REJHRJNjSWpVCsVlE9WPWUbSBsNgFjizidPPKqM5d/mL+HiBDOCupch
MU+h7qdZjnwbd0cBLmqQmqDyKXm0+A3QmTfBWCRGD1wJDFZvG1fQBSiiQKRyTJUdmdz5FLQraWO2
hHQiUkJQN5ZeVowK1Q3FQtgQLyh7XWDzqxHl9N8v9P/al3oMYhOCNIF2DUpC0Vek/icaaQrzDFYW
l6a6u6N0p+3P+oItmjf+9GCBroRkaa/MpuKcYWLsWJEMVduZZ6mbJ4dSLajbVh78GffY0UGYPFg3
rzEuV+Ay0Iykkd2NPScsVva7TZtThNshFlt1oWeUzFFZo+/5wZsiL+JnjAwrwfP2SH5JLLbW7u+X
P85kt8gpL9oImWatQX3NGjxwqWIYJPjLFPsDrgKkqHdO2y75i1DPvlYq0OtlsAUU3Kflgc5yOBBg
x9Fl1s3M+wAfv6l3Io8Pnm8KShT1TV8xTWsYvuPOh+M6MHeodFzdepWLpwsxOMlNeGoOoGes8pWz
j62oskoVqoSYsxmd/8YDVEt0OPIJeTDMItqLM/OTBw819/3f9FPjhbTsetCsMp07bmOvTlicRfrw
3V5QtsY4L1HlbYICm6jBhem4E92jxM+XkyVJ+6yrEULtNJrQ/t53dceuiDyoYxxov89lGG9aPjZn
iFEgQUlpL/pHDg+fLpt5+lN9Bn0o3lEXjIiJCNKYQtHHh0bUAgdq5YcAifwZhGwsbTwXr16Dhy0P
2UNt5/XNYLiPnnkGkNo3EOdFFg7eL0naZUaodLG3azz54OB0dUnYSgMjZgn3p/mX2Q3IYjsVwfW0
qYfsVBWZAWvNKl0+T79ytm5UqFD7DYkRbN1VKSDgzrcFP7y8OMkXYQoeC6NTn8w8tNgaJjw50PxV
myDf+H08NkbUZ1yLV5C/rWcw9Mm3By7+Y2sAHacJURmhOHeQNB6BKEmzn9t7kglsrYhnhdZQ6vCN
Q7UZ1Er2ynTIzxCYEi6FmuhXLrjPWGS7TGkpY+AWfv6CITjreDpCQ++yhNtwFrbfnJfKCJ1ZELfb
M07+vId7NAAC2CAjqs8ReG6cR6uKmJhwN0z5j5I/Hsyv74dU/0RS7oWPc6lBP+h6kc/VP+DEKKuu
BwpJvW9vBC64lATb5U2+69PUMX3FMbtJrPxXPvoHnUmdAsKhEvF4hb6Ld7kWqMVe0QYTUWcPKjx/
yw0uuuXkLJ1p0EhUQEdT5QiOjiSId1YUdM3QE5NaQtGSKcXlBOxtsMKF/gHnaurrXZ7M9Fd+DpzB
1LHbngZPueCz2LgDOlgnrGSkD0tP65+JXOCFqtcDRjgGDnQrxppHoa6y6CyExE/VdOwx/4RXbZWX
b0H+ay7YYNRxdT1HQkZWd7I+KRhTCwEe8vZxAk78o70gyzpbradI5AgHU8pmXhj5Cka1vk+MWkRO
laJARY/c/7FGlcOx7WVu6rJ3IBJD3fzEA1BnN0DsE8jEobIYAaHFITb5TFaXXHktrAE+p7PF28gR
zNhBo8cz96sW4kTgU+TVYy4sTtDSjbu7jZ3vABvmJZRXHZawdknbFB7a8CBn+JPG0x6y1rqiKi7v
miES86lXSHL7iofH0yl7nYGJ1n2gmBEYL5xPO4si0eAmSbFkmgOOKRHjJqfwJVrPihokP30hwmXZ
dM57nIvBUOOotPoS7knAhOMCDfzr49ITHxn+rJYxfxEx13wjo8qIRVlQqcONqU7TKp6weaNHNT2o
K+4YenfAj1hRbpgxDe4ifA6/OMHRdjcWY0tWRnkwk8KrckY95VQkDIRg/dtC3JAm0BT09W1wMD01
tggh0Wtp6xa4QyimKUEheLW6T+CeOaKdwYFi4J9GAy4bPQqhspe0y7guAaVdu/D0pvXQsCWQGCtn
3chVS/iCNEVGZCjXUCAXRnRxIPNAxdhawjlptwmT4+TcIvzoP8711d4SNxXOVPOu+hDhkfH3h9OZ
T/kkqgakGu2TojL8GtSKr36r1IpbpCEbK5kAqQSDHa7wi8YXD/9xaM8yqyK6RV4B0Gx2bEj0fpDl
+zBqtuXcpUEXxBgEEMWX+70O9eviU6/Yf3ly2azkHPuA5OzjHh6Q7fOwXlXpz9exaTcFoRLI7whR
/cy79goAyENbzRvwWgMHYfDI1zop+92cQYPBmOy9UBO0nR9dDuT6/O0r5ysIMFuoSX5TeNOzcaG2
AIgIazqzMXH+Wc+BOAGKQJ8+XXnG4HhEzRiypPuofJxCurGQp9R88tL1pcGQGEEfXoyOkKWqwhRL
Q6A6sETGEl8JJKkmp4qq9+BWI2NiaWKAsLdHmSxVosD4o4X1VBGRFY1fiswU0i6K3MfkBk2jCHMR
2R+X6NGsOwyWej3igA6onbmwHYVgO9xdMjF+W4u4Uq8wwtqUVioCYEuEM1qnWB0Dsie4o2P78GCI
lUm6MnpqaD7OI3cOQYMIwuzwu/3oL1MCcGeGbSk4FDAQIAdgUsFbKE1i/Gz+GA9eaf7q/Q6iNSGC
8pHWNiNoJxjytgAdtt2fnWGFZjEhncZlZ8a8udYcfS4uZJF6JL2y2paj1f5DSIr86wtLAlDbzi6i
Ir3uwaET7qRPQ7tZfJl1kx69mteKby+jCVcuetIJquyDMh+/B22l1zmof8ad5CszvXzwgY6DlPzg
q+UWL8Q3vaTeVvJ0lKqGDQrdjFr6ZwCv81O60nwLhJ8SYmx3AuCLcHTNW+bZrym5B0j/8G3cAQmS
/bsOUzyeUB4qsT756axrBpYVM22JsWCRUNUaspXixjak//GrCNer7xIDL6DmskPuoxxIiFQkbIPU
ZGpXpyn0+kniO5Yi+FoqaB3VzB3XhofbMiABWQTwGdZsL21WUyQ6vCXXDOyuDew1eh/3LRkunT3J
w6goCLI3iJaz9MoGva+18MshVaPvOV6l7yLmiP/yCMcgmrV4v/ZkXbksw6a8LvrLD/BK0xbCQpiD
gKkr3KGsMHfUEzmFktdpsFpviqGayKsHg61VsGMU27+P1uzRXZ0avqAXe7z3AWwSP9TeUhfhvIG4
3VQYUidwdOQhts/SOMC+cL/VXVQFA4C/vor4SPh+tibrLBNE3KD56a/zOJcaBAL7yLseMf5Bh2IV
Q4sz8tTbiiFvaOr7wsGrNjGAUTRVl7fRpSurgMstQ4Swt7g+C8D5WYj1rcN0YeMkcOG7tJU/31gr
WeEcDdGw6EuDga+OTintCmg3lu/EfnRfk9RgcPsG5mr7NJ5hodGzWAUa/tVD1xWQyhbdTnhU9Mab
Kz2Ei2HN6DRIkyILf76n+MERpd0ZQITZ5WT1pUZblhCZ4A5pXzumFWEalpXWwYY0mtcMwbAbt2VX
T1l21Y2BLIo44UZG00LXF7gPoPnh0DfxuGCwZOBBMAS8YiNhNsECHF6rXDoT8ZiengNi88CLoWEe
8WSLdVnfpxelbqmaAHxNoR++ilW7Wg9ptU5OWsk640oZGwxF3fb9izgsg7cRIyDCDx0I3iAj5/d9
OJClvEOAIS+gaVOWt8Tpf59ch4h7VhAK0g3Hm5867Kj0czJoggT1Cgzl5cYbs5tofMW68HfzB17J
j3k7vRbCTOjaYNNfpPNlqAE31F/VPQKoMsCKFZUeolIzZ90Byjr0hSmyWkq59PLleANf/PpGgkUD
rz+gM7oUy1bteW5q4hF2OxDXmw8XY+C1Ln/Dlm7FHCDR+ZeVm13ezpvVLb8G6/f7mK17LAHtS+Xx
O/GdpT4k2/lijvC1NcGtH3WJuhG6FoPciPEzdvjguRmVN1ENP2SuacxBfUVyUDCmWAw1TBjRjcXr
+mOzc6EMoG5RHM5WyYaApdvGIes1ddF1YmT7q+RPuTDnSl/CmiEOnERM7vFY28nAhBnKSzCD858K
6cFYdX/Refq7FGpZBKoV3gZPSDr+ivdQFhIxWk/KdjqgcO4R4Cwv3C6HLVAmGLXkAVynFydBX8Zb
IAmalvSbkQhlQQ7CHDplN6UHOdJRlNBXLeAVeSfgkuUFyRK5L41gl4dJN1ERIstnBCGkl0CiG+cC
ljaPr2vcjwx2zHKaqkOVr5NxKsvnHdNN6m3O1V1c5sQMFn8SpYgC4M8ZAfbvFrLR99OWfL8yWj7B
elYQ+vWXQS4pDkKJIK8/SK0Cw0tDUIsrskHh5Asym/sbO0DpEfTgTpAmrbgItPLpBV1Qr7+PGsnd
sL2GfRslMumqufF84kGX0duOqBJJGqMvZreqS/jPsVw1RKj+0EtaXM2KNYFQjmzp/mRN89HGLuaM
LETxVA8isSzxiEh5JA5BG6qsVTJwDsYzDoH/4BZYZM7c2rn/N2zWVnWDpqKN+jMzxvqzQmm7TFu+
6cpiTkXl4cvX+e1BHpp8sk6WhtixXSOUfBFdYsqGCtZPcPrka6qQoiZR65MkmHueFrjk0Qbgtjdv
NXWMWWe5qYoB4SmsLCkL21DQfUxePA/loLRr1D4otU38QoaOrczpgJ+MGidIxGG3XQTZ+Wb6Kepx
JroV8u/l1TQunNPi6GegfWqo/sgZtp1B0MNdPl5D1n/zpB6MSCMdHziJjmHpAwTfvqxZ0s1SLQ9J
LinKWzocVl/vFh7UQyaVqXspTNiqQkhNIKx1+80t6jV+gmJfXjoHz7dQAB9fzmgUSaZNjnbgd2CQ
l6YXRYqwa00Mke8xqnXQC5yS+iJAbTfjAjw7JEAW7FJHq/TPllgc4nG+Jd0gWoBgp15ardY3YOF6
DH0tUHoRUu4OaJqUKcEJBculoMNObmi7zH0lAMp7tbsJ+toMbJ5zuU4w2MhDJUIDQjwefAeHC9m1
x0WXqyYjtDdb7hifM/XAE4mofL1lA3GbJfjU+KGTA3Lb62gTxwysrGk16j97ybBkzktJPiGQcRB7
sF2FJ+OYNZczCJC5z38AbVjJZUl+H37ObA8rXzEJ5A64x1xvlWKSoNCTOQGKhDQ7KL/bTTP66Eur
W/BXxg3Bx0Z2tcpaVrPVcUYnl8D3KnBW7975byX8RtcioCydj5vz7O7+vT9f6TBayK4xh1cDPsQf
uSIxEfXkf8j87fHO3EwlnguUOwKaFqBAL3CoDB1OIaF3kViXY/kGAjBjuG+EK3+Y3AA38uzUKXtg
fgJYAmoOQcftMhgt0mBtRqrbmZdqSzc3M9S3qIIPXDBrtrVWkFyfWiOypmxBVBuotPKpbd83EW5J
wbh8RgtDrjstNUX0pMEPt7NtQWcf8g6iRsACkHI8kPWFrTKBvkQ/lONas0mnIgop9K5Rrpo9H5Vo
oj47/rGr5a2Rck+1kjtmkaajlt3Fcgr+whS+lLhkdfuf+nk/wVlakt2kNavoPC2UeoFX7joQVwrN
pX7edskZdQdNE8eIhxBhNgvlVUPKnTkW+2Y2+2sY1t/L9mjB8s4pQRRFGOQ4UG+cbxgRzb+Lmi8g
flJp5xteYdfDjYK2rot4kefeLk4QDWy/GGfO91HyxPlgBNx72j2Y6I2BhpxX69/SxsjjxMGhPQKS
aMSVbC+SaB9RJzvQULsBFB8l6XDnmB1kwgw2NcyDuO/orRoiMSOsR2Pi9lIOy5Ubs23/FLUvqghG
gL+1rZLRRuhspe1/E+2eUoX9vfqBkL4f+dVpSRf2YgFqW9Dne5m0A5DY6YGRvN+/yxSlpov5rhAy
Bpdd4P4z+TLlLtENdV1OTNTjdPTgyAlrJzUoyRArat7K5dW5p6RDf8Vsg+LXrLGMgtKedL0X/u1H
fQL/yYmuvut+AE6k+ruGasDI+tgZT6pXFs7tkjW/3tYwqOXH9tSs1Hn+XYvtGYMdxXjSNgNatoRl
xVT37dx0+9reidG9deHlKyXndMgBI14dj2tPwaUhQ+0/JWZ6Ui/++3Bd0FhbZil4t+6ME4TG2qY8
q/7SoW84tsQb+U3hobm7RX+Y891v2XT4OzLVM13CgCu2jhNlgQV3H/GfYg0rrttKENAR1H7uUwbH
I/d7/oR5lmSsIQ+oBbwmjYAJNaumOV9QUrE2qWBzPbijrbwql6MA5+yAdottcCF1sNK3oxLny2Pb
6gwRquEEkI9PrZRLN0qKg11UiHF7gtokBSXo5eOeOTmUnI0oMTRsIBIqvG17mB5/nlZzHjkiHUrM
figrNwrLrDDUxE0uU4QJ177LWW8jIJddn9G9QqilFAYrFnnXztxswjONt6QD88OE964NID0+7uPc
nsdqMZ0Ls4s8Z6YpMPMz/AzqOXQrErGvMzmPqkwLIRh8fWiXYjN+VlPmnkWOTIvmPUx0CxxpT3RM
1pHz42j4EPTooYbk5RJ/H/Cu1oJpTe8ijuWgizsno0MfwbU3wY7F7gNdPqwnswatw1Gvu8n18C4L
ogC71DGKQA4oEYmz3qOxysfoUijQR6VdnoAsRTT1qTrE80Lz144DDvobWEF0FoNE6PXCC6xIEJU5
V4cpJXNGE3jt0TN7BiWkaOUajCl7fwCtows+GAnFpdOHZqX5Y9/UVj+lUdxAthsNm3ug6uBFVWME
U+JE2KpQocikVaA8nivpu9fVnjIGYH9a1aEyzjQpWFDSIALeN//kYpmQe1piByeutvymogVdK6n8
ZvFRyJqo09GKYFYWNNWxUb38Z7exOuD7mOl5CzQ/EWaQQuedlrXt3pFmP1zQOYmVOfFEiGO6krIl
hMDZyPTzbx/A/SLMm1hgkUNIt2sFUrAQZ1LKCItWcW1tueHdOe5jfb0W4ZXrPX4Z9VI6RyAsuJE8
BJx8ZtdaXzaeX+Q5LYy6VKgN73uOpzVLVvhhUxK0madsR9K3Wbq1VjEjtEC66HXAv7ag5xlcNInP
IkzzmNzDctA9NgZdmyJQjmu3os8BFpbqTUinjqftULQIj8HeTKqTisRPyGuKlN3/U+JmzftvGtR/
gEVKAW+tEqtGREF0JjzpqgOrlxkRR9qEqqotpvUcghdPGveDFmBTPz27RRanoGJtOrNNMfgqMX1b
waflnPArt/2lKZxLgzYnU4gg38AAOf8Wy6eBJYX6ZG9ShY2ZENanwLO9B87UKUpqyBaF+iFzr20c
/Rc6sI+tGlmJjeLfNc15IavkG+evHPHWfUNb9YUpgphLGClB1IhgTRynCpZOz4oNkXFnaVOG9FRO
jb8LV355LLVb9MoEbXv7jwKCeIuCuU2gNjZD1+55+I2Y+O9quIra3+BOTY1blO+pjnMi09TEQZ1H
BhXOsUA8PW9dhnohhRU4YQNDP3lGP7Z4H600l8AiGMnZX/KmSZK8HmTLZweulh01fDfLhvaYLYc7
+uWYugXaNN10xMOaSuLu+/5lW8qiRjJFMbrZztir0Z/3f6pGG0UDvhrJmygi7NVh++ajY5jSrPbz
Z9bBEBnDB3uoqJox/QAs3uA+fDU8fIvbl0Mq5Sxo0/Zw4GA9n7pWdnJtb/01uuD6452OJ51Y3xAL
VsQfSSqUDxL46loW1WE3OUzXcOSJm/e9D6BlMYoBxV+k8OigzQM8QAE0JNxTiiYirevNaOPBfz9b
lf4i9mbkr+NLCleP9kHqmzFpKSSCHmLp3EZmimlCTyut7zhv9ex4CxH7NbdWc8sSa2UxibCnCWSZ
Qw718dgJCjTMV+wAZ0hVhU35s6t2zT0gs9IIQIdiDMQCOAnzC7ZmGgFBLKlp0MTiVIF1j8TxbbXa
TrVoBxfSlfGTjMcWDMN7lVnOmtCFQmeWMvdrTolg7KOu7u2EKLMfxyMPUOuRe/zHfy8dF3r0GyOj
Gn/hEEDOWgI6og2QugHQ+HzQkIAnc9zmHrTswrzGcstK0bsGN1qyESnJDMpj7QcvVr92wJZUEgJn
GuW3878IWpr9TA0yLHNiQuVpvHXLlnjDfVVKMyjm92sSOtwGCfkKOxF3Bt/erHwP/uyRX3bTo1uu
4e8Q4gZQx0kUSyPZVl6exh2TFGqpc8RgN+dZ9+M42aw1kRF4btnjRtqTDNmTZ1+7ScDpnA40i9v4
HDGUofQCC8sHaqppRq6Kc0AbkD8NvLSDnO4PU04bFuoKu4mHKRDPaghToAZ80vdfwG+eoUv0qfxW
buPcmHoAxRizzrJGs7eVw4TVuko4nx/TQCoe6PlKoJQvrgUvkXNhlheGCY8lG3BLPS1u0i/Chqd8
cvtS9jxFaBSzv1zmafj2otVTY5D9wWNWcn0mlPNWyoFru02VNlYCI25G/tOPrODi+YCXpld9hTwP
oAOF1UL/5yDciojqN3NafeN6OVXzOmyPlLWkyYOCKAxCnUf22jsygdMd/yWvePQCsfKh49vbtT2x
nVzXEoqRpDL9SQFdvVKFlePyLugAoH6QOw+/Zn/e5II2NXvvFMwjP8K6pj9D1qt6PMmVBP+L7ROO
a2Dm7AEHpicsLhvgFuNI7ZZt6SG59zkA+tF0/908+LVl0b2+CfE+ElQmvgvCg0jwosHxUjPOquys
d6Sra9irHH6La2YjgYrdAPrqamnQv3LBOH2S9Xb69mgNoNl8ZA5XACCHpxZvG9amVxYFwbrG6cBM
xHVZeumJoJJ6TsKUU/VXPg7JRduFyXjdGdbCAnECIyGfCJWZvqXqLNUgNkhK+OwOz59aqNHSQ8V9
i0Uzqbr/aGFCf0kgs1JwmnpYQED7CykfaGBf6i9s7yvsCWcEggY2iVf1mhRYucGnvrylw3vYgsrR
ngqhUv42pPW1xGCcaA3G3I2WtP22J9nP6MSpWhjsrLGncCL4BJB0+4OV0SbAnhUO/2VGDqdzrOgO
89N7eNuFJOm5t1v/veCyIm7xzwaf0omKesLvxV5s09w85gUByO8yOzsi5KhlsoWteQTGu0LfLPbb
myGBr2Loawj6YD/BtxkdAO2U0yGX/QuIe6nz42cIrcwy7dDCsw2mxFoOj+ixQYSv+mtnEYXQbSLp
tfoMFySB1+b28Gh2xZ3e82ikpwLVVps9GH181gMK4oIBvYGHhZLGcuoJghf3n7fylckS/MbriGzF
kH98LLNCZA56Wa3mKdQfVmMtIoTBo6MS8ZpAmOfdOTHOuCYFDwY+VINuc5lMjEIMEWSi5ALiXrDu
qftwkeSRI6TVN6pRAKhCvv/2fGCZfaHA2r4T6Km5JIilPl/P4HGR4aP1x0BdXBor0uZ8Mdc/S0xr
E/smiSUy68Gg8p4sEWIAWuQscdZ4Acex7NLXhc//1d36uD5il2KzsktBxSH4aVpDwU6r7Hovq/0H
N3uX8dDnILQmA2ipLees4SzG8uMZqVDIyP+5pVqQ3LiukAGWk9bPrDq0FhtqGML15yJGBlnXViBN
8im+v6/tQKYwMnQ7c473x48hs0M+9nvIEB4okwu/j5gR82suKlJ1OZHZNp4YSAHOqX6WPEe8LfJh
jForaAMbVDugV3g2fJ96QsjA4+/9JdWpIRZZzeSPB1cH4nl507yVGIu9f73/x0pzSrKjSMO1HUtX
iqbnbPOJBYeeaREZmVLnVcXGRwaXahqpMPPLaTaFop8khU3+Ij7V+FJvupvKtNvJrTtnJ7w/A473
RTO6q9h8aGouSprIWCGP5qR0Ua4d0JhUTbuKHXvGaf1ZerNa8UITg/OJrBWUrwOuvolgD+CjPgzx
p6jVBgZPXFlNaJrXQBhIGeJ/qlbpST7/KLJFq9sHR4Gpw0Rw1XDVrxX01tJNeCg0p4yN1olKjxwX
IW4gUzwy2NKUoLHNgmATN5Zq0m1bdQ/Y5vGH9HPAnsPAT/sZpVMvjx5KiZalTsNGtoYWGcpQHELW
y9zmuKQ0+annb+mJwg23G+EX2atn4/rqy5hRrrAMk9GDoG+9zFNX8KJF9pwATFsH8P4GNVum2yec
FVUPZ33Cmcx9XQBU+e8K0zOQ8bMlOmypWxPuH9vNVIKSNA5ZQkE+Oe6Y0RZD+u5u2idkC7Q+qL7V
BMtMvUCqr4H8dspAvnkmFW8arpNmTmmd6xJvjhU+OKB9/u+qzlEYSckrKguH+a2yYa3rtpAkgS9R
t24aEDq+dq1Wq/Cg1hrmlTSSKgwSAtUJUVld7wcoPDwHSbO08diqiDs/1IEw19BxaF0wSs7EfZh0
1EpNrqoBdydYBkaOBH9oLJShiN/CEXytW+5FIzhtAr1oxbMMo1r6k5D1xbQZCywvFMW7PhbOqK5J
nbh6TogsfEIS/yQPVB9Z7ET8gEyMWkGJl+mbhMyM1bCZ1MMKWrQblVvronxRzrwK7psv8MbByQGL
+yKyk/r5TccKaRCx0sxDzsbXsnAsEePWsg2hKyoMRy4zFZ0hCQUpHKsGRyV54b7zEw6k0WSH5Onn
Qn58M2Sa3O6MgbNfRxzVSDuu5TqgHTAK2PJKVKWbMTSLvyKTKcDO2NBglnifgQHKpM69++NTF4Ta
L/QJ8AzFHlpt2J2qLaZ7G+6P1eykCJqurQGjB4arx1EkFptdm0R6/gQIMLAZ0fEBy3QDYvzPI4rh
2eZsOZjkoaHuSpT18ZC7fNIApS5z5DjiaFVA27RQ15F35HxTuFLuWGqaxcEnVhL6O7DFIn1oFtMy
PV0/uCzUXGWfNF1Wfs8NkSygaDf5WEFOgHJjxiyYhvVqHW12dQdoM1V3LVSfjQ/PALAcFdG+p4s2
xZbWbP2tF7+i5bH9gXOhnHj43v7HcvDI+DMaP15EkaOMXrVRR4veNRPX+/Gm4r2/GF0uJfy5qKCu
gZP5iQ4KRIVbSFXTZpJdX3r216KktDhiX7Y0LEhpm+UzwldHMw0OI4DAtG+goHP6dLliSCgqmRGt
SoOAH/1/yYjz/CZGCyZVf99wQfeKkOUjZRs7bbjbh1C0gLiAZgIL4QWowabwhvGXl0V7didZsgDi
7DEWAAf+2t5le7I/b2eJW4YbdGW7bhR92FrlzToTqQxCTafQMuuAN3sqZwXeQ+QLk0t5p+keXBzy
KzbDxoFx8JVrCKhXs3cuJXgPbgZVFmkfa5gvx8rh4FavU39wUX8jbrsaRV6IPKkMj+LdiNOibyoH
RSsMhuB38Tgv7/cA6sDNiPXsQtDWJbw0j7lKqfUI0VEARv1ELZZOPmcS11Lj595tzFEhix248XyD
UvUUFcbOV5ZEEOJ2GfotC+NcOgd4lQz2UYcTAqKKJt8W+bFB/j2IiELkGcKAnvEuGD5anKTSRHAo
62RSyNUM0ac8iw0wer7Oo+chZJGmgbqpo3Ek9t5Ze1x2r5+qtemICswYz9R/X7ETan5fatQ1JhrR
MXg1w8MbQNJc25RhCQaR6yPX/I2yD7/Obbf8J3Ab1rCLncn0brW3Zh0eCxicKaLv4aPBNU1ZJxw6
pes98DFojU8+eey+9RLm1FtVYfm44WZy5QW3BXdi9OZdz0/2E/N6LqPbIMPO0OelQdYUmOTw2k2e
pyhHvGIl4MrFQ12qKErZeuBx6X323ftb/Cc/shFS7AJIBNqFwMCP2udTOxYKZgjpyEF56d5iVrQo
AG/syXAKlmAL3Un1IHnuzzscieJIFrDPWrwEiZ402QlobLI/qEvKNcl9ubHB2a9e1eSmUCJZQ8ha
6TaRkcHeNMgtK0nkgScFFaONxYD3tX1njw0YYh2kqI2sLI18vI6PR6xQv+F3LdEXk7Co5HBbK+jO
mApHSqYTcvGAh59lvzDPYAuJmdUdilHstTvZlxnD1DsM5ow14mb8pHzyclSCTfilUgpAexEPAbOg
4QtUgX97sufzKKc1fOiLitJfMI4AKfX8z57VhbHey0q9y0BNkuHorv6h8N/mmqArnRXjLlKovhDR
SLbgdVZsmC/NBRqrvnFmd0QtMkc1TtF7oJCMz4iB/pqVO9LUgK0Va+B3F485UiJLmeubo4j+5MAt
0E2Bp4gM+d+2+fqkRW65PTuWSSJ3xJa7VQADRUfu0Kkueg29pGXM6EiaLQD3paded/d6FDHNRz5N
RgHTwS15hNEgvpplR0BssWujJV77ItayfFmU/C/tSp9M7U+8esTZPzF+498sQLnVeOG+TDs0WqET
UTotmF4RIO2ohRus6OzhPh+B0p5tHLBPtXXqKpaPIqE2UICWrn3c4aI98IA6uVRTWPaGnHxAY/8f
5eCne2bdOc94f3RCKDLgBqWe+e8QTt0ebEuNtktTJoxnIFz10+hIS63q3uhKuHm6D779bNT1cvGX
MEBsO5caSn4xh+WcUsZf0TCoXL1TAoGn/r4Za5eZlTag+e1TrZk1tyyYWlwTipWQz56lUX5KAQ3Q
2FZhPkU8qbeQZrqfJZP9qfIWGDdFjCv7bVfzVUBHRZx2IsyPY+evFPkui29GHqhpXvgqCzsP4aHb
mUD15tzolojy2tp674gm2n3VeEYEljgNXpdF0jIw4UXtVKRobQ5RIa6qmHJ4kkFsQ5QIvzgcjmph
V7GsqUKJGvTAqOh+XDOXe979v7hlKfBkUQmFpR6tYp/d5yFs/CAtKPAgLyLTzuiqAbVbv1A75sNZ
U6pggFuKUBnk4Vg1DlTq9/P5584ie9kOAP280FlC0IiIrNpwFj/TnQ8TIXhjOSQOohahsMQ/mGdY
2m3BWCAhMOImz+A91OciL6ZyMCzb3/MGwTaEyZ8kcV4dpumw7YyASJM+Gw5XDBfrh4+bzpjScgRT
fWFVUytjJN8qbwSrqxcFZ+JFySeImaw2FSqhBOENcNl5j87EpN/jhRFbNp+F/78tZmOXb2CzZBmD
J5FVZNrOrvtASdicl/+knamfJVgHtUA18Uf9O9DYRI1sz3Z7eYOQ06KjXMgGXZL8ZPspPkyg8LWV
D4wshAujquTqT2/tXh91LimjAQg2XG+q7V7W/7BBWRSptS8wrpfrNlw8zRnxd4SSjE7ZuhsM1aKt
yQZnmgThO22ubGr0rpG1FJ4oUy2LwwT8hrjH6FXMErCP5NOniSH5ORe4ZtGrn3sl2H8MT/a8e+hP
fYIuccMqXTvYfjj8Bqkn8Aw03NOi5EEpS6A3wMYLZFURs3CWZUp3owN8g+WxuwkDqgIsSeb8EhZt
l0ZtHmETSDkaA0nxLWnRhY1exKDZAH9IRZsoJ5VJcHTuYVkm1yNVTFKNVpkQw6VzX89TDbci843f
oh0GkqJZfn4rpQKmb9IWYg6bmsXwcAew6ongQUe12ni3hNSMrwCXtFDgeMAqdGD7B7LZk7G2ua/B
EHn+fGnWHjZv7iSPxQYNQaDnJeanIi/OrU5Vpp0GLi2sYBgpdHQ5mJzFLP/1aquJaCJ8uBqy9kpU
2QtSWp3S16Q5smlG4ibvBPGZRQAnBGza8J6gAB8n5/3jSd6k7reInwV/UqmGHVmqE7mfOd0KzJsl
2bVdjJle0AEknyI8eGkMnYsKqMM3c+uJy8S40qsID3IC56Cm5PgIwxbR9KXY+7Zrpt8M9aKgqRyp
iBjou+ju0EwIK330pV6oMU1UyE2D7yOgsBy7e/iayJbbQMrhwSZmrMa1rokIiO+Xsy+ITJvBZswO
JOWuc9g8DlU+1ExlfcmiOiad2C57L4vsME9peufV6XTSKPf86LY7lW14LHu9lhNoXESyHbSDGITy
e6vtRr8dran04tpZYJo4/QiIlTti5y8eVSq+wPJZvBlYluTxpHgq6CEaQSKnJfj8ZjgBgoI6eUuD
VWgegTlmiyA8cei6Dk+lfUT1pyIxu1q1vHviOTXbw9uX5nPhfILfJnhZMhIiDW1I6qCUbKoBXSAi
5bDGTvikkEWjMmy+QeibPktEP6gyOpNE5+13bMoUanSb6kUMZ95BAoY8cbJnIzLg3nUwJdtHYSoW
NJiRSH0BThTqwyIqX8trAfajK4D8RWly2A7G5gWbXiEULhU7NKEKUskVIR4+V3KNCE70+jkRXvxf
fXnhZ+DxtBKI2syrt4vZbG9gwEmKfqWM/zC4GU7+UjfiXRuJH7Ejal2z6SUgJPdGW8PcLGvh90pU
dTS3+NvZTp3SpiDX+a6b3lBU6vv3AxJ+7g6EzLixr0ouhYPd9SXFoeplDbDdivegcoAebbdXs8lp
oRoxiNcQpi56FAN9V2qTDe1wBVqrPmeP/FnvrRNIbPvF0Mz1ZMEGGfgdf4jw613do8OEM+MlHIXY
qI4lA7D075uOeu1mgEn31F8f7EYb9zjs/AjBp8alYjoJzMQcQUSDQJXDrJy/I9dIkSCL9TnNaaCK
icxJss7w1GaJesvHetr2B+fbE6XdA8ggM1t46KOVq4UGLYvdxVprNkp+U8DLQ/cUBtEgzNJ7J8Pm
mqf/Tu6q8ZI1CVtdrwQ8sQc5YO/usQwNOAr8yh6J2nPP4NqGXryFCYx7pgeA4YWUrfbbJ1iZInFF
Ln5urx4SVkgRojtqu7iQGsylast3mrDdlboW7qOfSctLN2Mx3U0q2UmRcppc37hvf05VQx5VC5cI
8eUikDkEVlvXn/b//tHHe1NRgO5XP/8KJTbfNPJgL4dI2adeTbOMnj4+ftSauWx/k3GmznmQ3/TK
r67sRwyD8isM3ZyjNeCAUD+m9M5Zf0M/Y4IvHbW9022QDXzG3qAlK4Lb9TqdqH12Y82qDABtC6Ze
D/KLaSXNcTmhikBwyHEAuiRvfPo+7REqv93hAy6ChYIXxHAbGWc2cGowgg5nIldS9zsO8jpPbxyu
8bLo7Bb+N5o5KjRRTmNVEtdgctbPF1Qlby8gf654sPamUxlK5ELLdMqdvV6K4umdDNF5UmrlGviH
wm6f7RPP13Mt2Bpq3dkNQAreRiMoMLg6cFNCEmEUpiDt6Er3Y2+XN33JG2/UO/ibciZiJRfzXaBM
rcHMqCJEnnFurjNSRa8QSZPAWogzq/htfYbkpT0vXNoUOnSdr0faIZ9nCU9fYdVKrT97A4Z76cm3
2m9GqYZQ/M0/NbXVNy7MBjvxaofyUY5Krgs9xhdFKpSRHOmXt6mujOvxI3JluYhQccwx2vEQfIsf
nB4DfTT5KkJFxmcmRm5rjHL7U6uDrHfgHbW23iHNbhCfKGpRL9+8VzS6RQXsi7ma302SnWFIXIV4
BVCZe2/xFxsKAmmYM/cJtEiaYuzJYtD5lBHyClFwWzAQadi1yyN3S6NSzVkyjhwDHU6hrduGQ0U1
0OVJWQz+vqOPNZhFjNrUxICbU+lS/7gjmZO9UNJKJ95R4O8dUZPHZ7dNZMyLnoPDhjQ8aB8FtnBA
kR5kmMNBlJxdfoyg5wqxyfQI2/EcvcJbTmzG07Yxtl3cjIUnrHYsFIOgsZP8V3/EZZu509NQjpCS
eC8OeyAppRHB0Dj+JaVvw7wrLs4I7EYjTl8NwNQlH8X2uopxFgqaDq4OjqjMruPWQYk9PRW2CH1D
H8nyTflCaMroD5uMUkWGy7bRoX0pYC8QaCPOsfNjNKSyhs4FDi5UyC5v/ItR+CB7oRxpA/3h7yDA
uen2xuzqITxgTs71qEBSrFqXGOxKaBR6s9ePG/Buyg78ZaZPWqXFYYAP0o6MXQJCoumNqy6L45ZV
GeRv0OqRqGZ2JFSxrJeD8Zn5Js0kH3MhyDjm9/CgXc44JNxv9J14Z/GB8oQJLdDVYbDM9JyRBhbO
TY8rLIL+8YI+iQScbyLvIEOlQ2BZEIfH8G2qfPzdFmdJUU4G0yL9kJi4z8zzgnbnuelT7DUQkpIN
sjfdRNMPRvQr7qmf3nulzCMm3I7wuqlbHQY5EektG0Nfq1Dm1CTcx0A6kiJYQvuk+bj3kkz1SWgm
xUre07C1I+uQDSvnl6BAdmjalPVzfmT9JJsPkm05X4IAomkJec2ya8NfpcUAEKOwJuoqmzPxIWYL
Yuo8sB2OZE/4/SsbCaeG+hh+x4mHqDTDQatxHKyiWpTkGM9v8aKwVQqakVbIpLaumo/qXYBSSBN7
pkgUX1V4yUOX3fssxIRQi7X6QAar7N83AsSekVrfHA/y/krjRNKfVE0re+CPP/XcCAjSe7eJ6Rhf
M8btwmMr1IVJhcUS9Xdwua7MXDKECc803+xPFb+m9eDkCYJpDTw4kfdlup4erpI1ZgoKYrRf4E6g
WS7gPBYWH7RSLkTYn64FuizuxXIB+qztonttCyVL5Z9K6H1vVAik+O3e+bPCTRjPVnX5vPqlXSFh
c2C/mDQV2GOxIFswizhck+jvUmG3pDVfGb/y+EVKdpArxYXRMHjFKcgtcF0Fc9SABw2sBYTgFblT
NFSyM2bhz2AFRmsjKPiiiuctE+iM2X4o130cL2rQ9gavAIpYUZEX9YNqgSUMCkYvD2l0UaJKqCEO
HBis++bHceWhi/d3N/EYN71e0pKJn9e0Dlgx+DEfxK4ic9zBLhCA5ItGqfNjcwrkwLlD1hUFur4W
W4D96gK86phypk7ImLKYllJfe2kx/H3/J0e9ih2M7YC3zyOpqukG9K/kyNfGBB1diF/YgT/m9OrV
p0/TlCzQ5ARF2n8kBNHO6nKak04dpyyweCPpqk9hlXh0HqmGDrJjpZPYf0IZFXMK1RAubMmsLvRs
DsvikjKR10MD46RmkiaVQ7Xujfzroe5XWdqXt9jUtLhkLS+E6k3qyC02SBvOLAaNLhUn9uIt7/1O
RYBjSwR18L36G7MG6HYrCwBYtO81fZQwHq4IYjcVbqiuWjpqWfTGUdC0u1mkbNlXJiDiqMKz5J9Z
eANt8XZZyqvSU4WExBdPnoBufVb0407H0PCJjJypswqb8o5Ii1Nb84pkOScRFvlfeLUTHESXiApn
q6Iw+Z1+EJdJ4+r+H8fxP5Rignt3g/N7eUKkZ86sSVZZO055K5kbgiCNGHjBX2L342ROQw4ty2WY
acd8WeN2v7B+r+h7BVRislva2OyZOiqlekLHJ7LAxXs5z+RLyOhoxveUFFuTdlzuCvq6gRNSe/GT
i/H/jE5tnI33nQZ56Vy7bgif6KyJVbvXhypmuUN0Oe1/wjaZ3UJkgMcfnNlhAGj3HRmMP3YCWtCl
nNNuTZJXxdePYPPzSO7lWcDCxpBpJ4aY4w3r/CBDkMePg8V4TB46hEUaSru+YMVrlnly9rJ1AQuY
KgFDV/9RemJnr0qENHnwxQGHN4EEVeLLQKWyfluGlKOshex7v8+o+bQHw0b9vcaKa0GEpdFuLMsa
I+Qrag14PWaSn+FNSvj75py89q1XcCvAGUf5j8JT3V0doyrJwydMZBVP/WiEh+TVP0uFbuGunc3T
UxI3NfRPWcK8FUv7jEeK+Qv7sXVgt+MTV7PRYIaHVQYcfG1kODv5tKk+acD/azoVKmJ8wgbynC1s
P633FbkQX/Q2L5+dQySGCOIRrT9nrugkGxABOzK4+4VYNMmDuaMx9VyF/7Fg9lxBE4xWLn05UzlA
1Aax592sgnbz7uJjmbAOyHkO8lfkNIOI20DIQHe2O5rV/vfZ8Z7a3LbQvQ1bgwokKt0GvcsJ4JoK
iKlVffX6STczXJkXd3di4a24asuuCfUnL7sDdobmYzqX/7jrKtVWBvcfiCigMu37ew1P7TbPiIX4
e/414D6nqqTzfhXBB8l6p3bF3JhqJVF0K+yJltO+fNA5H0C6zQyfIs8CbZNvU/RoJOY8126ZMA39
E72mzGJvehNAO2zAVvIFPukxYUruHrmmd50KLwIAiq9W3JEz5BM/TnThA+J/7wUOpF2y79VP38XU
syBPO8PW1Tz/YHEIrSlHU6AFpAuKZ81Aks2F5fuEr5EhhA/xyLDY4vqB0ieIVLdbXEJd/4Oj+yU1
M9AGq3MIJfOLDzWIueCvkV2CxbxHt9XLJL7uUdzcEmnPRUKrCfT4o8j/OzsBdJ3G0K/HxtINhUEa
0tfaidWy/+pd8Sm/wdsrDVL9WdHAGHaK/Tb2OMR8pxbnz20wWQrZJldDta9heyWARGx0Et2A9Zxv
+GO0kRjR/+IpkGP6OuGxrEUl3cWRDYsCRJtHG1Es9IBTPT18FrEApHd5HwfWy//KMHJl/nuGgMtF
bogjx4EDIouRgcMdE2MSUVt/Zr803QA5A++hGh6orrUxpCrBntStrl9SPpJ4uQY1MJKsbBP6fK+D
CqT+niNctSwtKZ1YJwRJYDF2AVdCJlQK3XK2dn2i4FOiYtmRTtqE9QQctvG9KAVRNMA6AkksILQ+
vsNTzF4M7kTd26Z/Fqt5UzpsW4Dp8MsxpIIB5dSzpkzfd0+Xh6j1APZ4CloAeVG28llZcxn4ZMCD
D4jQoq6MrRwi6uT7j+fgWtH/14vFBZvqnqx2an4wlB6ke/FmFo7L9gF//LQZZNf226Qdn3EO/HXT
jA5xiS2/8c1NMu0f0tZpyujr2UN33EcDDYyWa8Kd3bPL8zWcEMSvIj5XMDi1ScDPAjVASM6PELD9
FWQKSDFQwBDQNvmL1q1Ds4q2XXEAHiHHp4X10DcsBLYX3NEP05g5q4FowbZePWImFDopt+unjuFy
rslfmhxOp09vxmusJHSOCu3bwOQtjk1fl9JItNdotkUXmGXSaQ8yIL8FLnbWOj7dMhUh03MfbHSI
uxvq+2d1S/lmbeuKk7CFvY6PKjKGbeNPi+smSiB5JfRGqtrAheAVYQnjabCfLpjTFRUEVvKPkk0w
8bRJ4WA7N0cZqkf9kjI+uKA7usziVmRVnnxwmiNMQcfeM1UQIPmF4/1MZAo7/Gx5gttlsvocn+ef
A2nzzscssn6u8FcY72itz1zD24ZGFitl9JMhP0fasc1bo8ebDKNnx1qZbIGkipVR1uYUxTxc5roM
qcbVMr/rSOAfp7c7C0fOjj7Lqwt0OYIXufjq3IAbltszNIA0vRbatVde6nZzKgZEmSo3tZFYtMiN
PX6pMAmxS/Rc7P8yYbPWMAceK3wB8/5jK4HRFlvV7C4e6y36k+43OMaVvLwknojnmeh53slhYY5k
ucg4cp7iImkPUGEEHyMP2eLWBm7F+SdUJjRz9wlxa1y7P0ORwcqr/G6ShHUF+wSyHc16+Uy8+qU2
BTbmM5fX6Q8HE5qJdLP/Hq74LmfkHYWX7IA1XrXN3WjP3GGV0E/WSdSFsD05QADo/WJaOL5o/6PA
rZQHQ2I2fWKw/0BfC+guEFW8Zt72s6krWHi6KEfhjy+2Hkr1kTxVAA5Uf2kjHKAyXbPRNbwmr1Zc
ox0P7iu26D5s7EcF13p+TuE9iYksaSIZ3chYMEbuv9FCmPOgmf8q47woVAeO+/26uOPhD1Q0iFDR
vRFRkyXFyE4IbyYpa17ljo4OtZuVSY9X7c4UStF5TayvecHPsQ1BMZDV7c0ytjRHzbchHpXFzZ1F
cuBz+g00A+MsIpX/sS+zE+4KMFvtdXT3OhwjJG037MFxvZTkjF2fEG5G+0VPxY33fuSlM7D+GS8p
z2dkkk9KCkNWvbCOdtbyHy0f2Rq2zHNZ0Zy2SCvRKWbAHDewgRoslaq+vG1xvWL4lWHJJ0bkSdF/
lcyOZndOBwwlKPAgZamyeferJFY+tT19ByaXjnFag3mDJvhUSLcGrMB0YP9LkbLqm88T137UJsb6
7dglnnwLLMt2VwsLo4nx7ssjE1MEzBqbiVEfh0K9kJrlSqnGs7/2q/XQPi8/E+CVHNdnZMaonRN/
qfQx3BKqzGOtxOgnQFr7vwbaTELqlCXSDKhuWApElZLzw3irxMpxGFLUkJ35T/RcNpUfX2Tw4HoC
OzMs8r9tdozZf2pPk3g/cDxIvO6Ep4syKHvXZ05DeWVT7UbWkbqerUqcp4uG1Qop9bDYArcHsaKa
wcgrgbpjrzZ+OzAugPIkm9kmr0Pqmae6f5aRL4BUAnpdMeHqTIoZcgiHphhmEGHp7/xldYqW1pbR
6GVbXJs31q0BwyPRJNdXvBS5kyhgF/y93hpGKcU/HxuW3DUP6PCtRCMVuWQFmuSBJwJvzU2fk+sn
gH6v8AY9EtV01l4RLH+S/uV+4FFt/ybhTFAXoJyWS5fUVwFtlQI/I/WfIScyZ/GEGAjICtL57vKX
Xfmjsy//5ZfKVuauTRYYVo0OATcxfiXJYgPCo6vR0WVCEVVuLBU/I4rSbf2KHEU+0RbVCpdgLKeV
FrQBR3cKj+cGAYX0uQoOLZP/oLDsyxysQMm9bdHsejYOFwepzEaBEV6dElp53LFLDiLFgX3SSXMc
6FgyWjRqz/h5v6WbZRGd8S4CZ6Cdtx3iB6og7pMfj8MxWsFMB5M6q2+V6zrQUCM584/ctVrdEu7W
ifGJfdqewXvA5AIvTFaAqRSnr9kc1OLtziQo77dINzNDWVkUMmdVvzladHJjkZvMpRhEzrcp6aNg
mfDk5piAmnOKbShPL65fvxOw0yNnLQarQyBv1ey3Z6zxyR0ulwuWMlE0Fx0x0BBPd9gCPVdQTh2D
ui5Q/2+mA+b0jfEZf44ou3NDYjcCwNLe0uhZ12sMMSlA0ZdQ8Tox/Et803kqESwizUS0OcSjJtf0
/2DWUHk6ZyeefM0pZKu3ZsD9BerJh2Z6tpaKWcz23or59/mZrxFTpAMqLczGklm3hI06FdtnCOVY
KROEQC98f2qgF0r65fkocEXqA5DnKFqFXLd04jfseYv7hUXsXFffjSq0dtBLXnnNZZCGozxfrHnQ
7ScScwURJNnvhxZ1xD+sGNTmyML09I2VJaQWdAEJdgEONLvRNyD9bfuFmQiV+42x+zXzgjmAEg1J
GlVYLQ4wl39jvhTNf3WtWP9NaJfqTkr/fYRkOwc6GGdz3OKdB8XjAKhKUou4dFX9vwbAdH8/l1aC
FLTSYILDOMwdvhUQON8bA37gnzH5ApN2C0mqitjnNKVFYie3qC8tTbrZ4bjjV4oydUWsL9YEMJjx
+dgPTB7dPvKxEI4xd5kZC/BXWkJy3lrN9VZuilBrfaPN9TmSaWiugnuvGbXs4rNHTlMv4oT8RbR3
21gwl+CfgUF3g1vH0VQPL2TzNDxG/38gNyBRVnsMWlSSCKhE+wr2ba8RimFZJirNIwuyRbyzXQ6s
5SfiQVgGXK3oTZEjwb0Kh/uDrp/sCXl8AkaibRkuLQfWIUNOxVybcEVmbuAk6VMK23GprrgqIx/0
KU6rKYWsmZEO2OwZ7juKjAOROr+bUWJ3nrLUF0DAXzD8KLELFhazo0jwQ5TLQp2OGlQiASUUNvpQ
kzPSTfnUAcZPw5bYjlosVkzECFUnOSMy4iu9yica+lax6VnbVEbvXkxHjDTl9vlwwS6r70yVJe0x
GHoC1yoDD/+6Xs/u7t/sIGjq2WtbXE248h8I1RnzkSIwERA5UN1wNg7Lwkk0HaHf/iI+LWZmZj9C
AlRRMwlqJKnK41wt+MYHr01QA65F59yDhQQEHiAqdU7FVx03PSPtJ9VTuE08VAL7w5k/bVSZ3kWA
6KaTL6HQHgzB68iSBC1zaNjptvEkdeDJJQBwcQ+NBV004KpmPSz/kdphmRs82AWQCgAd7kp+yVqV
lSaw9mh0g/BC0vppcEdCL2t/zK0TPYWkbh6LMImIf9nKZYhAqU86yZCieOa1HM5Qkrih9HXT73h8
RoNKslMD4OVn8pDnlXlqYxFXQX6xHuaQI3sDIK82zeFO1oXyyAtXDRuSLWdg/OmFota1HRIh46hI
bDF/VhwmTdqiR0/JrQJ38O1p0vBeXKPWLZNrPeQZPolRgGiQ5HJLvHLepmPf0zB9G8NJjNh06lTY
ksT5oShH7OTk+a9K5kwBX/pBKFzWl8daEw4IyTmaFD3KparrNU1FfzcGy1Le5lxpmuAcAKOk/LIZ
8Cel2KNx9SuayhaaWGZ70YG5zBiWDPIvEObReJIJVofd4OfDGf3zEO3FHdf1UuVfl43bfdDpxB3n
SNN3sNPreDecz6oL1pniOZKdVvC/jXiorQY2ErnX6/zINM6ywn9ArPnLbU3mGYbvRyC8GGXLWa3C
0R/bAv1m5oqNLBz31B/5eNOvwMH0wOUmh5qIR0GTdphtDlVI5NVAWOpHwwvTvks7VHcTx++A9G2M
wdqIuJ4revimvLGPnz2RgUdewa/mpNE+37hjOH+HXiaVAMcAxV6GoQQK5PeJLnnoEioYxIjM7ln5
IkFpAfCP7pJatWZ00meJ8EPDurG1niisA3NqbWO0EFMr0eQaV62hKiP8DGRJel2R3yz+x5K4bjNS
L0aCb67V9IxUqa5p/1FDKp3uTaVnilVPwuQheJPHEA/HWBUP3j+cCAh7ajvm5oVzTfLNld5g1HPx
oTU+j2j4qtZDrNZ0MiqzA98MG/lTFm/FK3mKY5ID+Vu8psF5kkGEMF4WnLIqNCo8Rszf1SH0KTr1
DL/I4/v5gwMh09XwAsctTML7Fg498MzsjCPaD3uGOUzfXdhNuWQHreTa/jZPNhKL8HhGatQ1LFFg
YEUbDy3bP9eAFUx/L4vIyRHGwi3Cqws6PUmF3aFOi+vpGp90/K0ppGbAQ+HXU34mv3yp4ASvh+8X
gWkuM2U/kfOIWkGUiXfIDsP2UlML43siHcMb5gs1sPyz0tRU9K34IFBTvm1CQs9ybvUAeTWU9wvr
F17dcL+cpOWIAJ1fPjbr6y9R/yEb/yzRJQIX9AQi+rBP7XQPzXFDQpOAyZlQBW0AfdlPgYNGgCWu
XG+1BL/pWW9/UVG5wFlJ06J26ZOlD6mGFQnvaNDV/cNi2SlACimbFHhMfkzZ5meUy2T40B2jH8jQ
77NRj+X7pef7H0WJYRqUtoQLvqa6ZoZoTwrz5lGxXFw9SiehA/agAtYTvyihlc5H3x55bIsCojib
r7jxt/WKNOmu8mQPfTaBS8XHqGVNYJBiwYTdei91fisw7NQWJO4pL9qYCuVXw6Rg7/Zyyp1EuOwT
UZE4PgWuHyBdngIaStqJ/dIaI2o8sxpDF6VCBPZqG9PrBEi+W7MKj4IDBamjWPZ0FGjMLMyaX/dQ
IlLS5gYmsMeu987es28md2/DK/jD+h17NuFN1lDSz9mEBBjT41yFwTUWb63idwxFdE2WGOmJE9IJ
vH8JJ4lgrsvjiM9klrAv6lq+vvlF8pxd4XpKsH6ow3F6UzsXeLtd3J4cfqLtHDhkLtHl/DrHkfEm
YczmxODzc46xBvytOif5dn0m5EhHbis1u2lkmvauVR0jfWPa/Wn/shXMzCwOPevTvVhMBHPvHnlN
NgtCRF+rJAEqmDTeWvN01iOG5x8LdYcNy1Gm4Hgtj6XnXJKmBl/5P9X3Msl4KGE1zMEcJ+0t4+Qg
QqXReErJXsgTwe7mSw/chM4UBcNF/LEurUAHgpVjX2Uq84jcunxdc7Ht2GQ85/Vjj/txehW5Yyb8
8mQXGkO5Bb56f6TI7AfQVpZyvz19ZuGtW2fdc3lwXiwx3IDsfOW9IizUV3z/UcnTwrs7Z1aABZ/2
ceQQlyOiHNpv8tUKumBhwF882z/yWKatXwMPFYdN4w3jyrDSWuuu4FnASQUNZcI4H4VqSfKuXLny
CQFmlO9nFqbptv7wb374+dtd/ilFcevAZdLlKtv/ljQ0F299Y3aMUOlV9GbugjoeHkEmi0xSg9TZ
zNgZrIYap7DWgi7QkssP4nzeGxatfe8XdCzBLSKwmoAJcdMel0gcbs+Rjp5KFb4SyIG+b8zDunMs
FDHtHXO3tKx8Wr7u/QGO4nJQFmmYoWa8uIFyaK/jH/fsn7EsH3yMhOCMnu87bHw9OEJY0fvPFXRo
o2kYSSDZsWyv8qp6zeZRykG5N3+mWru+aXrf8aB3HGwtG3wE++pZ+szo1J3RWPzQjqiecxJd0+kh
nETkAunEp9z6PaSoO53av+UiiGjhj/RQHJhZyQUz/Knmj8pxxWe6aTtB/n1fQx2C9Y9gNAdbIsp9
H3p9dg+w1S5uLzzLKsVBiaByk7FWBw14ZlbHmg7q5GOSC7jQz1lDH9gJeBazvDsl/t49eemAoySJ
08PQtjdDwEH+PF5dHyvkC3exOlFA+YMQzhQ7ANnpoztdb8o2DyXuiXsU6jcoKfFJsSOAwsRKizyL
oYmgxNQZ8kzrDjrwYfEUwwqLhf3IMWMFKA71iQ5qEs9eApQPal6K7VfYpUHYAI2R+KwdQsQoRUt7
w1TMYkhgmTutlBs39zyAztg12f/iYgutEugPrhvDmrfhXiIIEzphQfk0N27P3EOGG9r2CCbEuyf4
qMjTINGS0XiYtrthX6mCUOK7t0HtrM2x8ViPuroSBPpW6bY/UY63ZRS+eBwSdCc0LOEc63ZOgrGs
l7+695iyzAPukcybXehkebOykKYwjmJ47+3wkRjVbxaiLBNs9HcNvRBcv7eylMDXvWuTX1L29pij
vUjD7wmomkOPy8Yfn3yDoZzZ+dyDHuONo7Q0k5WWnjkdEhiFTLtZKtRLK+5lyfnH2oTZ7mIjIyAq
Q91BbG5rp+wTHQ4AsqZmNsMzSml44eBCWvcx3h/SMBCwKyig25ZYLOpFFYb3frc+kfaZULl6cdQT
5DRJM1qvxADrnxCc8NPqRxOOnaU070o6WNe2FYym650kroo+6AMaDw5gqELLCREqwYeobsPchwNM
8vXJb7gGJ/u0lZQM596cMG/UPyGEtBIEWfsuSr1MAj8q4CvhKUoDE6RLnsr+KBagsbY2HLflSa2l
wsBLFueX23Tt3yLzJSAYEocIRIrTu3uXbzqfLKLvdqSziupGay1IhNazhWxIwNAjxUHibdEWz9dT
HGUN1cGkWrPrvM55PjOyJNtPtMn3Z7KdUrnPbHzDCOSqPH6fr2VojdY/odME+A8rIHCh/18gOQDR
y0WJJd70iHesUsh+ArD4o17MxfRzDCv0rhDBaaaR2u+q6htUsrXaGtwsLnLIguVY9qcLDbpDKVdC
k5WGOT24U3AaaTIMgIIcDKM3BtQHQFq4OtDPk1WVbV5MEvoMiN8+vDM+rQWcAKadJ/4lJfCOaR1p
vBu2MqpkuRmsbTn5O2vVvw5gZNZzBSN27hW+UBg4HzaeviAirpceW9vXZVauOKO2OHOZ1YPJIzTx
AgbUgFMgji9c+zLzkPJeqwvRjRJRy4yn8MJqsBiypG4QByWbyEMDSl7aPhEWLyeG7An/kjdGizIS
Ql5xXJg0z3HbzPo7BHzTGcCax40oIxsKnRZRfhDZvTUczhwuu1OgZb8Q7jB5K6vqQ5LE9erv9BNV
9J7BU7E0ExkTUJORse71IU6MuWOFlmfeu6sVB4yBuxqh5tUWqZvVbOPzk5zXposk5BKBVTHWCVDo
9vwijsKgaHp3dSVtgzwzd3neIostNUY7tTrjncfgnIcq/vvl9f+A+BNc3naWon8/dXegcrdYS7IF
xv7c+zIFSSyi5sMajx6G2ANGQqkTJE6j6DGlDny6JDJyWGKCaxfKtBxuN2vChcBTW3OGCYBf1kx6
TBJCyzVJ0IJlmf5GmHc9s1GkDQf67XMhqhAl/CO2z7zPsnD93644IPziV2pRL34B3ElDcoh8zY3s
WxWE/nGVgRDXrGSJ/OtVIW/+Ss7gmkTCrFkEEiQvFs/wDyVuL70efzfPPZdycjqXPHEe3U/CDvcT
wtqQiX57THjRytMrfJXeVtJUvQ5GmmMAcdduFFl5EhmC1Pjg0rpiJ6+ctdqrAh8Bx/eIzBbMnO3t
fuCF3IuhWLVFmHG+MM7D9LOppnIHIO3QuYTKpUrKCBa9qpBboN7NCo0DquV1fwfLfo4aEro4bxD/
P9FbgJtp/9QQKXavbympEXMTUMo+Dace3MpbWm7Z8wrvsw0cVe0uzPQaxYWIeYYh7ygEqxE1MHhd
FdvvYuMHksfY/XVBXCtvmL9j6b9B8likeGp/+T/xpp6LNR9cSpkjQqS1V63QDIG9eCTsvmFFklpj
RBynuD0oQ1o9P6QHFmyhr9YoRGbxyGykYbhdACZWVL3ooue2LcZuOkXz0BfDqDlXSPrpeqd9tHFG
AxvwMbUjAPLtKFyJbKzPRpWsfD8AREEZdR/0Bi2pc/DVH6b32BbwfkfEI4R0tqik4y0iREdlxvxP
XGePWpapr1BiHutAC3OGu8i0nNLwTp48MLR8UCXckYLn+ROP0FqG0IH/SmLW6wzLpxw3DD8zLW2K
wZkkmWRJCJC27mjjbINLxch1tO2NkLBUO1Y9ZZaIxzZ8L0sZUWPqt3Y/ESFGqFXdhzkrBL4+iDda
QXzucEvP7iYmENVrSPwXTW1CprmuH4dDbQFXPj9RfShDhK7qE4es7Ch/H1B9+841HzFDJ1E5vJj7
tfoCBUYgEqT/CtrhKAwRJVBs4ByVZwDOG5YsNkn2S85v1GMMANpzUlex7xJvRPG6A6AVtFfhc0g2
vlaW56Q7Cq6E0T3MvNzJ7dTaqRtC0SY1lMwgL/M1Gmh4d6uh3n7A0s4alHUPIlMBoSd5g9QQCXhZ
J8jZy3pAqa7tbDteu2MXORYdD8Yl4klZ+See5KG+DoD/qxC4R0Lmlu7LoW7qAawd4m6A07h5VcuD
0JdCOmQn3kP5Yjuz0smW/bB1NGc/Cd6D2FIHfuufaMz2DSp7v3jiOdeptYzSJDr60DVYftzE7bIc
CaMMCVJEG91lEj6s8vQVaZ9E9R0Y8OgzJ2PqTon6zJtGVZfx922U7aRxGfc6X7uNHhr3vE78TL0S
yjGQ7z6GYHJ39wx4I0YXDc3xApDjxXSI1FIEHo0puTIXhLNs7NeiIrwsqRYyoHd8VSKbtya253k1
JECW7XRdCKfP4vOFWa9+SVtV8kLJIizk0dKjUCZ3RqRzXwDm+Ka9adhYNgWYE58rcJpSp7t73xdV
F3wqSWsultN55FF3tYhjH6Pj8iV57aPdXJ3gl3mWULGAsabW2Kvo6++Ktz2T7FylgpsKKaybsCQR
Z+OTyl/DOszaRiUdb/CI46MG1cTPzkYgSFzmfFxe9A9BGj0AULDSqbrG6BOorapOcdmw0PpPZscv
wzPW6WW6CicOSSabZcMYqc0neQENCcerd34vtlT1q9kWr8hS3xTOgEaxkKXDRgKDmS+da1TCSLVH
VzWdZi2IHEGYxFag1rXYrS69fEB79wqbRQdbsAOnvNRIRJFrh5B92/ocNEiln6aac18DeFWvpKfJ
5zNOqm+hOnttoFOCziRr1zJCmdfl35fvwOWIrSMasEF2o4MBC1V/u7eoC45Vr59xffMGnbev/gUz
0XpPm6bh+W4pSwS237/90RAoJbNBVzWCsG2aTbu2VZ2nRTajfBjyzHA/e658P4IzjUvdeq3qRSRO
LrcpwgMP+LkMLkmzJYxpqmyRTXO0hMqoPuvSDGk/AGFR3EEcdkLkJrZd+JeEG4YAMX9+wp1Ul1gy
Hr1u9e8tLv2ff+p2QySOo65tVzlYBoSPyPEs8aampb9KA8vd6MAJiXl0QVeQ2j1CdWko/1F5ZdVe
fgkOtpO5OtSvH0uXFxk8x+AnI+Q3xOC8OYVJW7llo6LzqgTUqVSBdRf7LKjl96yO182ngcrmM7fR
jgG4esaA6WQ2zlh4THitkhbkXXf0gEIJOHmWnGdcLB62A/LLPlDQiQdy7dDpbjeZ64/mLP9aa9qu
Llb2ofCjCSKVy08VqQFRTvffkvTZaPAXiCy+892HotoF/2v+7dd47EgZhjMEpMPZKPiBxx9dvMxk
PvY+8o+eg2WNJI8mIXDzByA8m1CKWuHn1NRuKbSyx9CycpeKiR5c8zf8Fpvf/p/XE++rMmHT7QJw
Vh5JvrEnqIwnDcraO8K0gXuUJgwnBBk7/rymfUm/CYCMdopPzGH/P4fSRvrGATB82JlpdR5cXDIw
ncasNqVtHYB2aV4Cg52Zd0q2z5RIVxnx+Og4+FduJRpOskeyuqfu6UTAayN5+lBLTMPYVXKzNlA/
mf7cIGTBWFQdmiZFL685sIkrpzGt8XZs5lrWS7paySs/Pa3+ERLOFgxhchJPUBBo5llpocJVHEGl
RMsJBkkS2ukcCXLl5YCCerx1mQbTuA/HZkaR67SGatJbG7mJHeo+1e/DTWTLlPYobQpmwSE6+3vN
/AkNJHXQliqg28YU9LxH77tud6FXriQAozUu1IWbDpLfOC9+z4yKWWKAY03VVa93m+CwbJjzuMXp
bK7g37xjibTY0/+K+BZPyMLGQj30XQzrcpsUGukBCMZ5ljkI3C6qReyVv7/LGACRrb+sje2G/osz
rzjhzMB87xXUjoyxsOvA1xpbOczt+GbvjtLzeAIcjCQds71uZOpfQtox34EVhD3ERukOPaPuSpJZ
Tsnkn4SJ+2/sahOk9d4yHo7ObHuIhvYsZCjr8JnonLSelk6HUsEn7AXeC8ghNlleUkI2sCBY8YZK
hB23ns2Ylnuh8A6/ZS30wTxwJ4n/ictVTw4sf7Q9X53UEi247fkRpE+TCOuEUHPPmzZuC8Q7FU1g
77uHNGjccml2ZHc83A+HJ5HjXKAUuEN43uBHYijwyeVMhrzmCRM5jwUMqPg1Q48+q/qXJlh15a9j
TMxPebi7jaQdyWK0G3GmjrKMl1Wu9Lw7gYsMRxFmTNfznWFq+fDAbdMmzFTZ0YyFZquZ6Iyeicnh
33LgyKIQhUBrXZYFDLdUzXBl0c3HkSwTPQhRpLc5NsJtHWmiEvZccPJey6ygc8OPZyNsQvoR5NoO
cLg0G3dljrk5KagcAqCY0vg5RylEWXFN6CvGciJ4RbA1CKdEKR+HMnRBoGbYDA/KPK6hagMQrm6A
cI93Je2s+ShLd6LR2KzYcgu5A+Flx4droFP+mzK6d9HOctBcOosm5WQV4KYXj6Y6X838UIPr/z3L
IbCzsntvc9fUKLaPVGBegmBOATM7YHlz00nnFAbPLu3w0S1mmNw7VEEAtUZWfDh+e8S78zrSK5kL
s4xGsUlduoTl69nV36oq6bAKHkLsFIPZaGnGm18r+HqFkFS+57n/l+E18GcDJJOtDV/BOBdrg1xv
5r0o8ukL8BzRZz+jps9o0wb5+GF96138XKs702/uuWiD9aqQGyGodMOA0jPtIlO4llsXinhXfX6F
ETyacy0b+vutr3gPXzxf/WtLXFPadTt8AF6kiderAKdp7P802KYiQJJn+IbQPmSunzm/Li5365MP
oLeIr2yL1N1/sBCJdJ/K9eYjNODxcbJjtKra06QhNPgCXUr8kuy6sO6xpf9ej/5Lquy2JPIIGnVe
0tm2+TJMylcuwrngTOOD7O007xCO+exAbEwGDhD1Nkq5JRpnO6Q6+DfEY+gDEyQvpuqXRI6i3C3Y
tCUxCEq3xfqd+AQv2WSfeg8Kr5oIPjjHJLCWVCMLXkpYejVOjN0CXDjv1UZrOkXpt9NgbkcXSfN8
HCUumothQQQQT1Lm8oLOHG6HiT7RXhLVB86jW8/MXSEUiiPHi67gVPi26gvAN0yNcSZl8jnMxGm/
VUOySc/NP3nLc+KTy3Z/AK9Fg2c7KHgvqOgLTOiw4lYmaHlBwbvcqycBdx5fomVvrmsW7y15FKLQ
4RRtraSiux9+XfaDeWBOI9TSDHQtrnYutgLoeKVLZei8+N4/GSzqCqroEXMXUqz+2GhSNXQwxHQC
zSc+eUgiKxZX8RNz64hEJzEW6IJDRHAZnAUnGnkYFTq36tgGkiHH5+/7N17Yr1oP5qchU/qhqvuB
bU9AWKrG62iyQLMcXsbT6kCKyVzcY9Sv/FYDc3WQmk5paCl9x0Gf6ogLQgjS548t+tetfMHl4dL0
zqoAzHktrdJIlnxyCNQgXUQGZ6Qyy/MkO+6zZxI6M7RxHXFsnJTKfxqySHAcIjLvaennCOotAb71
89/8f+8lMhhkXgi9QZ7JFk+LhkMeftWyRvkkYKe6ZpbdtOlAfBDuN7s2MPnL95eTSiAiQoenezJk
qzXTsbeAs74ACINHR6lMW/Gjy7Jn+PBzMeCCY4npEAzqTDYwYYQ/Jhiw8xjGsPjO12nC7mDGPgil
ZrhBP5TOenMdyQO5iON+MUtxZhGxpYK6K5kfTBPW5jSQ/rRZOOlB358gMSct5jzOBV7utQdMbgq9
COFZrP1RgTKtf1PezEmjpbSc93TeFZp7r9SO/uY9+0VcmHwpRhlWFLKHcqmI28TGerKaLWTUMywd
pAJfaNnIrzQp6tEWobXv/sBenLoc1xpCJP2UnlygHhSGjSwnLMBTRBMVbt301boOfpXhr/VEVrT4
7xLO4sAmuGA+OuYDL68iH+tZ6uvHpsVhUJ/FPHInSDOaDhtZbKErlySgJQQQ/pHu0y3yt6XFRM8q
8Bv/wnjK/bVZ6AlETVob5+f4z5C+zoAME2eiKM0FhSqDA/aL5d+wYOKkOZxRKbjPJwuddLaJM5Wj
JBbC2gRAHYpdieWvxpIH86QxTrFr577xIj96nKJqVWhbfBpUqQpbIeX7Jm4L7qqfUZco1nJ9+ZuN
Mp/cjOlwsw0UHuHs3sk/m/qLHHLwqJnk4qY2B84DmNHZPJjiGU5ZolON20f4pHgLn8lo6geFgTzU
kjgBPSbttnOdRec6oOJ7aRvpW+DZrKAzs5Gzcmm0IGtyyU7zUfqvQVbEaGAtGKwutKK+Qlv4L5i+
mzdbGl0o8Bm6DFWoJwXQOHCWEyEBcgj5/ON/ds2dNTXWop3MvXDVpFAwXuMzVSUCr23hw+hkH4Xu
QjFtaeYn/rn7cgrIctYrmuxt9x9Kc6phyW4QKM1qsbiFMDGjvHS0K4yhfPRowtEOJFCTkTk2Tyqz
fAhEFsRUZB42gLhyPM5VgFHmruyPzr4DDuXWwUX9ORGists7vfyxYLWHwPnRXyMmUFXBo2TEitG/
tU1HS21C7GrgNPhPPYG2f7t3mQ3gAcfIXuIc8hpmGgcR+gwcXiSAwIBx7q0LgohXbRLoofzj2qIh
FhQdps8AmcHZawecYsyi/f6ozy5wk7mccxuiidclF2v3KgbvM+GLkC51IlWWmkZhCSIXMXJ8iWfo
brpYrDWKAO0u6N6ODk9FfEFlaRUAuPvhK/MW8BlSGkibQUqO11xTlm83h0JJcz3N6jKcMquCJQIJ
jOflVSNdeisnOLDj7/hyna4wde4lppsEPaMARMXGmjEjZfyDbv5WTJVmxRHmLX6eC9t1I45MzKJs
FSpslx7kbCDgjhT6QbzC/Q1EgGt8hdEa26xWylI6Q9UEVwDFCIigiJgEB9do53JiAunitTAPzdHX
miFpNuPRX9zWnB2f4K0JSAeWRe8QR160uq8h/ZwXBwCme3tGpKKxTPvMWsQzlEZ20oXPh5SDdMVn
6PFfnRei36GbaKjIrUXsiQZtjBZXxlYZjL8NNhOucjtkRphU8kjShnpgPVENbhiG0k2kGoQAkiOC
hCu47hWSG5CFUKoqdsHYgCqB2/oQQa318UBPJuS09RNUxjN7bMqx+bLBY1nE9LDfYPJu4QRt5o2k
s2swg52jY84DYK0ZFs9i2t4NvBq6bA7OSIM0ERC5yi7HTEt7wQhio1VqT15tkcmAskiEpB4tu+Qj
YBt7eqVCJewNP+k7GFkDSvJ6920LZF9STOPQCl6Q591axDXe3iuckTVEkpkTl1IZFDxmo1WbYUa5
eC7tEo5sup+sv4xLcpPofA/xj12cs8fSQODerlxmDDAhKUBXEx+Y9f2i9oRaHJzpyox9Wfdyc3fd
BuX2nQOV+X/AtjFwJB9TQCH9iLs4rf7fB3MA7jSSmNzGTatriwY0EYU/Kcj0/OGgYtlK8ZrI9AjL
pcjzbdjP1LKQViR1nLNS24JsK8ETk0HvOsjsajf4+MYDdAxJKy9OZq+SFO9mZZR8r75witaI27KE
gXoaJPqkG0dScIwr4c9DVK/6RDgnKOqW1gfvjFjHHJ23vTHAuNP1iDNYkwWg+2Vf8qxlSgqBIyKt
fYiQwdVOc7+C1eaGdBceKPlk/SfI0PU6ums7I/ZR2S88W+mvs4ro/lKg4EdtHhirBp094+ZuFebX
gBwVAQEkv9hoOEFmOjXhjqTo5eEiYrrH0e84gLtTWbBCObCUeHC4wMN0Lv7N95XllzyIj7M2rWhD
NMu4RFUg4yK+td9KfQJBgc6rA/Z4ss34JxgjsXeuUAF+X1dkjULmFbuigIuFMjjDRF7sxxZDakVK
UNyrcggftouBl0t6d8ZnB8ykRpNpOGGOO/65a9jAZCkwIjLA4dAk0b3nkzR52tZoHIhnkS491ztT
xxRvJYAn0RlrJE5xCE2VkTJwzcSyz0FePpUcw4sc+3PUtsEuge2r8I/xydAvy9CLdxb7vc0vUgO5
TeM44E92BoJQkyF/PniUkwfj6TfJOcqbuYTm4Vy7OUvlnEAmvOCsM65mQoCzFVe7n2UXbWM2LChn
ov3HeNezVbVYPmKJKYTZ1oXPI3I0VJuy7zoFN3Nb+vx1/e2S4O7O/eLmak1r5yCJhjusvUvOBXZO
/EO6Gfdp3zlIxZmGMX2I7HknHKtVr3kJVAfe3yjrxnD+zM33sDCrlzd9g7LHCzP3CNLyfIrnspuE
xOPE+c+DvXBMhXSsZQ2KhcUBwRPndalrBKdiZ0pMM67qeGDRKQUJYnxTl0HJ5jZpgcIxxTo4azqH
gNSRo1mZwn4QRfedy+Q+fuYT2TCNjC1maJCVBjtAzKGB/HYFpUtrDaFcuBZ0RkaKI77lHD/Daxo3
4j7tGHJZ7n8rjywd1ikd0LTQug0xdfvo5MAeexmYHsSt2KXf95LKmokVsYoBaQwwS9cYHyy1r153
UqZcmoouy8FjErqs05whdTOtUyc7PCKOk/XEjUw62ExG2Mj/qDhz+lSk3EtB+HaN3oUen4ivZrjX
7Wa1iCSLDOGKTqPVR4UUomwGTSaxapI4YmPGoNGKNKEDtimyLGDerv7ziud5AsCCD7bRyFfdXSfA
2g07XnByPb4tCGLEpNZFOKvl9KmT9uGT/hZMKZL89y3OWkR1jkcxPGOCExoz2hC4MsN3htoqwHJw
x3OIluwwjN7ztrIDbNtYWa8/LeelrvZC2U3MqO6Wfqi4MJHR1Vz1nRxbzSjld7ByFfgpvcHYrecP
e4XxXUz5e9M0roEYS4q5U1YBzecEYrItylY5/IOjYMFMzJ7HHb5dXwGKKCsTONWgKKY8OzeFECjs
TP4OXuyb8pJBrvdpy72Myi3BX6YFZ7vNtEssbCN7d3c2M17UKH1PJ6Ge1iaYbHybLWfaDdvjFOlJ
fNUWhlXteCvSaAoPj2O6r6+GVEejvZKmaIo+EzDH4Jnn0Qd6+Tx7ZemMJMqTH2har3cRp1FDMJPM
jfte8ILSH/IygX9ukvdlXMg+yMBw17UHwXNsuxnwb990yt4A2vTTzbGDQieh5jxg/LaueE0BMavh
6D1GmWiQU29Nl2o9xoqmwGZ/m7i+JvtqubI3v4G3lH8DYdkf14QCpojKbE2nbldT2f2ldrtwNzni
j81gOLFrcT/yYbBI9qxmLvskuNntlBxUJ20ic92Y7UdL11fUY4stu58rgjqE635/VROqMn1BOTTG
MS4UwrIDXOSLF37fB0nY4P7GMI2pI2ecz8FLzU28aQm/Yj9zXTrEhcjW12gqClWBmBY/FwygY10Y
1XUcWysb6klU3BGL3Rn/ntol0ufum9PufVootljXT1ju/AFb+1zlRF2fPzLM+8NVLPSTW57HZPFp
khZLPB03JAaXs7UFbnhoJgGtdMdYEfwVvdDw//gm+RA60EjBw12P1eSL8V9KQr4UBiFQWjVepw4q
W3lXUNQqOQM5otUh+dhS2WP6L2zDW8CW1AfapIiTzJ5wSn5PhLesRtvJ+txD3/DiMaqRUulcBi5P
I9lv0Ip2d+DTmhkf9Xr2/7wysoZzdkHnZdI29nz5ZNbI0MPhrmsFJLdPcAr6V05Y7ahKx6HAv93U
h4enuXUJLDgfdj65n/urxuMH5wktOfFZ3iU0VwqhLPcZ0yX9PsBsbBxr0u0oe1l0Rtkg0SzEf/Vp
MqGZNDiKIUfETuCyWHkMIZQiVJ7ExQRkHOG1ShvgXIZWRYzy7ZRrbrZ9dbhItoT8kXxhEygfdbK1
iSSUc70yQwM2zqchQv6YSA6SwepxFjmtFMXPxFgKyB79gMBCrl91nqBzKtTch80CPlQS+a3/T3FV
KidPKzu72k99Y0B7ehHtydsChalLYhVHZQxWkzYUqFAYj5eN4dOvK3ofvXrPvPA3miOlg0nYdsr6
4g99GuFzJUMDv229gZWp2lZRDJv/7WGsQmblsrZD9cNigBC+rD5UyqOtzm4C6CcsP/jSybVfW4TR
Ykwd/bx9oqnJHo9jiwcIIlY5AxHU9ohbHjpBeisxR97xICNRZfsuYCNIPlTfgqEfO6R0rZL1PGFZ
OY58JT0WjCBPJVIGtdNrSCc9lv7MIb7XLhentrR95SN+RyJ8wRUkZv03vMebJh0sACh0lzuA9hEv
cx6kR+cLsyxvdIVl0Oyzmgl9bcZGLJWn8X6MYLBSqqhOOCQtUtbX8UFLeTtno4AzCIpKajCd+rD7
Hcks3xovhDO10qj68G49oLWrQY1TZKb2bHgZMlMF/nsvYWQ0KFovVvtcH06nvRt6jDMhfw2Lr+fU
t9NS61LfV++3REy4PY1MPQkRJpFhvqdQ8IvM8pBlvqQGjegueg0vnLt67NXbNHj2AMA7Taf17cmW
ZTr5pAi1z4INNKAk/w/WMBSf1JR/ZE3Ok18pBgDwtMpkA5s85JMqIXV0V8/cE+sh2IhblnIuFfA1
08v8cksGdbUukf1Fp3ScZYdc4HhRcOLZugobmcadowL7AsGFtGVaO5JAu8qNyE5kPXegemSK7U0r
YIBeqfXVqCfqBQPOQQz5U7hkxEFNUsnUoUBAii4g3r5NQ/sR19W1fRDVWvrAyhU/b7j5Vmw4ydeV
OV9XuyjwIBb26EFRk4UThdDFSOENv6AT+nqNUb6mOxB8ewonHzHAPPb82KEos6LGFVrwHueyLy1b
rNowNdp5vuqRAB+1B4mxcENRKXIOD9ql7wW+6A7YCWtOA9gsYwQtkoeFtXl8RsnxeCOAngjaWsFn
ige7Gnc5gIW4EiWNRwP6fLBouOXqF5319V8Cnh95eWxfzO+tWq0lXEQv6mTNPdYXrjEVxDkFFvDh
YyDr08T8timkcGSrON8xQS/zUFUKEOtareZIm7jZ/qfDzsn1WnSVDnNgndPPWIvXpxjXHYJI9ML8
gPiMid+tSgVb4J9N+aD6XOAP2upFynH+GeMiAuovrwKZaPQC/14L2fIBvBseiN9Em+zcASGWlf+y
N7z+EhWJ5Dwgl0lE9O1wxVnONKfUvdW/3KeixmcfljJFRcMU98OBjR2zCBdFAjUIqL/IvJSaKshk
fhkmftsUnBZNvkbYNzmf07gBLjLRXybnH+gUBqUu/OhT1TMOuRzns1c0eWmNY+LYuDkuu8tuDwyg
IC3Zg93L2SrF45SDZb+xxsDR0SJejvhRGgs2nJs4KKIoyS2AZO/kQz+qdOlFTrhPuPjdd4WOLsZY
vpNprRggclm+4SJ1VIJvgaJz0t9lilEqD4iF7k/gtpVq8/HjLMA2Xe4Vwt7hC4BkcQbIcmS6Ukpe
Gbnv2SePif3JnVz+1Az7Lx2AkJfIVD50I5P1zlWwuR0+JT4cn80kkVOiEzU1YwjDFLWZlzmOPp4b
spePnmOsXUfcGGs/kVNpK/f6wPXXHzSjgVRy26D+6HAL1jJQpcmUfxyFtj97W8Ymb/dS5ltHhC1R
Exc1I+55PZd8ilDP+SfGqXFTpNyd7R10F3DvERHcepzuGfBtLxz/XR1UwO3Dax2ToJza9U2+Go6L
BVnUjW+BZK6sMI48GZsaK1gEZRrpPpxvX/XCD9e5v/+XlDdDSNVHDMS1V63ZDIFe6eC98gmrtdcY
JZMXtzQNOTCDTIWP/AynSPOK21N8tA3pjVM1nR11B6e+Rd5yXQB3vGA/X9uixqmlnnMmLXSjuNA+
fU6i04lzsBaWA6Po+qSfTJggF+nztgSLhZl/qKLko6eLSJkzbOfeeVcPilYqsY1FxU5OHi2FztHb
fT0CqVGgr6kaq+er+8lU5KHDmkfwoJU50Xcm9i0W0UbulCPvelZZzDyMn5uL4JaJMx2MiZM751d4
c1SJtraU4Vpjd1GgIwnU3fOajE2sC2Bwe9nuJ9RigoKXpgVnzebtw/WQJBCBYa9EdenbG78FWYgT
5j6GDV+8PZMbDLwexHgjwLc+EGKszboAPaxtlc62VIdi6IWaZHH34EMFN8EbFKwe9YQ+lw8/FtJe
VEjkMcVv8jXEfBeg+RYsVMBPwPidmMRulUZzSfcCE7AmkIlSHjwjImkvuLLXTXfuwYFReBfJ5nXZ
dFzWatfsvy6pO9rW/njJDVKifwLiRNgmmBEUei8YSMtNVa3+NtzKmsZU/fVmwNoIzHjXNPLnVyDG
ee9sYFHBTxBt3Wb9U46Ish6y+oSZdxjF7Wor71h2ZcA2rhgwDHLDIIFs2pk/TQv1p201v86H2Ypx
p2OBVkdzMx3GaSxit6C6bfre+gapQqwCfkcPMaD3I6Zze6t1/dUxL3JgxBKlJrW1mWlUHvxHiV+U
1yiof/JLj5VZ7Q4b9aNCY5P7jew5/7ND8i1AJIL1hh59GYsWI8q0uGAwuX0h+9Y/27k9St1OXdeR
FUDu+s4Lh23Zm5P8E018L4ZVlhcOWsYuyPpn4fasfNEcXWS17FvDTJjlTbthj0Jp/C6aupa0UopY
3fM0sjeNqxJ7g/SenMy+OZcrPLYPy6BtXtEEcdQYzVavM81w2MH4/hsGw98sowNyuoODY9tz+Jsj
VCYCbxGLLK0k+64j/9sJmaK+21xF2PmZjBSh7YwQbjwWUBe71EMr3dPkgg6ojcd+z2TX5qOyCIja
28K2c9vkgdAzttdb51Ki8lKPbUY6FZhTEolUL9cfzz+sWzFzLDmm3p/eydEAOWpsTFy0oEUQ2sfT
5ZVlglCFntTdD2ixcf1+dZZ+ayTgDYs/dboBHRpgOV0M9qcv5AyEC8tQs+9FjnB/ySEnsTsbiudn
NmhPT9Jz7pIMlUHy74Anvsrcy8m0Av8nVJdY4ewm5AqPQi4SMtZmp5jSJIWPm/ZequfERfWT8ERy
KYwpE+IIYGAKwHsz7NyRE39tu2wNye7Nc8NT4hQvflBAn1/Nq4XJLdMH7reqbgLZCMKPfevEUgSL
6+IKdAkR3Ahg2Q2qE4xceR6mq7MbFU+b62OcZyzusqPXp3ou7cXyCILWcVx36Ok7eNel01htOD6/
KRj59ozRj6OTnJtNfIOeHxP8471WEn41ohTmwJuPcsFhbVY+j45MNlZUT20tpXEYCBEG0oO3Jelv
+Dh9I1I2BhHZpDRf28jH5auj3Gqb/jV3axjl9XHtuqWWdPkIYHtFZxA49dqPiXATHboANxugerZm
MBP0a0D44m82PACUuZKKSN5S+Aps23/dPUwl2Rmr4OgW8JUBwCt0/A3htH4OdkEYg2HaqP83Whvo
FEcxgXeIHuGKH2+TES/Em8V6J6h7v/u3gJK7Wjp5F9Ybkpi6HKwsPyiJifRp1ZaknA2Fpf5SaLk5
2QpqHmJxBomxvK8roux6iQ40sbChZ3riR/aYqr3Bv0yH7+HWuBlT6+SBrJ4UYJ2Ch9iLaYRBrQtl
Nf3C51S+lZYRH+9jedPWbUXyKYYFhDB6MifqjV2WxMpgRn8pSze6xmXEGozE1hf3HsrplNRePEe5
gJE8qbZaNehhInRclZ+C2py4ZOGshCizvjSgAFumlM03cvQDDOQuKy8ypUXdwiVuiwHfR9ypic75
CbfLPAj9w0FwEJQKpi/nySqiquA9fi8ZJdBnYor5YAxZO+6bwVdTDzyzV5yR4cRxObH9/ITaOFVS
FGFwlNxQq+0Ottg5XPcoD+h1cEDajv+K7NQBrnAk9LDKEBL8khDVTZAY0mT/GHStG+t55fZIXIgE
WTTX53oc4ODWXJt7+XE+OjPPE26WrbvMdCjAKJUAvonQQJByXBmDTmGnTZlQIiSjbT/i1ebOedSX
riOHRYPMCtFtCw0Togszaog1Lo+hf4FN2O3uaNidtOwG+wnJXyDu2Fmy/A9LOhGoCMvAC+UV8IKF
0/jVHJhqEaiKc06DeUFosMLOyXt8lUzAxCaAHrMvFRHK1E9tL8iCVLbGlYL3nuQQd7wZ7TX/R4H+
sB5tWR9y7XAtb4LhIiNJtxRaIiRMbfN0oWlTYLqb78ldcwOx+kX67sRoNFVp9k8pMUENkrgIiWwn
e9U6XoawietY0/9g39NqR7hh1Gnjcrc9qQyGcsAURb1TMFdKJLVZ2c5VvA3puuWj5dUq7Bl6Dvbp
A/TeOvi1X+nB5lfsZOZ/VyPnz4mJ1Dm2iEW3aurQmCroEwTPadGNFxx8/1IbL/IlaxUFRPKPEcXv
DHHo7+f86SIenmgXWi3mX4qKXdsst0W1yV/Xhyh0iwdNA8QBSXJYxJ5FfcRL+8SdVzr2zT7Yi/6l
j3rQSOxEPpXYGjh5DReKO1KlLHLblZQ6jm9I0IKs7/uukzst9+o4ZYKJZQDdWtq8IR6QoCrrKrm8
rdpzxY+JfgStR5n1re+7de9jjMEDq8nEP0nr9NDUSaSWNSZmdBLfTLnNJsq4/HMG5EadP1WQ8u0u
HoNrwbEEPsKMDUyt3nJ7DtNcd3lBi6ViStagPN2NTctXbOaw1P+pndxtUtcXe4xapPsFPCUOXlxx
5QqhRB5oOMjFKnx2FMlRpxdz6A2GbczCCHiTEsqR+McIpttuVfDEq/+rISnneOHFJRj4a1etzskn
9aYp62U+U5gJan9QcM6SyvlgDgnN6OBxuJkMUDia/LScRXhWPs0eaY9qPzqyRP7RSqHppN1MBrka
LQ3+d3tuqWJ39Ny1xFx7uY/iEmkjveJr+BgIW7GtTsfd6kvAIuch9Xmcu6qwKqpyoyEJ7jJinl6Y
hkpG4xScZwm1WPHbIAzqvCVXYJLYfNJAOiEq2wwDmkPbOkW854vd7FX9AQ8xxPp9U+OS2eMzQCUN
BOkhTSOdcbOhcDWmAVe5WH6omznXChFFz4xGyXDlG8Y/tklENr9wq+IjyfOpP4x1CrKcOXWR0o53
JKMQpzXEAvvlwVa3ZLgFlp+/0vZfYZKFgWWxTqSNvuhAZFr7+K7rhFlbynC/nodo4eo55Lzpj7DS
jyq03OLo82et/EKU2bAeoDsYMrJPZT15kCocK4Ssw6zzfUhDav9b1sbt5zp+NzdQcXiytvrBfTOa
EKCzkwTm1ZBQs87K0xeZPuC+3tx5nSWWlP8yvKBoUsFbhcSt1Wim5CxPhrvbIZsC40MtMATyfXRZ
GCteu5tbf3DSEzBII9T9xY3q6htORQ6CKcjO9GE3ZbJQ6Kmc9FsvE+zKSTqU8j3fi6VmD2HQZEq+
2cNii/lM/wKapLN0II0un5invnfwUmH/nvPEAAIjgJXUQRk8nysOq6OMXqDhKqCf/77VJ+oHPZRu
6P8HLAeqK9DZcKw7E6SbCNrMS4VbJ7lm1Kt8IDyxahgZo4iaRfMSK/UGpjsQPevsda9u/dL/7HOc
9FlUmYL/CN6lrry9/FLxCzoyM0L+VpRcDyYFOvN77hE2xvB24jrbDEw1+LwakUe6zXO47mEfXCd0
iZ/nIGdeaJLA5LpopsBbMAJ6O1ahtA5BN7h4904GBAxYhqHBFVRXCV63kWoGBT7g9QGq5HA6cLOS
9VAke/2zKpR6CQ90ZrsQUJ+AXmKjNFcD7K5pyyHi4iAC/Lg9h4N1hROaMxr4igXBCDslXAjIIdDH
aHClyskVfasKz2cPlRSzQAaWw+hmIY00MmQ2E0qGjB0HXIs9nKjsJrkq8Yay2xJW+qFbEsBBIqyU
R2RrHlEjOIeKmE63fDNnYzNBqaqcBlPRQh5oG3noQdBAOw5txmjV+vu8cF0JWPv0kj7kUi7oNCVC
V1wSfKMQSartXu0HEZ2nk4LQQsqbDSN8z0gI75fSFEejUzui2+FEZInWJtAkm0ltVlXQbic5wS1R
2LLeOuulPMWhJYTz55xECW2ESSQ2YKoz5HuJa6OtZFimp/e+4NdytHO5Ns3vyIPAyUNEBObhT+Yz
e4Ahe28icZZsg0BCunPNePXqrmP2P+UpcuHlVK3oZmEfkIfCgTuzMaXYy7c0glHliAsrGc+pE8UQ
zBJmtK0uH9GkZYqYXA6POqYuBTA7acTe/gYxTY+yvCWwJKNk06amdfuO13HRuDdBE8f3wRM1Dvep
jf8kBc7qX0Q4oHoRQKSBWTd1ZBc08N8ZvYNLfLm+LZHMTY+fJNbiTj54FBACrvtjgf4B2wtxjMrw
RQYgZ16rvHHszldqrSR8WyDaTPvTy0Znt/KNijmDByazLhrLEgHMPEIydKzRGK1SU6h5w7GWewGX
vVMobU7qg5C+GWWu9RivoiXyXafveQ4DlLWsVt7N1pG2kpflbPOiRSv1Ga1orWNVKm5socmM2ds1
pthFpK9usdB2lebi2wv2twVccttISS3q/8rUt4hd/CVA4uo+Y2FTL/uPVbDVh3R/8Vcgo6msaHRL
2FHRByrgHEEI3jsVAFhYxa+UV6JgLdPEEEfsTFMryFPonj482A47/JaVOjyhr+lveX6Fn+UaRMlh
U89lLu3cUSdQ0gjx+gEk6Qx0klCjuo2scZ0WPhYDFZAYSbBo7cCvh83zhiL5fflNWh+SkQM8Co4x
BfDdL8WkPrG4Xy3FieLwjmb5RmKrxv5qBSUerUNDOv8Si35wfs9iLn2hg2zqQ2Wjf70Dgxgg9YE0
twxe+CfurQNV9DZofv2A92pIazNWxL4/L3CSlhBxWaeL+z52SiJpBgNYWa1x8Tl+kQCKpr0vOeQP
GOFH2ujHFxKxuaa2zdpWTQNLXtQy4raSiwmf2GDLDK3JrtKZ/RbJuhUm0jMrkTnW+SaZwgK9evmh
R2QOHQ4lObXpto+V53QA1XOmTU9d8Cc7br1u25Rq6fIM4H9sIMSXZLXI1y1Ckri8aqmNRywVLABS
JmceT0dVnUU2d4hmF30GIa+oW2/TNiKwrOIf8LqcC+2hkGxMJ0Hv6eKppRV2oV+jPZBsJNNUcMZY
K5uR/w7qmh2mcuRceMzFz5US01oaD44EoJbHmm54bAJv7aUWxDgFaQXr7CdO+q1x0E6bZRlWxtzH
xQIvkMx7HovvXs9NGakuyK9jxodm+iuzD572d8dDWMWJhpXxEX8L5tILVT2Nw7J1tQ0C8uKuYq7W
sqd4jPL0R3Y+g4JSWOBwo/fUYZwUBfpkIyZilkj5b2NeXphGvecAfWJfdWB3k4Ftq80Wk2e3xPlQ
IJwn5KsidF/OvXFRRCGD6XUFrbiLDKihllsXYcxCnPxkDGmEhud289jvaTAS34iPBm2z08AorpJU
ZYxYqzgrQrLUI8SAE1SUUYX3sv6EcfL4Gmlr2RLjgxvzvicV/R1uJ6YNP4erUk0+EQHzSAMqogGy
rIt1ldR8bC8p5VLJNEzY/d9i+fOpWOVWHnOBYKpBWN8jRrQ/XnWpM8KYtijMeLtIgt2dz0Fzf9vF
ZGxIfnR07tN2nfopRhc1OHg618vEXLyu1UulDbx6pvlxv3lGKteqx80R8HvD1SUz7SyVjbSFORBo
gzIQIKj+RX6UtfATiT+++2VXmQKnp/wuVndjFD+S5dYN6jBk+3oa+01M5YuPSZOElmIO16U6GBz/
N7pmLh90WFFSparTXTresdvIB5+u2Lt6HkNZBzG5XZIDgc++pl+lZPRj+6no9G8MD/UbemYHdE6t
+a6U3oo23IOEBG6b95updVN2Kcl8bBaeDQyetuU+yImJrjHn4m+FE50ii9tAbDTNf4BQrrKq0ka2
IbfUCWWX8IeuTJVJ9TMHVjb3i72lJXis5JD+F+6C7+S8dcu2CqZcKYpZvZvQDMryic40TQRkq4YJ
eluV7ECDCtGok8dyqGexyAfLDIma842eD9mVDFp+S01oZM+yL5k8WM3n+mjBkdGM3P88wWUMn5rG
WUTFb9C/lMoUPjyWKa8OYHI+uF+r9bqWsMQWjNiBVedumx8Llp9QflM86HgGfXZRuf/OlGic+04Y
K6t2vrTaRE0xGlHKD6TP5G63cJAvC1Je9pmhspzv+KCblP/wyqIVZOdGhzz1y43YyjU0itYADezn
In1QI5xd2MjOxdyj9QDe3hmuTZMyThlxHXk1NwktntaHC1F24e9JpHD7x5h4soyTAv8sunRFpzKw
tzo17i42mhKZcOBiwQOLxej/iC/xyrrOf6vFBsmZfhQif/4HOKAXYLJ3m+YF8i3NMC9OUhNexOh4
IlYToBDBH48Qji8K2nKFhivZki8e5bjMPhPKfo5ZUdSMhsjP4K3Y4ChKcsruZ5NoEDoA8Wj+ulng
MB+th7yQ1XG5Tnw3OXyiL0UIBRtqKu3tmW9PbIY1tt00DHkKhZCbVvO8wMhyj+pjKRgoYr4vbRfB
lhR2NPS0zlj9K4+JCYlx6Rwab+GnbEMBFf/VrixWFJUhVlggNkfNqCK4FLKc9G4iD8NSkxbqs1kC
Oa3HGw8UptZBUVwp3tbwPn7ocf7y7GbifPe6esopgALw+fjztCrXg9VpIczqIt0Ipe9MOCWxShWA
CoD4hzqgMNYq5CXmRG4y7X+S8+4mluHke9vmpxufc0fXwNR/hxgsQ7A50TVXNSB8rTxxg9f7GLtV
N75PU8KzxJvuDRUYqJWAbxOC7mLbPS1Rc2+8hTOjLjOIGRYgseHE/c+AYy+OY3eXC54AC/5FfDjA
RI50nWnAi412MzU+j8aFHTP0SxHe4BmvYk/eHN1k6P+hnG0fiokm/n3kMILmD/ysUetnAdceQC7o
+h3aFS3zBI9MbRa+wivHk7QO6CiJyp8R00u96Wel2B8Lk1J0l4P7waVCK0lluR9h+V2zSanClE4F
Hx8Jg/52Fd7A8SpjvHMTCsxjRKxSfjWKpjuDe8GsK9/j0pzXkj++B713v26TTsbzr5jn2K0cAoM8
N6ZAHOTqej0D0vHNo6ukiBaCm/1X20qWef1MvzeuPTzgYW72scR1If7sTY3dkEePLNepub3lpgDP
jNsES3wezmkzUp0vHZKUgh92wBpPltNcxXhpLoyXM5BfE9hKI37Cyq5YbUSUiv8tv7VjGMQqyDG1
DVmdIPRJMiTs0Ww1Q0sJzZjzuKtaLg8rd5zHEsJcvib5M7wSziQmuGS/nO99aUTQ4OlMKexdHA3U
BMz+Z36kfJai5Oh4nFeJaEVmARrHvK0zpmT8Mn97/HoIFTLGXFhSesA8tiRSTyn+gb/fD3/ot2RJ
pT3EIjOJ1/lBqce3cOGZ+mQXo3qOgEC5AyZUCNn+VIT+h2hjeHMNWRJovJppEtxTayvNeCUM5J5Z
ESJwz5ZSuHfrCtoqeQNP2dxqnPd+4hGFgsYAURP1YqaWIkGZ/KDyyHHBTZm0IMnEXbYl41zdYnLw
V2WrnIKH72s+xyUBbfegAbb5HDszrpVHK6wKpRDVcxC5bjKc2q5KwQADe4uMU2f5yaGVuW6Lnkwz
LoHcVh5STTKDe8Nh5PNyzJbsbOxgIdxKQuY2V+91by6gROrwpzbGgz+p66DDUO49YBn1whpUCsMk
T3RKl3F1Xo0vOPdCwVbJAyxtRs2AvaudPbfjy3pGpq4DfK5Vd+uDPBBj6MU6WHYl1wUcEkFNuohI
cwrJ9dZLZbhlTU39g7LQA1F4B8tlKs8aCbgJFg1VHSpGEOaOEu0JnHshxDdotR5vYCLTvhQ4cbls
eHFGwDdHzzsRUmcszDT5/stryGqiVUPaYjcKZRysWa2RmC70Gt09HVtCBmwzt6iiffZx9I+FedOi
IGh8yVcOd0oloOqKKG8cKFC+L9PnsOnGFzROn6rLYXz6NFqN8G6F9KgFkGH9mcoq6fwthNEomTNW
CCnJ9v5wZ+/Agfgg2TBLJgh+itT36MWWOHtXh5m8pQVCAB3UjXWFHHb3JnRzerdVUnnn60snGfRD
afYsgbUA5cDzEQXL2OJuJlRmXa66vm1wBgwzQnNPiNUEKbAkKrJ8oncR6zPFnh+oBz9ZyTziaOCt
dNjF3QVda/54UYsvhSQmYApP7n9s5ZgSbv2bUnM+0tCx9WfVz2nY5K2oT5MTxiO8VD172i8B3dc8
1M9aOLC+h1cl4oza+YABW6726MDHVwc9tz/y6GgCnjczyNUHYDOtZgi2PInFm1yHJ+7SAQ49SYON
uEpBO2yPp9sQmNN5b0fQWFHhoXHawjdWw1zvOzalsKLr71oCiJ18zKpd1h8p5jBkXSCnC2aZGiHW
xu8NL7gvt9OwVl4Cy2O5gGTGlPS1G2wVhRL4VVJ4QsZgpcOEM0fxRhjMO+sPo0b41J0gS65kTl9n
jhf9LN5kd36pzFEkqkpXAmxERRUF/TQDgQdk+TAgLl1jmp7/TiwRrMs2qTNIluD3DWJs0Jskcz9F
oK4LsTKsNiZpEMyK6h7Xy4quXMFZX51pIs3qCIgGylBKQ6WxgWU6nnug/2FwKzIyoD3cUo5/ynrB
t3COIvCjYEb1bbO7Dl4+FIe1Qu2GIyDy6Vqq4MeQiq486Z4plIJUewlOoAx+2TW91zPtBI2I/VVV
Sqdguwh/OePRuqO/1artPnL3vO3Sqxs9DJG3z+7godcxfarU6g0fgLu2QFFo6uF3UWD/+tD7y5Bo
KRf1CtXIBZbcyAkQKHx4CgOCT7jSmJLHtBzLEkwt7roxLDAgDm0HXZRmIlFH5BsQhb9SbTqcKfbA
hw9GFZMQB4bg5vp7j382JEdIWBUKJBS/HoWMpc7SY/0i9GnteXVJqTeY1mRq5/2nTau7iE6P344K
WR9LQiY1imP1RO2nxyJSAAoe8Czxg5iHK3URakV/v6BWog/R7Vq+PpCbC2DNsNBSN1sjAtS1LVcu
fOp/LtPlL+qUzMGa94+ooGdprwP/maOoMD8na5WkGEkWAQRmHQ5+k0c9FBc4TOa0+g191tVvJ5Ti
K0V7tas5ykvKM9823SjsbYGIIrkIoMlgjWv4fbaZ5Fe2zUHGd0AiQDWepscp1Bb6jmt8HiPi7FPQ
qdrTyX5Lsvb1Ut26URlAJv2PRubQebmwUbs0jdVaOyDj14QsjA+Jn0solvfduAmeZtv1Ixw/s19W
kkZZCuQoQf8/RFnOmAT0gpb+rUtZEa+AKFMYUwaMZO2dVps9D4IGK3HXKUlSgbmuP1MGAXl6G60L
MDj/oWLTkzmM9DQrL+asY0MQQmGdZGG1ZExbaGiMa/OmcXuhWRvfjysF+2DOzpx0UOWNsvo58yJ6
AG0clmaY9hWYkkAOrVwLuQuSkqMaLTcciAuDVOQcpxwu22sHEWH6/HRsKhVwo7mFTpfaodFD6i0t
83FXAR8R8CFDf+jU14jWjRt5PyHs4MjnBgm2zl28DmTHwM29RGxyte4BYHLci5D7bzSSBvK06YWi
JDfFMoxyoYgOTzTvJT2hu27O8GT5dH2K0nlc3cQTwDYjy8b9l+52/ZLvSldGhh9BJ0ZPqvBh7EzA
80Fw+aNae5gx6LS6Ip7M4I3m1JOk1yA8NM+NMsdYDq6eWJWdXoaPkGclCvRO0WqqeaCtnqQAizPJ
lXjA4FxnvlW2OTpxWAbgkGVaeaclCClWAjtBxYFHfQi6xG4Wj/JoqqjWnIBYYMIi8S66qMyuzyhz
oRUSiRwhPR+A5aBrkiCQwj3sDvI0bqdsJJXA4sGiM3NuO8N3g6VksMBjgHEsm7PROlCwCGBWWa7G
/nSU8E7EhThZoqm81MPLAmEK831N6fzr49OKtLxudCeVmOd3zFTJVJGku5BELi6rr6TYShZtTUXq
QKV/DAhfQVi7cWEVj4wHVh99H3vimn977mszYtXvi4F+6WcfXr31ERhqmKjbOTFBeTaJ7Qfx4L3i
PbaASzs218R39SX6XTDqDTKimTvkV+xCWMBmHaBJZSZK8uUzuTmtTCYGVY+4XcLWwj5DMBUC9rLW
/VxIDBKbv6rrdQMsAeLktuu8An0o3KVgIfI/bh8OxrW3bqToDhOk6iBC4jx+ZBUp5iJIMtU7DTDL
B7PrbfYYgBy8Bh1ZqoW8CduUtxsrOv09E3JrfRQaUdfSTsZ2pMdsWa1Ulywk1jK0iuATvhrNR1ab
pf6xKm+Y9RzIu432kUnmxr7HqUBec4FAzUxizO8YP4t+QmKCauXXvCULFUPRvF7qE/oO7iNdWB10
DN+SvYklP5o5NcjuArMrul1T6IFkfMmvGX7TPvLr8gAE3xzR4h+m63tqQDkuiy/rjzrSnbAfhfV2
txsSODzvYHDcnkqwsCCivcIzo24M6EP4DDiM5LmwnPBfnhqjyNZK2zfHDc4SkCO6Laukwzk4bduu
dnbDgdlN3yf7Y0AjYIrSz2B7giAflPL7iroahkhyqMogGkklp311Ai4O5AMJUxs8VaH4O9mzrAhF
4ieoW0xmXZhqrmahMEAKZzuu5bNlc/uWCAyppQqMRV3Aq1LnFjim5tOH13OPcW+o7JqA1pogt6NZ
VgzItHDDJMgocJ3qgbVU6/Ti/gge2mWEAsY94RD9dHKnRmQMPJjBEyOAKVUp69dYhaVbaCx/N6UO
XWZ4c9MaYzivCoCTSYIhBYrRHy04t9IbGsPDxrqzpGwsX6ywfZk/87jVcnJ/76Lct1lEe/mpWwwu
kfe0InkABCJbhIGbqR7F9vAdTf4SFcWyq/ntRrqmC5D7YOkvOSkqA3h7TPzUn0KCzY539qLenSqA
u6wo79hI+y//lFF7pXLOJiVM+2allUNHafOY7HwXv2OKvC3Krr1W9Zv3DU7Bsa057W5J/OXIRrTe
/kymTp7GBkEZGHao5W96gpKE6qTdvZ3oKBDmIQITPa5S3KzKclXapX15rZ/TyvtSBGWCIbmTtmIe
BfnoS5pQbl1ipXaDVHUqQ3ypbi47v7F/Z1xr7oLkiMfdQDrePb/ZNvwZN1Xyk7uWQ6xKmZTrvyNm
QdA0nCkctUtJx491PO6kYPXG3qQURQNHyYmSbhp1U0QSazh88JIUjbSNR87UPT/MKdaciCxyE9gT
0mdIVfsz5VzyIFGQYBHJwSDcyulPVoc/D2kfedoqD/8m6xwC6nSjTsyW/kE9IEBDkwqOvf0xhLhw
0x9qgJ1RseWE+tAC4epVgQrqhedvNKdgB9Isa1/Sqe/uIE8CfS3fI6lSt9atvxnvuUtphQTzBT+X
fJBExWQDTFELTbjRAWdOKLL7b54ZUfY0ZfCc5m/wvydR7Gt6PhhslyScpU4jAbID+vCCBDQNvjJd
DLo9zMrSJn1krYXlt+KHejp6MgjhwW9WotrK65hAsDvs5FKF121jsPC3klgM+tHZ/Npve+SNXOq0
s8hHmyO0PD1+Vli9r+YHb4F/gcjRgw742kpeg1qY+MVKEEl8PUQTXxzEZzQIKeUk3hL6QTuhdQ7S
hBPsHpJ7w7exnGPlzmf3rlBWIPbnIFdvD5nAwy3yyzil0MocBXO8cgRZf1HBIMqvzfblP67lvIyE
vj3S41h+6JsQigTbOQk6nkJzMOQqt+ygC07OeMnZjiha8SYtPYdas6Kw9rWWGzdv3I8gMZDUQ2el
BAoCPlPu2A5L/viuCyncSNvKZSzvzyoCzALB8xnbEAeXrk4CBcjsTTxhBouIPWB3DW+aWW9nxDRn
WtIYt1GBCj6CnyHLY8ZcNRdmY8yhrrXmEO+UZwgj5/WzbDGE/N1c9/dAb610xvi0LVMm/vrYYlw1
yg8FQwuoQfbNyWQWCBCjeUp3RrV+2GfQU5dQ2tPuOi05sl/ZDjSvH33hoA6tLIZEFKui0K/JHUeJ
8RlzVcSDborMyzRNBc7eyV2+mF0HTMIbkKXeUtRY9U6P4zKRbCetRWOg3lIpz6DctqxayxgUrMEC
V9QH1kReAg13E2Lrw3jFR1LIibd6yBrHqbDmDIsG3tVLQdodYZ7WV6iuPsmhrkVTn0RLoVRwckau
zU0rz4UO1aZe7/3Y026VkFLkj1t0d+ufnaKljBOvw/cxZJ8O7wY+JhqV03wCQEnhI5L+QUpo6n90
dWGBbMlsaECkdK3ukOEgsm64pqTk1VnPx3ICJY3Eq1u3psocMjgfA3Mp4AH13SfRcw/eH2uI0MW6
cvdl5jr75VQz3f1CihNZzJVOfIZ3XlLFuesN2hHUgcUC1UT1t/+/pi6SLNS/PKJmw1Eme6JkbEFy
yEOj/MsDvsUiGaFByExVk7l8NFmTnzMxh8wDmohWhHEPBZGq0xI2mmHYzPBzbWB5r5c44ytrd3PW
fNFpgBYcQHa8mjcM3chY+lb50VyqMY80nwK2BtjavFcnIhH5SEcxFqTDF0JYo1ngYC5vL1cnHp+l
a8Jp5eEDM4lUQsdMRoCsF9++WJFb6ERipGPpgLTN5e8zZxxEr4TMAEaIfGFWqX4dkl7tsC8Mz9Ol
JG5y/VSlmBz1WgJ1GcQop5c6c8/hmWn6PJlK8Q22revdafA29JW2tRkgTyL6InkQHfqMYRC+jtMj
yDyzk0ztpUnFIFLxoV0x+kHeugNQb6zjTtRCp7i9hJ+IVd+vt8O5WzXQjEjcNXCfSc5XtJCrNF33
pd3FOdUVfOScbgegey1yzVz0rwym6+FyPHyszco2RhIZwq6SDQbouxOqmFTnVuRx9zU0XiYOgeDP
85AyBqNXORr/Rmn49kDSUiXkuRadGoBUFqvGNZbEVWkLPHQJ/Q88z4iUykMLsHX+XvdAMor7I0qb
q5oEt0gvGmxoOxPLP4Rkwn4yhfm9v/fuG/U15s81aVzM7K1GFUw/U7n3LEf3d97hQ2Mq9Zj5WlvV
2+VHYbLWJClS7vggKg4PDNoEXiWlLuao67cb7+VmQn9/kQ8kFSHavf12x6BgPHy3/gOcZnCy8RJ0
IZM8D3uxsKVu0FfLVq/9dCDE8owukxuZv9yAWeqqGWg5vMYalWGeRVZ1XkbQqotCPAZVLhTZP/uH
CrapBAFjxbZHHcVadKuF6R3921ykiibNQ3SiRdmmZEJti9M4g4Y6zG1zYESk3sOuktBUrcKq6Br+
OU6Uw8MDCVI0x5Olx7/wBCzq3vtbSUHMlgrBOCBN40xou1kCvaAYpQo6K04c8AyNEtlbRaV7N5TF
eiIJby236g0SjmTnneD/Wl8ngetQu/XlqCLL3xXR7/BFGHbwpiTSwzO6YC3kAPKdfbt1URXhw13l
pRPwwhuFbboWaQCkIUt0mP7xJXVK8jPLFNHg29SwUjBEv1fwcQsYiCr5L/DLSpugyaohOq50Fq75
Q4MWPmLLfvRvtYL4lwx4ieaQxZVClswbey9fRgqCOse0N/24maP2zBQX+wEOZRv1zJvZihb6gwwQ
dP3TZu08zjRqNv5auQj3H1ZkihMqlyXzior4KLeCtNqEfb4NcwfbxUTHtGq8w3zXI6P570s5+j0i
b6pxzBsfxd0DvW9vtxfnOOhs9flMOSpM0Slm7L5ZUiJa/u4jJBA2sUbOd971jpyoY/w47Ri8asqM
FpdTE+jgikobc16dWoGIkqIu4lADM2s0dW4/p8wp11vvsVidwpBogMpSLnMY7BHX1fi5bpBzNxfB
8FfMSRqDIV2091mQNkC/4cuF7w4G2bouvGUQJN0rd3Fo6ICmC5teEB1nMo2iu06Dme7/GZZHiA25
LDph58ZJjuSdH4oLe7D52r1i79Uq0xOgi2/BcLf54NpWkJlMERwiCjoVhv598pTNWy0Mm19I5AGg
h0ynK0L7nQMq36jNatcgCGuR6u56P3UvgSqlUHwj/sbJ0vpSblGuIZuoHRYBu5G0fQSeOMx6jZJg
Qco1CT/QrrUv82IB2LfsqyNfojJuYYHW+zpNbcm0qbVA493DHzkOn3maKAMZy8FX+ga9i0+zMCj7
GeuZ0PXSav3ZYxw176JtiM7kG+laHvEhGwyKfDRvRVx8KP31dC7kD7GyattErGlZq4wOddut1zGv
QYaktm2qBlrKshuVYsoTYJLcexwPiatOj7aMxPE6IgQp68Y/OsUpm7g0bYaZ31ANYWQDtzVzVM2j
ghhJGK3GIZdB2CWnW/nRLrpBMMUJ1msT4N4PdIJvYpMBCNPFiyBZlpt46oKbl8PqKyCw+pmipl+Z
IV08L5GcezoEQqgg+fRN76VtubCSWgnoQNex6cr+oHcvzU2fiiHfQnm4ikxv2X6Y9PaLYeA0lGZ2
esRYAo2dHoBb4atX8fCx5pSGrD5LZh1S9v6aOjbjG4W34+b636r2XOIcM5tfgndq4ejQrPaym0G+
Kx2tip+j+NFfoDISUcDDnEsHhC6cfVnOcXjuCsJOhb/b5tYXhlPSbXEMoSnTc/RKioWdppWB5yEZ
ny4NfCyZILWB8UnMEoOSxYr/7/5UcOWFgPzfR+exZuDl8mUxjNHMYvjZjMV+ZE31kKnRgM0NyhjM
FZ0AtBVNVsT7pgLm2QTo+ukMKKm+6MVgsUzQWSg3KnyK90OkuB5NePU24FWb7mIaoJzZT+UVygkx
H6hnPqPJaRAZ5h5yrIz995qqtL49MLBKI/aX5537IX9QIv0xA/R401Oh07LrgfM1071Uo45Ax4pr
g3A9z+6cFMX0nM1aqDP+l/1ijQg1nL+XcmiJu6miTY+tv+MDgWh04YDoVVtfNl9ROHHYTc/GTCPF
jLc+TdWi17X5ZArpnXRzPC723+DcTGYl4ctz36LwwGr0+l+JqblnGCkm3FuL40siu/xPxbKRFjso
yIA1xltkp4Sjf5YqI/mR+SBXnD6JT32+x+uUU/9JncEvZuYboN2MIp2S8e3hvMqYWfGOvJYH9vjR
i2ZpEc5njDmjjeL1iOnPBcj4y0kc/uhOCSILs2aXgsHrMvKcx/YrwPXy5MGfyG8cOC5sOLkvU2Si
82U/bOt7hYWJ8Dv7okIMyD5j9Xg6Oh4MXHYJud+Si9vvs9ZYYG5zYBtV/Xt0xqqVPKH3tiFh+uAr
5c8zoa3XB2zEa17584GDWMiGHnhSzwPcVfP4D0tdcKw07YUnADAa0t5Y7STIyufBIZ4q/66cOxlT
nYz5aROOP5beFD0K7994jBBkYGlGWPQMa8H5ySB06zE/J7hkvVg3mMBflVRfk/YGOKPAfDsi6gzj
poLmHSqWrPId80ZcNDiXFjz3kVEjwlPslC/dPAmGVTXNrblQrz/dKwrfVkwKhuVVPtUS5P+ygJIM
/hw+KJH/Tncrv4iR9+Iv4z2/gdoeqPWSjF+jdxPL5E1PBpDT+DbaidvN/rCPBUbgHmnbOIkbxwgL
OZG0Eli4y4EcWhZGkVa0f+O6zo471sBegMESAnxpsf9YdKQChmGKn6qs8X9lB68NAmAxKYKg9VS3
McOLaM/QkCkK1IG6d217sbzssVYb1ORTm5BZHqgIvPUHCCBggX9zhGVNNtLRzIGqkIqO7Ozi/ZUO
WT8/9ckXjfI/A2Xjc4YOU6krXSFhEyn0X3gq8pMzddKSgiGlXm2oPLELk2jaKH/gQ6lsvXYFdxIb
ti+kOiSncuzg0FmJYo2W4q6QOcWW3s/gznQuuUvcEQRoww2/rGTfyhfWLdeR8v+FxByve30MfQyk
fKzaaFW6XGxVgfhuVZjM8vBS4Vwq/s3t8VxJ12vvLfO8OO+NkLc8NZ0U+I/TeZ4jM9NRCCwa83Kx
S8FlDbhY4ILfigk1dgl0LZ8m0WppDfzJ1rA2/ogeKUfAZvZFjNPOw9L9USrQh3MUQTVsFVMZEmR7
4prcxw09MU0x8vSce9d0ScxfiPGwrKyXSOd7EQzPcVrMIq8pKvzymXxMxGUqmuLqAYYca3o0ZuEm
zdsLdp6Z7shI7x7dn8Awmrva7rR8y3f3kIPya+xwMDNpTQOodHuYWBCInuMNmwU+ofzwt02CUYjA
Syt0B7PTr4H45f2XO0a/ykProqDP9bTRuo+UKfhNQPY/qp74g9Wcq89jWg8DdQ3pFZ/iGBwBG9CD
8YsSZJMvhEx2QrptDW3owGQQILg6QFPnhHuHREZZwfrCPN0/xtDfIk/iCyhVTXjukxEF926WgTrd
i1WnZhbxn0n9rm1FCR1A+boQXl/V7HMe1NDplE1KPyEYOT5qMadvqPXnehUWPAMRBSjdRyXsrGsa
ueavYV4BmrxDd0enhqeC+A0ctbjMdH9RmRTx9YI0C5x2kiTGz3DZTeVZ4ZfP5uPDxiwbLRcTd/zD
k/bEZvS2rRLiaSx3XxAlqWPtcsKi9WbKDLbWdIWYon+0eTU1tknvkzCykV1IQDKJMEBKwvdbyZpI
uFbqGJOrJI/zbTrAO6gnBXOzN2GLchfM2+qMOu98uXHw+w/WnIaw1HQm3IzXURwwxP60qfXidbJh
ygdJQ2UBjWXYItxJEd3EuRIPbj+dBVuupgK2gKCRjNGF9LXFP0Rz0GazjQQNM6DKlFuQpxMn9t8r
q1eNCbt6CD27/A0HG3rZjrK/Y+kgYZwIPwhdKrmfz9y8rieA7V//Q5kPdQvYSO5Y37A3h8Lc9Z4i
BUy8jPapWJ/AV+d3IV90dO7yJQcQQdfUs9UCDnSQi9VAho2J79za9SB8L30y9hYSYAKKQhFJTwZl
PRlAljYfPY9r/GPqK9SbJShHrNPzK0DooGEy7d6937k7cmUtVRT398K8e0ikWU8Pq9flqgdpJF+5
K5R0MP8qlujFSFAoTvgrQsgsVTuk6bA1mYQkfxk4IGskILqiqHqKHQDOTpMVODLhYY8gTrUEjubO
rVCObbKqYm/soRewsECM3w7jUIHTBaVFP530dioGWkn/TIjfY4vtXl8YNQ9ySgcQXrY/QM+M7f8O
fuKZ87mnXVrFUI1uKeVZ+zwAdW/9h4QLGTadwgo865dt6tan3iCW2dE7zThSRdHke5BhL86ANXjE
VGmI8gTY/fHvY88JZsP3woNqZmfy6lQY0+hcgIDJLn2FyEmU7ds4YMCMzdygfXZcO/riDgOEMMFU
Zk2tVFA/AwDRzNKweNPN7GtPGeqw+YtFWob1Q+FUyK3RPErEjUGatEZorPfjb8tb8Lf1HGS/6es/
Z8hMeVjljRkgWAE/eTa5CTUCdytyU+NJDbXclqXiEFSlp7TdZbMYB1j+F6aRaXk0G41dtOYWDgLV
gSL31xLvUHBD9oXafTp/wvuU/R/IldbU9nvBfhttokInULRDK9yTxa8u/XUCi57VVtN8mIDXM4Ib
utoAgYEan/5iFqrxmjRF6/FApb82v8bJntU0S4kVUm5K6R4QIp2DiETx4zxbMv2JTS4or6vNUyfu
chLPYDM058z+yl8BNqvLUEaN8Woz4wuy3Kdje9TBeQVwmCARmTSWxBF0KKSSt4K6PDBawl942oP9
sCNZ9mR1jkRh13MXfHkLFH1Suf7zMeMe5oQGmleF8aFTHM1Adxl7Y8iKlAfi5zL+Wj08awxxvMOn
4osFRmlJ0G6RLG8m081aSptL1X7kMXR2OKZrinJhIfhNySMcHrAsvcw2ZHccJCpXnP2g0+4rsowf
h76+R3nnBPxJhcc9CMeZX9QDchLDe6rgzvYBL9GDVQ03U0QMLUMsJXoEawZkYwn0Wd3L4vYqsowQ
p8k7s9JMcmWzYVOLlbAL0iq1jnth6bA1Jn6raYh0emEHFDQvGLg3XWWDYVu0MZxK8cqShhcxPkxG
2Tc1Sd6Q/0CQb+Kyf6s3HSDxBC4NFF+TQ8E97J8949AnA4ml+7uoSxLuJ0fToGiJz4ZRhzdUtrca
ueTNsKFFouxd1SRwMmC6gWFjMoccQjHvziwCfpqLPqyVZsA/WSOxA+/N+l7mCkb+Qj1gIGbW/e2p
c8LJAw8kUf0WbGBeqILwYvxxzNemcFBypR+tk9Znv9NpihLjkqaTpvATJIcGWIrJwK8md05N5yar
DDYQtHo18Nlpq5SWwYfXVuvPSBG8cLM8L9XfTlT6vEuFkZPIbKQUInUE6V6y5qJwwcEcQCYm8gtB
mHIcJjYp+gcfO605VTMv+vnq/Oif2MkMCv+l5p7g4QPpgQMexpb8dpP08zrIIfB9NJSh+OcwW7Qh
TRDVvatyLax2biyxeFg2L+zXi8IYqrGKUWClBTAartGXFKzqGQ1Q61KVhpuDwvJAfiwm1MRq0L02
dXhWMBmB8DpgHT/i/APP2Q6wFqcT398+M/t6T/Wm9RMDPbc/Jh1YCODkZrE9e0Qj5oZv2uy3wN/F
hAx5IEaQdYSjopEMw0jrM7xQOC9wgs0jw3CjzP4Z0crjrZlL1SjKJ0CCHigG7eZNf5KVptDctlay
beZKj6/klVEMLdQakkAW9Uq/OzoAl6mdo5DI1oJr7XO3sIj1l33rCNPdfBsF3sWoeZoli6yyYicc
wsV2Pfmqv47HWxDx3eUUQ7hyaBDPqi9Z9RO+n4iBE94+29q+nH7638Nxvu5WyKHw/cXS50xReEI3
8kUgJhzYDilLZtUkkAjjTwi9DH9bcgZoiIGo+jqlxRnRbbwWC9MPivXEIWiOKWbrQRU5OptpQKxK
cDfaGJzcxtgH/6gvs8Rolj0pepv9yjA82wF73t+pRMBY8TV1ENX80xj70YwAOnRRJGMOag0eOxq1
6yxaWk/nUk6yaQ7FlFbT1+hHKVNb7O4dJMsFlZi4XcgnCpLk+rPMzSxSBd/wQ4S2WuFJF/2siW3S
Kj0vmK3dmrsqOZ8XH3rATJvqJPPbO8FKcpUZKP2vxj6CdIZo6p9Q/23bimDdfN6CB0iC/Md8JgaN
reGF04Gu/FgNbB9brrJMG7qnGCNAWLECAIEQ6ZrZGgMBqoQgiYMZXGSmjQN5UQ5z8jiuu1TcvFl/
BYWft6QTO8Jj6VCw4LQU26Ejy4IX2VQPPntQUpZhO2e7noVQQ+7UE9EmEnJle9jW34RSjUUB4nyr
A+pUPvQsxV8BXSL9Xux+M8foRatbXAO5zd0sCIZaxQgUbmTirvSi4/uxKDWMthhhZM3EH4ishjRb
ckHfR/m/e6Nf6yUhkWSHnVzIbTKgd3LGBDxOXr9rMxVI9dk5usdHGax33IOZZSYiQ7Wud/Qp0ylh
26Patnp49gbUO6SXXJUSOuiCCedlYQ8bG8bMVoB3vmtIOxc3aWDKCizK6ko9aDoWcnUljBMQCerr
bIvGr42Xd2ZRgfH2cM1yWPEFg4IGVpJ9GkVTRC/0/cyg/e2hlsCg3HxP2n2IiRI1LmJynHwoNfO1
DsMypFoWvcOIoRlLjCfEcRvEjtOMvcjAQ778QdUAO0tkrhLowHmMl6k7j6muKFVb6uqzv5Bna0f7
nmh1USbXHRqsRC39ydRw/s3AZCqL1bafGVQPh8UFktcS6DwAT12AQny6NcVHcCoSbN6/CBThmjFN
DN47AxAVCmJ2gXXAf0WIlEJZE+1esbWZSmHmeeU8MD2zQKKkoXyIBWpDcLV5R3U9bCZfIsPMlQlt
mPuksQLky658ZPasTsE5Pxcbnj5VcQFi9xumoHIhApCXTVAEB8ZPHgErn85+2v129519KHGi3oMu
WBHyGjl0GG0VlMiqsDAtKxqzVOWgpoyDcfF5C+AG0aYlguhnB8lhlyDvX4n7aS1HfaVJEbdY4dUh
sF0BEbuh7hhUus5DuP0L4JGVp/3xw79WBTzyN7fD1b28/9d+3YIUDybIiIjXXxxw2giUqfkXRlZU
D7RjgQBYyyu0wwGj6oNcctlvp0rvZlGe78TRsgVL9Mc3JDaDH1QZ/y+A2aGVOHAwYH0VkliLCMAl
szoigCUw3yxNFhbJnATOuP0qe4wsH6+/0I6b7Ci54X0jytT4rITFYTUyhwqhvDo/WNzO7Cgf/4kk
iztW51CSDE/JrHLnjuJVjuiNkR4dXkW3ZsRIrxrbNhYtxMNMDz+XXRCYwrghG90jfPYDx/docfa8
4fstp75dHUme1LK9GusDm+PcBdGsoknaeiR2Zot03hwMF0sP1ZSjRqlC+WJb36AKs6CreRKPh7je
r+3NIyMtazXTcaGX8gHePgqWAwjID8ysVh4N0FORn4/fWSYiYZscpMqVuL3sUICJPDJjdNxhXWAT
glWMYCKIQ0pDuNlsx88qnBoanGV8FH/CXV+SK4l620CtPev3InYwi6Rsbz8aHS5h0G6VRmkqNHES
r/rYiW/+CR+1kgRmEskX/mJKZEY3c6F8YYbScWBP9KsyhlDEBnWGgez5pVm1Q7WYe+8mBxZi3W+f
KFssXhd9Kk50Yp7Vj54a/+pCaVLuWg9I6ZvZ9jf9mbWk8zIxmroraA2qBim72hwYk7QTttu2hL8f
/GnJaSEHuxKyJK3YKXOkLMoxqO4P4Ff3iKV7IowpKshV6hv5Rn00UoY13EhF2b3aIWii2me7X2JT
zwWqW8sz5/P2JZk2qf6uFwkMedfTrcn2kfS6gcGtIqGVF/VJ3oDTVR7AIY6VLEhJiM4I/Y042EfY
O6JS5wIEiudXg2HgNx4fXx5BnpKG7YP+l6coqE/NVkP42rw15kKw50EMCMZg8c2MdvJowVGvcUxE
2LSQfOH70DJ/6IRG54EwJVvTPjZAyCLq3dAMiICx8S00n1zcB11rwd93hKqOhVYmdG/M7yQslagn
LUo7rEmoMPURlcY/2q0vcB0/LgjuIkAwuK90HpEhbXgyPzYGJI2PUT80w/6Rfq/VC5Mgr+U9I0Rj
ByQLg41U+IFFApq7UWJecKeVtKmcjt0xvFtH9XGqUu4dEmAk7DlKH2uIc2+9ng6N/f6Iw3JkVpfr
IxVHcVmjPhvwYFjxuet9DtG4+i/Gc3WtYp5SE5SmBBP9PUPDJOgoigXC7/RnF/FkqBlodS5zG14i
c4riToEDLoOIhDJfYtYd0CTflu1bmzXyKxPT+okPgrwZNkSX02ewUUTn/xZQmUP1yaCwUvOTcO99
y/rouYXKxSkZpH48d/+bsI/mihbqqGAq6UmAkZgsB3BjlW6+TOkfgAT/rHke0v2Yov34IJRB0Gd5
AQy0zO5bpjzIUE5UdwqSSrLrsdYHjnqd0oRHHQwGnL0RoSdVXZBhHRp2Z2l1Kvt2A/x5b2EW9bsz
kNzZqyyTWnV0EpHdLh3t2k9Z3Uyde6hqhEt4Y/iaTIuD479jkwAWs1jdYVkloNdfpVgFOb9V83Aj
O+h73xQ4UY6cUZy31MzYVF+epOeGg6RLKpUpqB905nMaanB6Rk2Ue4mfrB9SazNBQgy0I3rQNPZM
xzvikd4WDoS+ibSb6P6eB3yNkeMl+XGhoCp+yblbqcQ0DYHrim7Pd4uaqYkoCBB8EsKPsAV16P8o
6zNaFAp6hkHez+T6k9LshHpsT3ntw85B8Uv/KCA3Rbfez3Ypxxr7+JEJV+XwJVTMccMvfWvCCxFR
k8oXcgGwM555dTvnlc5Vce6o7x6EJbGvLGQnkG/JAm79NRS5ni7SaQGNLj22OzseClKrrbanFwDi
jKTLgqwvdOn3HfXzIxCi5/Qys+FshU+VL0gimdlWbbhNgZWr4Qtw7FB2hVdHPQ9svn9tJO1i3dE9
4jryLIVsfR02i+mNMCeraO/YT3kbje11AFOoEB/q2dcVC8zARt/tGpIuNxqvJa2mq5lBtOmy/4at
ouo7LUDew2LkUothkljj9HMX8qpt2Yyr4QAd+HRmNXtVJ3V2n5f4Xrujy0ujb00O6POZrhj0KOfP
qmFHuOXOUYtunzuYYVBV+iDqeG23NIkXY+XvKQYc3zoQSMmOZ/LaD7Oryq4mpVjyBt/P2Z4S2ihY
sYA7L8s1cWESeQAXRL8GQlHW7ZydFg2fKWBkpS2BAoMuOTexhLsIQiOTwYChiOfxgfNunI1RM3vT
h80lgxL7AhfCvvVvFScS1rWdsabU5dScbEwoKhyS21ok1+wY7JwoecEZXyXjk84er0DYLUb6c4zR
UNZmZnm3ze5nZ0b17p4QDYRPia7ue6HzT6y0LU7fbHgSWIsaV749sgA6gOi6CsVj+pnxc1YXMJht
7cwpekB6bTIdL5nLg486PkRvb5QQQwsuPm6904IH2PD9BPgWLyNMaEjpjnOXTKDMMMdwZh679hR6
g6D8x7W89cVOZG7bwC0pcPoZDSSFUwN5iBJhnqMVJ0nFii1iCHv8/+SIFpdUagFvcmmUGcaDADej
Ns/FV1vCmG4Mu5JlnVDqUms+ZvUjVJxp69fp9zctyHfXpoYNBz/MffN4iIF9kgHqbLwYHjdGjdpF
K6TCm4FDqNfGKfReP55w93RwMjJHIQhgWffy4XyMiws6GzMYYLk2iWM85HWQFZwkza1/iCCHCWMx
ZhVqan9re9rbA8xTave66HoLsrDTuEF7i/AMhonsMFSayHcCovMH/CAe+DgZksZJskWtJCwjBcnY
pdj6hHdncD0q10BYwBV7nL/5YI+E4icc2npz8sQpIaM1jgdvk9hzELNWVX+XbZGqiMjmujWoMRO0
zEc1gAcJdJTIFsvJn87Z2iTzTtJUzO3Pvrmx3hygnZqMJtafKqtEfQNbQmjIyfaRnkFt2utxY/6m
7iN/Ltkn9wFFFYb6FsapAKQ6FBsrisXIEhRcVfqIdxDqgWzt3+YFuVCp/3HuF01QzDznVKO7QeOn
9L7Hq+wjHxS+TmMVRDscNY8DDYBDbNRZOVUlQoQtgflcHyOEfcMe9ZBD4VHW9UzB6Ss/7LMuvoH2
4tnwunORKpzjFQe+nVZI33FbcOdvZxJR9NlWzFUrnwhNtnN55hsOgnZ6r7Q2Er9Hj2v/IoCiekaV
X7mvj9PFvymxhLzZHFPMESgD4vecmLcBzc6nEf1WPhySGtU7uk7mM/fNKb3DDQtDWIwjG07rPQ7y
10N9V87p3zkVDnyav10w1WEqr2zlBPvTTqnenFSsDLWmenSYbMf9tX1/04TLTQCoPsIbjLXjRYPn
QbuOZP55088MeR806dbsB9kumTua10+RghCLO/cwPNA4ueFINhnNxCAlPrTCd8EWaWJGsfSlfIPy
tE7qI2jyI0r6KwZAMnJNspVwa7kyPzi6REOq48Sx6sFcstnnjsahTnQsz1jGqLkWRdKBImq33fFX
SzC+vZL35sLB6BLBpqPK/Sg42l9h8VjyPd2HK11etfP1OdZoEwpH/APWTfMw4PaB1n4VmJdvuHT0
6mP7XYLbURHmB3ADxUWhoUXwR6rUwjT7YFOBFAIASbMr4QokCSztcmjgIBi5uUR7oGDPAX91cZrX
qrMJr8F5XbJqeCqDVimZJFYbcdYpBPUFW9posxPe/X3xmmHYSeBc/BxaNxCSk1PFzq8ioAf2DQ7b
az2sEMNd5h+cr5ZyFsyQoZBcGg4xHP2rCsPHuMnzTAlY5K6clxx+YiZD0KbXh+lwO5aDtehXoaTN
C40FaKA5k3W/fMGYMFExd3vVWs81ouYZh2Rrw2X/ENp6shPzbOb8erovRM4GTDVUC4Wnvq4EjyMr
ASBm5bmdnjmTThoYYwi15cmLX/HMIc3AtOA4a0hKOSiCMvoV8iIBvovQpPK8U+E1LV0QsgfZtI1A
9WrnnynUK0oWlYEFb5cSnIXekTNI5wn/kcdA9qqnraFHXJFoZFElQuK3UCunaI0EJmaETgu8xGgM
eOVfPLjTCJEJZZ2pzPGrf2Ady88iaNww6MWXHxDfp1g8LKaRTaY/uof1+JhES6w2yvJyttbotJP0
Flh/s6mdKBhWnodQ/2TnEmPHK1N3WAFLVEexCuM7wcvS8DXqlxUlNgjZEZDassVf7UOCvptj3Cf3
zl5yF3Qc0KLKg3AmqIQgBhfQEyxw1JqQQr9so68LohCl9YKy+nl9+QrQxBEnHWCRtR/gxCcSklOd
BkaGq5fiMOEfLAFnLV+7yieilOgCkmagXzCMGlrCCvr/uvHq8zzffZ82KEkxUhRqS2MzdyYR0M3o
V9RgOzdzXvgdnUz80gl2Sz/gwy2G0HbiszsCu0fbg8mCM/6lR3xDY9uBYJCQM+rz8FfbIvJmpC3W
UA5cdbz9NfAkktGqzqNpYpL2MPkdf7foFoLKR6Y7f0vOKXRd9OTI/9vFTy+Z1XgE3Jks8X7AB4dh
28Y/WwlZEuZw0DiI+CjdyfINohpk5PLiFoSQnFTt8JYdlYCAQxPmTRGHR7e95xkILZJAq2xgtv30
9YOrfG/b0VSPssWLxqIoc192KjsMRsG1P8cuIE+6nRydPScwL6VQXt/5ywJ2yCKEi6DXzfCXbLMQ
KR4ClzYPgyg2xSAROQJl1G0Vpd899oQ7IRA19TJqQznWR36qEHFP5vhJTSmjMfi7bsRJqBTG2qOR
E5gDk8AjAOqXhyi5rgGa40iaLqdbAGZmnu6tK7+YZpNMmFpm3R8Fmf0ziRYnY8zg0qSeTBGo5MQC
BBKYZy0c7+2Lc1WBL+UDrw/Uy1kY6ZiQMXZFVZH0cFJIJ8UNEvwOu6PjnfF3mqrukbIsK4hoTbaK
aoHse9HnHNTqu9+w+4TBEyj5XIfL3u+4YF8WMgXkRHLlOCArlfWgbHkzT2M9mIFx1zELtPE+lC5X
FNkaNDrKWUQ4Ti+RAwo1iY4PAcxTPQkh+EMNUq6GWmNGlu3BUR4Q2ufS1zYKFY/Uc4yHxdhpD14q
U6zntVNGFtVHOuemcx7HRjgVFEiffFvaBFguxgehzVN8U/fN8SVPH6ZaVqAL7eYUvOVHaw9m9LyS
Taq6sAJUDnmc72zkgxPtN8Q9Lix2TTFbPbeTRfdpZb8LjYNB6qjMbasBVPClnDwFCg5bSqEiLi8r
jySln+s6X2pU9IIjbsLOtCP/YeSjbNqjqy4zQZRFXaEcIg8ijUQazo00aDJNurM1Ptmqn/LQmMAP
XV6i2KN6YkwOu/5L6haZjn9co3TjZXSGR8hQAZPcx0e0Ddh0rwl8gqel8QcjSDwbktzV1Rm6hoQ3
uxzCNCrUdzmCDljVKG84ZgQgHlmmzsgZisPnsWhLCOU1glVQwm8HqSC2k9vANXTgBlUra4MDuei4
D1QC87Ux4S1taazRRMWGEZ9vSPDlsLHIi/Cyc8mAQ6JpiI44QPdhpmfT0UOfriUp2Rcx3I8Bv4th
z5iM3cs48mUmNotAVD49Dr9NQY3OygZ8fsag6ATgTnDKo92XwPglq586xcGeL4LElKhw3v5luVbs
XMBv7OzBWyTyiL9AkNa/c6Yj3O2T9jPUmQ236IdYw1YIpZjTUm1R0fLvJMsp4RGQF4A8CDd6DnXf
FuRYRH+U79wUmTDSoYOfuoto5fcuErvkiCntZs3rloosTVngvirr8s7M0QAmyHEeivGJvpju+3Pb
aEv4ZEBd64ApIP+SB2n9pEX9QoClqEPXecMbViq8jHWVrlIhkA5Gs5PINGFWhDivuEczs2ENdwct
VzNqoi942sEOFWl/h7kzSWnCuKft528lT3w5ONnNR1kqkqfl2y/68dmH8WtjMjfwNSVIAcc6/N+1
I2nICHUTpuCmpgb5jKFwPj5DbE8JlT8CuwoUcd1IOc74oqtn/eK9fHXX2L53LBno2UsYMkI/CND5
RBXnQUmje15sKXfEZ6EyAIvqkUPUD31mp3m8XhS7k9etzTtr8pgtL8yWdfR3xeBE+aVSpEAGm66m
K7j3QljGic7vQIlK2VmGg7UqR8ywi/7SqalanmGenQImZGYawhW2dD5YYJi+K6bcmFpzlIwIMeVg
tR+mEuDAqbGT8Ad1SFHGrhzH1MVabd5mCNHM87OUbYUUopIgtLvonEei/54I0xwWZx9Ebkee/SYo
B53jHWceMrBNlFjAoTKL+YAZZ8mgCXmu37WTg5U2VskgQhoi1GQE2vsPXSIHfAPamG8950xn1zFJ
pSpg0PtE1wN41C2x8hYL+MtoakGB7KukRhFt+Ah7W4SFuLgcT8Vpp3qfGot5B/lGB4k9gKKha+QM
YS4GvQWLWgXloS93JyJPJvJL7DsaiKpx3HuI74KQ9VoSOLC4EkcYOGDS98e4yW1ozqJ5P2MmNFYr
qsa4XIH1nvdyMoVH4it6Fg1iXYbwIf67y2SrWs/YUT/zvExIxah0zRcHgX7QQuTXVEVmIl7iaTXV
SMKucaIZwTFCImFo70ZCXxUszV62USUExg2cKAGpFDSzlGzTIsGL2mL/ULfzJVdaeAG64//LbI7R
gq7ZM5kZ84Ogj6xM9czxCaFlKPfrQ/EONCNRYQzGwNe5SVlX6KK+pNZrbtGCpv1uf7cwZhbd0Gf0
qKx+d2p3iLoUfxdVCrLqhfuOoEMGnUDfLuf9d1QfgIVnZkx5UNiflqsU5oWg4uOaa0gjcuzgJ751
IJ49C6LVYEsXp01af+EWRqfMavVLcE8z2MOKWhEVzBvDBBVbRyu8JyeSmi16AuGqquRiv/wCjWj8
RZdrk9r7UJUDPy6ZSJ+tVIW6u+EkLZT4N/0nOy/bHYYJJih1TEUKOMmogyx0zQO8x4tE1x7l+VHm
xfoncVc7AT+mVCudrVBui9bV0nEtkCfLJT5ZOMz8Z3NjakU433NC0zGyYJFagR4s7qLfjZ256uup
l4F0RzU0xHYpz3utbv07pPvQMuOO1hWBZmtnYv5QkBvBQF4EFZ+y8aR4JunDm3At5mm+6haByuwl
IU0hg/ZxjQUXHNtiN0CvsPmnWT/EvgHieCUCGLAYRuG9k8cGBgmp0N3lZajDrLteJc6Goyor/hIi
Yr2qtAmSPkkiFp6+I9vC5CtR6DmIpUH8Mw/qfhBHYQQKKAfNU841Zc/Y/SnAapZ+i+1M8XKGn6kP
agmOVskIEWomtNHdihRBsuu903zyLaX9e4Yua19kwU7UOMELg6mR6I2KhmAXX0lkcTbfa8UZUtid
bJ5t2r+qURIigaIVy8YBaaGwCclySH0ReMnNw2LJ18Y2YD1SHMi2a8nSH4rt+LYiQBys3ewh6kak
+tP1x/UL5sgAmKxICFv8zC0b+dSBge09cj6iDAkLk+MHAyluurPnu3OMUPlvhr7gBj4DvmiOQ6hA
oqxEpOHvjV7JQxgVMiV3Yb4qqaEbIr9abCom++Ks7jh7nDfsK6yJ9snQDnrN2Th2yF+LH2wjhmln
uOU323a45IhWotWX4++x2Mh3iXnL5FJekNHp0W9mZSGWnAOML3dfyAbJS6OVhRFRQ25SvEsOoj9K
wMwy5AbOM+Z8qa9+re9eAMUaGJqQdqJNvOYsxHyY0YZNwoQc0CtSaE4pMyXCgyCnS3BS3f4FCaPD
P3FH6ksAw4va3uhdnDnVNLDwausqC4d5Ni5mPfAvqyvf4XN3oIKN+SwhWQTJO+TdWrmGxpp9YB6j
7B8qTCSHWrm+Br5X5KwLSVuea1mkPlnDtzFNq2ZfeqCLUaFo/oDxNMlkluL70zm6TGI6/WQ7CXSB
LR4Idgc6s3kw2qQ1z6d7AipZ3nudKR6zkEXQkN2NZItmlqq6j/e0joeMMXZ5oUkxDOtxhSMawMUr
FGi9tGCBpM4aYuqGybzbYI5VIZT8M9yxLEsioBB6guJpUjt6Vl4mzLgHR2tiXX2BjG2BEGDs92U7
B58mHcLkUI/wymu6hRUPushRkwChMMv9Jbog9xsT5g4wc6uYhFK5NLcMWb0q26Nz6G4gmnbcOIwk
lwkcS7zy3JdRHNxsgzRzuFQcb+sq5FjSPcAP+gzHD+TYeylJdzCiUBXc3jDArYFrUp3ZW3YvtUDo
HqyPFXYDFmgdil2SINIG3c7uq6z6Di0FNXj+Q83RGP6lBC4qrn/3d0oWMPAOcsjmK46ZacwRO6e8
ve/Kf7Dyn8orPsB9V+Q+G13f69E2ttASksUG0W/gkjG2p3dl9C4zqW7bC08ix6gIKgNdz9VtNzg1
a1G7rT/+1VgPTN9mp+1YhHJA5PofhuFA5yyIgPPwVgkJ+l93obGXavZ69m5rI1AZthXKrJq7x/7X
bF0wS5PTcPoZvg0et58NDU0+INeeyOTsyv/CYokjx/+6x36WjaboEwGPUu+SJjIVGiAK/yOeFK/4
CZzR/IVaZGANly1gzqhV6zQ+r6W9HEGFpR7EMEGpNjE71uNjpZVQeyz1+7BFSxq3exRowSq8S/9H
MUEvcJ0P6EJxrC8qD7EzLq/JIOexpGCSXcq0Sd5Y26glfv+LkjiKx4a31eMbiOr8aZh8/AqF3rtg
74E51qiRE2WSUEee/t9gl5sr8TqZfVHlqvNnkLeUm7y+sznP31CWGyChqIz0j/knJ4eN79puEJWy
KsiKEJgDOyrz23Zljc42Td6iZ51PQwHhtD/2Q4LbQ+rH8VFqrE2UIl6527aIYmGZX3fjg7nJKhs9
7CPMPvrVOWTIKzElIvXVAdhBPM7spXN2OUSgitFbHKFL28BESaK0mtuRGbtqVtTXeYl6E61fi9eQ
E81hyYKKzLcZdCLMP68k0eUMoTGCLFWOOlH4GxxNZDRdB2mwHUBN998HJMAprszIvZc8/2FXM2Ck
ykbBMskeaR5Mt2mR9Dpm2qrGs+HH3LzpPAgGg0EYEQhrSOrokBpmgrX7oyrKVXLvouomvAoKRuFo
DyMuqW9BvYlw507nqeY4IRMbz6LLVfDMbRrh3a5X4Js8dzMcnojqj4zi0NXfOgZRpStjMk9FGB1b
k39TOtty3YCkAqIXJjfLF8wNQaOtFVXP7VVFy+vZqAONXGE2H8ACHaWSYJ2gcr4KqhJvXtE8zNpt
TTK8b4Y117uRk8vuOfnlUWqI4QV/bMy/L0nXgWpCT5cMC7YQtijwIimydneMwmm8TubLh7sspJlv
ia5r56bgcmg5QwdZaX3xJ5ceHYTpWXgJLqCGQm9LTxSAQDPwUTPXsdZPWM6mpcjtowL10ZBOmmQR
KCyHPAxZo0sTjqLr5bFgVKvd4X1IzHpCOnR7Gq1fWLdgmgm6Cw/DsphvK1TrQ/JCFNvculN6REdf
kDWKD2mX/lnjNdMNCQuEvx7KzE0HHJEd5WArUTj0yKLlf7hqC6qqWsdKhOBFmw2VyNYWVNO+cy0Q
PwIkenOomeg9JccnNhvLuUFg7BC9JayeLF4QkxwRlhm6FgnafUEXKNbv9Ndl2/4S4Qvpgj3OuzZc
+3MkjWGaL2viREGsqhs7MIf/IB83JNvkBeFOK08JDbMVj5NFk/UDgEZH5PXaGM5PG2pVH5Evu2cW
t3uPbAx1gCmkSoD4qxwDn90dk8tvKnf30wQhxWJ/zbtH01a/izPh7DD+gJQ/E+8UROii06g0zL84
wzQWi2kCWBEjxufVVpLGD4tqfPb5YI2LRpUjCdoEvJkMbmYo1BlSq4Y5DEzHV2LLclv2Ha8jYzhP
onMgj+jZHZ+i3F2jFmAE3HPf8Xd3KBmZsMcXlgrlH2cMigpY1AfRqCJXf/THMHqn4XPISCIv9r9Q
3KerVnS+Vf82rArTMphJqAh/a7KhEUU6KwjuL82p3Kj49LVnQHlAcVvpGuWUP9a/bmGwpZtSqohV
0WBHcOMrFL0hwbh28DHQNtw7V3Nf4Y5IKw6PH/W+PUIsdOssnXu/s62FXHgVnjsZfo6xvNlDjVrR
MyEdilyxOOkW6tHRslRCWBFE3Rx0BOB2ftUxd32Pgqq561dybvAwIWaN4jYLpoZ4cjT31v7p30Pi
WDcXsVIKhXtpxb1jFKLU1kjQYU6L9g15Gr75W9kTqDCK3P9/cQjZ52pGoGvsxKOGhyjgtjl9cqJX
SJ98JNlhJhu4XDNA9tuTnJ0CgjAdmjhsGZsjjEOS5SKfDMYWQ41IAkaJSGRtC1eeSgIViP/2V8B+
/0mpNLw0ubaxlRP401T5j+Y6I2F75MVF8pTOxS0jZRb4Yjh9PbsvjdomWNBDNxVJgJ4IPSUymiY3
D0SO7CkiZJbPI8zI4SYPxyTOEo4eZwTgCAYg7nA3+jd6cS7qE+v3X8jNUkJpUaQLndzoSU1IYXWj
4M+QBwUpHXL3WmsxHTIB/xAkRrhncjyXmR8btQR7Pz8ifnm6NVjmEr7VsEtHumBZsZY+c68n65WW
xQHhVssIplwL+Kb8qM54u5EoPeFCR5oOAZx92y+Ah5Nhv2wF6/t6H6mQEyHRP3Mm2GOEARWtXsh4
hOEDl8Rz93VQB3n7M6HkeBgj8ypGNynOwGBU4WVGXWfWy3Qp9eigfMVQe1Smmq0XR/WEaKlpokr9
kTtblg4ipvHi0x2VAGGVTiYQMYg8bPwxYNdvwzd2gbIvIb6y5CZMDbCDg5Y8AdjNy9wY7y5sv0S1
I484E4CySCXGFZk1AeZzAxvlvMGnV3u0JCm2lv/VbXMHrYbd7DlbaUaWti5pxFcC99lJFQBeT8C3
7Urc57a+nO8O5a0adWm6+Kk+KhcLWOU4k2vSIXI4k99BYki1gjutP5yEjbhQ9wB31MWYK6gC1EM3
zjinHUSuEEYFGL6bvgRu+OIBEV2MQVezgop2+4THrY7i8Df/vyH39YO1r6xHOqXktK9gYbDs8QBX
YkxSyOziQId8VenTLvKWhAr1TEzDjRRucgxoYq4tKmhyPgn5jqLUwxnb9flxK9cRzf1nk5h75p2K
L7KraTTXIHJjj3iEoTuJ0y/0d+sYEMK1GFVUeBDDZN7+z+eFY6YWSoxHg1jmxYUOJ0M2PLNvOn+m
OvBvXdLzWgHFv1HadLAgZRncnAo6rzOMk1fYH+w2YtEtjLKlKXqTdxWl1g6N+E+DtON0n/jP9Xnu
LSmkV50qe8LxNCtRKaC52wZqBuNIVP9WaH5LLeup7ROvxM042AnmLIXWwjqpSkW9RpQLoSZB65R3
0CcsGsQapDiCk5jMcTZe2rP8lP9hYg+tEsM+g/Xl3cPwrWR8Bae/brRchW/peIkOJtg414Yz66OU
bzYvRrK3wLB/YcJQGeK+sjDHnKpFgG0e+WEPnI2MPwmHMwoEMLd6vffORnA7AbMyw7sab9hkTFWs
iYvCBpjFX1N2neo+tb7yEjHhwvQKp4BxFeO7FWJfFLBgHXiEsd3JsoDGigI8jtJpS1fk5U8wI8s+
RpSDE44leLrLi4iq9b2TIP79RAVVKG+lg9A6Qw69xjYVFF1jml4oPtIqnB213HXbMZnf6fUbQeCk
2PXfED3D1zPWDc8HrPGL9eaVOOO997o6vCtu2CgJKkIr3sy8auwfqNgnpDiL9gkN8F3n6WYO+jgF
2TROwxJz8CWvxIBnx/bCqGmVcvxIRDn+C+7Kzutz7v9817uGUuB3YDWOMVQMlX5waTGN13i+jGIm
gElrF2+fzmGPxoajVaC+hQ9bSPJhhT/Ou98Y81HJBzaqC8b/HytUNN2J9ddydK9s1T9+YXB1lGbO
cZ0LAznO4Y42zDiEMjth3g2t1oyukjWjgX/6HpER+9D8591sAPSdWweyebRprPfLz3KVh5Lyo4GO
ZLGZfiZ6ln53aHQWE8ZwjFOafyAzAJ/f2kOvmVIqmGyvEC5A2gyrIRxCrfeOzGi1WrLyvPPqOC3d
dPE/YJ+WGH5KgBC5a8chAgMWUe908mYMKtpMbD8XfASoc1IAXFllCxT6VaOzXMBVD1hPFycBgCyx
w+UoMMqJsUqBT/f3uKGMeEJKVQBbboLSZ7Qz3mdj0iTYmvwBb0gdAdxcQ397yqbpFcaob08divHJ
7fxuVA/2681Cus4usKybjMtevfRSF7W1PzLcKAbYG2YKVHOLDETz65u3nwgkIziVU8Hywfd4uFn6
70nl3lOwzfIdxafhl9sx/mmtLdpe10CX12DeE5A9tG6+lP96eFa+nufXgqJvqlWU8MCz7QGTj/Q5
00YOtb0gStwkSHh087ILAda+upo3QcjJcMbkPE2GVGrPr3ldva25fkDrYJzsGlJvf/yeZupkuk05
PAU5hgpXUdN4nkHJfJU4YiH4SPKXSFn3xK/tcuDi4Gr4VjtvQ61l8+A/PSBVdB5skWTbM0WxvfEE
B40L+gLJgxxguN4ZI8WAciP8cCRwh74pJ+VXCJy4Jh7VQ77eBwcqVW6h4h5Jb/ZJD6dmps0qAE4e
uuBR/Ak2VyGMSC0JQu7eE47sBbXnvmKdPvGwutlrqPXte6m8yzMoKm5ob3mD30xFQRZVD8W1fYW8
D71PrPKcdCjOdO57/lvCqX31DN4IVtf56o+f00lDBFIkb/AQB50yQHOANi1pGAj3aZjiBk5y1R76
YVU517CqeVNRV/Z4BOabwecDENHFvq1yE5LOeMIgIgCqKlHWBHToNsiVWpDmVyIVZGS5Quez/BzF
9dkyU293NHPgOFI1r6+hjS0ZYSClHsgbbb7qIFDaA2n/7SW7NFhWXvTloSjCU5pt7XT7fUcapx3n
7hZEETqr6Atxs+Aad4dPZAy0JgBCPFaqsJ+qJqazS34o9qjqJIJtnxo05KreIf+32Bud+ZtNgwO9
KM5my93tzajw5kj944p0EoUrDjYZnFjYzcESidSstRg57blpUupS1+RTcg7EFMDh2/wnXZaRCkYw
R//vLGDBXfF0RkL8WaBi9PBaSI/H+AQwWNyv6pKULRMng0Fvqtp1lynFfAJYheZweC7GoQVrHv2Y
uFbmhauoLPDsu8yf1iLdyXPJ5Alz2joe5EkJ02GWLMbvzze+swNxaV1bqDtGtgqIqnnet6d5kchT
AVQzPtdIVIAz7Tn1v+IdHdT2+NHkqbcWyPhV4IExtVC+sc++1F9y6hlbZQOJu9SJcV5ASa+haU9j
zFoSGRSm9eoO+DRzH3XLBnnR4ubxjQQIQloKAP8qoNFEuK3IA6t4K0YJI2fn8mL1mQZ6gbef+0cL
yZSPfxfbsTk2Ek8TIKrhb2Ey8yIf7M77/Jul63vwghuMv7SMvG+Usj6nXLOzMx1M9xx/xC0v5AJg
pXKCWoJaFSF5IvaLXOo/ftnJ3RNG4KmEc2blk9/llfQ8d3BppTfV8w7/Bd4H3+WVQ7JTIZON9oli
cF+JspagAqFfNUIWH2pFCJ7sVPHLBJh3iBg5zk1xExme2NhxNPiKkFEBX1wd4lGOAUKWFrk3/Z2d
qdimGenhpZ1mjaBXK5N+82Xnvodan/BpC9d+9Jgxb/qh0GexxQKgRJmPfuh/RuGq0r3v7dQIBvGM
1DbTGR/irbGLQZS+glm8fU770V94yKqkXIcQmwWwg6x5lVcjjB8K+zYV4MYX3BeD34cE1Lmm/Air
nupq7DTgPUOjtX1WM9dLiT2YS8KxgjC00sizlMqVgKsOOAGfIUjZgXIHG9Se2PxuOfn+NzFVn7aP
9oroIDVPcuM+NXuS51yfAh+CUH4pXgXMwrPihYeCvKzJZJ61T0jHzs7BwGc8fuzmpR1rK7OkP4Gq
vfrNDO97fwzjj28m4nV8LRo8hhcEGoh9wo5b+6d2JzRaSakOSvkE52/jX5CYlc3BSdtz0PdY+c3r
CHyjNgqzqNwO1519IZvKMwptYz5vYwcxX7JjpdkvDnS+YAlyb9/Q0RYAZ3TKfOrZOlOK0+pPg1Gn
6l0oiyuOHs/qONqXtmc+Yb3N+F0xtqL+xdkrJDVG0w24ipP3WnnBqNo2osVZIyuVv/9T6FMWtWCT
I8UQAVExX5jCrHTnoy8y7Zd4f9OKSZ97MDQiX959bfcfhhq+Ya1p3C5udWAlteTuxzAafH5/zRXY
saHXn2nlcr9X03B/MKtcrTJ+/rtljpWid2T6N0voYjUA/ILOOh38Or6IalKf3gipOAB1RBNiH5RQ
d/zhRg7uKfP4Ie9iDq6twyL64M9I18rwevvirUpeUggSbT033ZnHLvWNGchO9qEbpfveFQPMCTbt
CcvVXT9aNtVb542sa3vcsCHZ5E9Amt44n07KJtd4G8Pho0ZBlQ9R0n+V8ZrIDR2WW7XazfrC7vE9
R4qsjex4P36VcqRv727irAxI0pBqoUpeGKgmBE2xjAMyV6CDS5J1bE6MhCI5lUFslTEI5OulYkqq
dHb/iA7T4FDifSpok2YRWpu59bTraSmlfCUEVFtcfuEKdtoOMEe9Zo5NuT7LxlRJzt858kfXkzJ6
2qyrBtVjwYnITuik4aFY5XO+yvRTgOt/JdRYNXgRX7J23nSIosm9lD8DEgqXDz54OkWyEI4IkTD+
Oaqnchdg+jngTbzplwVL0/yYL4qskKSp2GN9tmMSgsYoKtSPEEYqv/9j9AgMCoK9QWCTCnwj9zBa
Tm7v8UhiGQmOQWbYVCOY+pAzPuAo8JPY5TKQPVf4TSpi4tXC2mVmEUNsQQFLuFhFBZn4VwRmET9B
PDVOCbswowtqMqOhxRramCdqrA6ywF4Kiw0IWyVtV2+axVmKl+bBh8D6JdT4WS8S5bQurmud6YPY
6pivugpAalj55uBxO1XvXQib/UudQvQ/f5/fZzPpByYE3QTiimnP0e54rYkzjS/BAmYNKSJX0QN8
p7zgsMaCoiCeFudC3fSYl5ZhEFx8HUvnN6P9QaMLDU7mOcCo9qRyK3ZYok/n4jURFOXfqJYxb0/t
ykNQnv1W0SdsuEkDf9d9sRtx9eO1apvTpMF3aKF1Q9Dvo9ttc6qHkHTJRKI05cjqHo++9nlQWT2d
kNTNJuxVVGAQZaU3XKCMRGYA/wWV65iQbDLPuZTAGlyVX589MJDRc6zDtVuRuKQQROkzIP2ygKS7
NPjsAqg6wRJh01NqetquShrPKhM/1nUY+LjYWYoWCSN/ero/eKeN7pwUy6A3FUd1XqAYdSZcajX4
LE8qJdStTd/0WW3UmqA1lGYihybX7Owrge/rF8UVUcarRwS6b84jvcuxW9vvUp53oRnzRkOJgFk/
LzwU8ohukOHKfc6W4ONeAXu9piUP/q0dz02S1Uz85kDDNrlkA0ggrkBrHpFJDkrS3lW3ZQ80uGLK
gV7Rqif0mH/xVOW7D9ipo/C1W9Jbq+t95Kv61f7nED0e2s7H7mFRx2E5aoVI6O64bUr5ZRPBRmlI
Wk5qs80ZGo3Kwqr9Q2lIhdbrKK5QyOdmUw0hEZYw++aH+dk0LjQt7uFiQnWsF1yzmx0mEN2tii0J
235GaYYomYpTZPWQNdX3cr4bndR74qYqHTv2/HYZ55PsQ04PIXauQOQzdOOYDMKB+Ois7lbbhxYH
O9DtxZDW5VY1XkaZinfc17QvAZ37Wok3k1moiX4/Mibe/fUMBfkrnG7zcQWewIXgGI5+kFrMtjMN
sabbEeUIrfa4rj5V+uIPVbKBBjv1v5DT7G2mkbdAPuGCMixwSDPw/MFLfFpqLfN/rK8/O+EPbLkv
mJTn7ZsIXDkXVhClz52UpExZ1dXekjIT6I1m1IXHex1ltoF6ye/c2gX7q1sC6RqgOZhu4B/PSJdh
S4voHa11vlG+WETRwH4WnWaeX2NdRzjA60KtKI2fq3qkq6IWEK/RserGz8E2KgtEyZkZ7Wc0HiRc
3mxIcNHz2hRN17DlENOD5b/T67TVMQwKe8NVXCGuwzrz0xRi6KLe+3nnzNoGSl3XBApI9/w/ruCQ
AWcQBYq2Rn9YtCeTd1/1SV5J97orxXJf/MNK999Em2i8ZU/4hdbOr2NuSnj2ghByDHRQ0g1W5goP
7OX2nWpgg8nodsH4qDVaaxY1FfgTktMWYn501pg0ikGE1ueceQ+64qKZRHFE9InLjpnxdNrzZmTK
yQmUOzFjtJ1xjombT3gK8X6wa9Ycn0W4qe9vcyuyErgFo6NgQdwipMc3V3DGSE0agLZgTqhPtLEa
9HwtwUYGYEZrro6XGUcGTvzj7WMKVneS3QLLjhNY2gPZy3etuF1zWHOU+m8jZRmCF/eYqsPC/qs1
SR6bTnNOHcf0BGPRoC33psdeVv/7X/oTFsDlE2msjYxHsDbW2E98Mxlc5wt5LYsGh12KNtiy0o78
dvhpcKS6Gh9FAShLrKlclwDZURik9lWUhHpmChWQNBHmiS/jhl4QxELJ5nKPVCeK4fQ7NWAuPXLr
hHGz5qTBCXa7fGA+AQZzmidXSwR84tZknWEpKR7CMQe4uwjxpDsSu879/YSdqZpW3tSEmQFhexrF
rjvuqzpilvelNsWT+uEf4XmezbqIr2Fco9wo/B1eEJkWKdPRRgcI7Ivzxc2NDygnvcCI52fj0eWM
2PpSbY/3x3Y6IehtBJz4dUA238xK7BFVNZJvYbXRK4JlE33+qP038OnMA9tYA+m2FtLHJ+Lp4QZC
z7irY3nN9Du1aft+q4UuXBuVu6qzoeVtawm/vGgUvPZnA0rn249/ZTc5Oq9AApZv6f8Xew8EUrD+
BpA2vXwWVitXuo4/IvhelhBFSNObkJCjXeDD2FwmmAZQUHGwzgPO2sKvYhqWkMruDGNqytqofKLQ
H9VlycIy+5VIM/A+Np+JkFmES/YDUqg5dIqJ2t8Kon8lSbxAq/pyNMBQsAuTNeRPR+u3pEGTj9uU
0CuEFeajkLayUbfJh8IkJ9pelIGVCRYbkanzgGR8YiZNako2//FETszbqo8o7D7uX6R68LzgO4UU
O3tCmFJw5K9YxZ2aArTDDAzBG21qsfQJSHhyheKU3iSFbcZLIJu4j4FnGQ8HbQGcpqpDTQ4/HCIj
+naCmhmF45hpK5n7CILQENwd6Pe8uIMntJ0j1qTrpEQr4FtI4o/2ghLFkdRe1QKVtq257w0gb8xO
ggqqbX8l+3HYavKTjEu0PIZMzYRPo8knknJnPdyehNO4UwXDchtPAuI34tung7ob9QjJeKhLJ4Mf
8qigztR/0xuKkb4CFUpkYqsDSuAcsGmTzcNQ7UMOqAlwUBJv1h/1L9Wy79acgXotmW3fBSZKbka8
3qOCUmk17lmP3282O/YD13swwK0m07/fs/cH4SE+fj22Prvd7PQME3bMTiHa6Ecp+3YIyMtf+mnW
u5J8KhsTF8gxEox63OwFtti9zubXSr6RmeH8FQOLI7OeD04TgYCzK8KrJgP/XyjkL73qRA2qMXVg
q7Sv6dj0ZpMEJSUKnFQWkDCqTrx1ofoCp1ptzC5wCMpG8Jc3A1vEBy+7ZwEQIIS2qGRNTubkAy1E
ahuD8LF/odoiupruXbFlo6TWDbuRod4phnNqK14NU0oTTs4aDBrQ/I8VIuu/qanknl4FriBv2I/H
DCJ0gq0vpowOR0KJHTw6k1SWVjHRO08i3nI925ealoIBPW05vhV3kgBd6nEtjSPElTOJeBV+xk2L
14o9COpm5d2YN5XsS7MMfzPXXTw0Ksdw9xvrWDNzk90NZeVr6w4dCjx8BoL/OeoGXeL3ZZrfJ6Om
TTG4y4m0hYVoUhdn5iVDMQDyUqDzWNr0ihP5ASqDi4a7VpBTV4rB6KqIuGf2TZPBkPBDRRYMWOKg
tN/v8QmQOWT5EvOq5CLTvyhl+AVRMoVERvUY4hDANJg6OvXyvMlVL3gv8JUOQkGqBIvzewteQi2B
pPujx7h6BHudqrp7SZ/b75TJQdi6NWdUvqnI4ypOzCv+WB9yhXqklbhjH8fRuFyINXivL9gQi6jV
D2ucIwhlsYEb61RENbAp3q0wNrCInoHAJbW1spzpLhomhqv58As7yWOrhJaqLC5eSSq4WMllzjne
rbB23/BE0u4VLJzay13wmKKNdET3nOhA4Uz0ZBmgrnZZlsU6PWW176HaxDxfrueMjjVaH3GnNbcH
3bCK+/LmfKkwq9n0R2Fip1eqqmhIKEoSurwzDZBXCgogbkaQnu8jLEOMROipnAuMdOhsgNxXpe2s
n0Bn1nrCgWejmzmqdgpK5b7GZjRUMFi30qRiFDAL05G213OMfVf5fiyLe7lDKYN4Ke4m/8nQ0eKK
t8MKWU2JX/SYXpJqMllEotYkeewMM2y5YDAl7JscdVVMX4+N6sFyiH7+LVFOzO4jDyDKwZInc9QK
m6H52htyXfA5ZsmKaOFWDd8mU2HVrKw1UA6dvon5hJGHYkWzu7o16A3wl513jtw9+9sNP+wTdCoX
y+yiuzux33GwhcwuYvdOmQ+UHubj5E52u2N8o51wcyO6JD4VedojNd/ftbx3W7qh+KuaeEILCThq
5tyjF2EVW9Xgq8widB6xb+oXYQprO8IAPqN+v5k49Tvp7QlF58FRDW3WX/i2MCkRaL8Hhod8Z/la
Aano7TJjIvDNGuSIo5ignILjdvcBSEjiJ5IG573Ro4kHD3aeqDHgcc8YsQyVUPxY1ar7mf92goZi
cGOHxftbmyJZd7TWWgtTBiA96Mi/pOTRwQ/unf3lw3MF9Mp63fF8t0ZhAximay39OOYUrjSV7dSR
LLITLUrzpKiQj9kV/BAWTfsN08WXsgdrEARkzKgEzaqWg8890A5rvyxOscaC0IRg+KyKSAALJuXW
GR7jZIkeP2XtKiL5ReLb9oLn3uZ9SDuPhmFUUhnqrvPiLfqKn/eoVugiQ+Fj7Bu+a03TZ3ZXCrDM
Cr+HGFDF3MGRxqqqjhkFnEEPHB+K/ijD8iL8oZCTNzlqK3VNBWvvMQj5x8r54FxGjRDurBSq6RQi
dQAQ6LA6np2ifZmAENdYU4swZ0/w4yk8fZNrF636oJwKOetZxJAwzuhBxLUOPupuiEX+wIf7Y4h+
QbwMr6YTCnXF0aN2n68Q662AWX5BUE5Wi9n/5WaHgzPyrP/yP9TuvQsYv2JLv3C8WANLrhdKvMym
YLEjDtkw9CGHkPscZ11aLe7eVxgNL8X6F9Z/9TQOp05stGKiBEBP/Z9ih21EM1gc8amfzTAebZgk
CPNFP4boPwvo5DZ/221vyVQ4LMmoHPbGAMkVHG/S9EpcYnxMn1fnzQEgk1K+PyU+WCCk3qLRfRi0
HVgpsGlEvHkiQsyR/rZz1Qgk5j2U17BlFiBnmgyBOv47/q9DkCWp61mKTPeWRFdoeNELixNR69z+
8XQ+1OfpehxAzAgn5ERqCGPPsz0xbfsL0HgHR+hJqzAG10Z+iwrNfwMKZ/+nGaFbUENDmtHRJHTJ
UzhlNS5P81x1iT4L9z32m9unZVxqjWeq836tuk7gOROmrL4JFQHcd4tZNqjPItt4wbSGMRsvCLh8
DymF3TADwavWWPFx/GvEkUutMnL0r+lmdmCdPbP3YLapSsFACdE4IDOUSnF8vqeXWHqZbz2x4/fe
BXHWBZIAvjTX3Dszv2z548DU5j/aaAepXNCwuG+sCQROZg9k0qKM6AYvJHE2tKBBCiGf1d6HP1gK
By1B4kpfYRYzRTYZ2GpHhgblvKyhZSr/MV+UA4JdtWsFQVRJhbE903lgspCIptgoKPoNo9ApvqjZ
Qx8vUxqH4dsSmxTP67/jX5QZRU0nlmFGpHMYFEQsL5L/xM1+R9aE6EOizVEpSh+CElWYFmiRuKYp
31oLdnV4RrFrstoJexCUtHttdAaJsqxU1sOJ283Fv0k6NfL1RktS4bNiGX7PY15X+ydgXnXzXo2Q
3oCIYewTFos8xYuX8Y3MFAlUTgNhsVwtJx87512xMlq9Dj451KeljyWnC84VtE9iPbYnTa7ibimE
PRWhD1UHQp4SoUd0yCHxXgvIV4H4wGwub1wYJZZM9BDMTy5iYm17+Zmnkq0/ehmXTNzoYfvLCL9N
W9NBiTgE1rsBO57bF/hopjIphGU2qRou7q1yMsd93jOx+zgO/nNLdwFrsWxczghbXiFiiZNVqVQC
xTE1VoHIIg7xqo7naFe8berg3S9+P3z/ga2FDVmduXTdZj9j3pHSsXr3nVeVE9yE1GapyxpCdKcY
6vrnUKpaJrDeLYXb6IIw4QZxacehXwQ+MDIyGq6n6s0cU/71yfzH3khoSsTsLTvVfk33QkLNcFNE
jXljfbxIWA3wZVqw9BVzsBYOAcmypvL2a8IL5bRC6xOe+dNQ5kNulk2YGmmqXKkB1e5e6XkToAgv
5jzrq37x7iEWopBuvbpG0hv0zhICNT16XbamX10EjhPeHIPG+0I6Wc4LCcAd1UfbTh8Qe0VMEhAK
5iUBmnDmswi7JFTsQC8WqR3ZZvbsurrkSGozypcw/5Km1VAnPm+EEIJsFfXFndE6Y1ShsdDLWftX
IGZHpS8dAOHQv0pBBupAXuUv7wN7H8TCaALKaBigTnRBViKihRLe7mV5bQZoWe3cBZWT+Zq8CGfK
9eQYUkiH45hJgdX9Tmy2kaUHBw8wutxHKNCK++lC9n7410psbSq6Lgt1fxzQFmG7ZWqzvib6EQpI
+dWhL/EH8DA73LDs92/hUUdfshO+ajAjaO5DU9CbcT05Z3LvAxEgWneeKcUuCgZxnbLeUuqTBulX
LZ3hd+sQ7ZNlxzhnv27qBnjiBiW3nZi606wN9ZCjNsWcri/+QZhBhNjlcG2N64L7UDvWngcTh4ws
eIFsp0ki6mX/wYD4EcC8Og73/hBDNkSlLRXzw4pU/C2X3/bx+w+KwnIfIFmHKp+inIH98XMHDSTd
KwKg9MxZN4FF3IU3U0yYG6RZWTfoSw2WM++T3pgTpOKrl6VDT3PGu8neboNKKiNCnUWzf3bachGt
BABa6XwcSwLO2T+u9lDHW9d1NWLoItHrWXFm6orvpthBeGyONiX18lgzNqCidGMoXVxugkw+ur0g
Ta1Fa16JSFqiWWTt+/rA5MNIElbbDBKLK4xHiWg78L/TmFYSAm951+VMAnuEH7utihjtCuXO3K33
s6SGqirU2MsZ6D8NtPBUBIw1L4J1wBmRinsM0QsyqDBFexjmoLdLSF1f99mKIiABFD7o7EFuaDnJ
H8PsiwOnhUc8wGab5P9JxGbo/OtrZEiId0eQyytOkFtTdaRx9q9NyqCLMNdP8HrpmagQrqetUN81
kSobJnx8dh+cDyyfB2Jb1VOLitJX80Dpirl5/0hbqeZMinLiPjVwRYgHiJ7O6UOizE6SPxUnUivT
KfF3UDUCfNDQesFGbjmJ6vcB2FEUN8ESb4xZ79fQ+aBM0HPwfv0KPexm2+8hw0Nv4tcsoh65lKEj
VoL7NHY0aW0YGOipgBGddN8uqxXvX89bSL0K1E/HR5Q7albqPl5+Y9tFLtdibeiLMamIwICKeHpW
OvWTu2hbSVYhEPWWe8thI9QiLVMyU0x+UDJiyowQh5miF8a8MIL4SPh6+43SDEwe6noG0sFIieuh
1yzRV9CCngq7hpAPu4aglo1HpGPqeWqm7sVUgcZpKGRhCOXjTrRBSIV+H8BAEoc2GtzijI1rKXVz
Haw3NQyYFSOH9FWWrSBiCMuC0r6J6lbE6V7JgtEZFU7Q6ysnCY7AMcBYdh9HqHiH+n9XZCYPf2IF
b27jAzDeKpFjXIJ06RcHre9xHu8XdGo+T/Q+r496ko+YsUjJM/TzX5e1dcHlvYTotUToQlpqoHDD
kao3QYCRmpT5AwFJh+dfz/b1avN/Wd4ZlG+DHu7NsMZwKdEqqxdFHMYxRBpeeWXXBp8CrcTi5tXS
LEO7YsJEQ6P/fPlBg70Lpwv6w2DwdIKLUa01/O/jvs/3gsJ5gKUvGIEd5wytmOxLnHlwQkYyM4da
UxqLMHnfMVH5QBJm6pKV4dZvL95if/HYhOE7LHPPaIiFPUZ7SLeC3/VRmQDIVAJCxGq200xCGg9L
nPKY6YT1Yil/Nz3mRkva6AwbqzW82mK82Wfzjc11JNraypeDWlu11/+iwmD3MZn1edG0JrWLCdOJ
fxOWBBHtNuxSCKk381JZKkz2CJXQvqjnHDs4h+vStKvR37vgMnHOlV4Lng5BrAFAsGrw6/8+TBsL
8nrDHxjN5UEEgzjAnVJ4Dq5N7MlO4W976wehY1BLoCc7pyoZnm+Z+UKthOwToXAKM5YouhPwC1ry
N7wMcembqgwGcn3+GuKeOSb9/CwUbixrhYwQktzLX3co9foAYM4MUJXx9ssP2o71KCQYiPbi3EMj
NFCRakrPYuusPC2LtExc3Uj+0vUmHHufqxtjwA08qK31h5WQJoAcW5YaQ11/lHVhAanTS+8HI7cL
atSmul98lg/s+33Yuf4WdOg+mXDnF8hCjXcPLj0GiVHvgKe94gfkWtVb7/NZ9Nky07uSBk5j4zqw
xPC92S7SWGdQuNf406OjGah2AXT4vP08QtFMk16sGWUbH8ViAnw2U3OAh6Pi78i7PCyLIMyKQVTA
cGJ3k5tMpgQMGsvOWoFde4BuYS95eJGH3xliEwZy8+pYz0bTXGT2QG3JOIiouoPvCAD8iUjjMVj8
Xm/wblcY2xq/N0LbRyn1nBywD1TEj2a7WiVRmjMcSi3FeVcLVd6TyPmnFokDr5qKhVU20PS9xiYJ
sCl3xJ6GFAYZ/Nst1g69XiebfXqHcfO6sBTNoWxdxyiLaHYtIleN4iGkMjFd2WACMOo38TgZQLF3
j2wNEzUWILz63BJUWt2W6YdN1adoZ4L14sOB07I4FG2AB+mssrmRyGgoKzJ8bdgPl20fuYgaEsCQ
+G7eaUGJSRI7JY3OZa4JUuuaink46d7Fu0kRVmJqw7gJ+icApxOv8jQDsWrPTZRsDpQtNsH+SEz3
j+QDvXIQKF2DqzI08Ce53+ZBt90vIWst+VShMzzwyyY9mTz+yYs8faAzoYTtEaGQy+n0FmuWy9Xl
hhalLrYCp+OAbdVnr/WLUPVb9O13hz1nr94yuwar1o2tdl0SlfHXUUsUM4p3mBzeTyy+GYx+2rM1
HeNtkevvwTtXd1L7bm+MD3Yd8SYv5oDsGDjY6v4ErT/kg7rfoLn3SXNW9jbso4EAy0IDJboWCICi
CVOJa1xJxvHs0acseMaj4zD34bgAue9QyMKkGgG9JQYxK5CXmryRYcLcUQjRsednaV01PcjfBxcn
HH4sIzYA80HV6pIKZbqV6SPwJIlypId4KKzXQyfgXpqVYMsolmYGYnsKg08tZpPQmwZijUHanvG7
6L/TXk5VPpPrTnI0u9XGPDHQaYHyvQ7Fp0n5big/BzfAy3uSU9wb9kyAEEs0PRPzuIBlhf4KNYUm
DP7MC0sroqC2n8OTk+TwMdLgHyP3qtvmpxo9UiXDZBMBHL7YH2bSH4ndyjPN50ybTqS7Se2FBEk/
pw08a426h7GHwPtkKP+z7PUCct+PnqtgxFjvdjaSgjBX/VVMmkQa0YcViqiX14zmdJJeLS9sRiW1
PK1/bz+MfD0/d5hBKUlpQj/WbLJPBgMX+WYf35KcGkktcNY4+YBBNaiYRmzEwevVuRYwwMZI+Upe
0bQm6JWpDB86ja47/cxVSci2KPlY8d/wxCltVuUBGPSboF48BMRk7uLzHp8UGV5TsRbh1gB8L0EF
lETgE8o276stu3UbcIEc/AZ5PePcUoqDuM6sQERg5HXa6ey7av7pY42iZFhz/3FEseAQA/LkW/62
VgMZ4SMP4kpYAgofZ74aY6xmc6MZ4ODl0sjPGzpevFOlPVzaSfelfab+LcAenjE2EG/hz/l0uXDv
F7EW+Lx7xCccBgFRr5rqlfRZZEKdEzR6PI/scRxSK9MeWGY3s6iFsdrP5Se0phpvLNDNyiCvmBUh
7tgGeGx8aB+zAkcCvTMnnXgZVhVaJR7B4YdKqIN7AKMLGAi8xX3vRw3SLY7njrnRDhzrCl6rKhjR
bo08E3I7P6SvMVcdy8pqD9YG0656UVXfX5pHckUP07Lga0KNIeCEY9tXPMxQCoLEAf26gwTPJUtw
RY1Y6EZaOM6d+Suotops6bAXMuXWW+5aBgr+kxqEKhgVG/7LN7j6/QNKDQAlGz2bb+aWcasaQRmm
eXYIba7UG6MXT6MD5M9R/0aoJt8jtObmvEI6CRb2FGJIntFy6BZZzNEFni59+Mja+r4J245magwv
1HgrWh25yqIkjxrVgrhcgTmWin0tdFGvnuJaGGOWSJC97bbYckZjkuzn6btN3/f9Wl4vwkijaG+5
7rOIgMDL5yowLZCeH4ZWm1eH6lA4QMQOlmThRPuZpLI7khW7aQ6/SBgsAhD7xbk0UwfqSGKsKXjH
yRcSKKGkIQKURI+Gx3cIwaIp0k7umBfEbSUy0tahzqI9s8j8Frf9ftIlqqsSyav0MZr6sZZqGQlm
rWmaLtS4J5GPEqAbhcBUzK8LUC9HhAT010ZcvnnCNrQyB2u0/Fuu6tIMbrrtVX0R1ERCpKVpk8+5
P6cgThxTXoFA2LDT8rNztwB0UCes++HII/AkZs7nv/YwFYhqkhIPHZxiN4Yz4XgWwwdOsPOuiLEP
oRBxcumb0LtaDtKxI8E4p6kpFEz8ZGFSRYtJZDdTNDQ5bGG6l4tVezuguDtzcoDYOIT9mVBpVtvW
t3YVbGWXsC3KJAr6oQkp7uO6ew+P4cHlCizqkYHx2EYJXvIcIiuTuCUN4Pa7SB/It6niMo4/i1+Q
FF/eN1lFYCUpVhdbB+F5fv+jjSQ7/e9CBCfhrwbSLUU8pQ9QOLEM0f3lNxANcMVAxPA9Hhe6M/vI
4LB7EdGjaYSRNf92w2MMDhIa6ZK50xjyFpBmS5h8SrJhsDvKl02tNFqOJVattw4YyfIr8Zg0ccXi
1dl9u44/ZdJdxPvnALvK4p9OSm3YqkdSm9rQ7s12AULDM7KCweXGG4TWrCrb5XoN2J5hBQ0HCoVE
A1a+xjzhAtZ6qpCwkC1SxUpUL1el3FQxzFqaSb/3mrrn8qBwabMaD89yGg+5bhKb2FP7Uin6Pfli
xOx6SAp6X0LVzdH7J4+cmDWSvnAyNgNfv5BMFl0D3nV9V2QvVt17hJKmt5gQF0BeZblYSK8BR7Yh
Hl0LincrDX76VGDQcfJfnuxfsutMgficXDHcI427IPscj6HktjaBES+2oyOSRTChZvEZuja7SHhz
GlZSb/9j0+vvpJd4PKeqImOIeNe7epZ4J0pf4xEsaQokp/7l6QuOiIIk7Z+k/8EXN1piqoS7neN3
uVVfm6y3JR85MJtxK64FFJigeT78EWlPA7P3Wu9uUZEaTEdl+ftEocZyr99d0FMkC+/gwx/2kS88
65Vl3x5DgOJlMzorbXJjSg/RyRiHb8btjuPPhAGSk6/a3IYBxxzvxUCCbNlfbiTdJVj49QqUBqOZ
0TjHoY2rsi3y0Oz7PQNh9Akd1aznDOxHlZxkZGQ3VTkzTu0itORSP8r5/Umz6IWM1dq/4X5rdJXn
EUOUTR9kGLsMy/EY+2e/7WfHOd8r/gZEABjX7pR6u7NEZSuj1Dl+TNyzyeTGz+Wv7SzrXNu/B9en
MguxKNEbTUiBgWWjZ4uAno3L21scv+5efP7Xz6gaOvVWirUH58UOOROY47eANDS1e4hQMwVomzE5
qqt8lMkxn1D/MWe4KBepOFWtJZeHejFrf/GP+knpBLPmB7f512Ux2gaXDgmL8cUcnhVCzcPfjSgY
yV5MfAW4Cg5QqMrvyVDeyFdOzp8Ly94C4xTwYU52bS9WbxMj1nW+ByuaHJyYw+Tgz2g2wrotMAS/
Hd4qeQhoBevGNnEjI7GsX2ySWTqCblxDgKOtwPN7RWHcWQybuZo9NywqQ8FgUu/IHntD2zsGNoD6
cxOyFrIbtsNnTClB5Ez6whNA6gaPqWK6Bx3+394scj7VJQlQ03Uu+zb4mdCoLtypOPtD5qmqpq7V
s6ecorHfeZ3eIHJDaoG834v30UV5SBiNtWt+7s8PXrDhLlCM7Ox6wPpIRbV++SyvctbLbSi2TqvP
OefgXQc3QABSkh2XDof4GfeO98ukWoQBPoWpQIyXeXVqXwv+91n5DYvPdIWlfuMG7UAYX/AZw8E3
5pLAVX3Uj4R6RaxBi+hP6GBJ7LxahgBtY3J8J2yBoJ5TWiv+OWRlZpuL29MIC4w3JMjHRiw4PV9z
jj2We/CeZudvNBIxk7ILHJL/yYNt8sDB+pQQnzO1v1DrvKe8YdHTvTRlizaX2+ZV4+xb2dp3fmhC
KWuHCR1myXsxtsZO4K+TVJiqviSC4rqL6xmC9TUqJi+jzrA1T/y1s7HXbyB53VNsHBcOkzdoGSZq
UVi9fwIiVNEYwXboxJpLni0sGAcbZFbpBjz4SlRkXK2R+d6V9dBDsX56EnJ9efB5Yfc5jFhxpVz/
12l+iiwSbnFJZIsSafc7vlgWNw2iij7zteeoA8iSjKDGhnEqAvYIFi4uYYDE3eAt0e5UZTPL8fS8
sQJ40BbBeRN3Hb7idnTDpNkxBqxaE/6ACSqY3VXb6X0PAMvN4a71S0AS7l1GC1qkEVX/W4Xxk45r
WftZSUgIl46tV+c2pRO/gSLXsZKpw3nsqBFgIHbKpTnqyqR6s1eGOjtq3ynwAFtsQdQKBplX5E06
zCszCDiHXyWECJnfWjyetSGb1bFIg8CQzpAeAJWr3x1xzbTW9txyCirb8HDT4BslOKMCni6w1sVl
Z8pjM49fNZFrONwYi6d9PtE7CMbIsDEdF0y+qQer9ULR/hryIO7fp0kneu/FlajuUZQbl/3+vpuB
A3VaAP8oH1qLStBye1DX2NtF65I0HgW3zNDwIC7Aj3zNqb4bGA5vfSFINfofxuKG8vrSC3dh4Kvf
K0GjaW27Po1uVA8jwKtlOy30G7pnzOUx1ADAwZ+tEWtY0OWpr4dhJWOfwx93ZFOfeWs+xJwk3CxD
yGx3iIkoFyRoSbCMQ4OBPjuaSjEKvtoKGKykB6L9ATiDX+5fJv55S39EZUNFb26YzxrjEqbMPW8H
g0ntYeduF3w7GBMpw8ffn3rO4h/GjR3iEBw5eB7mmWLZCPRnypQCMwSU53cDpJZ23jEYbPt98XaY
X0ldx5yhvT/fv9wVDTpUbULV3/JTZYsJeUHzJs0/Q6akfhtrtXH6fpgqOL7xvWORwQCcyS70WA4w
MV5EanW2GMWB1sZOLNjw3i20IjahGa4YX1dMnwD8OmNZBkX9jXcLPRdMfR0DArLBBnYpd4B/Svfp
TuxcaB2HXuomiO1mD39L+jIjWwxC8rVz3Gz72ecvuWGzl8qG81woqbUv69BHcsmp2boht7Lzeegx
fyF0qSON/PTbI3VmAaUrzcT1Iz/9W6klnFyfBhSb/LC8w2vM6EJGrbVFF7Piwqyzd9JpTDgDUo/h
K7emKBLTCS/XQowst00vJqRNeS5IR5ovp4GhOf2c7qIs9429qkezifxvnn+2OzqSHuEqY8HlczwB
/scFBlmKRL7Pzy3ryD1jSuDHaPyKdOyFRPtMGoI0SIYHTTKTAty2nWxgKI9Npyrfctust/r1j9/a
iZZ+1qtxVemigT1shZSJNClS3WWORCt/K7FrJw2AqH2AEsqnuL+2Wnr/9vx6EQrRwOlORXlKo8JH
I4AXDoI2osgi0dU8wSHZUpHAzorR0k8hXuW0IoyqoHeQc4aQpqtu/xWIHSJD6QaYprGkbLAgBRWi
3nqfqrCHWr7TFxYJUXtKhb/aPF9vbwPY3ra6iD2Rr5gyOl36SY4JqMg8ISn+vgvXWsBhEy+nHUFS
A+O4QxmiLGAoNg0bG3TFeNgHKnR1eThAJ+vGRf1297E6zCek3INHOOSLUbD6PBPF4wPIQBhQvmvo
7WUIv5CSg4iAWuJriYc0WX7SbdGh4H6twmDxw18xK6fVNHd8rPyVqqVtaBR16uHeJXXfZurQ0VRv
gK/TvyPiumfasjLQP/k/SliweYfZYDjvxcWM9bsLkmAMv9NaB8I5MMF17Bo8bQleniE5JKUKJgqT
d5SZ7bRipSEGszInOBgsetY1J5yBZmbVljxEkmaE/FSuzEUnyXgRygmAcmtMK+1z6hINm5rdVCIW
w75UXEE0pi4EZrd3Utjn+Sn0sGbE4mwkCKlKE3mDw3+lTxjoJJbqVbl3GcLeAMxD3qOOpROGY1T0
KhDZ4a2H/aitaiJkpoiJp0nJhc5gWHqdvu3hDgII2DERfDOynVgv+/DeC/YJNIGD+yTQiV0hiN/Y
UXdzKMTq9e77PuA8j3838D3lhjhHbPfEBkl8UTy4S2w2cA9r2I/T31p9eejL4xbHJhw9Vl+wr+/Q
z9fdx0988lRvqmGBY+utB3hzmdaHJ4jDpvqgGTvlzoK9ZJ+msrgpt8mSWUexmSFJ8dl5AQ5irrtN
fJ7vAnY82YsitVNTf+bp329W6l4yayOJ2hTW3mtoCfLWqahZ7uAnfy4HmQgAL8MzZ92FWXAraPkw
QmUHG+OsC4EJKKPiPMv1GM5GevdOsJ/lQjsn0PM3K+TzTTVS/I96QuJ9St0ePrPwBPS7NcGDfpb5
pqFqKqNXNyH8a0ROFSKMVC6XY+FjEXQtVMW55/LmB+kqZ+5nIIO1er8giN07QlGzoCby5b/oiHiW
hu0h3umIxKlaFjoBblq8lTQMV2MflZQ3/8szairmv8pudclGV+Qpl7jBaHer+ADeoucS9VJDJfR9
S2waWUBtxwGYUHHPm1L4HJk4DCYoAhpt0Q+f4cU1vWX1oXpMuviXrqkknDdFHV2WVuml80rtlbyV
fHRixx+ek3PKxwP5NHrqBfsMejSQVXYccgtPa3Di8zZTvq3/GG9QqPGC0hg2DehHXXkO2IxL30fa
g73MKqOlvGUyXS5ZK4HUlXHxKpQWHxuEIosH5ctLbxPuDJPJk/KycZL7+BFd5sUbcpy9KL7POElj
Kt98XCICt2nLtFHwkBzbhNxI9lKJgCgcagdf1a4SzFRB7EZdaDynXy2iwqxEjWxFhIrKCqvHEmQK
3mPIU4kt/kCUNb+5iIVewwmwkTqVEipJ7MsFgZQWoJyhYPuHnQ1IOCy0l5ctRWi5qBJ9CiTI28Z9
blBjV4f0vzZ7jo8Bzb4qxH1bZ3hYvRonGnCCPlYVzu1QahSrCW78yN1HCWFZQOkHLPsZvMRJjwjb
6c3RdgefYyxrAESmuVVhy2tBHuLcMxPuEZiC0r29uHXuqJKUavlEV6qWC2GjqOyK+5IHHcXkVvq9
Vr5GJyCwoqXjcrQBHJDzPYr9vsitsUkBP4LjcNCCOUrENQ3rxsAj8lzlqPiQAkolgjN093OAeom5
VrDqnqTtJc40tTBOKspR/XWrv4vA0zBHp5lQjIg9yh9N0LDnkkvoccBUy4LgEJ7gEQSfihcZQXWx
Zof/TNFw8u8PUdCssuwekLz189kcgqzKF0dB08ABE1UOonGgXrA8wG2VUCxW6DKVq7et9HogToDi
YFNI8qQk9jtSci3mhVsrShnASDkmLzQumZVuVrSUf+ysNyHWQT5F7Ga0npKaNw1l57qwTlmoL6xz
3G+TW/wEtCx0H0AFS/lIPo0ywsmQ7W1pZD+8m0mY9+niMN93yGWtVSsUSh7gduOOv9EKew6dLAlB
6MijMmaR5pRYH4CIk88nIAp2UVaHHDHWuT8shjygE3YBiZ1I5YBV3MaquPPSYJ8Megn9BCMsoFlB
OcNSi1L27HEflOhzs5U+Ff6fKR5FABl5sJgXNxAAhC9AMNXbvlZvWQbxmc29c73p2VvZDjs8woL7
Qu/8/tA3c8dxA2EeYXkAPYFzRwBmkLaNz/TzSJFoQZCPK0+b5/vtJgVSPEyX5POsK6EPbwoSCYyu
dtBk00glx8yEviUWtOSFhJ4Nmbvj+P681VxpAE0KSig82g5TSc42/zGv/vDZCyov11BfocLVxess
zcdJ6YjCAbxmCRQ6IEiv6yXYZw689rbm0wEBN80K47NcrNicqecFcrRyp6QyMeviZm6uAXNngkFA
f4GZS1WIYcJw/JKkl5sLA6kgNvhBvSf7Ym62AsvJPogCg+LMQK/7h/czeUql22k2LqPrO+wbL/Bx
GxprMGerqTumPGo4mOxiQAg2geyTpLcLsqxipoYZC3jrf/MUCWbYKLB6fjLsJ4LFC+eadGEmfC3X
rznuQGK09+ejVofdx/FVpVvLiLXQIz0EjNFPMNEGRFn/KFygPqxMPQL1rY0O5T3jgS/irlnMgBn+
eo2D6KpRXd/6ARdDWYnTt049zvwBXtj7FtvtF077kPfqB0GW4cLoNcuZ6ZWuOmJMbzgDTP+GAa6L
viKCa8LFdr03YWfKM/7dyDzFsLuedttyo63ecHbbszh0PuX5DleYQEb2xYNmIf7xApUMw/dbVwm1
B9tNiuFmgQuAx53SRqc19uSHCy9N4v5an8mMeNZH/X3B9yx4uTmI2LYdte/NtomKxmtB83vTmemn
Ysfb773IVtprcEuGNUMq+TuZskNAFfbm4S47C9QxnFWdhOpgklSoHV1+ZBzhQzYMEYopH3kIUggy
F3qhcLJGxDGEjXfUZCjvQAruL8WG7IuWF9WfqWKOOYQ1iFeuuIN7P5b6H54peci3ENhPwfoWCGSi
r9eYYVGZBAPRHtAnbdx0Xe9b+0fPgRI+RkSaznw9s1aoFBCimQTEjgi3NpPcy13nJ0iHEvKr5Us1
fpj94aKLOBSwHaGnlqRm2zKS/YkhrU+jGp0pJPPBD/UBeaMUvc84aX5tqvQknyz1VKU0vl4PiNUl
O4H/kBvdxfPGSKzJ0reBmFyUCC3i/m561e/9mWN0d1P/3jgIzuybQRC1gVAqr5tOg5mbCKj5ch7T
khOfXj+BxGdAgI+h+R9taq4Ia8g9sXEFbEjEnoKRjhDZWEoRLpXhj6Ie38IP1M04pSGK3lqzlvxC
E65xkGXQZ7hjiAkdahDXv89T8hBTTnnHD/+3yTkplL7qKE1pB86FkHWr5Dx9NKDgxvLzkNzww88H
4aixluCWg7BnWH6vGsiG2puho5TTApSceFI+Kb3QTB1zgcgz11A1kBjWU3rpvKfK/uNtcDqSzLGE
OiPOYetCvWZIFw+D48JHzGrfUbcdSIVefr3FwNlcGYhOBZP0vGU8vnh4xvSZ4/i+J5U9vzD3+TdX
WMrDxp+W7durzbda98hEb8Nl1vAvLDB6axSgrnqnOAOmTXwahGGRmvOrL5I4PTwVlZ5sxQWqgwBN
eomhMuc/rufLEkckbwXlj+52BSIUVR7jeJhXDWk2BWjC0C99sZxEeIyOBeLRK74oahtGzxP0OFF8
JQssctOg4VjPTq9qB+Wkf4ToLz1sdaK38AlqhzWWk9ka5toOIeISyUkJvHSKWZwVk+nHlx3f4RxH
Cx9piK12lyVY5T6ekIqD96YhXX296pskd4EplwjX0BsvPyOmHYMUImG6BjVVib31bSbYNJzEyDiG
ZWVDn/GWn/zAutlUojVsWY9JmRM7LdWkW5nTSr4zr7ie0GvLAvHbIDNqySDiMdrOnrLvJuR4qgw1
gFXcNlG5zeeqDet778jSm3eLKyT54tsGZCiCHznl4IuI+AmO8IlEO6CTDXezJ6ghRm+lI6G676wl
wmJYp9naAg21zKVZcx82CBGGXQS901KwlkGldBDPitCTSSzUYr30i+w7tpp1GCr/7pOU2tTLPx98
ZrNEM1MwULfGou7dfRuwG1kr3aW2cKofhwiPzTgRF/CjXG2wlaKFOw1AdV3an320k69F7ZWG59ls
cUUDYX+2OSsL0A3vsEKfrULpUxRR/avTJluwsJdvT+Du8ztQWPfXOibnuih3Zvvg1/H4rO24nFiG
7OJrF7VFH9cuzvKuQwH8BEf8uCAE6jJGmSR26aLLkaZdQKgVwGQ0/xqf41w79qcwDfCggm6QLsCH
bLmkT0XmwNvQazSTgIzksGKVM+mEhZ0luhxQXmlpkEpaXyW5C0UA3Q3B35VBnZMmWKCxn7hjMAgs
C8XqSke+A2dy5PZ0Uwng71Ae7X6YY5jsr0Rqqtdg4EsGyTC42HY2gJYmkEjC+Fih3LWwBkNu7vkb
gVAiUg4KHo8/CyXRrnQ/yXQI4Cd3fPF61MZSMMJcHz3JJ0lXmiHkG+h0sVBLq215KFHfIr8FGV4w
u2xTYKG5udiaMej/3cMJ3FKTHrIHC1rZ8TsCwO3yVpV9gftOTXecAQcWYPwnjAz2ULzJ8G+0uhUd
UWpXEKlKFyZwD7Q9LkJsRQBPARDgPO5XeXD4eSuUNXp25RbtK0Ga3b6oglHGzzcX6m6FezURKIMY
9zz71H4P76pIp0RJFUVARKmRdS7uMLBL0eCn9DxSXE5y3PHyV5eitPUzRYOcL/hmxKDoNYWsEn5T
s8VFm+Gyz+QMCAwK5icyzxO8EwGzCHTCw8BdIH+mxntuBocfNIFsvComHiNfBoaJALUUfUey5vn5
aEhjli5B6slhEamAeB94mTi20s3kG63dZk+nqpkDrUaLuLTnh95FmsTWxZyYKBLcoZ/P7HEmDcrd
VNCD3ahTNQiFFroKKDgMR3LwLbnaDk1o1l9BEkl6fclUvAZPGoIWJPOTYpeC2xhotRG8c5RNqLFY
QPwZJeXOvwr1hCJFCMBjdJn2ziHYCCmwMrRVYdVQJRqig4HD0iXCHlZRijyzEoOhrTuenDaKBFDL
t2Ic8sIiYvDL2H5jZaEhFjbPvmK6XeXTgYLGN+golWpTL4gNPoSxCn5dy7PgW/6btJOc00fQO5mI
OhSBkxAgq7tpc9Dp1K/bd9KiR0vPd5qv84RD9Mh6uiwRV5S642FNzQyR1wtWKHbZ7X7sTlxMGZjf
Dv6oiERtwL7Yjacc+GHzSaknZHsvQhAex/nc3lNJHB6UqvjnyFSdMWOv/ZoZvAjGsqyTYfLWIn9f
fWHTlXGzZo0mivDcDWl8f8K0V/W0OepENJbdWJk6TTXew0PEkM9AaI+FZPPc79oiaouHbKKKjNH9
CUEBASKJ9v3BFYv5aoRBTGdV2DftFz7SMi9Cp9BZPvD4I6H7qYTTLuHLt8hpJ0kyC1a44d+HNtMv
jovmWXe9iG0I+3oY6WPm7YuUXok6A6eIKYSYItITKISHWPMeIh5pRpMbIs8oM5hdBdiyjdcjXial
O3uVgjjwtR2GM1q11e/7FqPZKw2FF4K865DOYz3jByIKPIwxe/IesuBDImLwg8e354ThtxlGhB7R
Ju4F9GUqi8x5mkyLkLqMnsr4mmtpqWL2bn4DvtgA/HSNF/wGa4U2DxYdjVDRFdd5Yq12DqSBam11
uyUiJgvmu8OS00ECjQlySgF5TKtumzkMgIhcmIniTZtxQCVLo5YydzW8aj6ZAxBxjjS85np/mX7U
aRrM8NzANlLSM7dTmr1vrB7hl7K+54YJsmXm3Dl3Rt9KmtFpELQ2Fbp0W9mvSE4rt/2qK4v7M39J
KozgXtOuV3S74vjYsKDUQACrEKIPldTc7GmzwMlXcBMRVLiu8Y2Mll/GIXs6xBBhyGjb1Vn2Hg4O
815BaHN+xVRbcQon0V/TUBf4mRCFuLARWwBWGCCviwSYeLHnakSckmnQVVny+aTs6HYYrrvSR2+l
Q5o3gWTGYaz9s+IchRBEdJx1KnCc4n3OTNItri3zB71g/XfRXeYWxCZoiRhJm2EoqIXqo9sQvd+P
YsOw6earoKWsnPQqWGZ3lxGNw7G/7RPTDDgyD2bc76zcglQ0qTS7CxSPfsw8UOlv3ex7wA+5vNfE
EYAlsqxCsr60D3Sxvs0hZDjPMSIJ0HtJXM1iOJGrcaJRHIFhq437x8SsSgjGySbDfp2Y8+hKzwFM
k0ZxEt9BUiPL10qxPQkGoOGmCPZCzFtNNfiZV/WfoLyWq1yTl3VHxhcJaLx+VRMW9aFn+acQfC8Q
EiUf2HyFkpg1z+3ebdte6YqRE/jmCN+hdoQw3e1q/WIId8jthjpJUXqNbSvJgtdsEZt9nMaG+sPn
sqMb6UcDODkJE7n6osD3AiHP8Rz87S9hedW7itrs0jpDpKBvU4ax1PC0fPBllhKmcJpZ+nqw85c6
AWnmch2ORXRSkTQqeD33MOZg5+3/mga+rh4Be52CgYnUdoAGpMnSE984yQNn0aqc1txEifgbn1Ng
3iRuij4dRydRlQy1OpH4uBrl+sCfkVj+JpQLR0zq/b9crpG0YzN+iIFbWVIkzy2/C5C6lYkvfIVK
E90wJHCUxFc2AsJPwVRRXUwnUZ//6PVjvA75YMa0megcPO4dRDw6iiZSZ34GoNOtmT5Djcz4N42e
S4qGTZ//M2ui9mRd8PoQrNzSbHKcerkNLcFMvx2w7nQiE6HBRDSnZh6FWDYJ/qdPXc5bUxG9XKBY
zeRNzjJ4GeNo+G2CV0AzstWCRxOoXxzpXPZkvoEnAh6DH+rxTm8tFQo4SEzqY8RXBFR4n9ijd/GU
IszwRUmxVgTDxF1xyhLuyJYmJ4TZswwMW355OmnZTMWpUwv2URpaL8ZldvojBmhInQGOaCuMpRYX
ld8MTfToZN25rrdS0b3+CJKMuC17lzcX52W6RXcU3xuLI4zz9PXPc4PFs5Aum1QhzUdjdVW3/HLy
yp6d1fsP5u7AvlufZpa9WrY+alXE7hSnaOVMttgi3DBIeuhXtN5yYI422XiUmCctfZMO3MHvsCxS
OOppH3GFhxiFSC5Sw6gH/4dFGHHATRKBSZ0PB+HsYA3LtCIT97/3ZA8bThIWszFJV9b3HjK3jucb
af7v5b26ll9CkD5kMh1Npkyudt/5ZMB4ze9DXwEfLIxK3g2qZVi0Bk3WgeFWV9oGteGACAC1ebL0
g/Jv1bmlkmk1BZ096j+XwDws6hyBV2szUa1Ubx6a0cee0VebN9JKXw9Fw2+I+psYfv3X0tjMhbzj
AGp407erafg4Y76NJ0wMKabBhJ3H68+eVizW/6XZjXWG6nwWOQ7OXjXNY9rTsQNVRTViNkleXyaj
d/k3c6a6zzzbl4PLKRxDbZl3e7McN6y/l+HmvL4YM9Rj8jZ7AqEQ4u1i7+LhkH2l+jFvbUmeuizO
abF+1Hm3dcqs0to1rXMWFenxrm90aa0xorZJLIZlnudy8qHqc2Ql3PXSVjIotnnUXC1KyQ8yQAaC
l9ZLFpTyBa0Gog87Lhvc6fe5M6hEvk+wINioTADFEVvkNolA/m54Wg/FbSTwCKeomiGhYdINTens
k9uepuPyMhP3WFlrK4KR5JpQit4YsAhucRgNAKUFXTAzuF0NsMJEHpXDKg/J6XLPDRznCoRXBsAR
PPTj7JU3LvwF6f+gImPK3kU3XIIoLTGl5JWRFoN0HvQYPJiwkNCPvMeZrQbFYgA8hHvaYkSDz4lf
lAgNamNr0ES8iiFDqUO1dTvvAcAc9EmVcmfTrDG7reLfJSqGEK6sf3k5o31mTnTzQYocx/koUpM9
smrrf5dPAC8NMsDY54qDtp0s33LFTAScLVr4Zd/z97cjasCdl/Jl5NbgBNrPKVMiAif26ILwnRB9
sM1u1ykGc6iZ3WiKMszNjmnnJFd5qFhIILQoWVXXXYyzAEv6lEOgmB1HE6/qCl+W74ujXpZYu/NS
8GLKU/xENofFxJsWrBzsPGNEklM4+1UprRqDYH/VtMl9YOcAyxCWTulIcg9uVpI3AP1Qt3RUE1dD
XGpiY1ocXY5k7HFVZEGNIqUxj3u2Q8Q7BLsUYD594heElFXN87l2ZPPkFbMYBsRr7v4yR7hTntSm
hu1PLumqOEY/Y17n0pHF1+aJs+z/5U1+qrg2SGpI/7mFbM2v8QQJ4ra7/p/hJo95aMlwUctqtVID
4yK3Ebds1bChpdKcMQj+a3OTbNBGcMOowwWsZHEwSZNv4dQE73JfiY/3+7htRQLpCQv3sRkAk7up
sHUz16P+8nQk5LtXk5siLDwPtSSc9scKWocTVozDUBmsla8215OROzSZlHqR0Y3h/nfbWMX9AX3k
s3QtGT2WTwutSzpQ8LEzTeSQgzfEzh4FggYtAm7bJtEhPEwNLF02YiZijoErc3geNWKJzaHD+ZSr
GUxs1vA1svgAU0Wou4FBVr1u3RkPv0ikIL8KEJyNt9n/Wkv1zm5R31E4tgilKPG79Aps0z83e0jk
Gu94USgZDNjqdre6RcAPpz2FVp8RMXCeOX3cEl2Dd/ShX3Oeji6RAj+RBrLN8vqzjrmtdRgS2uQU
fzQ1+N3kfczmcciLSKlcy7xj4nFhd+/oh4bDqoQiPGOEvTu2SdWdMSrR6/zo5JaE+Vw10Fr2ARrw
PE+y2XltdeOlyz5j5JMH2uNsj445eS069dqr5vAZauhSm2W86LSwoVWo8l3cBRobXADYrKyDKV9W
EyuA/MX25bsogRTnFNSPHMUZHkFZxN0tTRqByIB9Ql5rT3mE3rg4tatR31yg5/2V3UAKuxsO426l
l2lGRMwwU/ihGt+Jzt/H1WPUCdjlac1IK6v5dtKK/o/T41ce0vvOanG5npjdzL/yTN3tjonCD3yz
G4dx0l17hPKi4+RFTLM7gJkApBhgD8VGV6JrTI8m4ndToFllvnty6sdOZKW1uDZCcQ5vNXd5TKur
0v7A2m+D9+hYh/if8sxApJplO38nqY4vKh9rteZnZUvuA4Oyw5ZHQm2II+Gi1dwmZQ+SOhep3OUx
HyUOb68UdL/Xg35RyHuuALDC58mYi+EcrrnDKtpRoJL4qnoj/LOYRt0NGTB5mChRkcrWyE1/HX4c
3YzKCvI88hDuHu4N3j7D9uaQ9j4BkATE0ICd4Vmps/Ra2XfD7ofRL+YfudPhSOiOeJErXpu8kr19
s7yhR0n+JfXhH6pit8Z4dOPc1XTAEm8cOhxFLKZ15kWUnfHGPom4GkWtx9dQTIex7PAWV3oc2eUd
l9kCARgoqZ1Psb2vtChOwrYplAXvJD5j+JRlZmh37C4mnYy1cjz2/p9zZPybvy+iSJjh8EeSGc9O
IheTHhyFDVFu+gIgxJfh/NNoX0/wqOY6NZZM1tiqXNl4iVCJfvpxII/nqBHnt9jSgbaSzXgcBllk
6GLA6MNLRdU8mHrZV/nqe9FAFoDLkyiLpoEXQBllj7Sczy8ZaWZbahVeYPrRN83qY13cq37qEZAQ
fEypUoetsSrHTxCOIb+ejtoomuFjqWVQuakhhYOu+9nkwnH4H0vtgoUAuJas+2uw8NEtqQdJvHnC
VREfUPQqYr/BhqNtE+TGlZOVN99hHCJYkmyMbRjiULT1Ucs+BOhQ338aHz/leop7tBsyIg6ri/VU
lPWYINYHWVC4Tnbf1c6ABrmUNh8JdJNyT/L1BxLAv2EWAyjNwk9vrJOb9nOzHIGyd6ESAepjUeTR
DW6XeDHTdgpgzJjbXymZ7W4BdyELUODfQHR6E0iwlTjDc+sMGX8ij1LRNE8hC38dugYePrIMcZbc
cNKqJ0PNfCeyhfqCaAMX1f7SwuOX6DMD5Hw7hZx/uGbnHMI82IbaH0T2lD5jmOEYUV1AFf1TIsAz
y7ISQwpuwXz8D25Johs9AYYQPCsNzWJMRjRUq2yU9HZ9Ot8jquLmQP4DiS5Rbj6cwlPQGNmO8jBY
9AflByfnUkKAIplk0pqAMQvcoCh/EgcyxIO/dudeCwNUZfuc05FFxAgJyiR6eDfBCvzLggB9OTUN
dvPnCvUIZHyFCJArJ+D/50DdeCfDneZrxHGKEXlg1FK28tUte/ZZvjYlD9e9eiB+Ms/7p5zhg0In
mlITWMyoClb9+ez/9AbBG4TvSlDsicKYuSQ6TDQf+VfjIARimFovP/xt+QfTXp4m9y8Oi92Jcj2+
4ljlWq09Anb6Vcc98vYX/H8tzVrV6YjeGS2il+C0xcXGfGhxDeTyp/DCYzQf4UCE3WsAcHDKoOuK
b5b/20ISR7xQjJWpE+IVLUrA71M9guIkQWmVnesA4HdOQxlRmYHmT1fPEwARWLXRGtpwrLMcne+S
hcZ+xclAhBfziHWXUJCTQfZezwxPWH7+w1fGFIfUA89XOX7CN7IzT7ITlwptd6G2hgaeGRUotNAv
JJfB8e4u1/Csu4WP9+6w/HNV5eb6WUkmI5XCiLt9GFnEDWnEuRdYYfKSSAickFeDDMqJUCp8mA+N
/SWcnDTofHgY4HdXKJ+YfJh6WXkiKZ36IK4h2h0nXMXiSUQF/KeP0Mfjn2j84YIU+4ZTJYvP7wRd
KcismAzb0AB3o4MOxBtsUUyXEqCSIk2nMAg819X/qPDa5JU2OdXu57jPj2Vr1XxWxp+HvUgFInte
BSL+tjkIFCNu/WhoRfOiBL+jSbXvwkbsbPdUg16mhUXh0zb8/H0zXBF2svWebztiZr3YloyIY+nB
m2gnvjWBY+HvXj0Y6FYDTfSU7j0d1WBoZ1bFl4nOhRpxBSPJxyaEkj2HI8qweoZ7ZwkSWoTqjiCU
05qOQd4TvTwx3//SkGkDFY8y4HiqGfPdrAYTRVu8d8MgB7LHlrtbXbjXZk50cJgw0VxdNE05KOmb
sMzwVmm3L8p3CXAZ7HEx8izY88KJo0BucIyiJ3+dEMvHEFQx/EOzhkIa5RzBEJdP4I2KV6AbgNo+
BSdG+06Mf0e0abaqqNQAmWtApZlhfh02CgV1D0QdTuZGI5TSJVmp701yk7X8lGVsiwyCxnImH9zz
gqUv2XW4kWHHwuaPKlogETOVJcznMvqdJTFpGS6dQcqCco3MgcXlY6kBVhnwN51VLqC52qoECZiM
kqXvHoAwl/Fjk6eeGTVkaIOvoC1eGXyfEHPXGQJ9TfgMrVFkmuCjwFtyg73lzIXnCh47Bvc1RiR9
eYrMH3XYee2gw5IBpAKM/QEC5RVoPKery4RNVneaMyqeZtnCgRYjEt8ff+N2HKvxckFQqJHc7S5z
1iMQ+WKPLCFQUxP6hmFJwR+b/+3vXGNjRZo0fs7D/RJYozvzXPQ7GYoOsFekReVj6XE6OJOJnxSb
sGEDo2pi3LemTNbdYjFNe/xLVOTmkVWrcaB89j+cejsleoTJoo00TPTbBPrcUJ64o4/QPIE0OBiq
+mFTrpHrtJTrwIvk6TfWWNQvw7m5rLTs2yfNpoY+Yuo3rpbop/R14ajTX/Y87xb1ECEiHun0/nDw
aehcBcHEuR6K3CjCRQR4SndUyx3tujKVbNPgcKOE0wlbv+vlhkijZ20MlZOvmaWfxwE2i/SGL3RY
0Z0rX3Lo42uI2xosy9fmcmvJ6Tmvk1s4MwntD8f7faknJq/YEVas4n+EUZQngGbYheFI6HrAH/7w
TWpLh6LKEHr20VAFoxnGqFEr98fbM0sYQPMqWlZEz7WzTCWSdyd2KARet9/HlHC/kOTu71rm2eax
DwOghR01SGVkdeUIbNrWNfvo++3HcYOBk1tZbQsq1Rn4DGCGVOa0yfuhgRKUhDYpZ4Bu3JqKP97b
BNpG/W8M7x/39N5Yl+yyrOlseiM3YCpOOHqKIQj8xw0YgDDzbeBR9OCDkWZlfHTM14AdM8s/ps2S
z2Kfp/iA5Hk3ENOTaTmq8358Vlwdypn2mYDJ0uJ4fd6xipyHFhw1a1kgowaXsT1o9+oXrVTjFS0P
s658nIelN4XMB88rvZos7/Cnyh0xGPhDmVgzlDObd47ZVU7ftpZ2xONytqE/BOpnEzUIHO0oNIBS
TiRWATofgZkLfJG7RN+l++aOJBmBDcHIROmNu/MPPp78hsTgUTmy8an1jy+YT/KMiO9cnu4MCdZ0
MLS1XN56/VRHHeasbq6G/lfaUM5lpFinyZaj39RVU12TPBZopG/S7CVv0zRR2aemweIsdvyY8o2Q
Aa25nV9+94h0L10YyE170KhsBejCHBMWkSavryvT/kkSv/BG0zNX0jQEXuXjNcHNG5x9DIH3OT+H
PkQod1DW5gpnYzuMVnBRmJTpJaaH4fccLOOv/gKwG2wRT3a9TWlVuUtC0Ehr+3vE0sjNQYG4g8nq
sj6XfaSXl6EO9JCDY+wxQ2O7CAJlo5TRwteYBKOkOU5eMupmnqdOMvzmQB5DM56qkdg/qgTeESQn
L/sU+tbZ9li0hyyv55vBzpiiv4soGSs5yX+n12mQzXrRYiGjHhXqI5gsdM/fObPTOQSJh2qCTXhe
4SsUAJCxSFUNCLETBSOh5Jp/f4Hf+aFo0eDTvA4COcSU3//GVf4VAxd9t9wiBzTblvEsesP2cNcR
tQPxhID3m8EOXIvZySJnVbwqMj5Bc2dYfKpFcNo+q/R7i/8eH5SwMqlz0naTWsZguu7a90kcYxEv
odW91qoH2YtY2PWWlT2A4UqbKmlg7yIu+0hrEg5Pb++8aKCtOE2xdtg9kHIgDVtucGzbpn0LECr+
DSG+3R04/pFDm+3Us66ZxUcytsJ51av4ZZFpTXYA0Lw/AkDg7B8kcFIDp22Fx387kypFsXiZBjIH
LE7QVerrswUej14xbM2YsgpiBCh/w3WSjpsjRDMW4wG9B+a1s+Fdo0u54A3ltxVK32+nzP+H8ISZ
KGVZ0WRv9pPmLoEAC/VLE+vYWRC6GCH1z7GFsTph7a2cfrDs0zoppDNLMhRU+gefAdFGMncy+wqw
+MUuokuLFMlfCZZsvtyhFfgm11vwVRCgWmi4pKYdg4WK5isMWDB7hkUEYBEnpAExqaUsNGxzTKd1
BhSBByZva4LZUKgPUTtVOFIi7cr6G2zYVnc12hPEy3RyLo3SSfO76jB3VoqAr0bZDpW6O6HakWoP
i1lNYudeyTLKwVtHeGvE+yqBRf8kIK+OjY9cG1l29LvE06Vot2JH8RIWC0mQKgCUNDhGFMiQ1LMM
obHbg0sTPvCTu4wpQUbBfhKbRJ2KLYvaEOMB1AQihBls7beEDp8fmcf3gXvrc5rLIfPb+6WgNNk5
dECHvbKSpCTgBKsk1tDsdgFP8P3JrRrTgwAjzrt1gEOX38yq7iLdJAls/yUQWdHefpzKMVpvhAm6
pAfQKgnzh7ddEYBQZPCAlzE7Aczhkzo0aqjCrEk2UAFyTlHWJPkqQQNQQVu8wn89p00IZBdulDSP
cwN83CPoDZHPgb1iQUpbJ8bEOQf3sgNFGZp7OR1pfeZrfBHATLMtMRCEIyx1nbSGeu9lFv3QQzMe
M/6jUj6/bMFzQKmXNtcMxLWoTQxmud6bK8ivrKLi5epjaING4QbB5xtLR26Vsknq8QdIWZ1qllaQ
n+1E8RZzY4PUcf2R1zfcTULuAQmYH3OJ4b+Yf4C1B0W0++LuOOeJLz+hq8M0d5nEtp54ndW+7eZX
nXrxA1yMTDWW14Y7in7rYK34O80ORk5mHjKRV0ecCSqKJUUhjckWCLE6AVM2yzjvfglBatpnj5e5
jLVkwiQWIkftA7e5wWoy0khNAT8AV8I+EWr0MY6zA6Oq5FBOVRywFkXWdOlKw/Dqeo4lBJmiYLNq
ZOFxrK5/Ctpho6RBj+EQ5/HSACQYz2PNEbH+vmRgQCY8zoKqsvXLOgaBNiO5/S//Jq6Zn+h5c4Qg
+v2Pn7ldDULFLk8cEZgLPTny1gpcAaLvfDuVc870qUcNuEQUPuVXW6h6jc/5SmySZsI6YJ4rBEmP
Rc3MlSdwtE3mayO0onIPV8aJj89WPdWRidPPvnUVy0i18B5BDtVCuxtvWpHRYy+QzfdVrKFM6iup
x7Kg9+7tdy7+SF7iMYeAcKJATQLQoDGQZT+7vn9nwprb/jfHuCE/0KweAsQ/CHW9b4+BuMP36Jgb
XkLyCoKgfNURSQ/EP7P2hS8ukVV6HPOAPNZnJ83hu74/NLQgXwViisl7Da3Us1RMQsTyv0P6D4MT
UPit9MxBbNENzfP+k3lWQwb8bTj/yTx+J7kcMOqU3eANaY8cAWReRJsKTgoKBzyDqOt/KuHD5C5Q
RFg0iq7l1kyt41OSm5IxVqzxVgxpGlGWb3bLtm1DEM4I77KHgzS8lp4O/ndnFSKRcAyxy7+dLU+/
a8LU28guPZsN8NaIWLHDmIJ0aaTdGV6da5oIDOF8VyrJmSBaYtt/irocAwTJ3PwqD6q9WpQV2//8
nXzDOGn4VmuSGvoobU3vvSA79xT6ZAA5zY3h6h2yvSxyS5rLmvI2qtgYn6nPDiCSdw9g9YOD0CHh
T1WFa8/8X0pgterYtk9yhAiFz7zSTL3/QiSZUWMEyVAQPKTfzka4BWGchq/68jSZdFiIdz0XFvq1
i6yGE144SaOn3imAHUNeErjn6wCrnDw+VBjzxRJ82T7PzXIMP2JIuYVaiH0KoMGS5wjHQEDNeHpk
wMDIFZ4mn3vkA7zhT5clijov+3M7q0i3g0ke1xYE52ydRXMbqDrkCtZlIo9HFrGzoq3UCw58cV+B
Ded+PIWqIBf2gf11Rmej2ouZtghBMzW6R/G4mmkst9zxfadoCc5F0tsW4fbfGIBI3G8phEaqAJGA
m6p94xmTsvid0x46pvQljOHKsADm8Psksd1mnAfjs7NNcKvyO291j0/G7O0apgA1GDnoaHMr1Y3x
nfM15yRaBM6FMCXh4ENC33M+t00BpP8/CJ+uYQXNYbtfzHyc55rdsxnBpAP10ML1ut4VSLNThLCw
LsunsC7hPrxo8IdLrkVO1BxOEJlPK4v9PnRQ+1L5QacDW8i7zd7Lif3zY0NSqibXWRgzPA4YjHPL
Fyyek8E5VdcrZDwbZ1u2fXXuzC5qvT/MTA7ZmiT5KUj98kTkeUU+o5NjnL9Z9IaReTNovWgwzNum
KFq/UlO/bGqcZADDf4XyB6a1uMgj8T+DP/LNcj3YAKzFL9Oi9Il0ureCHeKO7GyLwe1JLQrzyy/U
DZ1AcgT27kaG5vZMt36bhv7X9hj/SxGUq2B/8vPgadrRvF1jKQvs9aOZVXOi6XpiiK9jn+YZfjWF
iSVZX7sx+a3WP7megoQLIQ3S7fvIFTfncIxGPsODXDip+kXQinOOInbD9x9wkn9zEmlURzUIROY9
ES1UI1hYTJrIiImBgqWN1a3wlR/r9PTQ5wP40MOKe5Itx1mQBXHdR/s8MMamCOzuSGJhiOr2Ijt7
m4klBGXuC4Vmr9GHD++K3sIONPWX5wM2qO9lix0nhHeiE6c0MKSLeRSR3lMFlJuIp5DjEjST/tkp
x+1YbAV2xFMT2vPoKEnPQJXxiQc5NgNWu1AZ1zDuhduWg7/6BMb3y6g8Q7p93IIOevvM3jeHgE/f
8ZKBa7bYty00w00o3jsZvrcN8HM31OqHnGKMbxDv3zGgsYjsugSs7iAD2OIX0qOR9pPTQAjo1IuN
CsibdEqci4XgW64jzCmhfUDrqu/ReTAx2ccQDOab0ifdLreUrRokPNyaop73FzcLOnA+VLNdDADa
tHgIGPip9NbjHX/AOHaO5qaAVrcqGqpYvyZKDdPu/hWajD2UJisQ8zaZgzd5FSftRYiopLJrHU3Q
WcmkjPtFGN+TZyTgVAQgKSQeuP3Y17l+5bkyt9L54KSFClS59FOYv9gaht6dSJG0jPfasddErIYh
xhBX+e+hMGEGvqcepSxY/v954cd0sbBnJ1NBHT1KDNJC/+oYBAVXV+26pg0woue3lTjLYYrHCSLX
DawuHToOdsKHvz9jdg3u49FOopc19fPeqKz0kYC9LZ85450mTWXY2NxrsSlNhv+oRF9OnOAMMvac
iYkERxdDPeKiH8UwTTuO5K/7buDnleZzBdO+KU4VUipbhtLdC4yNvmQAQ1DKf9yXIclST/nD0DtN
YNaIU3YYuF5TyskDZfX9fHNGRJ9JNDEEEOXJTHpcATXzyQlbidOa+TuLRg9++9k05ZP/LaoEZX2S
i/uVNYzZJ6S8b9cgP1Ew5Tqc3aIboKQ8SozQRWmsgWGpoJCxeM35deCVnOgMWo/p68xr8EMpeN30
HJr5KjMAbWmSrm4plrT/MX/d+q21HKL1+T5O6Klqojypw8gAYZT8TuOrNumMEOa/VAJ0NImNy0+k
Bqd4DOELudCY6kKL0QDMBNCCzQxdvGsKmhQeYYzelYELlG97KMRNp7LgJSOhUYp+JRIMglmSjNbk
wWdNZwmFijwINfzkRcKWNL6s2C2JZN8ooZ40UpBKTNeY5r2xpF/CJGvbr9WZtLspZYy6L0IGoz41
cR/iyzgMH9f7sTlj5S0R0Z66kc6miZsRp3dUrURd/J2haSh00Kddn4DlqXFUgb9ZVj7md51SzN7V
g7QudaaNaEC+yLwAuuRUnMHb2m4ppfRUB3oAKsAYAARFU3XoDHkMrr98GZCLoEMXQCBTxtyu4Mse
ueZfXf+gUEc1gNetlpxedtALJNJE95gvLydCy971z4qc7UjQ0sg5Fr0d+6XmzyYML5cG73zEM1vp
0gR7QcozKo3TnuqVUR0YgWtoRjjakYCtRJxD5ILQKCMrsnO0R8UUAzxyfx5mdERtZeNnY+krUn/C
WFYfG+yqaSsKxeXxDqNInOu1NLMo1YS/cT5lpQUaioWyLKf3ftA/4Y3vR7/5sTgYx7rFZsKMHQwv
fEvEZFSyfEZN8QNLZgFu89+xykcBzv4zATch4Ahn+UY68pwoTNkKB3G3L8Zbsp3DJlBJ9ddfyWqo
w9J+OTo4AQfl0qrVqgTZ2m55hi1E+e2Qx2kVrrCmh+s9LO48Nnns3W3rqn5VWDRr6fFxR1MyPTtO
5wlG9zieROVCvWqXgdri0m6XaLrxp5vCII0C+NSvAVt+NdEKvOaI47cimPb8gutdHdwkT5G9HT4N
YVhGkVXrfU+1GzxNsluStLHWEkKtGXyqd+2TtpmslIMmX+ZwWWZlLm1MbJmYg+mhlGUZnALEF8Tp
fAFHSudDXLd/JyR/Hm8BWJmV1E4vBF9UMTcYUX8L9OxRK5JQTM726q7AldY/zTxtsYLyCwqOwR6/
cpou+0eehvqWC0Pc1zE8UPAZQtJq3kbv8Ah4Em1DYNvFh40X9l2/7ikAbuJ5u1HYVxBBd+rtf9da
SxmxOYclk1WazXCvjWwORo+AEEg5xU1N7b7ZTE7fWwXKiUe1YpW8Uwl8VXbkVqDeYwVgha9jLVZw
pO8Pdo02jGCNJp42vCgS9oJhJwUs26I2TSZ0/MgWubUTY2r1a1R0ZR6Ow2MYPFfspzEeTdKiYMez
Rn52UO3w3jfHMPw/BXmQpUu/I+GYomvbj2TrNb6vrRJBDzrnQxloDsXvaSXnLMCzhT3H5E8hVAJY
LuGAYwS4R41WEw7JnLN4anHs7UAT1YuR5GEFXa3ZOyarrg9s/o/LJh39yFA4gUvB0Hu516HAux9u
kLatzZuRD5bFcFbyohw8RgMkjtBdR52KhjgCJ/L9TvsX15TaaPJ259LxWZ7yygCVoAuMFXD56HsN
+JUM+1FW04gV/jqHZD7sAV4wBoTrHpVXd6MgSGO9zG8x/T76Gn0Md/8iOrqH3+PHkfQ0IaAQ6e8H
7zwPK3AvFlnog6x2JNFns49TP/+NWNzQ0B9fhQ8UI+qz5KVCYRUGUZ0mL8n8umt6KTEQdcbtfMB5
/eOePOUZNeGmCB/yLYCCUr8o0lYoXj9QK3KEcQlV3dkA4AVxIQwIHRrjmkv9C0we9u/29jxTi6BE
kFIlda8v0LzoScQRnfMk3npWIClMhQb7uCSJMTVVAasuB/REUO2wLyHABmoglTbHTugQ2KO2qlq/
BJExW9USx2gRv2MAZ+lkRGqH5teWQSBHw6oBKBHJlX8ZXfAUkOLvmKhN5hyY2aSKWUQ00FJXlEod
abzZ1EJE8UvR/5mG2ru3wTUf/GeeQCwPktycAiQf8bTZ2UZUFaMzoZgv9OJKCtTCJITm3NvPw4Ri
2vpE5qvYI303YiiEOUVntdJ1TybojvBofWS58QDWtHNmzoOz5POMX5icS0LuyQqDm7Ilmj1MoP4y
JHErxrqMKKLRpt5Io9e1SrA23IJBvtn98cym4jfEsUQvOxDNAhtAY/5uLyZKnr82c8NsKj9mbf6f
GJDjnE3vxeba17IqlQaiQYzBz3OdRpK5T9RCervIakBbm+aGzt4DeF8rjlWaOUzhyTmnETsST4UY
M+1cnTYGKlhcDFW6VpSn+8ps/EOUSJn1o1q1tKoo5Or85hbYjIfV3PGhnOB7sPwWGFTgg/nwFR1w
5B/R87sj3d3NxeaABL5LZS6p2tOS2OWnZkTXI1IU6GdsXpNT47RteKdbyIncwKtupumqGUTo07pi
o35CPEi/vk6RVUmMFGmDHpRk5yD4mMn/ZZsxGKc9/Km1iZNjM3EgHUkA237wI2hjzrCED2rljuj5
1cGOO95QO0E8ifbINeFILXuoRCr68lIPat+rfbs3javsaPAl2b8E0fj98ViAfddQAt/e6yAGbmAJ
eR+36QzPzuYaht34gWoYn0pPfUWYN9f+UZqGh/uyLfTFBfZEnRh9bHzq6mN+1irLk5gbj9qq5yrv
MhEWq8VPNDXsa2G2Qg0JnKktPM3U8H6y7JcyA4tV4LL8gX4CU+EwbbgLshg+HQ3Yb71Ays0e8msB
lTBkyqDSWswoPAdufoq8bRbisoI/7QU6R7YfsUbmRrq9Ps8PRLUXuBqbfn97dSjKwRoGeKvGp7I0
a+lgazhFLiRdRdFDRoRKpDA2vG3VyzWycgSzPwd/t2SDjJZCSnG+TzWstYsrzIAP/2VCMWyY9try
M+WlmCC/VuS6NcfVe6cZ7KakdovvDnU853YBN0qcv2lPeHlcoylX7Z34mTNramaxNG2KLNdCLqrQ
SAZBxMN1ckvE0BLcquZIzG4kK/9y5pSp8L2VuINrA+vcdqPMNYOuKNBMJAnoHroU8mLhnXwWhNWM
gMT/gOaMoYuVYIIxQ+XUUYLolnsqWvjQh+NiUM0JWymjmTGU5DXAf3dkX2B9N9ovA2/AgEdTEQlK
CwTLzBtt/TFBYlqyGSLHq1B3Pn9NhBXlyVWT7GzO9hOK5ijT1jKgKHeGBqaknUnrLEVQREuK3nIZ
c6w1e14DV+tkwt0x5o9lwxfvKbyvKCmkEPSJAX5S9KIUREwU12cyMxktTX/+j+8uOPcXTUT09RuR
CAQBfRAd3osYI3GuYbCQA9qAiozd5crgWDz6RV/EKDgiexF2WnwetUl9gPqnWdlfSrHFlFg5gtJq
scy2dWWa01l2MAcxMcL5Kf4vkcLny9XT2gwVsugP7hnM7XJNW9y9qFH38FRG6GnSjxDGaI/urRpo
J67o7IKzk5sk0H5CDKjTG4isyDTuiUjKAmtFQHUAVfh64elX7vCQeoI81FIp8D52s7AG0Z55B45c
3ykSNCsvmzc1d3oppViIuAsBcbI5JwAntKxc3OBiyZN8wrYPuglJsvdcJ3rwcaq58dIyU5GhRVNv
0quZFEAs5tjHQlxzHuyp9/TpWJGb9xkgRWmTV91chQzPmjg6+cOySQmXM0a1qFcmcuyZQbu5079f
kJn+gjqmaXDo+K8PlnjPGSmT6XLxy7FEujRncIF48JT21YzZcIQGBO41kBd1ztGetjUdFz5B+3YR
uuZ0Pay/mKCnSFqaWwymST2d+nEjrA80GD+SMfMb1pupT5ydrfhow8ximN0cvKWOQtoc1x0NqliP
GHojwfZ0LW2VAn1Icuij474y4MO02YMYsw00PBRXdlOdNtxdoR69+oyiRIodkgWM9VbHpt4ggAI5
8tsBvBKV8wkXYXavvQj4U+sV9j+96oKCwSXUPV4gEOJoupAHl4xOctqLz8adRkukTAQZcLkvNLx5
W/TsvxrjVkTZAKp/6L+tf/0NuGO+TFy8u53Egl2AeURqbLpbY9bC/6y8dqdOXCvfpXnu264AGnay
eRKCLua6o6TxjSvOSv569GpE2c4OVZEsJtNCv3LIYn+tOpjenO7ryCrMFOx/IVIGi3Z5l/zxTE0W
Xlh+YtNYvzU+NlDpSdJ6Pd9SNRyS+/lOMIDEQ1aPU+bQsszIVapEdaj2bR5ltgb61bMy4pidDlSo
LhCgtbVhdDodFpF17zd7mouL1lDOcnL/c/qO1uEiBEdxnj1G8B6OLwggRGyHoLegL7DB2CCeHPE0
l7eJLuFTsVaCGCZr/86f81ULq3A05NQLuL+J4cWm4lmKzjpc+CDSwQxbIdgNvl3b8DgtzPx8l5Wz
mqTThOYqZaKRlpRjaPOVCtAh3Bx1lW0X2RBlTyNnp3BTYyuASfmi4+O42fpuU9bCudUVph1uDZPF
vokgC0X7IHAIjaGd7L8nZdtsJqhsBbyebsx4a5AziMXHphmsjvsdVimSd8BckrD8tU6jA8VKK962
LES95wSgQWGxLJzjFy2FMxIq2PHNIQ24wSyg+gtK3M+zG2mGXDJPxL+vNUvb7xkR6SpX6ygtDJPK
pciz8Q8rx5b781V9hyJHkYYGSsAeATv9LChLbOcasjVCG0wf/xOo5LdO+sbYUEpKokrS1as9BfG5
M/6ubHdCqrviTnIMzffrPGaidQt9A8AECtGCy2hxHP28M/Ef42ejMpY8yIFCK5FQJPpkhIvv64jj
v5wPeZEw/3e4tfF3Z3UMjb62KO/Au0f6kK+uhzDCEpBqm+tYqzsmkh0C1IsOTNqIiBtdn9snpC/y
DzUulI0uTiQQ85IDLzHspNzJV7CevKKqUbgf8Bx6DDWVG9py3Xmza0mZhG0FWda6astqIqFBDziw
X5chQJWwJnt+Xm8Dnv2ht4bb2uPNPqvccqHlyOcZjxnxIrElTrl1/fjRLMMuUKOhstqJHejQA6U6
UYC5yhMEy6qgSzUvUjIAUkRd0d0GRxCs5anZm7nPILe69b2yXGdznbGIh901eH1qM8heqTN2mmJb
NUHm707A4NyZZXoeEjc0sL8OfAK2C6uVxH0JJK3EoTL9hz+ro4Ih2rnRnSG7Zcy14gZ4yKVJSTXZ
eOaR3k9d3fqtVH6hUNV9QzhX3vkbxaVhYuD5PtZFpHwd772qu5jyZf2lTKkl9u/oBGr8bF/O2Q7B
utiGQ2i2aXXvLARpkCcsr55ydloFzMQ015o8epfHuqlS4jcA2M/U5/R4CR947PhmFtbj5OACz8xC
Wt4rtu6EvVbnU6bzDfZxswGY1yVh2aDI9DRbhH8DwHH5N6jZNGEARpA2lAKqz75g6IxCq+1XcF34
loP55DOB13pBmwEJakKqHbr77f41CM4N37TwFle0aYfsgJA69kF5lqRg9gidAAy+IYkzKBT76EP9
BsH7JwGpaeOOCblX1JBCYM2rA41Mk6p/wou/Ine+lEA70+dUlicLWoAortPgxzpMRMPpkcuyAjeD
mYP9wKZyrLnZPe2EHwzp2vH+xZwbj6e9mjg9db+6Tc6S4oG5pu0M7CId6qad9hDsfQcG/OizZ6Od
paOmqHskJ6Uy7hKM0d/Vhc6URlCiDudXeLwg/aDN5YvTXjuocoLrIrbHhiztSXeHX9VAMDaGQyFQ
QaCKgopVOfBbBaufgaL/wLX985f5YUJMaDWaXoYOQ2lGhImRlO2NDWwj22xGnxNDyrLcPuyaNlQC
1XpBNqYesQvuLmNIzCR9cmlRmpK/KhrsW0FCmUnSkeUEEZO+ff1LJdjVLUpGNk2n3TMyEgKN3U1I
PSTuGdoM4POYyo3MmXuKAPue+swk1rGNnWjyJZk9J3nU9ncZeIlO+rSBZ4Sqtbc4m7/rwtXDVLnH
uFQt0V/sRBRomVjmsikKI7NWk8JhCn4VHF2HnRyLAc9vM05Gyj/sDf61qgWoUBEr3/l9mDQY263k
AUXCMKU2LlGRZxfjsPZppkhheGv3wMG/oGsqJx5ggpg/mY+sZqbJNZq0uJjwJJl/Gd+l+Q1G0Y30
l0SKeYn6DX0tLbRdM2sz2GSQ2UJ7+i+Aqn4eSNDbSGm1C1f7/osGcpTkbmyy4M7IJ9IyuIcd4RT7
JQpExTGFtpcFTKdYqcIYbgY0v0aW2KDt4+l+PH24UPqA5n/9tcsE+tMnMpgOHrEQS/SxCQ0rdFxO
FavvZs3PnAem/QAhh6q6AInsQaxsfQK5Lu9WOk53yNN2x4nr2i7a/V/En19tNYqQCTDJDZXXTVro
FhyJPbOLLhQGqOrWz/r1u/5vyr/nP2n592mtXsj0tOpLnDJC5P0hXvQ8lbTlBwSp3UaWOm3S+BXE
hUEmQeC6ToesT8fejwF+GahVCWxr6GPHNaMntdtzPygJGk85o+GFpT5HagK4mEjXqP8FcdgPZo6M
xFLOxUBN2PHcIoAbfoyiJQon3VEbqm82vEBwRw0C6r2SBU0G70T52Imbh4CZ8Rp1uR7Vo83D7Bpq
8mgE4cR9L7J+I7DEillyqQYmcOuVIXmszIJWTkTqL8BIAPYWhV8ykk9lrdlCToN4EILsfz+mgcSA
YKCPzxB1RNBv6gHQ7SSGjPPbT7AYQQ4un7qJujTGgyaGaUjZsU76yqBoUOzaGv54+eFsrzg69qkQ
HiX1XIYZlYGBR7CMzmMX+d4LEyIwtUImKWDDmIuPkWez7EkuL7fkA4vUZhWQinQ1yh04Mw1VKR8U
CzJGDMEdAq1oPtwMqm+eMpaSg3VxBbA9cG9T8UodQ68zCr/u6ZkiTOh/w8vqMJQFs3/Qbla6lb0a
tHBolE5ULxJbjX8ZHHLpeJsBfjb2fvuXVAGDVdpXqDyoVhub/791n36gSpt5OulNYsLr6YNp4ngL
yynKlEDwApBSTglaTGl5NJ7OxnfGGXPLA0lrrVjHxa/Bd9Pf440NReZ3OQ8w1Mf7T4FdW5p9XTJ9
YW6bsepL1Ea9fe11JkzB5k8ktQO1DZvyz4Neaw/CXRzDDtgdYTdtwzeOh/wLHjlFNmSefot8L81U
YfQ/XUycm2nfvBS3bJHB/QMK25DdcTZ69LyMkwdByTMJfd5TO3SIIg+qSzAD4Q+4o8yviEiG+dG8
+ZYNLl6oHjtbRTZskn5MjDQ9G/54bRfTGrnjK71U44gGxKquvo9CPk7qleyBAZAIPvsjgHxImJqA
riPuiIczeRwmOFwvWb8+XBCBU9/XdK1Rip9tdcI4y/xc+bdX4OL2Meww5AJZVYNrwaTmK+A4ch1d
5TBuq6uHaWJDn6J+h+YQNp7sexWXVKygrSPW/2mPn22DHX+yCMpXP8hJSiwZhsLcSddRyBGgFkT7
s98W3/CEkHk4iLC1sw0wmYYP3tvrgYJSL/yjac1HZrVPB6+r4ltA+02rNI40YncLMkN0l1zOjnIz
PxGeMvtyUZ0tUi9ERiYYHOxO9+eACGPRcNY2DDW+aR3RBrioE5mPoiYpZOACJkh7Qsc1g3gmX1kM
9HrIxhOKKZN7NEirYzgIOHJE6t0T+c4bOP9DnoqQAHc0KZQLC3QLm5d+ltM/v4Xx5kMI8ajfpacC
RfoU1RdZ7cbA41UIGP56GyLn93kN5i5Vpso1M3wZux42f+mLo57QPuAao6z+EABH7zuBhb542TGZ
OOBwN/2/wjtiqNAkFEtvfedIpdQRMLGHXKXTHSYPVhuen4IBV+4sh7s2R2wHLPbnJHm2dAhad+/Y
22klhGa2UPTrxDN9xhdwbbe0pjC50mJ/lnFGDRka4nH0vmeVDcmEzrRYP0IomfaAY3vm7Gfm40LH
uzKSAxOn+zVX87+asrtBHdnnQhWRXUvZ9w+zHGVTjHtMA/+pV15qv9aFSKV2yrxRgZ7/1WTqNNcN
hgMdtCiYoamaiQ0xO7Ife2Sd7gSDnDHX1wSu9GtWEFhkxjG7YgwDF3i75LJnQSXqKrCCelCpTLVw
Ja8RXDOG+HI8eF/kTR2r8QPKNWXF9hwXTPTSAbZk8VFErELIvLwohqg9nj3s68DYMH3u1YLb0hnb
Y3bschGHDmlNUONiNmMmVKgUS1ZiqbTpa4wOJJtCJ69Vk7rafZJBQWeQBYQ1skPymWBW1YDHi8Uu
4C3BftIP0K4vpChJ+DUqLGDFug1r+1NQ6vH6BnojZEfjr1IGQgJwdL8te0F8xMMI4GoH3SMvBZmZ
Qj9rMtLqQAkWkV4O7TvFFDQXoZvi1wUw9s3vrQepG/UdBcohmq87ORWe7TzbJFLnBZmPbsB3AGmz
Fe1ZtxLbVXKr2kFSmSTnIJYbEcUlpbmSfUxkNijL5ospIKpCwM/2hdGvcbqroF9quBrKrhc4VERJ
IsWXYV00tqueS8EOHlTVCnUdwMRz8b/hfip3qsoVdaNc1Mx2iAqG21rWNXiypqceafk707FwYWy6
s1zSD/ikUhJFz0UDZKl4tuyQ16/wT5rWdQA2lYHh+Knq3tY0N1Kv6hU5bd9wERWW8pP5Uu1+ZMFV
qW2tkobT9mxOLYq0qzkNbB8ZwwPXjbSx2BeLEsCMvxjoYY2NaWpPNy+cDuqRsCtTrLx1JzNBPxgh
k9W4VafX4r2WriQC40HZAzUgyujDqWHCHnsomjJ8EXYHrE4X2TfYpEDwzcdw0qlApU237on1oYNc
mnrd1M+WQOGY17oqHJfhasX/AaUCdWc6H4Nj2eJvmvqfwvy70jGa3mVIFVjVH6CW+hyFa4mWnm/G
jfmZUnfaa+0zXaq2ldn2NKEQGum5sR5YWaPN9PmXZGGdc7OU6OZyZ2/2CFDe/3Px+k4J7PcSEvQa
/i3J4r71idA7Q5HyXfHioX7BZRXChspoB6Fc4So62VGF3REvCsnbNt4Ek1mkKvSDnXyscZqy+EZi
5FEJrjFuLJQIEzfOXS19tsYfItqMq2AOjFK6DbxhLV582tGs6D+ILwni3+DtyD+uBBznUIZzop5t
HdKhWUoiGciQKrKT8dh8oYBG8aquouxBHFbPMuUUTi3L8j8mnVUyGl5omUyRsrjfrlQqcewzd62G
GwoOoKfHWTjLgD2j4SPVfjXkZnHfkmg+Pn4a2DFs09Obebz0JQ6UJgMVVc+NSXE/G2PqGIf4aO1N
6wuCv2N/9RyBJe36ZzV5OrNztzKch0I3oSfk+4RAvyf4JWjoQXXknXpRiQVFaOmyaTREYKU8HCGZ
aNLcW1fCB4DjYmpQFGi3F89BD03Ly2VQC49tN9fm6sNPiJe2oXxR57aNHHZ1yhUDNTYTODNQY+qS
Ks6L+bzM88NcnKanlg1ZYL3t1YtFEYCT3yargPgStaWuTGJlasSLwqQvsVAPpeGgg34am6HvtiKq
ZRmTf8FlzBom3BReYVm8iFezZmTCprczUZWU20anVF99e3ZCQ/SXyE/DAGHaAxUQDaDn6Oq/060E
mbR0PLld1w9oXwD2z+2SbJ219mpJY4nule+A+W2MiM10xUfDJwKJq4Vnw448ewTdwJKZkzd2SuXh
1A3c6dfPfL4unWVLWWAr5EuOirdy2ByPBHBpIrbcJx7WeU7/acNzkFdfL6hAaYnCSeH96IPTPvo+
8W+ELYnst//cNgHr4MFxPzZh34/Mhf78I4NMvSnul/ZoBvlt/uWAHCRTlipdAkaVbjiCe2DOQo88
8+kET9nfDSBb5Sa6TPY7XxrCAhkiAVo/LqhW5sd8FKrx9Xjium2PVxCw3Kktvrh9TvkjZ59nrkLz
pSOoHKCbR5RZK3JQmyzjJiC4r5sbqO/mHNxtRnr5oVaKnit294dkxxSGYreFLjneJWjrG55Lw8SU
+a+HsYW04gJPIBSvnlXXtPuu0qOeXer5gnRgJ0XB8IUIhsDb1H2xkAaBUCeMBaFSJdss0FvZAo0d
6aYPrnJA2vk0RQtDx0Sa4E+MxjNpwyVRUrqNp5SGE0MJpQnlsd/5T38uj/L1nWvwiVDo3WkBsnvr
yvrrmfmcUuAEajKrW/GCmTElIYYXmbqRWUw5n4B6ug8Q3N1ijnvwIrzFQUP4QwLjts/KD3diN4VS
KBVlGS4rYxDcIyyCF3RIU2YHHrQkMKTkPhFSM6pFqhpkIUgiG/lq4G1JU5fQhEeBr0D04z1DVehw
fbN4IkFFkXDqXZCK4TUdKMwHLUtjw7DJG28Yhv1mWQtuHQb3+MxWLBI2uW7Tk6XC2Tw2o01T2bZj
OjdIXZvL3yOTBCcpNPG4S7aoY0KDjmWSp6mdAZywAd6Gl8hyH0j1wV4HkQmgw95KDRgbZhBmD4L4
BBgXIxjx3EwjXiwCqajdfK2eadYVAOpq2CbnFSDdZm1wzokztefae0RfcRcwrimvwCKnWq4tUrul
fpgs6CT91st8wF6MDMjGDcETA5JOEIxbN8nf/vewhvG1gcOctanV5zE649J7V6h5jt4fI4ljCoWV
bVrGW9yi/UhRkVROnVcPSsGA/9Wqb7aL1V1ekFRR1yPIC5WX+2GCO5CDhMVoPYjK2fhVfN/STV6k
lqleww4H7IPJ9KnIC0oSfTHZC2FbKlFnzzsHTCRA+hFclCWbWOL9lRi+lNSzN+TRughCgRasbG2H
HI9r3o+KomaF5S9RrDo7JiEHZGSWeU3VELqTWg+MYISmabkoTpdY3JljQzinoYJdKTdXTb9guhF3
B8usLcktBNwN4on7Ct+IvLx2xvfZ7aVXI3PXrUxn+OWPCDkFq8PdCY3DJ6PDMa+nHwKS3y2BFmFY
lC3EDt0Db2RbKLWbMKcoDCicv4P5FGxcQiRos3vMHcCO5lRYuZkuCXVLLgMh+WBlhh+uH+nNubLb
mjQgw9BZp2oxAeRxROANxqTPuAFKzypIU3VxrsYQ2JBGv34+pJIF/NcGmTuDkdmENH38jHlHBBe6
VVwVhsmcB9nO3L29AFiHuwI6xqJmpmB3c4c7QefKfdwm1lwRRn1r6Di3FrIrOc/+btmnHu99eAvn
YjidKbYVksiYXOZrakr/Sh4i9FjZQkDWNVIQ1eRaOi4fPuXNJU+i4ay3IgFuuVdmuq5ySWv9TDb8
1Gby5zu8KLxwTxDddrxCmdLFqnKeEAUD6D+xBWqXLsiZk6C/NbtkoyL8WItrXIpix16DB5j84SRs
+7sHJU0zRLloY1IQMsvrxPan7hgW78oRsodELsNSFHEUx6rlomZ6Rl24kUKeJsEOwlSsiurGEkIr
aNBBZLhX3qf05eU9W0s0B7xOema2SJTJ/JsQ8Cq8bGoHri68X5MYp5+hqTGOn1V8PX6tvKZ2jj00
2Ko2chj8cWmR4oTFq7f0E/CMuNajk8x92UxI8J7N60HJsPPO0w5YOucECdpuwmh+LhcHS8BO/gQv
yAu8t5kSzPWCPHClQ5Ppcc21zeTU+r3ae9IqryE6ZA225i4eoNLTu8nOsf6RJomRIrSkBOoUAV8f
hfICwed7luMf/tzpzfdUt8ol0rSM4zHYS1OE5WJyUVQje+HP/sEjEwbfmradVf1DO8sW/wPGZBXh
OlB9suZMNFdohYPzaxV3uzPped1s6EpMA+POC7Ve379EMTYkgQO/jHpmyFI+q8wy8/6FCSP53e0B
0z/B/y77O4xBlJX/n9jNfYSLKhLkBjaAdJYa9/EKFGAH9wPRk7nVuRWrlMl/af1S9cdQOs7xw2DY
BKjdzS4o+s3D6/DFfgvJ+75IsyUby8h4jr/G80KYt+dYyTcbTuqrR+Sze7rlamVCc4g+kRtpcWYL
ByHNfSnQClAyp5tzYW98wbZksY4g+58iKQhOt4p8DHLbPQOpvEbP+kJ3XDkHSRQzwzGo/Lu9A8mE
qqh0HV1+65kn1aUEKwh3C1iB4CtL0JV3mgjMlnDzi3polPskSLUkH2v/dTKhG8M2i4J1Bwx3InnS
YvYtQ6zKGbKl9hzbNmRu8HthaU+0pxsy6oyZ3lh7t3EC3cFVs2S52zCIPQ4rknIM0DkvTpaBL7lG
J8wLuySAdqBVFyLDYkpdP745IgfgIPnPFECsHAClxrajVqZe7n7ChnugWa2OX0N4Zr1WVdLcDGte
RBBu/7s2Jq9fq/AOGqvox5WjRP4vdWda0nIb+0KOIpMMH7JMyli9ucmoskeKkRTWNmjJ9LG4k7MT
f0hebkPGIFb/RkPzr+2+OeK1X4T8oH+o3pbt1OJmh2CqCwJrnxJapBt5rRJvaMULnr2di8LPA9OI
0furS4C0e/itqWXZblSp+lShkIkJtGdwddQDRY19ciWPN851UAl8BrAxKeILlgvuRuR8opzrS5Gp
YHTg0+bCtWrKudG+P5fzls/PdCbjC47K0kvvVKjCY9DQ9P+3UhKUHk2mkbxkiBXXSJo7rXnR/Ryu
HpxN9kkT4gMGZ4+qeszlQfmAJoXxHwf/HXyfk8puJvKcjc0NToTEhTEsdYYrMPe4lRpncs/cYO4q
QBKAqGOBnMGYQdW4lkSPx/+ngH3gKM4uh45L4Oun2eTga22NfeU2USj6pPbfohPIEuArIHkcRFZo
ATu+h9R0SbWer++yBt9wSwXUHNBkqX30A2XRkTcSNmyftR7Bm1jD0DwBi+FdMMqHKSOS2bo1eiaf
d6Njds+cClzC5V7jDLSEeQCeOqiJL6HZaPMWqXlKMzIyMT1u38/EHe9b/AlCOLNYxZrNxfvbJeyp
9WDpEat+7NlDEHkcpUDlGH5ypKSMGf4NXYMcBcnaWZi9hlu6i3hRs3Gvxbm5fU4/pxwib2yATYce
T6rWzFIxeToPTxrUQ/QDJ7kBqKsQbRhbTrQ5vjBQuw797yOU2xZ2oJxiDssuULifndBNHss+6sxv
TGAxaU/+KJ9JMzDUNTR+rwuGCVEepSGxBofRf7peY5X8YdRJ5nlQK569HDTKIcnDNov2GvCisxub
JmdWHahLbZ1onFjWXEsOaf/bmqQWhyge+Gm0TB5IU/mv42jSNczn9MSFMi0Zxt5qmv2es+/dGhxK
yaqAwe28yW1XoPnu9yOqIPGmRx8+SjsLmNMW91M+uniU+jqqkXSmKRSnmk6NmWZVTZnwVwvA6huK
ASoXiEzRXBO5YkKfQ9GveLWJLddEM8DMsLQBcgDtpA9RHwTw24F+Wk3dB4/shGtTXv8vTf5pPlZF
2QKEtp+XPu9ha9XK7mK+0oF4+ST7ZcOfag6X1bQUoWK1vs3YjGB8usYocgZ5GWkwBNiFrBSTGlmz
lq1oTICFV7gECI19shzTCz9/2ky4icdLC2CA3+IhEEMNxINiqADYZ/nMzcv8+QcXd3VltJi1QKbb
yg1S/hfHA0xApd2SMhn07YD62MJNZB6VetoGeCehPkhpaOom4W12MRkIDKAJgBa2bDYDxL3gIof4
N+QIHtr3hOjs/6mELaNehOa1NrgrzBf50eOopsg4PxU+hW0xXGOIxZAAh1J3B3PDT1Na4+HntiHa
9F3+dmPNs+09pYqTMCkxh02jc2/hn8NKp91Lmp01ad8Gs4GHS3sYhZBOZAeFcpVficfaT+fpWOPm
C1x3QSnEE+NJQZBWTyFhmVSpTXDrGVYWIDfxP7qWx38hIVHT8dvGV+zj70nu8DkWIb3po7/P1cFw
0DdpsXGUmmaQz04qYsdwlyaQmBGEE8Ilf3NLAinjwGUYQHdBB6i0dLxXjwbXak6/ISg0B5wX+Ve2
YS8WqOUsBifHcHDbA3G1XrAoXhq9/FDAlVvxvBBb4CzLgPZ0+n+nDgEATAUUOmE7szo+MgBGGj+2
VroHBkAPDIAy6QQUrrMzhK4iaCci7euVH071eUXZW6yknNCxNDR/JBM8mPTU2o9M6q9hy9deb2p/
2ccrFaSCmVVrBbl6E/v3T/TvCph9WILPa2/D93QmQTe6vI7d7QZ+jGZ5jsffXSwx7CMeZ6nEptcx
g9jqnH75oqYSoSPE4TDpRpdAjOAJQE1en/jGKi7a418CtE9zyiWw6HuPlx+TbnXFY05RfJk1sLI5
0w3i3zXJUZK1i3gDpdne1urLa+lpTtvtEMv/K7t14KslZqTI1ret/pfpdO4gK9wYYGnb97EJ+ki7
5+oivyqB44hLqSTYbrAcPhEAg9rvgHP+rDTfthOAT1WQOvFdH+aMFtcgYSxWcUAnFRva8tKgX9KZ
ttUtbw5C0ou7tYKKreKXihDk3095Cgoh1Q0YppEjMiN1z01HfRC48zZgoHf92+e3clHTnPa3duwk
FxW7ICe5EkjfJ9WFm1S22Xjp2G/mYCwW1tFKUUAm1+UBkYVo2moLEZW/uUVH9OZuum0oFjH6ZsT0
EZP5W0IceT75KR5qvzrAC/H5rRPkHuByxpY4z4Z4WL6qytKals+7qB+kZKotQGbbN1KOSTw5kQFC
cbFEqYUTX72Cz0VyVCrgvmP/lL58Owq0W8liMhOH2Ia0TbOiNcCxf60mtwkW3hRgsjOaaAYO+dCZ
yWwJRG3l578iGvXe4r+opqQDoAY+sSjShXBX2SrKMTj9LrAnyuedSCzHJgaPdL7mtrQRr1Mg2C0W
6eufNKntXrUUliUQDfG4psZ1V6q8Jpo/TyiawPoqkU9JHe3Ru271yWuyf98npPTlX7K5L9EgzxKB
NF38+KQlJdvgK8NWJwW0vOSpjQE+245/MUrUvClhYI8x5ao8aCsA9rT1nUnHnFPPZJvC057QIN6g
zupAQe2ll0pk3AZX/zZoy8ayv0dHww9P64Fw06PbPgS1MnorPvxrZyVLLWbPa6DB90d9ZyQCgwiJ
DkSiuttUpTEKSxcwzYwj5Mm5mTYocQbSsVVhc69gQpM3F+cxRS/MTWYwHZ/roPiyJvJxGtZtO55M
f/k6kKBrUhaS7tMYarHL7kjnYBebWdV08xoFAKWcsqnxBwlQG+vpW7gdqQU15F6QYzEdlqeE8hqz
pG8ZNJUr4sihXI4qbE7veXhszS1EVmyxcdMxLrV9/E/2EvsjvFhrndQQ0LxcDXFXyilrDgnacPUw
0nM6LVWrdoXShjNvpw0fVJ+dvPEHzUWz4LDXZVNTlUew87ILigkYmwVbghYWJvT7BLJVR7tSgqyq
sFvIgcv7qQ7pMmOySxeLFYwJEutZurnm7I0tfNd7WMp7LdLHudfh0nmf+9BlLxBONMFxliAsEtg+
pzekjTdzwcHfEZJBgUyscDoZc0aQ2I3GjHWfexwcIM4uk4wEFAkVEoAFGa42fe9kQWZZBK8QJEd6
UtInlLfpYj38tIvbko/gb0jJlmz8mEmI/Y4Ey3bajPJc6yIRvWtNWbO6KaZr1pTW/HWwfY0lQ6yt
MmwbOsmRbp7hK161vrKWIRrElofhMrZ6NWP9yfA5fVhBJKh8UVm8UFV63OPfH0tvpjk1nflAGcsu
W+4QmKDfOtiJxilAX0y+iqBEIFUlcZhBB7tWCZkNJOmuzJUktMIBzRQzm2y3KYmlF3c1AlWd1Eqw
sy6MXVrTo0X6gbFxhHtg/7t9dx2u4xQULB7hxmuf/vF1mMsdzv97CczuTTt3R1GgnHqzQP7UP/jq
WgoINhdlf6ziqOz6y6f7ZA9QYaO0iajKyOvVcLgQREpJc6OoUd7UjdTyVBty3LiN4pe1hxEh7idh
SgncpPTkXovF42BeSQZ4PTspE7b+EE0PoGgZqLJz3h4Ak8BpivBdgF/FzGWxe/KnaHR4o7qZuBfZ
XJC2noIOuOrY/EMdI8wr5shslNTqT3o/hCD4QXs1X6ay/ZQ210ZAzaGp/1R5+iE6UBilIpAb8+JG
Dcaltfj+4WcnteLtzLNiSJvFgUJS9K5wkpV+eFfBHc6nPxTJX3bdC1jeqSwFhQ70qq3TBD4mdmFr
h1fP8o6Xk8smnwb6+zI4ikCBtofY+Mg8oxzdrwB16/ymE1s4AhvHGkVUgerlbwQJVT45C4UCNt5a
xfJwCfRG6yCCJZeHisqU0CKQUEtnEAOL2Cbuqls3Pl7ZDkBFl3TEr4oQaYqqd1gyi/7yMp+lvais
LMtLPP1duUeHxBzKZfkt6ni5dUHdja3FYQcnNvsLCnrgxI2cXWNgEtiLJJdLCTOPqw4PHilDLnvC
zdd+BHXjNt9DG4DCE/aDPXOmB4fVqyw6uoDZ7wA/2LGhOSyOviRkke0ZPlnWanU3h+06KATegpCp
m9EK2Q6LJY2Y8RcDfJVMKL6X1kPQZwP4jPka+HwgLwmP26070wrWYA+0VFena5ZxYr4XfqOIUoEy
R37lQ43Z4A3gSO/2V4pv+XYtjwXXuE/YAKzpodDA6EEWmUXT+Gt44ghvM9OqE1Um8vW8sSi8pUh1
ES3OVbOcQySXwos6S74lEE2HguOhPYAR6Bd/RtXuIMm3AlP/3MIgVkij458r5QE9WdvockaA3YO7
/WuctuEt39oCmrRiyTmJksQ7Wyr7z8dvKaLQi/8DNWX2apS0YGuiXpeW7uz8qqVltRmML8g+hdHK
6eZGQhLSpxA3TD1oYgdg05bd1z1qZVuUCfbAoump+fu7M+g30FKlpXvISpvyX+2e+6DlVerNppYR
/zEhmv7eWWE29m1ilVsjH7epKAeQMYwmjZcG55rcWCWTP4g5qW0ITanc1BKGq4pspwcniyego9as
RfAh5ctdtnb+xWLq8vhPi71rUFoeGPZdS5kp4nPXV6Il6tt20kgHNCDs5wylV8UCQ2JG84A7JH3U
TuYwA784jEQRqJh7pdx5wI2FN9S0mb1JGnLlVPhf58g1cEGbYidZQWOJGDlF3F5H+FfPpqtz7kx0
i2UwoHyzeDZtqi6WEkHwhKtmHpINLxm81r93KwU09oaY6C0MKJ5ddnSMS1vUxkiBT213kWbWKzUG
urBdeSwcZbucrjmmStBkQWKdBOCEzk6oOaB09aZWvjXdeinGB3mNfBg6UqEb5kQP7ISC/6X+si+h
8ojD827l4ahqitdbnv/4q1Oi+VeJ10a5T2FCNBMIo+aERk08qiSxtn/RTuYJvsoIBrxoXMsgYQ8B
k3aCVOJKy5fnlpJsvsH7JDjFLDVGwl7uh/E9szlwuPYVLTJL8ySM0l02FwvBWpjYIlxL597bz0kK
Vx1SLFtQn7mfb8az87gj3nPClHStI/M1ODi8vwbP+mHnHIlxuYu0nLkJu/y0F7nsHR98GbqH2lb/
cQw/PAmf/LMLJ1W1Gft/2Xp9+a3WNFbzfsXFmsTXvuqLYrjLhSdaCOguNvfpESlJT/gbw+RKbSnY
sO+zlGtfwQ1BLhAOryWjSN5oMXaOjSPbzgChNJ7GICCxqE53E1DbMPrc0HguF5eGgIcHiLPY0xCZ
bYxUExf/j0f8tn/OGDgC+Fp3x5EkpkFbs1HHOvF08lp97XtcBmNFLbBt3Dbi57AOpTYT6qdrr0TK
/iBTTl7YOBBTSJxJPHvGR3AHlML6MGTDTb/XWbMPIPPtkSyZ2KnBAGezah2ZYeYOe9BsuLBU+Z0G
g6ghIsA3CdiUDsgqciYH9XPyMQpKx/WbGK2nmeJ0xiLfcweULU1Sg630yBHtugoOfZ31TJkFv/iy
skiF+2k0ESmjes6LGiMLaE7T0tAn3+ogCnokk3CETCK60a1yyJLYR19b7OhsnzzzLyjW1jT1j1b5
mc3PSeCPsNuxonISo5c2XMLedbKKMTglI0zPNiHYJn5gLX/YdyvTQFsyzqEYsZDAi2hpX1r039qO
7LiSJXd/rPmByRoxcqqN/vwUO+tiQSXG62b4l8eHstaY0qhtHPbNXPB1Utdh2O7AcjGvPkWt3JvY
Qr/pu7Qtd6dpwpee/hBNn2oleRJMGTJfJ/ez2BFq5jXIYxhAs6qXKq3Rg53UQJ+mpK4lRzCwVxZp
UPsrMmGw/xy+i++wGLpvDqIJJHxMviLu+j/lP7RXddSHxLIWo5TuRfDlsnEUJfT12ozbCdO5W8Hg
CC1ZK1HTs5AlAzbLjysB5cwMqQR05AJa+BoWZer4ViaebtF4wN8/NAz1BKJtjDQLzofrT7dBKsAn
V/Hy1fJxGnfFxJ82Y6WgaQPaKZ4wfGNr3sIlAX6PxfpmWYMl8pBNQ2g6xsG3Tlufb0AAX0KaIsni
+owqRhpk9TfqRgjGsl8MNChNKTltWqcAMj1lC6Xx17qp0GJI8Glbq9KDaprEaYkaQB+zlOcsvlDj
V0intSlK0qXR5bKB4Q9viPJt+vstWXA31277jBc3B0XwKOhpRojnduJlL0N5Ch1F3G9JvIlFhLo9
tAbtr8FV+mK7i6qxWYWBAsj08awXO/cznwBW5VtyQJaH+RiKn3zp6laTiTOawNlxU/Xdh1/DNMSe
Lsiz+IHocKDqvopPIz+iJS5nwsJhBqMKRr18rr+eJdB7AK1KOzAMBV2E63lckaE4r4YyONeRTIyn
buAW7ubuJCotKEMlf7/KczJ02Pqb4PoZd9Nvf44zPJPBq3i6wpvTNs6m71U8yMlrkHcE0q2/b+wR
9bMtR6MMxqhOnpon/PcLnXQHGKQM74rjMiJjVG5+zQJ3KPWNhD7GDT84RIHnuNiEv6pwNy+UAQ1U
GvrZOndX95m3iP1bhQkyH9/NoQ1CESHaHAPkzVeTScwHXjY7Por7mDHVEoliGbbjmb2BsdmCVoXh
50DU+9pxqZwq8vQPrOyPvmaraprgTlS8aubyUvsPazOS9ENL/4wHLmRIFwZsxPjCvR9tI1/Og8Of
SgselVxTbWt2o6pp0bFytSoOhPi2t4BjD7UrVd+V2kmCLpntXkrbCSDx1Fpg/jHPLGCsLrTzziYl
Ys7yWfN7qT/YpwkrtRQrCeUvbl2adPkcrQuHlo1pjGsLd2KjIa8NUy3C+RV6VI+LlSmQqDEi+G/Y
v4fx7wX7Bgp1qmg0MIFhJ4iDFXRW2BbkBgZT0+VIX8snkbDfAXBVFzaz7cs19Zzz9XLqoq+cyr0p
PvLYCelGFDedtqnFRPLakzEL0VhHijFDh5eRDPHLB0wpYz1D+qpfjL+/rk4xMWCKOGq4g5MgQbi6
WXanO13AFchsXdsbFu42tjOO7xMTVnjCATxcZ+dOla1vR23PYs21f4QdI5AnAJKnKxoKt6tPJI1z
dEhpK3a9bh4DNWPpInjTWte3SnurQP2jq1ICBmmgYE9IseqqIJGKQc9IBb2RJ3vNhHettFEPUaHA
g7R8Kn4KzPpkCY/JH6UFZbWcdMqINBVVlIFisU1yjfl5F0WWignRDBEIsucdpubxkcd418i6WwZe
MLM740Gg6pFPLMDmKcj4uO1KZ+OYDL/jdp2tQqUft1Vmgc3COcBmpxQ8xBR2Ea4m8RC7bcxZfbbx
5xTQQFdEaL7zKnHT50rYdQXrkldAo5tM09D2/wybxrba86mvQZU0k2yM1pZ74gtwyQH9VLDzrLnd
CfyuCDHrGx7XRfumWIq5urwG4LqA8BWZ0uzwCOUOju493Fo+8rpqclzWehSQs3hJac9Ino9KxYNU
yZP62unnntvsx2em+ar7DuBA9FYhacHPH+LsLjip9yfJwEYO0gmcNyDkmbQ4qtxw7XFMNFpw3OWj
2CK5fI0p/V1oBTf9oPNd5nVBQcNgqtM4Gaf/wtHWX+FnaWjV9mKul9x6ACmS6Z9nt+CS1aExUwSq
gQxYBlmk/i9vrQDR4U5ivhPHM+i02MGhO8gdpOQTDV86+qHXUmJBCBscw8mW2F3iNRevgYqIPD0/
MVzdrnVFsLkKizyjS5rIwSfkVlfAX8Sm5vvKiCum/kZxh1TMCwPlG75hKVrhmGaJm4EPP9m54qRj
nc6MEWqXRTZKXRn9V+c5gTbq+B6RLs2ygAah1kwx1KPuMaCvmuQhElrCM8c/H1t+rjm7He+xweG/
Pp5k802R/b+kMicJmMMILEW2wdjlRLjJRGO5eMGgklG3alriLQSw1Zrkgibke/i4GG0Fx5vAGT9Z
p88F2tqfNGf8kRMllW15XCpz5swKqaT8b43rSwJmsKPx6FmJozBY3FDIqbLxrt8zy3IT0xNlkV6k
aQP+JgftEGwcvOsbIRWfWNVUw8ClGbAnGAamq0/PKFN+O7AfsbUFfye4v6U41wBdPYAdq544mcPr
1le6A7Aw6kw68TwrpVyEakz8m6OcxZAaR+RJLOV8QWfcxkPwLhykohxVj/E5B7pkXFXCwOx0apaX
9aX9nd831EIYpU85l4Qi8VQXVP1NcKfsDKzHbKlU2gcM1oVrMjG1OUV88TYivMpuc+pEaYlNcEdm
0UDFbXz/EibsoTqZ5tW3tiYU1GlTYA/m9zofa3wAmtd38r8pQ4htBwqvW0t8jpuSuyUCvuxWc5Tx
CkVUUkqwa2p4zF6ivrL/Vfquh6SG3NBuZkyMVLO4e3xa0X+CrXEKiq7ofp9s7K55T/37i5sZxEcQ
l6qnHYJu4PC0nxTWO5W5mgJTNUUA07wv9+3bTwcAFvme1GcUnPFrw4Sg8cJ80VvFPs87uFDELF1b
9mEgu/xwfdu9Z98Zh+7ItR85RVgTjwGS98lT/i4bUePz6qAANl/VvCUpCa2zfrQDAnioXQtWmj0T
s7rLL/JF1M9Whkn5uDuUX1t3/+TYBhXsXTC7LF4iG7WGX6WeUTGLMLz83ilVRVAPeA3C+nD0Iz9q
py9UWgywpEC6z8m357FGQb30BoaOakM4udwfqUEoytgLGPAceo2bCxHA1e2Yy1y2KzAvQL5dXJ1a
BF+r+gfwMwj3U7AK1Lxvy7dUJaM1PDD8hxi957LLcpELFem8QTFKIvPABLCKWv97vY+BCrlKRtjO
UOJrK9Rj4kg9WGKm92PTOG3cfpRD9aPbfUPO1PXfkrRZn5sFngHYUXOJT9/YPA6iA8/Zf65r3gE/
88m7nF2C67TBWMf5dzRoEroDh496WGQR+It1VnbNTLoumAqOahgPzCyZf/bYwkvpvL8iyGt2lM/I
XabrYD3hqHszrWUaSyhp9k4M5dZL5kvOM8QR43NkwnD/B1qT2L4lLW6rBXCIzmgyaijW1vlNM7zy
4TKHKh4dSrwsFUvqcqJsuMwJeZpItU0KkVYcRA10BMEtOnREtdbNL4DIXG5NNp+QGF2G2IKHrHTz
CmaMij84ZhIpgDBVbInjC2kUcv++O2b4VfNrTGDsqBohj5LZN7w1I5qnEN37UsTSOsksrgPEUWd9
2MiHZnqPmWQ7PiRJ8HveEHkk8b+2C47uk6877u1BWDfu+KlRha8j3OR9KEfztnlH7iNyfu8FvJiP
Jo+fgHEOD02sxhfi8b1LjtPx9ZLuCNesEPg/J7wdaHvl70hSxB3fc+xeOJ5ZjeXDTBCvV4y+gzc9
aPOzPgsNj7g+gunk1EZHnIglDY9c+LMgVp3jeXGBvJLPlo5XhTAqgtvwjuT3HxeptTM/lvQ5eimT
7zcQf4mdjy3knKVinIuYfk+yWsJ5IkLQNbSrGxymCgmKbcyiMw8X0sN1M5/En5NoiBPJHre0UfD7
dlSmXPCkK66L8APmYiZ4nLqhY1zhZSSkZ1LSEVf7Osc7+BQPetWeutnm3f7jyPWzNFEVbSz4u4NF
ggNUmOV5rIjQ636zc+XBd/rtIKZhUpmYGjYA8UwYIsfP0bWHyElh4+etcKmo85Nv2e5ND9Av0Hdx
9YsLy+OmdYIcyzE6lgrPjDBJIVBHRjI+fS6ea68abnwFZngErZqsIuxdN7Rpr8DWhDaP3Lpo7W8R
3LgJhFhGr5wxF3X8F+NmlHkYv4T0mU8QKZ2xB0sulAlN5QaCTl1yiKoiu1+xeUIk/az9V7/OslCc
81dci2MGXb1FdsSh4DcaLqlUsWqKdov/TMRdaOgJXjUY+PJ4sQKO95tx0zDqFzqxYmpschgpxhxQ
xy6VHouEbKdsU5BvWWC8/htBqfF9kMP9GLKcr/Op9jfiYXvaPLkCDNGxfv/fy5JTHfruPrtkGRJJ
aZtRShiStI/R2ZRz/EKwk5vHJ6AIA77TNj8xJJ48ALNwt6I6l7NiZIoblspMTn9gTmzRT5TLpeSL
XASw/2lrlfbIQ6eitHpAiQFlOXRhjP0u+ZYeBWykuh8glyxwGQLSnCDQugs/1kVsRA+3ZgSsQA7w
9aX2bbex6vMojb4LuWR/edBfcG6A86k2fk2zjJ4Vo/1cpErMRLtru49tbn1gbn6quY/PBkEyXqnM
8YDYbss5WEQg8njs5ctQy9eV11diSVdiueTmp0EADgOkdZ0vcK03Te2gSCsWi3DRGLNnbm0ussK/
PQilYoGG33NcV4ZxiblO1VJ0RNLrHPRDQ4rC/88nxjTBaYOOacDFsVVYhmMb/tWPVQFVCIBNaaFv
1HzunKhYUQKKhzeUz5lwthGdu8gHfPQBfVe6tosFm11jQOcCWhZlLXYfnK+P6Ytl6dK+ePAfh/Oc
huK/RTiIXL5FyDdCOUnNExJJD3zd1hRxJi1LQ63F7DI61Uw9T5629rh87CpNipy0O6CSwxogpF0I
+qO/YqO+9MfadEzrBHTiRhWPd8VsM+PwPriDJP5P/DfrB2jatsSif5JYLzukfZk3+eYoI9L3/j/V
r+C5mSpnl1sPEX/o8ADYcFgup07PZaldjHw0Y0V+Z6jto8xVVvR8YHzvJ8YD8xw39frXEQFvKKZe
Vd7P22Dm6cjPKDtxPG7wtZiuJfOTfdxBbRWIbpX+ihWlNoPyfrG6VO0Etsu1N+sHyHDlRC2o//U4
ED/d7wOsVNiGYc4ruyUOwUhNAruRNNhRZikxNCMVoxtxD4G/CJpL/IxbG0HhBDEFj5cKdv5v4md3
yIsu5U5jGu1xSBzKkOCOSqavQibM/42YBj6xuBWkWR1I7GFXkUdO4RCToJuBkBUshqRLgf/ZDzNv
ADIccACNSRJuJnV2crdAQQHW1+bivI1Uc0Tkm7F+NlHm79Q4PXwrmoyoCS9Xb2uPTc0XXKKq/l34
tiCWdu9VIyNOp0y1f+OdbF/ID4W4IKi991ykZpM9beyc1HHRW9kAqSFasQpdtEkJ5L5QdAsDU6lv
WV+UlmCipgaMXVlWFRPjNrmOgp1cCxlIkp350ItAmuVv4kLVTVhdarA9m/H6ae9K2SOj08E35plp
jwosyc/xUqJiL/unl3OigHoXepWggSZPLzJ4lYoBV8X0oT518N2QpYxagz5aRvzR3SAlQwJLzamm
7gpC7ue89Q15BeWiTolIIboEkyJr75UTBhx5Q0lMB+H0bwa0FjT/mkCRp086dJBMSrT57wQhlG2B
z4oU+0mgb8VB+q46LpfPzyx18UGU9mGqNm+Ho+iBdQqMJ/PGXX0cGxc+cv3uuJxOfWtnVh++x69X
j7w7hzqhgRlTiX2mN60mP4dQZrHkq+TwprqavLIRQoZxvlnyptE7kJ/xiG11Bpkl2L+x5z5P1xsx
FcwxpQ1sEdz3Elq3qV9D7AUvaMfd8xde/RXVr6jBYSXRCeet5JIPbGrrUQFPpziFHCukmWcVjs6A
XxUoPgNtAZLgU8CY63GVYOsZoM7KNa4Js/3OwmhSrzBGmeiOTvX6UlCr+N9BDN+7wVQr2+VFhe7v
uPWv6Pg9o9E6Pt5hOVN/snIJ3acB3qCoYt7zjMnWD49o/ba9f2DnUJhiwlIdmhNL7iMAgQudTMBh
w/CvwZ9TlkSOO3Cu4SLxJ+Wr/6oEicVbJ/r5toDV1A5iTokBYekV/CdmYDqRjU7VDQAl8DUPAyvW
rwr2IQM+Hax/0fUo7r6W9TJWgeuHqm3bTE/2sqi9wE9kKDAqpJZWnnBfvez1c4gkR2PxtmAntdsj
D2UiUU0gz1GNpC5t2n8LepOhItNrvvi8zvhYEkQ9oF6K2aShBvTkyNwc1IHrFmlyLv/AJvC9P8jE
unNb3N2XjrNavx0PzRsFNPSOs7FRH8rGIgcRrN8yJvUw3ADlsLrJPsNxu+pL/DcUtQ8rwx7kcrdo
zlChW3tj4MVc/W8K2ybEhx0L7Z28QGfRj8lnC65GSd9QkKaDcDKuhI5BlmpIXxAKV549Qms6FLet
VswjH6WjrWdK0vqXSLkaWM/DjaXZ5WIixaY5Hwi82nNB7VRc03Tuh5L6gy9WK1+cB7d6yX/LIjcN
HB58CKvYXUHMPFPKfwqQXygtRH0KHjyQrRIuyu1s0HOjCjd9KC3pCoNeLqpdZsesoJtWmUgAx4xO
RXBhA+U0gif2xJBuE79ViOAqk00ims7A84YM3BXtyA8ZYujK3f5rVcijExn7RQjTCSWyYrzHDAnX
9ic549h6aCGWYylYV8/TFk9rUC2A5Pcy1zgXF+CcIeErNKI/2YRk3feNSNzSVAXZgdVTlnxjKMw/
y/t3Ro4mIc+gqhYnJNrPalUm3SAu/mCs1rz1SHQBE0cz8WEfRVTym8PkHdo/RfOudCPGgvoebwbA
6xA0H0B5jRcZgjrFbTCI1rGMvIhXlccSoAxGDZZexNngrXJHMULgZsG5GXWaZPzac6Mmr1K+pzJL
O9eU5WQfaAU2dkMF+n2x283FivyTGy+xAcA7u9Nak9eOvNPk6Itb15NW2TssRHBVQRVA7uSGleLR
+5VgLntIwA/VmVpOpj0uK/1taRXXPYcyCR6W4OAZ7ri0X45boLa4tnucJCQf4M+fVtRvunjhnI/2
EHJzNE6qCtkxZiD8EMoQc5f0jNxjJGuweDPV18p3cqd3T3PuqubSQal5KzoHCQ9h9X30rNNY1k8k
VQzAeMqklcUWPx9Hd9U7SiQ4GTxSPgQvtKpqve6X1z+wPUcZnoXNncdINCmHreF5qoQ+NCnMyR5R
HTn5oCe+uGSae+4/DZ7FF23vzf4RaGXwXoSM+hqQBwkKAGD7YAcugsm6ey4+5DX50gqSY7sCN0hU
sAF0jaQyOLmYqM39lUx3MRDyfWahHyrrHL91VYN1Y3Q1Hjc6i/5AMNgvHALAdh8He9VtqFVB6N/E
cW8spgTepK+dVUhaMyPzgj00RDRLrZNl4HWy/WNe7KqJ6UPj6AF44BtRhMGieiL+AVY0OmKCTLlG
JUWdVZVSzULG2tIuEpodyEpUc/X2s7boGibGXFMzosJdlFNCam42Dhzsx73LAWQgJI1XiiiSVQUN
BtprUODMIvkYzv5jN/VCvvnhb/7rxt/EGPADV3azqPpqtAZzt5Rnj3uZdBDWqpxxlDehUYB+Jyny
DWZ7VTbxeQD28RAntfPGn8LEg1Hg6+cflLbdCUSCKN4d8Lnjc9+hYCqM5ohPHQxA+Fbio/e6WvtF
NILzPF0FHUOZPHFhe+E7S3+c101uLhzeiIXq0Xr0mYHKQ0p0NqJl/1/+M1QaPaOxUs0eu5ufjZH3
O4aHt+rNyoKy7tJRCO8Nyls94iLRH0Le/Y8dte9/7a2J1JO02MT2OiR+q4tqkbb6/boSPWCC70b/
hO/hPgBKsU9bSggETjEQMxj9LRDWkydXe3nWID+abIZhBQ3S6H+IkjcEStR+LGeH1y75Fqf5FAjH
ytHpbSShvltZKlmjecW8jEq/4YwOglQwFFt/gKeoAF2PQIUlnRrlWj35xmTjPk6HSuHanFHLl7nX
I7Eb+Gl5DCayTALO5++4TqjR82L1gnlRe340cFJKY6K5bxPAcFKeeige7bSUcGRE/DRG8zmTQnkD
bb39pcQTIBfNX3y/HJEa+MBMdb4jsV/Ix/+ea/ehPjGrEBcJV08TAQfk4E/Pp6tjXT7RnprZn0S2
PVMjoAVdDTUGPx2gtUnGx6tXoVdpj78sTPbwdbs6uaIRRTybIilGxR4WxtbZTNXysb2XnV4qvtxV
65ZDFcGflIIPq6QwL10uvVn6zLPwY+qKlDEeqzSuuJLHe5b2rfiNOdO94bVAl+nbGYFeqLG26lUi
WndqIEDphGSBc+3WyJjcUtBsoGt/5CvqDTT6cyb+/1u6A918TSUgvwc2MX0LXl45sZevyFpiYi+8
IVdfxGBsMMYEfdY7xLkmpXDnGpF55ob5Uej9WwLBBhLanWYFuCWc5giJcP6x1aAC1Tx9L2fVhXnU
hUfqX3I4uwKUurmmMOB5zG5k3PckpLOr1c3gZBCBBES0mX/bdSUfK5c7NB5dljrrJYfiAnxZsxcx
DzjPbqLLAdkiREU2P3McZ1r9CfuLV2RXdBO0GwkF2RwhZGHNb0hhC8x51/ePI6uUkNXHV8nPcvR2
1QgN9PDMIZvt/4MhtagHpZxupDeQa1QxF55wxG+yJ5er2WlsCMNUis2auJOmqPg9vGkjL9daqwHd
VVOgl8PJCO+J1SOHmRd+lKgciykE794a8uwnqp3l5p00PXfZp1Jdel7Zsd05LATwTlAzAlHwaGZv
KAMI9jrGET65+pgncfuJ/o07FdzvX5o9kdR/EsnS69HVyXnSXbPNPy9rMkhmSsZH3UnQ6B0O9Ctu
4PabH4qONHcMGB+UEDnDdjB8AgVTdp+KAum77kZ0s369WnulPHpk2s/U9EEpmXOtj2iv7nKAf0fJ
9w4PwvoAykRJW9xC7rZxggTq3G7MraumIIP6vjqdlykRaHSuvaW6k4mmPrFZBmvvsmxOgvhNL5Z6
x9GSReSZwhwKyQjepVQEKANFK3p9uV2PDWAr1f1GEByyOqnIHcSZs+nFSb4sSOA9Jzo70vSW9rCp
LwiwtRlYDqOrXRq1xFivult4WPNmj7+lVvpDQj201b/awJB0bKKfTgH+twY1a7XVMdzkQ6d9+O+C
SLRIickYO4I5ZrD8Xui24Dusc7RU0sJOaDhXcWCTWYLI6gv04rW9feHfIOCAh4bimbDyampbjXm6
ruAf0AicHAVPdsMSkNtfU+z3gy1Ho8yQajBt1MYr0iy3q6hYdlNRy8igxpO8FP4RJLmcEzSCuo3g
EHar6l4nWNoJMtyzPxcnqZ0hZCZfojZcPqMQax8ViRVqtOZ2LVjRCN+sZzo3I4RRziCRxKAV4eEs
uKcSvT+46u4quzzZO75V/b/jAZ76lNve1xD6nrUfD9kbzkRE1fIo4X/tYpV8M/8n8B+sP3VYlJcu
s7cZLx99TQYRHesnuevvgrXa5+kVHytAv2eT92OPPidJk0Z0ESJGXbQbKwzgakoOfe+Q+q5VQbJl
zpgbukdypfgAWGdROf1yfVvpgqzRCC1OsN1byF3uQ6tiWhZCHdM6cfyPZv5oolUfqkxQHh0rr5G5
MpqyYGww9Igf9HdWcxZRJshrgf1lra94NycBhcrzQ0M4Vu208U4dgH/ETv9A7FIm/1JQ3L8R1TzN
aro/xO8enHZ+CLn1Qlaf/6JdDMynemFz+XnPVXrFD6qpzLh+1bd/Fk4MiOEMnSJVJi7oVmhCTTkG
TKUtOKhSPmfd+PLRfINu+7RsgjnpdbjrAIU6AJc+q9inVyXcpaYfB1lTtrI80rkCbs/8B3y6E1gM
nnboEteZSflyVqiSqYWiRdtkvalzBGKHU3P7kPFtWprfTlwdvP4ylOQYZRH+I6qJvg15sQG9BKO5
xwjUsD6QdZtHJIAqFvi66diRhlYZLjOGG597/Qwmia6mTA7Wl7+ytrwZRa+RjVOHkVzZXm4sxhDn
SCvyEFdjknN+oUV+I22ODNeXVaJr/hGx+RmfpiRdw3cPIQO9tnaBRrR/I7MJQehwKaUwHWc9xIh4
b2dSh7Zy8ibEpT3hFfGn02m8CM8M1Q0VHTBk7D5o8Cs6jHePt0igOz+CEb3WeJr5TiAnSYbEAndU
aJsBSw/okbiVGytu6x2uhKOpRVota4A5LilLhlZ1WIZ6ZGZ2w9rAkaC+e4CO8ThAud4k+GQalrb6
WRTj4W8fInIgu54crxYcZkRX5UYuTGiwC1isZ7E4sMvSwZoanDKg8RS76yMacp9b71yq0UIsCmea
Bug1aFK8X43IrWWFHsV2rdQXth0QUxZdC0sCMYLlxzOF/HwTeGYFawCiZY61C3ZR086dVGT4yRLO
4hpijajPYV5lH0raBVVUczahH6xufei3dq6PHsxMsop3AwWXUYtBqC6Q7i7z4Np+ucqgnV0Zt4BP
t9FcAkrbNfnFMQvaOSnwLGxTcGkcmeYvnNYRUZPH1PKEUvmpptA1RlG1msbwAqGxz1dOb56vy6sp
DeUJBW95AjzJ/vgUNtz2SQc8iU9W2Vfacvw441AiFDZUf+mbIaOXiXd9z1WlduSbwVKiqBGx1wGJ
AVOq1seeV3j8bNGRdCzbTRjfZXtkufCriS61C8VjlyZxrnk3oa7BTCfUkTw7W7H33B6YRDRU1y5A
I8PTtnmj04SH457+1d+g1OsxCxt3OWFGJGJ0iwfNvKdMkj8xCE+PEAJA93mw+PyzQVBPtoE7NC19
4oIsjfVs6I6cgj2X1WGMpQz6g74/yWPk2TQP5rzWx0oLc3DjxmENp2oqf6K4bFwjP3PMho4b9cPv
WXA5qMWr10EiZFaOppqUSf4RHCzwKmkYZ10zQH0Q14WI0+vg1T023bcmw8YmJKcjo6JuI4jD4n60
ThzEMRplb2tpe7mB35726U5tHCpQUWUl79zB9VOB/7TxEyQ19eXxZPqtn3cwf0SgxQNiycKd5dxb
4jFKcoLxyqHSzEj7l3RYF1pWqKE8enT9tyYkE/H+PeyKFuZKiW5Z7xuYuqlGwU5zvoM5kYfkoZR3
uz3BY/m5SqfArpRSwmEOfzr70zGNS3Ak+FlyLo6ZVqmLG20LfBl8VaonEiErVPuLFU2TU9/6RujL
hMxerj28RBFVb3UsDX7oyBYFWK0lZxIX2qaUYrCVGUpiBpSoH5Wl4HDECzPLQTgO33FiNuHDeeTk
Ep8OMdaMtd14vuuYummKqtrmMduZenETcl5RZe1XUDJK3AdnPm4oZYQM+28yAF1qGozRl16Ox8jB
0x+lqcuQP3w00L8w7nKlJNDbaCFAcAz65gdlpgGs+bIZmqwYDBArkHu5KICKz0coQRDyOf35hoqw
MM1MHXrLY27p0SgM4LPExi4nK7pYSaGvDDIZBDz7g2/rTwAZijD2utUd8UtTB6SEs71BQoU6rldL
J5tw1EFRJqfvqv8WxGWuT9AdorIwuKIaPEzl6CfL0xhwVKKDAd5oB60y2Y6vTJTcxiJTlNfOhv3v
bWSL0xTWECqCmyy5UdHsWfOCVMyuWF3NAcyUK19uyxge9I0mG2tg5TnVMpurm7PYYQTx5y12H+VL
GMTlrcyIMGaEo0ZCRethCDa6HKsKBWvgJX+HGrnC31tA2YYsK9YNmcDgwUia8Zb96SV2EBfX2mtr
L/bJ5Y2Ua0ucWHbLuK4rIjLzbHpTEuXXEnEmPjcKhcwt9ZXVBKDdiGHruTtRMz1kvvmADDOQY/yP
Y/tXBZ882Nw7xJF1v+5Q8YPIr49AaZs+/fkm8lTYo6b4u3MreEu50AktuwFj0mUN4x/k7WPYE/OP
SdEOrJk5J9kRgW+COIR5hRRRxfV+BuE4sGBXFX0VuQodzWmQGRWXCsf4u99CdL7DNowEPoqRDrNZ
xVTXIwatBQM2b69d1bkmfraPVOygqRO1uSuh4LYIRf1yPyfpHcK9kmhQJoNnK8kXMoDEtNBEu9pn
J9tLLgX8+/057xp83WYls7wPww6zcYw37DT57iMDR2B1gtOwkRrZ9PWgnqj04DFij9aKeYh6DTMz
xjshTczu0YP4jQJegBr66aAPOaC0gb9KYTxBGkMBlEKSSUlmDJlvp00hyZwk5lFz20+gPPsqK/Mt
lAFFwEqo4Sp2PvPW8qDfUgQBd0LzxdxMDo/tKxnuRv1snOOlk2X9NcGepJsMitwXzNzn/FK2ARTm
JrzstbXkM0uSS1srLcvGzytMu0iPpBQ68y705nY958Hc1lNyIfq7XQn64UeM2IqUFlTgckt+DUvt
b7cPm1E9ClQjWnxerwANgblbMyZctZqP1/zlyjQM4FZmPZYrUhgJ+fo7J+2ijWDLrZHHHVoJ7q8K
mRgMgZQgrrgDFkxPUieGzMMkkU2wDwpjhPYsg4ZghexDkXFodviBpw5azRa19JNauuHzJdKDBdL3
JlRTLxacljAQIrOSmlGjVfN45SNYxv+SZffV/M/DcOcpE6fUbnTkD/KmaTkLM2P0u3QW2ZuvvoWA
MP6wDeVGC1TPEU66n9H7FRikmzIOnloaimq3VZKw/2Q7T3loOxpeS87JibgZ67pTZribH5b3QCiO
gdEFuSizMIaWqFm+EGzemLIHMq/YPx9F2SgideF/rwj5qFGpnrxWhKcqUZhjJMp7ajgzBynLJPIV
+vglwKYxdLGTO/KUJpdlUW/jzSXyU13KZbLw+V6XOnAmaJhGuGWpPP3A6anKGwnLDqJCfxgiqCF0
P6b9wZ5TdWwRD2K3GiA5YuG6eZVO6Simq4noFTzqNpmvj0B1k8CaftRb9SJnRifndvIHIOyKViMm
X5p8yxYIJYVMQqJO0Xx2476DoRXOkd+NzrLwcbxCWBcf38PRv1aZlvNr1Qhm0v+whoOwjfL+5dNL
w1rBptePqpeQbhLtlrZSgiPtYP04SrRvbacgk1amTidALrL5H2EXC/gb2t7zsK66v8S1xfii+iKq
zekkaoM5HaKVhKAawWasXFVVXFHkumroZf+4/1gHsMFWwklC7824MHrgl8zTb4coWC1tfnonL1R9
rLjMp+PPvEIJ6aVdNVS55SvSbwufdajWiqMK5U79NdS6LR4fQbrkGYdb9EsTr0R6jKS7U/GSVtSU
ar4epmR+nRxMdBQ4IQp42QGfzB+hcXUz1GLtJSmiICYVW2dmS8ewNM/LcOyAbqznwpzhvoY8Dm6a
qfV0JhW7tT/GlJPHx8Nf4jqJY+bfU9QU5sqSXLOJtbVW+KX/2knrPSRgI5EWPV8kU/CXCH35e9GQ
13WHdDo3Gl73sun9OLxLDrERe27+VnLZGIDYnkqo793TeXtVAZLfNilyeb+SA2yXVOV3SheU1OsA
CuWabPAedmMXiiTSUE8F5ILduDDJ828ZJbOiQ47kaMfd3UjUQ52lCqaU4y4FfOzcaoKnO1fF4OrR
t3kpViewQ6edvP6ieq9Yh7c9IvHJblMDyj+HWSvlIpHTfHgAyj0CB7HzAAr4hSejDzjUhZKP3/09
urEgA3KxNSiZ3tnMB9jgjXW9OYk+hcV7AJ8gMpuPyRtZ2RL+I8HjAjDL/+gLXGW+x2zK0EcaE64z
JVaMcncoj3858Wu7IOTDGkPNqWzn0oXiuxFrRsFJiWgo/BO3GajUUWjTx7RUvGvVDsMkeaIOkk60
nXyid/J7OJfh6v9qHO7FRoSQ5OCrJRRTlaEol8RooR/YUkWYGZHtiJviFz5lCTFG/xJm4mOO+Phs
a+nEycV56fTPdxL5dK15ReEhoPzS52q0H6gLRsjw1lasVf8niADg+sRnagsxq3YxdeFXYKedDFqg
XlOqfBBBkuhd9yuAglRT7aVb8YGVoK1A35hbQBxlYXWIjZEfSI0cPfDF8DwABfbWAWbkXb9ti34U
ZWmuX7FVe1W9HTIH5rIf4dBhMz6uQD1TfTK6o/iylsDsrdYSoDy9JoufO2xKssZx4g8LAzTnd4GG
DR40R5VTbxr7KDMt/WaJ0ATp1iKMp0JNIZEWuzRv+AUAxavzD9Qvtz6qinRHaRaeLwTJCe2Lc6i0
botmZor7dR6/YJd+5vWc58cwMRFbaKCIJSWmQB4rRQutcEsq5sZXJtnxKf7voH63JDAaUIiFsmT/
8Fe87sENvbnkF8u27etDyibdyENN1GEFALy/95n8MUcdo9Abxk6gEKRt6eKVBPSVZGo64LXyupHI
Z1bf9JWlu8CMMe6K//ARP7a6IVVXLTzI/1GmhZR3e7doX/Qbob1zluBFNAHle9pKLT3lGT+i0Gvs
24OzPIhc6wqdqcyq6oauCJZaNKEdRRasiMG0jJzmTIEI6uinldxNs8uyAaNuEyjIIBDbt8cYmBEw
uHdv2b7k+u6ny5EUrGBEIXy8t3RfKNszgMSl7lwEEQzyMC6XcwjGBDztCOPZ3gj5W6r306kBJopK
+urKjDliwsXmHUqPseMJHn9PR2PAnupA1Uoy/k1XhMhPKYcJfB3SbyxZGap0am3kLywSwum42EMo
SrwZNb8PACCUOooN8R07IjSDoYDyjf4Wk4HB11fktndxPQWaRyQUIHJ/uLtEYPX7VftjiTNYN2Gv
y6FgS9M6lFv7cSklq/UzEjyheY0oBfrpOYbpbdECjJLOkGwe9vd7YGR0QU0bKYihQeNPbIXUNSg2
DhcG9mMhUHKBXg+C6BNZh1ZxPqRLjBz3yjf+OBrJydEsBRSvpqhxNx+DDQQ5y187CAid3xfomE8M
iW67aJuxCqRlhpyqMKi2RrYn4yxBjm+zSq9lqTFEx5hNA5i9E0HkN//7UqVT0u6owC+hUZ+4hgSk
c+YVoMUnIig5yOqU0rCXCuyR3qjK6X5LHdJejTEmCzZypSA2CE35BDn5AXAzojp8KLAnyU+ki8uk
vKaGL+uWWGVAA5TjCK3mrPMbC47+8o+ShFcsWTdxIez7XQ3DU6N0x7tsDWiXohTOef7zYgNrkuO/
6kDIkLVrPf8Fod5cerXSFNF24t7d8uDU6c2Prj36rogKcwZ3SOkvangNSsJkUp/SdD7YNu+Fbm/l
RqgXyzVK6GrZRj1YqBWOQEnWQqTdKeenB0IahJQVTLRCeEWcOngzHvTsDDxe6C6pkN1jnjBuC2aK
i5NVDt7/ys6OzCjR7kqg+zcQOU84pn18xiQkngQb9A4BuGp8FBkwva+4Fyc9GjgLFHLmlEu5og5V
xn3itSBi7iUl1N5DgcYams7bbvTRLLUSK9MF4Gvi7zu3kCNcqc+ge3dp1WQ6J04QOw9EeXS59n2C
7kxyfShfxmX2Sifm6KOcTK+beUFzMBQHfZYz+lLLeGCpuHzUQ4spr+QdKGB7XfJAGZi1fwIGU9pd
k5PB/MO8Pvm+BKb/aFP3PWUBNFuGX19iFUNDvQXWkyOdyffjtoXdYweRPi1gSw/syMwk9TMOvYcC
EjTk8HOjJqqfOjaPEtMQedIV31rdhdabg+duFMbuwO3E3oKKD14HueD/9/c+1Xx3aEMCtzPJORFf
nURvTMtl1Ja2FuhYfrfVsk1+j1K+Wr5dyWWTbyiq3IPd+i2JMurMZcCQ4BRa6n8Uw4nIdVgyJ2S/
58li4UyBGWXwBSyF5zAzGpEbfswEODjp4Sfd8TXLQJOpajrPhIoCONfg8jfi3LJa8XEx0PqKHfOs
wWrMjOKnkiRj0YSq2SIvnBgfk7GYoaHJT2BINpvm82QoV6iHdW+4nErR0jafhtpLs0daB6ug/Ic6
cm78QN5bFA4D0TIfoiHdhQ3StewUlqzFkE7sttTgzXUv0n94SyPjNztkf68OfNWW5e+b4ekd+gAL
XZswcPlbNGnYQ5cSgMcFQlbjeJLQGPigsYzQI6sWdERjYiyJ8+YcT4NADhu326oQxY5aChEbyJuo
tSp4vQ8Uu0+XH6RZxT2AusCyH9+KYUEnZ8IX1syjVddBs1pQALWrNaaPtb+9fcZYmXSQZyVbq9sE
Z8eKwyfcbpJzXxoJ7gdAysyWlvKNUqPD0R2VFilXS0ztXQMBzKQAZzRRk7cyTGy9YiP/UmbveMKZ
6oEfHXTljcQlLKGSdirY/UuJFuH4f1V7luRYXV0e+PU1t+dA4D8ZlsbRSEPPGl7CZKYQyIYBPeq8
tNWLOivPJJIlr1wxkQb3AXvBvlFyX6P6y8RO/uUmI+I9q00h96I1TBgFzlZv6TikpQvAAYiyrpy+
5ps4YiaNLYywCrHEEjJCbZwy30GHgfKkh7nJK6RMgPyJ05mu+cCeZaCsiKToMI2xfiW+bdL7BJM2
xjn6Eslla43oX2i3CBMrHZsxA7WnGSiBL7sZyprrUlWhKF9KOKXY+0ZTvpCeo5TGxAitrPDFfeiT
tSdjaRuEeMtYLxYw/qOazwX3hOd/4coQhBkJEGbqW1SxJmMTHy2vZSpwVR2RM/kL7obWx5bNaIpq
OJMuWix7imbSuasZEDzYS0c0SjOchTbali/goj3SfgK7kb6C1mQ8toINUwSHsp+JDLVZfCstbCym
trkz8ekD8uwwdEk3E40Di78IuKzXRwBpntU41YX3M71K9N7vTUn1coKavzthYpXlnazWPGfSxU2X
O/kuYLlom51lsZZNUXcTz8esklBzWzQf31M1WvOHgclRbwIT4Rz2h0ChyEpL3e4md3/xnINyYoiF
W708t21IATTRn0c3UcCOJqAJdviI8pfN82+opKXZ5g1ie1Un49qgqkf9bhXVb3M6RrstIGJLh+sK
/yL6vfraTrBQQl2xaZ99RzDuQZOIcaO+i8HGNgTHgzpL22k/SrJzfrFANad2OQltEucjVghZ3r0A
GY2O8qeVQzIZevglmGPLUknmOJ5YvOYT0xFftx2H6U9hk7ibKD1IBW7B2S7IOE99dgysIJb6smXI
1l5g5j5XoLrN0XZD5oemsAvm6FL9mofZ3Anc8aGJVJRWG7hdejS22+cShVmaoExCkbh3cKATtl6J
Ymxo0kOi3D4hNj8wfPXefj2KOsklgLQUHjfW7N5j9pWWCOjzs0NPES3atVv/m+IEw8tJtwaMiVtY
NMR7AcGNwvSIHdMGAtvAZcV1wgaHOQ+YFB6qpYIOD3rQhCW4Z049GuiTNva0JzRQCBne1tZ4rUlg
38JI20yNUrTmhIe9pndpWBOmAh5Jo53GVkatiJefkBN6PtWunZVd0EhZE0kb8Ji40gektxTnJPYW
M8j/gHAzGKC28wXAC/GW/8W6scvPhtSQKGexs0R2ydB0fCnDAJXqICkITp4d0YYXQXWUnGXZnnlZ
Vxl9+ECu9fzkCRLVjc9mn96sOvFfM+tLlv7j5WZUspgCXTrFPrRG+1Le9qpq+ug3K1+9Ych6Ya0z
0wzsHnQzbGDrgbQ9sOjkxit43IvETKXoTSdHejn7AEKsb/Yqd/wrovrQqNsv18VTH3oVr5x5tJnY
4Wt/pR6d4JopfgIFbbWye68xLgV4QC8rGjkvQa3mQFL7yQ50Ha9o4k/+KkB72gOWk1WOKh8Xsl3I
r4YVyk2+PR/WG2UlD+Wb30EOI6UddGcwU8cRliTCGQUrdHDpki908yfJO1clhEjPOKmg+WBY3gSz
JIRNy5gns6meIKT9rK/4GPpWJ2U7jBGL1J09hf6IKFs+z2i2KyOURKGHxJptXBe4+sEHVPzZVail
eJaVliUl1ollOUmf3/d4cE1tP9urRpCtaqpFNms5dc8Ylm6ptkUVmlpctCRntkI+GtPfl9oDifQ+
uV9iRcpCjwTQafLzA8CSlABJtDFtatlX9vgsvr3GUcCiMsPepTLn9L3Bb5BqjblqydfXriETNnwA
TP5B1Q9d6aQGiEtZblkEF7Zl3+Zej2AdfvyNDNwz13QfhWIU8rnBPA7sjMFaxG92dJON+H1u3tev
w4MHvhPBWjp+Ff6hn3JreiqmsSEo1S4nUn6fjk7wWUcrU1at5FZXmAUJ5BoDeEQGdRvqWvc0Jyvp
mx+kTpL+F0nlV3BMxHxBMFeqk5UU7xoOgU2CWi4MfnH7G/AvK1hhV8RbSM4eV76+kX2VzhBoLqDA
InAyoNGbOLtw1yGVopU0W11z+oQrbFm0vPU3s5RIrWGp1udQBcrzKhpkUi2EhJKzAvcQXgnV2NXd
uGsOWSW02je6ygXDZeQ2IZL1Ia3JcOWSd3WBIKzbkRnwOiDxbnBRTtTITw3o2pOA4XsCg1XmFZ9H
nGTVWEjYa5ndqgbNphQJZCv2YDsESQlWQ8l+ICEB3+K3ZXbnyWZQphfoV/0CpMVK4aia6G2WxHeA
Nw7R5KMcN+gqdDndPHuWTLj53eqI5HBUOAgR4+tTfWTpSKOBhXH17tCwNm8KfV9Ve9Ur1nHJEIey
zLskALBzhMPGd23PmRZhi6LJsAbCWpSoRaexGqAze2+zYMZ+a1otuWfM+UOTEWERasBbcDo1KsdI
fEbNCilzU8nFZGEIj45efPw+blUzkmioef/zE8dIX/wmDRRAWTMrEK+bF4sv9849RcSwC7g+gqux
sEDSviRFOMksABTx17nx4rAxagt2y+6ZxO53rlKO/BgBFKnhdZ8odLz+YCP582l1pgQ65343JaO7
+kBLUqjy3mLVlR/N9dOxtkr5a9rX2VGeFIOaABI5jy89h89Q5VEJ5HsqiQDm4KkXdX9kJ+DPhoJm
47tYRnrpEUY+UIc7lvxznd3zlVIPWu2pb6HZ9ebwv+9UqaPea8YLT96+Ur3TGR5BR6rsIPL8CGHK
27EpCdC7Tuszgg6+dCqNZFp6fo4oe5blEL6mZXYzuafMZZc2ylOE44pmOhq/mFvStila/a7G30Zn
vjLK2NlwewRrVBJQK3uexvzb6gp54a51O0a8Hu2sZD+IHsO2Hcz0NKaDPijq05SXLtNg4XAewZs1
C8u0ylWHu/1/HIonAANsyxn56rCn++UnyEl5FLm+bAk0YDrX10G6JxQj+PB3LVjQpDTiSrzyKNqk
yvRybVB6d2zk0Ja73EHIEhO3VcxgV9ovNihCqTGtV3nC5rbfJTXNmNzNAjmHtxINdnO5ly0uLMoW
xpwY3YXsf0dQo0rXKdTCtsZV3jvWQ/CcIlcwOGnOBOM964mbJvCrBXmXkeuOEuHLU5M/3c8OHzJT
ifR6KUpwhuFe2BPUgMyACTH0BISm34UgshiOuEtbGdGInVhTp/a1uDn+9mptMd5HidxJd3Jp5flb
d4ZdeGBxXW4qNak5bQXkNsf9zcObBPKvQOsI4OlvVPbastEwtT5arDa2icbh/JZA1Eze5Fbn7ClC
g4amS2HcDU4k5GEiXw+jN9eb/NzL/6mCC97iwOKyjDexZ9n3G3VnJiJD9dmVGMXhFBJ9I1BJu2Qg
tLgIlYrcVL4EOhcVWzp9obfvpGBBTmtXpKYgSQMKlSqb8AKLapRBhX2Qt4Q/9dvUxR/CWU5SJN/J
mACT33afmWVE2ykymfFlrWtZs35rne5VIG8rAlHtbTdZVLJsD7cpajUaWyoCDuFqd+THIPUFDwJK
JftJb3SzkWNT79ky4nPZVORsug8x19LKFw4gTjBEdm4U2+REgGOmuC3lnwNZRa5DVncGlKedXM8e
ieZHT5TgXLzk1WL+i+ZxGvVWt36rytnnP5zOT+wmK1JlwTUKUXKB1zrHOHetTcLtJbGGDwO/MlVd
MAN7FnaO5Z669BbN/wDrRyx9AdNVwnwM38/IjcnojYTtXwqt4ta7Gi44BfAW+v+z2X18oCdJ9goE
Xj+I/URfDyf0WvWmD39nhB7erQFaru3ZfeR+SJeSrVkx+EJpauiBit/4d2zZpZxH+RqXpmkr4AA9
P2YjJfgyUiMOALg7FJYgv5anP236wLCpGnamzbXPOYY3bqyqK+CGSQSNrWDgzLN/kDCqP5dUogty
7lf+wacWWF3Zc+cL4YdbSZgDubcXX/BNN5VwQUcLWrMY1lmvqnAYaCvJK3cevtDCguAnl30IIpOA
X8mqf3ONY5xB3mASaxc/frOsl8oyF3FvAImnVAveBJXS9TQUQcKueLLULkHQZrFN/quQvjTfvMOM
Za9/Pe/okMWnrgq6ntODwvcfCEgVw0iIVf+dnud3Rv/C+wnkDWoqkFMgrOiL1wQviCrmjBwbOXVb
xLiibnpTRpjoFTEETab8gLn+DTcg6vWOcoOWzobfZV5ArOO/XcaXFziATRY5Vjqwlltm4tl2zOCc
Vxq+82ncKKkHvKkuKh00LTUozN5SlIJODOAj9WKbluMI9k5eCbxVfaLBDOhk1qZelNEU7FEoR/Tn
0MvSJc6ZVUHKAHyBVSgKYzlKosRNzzeIHs1x9f/mihxkUlffQtWv3eJihHvJ9cqW9pgJIXDtC4uF
EW6nj8m6cq0jgN54tVvdTtC3ZuWqt18RD01mUVnHjRE88Zm/ZElXiBBFws4JbJ9MM8oPVEYuhTuh
mGtN249DwQAhi99MRhOLueV6avGuMxBN2gm+nV4srURfXsfFqhhCgHuGlByBRGl5+oMGjO98kvQt
Vrrk/YORRDSdLnt7G1iwh4zDX030lQ6/oc5coPKZgfwtVmpS7cQs9ghiOuVDCDYMO/V24x4cqrEC
8WhbKhhCyad/3e3mNM8k2OV2Dv5+PohrhEiaVI0oj+Jb51y/igLDq01Rnssja0j/XD9Dg5m785aJ
4jX87YcEzQ1uFdiqhdD3SeolSx/NahFU2vVsOQQSpY/Xs0hSST4U3elbkoqW9KOREAxhc5oYEMOe
lwfECkUEW5iIRZt5Q60s6dFz0vEGMAqwgeINEE1UGSIUYqoby2S7F8+NXIqLFBjZOzrHcHnLP/pL
7+ddS6PxIq2i8ARmAi30lu9VwVAsxdTqBy/sTBZPgpH9gsgUbf5zP0vwii7O8fQjPJ5GCB1MRwge
33rKE5Dxr+Xce+OHBkUtgsBDKOKlW+Gab++bB1c5a3lOg8RZ8xtszmltjSawN8F0mI7VQcM+SiBU
p5fWGJNgL80d/+llTNSPihDdoFeXHPMvsCOi/e5OZdHC4RkN+OBNc57TAC6mk2jrm9BiOEtF26qs
i6gc7kyHJoKSeuRm+XQu5iKlkH/HSh2IKxxu4/yq9m0vAhZkmDarH+6dejQ8xPlCqBD+PeOj6cjN
477YZf/XkA2/gP4x7dAktxWynZO2TlaNjSOrYfMjyUqeHFoV6d5V8Rs2lFUZstQIhJtr1Hu7OHte
URl32RR4n176rtc5vjmzSGu+sajTNSGDobDtmsuot3zxMQrmqKOhgdpw0KJ+Vo+Boe9bIJhpXFit
WV1J72LToOm0nBj0VeFfK+LUY+D5z3AFGyFw8a7WbcwL+EZ/Wt72qo2qkY/u/YFFJGXFpzzV54wR
k8ENZzOmVU+X67LVfIRY4DTqTNv28aYeG6WraBjChksfDX/F80IWkks9uWClYzzCRlY/K1hAr7SF
pIIIphKhg8nVuaU+Atl8m5XIygvvVtyeBGbI5yIwpU1UNadwUGzGiq6m15XNzX1kFeeQj9oMpHUr
Bm33/w955PWBdvB8bRZvRoGMLqf93IkRBd4H/XSys+42RMwZw9+ApTgeGfOLF278AVDxr3t7bxXr
c/BGlYDI0aZ2qY1z/cY5W5LMsV0GgMCLeKCYQCAcIpzfiwPGTa5KSnQLd4ofWfAl/IAUyN3iShZB
CUSvMpbbej8TNakuoE9GbevU1wdNQzJNSY49xBpO5o0rPi+0Z9CB/IaXqpXZAm2vyC7MQUJ5JBg0
EPlHlLtmfXQz9uv7gh7TTDfs2WeoDEEeoZ8VUCmf10cCJpvRCSSh8mVaozvDehKS1xdfjT+weZxr
IDnjNMQVKZnw9cklx8btOaPxLIUltAeLEybqMLp46HxAAmiaRUODfuGph25WOS4OCx3BE9qJKSUX
svZ2eUkwvQS8x/3cHPSsqC2dgaLorqQnV1VL9cnP8I0PH4sYk6+Z7YhzCuRDe2YUshjvAVFALvgM
n9qIn4trwYQWB8El3vOBlev9qEf8Pl9l+7h3WUQ01pHFEJKveKboCIzIBXyTdqVlVBV472F9M+uj
uO43Aq3byTKPuyLWqLri18sDnZsJeRtzX0h2DsDIBjiiPrJT5sZclk4YC0wEA6zjoOaw4GNiBflq
xdNFJtZwEctdUIuve32ROU6h5lapU1OJzhx9NeEhEtjv8jAcVAICZX1KMDwr2aa122u8U1WmBSbr
NgM+BtBKrcSYXBtXTNfzlo6CQo5AF0Gi13m+gSJrKLwwGpLMSb3e4S9vvSatutZyT3rz6KjGRz0I
9YJ21ix9M25cWeC+xY0rNvJekG4Mtc2yct9MeD+0PsvSaoMGSC1RSSz8YH3ExQnCeS6/OqZ7gwbf
zSJTnTDK493kmDUuxxPrg7a0QfC4aVvyCMmSK+8m8gr3FG50h13oi8xmv6F10/yyRZ6HvXLjBXYv
rKxNZQlNwGCnqO4OjNK8j7PwVgxjSYeCNS6ZblkKK5W8kRTDxJMjG/oMnHTNv0ERCUE4/P3t2BtY
Js6NN8Ml3964eSZKD11z0e6SFhpXIy0d+ea7HMFoHheasQ8IzOEC1Ims2kaHfDXuqss/bLm50Z0y
556loZfX1IOloa47AiOr9X3q4ctALDC9GcYm9rc1HDDr56HUIBY2qQ2lCdLyqzzpFAQq4GLl2U+0
mUdezJPM2Uv4L66A2u76Arp5yInp/fiDAk63IeBKM9I+bKoc5QdMBjmWOO79UyYCJHhPjgONw8eu
9v9nAXPg2fA5Pch5SIDKcIhXYsDa4EImnxpbOJ7pMYaj874B8zPF+qUXGys3U69dsileyjZF70Co
zO8BJb0qPjYc+Dzdds8Qs6rGrw5EJAq4+LgW8NGNLpRQekszIFHIyQLI8nteFijBY3nU2nTns5/y
RmQ5Loyu/vBzPz1hBehUmM7gsx5CDWwDpSJFHPeWj3pk9XdSWJzXN5on+cCfq8KxzL/ubfWn+rda
2k8XbAS33CdGUv2ieFlNi2MLhDbRU2iDFdOTmUb2/Tqflt8pvoh0JhffQfqonAiXlABw/+rJBK28
rmdx4yys7CgAABRmZhuxlDDBVUssFxDKP0PgHTM63QPOhFowCY18FEs+QyMRs3TgSTad9FIfc6Ej
jOegMrnNpd5YuSlObPL2K+YWax9dbhPFHw7rf8OnAEuNUsk8VW63U1fvcH721SkA8/Tf+irdnbgf
rMwf5ZOx9ET3RZPg4AtrrMPLezRg1YTHGOkCA/jC9W+Q2KR0jG/sAv6duRPShK3Yeu8fEpsLQ8To
Y3TrqQ+6YREMeNQXt0Uv1/CM19Cq9r0cJG1JgU770Xa2WKvbSWu3bJxtZgxXAKRFm98IiUpsp1r5
tErLR+nxj+/L7MT3tCDKK+qCKgaQ7K5JeAwB/DWQHRytSTWhwdF++x78xrhBoyRQf53CwGwHkRCP
U8LZwHOGdPvWqBoJC21IeRViAD/QjP1+vH6cnKMC518Fj3iGf6B2z/imtHy83+10lzI5jMmEL4ub
eVUAJt7I45Kx6Wj3WA08K8HbDr96oSiQ8H8ZA2W5MWX8zkm+AEabsIYlSn1qg31rPYiElLMDoA1X
4h2c5m5vQAHq5CZ0OXltxDHpo5LwxrlMQPh51bkKEscnM2QCECNJjEuACWDkerxG0/YsYAPBOe9T
wOmVK2y8MUEDC6A3vfXYEnqZ2oxNl3roV2jy5h+PREfqWc/udatZaQeYBWXG6vHBu5DecM/OEs8b
h9K3QnH5xjhzxF9Q/XY00zsdbjTs6/E2cxHwJV8ReADu59fbvxwFtzzRM7DxdxBs2N3npeSvtBLN
28AhI/4pAAxDfZrb9cP5JrBfu7ehs4jZJYjDlIDJCduKfGSKXcNu29OmY0qiJd3NfVn2EMnrdTT2
GhWTSTq8FIl1H+RQEd8O+xh2h0xPJkZT9f7FVZt/1oE0vi3zKBtJGq1pOKc7GW9CTT6+5YheEpzJ
6YBf0IJfag7yh3ZSxdXPr3zWm3x18bvZIf+6Q/nPakmcDJs55m9CS+fGfcCuXKlEtywqiuqfqsGe
9PRgH+zmOpk6SuBHnYsfqYfSmUEZoWNzYFbvlqC+pXuChKWYzZ6jgRu7XXrpAseiJ9uolPB6tBeG
utR/EXQC7GQABAtdlqdyFht8N5LckXr7JG3Tg61OfraCOntUs371SCXWIbwqyxgbEre4WUURPgwN
/6yvosSc8xBaO0ytqLf3iQJJARj0epl+8CslLHpwOoEXvOX8jqwIHXlzPBZ/w42EOjLNMh0iOFpM
0DemPHldaEGrWhwYH+33h48lN7+8Jcdysgro/g2wVQ8miV3ZuEQgAsJZqv6sYx3ujRKOQ6d5ytAn
mEkGaXnIMALluKtSlV4hni0KiD6ivQpwlJE0ZJZuFYk4f6EZUamwRgq0iDQpK/y38bar15tipjkb
Xmmwo7U1DUPBuHjH/XPGPhDhiDL0ZnumsIpuDLMqpGXp/5xuXNthLct8KqEuPLjveHknyGAaElTi
go+Z6wraNBYRZDIsTX2Z/FVZVjH7EqQ3eGxG9OFMHYizwBWNlfsl3/8K3Jj0DyqfE+AgHx4hKw8Q
r6pIpGLTxQlNf9UzQNZNu3BkpwLhgRI+MFyVsPdamiay2bpBWJEtLdPRzOST/de0Y5Gh7qZnDFmJ
UsFZL1qtL8+PbKbtOpuILXItpnSBlDUKV4hE0CIff4C/rDEI0NQNQ0NdqX8TEiOa82BcQIQ+Qnlp
m85mpmrKIUqVdpEiYAoYRNByz0y2jBK26yRuTCQ3hzcJcydXLVfT0L4hAzs/bxH3RuJkSpOrG4CO
jElj1c8J/xwH+f5/qCFXrjugQGC9KGv9/m+sa1f2la/Abe+r9X0gz50xWnvhcyA39niuHH6aD8Ge
waovQSrtniX22SJxzbgp8FW1lSnhMdUG3wSQ02UWTW2bqI2MxspRg52VeCGArFN3hG8hB5kXbydl
FOttFEh2GKQ8s0xnzogD9ZKn/BtJO8bMmR/osC/wTlAzs6tM/F0XuqYDeq+nUaKzZDyb6lDOUvbP
CYMQTcXLUwl+BAPMigVPz8pGxqSl5YWkWISRS+r45/Bp3okEft8+o6KPCqAIYdsxyqwxMtzcx+io
GmHR0J9HEK6htul5KQRtj4vZBCquDivPUIl3xhlUNERZ3hFmPgVt2r+6qm8S0vwPQQCAwTxCiu5a
0+H9WuvRcuqovimqFnYtWl6ctmItJ2GH9BYvWdiQeRHjXxrb8GgBlSWSWYo7cpf+KXg4W2etEZjY
hvHStoLRmt156E9+pnZFAwh8kfSLbeoOfh/aFicugoq3JVBiZl9Llt59kdOPNNHO9Kc8gL+kLMHg
dWPpbK8jywvHw/Csz1MEsgPlKKnZ/9W9YsYKPvonPZov5pmIrk2SuXJyXXHAA3cXYerW5lwlueOV
cm8fW7xsKL2WaltT1qVCMweMwUsBvw0KqVgxMFvGQdXH1AAFKGrZEMCnITP72DWs7lYjjIBmo9RN
B+Cql7hgg0QHE7CrrIQUw88fRkGYyCpf4xOkrsXQBsk5eOVlfL81lt5CMC6TpbKjHsabph9eF6rF
Kapr0O4MM+N3ex9hsnh995HU42lEIvd7fTMclef7RklhjGWMWoBVInDLtW2iuWkl/WN8Z9v/Tnek
wwL+CAIWJj6QptG+gac5nmKPbtAisssPdvtBxTF45bXYnvorc6VjqxveHCXZH0sqglgmXAS4r9Uu
fxHmnav1jZApNVPCsKXlZ/Qq8NpUjJBJXzPsog2fh+KljpGE9xDYkdf1Ea8wsjjdAi7UauzorJmc
UNrYqAKkN+Byg3ubK4SOuWF+n6nQ56KUx8c3u1KFAnCM4KGXOl4RakhWwecp4Ci1ek8997QKA1yY
4OniIMX7ZaHbFKxb/adO1qk3Rz50flCzfoYVZ1sg6kO4XnFw/kSCA2nXJ6+YTFW7EGrxqsHnDVSo
Pwq5BVjkKt49ozXe9tMdv4AJ7xNQaV+jANbwDAMp3RdHkoV/BBzksCw9hcira0bf77tpLsYZR+hY
CdS+zcEyQc0+T7+0uHZQ0QVLkFUBC48qxws4h3XkiIN+j1AWuYMKEvW4Sg/sgoRByodfURNbOFtr
mWyY+smLOLBBczjP4Cg9CxlWk+P2KTOvw+MSC7xx/rmT5jeZHDr7Q+/NiR9u/3IT3qWceQoOz74D
2554Zj1TpDLi44QfmuMZY6swTd9jssobrtu7GLk3bN0f6cjsFrLI71KbCTVCzRuE7+hLoaCTIz75
6diL974pyYAJmB61Kk65VPRf1ygSTDzoGPSCRmjNrC6TWLGMWqBtw580/DhHny7uWXyHYkB4lm1A
27nlllS9Fnj0OFwauqnnLZoSRuT/wve5Nx+PM3jZnHnVdIt4bK4+hbPc0nca/RPBWW3MFGmoAnFH
8Wb4KO9ftjoJxBCB8rplp0fmuYTBZhG2r9nGBTIL1JxXOpVABq8yRKDgohf3y/daTDUBwGyARdRt
KT6mcZf0fM9DY6pqlh9cHu4oTk5N3Cg9oDQ9E6sq0RoNRSYy4+PDWye44e02SJjet/xMZG/aRkOD
L+DOQ+fz9JHEyOww+kGM3ldNeQikHluJImn7t4E6GkstBs3sbb+fapdxsgZ96UNyyrJftwhYN8GH
RFv6LSTKJUH+5B4GqYBDa+jwLQejrydxCDiYUImtP9BFxV7L83SOcCD42uxr9lJXHktLIwTMJa27
fkf+g8osUIL4CFqAFB9psUlxEsF6LFzj/lSeBJh+s6ir6PxdEUkzjQv09o4RAdmZEAX6zbdPWzMw
1LhqLd0Ib8FKeYh/p9Go+rI8q3KFkTS0oAE9Pl2QB8k2tAENuS8qaqsJ6Pn8yyEYdMN24Jhj3UM6
N7AtjgnXY/OWmwiMBkEMNEB3Bi2iUW0ilOIVfDD0aelmzjAU1AbOEsAwwNx57zRA+vLpTNFIJUbo
zcythAvWmcSwhQZYDJVBuqvGDQRox94+Xg606XfEJS42vWXDVmrTlkVC0882AY5wJv85uPiZ5/qM
c2u+rugj9yAd4ZtpUkLnkjdQ9h7/cIP72PXGf/iZ6nLvKB/nG/87OqpzX2bPyYNZgmrptd40Ta0q
1vjx2EedyufThy3wo0o7AMgBT3TE/BvPnUmODDq+74EtGINKqa05hFZL97BaFQ+kAA5uC8v1dL1L
yIYJjxJVv0Ow2/hTvFeGxa6ucFPKCMnonxtTHILWade/AxH6gabgTjk9dQDiiGGc+LqOySEChSdP
yGEcFc6O28wzfyJmoVHmQF0Y4ZmKhYZnqhLZG3K07HN35h+au8eofKsjOEL/PPdnULG7/sjQGB5D
n1q8I5RfHxQ/aNiUbM4S3hanxegRvdgxPH22yuqKeCfmtC7kxEvGcIjyjkChQkvoYSkCy1rRgJH7
F9j5xpEPFMuiMTqMvTfRTPX9Drxq8AZ6M3maJ//h+DpZqELcGZFo+FivBQsHhAix1OPKLBdAiYKl
EqxtYf+K4ui83EL17srhpTy6nlWDtj8eWg6h/wmRj6oQXIzyPgPqujNJQxj1QU3DTbTxYpX+4vAf
RI2vO5MKJGkkFl0qoSoynvhvqCVXaVK1Pfq6al5gFdGTvUOMzy/uWTUY36DR6fsFO/fcnObOWrmA
LdiyigMb7QR3cDURfVhV58KtK2chI8hkGYCXpiHo8VGb20pWfY7PM2AAzEq9AzMOyPEEp9yTGRuJ
HAm8muxp92z4BXjk2CQhKu0KPz0Y/xq1WGZjXg6e7P2cp/u0N7+RM9P/GuezQZ8vREJQ0zJDyJ5O
64hOn27WTakzZmIfDFxjDcZx2HJsWTjmdrP2AY7khB0St3PtSJMU4qo40dHMrf1u1m6hi/1R3a1M
LQD75MwrFzaq5IDe2DiZ5FMOvXc3Ej9XdlWDpjlQrS5WmV5bWk6fULrSUOKv/bsEhs3tFEgfGE95
7ofRrVvulIiRKp8xYWnJlDSGoXfpo5ThOGDrr4xfMALV+buuyUUmMCUbXbPzfwyak3+L8Tuvmuc0
DojOPedjYxqEeEbJgaJbtw7rHyZCu/O6NuCaUpU3RYzcIPHLWFBfKVxu+nC5MU6OLNprLACoZXdN
263bunXsOvG7L/M3VIIja8W58sjXjUHYrEkRmM07e+fmmwokRQgaodRH6Cpu/TQcmLvIbm2CSpsL
mQUs3HrcKT6rwWR94V1Y9CkpHyRBe1q4601otj1kTOrUR51pk3btg5sGtZ+oMAbhMxIhEnzRzKwm
hjnNiUVDEVTz/QmkY9CamFbEQ8TSZxCtgWZ5c+BUt83bvZfYoByXDK9lhvgEvvNQPcqe1Mo4q/TF
JnVyFBKvDxCZYMGwe+VuUjhdKw3QsgX3H0h+F/cyfhnY8ZEYwFeqAaz3sv0wYkRLvKMdqZT6HqiR
PV5FmdyEpr5g+nCOg98DKcCkj9PZbDTLHV2i4cPHNrqUwzVVSc1hLaZb4kO4URPnF11JUFx5G9G3
ip+0dmqkfpsUyRzubkKbDf2ALDD2lRpmDs2G+jwpY1qmYRnAH06VePBnfbHe5MelZB6pW/camdud
sh0vBssWjZsiRl0PEaT0G/D3uNXG3Ql61kWMkYQNTORrVdnNRdpmwAMSCIPCO3ynkJX1ui+BMhPJ
gLa7EgUITc1Xfz1F5WoFyo9e6MnVpVLVGbxXCZ1WxxxJoUQxoLxE7lK5n+RfKqKIwH/4YHNaQAoF
r9J8uHnd/eLNwKfXTaV0VcBP/FeS8m9/tcUTwRz3vhWFg6ZbmUefFKsFh7FunoP8fGsbAGHVlkmZ
BLSTwr1HhFCsy6FqJqx/A7s272Imt6vLXJwDyAitaEeYMplXHd3Lj5zuoFqWe+pySYzdE+LsidBV
1y91yVYMfXhoeWVutOlrPA3NZ1WcGvKkKCTdDYSTBDd2GZWTNwHwWIdQpnAD3p6qt8qnx8twYqZF
udzf/7yCd3ff3Br5bJmStMtPpp3XR0YumSoWe2QRosBHRglAg7Q1J61ILM/OEXjBC+g8Qiw7EOuc
HmNkaeGJnqUBS/BF65K/0G2uHKGt25V79/glgHCM6uDCzdGa6ssOCmZNMr5BlvQE8xGxZJin+o4w
JDOgJdJMJnLp1Q8VEr7zVDUUjFv72QCeWTD/VGN1bxAQ9aR/hC1ztPzBHpVsLCgstoKYYAlx1eOQ
0MVJmrzS8JhQP2Fkd4IWEsQt0H4AV11A739wJZ3b5268y3+f2pU0WE/isBoVvbiI5Esid1uMVFGg
JkhRizKkOHRCMk7+a3Y+aCyKyvuyWWQFYcZ3pC04hi0de1TFA3ovTx5O2AMxBnQWzgmBEnPEs2yN
Fh3YEYRUDUr1UVrpWFMBFlQdFxNyKg2Hh7/fYF82nK0EfFSynquaBvHNBFMTv/uLDIfxdozt3Fct
Ji3UaEjrpqIvzg3J7yDPQY6jviZKfQx/7L/uzeQcNXlI65XZysP7Mfvp/0/oD0VzCwkohL68nnoI
Fuafd5MjobSzqDz6x2oDaXedV5/zAhKgX1yNzqhXMO5/agypALvqcUB1tsc9C+xDWZuaEe2SYPKX
nflV9IDCi8ZqibYNYbmEVIDu7tkEvsvcuAQr6RarNa0MS7iC1O1DFOWKcmbzNJ1u3Yepo01ie45p
yRCQzbw+D4360zCL8r1fHOFFVoTb4JDFaohIfmHV2jEuqL0hwsFpGl8WKQYa5KBuUfM9kWeMbVwR
MjJBrgMdFY9UPgyzQULiDILdtgUOqGPnplsPgUwM5wPCTAbzNW/ECbeG1VjUgiigA0ePZn+jxem2
7pNogqUwrncwp6kEDzKrMvfG88BYcx8qCGZxxZ23i3kPWhlZqFgJqA71EAsjOiFF7o/Aje0wiT7q
fj0IVMXESaD02/D0YqOgUqrumWAbNfFYQBB5fVLzmLrZA3c/iQOLhYSGwTkB56yc2wR4ctDWNL1u
7F6oPOCesg3xF4F+16q9AvAJP2LcYYbMW7Zq1ennXiITuNlIWwlFbpb7xih1Dm3zcA00FkoAlqG1
5uUcEXcVG9M5yqATx+I06+9YodGuIX7nIWUSDVTHF5zZ935JKIw+jgR64HZPjbAiHwvovnMPzVOr
d6yBkMfAGzuvtC9x1EQG2gvI6UMHRIP/bCwPvlUhzgLrYGT4fCVoOZqTzsDgK9OR2Z316zmMS7oY
B2raXaKELFZ6vRNpGHRS7HTjB3w3ZdwbXqPQVCpQjlTo+40yRp9OzLmLIYbEvLc3kOjWRVEN/l/p
fGS/KP1Uw76bMMqeOLxEalHiqyTvH31arkI/xvZoKmtzUpr7RTiEtv6Stz036QA5SX3/P9kAPXPO
x8GrmS/ThL6g6hIlvdbxOjKMB9oy19+lpSZl8U6zt/KDQ9u9A45NA6kfzK+MZ9DKjCEw/RgsfPIL
SGUFchM9Hwwto3rIb3QcIO2KhBkXI82No3P259zCioWYkRPzpX8XEg/Ul7nMDPItYm9mGUoWdnfM
rf5YVK+H7G42eKWM/JLcA37XfcNa3jd3spGI6oD+IgfKSmgeqWZte51N9GS4Rj5sf/3eJlvor8V4
n38NuvN2pmmMpiPJqcI3HzQDNTi5SePRM4aLMDbS2PMK0Pb9Q28ciD/iqa1ms+Pl0CieW/wudA+h
+P2ApEaa9uPkHHcu4ZJPC2vq+ZD4/skZsLMHCsT3fuxNpxZueDig8PjdIWKP+hV2BMUXMkkt/b2F
ps/8KQn6AzH+T7171MN8E9z8zgZ24xvMoloiHG7D/5PkrSJgoG3AfqMpB5YY9+DmoaqHtbv3TcIE
4J4q88dpAfhtxLPIn0+quvkEP4x8CSbwcLQbJGqeKG8J7sgB4WXtonSTnogsTtNEcPat6G6nHqKQ
2IjERvSr2bwwU93ybpHg7/DWxEbLXOwerJacMOHVI3xXOjqrAIaqv8BuDRjosjjB9/rdtriyTcW1
KdQgcm3uftEf7fcFqlMsmuMvC8DKuzN1XQz6m27cKEPevLuMm0xlmuzgTPL/Y9v9yDQbBgwsGELM
SzqZs0sjfLiKoFSC3IN/8xvotJqhmfFH/8Ng2QiuZmP27CNxjJymEG9BjY0XKQSm3HjF83LRymA+
GRc+U88gksFgVV4iqRRu7Kxa7yie4wM9pCetYQ936oqy6ARH6vZN/MejY/UnYqi4F/Zpvy9J2ZZw
leMOuC+4/FH2Y412uR/irtAEUrBrPPaYWKrxwEsBpJUCqr8SpRl+QPwMR1ZbeaY8wVgnfsqnvJhw
F1dz267hoE/liN5Ni0w8xNdgeRBWIIoLsUrunjYYvBKLvgSJuM5AxMwpjD3/d9CRRg08LPGjnhFH
oGMD0TIq+w1QqulvsLqYwbHzPGnoS67BT4aWJPIhA+92ZB5/mhlObrKgm03txHiVsv1TU6rWlKqD
vYxAdRdkLqFcFiF5/t9jqw+74G2MomhuJx5WHYY2L377/y6KqNPUO0IZqc1c6myNNQ4TOUTwvxJ3
i/yN4KzDbq7ZpBiui1+5dszw2z/xfipgLUS0lRxymvrVr8QJYO4dPm5Mq966ccA25w8mD4QC8mJm
Cwd2X+OZgHqlRO5ZMB1aBaXbA+BAj0AMUcjlstifqAoaHv+ttJDmN947QPyT42XdIveRLveidwpi
1ZegtgTWXnr3MLCu+zjkEuj5CcnpO2eM7aOHn7rrrMnKt3IhiV/TkTZ55xjbl9vP1XV0t2T5dCzL
2+5lAknliRmYTpH0x/0qSXVTJULN5jD6gWC2ICFkDPIdw10piM9GWpqTKZ6DBMBFYQh4KsiYi1zo
y326tKyBURahiOjKg4G+IFTMDUHEqfLALrLFACu7Ibc8h4alKsTXz1YolAEvhUR2TEnlbfkx/vQl
1LUmxAjF6Ci8f/z7qin8mxZraGhBMXjvGPk1ML9ZrhkFSgm6G1YlZJmIoNFiWKoZJ97QkPnP9AOM
xxm4WmNpyDYMXvhc7MGJi/GZw1FHJ0OTplMQTFQ6bxy74O5QGl12bpBrTTq/moB8kX9Rw7ovqAZy
R9yKSx01Cbo0HZEMilL4NSaV+mccjlBfIgPdb1og/WdDTCwHdFzztrUVFY5IqIKQoXXnzox2LOVG
FvXbrNS5DeB6er7HjZD+Ioy0+GLpWD/96PDm955SsN4EiitDi98T4UEkeQh/A1z2AOdutqyz1a0C
fSiSPUqjQVr/Om++DxSLh6g4JPMisIfSjatlDxVkeljkRYg4f9DpGaP3gKy9zs4MDHJr2b2h3eDp
fjhr1F6AXaM3CmYBfjDRdnyN5oD+lJcBMs8//ssesmAIhwKaMMkZTV/ahmwcWOfmslxmDVHJsJeG
j/wS6AhdOgq3CrwXMVoX/e5wWaJuyONzom1SWUZZyzHAg0DUxAcmnry3GKztlkEgt/pP70Gee5DH
dRq9+ga3/DyiJt/jOMSQANucPl6UsrVVDlaCTVFgrsTXbh/D0iDYgh6QfUPUy+EiPqOeMy36HEgc
Zuh213BhrpbH6CMVt0mmHLcZ0tXI5J6mw8qLEt/YQCljJyrIbXnxOY9PIo9+mw0LTmnXzWc7wTjp
vbe2yrAUImkDQWeRp5BtlCU84tqFlNRiS09hY6b7Y49qCquxXxAmznh3dXkKNk7nIhD5er89LzFQ
S4fOuRaS/s/LW///MtsUXxKpYuH4TYlvH1MXJoiHP3OmsH6FZhlfc0YCRlqTLNkPhQmdyOr4ojBm
Dh56e5lSh5GQyLjoiVMbzqS5Myl86aVi8GXCHF8YvjRm/GP64mvy/oAj0mkrzKetD3W5vS9iWVa0
zF9t9XOZ9rAk7tJiTX60w7aD6D1AImMJDOKooT/j01AQeVW+cRlT2x3AIj/rxmau4v9dqW70XgNe
ZN0W2mBXNU2cgQrsvMGu1hgu5k4x+u9ocwRU5W/5203+z608IXL/ZemQQ/nVmhH+9tctSEaODN7B
P4/IFj1kVjnHJSORKwo/SyAsaN3NE16AzMRS4X8ZUe3bH8PzgD5SepzCDbnTIh4nFvBnC1MwPt06
YGOUjfz8tNbbgt1Xjfh8kmqzx05bgllBBF5501qMJ8V+/q5h6L26Y3YNBKAik98bc40rd5y3HQEa
SToL5UEMyqaZ3ZNd77O68CPTbdaFkZPI1mYCnchoaleeHeK8gxD/BFWnyksF5ong2dSVvF7dgzvP
ow2fdqYKuhn/pAG/NWcTqtPSvPjY+e/Vo5Dwm+lfOe/UNw2+vXZuu4GJHfN+urbpFlHBpG5rIf6c
NtiYJCDHfPiyzE5H6X7kLtwQuwFVkrFJl/3yyn6cvjRvuhV2NlNdfrSO3xggA8M0IWLFjR5CMuh4
ygvREwdkF5WIpfPmvidM+i6mY01lxE5I9dtJU0IF65EGm6/6ZF5rzrmH9eJpcOVh1L2Bt3xQOf8Z
9kAKDXM5ErHl39a0GYBURD+CPwcz3OtYvpL//iOPG0XWmm9pKkAm/UMXA9tkdv0r2/FXLoL4SkSh
CBdSLHVJhptMLVKqK6g1nfw6KW6mASgPMcyYVk1/U5UPd7Dn2DRJHvMzIFvw7m+r7DJmgkB+tF4v
W89WUSAzV27qzGPdY1RGMqb6qjNNtVNmJ90Z3saKr/3Ls/5vNVvzRzG8RYrwBcroDpQliAxYTEx/
0zHXYig8kYrzLD45NmpEjwL7C3H/uFMQAXpiwbCbTzOKWcfnUn+AeSfGivFPkwSoGJKQy9DSfTlt
KrHWnynruq/jP6BfjAYexw37RKwBpNYBnxtkSesVc8MuT3oaagB9mwnlEFhWJAgz8y6n5kZY/N8t
XlvCIWM6AYXRGtAsjxcn1bePqUQifbDO8OhUs1VIBbu+ADLrWtvfCXQnEIr48a+6uMqcIzn+GHIh
Y7rzVviUguEy/5JgHli4mZWe6QNiI22xLKIpHrO9woq4c3Kn31R7E/cvNfDVI/95tll8NmfdpyFX
t06Y25HigXwXjsnfLlEQevEte9fRfDhL4E375bpboqsNs/ytNXY2u4/LnQ+TALzB19cj35yO0ihF
xYuSjMjkDs4DlIF+ELe/7Yc+QLAWCQSXL+wwoCYepew3DyxVbnul2RdOGJ3/oAwqXnPcUz2BJ9EG
GSovgzp2anjgQ24EQKMEqFHCnMhbeSUz8zA0nIe6aHPyp8KvjCYf/DgydOiUETimIOpTr/0QsbqB
m8rTdW5NodDMSLDCZlgmszNJWOVMFisFneRNb+UEF4NXgTpexJTeT+tLAKJGZ2DusG6KImZhUyr0
xUBgmxb06eED3YitSpNoztKQQV8AhUqz6DvkXYhV9S/lvQe9reNLux3qZ1tf8saicGTlqNrzEC2Y
9Rzw3oieyoGU5IpbRkF6sFEagOWksBlbPwD/xt1dQDI+9B+BJOLEz0FCqVg4XxgAvAOxsqbgqAzm
dYweW2TkcW6Jw2DrFWaT6MPWTIIrSnDWYIeqED4U5j9SLmFrPKzh5aWRzieCGO+MmpUcjHGHkHoR
RreTQg5MlAzDYSeBGwNGrrvtSE2BptLKeQ8qLfvqvCZRcLJiO/9kdoZMu3Qn1HGaIiS72rY6ZwTh
CRP7pB5PKGe3/l54F4LhaZdRt6n/9Tb12Lg6A2gmZXVAnbgR+kKllu5C0sGIO6yzD3ZS60NOsw4D
iPXHvwXRpxevrahlV3tA7g2bQNNWIYJ92VMPGPGvBo2i5yVf8V4+5U/OQwINMO9XAGf0yTbYVUez
XG3g+gK5A25NEP7aca81O/xWuH/z4yyLh0ESNqcpbl13DvLAZjGTDJLEj5fG4X+l/uMONKaf7rFi
sGMwedWjKjjz4pMR8Fj19L2AOrjb/vQUL+/GUthJ7IFWNnPYktrGOe8uHYSodcmWRECUFCNbx0ec
ldIx8kcpwD3EIYv+96QL7iy9QASJLd/SoTNvl+68l9fK2ftc8DBeftVbXUUhrWjIuLaxOSBzBaxt
lZJGOWFH8rpQE/5yxNMiYsPUoZJybDI99aUIZ9waLqcCaC5shNSwqOIl6JGLqU7xy4hUoPvkXK72
6lcT3qPsq1jqY0tmgXA+PPwgsVMErNw5qQ0fUEsUxkUplFO9eCAgtta37QkEpTouX4XT+SmzqJx5
8pssG6F0CqbiRUK01Xha8O4D7ZeYCjm1vub9g3WQsCQlLbuLmgLnPcKomuKRUGaDm073vCPDFyyM
prT/7uAKKBKf/osfTE/e3/s/wR9BevGDsDq1iUvT1vL5kHdXUZiVZluZlb0X30HqE7UDHlKZJ8gB
G0VQ72LXHuBUokHtNTE1+ORqSJt9SFimvHZvIhvbbcXnfuroQnTXL1YBrdurM3GynYaHEWN+02wh
HxA1UJjOaRTajx2PDNJGYIF7rWHgd/RZTivaJHmvNETmAwYLrOfmRR+5GZS54oSUTzl7klILordg
5FLkTrq4qomNrVRfG5yENcIWwLxRcqLxhIevAGxr0+mItFOLxKU/kBi+4dZ81ER16wjl6j35+e4M
/+kTIohniiG0oHBE1oddLOBLURpl3FUYlARvsYHM1J4URt4DYWJrD71y3hzUjxCutL4r8TpGGR1t
THKI0Ze7QfuuuiV7vojgTf2ah9jPRmPUT6CsQvXFM7sJ5awc/UEAFEHbSGtMyX01i9+fGd8v06KN
61z8NuCwHcdEBsLloAKrRYFJNqhggjVBn/+TAB7IhmfBaJGLdcBk49mC8/oUv1VEqIXh2MQzTcfr
LM4yEGFP5uw8KLe+VQ5anO8YUB438j5biZYNfrGAsjA+BLCVCUaTaSXxm6/lHXvr/Y5Nl+ntLgiS
qecjHYlQXXMvxgkUXUx2K5gjiPIvCLnsjGzyVCw+qn6N5MKChNA1X3GZT9I3+7mysDtn9woqiyML
m7BTqvN7m2fiJCxIfJc62Uu7kQiECaLN/ImbrsOviFn/5NFLEVFxDL/8DgnSynXMlYXKAWSvRGYZ
/gNoMOmmOZICSSrMf0z8GL+GidCkyzHAJGeIjTMgvs/QztAXLgOoIw7qzc34rKYAy4SNuYXqb44y
3DwGbalb825eo1UvwY9Hom66OVQxwmRbYX+ccnAEOTkwcT1N4NAQTlBIwC5RpLGi/VGQ1n+E6oZa
lPMe3WT8XxghcvzPDXhMtRGaI0LpdITf87URz7xgg/m4DbOTWLw8EINN+U/TGH8WJT7ADM0UlsGu
kncot/4eR1rCAYdz5lTjdbhIlRfLpKQ+eUX9az2XpLZCu7KPYZ4KUsJlKqawOkrqfaY0as50q+AW
qK7I/Gb3fKpqoMFlQXV/2uvL521ZAYj4jasV33PuMEubE3pKT9/dXpBIFbspC08vcuDrwyPaU9JC
MwlrqJuviz71zSIsE9TmIBtA43stbc1NuAiUgaEf0zoS/Ec8bCNRTJCNyE02xmUnW23o7RJ+elco
kTvKHhYCnpJuEyL0wOawfNTG4rlJFmqqUQrU+X3LDSoIIgP4OcVMoWjFjLVjK2DI0BgBOtRUjkbX
9oaz/JarZOW1Ug6phn2NT1OmMEa6fp3eYwLKTrOf+vR/kjwVvzuK7ClGw24ocOjNVRXQu6jSHkrd
F8LAYyCKDzEph6vfUJWFgilnljBW4RrOnceEmBnUw+m5QfCJzmBrVA2LvmN8UhQ01VtkWRrr+Kfl
TvelOEwT1IGMa+4gVrB+3ffpYfJ5vN3N0BYdkBLLpyvZQ+14MS4E1MR2yAGS8tiw2qXKtN/Im3Ou
H0KD9QEaefYmQGi9GxJ5SOwa/0CkgyzQGKSOMOleqIbXj7LXQS3gJukLDCXRZ9ZeuqfvQhHCfaTw
+T77FsQvJLYAaGEv9xaXVBn2QzpbdkUdObVIykkE1xHpKBFQ2LTFdztTbC9gXpxxRjiOBg3Sun8B
pTTCKqxZ/oM3j5mKZl8Cnr22Ji5ucc+228t+KO6Rlb/px9Ov++FtCgOWl2CaT3pJ0UmFu/wQqqtx
GpA4O4/Yg+4RbikRhqpTPZBW7GsOXgb5gUcyAUykJqB3jE+R+VWZbi0Uiuczq+4LlfJ97eDI4sRk
Gy6d2dt7YF4j5dmgfSGtFkpaCHm5h/MXhpJ6lCIwh9PDOXHO6yRyEgZhqUbyIrZjmdRUIxL+ObPD
v5YlabK8UyfbxmE62/Hcm+g8zMruSzOKH7a64+1DMh6Uhg7B9PEKu1bVaP6R7p7u8zQzMrOJpDuK
e6o8dCRHaWWiWeg4KqdyFfC2AA7fQUrrVkAuzlfoemVkqkQqarCOHZbi1t3k8RF1rbFNSPQKPPfG
i8KikqxYgFnCLThw33L2u2X/PPW6HKAwY9dWDHxoJF2dhbioEIh2nRcKdXGKMPp9jBnmEWprInSv
4Nm+Ua4VBJxGjtNahnss6U79CLe27qJNeIPomTZgSqh6PTCK+XBOV8BoOecLC9fDMSjHBIh8+5Wl
7RmLqF1J3G8B9oP1Tcq6BtUqgvu60rOHKByAt1R5VRiqi4pq7UTL7M074SVe+Vwaiesb1N6JVVT/
YAcf2vu/y3vWMk3EhDDLksvSQJZeuEVDP4PYhPr0ckwFIg5SXO23gf4SzPaDLfl6HiBTU6FTGUN6
NDeKDybAMO3b9QcjJcM21rsZSnRvFXlgPpvL7KjPKQ7XuZBWFZHEqdetRThIUEv4MshJGuE2EomG
AHpdYbz8pW3Rc37V9nRjK7NLPbxu9NAvDOmpXCl3bctuuLnOc57/BhNCjT/eI/o/wynDqKPsz4RP
TgDuBzoeGrO7wTwFfAspszhbk/cOCY+jrcOnqd/u4TC/f1CEdbdn3y32QPOIR0WO4GNQcTk6FkTS
llzJ5kl08ytOO8+dwZd11C/G/KE2zO9eL57qbTXEp1m9790dWquIlTQyMGEKVXjoHiQLziyEfUHH
8OsT92qBavo5LWlo3Atw1fPzWB96n6+SDfmFOBc2/ZgsIRVOXt/09kZ3pzTNYJwaCFdVs7EX//lX
NGnHlUyC2atyjL0m4f+flPvkn7paW1e3Hyb2GeMXkKewWaxEwFG2vx01OR3CV/OFLhaPe7kYktqb
uEPzaNGoiVzsxHaX/mvutSOFMvi13ynND3GjRI1VuGuMpbY6eoLJhmQjhC4Zat9JqKI68pYvd1sC
BSJ9aEkfL6/zR2m1AA0mv7elOLN1D4+69SJ62Yx7ngCl/uhhZy34AXxBKr/6rzdhTERpcpiU7TIi
v1zFKIXhMtMWU779DB8s11/GTeAeM3Ob854SbTeQTmEl/gs/HRg6MBqN1qupdp98G/gGcrZxbdQF
ibFeHH/Kjt0KtmKXl9gBzHYT6QN9rlxG6YulZXv9blu/euJ+emw+AX4+kZaod/lqLynaj5v6jZlh
uz4iCX3PIh9T7YzcMJr+vKPP50LiF+wxMq+Nm1MMs1anowAigVEX5RgSYrFlqge8/pnt9P5g5Xb1
sxc9H9/W6uX8r9eiQGvRSmyVlOKeBfsgEqCllisbAo1ye19SX98FXl+VtGtxwLkaX9dUXDOcu10X
8N8TH5EGNUQMVgzt+Xb6j4yr3Up0P71zHvlJUii8vypuTrxNs8iA9Ywb93Is34d03r0oI2EwcuCN
l7yc8T+pWT8DqZAAkE9XJlzTuZZ11H5Sm0NTp1UHxBxsQtr5tcGqo3Z2fWtL3O4cKPFNZfy19iEb
Ho6MK4Il912LpnBGIbPn4vo/Un2i4vGMNaU1Tyll5gtC8g4XK6I8K32W6+rHMXjSj0W7yCY8pVhD
vJ0TCAJ0TwCiKgGF/jGacvdWXrOi54kiI85uNhFtFr6vUyvU/i4WSmqn6V6Be7Jp2yQCVZeNfWl+
G0T2HQBB4egjedmuWzWIsFJF0knnVKrh6HEOJHi6AkkZLYESpbYIMpX66+ylgwECifU9FsLkNF7n
v8GXgSGoj0Kc3TWKFc9p7bsBACLJp3zXYa2f+qc5OAR4d6oWMDBRnUHUNJOG3SdDkGhwsaJbiBfc
qAqhFsZeeL6DVO3S5e44hL/QPtgvOz9JAiQvhQ8KQl/VEORSIHWcJpBewDcZThmP6wECS6cmjKnh
Z2TpXyW8LZu7VAjwRMohyga/s1st8zcHffGs1v7B8bKEhIf8SybjVWXTk4jgGTkTm7ORkvXRBWKA
rJJlL6Fzfyk+ux6tpzazrSroDOfxQN2RqomdrIB2qo5RCFoZYdVwbtNxrsLyWMfD8lK/LhW7lnoq
sQbEOrrb+mnVMPV5vWacwwdbG3CYwMMp34gL0Hl8SQKBDfy4ghAkjG7TidarKD3xUIOPfb9/EkJq
dK+Q+ZNh0dzypLmGtEsPKpX+bDLOzXIV6MNo+aGTM9I6id7JrmpNT953N5rEHLMCTXhwxJ8eFzCe
E+xWHrwvCA+LINdN8uDlFLt0z8umn0QoIQJ9J5jDYPVW9oNe21qyICfDYxsicFUeCVIHgD4iqSRJ
Aut4PbNSaTOe3FArZhjc5jTE8+FaSqpVAzQyrvUWvvdfaH6rXddg+xAqlvAVRKzd+cm8scI9KFJ/
5/ASrhAHAyXEeeEj3fgo/MzWsmXRkNJIoOqGiYl5W+cAVQzomKMbVkrU33zS09QJ6FiD1tEfLbWc
q7V+YgstNLEreK1Tb4XeNYfdjVf2KeG91CjFeKXLKybTPBsC2L3/BFrCkNb04etjNp+l8OjROJf9
ASIEnaRS+xriKnwQZBwhrBqW+lcqRD5OoAWoJMuTbdbIB5bPA1YwOfR1kaKhkRYFeuW4g0Aagfwv
SOoRZXnzxYwz/fb0FBQ0IoxNRPFKD+esnG67nHjWJsxB/rv5M+fCfxl0smnNmdIdIGeUwVr4LS2g
tFkN3pOb4wcLU05eIDyOQeDWcR0KCSSS+NGzSGlYvM+tKpUkbJ+4SmMHzkjWWXHQIuEg3LlvStHL
BkZKpFunLj3wfDHbaH1P83nKn/OjvKpPiHwGWwyGKFgE/0gjf1tgq24hQ2fVdtTDE0LjANAcl84X
R2FoToIjsXYVJQqGEQeGqSFMUs0mxvwbTfla94uHMQKJoAbaNTjg7nf6QjoA9Rwd2ilPc6ByumMX
nrnZ/xNfvEpWyFCh7zyw6Cs7kWMBh6apJh6XmeWLT924aw1xQwFYKM0Xkp91J4L65zS21JRDsE2R
CPtszJJxd5Z0oVZEVSUCsNt0K+H0BZjk0o56l/A85UzYHpmct1JQ7Au8JHjloKkmfvSRPFw8M11g
EgrjJ0lMOHpvj35dyco8tqGPHbqPzo1npFrr+hb7W0JWBKcvOn92IryFB3330kKkGvB5hPYs4emj
7345Em9QnamzpRGgpPNe4ReuMUrEN3iep9b/2m56HCHEddcCVsDj57AAtm4l1Sh+QkpmPqWHthR1
gckF6/fVIZgPW2iUwXbiNmAMJ3byUsWYGuQmdgkdTXmsYsjdRsSUd5e5z+tMCQuba1MHQ6UY3MF5
ugIHUepdSeEy5ywBJtSSmDXLy8xcu64fz4EtPOTGpj9TKrhSHgf/AQQMOfwrCTa9mO0ndcgFk5ne
sPvwFeWHG1Qs1Z+SUtYD0eR75SVsSmn9ZgO6aH8QsWzOnhs8jBMXcWO/O0udd0uJ/q3lu8kdj41C
KMRXTZBFnZ/G3whqUbkhmfhhmzsJ45H/be4Hf0lTyk3Bn9DnucEfr8BkOZd31xQLM2DAjnQWi0C1
YbHmEqyFJMubE/eqw3ir5jKXOPW/sqdmMlCaQyybkwy6+xQZGHB5XgMq93AlFLa3jJsm/L7eydbZ
sPtmmaY5kaN856WKOtOhOE5OQyT5OO6peiSUrD0EjMV9IZS8cx8pjI3w5U37l7jm/wGWKSZ5LAPL
RqyBXL04TcDzjqrN8CQvSmg9Z9ftRpL7M+14ezsh1LoHjMJGq8PpM6np8Z3f+U0OrRPZnQNZ2R6R
7cWaGC37gBB7euPRS5NopuvZ87R1iQTGXEuXXfMBqEP1l2EVzUyDruiKjJo6deyosgROsK4XYo3q
4ujcd1dc1+VGZexSeBPSIsMqeBrmRLZas0DlUDYY8T6WoMG9qBKKNW/8+9TQQv85wHWIJiUbK/47
tlOmLVODPZASkbiQPMMV3YmKiTAyds2yTbhR3olaC2H74W+opb3+EuDp71/HnJ1URqZrpfIxvVL6
HMIJ0QNiMyuPPJRCSSX7xR2c8nbSMJCflozLZ0ySO8eHkVsjU7//ckDvoBpkWwq9LXbeHxvMSaS3
pJSQF5LWEdoX7sNPXpVxx0v3/R4lCUT8qqwZXa5ZfONp65EQoYWtFeGpBgKKiDpd2xDKPDRs6SUe
AFVA0miTvYX9jSz6KPFwvmw18mGQp/EsdLA47mWyUFVpEpk19JbzXtB/fWh9p+JcW0jqZtPAWQ9U
8BLBwKnWkzgVmsHXG/ZWcoWDY8AoEb+Becg3TXX2UlnW9rEyG1FYIRTNOlcQBK4556wBGF+mXDlP
a/PQYgr9bBgP0IoVsS9dJsK35mUBy/XAINSaeQw3yMWRB8WCxG4tCno4H67s+vABpnyi+oJkhnKw
TTWwh+WY5mqmcYb7CfWR5kw7im/n/fHNwUxFh4XqlMZHdfgKuoJuQ05y9OdCL8zdJfu3nTQwmOI3
jlXbqP8E7l0Y2YOxfsNYh1WygHNeYOVKZHykc9BmwET27tK5oJrslWBuQkhgVb/KkPEkiEbJak57
hCYov1Lr0Z65X3JmIZbbJsR+ZxQ5SVaACWxjhe5qI/MxLwQAIKxyPlbEUTNM3ZXqU2yju1zmdXhj
sRTBdXbHy5oIp/jklWksCoAvFhxqp48NBYbj/HMqdelB06wYkWrx69aF6qw2DEfdCo0E8h+boJuN
v9+66VH1lgGaQvOabkIwasnjmfzltawdx/LtE+kCwF7J1HJO2oT67CiVVQ+IIoszm7Stoid4gRZ5
1ZjUuohwInkiRFhy6sEAK/+vlWC6h8ZAWQ1BK+R3e3ehNIBsWZ5jCXc9POOn9nQXH3JJi+y7K/+Y
YIbxzsUcZIgziOvxwYHcPzOdmFP3eW0cFFJSOEZDfB0UJ9O4mkxnWv/nsz3gjta2c3txZZdW+kRD
jvnpeicnIf4mqstgPDy+GxsVq/h0pukeca6X2oAnno0YhIDKtUGuBEhv5/qdYn0QZ9u/2xv5rcOy
uC0+Vg7mqXBYH9Rdv4pUTPfmIYr119Q10ySeT7HySgTpF66hsWblOL3XyJpkMAfpy+Ozo6POAiwC
ELMSaboIJiS0QI/0HKTOOuupAeTRnjRsaKh6pCBBzum+1LRLMsvU0LRmNCFYmTlIt2p7JMHdKCIv
/8PHSTPbtnCinIX0J0vubcBSksSf8yjZUJBgwZaDrDqR50gIL9NceG7StV2eAHfHd3WjECRH+FS5
AbKKoTzIMZB3ak7NINhjnum9cIGSPv96OjEWdnTRzxKeYV1OUq6rnNDxs6Itsi1O27oAwstpNnkc
HObWFTKHGZDRqldmfi9O0QFCZEFlXMnf2TQ/JMSjmU3HK9dzS//l3lp/XbHJ9FUiFKpHteDU6tV7
noyYTJyJB1zHqosrQe+WHCwzR6uRdX/P2rfYNZtKUa99kZRlTmBprlsY2Lo2Gyru/LHm41lXM8+Y
xMIvwF0R1Y50YEcDKqNStcLPhrTfUE/xIN4f1vW2x2CqXTfE0uc7/A4NR36twazyGGJbDXEKl7Ec
kZ8Rqc3PZ7tSvYN9W5X0NtKu8A+4HaRPfD8NiY5zCzPumkgo5Asi+IeEbvke9xLEHZbtLL/9v5yO
dZOBLh0/sPdDYQktOPmOEVVcV6d+6OrRQQ/7bzeebdqYQ2EGZtuLbYshvzww6ZvvUKV4o1tlb4/D
iqRH5a75+kKG8IRIhCm90JH+8r0h0VYCF/TWp4y0BFuSbZvYxFgrQWqCDY+y/ygRu+zvFADVJbH+
Kw2/cIUwE2c0D5rxxIVNLFDCGEzERErMP08E0aOId23jXO+4G64N4Dz7xS7J+ylW6EE7UT7LNNsb
OEuFlV650r6DEiNEdttE7zUMZn7TN6iwmRyY5P/gxwdpDEwmatXBr7BkXNcxzbDXjgm5xLO5RpkY
zrW9Mo0QwFDGC5XlEYOsoQFsyfpOEHhjUdiOH/LDr7z2j9KujZ+5GyyU+wY9fvH/CItR22TC828q
22+OZFOduddcQpx07L8Ob9gRjey4y7v/kngQY6CbvX5lYTIobelMDzTRhNMThMh51ZuUD8N6uEcN
IgQUqlvyo+iWk16a/ha2ixBW9ZhiDm/8rGycEEg3yZyy/K7qrIdJIMWOVO5sUSo2RYB1bcs0484x
sCC1owyO8ipDVPXf2mZWe/gGz4To3Pqwxhic9DoZWcduoK9kqZkCFxZPX4mJDHM4ailJRhUecFuq
tnFOGtpcWneojU4ZWLq6ttkHgGf7tKCDpBJ87URC8GdxS04lAtVE/nfHJ8Ri1jhtWGjFG+8IM0Hj
1mUOSBMkqZJ1T3s16n71nWvkevbZJ8s4l4qyYzmO6IG/QRWhVdOxqeFSuDRe3IdrKbSJcs8no4KL
XbOYEbQ+U6XuBO+6pMVbalGQjio0I2JA+X2jKHIu5MfKgrHWg05q1oPr2wU6fmSR4R5lxiN65t4b
GaqlOs2C+yt2AZNEKdwSDnylKoSgFZarFbKg4Uw0zlOYKwvdlJYzp3V1gy9exwGSvD47k6NI9zlm
XTqxJ1XIHdBN378X/s3CI+AG+ckfGv1luSAYlf1Uj16khpFbZ12UgpoHd5pCnzCrN7uRxj78qrjQ
sG10TxBkeH4PxsJPSiqclMNKNiEbrKq9cAMwb4cnTPglQTfVVrD9bwIBdQJj7reyj2qKLze+6QRM
7wOWYI1gfp8VtOjvmDffomU/9Kt6gwM8PRRXr0BL/bLSCdCzrpAVdEOm8yHrKwd2XctHBpq54eWM
OKMvaiU8Bv+uYarQnpBMpI7Gb6Yv57yJlnW5BWp8E/zjLixd8j9kxu3tHyCXJ5RYVSlXp2X4ej29
HXGruxwsajEoXJtYdb4cTGL84Z/MBdsCBYJvc1eb2l51WMltZcj9Vl6Y+fVfYCf2jISZMhp1+gHp
4nnb0zqaeJat0wMHD/h8qkqR0RrmoUEb6FQViG+/6WLJq3Lewc++sOFH9NS7KYVnH8QIwKZMcTlk
t9+Lb+yExvy7OBKLNP+C2J3Wg7BGnlzPU2yQmIo39/Ytn6wdmvt+ySLKB8j5gauJKT8vaOdEwemu
yE+5JnrsNmvLMS94iho9UVKu4iZddId2VnQXLdU1C+rSLJE+mSrdAjM0OBX0DB/Rzq8WJepGAwBI
XZET97jgCsdLhF00MOP9VAPskmZ4yazzj2FqKOI42mbXMHKXjdQqkm2A5sAqq69SbwEFPIzn09+K
wvG1ZwtIDInvsSVE+FBWmmI0GGzEphnNOr16hoE8CFH9wURNf5DTE47k4vUKuluOvqWPmn3EUwLu
PlB4uNcHf1iiG80HCCxX7c8+KifwFh/wtK6jdakDvO2sHLN81MA+/+MSt1b4jhBgJPNViEk1SW7A
cD5tYy9R3rxK8ly/FPoKK3ZiWAdjup0OGadfySbUxtD7GP5NK/4AWBb3RRjfbKahaT1l2EttBZWR
OREe0CNiy9achjRfgnilr3dUrfGCYuzm/bFx4wUyrCTbxRBghq5GhchQdAG11CLZC+HTMawDdOwp
0uduVNxyBJYLI8rXT65eotIfZ4Z4pO9d914bDtFPKjzMXtJ5SuhFPk8qNcd5sYCZNuyo30SRoSAG
D6g5X6LvBf8PbogVkCEIW66bI880B+peJsowiJb44rw+s+nXEvDyyrqM+c03bM4YgtdOAWOO2Orm
6e2ZPj52WJkxqFhoqdmk0+GWDp1fN0KJnWjtYAI4LVJ7UD75CPrBK/68pzGXnDmOiP45Lo0BZNDa
hsPSZ9fDlYTaIEiMouYsrvt8NdJNBux8PhhYqnHSanwOjpZ7Jx635V1JDR6aVEQpxHulDjfB028B
Wu/3ntsYtV4lt5YZ6ZGra8NdeAp0/I31qHC6NVPn7TZlxlMYJRi3/88ASPC/WhryWd0ayXV7OAl0
EaGc9FLzZbizKcnY1rnZuPkwQexqdDTU4OTHK6L9YFUdYaZVVFo2ItH+cbtfXLk/e/ng/eg31T2r
27HWazrTggWDcgKF6g7lesxG/144WMcMgvRB0zEEgaJ7kpG1hG/o4TNHSQ0maoHSY4mJJSubwnXY
22K3ZXSoZGYaKRsQpGpaqrdkA7FDWk1x/n6W1Zxy2eKsGCuxEQTns4Fd7bhmmUlStAdw3IPX6PJu
f0sshD16PSlRx/0VFOXz5OFLx7u409gVP0IDLUWrs290YHI4RXXkN290TE+UCWwAfRh/onmPOaOT
VvgmFz96et3oL83Ox73fT3AIO5958bwvQ2FVxWicrm5aKAaciNqGTaNem9Bq8oEk0oKAnGqlMGrS
ggEt5hYji1uylmS0Ln01LQsNSmgvxiZu+UJk3fJZCL+B8Uk7ZfeRGGDolYgqx9RQJaVII0/ZkzIM
DjBPkinUByQqAVE1UV8jIGrqNf1gxTw2kLLYMk1l0g+BSOgfLmmNX3rKgkrbyo/MY0LfFnNNlmoY
re2ZcNa5hGRDiwLVrVX2WQjADvcxvHLmMLRlB0WlEshYOk7708i3X90sYz0N4QnRk5Xx/hWx9zSL
ti5JvJ+jLV++CVWV/EMvys6C4jqgxIKL5peJ5Wpra5TR5sTD+gBWz1fx+T2TKL7d5dhuWvoxcyue
yUQT6Z9jrNZjQ+p3H4uNsIFD4s98a3sGzr/nEPDgcFGjh2MuZFt0yMrCussBmznwPqmoHPGTCuag
uHtGoqVN6aBnRfrUizVnt9Mvs3s3kyIHoT5x+8Mj2lMAo4wbmZutsajuZ+us1+WxlfeqYPxMTqaJ
eP7b9yhCywUn0uJXzh/9/GC3ELjeWU+hjkiN5k0jlSy+YaB/VYjnKoT+KiSfs7pIMJYrocobG7jX
7uxQ3xTO6aNBh4FpC0pxHu4tUIhD7Z4SjaZeNf/X1rjCCxM588jpxRLFaFINClOHrPxYUvy9bw/8
wsfSXIGwnM748IgDVo6dNP+4cfGWE9VQDfGx8ic6JcRtqBwYzNcNtwVmoNpj8yYyCKDstX37jgd6
DCdglyyZFyRe5ABABnyGCpyfxRFrsGkcJWDvoP1PnZjZy8J5mQIsFletnhI8j1lVuBxXZq2ZAu13
gDmImm1DJMOYBlKp2TX5upGmurrcscCorl82oJ4XIjX+AFOaDLDl9m8VeXXb8hTjLILJoPrmKhno
yr/+6bH11uq4Q15oAN4eOgKDShZTyPiQ52TC39gZermoHY/2ixq8+lrQFys40eb7z9/Mao3JRVlL
lPCrO2TylWLO6RI3/OruA9t4gu5F6tVpOin56pvQyJiKrg7/H2Insp0kP5PLji6MIeId0Pn+UL9X
lDQF6s2/Ek1EphRtk5+2Z9x8+EIzerA8hre5S25k61ZT9aLbSoYo34B7oko9nojKYfkXaCzWeGp3
uJF3tjmt1P/Zn1Vpos8yQ1qDMPjCkkP4RTJvTMwl4RczJ0rEV15lP1SeLd8wdrU/vd7ZZvMPpbeA
HKUGmkLRgihv3UYu1ZbtsvCX9iHxtiWmqHXo/lzITF2x3v3RsmWazcu10CDx19c0atpyuj3HvKTy
0u64sl4RKh/beNrtrSIFRQk1pYk9NUCJnh+u3q90Mv+6hk5nDy7zRmfVGW7UiYuguwY0Tb5K2Gu1
cSKgMLTA5ObwU4hJ+s4xlBU3zCEkjVB85utKG3uZrApLTCTSpYs7m0I9FaCQRQMdZmfhzk+SofHp
EjfRDyIHHs5uCc1plhJmttvAcl32hzDAR4WGNlrrcbMB2FOXc7qTu8jCR/11dwQiZ9Z/FqvuKXv1
3Q79pzArErp5+IplM9SBAGDIWwv/Kln2X6ByML3OgDNkDxdoy/QAuwbwtDRkSzsTLatkxlFNw1pU
NLbYaSWPq05fxSVUYA6sfd9swbKA+50MjmD4GD7sBJAep/9defkqXaffs1HyOYnmu/wGe71Tms1y
KOxdWwISEHGwzrwaddhYyrclZDUBqLFvpxH8Esyp3zNqSqsHJS6GdC8obdLDiUcMmrwgxO8CWf8v
CJe0TWvg8n63Wd1zUSe+LKYv3Kfj9x0CX7m7j8Lfj97pxy2i2Eu7C3682bppy4aVzYWuaq9ZnOD9
jcpoZ0Y8Hm95JYLPU+UDrwq4eV3nGq/ua5zwJ2U3/PkCZCt4RoP/IWjICnYhiZuD/I2o0QbU7QSz
4/cNfgqwYQOFqk07IEr0ax1OxLUFLO/8XOPUu5/Is51RzstlM9nETqC7X9XHHStUj5bBEUviVL+T
2P4l9MI8zlBU+C4vGuHt+L5jdZ4D/D+h5o+SIuzHmKE42j4GOjWIAQw8XCSZOKdQ8a/dpBlW2VOF
EzvZov8oyhEaGDWOkGCGmfVdwq56L2u3I12W5/c/LNJ/YxxKEmXXkOVbr1H8cSInhtK4BWCpb18C
ljyKRD3NkYT5tiMwIZBzUjXXScJvXvIAEL5ONGyS9GO0kZOdim7HDxenuRfo6D81phYAmk/5K1k4
7e6Ep4g2a33lBJuiJlaVI9wzA69CJv4vQjSwF6qAaOLLV5ZjEyWUyre2ACly3waCRsFkKCEcSlVK
XhJZxDquowj9mPBz7hwo/puUr4lgjpRUtaafn03Zqkv+1aqfW4YuSz9+6uBNdzmbM7SkxqzWWadd
6AqsXq60srnTe/m84+qRWMctt3We1aZ5qxO6yqeyA3Di77M2SfC0uMsGCYuPTv+ubQxDUHBPUTbr
MmmxGFy6IP6m83RVHE8moMklqeNE95xyOzYbmSO8cIOaug6FYhljziS/PGB/p5zrSgmlfdEHjegk
EKFDsKLfsZiPFJ0S19to3D01c5YAqX65Wz/OitpKVnFK+qUHJiFaHM4uhibUsIFmjF6I2W/yrNAG
3/dLlAe4lP5skYjorfboIczX5HscdD4hm2rSDNqCGhZHT3exTD2cba94V7yG+I4F9uOwZMOwkcUU
cLDp2n1ba93UXby9Evwp36+rY39rKkcKxRMySIw/CRLWfP5atKq8MiGVsYefS2ok9UPQ+r37zpbc
k2cDE1gQeMr2QgWi4pK6bhkGvnxlY8bN0bHMjsVfStJ9lpJrwepephFgXLW1uR7NbDV6wHG4FBYi
VObZYHkUHc884u7zmvK9g5Rc6pUDn9KCqvmYHSXdwgcECR22wBPqwxVzN3T+wbYG/+tjvUQ1aTuS
c6qVHyv5SBOwiFiyx57Bp/hV41CERZJWHt5gwjgxGxd3LhTHj6+p4JPvHFSZ+ZTXKUzm5cEAaR1Y
Yjv/PsMgobY/pb7xJ7QwswuSz11mw1VMz5sO5Rt4qcatw4iCv14Q+6YU52c5ocyLiWHkkHC12ipw
+nBnupqVrKy5N2MVPvlRbRrFwQeDgwTNMLLbxvsyAGhSSYNlpKPdi8IwTV3LpmIXCMRHgRJJtE2J
ZL6trz4mCsQ+uE/rHPO78EMjszIwylFzU1DNmgZq1GLuyC9W0lHs3NqfaHvFws3kkZ7Tnlr0YH5+
p134pCCVQYrvPBeAeem5DfbCUdrwaC8kSy+NPCFCcFbEo0t/1GiR7WCn38dRxeh+0zaISOT4tnlG
1MsKOMFc4EucLqc1YrubiugH4DqOtW00cjLmWyW+bhAmQqI45gOF2LnXTqRQPUICKCojM7xKCMKV
+HpJtTamvpuIK28fg1JFQXJELgfq87P/uKZmsOhTzIQJKFCik/nqdAZT6+UMT6T87R1Oo5G5/gxH
+NMo6uml5CVC0XhU2HYGVMP4B39pZTICcnAhdlraRrqM9ufNP/kJexG+XgEhsNh8JoHoJJ8vxLQZ
Fr3F2Z0lARSeGyb58YIqBrgm2wpPTQmEMXKUEV9LulM+yEp3ixkQXLDlZGACInWG1eRm1vQ6hJcm
RVy8BTn3FGrYr1nnF7Ljy5jzgYLMXru2oY4a4wK7bh6klvFEChx4cY5F1JaVzJIk0wf4aiuj9+mG
Q1sDlVs+WxOCA6dkABTvn/NPcpFcdqCx9VK/LURM7+tUNmiN9XbTDWDtIindk/Vdp282xdByP5X0
D5AiDD7UuNVPtJPOV4qkmjuO8DnJmGkjEr1Yraf6Zb1gWMU4KovDLAdEq6MpfWYXHteLDf2PCIRl
T0ZKaOkMWPqvDmYzfDFyy3B7OsOrathGH6W3nD7M4wmPdyGWR5FdXX3giS1bLrASMk4vc9+fdW8G
VsxRXbcOV1q8RCBMFK3J0uxE5+2IHfKkqeqrKrHKJBWA8s5lLVFVss2uipuFbK9ku6L+VLQsiQtf
bR9KhY2dSB+8DJ8r1WEiTVp2mrfL0bRzqk6S1iJxhyH9U/r++wbqHQQV0Gz+77DM4EuyFFjKhfrd
QsbrGKepZGIh2+t4aFk5s4CmgWO7i/w/3qAWyq5c7103a5CtOQkRzcIc+QIIesi0uAeL0GMNgzgA
Q1CmZxalys1N7isxHiab07N7wknkeL/twrhT0C8XgxgWHbahg+NpEBFINNU+xTOsJgqYgM7jdasm
YvSjN8DSfzEzBF8XG6LfNB13hVpDf/0kqeZf4FQqdr5ZF/RyZezjbZjiTkF2w+c9xFlnDlzeWD3D
WTzmnonq+UQR4+U4wOLv1Ym3/oNpTJ0eJWUBahk2AOUcbgSP2jrM9vyy/56fZ7noqHSqtgxRYyoJ
uOEvVRf7wYO/0tWt7bMHhe15er+rf2/aqm8ttErK/vFPxepY2CZMpO0hs04KFxMpXFUR4T+2s5QQ
4nIzy1pjgbJMKC7vS9U2wtESpl3DsyLnlcOucxQkZNc69ApGpAsKioGkwol8Jj0qpR4C20Y+32Ki
7sEcW2WUXND0/eVkZumzo9C67feVBXRdiwd8MciHDz9jCf7Q1vqIEak2NsL5ElyHBQvJeLBmWxDC
5pKmyPTK2rPDWLUYyUImULgCoMdHv8/w2eZB3gKTrxVORMq0Y6AWOBrOt7vdug51SorXcOwoFdsK
gF2lsKhZXQ2QQrnb0gJpm5Y6G/9ppi65arzoln0MLKmElhY80CKeo3lkR7QrTlYXHdp59JgNmWEb
OYbTHlYxPvSRweqlQJwd0wLW7yCNPLbPu+xcvRNoYe5EYyHef4ZUsBKPMVm5sOfre6hxasiAb2OJ
NgomUm60nm6ECeoUP4+404sdE74THOMB+kUpe9HePq/gNPA55jM6Qrme2v0Mp+VbtfOec7W7fFOT
GIbnt7+89LxPZO39Z2BL+C/Do9noOWfyb0Eh6S10u+JzUTWkIQ0KpLF6LQtO81QPMgQculMOju7G
JXF5suPpyjl8Yg9zyD+hIarW+YGJwNoCWYXs9o1u3+HUIMBgkXbi0SD/I4vhZs6nrmJ2cTFEOx59
PnsF+MqDm3XCSgyt6LiE4jDpPwp503IOe+b7D+DojSo6OPb7ocqyia2uUVW+g9WPL52u6jPW4nJr
eHr3uZ3SvjiGPw0flxdal0rFjDLMTynC57egJ++nMdltm0Tx0AG01n6gfeaBSS2fpGT31D/eLjUl
ogxl2K8oOfKnt4TZlRChDypP7tg2HDK3YEPOIhQKD1o2Vcb8VVzln1KcdnHqfCdnPmN+GkBDVnou
S4CVoo1T5FEHWpDwxEh22qA+gXLu/4Z3QUP/brRZu38TWxUiPFnhtV6r9c7FIgoNHQMA1Gc8ZbiE
gQv4/kDfD2XWr0uk7Rt7y2+sFJ9uyI14Q+vaKmIBRu+/b7WQ7ajXzgwKl8V8MqIEVGrCH0WRHzLH
vGgMaRHdeZoPH3HnJQCvjarOFCiSjafY43+eNfCgprUzfP+AoHnYoqqhbi4Q/cAlcqmGUAY5NUd8
HOePgcnREIyQUYDuNODqNEdG+VvGWOo4wadPtNQDBZ7CVNPuX2Ax+rdBLku0/N3fX25wM2sR37A+
d4s7slDWekr1dyiSc+xA9yPmfBlQYINfMB617mMCdteLxJsRK1jAoIOouStuwC36y3CVhm4cx/Hh
iCN4TqPfei08m39AvUJpxtJ2dgPa3fG7ctgXK1087K4fdjE8F5PQhtMxgrT0h47KT1LyQBbwSzCP
1Fs4kFwLHqxZ2bz34Zb6Wwh1SwoKwJk3bl6zA6UQxEjp9GBWUi/ZwNLdsVBDyH7YmEvf7Cb98h77
P+LXOYqxcMhd8J58kxPkp7qosk2bFTbd+f/PQy+KlYxOUr4PiiEMM8AUUGIw0542CpdLbxzGGfy0
PmK22iphTtlqNLdEg5+8ipsqTqP49XkyXS3fhz/F3OX597UGzBKnGZ8ccuObE4mf8vv87npiOyy4
FflgnWPHa52Pvbm96APb0zFoP/bRv/NlFohRneBXQmpStJreamVi3pWwLv6r4MxE3QYv+/T8n9Jg
FxjTummfLaUGPkkuoNER0cd79KkZAuBrq1IwJf+Aig2CD+FA5VKpJsGS55r/V5uPKuNG7HQomxxy
LTod8pp5oUQcCpIolzrHB2UhpJd/3gfsLoEv7V1zCSeNiJxDfMEsOcwG8Oc4T4JSkoSHLcTe1pG5
RBTOV/5LH/YukLXTSSdT2W6sda7vR+vtylSBnNgKet/U0DSumUrq6I/yqtzyD2gUffCNfbXe9gZR
kPFAzYBGrwdy9O1VjXy7fNn46MvoT2X0lo3kGwJ0LQZNO1ht4Ks+m8TJnCy350TpbudRMxlVrb4F
7K/BhC1nFLMFMl1LeuJ6a7R2hnrFcO52qlXFicprZCOcbPFZ7IDDeqxX1atEg97VAM6Ozyxrypds
GwZWSuWzVktRv3XEb/2pLZMuXqAXI8hcPt05mgTo6B+PYp+xyUEj5jj5YprVHbMCeIWTIvc4v+un
nQKBRo1NxqmFbQFJMdrgi1HbKV4wHR0qA/Tt64WjAk2ddj2gZh30YTKgiE+Pzx2UvtkgFKyRoCHk
HN/+zcdhZYsGvsmFljA4+RP4v166Cw8oqudUvZjVEwGXg12tsElW2WM12gzud+w7TkVwaoDtI+Xm
24NVOBS0WF2NV0Xfc0wHmxqpQb77N66hSrQC1ZlKpyFn0ONG+n69qKiCSza4nqqd9MLmBnfY5wqd
goOB5anNNgQbzJlzxzK5ajtzje/OCYt/ArXW7peJW/6ptMc1hCYW/xSEqnpiGB/XYcV6DqkkQWFM
3m76v4YdI+SVujigcyNAdRdPKO6T3j6G0/IzEJwcoYQ6W5u6yrWt6nPl1hiuWVwbX28i7QvJ1SBc
Z3AfcJclGUoOACL7V/92jkEVDEic8fCfm+K8+69V3sfsNXfsPrzzhzfD3/YK6+0Oup4V/+A2deFm
3vrv5JxG+imhhdtb5XJcXyUpI/OylBajWY0ilFvkr+itwrsNcWke0Jr0/vAhcouUpt9JaBnEb49x
3IW/QCchxYs8Eytd0DK87p1DpDBuysVRm5mvxOJYMu1cxhTPqPnDqOxS3NH0zx5WSpVCSrXyCblZ
tw5lgDJLhtf8IEWZRN0JZy6zwH5cdzCMDMSwN5jgKmDXsxZoc3JqGPu85JrKJq56lZigPsaLIxQy
0b0r/EyILH8mKwza2vOy3r5TYjNztTC5lXm//IUBEcEklw1HdKU8EfHuzryABc6LXQbKVksuMJE3
yTi8cLDIc+44uYG9U0h7s1B/2PaPG22pO0tIMDm30psC98OG9On7CGMoAYVj5mBwXwQtUKeQW4rK
xTbrtPy5V1P54P2hxvJ/OWfsH9z3dO4XIp7mmXwr3+ZDIImEttCBCCFr1BinTBZzHHw69jVn/Xvf
+RyU9xnMHAz7Nzgp1WfE9fWHtjjt8KigxycoEybm7xTLDhUR1qNYcvU0hdXjDy5bsbdVskklYM+G
gDiArEz4DF9LOq8hYYvqacmzaTcyOg4tdFs+0QdorVng75eaLq6EfJbSBl0sEradBx4Rm7ZOLn/4
bIyiRTL1gcpDO1p3wk14OdQZDFSOzZTSxGWxsZa04vtsdPUEYZTM7Hf1KSoJtz8zDgAfz8F73p23
3Y+BKJMte80NkhJPhD+S7voCyP12e+TnOMKkwuhW2R97RDUgaNj62VmWd7lKG3MmDzwYEAgvAL/P
iCgXMlIUmHmCmj2TaI0xCmY9lhKwJT5tksS1wWE7M6BjB7EoCcgob5zM0k+tU9Liz/LhfrWL77d1
hxaXlV1GLcu/UWhGx6aoQjt6DmLt3MtFLACCPBm7C/PIuFXkrfFswIckSEDE9TT6ISVyD5iYMjtF
MRNjLYANDlssKImHaV9aOjUh06EJXWCATqCl7ygj/a9H5bT7ds9IITTKlOK2mAyXSFsmGWkLNT3T
2pWnhG4b78nLlBrxp3I0k+us/NF1eAyKTMCW78zXS2wXXP4r27cP8TRwN+nXMpG3CBPN6NS6l1Jb
dZWiXXSXcgWfCcwWYdW62hxssoqQ/CRi0htzBWcm4kCQp3KzMQt+HYADM9m80oreUfSwf/D6v9W3
AXbMLrp6iXf79mLWQxIBalpKx5unaQyrysRDUN7bdtq3eVgpJh3RcOWxvl8EA2mzt+je8EyTnbnA
bBY1tcGOICrihR28yJOjkg6933D5Se/8bbNMZ6AUSgakd9F1IcbGR2/2lONk6/jJ3NPPqV6guIZn
2Ho0aUDTfXCh/gYjB3jYo3Jg+SYhKSrDDbrVdXFUJWu8135oifzJWxLRZ0J4EhoXMsTUtSChHA7O
o9Ul/m4n8TEOu501O6yaS4FiI/3JWkI8Qt5MjqK+HxWyDIVgA/4lqCp3RA3EHrve0qs4MyZYXDVa
oOeH+qHwKvaLDOR2Qf3/yyM1kiRMa0wEQfFchZUsUtOaA5FRurpFNvbkt9e9CPXd7dB9JXlTcyz3
tmhg6FIWwvPDV4ERYwanV3OudAh9T4+J+IiJwQeizp7be+uVmIhUBf7aR7hyAw4I6QVW8N9Od3mv
SzUZeLc1UCDKmXY2Bzr05IqGE31iDuOHg6X8d5SPQtAzb5Fzl4eByZ4PoW4ceCyC6hkMsgkx2jOH
UE1Y8JJyDPDqin1tZ5aeM9f/tc2107pwuDyy8peE85JrMC717MK5/e8fdy+CM0mSsr3dimXLYf6b
19aBRmdNRBVYKRr/bdv0L87pa5o553u5d5/RYeT0GrMt70nWU+XC5Qdu0c26sEvPAP/uXTuVvd0d
fcvxuCVRpNejkuZZj2/m3d1XSI1+yb3KoANm2GpJexKJnH/3eH9ka5GOucSw6w14kwGZWUbJ21ox
qyp2Uoq32HUGlwzWBgwFvjZdJxS6Ps6sMpNSWK8cC+3KBNJxvRMYawk0KvAn9T4oUnzLo2K0G10S
1NnsjfyYwHPES/V5MTrI4neluY/N2T9DqocY5wNDnsO4qEY5/PRWucOOz/UPh79k5sCxEUh+6R2k
8BD2IKG6AKOox10S8zjJDJxQ/I1fW2jRHIe3mGj/qP0ER6d0uOSEBvBBS7sdlb2ZgNB59jG42SRd
v9fM9nCt7yLtLykiMH257Zv+JViMvKuSTWoL1u8tvqkY7oTCFkPYuoM1RVoTpt6J22dYn6uiKomB
ggDdViecNZIuxYd77jtPHkln7131twU+mK6tr4MI9dLhGmAuAjYo0QmrUS82sBub3RxCPs4q0UCN
Md1+KnDTThRBRYwsdS+PaSy0ZQvRuZYWjuwljrPGJ2QyB5g3S3xUuhRex7TsRumqz5Nd56ytzvWb
OhXXbzfD4oi1shti+Rf7rh0UIbPysSdGGNCBVcGSnCdWc+ux0MVF3QN8FW8BjfFYQgIoy3smusbz
jKLzCgrjQ+ctn2/gSPTQooTl68Jz7G1hcV4OgIs5BA2qvUHvuB/Vk4KDt44tX1ogn3hgEzNrsEgV
RReSV8fLvTD0E3uqX+2OPaLVI75QzrVr9d5R2bdMh/5BzjLbCClNDNhDgPx/YM+dkSJbZ37cLQ5I
kduZWKSSuFXsZAraP96Q5lWFMKOtm1yNg6a3D+R4MXZHaQhz5JCh1Cqkc7F/YM1yN8oWIyMWXQVT
V2/M9d+FIpUsK9UvpC1CvSAevn0B1gVTUZPNCjwyqf6BpqFWpJd1bJLEvyBxOdfmr6YmFRtuKcOt
v51Lbm24qlcAnMf9pjujzjKXW8Cp1aell7SN/cUx52IMrdvfBbI6K1z0qBpG1FokcYb96TvN9wSS
GPhPmVbXwFvl2ay/VaCApbIyxLfVFQV9uoQalRXlFx+Ew+PUrioVU5II3PBOiAf0SwwQnsDGoFJK
VNs8YA1B9952laJu36g8TFEX3Lt9ci0+TmG1s4iqca0yixuex2Aik5F4K2SGV3KbSHQzFbeXXYd/
nGOCHgrWOeVjRoBXROZFJWbK+a/7i5gROSI9MWJOPxwKek7RGzNnVvG+jiUn88MYpJoy9m4fhuNI
pYyTQp9W05FhdyzQ26JLN80rnOSY1Lni6eJPBg9TqKgh+dIJujh/Wo7O1E9/ZGw1YqgYA8iBtwY1
aRNat0VxGFi00DQ+Y+Krq7ZhK6J23At8xnFgQp1Ehms+3U5OpHha4TKBHIIv7V5kjSUyg92MQrl7
+t1/kQdid1rfBJc97sZx/RImCFtQ5FJMg4QgLsKfrZBX4BL67URfwAXaALbWBjejccvhEE6+s2wy
B0IEYxStYUd3RI3eLhnx+hlhZPostrMwOWce8w+rxognu+hrXZPaCPKMvSW7Uuq6xkEPC4UBMvVZ
iGhhlE5vAfyVdAXB5AzZIyyBp3WX7Ri8dCf1K6u0SP90lsLg43CLAFn8NBdk9MvIkFMNQGwgbrBR
32w/rG8Ou6C0Z4kVr41bQR+6100NYFM3j9w1vbJxVpBWUh2nDRHqMeZVEdsne95GsYCgv9sHjeKz
hWYTX0z3ydHmS5KrGfQOeQvQT+6d1alZ7PbG5HsV1ZoQR/VmwrK0NWFOCJC+5QSIEFukFCvBaGp+
3EGH5WUKbM6SI5NspkOWIvtSKLo6vbo0QZIq9L1q5smFHJ61vC/9ZNdvTIbfN33Zx+iwA9jYJs9y
oZJ7bjeOQD04xmJCnlzL8mDWDLEfUs/l6BO7AOSuHiB61Huav9tmeB+VvAFyMhwPKjAoap3gFamH
ExSlWpVL2VmnJGpazDNpsSTSA7FALkQgvqtc+d0JGf9c45VBzb7Vi8VtPR2+RKP6YI9k1fzheTJL
CZgIR15zJHoVY0pU3QLmFuo7rPjar5+9NqNAu6+OTay6IvXq9BxGlwVmviw0S134+4OgPBS6Oj26
0+2NiY8fMrWvW7y4nR3Bdeg6qLI+GfLZgqOaPt0eUTuSu/O9+vzX2HDkVbqlgLvgRhhi1ScC/bl2
gik4D3ohWKb5FRIK5L97C7s5TcJ+Zx7tz1/QnEaPRdEc2bRAHgRr1RogbjEHgRpg+TYWNiMuVm9c
IP7nzZsXfDGsCBldzQbJ7XEB3RtQUVITgHjK66W1aHHCIZUuWvMcjVolx1T8DrdzKr6TFgTcsDBd
wj3bwCLMehtxzg5qW93ZkMunz+XukXTDxjttaMiQNNw2MA2f7Kjblyku5B9d9JfiyBfT130YjT0G
bHC921m8T+de2+eyn7voHaHOukg0TKRMIVrGVplZP1rjicECxKuduFdyIRA2/FXvieZLCY7n8cAD
3yk2G9ykk/lc85wP3VALLxt/BYKpoLM7L2OXbVtfA8rSmJy2F95grgzogMwGKyRVt6S3VXis+Iiw
yZpA3fEgrMOY1vHhBALEA3YoZ92Zir+xq6m8X+T6EPSlXcNMPSNXDwa7hJ21XNR0U/z2uJ3XIaFd
w67S71jR4Jk8YcPNEGXiHMfDfAIYXLUtZM/D3TbtJuFtZpM8IdJ10w3n40lvUp0yJxavQwl4l8Tn
MWfVwKuyBdaS7IFJCeQ7ckAViuiX+xs9ecD+/gNUg4pwlOHWJlnOB0Cz6+0jnL9Gf1lk2yACRcpT
P8RvWyJb9s4d3gghJUQR1aVWgvzF9YuUoLWQzsaWMFI+TDFK422WPG5srpfQIMDoKXK63NZS6/ow
suv8wXS9g7rbGXql1B9z+5rw8PSXtey/cRJE841z8u5g7EaikRemYhm/2WwBrt6ckesrvoErDcSY
NQxgmwoHLw9FHH5ly77oRLGMTinaKPO3uTChWiySmewIBMo51pg6DFi6Mu+/HfPNutVSQlQecgKg
KeW30c9GgO5iU7uJvzmQP9zEDlpeP3JWutfQtOX8OntPaBYbPXS1v6Su6LEt7XEuHLIZlZK8+wJG
0PxeElR4gbzHO06phhKwvfG864zdjcgoU/JtEae4BjG1QYx/zz3XHjxvaNQLMhURF4I75qZy5Cr2
cmmusqS+FRbh9jccbZeiSMpLhWm1K6sNDWHxGhg3Pt4a0UgQeT5xxabzpOovwfYEp1TRWfyhJEs6
cCJ8Qp7/IotSNSUAVo+hptcq1LfUQB6icBIwz8wnf6RMOUT/oThHbfZZvXWx+cSuMdpJSU7WTQ0j
Uj6HAthsFrfAHtJ1dR+UBYSgK14+q9Zs2l7e45pKiyBxpc08GLldpfkn8DAtLUZi+o6vYNTt/8+a
M042cBXO3aswkFwjZc+enSNMB/6b4kIbUofsJcyCr0ZT2iv3ESALaIRZt6IA1LR1xRes0w5y/Bc0
BfJtsWfcCQeaFJ/JPaYvCK4sq2ezb5RZ3cQ0fQWqgva/L8HGXt7FHGEHeF3xdloq9HNecVIfTlrF
m98UMje/NOrLDajEl7uWX6C83geaQj0h0k62FV4k2Vm1+BgjPVaEMwR+2rk7tPQkI/Vq8rXrEohk
ZB3Ylyr6ZTtINPtCLg4T7GSJRNNH58JMjMfuoRMcsJEXvabFNlNv8WDo8PKTaZi9eM0WTGruIn7+
F/rFyv+d4D4APKcJbAqZg5Kq8NSN40cphWH9CSH3aCTtUtWdhYmK+f2vSwREhY2dhTnV46/nEppQ
z+Vin8SKwh2VMgegX6JY3Q9np6fFEilEAPYo3rAuLGx4HNaGr1QdZioBLpf+z8bCgHijQU/4vsil
mCod6hU6O2SEwiBEdc+mX2zHrZ2/seoWAt4cigIRyGpjm1xgqRDE0wN2V2QJ1YazI0XcDjzbZsUS
Cn5BLKM+xQSp1IFx4Ndc5NmpMk+Bj1rMC0n7SAsJiAU+FQGH2K4NsXPVylF3l5w8SRKE5BL5k9jJ
j8PRJVZmM4e2Y4nA4NRlC4N7bqGYxi14AIf7tN7mFk+ajAYkHjhsHUDWkOVcnqj4sTurBmAeXff1
YWW1FK6Ow4+0jCIHuRpGwyvll0AIPlyx1jpDOe/TZ1CpwjgEX+iyxMq90UohVV1boEInbvQgrAkf
3Rwr0HUQ3ViLz+cPaqrDdc0Uh56m/pAVHs7hIah5ffgdW0IL7VMoVrNwk8uaGuIhRLnkkMdp7QYl
i28DdY/jD4Dk98jSkUebKpLHit0X4n/y3WfgXnjsi4f8R48bofFCLalWR1DRzv8pfkIfbek3Pzst
hIN55xT/6c69LpI8Jtd2d4UZYBIVWCuftuZUTI9OP1oSi72juJyUDvEqDZMBsjbl+bnv0/0qmW4+
UtiSO0d2vCUv+Rg306kk2t+OqLd0Ot+E09QbAELc7JwvXkKqw9Q82p9+VqWk3C3lswMtPm8gI+0a
J+Ma2RsRVaFJkznjvB+Twj6CgfDmtBCmAo540DmY9wdAQ+jSHrRsWxgE9bh5MH8DcCjU////tLGg
67MB8WXer8+YH/eIjfxC+eXsCbfTAuU508p10qSp/YTnnqPRV2VKnfVp+alex+tUq58VhtaflyA+
79rCF9tNsOuZ+s7DEG1ZOJa7udPScuUrGktt067N8k55NhMl314Qpwbx2LeDqkxgOH4ntglMOzqu
WTWdTEHxh9n1QcovimkEbwrEPzZPqi7yVonCfsU3w2N5y97sq/uKdxcqwKUWQMzKXx2uwLQpiPNE
CYN3P9fNnn4uEITiH5BZbAle6wpjZzpAu3W2zLNAx2rR7cinOjhTN3VmVqT0Hie8Phiw2cCLggzR
OpuqqH8TA4C3ri/pUO4MpnP5fyNLqL4DQ5x1COcqfe/2Sn4NMHQSU5gFi1R32QreqBR9Hl/hT/HH
7TG7X6DIVS0eWz5N9Wnc8rV+65/6Bm27SHc+PdbhLqhxoJJTpXNwBxdrCmB10358Vi3xCW6bJiQc
2eqLpXWzEoaK5TM0pA3Gn5ej2yfv0pAV/0IwjkVdN5F/JYO5ptg7odZY9gUVwBufGIn1PVELf4fQ
F+fFlzIGeV2qF6SPg3Q/NGgxW1U75nooUS0vCyJO32YAv07I0eygRiKlWyXiVKmdWlDoa7ubdNE+
RkBagZkZnQJ7VszVsKXeb/IsU0fNMuR36vHildAtg75LLlGjtn39pvKRmsnGmvgVGbI9P8CtObCI
xYeIIXNEn8hpH9JIfC4MsskYIxoHUvDYtFBmS1rz2u18p04G4H9gB3DxkjT6ybUGjK5AHp8XSH1j
0Pxb6yDEb3/gGySgU8Za/xAbzH4yB1UK8odEXdXC7Aal+znI/6BgzCTQ19A9p5aiFZ2G7alZ7De+
Xk/36kk1P2hadzuf4ojJ0XlXDc1ybSTldbDLJ7eROvGT4sAJcuc4HPK4qG7fz1CtSpP2nasgOz+L
Nu0sm+2tN7IBS4X8fSlEl/QrQouFMqPuXH1FAkiwYq9FND1fxCaKmS+o7/5owPzXevTr8wYHdO10
f/iY6xsm4Co6t6/4zbzka4sNRtPPJxeo5+BbdTgi+juyt/NafQYO4ab7/juV+YCb8vRjvC5b0Quu
eAx1hsf6dMCCn4gNaSgSsFaP0KrsDXyDf9D5jWGDMZYv9x6TARAbe1XkwFf8dx4s7MorcTiNjGaL
1XHSFTglE8YhiJniPB1IPOJLy5L52ESWlVT7qz8TYJDMSMz8lerpax4PILkfh0+S2gyg0p5O2y4o
IKA5c2QQmMDtqZNvnL7FUMbr3RNYYT9J9hO3jJcBkM6DcAJpQRbBWNTOq9u96mTPBNfDwTke6nX+
I10O6/5dIC+IRf+Ke5PQk4LBC1AUdYFFlBCq6vyEvrvYUUs5lxkdG4dXmmpV3AlBHza76bgHEffv
FRFDq7qOy9k8FCfxBo2GYaJjqLcnQ2EB3c57ekNJcChm28HFVpnijUUetuaivSC5EobDSIlYMRgW
YDJCImRA7J+jQR7U6f3AYKRi4XeA9shavSpd5W1VfTlpJI3h0BX+VQ9RYGXL5mRcofxvlOSLYCII
2rpF+168U/nJgrGAy0Q7V8oIcVHlAuo5RlB28BqAGZi/8NnCe1I0/itb0X9XwCjoLQXdN3W2dAAo
UIi+mKmnDYW6WpaQV+YG6fUnznbBpZT6hHXS0wllClcBhFoXMB6sVHNeNj7iAclP5pY/u8iU7Pxx
qDnSvzpRM5ZM35XHLQv+JyP43+TsykPa4BZLDKzzKLIyEnu0GkoJQdIF0jPDYjZchZCp8eUqVkTd
vljUJR86mJ2PQHImyTsJ72BrRLRj2YMqXWuhoYx9kx9LRDtcl9XS2hvmfiXdguPdYJyikwcQgw71
/xIkgUhEHp2Np1MVyC9Ir/t0WogSJMrL8zd5BgQ3zMgDE/nGUgnHN+K7ogUz5M9mJBwfxsO3LBbV
OP0YHmfQ9cNZnceTf55ENQzXCtyUrcRR6fevwoDP0c3ivdybGb25SkY1zcISLD0qqRmTtV8cVh3v
3KeumkE/ccYQ1ncyyNmuLQXho3TLbnPigX32BopQkF8BxngUlOgGYnu36JKndtEiwGAlM9+dDQ2C
mezS0eGt8GPi0qFmaFcZvzB9mEkMGBzcBMeVtgaQpHkQTSQ4Po1DYWAZA2IdxYudWUxipjyjjxmq
sAAfuDr9vA14Vmgu5Rjm8HztLbA4SKb+sHmLF/YDebsms+CYGEJsQtwDlLGwDPAu43bs2TCGS4aZ
oiUX8QgYlFN6shQ35xngsHmBHzVG8CGnvxDlqKbai6A4uUE4P2+099F+BjjTaf7+KVfAU3kEZt+Z
ycNFnM5bmdoB9eBbaFACGK0OBBGTavp77d3DPqgfPCC7PatYcKOtDEI8+/dKB74Yk4sSMV2BNMAG
RwPZowgPTAaizttJywK427je37TJtHHgz/Ea2j77nxR5G0S+Wujg5Xh1jdyoCJ39ghaT1kva22pj
1ibL8WZHxEH74+PkE+8HFKOx+3AYd0JVeXm19ysoHJ8uCUofaYVKFa7m7Vl5M8OBmG+u8LKztFkB
v/ZzqGojI9oPhIUTQY5n51GD8Kj916OPEkDZZUXj1013BZ3kwXRKfoimZzaVLmTDAyVG3R3hw/q5
1XmCxSjLsplDccdsqKrkEZAx34iU1o8L3a6XvbFhoS58Q0uS0Iag13U6IB3n8PuSKRxx1IGrd9XX
U3ezCZ1MWfJ5nBMwAuWZQtCNftBs25Kd0W4OhwoP2cTler7sq4bOYKymALn1mOZ/c+PxyoOP1ELP
hkT/3Tn9mRvg4aWrytgzBWtsOP8GeVlgYilT3Ib0tgw/GtkbxXrhy8YiKAaRyueuAo9XA+qXP2oR
8158Kt2C0isG+zw20NUhA0+yckehuICeWs7EQsqt0W58eloo6iKnCpzbXuw/5O79cnD5SZ13YEeb
8pENWrLXOfBhpOdSDWuQb7XscOowHKHO9LwmiMG0U2BwZEynrknLVp2KWFFOsY1OmPMhFWYdaSZI
8ohLsIW30727G8bPHZ0ak6GKL3Y2VkqR+TkPVspj6dfoGJKFkwSb3aSWOXkFa/fBAOHENxWgPyoT
SizOXR8QrqulwbJ3GmpNSYJWHYKvvyGWOvstSNYekAIiZJ+Ccc+22Q4frZhvSCoZkJV0FEXi1bUJ
KxKCaBhJj/XZmw0PuI4g0nA4rEXuRnt2QJtZoU+Nqx4ecy6pQK5aHIq2ZkjK8DsdGvQr4Rc8OUVH
Y00f54menOieXbnR90+8JyNX9Wht7Y3B3ksVkpAyf+03jReqerSDH5v462RZGBtI07XKjuhi7J1q
vygoU8jkcU7p/bY54i2VDqUVXcHA6pvY4bD9InZIzQ4VFaZjxlGFivBI0HaZK4ZFQpbWW3IHHkPj
BkrthZ4kxN7MEtsaxZngHGyn88Lcuc81I70wCXD0dRONoN8dba0mGvOXJzvJvuKUI3qoTGciARh1
hJNJtQBqeaqSdIvRSvoOvABkEzaCOjIVoypngKfsdLOgMl2+eHlbB1Gfc1RKbISqKM/JPa6ZgAw/
sYdQ+dva9RTOsv9xk8V6mS5AyqUSEX7O9wUIMsv4cxzqrDO3oQER8PjUPnKIfr9eVrIMRGRRcjIH
YHruLFf85T/TEXa5UFDegdlXQ1yofsmsLRjSzkKbWPiGJJTgNwVMsRjeUrCdSxNbyCCfkKxJTa2S
HpE/0vNd1gaCZD7InkieVjkdnaSdtWvXhcFmagFfpgV+amyPL40FH1qGoeHOjlU4jcqUpG2vztN3
OI8a9OJVR5ZPz9+vacd5mTHAY1y2fKMF992onPspENsFTPDPtDYSOge6SPkzGDlC9htA1X35xVrh
onLsCh9BJYSYMBqJdym+yOg5dIfYoWYenCE8l8R5JyahvXIjr6+WSNNfSLxkhJ+dGVtFfUccMJyD
BIONdL70x0ltdRZbWMKlZARa81Cd+3YzfC07Z5mtEn/6QxYjl95Btuqc0aUIAl9C8HTUkfYghr+i
FY2S2r/yqq3mF8UtFB0FCwHj5U94PLKOyoycoMECcfCkiaIo7ybGi1b5NyhY1qZoJh4TYVPsQFd1
QvaWjZ1qIdrqdcL2tGP31TPgUYILKzi9u0g3fiJ8VFGiW3EHzy+zBpfDKN+fgY3vU8D4s3eL2CFk
4LdC6R6c7eTytm7pI1HnQsphkOXW0DtUp1ExzhXvG2z7S/0y86VT1uTOBHfevJhnCjCxfXFufAdd
bxTn1XpL3Vuhz41Q0i6Fe+vSYW1B2k+dztd1fNoF17WyTPeTQEBfgJ7KeN35vQqXkLqVLz9wKWEK
nIZnq4tJ7DznwELCmcjT829XiG/8VFcl3YNESXUwTM24If+LfRX0eI2XTAQ3Uw/18IQl/WGF4x4A
IB4AVNE554JwMf9t88PbRpnYAqq8gzOsbGntYlF+ojibJyxWqCrQH4+tuZ5AKyxPN+Y9sI3RZXbe
T7gQeeTUGI4Xo6WERorsAK5V/ZtEQ6KGOWvBh00vUBxbyXHgJGdYH3rt+fJZtx/9/gKiJzMUOsDf
eeybPCCTPdDQ8vDH8XFnTyoZ29iFx4BacTeH4S7rKsc32g0Zx95GUc7A1uMJ2JOn76IRV4fzlvQx
S4fakpYAXRCTPIBVXhz6zjk35ZgHYU92CsE+3Q0sotNvPynjdFeR5epFPDjgdNmgJycSHU39KQsF
sJc+1EE9pmpVV8U8sPsN04tfT47Usx0XegxTvdpx6fpqrP7pGQCDUcDkMvf7ZuretuLXXbg1Vohu
HsVKUcs6AVI2YNvpIQ8i4H8VE6j9CCvwtzTyuahH9VOgGfVJPtwg9GlS/fGKcyB0VSB0nbZeJtOs
2kT4b8K4x+gh+H8W05upy+RClL5/StsqzEzlaM9HR1J5QR6ZOcE5XL9AJvzra3b/qVoG3GquLjvY
IxmXvE7hSMiknbpI5g8fdmIZPP98lyeDnHxBML98DQNU0yul1zn9rHRwKA8b0NvN3Z7nV+kALhNM
DbsBcApWWagUFr6eAj4gi/eREHFQTOCX4l4A3tvxPT6BzCznyUJIxwSKmRju4vQdh6vBHWGK+g6N
UzlKlrhjwAiUE/W9Shpz5ifon04l4Aecwq8D89DXKAfQvTicWNom8IwTm9R7oB0LpeJW4ei0xdm0
B1dooYnZQRwz5DY6XOQzTT4rbhEwLQ50zNjFMp4HZoCsT3YrFqTEIEA5UL9VErX9QFq4SJV1cW3U
4Vr+GpmCXiJNZpOw7DrAtdOSCD0v9BuanAv2Eifj2uwm/Ea7LEbnTY6u11CEQxSbxco+/FTi1ac4
hiajiQ4Xp9TelGn2diQerpy/fQsgjE/bbhNEBtQvk8KDveoXJQSB9sB1OK+E+I1yx1oJwasLx/K4
onynYUMrwL5xkQzbG5eoHHmRCDkH1PA9HYAMPKCu+ne4bnYHKyicKg1IjhvnAbt3gFnuKJ3ZGCrD
NkxhE7NRDyZk3cXNOMNingvCkMlWDErDe6RhTHBOLWmr4XwvH+jwmmvs3P1CLoOgGEUmvkPGr2CX
tRUPgg8mZFQkNvNc2HuBcfRaX92exAK1Tp56KNOWE3CNh+y/9vVrM8DKyRFpESDa6m4l06scSnqb
e+0IwKVJL9mcTxK6hYNsURW2E5x0SnwsJpdnthw7oK1eQoh/qteBKeg06djuQujOcx6op9B3vqhq
x0F7EXe21HMhBCtunolw3bD6c64zqdaO3ymMcd1/YkkA1cjfgsHQDGqiiHQNEsXSWRbi2c5jNNvc
y8ewgoPWvZ3YXqNOd5346fiQkEG8GiEc2g9GXS8zOUmNUW/x1u+Oe2VJcOha7308FMCxMFZIu3S4
2qRVXfzMYB/z7tOktLRXgCr9iI0psJ7QynHQV7MtCHTz7PoZxOXI3DH+tmqTdxnzBzVyja3u22/J
P11H47Q98XDMw9fRwrnJCnMrODeubLMHIFNdSH2eBN/qeh2kMKFmXmY2DXMf+RJoJAwcKFIn8ydF
MUCXJG6VDmMY9KSn8vXCbUk3Aw05siM5zHhJeWgCcd8RuLeDBriXu+sE+3zjFVfcdTTA/oY3jHb5
rJPbtJpycTQKojZpqkgNG4kE0LPkc3y8t0trH7tDFIs+ZeT1Evy7d+Ug/3nRjf9LVnosAxbr9kVA
6WQYQW4BGiG5Dn3KlPFEe9SbtW1FoGrDStkayr++PFUE6hyZQA+hNKWb97t8QUjq8rkcFX4aoSxp
jAei3fKP4tnFt9fD+mRZIOzidhL8h59F06ZfxsfxLaDrou6qTDbGT2BTKu89vH4OLSf/+ZZnsaqw
714n8R69OJMXODQtwhjX1+T3NmSDK9eiFvyW/N7XZxP6D5o2w3a4ac1SL/CR5JIgM3UaDyPEvppH
XD6WjS05fP//z9zpwj8LQgDAwOfYNWqCtGv4K2K+exW8St7XItsrXsHky5vFyC2il8N0dC93R6Q6
C1rmWwH0yb4ggfTY/v2p9v7bvoGl3LywenV9JMg66/YKiAbqPG24BaRb1SkNfnvUBx9XDcDGURc8
jRqBXsUTN2rJMek5u2SJtKfnTGU+KDyExRUa+scILQHDuO5RnblltjOjhAqqJnKiNkGHzRenycAG
qfgQEAUAFAixlpj9ix+u+DW6LU5iUYJKfmehB4EuHdNhaM4Rg+CXhXySddXwx0+b13uN1qPaGFKL
ZwUbgddHDWnM72DvYgKyrCh7DzB1E/xVgLCXSX2umn41Ooq9wHYuXn7zQowm0RsRxbp9HeSlxtpx
aEi9MJX/NQthHXsHYV7IclRY+6OslX6ldkJHtpfuzd1LVtXeNymQHhrkbremOE+Mv1rhxAYlDnmm
Z5lqfWIY+Ud9I/nb1Npx5+5P74QUGQW36uZVU6TsSjsLYVoMcE5JSJu7Sb52FqpWulttClE2+jAu
f+X8weIXQL7s4wrh69PHcpcT6GUG3kYrmMnB16zuggKbL9l7nDCl5iEz6BT3oINuF0W7tLWZfa1T
uZbUJG5/i+mCSntc7d4qnAaQ4HQJiOs/mjQB5SU/raYUuvInweSePOTakzjcdFwpi/ZJwjxwzsM9
C6zAqvlAnGP0zVBshP/yhrjRNV2YpUu0orOsDMdwdiTNDJWsoVgNr2zQqvMkLo2brxAB5D5YCt+U
YygeA0RczU3bwBOcjDl0hbqhN22znXjLDsYB8rAiMJaqgWQ5yt/4ESXNnG7Rh/77dyzKgEfSjSA+
nHsgGFXeK3QOsz3bLRabZiBN7eksIN84lKls37zAeAX8BV0UYzuSB+vKOh7ntCZQsZaCCF1c2+t+
VLqJVIAwd5AiFVfJ2VzdP1X4jCzVbIBDk4TnU5lEdCX9oFu5o3VjmlncID179Cj8eghphSCwGJzx
bnaZDJ5DS6h3g4p4QaPMdfDENeTK0QosxSiq52KJuYeEQSxWtG4aTc/pU9JY48WeEHh7+dAsQSY8
V1FYBU7L74L1gHFYWat/6IRKmVlOUzNuYO342HtV7baOkoSvHzRTo3wMXc+1Cep5HJXS0kdQtKit
j/iFWsNzj9cw8mpNQetKTMeMGsgwT5qmRQ1BWuYYjlTLcTJJmYZz7qIKS6KEjz3rzUwTR+cJ/FcW
zAP7n7DmFwLmYFS0RDe0Es+7ZZKv3b4jDcXBaBopRA4RNYDIXflNba9znbRJ3D1Qk6HfmqxM824R
VRxYiDbXTmE7cClkahUoNZyGbnMFSb5y05iiOgy80JkVuPE8OxR2VsshmCn2BVsulfyG0sajL1Ox
6rXg+Oqyk+RTaBXaez6u0DSzw4trixQLqswebvd1OmVCNfufKzZhplW8rvhNRzJzkbQJbO9SgHnb
EpBBaobSt4mowR2/UiBD9DxAZf0uy3TWLheVR3ZsYBuF3T2rtnMbKuX6SpNNYi90y6l192P/GOH4
Le+vPUBXAjG2ktJFdgUkn0DM8/ZT3nDXWx4258Fxdi8zwx+2nvrAKe9jUe58KSLOm/5eaF6LDQXN
AvAvJZ338sYl40DyZ2nU5vVGG8cA5SSR5LxqDeAMkAC935U1yijhipjpVJrGX7mwwNdM6p0SashK
bft+JraW+fzXN+cluoUt6gae53GhiYgdEM1SPlGSgvOg/UE4lrmLkovoaE0MbREOV4uPZkk3BE9F
UZzb1BRGjP27z6oPfU+janD/xTuIaKUpE2sHNJ0uzry5H6HsCnuzTTwFUM87y7CpN/KQC3sqi3vi
EM2QF8FBQ5/ugB+E3tWjAFXpuDFmYp8XKVX+5OIei3CdGtXz6yMFunnOuk3oXxlwNvN+Z/6Gpyxz
8nE7fc+M1mkKgg63i8X3xPpl2cRP4QbBALwlC1AsdtQOXN8OJ5Q7WFCCL5+fUCki581GnHDr0wr8
+DPDhhFKGgathWRuONmza3eSXzaQs34jWCgj2FcH161ejrUwzB63xKrcY7gFDnKq3RiwnvmUNWMX
98QhObJp4/vUAp+AGvF1QAhPYpYzYj1uH+xWqY4KwckSbjFhttcvLFG3PKcB6ORyKTK4VDvRv610
xS1CFokXnMNYL35Jps3dXKkxUGDZ9qZwu4dYXy+Na5n1qpmwlGumYbRcrysI2sGKJ3hlTZEwxSwE
gtl59g9LEGHeMazimbVWoSnSEMZG55HuyK78Fu08d5ovBI+jjJNwwELs864lWnxSjgKVA9VOSTVc
/NrjbPvt5wnfeeMZtKhMpLLhjn+iPLQb4zJWiZR+brXh7pj6cVFTLJOa93gb7nA3XHjrTWCahLOi
ptHRBmWQxBFq56G/Thfu2W65SNAHRGEv7E77P9fwWAkBKLyEjNTOycB8XrsXSAQX0UQQYX92KU3w
QR0nVNGNY5cRou97ZalbW0D5ghhiSlNiFJ/zj4U3HOuitKOo+DA1H1lVmIcUh8njpGoGpdGcDyWn
viABvdii0ZChlgJxeYq+86Zc1oWk+F5p3gkmbeM4gUEhMVQFNVVAORrA0zepuCwCouJJ5sVl+O65
AS472NOqcNN+JJJUHZYylAayc2xhxbe4s2zvPzLH3iKfW8kqIfnkDj4mOih3DRkEp/mYjGespI04
fo1bPbzFxv4/FN/cBIxDQG5+csZvSYNWpQ45JlLWxc1bbijfb8KEvO0HfoeLfsEbgrYd3bpi8and
0KNK459rtwe9ME50/01dzStn+rKt1b9MuNETW+YvRpKZUJNz17C3/5V2TvE9PatVssJSMHmVMQST
BQDZ0vdQ46nQeLee/0fxB53I4Ix8WksPVi7wmk2DD83K8huV5pYaOueCPhrqrLi+4NY4qby2Td1H
W8Lc/HFaHI0y39r8caHSidK/el1wpeq1vkORvB/Y3AWAw3Z4c+LxJv+JF2D/zoUHc8gwdZng7ez4
yz+KK3ONExSHPq+lAyZz+jifS3Nr7KRn8QbI5JFHg064N2SRKNhhmhH9E2qxTKJL/Mqvt+52bWOa
k4bubrOIFEDWFM/GpzyBJS9fAkdXs9toJNwhKEBXNzeV5jAbmA9qs1lBx4J2vIdRIHPSYHzQmXL2
Uj305xXbR9LG/RU0yfEeH49XyUKlgMyscKEZpu/W9thptLqsYodK12f9vJUOhMUL8lpte6bZ32oy
eVAEkvDhBju7NuqZltPfa+5JGmjceHporwfWboYdOEVdIYtwLEvgAV0pxPGUO2CRVOIGn3C/Bo9E
TuFcEek4iRe0O98TNBgwwsjjSvIAe3mBf5OSgrTOsXKGWp8W/vtkd/oDze6qvaT7i+eBnfnGw4kY
Da26zilvy0vn2rcFQF1KRiuvBPYhNECbzhY/W6row8criZuhePFFLb4K8ooe2sm8e6rJ6ky8VfE9
5HkzBTXO1i/vo2UHh7mcCC4cbOOuEAUtMr501deK15tlJlKGqu0wy1+Olac82mc0gUg1keUkAOcX
9I2tqnVzPTbdMgmK3Z5en69dy/+Q+UvaWh86lCa3ojfyVLIsHTbRnBDXqIS3U0YZ/V+dKIoscGqV
6GLxYBqXX2fPITxUlTSjHSNSQihfspi6ZmbSQmWvJKpVWaNlozYZEAEHDIFJKlyPz0F2TgA5X8NS
4bVJ9Uy+Uox1Zrn4M5mcX87rqMKve370YCrD1lzzHdCdbBMKcNyhB+r4eGpV9I5tAVVnBd4Hos48
VszlzlbSpSvBzdWKz7G+0ll8I0+fx6zQquNKP3NOk8eRCCdMZHpbABMbpLTCYjX8xuIfPshDjAjm
vDqOed4fJhmfqsdfaA0B918Wn931RYfDJYBzpUiL/kOlCoRfE2DhCv5MMcfHqCOsAzhPcQ8ktc1j
xH6Xyc6GyZzejeoT2sF+OQYiaoAdooj/+LrHpaK4ntzlxFI23HzhwCV4OKkpcnZtUkpzVkrxhr7a
xmxe4zjZqBKGlOpo5QZ9Umz/MRnQubQZX/6fxll0U2k2206rMFwvyRYcr/dj/UOwNYmtZZzYRAkG
4EVGql7ivoo4qtV3OwsTRxKXTX0gZ4Hnsd91szMlts1xdxTzIZ95vjbqvnWUhxQToj7bOhFu/5uv
BnkDQ9FX21MCPRJ341/yy0UkN6jDQ9WovBKaKWqRIq6t6/2C2sRipN6rCT/nIq0wXMQJnHnBPJkH
S2HUPhCjEgOIZimLEGRjTJ3WMws0KniQwKKzvn3F/li6eEXyzed7saIaAzDRNsCNAXegX1fikURn
x8wYPqb21sQmSKFdA+qxtopjxCriZ7pYj+WmrngYMt3EhxB5mhK9UeibSbsWV8GW1cheMbvNBj3Y
fM257LnD2szy4RKtzc6hfi6I1jPtRqSlEQEe1i85BsgjPNo6D62xkoJfM4ELJcfPBW+KrdUH9FVD
QBfw+kbbyUa2Q2OqQa+LqhWsqNbgirQphfKtglksV12UxQl0OvdNPU86yDitwSuGPCKo/dUUb6SX
MhRO5bQ6TCyOEgbibJ4WHQ267BTgZi4lTp6ZR0OXVpj4h/XmEEN00xZ7PjRzISk33nXgUy7ZaxbS
BRN5TWE13j39Kf4okHWskbrUZCZIblRAy4xqpBfvayiBpQz/XlwU2+EDxFq2uvbg/sVtUoL5jbT/
/3ISVuaI2N/BD8C6/H7GgmZOYppVPYweEOTHPR8kkvOxEDl6OJsOLE28WMdiNbKEDvY1hXgzIGH9
eRpil05oIUWGbZZYbo5jqlzBId5ODImN9TfhTGECE0j8RW0MpV8AFMwSJswu1mj0z8bXLRlkXqXX
Qx5txEfoS/g6nIKZIpoSPcSgVlaRwM2/DFzBRQYU1/LSkWSLKv7GtcvJS3qsFiy++GBJFxf6Jn7m
Y8tny3+8uPa9cjyTZpJTshem+XL9o2mjgUKH6Wg39TLqoNUFBsrJlxqMZuMrTsySQ1vDZSS4HJcV
UDEWQyJ5ve9SLu7Uf4rw8BCdCmWpaVxdHhaQttSwDfpiy2qtM8R9CiC8PyHEZEXKdZhwTrCbzDau
ZuNoerM4FShqUxaKNcZ83lp16tC+gqpnpFRa1Mre+ejeFCB2B2UHEdKl2VR1yTrxnjpVhPgXE/vC
CpXW59Nj/9sCl3qZ80ZrRfYFGjjR4JzPcNmZtdd61F1LwZTQvChAF/Iwtg/nybqghzGmMQ88n9hW
V2MJtN4qzFiKv/YmxrH/2A4hVU2XFU17QQuReSskCtrLwlSsIxlzC35linTgehglsK3fwbs9r4Ar
ymnfEBV6NJ9FEGvFvdnwNzNyYM88CJ3hXrNl2NHmBKAh9EFqH2cjyo23AKDKICkv14Hy8FPZYKXq
2prxPa1N/SeRMnPBdHU+EJIqCYhNIogY2kI3U9u9hmPBbiVEvFzIV2T81aENrz2gDGW22XOoxU/1
wCf2JkAe+bTlFi9JBLjd4ulepGuGuRFu41Lbz6Rt1Uk2TxQG18mvC+bTzuAAf0N/9Uox3Z2o5Vyz
FPS6nkD39RNrm0EK58Cd39xpnNpN+DzCTPDOi49tbLSZvNyp1FmJSdldbd234cGXpPZVO3btrfof
2tHGogv0WkWdLkALSM41mbFD9mzBkn6d2MEGBetcduUBPR1lGaCqydovK6WuaDVLEtGTpif6VpVH
/ZN72489+q3TxzqKLy1j8F3FJMRUDGu8NGznFigeLGPdaw13DGegky17MEvJW7TF6S8tOr4r23rl
Fwn9FCwqjUrF9Gi/cNMmZgjuxHxPZjrILkTAOGf3D54NtP0s3Xjp6DQadRK+vkpTT1xBqjFz2yZo
VeTOJ82khcWiOAMnyKhOlB0dBvHf06xWE7XW38NpobmgQpbMpQNnT9VBvGOU09RJVgufuhI0OOit
sv4I+jwvZPWvAa38pukkGjtvfKgQgXwIqeixbFb7cW3FCnfH8g2u37YJdgByCRrVPdwRvnJc25ii
V8AcbocxJVm44Y7vwM2B+eaXD3Nu2oDgAWbxXGR7JnkLjVBRRS9khQLeNrPMJ4nmIBZxf18lD2ce
43WXhwR5xtgBdhrSrNapu36dvQZ31w8xPMDGU1nj2f9Ogum5yxpD4SLV9YRq9b7XnGrOjQSK3xK4
MDTWlBzaJC1Zqk/AXaYqIUQ76yAtN0YlymNu1VKEWIazr0cL2oOYjrnlZ0D7KFq6XlNudeepASbY
cNzkGYYkm67ngImY7Sjzt1alWpLAMSLQdIImCFpU/vbrl7oedaeVSEYnmPPqTzeg8dsbQipCXpAn
uzeDpYfBx+Z+exs0NJn4d7CjQTxbe27PI+psEMd4fIU/jGZhoSM/lpk6ZOkDEZwUxyIp4fEvqoQV
i67Ut8PEsLSzuIeqaMAjd/KsJNRyKx6XhkQk0B+qarUBSsIKum3tBIpCVWRBE5Z06OGd+RCcin5x
+wFSldhmxMJKp+cF3ku1SG39sqaOhUWKqY0gw17LLPIVGU+l75xrfEojvOdyAI8T3hwHGAiRsz0Q
v6aYsqxybpTrV/TBae6/ahMBrITxU1R2/6l/dpk+wKJoWXvr2/akT83gPpW19vXYEuhdpB+ed5Xz
zdborZ2rLfcsp3pPF2R0TwzYKgJH2gs6rSFclOymHWGDiT8HLFPVZEbjRJENTb4+RHramvNSVSej
RpRhoFC+a17MU9sLpT5Y+gPd8WcZ2LrUqnppSoxoIh6UtogpvqoAWK3B3a5RAMpyuCo/0/qYstvf
bIMMM2UsN9Xilt+AdnIVKnOS1zz+6bvgR8ghehhc8+IgvJkfdZcYQiTZavtIEf+wXsVw8FKvg1hm
qGQ8s8m+AyQFsMiH8vxjBOw5F1SohK8hURLZhrd+IlKzLdYbjf4DE3AqmaAmjoI5lZ4WaVFOjSNG
AwvyZPRCrld532mrrUnsP/tEBij0iEPrkhDhV3JEABt23F7oYmVM/oNlu8vuJ5e8VVYiSBgIBLs6
A8pg8UQWt1/dPwp3zE7tD11SUhIO35o72w8XwcorR7S2mDsA1GZYrKTjRYJ29RjdPJar4nxM4Lkn
ZgrjlEXvxTCCPPey7w1rjkYc7TXOiOiC3OQcMrhAfHm1PSwaYvDBppNVt1eX7Z4nR1D8zdcuorha
E5mtPMaHSKd2vRTfwDC2cTsBsHsNzc39I4SfCt5g29UWlEECP4PvQbvRQe+enykhF4YfABiF4F0N
H+iiAjOydsIbU4L1j70N0IvAxrF+hTYHgipbwNe2i9Dn0+lS8gatb6KLEHAWhUzSi4FQ+bJ5Zz+u
gXduGeAAH8YJ0bUG1Og6fl2z2G9oVkpFfxlLkCZMoTvm2Vc7tT/dMipW11Bu3fbsxJbDZvs6PM9N
n2ov+5BVDAZpIRS9i1RVYDFOTd3FEh8h80QEFS96vxkX06+G6VPE1AaySR/503rJrL9dBAlTZ873
4H4C3jT1tc5+gV7EK+SUYLRAgHBVF5g0rTpDS3fmSm/2o/RVBCI7Dn5hf2TKryUFmMppaY7IauJh
ZlIm2560j121yUzWqDF+Z46a0kQGBZVHOEtZ6JB6UI9Xy/Mvmpe+6MMrnrY7wcyFHTPQL+sR+jIa
zlROOkzdVva5EyyEZNNADkPJzde1m6Tg3PjvwZkD2a9NZ6RHmGZ+unVA2FJ84mTywqF7i5pLCU+L
v4A0JubIEu6lEBluoQ4vzQiBEp+boiOZZi1iT7W5MaH9EZIbvwHQ78h9cauARKz3H5xQ1/PEE59d
LUJ204z4m0KV2+R8dDEDVSdBTzozUJNEagUGvUaZYn7ovvS+nR6cMgIu7WW1bbUdcuUj1IEk9GxL
UUL5uRWxNf1/lQyc6F5HOSls2yftjkh2wvxz0dfefFJOgssuI5ojt4pyUQ16cJ95A5Oc96fqosDq
STTUYedv2mBU64lzqllDVf6w3i8rB4nqtKuMsfzDmXm6cuTDKXzV5v7q+s65DThXxnE2P1fqz/yL
6kcCt9ckvZT1D6aXy0rF+VxKbG8zaJ07WQyGIbjI3vNDv56VP4+BTk/7Ixn/6H8Nv9LtsF5aX4lf
qjfZt2UvEd8DoCvbMGkJSGhQntG86/AH8ohfCAVhcoO4WefrVWDjp+2SM+f2gA5JQNyt/1lycOdP
lB2ODBWpqF/uhp6eDjlNwvueE/0hT3pomT6OeRS1PH5YNHNW7IsaT2S3jyiIXiXeGA5nsP6WScsa
ot6IaxY802W8kIGtkSEVecW1nbWuhflc5SkN6k81mK0uAI1xGjtyYhD2ZGnw3auA2s3Yu20uVAX+
+5MIMRIn1XimV2Zs1LucXFgtkjRe+HYgo2XsWCIHhH2ZfWfoQxhQuDxvwIv6UGaKjWBH9JEB0iJm
ecTtSjMoA/XaVhsr6gGOh1hSEDEOksibdVECGZ1DmESKjuTHrFfO2C8ukFgr2gm39p9Zy2BmpQaK
DOZdAv40S8AbXoDXLt6tK1THTpuE+Byf9twVHhOReBdMW9AfYKJFaneiBMhB3a1KiY0dz5Oc0fkv
omUh07v3b3WQkiMajUe4ZNlGAguzDjbx84xpqUmTgoQ38KRMUhyCH7HwRtLIsNueRYEyQyNTapN+
nchciQOXxpY/QGfCkbW9dAuqfMaW6XiYFX1YNn1FJHAiqXuX0sagVRmpz1BEegmFXmvmxy0LZYct
Wuy1isNIgItZnuHzcf9u0gXbpRWJy4eyKTfMiaP8uvcFlSxZ5A2kaY3KOuoR40F/Ks9e7nqwYbDG
F9UmLlXbBul7A0dqtZeefNaSAn5+hnlcnxuNZF32QtTs/XvYIaZKgvTUnm9WL0Mu+PKdAGF1LpJw
OnPPPUWOVgO/fACENNN3Ae6UjEpJ74GEINeVajvVppl9E047PHyOp+fNY/4dZWxb5fmow8HKBX6V
kk6+XLof6x3popvJG2N2NShGDod43GxmXYwZDHqeyvXF345B+4MS3EVxunqEEIK+QpME/fkkSKf9
8F+VttEePD1vCs2TAZs2QgWEwUeBTkRz0RoGzCG5gf8KFkuTaF/FNg/FHtHwNLJJ0W2tAzXR2aZ3
oO3x5Xf02mdS30NEmcO40gl83UcUEov1nj1P94t7wrnXSYg4S7YSqkUZdsZ+tVAviZ588QLzctMU
q8f3SoJqSEfApJhlSM9qpMZTzcq0Bfil+ETWFYKKyWJTNGkNHGWI59i5Jzu5xpcxIrVRnMRwq1Z6
zwvw9egn7E8+fxGUoSc+jC9ZMuM1fb8qIvjWKLW812lFfFOOqnnSas11ot9LuznlH7OCnciny72n
VAhjSE+5OuVuzVUMGOi/MRyP2RdZj43b9oqaI61jIdndVpRG4BsmMurQWqc9iABmj9kowzmHRzCM
RNlu6kSRwA66mQ6MA9YXM3ug/bdHCzhzH9gQ/bSUh8QiFmpGDkqc+LKmD60QUTiGQfDjaEJ8pwle
XJvLCWDNH3ThkqdYq5S7KZNHSvbxGmwMmdSmcl4fatS+TmIDK1ahKL/GxJpZruYJrv5Ki4j7nuk1
xnQ0x5raXRegvpqm5JuA5E/F7QT9C6zBoXxTbsjidbuSzt+kz8J9oTVIE+ppCFsNf/fYzKZu4rr7
TlPUWcDEEXWeErZchqMpHLVy21WALOBW/Qh9jX+/cvPaR4h46NtqN95XIIa7XOp34grcb7rWmtwI
DK+S8ss2bs+ZGjBTMaAhz7Pzu5T9nzjG5iXuLXM6F8X4GrOGJ8Rn/quB7FMPleDV/26gioeV5W0a
/18Ip8bpqT58tjZ59Kk1b4HaceMfGs7Bj3PK3H8YBETFEIRlE/mkHFp0qhTXu1ZhjsFCXgD+Mi6A
kZ1NyPG4DywL+6hhq5vWZCSWshilJTU74BBvAWv2CyiUa/CvyldGJfXRTcdCk0tA6vDpzSEcRaqg
2fJrSkYgeNBuvd065Nm54Gm6ieR20rb9c0LkIGwNwbNCCzBz0K+74YI5MoNRbgqI478PaccfDKb3
WHZ0O6s05ovsfd+9Eo6kkbDrmPmaAkqekACt8RlhH49EhloloVVsNyGstBP9V0OWrokPkffUiU1v
L+WuKH0/zXYFBZuOZ7S7SbO70/GBRZejtB/jEoabzKOnVXFrSA0jAswfOoiwLuui1Q/sTRk1FL8L
CJIXcEdWT1tGhx2yczp1TfAhVnXnhaJICeld+ITDhb6EzvtSmnrnfqC2gK5BDSKKcrEKW21Jr7rk
kiT9e6k9yrDGnjhhuSBXuqjsmQ93VhOwAWqBZc++8O6v0aO6p/VpoS4t48sITBNn9jTb3Fk2XSF8
ymyv7/J+x10I4vwdL3CQrs32FfCVBw1Z75ALHkhcXetXOigQlSRx670eVIx567+VV4sAeEN2Y1RH
EDHfW4aX5u+b+F1VmQnmrybQtsB7NeBLtTzksvnlrgO8/eND59jgbQRKVLSoT9wKzXDFGLvWu97L
+ZK59/ETGghH09T55cXoAoKwCC6o1ZI5zGz685HfSp1zLbsIBquFYrAr8rjB2hlp93vuxvuUJomQ
cn14cAqIslqi0aS5OnHsQ2hkwpxtwM4t+DBPt0F1sM+TALlZP1bZzI4/F5dh2bh+gW+UmlwY5m3w
cwDlFzpWyh/EeJRDg2ZKXARob5++u9DeC7V9ugVTMz2CcVaUfL6ly82+EDbul4qsiGhoSR1kG+cf
/TZTkdMrZr9YxK5/Zyv9Od/j7a39x6G5HfgwMVTAFwNzrMBuJhrLUTe2gPzcrxQuAdbVrWNwLB7v
VMFM3Ix/yqvbFxEwutZkpP+gv2w8bfAbC3rVTIEsW7wUyiCkVyYc4e1ztSbDsEIqm4XwtssJ/ZSS
qUI/iCgikJJ4nEEqnJfMKB2f2gJ7b9nviH3nso1V5zjhc2Vv7YTEcQ9sihBxvYsuMgoj3tjmP1PA
oJq62LH3S/ZurewFkLjBrdvHERv+3h5+NiIl2rHFAf8PRVmUnOpciD3MiMvmdzZzB7Do3vVrc52E
EJGoHoGKVvFF12Plpwe8pcbLRKPGA7YaFxh/++wqlRd6hQ2zEcP8uLFfFyvSMhUCEl66Zd9IIPSd
ftb0DYoA5GAZfa5L6I1pcJUGoK5eMhZafOq5A2YX5ToM5y60C2oJtnag2WYgrSqyYCoA/CILjGpt
Yp4TDcMs9HcgCt8V8zKD5lF9VlbAI/dl+7r7yIaMWGm0J7IBiwnxm4WLocZcKocIJXbXMGCK7rSZ
ko78E2IGD+d3UWfJe+C1oNaSmu9aAUHe52N1S+X1KXWE1s7uxlx4lpuDi1hRhvEG83jTnRn9E/rg
f2qKq34vlTOV6wdCBv/y0gpfWpwouYekfeMDRgfN0KTGuVupO+yEg5bb3a4pMoGGzKGWMqFLjC9S
pbx/fnlhxvsaWiKjJP3yUXzW4CcsAdwBAp5R6aZC/bivJYYEixwOIFLPPQJoTMUevFJR71nTRWAr
jyxukXjAs9NTPNW+QxhJX+a1RgNaAdWsM6tHdQ1ftnXzdR1lMw+DSvaoUuVyl6fv3TJDoclQFoSy
KfCZ1jKZq/M+fjIeAEfgxruRdUKhWCEufIT5AHaxVe1OZZLemNiJVrXDYDQHIm2n1+6iiJUnqFQp
pcn/Cg/r+DIT074UsTUo9LGAI70OBOr3vl9jiV3caeC6qg23SuQLWkuxZoNJkA2jOyiyWEOHH9pT
wb4BeX4bUhR/ESef2lDHw3wmG9rN+sHZi7ggrlakoq0OmNNd8HNiPuCEzvP62XHPot5OBbyOg4Yt
YrJUiYTDoWjDsPUas1s31Nc0aXxZcYauXmanY0xrm4exCg3RoeIOswUD9KdWZL4+nE0jtOnxRbyK
ygYtjm3OUU+1D+edUFUVv7xzrUEocR49x+Dcuw/XZ47BXw1nzI4TBN7NfsoqsoIIX46VcKyl3/qB
GvygKItHEHGSLAFmTrRFoqaUpMoQmI2M9ZF3Uj/9Ubdnz7Bs/QZfo5UfZbon9CjsSazpM+/DfZX7
Iy249Z81u/a7YCaO7H6VLlxoroSH2muR52ePoABojMWvygGlvMWYWQ2J9O98tBDaGUc9FdyXWfBJ
A9Iz0dbpBWCTLtPGY2KvRpfpKGCBVl4DCNzjNAttleMcaDMoHQs59T1CnAJ1U/tWwGbLK+bEtDgc
CK0lhRxPjGLRvMhub8Z9NPCtpZz4lmROi1WjlvG3l+dWvRWhZlxA8SO6+EdlexBTo6+4ayr+4Qmf
SNUAvCdthUbb3rXSApeAGsSp/0rDZGbxerbT87HGc775O+jo7R9S7pkwWAZb3C7b4h2WrIMnZfTF
L/ObRozULQW9q6eHflcukeZ0cBtTwQgDMwK0fzOI60vsiXrRgDz4GBRgIGNYPDxWv7of+13FClFL
MBvt0JRcLbLxux8sE4gKGw73Er4RfTWVv+iXeT+RX7RZDH2A7+aH3a4CNt9/NOE8qrDI7FWf8kDP
Nnm6SXRLRiZXFQHELftoLx5vmegYMWvKTYskFpoM+N9msPFDruIMAgky6mzITlfiFlvG51VkvvnF
seGfwNlYivpKRe04QHQZbZoLL9k13s19R6mWHqMqGbyqiK7wrPFyFLhnZ51tGt94QY/3hREEx7Z/
7tLV16wo1l34ZG63S7HH1Nu979wLGuMNwwNLOd3XmKrlGa5go9ntzGEEaDqKAmH9x0hzerWku/Z0
cT20PJtKte0Z5t4KfBBZ80swf7VP1B8HksMYOi8Hh9A1MaQ7eobhpKA3TysJBLXvjwh2ceqfZKdi
OjE6cVri3lKnotZPOlmfMRQ4Oh5jvMKEXNrM/eeNaFVjIwOkj3H1w673hjZGQ2Jlen3S53I8CNfT
YsclI6HEhl6GSlnuXQRPPV4vLfkSdGGYlLAyZO8KXPt4j0ZxuwUiPldnILaa6Go0apaXtOn+fj1t
xxoFA506UNKbtXEwxgO/Sh7wSm6c8jc6Sh3zdoyBcwUOPd4Coc1LPjYelBMP6B/LVRod1DwHOw09
8IhGxVb2TwNkFpUZ7sfNDup5k/YcKwoYzO7k+zQNTxmqy+bO9GIc1eEFbw1jRAqrl8SaBrVUODPX
7hi6cxobwzh73RLHSrauB+pU7Fs8yw/IhhJa671UQvNua0RDQHwOqQedCZ8DUTUd8pqsLRg2Y+dK
B5bVNgT5Somdd8IcOgX8qpgN+Sp5XnePyOlzyD1jtZqApHW7wt6w4Cw9WGZWcvJJlfnVj92NK7Ki
kPMgBYF3AcOuuBcK3HjzagTxu0S8Zuiiy10Siec8KpSp/5huVZrxuTf0PgRCKt8lDpqmu7j50FN0
NvJpAp2vZorhqIwVx6RStIHpLVEnOCrXlhnNS5dLnH0zyGVyzobcAsR947XdJP5iHVppwZO8gDNR
ucZe79Tm+cwnp7BbTk/NOEN/byUudB/IdLqHkBrtjPhjZZI1z2mhPAwqDZtdWg8m/H6K2rkqcsgM
9UfPsBlHW67RVkzxL0+KRiCneDWS30wglxoNRQhqyR61/0MZEtGjOi/nGJb8vcomY2SGp2QlCfkh
JRAtreo/odjHLh6UHQprUjtB4F4xjgDeSvYErlvUW29b8tNsZvpKYPJBCRp4xGbWpykB+Ou8ulVH
2GSKNZH4iTymajtKlGYWNx4BXWG/3jR+ICutN3sLPTe5kRHGNR7nDn+ZCRprZDkQM+lyL2v/4Psy
vmvmDrOiJnqHUF05wXq3JE3tv8nl40/eEisA+2w5x/RSWeb5OKr+utYYsHRfnz8xya9m9/X885bc
nupJEneesCL5dqLCW1tEF/mayaaP4F4THGEgYMwagKwNGCUiccHdgFJDjBI/HZlWHGgPLCrGzSTE
7iFZweyuRRm0JBp9/OAjilE7fAjrlKtAHN7qYXo9Eoxrxn1wiQ7c4hFMKhKsohg8joxoz7Avh1CC
2GaR16X2oYB0pM6sYX2jp6M3B8TO7sODY7NhKAL8YwKzldP21IvwuKhbYxHj+4EUO3NNqvCglPyK
gVfoVI4HHdhOJeTZkbOvl5vEDW5+BA3neVBpTjOyE1X3PKfbGT4b+bxFnHoRNnUZ62rVPT1Agi5w
V8FOMpC5r4A25w793340QhfAqSOcnMFP7YS0v4uYCftgB239+wvc7NgaQQOQSDQFG/tGF86PAyTh
vx9IakPf/nOiUMVB1z/7BWKOAV/xgttWka5UoxQAZAT4w4t4Heju1ALF+X0IVu/9VZvueqmJE5Aa
HGboGPWrTCkFuEQ10aDV7HagT5NINPhQ9cROLs7iLB1McvVIBZcIGdW0T6kISJd7PpUsVFZtQ/10
XfWOc/qsv23MZaqA1PleTZ3WrFBZKLKxMpe4ktMKUnYCCOVHlnEauXIFjoIZLNdSalqGmowwGUIc
VG04TOH1hkKV9JyZcHU5iuAUkI8rEE2DemvW1kOx7opcKB4TNfdeGFGu4sBBKmcRbEAHoquF2zW/
8Tv0ZhtpzfbB1Fr76ee08SQ2GGpDEoWdg9THujZbd3JK0GkRtzedUyDlkcGL8O/l3p79ikSuwHnQ
9oA4BjlJcMwppVb9yljj86ABxDtP2AWZMMr/Ri4R+t4BbK2qH1Dppvpi+rEQEw15E0h2Ql/Tmko1
U4j5awvE/eeXKM/97F3Mho48cAg12615kvcNTeZ1OaTw4RQpIxEDwpNviaNG1T7fuREN9jXAAsmt
LWVYtoBLF/PQYweKTUqt0qbq7Gs9caXWBk8ZdX+3nIaIWubNo4rIfnn4UTdIiRNVnTeAogYILTTc
OPoqXqI7muP+GAJlPmlPw08m3zgdr0lam8gsGpn/NGIhrUXJOdTGQdHe5fgPIFD5iSNgtF2/2gOv
R8nug0Id3I1ZiRH+9wYcRzvWwdMdSAjaSif8DUbn3mOyueQ0VnFK0wImHoe7ztkZsIPoiNKO8KAF
kGP9FFXC7yZp6AtZcx3oiLgxIrMosWN353FgmrT1nIUbBw6hbDb25cdQZ0//L3IytoXMtGXfTApd
I+11HL9dEeJ4K6Tn90/xKyXR9bV+xFg95LocqEpbHUh9mgkdvZ7YP/wgbii17BuL3kzwuW3lnQa9
09bxoboUcQsicJo0sGxdqJNeYZpIyvInkv5Jttd6VPHnydSW2hjwLU/ncnNXvLubnsQoYVMDTmtv
OIjLq+x0P8QJtKZ6bRBDY6GivMcPEeVZo16aSIHqJ1lbBvmEZIV/r0DwL46XfHfpvyJJwsxslZ5I
IGNVeK7cIrH9hOycxlvU3PGNsFQs0oiJlc30bTVheeoqpqjJNxzTaHEmTVG0yIgyabWIWwVS0y4e
Ml04sAu07UKNUHbclLEgg7b+eUO9ioip/xX1KVGWbMCCqXHDSTVkPJivHy036fXuN61FULQgFWOC
MmJr+CBAZTz1HVWuJi5o0G7qixzBMWq6RMC+nbpyZ71O4j7ivxhR+gnrR9pez44HYBICojvI8HyB
Q7AKf8vg4xyC8a8BZOj3R/iiKB6ppi8DPGcoCbv//rNO9mMm9YsTY5UZk7+VTYs8aXpVwiA2sG/g
rDD4OdgHHClNQQWdO3ygmEc8xo1qvK3/RitAxwvsETf2v3gbrmcK9lmYxpf6LhbZkvHrFIqXfJtp
ppXbP8VUDvig03QfxjTky4FIeYoZy9XJglICigYRt+7vg4RcAai2nGYjFwZN0VwkHMiQ35gGW400
eEfhPZOMDOwToiqejxC38aB+XSZjlZS0dAmD5MquFEC6TOlAv8292cwZwx2ic8I6cRFqKckjQzU1
R5Khj+72HqsyX7KyYMnlb71rhuC3HH0/DX+iBZPK+i5LyvOpLJw/Ercp637e2ErBpMT30TnHdzSr
BI6THxgc1TMHeX2YuymKhl3EusaHLgFC6FFUfEifLceZRrW8g9Nem0o/GxkVV1u7AyoF/1eeYKyM
2HOfuw0ir+uZCf/4DHuIrBmMy6FWHN1oH9lPIf6uq5xWDREHr3CfNZklDUafLeSxYguLzf09iVli
ialRL3SWH6/3JRHnU/F7mE49O5a7lWo68vo1g4+aXyo/JBupjOOKmKM+vlxcg0hi+5uDXU1aUg0N
wJyee3yPeGFJ62NIm7+djz7G2jcCMIYNjs8tFfDXxUdYstst6IhTpIBUc/86DNx7UAgXzu3B6qyC
7ckXRA6VzBikExH7730YJtcR3NafuKOM0OS0iagZZ9RyS4IT2oSKXaJt1lY5cK3daQC3cmR2vYfH
Eb/GFznvwpzQOacPQmsZcpw7EmTLnguDH8I0vYGsHWLgAsp/hqQW2UDWU2DrNf9aV/niZrSZT8MC
Ia//4kEAko8Fgdd69AQsjqYSYs21UfSrCIi8bTZDD89DdeAuGEPoepniBV0hDBwr4bVU13FqG7ur
piUatZ5CH1OComXxm/SNBFos+wjxZgnlMzGXQv0PcQ716qSIp6lkMekNfQC9EUBxRsWaXRRRUZ4Y
XGbAiado0e0PmX8D4PYw/t6emZtWkooJbFNjA0CAfBCmrhHu/5fFZubFfl3XL0+QWPSbaUZkdCY+
wTVttFTuUlx0O7lfHsTaRLX9rxh53Xx7qxySGCtP3kM20lVFbzHgJRST4+wgL3B5z2fn4ErUjASe
uET3gLhn7c7AA9VTcUWL+e+Fp8zMlqdPDaPNkArEFfI0iiXknLs8qby0EQ/DXbxQvennKlyQ2EPI
jwGyAt122gt6klahtIkj5cOfZYACiAQnAmJd5+jlxxVITIGYbtD2Vlyoycy3SkJXimB/B0++n9vN
ISX23XNOEwwMA/RID2Nn4tgd2vuAwJVxsDL5iWZjuZJSkFiAGpu/FGjcV/wpNpUh7prairmlqMDs
YzaKa8HW1eKar6oWBOVB1SHjdRO7IngfFJC/zv6YIfpppCFFBF7P2jMvFFQGScTycuK0oRh/k5wW
HdOJPD0oyeD2SRnyPmujsKHUujplnCuE5jCWQti2PrMJctV6DivEusOmQ+NEqDEOJfodcrewPGzV
+4tnqq4Dl/+Xy3XTp3g0uf6jm0jz3DBBhtEU2vs9KUVbrjZHehTchlFIOij/ghxqWIS/sa5apOZE
NRM+u5NigjqNXZ4HgAv8LOu1EbhjvE6oPqk78Z6f+fDYG9Pd+k+O+p3C1jGzhgcKVvt6nRQd0e+o
d0I33RuIRkRJr4Cu/AJ+qm4jHIbhr2PDjvqgCcFBjRLkyhR4kfTi+kMoOPdhnuMJc7noK+Zk+qbY
kboFEKNiThoqPi8Me3fmsHhwVq0T4L/Q6cNPWZwNYXi+e2WfCRuaX4BIAhoHnqfgZXyy7ox27vVV
QfJoxek60b8wWRk6gahA6Ul+I8Fbs6vudSftN/UpDpuS9+EsUrSzlME8xanUwaiwMaA7sv8RDveb
FAUe44qvo/goKS9Reba61LNBGw/t5d0rk7RShwxhgzWJZu56Ig5Lx35aZgsSXnffQ1+GHdF7EGaW
t/KGdWJ8ztUrfe++HftoBla1/pgbHb33cjN2NFk3dCUMOgSYIMn/zrf0xEc42CJN8d881XWKRawX
cCAN/PYqsySOeNOa3jUMXBZGbFaRlj4FdD5KcS3WIQUJuM7sPE1P5gIDxf2WfK7ETLJuGJA0/WIK
BebGpp3fsnuVmWaBD95Yi6sV8Qf2/rW0Lcu2bKoxyqpifYK6V1e9icFlT056Uc4g2QDlYyOvPSLS
XgyZCKZTYp90kd6eEBFVhPD8rXNLOkIoBZUmiJ6Df1olvBv9c12KM38j5bLeBUIcNMunTxZHFvMw
KKKdkhhTDxaX/2xNvPFMrtTrZCFSvMxnP5WJ2cjntDg6GyaS86YlvY4afK6gZ068TsOqLa92TzLA
PJF21dLvd9XcnYGdxYqFlkgloePX4yIn/hbIzIqYP9D7pZYm2bYNv3M575I7qUlXh7Jp3yZiyVy0
ubfBE/TKhcz59h3tiM9vXiWjTO/Ly0lR3dVIY/68KqOQbrk1ZKfVKX5yqUX7YCYUuCYnxISyaJ9D
9pggmZpEoFt7DaSPxMPP6XbJlg7T0ibC6KSXvYbRyWOWsMJg3Garn8LAz+egelSk/05IQxPjO7kB
YoFjqZ3HxMT4GyWwTLpHQUFyECIem4VOonWH2B/f9122TsmPk1DtFcjqckCaToAn0OhC+oSlfltk
MMJADJKzTvfm8ZhS7iYNG5UESdZy33yKLw6GwfG7iWVrZLq47QijAeqnLI+pmT/B5sZcfqujucyQ
nBpbBVyp6TEvmoY/X9PGk/PbPsWC/51FyYAFQ+7CmndfLQ3jP1gujPSFYbkITBC5ar+lcZTub2Ad
Z9S/DxSoQEu8z6Qkz2v/X2SvordkXW9Rwgyuis0U/FnHjJM3J4f9d6AONt7639H5xbfs4z7U4aIy
P5kAcSLxAeKCpFvI0swl/wEBe5pqdKXIAjKce1oj2B32hUku5IUD1EUcVecC7Xi5ppwvVLLe4XEt
0HC1IArT69gVcZGfcBognquOTH6fH/1YraoAUxqvWb4/irXwu1S7m1ubq4/Umw/63VKqkGE6Lcnt
CRGs36hSfbAZAhCoN1Xqpe51MsaLm4KFp/tpm7nPq6HqCoBDDm71/iEAaBnWK9nODudDf9o7x7jn
9W8MQQTIfibekGuiwEDEsCZvr12DXBo3jZlzuBRZyp2/c+itVOHEU2RvNwCP0k3KHsA8dut0OEcC
r+EiqPC6dGLKCxaNB16egUXajFsMUlSHOX3aI9Ps2mtJr+D8QNFWzuGrQcEP+yrMho2O23BEUvd4
/VaEJ01w22Z/xGHgNOa04vG5lh4KuNkclu+a98dLjMov3bslSU6lB52aYbGjeR97bT3ROOCw52Ba
qv6czkG7sUPyMzmi7TZwHe5p1IDUSIzd+VtMJLTSkgufAijsfLm9xXcGyB1DnjaYnabvgthcuhrD
l44qnZ/FrnRzkksHaJgyDbgDPis7f10yKADiwxaSmQAQEjfILJvAflbgr1TfUSIlpR1DfEtyqkO6
Z0VTL31/+u3dcyZMtSFdt38x8mBoVAVbwCuZnUx4APHPCjBDJ3trMtjNs1wE9W3Qz5YZsC4wkhof
c/v1Gg8hJu37WI1GgAHxe7uGjTSaoMYOj8en6lW3EzlinrLAIh3Klm9kP2yXgXXeUfWZO7mqHUan
o2Y24soNl6t44nHcWNXcwdocsry292z8JHChOFP1ySSBr3UmQXyU+3h3iykK7crwBqaRm6HYn+PY
F8riiFKjoiF9a1Tuml/J3LXPYQI+OwB8Xbeu5KFGcOiU786CaVnYQIXQTaA3NfLquYrNVklVVzHE
TWdKnmcVFsx1hAd8SVgGl+OnNwa3Q5YXfJ9JEQUBi5GrLesd2JH2wjBouKccnUX3gqhjxgD1pJNm
BwJpQb57VOKxN8gnqeQXatqKnMgS/MexvRHw87MGdq+9mzm/+huFs0C4KhqKwXgVMSHrmF9hSvhc
5tuA0sEka60+3d7p4YRTSPe1Xnn+sdWNTpusjte/Y05GQ7IhEI2vEihSpv6BZdFKj9qCaLaATHdN
Nd1I87+0BOZ6SbxyrLpOQ8+Pb4oGe55wXHd/lCDFdEwaXwozLyhAbRodN2jXRdQXU8hIgP4rwzW0
uCORGoNQD/M8kTEoNFakbvdifCUHdHwmkyKBYe5d40o2G4DyN2bqKWGHDYX1VJEDsgLQQxtL+z6y
Ykjr3kEz5QicY0FnzaqQ2swmaMLWYl/lihmCk5I70SUL2PdAPDjDFRQMQJKgL6rPPmrJigvfG/g+
M2O61sEpiINkZUW85iaHUDuIHXIkpa1FjbtBzEla+juYoJdBJM/6F0AR4laiwhD/nehL4Yut0XsX
2GgkgCrbEYtHN5SCvCnjUd8RzxRU6pUNvNxjSElo0PaJt61KtOhFasOVzz3EN/T9Zv9kKZE36BQN
tuznASnJ1rgzVlKjE8bCVZd43tt2H0newyw799HyxhtjX+pbqUyLdwSryw5yTzBNBk/0NAwGr4If
jQUw1gQ5+2IcUefJ00LCpVwrA/WdsQka1+lVsoQS+/Pp1p5tjlGF0vZOl7qpnJrI/HO9UQdpJpIh
aJIQPiz4kDuLIKs3YPUuLeSjViiHfC3QFgI4BlbWqBISlhtqsnQsavxDn5JK2UQ1uHM4AIuShBFa
L9IUKRU52ol5frHTtV9X6p+yabkIqCaeIe6Qlr0Y5LQggrLN1/nBZ9iNMvcVbwRcFagEV681S1py
ApqVJG0SN3onv9ws3JvJ5vEcUVBM2hmhcJObvZnZ+U+TF0Eqg/gcoyv9QUfOZiNfA05HCpNkgjRS
llLSbV+Sqjno7c/QuDKdNnTSIs+3YQq5BAy/uBGfKR1gTZlEe7GEzmnfWvPSlEQ8fWDPi9aKN8YK
Ye5gvf9CCTPRpYr0GSjQ2a6pDK9UPwS+bN6fP06lBsxe+/ucPhXbp6QA11IJ2udpHEMaugCtFATs
cfGOvKpJvJwwo0q6y6PqGy2fKmxlodhvkuU/BGd66rkl5Qn9kMhVXv6UFk/nAJW7sWepirnJUZxa
slkKePfoD9b9D+10mKQjKq55R3RSRvcVEEJ+/OwAUUvqElApCNy5cJ2wmD/ML+nuQXAT6PxWN5Bn
rRjZdxB5pqcFuXoWO9Dyr/S6wvYvmI2N0iIwb7dl6Yi3Ytl33e5rAYq/UL1REBlmnLB9FluNFH48
dcu+bv8CoxSZshcZ/rp9z918/F3h89jO+MoU9X63OzMj/V677k0ue60MXZQS5YTgF0xcvutuEPiq
u3CNsVySS3cprBcwc/mlrWwaAaUtUQEZ0O8r26uFCUC90gYmu7lZhzSA5u6lh/fPZarj5PlQTcK4
uZrr8g7XisV7APOt9/v3xGoiGBfwQ0fArdNEpd3EPu32ny+y1xNvwyrFDZMLU4he13Bqn6RQxFhX
0eCc+tUovXaMYazmOcvo2OxR3i61YE4zF9LsZSc29GYPLuuWqLHt6qVqj3nHM+S8y6Rmj7NIIJIs
wTKMqJvEZdndwJqoU6NckvrxREXylYkqstEE/paob/AiTrBSrc6ItyDTZRKEt5PVDLHSvFb/FLvB
wRRy4Nc+rjHON+gtjs5tNf/i7ETRZ0ASegp3lU4mOUxkC1lykCuUrAhmmoxWamXJjPZzPxLnjPEk
Vfdpr5CIRJ/OA5lbtfD/FNpRfrE396JJ4Fbgsf/5oI5uEki/y4LATtqXX/i+8UhoIubdJGbG8XqK
EacHQKOC1OrrFZXJTAqPP4kQvI0keADnsqTdb+NUN9jsDBd2vIgWIi0JPu2qv2NMKQKy8bLsp3rf
YV99Aq9qyvhspKDOOTeG901yMqkZ2LSbuiw+C4CgyOz/q0yQuoGeZhlQcruAe7ZpTImLIyY5yJtA
DWvxB0pgghF3lDvq0CuFkJXAdf9HZ18+dXz1gk84F2z6Ko4PiDbRG+b7aLVeC6NeuLm/PlFA5F6b
OzcWySfQalw0BUGVZZJBb4ouEl0GUDnaNO3YkHO3Mx6DpPFwwK/dSJ3tz0Isabugj/J54P+SmRnL
Y32invtLa27iMfIiu3tYZMnumE+zDLyWCguErxAGKg+n5jBhEQr8BjFNIM9HNm1iTMiKSQSIKM+5
m75CT8nqEnBmdzB4teun2E200wy8V6kcYarrjG6nuWxE/hrdv7vp7vsQmFcW8Olz3BQZZzdNJfcR
Uu6IyTVQ7XoXQHdzpMZzpUhMyxgen0j2pw2e/sdim8YkovrhhtMy5FL3/JChZYeL0O/8Xb6kBU+W
D5458RcZIG9m7pktJWCYIxh0kBbORstXRHGxSwPi61YUUpe+FUN8HqF2hUBYWlPhtj7E+B0gZ3yC
IMlaPwPAo06EoDGCkymYzaaj9SuAG9YfC6s3rEeOpPj0KriWcXKIsGYiEmEPJJT4okqJg0kuef/m
6BquFVNm5FMoCg50GW3luJcb85m8hIHcuVG6okogkM4ksBs006RFE/ReubINEDZMNrt7Vjn7IVkj
1c2N+YMKyIMhSjsLrSyHLFxQ36w2GIkOWh8BbHkRJ1/662qNvvGzb3zu1iuncoYMpApJzAE40f5f
dgFPZeC7HPhgV2OzJsYCDki0bSR5+1mY9z7xYn9MGAAkkrOoJWlSxmxScREInwiQ9mDAhmYKBeeb
GpS+oINI1eO9yrvHuquJEn07RNIuOFt7ob/CCTK0W9X22w9aCJzx+TMtx9gCqQtF1Pn9OtboFAdz
PIGG5Yh1u2ZWQhZbj4twKUA3b00IRVq6hov9RoLCPjcJGhIsFKYf0Qz+bYO/Itxn78np8CZeT4uB
OOFN85PCCq6F6P2VgRFqeB6JVrv4vh3Yp0rSCBimm3Hz6X+ChR+ktdcpd6swnCRlnCAAyTJadhtJ
fKsUXucmXq03N7cjPN8+Q9xkK2g2bLGvrwo4Snd9pKAMenNmD+lBRLKPtbfq3nIRlAN5NE+6fS1L
BnlF9e9LMxjXx1JQefsybFyyLOj1o3flMdhs7nlKdatDYSA0QxfE0mGMY1VwNWnaptCWe73McKc4
rA3fbOYKtk3y+Lvid8z7e0PPZ/HdSE5/w8bo4x1bNUJzJUyuxzUE2E2gkdh28+gs08N4r2n5jNWE
eAT7ozjqstJ3l9+riDpeLadxdRn/9VNgPudGgR18L1L3+/8+WJ9Oull/s7ek2zJtPwrZzaaPRcJ5
BZhOuuT7stA13JTYOb+yYtnrZ1l6qv5lCTtQ0lE8WUOnw48P+o168ywZZozk884VTdL340vL+W5P
QLJgJje6KZSfzv/Ab3DEFKB3fk3/pzHbtGnjbOU2wv57GUp9ysOOw+Os2a3dgliHRGHjo4w9S74n
j3n6j7lkRfaUVCulyi34MU+58XFpxKVRRG58YCwM3aZ/27mS49MCwI8Untz646yAV0/FfVEJCewx
dAZoExDHM+w5H6yF+sHHzI8/PCpcyHDPhXhQq/wOVQiUNm1qu6ZIKjqTmUiRwNy6KVujhdDlzt7P
ztZe1tLYjaseLKp5TGW4UYHEX19EumvMxfuEs79Wa1P0nj3KI4OUFw/jjZ5+8uKWnR+mNQu+s1kI
/jvHYvwyfp3fqKlASg2qA2egwkM4ln7790ZNOJR+DvFQ+W78cJTEiy0SG32CJgJPNEIFeSTy6fT7
L1CtvbaetV/O5xyIj7gzLTNcvZFQN7/qFZLAMPN1r+kOjfsUrync8GvSKsONtzjrTg2Jkl9weGnc
QMYN1gfGupS6+cInzbijaF8MgjGnRawW8SPOi9r3s7+/7qV/2ARjv0nOME3fsntfhJPVoJa2baCn
frUT7hk75RxS3zqVC3GrM9wT8oIwKV1+SBb58qdBHubmB15h391529YzLL0r/apdKfr2P9SzOf8P
79KXC65IlEuW2sW1plS+bnUg30dfWU+y8wMUUFzyiLiPpM2NsaOIP6DQcscQ/48v8VeoMvoIrDWN
Y8n1rGOmy1k0uVxoT9MMbSpHklYIQT2DtgNRSCuzAkZnNfX+s7KgIBBFsiX9SNNdF6sfVKKHmLOg
Ug18/hrM0Kpk5ykGG960J2AygsQdW9QIXSne2eh7zla2lYWmT1zHT8mm4wm5lK69FDXbgscrPqAV
NH3+rsYphjKUS79/WVGxepMaVGADAE1WsH7OdqErPAv2+gxbOaP3F0R6PaUBZ7TZMKuhoUH17lnv
JUXoE6pBZQGFmT3+DCuPY57rZwOXOjxuEy32WUtic91jfuvIOR/Ewbm4BJQFCPL8WOa3OvGX6+AN
QjSnw+5yvVAMn96ujSY87U9wG24e/67rQSWUe0GwdEPhR7Aloo1HgdgvoMAMIEM2NYVFgeKAzKdb
qNF3dPYXSco1oxQeknRjJgDPu4/GYe63L9Y8SMptbcgxjDF4c0ahNZyuM7TVLQgGjLPwSmnVoz2B
LnviwhOBqWYaZSbABMLLdYewuKZSb+vTbWG3PepnFsrCa0muYi4v2MfBo48iys9VvrUwhgRGtcOF
t4vg3XJ9Cy7904gQ9tyDPz8UVz+qLM8QrhurcXw1lQZTfseE6dDW5Ya3RsQeONUJY7QCEw5rwEA2
aJDUrTk/1gqmhRaCuxDCrS7DHQr079anTMh3xC/V0y/Ex4vLQAdnZkOu2khTkEX+pZV36cudJK9R
W4Dt92+jmLJuQZSwzfz1LoGGMQzoYjeWEXPiNgawpWonEnr0oTSFODzwktH7D70iLKBzH/A2LuPy
NpkO6cege0HBxrhBisiUrheB8LmnhmQiJTJHX4nc4J8QdqEMDjlUZLh/F9YM6HrUcielKL9rGyGV
qXQHDvOa1Nl/SGlYgwn7siTDihekbbcaCoVIo4x8snmiRtfR6T5E77za8H/Ja427RncCyJBBI3Ua
8Fy6Vm0t4VdeZfRq9O+6rEym94Va5CtTfuQbFq/hvrqY07cHG2tVWxxWw+jbhinqpjY6MavFF9KO
7c2hDoXcfCiYLqhJNQCEgI6Iq5XcAzyS0WzS1YTkJ+SzFtIPPgfTpFK8HmJUKRfsE2dxZNsUu2B+
bwble6bg4VAcsSMQORSzQvrTZ8kXYX5M4QPinTOQVoPoNszdcAOKmMgDtGxkBTw9EF9hjC8Tcvcl
y59aPmd/nmmeHKgwnlxte1xLTrq28yMSO9FWuVq2nhnmumdAKwuE122QkpCDOCTzNuyswZuKsA+k
6wbuPVNmdCoAI4YrBh/9jntF8bB/JAE6i0rpkya4VkqNx3Y2ugyqYnjMkTyiguGVAwd/1YNqCdNY
kCDBNwAQ6jYBspnwiXe9EmClWoTNNERWfVynt0BaRHZPFQgf1rqqeU9oPtzMKZeTyA9qNeBxBsV4
FSl1Lql+fCL0DJbA7UJ9mmGPj3l5Qls/fBpxWmkaHNShqnMrDnqJEpv5TYrOyh/DxQ9rOpqLHvVc
6/JLR2xmfI8orcp/EyZe03ApJNqSd/FdgVCiRm9+t6Dw2comlJW2ZoUwQm+stD1aOH72EEQQS6vb
IsBoptYg5YVA4PhDGwP9oEppXDzchDXYX6NgimxtQBjfANw3uccdwvit2B/Qyko4qFRRKdLP64mi
jBpvC6JL+UniVxP3LPqQNTg6MZ8HuwgbkmX9di9h0cHIJSpxykMY6NZrkI5pDyeHCJj1nyEcq7I3
xzLUjFIO3HlWSYbQ4h0Ocp5As46yu0DXIPVJaXgPme2gOIzYgv9rvvTiVk9huDgh2cfFQG+80ZMV
e5VnywtdlV/Fqmf4kZbgQ1fdW4Vqt1AoXD++IcxKTdnNmwsBTHEv1dJ6dTTqrwOQwR/mvs5Z8q8V
FK6+AOoEHZvO2lXr6glvxVQx6Af18kmIPRupuuYz61dOiikb/m73oIOAEY/6JXIxpP9ury/cxfhZ
YeNgPD46E8sn9jiPbC/9Zk3n33+6v0iAvfu/2PyJcobwDUiejJSEeVY6c8t7HK0yB604n57+8oVe
yeyFfg+gFtu6341OvJ4z1fAfOLnaIMs/kW7JD52e4SMCpX6n1aX04eNPVYw49B6HTOM+ek2j9CVm
61Z3kGrxstWR55GqHcMbfl4j3x+KwMCZppwYpxbstu/ibSbuX6yXtZbx8J8+J9PG40g8dmTAIMgU
61mqa+3r8fYzu5dzkd4cGtLTYBkM8VbGAPg5O/rdQrm03ykr7TyRt9/0U0aXFKWTn3SfCCHeDpD/
vvCXKYrKkSUJzoLAG9eDWWpdMh35A9+zPrv0L+phVeHTixf5hA6AhmY6CuX/ljW20pZr4u1vrMYY
DnQyFOZjouQ6iEiOZejUj7fGmMbWJ0uk739OnkZ3tAHXMPtbN4cohbGbm/fCchN66KVkjj3uvHu1
/hih5xHmMLMv16CxhuWxkNE4l/K39wAK/RfvAN0PEOcwMLgaDouptTiZJKk/s32i3iyNuCVO49Xr
4FGK2ANfCpNnZEbsni3iUVE25cGGbYXje5HWfg3WoVcykBrN/zN86VRghwoK1/uZHfRsYh8n6wHX
G+ZFZBRWTjSXY87hN8ZKII3gW2OXmPQWIYRGJ8Rb0ebCnhfKqLX7XQ8lZoNRkrc1tKcl6JBwnFz6
fHNiaupX0rYVEJKitRHuuF0yKo80p13crhoUgfyVkBI0Prvxv9O9SZegbjPHhS9sHp4CJe8q8VI2
eB43mPml2TPK/xFklrsOVFXSF/aYOnQWPeg8Yxwid79dbQ5kLFnvwcAtRafYL17362UAyXh25+nz
YevIWKlb/pApEql7BM2KOgG0g7bwLCCaOpx6bt0W22jH2A87Rn60FwrN/exk+ZdAQCRdYagsBLPo
7XAphhHto3rofUuj3atUEcUWMJg37iZbP+kew8GkjqvMXuDCxDPO38lj/omgB5UKSY/pw6baF+sr
GbO82E2QFW7lVrfosOFtVCriMtHsy4boFJG7QlFO6aq3wke6c3HM76moexH8b54ihgFQftGNxjDV
DEpfQQxQE9rr4GGtdbSlNvjGBVKZ8UIpBRjKEMLkn7FuryXWS3SFX9kINvkMJiGKuVkL8S4h/5+a
EydLrwdL2q3zg6aHsA4UzNZTFzK7pFzJbd5OjH2wHr/5FvykVjdn728msFkXaD8T1PDF338dYfSr
QRwhUtp6XP0OdOvcUglXb14kWdPenQOKEbXYDGmxaAXoCdsk71D1VafsTCR3/xNoLqgZNvWa7he7
NSCJjTVSp8dO/jpQv+dwMT3RrlmS5qk2yVnN2YTtdErTQdCVP+tqubILwzldR/esb8CHh2ywE9J5
ypVBVfo/CHLtFe/2I5G7C6DkWe+0BTevn7O9iTE1mN4nYdCXHyVQKk8LR6ftiWm1jP2d41kAm6eC
P6BaMd+8aMEsGpmvSp7BQvlM69rbTIJlUXDb/B4DKX9rVpX9ZGpf9gRaniJtEdyZQw+B20ulP76e
fJVwmHe1cspsuVGHPoTJWuqfJYkfEHuIvG3xZ93h+mDqWfUSlcn425YBlau0nThIbuhJodcbTkXi
WFfFA2qjTKavCw7022uHqscEXDZbK0JoTg30xhipEwfPks31Rs1W5db21W5vpmmGoJSoFqoG60kG
ZCcc4kw1O9Emkf3lISsoIz7vi0MOTksrR06SrGi7y2cZUUTeAtRjz7pLyaW84n+5dLqD37+3EwJX
s+NuZId33NQzTS7Sz1DpvKXelh1r2b6P79ORDDdQGwqoI58mu3ZNaihd3lzheF/YxmIOth3Xb0IL
SK9iZAUMF5k1LfOJrd88W9CA7E2Lq39CR4usfQxz0+lQRd2XmW6XndYjjT+nyzk4pV9NRg9vYkd6
Or1tzW3Q/yEbC6RjjuX/VfrHJyD6wy3PORNu388v01Xzqo9613WftNGxk8QcplIMRMPFgO5+ch6H
rgZQIrt8Zsm7ddvjca1Ow3G/ITlTI54vl5q/zr8aNHTyA8qr95d0+EUcCW26XuKWjFkZWQRNV0D0
67exgdkK98Q9dSo1gjTjmGVSatcWhxmIHvO3UtG1cM1XAutXwDDppWEZIhlbU2YQSg++IotkdsnO
dYdFL9TUcrBZbCPVd9r9BC99zf2+rEnn9rqSfk/5WUGsKzz7yL/LCSthpxAQvAd0m8anP3JG0IEw
RYhZ2WAGtBa5cnZpVaYbdI433E5dvMGAPFFjCbWYNXjac5S7g85NMKof+tjqeEkgRggT+CLcJe3O
Vslyis8ZnH9ASpc0CHuMgeZlyst+s54Yf/EAhmSpmInnEWWoCau7tsV4loNmGzHj0KjhP3ysYwwz
ZS4VI8XZKZuAajS3kL32SeZkLfxlepZWhZGpB5QeKYTcv7JaFlmqVkke/VoSSDSTINDSmwgwwa9f
dp4xtkRO9+KcK+26aOFLKXMlasJ3otXnP2ROTgPGZ+HCtQzu+q1WlpDp3+gzwjX8gScRrZGPWEBG
l0jUlMibbReRJn10SiBGu0mwhxKkbgraK6cwsge06rodNCZzPJYm2Pja50z2mp6LszVsbGQKy8S7
6p+ihfJVTUQKTwwIktlju0K7/vsdPBIASwx5AXc0PWsSEujEN3wXlh1oxpd3SBd1VEZK5eG1QcVq
4BbnXX4mvx/CZ/ylCgBx7w+TuHqaZyH5DI7+dL5XkhjQyJBbXh29657k23PchRXDNjvGv1PRJ5zb
+qEEFMqLGI1Q0beR9aTERfLpHWUcHc6SsirrJcVn57QQ67gGviZ2EVcwsa/bpW08HGC5AEuhBDh/
0N9eaA0I5OuBveL6Z+LCxpwpVF7mm77QKjSpWChofQbnYA8Cz8TkZiyxVuoMwzbmV7VfY74DS1eL
ITa0h7fnZ6+yN0R++tr7BppY21MwhnbbExteWe718idmwgquWTIIDfDyuLHtgi8/U+LYXIEraU7r
cXV9sv5jWbrBl53LvV7h/36bgjaZOz4vDHXZG2ZTcuCjIQvwS9tJ+zDFNl1kEL1neMrQpsIS5Pta
Xmbp1v9oMpL8hUWaApa4vzwe9G6Cwui0mZ652PDNdGWBR6Jvm5U0Ra+iG4fuzo94MRCOgHGDz/9g
RhmvGcc6dHcXHmygKm2KHitWC+P4SfiBwF3+nlnBtoAEvsXr7EHWVOsBniDuIykzGH9Mjq3vTwRq
gO/vVeSxBLV9BeBxUKe6DYFmAuapxF/Se5GVT3YUEHCtFSYBK2Zv1DS/y42TtaLegDnOMrUf8l0a
MgdJyDvaOV7dfc3QImx+2ng85ccE01OMToUHB5JzR2/Z3FU/P9ljrTw/U77oBVXTk3IT1lTzPPUM
tVWp3Y4E+3yXUypHbdhyb5SXGTSxvNXFklb85c2U9UqAEyzonHQMEvGJEwlDwUXHx9zP1CMx+zbx
52vHaTLoQum0VFn14RguWjWgtgLsEA8N156jsH92M3c8+uWmZdyyF6zNmh56FSj4Z9eONejM7hd0
nJbs8GfoiaIOcCOaS6TfOJozKXZrLmE6sOEusTF+7W/MDxdGhMgczTRtxUT69me1L1G9KIZhCxST
zGPBdhFatRhB8OesI6Ggo//7UHcGA5j3FLPRzTJUxFbwfw6EQLHObywzFo21AP7M4+ddEeR5n5UT
gDLNjaY+wYMt6ne4Hvf2s9EqfQPc4lKmA8nuJ64V4JXwiXYdqDkaTANyhdQsGxndlKG3tpoUthn5
vuo0khU/aVs++SmJXnG+aprNDDeZ2AeTSTPcUtJync04guYl3Qr838pd7jTxwsN1pcGyJIk8ZCZE
Ze0ZIPboVMYOO4MZrZN9132CUb77PqShk2wcN0tS7M5FNYCDFmpGEOQdWklikUT4dMeVTAM6DJEw
0gGPSTsOyZ+z4AMf2u5G0xcZIWwa23sb27Ov3lWpcNrqM/CYNBwSeK57t74MSfPTkH1qWurNVsPt
ThZdfhgV/uh2mn9TmMK2++53JmhJew9PvfiU2rSBnhgBvXdDtOlDQwACX8ndeUVXHjDfC5erfIAK
dzRTDWOZAhCh0+1SX9gniltDgbWHN12qf/T1/n7uymmGkaIxtscVf6aFMZI8gC+/rUghNurRabdC
S0dqdKGXG+jrIaCXkn7MnNZmKpMt9XB8CDEpxVrYy+e8agpj3a5lDv685F3ttzyoL/HCgfp9ydtk
Oql+fyMD7Dg2CBpcn17/+Ifw6uPS+NFazf0nKqjM19LfRcLLhkFNHRa7ExL4FJyqlRME2utdrgYT
MJH5ohUwYKweS9KvoDAwCQ+T2Pb+4oH71we4UOSeOeGU6QVXmogZE6idNP4s8SsEa9slbGuWzBnT
2LgC0RKWq9UuEBCN2ZsTnkDe8+tp6A2BYXbkoghZDBQFtyDp6QG5y7bcUV8cmW2FsQItSmfNPVIw
GRdbcQvTX/aImKJ14kzZS8ajGJjZsRnxhT8Q0/E153fwK3BGqMjhGvanGntswuKBmIMLab4oHazc
zagkAG5sz5cpLAZOhObegPKtCH97M2Kq7642gjn6neWLhb3ei07mLM621uUGRGhNLADJ+8u0Cd2t
GXcHHh6OOcEbCj0/XjERkR5JCfAFBDNnPmDkYu1j/u0Cw2AacJ+dKEWxOffZ4BXYaKx7jZ36f6iD
oH1aQAiD8BzE9ft3jCoBmaX7PMtmeh9SVkZRxxQ5C563tFSkQxrvIUHBfVsJOBRbLAZv2/qayVr1
EsYszWg1kCJaMRAZFFI5D/7Fl2beV4Co1+Wc3rUXuPXsU9yM8cmxkwePd6tANS/rbki/AJngauMW
LZMN9KpahAusmDhw1Zh3g3W8oyiEUpFbF8tb9fF5loThoqIPAxI19pGusfptdPJNIrn9VXZBsuMX
G0nKKNji9C67oNxQZU+rTq1bmfnDRrssdTJZQPJy1+aZZJOYK4geHT/9soKaS+MRCc9DVuh2QSpf
c0ETblRaluvwEhrNMm8kQiL4EXv7uKuWq+Ew/HoOsvA1gdFQw+RnJNENWADkdTimLZtrynfa1fTT
d/2ijeDdfAQXQH0SrRYbYEFnLNMVLwWKaI5SRTxKsoTgU78P/IodEnc9imVUMy3vHjaPbtIKmMTG
SkI+mUajLyJw+S2P3RB/dxxNrZY9G5Vhz+zO776jfF4d4iwqv55M/nKkPoXE577uYQc3tA7ahQIf
JQ1HxTwSi/oqxQ7gvlri9vOuWDYOtKMYcNC94scvVEmJ/yc4GTQ35xltRZvCjLY2Xku8P5/oeZW3
dYety1Zd8NRhtVdcX8G1+gq7pb14FhHSg5FxEW/jaroML/PLv1asyQ+SpdQxflJzLZxu1trk4Iu0
luPpKpl2e4SPBJe36hjLzckGu4guAFDBK9/HJybHcPK4XC1pno7ai/0516gYIqZgiBtxhImje4c6
d9sI4wxMPQOZRee+3Iy35x13WcebzksvT9Uh16gt4XmySQh4ODVtX+0o1I47bMWET/QcpQFITwci
OcC6AEKCHTYdnVwcVhgr9RaSPQoIg52zjXlXtI7ZmYYCpf/Td0mYFb/VGdtsK9JR8JExDn1ixotb
3p2C98dVh0yQazE0sxv1X5F+SCGOzjOMMLAFPKUZVvSwELAn2lh8R4T5YsMR7inO7EtVy69y402m
x7KEQm07ugstBr/Xim+yQY+nMjZw8y1x3M9BleuqVmwNIeXKx0bp+aadK+c3wSRSn5V7hZBz1Wrh
zLI/U4swuoFXSzF/livQjBJSmleGxTG3YYsLpJS3BUY/VnwTHOL/mXwCPozvto+4VdxbaAAXDtHI
KbERtqW0lLkiX9e4WRf18UuT76Gl+1Qy68z1noW5LV6KZ8YLJebXWXDjgppls1TcgihAGc6sTipj
SSpuGccY274nujsnhpeKgTDUEpHaSw08aCCKA5NH8RV6IEKJFC8ZJDlm12A29YfutDbthmDuuKc6
HyDL8XCTg5IJDwLoJ3nRuCvU9k2kaemdooE3SXhEMtaA/Tx9JBeraV5jqcfou67ni5qOMjWXehU9
5ixHhjv7yHYA7EIZNjxUXaJ5GLD3Uf9u4Jk0ALIQ8lKvBJaiOoMdhKjEZ2eWLT3E2MycEKvK2tdv
ay9J6DrO65oi2gCEzxHFZ+IlCldLweZJlSRog1otXXk5fNVxecFVGTXGmhLMI9KGxlrXmV72VcSk
q6ghamNMIW8yxcee05KDIG+n4DgWqKwBlK+PbxqEWYLtCtcvYlSxCXaSLiJozp7aZ3dfO1P3qgjS
VjNRebXN1PqNyOtuIg0KwoUR5Xz32+hwFwraLV3VeqJ9QNMwbjsSfmwyOH0mRP5Lf/SwTPSEpZhO
zcK8UbGmzbAondCXA6Gt49y7/HiVg38zZYPsExbhXNr3KW3v86zw/qYJ1hd/fYZztr6AW5TU/wdU
2MEdZAEQwcW37+iPJdOuRnm+kRI9GTkM4/UpRIxbk8PgtqALq7d5tZXATv3A70GEtfQ8ptq9JSIj
6UAddjHfSpSWroqmbhmH5esoLjn2visoEbtRKgO3cv90Odyr6zq03erBXn84qySaGgV50aNeE5PZ
eqzF+1kdp2/xneezXAYCcjknEF0mPvHjR9JH8PZW/hvXuPUuR1JUteCWlyJyy66hFf36Z8aPEIFB
2/Xs+xbCSAliAXSii5fveNfNz3crjKBX1tzmkf99bk2TChXTACrMF6/z0dTudyyGerymnctDNVow
Ua1kOASY5ShQlmHWP3pcojoTlL9GG6huv3STE9meC5yd6Tm39hq9SMlaZByl3p35/5kWYaQaaYLq
J1YBtL8DzItcaGPWwyZipd36lDeKSstWirqscTUpCZGnrdHZVm3ASUd4ktuAqXqXqLckHwvw6Sf4
C27i4x9TDHa0s4TBxaQVfXTTHFhXbMujhimSjhUSDfKj37zMzVFZDwzZFpRYJP3/vlH4f1YnTlTM
eojuHf8jyUuYDE5vGleCBXLVNeuZzFTyS2lgmA55HgKHviiVybKo3X5+Wzm3f5f5VGTlgJ1rSWUJ
59f2kgq8awZlA5BLsZlFiWq+NuD8EbnwDELlDJZuF2prWP9qlF+Le+lYWl9SkhXpTJZ8hAQRlS6H
EPfUpwCG73lNECS3b1nRigMeds/7i3TWnQdN5jbXTY0yrz/KhhwaIgpxvv3g5l66rVkBvWW2GEmR
80/gDdpbYjaEeZ43UAHvJ5phJcG1oIgjmkjv/JazJM/viEg5jAxcl5W9u7+2KoSc01Rhfcadff82
05DY8yzb945sZe3uprjFcJj6t/XSk4cSk4Ou8UAImjE4mgPmnE+bLfvjWs2/a2AqkONvlLjO9Jer
XmEMWTI3XvkwfI5Y9L/v/VKxOyGLZzuNMaE80tAKFhdI2bxrLia7llB9ddxvPwmy/TeXXMDcRn9u
BxiE0fnlS3F/PkvN2C4u2Qnya32uXNTRBvX50X0KmgK4GYlGT/F3MTz47xIEktEl8qUcBgCFSy7W
cMVAVpGBhHbow1cU4/b3A1RQ1fJb/C/4TWNDdC8DXbOU37KhrMB7esH3v3EL8q/LLomTwXwe/LIc
lwl7nTo0Tc06pnC9Ao+GFvWW0vcljJeLO2Km/uatIcm9TwV8TlQ23nacMxzfQryCrRUbm5o1GY/A
0HBdBH57y0feKPUL1rwRsuQMtE/1RfZzTlBRNSJlZgZiIZiES7+3lOl0O0ogQohDphTp3StjX/Cw
DrYeRQ1QXHvlmHoFsTsRNZR0eV/eui2VMJwA4D4HJXpbkX9SDMKo9YA7dKMc3//i8eeI6RWnI7gC
pGSTXKpDrHvplrMfIxOEtPzYaASzsGWAcnkJunXNl+9nKBOf1g1c1EINreDHq/luq3H0sUzKJigY
z29mnw8DS5Hq6j2FOedlAgO6s/XIfp9UTzVSffUJ9Xtc9mcP+0qDjsweZo9kuFl1d4n9GetM7iyj
0l5WVsyAOh1I07uEFYpHJumULSuRUlXfKvTZdatf6x9a1Z7fpUW6yXttQbyDK2Y2XgcCAT3NaVFY
v+aw9tdAMSu5KzZ3o4xkfY9p4eTa77oza/PWe9pQl90n63fsOdlAQIyi0EZwbZv2UHaxjCaRKPoP
e54Jeydvb1jt0HatxxWqw2kEEA7bZMgrU0D7IzE+ueSv0x3EPCLUfVkSSIKR2PQJG8Nhida2o6nQ
TTVi+aTsKra4y2VXF1ExfqsEUTQhKz3gv7e+Cza298hbSj3ZqWOXyMm2GPRrlhMGEZgxDtDgb4+q
LrCs0Sb2C0kktcm6vbFuRnvoDqWWDLMfj+B0lV34/vpbiDns8HZs6SfukexHLlEGUGlaRqpo0VpG
QAw+rJZdW+HyMalm0IXiDvtTBmhwXkhGPEuyBNtcGS586I/9Tbtwp/d3VxNxXt2iC9/1i6/jOYuR
cO2tBl1i35djNwVx/QBuBbPRg9LeJUd7t/tLrfnxrnp+PxlrCYjU0NeMy7z+raukA0iIwvxvnpf7
56JQ0LfraaRdR4LmWnxZiOUiEauFeUIRSM7cnMlYxDFzI15E+4zIr8dH6livGXkuZCyQpvVsNJyP
+mVUPTzfKN9fQ72oIZ2ajjFJ+0l9Zv8JFwKiahhsLkaqDMWcMQmzZxXTPqlIXXp2yjkxu+9ysgww
g22UPcsGyl4GJTk0lavoJwj30LBOgCoMTnWzvJjp1ECS1S9QDBayDNavC2K4tTsn6Ak7141Ti8V1
DtShdrrCtocqPdgvwfXg7TdyfwNGtDNpQ/WMTxj80CBvfjz+hZbhr/YAx5D7A5z5s3UF7fGgQyux
wCRxvh5OHhaaUcE4LoNxgWi0mm3jkExHEBcGFKaWz9P7E9rf3Z2MpHVH/N3JEZHLWbcxHBV+KtHt
ETo9AweZ+tgKtr1m8vxfDGoyEtX23LcEbYTa60nddwRhZhMjX1k3IPNBoF6qqaFvR6lmLM9d9OnP
OKxq4vN7vUoB3ncvDLi3pPExt/QLoSoKdf+cQ5+17Kz1Ha3BEfYOGBxmAl4ALzWXA+yN0IB5+RgZ
XvfwukJdm0ALjp92cK84akkUMm1K+Bi6avibK1w0SR6dQ2R3NImuWMU6pMK1ziFfAxv9/Mtddddk
dp5FNu5oOx0eSggvVTCd1WY53m7O43LQTtFFQO4Y73QnMjFn5ym5g07ukVIiZYg1Q+t6SjYjrtEa
+cwVSePBPaxsm7zakh7W2oCufAH9UgD2UupyyLzJEDYDwXyQjbpWtlUAxOpkb7intkDKIuIvW8Fl
RKJkRhYW6MD76Ut8pqeppQyqDDGGVXYOe7YGiEc7GQhNcO6msI2K7dWkl6aCvAR4qxB/V8ryqq96
msFcJEsRHGqpDpBGxpwyeQTKXPdr0Jdfw0ubKWo8RhdP4+xY/EgI2QKIRaP/CyoR2jCOutEXF2vZ
4Nbynf14yGmqLbjasMyylMx46GrdiTilb6jLb8ULfva3lpcPWm3X658+CtyLOb52Tdo16OHKJVpI
tswcXG97Vf8mHQhwjdRIuMZTWztoPQBVOHoLKEhsGW6gsNaKJtS61xuJClqrOiNiLqCtdP0W6MPi
9wL9hnZs53T04u1fF0QHhMKuBfiectnVhm8Sgf9BVwg/s7kTUJhBasDonnNO7yT8cVr8AQMYXJOj
21ZcZ3iCF3YlcwY9r5JKUbvCxMenzY6aYv2uXbqnhkxYIvjTSkwvlmAEqXmUe+3t92xL9GfhCQGp
ibkfis2j84Ze8Zv9tmhd205OiCc4l9t3Y6rSPdtSEdi2yXfqpxQ7s5fBD8zWMEUYSN3EOlnIgm7d
UpclmzFcuIErjV3uxADS66mtFUoEYvTr4M23KvK5TlAxnQ5OlrwDxZln1NnYryllFfP4JEvUHy+0
NBxMYujUaozJcF0wIH/8QMrzzZsq+jPX1VVEC1jvauDpXWhhfGEjuDLjRzyWw0lqGoPLbTejvX14
jx+Dr0wAQFqJV+QTPFuX3zMBNjFu+pskxpyFApM0KKiUTtFIJ5hDczkyeD/4ym32PSGfCgY8vUVO
yl9rOKryEZbDsMD/5VGHQ9oo5bAlnsE10ko27JFVL7mXuRiUp4cd1DIVMVqrSIMfTXsnUcORGARr
9z7ATVWhd4ehRo2UgCo2biC2fckcEQOy4jMU8azj/f/mSiOv3mUpD4IrD46FzQ7yPZlL9Dgzx6jC
vbQ5MTCApVUkV5tCQXWvbLad5i/TYjrb4tJT7JV7mQ+EhQ4cFWqTrRkIHZVoDW/waUi09tmKGNWX
H2VeJiNgF14hKXYrthcW1e83OEVsKUBbpp+naTnNIdMc5+nXvK5HOqlF5NBNMK4SPTVqp0IV03gt
dUvDAzCk3gZWl2vC0to1ftdwh0+wdgEojmDsoSnC5/xNTHaB0YYH2PkV89MFPOjlaAVlMA57mDyO
DUBKXzdCBfdQuVv8d2lt/sYqfPUhfv9eXCyQ9tvXN6h1oTJvjCUiLRqnxBTZCaCo6GjQHs7w1koB
xzEUR+Fv3kK8mNet+PY3CmvEpXOfTtvmJmj8ORSI+u+tmqUfSBAFMA2GeQhtYeC7Vt3v8x3Rrw0x
h74/OA37knqlPmPxPsh4p5UuUX10rhNAbeKuyNL/anx37h6FkKEP9RH4zwCrUo2DuTdTSOCxq/YY
haMugH/bdcRCaTcaSSRguKoJnxUhX1smZXM9gUIUlTKTa5+gS9ka0mwbrKNOCpQko2Io1TWnw/3T
9Bfoef8pcLXRulpysJHVxLiD0jjCirEZ3yr4T5/nl+OcRGQ8bLN/b5tmQlYdfwHBwziv84IL6y7q
A9KnOn6zQbPGYj8pFvenVBtGHCj9uYtCvRuMF98uKh4q9LE08R7zToUt3UAm8Bu9pChlGF8NdYA/
BeGsdr5Vmq4liIViyZhoCYkRs01yPOW6Clf2WGle4/7Ru+C/fXAnNh0vqFUWGFTGCLq+TkO48Gtu
vEjM1xnbTneGeyXd/zPNaqWc5o0cFhT6/OgqSwV4p4c72mAtK7ual+9aIfobM5sVYc4dXvPb8LE8
bGM9WtpvbgLreZZ13OwstZl2Wf+3CMogU51LPrEGwxOTYmUyoEJYAoq9JUTV+OHsFnaZ3KbCmDvs
1vgvq/0BugFnUHZPYgdS84EKh/w48lZ6NdmsNmVLEBpvrNoDglWC2TF/eJeABpsHe45UEWwMdGLP
mQ01R+ZWpT9A5LAbjvvCVetQaEToJVuT+GYS30heKpJ33wfPmRDHUEH7Zn21iGzEhjT+DdtcjMFo
5JqkxeEGWhy73DtZntZh6oJc/39SENehWkL4ndXoLDtu9qmNKuYFyO6jAtMnGzDwQG4fTMSxGf9K
7/uyW/Ux+zy9wQXIXcl/6rkNcZCK24b6WfIXGX1kPT06vbCqW+5lvMtpfxC1DMzxyBJWFb59IsBM
iSPErQu8LWBEJ1Y/Y8HK09xw6p5QojEN9EEzjEyOa5Pn6iXJnldmLNyzcR1MRqBgeRDyy1/Wh6M8
UE+MNa3RDxIaRC8L2egJjw9wV0v6nRCJOpGl2qHA6DhIK/lmesOGs0Ejja1BlHjoeRia9hh+SVOK
4U4twL8J7FyVx5tBmPs1Ok8nVrm8+9SjmsePbYDC5OWkU9eW5D0nG/y8y67LO+tpAOgTHZzRW0kb
0VYP7EL1ofrx6WF2eBHWdGmQGiVZFt0qz6IQaWD+N5uyNmOgk/6qfVXecaxmTt1ufUpda82xlgbu
fnrdJRsNJSrityWL2zRXgmTuigDALgRfsrJsS35Xt+W/gmuVGlKUZujUkj/p6fKIrSX0k9yf3OrF
Eq7XE/VPG21R+hSA2Si8GzJDU25L17BGoxx16EN7Jy99CKuAuwugN0Ds+BuIPPlFhtWqtsM7SyAS
8WHUmZnmchYpLTS+BhrT5lwC3L2LgX8x9Q9KFQQFVIAOIQvmLuDB9xgk/OZKuoHiagNLSq3nF0k5
D1+KaySX/HGQDeh06giAtWQX4CQUViz2uqrvGISnUjVZI3MVX6nzgGzaHIAg+9uJvcsbUDF4ApfP
hed8iNUE98vbYvLEluus3gwAQf5oAYlW0PTKgIfmQIu73gu53eWtrT70GkQqlO/jL9Z0Ll2QfuZx
IE1eih8UpS1MWYvgslw3Ee5wkZTo7SVwrUaWzXoJWakkmrYdh19IddHA173AKtOOC7FPmXawpzwN
n5om/lOccDk2RyX0QbzkgwgPNY1puX70Wm0mfmOcWSX5BLtqiF0VJWIJ1eSuhznEIRv2U0/ow3OP
zOSUBqgElrNhsqmKaUDFXF7nTUAuTMwVx7v7vCXls7/PsbdP5rH+8Oym1Vm071xZ91LLzZ+vaXxs
DVvAFdaFMmry/QLYkaox9XJwBqa/5LnD/ynC/Zj4vX2VOCqrN6O8NWuQZEkjjutQmJGWqL1OX7Yg
6tdyKYAAcsvK4kpwzzzzZkT9tHYmpK4EardlCQuMrhxM3kw1xpczhsMsl7gqsOpBGMqQy9x3OloE
bnPJLXxXqhQY9MZy4GslEkZNPhiAPXzLzepXiY7Wi999eXAYaDI68wPTs7ozvjRRNs189Ol63w48
OnfBQtbn4Z9Ej0wV57FrBH148HAIys8vEZyVBcbL5NemY6qz/SQO7mudXPuFRr14Ks6aI2tm5Tt6
fyoejzg48GIUEdWMRcW8eKSLck0EQ2QL70fkYIgHKUkzv5A0qw9rTwWYRlZMJxnsw1L20ofgGBCU
O0yawjk67HHxCDOK5olHOVY51x5akbMdAL/KDFoplDQZ9P9AUfAOMDn0/X3S5whGHECwXpcUu7xT
M28hgRNJ7T3J9C0qXG09tncaxIiF41yd72n5BVR0XCqXpujjLJ+HvACSn5hgNg16h5lX+q6sf6oM
tBi81VNnAMf7yoEOi9SowOlUxVd5KzlFVWd41y83unhNs31bRfh5+dubG+W4lPPsjtgLofe/XFTk
EF4YYkNZxBJXtmeXvVzq7vkic0/+e5SrFItvOCzYMd0K50h2Tot7hBBbgkxesCMj4ZJfYPOdImAK
xRBh5Ou3kgyJFRaCFssmYExpWjHmwUL0PfdZXZC+hubMzfvWe8eoH70p6rPj2XlP/e0JC5qtiqOs
ustuUTFFwZivnoPoRUWy/eQV4qmSyllpPrigTdK/81hjl1H5tINnIJm9V42U4x0+9o4O5cfDAXly
dJQ2eB3L431V4QDtPv2k9z6i8z50/uy2wLva3Kawjuw2iRnrMJQjA9ZpL7BmkI1GiektoI9mY7Bx
d6IOMnGyQR8bUgLyJjlWTNk8OfvXa9kUWdMnNPdQpCyWy2Zdbw2u4WoBWj5rimUU2A/NUIDyTmkX
HHlwu+qR+AJ6tiZzElonoDPpCjmar034r0Vgw4rrDAL2CrlIPyyAO/xtYIxpfVdKBLS0Ew3YFMB4
trx7tK2c/cjved87YSZrPrQ7sJedVQkFBa1NWPZpo78puNN29JGfe8AWKCdi2pqeHYxvBJPEJUPI
wa1natoFv+yUwFiVXVZEpwQb1ybkzuXW009NYSCIoUdceWCk5XFkK2DHWRMV2nEU42S8D95uzsJY
wDdhA8QwQX8VMNcQYewYwW8YliY1sNib+Ke4o8kSCuMSXmfhNz04TPo/0EsFuUBiCUrTvbO3cXbJ
UcqqgBNhWVpc7TrTjb0mJjUejQNFrZlZ+CrQk7sdHXWlTFlnDaSSbMSBKDt1bL0kWouVeMxegtU1
Jo15GqVF74f9go1+pvb+bbwaBVpPNMmMPNYYJOPO4ymgtQD3roJ6+b5rDtAzSUN7FCWUIJOXVFuV
e3E1VZ/DKIQaA6DByS8mPdl7IrhJeHWjc2PjD6Pfl5qUeij83Q7YwFa72EMoQ9Wq9S71HtFGFAvw
Aq/wpJ2yTu1IeCJ3Y4TlwvDO79yhXZTeXlhCxfOl4zYV0FuzWpSfrr6/91GyD9OAJb6TiR8QryXL
za1MIh4ka/86lCRWWBFAyO5LkQ0GIviDoI+vHhrVE+ToWO751rBD8JZ5NUPxrJHA/++IV1fD7/Qb
4ypFJ9hxVMu9TtUqkRIGkm4VM+kRTH0+rCgkMjLRfFqy7D7gGL9ZZnRZEhcCTelAObbXwpUdKzhH
on904UGaEHWebHHvGN+v6oPAaSBmBFKHltuI2kresPTil2HRhg0MqhXfD/LA7Z1srqafZT/oG1Z0
yCVYSI+QU/hhWcqj1ieD1GktxiJF82TYmXPy+oJ7L+uBzVNHRAAw74b1N1OKn0Q8x7I8LQv7XSxd
FHPqypnrDPjNEEUHuAdE2a7Tlbync4bMfTwqHcK0Us7fKyqHGM4SjVXuwLOLYBXIwjTv2wmBqB8w
LqWS+EQ0X9t1bMv4Rq8m3cN8bJ/j3dbQ0Zlt2cRvcl+sP0evRvMN/dgqhCIu3qaRd5jm25V8W1Fp
v4tCyZ7KawhHj6aosCeDCKvGcHKXVMgufwkdXwqvEpSUc0MtJkxkRtHF9un51rrAjZdPAfo1iJ1Y
vCCLyXC6AHzMj+nWgidbF6PNnDo48t/qyH0Pw2YyNV1LnNc0loO8d0nCLydNv+4KakfZXHs5wyXt
pno9ktgdlsU9EfwbZiYYIF3fTxFoeiZWc1ibjJBom9cM09ZyCa+VDVVTolzLVzmkPEQ5KV1obyPC
7jW4JaPCFQypIKw2cxa1+jKwRh0dFJN/KLYn4swz2JDbTwS8zHPq192WG/lsCdtiaUcsQJIykEEb
92G6R6MNeBzcKNfixyjnlMOX7fe2xC+6R9++G3LJ6cUZNdvHpf/C39XM3PCkw4huhiTKj/8cG66M
QC9Ow38IICKhWKuSdLo7VZF8aPs6w8asaG+F/7ifIlqdmQqwK4Y2Tf3OUIj+PXguayaz7QHKnQQP
UoI/cESQBaV5IbP4sFVpL9DoWMP7WS3yUpowR5AlWdEeCdX5HyAVmNme6LlGmySMla1hFqp9LB01
JAZ6f6Fg/GD0WvME/k3mRlMVRHhDMDUflJbs3MBaLhSCJdnTepxZhOfYoMsLGeiqDmr/CvMkJn8D
jcm7aDMIUZAwCgX5va8Vws9+r+BUnl27ew3DO+rK5zScQeiAXO/jRmbcYgu67wJdXci8IcHMTOsM
yg2xztxSvpVGdgDHq4wNBIudhGOFyhzIzCamY0YcRZjCL/H/D/UdS/KwtT9EwEvV2C56YDEUZUFO
GuesvyzYl/dajwYoaS2Cang7vFf8jr8fRcaVU+eRJwO9OxuvBpGgnRoq2geOaUj27C7sOn7lTMbi
b8KXH5m1WTkpAmKi1hxaZZalpgUshNovNzzTANWTB2SL2jk2Rq3L8RlsKdbx+KWsiB7sci0TVFiu
nG5UbUulB5M/op1aj7VXSd/OdTTXHV9x9t240deWGMGV3Nhzb8vtiLFna9XC8F8lyymJQ3CwVS+M
zDGOoDr1gKYINemr6Qy+GnDVS7Q29bfe2lXYJ+R9E3Gvo9a69YdacrDiAi2p0bJjnIhnBdWJuHnH
6K1yQW7b87ff3Raxx9A0UygtKe+0HrikKAwZBhTwS3Bd/bP5KsWH1CjyIt3IZt051YMjCSupzbh1
DOIniiPx6ehxYnhu21E6oez2dsYGMzhtXgAnOtE+W5GfhtEKL2RT9SSa7J/brB808O7TrnnhwKom
p4IfKgSCeFdF0592PdWlHV86NQFHO7TiGmavOJizMeOXDGlyn6singtuwzqnTBs4/wg/fMyN8taA
K1tOozvzfEfBbYuCbITCfY1lvRtHMPucpMWivgevWO8a0HgDFSlfi1EVp+lcD2YZ8bgywsftDeX+
YetPJd0rwToqmd61/CidHJnosraAOyC88WgsuASJHE//sxTpc3/yobSppd0i5ASPN8627l1WoazP
4nXhkZiH7b6yDBvBYQL0L5bhnzsnoYQcIyJMOFD5FuSOE+fKVYvjOFIkEzQrf7y4czB3fx7d7iIg
W6NFpyVyhccwR3A1S86+vpt0yLQraB2l0zrgo1F7qQKwRSD6IOzm32l64n+GM1Fu3pmafhfL3Csg
dx54tfeElMFkJbJM/mp42CdHi1RWvnsFqIxxT3MBfVx4u4IOXvZOObC9i1ZTZbarX0LHKylM0acd
AGOJ/yuJNV/AefocUA7RH7jvvMqNhrzMQLrd4pM3ofiAj2SsdjR54cFhPxuAJJgLZHrtvSstUMa/
y62atQWvB7Ts5ooL1Jw4I40rlokutql0Kq3n7z35aOnwnbpOXVaefs28LuIDhU3ngL4C2NQHMy33
pxBLwCIM8DiSS1XKlp2oSNWVMKaH3R7F0HotPatwXFfve0Pqg8kN2Kg22lOREPy8oCUbnUxT3yjd
ajxdonW3y2U6jLPlsJ3de17tEU5Roe/O3lX4kgWwS6wJKYlKBwLdeSfjisMlVM2sBoHJ4CmIMZ52
Ewbj7m7yGk2TZdBdQg5XDfY+7t/7C1+mbfNb4auEEyuYT2Nv4xHEnDpFoVhDEyRcHteou/ROAmH6
hOcirlLtRuY+vcDDBFH5wviRbexWzBd5wWEmbCQtv6X3HIIyP/DfoCl41sYliITvLjz/5Oo/yqph
xxrjBn0eX9wIltIuVAp0gahZw8jQNefpKNMtWVhkTOmSS/RZlSDj1MpBFJAK7RPZdDIhBCjxL1xs
HvaiRnFN9sFbSj3QhqxxhujBCfgcETJWgHmui/Na/rzT0SnAzwbS9jFCIy8Gmey3+RkLZEeF7DLm
FEeZmSAqBerekweKt7SuPfAI2ZuBBDVf1tqyISk/VcEvIMaBuARcSQ9rsY9iAwLLc9/ROcWiUwAR
6ig0h/LM1l3dlwUn18OM7A7IRuu0xYbZYyBkipyt+AcjH8nbpNOt4vHtNdUir2HMuOPCQ/7OVfYV
RI+ozO+vBMCs6VkS93LqG59xBgWG75NaM6xReV0zz7/g3gcQFWvkpO/Oe4yVwA4Kau0xjNRY7e7v
/+iln2vLUzloZ4z5J281lN7F4xh0yPlMGPhjvGXNmF1vBgdd/SGRppb3xfuOpp/exHyGIhGXR1Jq
UKNFcxNPEFHc+t/4ka8iHvaK2Y67xikbWGRNH06smxnoB/VT4MTETxGlWiH7tbsDJjs2xCX7griP
ZjU55vVKDlmyoBKhAP8gvYLAOFK7fGjFR2SosS1VR4k2WN2DZHFJJE9NdaJf7onCLKkKq7RsKzPf
FmOMThgb7WoqrnM9hN1sf3ivTBVIPSwl4EGWgyvW4S5zS7bGjeMCHwZIOkGBmkZ/YDhOGLSzwr/R
sxnZSWc6uzM7j5zdObNdbPcI+2htr/OKilHO3sJvja147E2uQHbEBJTFCcpjEyWCgk6wBM2BngYR
Vl4ssm79L9vdnE8IzRUETEZ62RLJQfotjB7vovx39l8f6cNhfYhkvnfs5Pvf/WjvZCPVmz/oDYDX
f03YYVjFNAe63MjmBthSGbDasleqbCH05OrwEOWZeE4i+hfRTkjqG9aHymxB+lonQ2AUaj/MY359
+TDeow+X9IMQZlxD7QBJU0Z67ePKEz+68CAOCcIbGXUtxl3DkLhXsgKa8AR8z/06LkOPpcZkJYd5
MnIKVm7vlsipALahg2lIIkAbr5wDtJsagydG7t8bHAy6nAVU4kSoH6QbjIpSXSTwTyg6yQcYEBp+
b+duTHCAyDfX6a9nXuKaGl1F/i76s+tXgORY6tIQv5GExdOsUsigxlNfREdf5QDFst1MkNT+j7Tb
u8RKjG+cT9cOfNrH3szJOX0+jty8U3CZw5eEfM5gweUEa2VNdyFajciRuw4C5egt7O8jAwfgMLlR
fHdm56i3+W65p0acaBP/dXBTOiStLDW3F4QWwCLkbVGFTCkPbBsyn/90aq75dZ1r0HHBufsVYIp/
VD9nx8FV+0/5aCvgxMC3ZAOwcy26oSoK0+2c86iNerHZwsJhGtIISzh06lDf8j42OJ6FAiOFjl3/
OvK5kT4PPaP5bGJOIEVz9EY+x/ci3+sGVU/MuK2ctR795wl6t/HcoS8AXNPICnOR7l0OICiDIkyp
0OwSPEZMU8YkTS4DvcGL8UsFaY8hE0fgetb2nEpJTo/Q17Lt8NkOl6lO9aLikMwGsuL6iV2RmOoa
D14rNIxYAUQDLcstPVqtyVTJfCqRYrU1mJSVbacAh49B7xGh7RZC2e3CFLCNiu+yfO6zlKEI/LIz
HEMYWqY4T6TUfbh9puEeQcONrHwUEQAh8kdZ/nkc8k6VMUJhh70HjMzP90iXzGj/4SoT5Xa+5VeN
RrvyWDEK92JFUbVTufE6/QfBoGXmJO62JTmAYRVfz9CzGihzjmmvg7PSh8AUTqfnRSIeuiNmsOj2
hCSyeU3xFnJzZ+wrcoSl3CCMD0DC4RzaEWFyZmAl/obPnD7CQ6yzCzTJIEpIS1sd1MmE7QZN6k2+
zRsa2sXEuUFD/lwykwhxHzJQz9e9LHNvoh3d7THaZqQXgvQstQIU1+CkNK+UBzjBs2wvlAFVLIJj
CgdC54SybmECrTjd7X/1wNZHtwrpmfcxL9utsuLqsEyRexTQFs7a2xbMBwLduG6mSqMQizcdXDGE
kxcUnkbt6xdo4Ppj8/wDefqInTn67VIanULW7pxuEp62IEfs+sPov9g/k8lYnr0SoCLoEPf2lvlJ
tGe4i8NZo+lJ45tF42/ZRFJo49hp82fKaYGhVnPsE8SgQrPxVPHvmZkS6soSEIHXeJPMWmIRPBo7
NcxyRldITvy2lM0R/LNIu8WSRJD+x8BBrBLV44hpyfewm7v9vvrJO8hUhbpEvWUOifzO1UWNoCpf
X3o6wLD59e0dMYfJ5gYPcAmtk309Zt5wcXQT6wvrgDNQO/PAGojFdRTnRmnaRDoQp1cEDdXz5MFF
8Gj3DEgdFZCZM0pFAvzFj/sgIGBmlK8m8GbcQ6j1JZHlWQ/nZg4eQQSdjH5ktZIM/0mgvd6SdglO
PhFVh9ttVulgUAPZ5gkBE0BXl3mtsdVcpj5UR3btefKTF8onJ2NL1/x4Co9uBU/BeoQI0Unq/3uv
GJLOVBqXGf5AmYrW4WuMcx73ZOv3SfkN5Sr971+3LIqJovNO8TKFCb3Ae9bJKWtRe4fe0Hxx8wXk
TvnCCOrwlssYhQn3cGja39+BE2Llx3PXppnbQeCAgk7+BZLuB9Hx+37/witPVVPwfkN7so3uAe7y
+wgK314oiRbTvf7I//ZHq8Ug5JstoIwy4Z+YMX8c/1EhkH5uq53jif5jxWaP/Fp8AyGwged22+xF
qYlru/MMCmtJ71c81/hLZ++gM7fHp+EC9/KW7t/vZEgM6l7Aw3r0crstt+0CKndDj7xVQtuB5TH8
XuFH0kg1glMsdWgFugyZdP9oypyEzOt57VIvyJUZwtEN/HL+YakCarx+IhQ787kNDIyWvAJXBF88
xEobtyrwricDlwOthMis96Wooyan4fge4ADzR1uXVIjkCpiYQeZLUnQWmfRbXpwg8LQxV6BkcMkO
YxPJOm+OiDi49pHmasVpiwkfG7k87VVPiTNqHtonzZLVBDg6Lp9SdyjjI7dp8pNMlqimLSglGSHu
Qmsj+4SGr3AmuKDLbUnCsXUDSYBqTwhnUb94T5wCpnhMq7NIrHMWIkFk64mDxcCWZ7RQ2h6+MCxC
H7d9OfNTU9wS410EFglI430ByeZDqVppDEOeu5EJvo6MpJxZSab6hi4B3Y6Vcy5riOhO4lXSccfU
PHQ4TBH1v3ExFNm5OU59ePWwz7ntbwq4/X8NsiMQOPlBRlK3n9YjKva40lfOb1l3L/+Eqp+ANXQ0
LH8q4aIXW6wLiAymapRWf8q8/ooqtkXKwy3chRLBZNktomAcLYfsD/oiaQKb90CBrmaxUnfUPBfX
54y6cPBDtwUkt+PvhU8nXFywG0PcLqqUabLD2TN5/VghBIuvWlFi6vYMXdWmC4FFYhPEPS+RvpQA
bBmlxuwwhb/coN6/bDYLRctpm9b2TbgZ/0SJNJasdMBUx8KxSQDmkZ7zfiZJxlq0zk9HuocmBNT/
pdWvkAyPSZW/LLjx+bn3aeUjuYOPeML0J3PFhktxQKqxr69kTs/EaeYsPxhe/iMEzOkmPyqgj8pp
mZUD3Q95qR+l0Gpkmq+voJbu4rtiuOGWd+LynqTZI2cJ7KSBCRbD0EwiKeQXem4YrOTqIqu7GCn8
WHgjcT0EN6DeUZ9KRDwYkhlfHVoeoTl2t+Mzk3i9fWzmfUoyg3afBuWFhV3FzEPT0sgAXVxNG8oq
T65t1xM/eAsGGaQuPP7bX4JyiEypKfYsrd7MYSEvsq5nT3yg1X2YufMpdgJ2kcYZDumggNzWxcg6
g0qdvAasadwMXBX07jxjFkIqpaAAO0R//keEqJkjaZDhv1PiS5fkVKVYb0DxzKtl1gZFwhzgXFk2
D2HCUQA1z1LfIgam7KsuRnRlfrbHkPrP/ocNks/3hM0aW/36BqGnHh40TjSeTP2Vyfs52mKuY1we
66tYZpmAxR3G1UrkokggJYk9/Pg996+rDnvZJFfpya61Q27JSOKRs09QelDGaKPEzRznk6xvMh+M
Y1rIt+SCb0LMzF9z0AlI65hboKnfz4QaNV1Oo7dLIXm8r5yXaorG+IAWp1Ef+B4O48L5QWLwt1Z/
kv5Zb8ApknFubsJW3zRsHdSTqJuZ81z75+6e4TN8JoHGSrXwLYAPdqpdwNZvwQVNoC7lY7HrLQnp
iGlhmBgRk5p9NGIX7VNfpaoIOcdONX1f2Fia/qekpRIDtz8ptqACUSzMMJavoKV6AcUNAcngyOSR
7KHW8/czMnLR/kI5JhzmW2L4pQXWR7q7rRCllxMXkrF1q67XYdMCmQkpLh07LPVxANzdZkBu81pC
6/xn4Chz4gxf8WmRQH5CVFvA5hVIM2X/kCI/aFZbUsKh1s7YPR9OnloDcTudT4jjVrbunBVvCIys
gPg3UmiQ+IFmVEDqiDXzLIgdf5zaaz/iDZjeQVCWCNwRFJ2AV18mqO+7JEA/7Y1MuH+gkPv+9UZ2
GW9utnywwFlS6Vqazha+8dfyd+4CDocxHq+nRfJrWXQocsPRP5BKavoiWeSRfRRuG/jA7Wgukdgx
CRwOcfcfhVS5mwzrTG9f3acViEp/V+SoryZlSsjv9FHD+YyD8M8YFTp4xgxlFPXBnxajYhNilGx0
OuoKSHZ8SeoSNZG/qyaQqpzJ3pIhohsjnOiqeoxsorsnWjAPBktIarxILsCGIWB7ptdK7t1egxGD
+fbd05Ss5UM56iSfDUn7PLmhzSGVGhkKowdUxBfnXDQduOZ9Ydcb63Fy7P8RIKzYxbIWrJsVKuNV
D9FbQTzi7Z5fC51gvs8Vi4gnvlY+eYApoQxn0rsZNZnu6X0D7gbO+A3fkfdHitM/VrNwUj8J9jv0
e3MlPis3Lmj8aodGXiaLCmQ3mpB6T37FELTxShb53FSpkfq5gWc7APqjDXps+ifWQ5ohtYMwaNi7
AZ07EhJpo+jD7u8jJK3U6M8OCuD6C5hUdhlSyCsAsNf3MqooLlF7gE6LR15IjsbZhguGnS7FVqtB
0ITqh3P2OS/fAL2mUHg9WflTm7oIX/YQSTpO/SR7d1SSZMvUbqtQKOx5SZjdOnFxTP2gcqklAEoV
EaE7M0aBBJhmCcCCvLyceM+qBFPjC9OVrRrW+bYzrOYPX608X+wT73ZIROUCNeoOByq30d8YEhCz
9UaAR5fZlHLPWUSGNJwzT3CwxSOvLsnM3O6CXXkFjddJFZiC/d0bP9TtyIvB9S7LyQwWaLRFvmQK
A0Txsd24xkdp+AzuvbVLkjrjz2tY+Hvu3xYFNKbkA0NWtxOvyFfjQPaICKkwDmCVKo1R9F1DE4KF
KmeEpHtlFABLs4WK4odKMYgN9tfo0w74XWUL/+nKVYSAUPe9bgTRXO/wCanLwZLR+cY3JgvUfZ0h
J7lFEbB1t1CnO7oxE50vh2XBWw0c60shF6PcpeCTqwONL8J/tpiVuua+KTJWef2RvSTDXWcoLBSz
LtRuzsMRKIyzq1X3kYALqVBW6WV8lE4a7mF6FvOkFqi0DZiAMO2Z7NE+LoAmfgzpFuKnHZ7O4Uhl
TXB0MYbitLEJW4b76v/vwpEiSpRi+PjVa0szTFEF8nNzOVKNIM5BAPtES0j8gVkkDn3sMSSmoee3
SWXZukL+4S4qGJKe1uqe3N+4qPf1aRR0W5qI97xztemCR2pCsFm/WkNymdnj2W6sDEKJTLqdAKkk
xs6N1FJIyDVwHtRswFljZmW/OywAKC4S8WWA1CdWQqDoWWkssJaaA2gWw2DxOcQ2R9KZKX+QKKEX
oHzY0giItjaOwmR5J5zwL8UWb5JA977rr9PFDn5200zhVz7io3jMc4qGHEQfQ6T8jjeoTZKmzj4G
B4xk0IieiDnLlkoSmyPijfFgvRsq9/79cMge4UnOIdrlsROLYyO+l2xml0fhOEDbHQsKQs2wdPQm
S2PxyFRagpFziZCUVOPNlE3hjmnOGFnB+VP9JZXpQg3CSyEiE0yns7ZFLj2yb07PALCFRpfgasyW
hx5DZMTzDmOCEuKzbLVjJ6q2m/QTdICwfiRv2ymNAHwg9NHhcIE32hLyh9LoG/RjMFRcJZyttmAg
DypH2ov3ZKql9m8gg6uiKk4Op8CWV8qJL7Pl+N1CQU8ZXjQL7aiczGDJW9LBQDkomKmC7u3CYjVY
mulMI7S4G/AmPeRJV8ANtV8gZatt3rjsMxAelzsjMHBj2dMGho/xYRm2AQV1MtNKXC87GwkMsGQt
GHV4C/OgmdwsuAYUjTU6sypvKMkAWmyiLlV00yXK8F5fEP7htaPAIsIjCTMCwnNZO5zATicGRMcm
UAIvi9GVgM9DUQgkl9jZ+438xN39JOb3G4GEIPp+m8Vz+OvOWcZGLEE9RPqlD44YYacwYh9zADAz
rBTw0ysSq5iAo3jVQyMxvL1cXihIzj2Sd1mk/CsNN71YJ2oteP6+gkMRuVlHKbe6q2ZXXhKeT0Ym
rvPbGfGOjRMN1WE8cC+AlNeVd1LjR+hjBE8BLHMXFvllZsmBvedUMNcNjuY3CthrG6sBC5DvMJq9
qHgttR4WLfG2RSLopuaNQT9EKjTRvbj8/Iz3RYOetkUTZ243L1C0YVwJDFrMuS5TS6ipPFDF2yMo
LDLdaExxrM+Y6wtpZsD5bhdxZwhm9kDH5EjpT3pm6DGQE/Ii7l4M4Cx1DIb509t3+E7AMV/5X1t2
2AA4YsNE/0b76H4QJLjUy5rPzzHpLLVPPIzYySjWogLeNcdiPMEj9ceVOjb6riXZKwLpLER1uR78
mYpqJczkA4Kn9TAi1Rtvj/AM+1qgLSvumvuC6scPbLcBojzFLDhEtvBxlEIMOSeH/vYM5MIHmjme
+otFK2IwQEYlq56zDsDaxdWeNpM0sT8gO3/gf1XZM3gm+KLGoMsjx/Ij48KxpHYaWilRD3jJi3Ue
rlwInAK9WUiHdTfY7VKxIqkfcRjBqbZMb9z1sdRoFgecrSBpotNrecYCe5kqLFlOt464olPXcWtY
x5IdmGqE7J/wQ1SeKsqpgMHervvmAV6i7VjJnYn9rwW9RIgnAj5uHpmT9jDhh9I5o3YigoiDc79N
lgZ7foEMs7rfvnOv7vphUuCThdbVk7s6YfLz4vvqe6qkcyptiKxJ/MGEs2oSm5NJZbbNQn8yAND5
N61fYCyf+/lyqjNCP5amt2wMz1mYueyyfP7Cm+MbFhEWiwe4xymfCyGyqnELSOJTK6BgiJUd9peQ
lbXOPsIBREIdTBoU6QY0NihOfpR+w4jpdVe9BX8R6sPo9kACAn9xPrdm7r/98MmS0WU49gPSajz1
sRlkMr3r+IHyrnV10rarfwd6gGa21WJZ+q/mCeSm8LjnYLxO9k4Rd7vuyJh0tePFEZ7rrw/OYXmB
KqgmELTGEzKRgnoGSJJf1TTxMQ6IPuT64g2oHG+RRWH01EXeg6cHqunFqZUtQSKdLB60+N1MwAXz
8yYXx88XvsNsFwzvZMWfmNDu2bjEnag1VEN5c80OH8J2C6OIBMrE3aBzTdKWtXI+mtOTyRYilJdL
43cvbG6deqnF1HjFRwNeAtFfCu5nL8RRKLB/8cuL80LrLIcU5Qc3jwZYH6pFxUXTAyCkKiHb9TpV
aoBWJFDlZF5YEqWQOADi1zlnVdusIVas4LKgwSYqzO9gWp9VTqhosnDKFmQ5OdSAmRCevbnFINRl
daYAKeohPgCJC5cUOlSuIn+K7YcBN30gpI46RQ4K6sGJURijSSGPgywfatVFq/0ym23bkWXqeEYX
09FE4Fkl6s28CJd73SoIV5oenDmUBTCzgOaVhyUvqnXnHJz0e2BNVR8FYu5Simhgany/EldZX74i
bCRBMMb76IZThtiZsMqDMDZSa2np7TjVdYYAoffcCRWL15mWjZqh8JXJF5wFpb0WEgH7coixqXQx
KSrA6GKkHgi5QC+SnAHrmKiQnm5jsibb6930xXdwNT//bocyTII7hjgeecmMh2ok/X0uq2wcNUr9
cOH0MS5+rbU6fjyMMe7qNqafe5QzrxdQs7sJHYk9uojHhEgl8ji1tB9wIoj91JOPq+3pKeE4sFS4
lYO0MsBxWKE4RGntAenGGUxEqu0ontkdznMoJsy75uZajgDiBkdozoPQjm+jHXcI5Jhm6pvFd7Pj
7wq/adevpfmP1YJ/1nYqQJ2OWwEOc6pmfEd7S+Wo/jeidthDH4n/STCyMWiN5Ef88NeoGLGtLuvx
niUaTh2eQQv7WT3yFFya63yuFCVXHa4xv2ocYrfckBpefsDC8tgQEw3UDfYsKTcVNF69v/FIOB94
CrOi8EQDlHKXsHSnKjgmrPFCW3WZljEhSkbjE0/SJZ0VJ8fGdWryb1qcXGh9PIQaKIrFSc/QOysd
z64GyHLyN2thMjQWIKICBvuDzawiCwMwCjIsIL6Kg9Ls23XBuO6lZ0Ku0WLyGc8moxCDQYU8PUMU
0QLQYMXXfW/SL38reyze1QRwdcW5TxuNqTKleJ2OLdHZHXcicKdXHpu+dxPXXEta1oAVLukWecCP
cBwa6LqxeHwu/9sBSyfSOF5UIbJqvOy4YNRRBXWuQT9o0P16sBbCQq/obIdLDrvcDmvSCor/dEqa
R87DPYlH1oRBlDjGOwWlAE0LjrgBGwPUDrBwlJKryEHTPiFjDpGvOtjqnscl34j/BU3Q/FhIp4Zc
O3gmZZCKoIrr9VjW9eclfRnNeahUp5gaaVFw5SbNx1NbXSaNwCjuk2Z3THp+H2ZvMpoCiNqls0OE
SQizVPsbmphtWBcAM2BOzF9M788RO3mN+ddXz0K+Of4L2gYQlWuvm85eTVjxTXGVzIKxt2qo+6Fy
OE8HNSs9JyYYnGE3nXH/Rx05lOMO+2E7RCYW5cqr+EHqDKB8C6OT2gEhBe1Au+1XT1bk+e+TcA+p
rQzp56gyR6bnIqCpahB74jBqGB51HzrsFwKABq03s9pjFZNqoZi0GW/QvribX6iqIw5NwYT7SIo3
aoqJIsMO65/orPkgHTMjxuVe7Iy5C7OcYB2ZMqcpqZxCw38D23NnEOS8ejG5IBy2Y42bfTPw9lty
hSRYXk/69ovFgWRuS4YP8CezLb2ztfxtNCoWqL40TGNnxE22s4pawg20J+teFmtn9Uu8KAAH4Ufl
DvdxE9N8NEAYc1Zxi719QSn7YHydFoiXI8vl6WQuBsMVRDK0icEfrh9dSnyoYGdNHrECEpxQUtfO
R1UxkMFYnjjurDnC/PtY3wuv/nojFrFIxO5/E8sURWrlpM1aK+Wmj/4/S9hVLIGvKlU0EjpQfead
NpHvrCdIZrNorSsdTs5VLF4MlJYrz5hShO3BNuzUVQdDf4k8oELpRgHb08KYjPpvZJE7zaeyjDzV
QVIbfi4R8QydyyaynDfwNuvkkTbhdXxPSnUHjIbei6djXWrbtP2XsYoRTJ/ZmutM2ppk82MIEVXP
BSV8uyQy2sa69TLXNJ1lLBlbGI2+SSk1bOdSKO6U2cf29cUxjDe11UQHKqsAqCedApNTPOyJL85b
qqXhexcGtfGpsALcGkztricem4xuh+tXjfnfFpXRcee55sCFZPHm85c5URCkmdKAQ4o3HpJHbY5z
xnmZ47KZrsJK0m8xyTasYGFyIXrF0PZGb5ARf7Ax9NlazoeFdd97unzzHe0hDBXvyAo3R4wFVMbg
ZwLdHDVN5NASwrSmsMRkSldWdWeKGUWF8mucPDTFAn+q1hcu/X0l1NACRkCu+1R/CWk4/cwaZQ4e
jvP56OMlmW/N95dfkAkV1gUa4HLtEO5wfafzFnaxxLYlHCGitP6i25mJe+CSBoS6Rc9iKKmbO7jW
z5O0CNUnKhS3OtXVLKcuS8kc99djTInXZqrwvUAtnRT0AT0xX7y7SzZekaTsjPldCsl4OXDqYunD
Vin3+WuSSx+uvXU+uRXSQZweeT8yOqdTKHIAcoJQqvMrrfSgI3p3iWn/3+fnrxVuPfwFtps2eQTN
iomHvPim3oKdX5FB4iiukbFQeQcDG3rXlZl1KvcLx6G9gWr28iVjME5bUaTCK9EkNU3YnKMfH4V9
GHWUkTh8c6StVwG2ofJuP8QJFYL5aALKeoT29zq+rB1AdTvAJGvKWnkXalc93eHhtJMBR/xjcNvA
Vr6BssglgH0r42BZnj9YlLfrr6iIHLNLjMs0HVKkFW6EdfqiYWl1yG3oczVGA8YQ4pBmNHFkz5h0
S5nU18MP/W67ydgdraddyhGDRYhdCtXhzVE6X7QN9X/Cf7jBbzDfO8oOZXejbWN3AwI1ZU/IEBRj
yEzCsa+radRLsOrj9JMc4qI1ABO7Sr66jm5C/YlgEN3LYYrdOvvYpbk0jjz68S5gUCm+6aYleMW/
UzMOjlqAUjhWSaKJEpO8j6rVzq9G3sNwLqnKW4sMufxIoNU0J9un6QcDPYc3KZDCyRpiux2gkcKP
7aBhGl6Hnx5WC0OKG0axLkb55MnRBmRAglvMA3RtOgMuixmdMUifq/dgg8cBapcGFrkI3sPSbdcI
ByVNxstn09d7bJ9X3nEQhQ3uIElJPlhoqMjWEaJtm+YPmt0gALHKBeUkEwq4ukO6P2Dccu8Oj57b
U+6uM6p4IQbMaZPG4KE/xVsi2nhZGHAtJ/u3JLmLX843gM2Ke7mQjy/k4ib/1OtGC/j/Dpm2MG3x
AzC6hZ+a6WifiC7C1ybesse+e/LS0djTuhCTodhxL7tUT+bMTlsWpIoZdLqvQa9CVjfeOuSR3q4V
EFQUSvo17sPQQktXW/qCUJWgeKZoy+WHtFOgEqFlB27/8tKXuHYy+zJY9elZqLEz1oBlGHrhjuBY
FY/VJFdcM73CXOmf4iRLUuVjkeHP9KOFL1J4ljEEUNt+UMx6hHD/smRPh7v86phzp8aa726ed/Zr
dhlE8PwdJageVPBA1oMz74+kiKUGlBY6UeVLNJxx+qSKRDEYZGnKS0mp51GgG/I7dekcPqKW1/J1
E8yMX3Y2xYH/LlKoq6itOOJuvendGZGFHOql/FIdRDH0zjxRFqHhCsCMSaWAp5zQ+zsW1l+iIpFE
C6hp7XMxUDgAIlnyu/i4VDpu7OJ3Uuwcgvsae4oQLAzD2CTA7HjHHSHTfF2hOJt9mOv42gQQLTc6
uqzxcWVCNXLPWHnprjPNOjDAAsx3+QzmpQxN1LMAyKjuKCKI9gMgKNQPdBAJLogXzvUqnnT9GiMM
7YGD+YHzfWSPNReojn+u19iwdGaC4hedY9YX8JsYjN7jcR/DC9df8UujlufzTSUOJsVInV3b9nT+
6G+h2QuG5+jQ320BclBi/o36NmGDQJ3WGsDdb5kEZOgCfIWzo5eZSMX3DYN2hKfdsuGIpZIa6FTH
zef/0si+VnhHrgPPBidrSGYuuvqev23WyHchiHIuLdJHcOgiPuOYaz+mn6u6AVEQrULyuhzC3tZJ
qMdlccVsAMZY9IGOdaMjYvyIpB5heJOwmfFnP7q2Gy5ElcuWV/Qjk5HMLnKTIny13BwMZB+xavux
QzLDdEXsxuATKYyOxO4A85dRE6/g085tEo+ck24MJMUS9rjaNIHAWd1vhqjFLrYtk50Xfgdx7dAZ
DCbq4MuLUcG8U3eDeDWJ4kzHEZxliqbNHM+R+duBLBe3gNi81rFBKBNec+feEQm+IVEkapYXhu6R
jv8piKDFaBHYOuJc8nX4u7q/xsD7rMNIeVtGLxp5RPlPFNtj5FBKcccKOJWUElD/bycXn9yDQ7Un
fLCwUojjRr4p2mgPKhxAoHVSxFrGX+3WmZ4iHE+DwlaeWAxAPzQdwQVotkPc32KGv0iVNOzrpyz8
bkU0n0sfCCCRQLP+0iRfUlAl3oGNb58jCGg6kFCRxJzlMHfwrZwoepPg5UJQ3Tl4mVP3RzOgkukY
kzbFS9Pw6Z00qvoLT+LbEAKsTREg4S7mWEj3gmHMve1rT8aSn+x6k88wj/rhh2g6CmhBNV4/4rmM
diK6OHS2dHiAqgQqV/4yblYQlvq56xk30bDhfsJBhHZRLYFBtldowpePtjWbDTMeBnhlf7Bw14HZ
I9/Juj772rE9cyzGSsRdTaJmSLKAKn7+qGQhagZ+zy2aAyDdyXZp1JILKc7hOi1B4i6Y8QowxF/2
pGDOdq5CrkDmf4LVCIB91mvtBlL8k+WHKVz/KV9KBEnchQHP0f6eauRwYxvEgPm/XWs5xlEz//l3
YKLqxL/os9MS/nd/ZOnzf9kMo2qbRASm2Neeffi6sgZYzx0XMZRAHciX0sxEfWhfZy2EEgqeVs+m
fcQMzlpBvrI0ol4PNF2mctusg4QW07m7wXugZCEGONH8kt0mTwmpd8zDKqCOsRjhzKQiMYGW4XnM
f67TuxaMnvVTO9dqOeIuWNy2zMEPkCDE69a6J3k+AKEZDHTOEFRXxQgRAbda+7eysVIuNObgR22m
60jLHJLycueTOAWgQpzhGQazyYEXR0weOYKJHewlWNzkeCtL4W2TObpC64/V1BEvhz4x72zXXVOt
OzrGYlm2vNNKt37AmHI3etfQemCKu5rqLUzBB6zyNAEBWAwq0uc30Spm52NtOfcdWa3MnF+7rQz9
tOsQvIlmzHEDWbQJfsTYqGtCd4dqVNGUOG4RWH+Rhz8MYEVdFDyEeutvOrp4ZeC1GCaf/Pukkmj0
f5HMxlPHnEBhEUKlkideQ0XinPZfoJ1q90xn0gvY9bqhFY7VkfoMDX6o+TTjIMWvKCIf6WwVswZL
snf3fgk8SRi225/A6FkWRTO3lJliphDgCprGYdV7xHl3cc+N6fbvjsr7Hww5kFa5/a72mtvacEf2
UeWerCtgehEiJ/YnLwe3HtIPcBhX088EoKVYwIVUp9A93HFn58b8PqRmof40sIf1IP5aXQccX35U
wdIRNAcvKRliBw1tFAx+8/CS18lxH5kalrKdXSjciAHAf7oYc26iyuzDm8i99nUh1U9ddPmbD01l
V5MiFsgYdiFCgu0urr73VdWm9bFuWXlMWFCueY+sXO5fPl+ITr3HAWaWnadxVBd2xvRLKtl7Nngd
wWjqP2Xj2jv4lxVYEpobuh83Fz5Nr9Ui/9c0AYFD8OqhXbpkDkaht9sAixSm7qclZ/d3vq5qLKWT
PHUe2uIcnABNqSneaYj8UraC6ARRso/QaMg69txwtIvsNfHm+LAJg2SDGiAk0Crqgk+eisdv+d5j
+elbbfHZ9C6rQHCMPHp06yXYjs0NkSeTCZrZmsr9yI+Wd89pLvCY5J3eFzTepM3vYkfGcVeP0qWO
fupW/Y3hB5jKG0kAjcFI+qmxY6Vc6qGkHtDjOmpox+2lD7RdIXwJJtMvh8ScsSu9J+Ofzcv6aHuN
lhmp7hdYHlhZWxw6RezNwg2SVAt1O3GELNleukDNFPbVLplg8fsPr9dVVXVaoz6BbAGLtQQc5G8p
gdRUqqVg9ts01oSEGjZD7WHnSEPJitMbWno4nbKEvBpKROC60zQwaWTSHjNe/V6qJlP8q5MmIqeP
sYoZAOg7MMDmfw3n1UDwz8lGEeI7b+nKzDx5CWlv+ewFRulRi+KwcaZfTt521yH4rYhEz+x3aoLR
oLrbUuyCpB7MMSd+NYv2sin5P2rCNGIWKi8sk/uz6rZDj4Bse4bLt0CpfAHvmhUo0FB2GliPV7P2
x2RmoM7dR6kNHfPRShO9Wp/jJp0Ofnz3Zdrk0q/Lqz+gON3qMUuNgBmD4UH5/NQa/kmExXDcBfUb
2fOI+fFVcX879q2Mbk/cBzVFeTnXfOv0ZVvt5ld3mx/XZ+6k/kFni5M0WvvTwhi89WuPiSX2Hbq4
lJWklABllxoxOdrBKHpDBJusLOnY8O+AjSj2JUonlEsgYjR1qR++KlFru637Qak4sJssc662H8EA
rUt0ZukDGN5qR5CGZ5C/T+c5Wh/YKn1icRzETaymq6F7rdSu/6uwBMy4N3OtqjnUKiTP5IfhghWx
oaYYS7ZIWutH+TZon8f38M53wJ/BrZBB/V4argxJKR+/3H5xwMJI+O/TULyLNklCgZfXAzaIe0TQ
RUPJoJ8WAr6NaQ6j8R8TVBPc4+Cf4864LHtszhj06/zjnKGcn0xrEnWgYNJvmhcD9p90/fBzbQ7l
BJfmNUunuks6XH7YhTi3JdaVhoRKsLrsV/2CJlEhzSF9AOOI6O8HTYJwY0WlBCAfP50QJE2mxi7T
bbHppW4uQYASXLOj3UVbWmZzzENldqsFwdtRH6b1CEsNMLJZoW5wOQMfhVM6jhu4gRO7MHGSpXsa
9RiqVG0ssPCKPwg/LipMPoiG6fLAfsMwxv5rpq+i5efCYTHGk4EiY+ZpvpkXY67x/zCfuKS7S0Ux
Xje9fofoZqWXs7jIn3MNJlBFFBjAVYdeSvdwU85cNvDubvZ+AvRqdImO1djD6XaLsGaA3T//6PHg
rfA8kpx6zs5to3NJWtBo8caDCedvkE8k6pHRP+I10PROcNpNDAZfHh8Pn4P88ltfounAcnNN3XRj
DB0/dDh0SqOM2HFk4WVKUcZMeInIBmr8qGNbwMf/ywWec0VyUz+NCbcxMnTACADA4Aie89RV7w0W
srPyopIfGD0t1tQRr9DlKsNkJcmq8eyff6ota4iQh2bJ9fm1q3StBxquaXRtvV3L31CKjeh1kMMZ
CLNu3z8v6C5xphmzfstbBHq13yJrY5VwjIya6IH6in2jt+SU2z8UI6wA8oDPrGpCH5mcNXIeezZM
+SyhZhUaob1ddINXfNLVvm3Afe+2xWF8teFLlfGMwDdqqrb4hkbKW2RBlaOUE+wNYHDolLZyCifM
XueUG0a9rXZ2PuELuLblrQRIrkyG0mXhSv/zLaf5pNIAYnnM/gtKfaGVCr2wqJdGOvjdpQ0KvkeF
eheYLAuRM0LjGniWkzN6kiVZ3RCXZuBFLvM/7Ky9EYMnvT7I/eaQ30uLw2VdrBE188JWVNNSrB8P
Q9KtS3xNuGxf4gb8Ypq6rFjfJz+jWvg3CtiuEHIrIXAiDaWL1Uc08+P11Nie4fHKCatUPi78QkWL
Bt+ICEsEo4T9UA87ufS+SyBhV7/+OyWmOocX4zpn1EW4SF4sXeVyfJlm2F7qwIrtbtO4PMLHpIyo
JcnOVZn/gIlUtEh9bao2NUx7JRx5r8qvBgzyTSXDz5fqg1q98/UQKSK6tIHAeWdWJPvz1NOmm5Qk
MdSH4yYu7ejkKxBs06KYPdSvJr0PspnMyUdFae00Zs2+v4Z4Bc0EEQBwC6JkIRq76v8RlZJa2s/9
H4dKClL5smof8jRaZ54zagkdgLA+k3I2ebV3xCEMsahIkPYLEb/xABBkNIrQJ+51lmJk/odNeAZp
oJnlS+a7blmEifUa6YGasB08CWRVAhVCuSTWbbocjK+n8Nt0Hvu/QKtW7zcWeFa6286wwu9aGvca
/5yz13sgl9P7Y1dHlcxke0PXhGGpaynOa2OAWpdfo7otWk7mjq8nhW5A8bYIhBw6y9HfQi8DrK2u
c6Me4mzE72lXvQkwuqS4Jvn1cOkaoqhtg8SpsloV1if4pH/qVDBn/fxiw90zqIn8eFqcXqBpfxDS
pAX/K4SI67CMdV4AsmBtZbMunOPozMFcxeM8N4gwow0TVIPk42Hl50z6YAl+qeC9G/3yOkWopM+1
gQHjyTfyI+y04pVhzNXTMsJbhvyOn8qWHzaLWMxUM+Q2OBmWH8aVaDUb2WIHib5wItfcG5wQI6QV
ua4GqUZSQnoZPI970UxqV+m+4Ok501NO/ucybJ5lJjwAGgVuiTBfq+QMJPWdyIZFfl9NeQcWhs6C
aTdtl7lxf2A91WAaKkTbVUrkl3XhKYNDNvn3Zc7U9gVdFTfBIhJ7IucV5lPt1eeRwVgt9U7GjoPT
dShUcpeEMc/Ea3X0E3pDkv3nIp2myMm3RwADEX56tlDB9wGSBJ4JTxM7dtIKyQwUxLUYZUaLJkXK
vnKidfjWKlSUCUllM7djvGDNCaNdYGk8psfY7I4N7/rjun8Qyy0Js0pDpHNhgbjAGARKtguc62ry
3rwlEn/br7Ax/Ia5Wgw7qhkwypmSu9fs+GlczM4zyDwdJyxpVdsnr9qMBZebzFyCFb4DvBau1mwk
c+UxIkDJklgdZA4+xR3mTVN0BINfkrDRx5m6bUuN+YrSUf7Yio6K1M5MoCQeTlQhtlAnOaHi0Hxg
F2y1mVRL36AjzBJ/p0mQbLAtosdXXyrPSj1pOC5G7O9H+M6ExkFfvF97LXpMiC6APKHmEz8iRUfW
XiSmR8l8huc0HbIedocaUaHB/kpAE2dkQt9QmXk9ZEzeUBDMP9SdEi7lEWZDVZXlN4b4pV1I0ijy
zkGKJXIWzPryZ9K9+Li1v0UXUj3zUst9g+YBrgeJ8RGvKDLBnzTABwcYc2t8OHZQ7hKUApRhxfOs
QhyMVD2mOdT5XfG28tLjhKx1dFN2xuik71vhuL0UThw06y6xxJ2wiJ0jJ9QjlYELVclD03Cym9Dd
fLJGUA4rSkH7Z+GcN/eDgoFZV/qf/JJ06/CW4U6FeDmB88Wap4yXnqEkaLTcp8uAisRO2evxJdSq
L6xGG/HIP46ZKtpTi/zBq1d4yXHmWY8VZyBJGlEPoBl84uoSuqTCy5Hb7ul1PL8s1BkfC8BaMpiT
OatIALW8R4J+0awUmoQ4iQxypi3f9brxEU2sdoeYKLV8ipRllbM0ut525J+U1i1Vm14joPPlEuYE
LlekV8AATg6PrahmMBFDDFTlXKZ3BI0vagOVggFNQgsnaM2DTGmxWfxWVpCC7lPPgFzQt2HgirVf
1KrS0KIVPWKU2M3GqI90i8nyI5KrcHhL6rMJv1t6weDERfsVD8NhgFpyF4Y9ksWcJOUAh/WBqi1m
bvvin8EIAs68fegkpisonQ78kxaN8jlcUYC4KOUOpbIbG/20z3BbNEfXo2txzKaoZEm+8Ca/+BRf
Gg32YsMEm3vAvufcyyV58mQn+JUL+V7JySCWZ9JCRPbGcs2GT+g8NZgUZlSBiNpPEaV/GQXWQuPh
jZ60sSWrNur3RPuHquu5311eqeUfDxlMrzn/IelQl5lt2Ptf33w1ylJDB2AaL+wcU6eLRtLtkWq9
4B/sfJ1qICNd+/I5JgzAqUZXUqtX4w+Z1FbBbV2McJaiBLJC5VVrMwPz5iOXl5/0pTbuBSw5C6DL
wBgmZTk0dWLLkTFXS9A/GLW6Tc9Tum9S2DmBXVWTNeZLxqAA4+Y2doFQBwnMFNFXbtUgHENuseS/
OyQA0p7Iar5cX2duAjqj08icpZn6ZOSq4B9TMVu/WFp2lYG1h934Ufap7Ef/A6qQ3Yhk0rothtVr
46XPeIZq65prgLpOoyVOoYrR8pTq3zeHN86iUqlALRFRkkLiw4iGPGKFHJSjsTTLUv9v11O3/Jsq
KUf7eQ6lkteGQoMiwnCcJZr6uvcGFw4sTTmPt/kkB7rltDDiGFkN2w6Lypx5Fhw/walhR3nTBuk0
ZW2KbNkvjm6OjlQT3ONIjJlDfI8pkTM2KrdvE+h9N/wD6GWZPNjs6ssoRLIcY0f5Y0LyW468f/t+
yr+LJllwHA0Wgtav+EDZv64828t36v5fD3+lCUM4DeLxLlobrzJdmBK+ZYHX8p0pNqYZ/HdE+ROA
7YSlp2QZLkmUfOdXI9ZjzUn4+uc27cCJ9hk5t5krXgQL3EoAwrLrvqCmgQNMSI0CCSj9ZPOZeOU3
ItfCONR/jrKJ7EoOfxl0pOOw1/jTO3GAby9eqb95RwD+GzJ/HZdh1WRPqO9hPTDnMBJkxFQGdEI3
edM388XOL1+n3njlsjF5ERVhPQWDwMqSA11FoHpOAP9sFH6sq8AZe0jOtEoq/xG+N2IgPrZ4UVAo
iKskkq+ztCJAb30XTzbrFgt6ZLVBnARuKKkTZ/Ur781vzcaoix9HKKuKuAp2ehnfzueqpY8R3Cuv
yI+JEtYy2KEFmIWGXqMLFB7/XUzmusErwRSl4wWrEA4C7xJZ+VoHcXcUTTJpSUDOPGcPP/ow0uKL
83CxwOJj+2jYWdxM8Qdd4YA4O6yh+YFcvaavk4j8NvFWlHArqa/GB8WNcjw3Vls2O8aVuNlk8r4i
zrCNbYoDkwfcm5UE6wezLgMJn7+fMLnT92jogPhtgJfl6xWFczDXYdKpjQasRgmXBBZyzKh2SmvK
DJzXu6HNRoRC8FrGIsQKa8cBZRKDDBez/dZa8vgDRacI++jdSTnB070qsHD9cGfkhALtWOtYl4zF
Pi8RreU2O0z2/tz7PzkNq1QgUOXrRAF9C9nSCInOKnmi5qxELTZk+s2CJTKj9hWcQur9/ED+kUTB
ppVa7/uudeYQFsohIPC48EptW/dZzMxaRX/fCdZpltgI6tpzJQ1P1WAZ+UNX8zN8h1RwEotIywTn
SPNS13Wnb8Os7K8deqSYLQDFHBooMQd5hBwjZoDmL2v8thSzpZVZ2lFgby6cyIItBUXMfYAQiyku
BFaDKPuAcpG7hh3Jqvldbamv/mMHUCsa8upnVSYzQZ+YzlZbsTJb0owYxL1rxrDYhK6Jxf/VIkwb
rpND55Xhaxgvdg+XX+jdfeF1u9/iLWeL9uHkaDJSj+4T/4QxYKGJ8hT7fcJseIwtRLHu59/t6zVh
qc/WWAiBP8PQfTOQv3k5OJFhlmx3ZCXC5S1cajQDYABiwN5ZNW72DMtoHgvQIKDx+x3N4fXdaB0k
jClfv5OOTQKF5GAFaoHdAAl0Mjfx6UCdAjW9olPk34b1glAP8vxUtQWsOfEvijfBXZ/fqs1zTboy
Aaagl+3xF70/njxQFBmdFeFFp9MFRu6ReAx/zR3tcifZVfgtBmQsqC53aU4iUQGKx4KdfEHVgUfu
e+zKBUVNn6DImZcz7iLbNUfddDgnqSCkHtrNCA0pxsQ1V3R9nYQMqW0njcMkm2FHYgO/tAGWOEqK
vAMLxZWWS4SrXXFmlR3a3IY1xaJPEyn9tRBnDU18LrRuubTthIFX/CmBZTW7eSStuTmUWzY0ubre
Rrugz0XqxUOwn1FZmtdjtlGE8DcNB8234bDyZ1+ZxbQbmAfZ0/UbKhk5qUA6ZFNzL74cXz5p4Mo1
SzagJ1tIMKde+iQjZGx1QUAvcofhOjskNY/7avNH7XNnfixiZXqn4hjn0pBhAWWSucu7JPppIGm4
zIPxVSCS08ll38Oekvsnd//y5KwtLdHXccdWRIpQsgFPpDsUfeHquV5XeE2FcxZHbtFHtH6X/YBm
q8CUEy3w5XrpRbwgPDBbZZJ9zlWdN7BF5/902d+SsrfmZpOblz++kECZiHjMYX32kyxReSKpFJeo
KXUU1RkkRT+MkLL73bcI3THBrXvnG0s+5cPbWcn2xkV+TMoAERfpKTd/ZMPitWkhKch2DUTM31Ny
RZCWvGe5RFcSWpfPviweMkjoIhmnhFF1fbQcfWv4mxHeyA+Led53VOb5exINYWgPojgAcXgdKUDw
9wj+K0j9uPhOXCA9xlagU1PSEcpaGwYGu6psg2cahZ3WyrFjDt3D3MNi4InUsT2ZfEdutayd5uVh
B47qsRsQg/lNjHOABVsWgDpg3iqKx7a6RS1HKtAuoyRTDjJMvo88m5spkLOEjryAHcP7F/QbofZ4
lRlJXDBDLgrti/DT3xhbyAMdHWNW2FjaoOfp/IAvGQFeH+PO+R7fIVbonyVUS7UCvwzFO6R0KQ1P
HZIAGdE6Yg3nGTV8ge4tn6TI2uW/UiVF1AkKG7DHkhrrLWWOvkTC2oBy+fi/JJIv+fnB3dqDS2Mt
VB1UO1PgcsuTnGn01JxdE2FK9HP7iGh+Nc/+TZ/rhLKfzO4B2Zo77Ojsw6TF0VoeG3LFxjXHNffB
QqyrWZCX6Xhcm757qAKsiAnDIf8dVbAtlYjD1X7rH1cGuCqf/cVdsRO9y0ShvIxaGvEzI2l552d5
15cOg4YSdcuLlZrVEgvOI+X/SOZyfjGMYSA7Mbi03jkfNiaqtWt4e/Offdiykz4XqMihC43nFPfl
TsZ7Xc8/OQ3z87HLB+/R/N7+rOYByE6Gt60UNq9eFjDCLJy9t/Ukzsd7eYIjjSQAbnbkW64hUWhe
KGvUhcwoWwtfxcq2Fp/NnZB3r0WswGTvsKDN6cq3qXnfwjUDy7zbxoqFqubDBgpDl8e0usldxdsk
igsS/3SErUcKTRgNuPcC+W2P3Dlntt81op9KHJvQbMFfHawfPe8DJIuB/VIok+xXK4AepxmfnuNm
tVJ+TWdWka/hfrqVQ8K6h9DvBHynPg9i2nbE0BtLHpZzmXkIWd9cdd4MFnyUsG05BOHkAEfaspZo
2+3lNAZmjpDk86dJCjwfoCrTpWpNu/Sau1HahfmHUklFMyeH1fgLgUuSJ18tEHc8qXdERDHP3kwG
4zorYfrQxBItjcq3rZ1n/kTfIP47kumeJ05GuRIK8S2X+93RsvMKhUsmZCBLbrG6PscBHrE0Roav
Mk8KYbOWyd8bO6ooalfs/xNcfUX6qglYPFavWGQdKlVpyAJaQecksFW7kifncOa9RPibjphXcXeL
5qoqDgW/33q2hv2C2qiWi1nXQRg5kidzEhbEVJ5PEuqMZGQQTkGEjPPPbAOBDBMLS0+uzp2CIC9A
WwbwNiXkDrO7lVm9y0lz6q6l0TCq+N313zRu4/hH6K0rCXhzFKgt+/sWbio+KgO2pKosIy8PZlcW
WOTbybzo2pvRgW11URg4l8lnO5S70L03o/Mg5CDSGK8IhJRDitPBX6FtrRvHPs9m9kUQwR4PwFkB
ZoO258JyfuzW5VUtblMXAmWZn5gTRTyOe2e5leYlcssU35P6YpA7K0T1pGSsnQnIZCbw49ZvzqIo
HgD9HDuZHH4+uNpIN1tZBikYd2Is8CENgOILSGzV1VbJK4+OF+9gEAyB5WxVAKQqW+hdTbYHqLw0
1hTcoa6NcC5G4Nx2V9EOoWALT/hey0I3I0W5mTCVKGB587DGamTOpyZXQV7PaIpIQy1qguG5SH9t
K5jukjZ9i2x0CH9SGl754uUbCiU1os1150ehK6Lnd/O0kXXJIPWLcygn79alDAdaLVmDhpY7be1+
GmDdFXhCujuPBYBDCupakEcnsM32A9ixv1zpzS7vl3xHSzexs/y7Si5Mv18VTrob3enakzg/RogE
dte9P7EoEr5nQm3gN8G126nKS+UyepQVStgejtqkRjopWDYwxQx6fXmahDxfs5+Q+PQxZAMMvqNe
ReggnphIzIQ0baslnKprU8c59uGu8RQzTX6zlwWcvzHAz/z5PVQdfilA5Bz9fz5bFfhL3mE/CafJ
1isyxp2kcQ5O3x1hVRH6aQP7r/KUjSgrgDN+NqOHZr+jrIlS5P+wWeKZcEOBMRZDERRZnl8BVSbX
V3pwIG7xujfco00kqDX7Pfhc1IPopvz7Zj48biruDhtcHmbASiUIivhWR7eNv83nPGA4b8FhWCIF
GsfaBHSoQfhbPzmgdi4OSBpPxwEyZNj3AC8NS28YgmfeVlx1og5+7Rw88WwGGKF+CIH865Lx3ARr
kx1y8paXTSG8r45VAL8ciaFhfglvjlrWJOAB9fJhgoOH8eRE3h2Y8WVMDl0Wk8B3qzjTNYvZ7+Mg
OA9SX4Um1Cg4QeNpExLmlSCGoKKy9EqHqAvvuMchxJFM4IRsicMs/5N7MDna7kkXXIkO/WF7rAqC
r8U2c7xTPMwVjjga+x9DC3hvL6nnWQQDYDq5QFbn0QWWQgOq7IktRrQT0Fg5orW91HG3HyhWAQ3F
mbORDWYyRGzyxT0K7N6veIW3HTqW1DIr2pMfRJYUHwmt418lx/kAHyDyUN3hcjx7PGEaVXOr76aR
gCYSDb2hvm0AeBZIX7cHbxmI9We7PmrRoqAxbHFhhY3gkJDM4aTaQ4lb8xN6PzSz2iyTKqOVmGZT
Qm2diBym53896gaAUCEjUeAhtgTj3ONSOOAsPT1aR2UhLP7Kajy/TfsadI83VSoe6/Y4ad/aQLUj
IDLggtxH8HDWDcIqtYLC/p5pwLckPLR4zZIHFZXQXiuWKEMrYjgxYpnY+L8LFKb6dFqNU2/3yjrc
z/Z1NfF9HArmudJWDWCRsculbYcKJve6Rp/ssuFrCp8LL2j2tx9v83dXRBLajJzdXwNKWWxi9gr4
ilEygBIDuWEukE/v4XT9bjeo81OFo2oscLRNw1B3aD8oGzPqDskPZAZrtghj81CwJrVs8VfIJL7M
B+GaTeCj9gGVjVEElc22Ipue+ULnp1VzBy8sF5D9WVXluxHSUTzgTs45sIppeqzHBbk8CY6XUXwd
uWhAoqaX5SgLQfCT2NEp/y+JT6vwJEsF4spSUrUbhoTpDOjDA3kW00CzMo9eb9qwcOAUUYaVXQED
k7VHH+3nO/VYpQyPEsrsVUETxcjUh1iJvYySozkNeZhRCyCkQZwIx+11mxp36Ha2OyTw2n4EPQrM
Wb3l6xKFCv3gh86SMarVdfYoc1qiZlUGrEhxR9/6Qn1WJFKZA6RsN1WMagK64w9TELkEd2nR5Ojy
xmywjKBU0fDIqLoJ3NFEF+sdvjkgE32zGaQX9l7CcaZqjJRiTVrtgJZ9g9wBtdZowlIWNOlEtAAc
xN9df7A/SQbG1aKkjnndVFcRh+jCrDK7NgtoDU/sIvB29EtEhrzn3mqhiFdRj0aHXKcqCD0oMRyK
v1ezFXyAchmxek7WyslB2kepDW2mZYIB46mchVA8716KNN9gu8vxY7aeX9HGbmWGur3wqe1HsQTs
kuqzOTLck1YKgOVKVfoS0+nnHTMUW3fXJbB+TBblALN8FCwsqx45OwAyySc7HUT3QrAXvVjB7V7H
HU0Ainnq6MBcaeTpxt6iOCBU/ecCb2q6Pjn+MnILor65TeErFF+Ksw0O89yzcApt+yVPLzD4ZQrC
7MeUbg94G7xjrA4Gd7Ixb+vniyzmCb4hz44JUqGHauEGbl3hGpOnBtjcdMNcRgRN/Us5JC7xYptb
LQVQAcAJN3G6ooSXzNe4HYkJzr+5SeeBMa9y2fJZt8vyXng8JXZH7MAECjwFvvJzoRnaLg8CBMgD
Gg9deucz75wdQPKsQynRutXdNfbWVmdJLLQn4TDtWIx8K2NYS2ZrwRuHobGVoJLdUljBuiUh1aRC
lfZIVhkMdO0gvRIzYfbfiDcXwDyZIFviNd8ez4xkFd23+8nh/6ej6p+c5INWpYhlLncaXYE7K6X+
1uy5GDzt5aBluL/uMShaauD8v+xLMzlNSPVlCBS2fIPdSD7Q6NdvmC3NmTPXR4KmHM2dllZ/PPxv
iLJLMjSdysM3yN2g05b7ogJrxYaz+TzIz7X0+x5d6Nfd70pAtW6OUOIdmyFTfewE6DIZdde0y8zn
36Om7d5aHmJ3Y2VVKbyX2gMhe3nE3BdIZG68ZqJ6cbC+AAFljRXtnsg2rQrI6zpe/XUcnmbzmVaP
2AAVyV/vlv75Kt1Tch9N7h6g4NCAfxfYV7xZ/4faCsb4PjBZY8TmODhjQyqn+63hZhsTrL6Lm4nT
JXrQ/DCLjSO/BZGmQgPXsZ3ShSnV6slCdv6SVLQ9q4lJI+ql5p8IYfb2+IFsAIslJD3zxdXeE3+V
BCG4lpccyoeAaajXEdha2mf+rVmBECEIbJ18RLLIp2BrDXrNhIile1WMVKsaIFwmg/Z1RRTiCr6k
oIM5RLrYBIeo9beKWgteskuDVmK2n4KTuPTyEieLlRFSSHjBfKtnVDtzjALplc9I5gbnD61kZJK2
++ZUu3bCcDcZGHQLS4oi9XoXkse2f1HpLq3afHJnJvKAlHLysIrTxKQ5mNE2NdtZMp37ME3ELVsZ
tgPHBrL9Z/ryobwHTkhUW2EdkgsPPa0NUacDLDyI9RtOpj2FXPdtYOinnGW9/+Xww0MiV1FbinWr
BB54oEXyuVBi4bsOqWNpkjds/4BmXZXMsDjIJwBRIAZ3JOiTaauV63H0CBEc0yZX6dA8XR0XweTd
0lqnqsSE0kKeEbKOCwhCPOU/z9KLIh8Poet6+3JtcwKkiAeF/+oZWsVsy1owwY0IsEr0ztVr4V8I
Ckz8pOoy4Hl6aCr/Ubbu6vYdRrBxuNRMkbQ+p/usVuRiSVT/XSYRPFzGUDjHRAf8bApNsdUBAlLW
zrqxCdGsxjR+v4xS3bqNI/Vhi35cjO6PcjoEqkGMX4qeglzFLMA+aWn9yFyVuGxpINTMj3U+uhYC
nHME/M6xKnNuj1MzhT9Ec4qqpyAkanqKroe5L/Q4OKr6BUi3SfokO5u5QlLq87VGe0iSBbRYMU0Y
Yp8ek7JVsGz3ocHFZiP+UmZ0DUAHJRdMl2ZhPJPeSyNGiZ6hQdy3+KnRlVPstSPhBmAC+4xg2Lut
KKft1UGf6KTLtNbI1RvE2ES7fNJ5Oh3wxs2qVnhb7gvkC6IpH5JANfEnVmasTpnyKRg94e0ceKsp
UMSpm14gp4oQ1W3DarjA1soDrFmo4+E7g5zwIDNM7qorSReJoeLHT7Zc0P2Cl+EDVW05jYqRGLai
iLqCJoMYkcE4RAJVxgVww8nfl5CSXJldzCde6UH56YKEBdZ79U30ZnK7RAx1WKRjMgpiafPCZ8mu
PUXapk4AeDh/5fSuR+mTLqnRMbpEVF9nNhvVTamNtao9hhMKKttaGLiqq1VUJvUBYt4ihAnnVE2K
noKHsGNO8x9n+yhcWWJb8qOmKnq/v/N8WLBLhSbFWbTRQOdS2K/0Pqu6ui1N3KsGVN8QneDfs+P0
0TI+qT6AERMKWa3F2FeUi9lNHRp7Txhl3HpVXUBL3QG0sRVT5A8jh2jWCTQBEGpTj818W6ImP4U2
wZl6b8tmgOAFPuZK3xdSMgARVXhKuLRFM0x5Eo1KNvl3beW3mDmTg81LxcZuQIzm4DsyBYfrPL0H
wxTu3YR8RwuuBpPb25wJEAfY5SVTmgKLl0/je7S9qIv8+3l7LwlBs/PTM7FCgAIUSF406JyqHfmj
mTOI7w6Ux2/bnn3Qihv/L5wzRXFlg4CDC49yezT1VZ78QnwICQcJYVK8wQHCLaD2pfvAXDA6sfOM
TX5743VMcmbx1TjvIHChHuwvGednyLEKYkwuTxS+8nXyUMYLpXh4kExla76Hs8NYz/yDcc95/u27
k1mmfrHVC54IG7U4zVFbD4c25dUOGpVSZ0gSlJbfvfBKJnJk0iJ1vjnPFhbcfjsgLefnVYFri2zZ
HiiW9KUiM0B+3e5dPE8RIzRJXF9oxt7wrQiSPPz3zRxjaUSLi9iGaw+aPmDjaiXR+MZtTOlHm9en
frag+G3uBekvq6fF5HSBqx1IJDSggbOouRiPq5RvoAMmrIeAjht5Fl8QSWwa156GnDCBXqI/WwIT
p01PbEMBzW1MLTKV6qdP1CWKiHKOe1/DEQV+mMW0xf3rkWiLuaHv316H+ZYrJmqD/LHyxQnskLAg
8cY5GgCgx1VIhXZrd7vQmbOHvEAZjrba+tAVfTLOr1X5SL5OT/THrzboCA+WB3eX9paCU5hdoCEJ
TDZ6+Z+p0wd2fTEdBOfbaRqLfMwmiPhoePZ3Lfinn37ee26OJ/F7Fk5Hx4A2IuoZlWA9u+bMDZtG
LAEBt0UC3JKap3cpDtXMdpxFAc7bhgGMB4MaVRPg3wVRaDKR/eDHuGQWEBIRi5EaTtK27OdDbc7X
lwO5Moy9ziRU00OW2gE7dDGwaAO/POKSH0kxCc3HAAG/p7iLL947efUQxBu7QrVPCgASkUQRuuM0
TDr0l6coWicBIe59L4gpRR/HC2JjqTmp9w+x592SZUZjlAlqZ8I+9c+pL4HybA/dJgzpVgKSqKj8
sFDU0v3sI8lEd3y8djk6g/YdkZjYf5iGv6SdXBM5uVpTzrfvmsvf1F2FBhohTRNMu/bB5yATC1pt
71LR/Zf70VvO3gpRSYcxu/m1Rwq38F+Se2IM716OI9eg+GXLO8t36y0EPnX559CampK4dyE/fUYN
0VkpWY+8qagZifE99HELEObsfSb2ruCxEKeCvGCL6LEecsTJxHQZAOtEYREXT3vxBnKEzuAPAoGL
UwVHmVYiHnKQ4AcisneRAw3HdyitCyFYLM7nwjCG9S/Gf80DQk+YhuvLfig8OJkcyDcMk9ZkgpDA
KCR2NllUtFccRaGbK+lz+x7z8yekhz2sn/FbA8olmfoSd+FXkdfHnrJ6pZYfld0XGomAdTBgw5kW
MySECAhSrK0DbBikObSkyW/B610GYffXLyBC39ge2mhqLxVOiCARGK5MD0e1RiJrQmMGkiHe43H0
ayIKk0d1HAyT0qkAqV6vyL93EUIeXbXHfVzCRyBWj6eSvEtL+WLGBaeK+ew/Vz5DcSsqJifHc8ay
cGpAjgx9HMrk4qTrShXga6bt7VJHvRK8vjAOKt6uJ37U8V1PTVVnSYDPIR5nTKnDdBpk0y+bHXYF
tHgvHQHz2TdaGoJVxt7CBQD0l9VxY2vL4BJIAWNcDTl+NmHHxgMMR6amz9VLrb2SOIrL2B0xgdux
XexFuY2Fs5x9sAjLDothyt6JlN+PWhYhS1cf86wicOpnD8/UQ1qDahwVmd0wfEk5RjZgbUrO6R6H
ymy4wbcHzX/DGqTxdkE2VfugHZIIy0YgsfZR5zVKZgnmT0QiVdGrXnEPjO2sWK2cmp6i73vz7p2L
R4lvm83rfu+mBqbPfCheLIy01zdChWMAVihd4surYGn0Cr6Og6elwkmw89V9UnsoI9KTd9JDCXNz
/ZvB0vbABHbDV+Mh/x592rYs//LusVIH88nd4C3K20/Wm7v6vRy3E6hjJ2wb4JVrPni0bE520r9G
EXncvDxyoKksioSWI7AorzHLHs4eeNeuVzuVT7T1jJXptEYgBNEI0Z0tZUYsOn24YO0wDacSv0hx
PAoeW4420iuS7Mt7jN27FUWJyHeATAnnzSXsVTPmewD6yO3SwNmy5O4/t1nsicdoYAAMN99SCQG7
51SE5iY8yXvZdZU9+D3w/9zO0/gJRs4M23OtgFiusyzNyEp09zB4wJrBHsMBtvod0NziHTOFv8kB
bJ7ibNrRAUYCUBrtTQBBETeKTTrlyjSEKZ7+kEbnctSSyTugIxR9RPV8oAhq6adkVw9dhjenbpqE
RmQkNLW5WzK+p+lNDULIZDKPFGVpSrpaG7FXfTHR9kr0GE3/WKvd9eGuOTnjSU8Eu0fQqOtaRmsR
nH1bil+6Ry1RlebCQlsm2WRMhmTLYKPQpuCSM4muvaSl3+cNmo3q6XPBKUooLMmFzzctP9IyjkY4
HSouF+SFENQ8egsab1LhKtd3uvG5HMwrehtqb0FdwZGLrmbxD7a3PC7yyuEQfWEiP/kRF96WD8jM
6ItCO7q2nAbJHI67PgPAwWVT+cPCt4IDlwTJkin6esLRzOlcobCPxQWI3L+DX3vuaMY7IHj+rSWb
yRdpkWNCdzG/zPEN0cWtAHc9TrcTcv4+WeE4pMNiL1e7ZJH9mzseAVQb8SdYdUcJtkEQdGtfDutd
6+lhO6k+e6KbwmkNv15pD86ysb7Vvm0XIMkwUy87z8/vL0dhKsP3PbSJJuXzjC5jnOH7ZhDyMR7p
oQ6UD0/+PFVQtQjZ2400ruIUqBc2qkfYwWdcgaJBr1rswcLUi2yL+xn2J3iylDAgIM7LqOf1cozw
ZRwGIxYYfk9apU48E2FBuG6ZXdnGro19HXXF76bbZR34tTF3ogsHs2ciiYs429yLp4SyBL1eGY+v
CH3p2XyWx1BJ4ERkUoKefzAZe+LCqMr3B1OCXFE5NO8kxYoj0dc2A8Zc6DyP9RsAH76qIpSkM+wY
gLDCF17F8rFAKuIpmIgYU0a4Yn46NR7lT+dOu5IBdEeRj6s/FTPTULnFZ41j3S6bJlEqbKBcGyME
0jf2/KtrmaCou2fPI3Y6+654hxxepjOlZ6CV794qJvgn7OHR8Xc+KR36CDzFsvn3ODuB2AbVCpLs
muSLMea2f/nqx8DgOvM3uztTZpN4DYQhGW0Io7aA6/CnGm3NdZ6iRQ+3On0wWZCaW+gqODBuUbrT
NpuEUN9FCld7tgktFPolUgt+m0THQRaSNiWkG/KOtPYxOSzQVZEW3Rc6GBmgZMP3PM/oveCe0/fG
5X4sVeym5UcKD/yBe7x0oQLxdM14UKU0UCMDLuZgSjODbGEqoi1bCxqhc5R2Vg0Qpgckc+cZZYX5
5eo2wl+mNVq3MZWkz3MJ4lBl0xUAklvyigqj+4slaOEHpErFGbOZYLdFW+WK4Pm8k+DHX2w86oSr
qm4QYDfIPy5XRGapKg9aMqIz/95O4nsGOMwMImo2sH1NPPuUn/4cqr4TOLlShjlt5ed3kD2SBGTT
2J/d2blf2ZMQfcRsxRMns8+H7XhFLaIVpYoKLolnwjWEcuk3HqIHzFY65Ux9F01ipyeeRAF9oOkO
Y5bnQZ4Dtto+CHg24wlEAVsvigoLd2+O9iN6W4gIDUsvyPSQbUQXzc5K+10ENXenMwF+KG+ZryS6
6e8RDEEbZOn+wt6JW0Ev3zeLJfXfqhzSQwFhtpOZi1esxN/Q6voxarmlL9rptlYCQe+GWj3cwnAl
KfxGrzSlOZULDYd2apokdadJ/a1hJhH1CYkNQGqA6Uj8DKV4agJVqpe+HzXrgwxCmTx7ZYSWaw5B
goOuvlgu3lgnCYmttRKpfQNQuAy3cvHQWOVyuG6NM7LlRMfXv4tIYmuDRyHHKBr/szwFCybvj+5I
8M1/v/JNvG3vdWeuXv79lSMo6CgZo007S1z/jEAv+dA5ZcIhoIG1BrLl8I9VFXd9O3stwPo8I8cr
YKDixEW5t/ghOmbboO8cWMAYw6Eml7oun6C/1yX9gpR8SILMcq5CUz0iNiiY/uYOxQucO5G9Poww
qS0Bj0u24xPbf9jjXeefaKD/eWHbgtLEGbrtuubOPmx9r9tvWgjPYPi8L2RKHBD/qkB3hxHPUOSv
wmjhbV0F6EEH+UgAHHDmka7GQ+ZMnGZYTDti5XyuBSu+FShU6kxqtrI6/ztaUD/G0sB3KG8mQLhf
ExVmZcHFLaNQEV+YTkKyUZl8FjUxjRo0JoUhBNPWEr8asGUcvMxQsbNr/m2VtcgAM1mV1Rq/iv6e
a73grg8ZhR7SaxScm6YD14OyQNLRqdHx96EZlzYqaJC6Oe1VjJtQAp1R3hLzMsUNEPg52Z4vvXvP
tqVo2tQtuYwE5Mrx5jajEmVi8GFBiwT85uWc0orLUGnfDqIZk4+ppBPMLQX9XjaLsth10dngJEXd
tv7D8J089fp/zA6RD6upKOMjltK2ue//L5HKKuQI3a1JyWXDbW5KabgaXPuogz/P0awTYX7ls0Lf
R9ccJQfeS0KVGpvKqis1n0ITIhRyBvIZCFOsGkuiHg0vEFk9hqDtkU+tU95TR6/S7kH1tz3UVf3Q
2q8umF15hO11mxC7Xhe3sjiisfMLlhANixMK2eMo5HH1/BrcnWCscvSbaHDu+2pDUn758gx7MUeb
YcZC/eF+pkuBdlwfi2BiCxNjrFM1gpOPreBMIO3AfZGGWqRMqX+2ctH1ebMVYUaiusAlPEF/rFMe
FmBG+BpaYOjO5rCyf/41xDBVUAPLB6GcMZI+7uRRuTKNRR2q3DkOQl5d4dI+fpWRS1Pt5qoRSKMd
wIenDqRN5zRL9c1BXsY8NKHfJXoT7OktimPJFJTIHZGu9mZOz8t/rzm09cZqN4z1bqe9GfRmMLsm
qO3Vb0bLwaLuW1QhmicAymDixVnnY8fyljNL+YhxEOthnLyuBL+DlLjIZDZvh7zSLThfvnOoiQCv
0wdnEctG0W03MHRcYA5a4cGHtA0Gq+pYi7UahjODjau2RgY1/xvcE2uM+TNSr2xw+67awu/muUw1
pd91ERF++znKhSrMhl7L/ZS3N9YTQrcDYYCYvaSpvtBFQ/snSLHyLdJ7WXx4XGdU+GxQsJkMjt9r
oCF1qEzBCks7arIwfJra0vUZC7o0qKjONdvwvIqmgq3jVCCFkQoa8pwSsk7uXAIhH5DHciqealXI
ij2ZrJ/SKv1uVNz0Fnx24WIZI7s4Um/hrIACuyUUYog4tdjSXYHafIXiyZkUItg3wmn9pw8I/gDT
8lQeLG6NsrbP9jZwmtggaXBTN5I2KmAAILAqoiGBfcs9oCAl4LepfaLRPSYnP3excldcA4puaynh
n7nVfqEeIHQU2Yt7rXtFneAVQ+q4oFKq+OCZMnldrnTUGHiZ4DZakk50YoFRZRQDVf5jKT+sM8iY
3OAnJVcb2oYbr0jHGM//UIvrd+sm5ClNCO1uxpIvvaDqfgPTyBZMdrFO+Dsm/pxFCGUkVHnm9cMD
cpy1CInRpgGK+G7Ff1Ikxa4daFf36iyAhKmWGBRYPR1WaaA4mOIiH3yVQRrT2AVQK+yfutNhkbv1
Gy5KQohTZtoEQnFF1NIj1tholDl/m3qZeAVMU4+jdkkt+1TzEAcFxLetnFu43umiunRg/7kLMvvD
1cuCqJMDr99452N5BTU4y+iTNtSYiwUqgBytUPiFahN3sHtQ4320UDRI1bz22NOmpgVpXndd9aNb
sgSkFKa7UcU/EwIeO1ez1tGTlExJcCByIhGRMn+/uqWgFIrFPzPFF4wUUw8BZtwdbzenIFebwzov
LPlQOD7obAPahtmDIKLpUYAsjpjHiLv0DElgXvETqtssbEfJsc2ylPGlZvW8/BmRrBXIy85Vq6Oh
fTnPghlWIJQy/66fCdLCyyXk/KYj/AQW3JQY7aSIxLWkcbMHq7a2mCnj09RQ2ILiUFpAEYbsErWg
TRkA6PiWTP0HHo8aV6Pax9IySOpVH6BCi1WgR3AigyTPDqGwP3fbf9Nbxzby6au7PoFmMskIejcS
JShh5xo/IRhhaGDQhtabP3I0WIk3DYI2gSm5vOnY4tfd8QHAHPo0K10828QqC25S/l/ZMo3/rq13
fJvn/VvwRlv+5+GJxox+YuiQiPU7cO0ujl3xlxFdR0znX3L0p1+n8doeXM9DcrIkrAi8iUtJ+0dU
/D6WSMetYezzwsJnPSkqx8Ir349jNLtlx2kaPj8wATq7BvJDR1LEDmbgybEs2lQruL/PpVvGRXVF
wKSCq/GY6gmQj4hkA6HQci+DJ1GB6whJh4VgcsXtKbeoyF2pjuS/h02yCKfGjAb3UHM5Rn+Z1jYb
RcPYltUnisrSIjBf9+F/Y7XiRCPuvyxhPzBYOx0JEGG4gUl9O9S+ZFSbkMl0leRMzzlpAQ44A0xP
lSX8aJroCGHxJxSbNS/O++PP42KkazJSik+U5ny0Fu5YQqn7VbdYNCcyOiDI+SSE4u6qGy1xOie9
+aq+Ylnl3hjKw1+l/LNPqzaLwUMmW9KU3Iq1WhZ8P8fduGf32BLOwJmJSWeRpa+HBFAqGDwUKwTF
xB4rC0jxxPnLJZLjvUoPTOWLz6Zv3QWsN9ebm+GNuuCEX124dq9sSVpxetKyG0ZsU3I5bEsUPRQR
u/sAKnxzfUYxuihkpABsuXpNwiNjAiC3ouzRl2WY9PxK0Oc3gFqS3kTxWNHFGxdpkJ7/glI3Hw7B
HB0Ewx8Ckg93s/4Bqfvbi97s9/lO2YBQ6kIVFC0tsfJCl22A1Ep+I94eugF1PGdLOItj3PJjJFkG
TY5vIhXxRAJNNktjIEfrRpIYr64n6y+imUrORxch83I8VR0MJloUXXCGhjlb5vCpsde4qNVItYJA
D53X3jCLooyYkMNwwrCtW7vTkjkYUd20VCO/mYHjSbwJ3qM63ydgLxCRssOXprAHfqV/rZ0oIQIm
EDglnl+0qwYvX9h0bkQH0IM1Yih6bmCLp/D2sDJpgmKJB1om4J7oABBb+4PEwOPABUOT4bhkpzpE
d9G3jEb0WhiH6DksJVw00R2O2sH10/EHL3d7xfYY+xZbqryKSvavzneGPhekOUnRBbbzS0Maechp
9OUzL1DTMYJsbsg/CbnGPKgQSPLWAfuoux2zoavUYUlUerpd+LJ2CuXjzPPNAtSE7uTDHzxus+jg
eP9HNp/RtbJaT/VwsF1rcIjCf4YbloPW0qxDSx40VoqOVhLdB6UxRjhdRm15u9S0ETQ7oyT9oPW7
Tpqqe2JlYm/EvVgEwI3pgTygbNoiVMYDZpgEJnry7R6dsgRPM+GLwFbNHCOxKU4w4tIUU5ZsBQNG
U1X+alf5PLjx90DCpAHK/AZjmfK3ODWp0FndX5KWgzpNFITxKkNNW1ZAabr4N0eqPQTmcyEzt07t
Zlu+m5BQZDTZOvRhUANNvN0LAKtDmK1+z+siD+rlaxP7Fe1iZTDefHxa27fa/Pq6qSVdkjRYqVTu
LEpwKxB88eAqa7uEr4850rd0pJ6Z3bG1YuFYG6WUT7WcteZ3ncQ7FlhVc4A3LOcRsnWaxiNQe1+D
8iDaBFNgKKaAHyDLiTYGb1CVmyFfg/k+NvK6AHxnl1D7DGNWEoWcRyl9mmCizV6Rz70fK+jfgaO3
wydizTd0rAnf/qTTyQIFMxd2XIgP0ZqNZge+nGnjPsbyx7Yh5IzbrBHXY2HjlXEjvprH6RO1bnmh
xOD5lXi8U3Fdy3n9LBEfujLkWtcbnv9knouCoQt4biC2q5u8QVD9+XqWmu+nRM6uZDiIV5jmDqus
nLq3kTFXEE7Nx6bRtU89eufVShCNWFc4eMESKWPNdM6bNki4o4hJf+rBXRDBp4o6mRQugP4GGcUK
cdtamMZIJ0J+PUiLxCl1p9AS7tSIJjzGCmLE/f+CPWHqCxA6xlK9HjxlDwxoBZeR7nBEDH+cJbKJ
q8AAk9nxkDCfMxq6yGoQUcsMKO/hJiZR/7f6BzJMl2xLKHEC9ZiiisfLP6dsAxnL7kkwffYzpAlM
w/VmWVcZwpakizZT59nZ9ICxQjCTNtAgJcUDMxiBxOoUZ4iB8Xk28Gvkc592nZoL7OYVQQz/IH3g
rOI/6bcY9fYA4gfzO80h3QjKL8TYTBjWRvAxkbzqzyea10wXgiEUxsss8CAPUlybeFfAgrynRJpA
8tQXLe0zTToWiz54s1TRXxUuU4Fj1BM8tULKQlWZGZ6st/nv0Xs2j/PKEBeKCPlBGIXUBAZPDzoR
l+zfX3DJfDzJ8IRsuO0UmNTOFMu+Z8BNeWa/W3HluEhkkLE+wRalHiKvUETZ3yK37AE5TYzQOK6m
LZ88mTo62sjZyFhUdGtCoTaA9d6DlCJT3rfCrQ9DHJI+x47fLbZVPvM2lnxN7nlI70iMXz2mBzhr
1KODteF/SNCih/o4Z01tWB8db1cKSHzZRJXJCWmbE/l68lSkIqB0NO+57mWAdHD25V9c8iZ5K5k2
ajuz3EGVC2LYmpfPc1HG1xKtwzAhFhM3+pd4yMU/7xq/owiWy5BKJwY0xNMBj+7mEXecL8gFmSYB
D0AnGpMAl6DmreaEbjefFiNE/EtzsXy4AonX6ZGMhKHv4B/XaFuTt+Q52J2Ky6Qu2UXyuPRf8D5u
5KENWvwPcNQGT/QPUQShusesRSLaaJMFws0cAoevb05b6HD4gKeHSxEjhBGv0OlsXIDEi0hL9kKE
pNQ3Fpp7Hv8WCaLRXwjAqUZq0z4nZlc64MgzWa18gbwK2nrbGYW7hsIukJk78NozHOsNHrnpmXn2
8BYUgyL7+Vj5YJaXz9cx7diEeQH2bRAR/b5QgmTpYP6vRafiajkyiknNJzjw2jVTNtcANbn/ywbW
rm5wvDwfcFemgqMHC09OpLF7v5EEStLOXP/k6EcbYobMroGdmMHRFxpTKvItdqxrTictsDexThiz
jbOt9waqGvXFovC1Rj8jHDcUqjdBAcsPiyKz75NK5LSX27SiJ5T7PTRux+fZL8lGFY3alg77H+Wz
Vw50ac3QSLuJyGdcs/hZx5T/CbmrS5nwNVHbm/gSjgEfYgI8e6ZStKtd99Uadj1oXuR7s9kKihOu
2QPNgGB5wCvoZ0BQCBxEOufZ9A/8ur/GkiZEnCNUWO0aJ+bcV29T5esxeBwJUQ/wCuf8I2HACUyx
5hHPEDM1N1xojeS4XX2VjeORrvRhNlYtC407e2PWJIgOt494UFVBuGg3U5wZb24IlfVf7rIygvqb
L5QgJ4f5rnksoAq7+HKQo3gXqG6y1VyGiU8xKhZ730vUlBmp4EMH4KkY/Y4JcwCIJQ9nG1HyxY27
OvXBOxpXCYKDT/Y2J7F0hHKYd1BaC0iJtvC/yRD+6tcJDi+dlLcQ3SMbF6KgvMX9ythMArsYQMpX
B8MShh4Svueoq29oY5bXu0uTVykNFiKtl0x2Whe9RDSM7EYawo986/NmiQLUtZ/8uI/Gd+Najce8
pKr5W4+zYJt4CtkqoJIY25aNXIeU9tbAchXFLVxw1N8UzkwmQQYkBZ8Uhdws9ZzI165xU3Nfx27v
G2V7cBGHPYf/XZsBYTgCSvhsE33wwHogDX2wMa2YtihXas2hFW1MVaZSvxtYe7XgY9N1dNi0lYOs
JfZAxvVKdPwA8XpOX0x6lHgf6uzPx8isokvyGCo+UFQyYFBRIteEESax5YAjxk92NuGeWAbsK6pD
+goEyak11/IDMsl7avTDVU2Vpfys/RZ1GXwufcxT+Tdf2Uded1C/XzOuXmoghus9dbW12ppn4GjO
8haiqEb2HQrDzKXbVyWNKVuz7RB8tE8pWHVbMF99ejDQRMfJ/eI8WyyMATvZYAWam7HdV2ZjGOSC
O/8FXCKGCuTRfxJy/uuSwiexrcpAfWKokyBaf7OhyF7an0OewKFsrAd3d9n/KF86NMgSgCqOOF7m
Gtoi7AXK5jl+jnAP9+C4jMvK5fPSv1Yejbd19de7PMqbFKGvDN1r8etYdCYpBrXAM9T3KVtSpwvi
ZeVr3dfEnZViskUte9Rf3Nn93qfdRd11fxgMit4q6swn+iAFwbGwMm9jtZNOum16TGBCRX7gT5TP
iOIw/BxozwHFu/Jbsiihr4c2o8lM7rRAmdt0+WPWs4S3hf21FxJiGrjKQxrtLYz2wvVulJOK8WQ4
ZR4fl1v+LmjRfJtrG9dfyo3Tv3d+xhbChpC9m90o3/mPsF9VwEHYPHp/0JeS4V1s7Y1FcJ429ZKd
4AOIMgXuNG2+Wqj0KgJUqddJhxLZz+eOwzp5ylhG14UW0UBC3JCjIhEk1EtUixNXialPliTfJ1es
YYYFqayUNPViY1uHbj1iLvWcqVm8tcdpDts0UFxEXkF+nLM76iZ7C4kvFmHHORYRPxkGRqGkMkaU
b8QBQQHSTRFQS7Ikq7spjRe5lfSgPYHxCEkmJH6cdfShpDhlehzD3104v+BlXnu/RgGv3Z0HOfYf
e6TQDmwAhfmFZEnbE15eJNBmmg5r05/oJNpAAHir0QyqdWgiZLlXJ6zFNePZTkNv55dEMn2CNolo
o8DJn6tUl/6Ciu29QzgnkStgaLmSfVZ9fprnjwcnlj+Ou1xzgQuocel6s0jDX7k5oecjmHr9QuQA
xGwRtM8Y7qm8QSQ/g+vTISqMuwR21OqRpxr9A4sLnbR2IUV/NIBA5qP3OMgw5SbWzBP0FuVt7Qbp
demUdMSNAlBS4oa2yZzQQy8v45CWnSdmPNVMIbv2c5QJxCfJvcjbVRV8B+BlaY2bsSK4lcugRQIb
YfMS5CptGg7iKrYUfjNInlea3Ajy1byG51Vqskztzs4U+A4/j0+lgd+0iogSreWAJ+/VTRxQ/qAI
t0iwyVJ+lVvJrTTV3nq5hhNt1JxuCFYNNSOiROQkUGe9QRrMHBZSi3tEW69qDWZMN+0Hh693b4Ja
uNjisTIIDjS5tmLHkJWIeL5UnmF+RiR4Ydidey0qODLIx8Mp8LgwY1FdAFK7iAFPHV0aJn69lMm6
mBPLqbzEIqKLkeFWgH/2bkbUntAFmLVMpEPDI+QoZvVZjwC/UYx6pO/Ub/dc4zWJMTme+fcMy4BY
4s/POZzG3dGUgXL0311QTNmafW+YbWUlVAudvLIVZJ4CFErg7AOf36eF6Jdipry81xhJfmrSONUH
vOKOF5F+9EtoWz5VG4mOpR90DSBCRg+dOt0dNPWCRBA+Cm/gCS1QGPKx1bBAUdXX2gk/7G25ua1k
CmYb/PnfwGaI9vITLHScMjyvGSuqiFHVAtqFxGeou5Ieh9fONCcBW9zZAL6AZW87F45rbym8eOOi
4xDY0Lqai3ezwR9gbcGMhEYmTVW5Pfek9xy61IKUpjWoIvQNhtbNTMy/raTHhIjdbd3JeJ4JOGgy
x1MgBHV4C8azrgL8Q/jK+7cKDVJ4DOUAPoeumGolXhZ1PAhNnbyjzpJgwQ6CkwiNkKuV3QQTJpzs
zuYo7SN5U6Ym8B7K59gp2sI6J5YelvXD7vLXgNkr2viuomQRfq9qkaZXTvzPvpBLx9YfbzE7P/bs
R6qYmmhem8xVIBiR7C7wrHEt7vWUImhpz2ANSNqGzkhDYxICQoFHE6NrDdh4VjVKzZy1GmWK18oU
tnu4PLmcJcIHHrKfEN/fEFhSzIJmeiuleozcJ3TJyLt+2y3HdA3R0bxoOa9mwsDiaqhw77mfZmif
/hI8g51KOdzoE8OqPY3YBd6ti4AYDZNQ9CibHNPuUQQ8gMDoMiwghefqF0wRQAjTMiYRo5PoBDrL
dVME5ikdswK5dDBZIwmITbdJZg4nyES+FyRoZvaePTzbnJQ8lrXBp3gCkX7+/9hPaScN7hqkXF91
2QbxQp6yv8SJwdueQkCPWFlI49ICFJIvZY3o5tzvp5VUw6saPjlNxOrus1Viqh/iAwpmQLZz/jjZ
3gClt6sftXd/Tx+/s1TVfV1eP8HfKuxMeVZZ7uLrkwyhC/ouh9wxnqwh8WirX6T4m/5qemD3qpc/
qWg+CwotkhXHV36JZDWiD2ybicKuPcJdl5SPZtOBILUr9B1DaqfUMkkz3MB7PbaXHSigrDQX8oQW
OIGRti/b+Y7UKrcxtVBsjCur902YYV7LNtSMGabbVDUcP7R+iasYTD6TLHYuImtCRPhzdjN5H+5m
Tcw/xvezJzDHr2r8hEPHomCoy7dtQfrmz2Ml5uQNDKFGnBrDk8nSCqF0gwK9xwcFkAylvJNu3KdV
iPcoQopMBpUAnH2uH7oLL7fLfnBDgNrI8jZlcDMupyWmszM4DIvv3cq/Erlr5F7AtkGFCRF5+8+4
CSEzD3v+fHFyeyS+x4spp2HAV1rf6GySYIDGWQAJTCCbbO7WqZ4NUaPC8vbN0RzGArofUyxOWSdN
lfOGXSpzWa+OCU9qFMaudqWyrBxdjPmIQGILZAAwFm3zCnfxYY1wv4KF5EB3xwaoFAeO+YGLCWRB
ft+e+7TSfw++WjWgZT33EaSY2PYe0pRz4ClSIBOxqEkQda0N+MgmGJGMhaUnwMmYbOZxD2SoctbF
f+MATsUiAXKmKkM39idM8D4L8brv3Q4W7yD9ZlZ/xer1ZYDFMuJixbkTliOk2A3vmYwoj19vHm4l
Ay7ROg+TanhGl3GMAGxBm4O91Qj8yar70gOjhClaGsdt6mucfyo9R7rmv7pEGI/656xJaZbibxfv
Vk48pAO80pRHsBdm43fow4mYQTx6AWHFO2PEA7aBcDrTdRdowvcPWAPC0AJCRit68htHWH++ZXp4
niNqzOf05G31pY8yQfKmywJW6HOOZ76M0aIrzHENBWNQWK6VvC/bTXX/890glvOd+qnrQVR4CmbS
V8nQQpTy+PjyS95Dz8oaJkqE5m5sT8hRxQohZ+wZdYNQT4DgPQUvJrJlSlcRPRUdL0Vudntst+Ki
pExAao7yOz3occw34P9tjZXdW/rKsbXhjmzibfPd/QxhWk2PZOgpsZgntzAGA1T2LawQAN+jd3Qz
C74jGy5bIYshxiwufFu9Q4bF4Hh0hEFFs/PtiwbeTvjDB3mw2Enejt/MH68Km+XFpJL3+CpIMdD7
q8KwToB986MDWAx4fzg3jrl+2eGxNNAdoBd2GJd1MtRh0o2RWKvG1Pxt86wLQaZMjpxs+UMeueSC
KJJbRoAkEf94exkwRAmTC27U/G+YER46E+fT6RLl1AOMQkC8NH5C6Bn3suLBJJlDjou7rmTUBLA0
nx75KbOkSNvvNK1QMoNjuBMJogqLl2TpJUHO1bkuoaIhyYB1gsEAi0I+mTwzuoGWgvMn1os7t0qL
+xE2n2eqHy7mqsVSJ97fTMLthVZ1OfoZyrZ31IoaPjYRTU1X0qRoTuTyk26DZ9A5ezeFonjLgbnG
ok0vigRma4SPQBXSNH/q9wSGG6eQsBro/2RT5TpkA13Z+5/AkxS8KkuvjHcAM7T7ijZMOSUQy/6n
UYDxGE44UV3+yO1xpSY6M61jOHkzg04ql5isLMi30PL/rBl8idcLxHk1+eIhlYlY8KSBQOFnWCnA
zjf9TrQg5i8EKOLmlUF4WJznD0YX/DnDqpvxDAjE37Hbt3YwZ6p6DoR/t4x3o9nZqOHMoi2bvj3e
EYELsiXCNgiIw8XImemT4lizMTBUCdaVxj/NIjoLeQ460qRVS98kIf3H25UyVEVjCTq0Uxbqb9fB
kS8IJnqZVuP3Gztm3Dpe3iFSRqHtMtuycpIsaCCAlv24gugyw7AJa3FjbGtS1S6prYqemjj6K22a
plofnuHRI7HhiuKJa55GyYnol7ZvFJBNYMNzeZc+YLLUnVdzAai7u4IcK0y/3Y2Ozo0AkLCU99No
cpISGhrMsboNetVBRcuW5fpZW/zalkojFkw/tN+aD344XwO3eQ+F4SFVCZPpiIhCDPeKiOoFwtLK
DcVhIQnClwgsjpUOtzNBmQFxK4vvCl+bh2DSJ3j7JQjGVwEL2Pshm0K0n5mlsPkZExWChF2bQKky
deeDscuab74A8qOuAcRTsbQcV+fORQib3wRpT7GRZH+LKJgcRQ4/x4FijyMedq50QuXjaOGSCsU5
nAmTrngHHaN8zshFk55oQE2IXKHzJo8G/aFiztxfiFbyyoJFuwGL+dUoxviIfUP11WwjfwEt9JjR
fg0WwLnBJbPpIlrP6Av6o+opI+arilP0AzfKkTnahGOYn019yUuTJo7fUVIR2+RYlVT2Dvf34R4A
kzfpCLOZF1KOQ+hd8zr5mGAOixCacBDztpsMzonic4Qc9+l3XdanQpyJv3pxCUFT1sUM5240zVLu
0JRmoG9ZdmPe8Ha0XR0g2bCK7Ye2trTrMGjEmiqNzef0OGZAbRAnpYssisA8Zc0n4smX1DfzwTUv
zTqki22DsbkYCesZOJ+RCDv6GQqeooV9TIoW6Obp6v+9y3UFCNT55nl5DlPpVBko1WJT+XlRjXfF
hhuCsq9inaKhWb7nMCMfrmMiuZtzOtjt9kX7sPLz8SmGr/Fk6o07cj9pGA2qm5PmqkxkTRrifc3U
uFZ2ctQj0iUG7TULIB3z00YWwdwygTJcwroFC0tbVP3CIxR7MMZKLvN4OJRtI7jWFmNnqSC59/uK
29XMoofJDnxoTb65YbSxVsQ3SMGQSFfPgGxGpxqq1Mi8j5k+Y5n/pRo7YiJ0GHZeTnIMFWfr5aNs
A54MHmK9KMqc54bNkcGmZXRvIIEGGJtBdwVsM/AVwItjiHelrDWoFQFYrb2lHbJfNGxuCV+hCvDD
h+/5cykZWY7hhAJ6w00lCAe/t9G8SbpWajzxy+qfyPydQ1rZ1Q1PcyBAeUElg9dCbJgrNOWdzKcz
elJn+Owelbyx7hho6Ivx6CvAvdqVdmitNrg0KkQOzTG3DVKhvvQPKUoJllX7Cg4yUcn4Y4k3Ww6N
cl1YcsONoMnRzdm75YyOxJe7vhZ9xSH/qTgw/fSgKgxl0oC8CDJc7EoZE8curKnhjnjR7NzqTRWQ
RvBQwb1WxV59gvuN3yblAaFxNeZnePQXXISDcFFmq3EM8vRiCJAbXfcsUSjv5RWHLWSrSiOZ75Co
YllyqaD8lsDHNGJqKbkXfJgXokwfYnPLNPU62FFk7znbTGTiquVEmM05q3Jvd1NnabLFtW+dtazy
1Gf+ok4ToEi5QYlNy5QyYd4JKSyPUUyQuadHsOJYoR7ubplBz9gDnYjvWU80zsLieObDVTdKVXjo
Tqenos+TjyQSjBxsiuetnwUhuvN71utZanbS8z4lCQrhKzj6RRKUqKcB8d2TLdvuGDezMd75jYND
gaLDggs80PWeLI4vp9qkisn5byQ3YHUFZ2N1pEVnRdsccAiAR9GgPh97ArnXWWrYU01iBpU6c6+0
I2h4ABy1Nqhkb5lEJ7DQ8YYzxpxpmdC7+NXfbQpEdXr1cFXG8UVh8Enj0Eujkq+Ho7pJzwsEdkcb
bj4dN2f5IjmzDdJ4UZjIVIS9D+gqyjogfOFH/74KjfIF44qLwqf5XW8nOcLYujKn0rFQ+iE/2YAp
4c8WCKm3+wUImtpiWhrfWHozZrz77emg/OBRnvJUWfD+MUWPM9TADkaIXBZS4xV/BRPcEM2YUCCe
fcCogocm9MKNT0hlwY5F0n8McPvUlUK6P3WTzK6TjcBoqL8u8O+rFWkUJizkTGkb0yuo9FCgbMal
3gxXKVpN13khyesGfZyAp0gGWx4HwZ1OdqtIDjHn9YUryM6h+E67kOnokzZIy6ZAvgNy9zxzV2tQ
epG3kaELEuESCIgCKYgOBEX97vR6GFG9TA+cnIv66vGci+HpwNINbHp+Rj9rotCbrQXGcIpyWWX0
bfvjI3+n63UqrP4EglEJEeRk1RuBa8tQM4rzvWsvvAuTUnRkWRPQyEC2uzFhuJXB5n6BXrDMOIC3
tQussL7l9YGZ6jF/ESSyKJp48ZG0HRx7UWZ9n4hQdq3zqw+dvE9IQCXxwMz099+msdPjcDF4jfAy
lPJzpkVWl3oUYBqed0cs4jrSiUG3wP9Hfq/QP4U1f1VyNNhhQ37OvXUlQZQfVnI2nYdAIPWPAvPE
CiJbdoyVz+olpvzT/yij2cYVOkfbsS2a1tGT+axrL6cRpc+mg+nJqkcc2P9VGIy3ifRLNrQRj2WJ
0spbnIXiEothdHlc09F+nIdMvCVkn7Klk2kAGTNQH9+tfUf9A4IwB9cstJdkAyLlm/OPn5+ydS+0
IFFliTUqYppSSniu+6iE/sAZlJndwswJZJc+q+K/menSTMxofbmfYR8ElGqAa4NXMtHLqs5BTWFw
s+46H6NIwIZ/NRTSd6mu1GoXeYaZ9EO5m5ls9iwchq0p0ZUyaco4cwXCyUBJgG2QE2U/DwEOCYmy
F4khnC3zqkjMAgM4QYvX9QOuCfIEYadkxhEstOI2eZsfN+e780r8LMTKJtnWcqLpJWThFc0/rU7M
cFEPdAKL85YVT1cEUFgIbXpS4FeKcPwymuBT/LC6ONJjI1/zgGnirpA8iSYRG60+eBPgwnlUqhdE
kGF0poBV1F4tXGzkS0Cv8G7iGTRLsQwBtHMvQ0U82Mq6sWawQCgjHmJw8ofWDsDZShxXXxHO9pLq
7X/ctL6KobvwvpDaBkusuqa/VdQcwT+V6Zyd1j30Eba5g/2TLl0yenruFe0gnnn7pVLku9Cj4yNA
MU9vL8pgkYEmCJOl2z2XkKplxXkhpgx/vq4olNI0QM6IGE1w8gsMqBXR82oLtk9RSwAud9NxoIE7
M5CUlVMZiec/CIsqwod9eSdZHCL0LHnzLFTI/DvlIMQycCdTO+WXiaHoBf1PcrqDODbBHWRl2Ea4
a5eL376aGRPBonZ8wa2TDqZrUT1HrLXjSKHBzKRFR5fXWaHHUBWJiXyQZOaQtQKWOMtNuw7rh2yN
F8BRqRLlxLQ2yzZbCMwXiM3t4cfDPA/tfgvCAkMIFmmoVooC93HRpdSmUHrps+LdSC9uh7MRdHiB
tSx6AXCqG8AgsMFc8EgnsWn1GWKddjQxV4g+40rvI3qR6egWpr3QIIt7F3kPiEotw6zWPir/JyV7
NvnLnrdQqtqpcWmagsLPjGaT4ILYMZLG20/Hp3mcKkXzIMVfXYFRnSgvpHqBJ/xqiCz2X8eDPnEb
zxryFnXlkMZmQlnRxYuADCHTVbveyd+eY3IQILreO/0fa/XqUZnewkzP9b050Tsi3g/s2qo+CV1k
1nsVxgyT3fHizxE5sqFXmT642ETEtKvvfCv2uyP7/dbGTLnKnOhTEFRnLbPMc1rBHulS8KfFNG80
NZY4doLjKhhxzpEqNs0yQrxek2KwNmOcniyQN2OEiDfsrODvNYqAaZF8QpI7eAGe4sthb/IQ7SKh
GaH5e4Oq6ZW7nwSjVjwy/Ox6nSTvxRLeCAFpExXWqcBMxrZ0+eg4pnrpzHxzuSRv33SrqiadFetk
DW5cXvDU8SzPey3pSfR0uw1fXkevuvY22+XlUtq7CUDYcac0gjfXHy3Vc4r6Ixgn/KM/NbZXfXDt
a9qVkDmOHFt1awfvSoYCG9iZBzWIEOdgBZ5nr22ftDMdduknV3Z9bFaL87dUu4hN7v9Lbc2RHSPh
H0Vhy6DCkDF6/h2xHxF+PtOQY0cT/0Cr0I+wODqx+0YboEPjJKbQNSuBURTKD4l0DJJtoXtI1Vlg
cp1+8MH9/GuTqmLM6HbU1SLg+EtAPh4bLQbxOfBobCDzgFb9ZWp8HNSuQfKorjzcJeJCqb1jm4De
AlJa/2ZIXcZ2cu1JfMXkEwymzUo0zMQltwY9NOjy3QcEQejbqJEABKZ87Py/ID24sGggqaC+iFz5
vST83T0zzx3g1ry4AGa2YkyNRaFV07hBVJ+DKtg0uclSgumpWmFP4xm46Ipi/B+WpV4zHDqtbXvr
E1Ja7CRU+ufiNkln0Ue9T818W4FCUkUATaMbMQRUL6NkUlaytmMBI0BwPV1T6hEDsb/RdFmp0Ttp
W8W/ejPEO2TwKCBjjp82GtOeImW2D6FF6Nwg1wq6nMVrIHkS4zqMonW5sEySRm2QZ6FmAxvAx42/
EYly74gRx5SpFyl74MI+a6z+aJ55xgEgKauWQl9PURe4Ch6OfHYeb5BjxEOXqaWxvg6MiABruVSa
49yLOcyCJi3QXuleTCjxqkcSWkv1jOHgT4QsKm/6OhlFMCisCivkMucNv1nDc7rUdR7t4QKSM/x9
0s8UE8ldVhpdfIx+z2zMd8AOdWget7cC7XbO26yDmbd+/PWK5evCZjd+LmHEVGJiwoBFHg7/0AYv
ly/zAp2wPB6m2ffwEhhECDfw0Trk492L4loZmDKItDa7apLO83tMCjNUhTq3q5evQUZO07+uLr8U
TxoqZopR0Jjc7a6j3IlPzcrLAdKGctkNUb7t/X+Cvi6X7eV5g3gC5E3AP0HXGriuG8wVQhrq1c3P
gKf116BQQbDm5V+WyBnwQeHD+wPauCgB2iRsh83AWzFzQX7OVd6nm0IRZA7eCVE4KTb501VmVGsL
5NslIAs6kCQpB6qA10ZUVIvdJ2QOF52F7QtHbXgisC4tXK4ZEiREWJvZI4RuGTU/0/fYRpsgdLKJ
E5M2abOHSB1QnojE0Sb1z00Cl4M3+gV7ykd/e8r0O8EWJ3W2zc1+oKYUSaFGWJdE1W4C3Ladm6l8
LteczZBGF1mkKzdm5bz8uaCKZuir5o76gVTWTFZ8PBfKasFFsmI8fGkejVCjUy83mks+S/tq9nJy
6GTw+QqBI3AQOS7i3G/J4rYIyz3AqsBWnI/Du69VaSBVkHU/3yYJsr82WVL5X7d0+38Gj3ISLtrQ
ggdJe1c0/ObiALVEnoT9tiBeZkHts1TEEXuVIVQPGZSOyxMrfBR3ngGG/L3IG+Uxa4PaW36hfYHf
3DAEd+DZWesCsJjNH9iR4A0PkuEvt33Df0rlcTKUSm535dMaYqgEyMUIwK+kRDr1mnn9Vt9x8Yxy
SM8fhtvKIhMBfGhHBFefCGWOvOXWxyp8M3QbtQNbGddXI9XawPmfnRFfCYJX53eB0u0dGL9dDkQM
RdWOP8Hh+oWpuoIvOSIZ4jPkf8yG3zPeykfqcl24hzyW9RvF8h9TWiadexdObj++DJiiRQcDBQBr
yhKJ7am9VcdRNWMIydzztq1LF2C4zVxFTnUMydxI9UdStXgG+lrCUh+tV5YKiXCUhk3w8qbpETdd
tHj0qJOdaWFKeuwcuJCFTid1pU5aKlQ0JIuTRNgUVjzU9EgPXo6ZXnCnEXkGt/O2o3GgqopAMPxQ
/lPMf+qalgqGwSchqWefGI/R/1sbA3qdrY2u6CiklnE1GOjiWlFH0lTWTrLAevns0G+OgsuGoWIy
aNlyTYBD+MeQL5gzVwIAtnyFb3qH8njtN1tubk4XZew4ObushKnaHsHxBliQO3AXwVsKEMyxJ/oF
KYVZs55Rd/5ZWEoXxqT3ahzN5XS5YqF7sP0jKxoRRlLDzCSohFzkBOi3rVxbtp0QG0MVlIICJ7u9
wSnMxVArDwX/ocgU+oU+DUT5pcSt6nAy2QxbfBOObxHHj1M8iGTqKpZzPRueDobdJoTO3bfYm2/3
IODOPcEh9C0anivSQRoBO3EQJmrN6PAUCdIxTG1R8vVigVA4InrfljvrR/d+J1Aodt4AZkSEcR9Z
CnynF2hgw4kTPqHeGOcJ8sVCDEzY6+ui8QesZKsVnZdtTj0Jga2Sf+xTKhUp/COY8YQmIFzMw88j
AMJLZxScDzBA3h/V8FiJs7necaKb98N2I/RXAD/1yw3sQ3AFUzPqemEDDHiUvDox+uYT5mLeZuUq
wLKDsWtu01xZCfJkhzySD96Jjj35h0eM42QKpjz5DtnsHu+QtC6rT2opfg1hEM8Qh2is8UYeTYk2
O+99WOBwnz1La+zLPqPZghDbvVvtNa6WAxBQuO7XT1zLhVysrqwymET2iBwW+aDszWzpKhr1Yezl
hAkyBvVYC2SD/VQ2U/QKa6tS6duj+Ihvd/nXxJXs0EuQgo5pwPnyYgngsUNK+5f/+0BUjrvmrKf+
lxcwBymN52pTOR+Ai/M9nMsS0lr3qaz86HuVd4vQKQejzWmJhVz9PSdaVnt/HBZtwzEAhaIrUyYR
626SDyMntsgIoB2SpEZM/KCqllC0OR2RwmTV/A+ko1qm8rVoustxJSIQWsg0YzWMnHhXIHt83Hqf
ni4cU5/Q0hnRAnxXK1UaIKeSr3E2QoUDSXDUcsPKtHJn+ZJxf4tinNH8ncDwICZ1lnTKKU0qFScV
wEx6Qx+G/EF4GVt39W30nrYZU+GxBu/eP3MRUVtcoB0VOrmnd4EhvvlJhS6JpsalEwBgqHZEPDlq
vk6xbnaiePXkurNW1oeLOuYXYK30kF9HpeqWRjDMpn83sij5o9/DmR0Mav0sHMi4VQZshB3uWuIX
r+QUhYZsvffzqeXfpUEkQ9FBjTU7zX9CVz/c/JC6M+fo6pbNYvOP5zTA/Z6JssZRB8H8Dyb94GMX
7DS705Tba+DxTRzj6ln66BGxouLDwmG2PRGvR7MBcX2vx/pU6d6AN80SRIfAmZ9oVIEtMJIJW7Rh
n6R4y1FldD52ayZSYM1+19soVAW/sYksv0nKuf95KbletdgKpBqLiwb9MDeL5rJGQhQqm3dvrRDK
1KtVEy0hsKFnvQjJwO0HrD4Y7+4GLJkmUCcpjN6DAjEpD21x6Xjyyewuaizv75exCx9WVcRYPP48
yxuowTuhXXLTqhkvEQqzVf5HPa7rSh9rWERdtiV0QSPWLrBCUaYBkfTcgMbcr0uQQJ2t2EHJNPD0
lKR6yd6GICvHTJ226Kdl+wrNGRQP06EXX1uMcWLc4zomJLjDY+abzR48FPMRqVSR7ucqE/VpkXsv
kJfGeGYddnPcjeOD7oRGhEwZxs1cCHrbGajN3xI1I0H7pKFYhUKt1e+Y15/yLCzVj7mICajVjMaU
uG0x994ps3bc6NjH7WpYSArWQnTUnqVrNkRW+WN4/+MI7ZNKLlk6tz0gKRyZ1krFtukogezYoq3Y
ThJLqDTBEMgiThf7r7jbWAhfnNW2vpx1xHqnc4Mf2ODWrLoj6/0qNrD2frlwfShegdlPLRtrF/7P
lGgWG22HCedWHO5BohStvju2H9sJCvAGtDcND9SuYRwmF0n7cVgIcKSIHOJGzOBrnvJaTm4FWZ1I
YDnATHZz7xXfG5QzWXtRlqg5lkfRDcJ0sPw2hccMwZ2sKuPCweu2SFcrSzKgDXQSClJbD0tlVOGx
pysIARoJYEfn9W4PKLDwkjeTSLqHwaJXC6yA3ixgukjbCFrHW2T8pEP3MGj/7pJaQrJgkOTyAUQy
icnDXubwnHFJKyndZqOoq99TmHPZ140y2FhmlrgqoDMexfEMCEmQiVGvKQArcmDDLal3oFwk7amP
7oYALIfzWzpzGRp6tzq1bw7H2TRUNMIz00izfNw9EP5xs4TW698E6zYpjRk/MCP7l0nq+UQRWrHl
KFWATstkTq37e185Jj57hi5kbeiYZyf8Cx1bKLdUbqY83eSRYnPxpg4QqgdSf3gJepp0I1aliNOM
urs3QMNevvwGRCNVDSB+M2g2GzDtsMEyV8Xd6x/t2YNI62tkebbGJKvDVhOHVpisT/LH2McbfUE1
fwtW6bdKx8vfZFBBFZy+ODWz9DVUvsgnPWEWTZMfuRPOukWCZEuZh0UYU2gisY6MCiryFlSSuPZ9
YL8qEJFIc00NoegzehiNxFtnuzVinV3PczNNe2WUm6/tGXcPi0RY+qe/+2QaHjFdgivP3LIAGiXA
LezcX16pMwNunrw5J2s71RrpPlwwyDnL/xgQhtG4Dd49UwiDhcMmDEfL1ZfuZY23RhBZD8zjGEoV
hiJall+1t9u3KF46uJmjIGRwGxACwmfzavF2LWDkb0UkbolcQhWipTJkyGFVcVHigUT0EyqJ5L4/
kaCo7RdqKoL6qgFPOx/gPHlrNM9q4Tcn8+HbOrtPkLlcofwWNGtGseRmjz9+7XG2lNGpKGMpLGwj
lCeChSCGCurYgwWU4iQtLrs/Z8VaDpjt7JK6UjY6ClTkTicPmluiwRoKt2cHhg1m6ie8iI4ExjYA
meuQFNZTk7KvNJFmY9S2Qz/GtwDyye6+66dmQpBmUE6k3M6ULOa2uktjJdfvzvP/mkZrjzAXnxhv
xgkwhs1LvLCnhNGNYiRoJ1yMNqaUwRWmwUmdtd2mrwYGk7Eqx6GjQmd6hgh/EGedDyzBEGBn46r2
bCjEjNj71WTrMzXVsgUQ3LuZHW9T0lkqnPc2Y4qqgwtuawCElmBFxkGGlY6LiIpKS7oQZiH4SpBZ
rdpeUaq4u9P0bzwP/+j0XPRf5KFHqqonQzv/0YUDtzM3TWuE95FYo4lEPrOxnEK4mH/UzEUrgEb5
+SpcBFGZiiW2HUISBLV9GAGkLnW6jQJ6EXnirvocQ6y4m349dLNazEzF6qryriyGhR4OPnhrfOQs
/ojZKZsCqoYp5STJ2kYhaaSX5nEUzq9mAEm4Xec9XwsoXC5JmdxRgQRLJuC25djOVMdEt7d0kPr1
I75nTJMDrVTWoC/bMEhetMH7fX6SjJVZpKXlRvk9jqOsCFFrcti7xlNxE1BtgcAnlTzJmtfebV/p
usbIBogcbn9Zd8yVg9LgkzdvW0X1GKcC/e9qGXRAF61fbOZHaCPn7+R55JinnfpGhvNFVd4c3WHL
d+ZtKOuw97JUPfcaM4ohEfdN7CDNJY9PVQfTfgaMROKWxeg0vacyMVQe84epZDBNxTQkcwnNcqNg
TrlSdw8P+GRYvlz/xYju5ic+z7s+H7+LdrtI3uBB+8GRyksvkI4JktWS6fVDXmtRKiyzd4/a/CQR
VQUYrvXDpOLoJIhligPAPFp+Xv6yVuvH+CQ845jD+McI/OatY8/dxBROTk7FwnvXrA7udsvnGYEW
rSj80Nz3ite2knBM3Lc17t5fbkIFhYEBBTN6wPhkcN/amQG1Vj1Jc2/g1ImIkjZ/1nsjztbwZr1W
4cJ8ZqjAUXy/ieumIB3jlWFstrhG0sHZqNyxUpN+IVFCip5VIsoxODasxU7LqF6DE65Ty3VjmPxE
/hSy1jdx/vYopaSncz1Kb3qnGJIjxgtQBxGjKvPp3j64TbBHjkFmC3Q3uBBv3f87F9bsc7XtxJMw
nENSxskGXISADP7Xf0c2JCOFQyVsDUZolywxOlnDsA4u4JebcsN56gSWuMcaASRNXNsvJiE53VJ6
Bd9Tp76k7G0TvJIH695SwqdYbzPKWKS9QzZmaevonXa8/p9P8U3bG/+u9ii5ir+EKwn2ROUJYcIT
2LQfgGzFjiyxgYWwGFZaEAFEfbzG9cF5qHRnX0SUKGdlY6VG4DqqJ83Ki8AqlOJ/7e/erZdggePj
EzbliBQ1mUXdYaQld8c5JnhqIG+yTMiBdZEMCS8Oi/Rl8xZXMj8cPeyCfl2JC9HAAeG97RUzoqrJ
1SdjWPrfkcif4twXrO9tLSlxb+jDx69Eoq8DizuDnTHELB2+irXFFBW9DNKe/uw8XXu8KT00Dqke
2Ud1WAGOF/EtIAqwtGgSiOMfLVcMHxm6goJZ/56FpDLLM7cpbyBadDTsxUIPxEwMOvwFEqBBGjxO
DkF9q4KoLEWMrrkhdZKyw7Ljtuk+0caCLziOHTYSM8GaaSkTr15gey5HTlPOt7P9bbCiBz/oLwcC
Au+LRyk8imuHuMtPEGhFIhXAPFdBIHQreg1cszPzKIbmRTh6Gv9np3Fw852LMYTf6UimCoQvrWf2
/+oYm+DPC1qt5WXpJkiz9GHNPWf1UHB7JYk6QqTd2k0CYEoAYt2sOS/EfHTZ5SZVZee1AgmSqsbX
k8LrVVT2nz4Qg1xKIMFzHLwNL9Si7X1yKqMxWzut+nCS4KSgXs6E5JFCoA0xhZY7aW6ro3WlWKek
wiDTMIFZjiFXm83dzbiGPa5JxPqFRzKnDVU6OgrXPIs7Wh/+7RLob6O8vzeptwGkVP0KZc+QZjEP
1UGxrcNhTQ/WtEzle/hQNB73I36q480IW5khVqvlUhmpn3LAmYWNEtjb3qZLOACagDksir959tM/
+GYbpcLyPeOra0zFIMNZMk5BmVOhPUFNaK0wLduzemJTZdx5v7M82sSJmsEyWpE9/zMEoHow1/ZD
iYIfWdPLCFe0TBnvQCsb/dRw1a69cJ8kI9szvKCJ2S5JCg9RzgJcA0vpbIuTE0C02NwLvBUrqmft
TNsaCmwe5WjR7W1u7eoJMbQYD3uUMe0aLjX3cluCJz6ll/ZS7HJn/iu4XKdYgp71KrEoUkyY+oNx
pA64PqMgC0UKOuDdV7YFlnsyEfbz8nt+xBIJFLZInymZE2bYebwW3qD19X8g2Nx3jq7GWNtu95Tx
aQNrTANJEkZYlQY619woE+LHQLNR0/qYuy35SEbruYwTjGhQ1tVQlQkw1w5tg/Uy9pdSPr1NtU/n
r6T11RjDBphhNaRONi6xwKFBNrPEC1+CJ3HNrc414E8oJuT+Tmu8DH4pXU3VjD/o0f+IRIYg7Et6
EWLTvCPUh0BTQ/Oqlh3n3GQWdwuC6qCPk2ULXfKADCZIsRG6+QyUy4TA+lTOYGwQMecV/7yXtKiT
4Gzp+GctiutujKjzr2K5dgeUMzmGC6nZNPFUPhKsqTfX7mysKXaj0aQl0FhYsK/vwJG4WtT5boEk
XRNdyGJLKnR9n/uIAyxRcyFEcDWvPEOp2wgMpfMNKVRjlrqbMbpPmu2Shn37g+HxbBNai76EAbN3
xbmncPsNZdsqiqwCRK0M5kNLYlkEG2IqNrJUsaPlth3TGfOdKYD9M2EIYPGazmxe03I9y+gFWq+D
4rj4TnpYfHxJkNiCG4Leva56Q3RHVJR2qV3X3u/AaNtIs169YvmEZaxS4KizUEBs5yk7uzDfO2t8
FxnVTx1eTrS+9Nhd7yf78RXBuPNG2QMgADQWHQ2B8rqrK+FxmRgNbcG69yvXJMhxYaB7Ebmdet40
j+DJcCbhbUuFU+meuYcom/TQgdbg6/llaMYkCLjfDpEeCBUdvh1T+9lcOjUeFYOP4DoKrJBGYOFS
85tLPj7rJEOgMkV9ktyNyzBV+Os10Am2hGjfaBGYJzlK9mcgwgCH/1wdQBtIDDqE7ru6Dh2XRazH
H9oGvgwg8RMsUEcPu4ShfH0jVBtS2bce5ZRErqe04gCJaxsPJ0gQb7/Ggk4x0S3UX07HkgaY8ABf
LTQFgaMWeIxfKymGt607OqozLs/Q7kHSeX1WMvTwB5iVgC/Pfgj5M0jOLK9R6swqExFaXgSTkX0p
o5QuLEGgTsuKSresPKcJ/nOQIzglojwG4ofxf1egdGkH08CCPWW27Ow7+ONjBDjLfmi8U9Fgfr3u
K+kD+lH+tCyGbP8TjZaHhsbolJ8ZBixHCeKVnmuFmdKh9km2QsjnZegcSsKxQFnZuxpc2h9Yqubn
Sk92Qpxg5XNRTUAkqSAnmZdvFLqt4UR4arTO71j0OPtGoFNOjkOFhURQO7aYNdR5ppQFAZNXnK2r
IQHCox69iVm73AITGyT0KjJZx/B8TH/OQF8rMwyywuaRnj3G4gVUXOch03K5HjJJ+kbaxgJX3Wz7
IaembC4sbyX14BPfwsff3m+DmhqUt1+Dp139sGNNI/rqXfJW5mPv3av5O6bdqVOgruPGEdyBomaD
tUW/pvAE6+RyAY3cR+FalSDm+8+YMzPNUYvwBFoZ1pLHTuYWrzRFc8WHOgvhy6OKMajychYzKHo2
gKx/D4EGHSGt6Li7V3BxYoX1Jon/URG7kcJS+Fc2cbANP+neEFedAg4AK0RcXyF5+jCgP2kouUa6
AxzBSlZJdl7GBJ1CS7RoT657h63avyXmEcVxl16CNCLyiQ3Uc0b09cpmVjVJo15QFyXZJWhfCrCn
UyR6urdsJTDGl8EN6rNn75NwTqkdu0gItVRj8aO13QI2znWtSlgpwMQewG5QXWCsG1Wb0SVOZZ3z
ER9d2qQqutfNLdHE/NtSazAsIsqbB4TEgXDT7AUlDNB4Wfi8dewV/ijf7OIA0jkSvmXPIDHKSwy5
myiT1LSSQOSy+BVJuOmjWUli2CnnQLs1SzZ0n1hON99LMDDMIRKQ2btgLKAaXvCUC4R7RIkQYqGa
MUioI7LueVtFkLpLsjGkvFv//CVUBivQ1PmtjFyqfK7jWnrupyfRM/skDeJg40AjOxGsvPmImRKC
t0PTnTEMmkxjKdREhjRY7mbfHnvoND4f0L5iXGwEuer/jB6LaqgMoBGnWUHw6DlLGB9pGjl+76Yh
YX6suI5IHI2CC3rqNH6j9jHFtlYAab7yQA5kQg2+KA+AVCE4rFQjA2NCIWaOlzFUnP2xQG+4fC5O
kYQ8iBH+7UGUQIIAz5da6ZETmiE9qeP05hDg11LHf4qbdL7X60YYJThhyMZOgPVvfgE++TyZ7yhZ
gk8xtJBYonxFDc7JNwU0BSqBlYsL7Cmsg8N8sTrTKYcTYgQU6CMECpYfy5lYyBn8zoSUvlT23cRL
4205GpQB2IfmH0knGkZaMR72C9safJhQamZ7iBEmJHOiIWfcJyGQCwaiCg+jAuE4puqvw03gXBO0
OyOBq1K+hfUr/8L8gdEEqO0ZEe4IR7WGaxVCFd9gbdZzUeTZBHEY0TOkG0ihxL84dEvITrC/37tG
btJsMMeMCYWy6gVZmyvRWGXkadVg883X9GuQGZ+7wsBUlVf5Dj6k6whoU5tdckcVKQd/AdFpgnD9
fnMvyBPmwlqrWDCqoY92756iwlr3l2fVsBCJ18vUDy/JWg8Y5ghs53ZU1BhRDGNUl3d9q4yBKM7D
xQkY1VsGO3sULi+RCsNrE9Mt839rtx9SaN3xAJNt4tTnu+BQHlakVW0O40kaa8AS7Lyie+NBIVnu
Dkmu/DA99wNdOBColUFi4qcvUB3LgfLyoh/k6wP/daleoq26p5SPK2aMfYSzeec+dHGMC3ZEGXVk
2OD1Q/sA3P8Ch5GWPcbQyMPSFTT90o7233iVdqW1V0ld+yw/bM5MWHQ/KhhP8bdBctnN9ySnDdp7
e5OQr9i6671N/1o/qg8ckrdMz05MriJOyz3ebyYbaRJyBWWwFTvDfG/JQ9UbF5OL7n+mIyfrlPFI
okaYP2IocDJ248fAqW/77B/VDrBPIOadVwEpPDhekKLkSDOMNdKAj9LVJTEMudPQ99VF8vre5sny
yX1qk6GGA4bJL08qumfPItkrkUbMvhDWcdLq1C48kolKy2bGccX8Y2CE0DpzX0I7kw0aYLNNMIB/
juNy92KvXll6TugmgQL9Cb2qasUaCkO6yVthurQGZqx4Bu1THy+BBe7f8gR433EvI53fw4Xb2a0N
PSHw6cGpSUca27HPjSr1V016W9DMlFn94x2OoPNvhmLFrMfYEk48NRk18KkK1OmUEpKsZ4svjIif
v+MxFjmWwX7BDmfOPgJBLQejmpXR9pwueIPd1HLbcaIWINI++aqn7XeBp1JVo6gMV9cv+GIUZ90q
joNTLibKjKgGDL5IVymy8a92qPnfcuAL03H+C5sKAL+J59W1dqApARTqnbgaCHSoJNmjTZFDlHvc
Z1liU6WYMGWPYnN2uCOnJS03WR83BBcE/pbMx/z8V3ZABjhnnKIJqC+HPo0m+tqlaqLC+f4197Nd
84gwGQAlv1R+8UxAZZPR+HYfnyzO3BC6Bw7WUueRSZTiRlI27qQP2aHbYpqx7K6gfV67T+Rnm9vT
KMZH4JEklpaQhg6htykgQ/AvDPA4nfNYqdx4FXQ5vP7n8Zyk5qRCCUSPNhbCYedCtyqmZbRmSLbq
p0PzlpLrhNzgHCuKJc9LdNqADgE99agWs8h6ez1rE7oa6S9+yhPVgKV4lDA87q8mP4PW7yv2+7zW
R3QVa8uckkmwMYr/viYqOjE/o+N2kPR8aFt6k0BOUA/uZMqwX5knbMuriEK+6YoMV5dwls+Lw2sp
/o80FZx3s9UcBvtirihvN4RcD/nEQskOIXlGcT9snmvaesyu9eeE91VZ4b+IoDsIZyQUslw19zZb
hzbnXO/fwbxcnFkv5Qw6/F7w86XtMv7Ie/nmVtbND3TaQ2/Cf9IEQYLscZSfb9tBnfl9koxGI/ze
6+pnOECpeprKNouUsv53lrQ6N966SdC3YnQXCMw9GF3oHjFn0n3LfLIwiVJ5dk1PljMphzsqr7F6
DMzz5gaFxvHskAmnDgLut6uFcM6vq+xiyThAUYf97vNmKFpX+U5FHIGYsoXbbDqL/H6BmDp14hBP
lFNXfLdRcM0nywNvUrS0RxIXNM0hPUmYG5uKwEwJB+O1lAS5ziEwe2ZnU6EqMp6jzCRRgHMhGy7q
T8dntR0cCgAPJhAjcR+Be0ZNzGo7CmVxx9Sa+B0ZMcl4WMY0tjG2Cb/8Aqiq8yKBrA/tDL8vpXK2
UbxGotnfZtqyrDN7mCR4gjXZ2c+xQW0jPW6oozUmVCB+jA4BhWm5q6V7qLDGhJRNz2NWJbAL7V1t
TO6e71wOzYR46tp/iawYkTZR9OCzdDocnRr6OSu3XoLAYA6rjK80B1rrnJOFjlD/7mrsvSnarMhc
nyBhduejcMWSaPfTJX5C52Pbp2kcyN3k6JH3763Sn55vrUdXsDojYZNaE5be9dnocMpVbjRK0hhv
OplEItivlnD45B+5eC/e4d2Jx1Ns/YwOkB2Xel4ARLke68WMWab51RtdgA4nV592xQO6RID1cSdc
KBcYF6TDR24SA1lyZmkerlXNJl5D2v4no3TltcUPkH3ja5ZAQq4gHu4Idqki5aBorwls9JHWWCD0
OPH5REz4low5tFHcb4wbaWGX6vNcfOkSXlsgDTZO5Rsnw0FqT8o2hWIkiyvI5/76b+nPzGlUfOFV
nUyFvf7UF6I+BtJuwz8zefOvwV9/6+yH0nC93OKStGniIltOrADYk7WyZcx8Zz/Lk4EkSRk7XK9V
GIkBaveihHgZv6XCMGZ1omYCmPyc3M7bmiqUoksRV0zJaoykalGEWoKufBAc2Z3NGUJRcZBVRlYi
9nYO4Oca3ZhHVr6Ca0qUgOojpyucyRekX10oxZ7j23XRtfQW/+WKPN27Y9lC+BuAp62mloWciplC
LoI92ffYUmTfTrFd2fgZkw7dfIJ6iRvYbIxXbzy/y180y0OChTbDGyFqDXyCn5BQtFj3FXYxjxNf
qgMUt21jgTRA8b2WoELuAU4JxeU9nFBvgpKdguQJR4wqFKrjWUGqrq5rEcrepOcgy16X15wTqV20
JTGlaG7j1KWfxGzm0oth6GP8ek/Q5+bWPQCIxf5FjQiFUDcVVQc3Wx3CeS/TFv/iGnTv8nKbuh++
FVXKZEVPEYIYdKu+iOIQqBEz6VqIuzbFywq8+TCgVp9zHIQDxV3siF4ZfnYtcu5zY4eyr+sWw4Zj
zYeUInkE3+tCRzJRfX4fh1TmgGfULRMzcWjhV8glFjFSHiDL6TchFe2Hghsh3m8S7vV3dnHgZPu/
7TdypfsrIjD8e01TEteIJf9MnGRULLMi/YEdGNKfoj2mGbGAhj2t6lZpxLimk69hXhmPKnYSRgyc
ITm+7BYkfTH+q6WZxz6pLxs/4VAsWllVSyZzQDuZ54+LH6SgKHEChw13vbUbWniTQ7MDP9m3vWZB
/h/wJ8o4fmaOs6LJK779jBYn5fiht362tMGha/OniVEGhJNIAz6cZ8Ro2gH+tLLXSZlI+sRtU0hV
UR761Ia7D+1b7dkoQAmJ90DBdvxTWUMhCZOfGdzAkrDNoylpD5vfg24K4+Yh+J/YgJG+QBBdec+B
IpyD86MyJb9F626nyrAwI2wCD128Q/KFZ9Cds9WKCuDORVnDtVDWm7Jo6bzNF4T49qEjCXvRphZe
U6kCRAFFSUO4ZT5e+H0JOUlilV8On3wOW2NQXBO2jyicPzNQotAgLXroc8DqFUgpT3RYPzbrBg5S
ArtKj+K6r+k0bqQVtCWLzur/J1szZ3lTPZRGWK1T6cHr6v2hVZznYqsCFrWvQPMwmC7mMwA/LUq3
QHauNPgAuNz3q3pBgprqCM0fb56chRSyeXNs/J7xFIrkuSEtexLi4RJr5vEzulHM1vgl98r3ZdYM
D09bg4Gkca4+VxAmMPe6PaTxO4Q/2DKBRyIzRZHA4glTuAe3y00XxP/IHH8Sch/2lndTm+zHATEl
FjJzp+0oDPlaVx2dfmZfuVKwCTGpcRrewhHy9c5qCRPRkkrThc6z/LbAwLiIrDpBa+Iw5yBckAH4
mTRbYUZHCylPh9f3u0/tHWaYhnXllPNa+sXMs6CQh1EmKdwlfAd/sIIN/Z/q4/wTegmWh7PTqbFZ
TQ2BkFutHuSOgivac09uJXfqNvorwEv7lojjVNUz3ENsSe5KJ18yS6kSWl3Hi/yOugXkLEZnv+D1
BMdqtNCES5T7g7VdU+hPyR7A5jUhorKgvydqXBMX8j3QfHDZmZdLcWKMi7rWp0a/MfpKWHDWazGA
xZ2i0GIRQzu6hev99hpcFHJ4tiqnUvJVt3vKSqWgrYeXsxM3IgBmSTujuyWI0ihIUjer5puwaEL3
fRPRDJjGy9Z99DKeq+JfHu7hVxkg5tXDnVTDP448a8xCblPRQEkGL29PLtv03sxeXcP1BJM7iP2x
eXzLbAwNe4hX0urnJQ/z8jOBuT5jDPM2w6pddA4lg5YWAcKSEFIvNACAp2LNWeI+WCEmw+3c1q9y
nA7MaEfBS0iZ1LsYeNa+IujfKmdiIJH/tvWvIARcIiVMdvO9mgSJP6noJxcPJ1GGkZMpT61eDPNu
n7f6/TSQjn3OhZlDMaQsp9P5lCsQg5QEQ1VmSqUaTOkhEAFh/DZ1cQldMKvnVFTE880GB/h974ui
isL3N7nu5g53jI6PNoMjOuQFxpDxUZuUUkYBNFQxn2SC/99FizobU22Fv8CSZADB+uUfFQd5urDZ
BikJL7qc93galYz3Yeoh0el1YKAz2d0aey1gt4l5G1bI6hnO3mU6mR3UVeQ2RWV7Ci6pI3E+gDHR
CnurUblpJk2323P4oevzn+sPE6OZ1PtP4X0+VHIyMFjFdR/ea5gCzm1IzXptK9yWS0ai5K9urRfv
JwyfWt3WIo7Umf8sxfy/sQai5BaIm0QxvYj449EHkOP7GLhtvZaFMNbpgrePiQiAfBqUNbTz3XnG
GeymalbMo8qU6swCberYB49ikzbQQ4QLOJ/xQWsEdKVDKEXwPMoyseEiU8vnE6lUsSHr0C5sP7HE
yLwM9KjhcYhzLbTwF01K/Oby2cFWcXfYb/bWWDoyX9KYKTMd1DqGCD3iwNgkGreeVEvSzabjXC+A
atDR/miA64xBoYrgc6HsveJJTldw0celrG53mL3xhmkwX/Rf0Ud/4Uy70WZWjytZSzwqIG8bGg1q
BqmkUHBx3UlEmdlM3Zw4xeK17vF8DJh4CE6bWmfw/d4p7PFH5Cx5vldem49G6mip8F0wPhQs9TOO
X77siFo5OAcfngbLZIZz60/DunveIxu2v2JNANvM14wD5mgygbaznX1zXYHtzs/qOanGvLr4zYfS
FJmAqUV8GEFDspULdmNpI5ttz70tvhQmcLrpXw0rintOEE42wEuZ/+WbHSNL1p+R7zs1U8amJRzF
XKOG70erBKM1lcOrnPlY7jrmq4NzN0RRo1L5czjYHLV88EErCNM3jjysdC0K+UtuzsrxDMh53IsV
J7bwRDyJEoXRLcdwpPFZOojdILeYqNB+Vx923r6x4hEDYoND84W+25WZOZ7cTiqqxjXFa5QtkyJD
i5qdh4nzrt9jRZ/YYbXGX46Ar5FN8LpA1aDd+wdjY8Oky0MHquxlytNoCI/oHlSDzoTPvkuLp1ag
+9EkGGCIi4DjiMS72ddxCtIV/zi5hpluVRELX2XCeTR75MqIsdZKJWCSqCcRx9WvGi+TSxsWcJyW
WNZlYM1ER7Ndbo7OfSQtbMTtCtocuwOcGt2aXrluu/BNIqt/BnOEcsxmuLehsOW1CEArihlJpnqe
vtByaBFRldF7RaKAGarkDU3NQYUlQEWttLlk8Ogi8cUSo1ElDqZJZ4pYTsJnV1Rxnf2AZ0Ejm8rc
VCZu+21NUMbItNGhqqZ+xI6XAMr4urV5ZsC/2H6GKAH2KOxVQM38CTmMEuSEjCwWmFD91J2SuNV3
MrlwkSyMJnd1RieRbNUBd/sYk2DxZex0XnGnCoYqIEDfuDpSDQEy5gYHBrmZoo7/VSEDffpxb+kG
eK9WJLVQZay+sWQ7Ds186UVsYjoz8dOH9xx9LgCzcjVMmYx1piMY11plnx69asc/cMp5XiF7x5sp
NyrDlHikimQOSFQaMuadoFrh9efZ2B7xbsvvoQMB+vNhjdu4GJ20HJcxp94xWsgQ5vDSkDZ9jS1E
y2a/0KqI1gkdZyQghg8fQtOuRi9IZFrZPG1Zo3MXGCPDiQTlwFELzbJ5MNTIwjkM0XSEEvlFWEDE
8WrHO7xF3MwhChrRSYrUdH18aYlSAUB7yAkHydiv+aVF47/r18Kjwu9hHH9D9eVeCJXOonuFwhj1
yxcuZruijxLkfUsWVk4PYJjPSpEKWZewls8elCbooUoynbvOD//v7dVX5LK1EaJXoi8bETdA+ZN9
FulQyvInx8Ru3G5LZGIdWil5mNJeEAo/bNANndXjykVmEUVIVemI0xfDJmINLvB5i6VfNEcAIvA5
peiKkvJA/IEQa+kQe05Q71ToLRL2ucvKS5TrGObUed33beH7qEq7jXn2d9Mxspimt2paa5XnIr5t
kZJMK9jWX4ihCRjq9/dpuVCTU5lP0gRAT48yePHQa3TRKuqvE3K3qQnGBJBovzRoS3zNrsb5ZZuV
KrbEuxYr6vKsSrDkWQqZiyJRpwSd6VihDVc1/p7wXo+4/zhI8NbIfF7PHmjG+tG6aTtrzhVffCV1
3RRtuTApk2nqhfFCwTKjT0GCYHfLk6iZeyFB6eU6iF4xz14Jr1qkNP1DOcM+SMvCfLZYeze3/lqB
60WCStM+oRhbbXEH8cle3yUXqMjAXR2Kz9HuCRIr1A9Smuq5JuTA8jwSnoQtSPz1LTklRgCz2vMJ
y2cJReQraoMlYOTWu1t2wx5SqLYmLdXNOE7NDbz3CdUds/dHe0zUWbz4C9aePdJJ65iu+RG2RU+Z
DLOxzohzXwNN7OXn9EcWfsDVJ2ZuvI+nOMLrbJttm/enxAAB0jZSJ8cTjHNEKWguyseCwoRwRTx9
F2V4vAuJfTrU2Y/e2Wz9qh5eyf0muQxOntAFwUo+szT6+SsZ6730HvHHh4BBLTcF6wEMQV5hFGAY
g8EsCQnv5FCiVqvJz4H2HlmxxdxX5CktrABpkhcWNXPVtgoSwGXubfpDSGOO8Nzgfc0DV6ss3/AM
vm/5dJdqoDjFRLWbO2N629tmz2n3Qjsx76mHcCQHi5cWWkIW56aZYb3Y0fQ2PechXF050heQt1Sa
eiGjwScgvkNO93PjmcWKFWFoKr2ch4fDvT5JMe2ozTL1qjFjumyDWDYUBA4/RAFqehDsXNi4M+xv
6pY7Ck7XvaHVvq63/IINYHxvazVWolMAZlwGsMFAm1pnZRkyigpV7BAZY2EtJFiNqaTEA/LwZmDy
r/pwv2aFVKhFpfMHM8UzzWBAlpCGCdaZGbRAPRc+wO652sFSkmz8u3BmkQqc5vKXNXNr7wqsu3Uk
V98MK7UHeJW50BPGY/lUQcdBbFsIVDadmVzWdHBuvYmyKWMFgzFwIubV8x1vucnqGt1YMaOrP+LO
M/XVrK61GuHwslBSbWBHmZfHDVbsH0rKhlUT6m2yI18IgLUDOqcc2HUNouMrJRpasW57qu4/Z09C
YXxymnbp3D4NvCJtB3GT0RV0+3L9T9xyP+RusUBDy0V69A6QKJ6yRVwQ/2AA2EJh4NdkAu0MtpLW
VbY01iZ2i6JF7eovfyZFQkJxbgDiD2yBRhm4YEcqs9XYPrv5N7AFW+oSqwTfb5Eel6m/IgRTr76s
yCJ94lS9r1fhl1faYj2zN7KubhB6g90qixRUPOzV1oOZ0HIUF5Jm6Euy2l5UNGisYptPw5y1tASl
cRpSggb6vxWZtWYJQ+vBm1udGMJd5ualsnbS0a/Vx5swjnLV9S2WNiCnDhWNkXIGf26Qv+L1jAfV
VXFuOMkcWC5dMxhcptGuxFfaVIR+lw6nHR4NMXyx1ldq8ywGw/kL9z/q9U3OiMxkr0Tzb29G4Vyg
5H8rDxe+aETPjaSIs5PqBR67zyoaUuuZulMN1mwNH2UkRtyA8xkDJ+dY6+fVznObFg4lWxAVi6qK
OdsYsacFqvHPBluTaZA6vZwp8SKmzTNnjQ103ktkp8xdV6kxAMf8x2Ay1Uix9DMAt4LYWpfQIGMe
Dj8S59qKZ4tiartnzM9l15UmxDdtmo4f6OeDzOiG16DpMm8tIF693zlnLXd2S0wVwn6wgmyhMqXa
5ddNeOrxNRCABAnO7I4/9X0tUZkcNXIS49As7StFrJI/DuCF1pmCrY/NK74qYe3e46MzobLJvrS+
z+G3a36ducnIQzAbNLL/cc15Sx/Gt8vSIEk99+vj4I/Q6HyFvwhfO+cRlDd0fA2L4ewUBwA6PpXf
wzbk4fMzDjHsg969KHjAPTmvJ2sPXjQJUqq8C5j4MYzTrxU6gfTt6KmvVVpZokgbARU2boRXsGOY
0IFMN0QWKRqAmDxl9/86ofgSGV3oJph/NYqwxz0u5puvQMdYKG07twkvhkD7gmW+wuaUpOI91MU9
SKZTQ0bWtqUIuqw2giw4jdDDcpS6YoKuF7Uqs3kD2uMw0nykQ+xv5X+gDQq6IheggFd1GgxLjVqN
mkrf6+2FW91Nm7z+Z9F9XAh06hbnYMNjhZZ8NXP+brr2SYErHIPB8h3pUG2qRI++WzciGZ8+9uGG
tZ5mXfIBNTHuXydVGX6q0BtqVVMHIUnhFEW0YanmDoAInAX13Q13LLK5mHqvGblPOTXoWmsmmz+H
ev4YfX0w420vQN7dLqlMTSV6cSdRNYLBfBAsjHzH26mGjszVdqa7do9fNz5tLXj1Nqvy00HmVx6h
Hq55G/kShqZF595vKWJbn05MGmFTAMqz/6N27tj26L7y3I/B2+cSeI1SX9zaECr0y4kt0mvRwRUn
T54VKOJ+IS/aKrpQ/KfxVxVG+HJIe5tUy07UCirkiHTKnLVuWHwiEdYtqALP1j/LKwanM9UcU1xu
CFG4Jjc+fmKkEzn14pi7l0f0z9X8AoXuDLvVTs7jVR8MdFb8RMkcQuuyVumsv2JmLKggqnKH/0nH
+09iDGbT627ghdONqLaHuiGur/om49JFR6G226zp21SEUl8X6BiTrBwfr9UZjOYbqOVLe132pvYr
6EU7lTTVqSIoUrkDRgbupBYgctBlpx70GjrsPaN3qtPWovvmGGCcxlZjoF0rkkwoE0TgeLyYAaHT
YtQ7IUrn5UtBEPUoVIuerLpCTYWi1cw2IPYjJkWCgcxEfmEi+gkQbrwGr6Y6cUTl9iaVzTAhavcn
OUv+8IwTJ5V+hsP/i5W9IB6O89Vxs7a6+lWQalrfgPDoqrRCIWAeogRrUnfj08T7uz3wM/0gn/tS
of252sIJtBbHjSpoYrCgd4E9jBs5QZvsfGyJaE2CnJJBn3Ls0/VZ5CankWcpwhA1OZ9QoeTkL1Wc
1AaUNWQO+CMm1xIB31z348pL8jqjvLDGhIBGl4d5FmlKO3Ot8URkretj2xQdzH3EoIIWmC5rYeR6
koNcHxXKqVpZC9OpasjdDO/thLQUFpek5+c8PjKy+Hmtq2pZX1B4Usyb2I3HCMsYi5uv0wuOTWrQ
OCTcWkbKibfVLxy4MuXmVnZlXMDsmSEMm6R9KStY6DYyi034n+ZZOuN5+5167iVtpgwDLwfIsrnb
zRkwmzGjazHENStomtu/LsK4wih0PT6vW5TrmanmeIVC+XkqVszsmyVICSbMvkrwdv+Sk8e1ShBX
HF5B//wUz9TNSmy0sA9khCncohevrR33zKt2G3KTd8R9wZfkWnqOyd+KRObav6Ac9xvxeV3eZSFl
k4ll2qp8scbsjQe9hDhtjUTosNUcMTfmYipO0isnqoSbBS28oTz3nlYmORsdBq6fIBb73TlmlPJg
1IbYWrRYa6LY4ea+nQOP956QaZIzdvxhXFM+XvMpdvm2URlq3iCLE79bBxc3kTlcQXUW5iHS58TV
kdSMdQGEw2a0sxBx6M8RaLSpIm0o8SNeMDdiVHrgMUXb1qs6RxNDz32SZ0TU7mp+bMUWHI0xfL2/
9I+3tOKRA3h9iIAza3Dia4V6r/kaN2B8udPsLQ1W9hkC0YQWwRxbVOx/RNvMvMg16fd+5oaurYy6
cKkIm9GYI8wMIGWwUYRSl2ZJjgw/3OvRkHSDx5UsmpPknQ5vMFcKXzThmfD7Ge9vQfsTopQO0xM/
qZTNTgv/uIZZFipwMbi+J775By5CBmnBFNj+h0who5ByXUq+GHYbUxVJIpn3TuMyJtNHpr8DhlUg
EKvS6RgkNyiUHF/AqfRMUFnTocq9aPNRVLXeAYR9h1eAt2Gy8hzjt2aM43Ns9rO2zLbuw6zfJLzp
7zEZAFoepJ6PwJi8GaocFI7yA8o1VmC/pK15kFlfzn5xY0GHNGTuBRFLKMwq0t8uMUuLi54Ftcrs
KSLuyPxx8Q9kY2fZgZ8SX96AyvJwIGZ30E7ZBgHBG/ZOGEgovmXF6NkLay00rz9l4vVx6ujysjJZ
++ndZ7QU33l3f/s3MeRIEQq0lZ34bE/xJOOjlbxXPYBkt/MIsLYkx6QOO1KoOeGQzpDEyIejE3SQ
wgNk4IFvxnkTOiUmheqIUx42tCH6U9L/a6NtkbrhzDkj/NemWnA2oC25PewrPBU/fw/QprMImig4
01zrIPVKpAh3pbR8cKRomI0Yw9HE3yOEyR57G4W7mtqvE8fg1eAZ+bzZNubxka0C7ZZ125Z0SLsN
5tCTGp2XNk8mV0XhvyjItExM9dvdBVGlZ0xBirSE68KhCXqHMSDWUboDmJlrrHAet6uaE3oE74Ij
8w0kjB1T/IsQaM9heeUj7nXnH75Ts5/K3WOsinVqqjxOsSd79smEspa2WRQEwgxU3LlD2kOQc0Hg
tv5X3PvfYB9r+np3/stRYwVSYK61GBo3LoOlD8J6OzzjF7TG5y6sn6RlPvfiWUl7bPv2MokY9fMR
HDG2VGfDl1fdwAcOqHtc5lIkL07VvOy4QDHvNdbntQh2iGRpZzCt++wyRNW4vbYgiU0iu+ZGrjdK
ktI4FRau72BqCtAgpuItJ6sahxf8GY41CghcIR9MajBuSjWMfIY4Onf15K2/ToBGrBdVxafML08+
GFpy6JX2wxJaTvKgwIrLkR0OBKzHZ3jnihxihpq7H1mcxEzxe8XQDmuxSScYZvZa0OKrxB/ZCFnN
vO8MXCIrw6v/GzLIH/4INj62EQ+5EM8bhfMaw29mha0VJYHh9uk8PNi55mclMC2bjvwGIwlxGuik
czxr8Adfpc8BKJRXn4iw4Qw5ymKhsRrSR8kQa8dDY86V/plw4QaRSwCenUvE+TiI7+wzOmIqH7nD
SQcVBxL68bhv/vz/PXHuMad61CQbHw4hKiWHoTJlr9p1VkRUTbN3mNjNtlpHX43EqEtCCFMycsEB
hf9KKTJyfk8SV6LVbqfUjWmuRdek+arvgNEp14KFN7GBCkpJMSY6gMYzMI5uJSHuiznjI/zQKUEg
oB2wW+4Jzt0d0e5mkWJc3A0OEuai9R30gWkzM3mQvkmAEuCdYNkWQ9R7ccjaRIDxumDQFNvDQ0lz
rjL2sWRX3qs4uD3Jyxpj0LdaWA4SC5l3/aESBh30Ww3nu5nzEqDPG37FQl3K4/o5o2ssNx7NA5Iy
ckb3Ct65umvC8Ktc9ADjLhdxLLQKLmBfsUYd4DTjx/vbGgbz4NUzfYBP0OAkQzQQsSaKvmhmQImy
ABupYiAShFi1+S5FpgpVpadicbXZRdOoHCqV4kZwfjzqWMJ40K6iy1vrAr9fN5gephT5fFsftIbs
dTk30eM7jzrMnb0CqwET7uCUo4PGLAEOHHirFMqkDFAf6tRrSVDmWKnNPrUHeW2srYc7Yu3SZAiP
hzjvt0ya9yXeAUPTBrduiwfIF1BQIkGuYR5RQWIdJQk0IMAVUeM1HCFqDK+MMetLuQnakYuKp0eX
sdq0LAk0dWXCrZ7KxMN3+mX4KqP9nocuaS33/L2o0Jb1NLrUMwIKy6w4cNQi+claIqahoGcibsrU
90Fax2tQJ0/nkReWwQSrwiwvONadef8qVPUCUBO7UREjY+ahEF5K5PCSjRay9nHDqulLdXETr8Vv
6upC6VxyGkmPehIP5f2YpGTd6b4zOGjjF+4RSARNKqUFBd1AGQRw182htCyvZdTUvjjf8slVh23z
R4ZmoFxMalhhMaCj/og4O0/g1Syu7XiOLBinPOYxjZ6YI8JKyWEkoh4kgdGi5TVXDG2QWqX4b/tA
9DyJv4QE8Pb60h7tl7x4of+0hqGYTxRtLoYFm9EuUidEh0AJUrw4vQMQhsTBJjMea/PxARN8z/Sc
cKxJLyi/+AG0WPq4GhYJv2JSKzkREKbn/9dNMpMgQS52tQaM7ZoNoZ2hG8umQ9SrTSLa+6iPXF9L
ikn0gE+k8pzcGoFZ/AGzkofogeHd9TXG3jVkbQI3UOvwWV3pdJ9+x2gd2seJ510JUtjck3ku5ZEa
62GMRbNgsD01rlip80mQpsQGo5DvZasN1TNjVhtM3p4NQjZlhOIfZrFzR7eeKc/yE99RtplcQs1C
6aTPdmADcusfnzJLjgWjSp8oZJ8H2nZp5MKPpIZ67MTt9H528u8cSEhOw9LfXWvc/Hf4XqgZFBgk
UZTTozdrGK6TpiOUUk2DsLigde6fiM7piiiGIz4454+X4HMgPpXjUE42En5a19Eje1wBRZ3eDTxi
dRW+N1KaNEW3uT5OBd4w8Y0sWBmM4l9TniX+yVvecvc7yU8SOS2fyfd0bWd3mTzkklb1jDYTEaiU
IK/OgUmQ3tnMgj1cW5D533o9HrhsZprkp0PmgwRBW8lsZjW/efB5OadhhltVIm5yVw6WHOHe4gIj
Mk43gO58a9HOQZaiSM6r6hWMJRGkzBto0MLVX48qmEUWa3JdVgpY634kHOC9rmsSp82OBfJ04HJz
cSzL7lPhsfbgdX/vvlF8fDYSE7LUhxw134i8w/1Iho4oDrd+Lq3/QmjgWhIV49sfquh1UwnBvhNy
3A/ygcStYisWLe7+9qTEvoiu+fqeYJEZrxo52unxYSJTmTNPXc7eOCJjGUPdOzqO7StakT/ULloP
cuORFt4BJTX36vDLSCSZDgNAIqtzv2K0bW1FAmPyudhsOc9zAg1cWTbQz9oCjCmLDmfC71cQDwMz
vJxNmZWIUKohkZ/sIlHYQJUAOR6qIed6FPdFsRiU/4eZ7g+pVBJ98p200FZHfUa6vSOISymokaO0
4qz6czKVphIPqb6tAFdbg2eAQoVpYi9j8V0S05yWh+wNUcL9BN1VXcne4RsElM57AveFs6wK4yKI
s/3/GW8aDS3c0RjO+s2KLvt6xZVBlk+BUNYTLfy8ldDJQRi1FZTUqf1bb6dEtKsITQ9hRhuom9w5
O7eCRRcKRCv3UfWkxr07dn7KyShm3ZAr2+WU92/49/8fWa5akGG/Gx7YCrduqGeLKX8rVMT5SWbw
bP8ecj2oMxtjoMqONQJ5UEo+HdgQ/GY0BUTyHBRwbIJvlxmAb7dlrAqr5jKPduFXm8E3cHnC2XAL
uIaCVRyL6P2viC2vGlFqxhGpy9vyOk7fypCLyxmTKqxoXvFa5HAJOiPi+vic0+BrVECR8NttU9ok
YpYnLwXts8bRUPY+LTlotWUFmh4qP9E1yi5y2TbTAsu4kRsJUzVts2zDkF0d7TrQLyvLww2IUGp4
PbeReHu0VNf6GQt04kAcJ95cteSFsuAxXmCgMKZVZAbKfTkv7qKu45it5sLZl0yz9vjtmD9GgZQt
zxl4CUPvj0/N+LehDhtxAnpkGnKnHyMqWmLLe19Nnkhlmu+HEcuOZw9+lWzbHZja88dsgZfVpzCX
bDqWJafu6aWKDFQvCiYBWC2i7e3+UWwFxykJD5Ll93TiAPz1HnEp8wLMxf1oqqWkdXjJwmRbiRpd
GYwG7uMy0nQpUoAhRv80ehflyQUMfDSG2KgwFUKgrJMc+nwTmODcg/M7e9hket07Bck95f70Ps6P
luu0dP83NJylqC/yeWpJeadxr8P2treKxuqvcicFJFIAM49sDKro4wTZF2Rf2EHLgVMj6eKmWDIv
xznxOqzJ78XwJVLoRp6/otI1v/BXz4vy7GfEvQZe7ACKeVZnpHH1BVWsgd0RnplTRViTYP6+zg50
9HbNVtIQRUMqp5fyM8KM9IVBg/gXlvyPE0BMHVHpjjkYUCav3qxzlGe/nc93HpHW3BdzOkoJ2/Eh
78Orq7g1nKrLGqoL/1ocmT9HEM8+FmK7TSsxCfvxJ+T1crVOfXsquOkkNpX/yG99f3zPtUQqyVGL
uYnmhsgl5nrSgc+HwJaVI+7+Ex4hCGXjRhgGPHp7NfT2PVnmt8ruaeCpJ0JMAg0vSYwlGfDiqBkh
q78u9j9exQCpn3qJQRLa/aeKjCbr87bodaTKAvtz86+HKkGL+VnY7G/XZ3kqIxFi0bpyIfKPsmup
wSPYo5flyQiPonIe6v6+FdRswWx4LInGvAjjrv4g34dgSkp1LKN4JG4hiTvsavyhycL1B3OZakN4
QjxET45uJIA1VQkgXn4qJvdDw0EoIFyCq7IKmfCbtHDval/7UaZtBG3ZWXyvvilST9voDaGdgcKn
8VFtihXuFTaomvhRyEWg8li45eaWZZfxJ0yEe53n+DW24N7FDSIpKxNjiKLIPBCiSNM0lFQuXag6
jGm1UPBWvPX/kB4KEcNa9KJHRijVgLMH171LxlBnJhaAeXq702P/2Mf/lXTUcKBE3cmxSQ3aPF1E
W56pi1bKSy5IrO8e5NNPAmgUVgxB68W2H20ZpzTOoTjtiIkWggZhlbyHusZ9teUtsC8X2zUYzqPu
iBttMqkeFY0/722jeDHmC2Obg87vPpz3iQYISLPSp1RhIwzcOyoHM0cFj/WPE39Gr3WRIJnqCPrw
Ygk/4VzrAkdnNWNUk0PxYSpijcJqLeOW721LKW1DsXpIS46/ENYr6HhmtxwmRjDpsdIEaKsi50IL
cnqjW7apZ+F2/ChQLf3Hdoi6PpvG64MDJjbPpckhWFC3asyrVJxmcs0/zq/5FKsnt76xHe05jLil
mD2s6+JRMhXpLCtPW8KzsceE4oEXTO6uS9eA4rnfn6ee0RFP0HO1bqU4xuLj+GtyyvmDVoqSNnoB
QE245ZAieHzIbqQvNELGxff71EjI9lLvTnGizD6uAXbJZj/jWuPsIK2nWwkDEF4uzqtd0NCfILQ/
kPapR0QBM6wOTLYmsnOpRG88nVY5YjT1d4jegWjRKhqTyhsbP3h1TkngEr1V7A6Lt5cUq5StAfls
yf1Az0CU1/q8MUZJmDf8um22Yz1GwCLvr3/lnocPrrVooUU216a45qxNrZ++TtZf4/LerB38d/zK
m+HOTqF3ly6u58fkNFt658jwVmiG2KQMWd4oXYOZqUuwIg5jbcDGtiCYKhvk2fwSnH8nmHvOZG81
EFbyLIQVQawdMgHCuXU+CsGPnLShL5HfT3Uy0ujeTw/QA0B143STmf1MSAljhqX+sAX+IJu7SViN
kpvfJw8EcTwcLGdrWA42VL/FP9nRrZLkg9JcIjltayQzhaNapi0VYyUPZvWQem63lDP9Yqo5KdtZ
XbA2Kye1tGm5w1R1MoTlHdjB6s2zmBW8/QXd0navy6NK8kqB7YlftieUTCBMGEM3FQ51+ElTlSVx
IBQnceP0Gc+HE+SaDijn+THhbgFUkk+tKQP9dI8xoYvwMvxInxyC+7SAEpqDVOvRPKWpDhfHaf+Y
Y0SPjfZFH+OqUV8sGwdzykbm5LCMjAQpeDKJmgn1e/hJcq3Taeswrj2bODcBGcdH3Nwjc5OC0sr5
8foaw6qxmE2fwUDStQT6XXDo795c4VkFJ7osAAKof+iKFHzvkKutSXFoiKReZ58lw4a6UwUmnBh2
bymvuAsSDZ+aVhlqqHErg5D9IeoFkyUHC58F28LZ3VvrLr5TpTO2ql7nRM0JCT+GYJlA4/mlSNlO
1gnQA/EzQYLGb+KVtdx+2AfW179YhvZVORhQNn8KfpaK1BtUD9pbTDXepG021aGPmwsno6bqgXgi
twGG1tJsRfRPfIl0Ll3k03GEeMXOy/u/9v394kZwPLNdZsQ5ToFSYR0HXFMEzy/JpHK1yRhVUwMG
LU933krdrtJvaN0pK8Lzea+2YSJWSFN0/2621ejqk6mGgAzikUoLX6u3xOGt9UVRSUbJHO+pk2Ne
4diglKa5On2rGNI4SVIeln0ms6UtKPkd6nvC0QfYzmPHyiLgtkv2JDKumkh950aizbpfk3ll0xIa
DqaB8+dEsmaVGj860SrVJdNH92f13XhK39td5LNfCAvNlW/iBF7TYW5gFPiHhCuUjOLP/ZAix5tT
P/H0jeL0iQOdKVUJvGH6JvES3R3ZRteWZSpbjWoQyy/44tk4Ir+N8pBgqko12kBbjtdTjD0y0viO
UG/GNMmdAikS3vUbdWHkUEZENv8R3djSFQ/8lBIxmhmojwfTE+xeej6wU6yEpznHMxoTju1IipbI
cICKC6i8CbVeNrummnfSwT3QwKcTS7PwlD1dNb4iQwaQk1ZzY4uUpiV0Jb74aMkrptOYyKlCbs5v
FAdvpSoz4qQFm1Ok3z/2zzifQ0awQlqVjlQJppDlxwTBVvK6fopTSAdZaeNoj74Od5r4FYgSr6J7
7Kcm5tQJ7YeSkUxyQiKlUT5jYUEPccU+JFWvZDLCVLAhO1gDBY7OO0UoJEy308kXndWw9aiqcmQs
pIM8mRm5Km5C573VyFxNFfiPK0u33bIeeahHZZ6bhApT1MS1DjcZBI13xjemJHSM2aGEifMyn50P
C8yPWUASXtmuTihBsagfILiRASqmSe0W18S+b+E+WdyVA/JUAwmzhxIylLIjSNmMesCNrCF0sZE+
7IP2kU0P1LZ6FHIxdok9NvP96A04oMf2TKDeTNuw8aYUqw6gRkM8dKke0F1H600fVoFE5iK9HzaS
0HhysLZbRLXeDcA1uehq5vbO0bhXvO6eEWHjeNlQ8CzUsv4c1OtMskDV21ZEnwpWn7RY/wSTAS6D
Wdr3uIJaf9TYR/y1X3joy14u9cEE47SoIMjkoM9IKIdLczLu85Dd1JhG9Il3s/pZPkL/GwA5kwla
uI3euWMbMc5zxI3fE7z5uqe1xcKzui8eluooQPCIBgG2pWC3WfAcYls39tkd+v+qIliVXCIofFVh
292wYDxinysqk0UYwa7H9/PUDsSvHMtspDsfIvPOrnK9I9kdA2J5dlIGY9kSDwVMZ8hPxsBeWxDL
BUh/tU6Q6UBbHdvDeeS5YJV5948tB7StSSDFJGEQqsjrfKX/ufbII6iACbaB4b/EkEPXqujX0gL8
U4yO1LGg2rBC/b/cukZF45AXlzrkfrWP/HpYUrCA1Po743qBRXQ2bE++04h5OsA/7OoJm3wAxStN
I3fqN88vDGEjE5mSTZMQxig6mh+KbjHKuL/bIQvtV9iVBHdvGlAlaC0Wup3NjyZSr3k4sifabNQF
CUoZvU9cEcJj1gZdGqfNg1u6DiaA8b21/ezwcCFs82mRpj0PDangdkHpVIXnFFvVTa1XGwyoQe/l
Kc1ilLTbqT5OQk0XdfnAQsldoVPzJOg3UWefNJJUx7JqP8n/UjFeSxdhY+GIrTWqkgoQrV5UkpCQ
WELyUQpQtnH5NpSYA1ET3nKJzP0dfUJu+EBXD9OMAxmRgs845V/+kCABYSUkEeLlQFMFz+smeM22
QuA9ZhY46cP8jv0aI7zuC9MhuPzu6R0D0J+TRZF1oRVwf8DSIZctlycT46ftj7gBUZtIEq6uDNC8
GoaIFdHg1rRStIqED6KYqGytRbv2SDM0YNvjhyQTg29pPVYKHBMJCNvMAsRvz5kpIEe37LwoNHru
f0KH59Ls6LRp72M1BQQVIFaZFggA8x3LEXkx75Fe8n4wTcnK/exsScAM3InjYQO7sHCgCRDWzuo5
+leh8y145vIp+6KucngHQcBn5cv7G7vVX0s5tW/a1QoZEX+NuIuBw8LtG7laRCspu3A3rtEFHVxn
vvvDrObqvFEFrJ0YVDdFzPT1iheGgTyAH4dfbx/n+hdhRWHBphFeCYeeF48KJhzIyJbtaiHKfDGD
SdNPSAbNX9T2iD+u+qPtoLV9hpfoifsQcMIZkHGJ3gqtmAGdB2zJfnShCSN+zJYk7LgnzEf5WtGv
IRIHt5Z+auNk+WpU4guuTyELDFkWGBqh+yUQzK70BKqPGoBwIGSC31iesmW04tlS79xHfnhRbzM6
TUPYPhSD2F1UIPXD9odNfTYlV85CdHmtNyYS05PpZcMFi0S6Pk0R/IbJIjtLGVi/0J4x4EO/x1MU
Nl0XzNlzmE4UlATAfWfO6w7VN/RYBJ7kyVvlvKksR2xA5oxO0Kakjx0tjf3LIjE+HZ2FlfNFT/Qh
Tdz5GwjN0W/5ui0Aue/FmoF6zB/WGkkDkiAHm3cB60aBK9UzRKoioyUuPPbm3kBygq11kQdNA76S
sC3gCB4ifnlNw4FRvIWL/fWtxCcIJvx/dmEsfjqhsNEWo13YwrY6sP6S8ogjC0Peu2FtJPNxXgpv
R8VrSU9dPbKmCl5jo6PqyFYa6Z0AuaUkn+eZ2fjfm94/RmFVjzaZ+PG1GxeZni9IhZfVqDbyqDea
wFgSA5VP7Ze9raLArPG7IWwlNOlxTeD8gs9jn18J0GYzA2pD44P0Xj6eMRIJZE30lBDKPUpkFp6a
Oe/9fi5UJ5ACYuPpo891qbsoXLiKzthtDg9IMg+e3k7iUt8yJ5WwsiZBQROwPNM+/qLUf2cbEJ9s
4UMVux9HRLGfNcCVp1EwO4cbMSu87DF2a5+MsUe/1rX4i+XRPv0gwgS4mSxVsO5Pw8b4oa/kFGLb
WK3xFsLT+Tcm5E0bEwwBORV1laoiFGTxfS7bjcX8aRM7XGxGWVd+GpCIlaCruMhg2aljzCNSc3nb
IJOARXdCXMLukpWdr8cJx4wrxtz+323jUUEJA8JiFIVSrp+kdGoe4E4UCLVSYkVXHUSyLN2SNJmp
rh+X3MA+gNwnf1ZXb4QLuWbfJWq0o0JGG76h3mvQAF1cWPUPafEve1TQMsV52HSSb+IWkXwr3YV4
19PXU3COT8SD3KTVeVkxC3lZSiNZynOITBnCGbO/T3aEWNJdCI+ZkH44jfAlqWlRb1OA94CDl9O4
pnzIgZHjmxOzMr0525O6ZaxwhucPeC1LbAHshlct3pqF3EcxRNGnxLqwNpuKzhxqGm/fnwQx93EC
wVdYlKIZV6j2Bs7QhRmEQsyn33B9BRoKoDuA8FnHFZeR9nnUin1Vl05h22URncgRTVo4oL0Sq/Do
4jX65eiwhqEK0q00AGQzpfz5yeXYuSz80uvLwKlUBK61jRGz349mux4dXwX5IvrLl2pHfIfEgBjE
X0m0TzP0XvnfvMribnpeGCgjwT5IH6t05Md2CUYPj9Louo270nuW/kJ97hpKCd0Ek2SdC0IHBXhR
ooUJW50RHvtH5XBXcpH6FcMJE/M9HERk7kLefFjbZtYPngrNPs3L6eX9S6S567yS73jHin5Ol8wm
xemBP6jvEEUzerYkPqrKDmfK0NpTqb9NY7STk3RexFDjGwG+guRpL5TqD3Ge0rhqYCmToOfG0xX5
UI6My+3Y4K6gQHWm5wk8JimPlvOKHfBLXvoY8u6Du/h6M/8EnaXH3S7HziOeW8qn9sPpnGWMkoeF
9DK8JiJw5tsk0LtcsMOChxm6f9IwB/weDjiXtX9M4oSg+xvu6bLYmzv9VG1KjSXAb0kroqeZeTCY
C/ljMNdoGasNPxvJreBE/N23vJnPMf4RoFvjTlHYLYtfu2HneLkPZ9CT/LJAyZpF3QGqVSHQLV4y
qO8qeAxVkzUNxDKde1qhnonCS8NimWZflVHfGp6p+zZXuYQBlW/kUMeqoxKdvryZTMQwXFEfH7aV
p/uCdIgBso8L7taN9Biv18Ani6KpTRYOSLbL5ucHXkUPNln8f/ScPzSiFEGqwae/PVyR1MqQSAh3
qOWbak1hV5jIjzalnXE8RXJf4W22F8Oo3nL1yEVASEDtfkdNsFPxeB6KQhCoHwNYGGi+ILqRQuhR
1YXyvavBCxJDp6qsXFfH/fP5QsSvVgF+YgOu/lx+taOBdSTdySDUQHDm2GV683UNsk5CJxLAflIu
wNUB9ZwrDw6TglJ1Lg8gJNKtr+ajL6BdI4rV9Jas4q/MjcLZVNgeiAQvQN9vOEaL/iXxmBT0ik62
RiefNeCO1POTLNUkUns/Lwo06FxGLa2fJ8IXC8bBiCTZbybifzCUuMQoiayt+nTfY3ewbFCqnk+H
ra2jWNB/vQt1elyiRhsiqQKyOfTFFF03ztiaFuMkDyPCxyLfWXJKi+/cG0MqWtA2UCRShAnR7ABc
B4A6WZTXI2ppRaGU6tqnS/sAdYu60oO/n5C+oT5zBqEcJkXAKe9Hv3Buz5OsGlZBksZFDs1+V8Wt
mSD9N1chgSE5RNNK9MnH8MrEkVWbGnublZUPYCgblViDrSxl4unKIY/wNBuQsOwKjxfGXErbTv8x
/trrU4sMGXn4fLT3A15/sWVC79shHfCQ5xtTUv+irHBI3yoKHCOs5YQomRaFuF+Nuac2sHJ1Wd4Z
2hC6L5SYOdj4BHcV9KzZAWei5FWquP8It+QX9TS5t1Fr5T8XVnvGYibPqn52cJul5DlND44KbMI6
Ly04LPT2VC5OSwKT+wV9eig/mVcfr5ZoB+KS21FRphuGWLWf2l9/Z2HkV96CvxtKU2Ayp+xNqkcw
kvQa9HU3tfH+NKz4w2ltkte7WEl+q5NsZWT0Yi8ZS3o3GRlsSBsVdaOfn0HFzs0R7fUNi34b9iWz
I25r90SL4TyOik3cUpBn55aGmvIYX7kpvr6NHl6ce7MpCsxOeLhzwI9atwgJfIp+PhJ0mwbNmFxh
Hz/HrQhVQiZVOuql3QKDUxt7fn+FEB799/b0y6Db0GZCJpNCtd/0DY1ms6usKO2Kwi4Kwa3zgkXH
RID7oFA4gSjGV7ChSrzhWuuTZsG9ke0h+ou09EcS1xyjKQFlzdK8pjZGwsyo+PaFKeMb6sofnsuE
3ZF8aFzw83k3hWQ3pc8cnzRBvGF2Xq55L4LAWj/pk+LwGW9pDzCtpX/XnYhxYUd1QP+NE4de0hNJ
RfZPhGrlBX1iXTg3QZNasWorv8O5Cph5ZB0zrmESzjxle3UvH3IhDW5GD5O+zeOops6FV6PyVZi3
5FfUjV+7O5VQkeNeE6Q2vTa/x/VsZQ2OWgBFpNe05neBXf5v5YhyRk680DuNLRkUQcLmrl2DFgv5
J/A4vhDnSXv2KpjDcM2rEaEUgsI93BX1EkxyhGsxWZKZiTFFaDuodsjU00Mof2Iiyl/ofdc65b/W
kZQfec994uvF+wKndl+5gx9Y96VKIIEo7te5b7b20xxoBWYtZ2r8pixjzhZ2lmKteItrvQ2jgzk3
riFQom5f1XTrCKaDD5ETBvCJgdHT/mruFjohxGtusvuUS/dKfjm9jmoRuUsy4shqols/9CM8DIGJ
cGzZRsXrYm/B9lKjdocPDIgPsV1FRfxlr3BupS8pxFhaBPaKyq89Z3VB9vSKDL9AzY0p2C4sbvuG
kF9zbpz4dVYn4L4YstWRfcf2PXOxFHe0vX1H6T+MudAPWo4rmHDfVFj7XP+JQv3k/CSf0fMDxvEj
71e21DMvPDwhPSM8Ix0dG4ZG6ME646PR48xbd/qelrK+ul4dV/dLc5j4VAm+yAi51Nyfd4I7wIJz
1dT9kiSrCEkdDkUU8F8F2sW0MM5/ZnnLNJk7Uevp3dXmBCAR6BSvGKLg/QMWG04UoKHbvpmiYjhB
fG74P5P2pLrLI1bu5YVainszwCHv+rmTq2yDnoMr4T8zt4QkPivgyf0UfTuQGZcWR0sxLkx455zh
s5s2ZptEDlw7OR9l9yJECsDcuCKT8Ool7gbbSzf3KKiYPqgzldpgJx/or1XWr9AtK63Cw8kHZZJa
u+p8cfp1ShaXjOkrP9cQV1dvAarq99DbRpO6Vw5DnUsbWO06HtxSFhNDq2xWwhI2OnTY+dR/SZJW
/eX5UzapuJN6CeBGvvzlHzFmRZN/fstyuPPjaut0fEubxiRp/T23dlt1Esqih5iidzZ/EM2RMTJj
NnbtaMf6OpKWaodQRxxQ5AEraHS8X0Y81WxxCQ9tdt+ua08C3yikEPX9H40w46Pb4ifNKnHSm63z
XO73eISQtVB2jCmlhxH6fbv9Q/s2nQc/xlkiNo06GbpkF8kn5nx8zE2vV6SfJXPFXIKiHJYrQhkJ
QTqRrtUylVBhNa1vUvqGLRgmcQ7xc4qR/3kw4L6ALGHgaNeHQKpSJUHLEMOsbZrddbzuWzGhNmv+
fxeqqRmwLcFGTKO97jsIgKr2jLE9h+PVmHqtn4DRs+mTRL0kX0cOG8OMwHnUrOrS8fITICCM6upr
MN0QTn9VPJEuJjT9lFKdeDcpChw1cgpSv2RiGEZ9yATc8Lxe8pUZ7FU1Zx5WxDJXAVt7z5ZMmuOq
m5gMXpPrWEcmQARgRLqzR5wbf4JXvV/FNGdSvbGLt1LEyqNponeRVTT2tMuR93P8NxX7ZylKhHgq
eEnb9PnUBIZSXh8/lVVUaldgjrUqZ+P6ZD6gMxVA3M3NYSNV09K20YokQvmmaM2ZLuQpZ7zK6P9r
YQ360wxMOFbCXfIdmEjMR7sGsSAQsFUqScLZ5qajAkLmLkgiZnSBLPIMEvS04AvwGifVeoD0HsuV
vrs9QxXNCdT9TmWZSigc1YNNp2inednClJv4U9ro2GJ8VlepuBamXtaXffESE4XxokNF+aYLQQeZ
qBnH6K077mJnVw1eCjx0LiCVbmQs0iYzKufLGR86bg8Cm1AcF9JdXdip91fixXq89kl9AgHq8BJx
tPQb9lButdykRhbKgNg+08k4g5iJuSFCqtLseqWxdUOBHiBAoIRxjZOuBwDo1/eXUdZGeMuR63jy
1Cui9yXJ8Tl8j4Gs+asuLSYREDh/I7KFymgN5Hv4Kx3e3gZlq5pB9DoVZ041XahlOkfuWQLMHQgM
P0oHY/d5/CriMZQ8SaSZT7Qsi/j2Uava+J+Y7cX43TNHGUu8t8bRfUwYPahkG8mD8Mpfo6X5o5MF
2gm0PgVYJdriqKniVaBMXaNqkUbbckqsX7LsALDnjxejwOi+0lHFKGrZIQvi3+BK6i7/KyqJpocW
THgLvNgZah8QQ6K1wZVDgIQB15XbSWIGQ8CW8kpjv/grgdikhbgz1la9HNr27TBy/X7pxUEgLLSj
yYRdp6ergn5rp7j6siACRvfhwxkkZw3FIx+CVEl7DUQ/dcc1CvVTsF+aVPmJPG87zxE3QNsZb2kV
7NxEojfPSHNHTqGxILaeL6DzRz5/SolS+rxfLbXK8CVVCw4wUBgiOztEPWgS6I0X+QA5r72DzNvg
6hjG4qXx4evsH9zuAsspRBRqDFEhHcZIFo7GBz+sq+dfc8WLjB1TxyNEvzxHd4ajJ2bQl7K99ZnM
nxGqwnE/tr2kAZ+G3y5y6DWda2BRa8wQN2nYfbpENOOHC72sstOLsj2GzJI08m/ugSbsbOx3RyU6
L9gI5TpZQbsUzZNgMUCxaiFBckwxoJn2SMMGotqx9a9itCzICyqEDrlbR1GgzfEvu1hCvE/93teB
uyJKJLguEwbPvxB6IooW2SNbagm7orr1NEKAihv1G+hdKtd1DizWbxRWJHY4Yk0fNfKSYE+OUlrR
QaetjP/qkdrUOmtgJvdasRkkK8OYq16+whuPSRERIZTZX0b3zXbgLHQmChZFCIp/Tqri8vY2kA4k
2Ku+ZoPllsRaHGvzJIrLKfBo2en4nTH88QobcCAQQ2xSBGDO3ZZ8r+a7OrPg6MRsSjOSTlcdSw9Q
yo2GGUGiQQQrrm5+daqXBIWyXJoN8plOVePs9bFftKtkikLCi/jZyGYr0/07l4Zzh0rQ8B7uqjZY
olTLoCqWesWF3by8xCsLnyq0ERRvXHbvpUy235MV68FujypQmbQ80RouvTFsXKXQRqW9AkWaJvek
FVenlUFHieGG7M7vDK4pZyXkboAYuAhDW478X0kUw1CxrlJvQTHcZDC/KAb5g2BPZqML3jx8nepG
nUetKOXCwzO2zZQMQOGmQDRTk3BH4pxMXTgpfn44CI5DdfcpriAZPa57PTZYzNc5aSkJ00vP8FDc
+URMs3t65w7S6kBMsfQY5Alj42UH19OSNfqLX6R8A4gTFtn+7MM4UtrjzvygNdyZdlxqNU8h7/yz
EEPuVm2UJnYPDSyJfR9A+jtAnk7OcWbZQWlVGOsDwUjTlgbn5VL4lj7e1dwHl6DwE2aU8mzXeu1N
HfTukuhLcrnel9jv9Gens4WBhG7d8fa3FUYyLl35L8rIqv/zRhIOoYgm6Shp4Pg3WJnWIuyHfLDU
9U9Psx+1yTOLBV3FcwfEeU72teLxDZn6KE1RJk08HA5Ud/+LeIz1Fo8pR8zX/Z68W9ThPMw5EL1a
z3Dr9QgLcZRhWAupubCa1sBSpAHId5mnYGNoTt0jsEnjLDC4OlUp9BYy6PAh0o/f7CXoM+ukNiYJ
2F6EbFyGpEfMH+GpOhAOwk8Pb3SZi4pIiAbS4MtaK/8AAuez3Pj33jADfjbdcGDwSOESIplGzezw
4G2T2SzEELi+wKaNpoZ9NQsvWaWHXwXGpL/VrUJS7vuBXbNneg2j7AEoZKiZhh5JMRn1Dosue8Ve
8tYRpdPrj9oqqxTCYmWtbvALtO7PTJ8j6mbay7jUOQQBmsG8d5onDZaviIopHDfDEPjCwrtfhgoo
+/L8Sl2+EQlzsvOr98FKRvKca85Xlv+33L78vaQCg2Au4mpLzX+Fjs95CAROx9EdxKxLeGQGqz0P
bsTmMOwX584XeFRY53N9w8w+jPbAtqS3Ibr+Ea88I+NGU09fgXv/JRh9+in5ELD9L9wnh/3JlHVU
m8jb22gdp7OpLoQs4u/SBqYsLz7QsajOn/byAXkfyhDzSUuhuD4ecgXrC5280sD+lHIcIok/++TI
AVvA5lFg9HcVUahX1UxPmCrgN9z3pWPYcdIS4syNWNf/Bd9HSJucsq/N/hmOUPSIF1ESq3PBIrO8
bJ1C7eA8pfDahxQ8NHsvg8uGmLgmnvtbuD19mCKIPs8KJd9joJLX/ZTtrOkPoFpTjOQKPWmAyU3e
vk4RbOaF6uOvbBe8xqTnUOUWTdx0QDPuSiqiwfek7xUG18dwuZEGTYQS67myPjEZxuUpA1OgMomU
ImlXS4uB6nZmqNCA481iWvam54Oc1G1wBsTVCsiwTO40mafaXfFZOOiAUtoOMeOKjfkd4DZUpP5k
PYXZw5XGqqWqbI/58eFtwkJAJ3/FP06oofquZ6DeUSgas+vIJBGyerkqn8Q56t8n48RO7SwKJ1Ka
5plwLoZvAbl110Qjuhm5WfL1SBrCGb0JMCoetH68MGgWXkXsIUneycLPz9r8aEHcH9Dvj5opyivn
2sI8LqkZ2HPTJdR5S64+fvBXCaybpRgQ7aq2/g6TLCGTpF9RFrbtbxn94q9AjE1mNbbifEzmrWhc
UJ0gruRZYh9zemc9kpQDqUqZIaI0jPfXOc2VmMLeHiAcbYqyBk/4tKBY3hsRBeGx57XW5F/C9Ajn
MvC7Nynu5pQapIaDwG3soQcYqDx6tshKWy0n16Wy35PMgAwdL21/DIvtYWMHHJlcasOSIsQDUAB6
JJ0g909Ou+o+Q0uI6YWelHGUiRdh+DswxnFjd25H8LGahpMsG/tSiSJo5S+lmYylEZRKsp0ET/be
ElgTsKMsW7Rm97JP/2vLphWHbgvl8DizKwQDyYJR/FnM6cmQ439klzUWq2VoOxHv3u/EXdeyYcDr
cqrOoxSzWmGGJtwAne/c4qf/r4ad0eMebaaGESmMRSyfOLyzdKC11QGmE3BlIIKbLjRdjZINfVbi
46oohqn8MpoWyGef74vzN/8+/mqVQ+1N91Pk4p+yjST17pikrMKmhxJEMZJFk0LoHsL+PRA7kzs9
TdXKmmqlLw9NxJ/YWCTbfN1D6T9DwmeE2p8VP54W8hmfuqc8AhgkA4x2sls+J89ulPifgI/pKnMW
n8V8r7kL/ZWTLGC56ptX03PRIzHENKLBktmoxvVaaOZJWuJR1zep1ySEfpgDlZyKePGFLZzoPf2B
Yzl9JID7JEShOZGYU2FHy9cVFJuguafzWQDNU/jfYhrMbs8h4AVyAUXz9UOcJVL856CpuayG/hFh
8ZJV+vzrZ338LqOTHDbUcCWA33CS9epK22xkkxdghfHuq5TC5chs8Mm6MGXvrh6pnPA0QVDYaO2z
RtMFmxgtRUivYbNXAooWL/CkmhPDcnm5Ge21oAMpFfJbKBXIa4wcJLaPJx9y/WwXXgCuSJUUOmsf
/Y6t85LpotKfCwk79lqKGV018wpnkWIDwTGVMnRrpsnbKEguMsu8YUY43+pbXZEmVL8pNcTAFE53
Jag3Jf3lDpAdOBTZ3Tl+TooHVPZk/zj+Gz7cevDAjeRYRf5lTzYJgPqJTjVCXoVYYAKAO9M5rTcT
VN/h6sKydBaKIts2TLHgfLiaRn8uQJ//ZRaIHwEBZQFb8qAc05QaGk6zaidCTaxK7+uGDlqFG5vQ
T2TMPR6UqBTbLE1koYtBZ9pq4imwhtLUfC4eVyA23ThMpTjkmo5MvABDLBrOPlOCvNA6S4kz++qk
q2jD93aqaRi7YgCV27wnlTZmwuGVOyHu+fF3ptH3EEI7AmC/1E1vGrJHfs/ED/4bPIL4xLvivaQZ
yd0XL+QdOyaXeo5pBgohWYnVFYMAX+rlNoUsxSabsPboL7jiV8URQqOAC8gN6CICzrHkRM3H3ZwN
/3cffktTr3258Inpu2M31NW6Kq/i1R4nPpke1+dlnWVE4ZAP31lszBthJ/X8tGPEfz99H2d82KJ1
UBMRPU3xLxc2fmlGeiuZtJBXsVs56vmQY0hBBcORSRccl2nwNqw/9IWuKyqHez97zcOrQ0uLIff9
p9h0LUMU+O37M9cMljnr/CqilxJXn6x8smSh0sfEVKAwUYhCt+jqxsgoqjZvbvKHkdH7b0cy88C5
vmVg6ZNSgO6XEWbZ3wJQcRuMIQdgaOA2h9X+Ko/3lSAdLonQwA1eM5F6U0ytqDe9CJPSDTZxZCfk
eJwSG126J/QnPVo151XgSSZH9JUGWhmZoHeJ4G1ywmr5sZXqQSWoJb89+Hj6I8C4gqpP1dGevmop
aWHLhnXtgOwB4SCl9vMcDJ+THfxs6iCCe5q04OMRY6XSfUmeAfuqYHLGkIjq/WUhwo89C2hliwzN
7fb+jsAGO3SGUmRuEykqiMXz9FNNBGk4pxOXUeqUhHNNLdoh/RjAO8KL0Y0CzakVNTbKnYH3VXR+
y7GRISSjo9gzbqCqj+noDXTrfMJBZMO6rTHXdG0CPkJQXDAzMl5aaCVU+lxRisfr7ZIxEDsXHl3Y
fkILZSBwX3n3vyAHIAFE18ypptfsquu6g1fzESnHeJH1wfkj7sKW5PkR00OPG9uiQdsUpvtYXDFW
13WSB2haa58faIRk/ve/OTi1hRMbSu1hUiFzQos0AxJIycFqaJ7skPozNifpIZ4pelyYQRg9+SJg
m0EIgYCgomfAkP5SYEQVLgCM/afHmqxiyIHgTyZFqNumGqoc+olE9qDbMII7uRUpVpKZPaDLTM7Y
VxX1RoFZ39hUfEHTLVnbwlznZMMoODz3pUX8ANdbqEJska0e4jFXAHLY7V5v1MunL4AHK5q9UZRy
8q1QlZ8HjNbgzDZlsLGXNue6B7FnwERSgOBvbZ1z8IY7b6MDRM5sJXsEyiUAo8PYb5ywxCyErHQR
TkoD6sIv3+tmDXCCa5DtA1lqW6J1ONUp+7aRqQ6VVb6DijTt8UNij4SbRN3jsWCWDMe43SXzkCcB
k7dnZjFajWU0vlKoIQjJXSpxQIYivQTNRUCNw1nLWZuORrEybm97MLz11o8xN7653jLpSzkH7pOk
jKutp7O0NuplPpMTUuf7vS1yyXueobzbFTSUiX2EC2hKJfAq1taSAdFs8rH/rjxXIWjugd90D/T9
/WyGOfUbHhbMs4PYN6vLjQKV/4ESVjXNUPVDskTkk3QfLe5+8DdFPonVhMe3KFwFCdokrWPJVWEb
8TgdJoS23YAALAKc5wGmcTCJw6JGXmMtAL7cJF35TyUJ4yV1FJln8k5ISUnmqtKIKvcb9HBL64a+
PCO4lrNIBHGDuKVCn8VvEbm0swMC6uCnxoFCdQLvjZotwQqMKe7w1v5YlARmRmRWa2Hn7d26d/t6
fXeW1sRyLpKytZW/SZVQC1J6MCQUWoKkjdM5uc6DGs4LdG+U8f3V5k7rlef45L7hNeNHuy/Kuc18
yha0lVWQDAEZ8C6eKl2TY0vu9lqFy5DOOwBxrtsTgVQtOpymL4+dYJtI54W7g4LWm2AZj/E0OqlL
/EtoM5UY250+o7f4Bq88lCqlUuENu3KjajYSHUiqMWCjbqoleVMznNWK7ywCATj29M/U5J1Jefyd
W7tLt284kw0kvzywdKlnTsFaL+9yryxBI/fNZWtYQqCfNExwhieTwvnvBYLfWI9kBdI0lm52aSx3
BrOQPhlvyyqd9uQXGxJ9heZtmgr51JimOdjXoDQ64nBNnCllL2e4LHXqLZoQyRL7Sgmh0XWr1Ixt
jCYtqcZ+QYrtyup1RDj91/YrXD6AAypGdxQc5dW3kdC0InWuFYp1eXBa8nWBj7gpx6GXlEP9Oayp
KBusVCpywf0L1jQ3DMbux5bU1e/bSo8XiJ1gg9yNcNoczQnQvBz3RcCdpi0JsBxXGMXBHoPpqD9D
aAecexyn261REBmFwEWbll3NjHlKVe53StyTEvo7lVEL+v9tSr7iSdWCDT9ZnzjD6K1QjJ4PklKu
khH8sotFZqUH4vQ0cTQnpZ9gQAgYJe9Xmqm28WSF+GD3MiY36HEz3qwHadyoG+PfnOk4+JxYVldH
myyaVcplBFvOCSLjhcrg4jPQZH7jbk7KUiqvxABRCQNX/B/nwInJ3/K4Jv86xRsX5cErx8ks+8wN
3cSUIU5YWwtzoNOs6WeJFsMQHXh196kShsRnAp9KuRfv3rPHG2Jo1gk7lqCnJ2qcyENXMpV9qwyB
nyfO4HYAfJUQIqd+lQrXYuTRRSYP0ucmuK/N1fCehlnpG8UOryjClFNVTSO4ZjTJdDtKn/+06Dl5
AgJ0ZFbaB6GtEsJ+knakf7Nf+Mov/fwJyR4HvPJwS3nZ6b+sZ/HNpMal9p3xUWzmo92WIvrAMdL1
ecMP4eOzZnzCJHq927/XWtBt2eAp8Wlg5laV5raizQiA88ci6YdvbxZL/c7HIzSS03NqHKvyPc3/
SPlYFPEDc2o81DX4igVTlbhEEESzRSHDPirJ0mt9BXOlSQR43HYka05SUBtD3JTYsf+6p8D/2OFy
7lzojbEHll9L3Vy9KzqUZRfLSZP4uzbXxc7TtZmA1hdsZExwaS/fqDwlhJl35c08S/Dg4nMET17P
UbkG5ycQwf99iQz826q1kNUnr9wWGjryIikiYXQwp6znsi9ClMQuvWIHU1NDYwThkNOOrBIHp3Ai
1GTnXKRjK0nFiBDCB8jxqefpQgOqijR90PiBgjdmt8gvXyEWKreDUTowZgR+PIgt6A5ZX+3KFvA2
kEvXxHFfajE8TTbGKjnzRSGnFIVYAuFhwREQuuqche+L/V/c4R+bZPjOBUq1icRqEdD76dIW/0LB
FvomaYrbLyU9CBpvCb75DaigKhYI6UMAZ8afyA9m9KS7G+0YuWLAqvXyT/bK9uWkyV5SazzShhdl
KOuKVNU/6/E+bBmbmn8Omh/uvRQcPj/WJzTr550emshWydQ/pbtYW7/zDJU0X3cxYb8vToIRNFXv
Ss2W+WaocEjbBg/ll6Sik7746r6+Qx+U0OMLx9MbcDH1GtflUHel0DqTzHAYGwmiKY4Q+zrIYcm2
pMP2UJ2XRtS1Elxr4mkMuWywTJvjluvgneBM2tUEcbqNPZ5QovsIlhqz3iW7mUsgKI4+n/919/el
0AF+tioG6XwCRVFrarw0ROIkCC5p7I9BhMipFXo1hmUJmBGU4vMmwN4ezN9t3U/WoK0XHMfCDys0
mTPaFQ5zFJs3G3ZhLebUQGUZtjP5LWKwfV4WeYLJ43ptYh9rHeE9FSyrwYvcPF1X0WNzfRI9yjo1
6atknPtO4UrVnBoSK286wR7muG70msSZ8JRHMO9zVAt4yScHpWippv9P+Gi7vgA+HBGMAQpu497F
ss3FoUOQkShmosPCSYziVD+lFWq5+JpLLSHUqhk3HC1a2Tes9gWbdZQHMwvEenQpnl3Gi6Q2TpBv
eZ1a2P7a5MFe0FqVPhBpOAzJpkr+6gf4PL45fZi18I6nOV38ev74c4+MgBjZTRRhsBDtL4dq190d
r+LhHX4k1zS+mCCEbED9QhI/ISgb3ETRT61+4Pl5S7XYwQsR1V3RcgXVkSnhZJ7KB6xTxdcvVveL
Vn8gRDtfAWICVBqd5Ey/kImNe91jMUvirzfJBvmCqOW27liJipYmAlzazMu0kMYLAmvjD78lSoQR
5od00xXgZ9FhLhUGBNiIvIFncF8gG2ioy3/46CxhYWEqtjh0p3X2wyJr/DU46Z4aV4Rc2q74tr0q
qydt0sLn72d5D5F5JIXW2jRCHYdR5Rd2YyVQapVcIJGCd/JtdlcpfPdSo6B2A+UHgGN61DBB7LXp
FP3neRIw3iv1B+CTq9RSG+lRl2hQ76JzMUWLUlp2Qv1T02Idmturv+A8GFTSKdap/U5D2I/yyBDi
9NZtWJ2WhqFL7JT4Ovbgc/VGhCQoFFtcDhwxRvuRvIbhxl5UZpf6GU3DV4cEJyFcSUpjP3KWwsEl
GMirtHG7p1Xg2ikiUmZhJkI47Dpyhp9dM570njl/OGNzrd/CawkHy9o5A540oW3j4bl69FhjFit8
BC913JMQ4DwJ66bZVS96A+3YvtwcNPcO5IKIA1Ki7irySwBRH7pC39MQpqE8Brq517lio2/M5KF9
7c41E+P4+6zrWUuGUv6R6vCGsOT9PlyzzMZgt0V2D35N8dqUFQpw3aIcOWZZg5E9rd6L0Wcg7S34
bFnIwXjuTOXnFkXfNx7c2KmbP3kVYndYp+KkA9JgJDik76kqU720adfKU3k/Vum89otwD0D+j3AT
g9s+dKjJpc3PVxD3KVVZkeJDZ8daqgMFz25axDn5K9IlRu2ws/hnuIo+RsEjdsXM/MFt8podRz1I
wy6PuWPGUMExPj0f8nxsey9fYaTd334TFP+kBq5ub1hWeKdr73dYxT4qIIgNMTM93vnmLZfG0F4A
cqfEccthhNL+MdCI+oPCWjMkTV7xZbEFCtvZGDMkyrY6Kd4MkapMtRlgGVXjWNOTmu6CdtRJNQ6j
px6uO6f7y/q4TxYhoE5dU3yRMnqQMLP96CG2o+fQ4/hSUkKfnJDrojxG2pTAskLQTZqW+LrkEkG8
OB/sqCoJFBjPS6MpThqWQhbJfTG7AZ63bBOjnDhYE465Tdn3M0o3tuwzLwSOw3ddnQp4xS5bQEPL
yhsgnN6wfjEUgH1yAqYGSRWl9Zlmh/VzkTA8TVZQCIzKbXub3ZxZe2Ts+Cz/weh0jOlwjiFuNOAC
9Z7z8/d0pQuq4Coza1mx5V9p0hGvlXxKGPLrPQICJgOGoi5i3GGGPf4qkqoDNxKEm4lbTg73dARG
DvHGRouvVR4ZylcPM3e+78mCMFchHrOnFr2Oh3tYaRnTr/w85EkeL49ekZA1JkhJ0SARph4eUEvP
OY3GyQsL4empoxdPKa5IGfI4IFq1O2nSoxAK1p0voErw8RM+8GTwAfVzKagQUlQpsWl33AqSr/CK
fqB8yUfd+X/m6G9KF1XjWkx9ANA/VRH0U+f6xaMzdV5rjk5/vbX2u5XSLQ7A0yDvPH7mI4nuvU8r
XqPhz7LRGByGMrjsIFS4TCLyhKCQehT8ILLB/6x9QbaawY4zA53BWatkgLdWXWqdrhOaXOsCBUqb
ehKogyV1URdjbmgdK/O975YVSBf2NUCgfpP0lmrEF/V2y4CWXRIwla/eujNup58+mLish0KoDVvP
EoBBU5Bq/uiKTU3wBHmBh4XYY6gKCcbwyxwtsTjXfvEHfhk4/CSEPacZ1GMF1dn4sDvQSUOrkYwO
3nNAhH5RDd0MwDdUBoXxO30GNEgmVwaR3k2i4thYJpO004WPhJ9veBV1miiSscNztUvjDfu3kZRT
0BXvnV8vG4mnxMWnOnmq6j+AOxB4lXVlU2Q0z6mNvsrgQqvxjbttYBwVuXRgiGaNO0dPAS6QVY7o
CZ/Mc9RTzsasBWW1Yp04tSCbeVQzf22NUL7jj3ZnngEZ14ez5JMP6WPH5crabcnk9/yvCbNzA7AX
ZJlF7eMMyg1ELzaN+XoP4Blfz3A+A04AtdHNk6VlH7Mhzrx/SpbTfpUnb99SFfnkWAbTPdjgAu7O
HKTETfZeH2gVn0MF2tmXdjBXoPJJStNNnA2Cp75n+TDbYESX+ty6/kAJrKGgdsZTja3ZLd8UkKLL
00xxqeudlI4EsXkjfNeq2ow6twlARDxwn7S3zZXbLjzKYJxn2XYcWns1pTp0BtYw45qBO54BfBla
y8eSq8cNFaONRyiAsnpE5AMHGWraAXoTErXmE8yUj/YP/YR2Ft7pCQdlRH+Ik7sMy4WC0qR+HGf6
8wKZ0SxatKbInmiP4E9ihHSggxFIT4Pn/xY3nd+zYH+pFQCxrm6l7JFs1b0pyh6Ad6pp6f1RT0sL
L+W3iSaQdz+2bUREPD1Z8sTf41W5BIYIWkYhT4Oh4zqWnXsUsReKQAOXoSTNhI+6FPiXN3qE7AaU
zQebLcNtvqWnO+Jy2fDpp12JGahtes1crgB8WLZ9JQ7Zpq3Kwe5M6DlQyESorkdAg1SMK/HkQxY6
QlIQ8AZw9AWKtjuRDIVgIG5aFLPl62E1iLWgDyqlkqD7tLbXbFSW6w4m14o6cKnb1/sN2lVDh78i
lEkIpuq2wksGzrX86Fu5Z3NC14+UKX3v710bQT/4+ONGWKSxpAE3P/yr2na7Q3TaNPVJty3euBv9
hA71T/wKHGjdkYdljV9FAttHZVZj6kXcwc0yiUbEQmeQoFHdF5L7moHhs4ROR3is0LoqKmF2qwV4
NxSzeYwLX1ThXEKWleOGo6rwiCwnAdEKPk2H9o3GVtF1XzS6G5RtqN8W25CF2Nv9qh86v6ZHthNT
acYp2Bh9Fsd42ZgyaYVVKkSYs6XMdXXQKHricetirduorrTh8Wb5sOCXifSLETLqy12/fgKX2wKL
tRoAdHdqiZh5GfN0MAoDPvkUMZou5mO8T/VE1zckVElz7royW73Uh4xzu7ArnK1of1FCOFxlYCjY
P57xUseitELH5I5qnDyW2AlKEw5xai7/glJfEC5aAlIi+hdLnUr+UoxnbqmCY0fCQxdFDV8rY0qa
5z8d3YhwDP7EIwd9uhcpR6udNYUpQYxw8HtMufCQn7OdNzUO5rEerMvQMPxwM7JXc05QkVIzuilb
XAHCQnVCgIfXGzySrNWtrVpTnwEW9HtznzOBfutm1X1y+SEiYVKLsJHywIkHjznPfofjvThGJD5h
lnpcBgeb9gakgjBvEU8yXj3YMotw6p7vHD228m0hNaj0Jljh/GhaVWrTc2IkBjEUdQcdPiVCoeIz
BENwoNi95OohalpSe/AsS+JpXl/tAe6P94woz30FqU80yDGh+9tXU0ltJIJTxhcf6588/31aX4KI
noaMpqbtpDZ2RN4eWpurUSyjwaZGtJVJrEK+GVToUESslCdDEw2AF8VqffBLwbDCjH3/XgOTxy/4
BPlb8+irsoAfh0rbqHRPW2Ae5QRIDLX13Kr2JcXeozhVZdUQnc4nURqjLfWKbpa5/6uPxX1JBDKM
9IYRydXv2B9ffMzRZ5ZzJREubLXBpbA9SCbpiV5wutbBbN/z3a8nnInp/uvcIiQM8A2GDtLS4wb7
Tgag54nsZW1H8k5NjP77FiI4prWoAGMhrMP4rBhQ59/iJ66ojiIym2NnB7C8lviNJPX2MMpGv987
XFk09ZFSJ2JYK7svx3rlEmoY856TFoCV/liYVVEsjXBEmIFOJVxjNab7JtymMAoQM9NjrWjxHeAH
H0p/T/QHLrbF07i0ljF1Ayq9nhzw1nyUqEHTNtM5V2X1l1IARSInULugiUZmA4aUs2dhjQ8+G1dY
Ic91AOOujQ1e03lg3yUwHLImkJhoCLhv3FbcEuP8j9x4d9cu30+GKzPIW7jWqrx0iYNrfsMdj3uM
5TOga2+EwCN/rQAB6dTkwCeCAb6If9PtFsfiZfBxMBPc5y8PuExsiyDnfS1y0oysoAHcBYKwO/Kx
gbcdHq9gkI1+tmHb2ceTOTdiwrf4XR0zJjsnBx4dHEsjWfJQFOcJCf0ca1iEljZNs7x52pX2Kopw
HDuDgwfPGiqMxIQWGJb+ihdTBjuZEIAmmtL1l/N95pFOZAXBzG4v+CUt7T5IDqYUnC29Aepj2M8x
8TAd4VeD12DeO7bjhKMWpp3yM6LlT4cLrGQjs2yikUGExNYha2sXsYtYsFdGkA6vYulfHTQdzOS+
zWJrlo9yLTddV0NsA7kGAJU6LhBvOZXW4x0Bwtvh7VK2ShaXS+YPWPDs8+nayuvYIoDKbFS+OWMH
DPi2vZqX2lyMIrMcKivSC1F+CXpI/ebtCYoe5Pzf+fNoDfDwqYUGkUPGWEaLHzmofyYEFfb/g/af
u67E7TkPip1xI1uuyGrMrpZeZo9uXJ41CP7phXD34fqP4npl/aPPwnP31U0g4FrCT7Q7D2P8PtKF
KBUE43n9Y0YYWwQnrhwPN60VOprY7PxPSwgis6Eb/+OIYux7wBTJfLLTt7OfP83BKlmMLLfidovd
wNRDW2WfzzxAGzfsBwLSqIkwTzKowkyoUYlZGEGA9rzZSoCZ6oZ0UeRrPLI/untFb+x6KVdZ74R2
Pndwob5K1XAUWGdmLgD8K2FdNjQRYB7OVVHoO7M09KeaZHiaTBaXQ8cMEfG89I9zv31Kf2Ch/ioo
yis/K5lmuuTJ1aiGAuTI2AyQR/LlxcH+dIPorrPpApRG7eLf7m3VDCAAZpO49vd3CAwSs0RLvyDh
68JlLH+JilyYmSKPooEB3C6bm2ltN5Ihh0pVRPPSePZl95py8/LtYjIWW4W56tBmnqMpemKstwJk
vzHVMPnWW//ow8mUm6ROv+2U0Tq9ZXrpezv6KxSrT1nellasGnjUdEn+qKujCgAYVw05M5mt+B/H
oUh+wDve+BV4adT0XcHeb0ZfKIoIOoMwTqUzd+hLtdOajBWsPDXW8tOHbwYVqOXJNWkjfqTVhjo5
y7YDXsUs5AZlL4JhbtH2enmC0G8rbi+cVZqNjtoG2rTrahsQac2y85D7/qZrGtdiXiL13lRdRfvv
DFh6oKDvAWKNtR+3AmHk5YUOSxHy8aEfsY/8Ngz3TLBlzLpFHmvamoEdZYjzsa8UeD/r8obRdCRA
KENPjmLmgqaMi0q3BtDwQLUeE8HIG+CqFOZbR5PAtnHtfFlYsBcjCsv+eBW0dRKAAzDeAEHXE5Z0
u6m6jlBIO7+bh2HmzIw26dop54M+8Yrt+uXq5sXKchl80SyElw2iyP0XdyhGYigfwrNyx0CARQCB
l/IywUnG2y5T1IdCvVYSVr8+t2jW65s5d21fFuJ31pSVFaUMsLPzuNEX663d08CmfWjvigLNhIP2
h3G355ZVpn202AVq7Kq2w9KIuPggOoF/xpEWgd3QSxxBxeuBVCh8rmN1DA2EZPQXlKX+QzGaaz3I
CIorm76m3ppH95xdqeQBbd8+mwZhxP3NOPD6KwsEaINeT6nPT2PQ20lkd05VzRfUaVjlx9hVbYOI
NJ78HMuK0LTIpxWRs2Jtwj5nTJWhHM7z9rApBakDjeIvhO8RpIUZlB7nxtCyPOGoaDzkC6r02Du7
tH2IWRx3smCPnLM6iBShfiMQbfUMF/6ryYr7EiHAPWQQ3YkYx/+KMt05tDPyczN2lXOCZM5lwu2S
7IrU/h7KdaDNNvS78NxXym6dmJLlz/9lBL3lj9OSXTZXp58jZ6genTv9OwLK7LS1+naF5T1tjVYL
ktEW9wO1gOuS3f1kZ87HM7rg5krubpPXbL638MYM69136zI8GEDtJwJ6v5BEdd6Ay4ucyVdjUXQs
qiQgDf63flF5zAi8wafTbWu4Q298g2h0NkhtF3e0MIEwmlzWwfewRwlWWwSVY/z9PgQTWb35y68x
AIUJwn6wslw+BHtfsiz3orcUn94XDcHk/nI+JdyHmvMRN4lObp91yyEBwRbM0ekziIZfgPMsdaKL
ZJiHYeXsDpaDgB+ZTKjnN0oetaFPizUYXqb5U3urBxIr01e464Hi4pAQMLMqwMAyZS+kNwkNMIij
zDF69Ceflm88/GllOPV6K0yytLVSMcxjNS8vsf2LT/lJ7b/Mm6YK3lhPrN00iWqaiaB6p+57GbY7
VHva75Fz8bfZ10wonHHN4ytZ4Y7OFz5IILNWflacHAEfm5SPl/ezj3WwwqYNCjMsjrJCB+ayqPQS
DfrYt4p7x2GL+aKcqYxoGHf+nWBmlH/tgau3WnEuhQLH4ec9P0Rcr76K8SC92iKsjRc3C9/pLbhf
y3Gf7b+q1oPfIq8eVL3GvCZPOJMLmstcpweeG9thf3+MxYhh/4umMJxzzNCu2Pg8v2MUKonYrJRA
JhjWKOkQkenYyGhrEcBhiTCdR7lVHrleq0SEwNuQzn6lVZ50Nl+aD5wbmzIUrDkqf7mgHaXBu62y
SAgRzjZKzx0O7QQ6W+cXcl539rqG/aCQ8ltsLxu+rgHVilTUsxtI+ftaw6Db5P6ViSwoYLf8H1wE
w7ExioGpdgG8z/mRUVA94kVQa2bxYNcjleQQ7L7q+DrU15Ka8ElFjslV5OhyQBuOQkiTwNd4L4Iu
WiYrR/hXvUjDaJTMVLQOEkalxBkCI78L/MLEI5zN5lm80RqgMbz8lW4H1x7tcfu2K0SP25vFND7s
zWca4UjJ6DswlRJiCPknSgVzKth+MrzE1X9MGPV37NFkwcFdyOOhP7mA7iujE3j4xmlLgpFsKVRo
m7OJbEt2KSGpvtn8CCWf+VCjc0jtGpc5CyblXDggcKxx6x5lvTVbw4IW29hHZpP9AUKFivn9C/yB
c1pOGJDejtgfUqYbpI9kvcmVnfJVYhlQ88FJIXtbz9G4nBTpC9ayhSYr9/ZNyx7fBBuePnnVVpS1
AkZm5HHKhhr+3Csa1HvM3cb1MYT9pOAm10E6kPR1e0ucZpLrVMp4iZ9RpY/SsdlVQRG4KsFQpUVy
3/wZdV/YBD8Hjpe5UiBk9OPaTlaQwUcPTilsF6CWm2ErxK5BKq+knqaCsUuY0qp6e5d6Wr563Wxt
a301+hX2qgorgfDB1iMB54uyFxPoRVCGn6AH6Elhm+5PkyvykDbPFAcrg3tHvyJEnlMb682IzMrV
OYulTVx3gGUmH8I+oEE2ZYW+6FjW+i9WGcmDSSwlsy2SgbDhpaAeB+k9S/c6AXDefYM2vvb1lvuU
bjlCCK52FHbZ6FwNmwVyD81Vk5/dMCbCGi8fJD7l4OpswnqfuEyKJqKjopBKG+2BKBVxnhNFntWN
XWJ9x1i7GBbm/Ix+/H8wJD2QRI59fXjxvwjUYeNrO/fFa+pvtyqPPxWd6IwXTZRZHNcuEg3Ehe96
MxEUUzr8uWG+MNuvDa0+Isu5AEspyzn3CmKU7uicDS9e99cLT83G3r9Nj0oH9PsYZasvzO67Zikk
mi+kabW1PlWzXzPUv6n2Nj1/dMRDhteT5IOcgVu6fJVTj8+oTOYsUmXMorDFQUqO5+AK+Jawjlmr
EdhIY3oCOSH4EgimmJdKdl81DaxnYcHYhWYtxqnSrV6FYlnwlPsI5gpsou9krbvaykw8OnBzWv+3
h24PQd7uzm1lWAPp7EY6HxXR/yoPM6MwyAAWCo0hHqdqjoLCMvobdJ3yHdrLEUoNLcauTvi1lzs9
RDQNBYcAh4cdFqQnpFqNUKXEx4HoHxA8kxJJmystKeGXyRQzPQCFeYfZisAnKDT/7Vag60tL16Iz
FB23U20X0BYtom2lxdWkSNXrkGlxUsG4K0K9vOUeKyM6UOLhZolLBeLpAH8Il5LwhBAJXnjPUyBJ
yzk8rCJKUKWzvLDsqXXUxxY5AVuSnxoh9F0if9nXKR2UJNqA4X444ZNsafiJoSLotGvItU74+MhK
O5p33ajdRRegyjjITeaOPnXM1rpTW4kbn+7JYNxB+c0ICuoBN8v/8wIsGtYFMNb0y/XFso4V7bly
ITshaSJ8fB0LCeWBY/EuOc+K3xCA9ZYB+JGbO3SK1Lq2e8kMsrR5tZHJfNrAoRhk7eFzkH5bOJql
RtCkF45ZZ91kIhEhc+fEq6Xw32KJRyp64/i1Dk9peB1HOjPpQOgAZYS+cyWARArpGbcE0hxcdoZ8
Z8ZOmbF20DG5XM5BphKR3/BVHR0W+Fza1T+3pEStt2TxF1l0ky8N9jVc867uNzVlHLX2rfNNK+04
wjypO8idQ1RKmyVCy/tCQlLblTfvcymsNg5W1/w5E/55NZnjdusFcRBu7Z9UkHSawuTjwpSin/Fq
g4G2trhcvfcZmfEkLnY472o6KN7EeHj8FxTWA8gli7M8tvnjMu6uBBIyvc2Y1xcdfkCd42gTPndo
0P2iiHvBM3iBh7VmKCh20c3JSr6rwL0GyNbBIDxdPxyBCItTGbM3h0oJug1hnEOTE5ZbJTVjR89X
T4sX3ZpdP3PWXPyux+alqASRDTch0P0p16qS9s/R8bJoutpiB5FdpW5AMbfq1JkTZVeiMXbsyObe
TpwHn4ArZnj2MxyVnbMfY87F14ZtTEYnJrIsTHJyxsXu4vr/TQJQo7eg47f3As7iyxIrv41tR4mp
8fL4BEnPoUS4Irl5mHN8qK/m/1CnlQ4eP5HqkRQZrluFiMsRstRb7J1ItPxghSD6xw96tQujaat+
EUAkdNvrI5oWbbzQG9KHfjv4uAGFhxqyTWj4LRFxUUOqrSMSDggcVuCvSQok6Plo4NlvUEmVLWY5
+F5BZde3B4K5OIEMoawPiW1wFG0pTdXJacORbx/QWn9ED9Exg00ZBKeqqMO1O6YQrNpHZe1fqbd8
mL7/mk0iMxC86sfQDFYMMiUjcI9rUUCPdC/wc+Ci3lPgCuACM6+YLkZMLaRZtukX5wvyNrdBb38T
CtSohUK8IPNh6VMXk0Jsdy0dPYG6s0AnqyY0cw8ncRhF1Or7PSG9GeKD8p4LWYaHXVyCyI8QZLMw
Ob8JXs7ReaA3MHnvuZeqvJqS9dsBJzbK/Lk33KAUMu+xQk5DYTYlgr70/AZNS8C+E6Y2tXK7Z2ek
SQjc5G1UujD0fCunPuyhX7RBtF3M1jmbYI+qqWT0NAknvuvhuGNAFqIMwArCZmUXZ+8ytdwbfaU8
7hH2cQevrb22CPodtpitpd98yekd+YJQDOI3+RGUlEjQ1Mu99gDCX2hkO0HBlbKwjTjHN+rMJf0C
WaOE6WTrLMOBIg085wBzotsadDoBTvtfTrKEk+A3hPJuJnGZHVpIEgbm64CF7Bzs2Mkj77LAwt8y
x+NQCftM7Z9dm9UNQqp5R6gi9RfaVdcnLI+Kgk8Vul/4aX9elH1rhnOsUX3/W0s78fpmYHRGBdxx
dFYbfuvWwjp4f2xDzUiPopuOVV4SkDkFSj/6TLug5v3yyCsZf8y9FJnK4QtFiDC+eLJTqRWWOewP
O1QZXgJyoqDLHIzmdgnlKv5zKAyxlT9iI28Gmj/M5LjDvR3a7TWtGpDCCiBLVszRHtg4bzOrv7CL
4rPNyjRmf+iukIB85fHp2rZ5PWvkIc9JmVIZdx8s25wu+rcwQ4Azyosiaw76aZ/LtoFQs8OLi6IM
Za+PWNuM2LBn/W0VfSW/EkhfSjyU2FRrEzFvCsO4GiXotMgFXNAuR4F2Q8GVMLGndDmWmluFfuIv
C+sgTu40BUI/KgxuzeEQjXxeWAdYmxleowg1pk8UmgYlYGm2TqAhpfBZaHKehDkpR37DDfz1JYBw
esTlHCA4rLckYtHNW4IKJ33eDx2bC29041sjEVjh67hjLrDgFBdyARih2BtcUPRc9ezGUH5gr1IG
QiSfkOIbkLF7Rearu429z+KjhqYnXw3dR5HljByLx/gt+LL/72Uo8tNCK6J/pWtCBDvglULpA8or
GzzNOiJe5h4a+1TfLc41jzhnJiov8wlNCcFiMRQJQ5npIe3/2rIh3mgKiRGIiedY4gMhbK3m8HD/
6kUucVPxUkod8P6KVbJt4o1rFMQCTHSneMgJ7QbAUQE3p43WZXFUkfPY0OwUg4hjFw/GoQywUoW6
suZIKz6ZLKgiKyeG99tRpFvDkFeGSsqWwT+gicnZWxQasJitt5Qyk74/Ae9NAr7Rl6cRGe0lZB5V
nCfOcEhHZpmrPg1ZUdOQxLpyktSiqz/6TGQ9V9im/CSDyix5Tb4jkPHn3HYAq5H1WyZx+Vn24aF2
kMeOg4KoXfwqCrKe6bcVJr/GvvvvZAObNBCULHV7BYbfY1p5lKlZ4lOpC9pOEDqf8UWkSi1Hflvx
hJui9inleS4ZXjLAoWxkA2R9vd0xyKLIN7TdIIfJkxtAtie3/NVY3khEnhZlZfv2KN5kk0VDZ4AX
uYx5aJLF4py0RnNgkpUX168ptVu+fDKxr3LiyMVc+kPw4cMA27BG36SFRhL8OY2kK9dBNpIons52
N+CtO3aYNuJ2Jwk5u1hDY9q7w7/FafnNsO8twXaR6CQHvBAwhh/xkDGR4Gjq6IJ4LF4zkzk7x9CF
bHpEusRSKH/yqF49tTwrmM0Yr1WekJLZat31rOMyZrmczu8GjL4BKWeNNSA+pcU8WEKDaX6YpYB+
+Av6hhHyDCm8Srblp3jwEIDNCcpkkdKTG9OJMcUXXRH2/1+q0KYsDxGw8TbEME3ZVG0kMZVE9bX3
ZgsR/NUJI0LqRGmWb8Y39GB81SNrtooeMPbNW0ohneHUf2ll0Q46DU/Gwj/n453vogtvWt4aN2nx
RopxyHT2a4xV90PTSkZ+y11osFMqdKMlQfPe6/YPO84NM+1pRtHOUjFgJXxArRmPY5NwObia4lHK
mRlPtmV8+fOmzB2j+V6t/iM5NFpdpAc1/BBXmt8drV1of9hvgzyPl74yHxJAOkMH5Xmcf49LPwF0
VKbmskCQNL6P3nMJkeqgAWIpLeHAGlKBiNu/76KhEStGT08Rc7xCvM4pihd2CDs1+8esDB/TUiLh
Q4KDkw1EVxil6oPnbUV4pWzLmHabC8JUy+7HgpXyRaK/kufl6VRr6qaHrT3VSvY21DL8SRjopcO7
1d9U1YAOVrP/JWHPwZhaDF92OB7zeuzApWg0ZCn2mi8PJJGvmIbhpBVuZJGn1Pi37ZkfDtwgyyBW
Ccsh2iWQssWJksLVaLHkmnmXWNzbfZ4y446vSEARGONy6O4NJBdEroIdQoWNX7DZKMgRMydqyU2H
Ue2aB/85Cplf2sE7FDGzA/uDDiGQLAtEg9+8APSFyTf1XyfoYz/blEFp4H6AN2LiPS6k3J0WJmBB
I0QFa4UDjNG8CL+5mw2zqClFiToietfFubkJaaHCRR3wadClEgsxHg18xIAzqH6AbU3UrC3qvmfY
sJcIDKTDqMaPtm8niYldmaSnbUUweAwwcactks2srsP3/Q6JdneS8EN/7zNwAIwoxTgCLGWaLnIn
OVNqdB8qvSOUppdv5tn7lqzr17yCkIDRfsfvESDol2P9JFsxCe5wUHb2b514mNMOo5NYHSuY91GQ
QTJKEnlZh5X8wxvqP87Ia1k0S7LH9BPzPKoRcdH8UUX4adtwPnhcXH7lIJWZwkarTv+2p+WG6N5l
IAHimvj4Pk0l8WK/8ndSmMcHlqyxYNvLG1qU6+d48SqIQxXNnt2i8GEXp72cnu280Vp563xLie2A
rFY0YCPSv4kerzppFOmJgXK+VbLOiU0IdixyyK61suc7Vz+A0scygaCYUonForRGQKxM8zAHMTlW
seOBFN0p/Orp9NIJF6zTbQmNDYR1OdXsnORdp/6sVf1NmOxiC8BOsIq13Acx/1WMD9gEVHF94kSK
5qfZNHJEPGKLWc48lT0broArowT/LQ+95nOxPUW/GX78dF3+b6HyZJoh/0ifPikCwJmygzrDJGJB
VELrgeSseB+oXcyYRaRwq9RvCrUZ13Ju+Icy5FOzNiERTOmnBTaS8N2ggkIYqM6kK7LcI0GaTxLG
3rXp/2ltpffY+pWWQNN9jM2CiO14LsmFW6sCGD/Menhbt/XCofE7LZl75HzWe4eWzDOyM45PnFD3
tTScw6agXneebJtsWK5Lxp4aN6KEbMXSd3f2I3l97YzUFhDyv6TsO7hMFMYkuueRTlRR5Lc6E2J8
nyTx0EXxun4UnuCQjYUDEXx8yyPKfj/C9EJo0iG/32X9CV/cAePE1Cg++KrgB0SHndK8mtHOGKuD
x2Lo7m+4lPCfyt5iZpjWxk/+ZfFuF/L4HSd7I//74pGEmD7uRoRoZewd6DFQVmUY6WV+5XCaNsRE
R5rUAaKfmhSU3KHNkWWabJrxr/1exvnb7YFkXzq25/y9khY/tRNhBEB59bne1dC1JCCSFPSckT5L
xnJnVceAD34WWoOw9X68zRQnS6+mvVXY6m5wQ0m+OgppmHnsO3mrgo8Hmr9nHrlIlOGXNdpdWALo
R4DrPo53RTxNd/gg+5DyrZP9eh4vBLW+g35McwozwsjxabbnzpFAQSQcxI1UCOtDC5YaYk5FT2mU
O+mnrMF0FjxfwFEv7huyBT7sdoH/SBPL+5SISMzpVOe9jdgiotfgXQx4roDRIQRLEWhgyt/v4QbP
TdMZQy6yEjVg6o4wt8cNHl5dfSVyMq2WGkW55a2yWkjLskg3KWtoKyZ5fwotytNVF9w2mnDZT/hX
wG2YaRABs+VB29L3ERpyWZ434dQ5AVV7RJBHqLdF0CS6jZjHMuPIrxDsQ3D3rwVrqYhLOof2yxhi
GAaUmNDoau/NgsjmnB3yTByKKKFv38pGY7J74Q/8cV5nLcUQsTs/5aDFbVDVspuzqeUzISWK6Nzs
XeeLtUu4X1IJcWH4h4YWfKfu8Goce2mtoKtASXcgxBuwZLDZn8Ml08dp4Qh6shFLLE/+9uGfBM7u
uv7G3JtEk67Itu88s5LjE/Moz4fUpuAgkaiA6nA5Ov3bK6WRnCYysFNHHofZFtN69BaWgo8H4EYt
0vxb+lADHCEPjHApq/N6n50b0M/60jFMTLYxkKpU8Xa1xnCyyc6O8vHb/q0/hZmcCGX1JgNM4pYu
rt9+kiKRKqj+bOrAflH74fgdmFcO/41hxbx+K9IAdZmbpBfIdw9mJ1rOm854x8leuP0sKye2gzWB
zwOB9n/mf2SXjoraoegocZrHHGYn1MYaaoSXbfMg+TDTsuYGL9lhHbGhgUZC0wY/ZqWN7mwStNfr
WA1pOm/KB+uhDHRqbElGy1K1vyEzyLqQSDJKcCwY4QjtKk5+fJoAmR1vQ6f6k5ArHMvBh2VmqKTu
5sCeVSrxH+o33ceycygj8t8XzH/DqgiLIZacb9/L3hpARc29dXUU20Urd/gBArcgmzxW2WxVBVzu
c+2LBN6CEX5lM3qHCQK5kRuLo99mPc0D6Vxu24agsXFjj6Uh1hLa68OkE3z8f+2lX+Q++XG/6YAx
5Xh0fm2YdRpo97t6PWH5m4oc1rKQ9+JZuwSoNhmSzrv4w309AZb7vLVazD4h7+JHil5N7Tyo2J/z
Yy69rp6jPOD8vsLxAQUMXK1vVkTypZ8SXUoBTUrEzNFpdOiVnx+7U31EIEXNDqF4KyIj1pNZAWx+
C8yn97fD89YpTz09VAtnbt+UFVuxO0Cljl8GHv1Ax1ME5GSdV10CWfQFrcHnkf8ZCr7rGG97djdy
Dzq3fhCG1uQ5/4ck9vxnO+mlKvX9YiRg1F9NkzeI72gECKdQJ69z98G6x1UqrTBKHxFKAtSjS15K
Fc6hvmG94cK3EuKLLQxZ6EQL+7GVel1djTSq5Ti8FOPZ/slgU63K7KC9Hm9adTswtD9a0MbOQ8aM
di/rb9hglPOCabwxDPjQZhaGEyyWqFI3wSD90iInVE3Pt20L1KGPcFex1OaTqYiherfTapagYhOs
BKiszW5XowrciIMiWE1ADED0iF7y0RUBajBb9/zeg+a/nG9RoyfxTgGsK/0LgWKl9TxRThUD/ktQ
v1d1GbzqdK67jF6vi+copC+bazsiTCH2ViedGZiio1UcY11fBq7WkFca3Y8n1q0xEgb6taNu4RPm
rP6bHEyAPAuFEwEzQVRsjZFns9CFWHbvmOquWYuvdVokkMXE7k+kswlP4hm9YoPbyN+KbENKeLkO
d/y280XlzqozxMcz1wLTRv+4/2xOmzkHd0sXXB1RvNhe+0E6NuxpfbjiAW10EYPtJp6lc7jriipC
uJMIH3bmpSvY9KgjbEDWBQZPGa0IJKsKF8BtRtG4M88KqNPIEenppT78OY81RX7Hxh01o/GC8Ys5
zoy0GtNpeoi5cijhxN2AQX/o14Sny3sexIqHfcRWoZMcRvsFjRIbeeate35ShC6N5OQ2UjUZgqUf
TJbEf/GYq7e4fX/MfDJmj22ncCulbb+YQtWyjJb9CxqkBxP2vIEe+AppX8ZnWVk+BvYDUbXG96EH
bPkX1qsXwc09jYveERXtfDRKfMKW6AxnVRHWxskLB+pfuJLk7BI9qLGiqsMbo3jLsHQB9G9kMnlA
Efi49D0AHsGwFaxNI+ELEHdMJ65WTi1UQ4hSIAVHAn9UGmdjCavRduoCTpnwYAcmtZ02cXSR6Yeu
FHmkygra3YTrdPt8/WtrhfHps33JYaPTid9veOCAiq/krGruUpdUXgX8S+gf5AAPkhv8INvL2stv
AgFpcMuOe2CF+xMpF2t+quA7qwUhI4Tf/WyHWIv3LBg/wweJ7pDW53v2ZvgMCtjicm3WRjPFIwuo
KylF4ZZ4Zm6sBrFCMIE/L9wj5Jj7u74c0QYHWDLHKgdy07z5NKrpc/PJmDf6HkW5Tvw+zVLXxYF/
8N41Igr9jN75o2MDUvkqyIchxCUrCvKiWM00jpESpugiOhnwnKewbCGB6SHQbRBSEAAqXctPmILZ
MlxNEk1Jgab5KupQEU9Guepm5Fxy9xZUT/z6c1N8mtDTApXuvaabQ5Yz5CZ5M1sNi/Lb+zwRou0W
oafOd+Q8Y6DwUVz+U/gBopmE+HCyC39Fjtn9KMcRtRxfSmKVJIinWe0P30Yn4fZvkmXaYfIu8Jf3
GY1wps+1UyBohvMVeFrPNmWke41GLQW50iei2QlFzs2MLf6Y+g9KPUXEOUSusUa1GoGassG1RfoP
gEM9fE/a9qQjV1rK52qTfaebLyvIx/+WHzUQxbytb16XfUeTignJXPEBTnsdr3QGBI6SNpJvgCG7
DOaWMwqHaYm8rHB/9nAvkx01o/+BnxuZIkpErzlYVEZZZZH19qMaBvIoCHuTRmgpWoTWof64f7Lx
anbNVbopryk9InHzCNWMEy0/UuXoQvXiMXUD2zcLeqr+BHrncJ9ixY1Se24IT7jtmadng+dHbpZF
2jE3EcI2JObe7Y1ZKvKXzGBZuSsIsnvrrx4UfmvBBPgpuQVh5iM9MszLEtxiH3WU6Kt12grExrV3
CY2G2+hgFP6+qW5k32SjQ+VtXARajZxBBonevOo4o4JqvoKbwBLCbAOqCUlzHhLDREbZeqRmN2Uy
WvTvUjGzV+ta15RKLLbUO/vnGByyR6+/Iu7TDpByxcKsic0HwV/XUTVcynGaLqZUjvVCJVm3Fu7E
uz50pWZ8ScqUcf4N5055LMe/34h8F7EBA1dwrHmFLhnWbAnKMQrd+/Vkk/FOtcTbo4mUrE1SLHcc
RsVReEYVunNEHF+OE8cWG/nyP69InCESWTwiMkzGqgHs58IfhUUiTqvV547Z8d4aXf8CDQBY6tMU
4njcIEIoZIQVPEyAqKw6c9aOXbcWJIFemTyNjvzyW4V8bxLGi/bC6q/ItMHla16qd9jO3JEMgS+k
R/gJ8i2MpvK3x20X/UplTYKzPHhXS4p9MgRn88E23OYZNBnCQLqANVr3F7FYjFrPIw2kWeN/Tb2P
8oVAY2Ta/QsBqNo2eMRPpNBRfk97IwENGUBJKfDwKLOkQxvEexYprKB9FCQMjTIEMBEuTi3Lw/aN
bMGxzYGdNANd3Ec25os1wNQcLbtKiC+UmDwymr0AHSo6aTz0dvIWFJT4TkFqBv/ZmcYPbs6bciwt
Sjpq+py0FbeAm/jCGhY4CDdzXwVn/3BllVjdFfpXwY9hhi8avHyuJOLOvB5bTmlK46CHssnCKZPU
J3QhQ6J1fkPeOZ+ck00b6cJ8XiJ+dIIVLZTxxp66SdadL0Xxb0bcbcJaUwtrT9M73dDW7keHM7sp
XJp3u51cqUW6tgbVMxwJ7mbLlGBD90Ijea1cj77PrxS8HtxtF5Dj8yEDrerZleltRYacloOeoDPM
XjLwD8gNeYvoJzEZywlNcVPLL8OXo9+9VTBjwdwuGQ9ldDYsNpVYMsd4lXnCcFOQbv8F1ZRrDQuc
QPDqNM0R6R38uiStsa8Uli7C32cElACRCwWasyXFto7BLmBrnCKhMctLlj1eZwpyweu7n65BhVva
I5Bo4dqJYFQCdERiXtDV2/ZipRWPNiU3uPwsDS3l4wBYqd1itLEBeka0qOjKfXDGu0zka8upx16k
j5Nik3XOnH9NPq1xMGbULPBSfJAp13PMC2Pq2w7VIAGEpOwY+g0hdSZn560RZlJXrmfWn4rjfggl
rpX7oFmMkICPASD8J1kXKY5+xKUAfst2oEvVTEgbbKNSSkQ4w7TPBOB6NNUgfZAo12iBhptqzESg
SQ272r3TnMVcRwEmdSRws1L5BXOTU4oWNMiIJwtO5E/NRm2cIDivB3dEqbondsMVKSPZd6pr2M66
cL7Ty3NDPwBG4FEW1lqiw5u6xceQsB4vr9LfzW4pA5Cuyqw8AYrHawCvcKTPFDf7ERGO5zbvDcLC
RZwgh2DVN6Brmtasj8VR9xHcy4WRp5GEU+BGsiFLNV7AAjfbl5o689dP0PT6hZLNiD8c6yvWZa2S
KKVyku2F2jD3XoVqU3DtVAoMBEZZigPuNa+D8wz725NEL3I8c9rEdM31bxbkaQU0vfqYcTNXiXyv
sxZH5LaQKVOQzGDpluH9JifvCFfToOQbOaCP0+z6rMmXONf62qceTLbpRfT0bs1Q+70WR8N8XsC7
+SxutsXz4al4l8nCslgjPUsGWpIWZQ6/M0phT196S7OqCM/UV43H+rjHUxQDDZet25CNmLYDr8yY
uUaUHSrMMLHKjH25OsaLUMMx0ohxymPITOVYnSHgAcBYhe9bYzB9bujbheV1se60tt+D80bl4gyw
xuzo9OlllzY2dDR366OAwUbKI2eQlNM8IIzHm0QdkDVh9HlCI5uhFyKmLbFxqSuniPJdibNgNkxc
8AdS6KM3U1u34j1dCYm7oZDmTrQpfXnSkUBh/DC9JopTDu/ZHB8X8/1M1iTPinsICFpp4hkjGK9k
ktZmNnOE+padydSpbbkOSnwr28QveF/k2s0cAIhIOGEKYJhuCW2Snv7FnSDjgopep60/8TAobDAY
OwEgInDgoeeh5nhLFyO5U0LT07AcZRuJlUNlJnHald7/K1gfjFuARw2zy7TJkUznJ/vWZKYdvPkB
zRZQ8MCmuij2oygtDHt9KEhdeC3C4M4pVtSPhnJv+00unW4WoSqCWHG8pj9PM4LSyLGs+FJZdh4l
gPCPqtaRSVYXVAKKHxf42dWinN8byati78TCY5N7A9yXEfLWx/9N/v8xinuw0h3LF2He7hfwRBXc
hyLJOs1v6k5GskduIEtduzEA0eAuG55QJbLnV/uwORbjlduD1eDIgzudCCKLqLcm5OSM8qwidwME
4kMg4dOKqqWBPOWX5xaA5laeT5yI+KhSWlNhT6A4PPr9v4RFfni2nuMXfhgzcoLb2eJaHbiy/4tL
fJGoVykP1v+zwpSaqqz15RxPZh/sO1VLNqLeRPTNo6K6yCoKms12zHTUweY++Xv+OHJ1eoIPRzTp
V5Xzv6THA3BdIrv0DNKxBQmTXmjNmNCxe8Acga23mQC7PTrx+79dYIegsbDdU/unaCF/6nQ1aEV4
O8S77epAHSEWVKHgiXpG9Z+v//D5Q/ZSrYUKLhVHWajzfuXkkUz/6bvQMsRFL92wn5YZBHkW0J+a
bk8qDAwaBMIK0GjwWlaVhxHLzjuWBcfPJG68YowH7syBTMQ3eEIAjSZGAYJ51xaBuEJzTf1e1g3a
soZFH/2ZIcVBU5q5QN03mJX+2fbdyp6rA3W/hAE8K61UYRyElWKlJ4jioBDhjaq2144iHFduib0H
fqpE8/cXTPpHJspbLlq5JT3Dq9M9HYFyFenevlTSPT1QEauQpTpHc08DMQDOcR6RwCBD+Mg7EWg6
uahpnUcnwkKpvx4F8tqdT2rOXqGNh5e/H3AMGLNDYhexPyEqGCCUGEbvqg9d1AbdJZWntB7twgHu
HS73ZJnRtE63ky7jnkO9fRKZGmIKqKII5oBieSte6MI2Zjh1ZJte6Nl070J5KPBDXw+NcI4MiNbP
nqZJh1ZqOYs0eqh/UTAeOYWBtzFVKmh5DWpwKZqVQ3BcInUPZlRJuDyVL8FJdtS5SFPWTyFYH4Pn
bRm5zr95Pef48FWOs0nsTNZcp1fTFlgGBP+dJU9GdtzujiCdrPGZRsqdSthA28VxatB1NJNZX0KG
1/q+3kqL+7/wabf7V0aU3KQCWR1HQwj+J9BiOfAc7GDmej2w664wo5iJBYQheGt/G/gSaHmk1bTn
sCuszjohaZb7Yh0ykmBvesX+PUUW2gvYT1M5KKdth8ZlGVV+OowU2sk5bs8SBEf/mriDKKKDO7Gz
z6VDrv9sTe4yD9QZoJnuYwGWCmH9d5wXy/nWZ6vkCXgbxyli+1dBioKlEt/I4zdIi/uMWUI2iX/C
yK7VPp7sjTsq7hh6rgWVDmfgKDfqR4+UZZyPrC875W6VQzgntPXNupk9RbxIEvKERixqtiGciYd0
1lcDsGTKktECYoS8JXa2taw1U+wK25ldqEFXeWAdQe2d7wQw72TfVMSPEwNA0Mnvt9udcZ+nvccr
6RR3ycMw4DtrJJrxgB97abewHrv1twjA22kZ8sr82FNcnHpwNb+SqeTkU9SVB2NXXt+ZmNmLR00b
VGtZVapV0ePbh3pgfDigG3/SmbdnBBko5QXKDPbDZF/5bZ3Kg6kUTd3RJ5tAF80kW/nETFLS9cX6
n6mqFbtaHl6+QtCS1CLroirjDbch4Ba1+PUOhq14ocuucA4Nxy+q6D5vZOFxAKVrdMhPuaR29dE/
erif1VKZ7k3nu2zMJ+zJzy3kryx6hBNt6LqhacWY97M8nRiE62o+BQLJhlaXJMcwSskthfzydD+Y
N9E285CpY9aD81EepaUc7mLarSbbGXYjEGzNT0OqcT+TQ0lMzuhMEgNuHzFOIMH2cde8ro31RcxS
7peHnILhUKEEkydlA635W7ifrvNc5qFQ9i/LvUIjBtrNTeOIkdc479FLERa8u0aBY3cVeCSPngZv
i/e7ijwH6fmcfueGsdOS0p+s02Lt7cL/8YPn7U7oD/KTMroxw68YwPVrqQFihy7Y3Z3OvtmuOMf9
8SrlzzLzepSxq94vM0DMIOvi9ZFM644MQxLpz1pbfFHhjBOYvghISeJ5fiDdne5AD+xNTkmW2cjq
YgchM4OQy/UkJMGb6bQP9WqJt4d8w09sV7wzy5j/hMtVgiXJlsLTUkk0BxAA6ysr4QWQUy9sB/3L
3kwGNgtTxl33wKhHFJQzC2w+bFDlji8xRn+3dQIATkH8xn5BQLaGDsuD79b2ITLgBpdH0jGhTSjJ
dryIY1OyX9S7YB4LOeTc5RCoEqj+B0nUj0GqGE4eCVQCLys9aBr4KmwvzGmoYvzcvEeMe0n85zuR
Bn5SIk0h8wbHWwZ3UeZYb5CrPTk+spyEk+MUC4Y82/2D2nE/y9ysUVOrhN+z7eFkfMS3xu8Xz+up
jjlo4yyKjJaaeGiMh0JVkY3fsIXgozAPgg3N9/yADzQKtByMqUmfwNKFqPp6aCCMkKnQOCPkenc+
7NXpQzRZd7sjDSdDVCRhfi6eVYdx8LWaQzGLBptlw/oVE5/DoL1JRhktD080zmXZx7qTofGT21O1
d7J+tUta1W6hxfQDQK1aazEdfmrTeReBGxhHCXympO8qShkDT1Lns3lFLPDk7CdYsAKlL3zRj0SG
RPKEEhkjjuuYByC/ErL4dUBPVNIrmymLaaYF3xnEa+NjhDBfeVraC8UQrcrsflzaElyKJ/16oe4q
en+oAQuK6zNLMjaxmWPMQUmJWhy7lv/hIFb683UJTM5o4gEH/jiphaM8QaUChsZYHHgciUBSt0JV
cyqe7vJKKRioTmNh7dK+U7CaY42/JeQ5EJVJCUctivFr7CTk9r3mWTXhsn57TYhvppMdLlL+lwi+
wYSZZwM9iDv4OJPNR7YziAanPotswEnUs3yEfNoMyDMzx3rH/4usmaF5r49vQzxiD52203YhgS5o
l3AoFAvbd8LPACWs03ou66ugAsWBVWe+d2PSfFJ4cLfxicUGbFZvz7skCcSj+OZZZwY7gWMey9KQ
8+8H+9cwikgGvnTVemErSAef2z7i2+XAhx5o+JpuFfzefDXKvhdJf4oApOkG1VoMgIIR12cQdY7g
weQLBZZNJI+bqaBPHs/S2n8nb5lrJQGWY7GZ8q59dkxK0ArHEcAyS/BRh707eKIlO5Am8Gg+boop
JYnLYbu3oPZhelWK5FiCTp6WWnzRjXFtpji821mBn+nhKT+2bYF3fbDaqwVK2TuQxsDhlV06n9yi
qA9QQsKjrbmviMrmhMBck4bMnERN4gbNipSZDTO60V4WYdPVGzywKaZ6iRDmbDYo/Kt+qqZs9Rv3
X7HYs6orD+wMiZLACQEOKQW6GxO0LEM9Hc5HQC4yaBxOk7gkciEDbJOQGJBHhhaCQRSzmTyK/uym
i+/aQsI2mW6MvhhGVkdUZUd9v4SP50Ca2vK4yZ9FrFQjQYn6OcYubi8HKCHhBrwU5sixMPHpxOgS
1zvg95D26B8z1BFcYEHboB3dzGPGyvMBGtJF+QDqAgfxZR3MVHHF+0NkTaFvNgEa6e3Rs6S9s4vv
jdCRMRwxuqtn0wpO6rSs3043BP4fVb2Ll5BYv7TnkP7NwCRH646YQ/mS2Dv8O3FMFjN2Ahtxq+x2
qo86ZjNk+Bxua/ds3StpQcRoJ2ynripJM+KVHJxi9npiuAWr9cjd7X668TD8cEN+Qca3aUhx7arr
//Ntv34xvyOhiRZsOyTFNxuAvQoIEHKpj4wFv54B8yUFZvtijpL7qWxw1cP+86p5XyNk91pshyFO
riproZUXA+jn722F+SBc2Fmf4cCwkWS/gWb1FBLISNB1zuOKYvpARshFRvAuMBKUzmALVXTUjSTX
YRCtIRlll93DmrER8csP/j0+aeNsYQluI8t0lVM3Sr3pm0ypzbuGfE9SOBQRQoFugK36vtbbCnH7
eIWYHbTHKp26A6ipZvxTTqru/PqthzzC3a8P3Wf0gYzBoDlIWlfioZ7kBpjUAEkFFyEV/l+9IXxR
Vje05e7HdS6ROyybuYMeLRGsJl2uW4Cg49FHJr/qTBqqz+oZB2qbctMa3fsLtuyElVtWP/GoiWys
s0zk4G0b00J/nmBf3zI6vG+JXcSi/t+e5znE4y4fkr1d0vZvw8nBZJtBXO7OJHiP1ZJRd4eFpf/r
Axf65NxU6FgKfZ0HD/PcJ8HlmlykenX0HIOgdkWgyStDuMadQw8zE3kWHA4sZPNRLg/EGzeyjCEC
8H8L3VXOkS2E9lRugTazye2JOaEcnsBT5/r4Hm3CmBuyeNMNx0K/0yX/NsvurFlXCa+mspJTQzM9
cHfNQB9d/fEsoixIvlkgFEkd91DKq6x+XNmKJvCYqpIlHnIpkvzjKqhwK35n/ZQO3EfERvDHrMeT
JNnJZ22a1lvB7ujdghV+4Fj+IAaNKHlfCQc8l2rH9GMSsMJ6WbEHtLKxEODsfc5Grn8KsxSFD90S
zgfxEl5XdC/R9jLG+4xmGoHQYbCM4wwIOqV4cVKd4mQRotWt9XD+936QMJvgokZuqe9gmhQg2Ck8
1JdDMZNC64Ukws3bLZ5/9ahnQkyn834QaZuPyVQZONFRGvTTZl/8CRG0dvpSg4ou+ovMdDhCj4Dm
sh8aHWvNWI9Mw/g1HBQtBuR5oBgmkQEyFysUOf1jGWPj3rY2C5MRIL+NC/bvW4Y48dCrtxaSkQxK
CCA2wiBs35z9mOYKfu5A/VtSDsKynNUh2/7f2VdGzKZii72oh/rV02X9RSkkeTeCkRa10icgQtZV
Tx/jqpFPq4hz9MrWYwzGZkd1FQDFtc/SQ4FKefL6dVqPT/3TsSZHlXsqm4TA8uxO1E6Ecg4i8T/x
nAI1+bW5o31Uq0BezN8y6rYHSNHjGt5PugbnXy60/z7ZJ/L4QUSfhGE5K2v0q0v6aPI9FLrBl3Sh
BTDGuMCymCEqyL9krqKmw9kFotv0jufJHg0C9BO4v6sxkGsMHJDdLgisGS9V3K+xN/+UCSK6CqUa
mei1+Lo3F2+mkUi+KYrsGyQyrb3xBhO62v7K7o7isPRES2I4Spl6ZZyhCzsBTqdx/vIv/CcyYIUD
8c1p1mBLGXETikJYRB3vnyGcGBK1/RArINiDsVMdiYbO8p9jU3qtupZRz5i50usfhbgvTAxXNL0J
76LF5vKt0Vmb+F0lGm87t5R6/M+AxRSbzSNaVTA50qsq2f2xQ7NtyOEfBEwOTxJjUGsSaAKciK9W
NbY2UENpuuBbm6sYjL55uMkJcE8Q5O5kzuiHyTYNpGuEY/tCAYljRqqHbT9fh+nnPpoinnKqOAf2
Mpm9JkndUITPRBKb+RVKyEzxJQ78/807z6UtD1SqfyQKLWvDh4I1GILz8DYz98uVR6CLA4Ex5Oja
AE3+zxra0H627x0KqBalJCW4BcmNWN8E6HWwN2dZAE8SbF227iUS7AEmJ7Qnc/97gzwNsJ+N35Mc
jeR0xiDjIqVGCTpjVJ/i9HY3BpOvk8cxJgXfhWufXeYf9AlxS4AsBZA0AwahHccIzZRqr56jhABC
SKW1Z/MT4wvCKyjl2u4REDNvbsTvtKgDDqBXnvXApKzmiuFF/aE2gpv7qiYbPolZFEvB0aLlAjfD
Y9eWw5ttiHGxu5KzHK7dbw+kwBfyhH/3W2zxTu8i6p0wcu1/Zsnf+J1Y9iJNteUsSgYKnuLtQ1U5
S99vh+NjhdK9DEO9fi7wCSZIDoDX3lV4gi8l3xeVJd3VIWp1lLSi56QlN5HMjRbAo4CCWZssb2Ar
+9rEV1bhWrYm/xh9z1RYCzAvVt1ZJJfvdTzATbmK5i2ZYSoEe8tnXLMG0QBIfx+85f5l0iTTEiy7
q39n7xkQuWDrQpVzXqrYVd8XTtxZRdQDFM3ltct6cFNQAi6dFVS1jv/uuyrEYb3XEhcY/FUGmcZq
A5Zf3XPeyEtEMlaBLVP4ytbWNWiOchFBjmGmtwwve5rDnwXrpfmihEY35CQPCSZ+JcfJY7hwI7YH
m/HsPxpFJU4sz9J7CIjti4Fh8+SV3wdZaLyPv1mfUdiUbqeDDveiPnXr1qoLABGfnAodZse0HboG
eKx3lArZqVYBRBQAwKvTo5M/iO7hsOzHJIjCW8ub4gPz/dnID6gdZQP1JdqcVbqSXXOqQT6+GYAl
U5fyNhGplK3kcx5Lbh3jdpPd7zyO1AUTQ12O6EDAPV+b7GOMeH3wyCXWWlpU8BZ7rZz5m2hcH/BL
tm/iKUi+GOPziWbZs5WTJqsghgk9DZX5K0O0kuOkmMxFyFdajl/FP3fs4TPkD6zYCNkadaU0R6W4
DPxxZrmgUUXnwE2wXBE4GKzBJKCmfC72YfbDKXqypsT5n42bJd0kOxLYiqPsARsX/bnAmxc1n5aC
VDZHkDlaKQUvwzAj7WXrx/khfTWNrclycUKpB8jAPXnmJF2H1l+DUQBBGW1JIif4+cZ41RxUWzfN
bmFJEEAZgCZiUrjUoirEqkR04+oeYD5XMi4hb0yp6WqtnnUKMucUTiZQAPvyI4SO8KrDAEWMXEwk
ddVh7k10skhS/noN302NepTFFpsRQNP3pacPUh/vj5XXDZLf+r/p3NQq8/FixIPOtVhFPV2qb08p
X8cMwrUuyGepCbdFyVA/dQdfKs71795r55Q0dw/pteq5BGs4oRlHrwqRYxSNt0onT87rK1LGNLIi
p1DcKNrWOWJPweB7H1vJlhhxtHkfsU0ENdt9//1dYU7hAeL5WZxMsIn60/WhRmceEbnUpVys7N5+
THrzWM/05+9VAqN68LXGYv+ISdbtBYBhmPjZiXh4XYBHop745Q1i33DK69UuaVbFeLWagh9Q+GTh
5+6IFrgvAcnqqWjvHPBdzNXhQW7QQwxd7IM1+bdxP32WWbqHUdzQx/mmz+ORYuRXfmjeRmfWfVeQ
WHSxzIob5lRfyyHdwqlxJQeuHM1+ByRdNoWX06hnLer4Lszn6YdhWrWg9RgbqeCduGNRSk25PQRd
VKbfI2Mngx164AHUwUx8qoq05SDGnYTGLGRfamc2rhxGJzwveErsbDXPIXfmMdxR21TCh4u+2jbu
6NAKeDXQQVrG5nqFm/XcaYCtBWYN2RXagx8tKXIwb419m18pZFns+cc5lTbNvBkyl7kWtGcVfRMi
O/bEisyzPfT8mDlmT9z5jxDILl1b2xVjNR4veamZxH3BrhzPXo1KOd0atYg0OpuZSJmWUlIWuSZE
2W7YBu07zisf3HjKNMGmaQq43ufqOwr65qpKvbuGY9w9ADPw9FEz6arrHZQvEsQ6I8sNT+/rFXVn
nOnZNpKTc2F+S4imuRI0KlxFuhrNr8hU3Z3Nr8D5WSjdZagFWTwxlxNRdnmE0Lg8juj9fo3Os6bD
3hpWiLTsH94XjqOdQ6jXMpHHDroWPZQ0+MzyHFhuHLsDGScNTM6Y0z/re8hQWnnAMS5m+Ildyv65
AV6kAbWtTTSKAWczb545bmIjd36icvcbPRrv01G+lhM2purkZwXTZtaEARQIiNsQwEidrcu2fhYx
E28pm51ybMVS8YbaaCs0H3GHPWeFBaFubKBo9H3/JVUCdD6OToOg3pGKgL0Vsq252ipv7Nj5nxbF
Ea/Uxdse8fh5CNvND3WX50/KxQBBrC5A+XybamZ1z6Mx13nWUE2oY/WeMaluaG+XYMjHt6jzNoby
WrwaqBe6/AEueHbEscTgakV77ODuCaMMPRP5ASFgXJ6jlAAj6Z+aksbiO8yb4LhB3trnTM0779oK
XgLN595NQHrkfabvx8w7kpCNeBrdvctov3dH2O/mYAM5VENdrs4sEYqbuzdNn/R9UcyPj/9bTg8Q
aTmMfeEI2p2inZDBNkwCCYRNJlnjnsBtmTnQ1hPxMoTC9rGSNA0GHA9fk/4l64oIsEarT0FP/jzm
zpvsZMCoIx9rTJyzi20O6s13Xu5YwV/4j8iRXoFN8sYdao33lzdfwxcX/tq7G04KRyt3YVQXIiqY
5+1H1kFF+rtT31PblGkhB/YzXO/WIQClutURWyfZJVJbH+/arxKfxX5tYD/9/VHGPYk4QzDbVeHQ
/uUy1MJ6YBxoakEMLPA2ktGICBV0jpi+KbHiCKlky4+olcGpReTwlvDLLQMIYGtLF4Eik4lSRAk1
zHn6jyrfBX03i3PNwWS/RsFd7JlgGEpDilPFjMpT1HSm+MAqSNHsraTk70fGpRh6SCd1LcWkC5cg
crNVMR7Qyo6/rcpbnExy3ZBQqQaJJQ7DCKe25Mt1mdPb+3Eya3vODDpRPbJSMV9tnMc1PXn2cdVR
D2PPLfuVzVRROxJlDzc1cy8jRMy7WmpgE0uriSCGWElVxKlpVGxbINJP9UB9hcHRpi0AT5cd8XLb
oLSG/9Igs5DeaOiQ8lwvPJbw+HoM6fqJWILJ4ave189srfUR6vZJQM8/MZtrsAuwQ2AejaFNLPvZ
capNrTemkvp0glPHxxp7jrOpyWin0qSn9k0unk4WHAbVna4Vw5vCpttPdfZbH+8cZT2A6eiQdPjs
Xkv3U52GGCaVu5AqiOO7Hj8tkXKjZG4FdKPIB5AAbQsBaGAQLWLLR4O9xW2plWCq3BNOLvvgj/hV
kYfOhghN8QPumme0M4BgQvwgz0aqWVJlIlAazpcq/X+3Y4MNUU6aAEPejUyLXX6HrjofyR3xRTHn
9t6M7G+swQPzA2xyAe5TGBRRjnaqlPRhkWHqAYtELJjly2YMRRE8S4LEU4thBllSdNpdASNqdgUe
GuAbIV0aQ0r5LBKzjmVLdIVLBcPMbhUh6YmOubNrE+bbPJIL4wE09JQVvVvmPpiRCoshmSfb9q7W
9mhi2oYmNQNotCnt5Qnf1iREVMeXNW/jCFtVSzcocMiUh6CN0J71TASMjGdoSrZK9DratSrmY/LF
IeIzeUxncXvkgxcEGsmkHJr/pIYHk6dYUYo37UGS8X7zW81e526YV84zZpMr2yQjlMuGJoOPW36H
W8iq53QGOyucyvYfoHd6xpIAIqP1NtLhS+NrYCfyH+gOiYAhq4dWQ4bwz/zF/q/tPddm8yHXk0xn
00K6LXAGZfug/2dZJElGoYkkntPTvfCyiObfhkPxLp4nnk1PlG66PmGtLs01g54xz6X7X5ULGpKu
lF3q9Dbu+YoXnkvJzrmeM8xuQbH3gHqdLkNQeqr5wTnqvC4sJJ+bJWGZU7UMuESqYsUPsaiVRNtx
k7EQweq64NCWyKDY/25LU+Z3CiT8zwrOFwpxvpXJU13O6aEDCIJn1wrKUbSpNvYXgJujK9Pl4knE
TEXpRK3EEjrkxG5sE1GJxRFMtSdxL/2ZUrHg8P7Y//zq9C34WOuN9sDHIncIBafZrF+Xr5+SFpDt
dGB74+rJtANar6GVbRLYrCS5rfniTPHZtjI8FGkokiiho2tu/Zy9XIsUPcK7UzMwCQxJ5CLYWd1C
O0MH+JFjjLkMoPu6wCApMbHy65uUVeDxp1v8X4YfrjRjYbXiRI1dLJK+ZYdsuXS2c9E+qFq7uZhe
dhKmaIUS9JMKgzKROfGUp1AQjBZLmmfiCJF3/4ZsUe8I4pRaXnLutI6yVx5B2E0wLnZZUvCFz8cg
Pj7IxbDlZhTac/gkGFL9Y4zakhwsGMNXYswPa3Wio/tJu42i66Y43+VJjKqAiLQauO8vSgP+5bV5
QF2tcg4vA/L1bg2ylJYug2/lkabSg65yind11/FHw30jy438IBgAGS9lSooLYYUhaDh6fg0Vq3tR
+k8IjcmO+CXyQASUZ4dm18Lt494/CayE+1edzfIgz3CJGbQfTD8iqSVOBLULe0UKseoW9GMtgD88
MKNVL1ahQUbnMoy3vADKzJHLwwvQotPQjqN1umPv0JWBgBQVhp1UBr8iV7ZjCXmrAWQY/9q2JYUd
ooGhAS1/pVKJ/qP/a4UDnISnplCExduSnpMztLsqGoLzfi5yI/mXQE1/BODOK+jCvQqHIVnqshxG
j2Mcr3YMgBkCtH7re8zvDV5v3L2W/6mCiYaLpjgTp8dw8C9KutaOUQleWsjlm3r1e9lvmh2L9v/J
78O/7MhkvO1wqMHqm6nWO//NmmU5iIDb2ImPqITm7xSbo4PIyJbs6SEfPZVZzNqvzJQsFyURsnZI
KjWOpvA4Chrw8vx9AFWqGI5yEpUlTZT1HIBZ+fnTlO67pqECHgfcUfntSr018BQ/4CqqfLLq0vds
lbkPCYWhTeh2BGhwYFyqcqdPGPiSN+RT+mqShXCgpobng3+91Ax3JBezT/DBU6QvMmvG0OQ2oISn
PzOakGcRsYC8G5LWE8sLld9nKDDyfLG8MA7SsU7hQQ2zk7Gr+58ADcS53AdCe+APszi32tl9ywm8
3EtVqSMBLFNfj7BEB25sObF2juFfTAvy/xnY9EtUFODXKnhRM39f3ptQm8T3bmkkypnHeXJSse3A
Q/LxDCOj2ms86/H73SJpEXppNL9jhEVpFi3WJN+1oglG8AntdS8svDtE2XoOxUyPLwi/GsQbeoqB
OTQQeJxhwK+inZDHJgcyKOAcXA3VGxL6XQ6lXxuG4KXjh5dmtCjdDD9hnIGNPWqFgJvV98mDLudw
HnsL01abEvxxObDTIgfnEf6zOilTBjfbJXNeJu7xdsKEIOoZKTW7aaJ1wG+uzEAq8b9+ufknd5KA
35W+ricuQ5aNxCNK8S+ZEQ9aKFUOByF9mbz8dsbGkp5nI6YIPclxKiCUktIUObwXsMyyJwgb7seU
Hj+Epi/y8EKdHV88ZEW4hMB9riemNQcD/XxkZa6UkLFPYm9kNpciQn4o42aUAXFaxHYz2pUz+kI1
zBmTY0B4U+7qRYw1NxCcz3QdTIf+sE+CQgo+6buSi7J2Rby8/XQOVuOQ3WYBlkY00rj1mkrkzq1V
ppm5hvexRJ0y2opbyTR1bPyYAUYBmnpk5+1nAgV5Sd6tOQ93UtpGed+iLox+1y9Ctax3CnhzGMW+
qBflkoeKOxjE2wWRhsP9V0E2LqUdPVewntammVSS5+40KGkPfj90di4MfgZeBVYrtCqJaf9W6EBP
pncRvoGlM55UMIXIcsrdwq57mqB4VTxFb7ZWkwZykT+nma557nfcp7EnM/+he3JkQCVW5UODFblT
pnTNnI5ud7Fpmg2CnWYribQIQQJLXCn/+2DjLnY5gJ/O5iJ5vcuYfB3O4ASTu5+RCZtwgpqvCxav
rC+3Z/EjpZEQoBrTZmEyCxEqZz1wupmf8EGcyJPkntUpTVTXnKBkanWMN4427cb+63EL7EMMynna
XM6Dq7UgvlXcNtl5C8w1HjICas49WdrDU/Fd0hJff0wv6Lg/kgebBEk4cpbzSiVbdi2WuqXWMeB/
0sTFzkP2Oj90BF/fR3ccey8O4/yirP2iPk6pUm/PZ8lh5NhE2b1p2f2vkI00FiDJ8IujuCoEbCGO
vZ2zkycdOIuphUdGcMvz9/K2ioshNCpyF/NlwXhttUlO0XQEt+Dp4aoFQWF06zYumm2yikgOF3ik
OwGRrfqhyPq2Dj8w7EFKv4p/iC3NPBKGJe47v4R1RWzeId6MIvRM6hVuYbMowXNzC8SiJCbFd0Gf
/MExhy7we5IjHSwrHRhX7CiHkb+fkgQogs0PdSC1RDFlNjU3TEzE3j9L3J9K8RrWd4vWhKqSFNuy
0ulnxM9uc3oO+Wds19KWJhiLM/4JWiesczxQhJYkduad2P4vW5fcO43fJcoT4gts9xugVd5O4K9W
hAXRUtY+a+RBNe/2b6k5nasdFIDdtW5YxCdujI3EEQ11/kLErK3slYzQRqYrMqRjs+SaSQ0Y5Epb
/FkG/Z71+aAlrd794LjfbCrBxnh1mcTOD2eRrvr9x1GIEUkiVmL90WhUQin+MgxjcYNHXq5PxDxG
FnZk7t1lR9BUsgbCoYzHDTj6b518UaUYEjITJPhOSZv7BUku77R9wDXzJ+0KXAOuMtDxQrgE1UDi
xHZVsNh+/aRiV28fizOLH9VGZ/XIUzVUkNUaVucqfzWkGoz0vgdQ4yTEit2btfpKJ7A6W1rjsnbt
xavYjiWUuM01bwZvExQQaOPfuVZa3DGrs0t3IwrVA0fKGGHCJ7ErO8qqXuLVQj6jLWemyAM5caYc
6m/ig4CGZzKEy22vrf+wqwOLwsQ3F07o0TlsGzivtwLBqCWVkUYDXUq+ngH33KmEkAoVvNw2J54f
ZxAMXtH8ke151LFwSwUZAPxBh4xsR69Lh/opuVEZW5CwOI438GoAeww6RHcq7pr47mbcnguOYQGN
FirHbKdeKpZpcBv/oE13PhQgXaIHY2gUVaORWSqFbtxOS3ZgfkvBrVXEroFJVI+I8yY1v4DNBwPC
eZxAlFR0xYyFihPXZn9Enkha87zSv50p84ehDZ+J8d2icgNKJZyTNAJpNqXE65fEYzwiqWOu2+AJ
xWlUKPgzB9pA4f6P4nfxLoKc1M1McijoXyvYJNPpr8pOUe3J1tCgDYw6UXl37s2//FLX/SebIgO8
PU7ihhe26BjOxzjV5WbMiN8CvRkn1xCWe5y0Jx7Jm3zqB3x19MGOW6jM7THerr8PlqjVpxDTVEyh
TdoPerSczDNA4CwGxaVd7wWMGPcQASxNUKQZkK8qDumP0F39OJ41o1vsJctLqjHIxu8Jf5Zitjh9
aLnZyncijkcBto/+nzHAeTcJJxzkjcRy7SdGmHXZqjIxcXJIBjj81KKtccFpWh6C7bBOisItF5j9
VG/mWLth9ltQ+COKOwj+Ees1t2dWypX9EK0X7DqbA0LjGPB0Wlyv6L7yPVQMVucVCYunEK85WdhR
gBoo4HuN1zItLoWkOPK81z6vOG/h0QKuKKhyQ1amRmwEFVnt7h0CUjCu5nWb1fP+Kn2fHQSnobq0
KSyxe1UuwmEA/cWfW4eORvYt/Hz0NpK7rbnz/PWFj1dYqnEKiuUlkPyVGFuCOkTUtu9fvCs+qOZT
qRjXty9kPHdSaxxJ0jCaIwHdsWNDI9Iz6shyKlvEKaHcoG75Le4RMesYQI8jJoo0ooJC/2i8fDE2
vkprb56bSCVsYNH1DS01X8RmlhHnQT1APpkdzQgxCnbBjqVYEeOsHiU3RPYI+FSq2qu6k5LEXjMT
sWANn/TWt66+MolhK6czMqQja9ygO5UWwQiOIZi9O5C5dArtyK4vzGCHPAFLtu49ufmfkf6RSCgb
ay5GUM9+uwEenc05dvDPlDZl0Pz+Yf8o5BH5xF6NtuZ3PzoHGbDFHrJRh6lW1LrezdmQL+NnR7pR
bafY2UJtO9kIQ05SoRn4cg4k1px7vzmqmClY7opaFX947dMJrklDnMET60GyRrx4Yc2HlfGEtpbj
wgB+Ougg5RWz96n5+wUcsQ+5DYEd5Kwi4rmQxsLDeJ9WabClys5xnWeyHUDdzhERchJDBLU/miN/
ZBEwqUHPW1ys373NXDZgNxuQ5YTxnap/DsNlRK4DZGErXH/LhILZdBzQRKRXb+C2jQc+PBTHBHP2
dZCoyicKX/hTAAmkNVcuSyA54OiSwtOlbXb4fGbafQhxMXQOA+bKNFq+d6zGpduqusU486MTMZJc
DSfBuWpvCFm5GTfNLlCJ/GhvKjtArIyWmDRQ7asit53VN+9I3cWcBTt3Nkgu7CYzVjcv2BauuMBW
Z3WpEsms6q7lYXWoLeJ1YkriB6arLgpeqGpR1T/lgzfKPpI7dXKT8jbFHHZ/h9NKrsZVXc2DNSRV
VqkYFPhCeOvCPuYG92v3P33vngIgLzVjgmTmcfnaT7jGGCWS7mVZ/P9PtdwwszwteGcZ5mauZcPf
24HPuKkDJj4X7V3rL1GVVuenwC/js/er/YSl10stvOu+kGeAC69wBk+W20gnXsp3gJ0OZkzkJ2pO
JFkdkouYeXU5ogUeSxntySnVkCOQ7ejmeRRha0KKkI+9Nggrk15XLugu8cWzHHa8F4mQt/dvGJ3S
ieChvpVfZWBVTRGfxL0z3ForYIhlOtzPWVMSSde8eHIxlPJWKSf+grYe81d+h0vFVEoc3rw1eBGz
GjMkyLry97DlC8J63xtgJgu5uNoY53YcD7cB9aL8gR2aablRPEllBzl7rlyW1TogivmX6ktQCvDz
Cgkhl76jk7zhQB1lOl8ZoVhMRDKEWUPRwk7nWzjhXgSzXKkUsZAVzjywlRZ6UgsJ0EVN0tMB+0N4
XYSHxR4K3TJECazarRFRMbkgG0/O7MdaL1noMYeHVjc74eXFNUP6esmBpbKOkGrk95fEMXV0qazI
UXL4VnOJjn0fpHZZCBB9LsgMCnNPpsxdJYU1A4Mzp0EaIkZYaAhkH3E6k+5GP7DeOBv5KC1WKYAA
1jq5B6UPoBT22mEczFNTc/6svQNvCY2YQ1TsngNuzrzXtpY2/tkGhGfE2otfBeQYirnLdMuPivvS
fCAuM+nkuzBiv+9vqSa7RLeHyy9QiIP6vQhTxblV8CoyI/7Uo9T4PMLLUfjewwfEunK4JwA7jQA/
oLTXaeRP/HyAgFqCEDTFPynIJw0QSubmuYPp+2FgnG7dfCjNQRINHPkphTnxLJnkFiN065Y1y5OL
lxQrMxLNVSBjXwwJd1tXEiuzZlBZbTGqA9AaKZTTzHqZk6yx5tOpkht2Ql4YCZsc6P7mPsLwtAot
1fvbQvL/vJXCyiar/rUh6keKJBJdSPQO0exUrfPHqK49bttVd3F3SJpILFcoA7MG0qesURF1TR3a
JqDDs1jS9JZKM+KCBB0eGIQQr6u+K1AZMeDNlLQ1+RLtsOnprWYwswSnq//nSz23aNhBeqyO0evg
UJt1x4FhMsuyAdZKOOngHsIylid27SVe3+2wM9YH0fScBTwKeYobiX1FyAQhoqI10euCK+o9OPGY
xUKSxIMky3H54u7J4ysO19CmbE1cnq+7JpZbxLgxnb3Ka3JeU/wBqjJA3M/JKv9ebksItnLyz0Ze
9NUprNDa+xmbzCuxtNFG0hehKnvi09tXLRFWMUzILawxLJhG7RrYN6D7tbMVgbpeLVBex8LaRJX8
l0Ad67YN2mm+2mb548YKdUetK+ywYlMgmYBhsBgnVfNzH89zVrEMGbHJW+1C/F3LdQnIZR5f38RD
toKU3FqKqYIII6FVx25Z+/qH93LpAz5oVeC31fBbk2RAPwC1FC5NlqwAJU7ELCuZlZBo4kFVZFpL
fBFO5DOcau5Iy4ujRbG88/UxBC3fQ71iSK7t/DPL5+9opM1krv3RCQkE6A8sVxKscBY1EcX1lV4f
ms/F9iyLSfsrbjjd1jeWNNnbnYxE+4bpvbhS3TD1+5TdVlMva0e1TQEk4qgW409rHaF/YvO/PFNI
OTDp3a6JPI7kL7h+7CoYNEYJ11WzFIqe/eekRKyR3uYyZz2sInk7IHqTchT7cynUR94CrhrgLBA0
iBAyJYbjyYo4RKyFXDYzpepDkv3/xbjtG6ZKiesm1iB6P4nzylHbJz0TO5HOFeEYXR5CkiLF1d3t
DSLRTfDR4/dBpPtVFsuB56Kao1AQAmtg99oM8UKcbLEhDIifZzZ2Unke/L/u2CM+6E9YNTexpNks
Jy1fITOnjXCSH7sYrrcq9+tRKeisZas+Wg5D0arakJG8z8RGOYp7gcVTiL7NWQZFQgDpPzn9LPMh
ytPCSubZQ2il1FAJVnnA+DJG9nP85Ux4kshtUxmrxAAJpBz47bQzNmjOd6yYP1tcLJmKN2joxHdW
DgtzUOFstYAcx3adZTBgVMZ9CGvackY2OokGWxQhOYMs+hm8ocm0HHu59NYqrU+ucpF0cwFKrUTJ
71WpMD/l/17hqf0Lwicw8qSTxEJ+KrrjivLL8+O4lh27GSgnKuD5ibOIouNx1jvM7Wfytvr6MK1j
HbskVLYq4uD0nGXd65Tyr6Ch7SCEclt3Rh0Wzul1sCdv89LeBskOtdjFc1phh/+4VXGm80k76FwS
zaZ6+X5A4mbfTDbMgET4HgQ2fS4eBlZUshayTAYqBZM4ee/WF4pHN7oPiDzqYb8OCtEwej8rIPsa
g2gdzzF034kSkQwDd8FjbvyH8d/6xKuG9NHHZIG1wPVxLybeZOMDlfWw3ExxPvkXhCXX22SyEdoA
PGc3kqd93mu/RwoHHuh188U9NnQYZtg4488XkESi3iCFMVMYetWeHNb+HbWgd21nwtuB1/ALXT55
1DiHSC046RbwrJfZvqizmliSA6/USm3mFTuTMz9o+KF384f5WnMUbkqwmUqH7Ui6PfB4Tr5K3JPx
Unqcnlcm4dT7Ut/I+U4QnCbVHPUMaRJ4s0V1XtHtNN7zllpXrC+tzlt+OO9UUpjghgEuXivEqzjj
3RhdP2qr08tvKe6wMZTzjNmVmyu7MY4Hz7BT6Z//VFgQP01A095GiDrHubuJ0j6ztB0EZr+tJydF
M4UxCzp/DUrDtFn+W4UsuzIsxhomELJ98WO/rXw3J1tvz1YJZLswouV3wkvgvd8FsqLgQCO9stA8
I3jNUxj3i9tkg0aznPGup7RVKuvqmGTe961MJIWAspmqgR3ytdli121JqMKHU4JirFikRzHhzOmL
hCgZdnca7PkP6WPyJPHazjnVqt3N+xk9PAlGEsdInRGPHewkgGltOddKBlPKlk52vEQAX1jGBPio
zxiW2pIKfLsF/HG0gyOTs/t6V+sU4i20WHbGTgw3dVMUq6xOmgJG48Mq2aFIQk7E2NJQo3SzvrWv
WA/J76hmXjr3DnaXh+aejAI3JjAMOTRjK81E0aQ4Fr7iieozDX8mye57u4eaYaK0etAayJFSVnEu
IXkS4f7yxB1folYYVfAmEoYsiGgeFlpV5aZznGBXl9/Pzv42wXNL0htIJNNeoU/Jww0QZiPUjLIH
cXxsCmaPLm/zHtjnz8RPriPDsSZ9maNrYDRpVkKATuPxltwrJT5vvhepWRVOliifZ7HwCz8I4gIF
89ux/omqGJYs+MTKpPUZ7Yegk1zbHoac/psL0hC1kFX0ZncamCg1hTqR4yiC84ejc8JCiRRjDpt/
xaICsytUKRAtfLeUOeSAIxaaf/cgT1GvOjsZLV2inxwMFqmF3GxQcmnGtExypg3lvkAOjIeDX1sj
bTxLTWrHLmrYSHY0kK8VDiOaRFPbMZIQknYpoIaP29Dn+Uuy13hx5YnA/QNcpkAwVwKmquTKZ7uX
sRAzX2R+pqzXlBwT5UkSLrHYSZacfgC+5RRCbHJUk1sUyXt7WXY0uscN2+zIDJRvpsp4K83zaYQM
FUd56L/RZbjls4jw6nRuVVQ5WSdvgh3fyWYxN4cgJLy2k40uCOD74YES28KtHMBfbEfBoCm7IrvY
Qkr3XghTJdlLfiITPm/eu6ZDEBvYLi8/Ykh3L8Dq3+UmaZmVfCpk2SpA6PnD5gAwdSVhn2XOiN/g
/5BrZn1rmYAuKjtXu0oqhxM/AAg3g+w/n7+3Vv9NkV3hC+WHnPGHvVhvu+dQzz4ZYw26Tw/GEkzt
E+M0N7MGLQ7uU5q0Rw4MzAMffHB+s3Uzn3+fWN+/dUN0fJUSLc99OryydecPuV7cfQJOaNJIO0I5
Z/5wh4SjM6ybBNQ6mvc/swgNZfvJZSMUmn6p9s1jt0OrCmC285NLrVwFLKZ3qI2nmtsg1GJLtqyZ
J3MfpKtiGEaP2jhpgSebKtTa+2VELn2+oVPO+0uO99Py7uu3QShAnf8mncPQEp2wjQjQf3E/rEsx
DrLKjXR0wfzj4T25j61hNXBlSm6foRl7nNstWEXmWMZPl+BzKYfnw6vsbu2TLqOu0Y9Uuq+1CHpl
7lOjDu6GqgvEodrH6n6yhCMpw6iuM0vKTIpGUEJ9GG0mCwe3SnG0reGhBSJL7IDMVRTIrhyfY3Zj
3iRgGzQDAR8s3AfrR1PPoGkdq+Qrlm+MLzp7Wp8zTOyuWyzf7+oZmjAiYHxXRiPBdJNH/V6j2I0E
DWqjYGJkX+MSYE00dWFzkcSxek4n8P92Lzt1/7kk5OEQjKLgdY/2jc/e+5KoxNgV6X5lJWm5hZUu
Be/k9nRNPdRTUJBXv+hHF7IChVpUMkz3hkhKxWKt13ysaPGsJQBM99COuKvI0jifPgOEtMmIFdoS
LNrdp3W8to0VZkbrCFHV3aFqqYs8rgzotsUia41YSWHqWO4FK+/mVJC75+AOHLDOv0jYC9piGRrH
6DS0yjeJjODQE8K6kf43eULmx2aY05ZPA3gXSxo89Z7S+S+e3ktLEE1swfJGEruBgFIoCH/OHw5R
6aLuUJG3wtlTnhksxXeG3BcOI5CDSXI281uotse6xrRIyeJZV0oz1ZrYmn6SiVkhiLzvjEH9jooy
n01dnYYQa42H2faEqVxctUR5cu3OYh11z4p9YX+eGu/Pc9rWwCquk5ZNEoGu9OSA2wMmVLraWotN
bEE8NGJisgEDt1v2oym4kHgYsVIMiYi+wv2YUI5GknkaeY561yZvqVsoNI/vcYO5+O+Yha8zbg0Q
t+3iB/+Q+oP/ioS9JfCuQydAgLntKRD7TIIV8Bz46Y+VJFfeuYIheNFL1AR/L290X5LsN6Ejue/i
LB3zWDZGRCMnt5D4a/SjSWQFAZtyJQVMlJYatipSoxzwbyc1tdAbC9JgacsRSghkUYmX3/qvxbRz
2R5Zd8Ie4YsiFyNe1AuKUiKssTzvLWR14fizJ0OmNsWr0nhznwagwMtq1N2IBu2WXKMuPYbTVbvD
zGszsKUt29f6+QYkUqIcyCibVej2bvOUdezWBLnEcQhA2M7DePgfX0vAV9lE6Qyqa1Yu58gPHj/0
ZRwOq+PC8foRclKP52MUd50AmU6k7xHm6L2r6RmonORX4UhP9h3zsKjbhiJ44Hcvp9YQcW/mD6wp
nYgbI0Z6B5t1HGvWZyHj2PvgzkZ+15S4bEEqViTJwpVCO31KzzVunb5pjyHabD2ANU71CXgii52U
t15tEVUbOMMwh36S35MbAaiReY4+q8De6VH7TGBQCr11q+ZaBQew4igolPrrctag5qRG6FHRTN7S
ONEJfH4VGztW7HbxrTxOt/OlVDH9Ghq5sETAj1bD/xejJysYEAAOPctoqjLloqIj2GvOuoGZbjNh
rHiertsA6gGrm5MLmvPsHCu4PL5KgRLjjsPvpx8zdiHPTay4bDCkmOaG91tN70Py9p10rCUCU7wv
hPcwPn5eZhu62Q3hrz4UzYnSaJURshNIyyJlAmWLfT0QmyxHyhLUI+pGXw3OMA8GWssPHrErrH6q
WrDAgmEwtzs2zaDodxRBvjFcMbl3KeK9G8wdGf2NhI/JEvttC/nZYeeeuD0cSemlLUKwUbtUprKS
t3qV8REIAFTlndp6LhywTNAgEAbbzaoSOEQXu/eFR9g41HLlu6j8fMX/Q8UyTwl5Db181GY0iB1a
xImUINW+tXDeh2WlH/5rW7/WPp6sdhf1DM1ulAPqdE15QnDJgG9BsCYfgWtsTJJL1zPY9xP4TMzM
iwdUH5eaDyhhlymTJh5APnY+GbmLKcuO5q4keWMBHvFhJlwisSy/+eBFjRZSmi8w72aO5db4OJ7z
e/W7D5aqeI6hVIFjpgIM4+6T0Dihji7qPawgo7NjgcLVP9VrvKF23PxmB5LG3V9deQg1J0oaq0sW
mL2RWdzX8VMtvAtGjUUwVXH75fPyk7u24aeITYgCjnKF8npQYPUZoYTCnGOK343cfkjRFlJEY0nZ
k4yHA39Nba/dftpPxm0TDD7fwv3rgFnDw3/oPf+UviSxzG9lnqQ7KJ1Xb/fFwqUySy6vUX7ja3GT
6IxiXZfnEsL1B73WH+2OEon8NIdN0G+L9o4Vi2ZtG7HctpEBm1/7PMcq6L5sE6pXh5xbLceeQfgX
K+PEHwp+RJIrrIACwGiYkMzb5fFpnyp6Ik9BrN+uF+/WkM7vclzAAMzPCAFXpKQG4+bP8GKumFJk
VtdAWsmi7nVgCQ/TZKka9gRtk/E3BG1aRw0NGiPC3rnPpvHHEmIM0puCL4tcmy93PZ8TfGb1IsYz
5oUnb7ikm/2q+qJllb57dGsfJ6bue78B+B922Ptypp0BnOBDkDBqxZniG3qCiLP34JRP6v8X0Cb6
ZRMZXrPbmkp2avGsyvgfIW9e8xj3x9EkoXrFZBE+QpsYNsm9y+RvkW3fwdiliwjn7yGlCb39Y8jd
/ho0vBBLge19PkyQLcGE3D/N3GczDVnuAap7KrtA596KsbFJU/lHv7jlAxahbtLSVO/Bdudxw4ak
94+W8agWvUUYk8YBM5rEgYrU+yaoKAnsIjs63M+YAK2ulfwyK+MurNXrFGh+bCPCM3saKO1VLuAA
DS+hzpKDHxuV5j2783vMpIOYd0ZtiP9buhsWPebTaLZdc18s2RFzepArKs8XLAxBa8tl7eDYiBqA
W2bmC9TtSZEB5ZVB7+BV//P4VG5fYIEXMkXHfgU3hemncrcd6TnOYRe2R8Pcu8wEo1ZgZRHVtVXR
aSXwxIBrjtHWYOiEBMeroxtOA3ZSgehb+hacg2mKbICyMrvofAb+NhnXUVNUCJPEPFWviOxgzP3z
Cb8Jym4Mj7Ygcg5w3xJxrtX1aYuD2vhK2mBaKefprH1ead8IlCSwsHS8Iujx05P+/4Mh+1SLNNC1
kJanfRTtprsMg8xc3dsj3DRIek0DoqY2nQbj/rKg1Vw20bPOLn+sVqUWxiPIVRjI9O8we0vKPJ11
JhfS27xeGiKsClhJuJvgGILa5rbOJUccj7j8VvRrSRNQr7tL8XAdZGKQYiBZih3wDvEgpKZUT5eC
/OZN/5vkNPYacACBniJjjriTnPVqjd8k5lJZaSOlQjTxrNR3EQfL2lpmHMj3tly8XCo1knw0ggjy
DqP4L53nv71+NeZ/1FzhPvpQNGF61NqB5QhfO0Xv+Q2SFvRHb71rsSs2oA7jZRNl/giVRYnR7UKk
6l8llD76v+G6YtTrvLsgei6N2BOPwxXQd0zNCFe6dmdlFzKMqAzERcAqiAtePXrUQw9HGDx0Buld
eKLgk/uKw3rD9ZhgoDWsdybPEmvWfAdLfpiid1pdhfRkUUZi2kPhxT59rwvM8b0cT2FKEWW9C/WC
GZqW9XI2uxMFg9EXRKkAHIDw/0KtRFDNHH2VaclRkmC3aMXGwtADw/fSA2uS+f9d/2zCSGzXA291
XfcEIsrcmnnWzZ3/GI5wFVDm+vWnzZg/WfA+nquU4DG+tRAkauDxWCx6k3DQT34wR7Xocb+mPofp
ehbZ5zRX2VWM6Rz9H3j+4So5VVVv43kDiJXesKbqb0+gGU6tOEPT0T4K2ocCzZLVla/8BDHRQf2H
Gf8aGJ3rtlgolrEyJv1QuXfosYmtc/m64w9RnAINokbXaEJbd6ekFiyO44X8PDXNohybp9MjUewX
ePJyTCaxzxp9r3UdotDDAHZB8bg4OR8ecGUFbwiXagMmRrxGFTCbtETDQUqlJEXKqlm+pD/ERFni
upIC9YVk4NZf//+Eer8hycBkiM2x47CZAMMkFtzJxjTvbceaT0iv+r+TxkxUWgXwwzi9EA6Bkfzo
5j+NfM6ulpQtSbQ701U1P8bZlmKNhx/wJW4nyesOcKQcZ3QIJqg63NdPBjAHs+M39vZuzPZtkdKp
oLky+u/FrzdcLw7vbQXtfuS8qkNJ+zqdUILeYc0OlY5FA/maNOKcHE96YCrf884fyohGwI9gdyhm
Dr8ipJP8QloAirs/FQT70Wca3fzdTvvtiy95qCecSwf4P40JYpM6+Ou/c5W2YrRISSAkNQ7CVKCw
J9HIo+FEcEZBuQ8qVIDps75BM0Ni04AL0Z3hP9Kc39zuXzNeVOw7nH+E3fVIMK044PeDKPLUih7d
gaNKVhyx8//TOREmEFEeD3vVS9pMpIsyhmCZs2i27AEAM2MSTinowDUpdkc47+SGZFDKXw11T55Y
b9fpQnSF1GqVlYvyMD1+WwcQaTb6z4ZzxzQomRwjFhPqCEknBfr0vhd1bFibSNTwnA7EIJhAt1u/
4ZJdJ1pW6pBw8PNoyol5/wnPYXH8S+gSttDbQLawNS2flp677WuhD54AKL5RWCcR17h6ZruB4kAi
6qEXw/Y1YQRNL/evsVTsqr6NmHxPUuMAxDlCb5qyJ9Kp18BpyL2LdNlI8Gm57gRSMs6dCbwqqGZP
HL5S6uhhUkSrrY2fB6c73SAqujZufbHai4oYoesRMlZ3FkkXZvU8wo1/kcobINLLRw123SkoB3hK
UZS7xPIVbxObLqXn5WV2r1eDNZS863mR9C8b/d8VbJnalDeiHGxAApUnIjCJzAVsyqWGs3lCSOOj
vtfe6Uj3EEDFtnLdNlLlzwvQ85zsV1SYwtS2lvusCgOVPpqlucGS5tTeFUpOd4shAzcwCIFk4cEa
GDU3DkYuclUEeFursmBsSIqI27lRocnGGkkpvlhaXtUpE6POkV0ShJRTBc1G2rQ9RDY7qQ4sJgJg
7BaU7tPPNZ7KU6BwA3bHzAKPSh4zrQOr+c4kcmsCU5Fig83DC7CRNkLSrIN1xnsZ1h3w9ddXswga
l5VxtwvQYkyIE0tuS8tlIbbWrPsXVb7DDZegOzv/oeeNCRlbs1sWLQA58OvTruA5os5iJOUWw7XO
7lXJZsv6YvKUMkIr/fk2nHrZCA8we3llnorR6wlLSuNc0yhE/8GEH6Z25JuI1wR19bHNKDauxuH0
8DSWzBwxfDyKk/MjyM60wjLwf8wq0qOjcHIwvoUKg6mOt/GtBevzuPjESWgkBvMRsXrx8zCGUypq
2rlIKjCG7/oEdBfgtLIrQfxWP+Bs2JzipHc/aAk+CUl84SBjSQPvrMygmTItBG4thB6fCFbGRjeU
Nc+ecjZ48WA4QmSAYsxfybSwPOEMVbvY4QQI/eT2WkHooDmkv0bKS59GDAskcJrv0njDoTlX5p3y
HbQ/CniAxrQasomXCly2T0ytZjNhXlk/9IbUC1i1SrVYioc9mAC01dUXl71gfSv46IMHP5BX0ewW
B7OFVWw8RZXMKFjR2cBqV65VX40Gz2UJY5t20kENPiBtnfBiDKNMeuSgLclLqNDOLgUxSE6a3cpP
/k8bPHUUounZ1V/oAxhr1uGMNqbETwc5P8bDwT32j01zH4eW7RiwS8vuxCNIDNP7NHN8yH0MKhaT
wtdOz3Koh48c6/IXuRGmB8x0EcuIlVl5SL76fkSEVu0S5HIxrODYEnH8YqfxOTwg7LQcUYPCn+uo
k3pWgmXO6wz6PAxOF3fbk4XzRaApi6R+GEOdv7oLnuKqrr81C3QqnLeQ4aJE+3E1SW9pQlVNMWI3
EQ2fmlhnQgsXRYfIfBoyAKQabcjc3alkjLQoei9BzycR1E0a1zCcEmJHP7NoScR/EgFxJh4o34SE
S5nh7RFWzOUJfPTodFL2fXB/3lM9aTtaDdfUBPT5WLPkHF198wjcjZCQ7tfR6t2OdwZoS7RFsBk6
SdawZuUHh3Ba6Jq0aZB2KJMTUYlq3/RcNEx9l2bQERIXCLvX+sPk0lRAqr0n3YlsWwN9J5z0dxSj
cMnkbc3b+OVClRXpihgbVXRYShCvwaWDIhIwodgr8YdZAK9iMqKQVadNHbpEzooHhJlGUs6bnvih
koOGoqcMAEL23etcVme8UOgQpZszFN3Ac9gycV59OOxSrhI6OZ289luI/Tp4mHDKdt3qnyHyYswP
bxeyfA0cMftfgJGYRi33q1STbjq/VSrWImDb398n65phVGExc6ul+c8N3pJU+gt+oCnc3I9Hayph
9thUzpWG1aRraY5RsSB1hzmXQauZlRnGzN4QlpdlnZLfg5yDtoq1x5WhnVguyTpbjFwTheKcb6Ve
WqK3hu6sKcxOQZeFf6DKr1+mEFDDSc4yOsLDx+de2cNdQUY6YD6TKxZhQ2uncNETZEAZYdzei49e
IP4qdc5R94fIJhGXnrStBanBTYfs2jcuk3gYksEolDJV1DhdNMrBdznrxGe4a52ocblOf1bCGk+Y
HTszJI3L14aKsDvKx6TRDZoXqUe80XUVmrNgRvce2w4Q4bBGXs//ieNrIoQA52hmeGCMf9V1gEPh
BN9QDXdOGCWr08HIOtmagqt5wrR6PhiqzChjpUCZzis9zdpuxCB9O9qnaqHJpYF3EAHEKjKy/dKU
1HIOsc+gHOQp9ZwIYQWH7JYHjWdn4lTkj9CzfuWLBOoS5aPvk9yI2URbONvz7T0AV672lS9TTLVn
4Ku2JGG8ieLsyxzllPdO3Mnp9Jx8QwY9uuoxWOGHd5jJqmbVsKHyGphD8ggyVvgw3BCyd2DBjV2D
WHyfAYR1HrSn/4NoBlGDWu3G5P3Ag1BUvbbGnAJ2HGfIMqZ5XFh/naJCMuJemmZXp9tk+wSj9TPd
4gTzYEZ1CnvMyT4J1EKPF3OulnsOflWlw8Aas1yXMz0m5vN8eu2UMs0NRx8kxmS16hzSaBOQ7Yx9
dnKiJP9shxiwfgSz0wBuVnVxSeJyZ3rLu/1yTqDQMsyuxqm7N4nZZOVeWSlBspwZhs/YboqcxNTH
gpN89RmAyjqYUhsDbi8MwHmF2y5+FFGFNfB9N7fl+Klz2wP3s9VppVUCnEg3Zw2abonVytazzcMv
y8XHi5yO5kkCQheCcHY8csBW5wbXlo2muEMXER/yVl4ppjBhqGbNA2VkmeGwq3yEfUXsvc1p0Kzi
deQ2fQ8DkiXevHHVZQ7CAwsaQF99g87BRmYVKVtQz/O5YcqwURTyPR0XwmzYMfCmmEkbL6CzjKPx
DjX9CdKHUMMrZX+deyOCfzQu/Y4Tt4LK6CiQjlmLuCmSPAzMLFocdMPmCe9QsdXzYWOp9+firGU1
AszeQbPzV6Y7B2E324i/h5YPXVnmy81HOFTO2j/5T/XCYuySpITN1hjTviUk7XKuxr+GQAZg64r/
jGCjNc0NrAcvCxoHLP91IJgYy+ekilUiXKCi3Wy5xizVLL6rDCnKAa8e9UbSX9S6to4MP3ODKndL
PmJp7zs9gSM4RgkBb0byWf+KruFdHDO/6fYngGDSMA9gclc87WFzLoTuE4KV7z0kr27wT1s4eWbh
kbKhmAxFsvgG3ozCdgwIwHVi1AW04xzkY39TMHKBa/MhfrtK1pov3pqXNSBoQzAIZ5wQDQ7uQI/h
kDBaCnkJjZ3bCTcv2neN3NMIfBYtnywc5IWJmOdDe3sN9e4qg715h0zZSQQ7GEo5yIVlVwSMMmyB
EJiYswvamSQD2spaaoCdnGGugkLbBphNvtNxE+xfRfJeHWzEFl2WHa35gEID5/RtwUx8qjGzDri5
CVk1z6LS9g1sllj60VoR3PQVCnNZkldKiA4df6LGKiNLsiH6R17d4e+hAhQbsG4gxc2FKyHPEZmr
4KkmQb1DLyN8h+v/kqTfQpfCg8lFfiIIQmhZ/f/0FvQATKEKYbRVaJFAG3S8Cg8VFTBXRaBA1hrj
s+Rrpw9exqrArN/7M8gkKWRzxEZqEpw3pq6hEfrrmeiTZBdTwIzs1vTZr6g3Y7gZhNHZEielKTMt
+eM4o7c5f6NvTEPanQRE4bsWwyHr0ssaTlu0qWYmYdDnQTLzzMYFt1zeB6kECJBevn2Y6p6maCil
IDjiL7UqCcUyJmyPOXQpC8aoqlBTWwVm1ilxBYI/CVPk5e91mYZVc23hePy7uXatwmltdu9ACi84
O0HF8oVjItWw4R4CfMGDCVz5ljdGSbF/XgQGFmEcnnxnH4w3paoAiqB5X8WzVO/meqhY255q9YRC
ooYAgwRr4sIsl8Ndxm335lgGKATrOmU1Kr2/6yKpLYJpv5URYGpSAmPdND0oH8nOg05Md8hUJCPp
qbYlOlfP0S57p9ghNabxlfvCVldHM51ZIw3lsyt0uJoQ4GNUb6txcP3NFmURwmprcqg1biK1IBpd
ul76upTdyiE2RzIeQBTO/zNO23AiOr20J/12sv6Q2jn+X+zDR+7tOm+WpE8dDCkaiejOJa9HHwCi
WSJE+SKoUYn55v28tw1zd00EN7mSxbBCYfX+Dmpno70BLKCU5+Xh0yVyzXV6Y0NYhNbRdEPTgsG8
LRqiwhgNZaq8jb4z0qRtFfbqVxBeY0dLLkqYvRdzbdySeQoSzYGlCV3CXcUHNv7L2357++s9MHzp
LsfHNFsXzcQqJVTO1ke6y5cL7AR3hPHJKgIoho8hZg+9LflgyQ2XO6G3amnioOQzHWoBPAAoYnpY
17MB2CeVaJKL+tiyA7orB+xr/7MCCbv9j4cphotZM8lM7wv57UL91ovNAoRnJNCtvqryFWhqFVIT
OxDsNTc6fTtQrGE6BLmRRhE+E4llRy0F5Nx8f7JkV+cI/Ui3ITeWv+1Q5ucQ9A5OvDuxhjE6yTJc
sCZJ7YT1JjQ+kIIF3bThg6TyxMKLRPQ6pjcL7a6HJgy2X1+5UZzLB3ormI2zB95ketvDGFYnJOQT
C+9o9y5BVEN3ToHGGVHKABHGMtTCvZ2ysn+spl3Mz+VloV5rL+0xlkTHkRhkbcbYDlM/ZbXmnZCw
aCMHT1/8M44SBJwsjG7MPY83alDWwrEaNGSvgjdy2Kr4SypDL/FPfnTp6fkYhmacB7czmIovfWWp
xXZHqHD9+dMzg4ehaoR2GpxfKrxBxLyvfStC319KgeXra5ijzxYGPsTIUUjM8wlXsdClKTJPqMap
QgscVXbeleNLdvE/fa6gSdnu5mHA/h6RQp39lVA1db2pIYsNDkWTHW9N8TCmHCog1fAh/qdqZUQq
IAeNduyFVp+k6JKvFa0xnVXDuG/vIOS7Nhs5X+5DxBWZvoUeOa2LTaKrOup+9jU9zUD6tf0vtu2b
2RZ9bbQVsU9speUMlCrUm8461K5INSQtHT/aTxPa0b2agntFHfuDA4SGevUFaS9nijXDtiKIEngj
7p6ZfhNUbc8IeXyX4PKChXvf0RbFnezm7PUFgVNY4A7ahpfeV4adTDXobVQAVspaJ+kt1NrbRnym
L84jiMcBfbRiByVbOSASLMGWewt7n/5J2/Z6JPkSyGQWY6UiyRN+heWaDt8qM7hf+YpNJX6G21OH
N2R6Ky08Gtv3yLFsUtUtP7LUoVer3U8CsZdpyAMgPGA6sEJ09Kin0Yj1Vzydmg4roi1AR499lWNU
JMP5E/jcWyfJsu7mDQlahG0hn1cND4Tc3ftheqbqlx7Gnzj7KEAas+mCI6wiTcn0MOVADw06rJRV
sNx1zxA8n+pt2YhbexvUzdZv+Iqba4Nt7ZiS3UAxCZd0aAUXWdb0oHgoLpeq13NbLwbkQDQyaqBq
ZUGAQY31WMacgDbltleJkmdOagP2RvrQ2JIruBSTccate2YUmm6z2Yb62hX27gsziqKmt7NRNlQ1
ypDtjLUOwTn7V+WZ042wWETDa/Eh9SyPP3KemSOJS6JdTZAGY6qupYkTQv2m6vpI4r5vrjnfH//O
ZbK88VRkxtn5NVXa2fb2h52LXDYc6aPqhpG88RRmQUGtFsVgf+iQQpP0bFQkUCCC7MHifXNsT36B
tF/FVsF2bjreiQ8gyS7CdcsWzDKEULLMeSy10xKcbGZ2lLeESoE2IG04WOmrtO2MIyYwGq5qLcGA
Y5+LBjHtRZExH/u4i0E6kwJ9qBaZppaDDOHwFndAUjcRzNq1uhNvi7rP5v6Re3nZl0gA+vySWYkD
mnazfqoDL1azc3INWO0fwypIll3HsEHWizwH+waJGziR4hAonlutUB0poqAzKG9iDrOCpUSvb9sg
FqCCd/VPZcVAd2pYRo+ykvVuhWnnd7tnPHBdlGChdARCNvOVKGfLvr2htxA3rEoNHcRhTA+Osvjl
LxkdzyZoncOlhtTkZcIMSuTOQ4SNl3/IgrgraCHO/8W8ww0Qvb+hi44KEi7Ia/JaI/xby1hrtMsL
KfrbDSj+akbPMjvZBnA+fK4VsLlTDANCdrwioKafToxLnnnUBUtXY/pgQDQ7+N0f1ArORRkDIQNF
/9+vvOTIVJwbji8PTm3bhu+qTPzybAAdP61CHO2ixtrvaa3MUZ+dutjJQsAh68gTGS9zfXy73HAf
bEZnnKkTH7zrhVBOUa9qVAlV8202a3C+3Eq9+BXvutFGI8eapQ6PnzKhfB1wjjRYomlKtH5oWdVY
nKYlG7skFe5wM6em28UzNDKjrTNQ6y1S5nhM03rnKJyt+v6OpME8SEFW8BaB9B0ZcurnZjTJ2wcr
WR4FdsfWGlhqLIKYm6u9ixuC040Tfo5QgC94uwKAWxjT0/QcVXBKz+Ah8B9dmm5cXRTt/Um4EHbU
Euvq4JYgk2odSNLIlkP8cVlpjmhWkLu9vmVOZMK6LC6ikqSgWGbv24LF4PDKyGXYMd/AtYAmgf+C
daEI5k0lcTNP9rH7TqIvbCAKlvXIlZrm0QeijoqyxKTJ1JAQKMLha7IQH4FeE5rtqwNYRZfFlvK1
b9EvTb+DNwoVSynTmQXcnP8XkOc14EfYpV/11uWncA/KHqeRz6OZbBWk9NqQCY3ph25V80c1/j7s
VYH7McuXNtPC7YBcpdUZtLZcNNaYd0Y16xgIVsRBmUb3LeNRmVkgF8NAH8pi/zdjc4linCQzVUjk
2Ka7gmEmZK5I+YOfgmpLiE4k8k2CZjYFlbVfA+wkArKxGJEyO0QA2uuTxXXCvzZU+doPkiykH1tL
pbQZUf8eEk9U1hH3DmRC3vjRn4cTAt3a3GURGRYsM4QImBm9NchAqOPYGxHuCqpnpiwPdjHhoPlW
aI7Ysa6bLLY7cLgz3B/pCvSeoYKO7TTQt2O8KV1CuuKtRckLn817iGf+NmI9rROBqlGSP/I7WzVG
MnM3NFt5/XN61ocSrymMcPycT5CyfbujKauGtTy9h8fP4J5UZWPk1BGlboxY5Ejul+IZhMpaXh6q
xmOl08vCrD1dc2hwyrLGdw3MLspILmIhsYBXNk2C58M/w9lqvtpnzlME+g6JqlmjKcOItohJS7uO
Uw1r18Yudl8EAkKWzJAOzrtt10SG6KmZVFeJm99tTDzP1/swfwUX5JGYqgKvv06RNtr1JfSSrH67
UTQP6Olku1+py99wh+fGggL35IcUB4dKg5PzgrldJnuepHRF8yWWMVJ1/PtF3Nq043QNPedW3cUC
bQadUywgNZ4i/fHvF48cBZeonIxbp9YygtYJtMTm3PRWO3sqxLzfWvmE8tC01shMwCy1HlePFhs6
wDLm6SdLxXP04UQZYSiVX/Ag8Ei9rrR/oVJ9JUh0HuyfKIY5IIUckUnDjE/vxU8KSJPi8C9SqT+Q
yWNEWpYssHc7gLVB58pgFboWSSZ0q596qHu+QC/FEIv9TaDFl96cwrEkYufRq4f9ybOhP/6VJqwd
vy4ASRNpqB3LuNFnaPh5kM7QLGeEh6ZnKhfwrO8xIGD0S10AtgEk6CfT85gXJdtHyWDugBCkAUBe
AGy4CJGEEnaiziBoooAkhRLXIsFJ7BdPjCFU4+HApyd2hDGyRl8TbB4JEO4jOpmwPQVKOXkk6s4T
sRdWbCb8GNUVBH39PR5T2gZAR4llOW4ZhYd+aHisGKt42W8syY9h4wasJygkVurpsYeeGF0N6XAR
7rUHXOoUMbrBae/Mq27D3YDyz1tDuN5ozbBtuMaOs3vYvX2ZnGacumAHpDIfFKK5dL734CulV5PZ
ZA1Kkvw14TEDj2Fp6TI+Q0lSr2fB2KV7Fo4Yz7i4elVfDpklGauJ5L/TV3m+tJEj4upDDMu/irZo
Hb1xIpyqPS6eqD31eHM4XH5Y8YAOdVpZtUwRVcSmffl4Zr2QorgMTw5AlBG7wFgyoR2HfmVHZOV2
g9eomYwupy/7EbACnma9kvuQJZ6m4pKdeY6iO0jXi4riI+ol/6dvUB82EKIYb4r3Slg+IZmBWEbW
OgDm2Qgz8cSUY7K+xlAhnB1L3O5DzLYFTx6RWvBXp/lRDiGdYBMrOd/tbh74YlhRtspY3s5yAvXj
Ba/uOKLkQVbnFgD0C1gpTcjTpKIh6m+D89myr3EHoIwL9fSjSzSrLjELiJBEYRQtdc541kpwXonV
tB9VDRnUTRT7etjpNakLETHKLJQOUGwChnrFPT6O9AjpzWSGB6mW5kRux0U47ON7492sUY14kupj
i1fZfeyjcIOequSOaK+cjKrLUe3iRt/nAVy/0sor2MPu8dbmolKCXXWAyINNqVvItPi280muw4tv
JygGfrokCqZzbCPvsJWX/uEBpyBSZ1FjmTqBYcCFBzQcsgByFJOeZFiLQJUmxwfy/d1OLiWBUp90
xIrlk792ngPb2iQkgbi0z3/CrMzOZLDmTb2eAmVQVR5kDb9Nm5Gf8GveNtKGGomtepXOuU+g30+6
mc4D4bqiNYuqgy6cHJtunjNMSbk9sKRJZoBxxBNbGAtOP20kZ6qXGitSVLvue2gV3xjIrecdQQEW
cYem9cHVPY3x7UrylpFRZiNMwWzXHJranlXoxCBUECHNBN2YBn17X2V0JWWZktkIlGVMs+CO7f7Q
6vIKYmnPntvwb0V5az8iKgvvskPBbmZcdMEsxz++/2BHOxEco504Q5YvUx8neDEx1+Rm1eiL28Yo
B1VL8yprI1qfOlVYPVvWFxTslEt7vrPNVNf7n+Mq9yUFZ+UygH8pLbQWQP+OFnNXpB8bz9rCRF1e
zdhK9e7Q6Lj7gfiq1ceKcQoUQZZ00ZXIcaCJjWQiEtKaC5Lx5Hho1bWSqqGTNEs48F60bGjfR0c1
vEDJ9KS0pey4h2qrUqTUDTUgp+B0siNJL6RF+dLLJLZf2oHNE26AfYzd4N7OJ1tYklMZ2/gPfUu3
Pdlmy4VR8XwwfdSGjGU6/bjUMdYOx2HrG6cFiASIKv5OW9e2dCnoeXN/OwprOhf0E2NfoGnGm6yR
7eeEwti0YPyTXYYFYlSvuL4WxZC3yRuUHcllOfdwIswVBqj4Gc9BGwfsIc/k59JJYg95j2qGfR/K
8sQ7IhZk2wb0vo9/Y5ppfPL2QASXnAxSbWlILrqKWfM6CaD5sPOxYR/yetFIAza0phikL9Ud8hLl
xxKlnkCBjLzOvhQ8LNH49CZBdHmJlfg1lgNV0gsfOSGmp9UnmzkewmLokhDUdhmHb4MpvtD7AXhF
GgnkNja+xkD3quE/ZQ1RbxJwanZEu7XGohyTK5YlIMQ/ho+G+LMcVlwDYG0TkdExFFpk2CIZdiCM
ssYq25y5FsEJWID3tGk21xlIftJq0qJbT3PUEjgeQ6R9w3XdXFEdqB1v2EtwOzAE12KTdUR5McLv
99z8BRvZqlxZNEzx+b2eSW7yo6jEPQekTMiVlDng+xequch1wyJ6fNFUriLL4ZP8sSJ+LUwkj4+m
rfpaSh4IqzsE44qHMUlIkarhE5C4Eh60pZu8LMeuw4rGUiZ2PP9xgRMUCHr//5gueYV3Kmw2nE7m
GrLDwvqFcZpM9EiDjLSQFIGhTSUQ0kMn+NdO3LSvSmnCPbnm6rimmnGHIz5wqZU1qWQ4enm4s+fq
K7uzoA6qEyLLHzOleiPBL7C4HTBkU+EizL36wt+s/i5OIxsODQYiFZsLz+u6DcIxHQeQLfFw/BR3
EOh0+OHmpNonpc3XU0oOudHqWvO1CGBrgMfD28hF9nR5nEEq+0O+/iuVwlXphdrPfmoqawkZLoGz
cFkr0n8DdyMjJUYNDr7QFcqzhykC3Xdw56CyHeJzqit7wcB4AzRHkyZmUJnW8B3rB403LWmq2spi
/UCgxFftREm6SKfoDMJbV5loPTGchldX1dZaLI+bikO0P8x9HGc7yE81Me00QsskmMKBFCZ4SXty
SySVYuHlJT88TEeIG6+xGKMudbEQT3Y/OdkMzGE8SH7jNTA2vmqG04ut0qLwzs2XzH7ibKdIBHew
2+Cb0mYDNeYx3ULZWaeTSaYaSWlvoHbi6kziAQGjI3cB6KHmvu0+gEtgn/4fkGwpbVBoByFES59H
Ug7fkw9Np9f1jKRqeCcrhm8Iq/lEfHvvyZkNDFhsMZsJ93Ot6YQdLKveagidPZXs8CFgN9yR++ha
VxyDJFmYwO4gNrE/56cYuFqxn/yZGl0eVTr+66sk7Q90bU9Ywv+naBG6r7M4QKyG/mrEzM090vA8
Bf+QuIry5xvC76qBOSmVSVeJ4rCCARNsUSnLwLyPdhzE0/rtp5wOOS/+aqvDaErAp7DiC/mKBcfc
4mc6LjHigtIU34fn/HW4oSvTR8OdvvVNiYNSuhJueUup8pbSbTdjk3MhX8yikndQ+pKDjDUSL5ID
ZZAa5iptH96M89HOizm63B+9ZDC501nIniZPpUb4KJlomOURe6RGk5FoF3YkAqEXnR3qBF2C2qkN
rQuqt4/ulMusodUPc8spSfoGeSI3IQa3N2XjWxmla9CsXCC2RpLBwA/ko6R/a5QTzjk8GlzW0ufR
ckhQZSxZsLBQA72nxXtUflLGY1XdwCoPK2SclTZS55XVkq+cVnK7tJAkRBvIXRsKtQ1n3HAJFZev
lbOvCC9OsAhncr7hxPt8KbENbarvwbod1a3WnNlEDoL24mJjqHJ+IvwZQ/L9//b4FqCw8q/FyAR9
GWaKTvpW1t2fGBzdwQ4Ac/npEELDamhf/Lzg44/+6EPQYB15QfN72TIGYLJN0e74pVCByjWb/yPY
XsaACpBaXak+NoKpI8lwXlFRcFB6nESiusrJX+E6aqpYtppIILUH+KqqQIZ12mWYx6uJn8jtd9zC
/asDZckP4bAKXl4ragFsmSfClgu1y+BI2F2OoFBD/0HfbX6+J0R26LSqhCZzX1AQ5bASyCkJ8Oh4
2LKjJI3Vk/gO4p0Vv3QmfXX0L9NvjJ4hCmBhK2A/HCUW1Q6hyyrKxVPr3CLFQSrQONTLBFAfhi+V
kwHAaCy+1LR9/f+dAaJU9rrU1iBGV8LiHmYjj6uwk5vJc1Xyv2sYnaXfjEHwcSHIGeqxqACrF9pp
Wq4Oh5LCiowSD2zb4PJisUx5Rv7a2GFk9/VBkNlaeVsRflEPd/DxWCjpxRmB95eGB250xiTohNN9
1REXldVu0/rfcz2N/Mv/ol5h4QCfN+He4u2obAOmyAHD7dlbfqlcEeKEXvz7suL9zKmAtuK1w4Uo
unBlz3TTwARRl+MNFrBRDYSOxpX6TPsRxwP/pOds7+xIiokUDDx9cdqOsCL25bwR7y+zAtlLwAU1
Wjz1AWziRAiW/DmBfGIGXCqNABqXOzg+XPUNcyUWCva/3t1Mknw4ykgPMR9xhNbbtEHUKFZbwf6J
hgkybkxYdFXOLEtyIuSaUYTYTH4BLmFeObZkGEX5WZMD3pQKOYvbjZEBv/S/h0IOfMGLXz4E3mlN
K+wl76uXKPFN7qdbA1+JK2obsuPW8d5pKQSX6ux7wFaYzUkoTNsXujUnecE3RnNor7G+Kv6opgFw
PomlVo85QRDY6P6tx0mJPAA31m1hWs/sPFLmFxYbiIpJhTyESmKSrW/q2FQ2APcWYGG5+J2WRrCM
bX/417/v2NdSpRpP24wUHAPruKTme/iJcr+EWa68Et1fEtrVFz4VSBNe+Jb9jt17csWgenHJHgrV
5tVY0tt18tKVlfQL2mYbZRli9sRIyCWVP++a6BB1OTvDL5GLHdrhcFbImsS6Dw1n7xT+Mc+nUy2g
IYjwWmRBqJf02K89F4xttGTV2nV1UNKOgwkqbPZUI3V+vaLY8LcUoDjsMX/MakdE0C/T0NkChbj0
ZP1V6ManCKGZc3JQfTAHEwdSMLEUWHyles6U3Cf6ighOTi5zLeqGy9TKA88BaH6YT2ary8JhAMFf
v9+rpeGyp4qS4pb3HjODgpzzblHqYg1HhQC0Dzii5FByvkom03/wiQYY8vxIwr+axxxUeQOWapo9
IGo7EB1NAJSIAGycpxBNk3CYGk+X6Y19soJXGdmQy/d9kUvuj/lQNWiy9HGtO5wPqm1Ls+G0vE+D
EdOhgJk90r0fz3kMv+1uijYAPYFtVJWDUH0HXZlRQ+tRT4y2HF0YG/6k97+ZLNcbWp7TWOHJtkzv
A6I6tE9SknlyEVGuylrPN5PwFBqYD2NhnxPGy8ZxdJjVGFteV2Nk/WeEHU/j1kCwaesFmAfHlabr
M97PxtRGeRdbQhYmuSCk/QiyJIyVS8Udce8pzKDlO8FNCK03oFjFk/n2QaKtL58UCwLAszkB2ijC
ZEfGmsLEYSlGaOtJMgTbWr+6XQpESIF15XEO6WvPiC4KB3fNGNkFEFvbtiyp79M3lP3DDfXiXn8M
oRsQT/Vo0OWpWIPo+moCx4ZMgthxcX7cLSIbUMoMjz42Vy8AfT5DratGsq6OtblbjbSN/LZ76vz+
jO7gDu8jE6b2id0kSye6Lmpfny1rPBqk75tm1vLyMOrr3ZUNWvRhIw0Lnn6RDmLacYKInrKy8nGX
Q8h9e9iZA7S13UacSgQmI3TamtZ9WBngUwDQbDKSCZQDrETdt9ZrVEhU5Jo6uvnpn2yhXrxl507y
FwQnmmHFWZ5mx/ATzjc0xzd8WEzyN0KHzJ0UYalS/IksGEDrZBq7SL39Xhkiqz2cD6XlALGT9pUK
NpFtks0kXhQCLRSf4StE8TKNu0qY2d4fnlBDkPZVs3BcNgwHONffi05xrwLiEqMdXdShIBblFdBV
8j9T6B/qrRlaIvpXyKyjT/mi6+wilo1gczk35tyde5PVqo7z96B7rEZWdk7hilaJzKL/tMtNF8SR
DjXL0+m46a7VHu+6RuqoWD9LCYHiUBFuGZZ1AnC2FHW9fkhsiH4+u8eynczte/edvTHE2/dRdobc
DDs1bvUXXhLYtTDEYQ+N9HoaRm8lLPlVACzGZLK+OhwEPwAunmnFCUPN056jtsZjK1xpqVdc9I2+
2utjjVsm+h/Oj+NTv41p2kqB7qdREzVsG83TRXHKXpBQGGL5nd+X0gdECp3j0603T/XhtvhnuIbI
Jau0MHzq5O5RkwL2gJbWqKot2cTmm57+yF/+jRpZeI70uFxklQLqj28sRgFX1hNN0QOacglU0C53
UaOSfu5Q5sQhYMc89Wg3p+aCl+2uIuswqWNQBrShUp6zhBDMUE2KXhI2KyBrjci0xjsgfX1+QbVD
8sTraTg/wMhokNCaEpGPPv2YV4CBxL0bdAS8kyk1yHyveUA/TKCLdDTWpTtHUBF/WHcc8nwgfqOY
IGSsak09BcaxtND+SRWxsypMc2hpZVp5FJAqEqCrAWzz+ZlBZsh91xxPdM8O1X1DR0zSFhbamHlf
jSmYl+WEf5bADXMD2Ee7S7ZZ5uDuf/CJRzV3Thqv1dEFj+8o8z0aP15IlnrQjg//zRm7qYUID0x8
wKF0GCg0RbEDySVg1ETRXS1NDZb4WQiwpPZSgJA1gXRWu+bcbQCzktV47OiE4tEx7Kx03bd8Jgcs
RCamuoqF7h/qnzzpLuEdYe/tR0YknU61TRJ53RSNDaBIO4S9ziB4by4RtAgU6wSP2tSBGPSEJcBG
IkTC7hO9n+kE3pzjBA4wsrvxe1wP5R4iSflp5vQHUuMut7ft0AjZzcaCwo3Zd9LUYdsQXw0DGi/4
gBR3Exp4TWzGshfJs3Et3hkxwutkIgZJHZ+ZGnGRe2jM+PUTzXNbkptX9iMqkf6JGon3MhVAU4Mv
X0EcFAH7cldq4B+D1FyR/B8fq4OHk6QRcIJhUihS4Bh4LLBGmm5VvNSBWj8D0LPO6y7H6mvsGK6V
Ps5MwPIKmvPrhYqgfrhWQ7l1mWlh38bOOcMjveaESQbeLPSFK8Y92zQfPcBO2wLZYvRDWWeEP+l4
8ivmptz6ASf7EoCFCJXfdeKBddvFmP2IEeHvyIW/qkb6Zl+1elylQ+1+fYGupSLTzqBc0CJLpgAc
AG7CU0QbQ3fA5mvF4K3UbYwyyT94OaLoGoJhPpoeoUIk4xLTiGgd7RzdY6Gf4hmg5d+rysfjBR9b
9Uy/5MFJDVfj+12DvWKvzF2q0G8RCCemsvCoJU/Bv3I6xJ+A3AC/GvWuBebjQrqU4Xd/fLuzURsT
ggScJnf/Ih7XsTDTvos2UWImntLqcrJpmLhcfkOW+aXqmmTUS2v8+53PNfEPx8iR3qe77o20eSgR
dre3wEgisT/gKpc8bv+MiapPL6qdryCBYEdmRA/KCByE2SlTBlMsChAo88/2/LKaZVD0VDi1xKPu
FHexh2QHkdNLvZX897KxrkmWslHpGU/mroU0LPqDr/wGXS3cXI4uilf1uj1cE+RzYXR/sk5bROOz
J9l2z0OL0UgSPQvHzmf62yzajGaYW9WbiC+0w9hJXTs2Hol9n8gY+/1N1WA/fMBHV+t081OAcTSh
wAmk1wN0D7pee2uNw4reTQ9XIoSrSMxLzzRcNrmSFImDTSzfZ4CIyT9gfwl3jaOg82JK13uc+3Wz
73wNXCXzEf6fwCoMQnpccq+fluCOuGz2eJCUSx48c8rxxTOokkGrtwporBHiv+EsHy42REJ185c+
68ZBUMvKs7Q7QzJO3zjy5OXPQL/bg93wALRg+vL9GU69/MRptarix7pyFTh4NHS9G7Aitcb3q4Ha
l/XeGfL4ccvSZBTNG4w4G49EaIIpQeEI5wcUPPE7cOn2z8GFy9HYkVj7ryFWNN8ToFYiQ4LvUp7Z
LTAD95Fg/70vUEsxKE42tAaFCCqSMeo+xLXMEMJOpOcchTYPtcS/0AGftGRS9lTh4hqXHDTTW2o2
nOcoYvzelDBI7kaZd1C6ByCf/Bl2m0neLA29fZr6pD8uX0T6Q2XLYZiGpXUYds4KG3AvwkqTguWq
3GPKs8nVnPIVcRK4ZWs43fxCLeS0rEXFrmmqdzaAA/p9yw8Ke8PSIPz/P7LL5868RFaEZqvKNIzx
j65DlC1Y75dRKiNv/NZ7peg8nLtakq2AUXfNRVY8pc+3N7oij0gT5KeNuczCbVXXWxZduhxYXkQ6
p8/ViKcV5xoN7geCZMdX6s3YOwpPR6pZeSXB6x+pY2/S4DiAOWuWPUVaP5uc2NsI4/ylCeVfBxgV
oPRIvcGPsucFtsK8DIFocKa8Y5zbnu6aiYdnZysAeA8G4ObaPOUkZgrrUNSyzvPrTaUHh407HKZM
UWAt5Vpw0wgQpTYIxwsdkSai4Ouj/tlf1eK5frR0/WNTUeZ07xxwkk+WO7fuiqbIOlo7DjzK5OGM
xx9jvbY+iQcEJ9Ut7Iwk/GNCxk95LTSJKJQayFQoNvU6Y21S8bFpJ7DTeyXrL+0jqUUVWpfsph8L
zJ4mF3FWP4xV0sIYfJIcUem0Yxjxja3TXkKLwklmDdMs9NNWFLNqqXJKb6MPzZIy8FV9XWKK9g8r
qchwgqTrvWR8/yHmKroxd4e8wvcFKMiRrzTCtFyHPd3CZ9cilxfLsqsOPKF8BFpud0ovniytiiBz
E9ArBMmBenRLewVH/txCNKVZdD6lAWZily4Zj06ODiOBISomvLsmk60yOnibCtyicko8HUrXgbev
oMvZOQLOmfw6DdEv94UxXmGNrCZ2eZIzUXDSW32Kr+BOq4mApftNhNU42D2KlhQLdWe9OUq3kxU3
t/mL1ZNmubASLmQk0mABE5UXQ7eFrTpO2N/eJbZ2ACnNroQQI2CKS3W5fbabPa8vwuCZzAr5pmxt
+elbUjUdmKHAgzvfwyawcBj1yfpwoi0yTQoRrcHiwCoGzH8iQF26nq6gu5mZCxkaNIa0QyO5+Wuf
qE4R4uHyVKq9/gY1poPbvro8GW9kKJThT4+EDgtCuh+3SXuJfF7vGa+ze9ZgyDzXzVPTLX/s6kGf
Arsd90rZy988pqNdMTx27NYDgEYOQd+21HCCfqbhVCjdhv7yAOyy+D77dl0saAiWuMMaJZnUYnCL
auHyCLTHGvmqOjL6s3wdH5+jKYmqQbYVoiQbcc1HxI15fGFjoa/aqDUM+SvIMuyWrlnrvBZ1xnv8
eF5jidyUK/7QvXM4nym4UqDiEI5yzWf5MYNMB0Q+b7JH76uPnX+XVu/EgyvzSqLwICzYAameiW8V
mRel9JkMg7FmRHheFpqLo7Ovo/VGDb3HsAoAJksEFxir0j2tMPjLv5y1lbK8mba7XBGcSivdESQo
R0ic9cHHU+4Q89r1Y/wzofp8yZ0Rb0Ql/3sZLZJJ5VHMW0ZpNYS/JqFS6VXCEVZqPb2gchyhhr1U
9rZeUmwc5wHkiacxULDgv77Nc9fy75EfNUNlVTnN2V/yrUhgKs1n0FDMz5OQFTl81tkS+uVjJIET
AM+sNNq5rugK2DZPkNiCgoqLO0rG+cEwReoUJ8Tf1A7ROQdEjtRgR/FSJB6+YxSdFNogBWDfTMuy
mWWGlffmhQR6yJE7iQjLG6pwC+l9dIaQS1aCmAmQ51iuao6qgPdpU/msdnrHhzGpCl+UGxXXqmc/
OAUKssbZoXJrat3eSpX2mV9dexW7hLs3lFyjwD7k/02eWULbat92J/kb9nV+CYRhxXyNwafX+nQZ
EUdVsng3SdTaxWzxcIRKW3gRZ0fj1GmM3hxhJcWmxqKv+rigffnu6lYUr+JEs20u9L5Bj4s+M2E4
xreVsfzwMTxWY0gCSA/DqjG82vG8EEjs/QsCv1FEFd4UrZMK1p75kYmNn4XumpwUcdBdUXxUugJ3
iKr0QcERI87/9Os89r3FFZ82MhTq0BFL7kKmm6+USkfMEG8+/ExCmhGPseKS1kwTbIXcJY8lHsYp
XiYE1SYmP+KRw5St8s4UseY42MBXSxSc8RnNnZLTjgXdM236yBiIO+aSyHbpurDH/8B747RvozjG
M76QweqLLZxR3rukIycpIq4O5btpadSV+K5ZyDMXqAh6YENQOLRVzrNmbLQUosiAwjLZ2R7/BOFm
s9/4plbbi3RJFZf4XnjCMlbQSluBMultxdD6quNcZgM5x5IHzCa97uNOmru/CMQtbi49kexd/nma
Y9LRAyL6mc68CDUOkrSIS8ovvxZRqjmjAs06T6PZaTPPutE8KhN2STbkPjQQw9DHRPRf9rgKtShx
0/HR5z9RjlXbK9Zn+ttPxAB1a80Cmy8u+ciT9sPzXp+2czj72p7it3noFR2WsS9qj9CuEV6x6K/t
v9/hLVRaDZ8vDMV2IpkdwikdpyK1MOD8PVmgViOTAxVPdz8EqksqNre6bgW8JUYSR9QcrcOIfh6H
LBaUgae5FPeED+03LipkFY/vE8C0r+tiNt1fcnADQnjTC874snkfN59T+tsgpO/phuwnLWl6Jfzx
3hoR8ftaxQkKsbaOfc4n0vHdMaUihYMF82v2jIZR+ozTXFywgyYOFjtTN9GriZX/vu81BYPl7KZS
b25ghU4CTdn9zsepA4otLSAuNi0C/lDAgbzeTy7ZL/JP6SFC/nCR7CT29g7qV1wWoK0oH6IF3JCa
efKleYzION0lzKPGaOa3sU7TF7YwjGZ24rF6rkfhjU9ULszI2a692iplB+PUdVCM50SkoGd/Ix0t
vIOR8OHSHyRcTu7VnwiZVb/eL0iPNmIi3KyMQi9LTz6qMBe0ovWTq3HBSKOqANHs9TE88LaYjqB9
VkTqq8Mf16XuUIBKVVJWFqKDi/kSRpnzk41ojFa49shiYuFNuZCiit8irEUda99guYZFXYBD5xY2
d8rtIwEqCsB5FH2J0XHg96Oio1SCKmlQlUxI124FaT2aAc4cPTI9+Y9GwhhY/KVBt9n5+Yyx7vdm
b4RWdD8SdAfi6HlIVbN0nvSydHS8qYyRMTIF+7RMStXzSPUWUWtswTPp71ZiODIrzf541Auq9+yK
iXoyn9jf8C4+smJOzzWRLyT10qJ6g5XC8ADxdOgcxY0J+EDcqU08JCAeV6UjjQTsZfCxl6uLTixS
MSlb0C1D0jznXTHDYMq7s3+Y5zCcqBp8jZfyf+VhF5DlD9H2sNqOja7jf4vgjBVLaeWKcjXxMuX5
5Gq8NE8eWW0AYIfCSqRjI3Gemu1msUEqroLRw9zP41ycZcOMQwsYViYSakNYpBPy/Q3tf+3vsJPp
BsG3PT8hue6ISm+8LlPk0Qajsld/DzRT2xVKlR/11CQWz7m9p4/rHxo/hMhLpU16F+aPeLPuaNAX
Sy2ooZSTvSZN0N5XaQ5BZRoRxmn1gl91PzSAj+QGXmcqc+KAm7LBHDJXesURo8d3TWPf04Yr/P6b
Wo/NsUCmamNA8p7fcNySAQiOmSIPcPnpLwD5SdDd7FikpHxpgB0zBB7orVELKA3cDjM06caNsXvz
cXMBajAsUPVtIHqz6RwvjVYxJSTZfridP0zwkCPC0IenfpaxudgxdxRWJKTwWmrvOWjJFkxM88A4
GcUFrrji79bEmqp9uj2QFmQXAcNx56aCuyPLT17XPBW/zZx9Rdr/fdRa3OQtoYlvLHgwC6MPCW1E
ep/eAZZ80D1unajGXGBWo1lPz/eY4Nxn4A7Yih+P+arHwsppcCeVtUFpw0EHWYOKF1L7+Gamhj7L
8hQ3fJ4Klm237xWSp1/jx6HVuKbcY303YgUCIQHf2xzdRaHVym6ITt+wE5/upuVtGj8q7obqotee
BZUgoNs7dUZ6gPZh/DUn/DkV9Y69ZQtj7v8kgR0K7PwPTMYt6/6RE6499jN810mV9XRP6iwRiDYO
0ee18l1udzvua9gP1koZzmCZD68q4IAtxy5XSK4iiHoZDaHygwQ8Wde7fcVEGbdp6mJ51kKY/hmu
edyL7Y3A3UzPB9Kz2SXH50/x0XCASlZ9CV3f7n5DVA78OdJuvJTO24vckMVdOEaMA7gaUWbhH2xB
A64c1SUYKZc1vprncaNIwKBR5ktBgIDPvVCvsKTJwNl8M0spPyD07C/IQz2u9zBq6h0I8kZhGo2V
mgs6PYA4+w8JXvO8tOOtmAEw61klCb/HuSsYEJ3OQrWscMvbSmmkRnnEKg7OWkvmwZnv4iTBzIOu
IfnCMQcXadmM2DqYfilO4qYegNI4gPML9eUXGA3jhJWq82u9l3rd8WH6lbNlSMcMG9xqZuDqJR9I
LxcfwwRN192S8nKsUPYfY6aLQ6F39lxagZGTSqUZLBC4Fzyau+OR+GoI8LPOJso46RBwWDgIPVfa
Ixoivoc1T9kiEJsbZcEiR9BhC8Hlb3aeLQwl108OK1/D1LKGrJG9q9PJJph72meMRLMrJ21RO5oE
eqYUuQ8b8Pgtz8ep705dl9YmFMYpzyybpmPUSyCKIW9zNxAMBOpu7EUxE6rDYsE5RHF4JzPpii+x
nc7A8EfDOi0WvkTfk3/bMpbzd7W4U/4IMjDYooQaRhE2gATvxi0MCTo9IvYv8lvWgTc2wdRLI8L/
SYQ696XkBHaM/gVo0UdiazQ5LrVEXd+HeA1BjQiEcwWMjTMBYiFoe8xZb0NIdZAvwA488rLPKKe8
TeoeY9vfHaS5bAfb00CDbRSFFVj4Z1/PaNpd3RIQWJ+62LXRLjp82aV2LK28NQUMOi0Vof3hPxEd
mERU14+1iFUvsOmcocsOy6nQ82w/1uK39vsdT/5Sui17DDy/bBTfi3xxsc3Z4h5OC1WQKKSdVKUX
G3tL51FceZmGyZRRE53/ij3Cuf99d/TxxZrvf6Ttj6CviVafgVk9++EEcWxyqlk8nOgJDv0pIPPw
EUr5ljnfrAsroa+FjVzYX+SiI6fz9n03DUGQrAjGdwZg4LPsSh1GBsv3J2aAwS8Y+eCtAbDRdUpm
eFqpQ6TItC0Lm3qqT+6AVRvxV+UdTaGmF7X+RGGRmAU2ZLKTsBi+tmhI4tA2gdo721VrlG4QxKRZ
Wmdr3LdOImFHlR4dzhNrOrI/eSuffb9+mH/TbEqz7Yj3XIoNK+5z5QcWKfjpxWwBO66l3CbDzTvL
Olf5CkNlMBTHk453p0L/RymXea4ytsS9bM4j+8MRIdpLYydN8mTdfKLDBQ1g2LErgH1FtUtjqd1Q
IDuNW92jfOm6CNlIqquDeoKKNxXgSE5GVTM9TyEMOEFBd/U/Woo2mnGgjN/aE+YAFgMdUza5/fHf
y0baqeDiWRykqOiTiG3RJwy0AC8bLSHNWAMZTzSaRaF9p7UwWoLny42I+mls+db7ZzIGf3YUJb3N
EsPsej0k0a+VC832vd5H4W2kV02d6Avye6WcDjaVyqmC0dZlKhAN9/W2Au+VaZV60Zy4a2qjbTDZ
SFvGIr39GnAZg8X4KLm541EvFMnhke0Cv30u1Uyj2vVwnV5QKLkEBIHx73/fDOHk/cGs4LCFvsTy
mey/iaWJmr+LhSbu7ffZxQ/AIrCRl33FZLJG5MEN/liTGk8LureV8+p5ulf4K82qdrCYguq/CTgw
z0lz7VKwAgR0cswfeeoB3zyBRGUa89iCaP4TzyQOPvPHzvpsfBsr6aTGjPqiM6NlRt4faZY2fhsw
bSxXSFcTz9ODx6m73Uc4WBJ2mFtwTk0OSR54L03UbUmH+Cgc/PS+9HbSB1aKtZxvp3crFOXd2kch
CtEydgdSEl+oWgQR5z96JI+GUeQkeXNXDpf5DVohT9GgickQVbhgS58oDKgFxzuaBMBAEPiqB7RO
Gi4AuYST+V2PYnSkjS357SnJ550e6tDfB3Sn+BAj50LsQc3kgW11mQ8mRsRKDo01L8/kaMrxIGbk
USoR2TJfWoEEnOaSGyzm1Y6cGiC0pGZjyQfYkdt7YiANiQR4AYzIieGKEukalHMVQ9ZGHeh2IWZE
V2K9pzwoz6yM/XqNJEpSuZPoZ9hk6ViIah+zmzcGeawaj1SzYeLWFOGTavGFz8ZB6VFmQmC31wTD
LrI1NXTMXFp7hAcgKm2ldNGtLOKHZS5RfBl/X4LRHNf4wtSNnGrmeNHkKucESdAg4qaepWqdv1QN
3D8NgYEQ6rekKbVjfN8/G13mzaRfSRv68z7eA+iJ4ttqOOFkEHOI6544QyiQUJ4j3DQVobXuVKLX
bnhpUVjhY8XcR+jCz+ZpVF80L7TJhnyYuM2K6ld+7mfDVjOGQlZlRC3XF9P7Nq5DebuMf8ypVeCb
xNyqrOWPWb06k/gI1ztdAUgg9y3kkZx5IEcq2LDei/CkZBLCh0sBfAkT3nHYvCBl5p1UJ88O7Wba
QKsRhlpVsruWs/wF62jSzY/5GQqnIvkfXPeWZrfDm5HbZctWyqPQURpAwAhX6aRU4GpUWUgIe1aW
FiWmrpQ06f5aV/fL65n6cAAmmQq/4Lb5P1GUwrvgzBrOFWtD0gOAd8DG+DikpjYv5W2AerWIrFii
varriWlwiyDL/BrzCpRusZagXljo3UhFOAeqQTs4TrMWXfxOSzeDoIgbgckHdd+ICEY9dYjpshPs
YF+mQXevcXdoUdfb2on5Mb6XS/bkxHe2SSHhTaM/kd7lLCN69uORj4V8niE/JfD/hYCO0jKhqSa9
y72W8LbUHOEIcSec0qBYGkxr5eLpSwVtVvwN4b2myjwTYC2JEJ+uuixfq2GK/vpyG3KZ0CjRmtxn
TboHPUair7h8gwT+ilMsGy37bwjmfwbnYIGUA0Nk9w2nHv+a4a5zV4Bh0bM+nAGTIRzVoiA1zNvB
saYruQO09RwCB4tXKSX8fzpORFuiLzLCqMh02mSlPFzT6bXbZ/ueSnwoYO1b8U8MCWdOxbxqpToC
7qbV4yaUlXuqsxeJKkCjYGZ0nU2QcsWlCjPRfRCVDb0+ZD7nccKNsQTcb+JWcGRhRg+XzlaYqgKC
I+fnjaLAzHN6AxkOTX5uS0e1RsEzjqKqm8xSu5o3MauUldyMHWSWZLdG79BLvUmFELGNqNQl61hN
GzmEiN5f5oYd/qFUEzw7b/E0PXcbc2FOIYjSJkmwgepWxAo2mLhmFClZM4f/H8d0Turc+4HIg+Fx
7E+9PDLoyT+SG6Ekp3+KT0E9rv8cwG26G2b12rqu1a4upuBDjDbvd2eKshmPqkvtfCjtLGzh9W1+
243jzLcAk6ZjCRWCU4dhWKrC4zitUWpneQ069Yh2mgnSMh05wQjOnf4ePLswkj7ZnivnJOWhYxaK
A9vZ8dk0YI+o1Mw75Rmk8vyD85mbP3grKiao3gm98oeGmRXemXqelyVnkbpjKGEpfpDl7rSPNqmV
efFg3t2DpRVCnq4fknmOLVWsbQPLA1LnjAxR40NbpoC7j7leHSAwl15eYFuQ8wnlIzwxz4DDV5i+
of6/OAVHBWGc4Bd9MHtGUnfKVPFEcItrw6hojJrouFqiihf9z+nTvAnpTCHvCxOoIU+aNI9h0bvO
QWX/nHhmZQK0iHyoy8Rlc1bq/bs8Awalfvgiob6d4MOvBKHmL+HSmPXlCIf2fmNKdRooA4dOOLvw
5rcGAVEHrXN3EDHIYePGg6dcq67B/XMg+oGO6GSyrUJd9bmo8dCp80EZBmfX13h5VcOI23jrKb3r
N3Stxpk02iRiko8tx6nq2L+XXCP2DgTqou+LRBY0YBpxVWlFLCZpqPPy8nWa4VmDZTABYKimVC2B
TO7jGaDy1/d7ZFTquQ5ujKagSBmMuqjRn0E12/xjVWmmrEORFtwFqB90aoLBnHFcNLuD01d825cY
Vs0P4G2AdvsmEhLcQvHZHDjanuhHnGkfPC3b1+Y2Bu1GqtLKaJvbz+42N3EqAClFIx8wv+3T1ujw
jYxriFwEba3JIwm0YP+Ys7hwMP8NjoFFOykbEo3PZMQ36mMKjm19JVt7vH2YKVqEmXBDrXXGzRLj
YrYBJU+kAU10Eeq2HybzkF/ST3OEDO2y+1xHb5Z9L04py66/JRBdd8HfFRh8SuZaX97vAI87ik/B
On/YOJQHwBqptgbQlv6CTzuoXKYV+hgWCTQnGhoTEXQTSRh9F++uCd5GcLG4YjSSquVTmRbryrFo
hheQ4tmJw9YX7p6uppsvtSUzZeEvKPQdfe1wRg6BbIe/Boy1XAHJf3pLlTt7Q7TjonAhipGazf2u
g9DSx8vImWE8C+vtw0Y5TZBGoXW8vFuAD3N4YkqB2FXLQe2LaJ5RWcdb/7kBEAna5CqS4It/nMCl
cOOr+8p5pNW5WYvqTsfoRZcclSsXALugruYt7dyv5hTmX+zPG1OtUC/XSA+5GzvAZjIj+FVFsdyq
4Ml+mx010WUVln2Jo/2gJnIhPE7kEnqDe1eS+tL4jtC2iyukwUtSz+cDirpFaTBaoJOU/ay4Opg4
w2MBNeS4mb5kpDXaagQKwbpZDRy0KSDXZNYWp9xnneveLY7lvA/ix2S72VNbuPgr24Hbcg3bR2EL
7/n311MJBC/bxR5CWR7uiJ4YIVJPfczjqxZnko5AoKkiNnBAaVIJSk2a5td5Ufvse1RRpeJbEp7/
8Q5gqxEd1AjEHyhGVmbVHKajbOHky6CeSGe9yNQmaIR6lxmm7cRzMPjgurDZBvmhm/ProZYC6Eyu
5085H2CjKEn4n026A7abFd7biBjpxgbiKONLmDiFKIcTWWmGIDRPfx0hb0x+ZzGd0uJL84fmJT8/
7OJFOzmImC71efWNOjzP5mvWlhz5Ge41U+Pr6E4V7V08ml8vb2jdpTpirLIRhrFuzEsH2OSseRNm
g0ckRtCR9N3S2AbT6FciUzxjt3uf9uRNRVIFNvRLTxZ3IF0zUBUlYRidq6kLb8+dT1SAQhwrS/00
rQKrAfoPRe0itDxAwVebjuy9Wx1ejh5JiNhrTXHZAsrwhdvEXbHdoqjaveJQS2W7QAVfNWVqnpmE
U9O8uxbCPfxV48RtFekHabhuDPdarUhs2AHza8edEhn8jv+JIU7tYeycutG7U24hJDJrwTtaPy7e
PkA2PxbfvJdV7PcP+8iXaTR2bUsYJYPE/g2Wv6QYSfMntbfI8PeiL7NvGlUBS1MMDLVUBVwz08P/
dcRcBDFrKnGp0/jjw9wR5/k0lgRtWgtKB8XoUYTBFZTcUNWED2vTOMuhMgr7vfT4HdenYiL0J0BO
nsGBfuhxhKeJcbnNrgf4RjyMvCswaoi8ONRNdCdW2y45sFaMjmoctVcF+eScb6anYIkIvfOjLJv3
zCbG1lTz/QsGmdJXFDyiVI42DyvIYsM+UC8P6fHqCJDCQu38uUd1BMosOa+v0rMXI74p1fHPtnMt
lefP6DdxNeaoP0BiVJP3AoS65CdslYfTstSwWEuutyvEgcJaXMlVmDLVt5rA3CBax6UIEZ6uwj1R
RdPnO2eWav2kBt9XkwUnVqoMIK3lXz60lCfVaEwLrSLypL4Sdbc/HmZCheV6mvPqD1DdXnXvr8Zk
pai+uwUVtQbTkDwUUvY9dlxOFHwqFn2uODomTAFtCCtsgmgH8j5KePpMorppTXYWreptsoyNyVGg
pxSuhosBUXiHuK+zm+LQV1LoiCsM3mmum8M3rP81JrMK//o/BsF8W7nHf8sHcDHaBZTzeReIa/ER
Blv8n9Se8bc3bwP81ktEtW2O9/BHZkoOTS9oa0z0/ezSNnQe7PbuTL9mdk6hxzTvO0khdn6SHiOY
CwJcRvu1h8J7TmFTFIybl/2c3+H3CKU8JPxnZwaKmXNHo9Gq8+eenj0ME4HozlXXQZ8oBy1xOkdL
GJpBw6YqMDamjhUL6C3L8RMxefSni7tAJEjWu1hK9lD7ExyS117hTcgMUN4kdr5/vnb3BlBmQ12k
5oEcZL4XXNmAN3T25Hjh9mxwM6reQKR740Q4E6F7WTq0ARhz394QtYXwwcgB+axVxqPCbR0D7aF8
65E+tlGzWJDqVZnlhLBKidK32e8KEbhD/cqQVjv84AS5ULBsoyS9X6FtkDZoYbwd662arlwQUzEK
NPyEaQwWwbT/prtAXts7Ag5j/tyQP33IRe7Ov7X41FYsGjKdaxh8hd6b17iZhaXvdSlIukaVnklZ
l0SbII0DDPjNrOCqWc6LWkIg6eT2Qho5PpYnFYvQssGa5mZ0acmOz58NlYjRfARGb9DoxTX6txcu
6KL/QL8W1OWyw9YPOn+++JM8OjXWy82lnOKfe1M1DAr8A0NEtJXxEXygUpVUkWr1OUx3jhGtg5Tz
iI1Ie8gxjP1SiDnlxCcvsvK/bp7N6Y2tQO4Z3B84X18HVNj+OsMviBvXEkfRW5gwdTRZDZjCl832
Kw4L1JzaeqSopTfImtifTYydw3VM2qwDuTgtlqz0k2g+2whdeFTVOrIo8HfSv8cXCKHM6NX3clws
gNPUVyfP4lQ+JqlYFKlmwPpoSWTo89bxZmYmsEPi42B8yfuZtXqhJ67vdR0+vEcQfaBZiS3Lg8Gx
h6/fxSLcLLCvn+mogzxA6o52MNcHP0BxU/witPfNxM3IXlJaekouSIkDFEQ3EsVk2PeiQiMZ4ieV
rP4HWyY0xG9Ei8HdxoYPClf+fqkzuuzhzTIpYgvtmjyIt+W/P97oDBHA3ntQhOgeED46/5KCp1Tr
+hiiME/zgbW1tqOpieZdBNwofpYyzgz3swmhaNYK+UDqOR3CvddfO0vhg7R12uk4JxCE9x/YI7C0
drL79ZcaAZw2/afc1IyidjoTPNLfU5S4riAIHiw04ybf4XZQCA+gH13YHn/Qzn7gd6J2SMPz7pw5
AVojlzg8DDOpFsE0NBi082COJ9gqKK8VlXGR78Nt3G6u4afYazQYzoUYSeeszN1z0WXl+RokUtBd
tvnf4REgnHWDTUWZa44NgkAQK0aYEse6r57VIb8qTRvXPgQFfeIcDkt8Fnkdazr7J0esar3aJD/f
GyUOSXwjgcMhi/P5ikC/s76eJkfIGA7TMQSChy8C8iSIACWbSc5IenBgcNy7rFoxXkboCRyy6s5T
XuH1IKB0CDyH7VkCFHefEOfv2vFDIPAPythAaZY9LA1XphrfNE9ujSoDWWeYztY7J98MAy2+Z6lC
EQVD7cvRBE93D1Y1GmQA8RGA7bFElyiUtvuIyQBcfaFge2Y/qmVAXdmVr/zSFaIuX3+audmuvWND
+Wi7NwP8RhdSuNDgYolFo4+KvVm33DZcdB+V2u6QhUuUxZSFxWnz2CASJDKPkmtY0K0mu7e61mr3
ZZc8qgOs3M3XstgLCkFOWxxMZ82OkZlCDIgC9OP32ew0/ON4k5TGzQ04q3HgTF0iVYrm6W+xM7EW
4ndrK2RzLK0BwdJ5ROzZIUn8wGnXAs9pntKM56U8bNeI00H8gL471Lc/JE0j7zTLcjFRvmU3KS3I
6kRSxm2I2ITM6WiurAUyrYyFg5jSu+bYE8shSZ8W3EWkYl59L7oqxAVKCCiWeJP2gfCsZNM2LY09
e5urSzyHqkDcF9Ydj/zsMhRo9pd3QQLVm7mnbqXlw3PVAeqFfCGEDkzNUor9K/Z/FZ/tMcAVAsj6
v1bcoGe/Ah8FTfgBuJd2LBgEMnMIoZ4p7+LNUxetoFBZ6+FPapKl/s3dqn5uUskN9sg8S1M2Kcxz
3JhO6cOXP6R+URheIcpU/gLryiKQ2omJWcA8GSMcW6bYeX14yMqtbH7h/HuKwA8arjlI26urXd/s
Jtxy4hi+prKkzmbb4OS4M0mglSJHbK4jm9ZQ02vtsyoaBMV7m+w4XpWi6XCOnthr0YnySba6jgEf
p0mrIO+xU+h+ROC3JuYk0SLBnf1wsd8r+V8EYHlfzEwGYpmRRGEOPccMI1P7/2SyJuCi+5CrGZk6
bnisj+0gh7S41JMoNCoMBka99J28DL5AC+sEyL74BtXkCrgizdkd7M3uOrNf5ihFugpX9W+oLZBa
BXfi/FSNkjIx672oO+FAft19toNOgeKcpHObbaGjtA2lgTSteQlgCZJ4FOEsGHqUOlPgBwvYgPS6
ntRVAaQX3f9KQhczRhxE7lmMMZyuditiVyYQW0a2RWxAUrmxjmVI72JUEfM1UZFnqFrQHsV1R5iZ
DyckQ2cfVI6K5q1WWkbG6R9ocVi0a/6ICQaSGPV1RqGuuopeIcCQM6MGWX8uycBpbes6LmttAc3c
nHX3uYrbqtIBjZ8XqNU0WYXRBpRjGKx4f79vnnMtseAMu9CUVYLDzxUTz/lQLG0GYn3UjLFmpseC
wkmNlcwn53s5ynUBYL+UdC98Z9hzTwXzr4mgfYLSTN5/E1hJCdut+xTQvUBTep41FHJe3/FP8AAc
UgAbjryOCu+30WGX4zwOxDw8pbEvfm454pahUWcKKVtkf/E1fL77pnzjBuyi9vl2EJw0tJBEOtw8
6d0+qjLZyww97O/hgybf9dFwDJoa+IcuFTxMA04VKZKJP1ub+G8fpomky9/N6vGhhKbBgw3S7CV5
0NrwjQxipFLJWYbuoD5o9Nc7N0WAHLyEqWMFGP4BRcuzzk+0NKLPVbXBYtJn+1NBVG6yTq68/X7j
dtaXse9sNGUTxk2wa0VttQ5iCxm+p474p7ak/V4qTGOdQEsaKs9xoipar0mOTx+HbhYPRex3vAt4
yOunArMOFobnbMmkLGXvx2Qaj96VJaQudo4GuVTn6rDLa1qFHApY4eO0vrf26SQSl9zbq7yI+LUe
C/Vw3G4VDMdQZ8wMrJsjy8Gj84W52EEJ03GI43hk/eRdSGz37wxmgxYzCN+xhZQ4xIwyMHCsDwpO
MmM6BI/TGWX7EZ7H+rMylTe1CVPrCDGod6BZ1uQOIqm4LqQaGkFs0miu1ujUtAY5RbsNJuQKOKve
ARWylV8VIrbBU2ACvtNfAYPy1BP25TqrJGAVFJ4sjBUx0jaxKWoGY3JAGRw0V0gfPvafkhWRmazy
iHBRgyLqMBCnqDGQlI7XNWjf5DYpLgAntBvnMgMoNb/ia4i4HZIAADJvDFSyFokQxOJt8DBPtht3
M74nvHtd6uoYj00ySlRvmg0Hj4hILhlYr7ecKte3X+4tgU6c/5sLeMtT3NboVY6vVhRV+NwOZCuU
nJPgqfvFVR66wcBosC6YeVhL35v4RRdmzsp9CNKh/Y7U9EF2BrG3rn2Dk15jImzJEtvg4T945hes
tf9VKmSIV6wZWI2cZHwip6ceUrXBvuRqWN76F2bEvEteOJrQTV+gyT+tYm5CpouBOGLRvP5CKm0z
7iGoZMtmWwZfGKVnt2X9xsfdYvC9B8xpjv7fROITQXFoIqX2UU4p/L3k8YBWdfEbBda1p6H1f6ck
obPIkSdg1elSIg+/3X0akEvAD6XKbuDk/qjKv7R5CXWIoEdLkOrg/XQcbpseu+FVEOYgucD72KKr
k8FUdso085J6D+9+jasVcipjOLG9HTky5WAecpbk59FKAwvKNIldbiFLEgGsVmGX+Wz9Y8qlM7ek
xmb8Eb17tfUYjuomYlZs4h5F+WYDgj6waYVKvE1U6d0hofiT8Tt2O2nDLczBlVlfaDYMOA2lpyZI
j05YVVrcRhIl2LaR2cJ+hp9IeLgzY8mfpoqYupgaGCB9D6OdSvi19BaeLfGCr8KbIh4i1Ow519HJ
ERswsgCpTxy4cGn18e4wkHxGOlrJcXCtniwetfkxhvUcP5hA0J76QQ3KL8q6yeXpI9+ohZvf8fsi
1EArtB7yvU9WR+W0s3w/CVqfD1DPmx4M5l9nyrgxWQq8MSOavBUfYsqdA7b4GyMrldz2wThM2iSF
7aJWWk46+MqPYKoH3K+Xj4QL9gFGrYFcmEFMGR+IJhztGhsccqxMHmjEwQAWiI0aNJkFPexWr9Vd
mEA1LTiQtNLLTD6cLL/dfKeDf7xqTuwO+Tc8cdCYMTxMvpIxGnlmc0pFs0wsVTtpntheL0wTlkZD
OEha7J8pm/nS3Rkm/s9Cq1C+zUihnY68m7xAJ/en7DaFGNUEygNX04CWJGFqhIwcLubsmzoRBK9+
+V0GmgDh3i5MR0oQ+L65n4Yafb/3UqQ2zKOoJQMmhseL8DW8wL0Cja7cF1zTiBGCz0968n4dA52b
DVAe8iS7SfhS3kMKLXwChjIYcQYCi6FG05wRi4LxmqpTjrn/jQR98IKCsbM/rgHuRvTUh3zPTB8x
/acCJaQT2P+BdtmhbSjtFJkTPU4dmVF8J1/7rEl+6VGvCOM0x/0166v8+7TbRMiukVqO2jHP8faC
62vpmkziZ27bA3/CZ+L3e2DxBw6ZEGsrR11nbR89r3b4Giqm8b7jO6GAw+sUCrkwG/sQCBOd2bYp
OAXxTsI4IjPJc6fvH/vI8bjlhrZfev7lGkqrZkH+KJ4l2f+2aOvsP4Nmywpj0f92C+PGO2ifmQXA
VB5jKaNxUzjV8cTboU0G0830FKUiPgB9y2LeBXmeP6e3pV+UdPCS7yZBJOW0Dwn1aXNrBtjOLFWm
gAdaNxsJLLMfvaFRux1NHyFRbRvpCQOFONAhH27sqn9Cpi5RdWgQUekiwA3dUzdbdbNmuAOe7HTw
PDq9IN6UF+IuBW4zciT7q/YEnPGVVkm2iza4satYIMnaJ3Z/SQ8hRWDzgLp65rhntw6BxE2qv2mV
ridt1kezW7qFDzNhWdZzgRQ5D10PKocHqnbaievxHNcEgJ32UZaKB6uDCnRt6I7a8n0c1YMv4jxH
kXx2B8I7e4iXkeMIV5cTtqRwg6oNGz1zWmIrjpIZiXvhEBzDF5rA5SuVNPEJ0D4CkgdVF29DNtJI
RPzxduBba2xMYKo27A/THK6Q4qJeqkZvacRsOt7DmAczDdyBBPwV1n/EVn+TCV6vOEQDtjRv+zg3
e79REAWSoe0nRCGURxyFeiiGCR5Sn/fhVpNOTx9io04r/kkGX2lj+98PkG6oNb+npGWvwroA+Ov8
OMmmxdPPi//z6EPRlgZjJzBAj/T14Xyb5CC6oFCtRvh+qySo2DDecOglDdOjHLrbAPBOYlBRXdI/
5OH5G549hazIY6vWKWC/db+SZh8f5nzBoCFQHrr1gxf6G3Z2to1oekYKKpIXzqryHWME2g9kXNZ2
BJ+Dm74gZpBQz9oOKI6IbtfANcmN/D33bQ1mSjYg4U/q3iO2T7JhEnpf1TipqJzQfWPrb42OzQwj
U1DCBa1QYS9DLCLQ+vn4w9vknVRgDhnbD3mzNY2iuXCqKQH6BJYBbGmxC2TSPyh9N7Lg5nOZcV0S
vW7Wz/m698nNY3M4EkC8+n26vD7E3H8QPMtfy9UVsO7vKmTITwBc1nO5ncdD5MKzr0cZF16IGmcg
VjdjWPA7P7cnrogxWqsVS//+A8VwtlGN91xcvBn+GQyuA2egSAYcxbbnBHIpSYp51T5/0DVAZHO9
WScjPjp/uIB2conoY/MnUhT/ZZgAOYm8rm5uOi5PdWf1q4449ER0xN6gf70r9nsu1aSRAmMsELS9
ShnElQtCoReUwd/FyvyTeXTIZf06D+pf1ETgXxQ9WZdjFMqY5j0lc1I03UeG2Ta/9LCPS6dgqntC
/S4Kpq9+zZTYM4wx3MhBMRqsU6VXvBXjJmaez/JEllWOFYBs1+FAVrj/F3KXbWBnUiPCo0j9qGCG
Pi9FhkYwXKpbbQqYevKjdBh6+wuL92qya1PFvskqXnIxhuQD097Ri2GiqafPwYT6Tphl55W+mtNP
xQ3XK+7gQ4uDrXWkDQjQ+2yLZx0UEe+UVGEg9pr8MNpbyWC7Dej8JedvoOjaicaUOcIC65C9F3BZ
5ENTnZ+n5FR9Vz4fkdKxpvWabWa3u+mdZFw8Ipqx5UncXMyq3+tuO2GbQAO4obv3NiTfAJIF6fVE
u81shROAwzRiS5wtzT+kV6gT7RJpHnIcrTZfZDd96xldJg/uYRFoR1adVrP91u/ARKLwoaHnI4rq
/O2ntUV2QRcEC+PLH3rJh4J9wxNsYMoVrJ3i4+wrEWoevtcmTBY4yayy09vI8YYsVjv9SpwzwBql
iSgSzFhtg6pG7r424Fp7I8ho2+AbqJkvXaWjQuLYe+ROcZfPp1ZQpOwolZ09LD3ITXW/0xT1EUTD
Cii16nh8NasZgg0Z+eqSoMX2z7lUxLUgmV1y9NeHQ+FBzix418eW2MpAmu6g4WRIsmD5JVYGN8cw
HLsUa4SDRsxRXrWhrXHW0sKn23axFrYbtkXlH8GHmDDlF/e0YA7pJN/PmZyufcq/15sqdjcJxA73
XirAH8Vd/S0uRLfIeKn4xIkPl6R3tG5aOm/n8krc3UZ3GA8ewUbS4drvX3Tg/9k9ZC99TR4rQE91
Hdk8i6YAzjBdeay42cR6bWmA9YfteyVYcPDFQ2YoLT8/zuswYLefNP2vKlnAh9+OucPgKD7b5oes
rLbfXLDpQsPgZABDsbT3LOD33m/u8X0zI36Zt2LVJaVebP2HF91H73tqlBw6JmWXejQ5DKhHk6kr
Gu9BjLixu6sLScKqzBgmaoJtZ30+hKsemknXHNYL+/6FETl45Zlez37yuMIgj3BhLnQVH5bC+5mV
pVfRaFwRSQstm6Wr9fRh7KaGUvCoUqFv19ZYXLSJ2P9a5b4vbTNlgo7WosF39L/R6GOOgHJoWx/i
Of4zu1ntCa08ABWIJBcKclkyubk+QqakA1eX6f2d2I4v9gpP/zqqTkx8dlvJHn4a2b3KiaBhSVKN
5pbj7zm5MNGkdpFTHULNg4myTidfXk836SI3/rpE/E/xc1kIF9kN9ktIuhCFKUMCEtrDHnG4nE3w
kwdpjHTzWWW3WCMfrevfSp6xr1hojyJOBF4nHrp28M3yXOAcVCN98RW2fHrjMnCe/MQ0r98vc0wc
5FrMO++O6sxmBB/yHt0PbsXpShDAHRjnf61OtoT024UTGaukGNAaU1D6FCyyvMifnUV5tVp68KM3
3s0ARzCWK5gDvynesI3lGSMywdgjr+ef5vG6RLsAXPUqb3bqVp2Q5QKhMz1can2S/CM2TJrchbqc
9eID1sfj2Sw7/2Dh+IBKHcgWZ6V4AA6HQ2F4iWBe5REqCezpnpYnn3NhhVBHD+20OzBKuxD0IDMS
0uQrGvdZWB1VIlsTMorx63dMfse/MmNlNDA5gPUHsONKxdIcIlr35Dv2QCoW9G8bhzJDYbPWzeVM
juPApzYrnhbxd6XFSlOirGeMckjZABQZAx2bqLISB/r+5AcW4aCHdlvdd8T+91JoJQubzQLh8e80
adZUc7dNEY0l9O9lAtvJTkKftTIsZxMkfkmvvLQ2pIkRzfDXTnEbwKp1VSSxNDX9aD9Z9OdI50lQ
r+Kdiedgq5wAvNPrUYRKT20MCRJm+moW7mgX0/LJkf2AyEI/Klwddms5uHBxsfxgQIPaJmguR5A+
YiSNZo1tAM6aLCQ5U9o+iLjOHgAse3VDNB7HB3BCI129OiuZ6aQouJC8vSsfr364v3KKfowQq7u2
yteOLoSWNlEqQ04QCsHQYftLARe2NM+GB+68dtUnUHi7c2IBdQgVGuOWsVd+hRQX/qg67SvDUxOe
NczGPd3rTr+t+xLYjeLJbH+RSat0xPvF+7jwiW1NPOSEQduGeOMJObKTIJzH82OEPn6O7+6pExz9
gfgxxKwwn97j/vfagG41gbtsCEvk/EuEDIfkzHQ01xFvWTmPCwRKBTW+ktdFuykjINj/zDLPvNgu
TLn9nzuEEmqSxvr4tREVT4jcrFyxD1TdF0wkVTrm52HKivUJ3X8vR0aOSe5xl0pr7c+Pys/9NEED
jFhjB9E8PnTWQU4O3Moh2+KBdHg4eK8V6TtunNBabO+kvai+7Ph97PE6xwfVf/9mS6D2MNAtTQkD
ta1rA+bSuczr2DpIiRVKeH+jcI9F0Ud7tCnIUbvuwp34wYZMm1Q8dfLXqq/xnf4iUf6cnLROc5VP
G54HbHq8i5dLwf9/82LzZ1Be0EKjZ7v6+ijtyOzv2uD5NusDH4iVoCBwbsh/NT+EABen1YyrTsIr
CVlEhTJA7eCE6OwXPhjZ0iL6qU7DDTql9BTIKNmIU4h7pxCXUlIgsjb1bKsm6W0TpF49q4d1C1Q/
AyOmbQeAoIc0hCKTYr7V5VQvwZ2SCIzSQ+3O/6SpXM2OECW3RzofiYpAGrUFfePB5lxq4frjpwpu
4ZeUJGmv0pFTTJ60B5t6ZZXoVsbdgLvYvKg3GRxoDiAVIgbecYxjKGWrPUW0OBfkqn+dDih0I+B9
I6rCkRZRuc6yYrlRtdE7fKPHmGSMgBQU20Ld+klkd82/tWc0D3VXHJrGd6NsURusO4R43GhpYwo3
LdPRMBhDvO47bLEp9Cx4u9CxnZmnjsGBf4gdKtdrWPkzcAoJszTJnhTR4oHrB+xxLTBn4maYCGWW
FgjdADhjSmVUj/1xf0CcZQjiURLS45G7UdToIoGfaBkhfJO4uSGz2UZexyzAzKNdfee7xCN1FYJl
h2my105Clze1flu46iG9Dz58VdVVjrHUcqB48YhngCZuYkNzjxe/gdTPCFQwYLOUY+2Z2RPG+kEj
dHYeIlBcAhsfXQ3rILiXpDpgMVFybev5n0BFL8aI88NpMiMObAlnVf6sQcDK0uoEocrKaZ9zMQ9V
jnSU4OtWNpGjhWGgrkI4qXmx3ISb1+UK623WNR+9MJedvUACbO8MdbGjZ486im84ZyaTnvj7Vhsy
I8rwqI0s2dvSgxNlhsWrY0YLGaHLT9QeRSxmTT8G7ct7JrsJNLfsCC0MCwE325ZLsYk7VMD46Mre
2DPe8n/TB5JcVlVVmsK8o7h1jEv8jGvvWx8YNC1Djf6Oz2MUzDC9Pud4gwQ2DXrcZn5Nf1rNNPeV
7JDLbxgQ/s9hNVVJTZMAKKsuLKEWV1DYUUsZNbEd9r5fGZF8y45EbA0PqNU2bh5cEmUH/d0+UJLP
36et3gsUYsd+xtR9alkS3cPXjsBjDUBT3VOVp0a4YxoIM0CPIYBhJGxzvnvi2RSrxtNxtSFTnacI
sAbuhhoz7cxDEqfKLcBFyOVNkDzxw2bgh8l0EQh3xmBRLBQ6VSGZYq/p/hEEU6l7eJsT2NsNASd/
MzyZUldphn8XK0Kj9HsZD0gQCFc6znh9PiHp4amAxqknEabgwbupU78V7rzd0xTyCcjuFk7TUGxO
641HSYT4NVMyxxR7pS9yLnkKd0gn+Dn5w+9qdH6RqYeTvc3jO2Q+FsicZzAlb37c0EcrzTUoPJbv
6KbD65P55IZ03Kn7MZix8w72e7DilBBh1V1+IVBFfjTrdkUv3NiFTh7ZRI7ivrBmUIIsQtTVitzD
uReoqAt/dEez7s0AdXXXqqXuZcPJ1X4zYOZUwlgo8Y5oA1xA8/A24YYdX7LqOIBIBue8KI5AFOrW
DqOvux67zbCfmYrxPC/DK12QjqfXcmdqgXOKlYXSQ1HYRpGfFH0dzZXq1Yu2ETfpmzrCb9c/9ohB
yaBWdiQwnAcaJAM6iL8h5S5QaIPtGw3Fsf2Ba+kWkKOtiWOomg8KNlCmfI6UN84rCuK6qDT8MQiQ
XW6Lt2aTN9H5mOk6iP+Tq0ynKX1DPp7wvzQBm6g/o2LosPKx562thZDA+bJlsBWtOVl2B1LLgev2
aulOg86xzi1fLBBenvMhZcY6WocIzP3wjonRwGBPU53x7R+LxuTGVqEFexm3HkOdLt/V+jugqsS8
7vw4rKfXKDwemsRE6Nj+yDr6bNYT3ZTogPWTM7q31Lt4YA/DfFIoQurNmSoxuhLt5KxcUwPUD7AK
uaoFLJLDKBCrQDJa0rGgt3jq/3V+4sUXbj4fLpXU9+h4688IKwayqPSZSyxMmTDS+Vn/3fqq/jGc
1/NIjDQ9F6fsIYfeuJMPM98YY8MlpqZCwUHh2AZ7TYk1R8OVGelX6E8BkO8HDbdrnzT1ZMQBO2tZ
+G/86AS2bODdH62w4uPTCOgi3Hh75i6VWkOSER/ns0DXNyRNJbI8WaWuS8HNyd8yohgNfkDrZ2CW
S0CJRiImaOouYnaqX1Zw8T21L9Ewi744RByit6HDNzZIIPAyKizKgIaB7g3qqTFAeFntrmEXrchO
NvkKn/+w4k2A7e5zM0ogp4uKvko9HZ9U3kogxgMTN0gSh10fb4MKhkoPPtyhuFdCWU5za/upN6qq
eW3dlwOj3URtuK7hsMeiNWrLJ8TaFZLhy4wdPMKabc5iATuaGIqXhc1/0RVzQic/7HL90cDIU5c9
QqQORzcGm8MPXpx4mT06Qtz2O6g+8Rx7koPv5vmfBT8YO7ke+EVgo3Kn3Tk/veyQPp3PgLwRpe1/
W4r2WXrvi9R4e5dQ5PlYQ4VUm9dx+W7ezf36xmHsmur2zwFg9OX/cCde7tdrLFhRQSAqoA4JQun0
vwxJbNO6pi2DklKtCpzh79naXl7sdew7+lC0LEiqfcorUpRA7v5CEyk9nMc0rcB+TjvewPUqvx4f
F1p9jAMzi216Gh0NaamGxxDc04jo0dkyaYb4sKT3EdH0aXXfe9nEvxAWUKucnryoEc7exlrsU8Wm
CqoupkBR+k2gKtVhoAdPLZuJauKvrFjchI3FK9Qw5BccjDiJuXfSmCkvh6yV2ZA9LSP7SbCyUDTV
tYelHGIp7rq3qaIih+rw8osBuPhxmJ8LIjsmn46wvfaEkmDE+NbrqdTL2dzbf0WsYx1rXVyU5KkU
oak1KWu063ikfruD9Yz3Ew1X4L9UGMaVq7ovBS7vWsDK4aGdsiyeG60U8xwR8bkMGd8sR4bF5teU
1MDyf0TIJp+eU2+5t/01qUZANNZbrmNwnGxMPIRCAQqg7W/v7DAVAR2eL/reA+vt4ctuswxW0gEE
9MZ8PlgHXc18Axx4qbLzv9MbHKYsUeyOCo3ft98frQKvF84pHXRNfD12dBmMWvPDS9615rQPiVa5
U2F6j5/+UqgftwFZJkJxjni191HX58q0Q2+HlL8TxV+bPsB47KG3/VqYW1jkbtsGRfaOP9nILa/8
GB73WVzhIGtHuj0/qMfGZNHWyciArBF9i81++m3KqhI7fvIdw5JuHaP1ZEDbJmFi7ZNHbTnD7ODo
Y+Q8Ft7yk8R32iisT5AiDyh9+bh29T+MhQxLWrFJBWtzVHKVRsU6W8Ph0rZtEpsrpxC0LUupDO4h
Uh6ebK60rzBzq1jEVnUGwCt9Fu2bC3jGb0H9wo+pqs7rQ1KtT6eKk61yRIYqrmC1AcB5A4s4+/lr
tbSdbC9CfFImrnNDXQ1J10TUhRVq9RygHZeXPbZlFeBb+872z3y/AHKBmrg21Dz/sKXT6aKzVsTg
gE46Uswf5Ly83PkijFYl2wt/mBfCUkHDOShEhkfwj1BraPSuU4xt1WSULKn8Uj8eK6QrJWhTrES2
5URRrSNYwsKUIyq7iMjU+7pUdf+7Ypwq8iZdv2/ieQM8kt75trcJgGm5IOiCLY7zBlhYZK/6FsDZ
O6w78uFwqMDxnBbAiC+NMtGEVLqEUpDxwV+qU0XFAVLVR3WNV/Vs9dGoja/ZfJX0yIi84/Yx/6v7
q/Id7TMSR03iUdN1lApopF3/nBWbVRi8JmHjsGv61jtPgUunk4ybM3Xu3ecINPZp2tV9OvbQIm0u
vCnnI9XYIdJG2PND5c9ghXmPEFryXzt4ij+R1Sm+cvmavDM3H7+PegH5NATIckEzqjN1ni97w3Lh
G1HAhcMcuIOlSHXa5/s1tM+2MCYhPsl0EUTWVdnmdgXSw42PGC0+XmHN5Z9D0SinxMhCNLqrBq+s
64TMBq1reUTUQNoEX//ojyuDAT4l0EflA1RPnQqasjSEeM6OpsupzIIVTgtfpydiRZAR5R8sgjS1
YPz8+8+KdXDAe8qifB+K9hnbZ3zoluYH6uGuc6a4wux/bAp5aco6aYElFCNVhYLZWR6ewYarhvnt
qJZ/pO+fUu3Ui+4ndk530ysy7b4Y+4cbMP49B6yY091MjLap8CQeriXCoaTb16jkvckhZRFJCBk8
CDhuPXCLbpcT2sP3fKp917kKgCA4sH9jYYZZ3yuEgw/m6waRJWsyu+WKxe+45J0lH3Kds59GyMx7
KWy/ToFHSG+AmJOhjEzu6VeS961sWPVx6UeTKa8v8lHN5lSJamO9iwVer/iyIxzv7OcT5GLQNghr
zpVdqnJg1nSmndPFGvFVRpFxMr6P8ROe3tr/tmdojghbV8tdyiPW9EO5KDkXzWkKct1JBL0iHiqM
Ky2zQS4GeKCWmaFaX9XeF2qasOxUqDVmV2u2vUJu7esB7c68rrpMdAqv4qp+hCalvc0M5yPKkJ5I
jnu27KVVeKnsrTAeA3rO6wmcnQ7mwtAJGWHM3KhR2czmFwTz0ygiaAmTaBy60pMrobMR+aeFg+tN
Qszk3nD0k40V8NA3iuWF+iNtDgwFb6+Ic3nsIEtD8n2Y7Q4kL09znTWXL/qd+MRh3yCqy6cJgWA0
fHyrcUp35c0Gor5HlJf9woO7G8OAhP17MT3quiEP+C2ZEWB0jazA9as3TgiFfAX/LQbpiO0MHtEa
PaV0t69PUCQ6MDkSB2eg7YesEGidP8svt7Rw9nOsqoWG99BIe8m28aFkkgDdlQm/hL3GnIFjblvT
ga7O8yrIoXzEETxSVTysnoxadEUSG7BjwLSF8WV42s2k77XhN3EtJzqrHJ5xVA4UKAAk+fbYmwBV
Tz6TD1D9lHNqMjvKX7OU/bQiNT5+AN1oRSLr8VxxDBKg1bpx1f9ZR89BBEDOjLDY9OHcn+0jgDLb
hqicsMzRldw68gez1pRJja7Ewj1vHl1TzjwHWeH5Ufz5rwlufeFnR9eRPWwpqbAreAO6BVYy1fKI
QRsHHbxYGj7JDXDxz7ParaYxF+qb7Tf8fITdNEv0HmhW8e0guo8ZLopjZau819ePwkcatMVmtMMd
ZPGDOCFKKfaUXRFJ7cHUpsLIsbtJOH90LO9BVHLeHJQNCrm9DpQnUxQoJhtZgf5xM44caIzSXJqg
mwHwHLHj9+l6URtnA8AMwvYvAJ0OlfNK1w1BaSTcLwV82zIo74EhiUPdD1D7wg/m9e0KHDptv4KT
E1gOx2zkGa/9/0tQ+rWs/iCGp+oi5+i3EmdrolVdVMIZuMiwJDPToige5WZ7aLccVhNhZL1+b87x
rXJFVkZvjFZou8pTD/FMQeFpD6mc4KxwO/Y1w/2TrZkplDmoDsE3Bf2jegOhw0jq8LLY4aUidTDl
qwmBKv6BXtO8c8MWd08IkKCecAeajYPRKoe8jzm1dRR4Hi9vhiLLYgpdH/3sEsCUATdavuYIs+nK
aqjfSGmUZqGozj1h29UXGeF1dN2iBd+RID+yhC77rh8SYn8nK0yN0InFrHILlm4NDU96SHqmgRT7
0pd/HbWwRFdvgCiGtVZXJepBDx/NkaaeinlClRHo7IxKmsW1eS/5EmWBkhqJGrs3QUV1NzCfHxLB
n8IHV1abgTLScu7aojzx3ajG/2SAHep66ymJplxloRd6W9aBGGNuz8pQxWVUuGdKtEHxpogZmSgh
kUnXkYo3jGDtuJydAA21JZPmc9Hu+o329BfFXdc19fxNftO9l+HEDK9s85sJ5C7qneT3mCfjbJeO
xJDCR7tM4XXIfJOqOdBxI/LRTX3dnh8Dh5ZZasS6LRClV5KvEHIj/PHA1+AlCCfXyb7UU7dNrgIZ
24yob0d/63UXg5qDAa4SBL5YObCXniNuoWBU2fbZ2cmOkU/UQGDYkyJR/Iu9eSCR54Bx27668YuN
9Fx7Z2BHA8/St/gSOm2lRASqAfXn2MbgZW809nxpo/qnvBXH8P7MJTihyGhdOkb8dyCGvJzRvyTK
em9lOCtmQcWpXB5blwXF1fc+eO/YvoV8QaYnlINsNO9h4LkH8IlIyzbJGsleggGc3A3nQFZtoTIb
F28F+558ynrOivk53/pfh/Rpj/S0WxUuiktMMV7GA8sHt3oXeTk8oFBjlCVkSLL7NHFFsHL1Yx6w
TzhtOzU+eyMmm95RM2pyymQTpFLJ3Y+m2S/itlGo3t2PreAmXQVtXE84w7pFr5nWihzd47AtfT/9
9FonWdZIrXrsguV6cTgGiBuTUGzLudMRb2Mo34eXsbCf33EvL+iFeqTEwB/KWkEKgD89jSyyVP+a
qelykgPUj17MWy8WNeGMLTGcQQ01Ui0DUIJfhnx1X+6vKAeyBw5lpjai4J2cdqe/4jzOU3LKO0bN
YxwOF+Xza6f4DaujaXoqKF0jKZOPneUgPQ2YVOsU9q6z+YkEXLbQcv2mtJ1K+jwnVW8pvUSe0C1B
8h8UlT+Vb5I6b0CgfL8oeCK7hduXFN77NlGH7E2XiO4J7EeeL2YX0s0M2qoMN7I1dlLBBdXR2F9U
IbQ0yEOnwF3Xp/uTXYBI1uCeKjvqoY+O4PnUeaOiFQtopIw7Qso7gkaeJfd6OchpR82U0czCdCWe
bDJSI17l/WVCU9ttNcN5Qz1ZLhOD3hphEAm2EV/xYqAKeztKNAJTXSA/RqiiV6L2HKuNLdPHZhZo
UVKqJsijfL/j1QEopXW2iIsI3E3LTzAE8mO8fAsJrFnS3qtvxfvwWf91G9Jx0SKDFIiSftm4PAgR
ER6AeHWiHyWjZnRf/kjCqL+ryBKN0foxLMpC61gxNRMzpoJiraGNlr7K1VigJV3jMaogyyCI29Bj
nfyf7b+4bc7Ctmudy8jTY1SYcN3jRgpoBd9/j8Ta+JdCGJrt6jbpZCEXSjFe9o5/8iin0+Hc3D+v
o2/+VajvKzd4SuvBSshWIm8bFulGZwQyLRvNNXlXTDRiHZ5loqiPJeiRekfe4VQQQ+L+ngoCdg4d
bLpA5GgCDx1Gld5KNKpGhN8jDA/OKPVbjnT6ImHMpI1841HgYRm9jg32sihurWRdKC+nmELceAZU
xRVbq4WXVZeMj5PHlp+lyjIsu2GSlScRBcXNYNXfnHOO36wROt0m7hSQRHG6FPERWtsVVaFK7n5Q
MCai9nko92vgV5k+A3R0mo/jueQ8cDGGcO3rYsP11nGzSAP/aUckLf9FGbIldjwvAjU42IadoMAO
4Ehmi21B+Oiqg96TQtmALnNi3tua9OVTw+UxVca3Ym51EONBCD+EpicaxLGwlFzraVxLoJmSOCJJ
B8OUUB5aF+qdMLSoxaSVEVNgmZ3q9MLiPkvVZhSCPtMBcQJjKzDohUSiLhwFGDgj7DUWMahZ59yS
iS05bLClQx1UAdz8bmgK0bvpdGxyog5IAYpE+Mqx+4nC1egRRt4qV8doMjHktB0v7ojSU14N7j09
jYLLWfTg/mCR2hiSGfttJ6aKnFmyTx/SuHcge9kwzEp3ohlvyIzcr/jL6l5e8kgSfWktQvRpZADO
O9Ky1Ms+ovtYToCrL6fB/JkOEKG6pi/JB+DQrC5BQ7mXBrmm7coHmyh7TCCmpaJQEZBjjiSV7/p1
o69wzMCS+uTbnXwVWb5vz115udAXlfRLFA/krwnLDPNThwMEOPkPc7vcDc2CJyreuSFqnnXczQST
dNUVQ5ZlKECT4Ch2xoHpzfYAxM5bWR40+Dorr1Ei47emr7fZ7SEAXJOhVuRvZUiCagkPj3OHXj1X
4vNUV+ANVX5LVk4IZ3WKh39IHmyVuxGfwvASQxkxrgCPj3KmbrrU6KchgasuOKW+Mjgxh05HCaPa
QbEfbIjflMOCEoMImzPnJbu/5RNlPiaEd5SALDu3a4fkoGd7CvvcKM4MtgGk50mDxOetHkYqcntt
vGYXmrIoYCnC0TOeV+G2YU2gC2EicyQ9fPF9rJ4qlSle/eN1XfK4jLvvzgz+fCNXxqqodln2ahDW
DY3FDLAhg2qZjqA8zYr3UqLtO+kEEM2U1zY3s3d84BnTqrjMXoT9SV9iAY4BkE78lYNI1K937Cg3
YtzpBW38OqZIDU35pVz7fgBQFsuAxHe2Rolu6u720G7lTid+2r5XqDughIb8E3ZyetDD93RR27KY
/QhTyIXphliCJLvwpTo4Kasgq/jcCizuyQZjPcJFJY/r/w2zq1pwI/OlzVRetAYIlomXXAXnBigt
pbqcq0LCICbgFPhhndn85glPip4MWdBtOnccDhqn6bIn3X/EDfwMi9qkfXXnF8AgjZuGls6LHp0q
+cxXSFx2USDkyd9VWLN1jhTxHsIczPBrFhFXmH0jzRptOb/jmew7MEMqBJxXhbHFl0DcubUPjQEC
XGGeGkCIzPAzcX/O48FJUdONWWoV8jy0ghvz+vi9e1hgz50NUaI8K9Ao1yANIj7LTJjSpDiD+lJC
X900qAh0K0IPK7aJu6wtBG8JFe3KoKtt9gz4owyLOMedZijW63u6kNYX/lmm6IpMXkT/8oJER0Ew
yxaYqGa7BemMbZDGx71RGnL6DbWalOxPBGMvgQwt8jRoqmq+hNPSFQV3BT+U0K8N99ItxZw9xlZG
zUrwXjWFXLExWY2/jjM0w13RAtx5PTXSY6cwg8VgqslDfR4MZtVJe2bN9HDtxMCwVWQfW4DaR0X2
z6ls3OM0PmPOO45gOCca5kOLQXaNSj9RjZbaAP35lIZR/8kl9a1i6h8g21BtXCGDQNkmcI7RXMk+
W77eIm6RohfNyLrzKJHiot38/kWHQiF0sGnSowkrXvzEG+ZoAqpUesjyhwXFjrOaFZlEW4Xh7HWL
JqfRD00bsnNQFHv5oT1861vfu7LoAcDpHc0dAxHgep5+q5G8DHdaZ1NeTguoeTf1kwn+RxkJUaQZ
9n5gFt/RE+wq8OI/N7wRw5JdEO2trUZPQD6oZmELLeLjv29wQ7j4IwEL1KwkrBqV+VFbV61y2FlS
uenoq79Z+KBUXS7SUicdmQmJ+HwS12yXtY+nl3g3XgmnKj3YqbE/I3ZC5Pd2BWg5P1bJY2gP92nj
sOLDi/BT6CJE9r94DqsK8vajEDjju+PXIGs8UyKIBnDG5q2zwusfRFhofdzd2T24gQOVtxGR6ZoD
b/N7MjKN7+NR77U2g40xZMqbRAMNyVIwFyBVMxTLXq7x/dw4BR3GHcwEegoF0gUfeMOzMcSmywDM
njYipPYpy2voVl7eG4w0VIunvpegcAMW7uPszWg2JnshQOfJtot1CNZ77Nv3R3A2EL6AHnygcAJZ
C49oQEOseoMEE4rYatrGJKPFtzcNPG9+aWz+gwqWwylMOpJhYh4F2eCSf7+ENj/MTy/D7az7Z8Kw
V6qdLW05YpqJkAfOiBg4oOvchOX8sLGXRpmLCoCEp/khK+Pa4afu+TP3Pw8ZNd4U+JhZVAktW8W+
FU9KxF3OHkDz1Gf8mhdzMclnL3kj5PMapVPS71c9cV42sMV3qwHOOdGI0F/jxkZBA5kbCEyV0xVu
Mv9QQPeiOgEsD2cYRrvbtHmbxLfKrLw/5jmp6J1ThvcRDu9uYQ6IyZwucLidxkG8W0vK6gSmY30m
Mz+ZZod/lbdH99JeV/IrDQurC9jcojlCfUHW8N5EsTkUBA8bpE145CaK5SwKkp3wKj9mo/oKB4sr
Sl288g3F9lXdLOvr4PmqTAbtc+sqf4eQBUgSfv2mh+K7S2FS2GEeHgDiiC/18jmfxE9orecq6ae6
c2v+k+8mI3wxx18uLv6RBTS5JcqOO7TsYklbtbteudn6PYMJZNgx32nK6WdcVdi9KStswo2VquBj
mVxXD144aikGTHg630NfZuPRJKDS9N/moCOxGlD0zcmOFfexzhmmSrFXVlSMNJvqyK9rQzTrrct3
YFTVEbK8T1MJmMjf76cQv9QtJUcvfs+Tt4QzDnjO14RzbGE4mkqZmBCKwjEpJU/dDfkc5wakJF7c
2+RzPdLaPm6kUEk2zaVvxsE8+B7BJ17UeZmSEWkK52l/kYfj6EWOD3v8XDX33EWTKt50/uR9jzJP
QzGgq9bgWPzXm62KRzZOSUvjdyDWgQjjdayu7qmtskeYs+80pXHm4D8wBh0rTwkv16+xhzcPOTLa
/5g9j0SppK6BPTzFmWaXClNCyzGk+lVN47NDk4jdnD9LA+cdVCwb2pp9x37q1qzfIpFGS6qrFakU
uY9UAaycBqbbE+mSHtkHgeeGQroWvzP5iWSuvRUfvy05A9GNymbJp+MJ/k5Les4acUPtLmwsGI7z
GohYREpj94zMwFV75n/Cfs3DIO/XgDmet+1+34Lpe03gg7So1QlsFqZyZFzZY78cggXL38H/LtQu
nmwWj8OeZEsB0m0FGg9XOnIra/bwZmD/zZYp7glo70RsAYItVpgZiAdCToBWKxL9H9fbN3tmD6Aq
Om62yuKEYoN8Q+vI4tb9B42aHMvag+Ar2dkiwB+bPGZjhRGDIc+7pntCCHAIhjx1eIYdM4N7ryGa
47lniCmKOx7CKqIcwxiX0Oj+GkdCJe+m9+/DOA6GhfSdB+AUv/ABwtSzj/vFFW7PLLCzJWQSwVmU
ucbmwNJ4APE6sauYP/mtOAjBskrr0CvytgGsO2P3WRNV/1bWNkr9tFnDbnsdj2RlRWLg1WXNBS25
e2uFa25hnBoJQHEgk0PskyWe/cJxoQh9X3e9+zkAVC1jaOojRpJcPn7Rmp5jGehPDvLygL6bMzkZ
beJgPe525pGz6o98+OOHZVJaUwhQG7AZXI2XnLg9ujPw/2EBsbpO2CeHVwOyZVxR1ViwYjeS57ir
LT8Tfoo8/SvkcfXgtGTOCmbc3lC0/jxrEFZ/WgdsDbIYtW4LKdwlbDz4mvRbY2j1a82M+nT/QhU7
bJOVdpmmdX3L2p1Xn+OdhImvSXFbe5OY+Detx0otll4MtJKkK++JGALKWBboX/yQ/npTkSn2BD70
nSSvAk4tXN6rUuWWzndhQ68gHjOvaeJGooZUFOM4uvBv7dKojkJjQJ0rZoAXeIchq+qUJrT1JTDx
D3peX2Dgt/lnY51v4kug+9TZfax7Zwt1ihsZl3A4v5k4ngMJhyJGA7xmSrzbahrj/afst5xtymf3
q+2xtNmaNZPXD5G1y9agKzFGegFMw9JcMwuYWoObuNJkfzWJI+P+8wW2TQNMp0Ce0Xm68Pwj+hug
E30dGNGF4evQ1X+lR3ZSacDlyPTXtuqY0iApsvYJNTXdHVDuhGQkYcZuZyNhDzSVM9NZ/TgGj0No
2mLFVr+zlTbBjnvsMyzjoOgnxIDeicows5BuUF3X91eiM5kOhVa72YaaT8iVFIi71yQdeQ93UYyn
O4y1w7S2BZG6LfbtP2e8QODW3JuRi90MbSoOiqczWnlXSUfa9m2SC5+3IQM/8n80hLGbAZcE7i+k
1/KIJn4g0NKUMsPZziKfFT6KsYuX6qzcY3MXMTBYGyo6zgvR46dSnq1u+u7dBQmVpKlkUo2qxtD2
Bcc14/8l1QNNScZZqG1Q5yamfjUuecEtq7OZzYdUReZkGrdgovwzMi5bPu9HfsmibzlTNsbmV9Lw
rDysIPS3WRh5/Hi2wloKuAa4z7iYv+4M8hpVKuyxJp1SEjIc3HRW1Z52tpql9g7nPneVr3avn7HD
zZMfMs4Xv5+WqkGEjSDkwDW647kppHQmcxxIw4RxeKv1y7Vip6354rdRW/t4Jru68fAk35F3TNMO
vG/njUF58eIVl6ZBcUWg9Cslw9DmL8PCmk79we6HA9zarMeguI73iESUkS1Y1Xl4/LAUUJNbu5TQ
HL8Gh6mX87tv6l5NJQOVr2qU6mWovb6bwiEwOchI2N9gYJjDL7582QDEG8Ff+Eu7vAl0BRJ3vlgY
Y9OzMD3iGs7AGxn4ydFiSAZnlcXIbyoChDnjJHRMdHGh7Jrp+EO6fvqiValH1vSSD/xbbQ+ixrzC
IVxRrZkb5XSH8cF7Ym+bDebhPwL76LfDa0JNzJkv9lZ3NxVnEkHPDT9OuFVSwninZADSINOsMRHu
C5lvboaxiqCI5wbIWaZTDPN1hKyEO0DTynb50KLFOJSP7h23gTNbu/Z0QpU6cWtBNTjVUgjee7Za
1wjf6usYJinGVuvbgTXWmcx9Y6/MmR6CCUqEjHNrC00nN0uANKY8FVPnSmh4K6HaVIdy0IhRN9wu
LM3x3Ksdo35UVH/nO+b8Uf1OYGrDkp7d2hm3gGxUYT7uKLOdqfJGePSosahvuxaAW5jKzsdnqtcj
Y7vdPDPkCXTVnriZYKxkAAtiJBtgMZx3sl1JksCtkiB4QkZlhF+0F0oWyNfFL34I+/Fpfjo6HlhV
Vt6mxP96gbNYAxXuVefqcYnpnaZJ4z6mttR64pMgkaRnexMGYxDX9C0lcOhNRPTjA2Ju/6vOCpMD
1yiM3ZsxHU90sX4dfroKXdH0uItfotvPeXxeecxgpUQfZbYNq7rHTu+I7SAkUAAphs7DUSCdE6R9
R8C9F6+BUbLZ+I6w5GJkKFczxNBTkfcgo6FU8q1CaLR3cwoCRFaYIl1z2AG4m4qdr+HT9LxKjty4
BWbRfiPpoylUoPUIeaBMiUSSUJLL/waUXUm0p4DrTV0i43Vcb8/+crpKfYMt39p2OMaXNmIhNm52
i/c4VfVKmXLo06rwfX9oy49v6c0yQetPWlhstUh1qg3vyjEeUR4bSQawOIUgZhzO21qxuYk5Fw9k
cQ09Ki3SX/a4ROWNMCyFONl3A84ACgyoSFlwPejgg1Ygj1/bS1F52y5thmWMrEapN3ZDOWy4Y9R6
FvKuVLw38M/2+vsi3F8gdzzOCXxCLqmZRAfIpdRV2j9FwWu8AUb57hQAj0yxFld5dN+4W1NL7/oz
Cr/UiujQBHPnLmpZoSMvrPeUSUsHc2fv8pVe47m3Pt7Z+GC5wOTFdrKTpEwreEBi2vZVxqA8vvrb
VIklCeVURAmis/Ogy2dS8t4rq6LCEAxA2n+NpfMTWJPKQriUqdGAjtAuTYysEhwrCSw1pZ8Qx6Z9
+4cTCUN+pFRWy4Qu1UoXN/h8Fazn2bo6ognw9AT9n4vE+8nKLekaRg2yhOo95UWKT5VvwMw9Oif+
Y1oIC8StQFrTlhuQI2tsefQtB8RMcjCXGFpTyiIRwoZ0J1P3ywX1u/09W1xZN9O2soWd+BWuSzW0
652hpfs22smhLJ5ZZpO0s10yo04fTNEkhgZg3SgKVSesrhcN+RJsuwoExA19JhaWA6lyVw97RoBt
/yO0pHejZA5vAjnZFgmy2Oihw5CxwGr3xP+z5v8YLJ1E0Op/6roxNcokISBN4kxBTdjibjjEagMB
pqiN4Xfnl9ckQO0JM/PdankaXiTnoeIvlhB2spjro72zNvK/VbvFekncDgBLihFP9ZGAALZDqf7G
W7uAV0Xr4ltA/27Jni5Ev1VOSb2ZW3hdNGlUAul57sVDCAOFACgvxslE3PBBC9E5r6G3bxt4G87h
r+Pr0BBrl3yYmXiWJtOd9+EESakWEe3QXTmV5Y3UOdmOpZxYV7eQiycmOIIs3j3BXDGA2K/M3A9P
hU7MEqr+g1W/6VWMxPJcOKp0b2E2Ji9xOlKGP1JGmcTtnp6CSCHy2puNFPhBMi783aGO1oOBGp8g
zX8OKJuJ44HT9COl875SZSLlwP0v2PAP99Gjv8DwOJoN4M2Pl+Eu7JKJzCSSgxbwYsIWqeuSEbZk
E0XsqG5ck0k+McOOl0ah5KN5jyz20TTRKKLeWB3ynjJG2MpRLpDtF3H8aKLnHPZybGkAJxshGL0w
w+K35UiVZfHtfldO9l5pKyIzBpYnKZLIm3+WHhn5i8zeJTiFcNp0T3vl68i21n1aRina2gNyevcn
P0B31Ba29wKmOLF9qeotkaj0/fRvq0POJFl34AqA9seLBBi+yKAjt/V8VAjPLyR6nlk+XbFcVkKK
j0A2rnpps4x5SLkrgGyyQ3hp08AyZZSX7NCHnaauRAo5FPA3jFYL/ynYgQwKR78t1XRTqiw47zAC
nHDCaIhEIs9W5BFkMITCdfZDAHkmR41AlD3eOeeJ53mdWHlxCVitIPfaWPqwXarhg2ivmPiicZAG
BjPbjD0j5OArGmTVCCdMmnAd0YNAViH8XzcrfDytvN9XTEq93T0L/AWTI1zXKmweqxmPLMxEbPea
ShJANdKXwLgReNvIToBTNWWckdJ52dn0RkDZnlQTnrusmfS+hJEgNWhzMnEtw2pa8mQbB89bEcDX
AmI9OBiF7gUZCAKN91gnbMvaY3TqXewTaMT/YFeApMeru6xqPWjNbJbdSntLgXqWpGJ22jLQ8RAf
tjVlkR3i6uCVMhauSViqOV5A5IgnhMmtoJw6jM7fLb2lQG8y+8I5S8/dBacb6XfXVIrjaTWdDyv/
L12n1Xci2HqNEEuliXxg/Pi14LJgvwrpS2HudgLQ7xddJPuxU7Vta/CWi1RBDDLVS7fhWL2/maO9
/86oggD35AXI1D1Uru+wCQyBCojqBqYrAA64oPYAbtSLHK4b1gXiNCuC1Qk5MwNbcg8CIxGOUxgn
gktbvT9x8jfH82VMShDvGXyJ1sSTALWzLz9ukuSVR6c9PHV7GlQm2Uiqyn3Z/tLA5yrXIvhRMqyd
bty9AnDusz3/EM4kFJyeEuStY59D+Wg7zXut0vUZrt7N1wt2+DYYEDdJEDOyIToFlcPTyv0F5u3g
ZNRzfjBpeWr1SdxsHuwOjbHiwEK6cUmCHZwD7GfYiOnLDaIK9OcJt+X2XHU9JPTFuF9dcL4RTZTt
CgyzATV9ldPRiiJN/1OB+nlPXiyKfRFumg9o8teVVKs3vPYnWnlNhgi5LmBF5n4v1TPtzlMdNzwE
4nJb+xLz/kGUU8JcJoY4HY4VXmYfoo6YAMsW2l7Imo8ELCdA6HVRsxLNJfzZT+Az2tb/acX727uD
MKjdzFWAfwS1GsOVAAd27UwVnX+CJ0BQ2eS9wY+yoiXlgGqpYGYJpxe0jTpJrByrFFIdJh7lzsFj
CF2YbnqvOgTbwNVTrsuT317QaF6fXHE9fpgNfKajzWkn38EIdkglR3tXsLCD/9SWga47oiTrV2cm
aEld1NTIJWuCeIYwLVJgOvDVomYda4+CndJvZmKJtuCbOyFF1U3NloviEhZHkc9kpcjYWyku/BJF
lq9t18V7mXBuQLHZKEKr5Yknul4A1bpJNHhf1RtY/p5jNhQFj0aiOeDFaULCZo9ngcav1R4oUdIH
8Y535FgIbcKUPZrZVvvAfdOfi3XWj6grvPzwT/ssp2QteI1l900195mdaXYOWMk3ZlyEx7pkVzg/
0fbkyZdF6EKcqvCzVs4qF30C5RlGRYhnPezRIReJni7VWlDeqO+7otjF6EZW+lcvp2VDjmxuBnpc
2QufmH7HMC5+77ssnwJx/h2G2oKUZxRE3anC4nGlV8r0K7mNWvAOFZDsFWBAPXtobYLGZc+ZJNF0
2tfr5ccA5mjlIQcdu3tqmxsC/8FnHfY/k3dVVJ2jhiKAfiAfMexnrHAsaltcow/yXErkWD+pC0uW
k0aDnzMqkn2lTtENXINy639d7QCYOz5YqqmGwDkE2xYtDaLthgpouRCvH98zEy53EHav4TI9xY2d
HzrkKalDHnRCQaLjjofxTc6Wi7I3WlCuxGyOu7Ri5YlHAzG9SGP9L7hVcqOEkPGK2dzL/GBIrA1B
IwUcmYWVscrxMegl/vOXY/558743AE8Y+vXFo6al7Tsfh9QpzoucJUvdm2iapETzcwzrY39pfm3b
n9p5CYa/VUySTwf8BNq7ohkwRBnRapvbTpdzkiLhFMfYzYzZMZHpeRWSzF9BDUVL44ZXwnjOWY4f
hTaZnbqGfi8zPpMixWPTDHq3H5bNoO3E8f40U1EJ3U08IScuVBPNQWQ9QYvpYyTki/zkLz5BZNYt
4Fl62oQ4PFz3L5tZ2gpCSdxAViH3ct2FJ4QJJ4RGYOLhDjibrHnK8cOft6jKMHVpCtdTAa+4hdER
QNdt8XYvsfbLFrbFDkanQv8rq9GxULO9G6dCdmxTYr1TNCr1/LHOMyRhNLlhiTUfPWsw9obr/frQ
SYMC3eR046HZmkphObhJ3RmzOlkqGObF3oTF/890wcboJ81Zmfv+f2JRhch1Ig3euPRP2yqpw/La
k673BzMptAB84Jj/uJv0W0/1VGtwXPb/aCk7qBRgRGKpGx3yatybcCIoUcmLw16j0Th35zNCQmD6
V2rZiAbx/1/9YIWEgwbWwJQbgKZeqvv8UXwgbJSGzGJXeJYDA5bkwC8kUfRKQFKc3Q4D8KaAcovm
IECWDsIRNnUA0sgdJpJPY/QMZCi+MBfK+Z+yxQVH96oVNak0JrlZNznpgGJdRbkjRFaHY6GisOew
ZhXPtd+A3iP0rM/uSQb7SS+tVKzmMqVgP24FJkQ7sardc459pPCgRzoC5OEqfmIwd5Ez5qsFsdy6
hqZKh7WM1l29lnn+QC9pqeAPWhyMT3NcHgNtl0DSYaEn8LsXwUCrPbXZnS14C6buGYMquf7OnExW
oetjtTkraMyHD9dngOnhOIIOzUqkDN2UoqcCqUuQaqVfSayuCvxPwgzQqxUVYbZpncsmzeY9bRfI
Ti1h+g98HUkCgRcRtgXsnU0XRRRzFxx0NVsETQK1Pji4PXs1Il2Wb9W11P4d5j5UlVlyzP0dSrNe
GCkBb/YLVze7xzr9Zn1vhM39nqqRus2mt0T/Yj63DF16oyPc+cwVwYdAmt0EBIVVAWXNLPKSaLcK
GRnb/kBPA9gKoCj0/PucICfWDGan6A4JUCU+SP21atK/YbwDX6Ya4oQN8NEOI+MjktFIs51FUZ2/
IBdqQPBjv+Wt1xPCmiHrf+JgIH2xNA4mkr+g6nrwfm3odvHmWOT4XHuVTUr/47jfba1C1DIsJGPU
BhzDslOt6IzRFeu5HfBpADStUyFC+y8QrThG/GRJ+AHxR0mD14ubkhqXGTpdw1LlMJPNRV626qx/
LM/PUj5uImv60tj1vB8RfJD1w/8vGD5J2/IdFySY/WyERH9env5sIYl1d9q83St7ReJ6JeLWODCI
DCKCZoQHcmrBuXDIlY637oyExGHDyoEye5zuhLSp0Kj8lEKbLw2eEJPTLb42CL+SBmeCnaHCd5wK
wI4AqVuuyO0z4l1+nUmLVEigeHvLXS5jdDzqoIzal1fSRtA2lZxrmo4joW3KZdSFS+wQwjpztMKB
vUc6/xZ442izlW14HzYRjoSXgaKOttMqnFrPDDCO2GmQX5NZAylfAM+ApUXocncy7Dr2Ps/UvR+Z
06QVfqis3amWN4qL3TB/CRWUhwxWYbThsDEzEZDJlmDGtANNYNzQHyfqa4sRz7ifCUorno5GfFOZ
7HBMrfOPPWAIFIhZuWb1Bz+p6b0xohFZnH8P5mzp7PpjdXKDweXHG1taGrdirkb8pwD0tSlzPbS2
dzHyCpJmZhsXba6r1l+0chOdc+N9iyeVLo4QI0/lkSEg+a8D3zXWvDYIaJaPpv/LzxMBPlq1vd7i
WHLhF8qlEPjKnrCz6Y888fV/wsifqw0bke9IoRqV7zOwYZYLEWNQh4CwS3gLUmMvu6RAoh2JB9yM
7Y9d/koPN/TRiuZgboOCXS61gGgvvRye7sR/fitVhCS+FhORBU0PcDYA+bsPlnARjpDTaJKkjgb4
mrwtc4dLqxRTQdchOxdd9Pzs9N7ZUFoYbPS8VjN8GXPzpW8UYRE3Mw4ZZ+YPiEpxW65LMHARH8ci
V131spdhvxE+oxMvVazf8/flzknZhY7kt7LXGCHhX5+j4karSCXbc1RR23Xl9l8DBvPYMuEpOfWY
TGgib7Cf2OSVczgrG1Aioq9uZg5joFigDhQEKSQ2onEPGhDTyJvjrg51HmPiPGLg1RMn5n5RBW2t
lM8a3naJUZ18Ua+KtVUEjB2NAbZ/iihMEE/jlEr4j3nlNsVgpCtFxrDESxYm+kp6NyVj5g18LQJ3
KAN8aFgaFj1SuqWibTx9xEwxRMv5QIkbCCbLFArg9BnmwEDqnb6nYmmtPGQ75jSxho3nofbaqX0f
IkKmDj+aa70wngYjvIFjDppNiJYNysKpvRY097a+G02A1EaypElBiqHA8hV1nnlEAmJVCuPfii1r
H1DQbCE6j0AxakaWc3+2106qTpyk0XuSUvfcae8eOzPhfLsunyGkDBMI2spVn/jtOKpevnseEF+J
QwLluZkdLak2Lg4hpCLDQtjHzIeg9jPe+mxsebFNyInoBxtW4CErxK/Oe+QoKxOijVT6dg3m2XE/
Cd2KVUjwJ8IEDdeuvQE9BUSn9QPML6BMXUiuRhfkz4GylQJ29pboOobODbnUyHXZGLagjDT6Qbm5
2g/w/c/O9Oo1VNHxSr5mcrlL/PXtipdlvPsxaZx6CXTNTuxOa469lcLi7pqfD88j5xGVqh5F+tRM
dni5FPB+rqNCO8xmrf57uNorGDohBE9AgTvKIfnHGGOAdZIfbcIoFpu0jloPXQWE8dJojkRNjhWR
pRtKO27WXT9cUkZj1NnaHP3UifHDkz0bGAYKcTOhUOW+1/oX8AY+9fq+onX97fWgOgIrlEDsATCP
GMoK5zNNpEfV1ObS7FUAIh/PDPv9H0KCv6ChwUA8m3AfaOy5p2g+kOkDG6SxUUrebNxcWa4560s7
Z5mYjnRySbJuF5+exX9n+H71On94L03BV/JpzqDv2B2vSjVeyfB4dXiR8ETPO3B7/zNktgVBVgA0
gIBUsso186NRXAHnmlid2GleAHZhF/tRYm/SRkGNWjX++AsyB8/T2r+mTjLclAmuJeaCXKCpdwuP
lieOM+GndVQxPS/dNd1LZS0IMMBsz63oULbRtdJLAEAA1Q90nF+canSbXlQzPcCFar4JS0z9xTdf
hmO4WgbH1UdH6maZx/rjActFvSgf/wh44dl2R/FClElCf9m9PcywWVkgTCYgoBjKwI1E7iV3TCFY
fQS/5KhTwgRAdyuI+pWDRQhD0ciol5W+6xYz8c45kFZkSBIIIL8uIQs4Z5vW+TjVO2s6RQqoI8vk
t9irPgXDFLOlmOmZ3w9xxUTr1oBttg4hd182hkVb4IE0IKumaDuFyDiAC8eWqA12wYm1HfdXfNVO
jxjeiKoga+2vmzFtu2DPKvmoy+FMJChiBvuHNeFniKEBgae1fSZe0WRox3ebppSLYJKqbsSTd9QC
PsScJLvtT7STKELpHs0nnf+e/R0OtT3W8Kc31kpT1VazXya10DyKFCyt41DCLB+WWWAlbjkQcicq
SJdqRscIkfrUCKD0C7MwTK/JZPGovTArGV5ZcfxaRklpd5nSLXKLYIOPkoiDM8GtJJbX3IJEY5QQ
V9EdyTrbIqGsPrETVUzC/zt08JoFmkkUl8VrSBjYH1GM6eo+uW5XYWCTIAqyMsiNE3/w5lAxQGGY
QODnuBCb4aStp9W+HMopsuQhx0RzJuNWvrIZcptevHuoy53LbkNr+DrChbnQSubc7RLn4NUgbqe9
6Pm6pCSfFBl1jCkAmHzCBjkXvWBxYTLcuu9ehsDo401mA2eGn2aaKxjsFAUU6P32ejB3PYJcUvjJ
8jPK73VS4zBT707y88RIjZQYotzOJNLXTc6UXt/y/FzQ0kFOArpSAgoFjsxDenuS0zEtkQbclowG
/Px2tWWucGuyyPUyB+/RthvTfNlius6nZ40YCrSeNOJWcFA7FySH32jLJTZ05i9rEa3Np0R5op9E
snOL+bLZIqwONKfXBK+0AXThOfwpYNof0lty44rntPFLQ8LwlCSFdugnf7L+bSBWT0yjnrOowxao
c1loB8aHAdyQciTF2MuXRCjpD0tcw7aV7x3TrEUxKYgf/UPHcq/R0mvf1XV0ujvSyb9b5Ncqo3Ei
33qyn8sOuwi7r5/R3cFQoBHJFOOkh68cLvyXHjNyy3paKvEky5z6K9Nib6UEHWrWzaBdmGLaPC/b
wNyqVXYPm/1Zj7XefMz81gkxBbuHMpZXZ8Dnt1YrxWmPVhgitqwr5tNL6oQn8T+wylEncEufWNkn
EFFc/OH0as7YXOzhB4jHQsgvC+xIxXLVtj3wg39XII0h5SjdsqYHLDEW3gx0xVoD5yWLrEbG7szK
AvYRKuonVxgKfivF6aPrq9m3QdPxXO78KbyQixVgeUt6M1fWAPNouYT1sCURHQSGeYm/RXpPfNso
m6PXG1B8JWrI27Pi6pkMAQK+Nq97FpNJqcjyzbRsGmg6pz8WPkZJh4966prZ4E9tCQQwfjNz/pb1
HIa58wikD8qUILuCqeVP9wBNaNo7d6v1NK7LQqWkfGW7zzInm8riwEG2Ln7eZkEfB3Za+jMXYsMg
+aKYIPynbsRtvUMvdaQPB15K8BaQK9WIv0lmd8EZLzW6zoAjkzzOUVGu5GQGLGx9f12F6xAi7yom
WWtKMfpoL9bOOSw/3NQNXrMfxrSyb0cKP/YwUVIw+AKIUnHpgUvHQ9WJIJMAatQwC0AIbJt0YIXc
2xzabGRer/IBzitP+oA42+imthw91+/5fLa5rPoYArCc9f9E9Um0TEAg6WmWzaZMlzTBhjRrikRD
9lFqWVAIBkFf3VnI7e5LoFsDqkwLnjUFDtvL4rCkOBNbAmay++IjbY0m7ScqTqnrcPQa6Gsa89ZB
ccFpXTCd1QqPNXjy7tqOmstMavhqetoIAWE2PcjgzEk8uesPZioUCxi953s4Rf4520YbVsR6KW5J
E9UFbkgctgoZ0nQUYapGUEYFhYtgXvBUnUwvjbdVrHv3PSjD3zUBfNavh267K4yg60N+hS97L4nU
tC5QbYA7qdeondha7xRdc9SwgA/83Y+p8OQTd2Wi4j7AZWFX4jsnVRgIZVIFudZdUChkm3m0020J
n0JBUJ1Y8rslMdg9V//IZPKPnBl0eq7X3Uo+sUpzjhokN91aZ8HwUX3C7c/RQEWK5hGiViYzjUdU
w5CJ3S8uQEnlObe4pFZTqrjv1C1HB5HBAgCSKVBiiDvKuCRPE1Xt0tXO1qbvIrBDtpqZgBIGCB2U
Yg9Je182mUt+ISGsh+4JL6T/pe4q/qXmc2F++Bn7adJLH187DiXrQYj3b2z9E9+sMb5teZ9flHS3
8fptOVnTXxMYz0m3joCUcgd1dq7rcV+/xc3TgrSB/AzWDv0OQ+zA/oOQ1dYtU02Iw8Mj+k6Vgfi2
GuPf0unk5itccNKSRiUl6j2lG4CfosYJI9oyvb8DAQwisqChGT4I0VoofB8A1Q0T9+msJR+JDXoQ
t5d3bmqIUBahObUe7HwXr1pya1PdgZNxbsmHG4pQayhHsDyG+kNJQc9BwzWY6VylXCtzT0evlS7L
llxi23GozHGipAO34gdsyUrz6hObRilrdwFBF1slTscsE6tXSX/9+oPKa8waqrcVVEEdATFojtHC
S426hYbjJRHHg/DsGTI2bmEDeFUHVTrrss7mJfOfODgFfZSu7BWViMfc33JvyvvgbC+LX02MCdLp
Qp0VSSFhnWPFmbOyewE+Mx4tDgON6+CIDz1jNhCkW8ItGt1Jk/PdAXnfsgRNkvieRjACvM6ChSjP
O3FlIjdNnnK2AqBnGyMI+e6lJq3Gy0kovitK3PkUHfrDA1hKfvNktRRdZmRbpGTjNnCbC+6DAmAL
OZ+THNWYzlKm1KAfc7n+xduvO9UukgukEP8Ygcn7fJa4OCc0nnoLVDKv8Rfwkhv3I5zBT8CJ83rC
Jvr0yFx9F6ZnPwe6Ns/rx26rKjEP/plZE5XcwNIXCbJvp/VLoqRZaprB+vTPMYN+0rsLXqVykrhc
iQXLIaitado+KqLdoKJw6do+kOEzXzsiAjhtQeEkDmzjoaMSBU9YmeVWm9jEih2IhALN8IZqMcA6
1uQxFQhImLArU+x1j7xpVbJ4gMMNTmVj+kAxTlKOWQiXEkxlV6857C/Xn263QmpB2WFjSr9/ae2u
TQvif4xYWOah/hdMjiNYtCH9UfLfnt5AeSsYLbUrIFc2Xq3Wo/bfqQz+GEPxoknpqkuIay3VL+qr
dRoBgc0a5C4skAyy5sYPGGviSLHXeI8xme91cQAxKmjCGzwYXqW0TZcrROb4pWoxVhPDz6N1kApu
pd5dWgtdLlY2NSrMYFwM7jL0sh39Jy134Xq7HkrjU2TtmRStV/++PBzVYfVXZlzmaubTbnbOFilv
1twZJg6fiHEjDVgbQOdrypcnraVR5V7Y4I59x92dFHQPsxJuD5Unk0++TZWqqRuz5cFLiprbBZTn
fXvqsCLHA51KNQIE/yrdJfjNVOjEd+oabhktLEvLr8nKRsfapPXQcOU5n13v2JTGSgdwNX2BrBmF
TaTTn+mrwEavbdedI1T4N1p2H6r1H2KwBMKJMTmG75O2wDxgQQj0/G+usnLF6v4R26Ob4sOnd595
I9helSsClZybFHtiOKnGkJTwE0ZETLo1cIW9DbrP43nMT4fCVDwWs9nvKDvOwMAA+j5cdGX407Zx
IBG0b9H/EwjKEQG9KFTkwsf5e4mFYZzP2WSZZenMHVMPmfbr7+xrpEru+c9UxKY9LSXeBrznM3QA
8JPfoZ2i9WqpKXUSvD+Gsto3XEf5jafXDJ6Ri5gfYqgBTVSasOsVgh2hdmfDbjiQbuiRadikLH0u
plXaHG52kMg639/gXN9KPLM5GVs/hBROhhJZuH7n5ufbdLGKtflhNVAlarOWyY8k0rDiuk2nulKz
rtgMR1JZfrRZFDhEjdcb1f4xPmcd121/XeNr0lPQDMQS1KBtjIi8ZKw6A0SChaKEF5PFN+5El6pX
MS8F/yDsvBMeYe0BAMfctCcXuFUu5BAObnEmHUjMGcbCIeA55ZvSpEqpatdPgJRMbkqHpSbphxeo
fECCtmG6V0sKRDqC9naXSScjpzsQ2fDyAgRnV8rLf0XuAdooQZRJvk1qDmxs6gU5h3g3LYHFfK76
+wU/sP9koOKknoInVHXWPee1eFPtlB6Iy108ETivZUid6dFzKTLYLh5x2/EOccAu1G6CvmLsN69P
p+9vUxqtvMTfgBdpr1f5o0XlheTAPx92z701RgfCkzTdUdOXG4gIFEHfMoEN4N3eg/qmB3zivTBU
0/VaL1q0nMW3MFBlCIoWGxsSbo+Pr9WyRwFwp/DAmTnS9xBSb6/sz6/7xxBusqQlH2qKrVPCyNCW
MZFAsEUwwGqtHG36nfVxGmZzuPgDQ+moGdhUWK0YTcRJaoV+o/zfquca7eE03kgp2I11uNOSKIl3
hjjdJMTvI8Uh+ppEBXNEoL9uDRiQUafZTvtdmmV021I2dEoRIhyQybWfZQmlYM+ZNNzIFed3dDz/
uzfo6/WjVL+49cTz3aNo+VK0AItqVo5xZN6sa5+NlGjMyj62Q8+EHwxtwkLjeJ95kmO6vCgBNPFn
IHHI8ttrnKKDrnWw3NpOK+OwibSN7glR92sBrSDTzQfxq1UKhh11jAknmMmqxaSJBeCU1H7YcnVS
W8a6Sz8biR+ZMya1aFC23hWFmMSHM2HOzlclaXVfAjRkX7t+zJDFkRMkyrVCNKLE/iegPK5qYQTl
jOArBhyPgvAwq5fsRB8iqEpQi7Z4cOLrPQuJGBSmUnykibrQNbX/ZvvTFUkaZY+2Gr3xQztOj0tJ
ASjzpE82ZhTdEsKYOBlPe3AOS62R7eOMKbxBgQKtp1BPrQzFjadmoBYVL98pNBe/u4GFmeh6g2sR
bX89cnIpVYxLLjqIFupYYvGPtl1J4HgYkWbPuZdvrdYE2VKgqVD7ha5+viJsSQiJN5h6SpbDRo1j
tgCngFaymajA/LZp94f9fGpakAKb3bZ6D8X3Le1xBxip7cyd5xug0qU/aW3vH6muJik5S5sB7iHI
Vm6uI7amLKEe4P9k9KH9Z2ZT/+6U265ho51B67oU1AcBHD1RyDCp8wcDiGdujzpVvGZUlanE67Z+
BzfF33oIYgexDC4Ah/9lnNp5WHGt0sHWFVjbOuChWcmcrzQ8IGzQKDLnCbSjUMXBQx9ijGHJg6j2
SxCaX7fWSWcZetFXnsowN3S+/88aaWXv32ZvACgcIeI+H4SM8ReHM589qQUipF6Syj8FRAshetQu
gTIVaug31y07j6k129A6ks0oKi/h3DSLJKyIl2EPu+9Mx5RT/Kx9UbRvPeTVUqZN58BvlfJ3zeEg
Xv0ZvYBFn5eOncNG70YYCT8YUJHuhxhemTU7aKaziz3pL1IQq83KhSeDZURJpRH03wk/VdR7Z/c+
0zG3lSYOK0vbiD1EpSBy4PXSta3e1fjhN0G+FWNilfnwTAOjlOzo0mZJWdadIrwsbs+8SKemUoyp
MykZ7F/11B9EezshzsCSlUPEIVHdZrQ4Uue3gk91yK061B2jTMHZtacLm6F0fTgV+t7eIkP5T0At
uQcwnL/NKMQKKBn44YhKCBBA339g0ilDmET4QW/PpbsWTi8Uq1c8G1JfmHHWnFyvLcLfW87LbkTH
3o2azlovP+fePaX1TuIAbhsB2BVNCp969pJQhn+ZmWiLJohCCUAwSyfo16Y8gCBp7KllA8SniTWw
iY53eKD6J0cgWFftysjdl1e6vOzx9RHZ9vTLW7YpNu68VN6oHM2kWc/tYH05QwP+Bt0dVBlp6sqL
QwmGJPuwg6ESNWft7aznGQMgu2uIutrUwtXpOXsK57y0wHk2kBWeO3rG0oW9/fhsFDw9QnvE9xI9
Lulb4jjbaOihp2NcY09pUY1YS4cz/TzctNxttqbrVruTu6bEob/SLFlv8DWIWHIUDHDJNTHMQRUA
fUMeD6OgY4vk/g6xT9fCAxrFhhADWdqZAFrGLBqQ7IxTZG+YzBFHBmIMS5XYrp/jiwqES6GEbxFV
TsCNsIdCGjn7TiMl7AeDDhjrPZ0jUIEzpsnanruLF9J0E/A37hwjTEHYXFolbRUYf7YsG8xE6jkf
5FhU4X0XQpEDaMGPq22nph3VfKXQvXZH670kBaclXpZ+T/9VkRnIzh8JocTIjObEFaF++TNuEKfn
AUq9BjPxCRr1y759J9EJ0xmfACBQnRXQNvJwZ4MFBuce5CSHpnG/h1QtxGCrEWL4A0A9wmwJbnTM
p9sVwbvJiAX9UVOup37xHq4+HWyprefbgVvhKcWSTACp1D2LC7p9u8QJgs8WCucv0roUHLkAuz+4
ZU8PKkEqHPQ6r8iIYBRItx60wiCc6+/PYp9MuStki+Tw39HhqCbDtDTmKenPQb4DMy6IM6vxC7J9
JxZf1y7HU640M9MZxcjQ0F05WQ1mVjXLxhKLXjpjzY098eN5zzqRnQDCGXIFC5nEqJQUcJ5vf4RB
D1ovDjxQUUxG2uMIUAkniyQ6XUwjuQ5HDQZbIZiyd42jfOey19hEPiFNTlX0wtES0QPiFlY389X5
VwDAxFUvqmGnTxm8B2qKsPy26jvTkPTQzthO6tmgGKjcSs5UMcMWWfRRg5/pXYuVSCqk9EIfARk+
aLIU8XktuwK8rpWcNMEFhCbePY5tKY1CsGlD5DsoybJFigBaUh2mmzGodOSBC4B9naSP+7jMcxB6
uFR2NFaLq3iSrqZtszzo6MEQg88Sp1mAeJMzkTXOfgqHPbt7ygDepncnfb4tjnp6guZZSCcEjdh8
WXA8ENx2eNKC8GNoX3vOXc5a+z7IqRdgFtJbSxRXNAVCgJBaRuMtgcn5op/4EYbNNzf4Q660krxy
8t2g0ncanV8jDAYd8kvWVjtc4fZuVtKsJ4KRmHwqBr7fatgOAC/s5OfeBZMXFZSGK2/GUsx0rAk0
DOZf183LYs6PPWX7U1GX6yjhMeMEWpsyYbvsuPUo8GbcMAN9z1ZQDMcu3x6OoWDKWrRT00mY2Pcz
J5LLzVEGgdTdkByhBIWo2zHzzImQ/Mbuj/EVyA8/8I1YVxt8uPTHGVQXOpzfKlrQ3wF+U5B78GTu
S6zqNMtDGdG+EdVNdvJc4YFcD2E4nzcBCxetWXDvIrTJxc7kEqeSAxUPRBsFA+sCtq0g/6Zwlcjh
MJerMhJWLBi4LFuxGRUoAX9Ig7b5Tp4r0/6fv+KPPCr4y86rUktbD0Tcmku9BzW/pDQ/94lAG/NU
prVZm0ODvtQHA/+GCz6MGXlTNHDmBc9oZz7oYHmJVk7cfG5NJicudIOQ3hTns8oa8i1HHtFE/BSD
rhyzuBVCa9Lbr42K4rSI0fi6b7LrkIb3KhOovzopBIXw2T7v9F1so0ON9nK5zQKMbXHRCw2zT/gV
jm34y+3J1hsmVUD94kLT/K/iP7xRvwu6Bx1OMyxde968RbvQE78CT6Z9O1CIqFvXnRx4I3saXH9g
4wTPQbCjJIhl+WqrZdHnmqvV/GSVJORvladRxemHUvumGlnPF1tgHCqCA74uo9JfPfxJ30Tzv91C
IPdZyDv3LJYXSk8VzLvtvFgV949Tijp+P3IkMpx4/JUm7hYeEw2CLvN7SspiDd3X9WhRSgUitpth
6XM4ZiYwZrM5xlb2lsjwnp4lGEmZqrJHxWszoRZi2cWkhyHx5u9Bz1c1LfhNnN2xZy5NyI6UbKEJ
CzH7x0nuGCFXZGF9DLay6ueM+NFNqXMvxXTUoSTesn4T8XDhiDpFwgnMLz53Yl4VN+Af6tbJr7Eu
ABmo9wva5GZX7AAGi5R8U95GAMxsO3MMGCXm72m4H1OfgAru+oCtchsRCMbCA+RR2O9Fg/10unHm
kjDhllP5nqfgz7fZqU9W8m4Gpb1HxKcApAiXZ4CIujfF7OW2Md9wZndaYLRIuMfOc8pA/wzRpkCi
AQJsLd/+MAPeIKWYQE9IStwFB3HRGT9OuGAwUoYsh39qPh+/IKybxPu1doTO8YIB5NRIis5CvmrT
s/NXAFw52S+rXYrD3k4iWimrKrcO1QZbqh0/cxCTdS/icgrjG4/HwJjAnKoqQjZb3o4CE3yWp/4r
rHIHSSNR8NbvUKL8QHks5IgNKnGTPvEbFfsdJ+nIOIUlaKEJhz9bPwAjQO/DMQiUOepyiDM2URT5
kWFmgutwFU92vfqsNHiwPu70AGbqpLfPA7RRzm1mG4haLbj03BRG5poHbdkXkIhK3R4rWhHvcMdd
4zAn8FxcbSoW0HdhuHe0l2xPQowxS8JmF1uQ0BMAAuD9pcW1krx0vq0HDI1c/4l5xlS/4pJE4u5N
iLW+3KM2/wXfR/KTGYoXJD5gwMp5PCxLolBYmT/s9G/n+1CXMRR+K3hjoyYrCuq/+R46IvGsWYQA
HVoRhWJGs8fd0orNpqSipZ1uecjHKfWLj2UFvBXOxSTUCahDfrYYTjUSRnPiGnig3RSoxnlEUUX2
4pzHBkN/2q5KSall0eD6G/7B9VB70bQV1JvmcNgNombYgYpgg1PxCGIyyVfolsYdhsKJwy5J2ujh
otjmDCu3OIvF4C+iyeC9aRiCh45x1ll6deYn5xLAar/y8SD0YCY/2xgsPRdvqPZF3mzydiF6dzze
2s4BownLa2WvWIFDhjrQ5G6CYv1F8tgcLEHVbJ5GCdMoH8WkTPr3Qt4Uc/qcfwyMZCjekTIhkxb2
JAgtqsPM1m0x2rmG3rOHjebgwx4NdqsccrWhFphC6cMjUeEKuCyeEySIeGCMVAnhyzmgf3hfq8ZW
4ul5Tvsqkh6YfVH8IdO1wajYrP7Ej+LKV+04jG37Z5DMXNGi6BNaVv4WA+nQP0srinpYfY3bS/wH
8iykx3hhrEvVTctrxWOmq0lV5BBwldoNkBlqKQ5AzLBp/bS7F9XO5OFm6GIz1vVStdOq/WrKq1U7
TbLRukZuGmuEytG6frn7bb7dFfSND4bkOTK1FnZOicfSGCaKygi11fSZYqw2InTNrj4L+AO6Kk9/
EQ2im2IyvDdyU2/q+znDvIZeaGXFkYM6BOxXuNsZZ/o6xFanQcS5KJ2ueZR1LKGLOEzAA38zECmq
IQm3/UjRIqFJZINRv1cMZqDV4/WW38eSy/9tTUEPVzcyfUr79gY7ja0XEeiovZtUMVbLMUH2XB16
5JsTsYlkVvn2D42XlbAmCktxTBlnYlBSxuX5JaZBoz4qc9Zr7daysx+w+m3hyLP0BhXlRFztN/ZY
4wl3+zmYdiIZ08p1AvQpzdmShW45wGct5KVaeeosKEWgo0nzRM8S0wgMEw9+tkfG54FcpF83sK6T
VaKxa5yQWfumTAcWxsxEqMIeGCL2KlgAbBP/lySmmwSllrPD0MtCQiqkcmMHct9XxsItHDxFrUT3
4/aogNhhusSnIuHBh2lI1AySdURruaTvp5p2EUFPRZRWCt92cHh+O5oTD27Xoe1cqEEQLlU+jwND
cef+BtTkLhMJyTuyxjhG+mk7WG7IUAYG6t0GDY3wDeLVV3F2lmO/Xbggi6GHTBNWKgWqOz815eY8
P0WTwXKLoe+mIZjiJB6vtfe4nLpXLqjyp3niskCmab4yx2nuhdNNqCEPINplliq7De9gQOZQlh72
De88oOdwKkipT24eyHkMAdja5kis1ogSdbvVurgDng1Jdsvym4PUq92zXGMxywb8ixvA63pGL3Mn
jw6ZEvIUWgcj4fE/9QBfr84jFIb9qweKcNo6FUxYLUyJKloPtftKh7OiNAF4WlfPzipDgVSuS+4C
PYTocC2yqCuiQORouoGYVY+0CjtvvRW/TYCOeowWjBbX37fcWR9jV79m9HbRjTTgfmyDmHvVKFch
Zosg6ozPfSD3+2l6aQ1ans/wyXL63yeg7lXPSamaUShZAj1AW4wp7PebqhUbOdzj3qUlnJ9OOZ9q
CCUmfC1+wPqtEeq9AZN3/s6Xzf0eOMym0OtsiJDJybgyvTNVBRvjT0mDeOqb2Q3BQKgwiHm51vBP
w6YXXsJCAIl2mh35qrrpXlwX4GJR64hV+pF7CM6uqKf6shGsgwuJGGRQYqqtkbfifMn73zssEibj
ZgCRjfhKSpccxXx/gnHM64r+mt2WMyrosg45HhaVVDQ/OVkDPEmv1RkTHyvy9wMsXjGi+nXk+eRa
IXmHVj1+i/RJgeTpbHeaREXHt/rj4LkXHozM96euvgDZEf3+qM7Mtb6qmSJSuvisW28AvCLU9RsF
3tJc3sgFSbrcMeeHXFLXhDztDmK4ZW6XU5pffurJA+JsVuH3htGNGlEeJSz4aIX5j/ZCJiH8BRoT
rDsgEGDW8OeQimHDkIvpZ39Q4nbCB4JBDail5FxUfeb1F4bCfy1IO4yuDm6h/gP8lARsdIAG3tzg
IOa2lpsradiq/ehgHcnjB9pB2DEqm/6tvt9bFWSaz3sFog2cljrYVY/tGEL5noGOOxgVaqL+vmXw
8V//+ft5wBMKgWhZwGbvAsQt/OTDS6EKyZTpH1W2oK98VB9yhILc66ND+N0jzsd4E/RRUoR6OYnB
vZ97gEf8rmZ1s9m5NSXMWhnyXAICHJD3p4gCKNPpel7c4UL55IhPLUqUcCVkT3DCRKKQkTMOF4bi
PfOiQ8Xb7SRqAOYyuLsdrFprGrkM4Ts8DUBFeijkppI9cbWXv6kOsBKYRwZhGwPFlWZ+ZXasR06T
axaSpH3ukHOKFUWKb54rHlUKWyJSsjXtuDmJHnbgFVo6jnrK+XEnYdhU41Mznws1vjitsUkBaTYV
pC7LVt2j6BgwftRUSD+B8DIvyb/fX+v0atMg2HLZ85w/KkmOv+jxad23FKjWoTmuXNyYsEopqRM5
h0DBhYnF4eH8prbmqLwHyPI8ootFcDl5xUB3fyTXP3dQFSmTApxNlPei5E9sg0bitRU1qvqQWm2c
tim4TmI+v+SG1Iu1sYOKhzughtCAV7VxAMWX/Ekibiy3RmpMfMNX1bKQFwD/PJFUKJd7RKQJA6Sr
/147Xf9OaRw0pibkUukyJp1hr8iLctpbZ58cWkUZWBh06UDlIPBzkmuWWDTwktI267cySMc05vLn
wFkASZmbZWnZSEjsKe9QXeIanhBMEb+gIIjs7DFg0NhTHOyQ1o5hp082/piOJEPBrWWkvdFEaDsF
sw7hV6mW2OP83+VKa2mA8DguUAZEU6QlxbsSBxcTaYFcWB+mW1/To9tUv+D8vMW2NUIt8okYOO7y
SL4ozLdhsHb7zeDR5PbN+Xgpc7jpiFDBgRF6HjgY6xWEPBDHPpgBxbDRZWinZCkn8SmTdO/CzkV6
Pzw4DuDdsj9G9VzZZyLc1v25nNJxO9fBiabjqXs5a6KeMgjg5suElIDCLDGzNo5N7QHPcd3ZcAg5
q26uEIqiVzO60jUxFxCApWFKp99rnw0VYlUANQloAeTy2kTgGwamFfT60lKZghAjprnBOLHNxZum
o79FLsf8QmYxqTZSHA1258ZEZQ01efhttqMtgMXaJdRzKsF9dw59QhtPKz3l9J4yPKNakmVmlByK
dyI1gGbranHRnhEbBqC3Kmj7ZupAp6NTh49fk2LoFOB+BPlzJNLFLd007kDWe3eadBIoYSBPjyvY
MA8nm4u0IqhEy5bIYPOJSlVwwrRLieURM1GwWgyyoXU0s51kLLaQ5y9iyMXOuWZ8LllNdIJjc1j2
7zKyX2fRJ/C3TsXKKuz5qp+RGIaxCOC5ilV3fMuMGgNT/WuyDaF5le5dqd+B2aJbjN9LSNophdzp
usu5aaWm4tJ/Dnut/vehC0I0T73wV5XTKAcpv3N5gz2Q4w8cYon0xIvlSWxrxapI0S2h/J2zplaY
6l0FOY2/61aSgms9nvh2+EtLnkH89aQ5kia6t/xNFixtuNdVXRE7SVsycMQP7Az464PmKLQlJqd+
eSr7bFYRQ5iTzXtOodmHaEgElml8DEcEKV6ioeJKlGSdjbZ1nM/a17bLks8cUOvyj2Ht7hMcITzG
xXD2mDNP0Na5Mcc2/AgAj1zLxL28KQOPYfuzoWZ65DfTG0VGGNWErz/ftvOG4a6F5t3kqg5NkRzB
o1oZLzbTyqN5GzzncpbwJCsaFAK4Iy5sA+qKpUhV775VajyyMvF3B5Cmsq5NS8+QBKCfLDGHMpH3
gZMKvu8YNtWNULbYkSxphmYgOTUgEo7ZJboA3dYqhK1KdUh2wqDvvTyuPbQjd+32U37hzit01flL
oenhDLSUji3jh1IaR/UQbN8A0TGjVH7NYNJc0RGp2uW2RryBG38kmehLQFAIe1WAKeZvfgGrK5Uc
qocoMudiOJkAIRbcidql9VRIHvXZBVBtFd4yc9LIYXIP92HsELED43eDGTFo1H6bN12+BT7PuGX2
rjuGS32P1osndnDDhAI8diPcHijxR+LJ9ISJkDAVZGWNze8XSC08lDZZuYyDmT0p8eR81RX2zPu/
KHu61/mZG07w7PFzu4zxhTDAe4IHTFJ6zGndN2OwSNnxXVdLZcjQ00SRi867gYHAIJWqa4axlFmq
kPYf1/gOqFAyAJbt+9zlAniRfjil79aXEXYYawgTv0QVrw2r5sKTsl+5iMyOxGsNForsX3nC2SmK
ykvb8tvAK45hbSxgkOxxBdLNdjHcR075NlEmKnLHedy3Diz0uVnLgIXuflgNNnhIDJep0yGZoPwq
flU8heX8Sdkz1sUeM2otRO2IfmMb7c8rrKP3M+SRYWJ9gcWET0rG2XG/FwCB4J9OgUlyLeZ610lh
ttCy9f/1CXTpkZ43hZJUdVX36VVDZRHok2wRWj+LYxckJLUBNFkupZtBWf9qfSFWLRYwVR7aeB76
O5f0CuY5J55GwdO2BO4QrQ8tfnpk6KCMgH6zcoi29eYw6/ZxPfeui7yhw3FI8uTCOk3TriXGOEMu
PWi8e1ApeiVm8bDn7aCh/QcnhFtv+//rtmauBCQARp0lvSsjkQ3CkZLfJWn0DsZXcvrrtng1zK54
S5J0ImPiaJX7Sl3r3B7cdjC3coqBnZkR2uTfkaYzIt/QSDyzHc42vT/cZL6Jaxuqit+0jsisRSiQ
HIzZt/rbXrELMZTGGMl6shYzIu12m+oo1fP+eK4kt30EzMndY4npSCWMe6NNLvG6iT94csQCZWRo
7zsUggr8+EMpMnMVLC5OCoUL0r2PlpmDvWRAxVCe1Gf0OqLN7Kn6nR0/qAclt05/mD7xnjY71+NB
2qGe6pormN29MBpPmUl7jxcFcYgfbKYeL96flEiFRgiWdUt2IcQw8SUqhmAD7UZVUvBUCyvbXI3S
WCDAIQfa8p5aU+y2Fwb5Ctb+O5j8jRZiaVAGmVaZHMKeHpvPIavFbYzwziVZBONlFCRTXJs0fUFk
0GErb8l9tQTFzI8zKI4AQm0g+wzkVGPk+IhysLJ4ZT4URf3kZVUUunuQYqUHPGDZlb4jIGIPpBtI
8Xk9xCVKUnj4dPlOtmf9EJlFlyvxjnmsO/rzfsgR1Aova1qa3dJRbbAqCPPNB3nCQclXIwP6K7YN
VFGJOPOKJRaBkIcqRPNwNEza0SYH15pAC37EBLozrRmpxRQMBuhXM5BEdxRdRxRV136hfKEGV8BR
YIeeHTx5eB3tavZe5Kiyisn0wumVY53OxHmOb2evo0ftU7ipMhSekIUZ2/tvlA7B/fzK1pBPzM1S
SINh2/sbqAuSRsUm6knTtmLTUjWsUBFIw9r2J9q4hB6RGWM8GllaMIhIO2CpvvcyC6YMK6Nml6Zp
o2/m39PhBeCd6AUiBzMKfW+CmJEDASWbC0RTGZTtkzAUPRJHxyUETG0b61HN97DvrNLhXRSLKjY1
YE1I9clZpPpNuaS7KhCF3MeWmPWY4kakMbe+RYghX6iobd8YoBwv1JgqtdsHIrD/s/hBSaa7WIib
vSLBHykOZSeM02HiM7r7lNazeHlSVFPvsIHXDVJW1ZeAh8KyEpt1aspDC6wdZbtOZQooTtlR0wZ1
x3bQMQrQEqN93pfffg6It9PO1dica8KrmJN4rGxgUzUfBsnktt3ZMhAmykD0sNwBSeR9WD0/BQnq
cy7mIGC0N+q+WtHVvBSBxd54AhexYOj0rcMTaWcjK8AcgiHSJ/p84vKoxSA9rl+6mM8ov0AVp2oL
tC61ctq+Crpfnq8zcOD+O2DRaYWoUKcSV/68GnAijRUbufdb5cq1VZklqSkw2lI7jxE0YjSMlV+E
GIcQNp57c6T3GUZ9wDgfg8X7KB2IljDgLCCF/t7QEnaRKLP3Uyse5BSEWLoPrTfIuG5N9wBideFz
vH1jZCM66/WlT5PC047XnTlOxmHs2ox2vztrqDDBo2tFAf8aTBBGuV6o+f+qecgVWwYNZiDu0rT2
Y627vdBWkQSLMy3CtsbZzojvQf5Xl6HTEFFem5ZUqTZISNgzmy3tnq1Glf+dDgWXOi4iY/09IG60
z3NgmwGR0mg0ndTmcXrh8UjwpOdj714QNYzcVpJA7bynz3saAqAGNyy6Ok6y7sglARJKCIVd1KxA
t0o1XoNKx5Hv233ht6VCCGAQ8FXcFLO9PdGKNHhRx4ZhacKrTfQ9JZcCeK/PVjhG7oWLrPZO6jc/
eFMIisAy8PY0xEcS4fVjtoo8LkCpHfcPs143fsZsTWUFk+6SXosWUG9hdNkB7pEV5AhmP5PgwzSb
spJxvqWDKYzN6sJIpsAZGiwPRWImpC3/3SIsjIYYboqHz+phxLJ9AcEroxvk2kHF/41cOFvUuad5
/QexeJ/1uBGkMFTSZutOTaaD7qcOfZHu1Y/ggSgMT5VxtORfzhYL1YGbbUOMMuOiNoLET97YfcMa
DhfZEYAdOyrZODOIHRNvKRQk8yGbhNUxlfy7wdpQgSLG9DXNSSxgAo1Ah+x6LK9MhFSleyX2+hPu
pFtKyscPne4RKm1H9xGJKxDZFdVOl5tm/KZU4udcFAZHy+a97C03trC+qb1UZAafWBcHNWEPs8VG
ONhWny6oeMdmcu3rOrpPSxzuQIw2nWFtUhLbSoSMddfZr+8IYubnuEKvdwpPi97ip3rRgK2KdMgQ
rGKKOcIoRb/EShNwxwuVN/6TuoBD7Nga5LpiHsb5QODXQ1nbfOihDyvA3dbCVm6PweiliPQZN2II
1VDYbuS5upPIOfDPW2jAwNR2vVfV3JrkWQDFmKoBJjNIeD8Yfyhbvccx8cn4WE9Kt0RSrQN5TuCZ
u8hGHOEYDrn2oNKXIh78TdKNtTs6GdEieDkxu7IaPN7oxotW0cO8MB6pHk5DNsHsdOq/Q905unbq
Chuo1vlJU0Enhol/xAa00UPd4yE8A2w+vRaRvqGg0e7FvWVD6dxccsUVJlw20rO3mPn2Oposqmsm
OCjJ6WlyZaMVTcJkrgk6vdsn7Sb3uWcxp47vkvuSiQXiJdnFNVnE9gskJnzXzCuRQi/TW2WyM4mM
vC3XplOyXNwjUBgI0P5cWr1oAgF7xNPftN34p7aeTe7eDn40B75D/mi0QiYK0Pzzw04VlAVr6TGF
6PeeLyUi6MrO4VgZh6dU0qcziJzuLDd96yvN8NNwWwdVo9EVM6kifoDgefDhlEShsOBi2YZRa9du
dXZeS0jDjlLIBjIxLPzxtxSf6kwIpJw8tWTrrDb7rqi6eLmorlOnQUEfzU3TNSu4iibRvEeftFMG
N7jZZNUphcL3MRuxxJoRvN/++6+K/WzZiUQpFTqbjxaxjDqijIW+oP9+05zG+nj8SN8q7TvXpVeY
6/+GlhgVFHRpTnz0AdR5BA8ggmGaHsvBhXrd3gloVYnVffLtO5k2lMTIjaUi1mQWf6J+B+SLWvYO
quJWGwALpfxgROgEkBbuBkF8KnIbeDMGPmL1Lcb1MUBIs1n6w42YWSCSOL11iAxszZRnTgSMzWOv
8zCkYTH7NihOud8oatq6zaXMYFgpAw875TiQm5xtV0Auo7mN0lbonZlZqLpRGK1G5w5PxaNl1h7l
l0M/B6/RCVW0nZrmpCvSdhgXHRUuhmsVfA417ocpb+SjPj3qCj/Z6XnXPIdpuK+F2SA+lbNQeGnB
Ekaf/x7dfBRftviK4pHSmKXPHXxIdK4ulXOEc1Q0JqH4NUWoerl3aEdhZ+nOuDmbqYvYBrfUT9PZ
sth88UqoECnhd0NpahKkZdSfw0NmvWr/u8I3Gvd0G1zVRyHMmBoo5W7jkkwph2O7vkdKaOEwZuD+
ORX86V6QlvJ9vXEjvIxyXSLBUKetjOWh2u3Jv0hB1capZUrptaJRVpYnyU3w78Ehtx04EtIMn+2j
m/BTjhI0A5HuCM1HPBcFuKhpTXwWjh5iTw2H2H2uTnnVgEXFVBvUbaqryJqkXPBrlvYBY8fbGR61
+R5eu/iuHrMQ42QmzSbTcLuS9br945BwxJ2bGy89Y2BflFlt1Z1Njs3vxgt8u3v1yieBrYcDgi50
7E30zPgPRavGgtLFozMEMEH85JFZkOL6cpP03D6iAKUFbrUqHVt2y8DEcCchrnzunia70tryoYq2
Hpui4wualrw+odPVzbHlFtBsrJB1v7nk75dm0ccFGNi03uv3b1BBR1ryysuQtMyze2DvVU8xqq1P
teGUv6MDNRXHs1xg4qWoj587Zrgaf6Lf2BIC6u1VwZ8HPT82OQKoBv00OJH9M5sx8qqn+iLNKvwW
FaD9NJ8Ed/xNwhQd4k5tRllFKCAZ0kka16FOxhp9b3lYttsxmrlUrAt50cjBpYhLzPKKJdun8wgn
gp+lrVOkkRAOkws6D1xvBet+oSM9aEYwPZ5a5UjPBC7vPjx9aMvz9g2FEnfcA3nWneTlioMXgmkz
/DK/C5uIDcyYH9zsOAdjrlziJAvMD4rVcgHp59kbNHhL4CGFI++5lzpo424287GEyJV9BKyMygAw
dknnhALevjQXcqTqrsw62I27miszJe1H/shd2oZmtMjkYRurid6S0iJ6uA+pm13UlsMTRGjG2c57
q6JZD7Gs6iwwgV329CY4jEjypRk+SO/QAPTFdhsbzDlc7V57dxv9vqMaL1qR7UisP4x0PWPbPchE
ggqw8oTTcjK/9dlFsibpJ6tuzpgHyEqAgtt9yZwyuCSBs9zTpDbOKP5OX0OPUI4QNAgPMDPNgeuW
AcQrj6nHC1MtIQcMQBXNSQyGw1BsrLGomhje2v42JU1zhFtlNgaqck4oHazY7Yckd/UsOIpwzos0
e870v3MhTcWecO8X+83KkJyXGAmP2wmnzh9Qb7SDiuepgXAycwKCCKHEvnOqR9iw8ysCLDoAyQ4X
nYKluT2Kj0W2TPTQ4uydeLPMULMa9EgjploOgoJMyBAsFya4KwCkvrO4hggWaKQmulPRoUUzZ9pZ
63HQXwom7hpz0nMdWDZ0ipcsdE+9aZL9KxwAN4DqIFtBmwMvYGTe6wwEd6ta/QtkEpXxoJvF+eAi
EfZ+BO66IohbNSeGGlHyLzMoQkO6E6E6rnYKwhWR9yP68HoFS2Mxa/CcIOsTYu8w+/VI5FIm8zDb
aNaGEFKwHAuAXr2Yfmr5aM0OqiEbJVtHlDoD49T414nqU9fGnXRJ9HgxAyjXaj72m/N1nWpcV+ed
euHSNy+5vZDcsYlQJvaJzXlNMOSCJ9SQxuoiRXcW+FwhAKuar23B2jAJQn2yOldSYDtk+XHk1ZR2
1/vfFRW4VDX2ibYHUY2PXKM4QJsXJRqYHGy0SLBPjkDREEMCoyrBNNncgUmDxZ9Ha42GsAFaR4wV
8XH4B51A9k0cI2Sxja2MkxFKr0rvfilqKB/HsM9PbrHT41lYl17P7sDALyrjYCtTHBEYQ9/3lVyz
JoPRJdhiHYOdxUg9W4YPm/i8nAY7dS7jyvH5+S/vfgbN0X2trQjXyrIP4k2pHsv5HgMbv2AEhv6S
fjjphWPLJx9qqEDi/xmxNEwipX4qsDRy9Y1K5DNWmxQnMf8cOPR6nTnCugABow0nOgdklX35CAfE
ek8Xnr0xcahm5ofNuu4XS6IUDVoqsIudH9CP1o/dDVSKA43FsTHKFK3VYO0u+wuWTdWg3cGNek28
sBpTjpbJV9H5SpuocMfhVfCxgK/iMw/KnaDytDEOG+TcqkJVBDaal4aCKUfEhqdQegNHiBJ+CLvt
bLY633Z5EwMP54HsWTE51/mjB69juO8oJhWVDzBKZhPY41AbvWZSQG4NW72220s+fl2U+7RNy+or
JQNEc1YJ6C13FuABVIPZ2HlaNI7quRyXC/MxAd33g4sWHSwYYx7t8gP0yYRsIqP3QZ6gy+XbPZrB
0y4+E4qYc59dZeLIq+c3hsDNo71enjj69ZR9P6rnjX8UE2DZnox168y+BMSP4llykpVOlXtb2gP7
rPcNpvmJj/gB3/xn6+Wt7V+uLChnbG63gc7e+dKIit5t14gF6jFKUT73UlKEgWZKIercJfTgPkiB
ng4wbJYtRRVPA79vcjRfKoccDewDoF8p6RWbfGIJ7E9d3NGdUL06oiFwmHRj8CfbY6GjPlHmt5qm
ABHroq2EtfBpnqRbJWjE4haVBiOyucFI0oauFXr5jm9KX7e09cOpLOu/G7q80i84J6dcSHielQin
LSx8ZXQtTi09cTt/RuJ+g2KPUdwBOYY5gmSAizZZdukrCkNLDK5g2tn8CPGi+AT+kE6xnuKM7gLr
1vOUWSAF07G54qBLam6v5rYj0BF++7Ao8oXHgnqFMUnMOhXg7I3gwvoMdf4ETCT3/SPHpldbPR7O
AXDHXzMthFa7hPAeJi2UzKEe1NrrB3lgZF8HUxzYQluvzrxS7jX7pmyAS8hdsq8F9+RAwfZ8pYW1
4PhZLzWXFmmFR6U3vI65IS7q4CtiOYPkeeaboOOQv+jCn+JwA/Ij35m+YvA6PNCWHNz99gHD6JEg
NI2N/g7t6SZWHOiLewKqvEfUQgz7Lwy9anQJT3DGVLJb28GMgz25EIG5dfiCKDMsqzC5aNiXZvuy
rxBw9YoxQRbUp05w5fs0b0Osx/GXZYAdj5zWaFxhkJAbUn/6o7mR/WVYaGH3ztoFDGD8JEhhBoM8
uPw/hV4gOpHtFgMRENL2nJAF7BS6tw3XNdCcmd3xNPy3osdWmLVtAg5YltNSh+zd9yrmzQ4bsiMe
A0RdHdNH3BUX6FmOUs1jPlvTtfRKev1yDyk62W2azbiCWxntmjWe1M1ULoLo33ce8iWpl8h0CzQZ
0k9JMpkR5j9NA2BXKpS6NbgmL4vpYu7FWEoCczvpZz4ljvIdE5ROCxbM7jtmZPweJaVD0/KjMgMF
9OV8YpNF065/8EmNoxejiHP5aWCUOIRTtCu/GH6VBaOmoQP84pNvaJyxKbOhXc0wqrlU51JJ6LPZ
W6i7VM71WY6ulxodl7o+p0YMmBU4jbkfOY/kdn1ssiwYjW0TKhKl+udXpwl25mpgJuyVIPKjiJ2D
SpYt2vYwkcJSjWri0EO75+iICNGBpX8f6djV35lA6OVIuxsVnEYjHjXGeydHs6KmyOoUVgN505fK
weZTIG5OgTMG1nxbx914HmuF5zoA38VnoAcNxXDU507OWZZVqCsBZW3ghxT8fNo2oHr4GzmmFmfD
Ehe/w3JOY0b0EYNW7svmGHMsGgV/cUY6W4Q7RqqtslWZOfkHkfiWwz/uhSBthpyTwNVjKPABoOsF
5SFoNB/K4K0qxu8Tdjc9uKFYDo+k789cb1lFL3roD3sVsDjvicCd67iTvLePpffpc7A1BHl4Pfhe
pxJpt+mjoYt3j4jY/j7NDQLwUmjpBwOo0pUYxs/dPW9hqd3CdVeUTzFclAvBXzxKkpm8aZHHQQk1
G8Yb7DDgEwDrLoVWjkU4uRjWpt70ApnyZegvZjhCncWfh1In1m5d3GPR1Kr0yGVh/Abu5vi38AQQ
olnMpCpA7ga7y+LzQjoysoQOKUUnB7pNlvT7txk/D+rwqnd9oyQhx3NOJfJpKxul2ds5qoWkfoKW
NyJ6d85pJ0Q9Qz6edkTS6U8XqmJJVvarO4yLVPzj9HhSYZPcqKAZOaTUAiRkzHyirUMXWsM1oNWH
sYSjHIkM1L3myyxhec3rmFjkMG7D/1HOVn7s3kjsCJ9kndINv61SxJaM/9XDAaoR2kBYRyn5eBBX
3vSW81OYjALOWbTm7+dcAQbmBaewn3WVAhUtiBS+Wa6dTs4dvVcQX2fUR2X1UjRdBu+btdqo4VnC
+ulx3SnyUnFsc/2zSL/CydntUnJC6jUYQ8FuGsXKFBonawcJUDvdAl5BsnB7IReFjziR/5cLiJAn
6LfJ1VWhg4YbJOpIDT8l2nHEWglMMBQKAQ/EmM+R5/N96oz1HJ3OAQUXL+vAT6lqwJDRQSURebs4
dRiUbMXoZ1ol2Db3z0UiFZjGbiXE8c0zY+Ra9nJhXXq7V8725LTysx8yK6S2V0dyQe1kvVoPry2a
J1EvB2w37AFPApPoJTln5xxQ4GRgpCx3nkqeqhqmdKyE249ZX6hKWcDGNvSPD9+MU/x//vM+C2fD
hNi7r0+IC1aiUACA6yA6X9ix1d2o4nG5+Rlg2JuN1p+jIw8YvfyOV809+8ahbQVDatwsiECYfPCp
75BXJORmsl7/KZ/GsBQoXqHuj5EmpW41WOpiseG2S3Me6graIe+RsUslBa/em3xL/+KqfKhCH/Hh
EW7lQDfmHzL3RatDxBZHaX3LsfjiNdJxZLe7cHv2RnvstmAXaQ8KGyxpC1rp8vxXgA/y+y22TksG
VsULtGlqLlPj48FNWOLzdaHGdwnZxJRtG4PnGJWnlNoLsxHN7iUSxiGOzaH2vWdkDKRnEa1ac/uh
iI93lnE/h/+8yyfjuzWA/X1w0W1W2+LXiYst8fpCH+0IEsntgHDp/XJ6SIKi2IfW4OHV9Puz5HGn
ek3DF7w5faxzYW0xwf7NAhXr7f6p+bNjmNBSSuvWKFwelgn8u5Aa1ISFXShPB8VS+ILx9+9ZWQXB
rrv+nFROXEodLCkjQYy7oxbjVdhQSvTYEpP5GaNhsm2SZ/L29T9AwwP3TmYd7JeQ8n1vm8qFH494
HffiMOrTE9HZZDAFZQyF8dZIDWEH6/7GC1GaRjFY89S2JSJbsEzWdtPtRphvXqaz+non9VDlChSy
n+2EP298Lh5C/jQTwGEwoDlReeC3ENGadZ+iAlgEaIusDKqDK0HpaZG3w13TAebb9bmBo83juAC6
WZcIyjg3Flvq+s+tMGhSBbKAD5PMZFwJAb93TYwUueYNuhevhTk+c7Ul/TgUbd3YvpjYR92Uj+zt
02/+8dx/HfX8s1/IUZZS08kHnYnGw0r2P1EJPah1oN9FZv7J0efubncY5EgpIWsBNR0HeKyq12Ji
QRzgXInk5/F6AlKxTJfxBb9AcEAcyvOq6FvJaB62DIz+c2Kd8jGhzjfDf+5EhAX1oyfewBlbDulT
YyM+jyT8eDFEnrzWQTNn1rGZCkvU21H9LNwyR7ZvEULzhKJ9eYVR6nm4IN7PyOWPEcBmOLjKRkUV
gOf+ocuPKxNvWs3LYPwjZTb9Ds+OECaAdPQcxSn+nXuTORj4Vhtj20J0YCytzqZpkAmFVpwtIP1T
qS0JnSGmYaj3OIqGIR4WU/E7mY4JVoUztvBG58rcUHqqe5AT3WDYqMNSNsvPOCge2NfXHLJWhN3p
a+lQjRcqq8ABq1H3Iu/5YQ/U5NaGTQ7Ay+mborNyqun4SaFUS7UZY8CDw8P7Ttyf1C3Ql+Q17nEe
349csSG7/BCj3C9joHD9bPDfri6NwL5Ax4Ff2zRT6pjA9YbZwLxPWF0/rRslmfBRAsblHC91Px/O
QtHsrne6U/p1fofPQV5oUINRnO/U88q/vbubss8RV88VlXgNnzS84wGZf7rvxx7I93eFUxYQWtAI
gFwQ2fMyAZhDRlHrDiLlDSC/x+MRrydFxC00zTuG2ub+QauMtLlWiELPcFFSg1EBQnfOlgsSL/Ka
ZIvtslHbC4WgXnvsFMmQPHocO72RGl6SCmXdIromJQpMKbk9aQv6n7UIQYM0CoStLqcCKIAosBeC
7vYovgAXzl1QE5RLVto+P6AKyBs4x/BFjfzdjeV0IMg98RmbPI9EhjR5f+94b9HLH4AR2dEfmxAR
AxYh6H/sn8V99BreUKaH2uwHhsjANRG/f6xCHGvUT9oI3KVaan7YHK9PgkZ27h0oBmT43OkLwfg+
XmP+Dt2OtKyDgUihNS8EOaVsMkMeBDICE8dF5pGtXDvZx3eiKKideUqU9TUvC2TiDZnn8eW1Jmiq
Dp5gOp1hswInglLo2Pl7Wiu0suExykkfLdYoAcieApmkN+xQvJleL4zS5/xzUfv1TwefKtKMxcZv
YH8ft/w9P7lYUyxq/f6Pl7k1Iwytbn0IQ7WNUPoOTcsQ8tijyiD1W0FEaMq96yF/ddDodZQlwY6S
H2L+bTKGNFTD6WX7jwD8tAsohSskHrMZN7TWLen2nG6VXL2XASAaMglrYOghkdWo7PMV9UykGgky
ShLfBl7uvX6OHmZgduG297g/o6WDpDW9t17OhvKLzMkHaPj1hotqmDYGpl9wOEg8h0Pf2l8oRXbZ
f27f1Y0Zuv/vXuMb4yoXzkfhhc3dobmoEmqK6T1o3UzTQs1/m3Z3lWNpHgeX3qkpq4mWBtSEhXdQ
WWgWu73a2qN0CAg5XD5RO6eBb9ydu0r59269sjQ8dAhNug+ZNzm4YaHFLqFuZ7gdsgnqW6nmeqSd
8TyHYOFeNVEVHSVbgAFoWWutkZ6qEbECye9WQ9L1xSeh4sX5dkft+NNIT9Lbv0j7hCIWVEy3A8xt
f1a5SlTqgZ2aVsOmd6JHwyYdmyPDLNt4r1vZ2UGBqKXv7ld2wlZI6d1P8d9KdA4xZMDbu6EW8SOD
bH6ARQ1jwySi2mtE8+rAntkvaTZkbf/gs7n7kNOM602FSJIf72u2ac6DVOMtyKZac0yb+mK/DAYD
No9p9HHKcdhP1zskpQ7o6ewtjpgX1TKKWn7XKE13cVBCXbGCM2xKlFArVPrb+y0JQGeU3QM6faWE
uraQwtrckysDrcFr0KKvxRKPgXfRWYdqGThi2kWRydsb7CdrfwzDRFEE8WiaYWercnmhrYT0pJ1S
8K9JUKte9ajcHqgueHDC9dP076JINk4UtgIev8RLHiK1LEhIhnsson9NhVxxCXfROUbMnwe/W8tQ
nQ2KxqNdiCv3U06ZOHQXrpSqlUmUaqdYMFrYCCDU39Ij/3UCaxpp2Hzw1PhRD0vDZPyHrQnKi0bh
VpWzq4AYihud4o+pwA5KFvZ6c3W7AznM68/616ImEbDiL3b8ZdwZI3z3ZK306fq0CGUyyRms+uKX
97fZgSNxdPea/Ji+qGFC2yrsfMuXXlzxasne9t7kWcn68c/pNacVJCrREL4TclYsK+dmY2OFrBNd
llDMbWogXSw55emFpDrHoGClSJidKWzB5pPe5RA35F2iYlUO1UNIYzvPWfsUiE8MxA3ngPGRCfqI
035HsEdG9I3WwRGRR3rGSCruWFTUqDdTGhYgXCQSK0OeoEQmdORZGJHsLBw/c2YL0OdVEakhUlMb
hzFk2hQ1RZJ2StYJ0PO8NISRy6y6C8JRp7IxGgzI9WjPc20GIA9DEQOuW3Ns7hYiEWdsWsaEytFH
ZCQjHrxIzoq/hgM8vi12k/hYNKPB7r4S5BP6FTOutj/PTSRapWvgysIersyozWv60QUzl1xYf5s5
t0uQ+MNUZuwZBIzHjwZQT+Js57D/fg41pcEhamjx8XTeSo1eI8qL5dueKcbpXuFdna3R1wLsvnvY
aiP2xAuJTcc5q8o8c8ppAE/jwkW8y9QNrYdAe6u82AjoQda5RYBR707/f7ShutiBDSacPufWXZki
4yxPGfF+mE3YeM6Hsv49wwET02Xo77WDTyG3c9l1xYo/p00rS5Wk0x5t7ZLcq8qV51lmRLJAw76x
JRbr2DafWOg/+C38y6jI/oazeV3rwyyO/Vj/egKTlOiC2xtvKTc0EQ+4ObIS5zLgUpEmln2uDGtW
H5D34w8g28nn9dQcjT8ShoGirCkRMf5cP6Nzh86/uvUR/j4H0TqDddPq+ByRn2t4A+e0+kMxsux/
Fpol5WBKUquF1DImRV3llzwTeaErku3jtB4W9wNjytko1EfOJrxDvbiuxMVJJeFCZVcpsV7HiKdv
n5Q43xuXWERlGqj0ph5D114cqPGyXeN9q7kuLom4ecw0mJvtWJZa95rKloTlKtrKCcjjxVrtpP4c
wM5SKiJOLPd5ZiLhHXu0mbSHJGmVgpbrv3ZDE+VQtSAVpPv+OVcU/HjqBzZLhRRuiGwn49GhBUpo
QO8cQw7cytaMShk/v/bVtL4U0LzLN7I5oFSmDfxu0zGWWXpWr6nxiIvvSRg5IMhzYGtQKIOs40lg
5OD3lTwCQmYhhfBZvt5yIGVkZ1vGNEpmqLdwUpPdQOUZTZVoo12/vjLlQaHDvIB1Hju+8GzFoY8E
IGG/JviMTnyps+5temsxa3jSkRa7uWDi8lE10LT+zm4zIQZTuDH4ja9xB5znmpercYpDPZNj4qCq
aJbQzTm4MCwS5SqPxhtvCheHqCtLkVjHKNGTgOmWRTMXkAy/oyj6ejr+LEjaB+c8qQjBcsY+3NEr
IqG/m2lolIpN5QYkhP/YqddXy/zvT3/hlZ3NL7PI27YSMT5rKpl6773aLGcJE3tNrAnMFw5VZqGL
Sjrv+j4g4lDUKTzKjTCehMxBzh0r7f05d8gUjwweFYKFru7YaQMP6GOTe0OiYJTJ1mZZ8TD3GYwW
Ejyj5g0fHIirpYz8Mx6tRJjnl7fcKVzbylOFl9ScmFGq3PKXr2HxGl48YI6LlMloE97b6Q6bi4qQ
bIpKf/i9pjv7EGr/UMu3c+7ONKEdQMBxXj3S8hQpksUZSAn42rnpVEJIydE08l0FQM8TBSEOIBPt
MH6CLERCnzdc84+iLz9s4mQGEMcliSpZePPZKbm4EK25DH8SbNElfS1XbFrRUXM7fVIHzC6gnPev
7K/EQmnKvpd36XtdYP9IfLUfajl5HXy2z0LOw8HSilX6FRWXqgpwS85cY1Oa21U4lUi+1bP3zEuB
7dEVns4tFvh/clZRd/lrUAZjHP/6YDlMQaSBufxSpiRjW5ST6uZPxZeN31vYL7v48JD/bu80wnw7
CN097DN1pHpGlMlcmHppt1EoKIG5uKz1CXPTnYAQX7VYwwxkxYWfTiP2NOM/8adUfpfClx8PAo69
zh/7ZTC3yF3aCoYwnVLLcwToJYWiTCCNI/Wqr6WokoYdem7NSHTtLZposeBd2HwyQVpT1aHiH+mo
F13saF9pb4tMKBaONy+jf1VkSq+nEVIcObzkdMtrrE6bCDCBikUwAJDIwiCBQYEMpyUwAgsNK1hV
TTpPp87Ln20gP8Uk8IT8IeEOKNENAgWn+0VYJQOqdl2YRXyW7mRKXT6NoRkyYZ5SyDnYtWv6nCSf
XJDwyKnGyY6eq4XL7IQdH7PCaR/3nf6AObVzWw8uXmRT2DdbKKAE6U0oO1o4o/G+lekwN9dnLdM6
2Wcx4zPD8AIgAmSbum3FgqGYVjTuNY2vM3VVFs4a02CyvlUQWVMTDkEiGR6K2JQNsKcQJLVBILt2
vmhe/HL+GEbDXcsY8Bjos3xJa977fkQCNoUUlCVh8Fx8/GgpOWld3X9AZcwzsxGQql9HFARGiXUK
eD3zAUgn2B/IC6atBuA87qYzFgeg5GDZgjkwNB9gPyTrlmxXFKwAcUw0IQOylh9xLHtIoJHfpJ7n
uvP48WAQDE7xQhlhZzBgvMiUNW8RPmLfVOUCZPvd5SXVuJJTPqT0e34YtObCLxCSkNkpTr+ZXocj
G2O632dT9wtN6EcvPe/Lb17mp7L8DeaqR1vSdaibtrZdAjQ07cCu+xBgFxkM/KD8B/1V6Z1KiIRc
Myo0DhCKh0PocPp/ZzMnTADOlYbRI/OLa4ZXHGss3c3MJvQOWWByJASHhBwsQN0Pq+DOXj9l4Jgn
YxC6ayZmpYZQKQlOr6TpLxxC8tz751rx2dFmrvHmAsaZpUGks7/PEvROYZJvFFpB2/OpgFzCNIMj
f354EUB+zN7gp+yt59SoeX9Hpy3O5aqrK0bZJqWgqRG8Agt3uZSRSlLpV08ASciyuSZyr9pSsIDI
0lxku9xzTx5A8570vKjp6SLs8vUo+/wyJh49ia34kYJkk+oy371Haka+uezUlz+dF2daECIevHK5
dxlpCXeC7+khU+mXWtPNkgPn0uzymRlz012oBIUy2LOX1jBgvb2ZezHrdvvOqSsOOqeo05s7721Z
r/pxxKG21zxGqA03kRq7mnl1Nxc1i4jm5TdAFHB5ykwm973UcAJajeI+/5CPuKLG0fAU63vO4J0V
PEcwGc+trI2hO0Rwq1pV2UAf2FtXrCcuy7qhRr8lJDYMhQycDvPNwfeccqL4SWout30HLrmp+Iv9
7Ampi2TFEUNhbYM6hbNv0Rjc0+Q+/cFhDDenQJklDc+VkHTv+tRqkEFYaYAJ63fs7Uth8tS3/RQC
9DLTtLxraTrX18Vu7L76cv1wZFtwvMNY0bPYAxJba+aPclUxt++idNJManI8o7izF12VwM4nUU0L
oXATMoa4BcouYiZ9cumWjMWB8nOoZWNjbAtfcmDLDQ/LkOs/eO2TktLLwY29HysqK7aubXmXkObX
ntHbgdPkYviUuYkIAYCRz7+tUCc7VSJ28hZwMtl9yQX+oNfybJ1x0mK1znWSciCXnTTXb2OVq9ao
qeIefTkNvvTxPLpJ+zZSRkK1qMBk90OMgM0QO4HKJ0tMZUZMNA/pn60Hce8RAM9uFfJ99JtCVeTf
oQAdIrMMWnUrlliOBgsotdhPFes6onXlEax8lKVOwglgsJ+ceHWry3xQWtJkbDpjpZHJ3/JlgdGF
hsxuvHHEdH02Kjjm4+wJtR8KiMj9n1k8nHSr6FaWM2g9uDtrJHfX4SmQppfoAdn0O+/+BqHIIwGg
+YAuW5Ehl4z/6Q1HtmuJZrgMhOTr5SW4RGOaR33I9sqfWSLhX6tct9CrtTiwbyPKhuZi1FGW2nNS
GrXhPwiU0XLkxGZShDJ9il9yjH8IzSi7/Y2cF1W1Qy4305rSepRJhd0xNrFd2xeJmWhwD4sk+noP
ZIh1J92PTfPRQdJ4WcUsc6V3BIyI69FzR6BpBJxX2lzfXdoLDzAgNBduQl0m88eIXkDsnYmE9SHA
V56Ry0Rdd6vd4bTHGTlAJJQwsrFINhAik/20OrX1DcqmYZkE9I45oSevyS/oyChpXva369zzW6JA
MZrGtx4aswfQ0ZGDONDo8Q7NfLEad6lshERbzBceKZ8Wja54SrO43wX8AzBI29DbqPQRQJfq6c+p
wACP3oMMXQQOcsHl/L69WzrhAyOMBQazNuXTNU5FGubuY1X6/y6qsvpQxYsyBDjcv1lTq+pbchhd
ZcLpOgY2ou03CXix38XfuiWZkcXk2An5WuaJmsK6z4iFfD6qeygUvUJArDd2RksShGfJv3ke7fkV
UJU6EHwy9xLt08KLT3ihOfyULckGhMiBu+6x8In/lfmZT1OvwzfwN9+j35oe29n9F+ZTKyerZgK2
ombaodCeID56ZjazZBptcL3gPbcXrJo3GS1fzOrfleWP52lnunRumqDQgEoVOhwEQgP6HUwxyYsI
C8Yg9pgeMEntwiVC9HAKethMjJs142Waxk2a1vsCyXyHRxec+IXexpNKCpLuxT1Btoewh5wJeyTH
eFcR2PwNprj9DFZzhizLl70k0fkweHYTmktnGyhQTKZu0hs/oUgL6Ux4M8fBvxJ4k0BrkE7bahQc
KuvZmApWtXrV2DpRId3v2Ek4pHcwroILQqxMNxo3nexl522f+lqDIxM9HqBQ9/4lpmzG8fnjRwLU
vnkcV8zVPY7T/UeYqu+oHvgk+3cOaLDpSVDcZoy26iinU/bc6/NOKlK6FE2cR5p8AHlaFCZLLSkj
77l8mH4U2ApSNl2veKUM3k0IeG7Bz8xfK8xqW0uYzHAgf6gAZ0pU/kq1uk+KtOJy6+gklxr7Ivf1
uPJy9a+Wm4N1OfkYKrhEKgyVWiNK+VUrpCBh72NHIvua858tw6sFoKAlCjFIxHCYN4eHv+wJu8VX
nN4WhIHsZ+JvY1IRIm5xSrgC6H9vBO1pMQHORxa0kcs1VtZzdzCAA/JWt0NFGPWU222qLfD3NyTh
HC6NALy2nWMJE35jxVW5Ok1QGEt5GQiFpA8NrZ68FNFa+nsPtQxCe2DaOv8+qGllFvFU4bl/8ltA
bHrzXjeAQ8pPz+aIMAZhpu83hWu8TqsJddhWaVvpx/nrX8bDYDdaN1mKZJHDIXGqzDWW4fS2TAHy
2BZNRKyS/u/FhPr/BFo+ke/U31RXVCZXkwnw59vSli1IVwGw9+H+lmiL4ibwLTOTK0cD4FM75jMm
Nbg5u57r1+1eSDG35B6z+5WzGq/EAJOKjs1r4/F5eIAGD70xkwwT1KKcphUiIXWAGslwSMZdZYhI
grL3ZbcLcT5GJwM6+jdZybkKrAP+KvXAkMPcKaw2qp3k1TZlWPRtEaFqkLow3zJcl3Xg051T7GHc
t4Fz3s9V45dkr15TN31uYS03J0LeYHcYVz2ynZVxYgkSEHMLNDCbG44g9z8EjJIhIWzfMx/Tk4OM
s5bnM+MI9gCLWfHCkCe6ofSPyWkKAeVGadSgx2Rw5nQGR217Prjgu+7dqTBan5mkm0h504GHQEd0
AVFTWW/3W6r3lHC76Io9UxnUqSB/DkWL1xBbQ5bjap6kt+EDeJLxSdI8OGKIQ2I0xkDIHYNgAAEz
JTOBca133wEZ/v0PKUbFDCWKwfKs+cGVsy70wWU/nHCAlWqN5/cVaxbyi0JA3VCv+yCJ1SNmY1nZ
ZuWEsb1c0CVlyER9NKm0G0DbMyJeRtERrmCF+MgBFwOBz8p+RINx/ZHijt9d8OnZh1uLxfJAA2ex
rTmA8DmqPxWxHCQfFI+OyRX7iRuA/pFe8/06WFmvVaIwbA/s3qAZ8sHtvVDc+bYCv9H+0/c4dJQS
14Y9ahmV0FZ0kbgOylZtjhuBgRzAftqj8rrVztQbkfkqNjQJyAYXe9MlHAKSpG3mLOLvg0FilLDD
C3+RGID7W5zYF6DSxOZBQ+2Fp0lMbkH7Yg+8UTyC2Ste3mhIaOQ5aW6sO8eZRnJYGFa8TPVUu5HS
KXku4mj4FAWwNX/Tppq5mZFMCGuWKNQLfUyTV+NCx9ZBYgPmJD+zqwyLKoxK4QypcNbtRQGMPkDJ
3VXI7EpeBmPYUOP9yoVD+QR2PirCbSz81Jpmc1ivlbhTj+B8nYCAvTh77ja+PnlHkFJKNTaundwU
zlG+7viVzH1KPl8BmWBTmLqQQV5/rNDaZu99nd0ktamHbQKE2yyhJO4EypeKG5KigT/f+exxM/wO
obHq2UhH2ZlroepxYpIwk3iLs6NTrFIlWM0g1V1UUYvBbffvozOMZeBCBM1FJxRjwkXB/ljT48b5
87S8yohOaHntAZL0CEVEC3j9xdpaqb1x36KPRKgjLEQK0Q2iMuAZdyA0EDMVCym+zrIppJAR0CHJ
r+iPovMSk5jl5t3/+PxdWJBpMWUJhgMluJYoJmdgoBBA9ZChrJThsLF2j20yeKlbTnJLg+nCwG6e
a+W/z4C+7gKwawRfqtzLYrQrMOBprTi+E4ny4nyXTDdqTMHUelhrNj8XfpeTwFrm2fCQs9NoPmH5
l5kWsPb6ALdgBTDD56ke9FgZ5Mlb0W3V1rZm2a4d6Zx1JTcqo1Dy0JBJ62QMc8ekBeX8Piub/45z
lKCcqmNlMr56RW9mLKlr/pbP6JdDd5WGg49oe42WvxBzra35aXivgHG+szWxarkbOOtEFmBJWnaK
1b6JNCVXuZZE3Ve51rnE6qlEr5GhLRw+V4OOCVkGWG+d1UKIOFEMu0pS9ITAA9cB3zDhMhY+hYWu
YmwbehP4DD80WmwK5yd3Vn/keac9zH7Mx5nV5CiAgvOaqdiONVFKr/m2B7K16YojgapyeY5aCJhG
lujyE0k1QIIrjPjaPQqXS5e4c/B5f3G9k3zt6JtL7ZsvdUMMvMTTMXSQ7jl3gK7UKuNiVV08zk1e
PZ4FdVVJk4pIx/5S37ESCFqDUe3abf/gyp+wW5SnJGjng4Gnkq77jqxgvzJJ2rXo/iZKNl+ly7GR
N9crguVcIWiPtzS9IHtz7OAn44ddCbtb6H8NkSBgMwHOs0NdRMCXT77YAZ6cqq0PB2jbAb+kiAtj
vnEED0wZr7NkXQcvswLocO/Xgz9/GEu/t2q4PrYCWGHpm9Hrc1nS6R5Jw1Vi0L5cTBl/iMyk7r+H
IbgLTYJ2bZfEzDpmBO7xWSHgbmP9+eMhdL3JHJn78SUBcNpbo/BzeNEgQRBjiOLEwDDb35U2aXeZ
9dn1aSJZRJEuU8zcOvVwwBH54AF/aisXWR7ka+iH2XfdO/QjzU3geUZk+a0SV/VqaghqKWRlS2Hm
ma3pPPwR5plDYh10V2ifFoexKy3I2VOTn8zlT6/kKDcdyu4m0884jCa/S6O3Tz/cWT4AdQE7SOuk
VGLq+IwZMT7Yq75kaZr1Ijy622Y2e7Hipyrld+teDl9e8gmSVtEiAh3EeoRS/oEOVV5LZxFD1Du9
V2AeM0iBd3/wv5KHZclp2sPTITYHhYNuRPJ6+jNbDmL/bzDWekHMETjAWk/RygPTX7yIuABAnFvU
VLKLye04RUKGxS0kOhX5sA79AaE5XmFi6cYG87amLXA9MAXmylYTMIi3gSulbdDdPWv4eIeGnZBU
mOleogxJ4QFcP/w0AGgR3L4TzSPKkrUwa8HG2nWYQAswyJniFyli4XWHAS9S7Fl8G1yTbaREfRiE
3rmmSlAlx4saON4k96cQdzIHhonYjiG3syIkOVTPyV3/tuEbq5YK8qAfrUaneDwdMEaG5TGYLjzx
OLksmxTAvmFqj1ZKHKeGiJNfI15h9J/bQw2oE4RvjYvC59InPQ5FFQ/N1g5PoFi+/xY/Q352GALe
1ImqB/B3vOhVBFQkUXQyYEXn0Y3L6E0hWiejhTot2rlJiVtSePEfE+R/yDOiWx/3qGXDhcJW/7Z0
fFe/CcZ7svTiWVlqydhaqGjz5Os5ch/gC9Z2UPuCmTaO03JDISXKZDTQ0+xiGBgVTtFXmWGVIRxO
F5SrLhH3B6Tbr6xrfJHvkbRJ3cIWTKXRhOQ+AWAu7G2V9AtGGJ343c3T2nziZSbyP0P5R3wPDJ7w
A1qX/COvgq+W0aXM+rTc8ttYN0dEN5q+ucdoSFOT8b8sEWW2vj4b5WXU+5jBoXlY8LB3yvIB1EZY
0nKTjnfX5C8oZ/4TRi/V/4DFERLJCpjoZlp8jv7MCeIDT+8i26bTdIEfPlygBcYDT9fx+NqKnnK/
zASUU7BYPrvbMhneKsmrz1zcDJKNPnplqW35G7nMpJmX7V/9YVwOI34gB4zInKd2eGvXEvwuX4qp
z2N/b6cRu7lsMy6rqUDYDpD+U1MuVrhdJWmDdl6Gcf6nrTVW/dKVbLDSFweUPab50fdTK+yEWwXK
gTc3nila98lEbFhjFY+igsyq/aXKMJN+4IpTyqpLPA2K36/bSIQ9n4CTCJvzpRyG0uaEYVy74eqc
m8JCXTr5EMgdGN8F2oqj2IrcLZS/EnWTjqiP1FOsYaPRQTKr/WS9Z8f+7WGT1/WfH9S13Vix93LL
Ug/29CBgxe1fj+p/CiKaHxMh8Xm1GWqMVsukE0LHW9zAfxwua+KiXGZZRL6u1MszvlMrxBcvZQVf
KBYSRb3n8VWoN0K42mQYpjc6F9sc94bVFb0cQOZt2BnxUbo+ZGtNtMmmGt2BjJm5YT/l63N3LCVU
sRAouPCkiiR7s92jNoRguaXs3CFPmqp2cxRhkXNrDjo2G6QwQO01l4Jk2zSlivot4lFExmPaFQtg
mjdKMrO4LHby67j0zIuRAklCjvVpKvPt3s5JtUSxgEPjw29K/hvZVsnkjPbeSS5AOdojJrK5+bnX
Im8lFt3kl2ogF4LaMFbP5fUOk1DtbRa+sO8Dcty17JBoCyBFXt5GdF7jevsU3aL8AzBqAcdtrglA
3mNBxT0V85PRiOXVseNCNCxvVj4yAuOG9NFCpbAevG+cjA4i6Vp5H6uhqWPBcsnZ8VPDJY5q8wCe
jphpPKMw3sPYAYEbGDz2LWypqDObEoC7RcpqhhR/D9WMSqFS+7tQkkOWGO9PY7FeR+cg5Rr8Xb84
IeSNiLaGw0rN2zKKakMMNCotXCRbPeCkqqiTrwbK0u27aIKldkBodteJyRiCkGTwoUV3FFnqdO/1
RP3W/jujY6WQnMvpPjy+Lwx2BiA9HNm5hfiHrnqQWPY3QDvJ3ahfTLEEyumGmiDYlewUtLzo7rRv
VbM7zD0lai1kbv+vpX7YLKmjt92Ovg+m0orem3I+bv+lRfdHTXVYw4IgsZyzCOm+INzhEMCqlFQN
938cNO4cMroXvxPNAjwTs02OPK14EawDV5Mf9VbU3w9dq2CnqUu55zR7FEem1dZ53wIpXkTyLQX1
mhvqKqem16M2qychuk4AH90PLhpTbZHHxP3RL6HIMXFlguB90RfCjongwRPV1iQG0zAsuzHlKATj
GQmU07EaA34tbUrt8zd+2YfFFZJqMM600J7w8N/52HekD3CYZ38WN5Y7BUFpirB5nUzJHq2Uu1Ca
FbLyoOWFPmbRGQSxihczf3dlon1LdwinoBGGXWvkLZBPMdgNO1TxMyJoIaPZ2Zz7F7jRRmMv9zzC
iflwoYXVUwa/bXnwWEdpjeSoJQsnqCP6OAB3ZEhCVtKifcDjKMicFTLWzWbF0T+PfW56ZKl+Ulc0
2usqQYWJFN4ql4yadxBFECLUKb4k+oqzFQB9c8KVVIeFZCUae84gfdmlhnCu+3aDDncJxTR5ujq6
Qgixp+Ci/N5U0q7QmbOR3d08kk414XiHVthVbMfRKhTBWNQQ8d0NURXbtwBgZ6zGhonaDCWScCOf
im5uHaaWg6d/ejv4dVP7/D9jAHk3mXCa5kdUegUNkM9xK6VtYbMGelDx2zezY783xQvSy43YrKJU
DII5Nyjg9rIA6i0hfgtQv3GtzwY+npF7N+3FKnX2BHq3DB71I1MwE7GmMFOMnLXIjbRgNN7cZPA6
O5MHJqC9yMOoGp+UjLqi84mQhDLiGmmI4G+I1Dh6hqcm8H2vSkQ/d4MjqsXUILfW5ymYKKOIfkhR
ra1dgpNRk79kYVxKfvUWMkeWRQyDZ6EGuJ35FqFC+uHOO+uySxAwxnGzkvGoi/GTtj7XFNu8WKYr
xlLAc6lnXeE0LAXnZ8FAjXW0RBFEs4U2Gm3JsQkZpqlY/LrwqTfykzOzYAsd0wRNJhdxHXIhr/ES
UKHIIepHG6p538Ti4Cs/3KFvCMoH0Vy2MqnbWMd9y8GKbdcP9i7h6zCvmoArLnu4+9q7G8nA6i6d
EfR/FDLevLRxBWv5amIRSCPPVZ+IZzfVeKXdCcakF2OucAx9lDf1y8rKhQkfMavgj8yjbbpSqUyE
yvn8d4EhhbQL6FeD1t51H2DDylTTeXfOy9cxue13xsGiuX4XWEbWXKTNP5xP6u9UQwOqrAKXrRbU
ONSUf/eNDG3eQFTKsl1ZCPs9uMqyx/c7hXfTggaWdzQh5j/9RMfdBDAU8kZsNCZrkLcoihbn9jNo
Oq2WIkzze/p/Gi52CSQA/UlSUxpiQsJoYDs1VyoVmNKPmSH+3fzLTQvjHyVkBfVuysWalYBgbjsL
x6aAetF3uXleTfH9Xo4ku7kOCLIQUwBBfpKnHUphw3J7oYGZ1LiLE0iptUmhy8vnTtDkTMfmvRdf
buPwFFZiddZwGA9xUOsscLCI/Pb4ocimT8Wd4S1tcuZAxlXXpAfJb3dME633C6v6mOKwWXBRJpF2
OV+PDh3kFfMkkkaxbY642fNAAfVtegj/tf93JkgZtQgzodQ4dTSQJdQBhKFtqRcjzuI2ZGx+cO0u
ImdrSdf7HpEOrWHX29o7yMQP6Dk1VOBPSgj0WhyPaVJUVZrz/rjfhyf/SaPxjRSDVdc+Htg0LiHi
KmFb+rORJKTy9x6TYPnwnkO4BqPKPt7VCPTx/EA2aCijhvU5OrwzB+g5sCKNA1JwMpbC0jdWK00M
SYLQGsvfTmzrr7CjQpEtGycgrW3d3qZH6bZr9ArwFFW+amrAB47EhRQtqgS2omEI5ubaFJwRVRav
DIFwRw87XKBKdMbkt1H1+Jt9qQ7WmmZGcJDppwINqCqIx76SQh0vbipzVFFLcuMA7ROtTIqOLPUM
Lil8Owt2mtA5wZlpWWvNTc1Nye4mt2G/3KwxHD8dYu9tTf48HnkHhJ4amMJWWnWSv8DY5DinrHzI
7LwdnZqPZ65Bs9Mpzmi12XemY9pw9w4LniAZb5o1KFQfUNuZoWo8zMJgszGlbj9UPZ13r4bniR+v
xSlyTb//8JDAZEQT90mjZmERAd5xOrECwDvfkUP7RMq6Vh2AB34GyMAZk3CLNfh6+qQrZOfqxY+i
X+BrJdXZSX5NFs6sHS+Z+KktR7W8hxQb7jmLM0yXT7RomilLgkrsSc7pTNsmx0EUwLh5AvUM8FiZ
x/fNO3op591F0b4cbaUYoWEEF8bMYJHR+WHMD7MJP60ve3coBvPs5/gWiile/bd2D3RHeeSJoSns
MmlC6xOQv39O8iS7XYi6TaOfAGRMfeAu/vruaJboGnVEYqHue74cCS7DAYiMgbR9CqWpfqlD5TE8
cJad8dQsZpGtxyxMsPxP6jk4lXHMor1dLDkN0lpvYC6CCqcNyGP1oQHhyvBQrcZ2PH92aSGECC3U
Qhq1nVmY0XOyLDqVbP55gksTSLEYZEJpf5aiBlCTqXPSGdLXn7VjGNrOLKQFdHqGnRsXVAkqEbSd
72/XF1xmmvI2ta/dcKBMI08RZsKW1BJuzCik6trrtskWK7oVEbhcLqRuCcbvxqkw7KTbtU1e+f4W
RXZWpf7gTuDvOhVPqnRPKJfjL4u1I75KPrjpVibWZsX4EML/QW/tQHkGtVkOa4BpBsWifdtUhtIp
gGvowY5euLt9XKgatfXIeI89Lul3fjnxvIdFaJhGxDNveDqbzpJSojIavnRnqbeCS5CAmt9Q0rSC
j60XTNxvyXIctCApwrx6kJ1TTm3FuMNwjOhBI8Bxqxb2F0wo3Wuc7MGSIGot9qwxM8AuPo7J9cG6
46DjjVy2wQd0QYHP2gJDvDdImVf9fJ/rtDpNplWlEygm4InDDb7K7be1HcAGpJt372guSCcsjWVJ
JrTGmsH3h554LYOBV7VRRVMPfA11s5YWeuabXMc1ZkkrNoLPKcFGj49GHCQdzNrHHDDTEHxzXTJ+
0XNr/oYgOGDAKh9c6D3l8OP2fsOdF0cE1VIak0Av0wMtSQBVyCQ57nVN3jLYiZ2ETmfEBHa6LcgT
kqcjP8m/adkdGjJvZh7Bu6ZtrnHjKiwCQHyl89oTh2ptgg4163iUnh8YVZSySKuMbdWTH1HhphBo
eCTOWxG8DNBaKuY5RVL429B/HxSCt+9gzi/HlwigJUYXBIgA3IdSm//fjELiBYwXDzL1l4UOPu9A
kwkg9foyohqsMk5f6aaMvoyYgkAJ9yWQxwbK/zzdLp3ZOtt/rK1jTPkZUzI9eYMGYcBt/x9Opz5q
vYVr6aW95nNrxdbVViiCe5Nk7YxRqsrOK53tT3FJ0iDmWGTTgiatA+a0Ol8fbg/xnI5I8SRLJVNx
1x9HTNIsTxMQGdhJyFq3jKApvZNK7xmFEZGFCXIHNv6ONGDp6IIV9Nw4ppkM7dQ3oDCGXqW+L3Fk
7QfdYYzOvY0X84p9q+69jYRP827nnnDbRZ1nuus10QawnEXe8muqTc5WdlyGuEA2kF5njcNso5Ru
+kNWiwUvAMsx9uMGrpJR23MNC0CgBv8DUiMgGC7YJm/dACWuatBQkGJtZ60gQ3s4va2p90DfNLFf
HMp0jpNs62nQIuq3RbGV1EQ9z08uDI755BLGWoihQC71i7Pbtkwn6i00LcoJ2/Chr7Gqpbyioeie
E/2kVsLDUcRccdp75Q15rC/8Y66X4qjiTQCFdYj14u0p6ghRIkNooXfQ0YyZtwK4OlEqhkXNpnBD
uoUhcLjsX+BYFvQFVyaUCzBtrSLUgsoVI5ShOH1/9gcuMH2UNMRJGB24UvXJUtIwvPduVTE7kfMV
Rr6fRjsQLhaflbAV0g45jDovd3EQczjxuEdrbPc8sJ/7lDui9nyqex3oRZSGCOUH+YfuX46OvsL/
k6Is9pMNrsWbaMZ0wwy0TrlRA5KYxO6W7+EF8tzHvdZaM+X52zedYO9B+eUlw3Fpnvj94LgnHEWT
0a7MVbqTXvs/u5dsIRT/N8RRDkM5+nieJxSxE4opVxDL9i3Vbt2sJyflGwsSu6RCxH9x3uLj+XZl
ZtoEBg5GPqmG36an2U4FNn5C4j/+sMNkCPa3Av/0FmC8hfzswOb+x8Ei8fha5BAi4AEFaF13Rsum
5EOrRLudSm3EmxP4X+K2pmMQdzMadgyjHtqiEGyrTah6Ur7kkZk4LYuDW9t8m+taUDnmVWMXIAxt
YNaOuy4M3gkJfCp6UYBCUF4BEt0I34qtfo2e+TXU8TGKWZDVTgjg7PG6hvZ2O71BSQ6Y0uiF1ysZ
ERguI2A9teNV/vTVTM4t1tLcnPFE3p9YJLWHB81lId0B06r/ipOwh/xnERsYyNSB2ytPJI6oaQhx
Lwlh8p5m8zdAtiWbxRosb/kMudVbk4lLN52UgbgFHQ+lixCLvxACKnKkzdOiRgixdyvwIUwd2wNh
3X5H5pH2d2hSbt0EotY5md+xnFUbP9s+cpDg4Jgnt5QwWSwZ7ac84nuVdwHuR3qkBIQkqJkRtMX5
5m5LYyFLoyfvMJ/KaZ6VKwc+sEg0SMuDpXHWI6FDesa+pSaBrA3y0/k/hexau5KvI6rgfvvZwfDE
lY6BMy989s9Riw1mCxHKrPsgaampNljVzsYiT+tO12ge9W9Q/RaXmty1i3e5vWeo6YuLgdMFkWlF
5gNLW00FbguAFV2iccm3BFUfABvBRzMQHazcBgJRftYvAFr8a77iVfxgcO33JSA10GahkF/aMhLU
dnG8+B32fHECNkmjkTzMUAbn/4w3kxwSkAH4UFCckEzZ7h5B2EpR8Pi+h0ZYwyVr0kSIj6OJ+soi
7KhYN1+QbAy5EEacG5tvTEtVJXLLT86byIy/gbYDE/NQtJz9uYcQpvA9YLM6TnyzJ25LmcO6hcJh
5hqkX4q4wuw6LRrfzSIW3JiSLQdXRQAk186DQ61CC/qCoi27aB3otlGm7Udrwo3XDCuT1fziRk0B
iNMZQCUcUaWNevhmmyZtFpM49RACATpG3GTgUSRLlyp3ylJ4w7eisUfWd+nLdd6Fc1mYHQ7z/cOO
H7E+GhUbRDGopP7yhUHEcIQF5pbLfsA0GQA43O8uyhwdFwDNGDTm6j96DuYjkmTfR6oVF+1xNgu7
1mdvXxy+9bFsTKon3rNN9XOuaY8gsbjAK81ldawuj3bysUJK3VNlv3ggCzQEZ+7KEcuhaxgsevj8
o+KAAVm2Q8nYrHQM6fabnqi/l4wOKGzkyDf5WlAX46VhBEeCoPJHZlnBo081BE4KmBhsw4kQ/Exv
oxpEemtI6DMDI87eWW5tZG0KnvpM/UTRYIv8RTsJPGe+/rxl1eLjVK/mo1MJi4ot1w67uZreQ9oZ
3O3avgDAGsjA4VVqiIFSfJ2v5Fa+p6grf7EvWTuJVclWOS8dLeCw8Kx6F9Vi/C6hZL1m7HcDFHfF
4xTx9FeOeKmuEUawomK/eR+wHHS2iKVCEe+Jm1t22x1OgAdNHj1PXhn7boehUapS7i7vo17rigdR
YkiLoi31Yi+ThTBNCKwVSsjwPfaTLbMb09GLn8KRAZR58ww+Fa6Cdgf22BwlXhlPZvNtB2Svlvs7
LqjdWe7QwB8Nyc5iRkVIZpdtFQqiUNDivdYAHMbigfpi7ittRQlFn45jt8GszM8lE9V6vpB+QSEF
K68ZaMLvWuMVgLZINTVv0Nl45AuyuMtUq7JjdlYuC9cR0a4vxOquwnUcbpwnwTDtG6oEzUJhJvNt
EvtFp/EeF1awiudBlsrmp/O+lFwJi/KJWJue+r+3rfjoYhZDqjOqUBrZtFGZL2eGVVJ5rBSeeDCz
v542YbAsmeTQLfcjunz7Yk0eJt6SdKwe2Xd6cksTjCNgZ2Fz3e7jYMh4HrNhe+DG3x3IAXPEkFwB
nYLiGb5gHhNvpJozXyWlCvk+7hnkP66OsBCDQyulH+VP0VezBtfNOlIjcSv3IKm8s/OQYz4MI5i5
Pzl46lXt0aCAnOgb1IwtQAOj0slWE5MnOT20JHmCaemzVEUZHprXf2vV9yEAEvtdB+UBmIJtWEMb
04+A3Ffxr0GNB/571OV81EGx606rM4fH/Nt8XAybAKVnBEIjAg24Umj8sYp5PlG3OVnUT/6Ssvw1
cZy8JhB1+4SJdgAbO5HqSBHXosmG2mnT6n4Tgisqjzcv5BGXSg3xPtCseaN870NU7ayGWyGYsG0G
jjdIW1uAcxE/6fOSKRecnkjBWAzfOaHzfjFiXa3eIilhMn+khIbqOdlUtvZ8y+1gGp7+0yXhtRxC
xuoWIjqD6aERwW2yHcWFZKI1G4Q5lgV/WZj1AZHUKV+q6vJrlM+tHlb1KFTW1zK+5n6hwi7RvkYx
udAuUxgbU+LP5SmO3qPVWFgzE3IUpwJZ41kAt7bhWP/eJivzz/eqt59iGtseRh6ZghOOI1yW1O0D
WqsIpxpD2AMkhT01VYqkSoqo4yu8eLheNAM2uq/lmGuqePpmm/AtMcq44cJgseE3qVcFBVulp6xp
lPevXEBebWJ+MdT5X3jcuPsnpe1pW7hat+DbvtTwt8yq3odx3W/KTwQMZwQUe3WE2R0XCcr1a80Z
GmnUyiHL1w+rZch4FdnIHqTzmLKtICfesHYvpkcMTpQ9QROHvi3J6m6l8dMra49CGeL9Okm3hR1l
cXht6GKLUBJSymT6MowjvTFu4tM1+BBMn/90RF00/NysWFM0mbdvoKCbrkWtCDAu6kpVnIv39R/G
f/+OpCZGJI2oG29zgbr91sW2uLxJYOp1ZVvYL0IIkyek25O4ZvZzmefAicYqx0iQ7Z4JMFk1VHgt
qWE9IgWQ6jglq9rK8fKF14aqCCXoBQW7x+Y7VLY8/47B2cXNtDPLavamrZsVXLsE6APTzkRNispH
1G8+RRJa+ujfm3vnDPA1C/WC98eoRZPDne2PrG4U9zNa3BtScgpINDagAGayrtw8p3Yii/Q5ev7Y
2dTWbOxgcykBVDlo/QA05cSEnx9O4yzi3VDXhivukw6qt2TTn80rPWwAg22Ttla6ND+OxGg2FYg4
YC3Ir+O1qj3JM48clNgHUkXC92pNKBfNQp7+T/uZvvFEMbpGjBmKAtgJZklLfDoS6PU3wEP/scbx
iAN6jzpm7Gw8wN8pZO51xgYMNKqzWOSMTRhieHrr1AHjhgH1vbSd/CcTn4nBkh7j/v2G/HOWeX9C
xy47U5gV3L3YHIkK1ghAQsbk13jRQL8RPrdG/01NrSQgwa0lfUVkxoNyV8E+yeyCTEY+DT2YAY6n
ilsWrBJJf435w1ong7zfmAkB30ROTGwxeFa9cOmW9Z07aJxcfDolQb9xFxb5/qkQZqdUwXces52N
YE6G7teSneEtzGcoacvrTCobkueNDZSXwj64Y81g0Diad9kDktbhmmxMSYYpxvE3CczZL0L7DDiQ
O1JNekffW/iRnprHbnJKHvduv9U+sFJl3sI6/nLajYTeEy71KtqNdFMoHdEqTviT4W5zPoonaIPz
axVA0ZxRgpAoIiQm5iQMJ/eQwtzkqzO/ajVmQB/PdnWWA78Y8T2FmIQh05IvckjwN6MjZm21qKFo
0iI6c/Bjm2NbXmxesU24gFHG4gEJn4vlYHIfPIWcndAEQqXGYsqJ7R1BadGkKb7frSzVQbJTsclU
vpZiIFJU0Elg7IQP+jzi7QqKg/ntp+DTr8zYKNDvwzHLgAR091C1WPZi+IwJe5/iQjkrg5Cev6a9
bvXnnl8ai3esHzOl00PS38pZJI461QAvYrDt0wyl5FOGBknEtQPjLgZDBS1XOjjoL/hi54kgTYG3
a7moZZjAL1OQte6MZTCP2U/czheWphWmpMXHYEW+ZSZYRp1/IQztQEQ1Cxlrbl6zFOVlzpthtMor
zKUWtyFN4CHStWoUOH7QwB8rcWbiwEHXaR/E3H6OE0p8O8YhlQi/kQ/wRfK0c0KAegjcMIhr0qeU
QQJZ9VEbXORH1hatasCQ6dCN914cazDdgDS1cTLMCxONCGi1beBVK61S54A68WFHbxa/gCZPqPYR
zqlSR7aGduCBHb1TbgaPEwNgnWbquYGXaih01l4zm+mhcHsuYnl/O7YGHKssg5RgkUWkCyghtxrP
xOCUw+Cl565hoGuzTqeCJQDtBGRZQE0U4BazDj9L/AQSqwM2Y7m1S+MZhlXzIcTbc/iWhVE9iocp
Zc8wUhe8TCuRL6267zCjAqBSigjqKiiZevUpwjmuWL/yoXKgbag293DTIg8Wwm/3MTef3RevOwZv
Pi1FIGk0C0HrRxx75pBdgjHQQIL8qYP+1kyqDi8jjiPrG5fJ8wjtEARiPYAE2dK1jQtH+EcbWRH8
H7bA3po63Cs8ONFD2YdBUDUoFy1Qp39pXP5bmr0u4Rs+kuH4sCh9Ld8Ac8chFZFY035Mz8BlTOTP
NYqBsMIYV1YAKzZTqX6oGVPS9Zpw6q+UssvcpbUraRNCGIg/8johUYNpyAdwIQc8lqPx6NzjjE/l
bTQ5XCfLztpX+kYj57uBJYOxGZAuLaJTvggOqKpcFNEe42ompGwWFF93Ekb2vrB/ciGtO/ouOwYQ
k7XqiIkw+Qwa1zG2OQQ+aU7f36BL8+F6sd87pwMg8N71AZ3INkfbSfCoTyAnWwfFEZf5c7BOpYnb
qzNsdBg45qGXJarOSFlWsBNNtS4vAWgenHgM9NZaZM6TZrdMqSKWBRDNNr40e219qTv14J0sDbAy
qu+bgdW7y4JMq0u/xroJIbB5JFSYUR2pcCWpys0HOQ6uDvdYLwjiGJ4nDTw4nmU7e6dI/LC8QJIK
tmfOifqi/0mUcfGj9mE5LLYOC9IHdSak60Dc2uNJmxSOaqAZHkE/rI4MpjuTeKSeVID5fcbG9pfx
Ehz4nYtNnox54TfbmNDSK9ohOCY2YYFYiJc7xABOkw9/IW+lmuOjrSUVU5O/S8FfOCYDm+Jh+9er
FEiSXreUTloaNkQKGhBtCxHbNR1XMrRG203iYBeVvCn4sn38D0Ur3z7JoQyA+dWY/waErLLAr1zk
0qIeAGtnCKRcVq1NR0gEDrWiq4Xm5tF+yR9FgAIvR2ymUbef4qFRoHPxLgE9CbvvHmy8XfeSraps
On1lhQ8ZiZdbx67inC1GutPQpQ8pj7Mppz3JFQz1P7WeuROeKrXa6qp7GtwXJabqXDUtA9RI7Saj
yKY/tx0XlTK8+u92MsVf3LCQcEbqWD4Dy+ftQ4UC3r6U43eBKa3IkTyXIq1UubPIOA9QFIvytsW7
VOSdTLvH2eFfJW1xK5dQPajpv6NFyOJdE/1RQN/+S8rHUo/wL7Yzh9wcn0vxuy6ICS7BQxympg7Y
Hx9vJaJUBBTDR06WJgchE6fy8IMXcZxFWindugkRgFC6vu2TdpnPvy7320dvl14BXlPgogSTDPIw
vfui+dWpy4lXIE9p2nlX54bELzPLrnfACsS4r/5bfjO01DezVDkSEc2YbE0fPWA2lrLMkVutel1O
mVNsvsU1cgAnbNHKWpnjQpRN8ZHHhoYNfCIiuXYZZWW0GPMC1eX4r1ocGY2ph+wodYxoDIOQJdAZ
LQxQbuxHLc5s90Plw2+gQ+Vo9q0OgvlFgQoXchGtDK7X698m4OTtrUpMrRtz/Xn1g+GxeKuP9HRv
Z2af/bGHQQu09mQ7vln9IvWTuL1vIinfJGLdUYOXDSBoGdpmYP3nRlWSxyK0FmOtlnOATihe66c2
EKbHa5oqXkOq+8xANmldFwVGxc0FQbSJAZXaDYWr3AZD5mtRO7v6M6ulFLIFYSb08iEWZ5EcTWTd
84D9G+j7QaolZZS/MP+ilh6fqnq3PlqIniGoi7TPAAE15r6IbsVLXQjY249vuTibZQP1AghnzUL9
b8atfDl47VUr1Nft4YYMgqj1TxAt/8kyIw1VP9jr+ck+4fZSYF0jStjsBrddSAG6pZs21qD4go0r
hMlm46TemH89GMhZ24bDU0TPvmo0DoM5Lql579ZmU+dNm67mGHNGV0sRmD+ptSIkCR3yO+MeplT/
Nb6mSXe75TBy4HW2NhfIwRhzUuzicqy7B/Rm3ECnaoh9BN3uZ5PCNV8mz9hLFgY8puJcCpy4lDd8
gO+q2A9ZX+3mTFc8R2HnVAxjF0tdY7ffRlNuu4/EcmyLU/LDDdrGLP8mGaHPHmDISKWKkeujS1Nk
SuNP49t5Fm2RBE/LROWgWU1ipSJEjy+kANvq8Ibcm7DDIEwJCxvsPYoYWMwjOp1F2YvKdwjD4ZyK
s1WqN+DB964H343aKxqBZydV4yPB6kxHntNitYrEXlkrsvhYdZZLN0I49InqrvPOKPFXDk7aqDCs
i4T07LKL6u6JRz3waeVLBgBkiLTHnCkhfe7FTO4taWbQc6LcOJg0IPnnVPNNnZzoCKCkAvK33gsP
MBKhtUoWYB0+gNOOSWGqxnpFPE9oN/xx9v4PmkOT5QsayA9Ita5B7TPNn6ks/jez3/KqapNQYj2S
31n1cmwQEuG8S00ZbSt0lMN6T+SqIEHtTbxmIE/QWAeL7jlapRVvXYXD5eygZofi5IH/5oNEJ8+p
+XlLXUGbrTBcVkjJK71AcRqmqeuRXGFg7OK5qL5zPOhxo+Lm1L086yF9iJsHog6XQ2apEFWzoeqk
VHziKaMWre2b/7bK6Xtbad0ejJiprMJZv32caftPS6bx4XS4yPGWS1yiqpwl8o6/NEDHIg1IYNqO
vhizZCdjxn4Oo0T32feRTXEDCeoGMFcZlDWyk+YwPK7sJw5Kof7MNaBVq6emuz199tTUJL2CgYpP
khTAQsg4TAEXWSkidyuJ0EccTGGHOd2s70hlVRPjp3N5R8+wlbuG2+m+rp/FQ5GBT64JuA/YWsnT
Qce9wUN2kUfW/4xneE7Azm8RNjvux/Gj/io0CJTRPFdKvaFhbjDNJR/J3dqCanlMjwTeSpt7jVeN
gVQJzoHr5CHkI2/4b+s4cr+EdaP4oe3uOLKHAZX00aCwjxEr4Q4PIvgi6Yy3sumP+3uWa/L9VFSc
b7+9cQwfSEH2zyP96Hr+8eYRPf8JVNeef+RqKOIB4iKrSlxCfOxcjNv9e6GLSQKZzSmA/Ow2Z3om
NVWBMQ3QBi0wVSWjkcCMdreAKMicYGmYxs5m+KTcpfrtHf7PanA/WeBI21v5+i3tIuzKMk55jGPz
aGM8Gvn+o7/TTtjnzqoAWqf6kwSIHK+rNFczQHIYnNRq9It5hCNwToRnJ+B6As6bJa21eUvIoOfr
JIb9s8OZciXlPAHE8z8+9KiqEDWkHADia/YDtkK5hrEYJUo1bluFtK3Q4ATh9BEGayaQnbO+H9ta
zJ+k4vVqVG1o4Jy05z/R/sHWm2PEpJD3QCfhBP5v+vB3diGmakEtRLXkIsz+Dtpjl41dEq9s1CKT
pHLTyC00+IM53nWAHXyoRxmsCQHGRuPWVDnqDyTgVawu4Oi6xuXKqZCOEMtwY8flS84Teay6r1OW
ZQGAqp+cf53pw9Ek0pihYYcwlNi6+OPULmjyJNoiaJ76ahOkUBKWyAIUOvQClILlF+ffopgtSSoW
QtYLLX6gUNS9O7hJY+CYoTjuKO+y2+A26HgGl5AXiRMaV8enoSPNN4Yh9+Nj9tss3wR3tQCUBgLf
PDqhdEdqQEogwdktyNfhshRcerNCxV1KpvzSQgeiBrrYRXQy21Ui9SV8tnYtf+/m9DEpk4Gs8ZlU
BIh/Ibl9Ve+QRb2cSfhvXo+hVrtNuvq1rXNhKK422mP0Nnt8q7Kz+D7iXZpq5jm7vX/NS86rlrh/
WxO2j0zJSNU3tc13BsrjJIcAt8lhWciKleKt0DD8OTOo4l1yd+hRyDw3k6WouRlKkmJS1oRPzp/P
yty6RZqTdZyTA1i7KGDxyO/RHf8ht7FSwKKGf8LMVCS3UNeenM+10Bog2RteGFdKdcg0J0yQ72n4
1Ea/pGnOhQf/mzYkpRgmSUxmblKuELJB0TSj/kkpjPBClEmqMoh5J6iCxVsXIZlqq5KS2gRbiLu7
l+WEQWwfX401DRF8NhhJy+tss6jOolpGgpvwT4TL5Sq7ZfIoOTL2X0vwhGlqoDPOog74hxvVDxrM
E89mpD5TX1vOZzN4XYJFiIdlLC0yJPlXRR6cMXyhKl8eWbWu2ICD9U4ZgLLZaugLkL40p+1OxS4V
opgaJ3GP5i5olqaOTz2NwAdztW7NzV+ciFSnu3jrTaBcSN+fztNmnZ00BYQxSvmKdFNlNl38GzeB
zEh4tCRoKRA71OFlbTkA8LvQJq3WK7aSbC64SUEQGZafTuyY9ZXV9A/eVXBcdnJ9SSmnbTTxqjZM
Uke8v8Q51lt/bF9SuyJDSiabsOkawakYi1agzXstmSHxRHMkz4eXQR14MP8nG2YHDBExWqht84v1
uUaLoJFdVSmF8cYigV2Tz1cbMcFAQPm693xmmyXbTIRLPAea0uqRL1Vb1jRXSB/1LKW1EDFWgwVE
kCW1x6VpsoI/iZuXUoCMO5vwlr3ZHVhQZ+HOUqHDaJ2d3+8ziZu130oHACQoehVVG/c8pYMJUrX4
6zT1LPfirYOnRh+3pfsKq6M3WLxKjaWLpRjLv80jPumKX+TzPIscbzJE6BOKVL1WyY9UqgpsC0MZ
NZSCfGhlYkvsWDV0GW3oRQ5y9KHMZVyeg6QDdkEBFtCOa14kHcChS1gz38aCsN/iu4yydaqw/P9b
g0605kEH9JjNcqNg+h5/lMUtaH8P0/w1R6je1HN9R8gUUBiy04FXMqJo11PbJ8lqHSe9eturBefu
2lj0z3y6Tc0W0IuG/laUuWDBBiIbx8SrsNVsUzL6J678fd3BXAz5MJuWBP33/YciMRKpwikXeJHi
i0Jal5WlBXsGMLodOxsj+Pczf/O0F111m5uxbFvHjyZLRsp6F7PA7QZg3nnfWFUelFq5kJD0L6Ny
1cAcIQM1B1c19HaI+FeKI1Q5kCW8sslorRWZpvveF3WB+vHaxMIBW6+HCUk/IJ9ljVipUO8YeIlJ
d1g8A3/hOdpN954BarbD5NNue/ixFlRGX8eBoDotQt+YZU978tXpV4doAhVVtM6/EpWxCCJVcUGJ
NkVz402w7GpBPDN4M48I3aZmoBgQrM/GVlFE8WagEpyF8ifUNlYq2a7QPUXebd89Hmyum4gC8h6f
NRmpAzTIzIPM9zsBbIv0B+GJpExUVUIZJ6FjeYoSCg4nDEZojHHNDtW98YKwQeZmnUEiHqldkil5
6V4+8SgUCyp928khdEwntWTLh8CpkLpNEPr59/PmpriHkjDqJ4RYd2mx0eZTB78NpbAC22v4ekVP
3vDXEqCKNG+7SsbJ20BzCPhCx0A9QByID5GCG3HEbFwoqZN8FY6ROb4RGtJcgE3Er0QcZrv0jnpm
y5gMsJfcSNZvOe7/5Go69Os6orONB4UHtZw3RfYK1sGM45KUR/1/KhQR6vz+6Izyk4h3L1s3/PLD
c98DXzoEXZwBQ65NpllJe0MrRbmibGBz9MzymA/tNqs20h9wieP3RfSo3xG5RpYqXv+3od3CQLW0
cqTqs4N7Sxl5q5wIVTeQhXByB9VI0vKf6A3eYIRtUDUmgEDs88bYYz7CKbMHscjsPu6Fl4TBekmE
shir+ivpuPuHDgvBEGntDuN97Mo27BLH5JkuSQJmwin8HuR41Z1w6os1YTYwlhytg/dzu+TAgAkg
uoT0ERrjC4RmmR+ygBDNt6kiagB4ovszX5jW2RVLLXQjN3zMfl4zp8Py58toEqXNW7I/9Sj4c+nh
r2SNTZWiySJcWn5FCdjOhuuv2sgfX4261WPDeO5lllnQmfwOXw5le+PGfHqo7H4LlkS7zc0PzDaq
5dPrOF5cUTHznzyFwOFGpZq3hd2uaW68gt0z+Xk/9caxK87Ahxu4V8MF2nTSWObE8JjZq6f1DS4u
Z9gBkiDyyMVc91gjL7iZlfLS2a0tQrFScmt9CLXCqcnWf+K/pWncTGlDuHngXS/GT7NthSV5RJMP
hx1PlzdSknU+cP7NZnEomH6BsT7vABeedbzoY6Z13RHPHiQ64fJFo3cEwG2uXZdXsNFopUF+Hoxj
rGAJzt8jtiDndXvDIRSKabi3cQs5ku0oa6+IEVWC5ad8c4rnov+QP3+gs1RphJUl2zDMS9qAQxNW
WlIBgAcIbNJO3zoZEoMwMZSYaFL/ZGO7DyZqMbQD9OBtFeZCOAjxTZ750WTg7l6mUh0n1vKfUCoB
gyyiFmPwaI1hNIcQxjsEqw3AyyhhgAkUzHtRGafDhQnOOERFrlyH0totTzommiQa0k/ge/3JRHJ7
PwYgvHYQCwt7ZQMGo0NmmJSkXwJwZVNkjz9jUSZyfAq/bKOjBX9X7pgFJIAbWridMJKWXN/Y2cN4
lA/rFnJNM+7vYwLz+J9yC07VhQsnpczpQz1apdfTw8rGf4Jt2fj+RQXUshQan0rTjcnDd0JzuIkz
Uyp8qDtGIc27s9Gv0TuB9vIQkmuLIc4tlOSnLupaeJaqL45oqKzOUMnZRXNyqL1VP7s37HpdE04H
PKptme8apLXThFkW9Ne0MiHvb38rQ28FWCnduXlKf7RLzPbrq9Y8XevlCmKPbmr5Wrxo/ZHZvwJf
2qwMWUrYBDmNzsK7B8dB+SYmmIRIpAGCJfSFa1CfuPA1GOKr8RnSIiV0yMYvJKZDvdF54u/rQ2Ul
TL2VNdAnHAEEap6SYHUXdPjMHeN+K6J5uY1UQBP+JtfhQBLXY1TE+/4VlOBjdMK1gmTqNzMxSZLi
/HwBSGeyRlMont+B6+n3cgmYOhw62HD56AvpwFVWoudjfMaHxFa9ONLhRQFi5AXTRLoLYfaKa9EQ
8O5STbmHpO3E76M/0j8yMcrAOxGU5uDd4WmTewlFHWhtw5sRDDg0ynd7hloLsMZqFLuoY6jtyhNW
OTj4FpkY9DDvgCQjL26lnMd6sUpeq2Y8jhtFtMz5KNWuWx5CY5cUWHEJLF/2mAvhhy9aL4u7USoM
bGE2R4lsjRQtKqOkfDdlHoaie7cqcJV5W2qODJDP/oYgaT9TaBhALBx4kKFMJDH9OfAsvLk5M86n
oqZ/29tLOWo/qYMQUPrE2nI1HvoXEDQGka6XwcDLJcHot4iMLyDsFAg8AxFKIzHwePDnGUoKxcku
asAemd5wMn5qq0NP0btqog4n0YJuPQG9Z5vlPCIYuuWKwOSg42Fn5CL02gPHtw7qW6T+Rdao9bmL
nxNrayfuovIjMr9PbR1aSF0uk/I4MvrD4SxFl3JcvcGw2iaUgmHuPRZe/R9uwRPlmMjjbCw4zzHo
LaWHg7h+w3FS4eGl86af04LKsy0IEUehvunjxT023CdiqP7Zi2pmPjU/fFE/uMgiJM6lLMEwVnn/
SnIZO9XpfVpUZ9Ix3h2vsGwy3ksfjg+SzSMYHMY9IjG34/SeRaMfnbNW3xRgFq6qOL9rGSDkLsAG
crXbhcl/Ansfds0QhoFT4WLayXmHZQNGQ9Q2ObEqotRSYjBBoczFuCSsSZsvaednpl4aGXo6Qcm+
4Mmw/Losqrnzy9sKB4WGLOWVQ2V9jROlOhAeje9AZsWdsWn6z+sJKXokZ4EQG7kgtc2JnOs8lo7h
/ifyL+0NZmt4rSDicylFW9gJkWEj0ECoo6MNlvT3YlMFAiaiEu2VQu1xorQPQ47tVq4DgOhjw1eW
16LtdD3P++Ikx+nQTD1hadrtsq6BG+3jXseeQHu7W5abM89fTPLDdrIjBioIWhNGmN126FZ/daSK
ZWHF9lNOmHaTdBq4OoOUjtl/2xFj39156q6QUAxFdcsgIPhbK9xAQxINCSr7ROVz/qmvraQDIL44
tyJ3JW+Ij0ryBpY0WbuGuaCoQhBrw7S/irZFS/IhuoS97Yio9c7+DpsdH/LkGNnUzAypc+UKdjT8
wOi4aRSLwxeZQdch2vEq32ThdTB61QFiIbX8XY5+HvvoEduOAjdW1d8SY4cC2r/atSoyrXRQVbR0
YtDzW6CZl7PqfWjt3XFT5NWkC1UPYRUgq42VT94b6sbz/uQb/fln9p21e1/1RDw3s7/huD+5T4X6
DApW2DbKkW1Q5U+EpxCSXqEzkB1gZPGcC4agtbTxnO+Y3mH3bnPdGcZb7gVOEA8eG8dsKeYX2vOU
zVevlwItl3A6KrMWepsAwGB/yAQTjUdN6Xuj8KYBT+i3SSJLMIVD93WnvyP1RqGLkZT+L2blHhPz
fPutP5OmNQj6OekyohUc5kNokdXflH8gpNYKzN3yC9T8hjWQPrH2yk1n/aXvxKhf/FS8pIiFyf9t
cDC9yC12Dd+wEMwaaa103+W0vfw6uEaYNIG6Z8KBd+LKklcymq86NxokWZXsQHwJ8XLkh2GX3SSE
SsRGTE4ynTiYDl/sz2/uUyXQphOkrg+x69Bj3VyDN8ST7akEdv/LHoPszUcqsyjCPZ7BReoEdYQp
61MSXGdC3ZCGl6LACELc0Ve8TvgkBcuanBa6undeTUViugrBhSHJKsZiYqEaOoX2Yu2GRzFs9Za/
1KfF+cpo4cbZjxMrue+FjQUyaZDd2DuqUCxJQ4uCKxn40xyZ/iGa1slEJ55dH4WfpMV2Lrcff+ir
FM0LjpXgCZ4Z2NmfRfEt/HFCsoPTWcVIvNbit7a8sNUzmcxH4P2WHThI8NevTnSoHmiTaknhAb85
jYk7ZUxjkoaae5P70r3jNXXyOunGHlO9imJ0Qr+yb15SWShTFV2kRmtlusuEbLJREzRuhxEwSmft
iDNmYXQ22Kds1XtQdpASPEEeUt2avV8lqt4LPAY7aXKDvXlVqQdsr9X0RJos3CesxlRH9ZOZGEQQ
ZGTPSUms6/x6JnPk6QwOdSx6ovyQt5Pq63+pVcGpdBORhxGauLBtfP1L1QQxeNAzmnJDFl9V7cg8
/bT4XtlqT9ENcuWlb2/Y/s57ZXM8Rgu0ymPBD/M84GYyraEobklSebAbySXFB/zvn0U2AEEh2aCV
KVPvGhtQvlD1GCZOLnT4y1W8mV2GEs2YlPIUTTKf4m4SeiCYuT/ql361GNF51chCTbErmUzn2a9c
no4vBYIKgZi+TijOKhDQ+HmwLYJSZZ/9H7oiBfJTYt3qMsnxo8xklLvjK8FbvLWZSWA94kV1NOWj
3gYWmw6jOMWAAVTcRwFj430dUIkaoxXVH+CbDh6Lg3bRlli0L/30GJ6hciWAr4+lKzMe1+mEzEWF
WaDHEUfRkoFeJwa7+/gQoAoWobR22YwKs1jQllkmmF9vkYJIB8zWB+dUe3zZDje4ZSJhgoDfIKrX
9VSe30EnH80L9HCkenB0HUIUWtflwMLgC5ukR6591D2NpfNkuWPtkxmg6WL1Lb+xcrI/wFXBO/bT
zRMQe7sk4I1X7Oq1ZYL46kTYFiKZOZwUymECkEpwsdc1osw7rjp7erSIVVZ+Y1IYZf5DwP1pzU+N
to9qhze0QTm5V6YQl+W7uJv865jd76MJm8CwRupEtxpxdibAdnfbi/9xxsUqkWkaxqM4IGcUyc3/
6/HdprVPp/MHBLK8qT5BklV0CjdzgewrqcxuG8xhBr2A6eW4SxPPa2YskYZPCKiG1PdUKSX8xkuj
igSL7BUdUAILXuSECTPjck97HIC/W9ZL4018QdgPyAF60IaZ/zDP/4dK50Nbw+laGDSu7//RKiwt
CSmZ3eoozPb7NNeW37+IBI81yQDsxjKVLIz65dU3YBPEp2XxCTTwlcbsCWmy9uT5/TDqTV1fM2tv
ygPx+EGzpd5qdHfDQ1h0mb6lhSQ6BGdaLKsws9NMbrrDNr+5x8OxInvyiGcDf+nMKg0Pgb78EzZx
fdSiSASuDqMaTGRFgDNdq1YEODYOmodM/e0JNp5MTk9hOzsaFGvhIpBBUx2Q9V6P9L3pO0crO9FP
Aid5VL1dh8LhitjfdkZa+/JPIgoEnX5tb/PaoasBvVxv66QKk8RO30PfKO72iHltNXwPd0PvrOhv
cM0Nc+R5mRgVAw8JaZn1VQJReJ9k9jkQyzwWIx3egf0WBpp6WxTxcx+eAyc2AT9gRp0h8dQ6rJ+I
xzktbJ3zQUKu2D3AHPTpNYQb8SE8cRGzDR9q7I/+qtxIbW8pF1IwNy39j3x/gOgZ3t6EZ+/gvcWP
X9D9xgcv6poLSe7dNGKJ811JosuCD6bwunHmPHYB8aKVWcyBqX1jXqdEgZk1s/DYTQh2cIww3DU9
jExVsuXYBomrVnJlHDOsBn+pPBFPlpZGN/lpKlHoDODpe7OznGCSB6NuhRP2H5ONm/Tjz+68JBT2
awcYkzX9ZIhB/FdWMfqP+yLPdLFsaP7LVxYw2fLIv8aSsdpAp6a7CTwLCq/s7+hH/J+NT9OM8js7
1QCCb2Z6y2/i7685tnR0TH1u6G7tHf7xUcpzir9VbgU+3TtkHXEnPts+XW8Iw7Y6HIzC0p48xJUm
2T65YyhnvwtXBbZ5e3IxENyQYGZXVQwe6dGrnyQkTf7eRuFynMmBaBV6jO9hvDMMICNyPnzzp2Bn
MHOYqdiRi8DCTr6TUk76OuBXhfOzt+z2Fi5ZiCfdhT7gR3LfQtH2CDCwZHhSnywfMbsN+tBdK8MX
0hsHQVOckflFaAklhig4fyJxdK5xO9eU4obaQgCwjX+3zXk2Q7oaJutp+333rBDEaXj7v3EnJeID
xPGk6Ci5sOvoFACVMnc9X+imDhp3k/5FDfPN6V7p8zNMXxUWS1rprmGGSqEDtl8V9jUpUIdOqYXB
UiPaHAQ5H1ACSfIzt680qBiK6DWbeCETWuFucXaa1o4MvtLuiv8j+m1P+B+6tgIubl8nLNbx73mn
x8A7cVN7e41GzBnpSKVVOe/lxXS2W1MxZnVvQXummk+b7punT/W3EIXi13bPqzTK1M7hOmIWxG2u
QlIpO1od8RaWyw7fW5WlIyekq/InVPQUwMcDxT1XdkoRH5K7cl1xLa9K1jIeINdu0O/qrXkRsBAY
0agxjLayDFdYqM/ni7zNI3NvbPJWSMe3gg+V4qs6gyTnznlnf74f+12Zl+qVKNM3yZ88h6uQcp2k
jQH2bVTfpUZI7NkP30cyCxOAQQo9+TR+6kFDvie53BjNhQfQ/l3l2QF9tN/ZuSXuREDMz51BC162
BTc3mN1DkwG9UYbVJf88aDuOfTNiWgOjdaXLiy5CGj9K1V12Em5urP0uMMqbJ9y9dnrNAd3sh7+G
1ZpZy38q+tnqbQ2wGRRwbc7j9+YFyRpISND0ID+uHy3RgvvLTholvvSRbZTILwtiZe/gjSP1LMg1
2mcqLlxgJ+KjtsiSq39mGfYRL5A4LQNH/+Gj4Of4naqjkXn2A81nI2I/XQXS1c+oyQwT8ZUInHvi
3JnvHDq8PT0JHU/zl1zafRAAcwHZSJTNfct/swOfBPbT2HWXlaDW2T2SF7iv02JS1XtrPRxa1TVv
HvsQ1pJdBr4Bl6DxHejxwMU4LURAOaXkXs6ICPsGsiUs6lJD2ol5tg4Ed3nWgS7uf9+bLMNEV/n2
WDgo3ZQlrlcG3VWbnlLGN0kId/mI1T9VOjfC/e3WqdVSgtfDMvrDHNWxiS++MtL8k9jdbk84jgn1
NWDdDb3+n82SGfPk7EJuagcySGHu+5W5U937e/MJFaX0esr1cFQkOQUFtj3fXBPOiCsORGmg9iIH
OV9umztfS2qXJbtz7TBG5IB9l2R0o1IxtfX4MIDfFFr6lJL4rWVvvqfN1l8UsECtBBo6K1UsM68X
Ph0HVSvWAFS0pQjC++ogPyq2PqtPi5XpAK7G7VdVlnO2gFsk3EIA0ndhTcKoYOD8DZPSFtZMKNN5
K2fnK+OsDKkm+9x5fUfytAQvohMt9qUoDbAy7vuLWK93+mTec+WmkdPUrAKlXzN3BONChqi14aJ+
ME9bw1RYECx+OM2W1JScNRtx/Vurw5kTonvIYqB3P1/wUFOojWQIvut7E3+yPeGAdSV7b0GQq+jU
9p5Z8ZfxmC9mH5M6RdEpc9p9xu20BwKQyA7uU+f2sVqllD4Fy2ZBCJ2zfXT76Z2kLsGZW04FNUN7
Ig13SR2kmyCnynQJ00l0GhNrfS2gtmZtGslGm6BX7SS+k9cPpkc3msfD6/XQcrmXos9yx06halKo
ga+uzQjE/paQ5OgPNRRlSMsIRxtK34p0i0kvidqH2qk0JVTgMPPXdF+QlbY4AOWFQaxWoyv4KKR4
ML02XE53LjAEG9DpC8GD8Q9XptVu+idWnUFUSarQNk0bSHRveEWEwyIknbOfXpCe70lKaBWMjUt7
n+IUIK0c9ZJmWpNHHCDQYISjSIUeZbX1D0HvXcYY4mFJvlJPcUGKwMSFQv2aYtLT4THdKXRAr908
XngjSvo9dymVkYIRnsnLA6V98YeddBY9CQvCFJX994Yzry6MMtU6G2uUWUkZh8QI5E1gM06Txqg+
uGCqDyrCKIhD+zUOVxW0trO6vPDUn/eKCTbgRqlFqB1Q0esTKBOYFgLA4h+NDl4SD3edJ2kD51ip
lP6OZcZFsAdh+df7LH4tKZcIrdv4OJh407RVSKxLVa4Gp7GbgiZdUxrDAKl9Yuns9D22SWe0jHPT
JAB1+UWm4zXb9t3f8gaWxE4BLV3j4L1xhbFYwIxjQAIY17SQ5SUMuzf48LrPSSGoWcimuIzy1LoM
LpChS2T/WSEG9YZsbjBtaqYb3JtsB04aBUH6uIoz5yU/4tXCkGJ9epmsgRE6EdyTC8JpT3nZDSfR
wgZWB0DI1vgE7kdOX2mvEO0+WFEjWDMwFkD7snURBryHPdyOxDFe/9Si0jNorQK1PI+DeHG0TOFD
+AP1QMcGoBOWnxGkP7m0VaOo6cjfKduwxmBFHKImXTu0MeJCqzd/sFKi+dAyZIUMjx6ziPBtdPkJ
wGGhltCwvNgTxPrfDU8MF24ZuJDJ8Pj5nSqpSnh18eXRduKSwiVk/E9vJHC9o/6QcqBS+VFi0q6O
Tzp9PfZiYANlThtyKfMETLsCp7ggfkhPWykWo6Vq4bwbuMrsN9OupmZqnAug1jThZEjUtHiAswZa
hZEIG8b1JaqiUlo1grVrqoRqHl6d52UDxyBWx2MWV00brCIF1Y4hcOJ13dlr8CXnD3VB2pjnA1Uv
NUaMovyOq2NS92+K/BApUqY85eIYJrH+pXqFton+CIQsFzU0GlTwb8C4rSo7I64Evf9a5SsNFKZv
jvt/skMgXffbM62xfdVLxMBgpZu5809RIaDpIO9VmgPzSUj72IENKYQPuJb5rBTbuY0Zz0ZE26UA
0lHGZu8SnpiW4k65nzWjly0rGn7wE8v9RJw1hAENRRUfRGnav5cgGEwWzGsPu3C8d7dBJnF2KMfF
kxfVs5e/DcBFBUt76WM6iX0umI28Bb6M3BTLMMz8DI/rUs41U6bNnFIQFsVBPj0JQvoE02GPxx0Z
47BsZB1F4QlgXKHzLw6TVBT956HXy2bJe0jYA1PYa1j5ExqC3mEyPeTI7AZkmZ/naREpNJTyTOa+
nCP6q4imJBLipPglQRanw3m/b86XYhDYj5wgRk1SM6uhFsNilQLO0o7Mf30epFLoRsj3mxyVcvBl
qp5vu/krycJqQ5yXpRivRwsH5V1HcKBivBgA9g2jLIqNjTwdAi7L5krdfIEIevcFif9X9lR3a5f1
daX/7BGZfLVjYX1451WHseiMBniW3O8onxirDFEBqCVwGJmKMTGeZJdomoLcsQEwXGdesz43ufzE
oNGEOzj9ak4UdfnXvYeaHzysEM8rOGWr+l/yW1LOFUGa6qg/7DgMpVjYQVXGCMsWz+3EHqxYP5eb
knQqmsC8d0PjH9owE4yFSTxA9GDefNAnvOXqLJYCb9GvdAKIa5p44bnAu+/DCMp+pPo6Vx2CtAtK
KpX08SR49wR/ylz1imcdndncqlshZwHniSiC13NTsch5MpcyIyfolhffT+b6QrCYLiZTa0LGa2WH
X0smesM+T7YX3uXbq9ylf5wN/D3jsXerSgUZ5oQqc+I7mLvFv1/UJh4jl3pFQj2RLhR7DJob1nJL
DF/qDSDwXe4Va2SBJvUn3PlU0f2QqoluTcPO7qBL3B6umM/JKXA5u+eXir4BfRTudREpaSiLZUbn
8Or6iGJgHsCHaUTza0fYACUcwpWNE/+UZJ1Pmh4PkW2rjvQR3Y6shw0Zz11sA963B1YOz26kXRJb
Ag7lmxxVRfJ7+zzsG69dK++YzwWjH7gK8VzvYUOBxHjoOiUkyr8Ea+98qxTGnvIFEvhKb8adc6pI
PQ4QQmi5qassglgvQBSI/A2mM9D8jTktz0LulZtQNaYlufk6AKuuZNtOR/IHVNwOOYHCbX+eftMd
LWClv2c32ElXRaNOLQ8Oic9fAnRLNCOG/3Kr+Mv03cxDdNRr1lP9a7j40OvUTFlJ/3V+pcX01i4k
INPgeR4lH72ViZetJd3x7C0OuoitwOGd3Pxhae9HMRKXfHSSSjYRWVItEo0Ez3C+pGbCwabyt1Zs
SztG9+k+DiRGwbAdw1grHn1gQe9e3hOM1LYEZOZGbeRiLB4L4AKLWyAOzWBVKwY4SqIBbUMsVIHa
WHKK8DUQldjQwk0lRQSg+2DnJRQXIt5wPkvSfxc21X+L1JvW+NOrs0V1OynKzRA8YerL51z1ajXA
R1sRqtSb20Y7G3XcPjpAGtNRhQk00UkS3GJm2Fcntt3Yi7lejOU9tXZ8QjQpkawZujEkVudSF2DC
WvqXQ4Hb1kitvEc7NMz6iSk3zmHLu8nWW18AT4m6Hxc5ttkUw079MPb1OMTEKKMs1XLH5F+ZA6de
e3zM9iY1mV9FmArpuIp4y3pgSGC4t9AuVf/L1xKMod2eqZjg8AID3+dU11LDERQnZjwGLHLWa3lP
Rc45O4DjgMTcHJFxyG3mkZG1xJSE+Wynh9vdkng9KUzfgnGtmQBXfgSzC6a2m5oDgh7cqMx92fpg
U7ueje1im/l1nVZCtcJYJzd1mKxZmRzkVa4w8UN5ybMEMrFRjt0yDb79rO9m++wsn4VpxueQJ0gb
czrvtC8tJguE7/vcleWb+ak03pnHaaqZTtpK/1W6AJdWYfCvGRHhmuRoDfmvhL8w4UNjzMWq3OLa
Moz+ud2xAV/qeGChsy6yREoJvFLjx3inEggv0sFowTUiz2O+gLEa1sdeZn3SdQ3q2IxIXucBo5zI
vtq8d94FIppr8XdVZmCipG9oTXFVtuE/GJ3Mbpuulfr8O0FzscTKZvE26yFXCkH+pOCOfLRbuurr
D0Gd9ommqmcSto89hx+PLsD82cjgRfh3jeEvmzSG+zVaA+tYOne5kXDVk75weYnny65ApJ9n5FbQ
IdkIJpH3njk1iY1rKda9HjTKyvSWB7ZvmTYE9Yb1qzKG2DMqegRGOpNlYvG0Io77p/W9eo9rPTZ7
LSsMi4o6Ml/t50NOJK7t0J/pnNjABU8bcN++xOoriC2OCWEuCHZCZWKO2R8bqdw4usdfD9hR8LFf
DxOtKo68MAfMiVPKitfNbvMGi+k3gNkYjT8Pv1WO1XPnqZVy/hBsLvQaz1OkvwPGSXhSnHGmrHFl
CrbfC3StRbvOD+F740WFthK2UCDYvDFLM8Cv90DiK+OhH+kf3SBY5F1G2Ut3TH+hEWuyTwIu4Fg0
KZAR5DYJvYxv/40JnDUeZ9u6uRk2fmq6HGIXl3h5lB3PjQVKZPmA5ZRKoQC0/NoYRdfQh57zw9a5
/O99LCuX5WBb23n+WaPTDVHE07nFsZB4fCnBBCGBinHJPZL6LuQAfSh7rcZuwv5gC5LMQFL0W2sF
/KT7uOxIeESjbofi8h+kca4jI2gjTkB5JTPGXKZYsltIWfEPWjBDp9dihxhD5NHuNoGDfE79gcbO
oZOhKcB32kH+HoBweHOiYONOCEbpIu69E3RhA8zIZdhkGzs5F4yVm0NVyRn0N3zvKq3EPds0Zel8
GfY9zrOpAF+QaHxJDOdVz2SjNu4CvFquoWdw735xIhNfInR4sSgCDb5QX/flG4O4Zvwt1x5jDuvT
5tfDBw6cz45zYWI7shq4vjiYrGpP9NiJ+NO3NPWaM/NNOdPW76sxsCqE7eIypUjNYXK78jCSVOxm
xTXTBfRLGCm0dfldPw+ZJMTT16jANvtS7wz/5LrEfqkTQtk9tvfUX0eUBgInMD2hMdcC6ln9VY9Z
0EjSZ8HjGSZKSFURKPqFR1TJT5LtL/dbpwZ0bIfWzLBhSeaFp36jX/GT8St/9ytOFOQhtc42mk8v
+lAaQTYpqo3rY3MNvF8fsEiTS0H8NfV9ida5FdHqYUoIMayqXOBIrHxdmf9K1jiMRQUmxwwFdn0S
BZPuEZeUXiSFMaNenOjtF1LBppnukdm+JhjhjYlYMY94DlifKTsPoKvrP1bEginre507Ki0SErgy
80GTqApt0Gzi29yOZ0q/kk38saZeSOC86cdunsDKP5Gd/aWXkEsr0kV8ftCkvEjdSRFNLhD8EJsu
+VAc/I0T/2PMj0hMkySNjQ+FR2rnSfoOolJwGlmecmKy7LFo8QkhIkasYsOEe/LOegJkNtFJFFQN
xDbpY6ddXCW/EFLrNBUToOLwRdfeI3CQDkjbIvFr4A3r2AhwDYS2uOFnf4OAkNXj4f8GbvKJSzse
wCHgxVdMOjdrcUDzyCJZay2gMuUahko11cvu5Es7VFtzrvp990HY25UPxqCElLdAs+1KRtx6nrFA
7QnyahgJXSGRnwUq8Pw2dsB0NlqZf+THrOlbgYTi1AAvlRf7WNrW77GN3oGWyT7deMWRD2hvwBBe
H/pBmia/RlicOXHMGaYLTon1Rc2CSpLrpw+H9d62CP5dS9IQ33xx6Vp41icSVAyUBMuVKE3nm5VL
WG1kr2Sa0loHMeskhDYa4boQvTKQ01mbHXeBgdfg9BE5bUPA70wofB5HxPYmma6kxzKqnb5ldIfO
ZftrodfRNBDofMQWKybIp7xfMpkig7eo3Xhw41iX1ymLEG3jAiBGcLTkrxKvO+DHqFVBq2rksGid
V0YW2glVUxeZFI4j1KgtDONQNn6fMVDQTtdVdGOKt4KrAIo2FDZkZs5h9JsBPGHYFtmIy/nmHC5I
BsRU6+exZ7rgfHVJVLsSY39kW2auSFSWb8LCQQhXp/pdT9rnM/vYNp0L8Qaj+zeK/Pi9Mz7ZVSBK
A7s/hW12bnuDfwyTZPQb1e3MkpxbBbPEwFJTUYNlJkhA2YBlQ/VYtqDmeFeeMJyy/NIZ6+X6bzjT
6TKALp1UQOirdekQbRFX7Y9fKAfTEf93qgAlBXERW+2n64mOKaqYbs39kK3EJMMt7RTochT5UymU
3u4Yw1R4Y1MFLh6NRiyr2QQ4FqHxvVnIzAK6oDStNYRCkHD0w6HIB5tQoKAzS+GPFocrhRgznedo
6iajUtw/ipOCSope6A9MWiXFW+dLYC1onlpuxFb1O4mwAG6iFLLKGqxkNTsyvxpyXqoCC1mcQFm5
RDlGigISmRFPT2eAeE5QsStLDG9tQ12xXMBBS6zfYsntByD8HRNBMisw0gXwvyB3kmIYbBbWH6iT
GV1NTsEV6XomRw5Pdf7NmKVv609kMp6ghZ/D/rzpsP3HCszDqzX15H1eC8W1tPk9/E/o5ArPxJAX
s2DeduZBqU/+n+Xa7nqhSpup3HwRySFemxjpzvj9AxzuaQYuRUFKTmndUEqApPO9Sf6GClOqH8uI
+BFwhsKllphKl/Hco9pW+d3bdCD1VPB2DaH5SgmxstSDI6Qcfmc7VHnugRd3caQw0wBNH4bHgy7S
+364+EDnzJ1teo1JJLRjB0GrGaCS0Au+3nQO1WroHLy6wWCQphpCsRqBc313honB9sMVTdllTmAn
CE6hpOYaXiquU8R/hHPYPvqlKGgIYmjFz/0elfi9l25styiXowAuJO1BMI7rnDlytQi6P3znKi2o
MUYZsHH+AZsNC98vIg4VmYuTc/kyHRxFGGs8F4/7ov4470/tEyHM+u5MBJmYOb87O50b0c0JSc2Y
EVbZdFBO4m+X+9I+P2AfjXdR+iLJOeogeqEhQTeFeQkHHFyuYMEJ6a5eTjvFMauJRUhgC6p5Jdy9
YRoDfBatV423by9eXM4Oc96Y6bhu2MrXoAwvXZ7nWvwEQCX6//F53yIOKqBJnXuYwb+i5aCA65Zf
yw+C3zMhA8JHpQpgDlS1EGu56bly/MRVaSKVEWlmdOuVIMvg14U8r0NYIXfbhp2pZibYN8ZBZowc
2h/XBpobtD17ZWN57l12M01wn+k4/qqlaVxLwsDhgdfsvGc2tO7obnigcM1VSucEWo8gVo2Q3HV5
iiiD+c45mLgMPLeIz0LNyuvqoTVe0qNxJfcP/pswIIfH2PqkdgUxOXqqeh1OZtMda6l29rI5FJ2V
JLpQ74zeXwHMSfAt51vax0DozD2//QwO8u0TadfoHg2rnEyg1k9kvU+D1cN3wI2mUwIsNcLyqF0I
UU+apy0h/5H5qR1k/ntxkyaH2V4baJrlYtA3kAUlG4y25pTNNLGTF9qZMZv01d2DVvnwZvX3uivV
YYgUvmGZ+hdDv+TPU05o/TqiUYCDar0y3Yf1hD1cUny+VbdiA0rLiSCq1ictmDBmFC/e2FGrZddx
3db3glNW3I+9A5DaLHBElUZvabAgH585YdyNKp0+CEKK5Jlm7o7grUIazjdBuUB8piWqE647Lbm7
KGKN3rrD+Yyp1s6yUUURZdc9D1IZ2n3I2vQunf6PQzFbc6oFLtesPj6ilbw9z7BIA/CwWN+iiVLu
Y9LOMyVEyInVhAn5O5CQ+Jpe3cHDJxi//8kllkOZ/e9BsuXJnOzqHbay+YesP2oU0B3Cr/xOIsmD
EqZ/GbYSvYRmjVIevAbz26cqKPWWrKh6p0//4p1huihIP4z0Mx4I79V6WJn5XJr274PoqiYI/WMp
inXlUWJcPuA+PtelI1bcRvGTTlCp9J4H0uj7wXNekcvzJoQwR8BXIAosoTUbjDMIZLZMLbIiiuGo
dAZ3ly19At9VbhrIRbC6qqhc/BehaHVH6Ke4F8qJrN3wRWAa3PNLopNM/3CVJXFg4Q7gshnA7/bt
zLzKsmtEn1AuIOMwZkRYt6YiYRafUWSNKYmm9RJN3kAy9l+Shn9KDdbYebOtsB41KIrsNMXb4xSo
K1Gr0bBeXVV3t3bMYQX8ucNiE6p7twDYoUxNWAg1l67tEt4LY+jnBgf3Ptv384rX1iqWW6yHEvpZ
ejnGmq7AuvEMLFcql/CO4SbyWwQfln2Sl4u7YajRCdP4sWuT8U21zwaU4CF8hDIOXpb69HhmC+Zp
G8GErQbGRN+IF3fYdvO2RdaFRbA1Jkvc14X8vsHYuLjozImHOcE1UHt2VJ3eMgbXuq+52I+J5mwb
+fmfS5EZwPAv3l8JLlD40y6CHf3pdgTUOX07UWF5CVALI/h5M58LlPpMLhaoPDvvJ7wag0qY2Chx
aZzbUDStqvv/2MiGyXPCDKstFpgaTbIUGMFXROPc2uV9XF/ZYOovjnOhNNrObKIw3zZox1jlJyp+
6OxXHJZeTvh7E1y3S0BUTWPvwfEaonWgSPu28IuPOF7nfc7gTuxK4XcC0xgGMV+D6jSYHi4dzddj
WFzs/sgZUlig/mWy6d+ALZXmQg+CQ6hpipal5HiKZX6MMTcfMw7BLxBi901mPZKLU+u6hTY/ymCc
5pT2TzSmgcJLoovRDwMD0myuQ12TMI0VljgfAnreik3zaEdpBPkp1vX1etYwoyYbky5Mg/gSokad
0OGPhXyK0SxF19GjgeyNIg50zPP7qSyNdXKohrQUVARBXAxOB+I03SZBTtahGv7B3qc2yh4pN/0+
VsPqNQ6dOqo4uNXSUDJZwUFCWxSipxA65qSbXHOODNZlthr/ZrIRljzCt4g/4E19L2OIfKXa5N3R
4+gP1aHhIgOamt93rcCtEcAqDUm8zULj/js2qtTYdSi2zdSX8f0v4Kfcg/AZEJg3EGU82Vz+RO9c
X5cumv5nLYJHMwHMYe36982LYts4HvLtPh00kgWIMg8fNvXwJ7qFqxOv61kDyqLjNaSbf2oHs0zW
2l5R5P+goWEAAHGvMIjxT23Kei8dKLDLCe/Y0KszVov1i+v4BxckNxMlHuSmn9HMeG8JPwy8topt
KvAXlyHNqcqy6wbXEXVFVc4VF0Gy9kpCoBAAcasQxSCfJYkodedcJGZNc6uYylmocsDjna4X2hf4
c+sDZaaF5uYx9EY7EjEkWC6e0j+pFUBEpMwHFXe9xxA5dDA3ghEEGrjdD1vcA/0KuD1ZX3hz5V00
J87Ox8dvPjTlxUHGJM8tVMuuGwurQDC4WZP3QUz50vrmoDIlbElp8n/lfPlyBQTQjgqJnvMAE+g3
4yqp2s2N6jwVBVCS13EODfVB66jfkUTv1VNDDX4xfh90UlMik1Ce55jpf7BKDS+3uwQUYIwA9FoW
txzrW0haSoIE63bhyYD6ooMYpRuqLTOGwOBYkUhD9GtKZ0mWybr+qD/9EZLYITa6vee+lyx6sgHs
E580p15iKvm/i+DU3KpRH+8SspdyyNM19GChCn1u7s+jJpg4lEikY8LDQTjxKQGGh3JNwKg6uWxE
ykyYeGROToXQFsWuS2yNUC+CafPYPbH2xkMJ9NJkBzWc1dwtmfLiH7bsLSDKIuzZD8Af07ly4jVe
o/jFXlDW+JdP77XAuXhgxPVYfXFkc9GnLho/+CmJpPy6+R3d+fLVwSHMEbfuJX8GJ2i1kFl7a3JS
+nds66sRHe4hxXMpV28EA+11ZSDxDA0CqTqEwRSWDGt3MFZorfIlZqKTnXSP90360x5lGjYYqLD5
XPbQipyQnsFcU1dWoJDHRw9HpZBiv4Risqqv36PACvC/BypV6BHiTLJSb9YMTFJ0oYzgBqwslUE+
7V515vxKsyFCfW7Yd/JfkqDtXGCzLpRm2JcjBQI1icIqHwpktO9oCnexS+bCbIc7EiDHB0KVnRVJ
UD+ZNOP4WuPfpa4Yp2JKSYMBhMllUrxucuq+2mN3pcpzYgoE8aK5phfLDN+dgUDYIgvdfPt1SsQ0
YjHPegqw1G2n0vWLCJxgorhmHNeXf7ERdIlmU5EC2w4bUb89p3kuiEWJqJvFiTklIdVNkzhF4TEL
+eERK+WdR3O8wBaMzsfiKeglV3z6Dr2HshHZAEyyJ9QGg7DIBrkEvmmQH/3AGXKKoGzoT09ql8Oj
NxSHriTGfvpHuwVaanK7LGmVV6HE5rcuKTBZqyMHMxfXBFAKv4qBCosouHRlbgEGZhXFdDxufXHn
gN9ERR3Cnh/aDaDtrjdnCZ7Xm5C8WHcNI9o9bs8VtQ9tKp8ymQ6VvmkN4kcqSeOBIRuhdB8qbGag
JIS44HYRX9doM8N4vGK+YeioCcSnkHkBi8c0WvfR4oq0NQUPEwxYh9YgiMglyBmIs52FD1K+PT09
ov8LOg5hSzTZnmZZHM6BXBGaO3J7opnYW3iVxjBM6R4iTTS4Bt3+VlgUmd1XNeLZrfv8LUrbbqou
4kuJCwQ9WFPpjMVuJ/YvZJ/Q+kNgWTCUZ0aw9eu2QKKPHYwwSKSmU1mtI2jlNE1+Ugm7AtiQd/zP
3JozRVZV6408YbtpucFBqhvR6Zwtek/vHXGMETpoWqEtZii8JBvxhbNLZnRaBQEEzRZysZRv4WP7
sdVQabC/ABuYMnbBCGqq0isX/EemBfLiCTF1jRp0Z5JpeJBD5xjEMnqshcyDO/yka5hSVJ7w9LiD
AEPbfZdnPRZqB227ns+vVcA1UeXuFxrTlA8upNu+THVLQPf1tQpEKOP3PLHv17QVmSNlJryluaWD
XiE7awMr8uK/WH2iiZF9dtZLixoJGT2NOL5bH+GDd/FUCt0V0Irrw1QVBhvryH7y6lyfcNTOAFMQ
TQveUiaXtRs5nRaS253sxiCkjPJ+7tWoTL4deCZa04vK986GJoDdqLrwGOtZqeK4dZjJs2Dc28BL
U3b8NeONpaF6pkt6LDJ5Uv5nYTVDpa9eFWOA4E4xTg3jOAiAYh5nRrVUQX79rLxF+9Ul1Qll72M7
tUco4kSzbsEyrTDb2KV+v11R0JC5fx4m4+dPy6pMS5cUYsVzgBi2LBobEgZk8VAfLJxePXDMekd5
e6xgNPElxTWhkY2VUSqh3QoVd24eoJbH5JAL7WCGnHjZ+4OuVvrFYOd9z72y2YfZQx+EL7PsEE0P
pco6iWJRKIcmgaPYSY2AHzPxsB1fZ2BPCxZSpkE6RemU2tHF3GGAZClFVLOt6LV0dKrg6QdNgGPy
pP0kvY30wD6nTESBubtKRcdDZe8xLDBM4wdPGcRbP/E27Vhu5nF8/uBOl0ReoyreN6BR73HfY/jD
cPfQD4g+qw/uTyRGn1128dA25LmgSXCE5b3PG90Dbj/gNSeC7kCQGkL7gOtEFVNO+QMx3pK2LIuc
h2p8woGsZ0t2DLhVtWvmJDWJhErsmdnG1MClbq1Q/yDFufQ+OQssOTT/LtYmghzirPPJeUgeEkbz
gWPGhvbSKsTdmz/SmNgl88tRW4Rf2Vlmm7MwU5HJbFO2e5AN6FS5w9Jstqzi/fb2vuXiAA5njL+S
w6lW5rC3+l7PODNUQOdP7+/DIlEASjPQOkgGJgC6llJ1sMKp3TtLcmPkp55E5hOESaDx78fjKiES
cUv4pjhPHiTgtmO5uWMqjwUcMTvDhlGKMk5o+xBkISL7aegpSEN0GyrAkyGuhRsQ2FPOUHQHdSKw
VeQ7pt1Nd8xxwikahtm2aYRIPXbEVeknExBkuK58ahP0D+xMC8fIzyPW6vfukOrRogw2QaOIFUmB
s4Dy8yh4o0Yr+qYIC3t01W2GV4Dfvmv/PDt4gEmEm1dfapqAyM+uVrPspQB2xSCorFwI+thIA74a
nEt7xxiQNML2t5CbhBYVAxFOwTQlnl2V37MIlpqFkx6AjBWh4IHUoTS7wxYnUsxtIHbX2Ny68kXJ
RFYCFqhALBmgrPbUIiuyygfkPkF83NYQXevYFHEXYMph0Qb1Re9pWJ3oOowAlyZtjaRGQy0L8At5
cmJeYvm0s1Dr4OdUMRSYVzaaMFoRlEj+YH5P4VMh15SR8BIiOvmlqZ1puzmhTBkTJ2pdiu2detAY
wLHUtrt6CmJ1e3EPPWfiflsdR6IjLZz9tbxrDeRSs3fyTkiyolnWjK1ellUqY+JOzMP3ZNJcmnoZ
jqcvn9QNTYteZHirlBDtSCr4fCG07HfFNScBtHVYgmJDVDyKM7U1i/qVV7yT2+DO2e1ioYsa99lH
HCsJ4Rr0w3T8x+e8p65OvSe9gmrAio3k2aSv5I6fFWIl21C+NuhgZWxrMoV5UOtJSeK9QPkPbB7L
/oUsv6r7NU/SSpXBdaRVeSRzlIsNm6rR0qbRWa8wCcsFoFvIKpDzCWT2/wHcyuVLiG73hAKAnMSY
LuzfPFeynF9vTx76AI798z+DcoAV17EEUO0UrR3goZ6CjKbAZ4aPA77E8retRq+JUYphaSsLQa3F
cuwpFxOymVIkFHxaBtIiDq67TINnwEEdSGFlufOODlVxksO4phuMr42DMaNeFPKXxdFJRCeyHIwV
QDNLQw/mFA2+28z+pM30jefj/Mab9MHb0rKDPE9ixe/Y4N99kVeYZGeN0AvPElnQVf6U58gp2DCL
0u1OuMZVkre/WneAW+Qn6O7X41wefW7DmozLwDXTvRg441tFOJr0aqdhUPMV9Gki4h6DWG/CYDpS
RkZg5P7MyXRU+W+sWXzmS7K85GDouCSYaWQVsqDm1nUu0fYt6pyFUG9sXt9pof97MBJrOB7mVeiH
TMkRR2RnXMrF8R/sgnNb5DEoaJ8gAJVaodiSN4QsD8Jw27wQSGVETe2q3aUPTKygxxzDW9A7baKc
j3PsXnNYlU/rvQPnqOGfB6t1ijGR9I4WibgwzjRP8DVwKDOsiogZFyAvHCSWKlX77lqJ12Gcu/qi
TJgp5oQJhhqn+JJHaa9WYLPXIHpiD7/gs/QY0tmNbSo8w0fAGptuMKPFMIqergqxzIzl6jBaARSn
A55QdbdnKEjyPHaLyS78bLfMRZXKosni+uBm9ldqagtfAIn+jJtU1TdvpxnZxtj78T7rr/KNdf0z
LGJTKdrsSdrTC93lnB4Bvl9NbeU6LTY4CQgBDv/73yGjl7C7O2JaZyoSPs5JMFnIJiD+A7Gi7vLd
iZWTraTyWWwmcEzO4bhKr23hlDQmBfo1x8+Nys3OGu/QMbYrYMEjOK9CknwW9i1fFYpd0+/ge0iZ
vlpuMYva2U7h17GYiZE15E4amJIZWoDrcEM2yMF9r17VM54ok4/tdj81pQbG0n7ZrSz8ZySk+mNO
SRgIP9qZOpQb83Dod4ACYQESznTYfsCG7t16DEqckAhjvOTsttVoJNmlxd3XUPcPUg5CJL3qPwtM
0k9WwQ3zLeW++08UgEt1zV5kSXsVrY8VDYhZawV6m5543lCSn4f3OAGMdZD4HOMOXgwmmfJTAzSW
ZQLsgkoXmfneJcMFfCEe9C5G8Xk1UfVe0viwYOa5xQfPUcA2F43FAgUwWWcfSisVmAffHHBW6pXH
mWOr+l7ctn09lFk7D58Axd7wYYAfXjcYMZdCHw0IpFWygsRpjkxTj44KQ7MurhPskMEqk7INDsDI
TnSN4Ip/f8HE2j13FAYvm2awNRSEi8B4ZtahVNcpVbBhHf8u5A/L7hyDc7NzSs449qyh+YuWaWkT
NZkFxBjP59hyPFnEMS6wNZ/CoVAxzKYJPOMlLIqkW6x/lOaP6BjhKp2n1D3KOLRStgpacMw+Vtd1
FMyt6JK1r6k7U0hbuO7+MPmbJlz3NarTYVhHhscO4eZupvGXSycu7YI3GTMNpQ1LAwI0YBGgdbzs
0FaNNvbQGScpAs5dXxNyMjEBVhNm9POoUGhodaYVFqhk6c2Vj9oZ50OC1kw1jP1Fgupem3fWrW/8
Rdb0UAF0C9NQ/NxyVevMfwok0Am3lpjnAyCFKebQW3+JTciCA8Bdefp+OLn0ekkuu09T0rA9HAlM
sKzEwZ7l9xApwzr+Ofht5t5mn49EL687hTY44/rxuSZYq0daafo0h/q/0J7Vt/FoIKZI/EbJ4fpi
Z0azmENOjA+fBWiX0iRsTE7/Y2wJ38sYcEqFAAhFp6EMNXteU5OaRn9JZ/POMiwanrd0d1jj2L0H
/0rjYzCSJfAnisL1S4XYfGyr3Hk1xfolTzxu7eFN1h7+fXUNumQM/KMSsfVJmvmXBHqsQkFEnNwP
6KoN5/TJu7/2aKOVRgnG+nGc8n30w7x2HHmAY6WtnwukRate9IFITt6MdRtFR9LDGmpb83WUkJvr
51m7avRlHs4HoO8akxs4bEfOz9ilFjSJ/AvrcdbBEq2FK7DxAG9FdGvrdUU70eohm7TQh0bqzekt
MOLfOAjjQ6NdWLikodcuFPI1OEirYvEC3tS6czYkrkyC7my9z+D4tgSDWLOd1m6l24XArUeVjjUH
bZngDp5E7KO9Z13giMhp++xfLEJYuGOgME0sUInxBcCnV9oKtxwSRw7vXez2LApiFKq/UbxSJPdf
MW+m9r5o4ta5fIDivd0lBpLX9HGyJozI7KCqQQEij4I1bh71S7DuRY+QGurGZ41AEEbCPeYxZbmU
aHtHLHZrqJ45nqvfIiHCGNGU+fgRnfP+t7yQj9qECBe5uMz1kNQLCLGwqx0CpYmVnt333uM0D1EJ
gZzM8BxrKlrygAaHnD6ZBKLTslXt0S4tYYQwk4blJaINeNzieDl6rKj6CvMW56XcaxVPIM8/VKrC
nORhYaTqq3jrxgSz1HQdoHv8EW6CpnB2WZQppDX3By3YXTA9saX643N/HtpFs6cxbPrMaeDXsh7T
7CpqUqOblrnMWZ2Zs/HcJGuhoCekQouFVF3qZNL81/XOxGC1rzWhgzpAqHOO1PROWFN2W4jg6v1X
lRSkH3OJKVpj4MZFtlJRsehdbDurqdnKaQILfqoQ9fwN78dqbGHyw5mW4n7z+KNtt7ayK/UZzWRY
2Qg7tuFMZH/36VIhfR6U0whNFzVFPUa4G+8grYAmKqeXcjnu0Nkj79T7Rx13EB7oNUXmHGL2r19W
586c1vD13TBISs1Byeaoh9/5lNJX4UAP8t49ROTdBU0RBT10TK3Bj6JnaCgtr3nh09qLnrojFo28
dHI1JWMbfy9QPes87g2DN6pz8AUzdtYeapVXWpYa2F3+XHz9iS4e1gmtoCVNQYxRLQcAqzpWTo3v
lTCIbjCz1XShBSDb87z8Uelnp8hbwak/xrJChswO1jN8Rsk1qY83PhnUUb57Scj82UekpYKg1GOK
gcO2Jn96dRnOYl5a2Vlm9czt0ShBDyQU5e9WwA95fGSKKCK7+u5gR9vV2s1bNHZDzU5sJQKxKHEr
ZDnczg+YKWcFyS6P0doUY7WbV52QaoiPU4h/d1ISiao3u+13JOjYSduGj43OcZeIXWuuWiiat16r
Mw0TebWm4DuXhlOm/6WGXHe9HOok5/lKlbUwutghTF3D913DIBIdrJGqu8ui0VdW4QMZRsaFuLRM
IiMpK3VZfYgUnMc8xbfydcq7gGUt2vW1oVpoxY0cUoONmEdJ6LU4sFPvk7ljv0D2AKigxg033ZZW
nA6R4sBb5LBQRhppF4iPL0SxKi4gBq86e75tZQeRuJrOTnVrno31ZhP4qoBKLfjtMdSDHRKPmMqi
Zymw4Yg0yu7LatjpcHPsbe72m5I48xOjSzmFcnVJzgXH/7vMfTtwuv+LASS54R5uO5kAtJ6F8xBU
GRLyQfFz2vTdMkwj8Dk/Tuo2ZCIwzOZ+ZHCA9cyexIlozzXbEc7vhYeTo8IsXmefNlWlB/TeV3eg
sZFOPSM8P+Tzb5pltiCLhnWQVaoBq/wBGqD6GYLlIKmp0eL17aRcBr+T+xVVY7VxRSwqgS/NC/cl
MhmZl3hkM6hJHZ5uWH68OtD0q3j20Bsyc4TeQiDSIz3daw8HJcwEnEb64b3+YN9OLH/7fDp+Pilj
C1d/+jfjH9OGpKudKL/1E83Jt5uedrmCxShUd0G6D7Oq0xZGdzaBGZqw0DiMQn2CmxidbSuWB+fI
waPe/neEW3z98gLGeTfpG+TjDgpNKW9ds8aFkeWJd2m0gG7rpXS4D90xN1p1/QCn+n3O7QoOtTbr
oPeQfhJCACwo54NZ1ji0s9rQ540isaaxiOFlabXma4TE/3onXPNqGb8JnJt9/ADxu55rRUUNXkML
Twhyh9hLaQwMHOahZpKJrry6ADn0trwHHKgiJ6IfwJ4nUn5j4BKaRImUh5pQJpTEF/cNRuAxT9Bu
3j8Y/Agqag4zWkxqknPyKuzHN6CugLUwmStEJKDzU+5sqvCIvfzcimMzIusCFAUCtwktr5CFLKwr
nbyHS4n2oLw2ziyCyD7olJu6r4bORrGulRiNjXYV64n69ai89Z5e6JuL4lncWqvs931Qo89bfTIH
wkSNMmsqQWo6/r77EI/rw63AGbJHR+SsiB+akHBekvZEXJWWfpa69LNjmHDoK2RhM/nxKEDUtnSx
B2j17QyrKHcyDYq+TClzRocplWWHx6jnRNHqtz6QMi12ZKkfA4Kv+UUpoTeQ5BRNJ+TTjOvn+9pH
7ktXiVAQdIWfSIoE2gJNo62QgLtzvDIYEn7M4NyXuyJ4o9mOPSZyi7REIF9YV+jDub+VlQE9GpzD
cbYbZyKTbCHn00+iDld/ryaqapgsvrXGFumUhhQoa+Yda84JwhG2Z3zuE2Bps/qkQPkTq++Xxi0r
ctx6i0dnrOxeBWbSEykx5xDaAb0xO0MKBSRgx0uzVomP3wHZgxsJOsrt9KbxE3A/fyeY1kBZXxFN
C2kz2nogS1SmLFld7koE3n0jb/piXuFi9ia0SPc4rhlRJhyvWIDcI0nAdYPM/9pXNgAkq3VclCDi
GShA3NqQxDkmbVNZjuOG1E8MsNPt6Pup6D3WnaIEeHuBHWYZlQcUTLXbNFxQl05ZeAFppv+h19a2
LGJXXLAclkIrkU68QGtp29jCwr5tSj93VJy2Vg+jf9KYOz+H7ZP1dhMsNG06i7HcZCIsyqAU4n4q
kSnsTOfO3byks2jKZu9D665wInWjYgVvyJD8RVH0ifG0VgHvsJ8HzNQPn7Wm6ZZFWv5J8LXcbdq5
MDYUgP5p5+EgYcPad/DKr4MVhBWv49IwSTr+fpMpquhnp8Iwm40MZKFfclxTjfsYO4yqwU50hX9U
bI2C9jxZm77+sSLSRT0Iq8abozddMtQ5q+ji8dJpsk364z4eVDPf1ispz6FVGt7BfUCnya2QeKez
TXLU8cpr+S0UAP/Xw5vuKxJHzxBn4hQMxY5OJqYvSyw5fOx42JrybWU3rW4yAWRttIm8GAjnu/SM
Zm3WhkPc6ZphClv9rz+n9Dl36c0+bhS5kqiualA/UTcyz6affen6NXawkCy5OFJZOxPrRmsjwQqc
obtv25u8pWXf+gBWAvx+2FRx42zhrU+50eM5d+RIsmtbSYlQpNQWwRMOd5fEjOKM2cshHzOhqQfI
ofiMr1/MrD5BbYiivZef76VOjXj1+yEreU5VJFtkAM8H7G/MKYnoMFzG0goTbP6cB78qlVVwnL8e
Rgue8YI6lBkW45Lc2+6RMQY2Nfkxq48Y4SAZAp8W9CbsZiF1a536BDJSCT3t9HEN81bBzzIoyuxZ
dyDHbwU1GckprhEmg40MB9j68Pp6RmHXt50SmYJj9uZ/QKpG4U1+NQ0RoWnIW+nbYOLyfElIcrCc
sd1d+SaP3D7FDsO62V5xjAr+F/5Og7fKiLHjPDWR/6dUfIjmXbOY9C/lEduWh3qdIFdagUUxFRBr
LBAFNKuBwgKEQO23a6bDOqEYkUgpD880PoUSpFwh261pHt8lrwerYNKoqJuW4m4vD+2FGoI+e4JP
pdt22CD2UP8c3kwYFs9H6lJnuroqjdjjSwxUbkSLOz/uFNeqjH3Dpx98nqI7MH02Fd4GWoI0luSe
sectpZYB4xO3BdaA/z2b/il/V9qA0y4Id6CSwVOhTYy25R55z2efdKiP78F+Uko30guLLeyy5Bga
Q15sVGF868994JH/pXSm4jBXO/A8iPvYsMmvcnc1VrRvpbpT1q4A7FItszhLIdX+G+UTI0TmtaXz
pbKH3nB/zSx8C0XQXKbYjGVSNwuT6+gCxKNJS2VWdO+Lny+IWN9W5kTiaNGzrm9hj7O8fkYlgLNO
v10SwnaQK1vwc2qiWi9iyR4UVQ+5fIKgLqZ9YdZeYJ9Y6paiMryNhX1++7NAo2rM20QMkCjWXPlB
/iuySE3JwusmN5I6/AmjsmKAJe4VGReoYukO72VwTy+AJG4aMFQrd0YPeEqxft9dDpvo1sWSFPRi
5eW/94Pp1gTtAdP30izJPtbRQUzQWEy0/Sy5pyIqqpgJTDGlmWAHinjgx117EwWieGFm39C/wcFf
OciIvoSVv/cFFqG1iuFsFbDDb9QkR1NLUV2yHpxxqcLMNKp2rcY4NZbOXFRdDPCBF8yVFRn1UG0k
lTIso2XKh8bAeu4h0eTIebqukqodx3lfAj8u8WIEEg5ULb1BdmWOAEK369k81NBjV9cJ/x51Ar+/
l7xglcsbqy2Sml0ms8ovQBfrwZkXWL0CQPg/BBAZr60lxcpKnYb84vH5iA+SBqb8wrYHOEHHMY1D
Obye4+41P+u/3z83aq/qf0dA+s/c2SXiMz6JIqdqCFMNeixM66mdUkkr1D8jjZNrnj+teynGVdMl
Lf3hLLoZso/bNETYgfQxw+fbU2MmMcsRjZCuSmWbrd6QTaCO1eeS+Mxo/X6z1ByCA5GIjorUBjZw
GcIPbwcfuU//+btwL6imu5InGBpkKTyaIMlCpCRcIYlABkIAcLeoii4rF81KMzcKnShmwK20BfXg
6huAlwW9OiEM2p/ZZp4+yGKXIrxv4cB20l+xp8Iv+FMSZs62/NTMs1oTdssy534w7fC/2ICMqLzj
Aj9t+lD8f5JJPtnp8aSV6kumnmxkrcAHA1drW/S+CkHK332vj6ol0yPC6ChF4FOF4fsMNVNHF2Tu
csIBLvJMThAZB5a5WUqaD7mkud5NlLZ/3oj5KBTM0z2UlV5MPMpDGtdF8XdWWdOavl1qRxgsynU7
8wY7ag2M10CfU6OWorzcsL/QyXKkdraULGyHXN71VWAJe5ZfxuUxl5MTYLNsvO38/Q26KudwY36B
fOebwaPISttLJv8/HnnfDNKoiSb9WGD3a9shvdwHvO3h8hwHVxEe5UR9cAhjONpYjIzSsk2DwOBU
YlS9AFWAsoxA8VO+u67a+U+OePux/VmuERXykbWuue7fvu3TNkWh032JlhzihVfEvXE3XM4OBEiw
o4QYKhCrHQmnU+c2hpb4f25VwEVGargzpBwbZ80lzIRqMFL1Zk12FjC1iJxG7llBUuMr+czbq1AZ
ERcChTwc3GKahY3zHgayOEqIkzGF2SLgPhGLZWLG7hxbuIzo/MgkreEExVgpTcznytrG784vMy3/
KSlcNQxlCPxtuX+jGITZge0Wo2i0PwIlbe60RR9DHV2UyXq74YSHSkEcpvnB2v2slgFbUIwssSgc
I2MP/yEqhCvaNbjtQQxaMpvG85AD4dWtTLDHrJoa3yyrjfhbcbbmf1HFnNWrXodkoGqyybgWisgY
k5Gc7NwUSjGHXmYb4Um5BTuHhuGrQsielxPnDr6LEKKyRujjED42AppVtY/ocpzMrs+/blnWWpRX
9a19VH4gWX7OcUpxDvy9Db/NHf+wzL/kK+z9nrh2qeuIGVa5i9kUQrajYBEh8b7ZVmWdtPN+Wxro
Z6ON947kpAg5pqyE78bqJAa5TQKS96nnKuRQ3NOtDMZBXv/nstkGAWxQnxyTYuGTgjLVF8rvYmaO
qXKt0d6VinWne6XK0+JlJKpVxBuV90QaZHfA8Om4WslGtfVg+42BHFdtzOSrYOBW+0D5DnnrNM8I
y7OQoj9iFRQJVfxvdLZagKiQW1Of9oyeNw3N8+2h+Gdsn6SrrudCwOeSyC/MY4tMkhmABBumHJGu
X1KD3pYzOgPEEJ9oSlDBw06fK0vKgfvfaZXNpeX+ITdW4GulBnSTYSbKww4xtIjys+LR+rtxNDnQ
iGqgPaMB/bw7VupeMxt4b2CXsG2MfNyAFy/2KnmWXU/+E37hwl9m3gCJckMJSEJISoKyAxpAgPDP
E/WPF2JWWDBBJ5VFr9ypu+k4S91yNCdOoeee8zH7frbItUxItOsHvLfNwo980dZxYdYr4/xpSt/2
kRoyVDCwhQ7pDm0gXnIvLD4ge73tuZRUid6LdFSd8XyTjDFD976Kibnr2yBq6Js1bqgC4/1QPlRN
YqgSSw0vlBHfd6w7cagQ5JjH9J2Z+6VKy3vNvZiM0DDVlrMIft/h6xBOAyAelB5XSZdbAjm87FWW
Zd3JpPhuTV9gDsT317Viw1yeSTN70m3DkEcdbrvBZ8Y7qO1BftWkNo7Ihs/cfXTV9NViow2gIhJW
d14J8gXpyr/XMZxCyDdhLsu4bnul9ybfRHmRa10M4Vnpbetnxyv6H5pWgJdDraeMlwad8ptjuExY
ZEznb7V/7sR4jrNLCCMfFcnf5fsts2coTYtjjpyyl9YYUYUtj3qc0wNgOT1BV4Brk7p0sWyKKfTH
91gTbaRCpE3SLTrBk4Fpd9W5jnSev1SioZyUTgzgSByzc4x+gMRw45HwNRnwQOuw6n2m+ZEyP8q2
2JtU5mNH1Bfd6JCs4Qqw2i9sZXxH9WXhzdZbSmn99wB4zwxAijSr0kGUJrhZnWmQa0P7rcg9+HJA
5+g19IqpO5U/Mu1Td4QPZcIlMXG/L62L7qzpJrtOuWxuV7hD5nvS29zjC3A/VgXOD5bj+cMnE/8f
i9cR1rEO4vIhDNdD9hiRfjICkgjW3rAVTILeX8v9+FJy+YClJomOLJg6/9AxqwVyQ/cY8+C9Eo0M
SHRGRA1LhvhcvBBoIZp7Cw4/QKNYMDaDPi7NzgaBuT9s3C5j3yUuxG4pmiVW/ByI4Q9Yjd33xs9f
NYYMASW5NU6XzL9LtukcRTxm4n1C44G5ylOF9Bm+2PLNYk4+7nQXMwJv+6eCIXTSSzcCSFJVEWhu
cJmVLwZjKGq5/IuZu3niU5Bl8nSrhm1xRHL84YVX62MbSpzILZ2hH+KhJmxCDOFhavnwcEe+uMbH
gL7JU4x/Sl74ukbODZszFCDPXaVdin1+CjAs5a80JPjOdXXo6SM4hc4URo/+iHp0OGetfY7yx7Vc
6+cohBcHB2Xnsnr3gwdl0Z4t9WDxEXkR4qfCUNB/FdeFXRwZ61opOD9VnTnyA5x6wMwgW1wwaKhK
5TeKXmRzeLmqNeQWu7Z4rbZHsOUmoqqPmBQj/Bz7rNwNZpSdbM3hFIeAYBqzX8iJNBOQ0DK1RwCz
ijeKygEAcK41oN2TDi30R49ChExV3cuy1VMiLR/KxscI6rHojNDQqqP2u4B8BI+SKXSYA+uOUsjl
l4iqvNDhG2D3jH6zXyW+Z1NN1oLFZgzm7NGk5RRC3sYD1E9xb6PqoSeUzevTHWXIkOFg/RrK8Ol3
d2H0K/4MyoL42XJiuKeZTCDyQQZYq/QfSnN0jkw+Z6p7EwFtSRIbec3xMvnlnK8aQCkgbD+ZfUQd
GfBu8kS/xx1hnSbdWpUk31FJXDZ6QhmEFLVezGQVC2WVDqEjdFsoLzcWs005n1fTiigRVdyxWeLn
WXa91iJlz5hQVqQ1jtHBU13nPRgOf0fB3+PJW9JYM8DTh1COqqkc19YFSX5cI59YqGkTP2Q1EOyZ
jBcfiHAuuFXCaCqsjzD2Vt4oOhT+8Jhf4mH9gAgAVxmGMp630JghOpMRtgDcIxdGv3INBE4FKsRQ
anLsW9qZeAkpyocerPlbmV4CSxchu4cid1RAvwrIaGQ2lSMs3iJeawKkXyz0H/mIN3G/il1iBQCu
8hzf4/E0PZuEsHfcYeVDx2iUgj05gE7QUsbVAjCtzqS72yeetbZj9qY/oCRzEpjSHJcb3oOdIm2Q
azY5RdFmKh1ynJqYUMfmTdgH2Gyv8PL9W3n0pxHDKfsglPbuotXI+EoYMON9fKr9esIiunVaIJiJ
GA8ToQxbfvulK3+ArZWnqtT5s8qmpnsDKTIGyt9i1LOwbvHGaBXht3NJi8Ntcl3EI8PY616UXWvv
1qXNSW5U954SOhquZ2oF96rUY81qD7zZXbecjQnIjzfSaeEGA2I3nkXVqkjeuOJ1ICNESKPJKMpO
b0aX22q8O3edIRgHIQY5g9Z5MkMNSWxN5zXniAXNZHVp8TaqPduxi4winozPFGZaT+N7Zv5UU5iY
GoYUpNNQ8lqFf2QKlltRjP+u9JoGh0LXv80C67SYF73SO9qoo2IFfKTAiS5pBWnWPZ5NM2oMN/Pz
TH3aE6q41UIkDgnOU9HWksrBUXE+LT5TcjqoGWtaGmsZse5EIaRpM3cnTZ/8n+oQNQdyC6boaLkH
6KvlwqzcPmQhlmEG9AKOFoOTec7GtZXoyOM63IsKd5eSibRXkKAnPKdj/6jVmDN7uMBDkrnM/kHC
1X0362fh4+Ge4jgPXIm7VJ5Hi1kZ/+EheL5mOpAYgsD3cb7MuqOEF10MSq7sr+BLsPu8sIHm3fK3
eHYMAplKGbBFvmeayoQgi+a/cAudNiI3TQn32uC+Sm+rHT9MSBrKOmikUeENVSoOGXAVf79eM83e
abzrGGf+Gca00HKIGJVYo22VMHEuC3EShpsqkNREJYXfyTR+AsGSZGYxdaVw5EjGYTWujsx76Vsa
zkJePVvAjyeql39YB/LJhW/M3zdjOK2veXiYCwEu/qy6v6EwrCGPA+DDgCXMFjuWTd0aq/YxSLfk
ZkIBu8oxXaWZo6WQPVSogpX2eAkyrnDrB502iMjzOixpKnO3HQEyidPJr2XgfSZRzWYyG7r3PS0M
RtJn7XesXOeapSPyk2MZHiHb5qHst6jn7l3+0DSmnFFod2GoKphlGyZR0NftfDmQLosV4oO0Y1Un
IU2tMQ0MN62NbyzKxdUOFvNL4SSOWVpGZu5hHH7dV+A7L2miwI196bnlJdo3Mw93p6ERfP2KG7+U
9xifGUdmzy7c1nPBfVR8t5ydjr+/aVhKSz0RORjTnKQ4L0w2iBhm2h86kq6M1ZKN5mNV5rh4R+5x
xDSFnIjlx4IUrKeD4PqRvKnLSZEG1OI2KMp/QkimhN4+M9JyVzBrWE6CKw0F7btTL4tIXIOBcmvm
4VxYJkUIrdnC58oj24yt8geoIcvZZiaJYB9f0x9HQgwCMufr4IdiW2ve3s2HpopxOp2YQJ1J5P7z
Qi2WwTC9XMHR/69i1Hf+of5mzcZ4gZaKHURAYRcuKL/IlPmkIThFirNfND03B4v0ewpUSF50C03u
oXy9NixhDaCj7FQvnhqQOtsP4Mdnr/oLAD21I5RnAI5JdSCUSGS7thPMlg5AJeOPeSDJnHA/Cv6q
BPns9VAUEOeMn2tzFbAS6IxjDkDVYUq/kC1NO9M+ZZ7ZN3bJZaqdBG1b5ymwz3DJaIZNTEYNaSNB
/h18t4XLSjEuoOAQ8MO4xYyN1YuL4CqKUzhdhXi8LpHULat9lNgzAsOwmZOH9yuG6O8i49J+jETl
9OUEviLEI1vk7g857kjyRofHDAvZ2LdsV7XNBk613Xnaav53YDdh+kXN/ADOOQloLTsPV8/tuwLF
PVoAob7p1tTdgXyWPAS2rJfiz99vQNpEQv82zqhnrz94EWYWq7O1V6gc07PUAJykB8yZv8Vug9rg
oy6v+oVJ7zNRuYoqr59FfbZ4XUac1Zp8suLCCD+OSQd0Snb6L8A1Rfxv8B674hdM1iBjrIX8UsBu
DdWHfZ5bJbyC1Dz53ISYiBTPju6DNNB6u1usZfSpvITE3ONOwI9QCuplhYHS3WfNgwuC71GLFNRf
97u0IZDW8gpY+UHBFMvt50ZJr+FgbD8JoK5VnD4dO3ASmOgHnKMMelnUW56Qd6wFC6gsLj2Fflv2
WVoEN4lqlIrPvZCxZ8Z8c05lEiMAjEofS3JP9BcNu+62vyyqiPW+9Q+UcEX0ckI6rS8K4wzJ4L+b
ArS9tczekdBoSD+nQH6jOLiawbNHVsRDRFdjB5tgprEsokbr6p93eiOohX8kjANl/rXDkixtWwLx
zSTKioeH8wGik/4av3JMEZAky6fi/RmyMJfU0ynTMaWUcZYPpUkqsT4G23bIxKtGk+sWof1pKpzT
JxhC2FmN3wVa6NDWtBavnSnmCgAvMMYXdup8FIZYlUsmtxI7V0l3/esouKLGy7CXI7QzJkRNRBxH
MgHBLu84vdE9+V9XYJXEFMtqPOUubZ1oXtJsGQ5ihou9iC/JyT70GXnfPcK0O2DBDFb+XzlkS+1L
HvKMzLS7Hy/eueaiSgw05Il6s+zSE5yTgUZxG7FsiELMjbCBGRo0aGLzwZofdateJggdYNxordHC
Nl1xn/LVDeAUpla5JEulnTW2jiYZ4IpdE6jP+jxALfPN6Z95DUH5t0b7uRV7UOLUi21XlIAAsqX0
jufdPH02hjwWCaBXH+0LKSwyJNsIylBuyaL9LOdkRqA/Y604k/xrvqPxV2Oz2D8GOSr6UmlzMyPq
HMHrWoP92X2qFEw94+gWv8nwZgd4IYvR2QpP4zYdqfs/d9SSF7KC7JRnxkWO2hFhigbu7Lou9ntk
yyKxAMLwoSu3Q93V8m3htZDGHv7SOP18Dwa7kwR8BPgabWu1Bcwn2v2L7r+fGZX3qNx9l8JHbSUU
hV7EbaF7UT87ARCpb5OE0LPQYUYwZGsAVeZ7xjucTOwY7eoy2Iiw+B4Z7ai7u4PbNhoYL+xHEijo
HysRGWGX/BYCxN9HcngrlqPmz8guf7FTLivdUrh9m5PyEM9U+eMY8eTFXlSp6EEWmLwqh4hv6C9k
SmgRLO59uJkKoabcZ/WPtBlliJ085DDw284UERH9qxCBp/PQ5bLb5jWflhPYLa6r6znXoAQhOfO8
0W+RAtTVxtfo4thb1n+FcV77IPpBUsMwXMmPCK/RkP91vTfg/C9yawgZiY7BpSKqYyfG3ICVRCSJ
AZXg9MjX0L6bsAyNKJtIuaJ59l5QHL4/W56V43r5X4gi/swrhTOYJyEY33TgTH1b1UBQaK+v4/6T
QaP62BZ80epk23l1c6GbkrpWKLqRELhBPCY/8Igog22DuallE+RwKaredI0zwWqTK7QNzVivpIoH
Q8Hy613W45dJbgmKC8i7ou6rWjEc4z8xnbCV+WZsasf5/Bih6H2k+wTvhYc2nMcfS5SSQWA6uWmm
c4vFSa41nPcaHNvHSgqHtzJGfJIDuUuFj1esrkyt4KUtnZ7IZu+BeHAx9LvWh9exkBlsHahjLHzB
TZCUrq/bAm7jXElFYrdawDJZQH5ZPx35oLob9cSyCSLVxVXKCkeXtQB5owZoaqipCMNA0kYGwksU
jZ+nequvp/WMjLncANZHWy1Z57U41YrpV6+0YLC/R0vkulB8uDfH+aTubXuTpXWczTxZ1s9hVdth
YxO5KY69T6jf3w/jLBVI+ZXB07Rnu86BzmAapsTOUtgfmudu+mUMulgYq5+ZMLk4LKhoVvjwZUUb
x/5sJXNnbItC0EfGAF1WevnJdUNy9Aum5GLxVAPVTlxPT+0lgWdMeRUK/Qcbq/kcpxtVc2+j/e/M
3w+LGKqxpIDyG8XAA4xG5IjEyMxMrJIFVtGpMO9SzL2jTYRol2Dd+NzRgNpJoWspjFrp8N1fP4Rs
grbVJdUz2x+L1lragpFMvnAu4yEvNDl5t/AWb8puJ+c1Ki9QxyAjmfF3QFmiHYpLlw246rHma8/3
APQEw7VjU80QvCY92Xb54px8fR7HF+6pqFh8QaiQ0PL0Lw0/9yMeRVFlb0l1g0tK/aKT0CJXjNdp
QPU+Z9fM6M9+pupp8KDji2LsSxTvEnEXLRWahHiWenF1zG8MJlYld7j75bsh826YQ88Y96vpEJcp
ANk1tn5JgLyJ7bql5NbOm7ahw/ecNIko87nkXieNUHQ4UZ4WuA2vT4Kc/w2b1kY4s3AEE4tTv7OT
zElLi5x6CfS/ciEksyKKbMhH4PT/SNZvMV9OKLRabM7LdTOEUGeL/6of7PKti4SXhmsRXA830Ncc
0rlJ6dI9dTEnBo/SMAWiYUg3I8rJQrX4YHgqrAwFHbwPr07VCjSekU2S93ibCJZrhxqw1TSaouso
cJwBFNSRTPF8L00s3dGCJc3jsSSCzxDVHjBbM/ziQ2jO3Cko9FAg06CiRLRheSxPOf1rAol0IzPd
df1O8LQ8zyTrgxl4c2nFwqlBhG4JTEMpY9ICfD+IGV+MNlkCN1Ws5SFSMUpRckOq1KjuLKMYDWqM
rCM1RMuZzukNgSmyP/9c2f41a3owpcCuNfCFUig0dL0fZ8YbfiauUYOx4yAB+kdxKktkRjv/hRjW
CRSj8nv3/Jc3bDKqM1Tor3+3xNq90y25/N03SRahpEaPjo0yRYnG2goQZsUmdWAxtSrEqM/WeHI9
vN8mPX2DpzKmUs4xWQvwAo8s8tH3zJmRr6e/7WK9X0kaUAA64oAmftfM8d1W3TT2tWh/qa9HRkJf
tPPfg23RLVs6ExlH9OoLv1urWodp/oS4wNeFWwMVBlJpRRmE9btjhtnyL5Pb7ZbC+Xum9Lso42xt
l+wb02yKEO9FExFkEYtDTr8t9zTqQep4pNtSkgX/C6FiMO/meG5HJSEI26USdHfG8r6zB9vvgM0X
7ZsfC9Y2xwLI+eD81k/FBtMkFfn5N7KctRmZQGAdcYUkPlC1VT9D5hPS+ewFKcVMuvFGrJWJznug
NmzgNCx64sfOYOT6YZdmeKwesmDgmUCCqZW3IjEWTbHrG+iri775WSc51fIObCxitooGsWGfDpc0
NhgkhxxMDr7t+8ZvXLrd6tM1Qs4JhdgQ5Qn6BygifHJmWFMZgAmgV/2vLm3kjg509DI9M5w7Mhh+
w4V34rx+eHdXRFZZxQGwwgo8Va49VObgEpU1BcfIVovIVKxoHV1klpg0FcLYDZilbJ8uxY4t0W+b
BCH+aZD+UU9RZMvEVYQ3Mu/GuoQ73syKO3KJM7ymfaIH4b284CXwbbrnLGmMOI72JWPgP1b7MqF8
3IJ4huf8Ml12eFni5w2NzCpiUm9U116BUR+wTSQ+bgZJ0fhfvtHgcnbzn5aMWOqurQkiDmLR/7Nb
SKYQauibJbOaw2seBhxBTH5hLETaNypMfR3EVtF6Kk9tRiHK9PYQx7auhtxmDNZkqWzJotZINi9S
7RFVCgSO3gCnIKQY/wTHdJR9pmlObIPF4yUHEJ3Iwr6Teu/ObN0Qjt+T+1vPaxCrAJyZIT5Lu7jh
GR1wENVLGWul5uNK1kbM+VgOni1qg/OQJsn/OQLC60ViX1xs3YWFDqVOjrlBhUDcWE5H3h5k+YmR
PPF7sg9tSrlA2a6BfYSk1bHAncfSY/1zb4T5oQaB5Ul7k+BDQf7xeOSbStnz29Wf3JcgT6OUlxX4
gly5hXZhQHvTtInBNYJZVFim8uBlRD/jBobuJ7VJb4t2xPZfELKB59894E8jxECa6+xP42tOi6jy
zYyxlj0BL0sDTaZuAbCrVmpVl+gpgmypu7Cfc91IP2Vx4ErA8Me6+LWUkJDrIu7po9zGNsneD0uD
nN9prE9lh82ENZJ1MjKgQ/MB5VT3K0qGuWrezFWKc0H9fmedRTdTjDQlBowcwI+rMhqJHT0fzkwC
FttwbAKih9i+F8+jeenn9qDgNjNGxcmiMGAoO8a3+ysy0fRr1HC0NrLpNalNza7fQjRVDZpUaZ24
6qouj46HM5N4+8KFMd8c4HzNoNe4xKxnA2ouOQ4BFWu+MAujXYeMTXfmKW5Q1PcwHHIENWx2w7oX
y8bFgOeTlE/+uDIMpm0z/0mCP2WSdAKXBf9LMTYMPbgZyxVE1XNMRZK+i6Kwvuxd4ckSQmzf/J83
1sk2Cc/dPsD4ZJdipBHE3V6Smm0r4hiA9TsEGau465mO8ncT2+PhUn6Xm1uICDZglPL1GEGUP8pR
kxWLG65ERjlmv9siEOJveLVSYCxZQY4vnHVPhWfeW2fpNHaYp6DP4irzYqe1DP1hsNaRZrrbJXCs
iei9TLWV1L4my7l5KGQWAA06MSPG2CHvxxUpdENlLBwLYflbABqOrgDwj7bkVQeqxDJ0OhD+99Nq
VXGj3NHAI88Y/AasEG0KpvIbM8TIFy2flDzt7hrGYPRb78WXWbNEqxGNdP8wQwO7nH0X5HVd37OM
cEa0QSOfkyCYd1ruxcdyQ8ZUquLmh/MTSC4bpeV5rK1crGeVZ8XLWGov3nQkPKXMKTuabKRTqno9
tpk7mCHbaDv0fV7Kpiea0d7yqi5rtwAorPNEv7Obq2mls8ufmYQ9Enu9FMfSecBpAbZveVFrAXlr
X0zKo4syNs4XYfRerEmElW3rds1E1NJrjmNDOkGRZu49T6j/bRfD5fY2QPY212aTUkdqgeGgp19D
+X7ez3zORbSFQitpdcNqQ+Pw0LqpLvo+5bExkMBNnC55MYrH992xw8MpIVSFBO7NoD8QoJVNdxRw
7ZSJT3FakAUDrpivxROL2cSsExA/AiPiv1KT6f20TtnlrAj2k4BLyig80c1TppbEW9D245AIUJvo
Cq4TTLMqOZnb9Kq81WWHqPOYYBg2EZuKCr0FR78eRJcIIGVGVHWbNqYH8ygkOTQK4cVx85P+k9Ej
DHyaBY6F6Mc6qzZsMliMPUnJzm+KCcNc6ex+gPGrjhwdczGeegbuE+Jm16sDXrY2kVk6e8fHMeUl
kckHJALKKh1s928ig7k+KfEGFNniSjpxF0Z0pfQFZIoqsFttazXvGbW2CrIYoGcCxcTzhE1TSvSL
dhVEqUb0Szo4h4iSyqSL59imqmFtFCRvAVrKe32RQNGzBb2JZT0J5/96PGbvH3bLFubAdYHkAEWk
oNUAbr+1yAMuA4nAM0q4P+WKo9zhA1nytJcPUtF69T7cxJamFD6pIxsn45yGNizw9oTOVUsRnfTD
mRB7evDtpl6k24Vrksqe1ytyuNDXUcSSd8t9l46D+c8ORQrXp4bPsAJIWsI9xbU8wGvlYTLQnWgA
6mKNT8vLOgAxrdjbq+wdnTGWy3UYVIMo0M32ZRJjpOMzy8XgCi4CmKQdnjD7radQ8g1oLbz3wmGy
27yIaSXzYKX69uqUbmTH0vqGrDG1V6epxIR41bBPqVlJUlMvq4S2flwkPJW8xXrvbS98nG2SKKYd
b3VcslBlHoshx7K3PRjkfZWVk/30Limu7FxzaDL/o5jUYfMyJQviPqsBdAtsQYY2maNklZRpAiyu
lpt77swYsnY8YR7XijfT3kfFVh+Wu70OMYP+EPi62SNIQagYsL/MpJjAWDGbUpYyOx2VPC/I1bl1
yEPgDYNBfp6b7Q7LJHEaDkWOxLeKk49pDYL4uGwaDQ6FauLjCWYWoWhkH5pNRRXlUO9Oz1ns1glf
/edkQ6cp1r0YjVlB4iVjpROfSAFk1ak7pHNnr3F708ogjbeXyyiLYUCZLMhhDnQUrUaaGgzpOCgJ
8hSVGisZkNA+9lri6MW0y2ymWUfd6Ujv7GZgbeTYKMdIZ8vLaNO6c+M/cVeS2B+jzQS38fWlV46i
p6Z7sAsJRRZr5LeYH1trD5cPQR8tFjm+RfBR136tl7DoNG/DIpHhNzEvfosdRLeHOJ1Qp+ax7lE1
d6PQu+GD0wVvpNnvw2nNxegQm99zsOzo+doT25RYlD2nMDAOE2R7dIUB1r6Wn3GOcLntDOOkxeQT
V+VndEBoRCww5ij0hvvZ2e1kL4x+0HQFP7m6T9fCWVWG1q2d6V3tN9q1pgPM3CpORurphvXWOFuC
aUG7iKMyTDXzEEZri3yN5Vs4XB4b3vTgJnn6nO3d+qBCYlIdErUrJS3xzYn4cldx/Ordxoh80JYP
oIz5TuzmrTz2EqgcMO8yBLQTg8DLNWgzkp5JsPfkBHrFLdWuOAKe52cziHJawMAAhfYxbeXvr8U2
iWsT16ydkxK4ICzVFEjIXmL06jwW0gzp7UulVDIrCto2BzxA9lvwaz6ZqAYAdMm7Ze/+E2ADh3di
4E2KfaFFATf4fvHTyOtV8PK/CwosEMF68nGEgGdb2FOXNTryMgEOOvVxmf+I8dGcHrIoD/yuJ0Hq
FsaiSPkTVvICRrz+BTbiuc7+/AEEbvtzUpacEkAVP9MOKGyw3EbKUrXGRpKZ6m0RQPViM4jOypay
+NYK+EcPWX0egA5cr2JWioGJUcqIrXx4rBWqxJGiRwRnUhQrR/S6LUvmHp8rhE1pzffqhTnq6cqX
LTmqaf/GuvSYfi3F84cJEF2p/fg7MvUjir4L4eXN4iJ/iwDCxIT8850vNnLh+o1+kpuQ3IXDNpAO
48MgrKAyedRE2/Mv78J9Jtpr9bKncRUezNMPxLE95ynChKHKBb6WjcW1Pp/LDdbbE4WLqyeWyi+r
UtRu7zH9gAN1XYdAsrhYDuNRf5mhS/hoRRHMb6Tz0p70JFdXIZMGUQJmlsjSU9mN+kOA16FrR+tp
XI7UlQUJPVX8NpTqAqztBIUZL7ivbO5HREkUomHoYFdfeYMBy5BBMzXltECWwgVK+rhOyoYhjI0E
UQ0WDMnFEuM4J6RTBdp8UxMILe7LPQ6fO6VcEein4L6zRCzJUcD1cBdns2msPJIVd0yKsitThl4g
mT6hcDxJHnkqCb0zsr51mM0sQaz1+Ggaa2DcSEeS0cyojIyDm0vm6VHwMeafluYdx1r/5XTlyW19
MlRKa7AdvHlew2ty79VkI/eMrAb3/YT6wzGzFR7LlkmNG69gf28Dm6qeVtiHMQr9re39YIwXoJ3+
thLeZV8gT8E1jU6gdoYVQi+NRnbtkRXl5Q2CphrsdFHTStG07VPZ8P0TdvLSCx5yvcxflFPKPB1j
/PiMHwH1HQwb0Ahg2DdDZcoNzB9/KBKChcaDzl2N+AwMOjMsgqcj4mz+wj6YAMOCIfb8mip+vUlJ
zRGMKAHzh59eW/s8lsePEyZon7BMW6ShwrjIDv2hvNR5/v6SIuR2NQJw86VMSEk3fRBNdVVnc8dw
o/s6zcRt60VQ0b4klpXBVvZSUw4YIsTVLsRkXwKEJEtxEzFNeR4JIDRrbSUd4cMT+13TU9RyPsF8
wTOqmELRmAn+T4tpF35/39PVtuyZmmjLiyc/hdROlWhs7sK/lg86P+GIjhBvOQ1nGyPGTSNICrvF
J0FRji5BBTkLfSPwty1zNjrDwuGnYF0Q0G8GRz0DGKMCRBCSBi+ZS1ac83D15n/sQ+61Uqv50rGE
Jh33FhbcPaj4TkdCGk7U70I0v2CNwjos2Hhat/r/Kc8Jv5e1L+g4xuOtRFDpRnhO5ExeTy40pNg4
36msCFHiSzB8VLc8CRrMF76gefVOQDxoam3fJr1tFJ3km8t5GD7sfBgwyR8L5caZVESaRoPG3AT3
Lj4qz0YOwQyWBhRKWlyGKj+w3V7p8K8i5ZWeLsNLQLxYPDLzfTukWHri/EZ8kFqCvHBpB7KH5yej
6wvqkSM0bdUGMgid+sW6p4rhPlHpPJDrE3DVPgsBQMxrSjMwRjwKl1BliNe4pMH87YZoOWnNy+xK
I/RpIpeOpO5yh0GlYll7/5S55r9+0pUJ5ZkckjUcnZ0MTNpoHXpObNUmkRz8cABpixh8a4LO2l6a
DMBxcTgCobpoTeLBJ3C+terzIKsViuscaaf+N7OR/moV8wEpVs4iNFxSu1ltf2WKrfMjMM+5tSEf
zXSX0F4YEOpU08M7rB4hZfPK9ADImRyg8QYPy8tKM38urR30BR/u6CeZi1tOZhU9CLj/u5u4yXNU
CaNycXi9JY9XfNVd5m1yj485vWn8bred6SkkqGA5va1ud6ZLOGHNjTLAlv9JI8BKpHXWF7O2bnND
WyyH0Jg+GmFYxJBlxF5Bx0ChhVy10eC1ZZcrpeJWLuZETd1UQB8guoi5CG566ScZF9EguBXmmFxc
Tau/gvxKeeTpjPs0OrSgEsm5E8zK1Fs32/Opak1RAeFLefZ2e57j/OvQVuEVkh8BqPsnH/9DebCm
MMfgZnf2ZIY1nJg7EyPj1SPLAmiK/vzSLlnNTwGy0llPkeZnuz9JR+8anHP86p31snXSAOCux19A
S8LqLJuHQ8dL/gMWPNaxinNHm95bGju5ms41dQ1ezU7r4FTYxNkD9Pm/YB7CFneOnvlEPzH82EIm
HqiE/Zbely+FsJjrNGzZphgux3sdlHb7fxby0nBaNv62mSvSTzbUqGKs/VY/81GrVYjfjAwRDK0T
oY/BxMO3F3+iWmuQMznkKA65XKo52/jvk2R7OHS+jVZ2/WudJ4wX38pQoFHUfTUoKLiJSLt0vFID
cfVwtxuY97wToGZeua0ISb+CqcsdI+lK+Ms/+3qcdwwivkN1zOUHd2ikfvg3b9AaKcTsFXudxdKr
STtyUz+LYQw8yrEDZ9u+GBAemUcur/5TE0E41JdBBw8nfFanTlNLN3SsoGhOtd4JwuBzT0QFndVN
aEaLlF5+o8Dbhd+UUGaUV2LfWlppiyGNEqRuk326fTNdZ1pmSGhfRVrSSyfecbA+1Zg+ITWM7XKT
rd+tQU0fE7pVezJCNeL37HjFYMp8V+qZ3Almt/mYioFE+c3tZadEZELSbUu13EB5lCYHMstLsDKO
PVoLkyKi68LFJ/vO7Xx49eJVoO5yfpXOzbUhtyk1AvNU40vjYHH4pbVmjfVXPh62afatJ8KMJuKN
Qcyi9N7Ea+M0fokhi4eHYze7UoSV+eD1q0RprWTJKIpZr4J00lyWOX2oVcN7JXGQ4iZlefZo9lOq
QK6LS7Q0HpBuFQBMCaYvLdNNBVLA5bezRDZaC/19+p8zDoSiykz5lJwUoyFLXEatxoLXpUq/sjqZ
VUUz7HJ9tGH/VylI/Ej8x+gz+prCEh/DEfkhl4jjPvM3S5/aQOuPEc8XZapEWxX8abeGUqjlzQ/0
6LnkIBhzNPl0AvDG8hskLE3BdhbTHJsax53hzmpUJ/bFib8n1w7iHVqBY24Xj2ND+yQoRPitXrQV
lyx3T8GKdQekUGCtThq/y8ydzmgePukdX1K6Pym6L/JZUfMkYg2vw0moHyzp1D1wsS4En1joiQqo
d5QGXCcS+FY5pEM1czts/DpiHiPyvibdA6z3axqIVFIqEeX2/k82b0obWwmdGP/cc7hTI9KedaRC
298jFlSwGGJa5wMozpG8FZN/xsChRro3LWUxTIAanJg1nMhNLoJfAsIrcvU17vrT+aW7BbTeM/Tf
qnpOBiXasVaRziYExxvPwIEVKJeKUhEwAjXJioQyh6oHYzciSoSX69pgyGt2OYUFKIJ527+/Qwb4
btqh4tO1Uc55x+bdUjZFXBAohjUin+ui5qSJFE5pKf8EdJzs4a0pE2WgajUMrNivil7T8Mhk3Ev4
K27AF6/86Wwh7x3777dFHwf/e+4qyGNJ80uhpE438HVdkM/yo+025oz4TuE0akz1SiHJcLX8db7H
nwtcXb6HLlQreDJjONlKDBqqXTI4ldly5rHia8K0f2yFqMrG2Ew44tU+ZtPq2CC/zgSDlwz0Cr4a
CV188DlG7Z+b4qDOSKlrXUGtZjHncD8/NiRDfVv/V7sERS6GHqPjtDOSKBUmVIiK4CLMtSr26NIq
FOcVf/DESkIG/CIXICGa920xMasETlEANf8Nf3TSD5bNVh4RhyD6GpbdqE+6uwTZk4QhOeoWrqmB
2xzhSTIXNCKMfqEuHMq/rOp6dSDgQj91Ofgepf3ktfjkPGseyUUOFXK0qSSeCKITKiQ3AsGSRN3h
L8y3FJLCy8a60Vnt7lqPrk5Ieze3RgqknR9hlP8jVLXg1Z49Aug2QUryHyVrBEdNvmLfN6GGE7+G
rrfxrUe9HkwPzlE5BGf4Ktx0DcLDu1CYM8wTzDdVWH9PNzwZRlODMkwqcW9TjozTpF6/4G5W9PoL
Z4MC/dJsTV79827lLRumkqQof5MdbsNv2TnxcwES1WheOv7OZLnbIAufklTGsrrRCPZ0HD7rNzqq
POJVZW1na1szDKKJHhVS20DGghk/eFN8zFo5u8OQqNOUlM56igdTFCMzk+6pJYaaKQTFTyRyKke2
ZlTszh9gNt3HQRVr7Sln44dXwdrInVP5aUMnaBsJ2swz5//sqCSJ8EWuYU4bFAt3QLdDH5jpmzPk
GVbrzk5KuVmGlf0q21JIBHqwaw4SqtHO2hX+2+C1dQrg4YooLwScy9HnF9eIGEwGhDN3AghTcw7R
RZLFuO/aJfZsvJstHsEan/7tpq9W8gIRdKtr6TDcvPn7c+IdEYyz1luRRTZkIZOK7XvvTZGWsW/g
jHasTVNkT8HLak6FfVgMPJugu2slqUCxMOITPe75+Aee3lSKDOClt7N7D129lMs97rWsqPeHe0uv
aNijFZ+xm7zk/FjYwSitXrDAJa7IQNjoS+Az2RjEGVtLNbN4BNhItqV1JIei+7iUeNOpqLondPpU
c1sjjyAfCSrvSlBADgs/Z1AFCrBImFqoBKISNr0hrXov3pXxnUGY3LIDRud6ee2N/k2wwHEFEDei
29eLIWEuMDb8UmcZHH8BY1dngJjrJqFLEoV/2f5F+DfzDiFkVoXif6YgZaHu/sZA2QjGZZyfS/Zb
yNcQFgSJd+DRGp7BKI9vxJHZBQDPPqaYZoeO6ncou0KhJvq+b2U0mUz0qLe5lMBkHg7hxjavS7af
bw0CowG0rVgiU3ijyFxswNwT2xy26DP3MCEYgG4g9obolHv3MMXJgzOYcnphJeahGbktJiHDxGht
aZ2lU64kTh7So5PfGRSPfNrwxu8U5IfR9b4IE71w2yS8CVCFNz/lQOZumIIDB0ACgXVxltgfgf20
dXX9TN7HIAw1e76WbTuy32XROLMFyAFE1lcGWpVgevHIscSq/KofuRYvMMjA7x/x9GLi4ZSTqlfc
q4zplvCd8pmrQMXUFiGL0yNVvRD/cY60TSguW7/MClaHye5dq6bYbo6AK0INy0Bpu1A0ynF3HPzS
c8K8vEDFdMRgXCTb/QjGPhXAGCQaHQ5i3apmvGjumxPqSh9d84aEKRQVGyHn4STgaQ/w9vJyacE/
JdijGhBK4uelSEJnmpWDVFUOZjDGDYC1YjHmme43ZhM5xJ7/j/5CBhH+M2x4ja9xiIze/MefD+kY
CoLtRc6SRzrpAU1lKSpn4X3qn+E62uTBbw5kSILqLrBWvTKolfy/l2BPQ3oGXKXlL7Qdq0lcRqWD
Wc+mIoX7b+LPR3KoBsMTe1hQHECiVXLXOAL2eM4bdqc9un+AN9ShuU5300X6Vr1NrYY5sAaUscPr
9jXWR/BZlit20bXOzStyRiDTxG2VIWalxzo95ilSHU1FysXF19m4aIMlAbFcZyMusUfyDjx0cT5J
yxd1P/2cMYok2L17tu0OMFd5I76qhytK2Vtq33G985PsqV+hOWSfv2eMgWPM8Vvkc/0dkijijmRI
NxLSrk4rruxLy2vlDqKlZamtGat1YulPhmZCgNiIOLtdEbM3R7j1pfhmI9+7kJPkgVS6oGooLiK1
z1/WKuE5dt+7sKYZjG5kGWPhFT7HHOWOySLUEYvoDfJEOQp1OBNNDGzbAppXDr/m6qHAR61EQmY1
cn4Snu4m1ggJIN2Pf4b5aGr1ErVidJvKJedAwVwT8pUrbPkF0iOyVhc4alk0cG+5P3XYZ9YJtSH4
fwLnirwiqWuTrBxXmUoPOGEOMazBRPra01dJRH0PDvq2vg3SP7P/n2QTXDxX6BrfiRcxsCHL+QaU
G5jhLIcOWjvlNVb1fbqsJEL2L5JUkZrHuDtguSlEL1HlhkIYiKtb0JYmCUfFK0sIQh6oxv9/LT/x
qq9BHI69XY2OGCNOJ+jEkLayr+wfeJ72sGKhEkvVEPqzSAkSOIHB0TCpntIv+m+QVf5EfRuR4HS3
ILyltqCwdEJ+0tIXpCe3QaBvvyonqGNIlutcgrhPtW7uVCrGmhwU9rFhkwr/Iyt0Y+4u2HNphQDA
Mvx+8e2Of6JXr18U3QOk0U6781Z4M+he47HJcJyJ2m7D/yOZdSywyQ/Luv/jNuaIJdp9SxL0/Ebz
Nl84bQz4ohvNRYiLDHG/3xkm+D83aSRxYXKjr/tBypbVt6H+pvcDE1Fdk+rM9fxRTLp9pANHU7V4
WGFbJx9QabQLgTdlJjocCKCuRYLBIwwSjEj7Jgwa3zJt5iLxl5O/70B6Z3/E5WzHYiX5k6LOfte2
mUk3DelZimrf6E/d6MMeOSlLTSVPOoY88ovXNyP+uec/KlDNsD7D0Ol88c1cWiDGGNSk+u9GPoxu
7ZkjdqcyeDIfWHZLqC2o7IPT4ckA2fjk5LpojrunElZRs9r1UfyeMQWv+12te6d7tjh/qnKIb4qo
opspmODOlMUIHtnbWd4k9tCtQhrsANRIoxwHptl2s24sDuR48ne9joDveCgGqYrCjqP5aNrCbMIH
reXUSmkSwvEOv8EAtkJAzw6NpNQgMAYvx+k8zg4aKf1bl7k+4ZHMW+63qkR9nQeF5VIqw4spQe+o
3CAA3Ytps7uQTYKAN+eObqT3u2/GC26eUphgDG9NO7MVrnUKBkRlN2O3d/MT9IalWNltvXvBfL2I
Nr9HfkKKMcgZ8pguehSsRc7aisPQwm8Ox+gxjtOemlRi9qWVcQ3yd4mdMqxwDaa397hMIOWTuwL6
CJdZAM5E7zd1BYyjhp3mI+R9gtVmkbFGRqL7UsGQamC5v4wwrEOapIPBgGYz5lXIo9DQgSU1u8k5
s1xo28KjL92VFjROfOuvupBBl5HI9JvqBIxD5Z8aI4Ju6WxeaiC5SIRJJF19xycVdJZ4rIKGwQwc
gGLgDO0Wv3PQwubNbDlBeWUy6kGHE0WeANHjuBwAhKBXByxeOvU25eVCSeDpxvAqxrKCxs3UyZ6A
4YMHWhFeZNw2OoFETRX0lQkohJrjiqNG+n+HmYKvfDjFfXg566yTHySb5N1gxaP4nYgA9u6v+oUH
47x26Dh6oicIVqIInY/sQxmsJO9dEECk41EmxJboTbpQQbnSU5qThcS196vlq4EpISKHP3TJtsVW
l3GLrNsxuUzqMjBEzlXqnqSi3PxBhjqKv8Eyg/I0utQx8rgRHaCt0ZKpHxXWXL/hUbG64uj73SX6
IdnPpxuM106DXUSt2P8nnadTVQ/GMw2fkBIW7ZiI33Xi9TQzLGMBdem939XS3P7OzF4u+DaR/Mc6
YSwaHQnOxzfkthq4paELFyeCzQ6SdxT3Iy8zbjYhZ6So0MYyLPGuPltVp6W3v32OJdU5rwuoDfWy
IJDgNodBOjR87DPEyMxeo5kDrkTboXpO22eYWkngXxxUxS5oywcfveSz1FeIcXXUE4Tj1t66SpKa
dnDInP7aNzcZc8KKD+4289SW0J6TcOUksFHHeMaHyD3iSFbvxUyZzSJ2t7SjPvSHyUbo0hV07LV7
hRAJ3nutE+RZHCAHPuQJ3HKmJ1yKoa7sScqklt+6tS4L1c8JOJNT5xPH9pNRb1IEf6Ju30FWJA8p
oteXxFb/NTQ6CwDbw8EIFvHYMvPYftFJDVNMg+e6OOFGK6e52b6ocoiasv8ak2BxiEciQTs286W7
zbzF3mNZyEDX3RuH2aPn9Y8puG3SWk8SPnLZWYhCMG7lrzFq8SxOYJTq9HkqYYxbkz93YsNkdgVk
j/edjai6PQeHGC2tOhTljPsRYoPkHzGYgQVHih3PrN9PGjcMeVnOixklp6HWPtOdBKqIE67/m89n
WQg1sL+pfCHA+tF1oUerkzJP1oH9qA7hZbYWdcM1iTimI0LEeCgjY67ee2DEPoVD8nczc1ofdTl5
vgsiQrzQQ4Aju5J4rWPj2g0qHKT+wnS4ye2S/775D7Z6Xw2wxohPaiin3tgcqAErKjhDrFQBfGBX
csw1go7owDFKpm8PBnGZByxLjjH9CGwLwIwZ9cZHoPWzsTTkpGMmASgNPHwC3czMTMWsjKZh0wm7
H4w4ZDVFjjG+QIhd1CUbzgz+JU3cjLbAMS09cdPgMFW3mOe27wvO/Ozd0GObZQJoFJjAfwt1J1yW
HxonDTU/C26lANsCs+MYfbQ7bJngUfAdGJgktNIae6XZ4k6/hoVZ8W4D1vFjRlGQZJFRhqtm5r/F
P1Xz9DyAz9oUu89AdCg5PfgA4Mxm8Awe/UBXyb6qaR+IJ47fzj0GacKLVTuMkTXV5UAxuaxQ5B69
3upNrduSpOvUDOJx5ny/B7qbRV8YyjQUI6u1mJS6MUtyrdsQ1TFCTR5JHtUF7aGUuv6E2rFWicmb
a2fNNAi1ZJsw8a4knCwOHLRwFUSWi1xZ4P4ZGvuM0o9JEdzJCz+zLvGLv0nGf/+NH+Dnsjoj5CDt
Z2gSyPlpBnuG68eaGt+vnOzKCNaPOryxuoOVI7Sy0AJrcfirm+UI5pnFnwFlPLBvcNoEZevp0bq3
puFrFm1E+AjhqMLvxlvukgAwwLoq8cXPVBsG21hS4J+jnU+k/tjgq5cbxdN+wb2mVGIYDE7B/ly1
R1sDNVbGOznl0Lcnh5cW7qpiBbg1HlLkPXjpvo8bCY/DpX8uEcj85XCZ/c9doqmmO5FdmzwPyXBX
2PwlOBv6CWit6ROzfFQEty1hDuFBmkzA/93ArKVM05NltQPhc5coX93FuOYczBD+EsBgVqHgK07H
jSVhfqTVw+2ye5VeiOPw37pBtaM9KvJ5pBiBPc0WmB3t7J0uix4H6XuR1uvy2jzGYfAHxazIKRv5
EYdGti2xHl9gyS3TXltVPWSB3TVIb1mbpdiNgUiUqht7ojFUK7pzjzrolRTNiSjVerGQqZmkJic2
p5FWVdbNLclH6zie5hNj0WnegkWSdtBw6PVj6KMXL6V52DKjjZlJ8ivU9GA8MQxERQK+sV7IlEcM
szNriCsUlv+hSIvQ1WAmMCBobVifycBFyX2D8cCwZRXp9pUc35lfaxqBbjsJRQWtj72/wSCi3UYs
zc+N99rNHAnRVXyqngF+YCG/5lAf4r72yi3KNMuPwgm3NeZW+CZP2Pbik9zhM7Jxv6HIckqDNlwc
KnFz+J31fFcqMZLGp7ENxvTilE7TAi1gIZjEuBEkE+OxrNlpYzf1xBpVugDmZirALrXLPOXPtt+U
TdHaAbBr7UYdFNs/ACBSbqa62Pj3svzb5lK4UpLjDTgxJh5jiGo2ZiHp2H/4EE/ZPaRovVJuDALO
4GqgqWG3JlC5C6I3MqiDNSIoenFX7eFKJzOAd5/jMILkaK3urB0PIYfDU/oZLHsqXxL33gEPg0gJ
F6P3eYFYEXQUSyzhw5ZJq9F+g071D+eR8uuJdRuMrwBC2X7WRsPkvEFfnuBFVO6fLJKUySQQT68D
fyx6brEIgibkgTxSZs7z6lBFzeH+yQEaFUr1liy83SYv0NmMjgIbZ7XJVZnH0JXxKfylJPQdszkd
p5TqvULOjEpyMM0hUK+BSnWK0EL7xbYEUfEV8e+L1E0ulg1dFZo7HH/hcLDqumPzm6L5X8Evnfle
isnE59CLLVGhfUZmWXObUUFWwW73FFz8cm7R/tTBs2a7uRScOn3yqC6IylowjKBPNDR1lZCwMCL0
QW2m33DWvVY06k39ZkImQ9B2roqLi9PVecj54BpE7qUxvfMAiVVRTKE9EZM6hEW+EBrshHe+PLJ3
5AnHitdm+Zi7Z9LYP+H25FyDVJ/wV5wOiSH1VKIoopO8wSKG6BIaXRgvej+4z9o2VuEkD4ItyU8f
thrCpVTg9wcGRSdUIS1nSEiw9tvoCgirwCdWTarQxppOrBuU6pzr12CGngEUFE+/7Hr+Rcc2hi8N
o6oJiUrLWse8a0DHDF6FntZkC7d4FUaU3DS/Fr3Za2QBRvnoE3JxfbnkQwjOhb7Pe6yE0B/RfVy8
gvpco0dyO3fkiSEnRzxymdfFsfUmR8Nyyizd6BzmWHoyo6DSD8i7qLwyGolaYVJu9TGUYiZtLMJc
0SNEyQR9k788ODZhD3MDklKPfYQH7pnRBZa+XxQtsRXC+/NtW5SbQOschsIByspuRU8xgEjX+Mhx
bHqopnSPctauwrWHvbOnZjMWvjk+vMznlfNdu5Kd2zf/y9QKn+B70Y1Vl3n2wIa1jaOfLdHjWb37
WPqA6aDw4Mhny+3LtpNwclWfKjxQzsg7ocIsM0ar1vbkBilsrc3R/on07AOk3kIEwjx93fFkU81k
fzeLXA4pK2fkUbXj/eZ5l0cRcp0SyUGC04h119kdU87nmh4ETzvbxH/yHvjH4S/W9TrJ6ejOi88B
/5uoXdoA0QuL9ZGWAdg2ZIaj8AVFPTAYuygUWSyltiaETtUVdpyErN9BXV7u2NG4vfRWnhmgu9uD
+NB5OKLPPvziav8zA1brsJAErJqPEtLjIFcJaNcAEtoai7X1pfeVw0hStH6wEy3VqxdqpjMvqijF
wxFRdsW0bUC31FemzsSo2X2Ic7urA5nUAuOudkHEDcLeOeAxcV0WD/+mvejGIHrj8PBwOg1v3nrx
VT7ipg327iZrVf9RoIPZSe4fWg8sWS08rmX33u/TnxOxcOe10KTWiqlQJaWvCNnkWSVM8vu9FsGg
JvZNvAqQXzw5/jZLfdcZbHbx+O/Vwhz1mbMx2iSxX6sVkyPHEBXjaBfuVZmd037hRRO72Hu8xjeJ
z6f1WY00fJ2T4hI/BrJEuYNcr3dYkUddVIkHoRt1MOHpk/JCvwF5cLwb4dOqO24hFzdN7+3/aJ3H
lut1rM4XW5kH2HOKTNLRfVBWvLbcLooE/mOwp731fZ93u7bM+VzparYzpebT6gyKnWZIWARreugb
KFe7N8Tb3APFJ736EDrHTDvveZL0kVYh4uvH0XMSw/sFLR32aSyDTz07tZtgCHfpS2xJiEpmLDHq
zSsHlHlVOLhmf2KdwOPG18BNH7GjsnVbixPEwA3Ii0tzM42RWYGGliGBOOUMxgXJ4X+eLKl1+YCt
YAdqVSSX5NDWjpNV4GkmQxtucV9WVJBXxaqfPCNo+9aI13Wt9LFsnQtZHC9du5E4USEONmohUHyg
0gOtA7ohvdh8UwwYvqSBFRdPVLTdAuDprIiFpBvDRfsdn8Esmv5XGojy5bBG/HXWsVxS9xorLz/2
3/2J9O1T+8S2fb94mxwoyMLYd/Ecxz/ewA8jb4jJVoFCN+wFPOcHelQmoN8Uz2mLW6sO1i5txsXe
4o1yBXeN3vOX1YENpV/CtAyhmIdpK2vaEH5wMyntFAAK2SwUkglOd9V9TBEwrcvIHp1n0vOZDzNe
ZYT8ncelqyMO52CHrozxpLWEahzQhAX9i3Yhd0HzTJGF3CG2+7fGutjObL/8aQFpyg6y2itoonza
yseos1Vt2Z7wM25NKPm6NIm1H4LNiWpB13RHYvMZ1jv2PMQJVNmJIHIhxT3wTppwULNSsOYLZlCa
hdCrlNZW82A+a1De8jEFOwxyN5Gr6DXC/Yu6sXhYeKdF1TfZI+nl6qA+lfJjfHMQo3+TOhh95QpQ
BUfR6XQWnTPPEKSZ/xY7n6i68BhIKk8B1+2hr7cmQU5dn1x1XNFo6M3nQU0OYJVpta+OEud/xzng
Xq8/wr0OB4dVlXvqIRXGtNFW58g+4mFX4SVuxb7aHVxysCeTwnipXrndBcMuM9hrIsQfM0zgKaC/
T3lfsXaAPOhG+Ir7mZ8cClkwem6qindyhy+P6RsOAkOWDi8esQOyyNhZl5Tj8rVxXxSD9Bec08FC
3nyhJJ9tGssrfNrBsYr94FQ06euzTmPIZLFrc+0foNJddx5gC9qq3JcyG/VilA+HI/XvVhWXNWGz
UPuvb5uRixnoa7DxOIHaaud5S0K1C2UrCD3RBX0BzfWan5LhT8qn2ju332yiJQD3MO1VaQrR5NZG
xPFj8siqSd/tWD5PNW7iLzo6QQ0+p35gttBIbKm73w01rhXCiKOg0JmVxYDvfY+Uz8Br4H8702q+
OWOuBJ5JnOH+EVu2iIgt6JzUP05xUzwd/uVfksZjo4mGlfcLM5IYYzuskZEBYIuFnqhRW6JWqQ2v
nFJWHFLdWbMngYGVVtvnPOGPrK0Kuz3Tozrp0uqAHAQCQMpDOROv9Mg3Yp2RxlLMW3UbojWkmjED
42nYtQmY+RX5XjwVKAQKZokIc0Q/kYZzlZFCyBS8AYiaZlXc8T5qadWRsEEfIWB/c7sepdDN5CHb
6ni7mc+2GkP5M8AGJcoX9AFpzvOECS7x8LY43+PhAZxbNMfrO+5rYYqV6Ieriz7RIJRW73fMnErn
8EENVFW95/zYr0IQu2XofLMe209lkJA3oc7sJlrQ5cCqZPTAdGHxg6OUJ/rSziIb+JnLC6ZNavaY
2wrovhgZ6nbHfdBfu+CnnkFLe5mUJq0BLeAXwIfqFQsA1N4u51kWa/98kttGrBSbQFZTFh2XYuJG
PuDKzqQaX/dLJRWbrY7jmPn5SIj52mHlqsaSBC8XDkncqO9OQqQW+fk2KniZ9wbwi47nR7srMqaI
F4ps5gWSVKb5MPZ5QwgmThSGm1cyzRBFhnrHUhAbDzXY77U7gUc8/J33Z865YjECoWOLAmIViDoW
5RLdktvPZ895wtbXTKJ8cs5d1D1mKrWUC9T4Udjl7arUKUwFFg8vEEHk+6RmWEZWrCwZpkGior9j
t0wObE/tw0JAGAMSW/R6jJB0fzuzaUY+jIvviDcb/ooenNUTvsL7AA5rCOTKd1TRRk5r8XvyEVgX
FI5NMHfxwD8bKEq8aWoq7tYbRSUg1J0gPGr5tmCXpA8aRGGM63ivNQuspm8RgnTUCl0F3RZMKKAB
TTkAhh7qfkvfxqF5wbn/eh6KGoKYG0dLAGSlcDEjFLlBm6wPLpXgitAd7CNq8ch1OtqYCYPb8CBt
pX53H1rMAR/+9JzRwLs90rVLZe5P6NY8icuvi/WYHyPVvyrUBjREXARV1jMl6s0TFtk0Hmb6Ajkp
swyVoT/JReLaZK2/Dspb6t+Hjiuyvmw2x6NPBhqzm6gAjNOQkEOckuJ4sDMFhbYuaVymbChRUGwg
nVya/Lq1vYhAQnGXAclBzRqOEZ2gC+rwNnAw8X19yqr4sL4c+upWqpNafY9Gb/tPoWeMdAfRPeCC
zrVzIUZNjmS4IQs/8NQtQalMiVgEQsaX+srhXX7Qgggx1TTPPIXSbi2ZfTPMl+ybFt9/FEo5WYm4
KdI8brR5GA5f9wxIyrMt9tvIbD8a2RnFlXoUalHli21DrO/aqgNeyRTRE2cqJNUqUqNMO8JrBEK2
6xUMS1d+UVISS/2X2Uq3C/2BqH7PNgskgmINPPdn1KHSiv/JI1wwSHgAPcNjQByHWosu25alriEU
wE0dh59YfDtrsT8bXVqdcsSCJ8TQ2lX+Bb0zT+2VWs1PlMtx2APdoeUllUwZvq6DDLqMwiMyRHr2
NWbuhVSmDISbQtIoYAhG6T1CUIQZA+OXPxeK7zbqEQlInWy56oYbU7NC16Gu+QYY7LGK1Zb6yQk6
uFaMIy2ENug2Bz/cQPvbLGdcYVRT/IEOhqW8DEkQClHB1aeAps9Duu2wluVu5jeLIEcOPAnyijwi
dvFT95ozNgMtDY8bm0lg9FlYTBAFOjXV7tTY5ly5bJ6mqPf1fs36zuyzWkCknKAR/23RRgYdssHV
L8H2MWScV/ekNLYbVmbCq+vWoureivI2m3ECrD8KLsd9pPoLQ7Wdy9rBToz9j4nM7r7D3hBOtZjn
Le6zFRHK/3P1XoyZJ2Waq6nyCekZ4CZ1sApdzuxj+i0DR+6R8/qRb5wnC+uY0aQIzF5HJqwyPiwR
PIbcxgdkNDMr2qY0OMU2lOmTCkT8qTfcvRL9CqDmvtnMkskZP6QCJoUoU3gKj6rxlLjKWAiBWSKt
c+lDakePEL+jRy3y5PI3qfLjrAwH9YCsp/KNItxg1n4Gj1TxhCJizQa5Xl6RKb5LqJr7VpULwfPy
JgN5YmbFwoAv2qfSwDTz9TAVDZmyPgineEIuik6fkaXFrcchUgvZnUAulkva7i0CnfVWeUuk4LnT
Uu2ulEwgAtLocpbKSlx26sIU1I6ZjNi7rZ2qWUX5WcufZe428oaI5lZrF52ydDI9mtpj1PhT6a3D
ptXAOgcCIrp+1JBTc6UuwXQzInUw/s3+h2kMKYTW+Urjuk+ICRIN9jubf+dBRDsDbMihVFJKzdYr
MpmU/ZVNUvOiwJu+Iz2hax9b6Lhf6xx1c6KXajtgrWgN4XT4BWnOLTBMHDnzY7oo57I/EY3djUE8
ES+xkVhIDRDfwxAE9XRKQU+LrE7pu5s2Z1XO2dkpVMf9GTJFbQ0LcR4ya9/b2dvN1gxDzlAEylW9
ofSnloriFDgbtHh2Zjf1kABHrmQrTlvQ3wsmznANUuDSFiCWkOBD5VwLmnbpw9eVHznk3n0mwVaJ
apNMBJUpg12gINMbcm7EMqnmStwZ/amil9oC/Mm4Hy5e3RaCeLoOGnsk+GHdwntLbuS1uvIAcYSN
MV7oTzsBzWKP4hmOYxC14aLFqPWQs20jwx3R8oSUTv+373LjYXdkVsIOaTba3TpNwnR3H3MJhuAH
2GRzHz3k91f+14EqH5uIiLPDRZXqhc5zq/AFY9EGpF8tcZzTw+RC46MQ4lrNz37zwhuArldhCex6
0Sbr1/Rr1Eyoq2UZs/bLZD0s854061zgOILRYcJoT11nS5LuiRNWzMhdP434tngkpn/w+ieNNrpO
94EZxIbBqroiJIupcjR8wyhywVtaG1VaAZvE1N+WWwx6G5ENW1MJ91iEKawHQWkXr3QPlW/Ni139
Oa2Cx8FO6FoZQv6ePxuW3nkC9XfRznn4alV7yAjEpMwsY8rzRz3aYBb8iLyqNq/9aYqBYXGtxso4
PA/y9EcFpfoRj8QQmnpk22nRLpXxbjGAl8muAFfKyw5bdJOECeLwZQulXpzcEKG08DyIJNW9n7gb
2wvmB7Pkxq0eoNPvIdrUE2xuBw2bc7JGFWef6H4I1vAf2zpbXoG43Dc24bclCDNfrTyZAmJoCBt5
6B8PBst9hNKDmXKcs5Al8BASZgriHsanSrt1zSfi0s85cno0ajwHhI2/oWi7DVnWIksPv5GFaU8s
i1R1odS+XdGucFtcmYcqhOC/MVeUtAktaRiwmL1CX0uH2c7NR+IcEaYwRsBuHk31tz9pJrBk+mYR
45Bg/G0a2AGg4IQZc5iFLGAHMbkTBC/k8Mu1e5opHCCCADWBfeHrbYJDzCS47DaE8lYL80zwnmwI
UBKJr4qk3Lodl3UDCP2ERfoXvs+BrETzE0rNW+Kf2pTa50Q8yXjnVHSicoLjcQX4kDesJoMTIbNK
F/xJrXAvRS7SRuQZs0p+KoXgISm6xcvEjd6IVcZ2zG3WEn6gN64bhpbANWNB1vct1UZFLavz9ogp
q4RU9IAGRlow8hAtiI3X9KzLEGVoj165hlgCw/TaQ4VgGCCvDHv97gM5E9F2HsnofIpw+eI8O6j1
EanDMNxk4NpiYLJEQCc2GTupyMlRCQAhiPzQ04VvMxud3fMz50NqIy96ViEl8eWiScgtiEYOkS+U
/Cm/QOimyDoJUEYgeNUAzNozbwO0wfBEwRX8ZxKADDYjWnUCr0oDxca+96PzH5ZA8bWEtbp2Tof+
BaV5PdVFxaut9/Pj5kANZJRzruwDibJTSsiOi4vJhYAmnwOmCLeJRbb9McJr3mc19ZBWuBjqhkY1
3pAxddBrfB9VhlARyytypHmRZtLwSWzPsFdCclcScFb0ak3ku8nHRkZH084X3E682gsJel5ytKJD
7PEaI4pKD1rl3BImdNd5AD8XQFujtqAWRNR+m6g2OrBznTCiwhXWlSIIPbGXMIwr05hEOhxKP2nc
JgRrbZPEHUcpicB1yJqI5cbNLlV0cKpZyYtV1HQC1OLa+GIvKiLl+vUzEHZN4SBiigndHyYwJ5sA
2g/ZjL1uHntf6v7g6DBYSwDuCksqCbBtVrGys1C2iSOCMCuOTJrlymS6J69w1PgU9Q2gR1pw+4gv
Qrp/gfECvwBIInm5DxmXG5p4zDYQdpkGy3uIrJyDUIHdMY2fVLzNEgDgEbpml3fa13M1tiY0Xb1r
Pyhl0c5WbDHIxxNATHRF7P55wdwbMLbocLigsuhWXPIlo52vPg6yBrykTIae7mcdsRC+oamrO51Q
LbRUvvNx2N8Z2CThhjdSP3kpTuJAZNwjinYcSsFHW6EQBFkj6K18BEHzJ0aFiTqEMOtdIs4NFyzm
tMSiP/SMd4VCwQ5OR62GXhjDSX1bUf5d/I6lcygNtcn6KbigvrbDseeU63C/805OGaqhJjcNEH74
gTKZGxwp7x34CXaqycyz9kif9IMD407mB8O6guEnDl4RCHL8MviJjCk/CXDFcADlWzNw453AApEW
vhbrsAF1DNhogoPuEBbjmUNBoyNvuWOiqszb1WdCKR+WJOqNKYEDAU/0lcXwRkVR3pxhm+SlPkBA
PovUBEqqM64JHA+NqaHFYv8gF6WWcquz5NY7x/msL4c83+KQ8M4KtN1UpGWneZFqUSZPBB4XxFgB
Y1xYLW1WDQ3Q3xUOn42oexocNCF2Xo0AwI061pSu3+5F0KymJoZIhI/9VSWq+V5Hp3SXD5iD20UQ
UQ3bV+W5vrlZHiKwlA/i4/BIQ9DMYSpuV/qDY4ZLzy4WsvQhrFQwq+2m784q9Sn2tSrTY9Cgqmyl
otZuIeuk4JvgN9tgAUPF1sfVQTjK21sQoLm7tXLc3/DiFgXSzOdQDRnGSzILXhuSR8qgxOiegjoI
Oe7LxhAGejc2J8LsboTK8tBzposF6GWDkUyYTqr8BIMsjTCiEv+WxwMJ03qE2nRGlSNH5ukd/E34
UXWIy8eFWmN1JFYV2dVwQcfRK3XQIa4PTat/4ezBXWXEf0MhjKQJ3tk1yizcx5VHr4HOh+vUr7nu
Po94fqfgRCDstqNKRKUdA3AmwDfjMzI6/2e49+pMv+9r67TpDZ5OWCdWkgEHAzZRbQ4wiK5vy27G
kJ2/EN1HK5viiM9cvxSR4shMvLXoXA28C5v0kZmtrxtfmH6YbBCVPWR6m4ImshRRUarHAykMeoKK
bGwCGDOAzxJ2Tmlf75FMexJ4JJLkMB35Yh99WPiaOaMY9SXHr+GTRBiXg0jMsFzmjIDEKI7jWG3O
TBtFQi3LEnOdwj5qgVjC7YjdtFAp+9RDiEUqvxwfQE3FNAuzslTI9f9AD64zatBk97Tvvt4it3pq
H0PiREnVo+vNPMYifBiXS/ZFfC9K54Oh/ZCR/4njsZe76CSnIq17bejODTa5ZuyaWAt950OFOhnB
6I3UnrFzcKto1bTrGlH0qpZlNsxXanuf9Z3Iku1XhaLaM3yBqTuXG5JkeONEYtIhjG+fJpkfRcIE
25U7l0MpN/rb6LmOBvb21EDkOFo0Faa9YTRJPkVmlXQbhWjWt6T9OfFhpspkUAJ9C6rhJFPzVybM
2KxX9/dGdaneoqAMKHdIcJbSA0pHjK4I2myiWCoqlAN/x8IfNAmAnBHjoz0zVU2B2FppGs8Oyy8o
r/VFKUz4FgLXJRr9fAoZQEeRvot1qhfpmmgi3is4JhR8/ImjdRz7LxYqwfdjbCqiPZUugv4+I9rl
zzKsgfFxH4Fhh06k47zLOjFRHfyPPEKgGfXC/2XdcJWbftD1oGvCXtdG8QsDcDkNkRnVO+7vhWVP
Nnf1erkjtVSsbLOr4N5wvWsQ1ik268bZtPLGgxDw6u5tal3PUMopEjuvxgCQZTcghO0gVmy/hvct
yAIGlQAr31C9NzWykLr7fxJ3Bttq6QNyuS1oveJY4UlhXMC5xQe5VbVbHmOZ3mrSXic23igXs+mX
TfFsQ2AYv3eYOFMB6tWKkKVKoq9zS6AEFCwy8visB/ATcW4krxg2XBCWjcGwouwnRfLG2YJlRBzi
yESNhDLG++a+CteTetp1VBlKmYycf14eFQ3eRqtGgePwJQEZaPj5YZC4Ob7PLQaExJBEanLKmCXo
CUV1xEzEnzAlltl1/JRHxKAfOyIBG6DPM8VuvF6MCISpqKTacaaex/fGvCG3Fy+RRUYUyVxq/QUJ
IlTy01aNu/bxwxOGtcFKT9+45A2b1Y15vmqj38Kw2Ba37Kk06OpwVuqgvjsgwjmgrEyFSG4R+FWU
UDDIlDtoeoffWPlU+SqhmeTmUuDY7oDAvEORZKZgXPbny/S4MjT2UhBlNNWiTlBTDj6ltMnS9MV2
OEzu0gqTdsGHHDRcJhFZIxTbA6xkYZQfROzQLEdoKlepHzzRxqOoP+97sPfP14RPRxvWKoDmlmBX
ftTi1w6sJqF28C/4nJiTcA+X4P3eMOo+Ae9UFugjq6GAEO91GPWpNGSAikFuDsJvc+rgb6xo4NdQ
wMKkdljr3l9HzTYzI/NZd+u8Ae2uYopSyxNG21qO012wxgm1Pr3SELoH2fAis+mydDOS4BXzGjR5
1m8OazigE/YmDLcXSqp1U+DIo44n0aQf4MFmsjjonI7D3jhjxKCA2pnmqAEwHpievqT5cwMRQ2CS
hHULnrcWnq6cxqv3/az5xSsaTL/DQako63Ge65M4tFobL+dRIwuhO134L33+vP7FrIy5ZA2LYC8U
fyOOM9dJ7y6nO57oNdsVu2oGJ7c8cFp9H/C9283uef/CT2y09vtxbKEw6L3rWYpnanZThMd2D9US
ijZAUtqxHirqK9b2t8ny8zQV12HYORHoIF5g3Vv3ZgbPbWc3SW/aNoTYXbX/DpsWweI7KsbZt+U0
N3+/W3lZfX105Q0pGnW2OHn4dJ9Oe0XGxmTiKPca4f6ECR8TI7MpnZV2S3tZ6PG6k+wn+YPdXfG7
zEY0x/CehQk7KR1E0giYlvIg0JwnAM86+drWyoEfPkGo05QQjBrMIlLsqtxIOLk3PRDR63YqlDGU
hTzcq+nRM3EiqFfZINj8qmZJ/XiwOKCynIFX87bGFvj4axQyePeN3v7qkLClskrRCpoXU3HM1vtg
rGCsWIMBsPxnMqO+iK35exKQjnbFeHysWGXShgl9ZtAFTT7j93ZoTdbP3eQO4K8UTFhIHXqxqNXK
Jt5BrvsmRwshV1ZE3jBa4/d3Q+EDZslcyYJ4SRIMWRnVKF4H5ncBjjCDUC2TX9b2fPhiYwpiLnhe
XJR9JrXDhATACmq9DDO6y0uhiC6DQ9qnUi86GMrNlbJAVM99SgOpwqGsKxq3nqXBE0M7eKG/k5fn
ewK+xW44JLWrJ4na1E/2iTYXHN3iCK8Cxwpm+OmmK61fSYXcC8xfGw8s7zaZoFT/ocT0MBrlj9KZ
ztwy6K4bQpGHieHTClxfqgCbHZDiACb9K4O0O0gHgiXTraUv7nwunl9CZB3RrgyAM+GK6e/zUIcO
q3hJ3dcM8oQEbVHzpMbYi0AuqUCGx5dQpF6SIJMVbLbstEkUrVHeHulw7ApT+j0EDV9YOCIrMoER
F4J1DjCPE/6iEvqEPbThqw2Sju/3XnWEIBUOY9ePvR8EoqGcn6gfwEAzXvMXJFQzsOdpe8noRolJ
paRZRDYNSYFYYoGdKfdsVnxA+f9jLc8TSwb/nbSosIVt3xoZfA0WskD8Esx+GpbzuxCbmZN03esh
miPdLks3d5O3easvKsJLL+axxAQ+qtFDFeWCy7LfOZOhpEDUkyrDkvC6Vn2BzehLS2+bvbWlUcq7
35Sfk72Ld/6m313HhBpUoyA3JkDqWVr+1V+yn5wYH/MFy6SnvZwSM2QmNb5+UI1G8Mg3YiGwVasA
lFxrHEicLOd7WhxDcLKoeTMoqwXtl6By8QiMWwnX2YuRfUr/AS+eyis6xC0ZzNYQsyQkA+jxQQHj
WI2LFARGCNK20mwhw+V6iMOFz15LdXlVXbRLoI40+LzWAWXVcInGrARYFk6bzosvvOnaHKBgUu5l
xI2+WM00/F0N34i8WDdZDPuZnQUQXJAxI4qMxtFW85yPWBDDTlCNCHKeAEATzFu8RuJlZtYqQeVF
pHxZ7ulLXBInyx6PaQ180Q6RWXv7zx5rkrmXBZdwKzxpNe1jFUaGo1n+g9SxcbtC8XIahYluCtVP
snYFH0qB+qpeJxq/dlM27RkIPslf2f/OJDmc0MJqCWFv8xgLew7hgrJIOpKFnJxx5tSLfJUoOPpv
Xf9ZsRsQJXHijt4jv7ALZrWCON2M2hj70C/VqlUxNHVImn9ro+sv6boABwOu623wWQpYj1uOulIE
nV4OivYXhqp5co5wVnHFbEUX0SpJSnt/2Hf3qRml6X9xqTtvt3XGdkoKOpqTB8lW9YzuYE8JwciP
MN03kSWglW5VLh+mAfVlFShS7LU/atSyahpchef6RP+x5BbdEh5EyDCnZHMLYltfkihna/YgoHly
ptzGWT5Ey4+kpZWPcQpzr9VJP32ECcK/ifr3lzihk2BPmEkWwQGDUbB8tL2JxeDICRG4O2rviWl8
oiaiNlnmz7C+HAXzMiXrGV8IeEdUtEDm1hum0g8ETaBw14LzvuasHcbWEhfbX+HyPZCH6U/LB9qo
HGBsHnHpFgrrPw3CrgnsuuWCOxhpWbCMXU/XvxFgActSg0CeHJbRFJtTXYXmJ+XH9MgMdeJyeQ/m
NlUS5o4msG13Gv4p9/VeXbgTIa5lqiJWlXihtPATGEuFa2yPar2UciBCh1cI+wsPCUpyeQ/SdFMF
7A0bxq3Aq0dZoC8JAC+ACtxfac4gKPpvobA+i7hkaJDsJ/mu9tug26nQKI19Zwo0RY8BOltyTyvO
m7IFEHXJF4QSsEyCraIRvO+KMaPlK8CHFKhC+AQWpc5P4mpdUmLeN/WBoBkAW42oIZ3/pMKJ2pzP
lp8jBab1Ti3kV2mNxf961abe1WjiOddw+OwVpg3QoA/U8KUC50Cfi4a5hAH0BZwdwmLDmdU0TgvW
6uPR20GFa7L+NneT0L5MbCAYqh8Eyo+QRJlZQAD5LbmY90SPaxbqmg7JStk7F5HCVMgY2ALtlabx
4/dxReZkjeIiP9n1eimsTZXRSislNTY+qzYrLc3YHf+mLIBaClgFd2zwsf+PM9XEl/tyjKtNgyQD
9jxsF/ZX1KwPagjRYgDHkXcIa1Gp8Aj0kQ1N48jqM1dD54LZwnCUE+z/ig6dvofNJdreNRWRfLdM
e+0UuPqveLqZmXrP+28ylokVv6AnfCLIE6lEWwCGXbZO6jSdJo+/QMZiO9E7qaq90UDM/go3ueVY
uh4HZ/eI2VPQRqDNTHXwCZJCEL7m+oFcilcjHscCHZrEOuRVA+LoocPWVy4bdszSio8AHoYadCBs
aq7urFKaR6QRtTUjBd2wxMNU1h9rP6E0kU5auBBo+8RlssGAJ57eL4C0pRYhBNbfcpeg86CaVc6W
24Yr2GQ3mORwTrVS7qPfxLscRiGbZyqXEmitHYjhWTnsaatWCqYOPy1uXuQRjnL74HxG/HhGmNqD
CWeyb8ijIsm615Gt8oJkRmd9VKJxi9aiAccJ7Jx91h1X0ptt9hn6Gdjl8gm22smVT8tzsbe9nrCl
JAtbiTGcPG4TwGVBL5YIVHcA/2GwK0raCW3E49ndFpUvL6b2uR5YDMwk2VGYuriT3J0nF0K4Uwrt
Wkz61y47vQMzMKp+lX0HXSvGgyVcILB0L030fd4qhweFBOYjxcOZ/QB3zrKw6Efmh/HL1lz+OfRu
eJB+6hB/7pU2dLIXbInIBZEE/kG6R5POdrnTpDup4UghupwePIzzTM3ZR6Ul9tHEb/9HtZoHQ3fJ
GWzJRHFCVZXoy+shMtkEe+Bw38wce0cWKVhdQOUpE9sqnh7UZXBC5v06pkOqWBOvST2jZrJrG4HN
yWPt4Vxs4bnf6FiD6M+CJmiVMuLDJ7zeBxt2mvDOTKa/qheifh279BUa0+hjOrelUIgoKj63DIo+
ZzWrhXMl3tzQlmxeR7VZFqJUZvwZLz9QIsR2FnQymOBAI4nl+uMc+KWxGI8yIYaTj8sF8RWeXMfR
DjnAdYaVizVyGT16YsjYsadxAbQhPb7OdIrzEFctZ9hBL0yP65pQ+S2DnlSBGFyzLDzYrqF+jDgE
LYA5jqdNCo9hjBvuvTZA8ZU9mfbFVW4xJ2oTPBVmPEyHCoUptpDEWbcsrcwrrQx/YaJwJlDAhSLB
arIxCBDbPRornOUQrOspeiihaqBynHMp13EmtVT+vaXV4uxLyEcKGG02RgKk4ruoikkT4xeJLv69
kcbyn8S4T3T0cR6rCKcq2tsWcaXBfJ57XfURIwmLmG6jzb6cgSpFT5jUZck+iDGN/L9jVrZK7kMD
SD+Cwyov5FBgYW/umkU5wu2e7ukz4YmqGWTUgz9tvgwqqMKCnXvK89UzhwiaI7/DnS70t3YN0sar
XE4OiregeiyGAc23EL5z59C5m8aEuwzZ7B9BiUS0Wp9E/hDcGUFtx+eemOglOlHKehEG1AhGf80L
ZFnuGeR0H91tmFVTKCNhGmTVHMiKqDe1spi1gI28pbG6BjWrnJWQ0FU2H/0R+t1fruxu/ECi/VEV
B3c8t+MrpPZL2RGzZMl2+d69xMYrYzSL7K+eSGmebciATLAxo7Mth6VepnxHcL5z+oLpqnLpNjvk
Uu69mKqxB0ZOFYwy3dTnN+9RWJXb2Z+WxInK09I8XmG6/2/bqu8tyZsU0LQyN6Ebyn+etn1wBJ1y
Ta25aRuMHJKu94187XZeWGsWdAyKewmXUc6OU8MFv8Fquv4skgopPEsS2rtOxhOrdV3Jgt22E9wU
VrpoMnCkWDDgunLDY+Jh+7WLa6NAxBB2VU8SXQQ3QcB0qKjlL70DoP1HRVVniAGzQfU/xmFyvWN9
dTNw+wKczCWWpySPBz/Wl8u7U8jphuKWcKD7OImAAZ/IawDDSQf0ogW97vIS2qN6HDr7kDp6jVEK
JFuiHVjf/iwQBWItETbLZomVI0rraTlxp0Zq6ueqnBvzWa455etZ5JfBDO4N6P3dNl3e7Q8vVJ55
x87mOrAu1JA44o+7OeKjZyBpQrRqcOP/h5eESupLp3oCv+P0X2Wq8/XUyiytrBtyqEywYD8ho3Wq
iJthIaR3E/c8KLJugJWyzlQ7LLJC4lVhWJS36m0iauq6336HwyDU2zUoDWOqfJ5f2DGpaKwnV3oF
yv1TgKANHlR2m63HOgQ/5jUf3rt7w1BcF9jJedwVX5xFI3hZLYG8G5EDiWJtgI0E6EoB7NsuSiXm
Ft01PKM1ie3ObrqvSFzsRMXvWF8XOoBmtBNqnUjjhY3soXPqKRE1FqBXF7Mo6316COQ9T9eWQrge
+UgG3XHkuIodeIawfkjWYgFypY9QwRkCFyyRhatQTPq6JzAPt/IZqw/Z3sGQC9RhK0n/8VmsffVX
+Ht6oSjrV1em6KX4ez/GwglRG6NYduVYrRgjYP8i4mRoqoE//kA8fp6SIPMqvXduWVp82Tks1E4N
j3ObC9F7Q3rDEZeI82EVk2cV4D/FU228Ul9LjnDCYnJLqDzY5jS+rsh2x50PyhGMlMuiOBl9G+fa
23RYuUCL+z/OAaokZEo6nOufo0XIswUiim13wWbL8JvuE0tUEBnxnqgHG2ARlX1x8/Mf9rMduqE0
gmF/3jSGjeDkivp3PEWpKxYSS7WFeGXkiXODhFxY8vWfGQzdy9+9ApvlIFNlIKmOyyav1T27NTxG
76Jl6Y2+D3RQhzMlQCDYbERDVwXrFmpZ/acXE1o9UD9BcXvxPH4rHW1T+tTM5MWWtPCXeKVhMxu3
J+EQ5vKiy5rX0lfZ9FfJ+s+RdTqzFrDaMuSMcwYdQFNnDFpWoIa76qESHcvsUMWDp+eL6YvJDcnp
L/oXvsZXJADAck7fULvY7HyUoXhx+IT4r3A3ZeiLgSvI0NK+VxgMcP7pKCv/KEYUVlsF3K3gCAXo
y3t0LE14OvazON6mgRbq7Tdywf0nrdQ7uJ7r91TbTfT2nrN3h9uven9PFSb8gY9HaVVRXjrDsYhI
Fmoy/WcP4/uSEr9kpZdBHph+VW0UTRoLJ5gS1rEwGekZZuWd/VgOTkBg6LzqOg9eHzS2H3VWA+X8
txhm+NNtPlmL9tFa8C9fZZMaGYv3fDyDzmQnWu6GyOpvbQnoxEdBNIymyMWSZqUJxlvHlkcPnS9O
I0b3tYw+gAtDYAgg0gns1RkI4ECNT5+jHGsAuVspPdiaDGTRVsTYh8FrC6luTKU9p030Ap7wGb50
tYRCUBV7cmxT3H9JBvOi+6CC4Y3p60eIr2FhldaXweDESm4yUi7MIlfIuMtK8gTVLCcYtx9iVmWG
73UMlbETpeyuSnCZxnF39Tv4c5XMjNWtoGbTh/JP77cqSel7Xy6e/bHRGFOw0B6pLQdufqPekvyI
eomJQzLdkTo64bsy5V12+UTi58QMr63wI8iiEv9sWMkN1bli9dv3/Wim3C4pxgdv5OpepdQ7ewGS
Hta7tmsVz8RuERYOBqxxaBW7w1WslrpeMPn4jC/vJTITdYg7ZJfCL++z5wdwMrxRtMgUYl73jjDu
eNbnY6YypjAdFB70Ekf/r3tjysxlmjGOB1YZ5pBDkRYq5htJ21OqeVDMSjdNo1k930HvAHOcE79q
kOwx/KgPwl97Rz5wJbpxVZTVjly3Zo2Tu/S/4scuhWGxsFWCLrNiQJrr8soEdDPOetB0/ZL7RNSd
iqbSHt6Wbr1oLfSD7O9lRFWaw3o0X72Uzl6Sqh9TAU193PS8t8rmaaiqV0YM/V0s3KK9V/CheSCZ
0DrIEPVAQ0Oq6XcWrBU4iTOtF0US59ayTTb9587z0n1uLIA9Cj7FubNiPJrjljfVyuPEMD+8+4Ni
ld7bEIITNqrCnvJNUs8v/64QiKQTthzlHf12AnYLieR6q9Nwczt18ZkdHGjRwADWaeV3Rzs4HP4M
RrAX4wjP/tHkDDvzBX7kAwIZ1ISK7u1uSx3DhDQwq2LX/Sn8AnxE3NwNkpVTCNyrdA1W2fGOY5zL
d9gtH2sh25FaX6RV24P030ndzvcYCeoHDpOwjgflWVJr+5DzxbPz4/HqOW4eYVu0EbsZGYNoOWTd
rtx1DePkyKLG1dhLva4t8bxym0TJDUrINDQ3x8T2yCzyTYl/W6bSZPd4eorRjvYycm9fJa9IDkk7
sFsV/8FupbYWit3WTTvj772TZ1zLmwPqjXbwIcmLZXkLezgBWYbykBR2xoBDBf1aqT4gsgIp+SHd
a1bkuLb7HfwomfuWnt3Ng5q2DxErJNit3EchMQpwngK+YbrEiiiAJr3i3HHT4279HVEnI5JhhV72
ir6KbIF1bq5a7o9JBOfo4iirTCbvoU3Rjr1qlat3cAbCGgO479B210yCrsaP5VdXs8Za9Af6vcWh
Hgroebw6rHDQhpoBSJL19RHYM10uTzEtvSRra8C581ZDhi3bmic9yRVy3S7bbuq07RtMIKTi7b07
YJNihx39dVNE+x1vzKjnWghe9L8HQO9OQCBSCkv10bhoeoxYK+YrX7yQw5msrU8pDyz7JNUEBcwA
H8eHoO6HzSjfJICOCWksPkv9mXm3jzwl5bAR1tQY+11+jDSo8KyzeGUeSyhRt71Y3+YoL5KrOmVq
lO5/YHJlKSOPZk/gjfGQEqz05N6rtoxKkDAYXjFhSlmHzEHPhGN9q+m57SFJsw1cG5li+h/2pTXP
aflB4eFz3I4WceCabAQeI3nFPhbxvV0CAKcXloxcVg17D7afP9500NMZ59K0pWRmQ5YjD81I3xfO
Aiqh9P99fd7zrSxMd6JWmj0mnGU6dB/q2LMmbtb+YqQjRFaIXkiqaUk/gEJY9qezSLIVTvvc9+nT
9Ty86H1H6mNm0D/axZfrcLOCsqNNCtPxCAG5yYD8aNDJzNK6tQKEtv5IGhBat5eLkHTPHGYJ6idM
E2ZMO18U455vlscQwUAyOKrBCqZzQ3AiGl3n0XaucENa3ugipYiW7UYZHp0WCVBbIn1CuUDVZ1ab
IjKBIo7CeeWucTvuOK+bKDujkc1z+3gG1KK62Bx2uuH6nbJrZOx8NSH90im/ggl7TK90fumHjN/o
ecAtQdfRGM6FrAibD58XgVcoitjdK7qw4jLfoQFHwIpFIIrTsNyiswK49P5yE+EDCSHoSPGz9Xyi
LDELe/Bp+Znlv/LxWAxKvvHnvm6oCps8FXDJ8rwxIX4mrexU9epKrN5PkrWBGBvdkUYTpDY2zhms
PAxWzGo/n0OloY0ME0mL71e2VPahmb/TML/otjd3ThrCbzQxyABgtjPHVX+J3IXeoAqofR1rLLcj
xnsLk1kJWMKvlAUQp0jQUjGySiUChsKX018TA8hgJn7asGQePq0ngaREV2TCtB+ZAQfQ1ae1AmRQ
mdl4qPWfLwi7ikxaRjcmmvRY/OSC2PKwQXmmfYNxt+dW9lX91or/X5xr50MjzhKyha1k1m3SIouV
gKML0m0xKj8+ZIvoMXJNV1KvBj20xQ6GpMSl+BU6LzjhoGIIWMO3mQk+Kh4HqGaikAAmPZpSRzrd
TzvzQhPxr1b6cfW6LLjL+K8PvUeXs73ZyqBAOdxToKz9snHcxBgtEoeiIwqYg3hiDKunBoQqQjj+
x/u/uN3FbwKS58jXEtE+w7miD7fqOL2EM2/lRmBZTytJRRAH0ybQw0oVj5Fm/+xp0Y+zSJdHSC9U
a+79CchS1YL4xSf05AnLkJASEEljPKeJYDEGiTWycuGt4Zn8A87jGF6CfN4ir9mNk1qbde2TOyte
h7xiDtBI2YY7xAAGZIhj0m8dWikv5gOcYomx/7ZRLSFPOVonUDH2Hnj4ZGYGieY58LeGYASBMCkp
eB2tJ0T/i+gCEyaH4n7EGgkSi9U9v67Ghp0Khrf8+oIDcbKEw3zSQcImfoGYPaGpMgtBPxFa/2jR
zaralUmqtGfGQaS4RB9pLQLHIxPurqq0XW0hO5Ht5UnXl6PulatWpNivGgi9bpT1hR3EX4Wlhwer
Zjgg9qB2SJpSPCuEJn/2+qgPfNgJNdtTAV99R/HdRzzRZKGfANpjcwPVxZcoo2iYXcxnJI7Yjm9v
rbWvYAEeLd6iauypLW9QY7B3KzvJ3vF8fWitO0+XIWas5Kuu5FuSOtBgqkg28/o0kuL/GA4zkfUh
z4cQqHfS+ZFZJ5i1VFsqgc8xpB0JPmkU2YXdZxvAa/W+BmuE8Y7SBdp0cXlHwhpgY+J4qepm0v3M
BylG3gjdmxGwgt+GMHTjXZbQa8+p8yP+jYFfQrF4QfVylLulgg+b4fhLS8llR1m6lzJ6Uraup8IV
XkkdsUgdTo+ozIQ45UwrIc1AfedU/GjXJNZi/PA/3+J83yyWudTPYtuqOF82Mo0VvKhgt4hspKSX
U21sKitU+nFN1tnSX7g/CNkis89XitaHEJtwQosbux+xrYVPr/W9C0/TRPyiF6hiF09SOBvo8KcP
WW8KCMPB8ksLLY9A9LCRZgb4+wV5l350kbSxTDfGF/h1V6raqoLUZ8ITUe5Hn8HGQu2sKM4M7lw7
KK+tKC7QxEiknGSjGhzrVeMs5q5SI1V00ND42VOTy03v1YngcgvaJl1of63JHm6NfsIJCYpAwmFA
wgR+EMSWV/eYcbGo+kcUU2gNi5joXyqEEl9PrQOjYBl6qMv5EmBB7wBDhpXTc57jUkxfQ+81Lo5F
4MUfMT0sORVQmtIbTFOBliPFYkWJJM0IsLCcm63CBFAlQJco6ityHW/FIxkcJ6aI9Fe4Whfx8LzR
s30oM8sqiEYa4YfS/HgzDf7tmdkj1FLfC1LTBXnCBFGLrHYBRoKpN9OU+Cyr9BKl+TltshTjYP2s
VYovKn1b+Rrp/iThrgtXgnjyMXJj8TuMef7CJYK/du5VBgQ0J2IPFDlR7iwgl40pRja0XuCj6Pi1
2OFCDnRy8gU8H06U43DVj90mJTV3v9xnwHwLGu0JiY53yBBV3noWoeXHF49j4RH8krFMGhP1sefJ
Jvg0wCeWJWId60YfkHB/GrMfjxOGODD4eskDoQhkZwlyn/CICFQqgq9Io0053ws/xai7/Ehq6GpW
WSk4DhycyLe6RZSOZySQRfJuXH+CdHjXPhQuUGex5g+0KS/VAd0+5ktq8xqxtBEPDdE0t8QkfaVj
Q0hB0w+GZsNJys4qStNxTRBEp8ckp9l0tE5rKQK83AI/oEsFxGUvfml0zvBLjrvZGkahw196ckO5
nXhHwN+hO8slAFWnAV2U+BR5uGva+2p2KZWWRrjsbWBn7KHwY8aQrXyODz/r3lZXETDkknwDTqNr
YW+uQGea+wRmtGrDxrKJz924udCEjR6BNQQZXGdolLkfvoLNbsS/8juwBk/yHvsrKlCReeMvBxRX
dI73W/duAOyCEzYElTBeYyLf3D8FmDBTYwNvkilsqJe/wk1O7sIiM26C4vVP8YrfW6AcPP4ZRBXo
aaToLUZs6D1tweHUmkAPZC5ljY8vznPFP9TyYvgKpIGgeb6Fy0ICDurphOs9lhvUH3B281/C/htR
38txkDWWvzuACWVVSyvl0MlZt+4/WjW6OdgebIzZxlKY0K1/ek+hFwVKqx3gOYSukDhox8xKc1Gj
pbYGG7iQWywpa8Z6EEde3NSqsVpy0DU51COlT6kKPFoVp0wcluFY5nlobrFw5JMRbT/7DdBQ5y5V
H5EyTjCJikUVCUt4VHwxBlK9n0dQqeWC++GKzoYAtUFhLOlx1M0WO+vY6KxaDgqXyNC66ZAlTVS9
X16lnvuykFBEDcroDGgc+pYbzfGLy8FiebPjZ+z0utiv1uwIg+TtmwdKuJMeWLBEedayZDB9f4xm
zJm8fIVdPeRBMReD5CH1oUPYwc1rCkEoAkT8rcITRgOcli7JgxVz6AczlDBxMmZwfbohpd88lqgg
vaC0g40j8wQVwtnAYPvmjVrfFBHaJFE8nWJQAFCZQt77DXAiNkrV9lIGBAU9rni9GG+Ysd7mm35z
ZeQqE54X1psZra0krlVzNaR/1RoXVU+ZwOcXDFQCfzaLw72+cFLYU602ckB27avwJ5FMQMXv3x4n
4bafKcGK40XN+tdTPoFi6U9syvSwIhRS6uzQvm/USF8k0DShdQ+H+9F+9w8i90hFkkxejI4jlj4U
okPhgSXmj6YoZJ0+LPn7WllM7X2qmGfNAty+juPBaM8PN7i7ZNzlPYVh/EKKuomgg/lbtncUCEqp
RyUvRw915JXu0Ddpp4o5Twp/CkKNjE+jnxafnW0OYFnWiLalcrOqEcIu5aj526SybMeNcOrggbuq
ia1tBy6OEww9wrBaZu/P/I41KxMdsnkBHY1+VWk1uQ6fLky8PwadAq+RV7FWOCTfvESVT6nJR9hX
V+6Lq5NnFh9os9uFcjmqVaCVXxh6HPHYZukzx6SgdvUoBNl78hS5J2qws5kHV8iE0u8wdVbWPs7q
aEAs+KlcLcM3u2eg+/VyPRitHpMO+ZNqNs/EzbZOoZZYfU+Cl0rUgcYxn5+oWTARE/iLCARlve3u
rVAHPWDtwipcLtdsolM85+q9Z6RjyDlzKevtT90ZTcuLm04IfQ2Iggh6SQFqDluodnWcdA6ncTS/
3KVpXFXqjF7JhtVMoyC1CLBZdcyRyIUah4AhK6F8IP/81ir8Zf9qLk3GABZD5wCxs9ST+ZxY7xdN
/JlZm48AAV45yymnFkyJwYGMe885rwVLnt2ZfYC6Q2SKawfuVb/FrF6jdXffcNS/ty/xmfRsfpKX
mIVfNjhW1D3qt94cOjymmj8ilegNUFZZQQUe+gs1hetzs0k7xEOoDuYeXQF/HSQ2Difvel38yYX9
hjTON5n+7AzuXPmS1ED6ACShkjKVCAGjPKM95NjC5w2cJwegDMd0uOhtmv+1brcZsFNrpmaWruib
lDNCPaTrvcvwFJmUGdsX6xQ3mHDvWzR+k/T8N+cP5R3fJaUkWaJeHTQ9UpRx3PABiQ/VtmHQr/yY
KNqtuRzdjVxnTibRfe+0gsCpi+xLHzPraw+XsQlcC5VjLfMsb2XVqIndaJY19KLkYqBMp+eNCZgs
p7+6oGOuJdkp2dmR6I2eeDZAC8FcW5hOO5Fg9tGSNGgLYPK6HDd/QM7qufw7mzIYgT4G8UsUlkqE
SyRSzevUU/l0A7zN1Oj9TvVU8QkClna/NQC4UGI8Hvi9h8DSep5pVz4O2Mimowyp8XmJp64Cdx76
moddWEdwpLSaeRnMI1cb0VrrbDoIT8AKKUyajk2LiY6k4n5BU/0TJqDuI+2C+3Bd94E7d1lnHd6H
7HZU5z2cyNNzAQjk3IE3ndfm10BRvzDXKNGF818aUqHh11fjFE0XMZCMyKWv1vHYLnngJzdNOleq
DEMLlV6qAINS4FZlZ3yizcJL7oQQ+AhU3vE5qKZZ6QTLYNuxjKeYffm/F+OM7OxfmP7xXRW6OWGe
fKKhCbxqqFWCMy7PKpYYUEzdqfoWorygXap6ltfb0dVz5NDYE9rmdOOmuHqHQVTyNLBOxQ05L7O0
3liUE+MYa3mnvYVvtwS3VNTr7dgKJbnXIjuwfbGsMifMN1ZmtjysVeWv8s6ZbdLP2hz/vmtS3VKd
+/t1eoUUzBMPQPzl1NDJxKvT0X83a4WcqXGdj0EPaqO/23N3LdVkHmZtDZr3n3pYAxhtCsjwZ0HE
zy/ZOHHp4goUClHKnm2hCJc5q6bwOPrvELqSq3JD9hUw+bM4pO5BD6tABLuAjSZVjtaO5jGJFjx7
FuWULWnATkpaK3nK+ZqYXwnNIUprQQTjyALLSAnoYdmY7gAhobbu8vRe7L8zZ5VngpSvRkIJPQGD
Mj6lgsHQIvgKSMKeZEwtOJtEMq7kW8bFUscemSArD1hqY5F6jRnCfbpxUjjGH/05i2BGZjPNa+jP
AU6ouToWt26LwqsVU+anZZUPCpucw9sXmf+9qpFgu1mbHw2YHv01Cr2mP37RCSuLCMa2V4LRTh4S
T8FmCy5KUQ8r+bhkcdkdMl3Z/QXA/OadJyr9JORRkKp0XRjMi4vRxm7IosHzdvyXCUEp8kVRyUPZ
zo3QLVZLC9eAyuTSrd9whL2FAJNSeaFfR0dCNEdr4Lebc3io8je4qVc+q1cXukE6PxiutI1Qjci7
2SMsJ2MvIz7S7rJf68b43qKIagQcD5S9UXOKbi2/V9gtHxMgGpmzxkBOIJxp9tSpxjKXKPVW9XVj
3YMnGJq9ohq/SWZVUSSnC7cRJGFmMpUY/aZnm+hc3aHJGkDJDfoBDnfKgv/TZwH+WB/HyFMTyh5r
ZIYlMJxNisTnFlTUT+dbQLRXyIxzKgipIJ3OnVO93Oq6lVo17MFqdFstkrpGWH4JP5qauIhszBlr
iSR8HpXFvCpOSm8pHJzU4ZD90mnGdcSLioQsMpYYupMbykSs3GIczXtClE2PkPrCZ5fCe84w3mMR
BW/Mz4/NAL4HBNMgI0k2Rw9c7TDPebN4gSuywyEfjnHQzWfZup8pEylwvyb9s6Rg2NBlSSx4Qgen
NjURe2k9dtZyFTa9PMTNjZ7ecO9akJRyubUIEioMpsdun4LXIFlEpmRK1t8D+DcQ0wvAaUu34TVL
gJ6ftFzv5h/U3KRMINpnTAg0+Rrhb2llGAAHjDRqw0K+EJypIFTW8oBbJyDZX7PwLovPAk4yTk2s
4o3o6UWUmfLpdJQRj8eo6aQLhFOC2LlTFUaSYpce+iY+2WnBZfmwgao3naO2p6fGVvscvWLhZKr9
TLFZlGWy4Jk7SCqSb/ivD6P5CDtiA2cDeCw9amiRpk94vREV6XQOXY+ECzfP5KCmLTly8bvSPKy4
C8X83G/wGEInAh+DSgjy5rgk+tjnR7j68p1LfD9x4TSz7Z2Dg1lhy4Kp/XrY0hLJa/F+zEBlAGB+
uE4itP6UELvHbsTGR73pKllXR0D6YodDv02eUs1ZxJhq3GfVbyq5yqo7foHDSSCVOdsPVSvbT2/Y
aFAXyjsJ3HEwYkjxW1+xC3yE3qyIhe+DwWULMgo0FQZxzsHQlAh/qWaMnZmYVe5ivsNnJm8BQ0lL
H0bd70TBmkAC+UGst+0JdnOjsUPyKRI53W8t4AKl/BpAt6nXubZLy+iFq4s5pQCwRU4jc43ay0C8
B470PA6+8cvbtA7o7DORuHkqYrJDuLrueyrSDMJX0WM/f8F0UgWV1pNyTpkp4kaHzpSpUEmEv6kd
NkdnB+3jlZBfKZ8JO+jJPw404YTQpdurWj/WKRo10W9qdsf6WV/VvmwzyAh/9l4THh2qLN3a/NKW
8Uxr+5TAmW0lNVLIcvEnDwRf3zdqSBpvk6zDc/mkuEU8jjKmobYCwKiX18Sa0Lltv35wb2Kv+sqw
hBO5qlBUvhoQhEQO5AnvR9eNT+7SV/uNMKyYPS7OUwOIK3x5GKt83fLUQkNptooOKUy42C1iwQu1
oeXOzCUeohN9jO8OFmcmqdNPzDNDW99tvROvMkAsc58ArHRUBK0UOZbrHVzGGaYyEsfZiLuQjJhi
G2NU3AC1yDk6JU5M+y7OeQraMa0gavtqOcaOqvDKBeXLGMerJRWJa+l15rXl3Qy7cIafYNvTCLL5
ZHK/qsomRWzfJgX2Jz8KfHFmH78qlWEsCCULhBHhf4rcmWjTohCzNm/dbeaLyMUcPtleitl7aUGQ
oblVwuRI8lxVz6zHhAbtjVhh5Hq21VENZrNbmaZKtzJzuLJelgtXbsgcnl7q1WJ1RNGZWxHQG2TH
uxrMd/EzJF93/reu4CmES3ORTmleUK1Bfs16X6jCxfDZymW4e0uD0p3UKMQWMmu0PJTv8tUnLUlV
hwm2DcWlYt59ZRhkI301hDEoR75M6p6trF6IBG8PPi3ZWGSdXCeLzv31F1BvXkLCdg//GNLUPzbd
01ybuU8IGbRxiRB+ed3u9A0nTQV3uxq/o8vT4dG8kJK9ylEsfbhaFcGU/faWzBtlPTciuXNB3eM6
gMnCWkJN+/xSG1jZaFp9AIj0Cccq+sc1WoARu70uVp7adADcevIjo7XNl+qmtkli57q3Q6X/ho01
3blRouQ7NTDq6/6TfYsIIj21Sq7g/6eV4BvbbQu06cOcYBoyNGuS0jkdWCljam6JyI2PllrQ73Qv
UjQL4eHYv66m20Z4HYJwkfB805ZzMmmrYKN56ZdFBtCvWp4z4fv50TtleGo0gKBdQafwq+SSwmMv
rzT4zOljE9sduZbhOUEo70vRDHQUZceFLgPQOqBHXHZplqtOf2ktEJ6UidgKPK1j5mGIf1FPLdtD
h62AFQKMZVr9xaf+K0fsEKpJqeL59xBnaKlRn0lrznm7uw8HZlLS2Q71+APKKX5HogV0DrIkuaKH
NFEd7ci9/Ybmxi7TPDFEz8lU6Os+mT8xctzau4PXjHo1ZSXhlmLd1h5ITKkrx8fHd8l8GehXEyuf
H7MT9RtIHeEbvhuEg5dF3DeFZjry7bRqf06SZpUybywAEZMN+AGPNm/bWQmRhw5tYfcQhXeOJFLM
16oeLzI0fu69h+51BIIOEClzR1ZPZ+GnD/N60BFclJv3+L9BGNhchpDtqQik5bgxi/v297pln2wB
WKHec1QP0xI/iE/5zwf9PPHwKGrXZ1bsnrE3N+rX8E97EA+qlD0rg8szh85oCYncKFwxz9Knh9Uz
Y74yXW5xbtBZWzRJLHAT2Dwq9PBzfa4G5sDUrtPV0DrkbNDB/PehZLqZy17tfTz51pjvizq28z7C
xSYFBSv5tmf1YdCRjblHD7plbPen3IkPCggvgP8BR82UDFooXLA7qIzUkpeXWDXdZaiiJOXjZNgE
dJmLeQDl0TnoNx1ZaGcEYsbGU18kreGv9Lp4sI7DSp8ZYRDW50WLFkgndJCG4iv3uL9FV+lDefC4
TSewX79w9PAxYIk3RGOk+w62Y7J7EicC9IzzOOzu6YbZdoxDaGcYYYntCmAZFe35i9t4tTtPAi/a
omg4YC8R1P643PJkcA6M9vehG5c5FDUlRoM/v3Z2b5HU4jRjY06uQFn9So1+gZd5h8hlH/J+T331
0Om9UHRlwyhQhaSbcRYUTz8nf/K4+97rKnObZ2cRhNbnxvZ+1Y51DuMy8YwBPZy7m4KlFHpkdSNx
Z2C/uY+6K3hr7zBcujtEF65K7CLoa2J4OmkV7To1+LRCCPk7mMFyssdAY82wJsAQOD5pdu/0+Gvr
BkhdoUOKFPrIzUb1YEWfru/BnEaiueIey9Afpzr6Tw/I40ZONHcV/ESjmNsSWKVZ7MYhSoJUaD7O
kCS/Q6ciR4RL97Ad39J3tOBI+xazFdW9STwTfbzupaDodGAEohJBf8yDfP/LVqoogo5xvXHs09pJ
z7l5LY0xUW0WsKHoB+8VEvvuCj1cNFz/BZVEiax4zR5WLdE5DrfssepFN+phRPbNkBxTBv0lQ0Ro
Qwb7w/Qlhr8sZ5NxMSmBToqdx/MABkjW5xQNUAIExq/gZltDNT0z9c908LwK38nXK+fcMYRTeWVQ
CxiPk/JjkvMtZHMCsxctPM0Egxa4HDnzvK3Ce0rrYjVJqGkBSsL+y5ae0WKo84E+y7nFh+BzTBb3
HvNh0rojs7RyGiYzu1rnw3gh4DcYBjElwUb/B10ES3kwKEpVLakCTalTpnT+qM9XFR60m3cHIlp9
HX731nqxg+I4Vfj1G5mk3bx623+gm75CQEuRHSRloPtfOC9sckQB43R93lM85YoeBrgwfF8l1vFC
SdaMHN41HWHGX9EjVxRrEWZQTIAybvXCUpdZUVNwTBjTdlKRnXuZSQ9ySPUu0AKLFOnQOz/1lQIp
LJKx+LMFxSNH98so5X+FdjnngPXPubN0Xt8gT28VeiZHjJwNwZuODahzzCy6DAW+D+5ttI2dk8I/
QLXqohAMK0haTVS+9VXJn7+Brny2X93wZkC4G0PfGE78lsDl5b13Oo99G2jqcsN+sB3ggacV1K3C
I5VlD3243qGjV4RJltxo8ELhyNNepPMKgbdET4cI3iybPE17ZFgRMWgJ9uDv5nq5lxkDfPlx0YGY
Z3ZumwpJAndLvrjIOGS6YheqpLRxNkKgcYhmhccroYFrklISmgNKX0Fu2uDsK+ddS4OKJ9XWM9RG
InjISzvPN16EFMRQgYrrec4g68IZhpJ+RdpPtrsuOB89XrrhS6QnRnHF9AlTfXY0giwbo6fhkZ+K
1FbQ7HGe5PV9nhP+6JtvOvBmnCq1mIm2l9+6HwJq/z0TQuROlgUVyASTT9FOcnTpiPu71SMbUquA
+xBL3RbXe+HGfllWuii458tXl6jFQnjfTPXiHGtxw1fSn/YhjUvVSDlofvIEjMF+1v3b4A6cQntV
wltEuAjvwGIoU6hmLXAYsSAhIAhrNpysMk8xH+3AMarBP0c+WiiyHYE0mMXi0joIeFyJ/ID/YqDq
dBVmJMWqRhHp/3IcAMRtkshGDePYPyBqXOkxFiBbPGDF24NDqlPlHSyApPVMzEvL/XMwprPyjooV
LygcOJnNk9bBhqJGksFqAfFIiDrZ/ikOnVAv2H2hQ9PXCDaLe7Bcj4jLvFrgl+XaOx5fpCh3bUhh
jYnnuLtXMamNWcwmrXTgWdpYNxx3k4XSXzc9gAsIgy0Rjk+vSLajMBJU12oc22xOBNdWJmHm4vUh
YYjJ6oJQD8mD6jgFCCow1eQ/QeDnXjqSA6eGqewK0zW/uLNe55tkb50XKC8m8ejxbwmynwmaTJlV
CZgrZPq14HjnJrY5l+Pj2lcOT8sjQ3KrpJl8MVBJ8AfBjuwY3bV0PDKi0wDb63Vi2Tyi5+MsR5wM
ENjCf1OYSTavgv0YAhRS9rCRD5++CEdEAmNT7RAj5GVu7bFE+YqnOKQDD0sJAWCYOL/Zbs6YEkD2
bu3fXt0UVM8e5hcUqd7Ff4RyEJhH+Jj5YLoBGxq78eWeFSCfUPdRJ6CqR8L24sf3FV4oiM/nEVQf
6mom1C63lEzKgvX+FPC0UiVZu1U7kUwFWczQjssEoGp89Q62QvBOHgGZU4hsj6tzKmmNK+eP4p74
hqPSxZEqS0QpD9Bj3CKTt/JOeH1p0BPnGvpF8goKoGSWH+WgNpUKIUfCvGtawL3vMjIA5wn9CdTy
bFJ6MieuTSu383Zuj5UTi9ZxxGYiE5PrFf5r8wo7ijpy4YNkgrg1WTqQUwcHG2pKRT68eUEf00Gd
Yq18X5sygnZIkmVkroOnVrKIVUoeti3lvGA1BR3tFg8/aATrpBeoDY2W1mwHnNIn09JKFkqs6K+9
pIC89bQ/7DMeq5J+Yj9MklQRtQVE+XHTz2v3iyinoihEnhPZ8Nwng8LccRIkMY5w2FhancgDPv5Q
Sam3kfi/2jPz9p34qnN1UrQ3pNKevl3BPP/NMnLoov4NQNnjXhZbVQ6Ixnpwm4MKs0akKmudKcfE
yziSQk8myc30sBmrPEFlO/wAumw146pDCMK3aA77KXSwipIGN9IUG5okNQEauaymHnIbmMEg4FQK
X+8U9uEgLg85/JQHq/xWbk8dlbqcu/RH7NqOWkImBydGUxdFAb9In6LDtWz8zm0UUtYdnpCh/cB4
2yj8UmZxYjsZ2qFTkJmkRksjK85qDjWhu39jbFCLyByX7S0DsHooz6DqwkGm7Da7OBm9h+/xUxb7
9s+1VwrQbLqA1s19o8xg7q6uKMZkUBJy3kDGOAloRBGyAUG7rCSn3aUrtApm6ZCIJ5eUfPerln9H
N3PXgIXPSVmv3xckrRqM57GphK4IknDTRwbdliLwpz2MPr+0hnIZ2zJoeMMQK4L7fwl3H62WVEXT
kJ1gK/e0q8WQCH1BUOg5KMLiLRSkziKHBq1UdfsS76RPl49pDW2a1KpK+HbIr9thgbQ74RqTBFrd
0jDYTNBDGwGRLqC0yUh0382KCc4nFD5dta+SOUbXodaB/NLBw5I/MkP8wR036qqk15KyeKXUrmZb
mk6nM7sVoyINsSgXOqMe1WuR5AKIhuksVJnj4ei6h44gJLUJsTI+ZUjVGkZVY04OyASQhXxTSt1T
zgicnHL1UOfqORpvbxJ5CQmaxeu1WKGYGezSN/D5Pg/IbgwViqBinNB5BaGKXDKdfdAn+PMJLX7B
gFaSKdMi0+xu3btnJSoC9JQ5zujD0poPFwV50Dtx+XRW5JQLj+Z3qjESV9RXa+K4eHHJwKiozUpC
uZ68VZnG/RTwocvFkk2qHtDIc6Zvsmp9fE7wYwa0An//gXoj4lnUih7ltLrDnqajklR6a4Dx/VmV
34NpFGAwu2XYLvgehvua+ymiyEXVk5GDDHAGz+5V5u+YG/G7xJ4bSQ3JXCP4vYCdricHkUGe2Kwm
v+o7SpBv8PL5J8Zwxy1sFzixWGqWLwuuKECfBXnZxgsL9+9zG4xmieCccUJuLtb6UAgK7VCbYQBj
j1E7zoR/rKuMsx4eF4U24r7Jc05m7zUSwo9WpeFvbCgrULE0bCEJIELhOD7YLzWctBLIutgad4Nv
p2RM9qo0JiIh+9xMUkE3+Jj+Ad5FqmZxwRdw0h6n6kercRrZAcAV0MlEsJhu5YHPsVW1nW64UiqJ
M7ZUdTcAg+Rk1wRtkx61jx7ipRgN/+MRi4mJSoTOUMjCvVVQ4zc4OD2x3jXs7ir+MG0+C4BFShDz
b40fIKgZNwoLwWwlQLhc797QIbE3ZJsvo/lqmEiu8ukk8TMZhOPdGHqryY6Gou2LW7ohw/944YrC
jAsUMkXySnQQlIMBCCdP8VPuMn/0F6Y+1znNf4Opz+B2ejHybFOeRfwBw9K7qndGf0sf01KhxJwg
uQqd/mhQQVHyK+gQRphro+aWIvOM7NmKR678Tbzn8BbJAm7b2TZ1dwUGlel64/Lx06DwtTF9+rfy
lFyeU1lDfNhQ/A4WlZGZP5dTvKjOlHVF1rbVn4j9t1lQJgLJWkgOejLKduzkmZCq9/eHod0aWVYT
Pwb82I/YdrnvS9C0ZCWZRsDAthS2/n4uw/gRqwcmn7RmydM2jssQ07ZHaKKp8udVFN8tmgLUdaWA
R+SZrRTq9/0hfBMERqe0dzncCUdvIl6F7SaSgefp1CngkGX2rNmXvbNO73zso9YG1rtyuLSkPvwY
lpQWOQdK9454llo7B6CGnX4ViBSYeQqDSmTVViD+hhkiY232STMiHfs/H2nmvmHLnwGt7FWWv3tJ
I+Ioj35R5fofyHtp+oZYRPrlZvJmJQh4AVKBFxIP0DbPQyk4Lu4p1zIErRyp3dQGuAmybgxPY1Xb
qHAJr7hhXa82AX5pv1brStHoxt09ENBiMRXDMvYFmA10OvEoErcz5loU900Ok9dK9jzLucFh/nFp
BE3oOXovfKxIe3byABWig+yaXjD2KvNqXJWbD/Pt89IV6bhL1iwf/pU7C9arjAXYc5yx3G+IFT/U
/lhnWzIJGo6GPfMVvHLO/pLAQDfz4ggRgqhiXIumHBLlWuu/CFU4FcOAQFNRjtUwG/ag9beQHz3/
OxvaRKG/8LkmmV9SN4WDycRlhEmv2Fmyl8ZjZ9bYyrrgEp0S75rQJpnwoGOmYU5MfRiksgxk/SDx
Jcf8QIUppdT/X4efBglHCufnVllgcfOBYfVp1viiguWTu9Faauv+tO3BmP5M5ilY1aflhuw4VrQ6
RqSc+hG6NrL14WqaTbAW1AlwyH5l2tI2aMnHMmvg9ZMUQtIy9j1DC9MDjA0O30nk9nhrSwOM/x+h
8pzrOp3BsZvRD9O9f89DppODZjSvz4iHaHrvwgoJxlaWoQGA5r+Kih+hzOM2A4Tcvq+d9vu68RUN
LZPbk1naCEOwkABVao+dfDfqATxE+3WKKBzFe+XpNEEMnHd2OHK68fOdN94XMNfmvdjleoYX9xME
LJZXYzgH8iB/lVpBV/z3mL3nwWK3EqrAB55R+G5eUQXcmN/o/3OtEi67L9F1WjvEGEqpm6s/jPL0
50MZJvehgC91KC8s02YA6xgla+QOt4DN8KhS07+vKv9ktEDM0dScdwiJTeE1tk7rmpTWnY8YMPft
jNgsxFfnbUBi2Qldab50VbmcUEnkuufzz81jBNEw6YZlSdEnTBw0IvW75kK9RBDVA5AoxwB4POk8
qQr6K+0ZhJRarwXwcJdz3k9wPaBbwta6gW2qafGkxb2lFBXfQ/zl/MlUdFCeD6YoOjSI5D3rzvT/
oVoVvYTTN6q0gd+HtDQnbF285HPiTyRS24W2pPW0DmMHVtTNS9ZplmIe/WZDcdpUTrkXPkOPC2Fr
kySnnzLyVuH7R1P5iLIUoRhpaORVvLXVdqh8A9U0Ekx6qsdBlPCKq52EPujdLcdwO9szkYAMD/MC
CaD7R2cQjgem5XJwtvFzp04c1qSxTTcdhTHT81+vvQcmovyoAgwf9nj5ZdBJ00TNYouTzHRwutBt
tEn8auE5KVBRlD0/cn9AqD6q/AKabEGqY7AygiZatg7UUd+TgaXhA9r9LaPpdebcas2G9wXZbO98
UQSZjCSF6GxIoyTJdhDKn8wcv1RPMFULT9WR5yacgzdTMG5Hm57zmI54/Gq5tyK3hmR+vAWHwS9o
friP8x9e/MRsm0C6VISH3QZ66C/PrGzy56Y8MgaPg8Xw1/ZLY70eKx7Lst2vIuCDtpZPPiOXoEVy
KskH3+WnowY8KJ27YXRURRayCzshj9WBgf2bUmxjATxf3pHirWvnChKma9uODR/8JNa+D+0i/jHF
6hteFgiiMmXV1zF8sZxmyZQFptW8F3DD2nGZ/WlADNdTggE9txAOs6ADNsuvEd5eBl5QO3fNHvpb
Xf9Ry+uW+ucp/RPi7RNxwkzqKKwaqH1TyY5uf5dpXrDOiT5zPnzLBLHoAhTQlOpT4JmyKqOqEJ0F
gx1wxYARTKkfOccE4TjBOFOSqaZM8prH4v21we3n7otklUGOAor7BjdS27qWSAN7kLBLsrYy/xjr
Agkyh6O+IPRLKxUklWBE1SCDo71YnAMpgUlEXngEVm0o4FTUlKtoZQjXlQtNT+QrVrap8G7G1pwi
FGJDOKyqwiPavVX37CIgM6f0NC4BuQ2aC34b4SRkiBACkGcSjYKcpIkim8cY0/X8pScQ74Z5qfRo
Bh4EM8xr5CYa/Oz4CD8xEurGYZAsTo/q8ChGe7cNmhH9R5hc19yaGNM9d7sKO+tD5CbgzOO/wGKU
rgff40a8ymkHzFEzPhGjioLyHIy790G0o7K/+MCKkxzwBZ02SA85XGVAnj7fsugI3gWBsNcdUFhr
HwfuBws2My7907M7rVa5Pd3VAYzgksp/sOENpIqK6Rje+CroRfOlG8FkV9kRYULWtgaT2cmggnEj
pu1UVN/xWDKrp0clMu+HJUmFQgdAlBklk/xA9z19cPx3HbTrJGJxz6WrknUzIwbjmQs+8eZ8ku2P
821pwZx9IbN1cicvg1fcK5+0yVfCZqPr2F8gxZij5WlF/SwpQooT9MHupoxMbhb2mPggBmPALswW
NB2GI2h/4MO1Dde/47l+oYzVca5sU02kk8upGasj74D8jrHu/Npz3ucgA0C0Oh9vlHCsU0BNB4gW
v0n4gIXbJ6KHoXDmcP5yaR2N6JD1wWPDmcwjXVPzvfnNAZD+1pbLErPY+llg4MfqY2hAORx1521K
BQr8zS5eFOl+B8mtlUXOH5xPMzid97n1mz8XuTCwiuivwOR8ecPhc4JxIST9iZ8OWwyfs/2pdhRb
IsH6kDHGAyiadyrhetly7+IyvlUQvrgYUi7yMLblPHJwivFH2K3sYUCgtS6vIhqmD40eyKp05HGE
kS9ItjcBJbCphE612s7K/yz8JAsHdflL+XEogndlqnHqTEIvv2mEfavxrq6cgW5awUYQ2gGNZN7U
AIYLjsHKkT3slzdszMscnWotyV618N5WGJ/E31xtC2IolJrO1/mq7tuSsIALr+sYeZDV3j0ePeSE
3YlTK5NG0tirBnESWkatx9mTOLRfOsYaiwGZPWC7r0TvgV84cBGepF3JEjTmUSpNOVL6O2aYAKgy
+YPrc/q3b9Mbf08BL3wDm9D1fzIZVPMqyatKi/RIDHbP9n0DZ6EvlTA2GalAuE+qV6+NXwWvuvoU
i+1m0aGyuGAgwFL+MpqAHr14qRI0wdLMh21+rp9avj02YqdK/awMmBb+QjdTJ/z3aHmAutL2L4Cw
p29GNgfB9gi+tVoxZQ04ZQWIyT4DoETWgdV+5GTUQtwOYWT+noxS7Xe6PKCoCVu671HlVsJ1MvFI
eR6d92Nn5IjehKCeRrvh+bcxoSVls60h8N5GjxYebgeTSfAYiT6gRHLELnSN36dRFMAFlGoVczFE
BH+yCrUNpsL8yf57Uvmef3u2+gTUBocigS4qLOW7AMLRyhNK8kthlwO0xRJJaZW9RTchdCbe9MCX
euH1jTyS/yfRSQmLxJF8gDir/qSv5yfhM+KOfEoeDSf/w/k+cOWizCaEzq54hXUq0/6tB8D/2Bjj
qz+qz2YwoaU70FUOqKcwTQBouKMqlKfmxH9hnbNnBfL6mCXfZc3K1dAipF5AU/BExThodE6nokT5
5H9F/NlvghwWDjyB/DbafYfc1LXw0hUV712RVBg2++YGteVzTorFdusOw9TPxES+HZ9BvDKCs7UW
+8vLgpIAa2/J0DiePrXRP931EvSF0EOzbgkfyH5LyU+7TsvKenPH8o6zvFM5BReZrgnbnyerMofu
XAjahyYsKIuJERf3rZa57VhVC5ul4zUuvgs6KiQCE7m/HpwsM4o18wCdvGjDiq8q++S6sIZBDHdr
/1RsSv8vwMynDUzyVOXWPZ8Lar5PjeVoD+LfblVIH2sD9Tgfu+opv2iWF2ag9anoCrjw3+Fgobmy
YXWBg47u5LKn6XVyLYR9blF66ALJ0oDOYemVrgVm3L3GyCD1RxAjmhcExW6YIm0H25uoxJU5l50Q
FHzz9/EbVyLqGrg7YwzA3hhAYgzpxf5lfDVnG8cNOLEQQf6nrrJg/HS5nGAh10Jea4byWRd2s6lA
R8eBig5kfyy1TlLAf8wsmcerVCDX0ZBSEeCyEjotP+F/CdHyyAFlmIlBI19cj2xTyAEU8J5YT0qK
ljXtxCsmMrJG4Krr+kPKnC+pEbVpJqwR6pR6BUXP95nJdcpATYIulIcOJeVlvV9m5bjTHRUdcwuY
OGvWWZA3vkZTeUlekoY8SyGjRx7PZMEpKi3PYEOrNnqOyLm+bK3AXslkjZ/wVVdORlsBn7dAnrVj
nOSSNRJpEcbXmwdYxgfVED8uFg0lEFOUi0zipTWiGETy/r7F3j66i3jBVNdIcBs3uaSxzdOM9tsK
2zFReQiGsQv/sDONpe/0wYEvROiqbi6qnrdAlzgs1OUGKh6U4A0jKJVwZfUrQCG24Ml+Xpl9mPbW
J652mYLNgOo5eMZRFh3mey5qHeUmD/+CcEbJCg8IbdRv0jIHfVWFp2z0Ec+QABII1M2HMAEPc2k6
diMLCPOYSjk7M6xUL/mau4zgiYs8mDcqvf+U0E7xUKX8NQPd2nLrRF+eGx9x9FRqCNx/E30z1eqY
vfgofrwX2ZdbftWjj/Q5ePNndzj/UHjDxNYHj07VRplmq3FsH1qpW9euNGCrQfmrho+rrS4YMy+d
7CEGw5AOiWwfRbV4q3h+OvYnZD35nM6+aBYOLbWjUwtEM8mfcEha20DFrxO4CHfOCBxmWvVUpZrZ
spuB7IJzrMRGPJD82JQqf6Mi8rP1ANUGqH1XG8pnnGMGHU1xb8vKKdcPgR2d2mvg+1ngxssgudd/
QIOS4G74bd7pdjBziZIuLApvMTe8csKIK9rSsWLxQGvGzq7lCG0Sy2aE5R4+96HIckv9aGsA7w+4
RlBHolPPiyGh9e3iKm0ViUiQHapozy1JCedlBYVDr7u3i9icJY3bGkMThc+odK+RJcrjV+R9tvE7
FXnnExWhirObI0LIpfUze/6mx6Km8vPTnXC0JiVeZlwy9QFNMq6+P1DguRuLIplcGiFzSKaEXHwy
gl3EdgdqZgm5WDnNdoSrFLlrBKUOf/D+OhsXIOJc+VOo2qK8RSYuYwzhg8RgCt2YxdVGaIYGlQdY
5h5eztJa+MGdToeHKFYyY0ASAv3FNLdsQRVmq3oCuQsf/kp4DpvAx0bQ0BPddDKOfVn2/mddZt0U
+yIuY6gwf/l4RXT5aVUJ/49255qfqydDpeM/TV990lCuVfRvNKqPKbd4+nXFtTC0rH0VcPPLHuow
f02mS6P1bWDuAGuMEXcEB8I31OlJZa8JMgf9ONF0IIuKNTBVKbzmlN63r0FQHECNcTJlyYdiWggd
3jsEpMUDsKUesjshUv/EWlNiIJFfkfnKl1RiBBd2x4Hpdz5UTAfiWvp5lkT4rmux/ZyBMog1K7rB
jzM4m4cWyaE+X/XZCi8Qx9USXFw8QgIT6+fKzxYwgwIjbXnb3GYUUI8+XqavFWBJ7AAOMQtJiJ5X
9qeDvAoc0fLk8WGibSRmAeaOC6jQXrPgZ+5NOmLBoqwqrI9cBj171dQj1PsxHJXB/GsQz1L5FolN
fRw0JSnn6CH+C3VJUu3LrM4rVOkYMcuMg+j4Yg0/1foasA/PjyE9bBcwLE4vGA3ZBOChmRpQz4ZT
VcCICLVJ7xGw7FhZBpBBSvokU7nvB4Z9KH8TN5IHGfEDkrw8rUAHDkZrLGXDkocfB6SuNgvCzT2E
xwnMejbC6b7wcuG692tmF4nGIphADW0RQsJsPV2FCr9266jLCKl9vbdlZMKEv0LTR43J3iCnFN13
SXQPKlNNMDGSsNXlOH88E4tYTx0mK3BWtN0XuS7SlMK1MEWZOZrb+4j3kJIVgZA4GryPEc22mbmy
1w5nOnQmfTlKpJ+8RGdvUaPP6JvHu0TLQe4mAhYa8MTYg7qIN2ZNQUyIW6evsJuINRtownB74XCT
zaQ3+E/GzTa2Ejhchs5Mw5fR2lvI03t4xSAnL6xviWLpJZ/5T93RdAAmmJy7b8MSHQuqtWF15+rK
Mn3T06u0nUgIFP7O+YCyjPB9VHCDiPoNnxQnCl+RLHCFnUe04PndnhRTV1YJZTb0DGAO5X40Vtgd
gUDn4dUQG8nGUL/bee7dc85x1F5gIzWYubhhXxqFm6vlUhiBtAGgJ6nmUAtDJVeed0bVtT2MR8BI
qYJz0hNEOto2eGDr+nhlHsh6O/wopJAbIGYNI3SEao77N9D0dsnkc62iT5YAqha9Qgxj8opJCjI/
UmzN4odfDBK5j1sOtY6lHT3fGCQG9vD9UMLJrJiXBjoBM96SqRpH4NW+5RFs8fb5LMm4gME8wvVe
tHnfA9tOS9/peZm1+jol6BtFeYq09yg1iGFcpuD9a9VbT2W/NJlH/L3uavsKBopeRHH5qMUxl8s5
64HK7fGeOHDMRvE92ynn31YdYUM0x+Tk1tunqUBmM0Y6kketz9xZlocKYGxUIgHfhnOv1K8mYneY
3k9WXtpD7grpcT5BHHksfAnYEDLZjZvc9nQPnFIYYsfIyEDh36S+Pd4MZKdjw9+jEwHdRlwlKIAF
QeqRjouGgqxGONtaL41kApzLhUmujyK7vnJe0ikaW0t232Ef1UieJJqgnT3jkf2WtTZV/PTgLRgG
mq+d7FHz0WKk8zc7M9jAgB3OLEmBVv3Ldtpqe0iPgFoAWpItafFjv7Rc2B7dNnWyX6ZMDPK8aozg
4e7cosTpGIyl2KO3QuiRWWtrSp5fUBIssroqj4TDVe1ZG6QB4K4EN7e8WwDmeFPwnTC82WNyh/hu
dfgZbxBs5NVoHp2uThMiPRq+9w4o11YttPhVxC97ZfkzHNC2fOS+4Kms/9xqO24NiYm+Kh3+tpiq
m2fZ8VYlSooZggOZ4Tkc5SwpvrX1Hi/vdh31RZvOHFRfZ3X6Fq6CziAy+AdvTZ3tite0oPxPNYK3
JMMyojc9W2OPrvmkQHi66XDXQt2fzETOcDKW10+kj5jjjbFO1wNWxGlqcwiEa2qrgk0lQtRI27WT
/gTchKrVA16BFWjxGAhtEQJf9FZR/Tk8eD9tyjle/u252svspTYA5CHPRleJcRVfJimPtqGtX8jm
b/qa+jbXRmc5JwCm81sM7qXHHxRp15mBInOo4GU+FfE4rtbIZslNWYKXFiKHmA4s0PxfTvv4aPYu
KanUP+uQu6nwgbDnmKDlkAWmReYwuKj9tY4LuLgTae6IvCwWhLIkGaj1M4ufyolfekWuWnIqjqqX
3/mkuSU7yKxtxC6o/b5CIvBeDmbPEacXu2q28+ItjTpZXlFc7zTbfP1DYtdQetwU5KUWyrsIa2hn
wPBEP5Ogrt+/xF4Ned2Z1RDILQOLIAr8CgLHKig6Ldya4h1ZtDuAQOrnGVT29xayadwtNzFhYFBR
2reVsMfLCj8L3TCnnZ2OT3wk/unL7YVSl9LrpzT8sxugtGUOsUkyIw1qi7pVNq1paBgMoYyjPk4E
AnCSZxTjol7QzmZw3SY6zVYjArIo0AcKGibaQ5aXq5sIx8sI4oEbrlWQjNgm+yxp4a/ARH9KslvQ
LPqgwW/35yiotr2GFjznGCY3RjrgOLTo6dsmmHv4pSG/xrurV81Mq+WrYcE5c7C6v5nCiPcvv5EF
jRSEX1cvLII3V3K+Hm0cjppPUEod0j+KZpPTdu5NNkQPDhlJQx0iap2n9uOStPM2Aswdu+fyNO8h
kQDs9EOcHsTq/TKX0vRUusgstXq8FJF3GBM5T879LwMQ5ir7sxmHtFov3+otwtPP3Gx/p1iZcTxq
afRFzOoRKRCsFlof3FgwFNeEuWrFVpG7nGfpExY+MOCwPqA5Iu9qi7mkOyzNNcGhALAxcFDk6WPY
MyYhmcHfOqIPPzwJQCCaA5zqsZRZ32yV8JckKoJmTLvheeGRQ8ckb8ZFZoo3kBdZPC+BsUO9cRsL
Rly/VS9YODHPquwVHRR1dIxyK23d3qV3u7ufSf/GrFHehD0y5SnOz6k/J0W5FbOZXNj4y6knigTY
MRcIgnKJw6cZbweSJxMI2EXIe+HRMKenhetWOBuJD3Mfm+JH9bRoGr7d4fT5RKNndX0pr8rfURXf
vANqQ405S6U7wGQJc/6XUxRlqNUkFvCLsAUjRK2VomQOoneEIuBNsevg6p4kUuLXbJ5ZXCboZOQt
3dPdZzpcYOFm58foOnF2568OdKLIPRLIksy41rWxUYyHeUgpelN2q0JVRagpvcE/rVzcSOk+nF6u
YIhMQIpHNypnKDQzhjGOKE3s/SB68R8pcvL3N/PULVn9CvmO4Od2Vwa0IGELhtIK0HEjDOIgWXQt
f/humIj21DaRyxs+UDDSJfUz1P1Mca68+RawWuQP14BBEVcVmULJ7wvKbWRWwqAeTUkUcvywRxZt
rkMacsffQYz4pxC8QqBru+OpyR5YM5JlFbPBeUzIOoeHjb8amEzYHN428J+rukp5YP7g8Hk1hzTQ
4VkOFNREeB1gMCYL1UdPiSoKYYNTWiPI8CvGLlLDJSL2+23yKBpgntckNmeZ1Tw32eh9olnQ7A74
Sxh7jOwtWYDIju6D7G21W5Rxzhjy8UEes0D81MWpzPjlSPvgrkjM7lWqa1qRCgBHAzDMjg1IjRou
Zn/GpCyPEyJuJJTgKN8F8K38ZobI2VYydIO7ip9PwzDPQXXdsf68bcpOvxGdclqsVL5+QQIkUZvj
fXa8Fc959OpZZrJscmhhpd+3UsfURkRtUkSkG12GAvIwJDYH4GellkdDzkQnOvmWUSEifj1MriNh
trme4tJB9tuaQWTGmxx8mocy6hFUB73Fka8O/HJE/p+bd60F/cxuLPLZ1SjM2x6P3OIfarXDF3Hp
RdHoQhM4kciygyFysqm1nt9mw5J6yLayZ82pVCbt4eSL7HmVBeq+X3MaC3TIx5ySYw/bmFoal1VJ
B0o/3QEJ/2XUEgesYEV91e1UMtuFHwoANwvw8eeuCvV0Fj/shKgFhhDiI0q8f5s+huvQrSZid4P1
s1iipfZ2eWTiSujz5mJ8pN4aeb2nRec97sZ8aDZnkWcwxgxBaQf+BGoqUsJpsXgzUrQN901JGXUx
J78kj0Iyx2fVAEI/JxbgRDkS7v6Kv2cC//k8kDiS7d9VLetHn8M7iD/TDA3/nH9kYKcDN0nubP0B
ZcpN8COU6VyASDRlhbi4upFXmC6itj7ZOtV+3KcWPyHAL3Cb+dS8sKlfhbbtVaGFBQEVBTcpayIj
QyOEv3BXLSjYapG9Ps+IOgWIONsqKkdNEQKt6G2zYrnRK89lYNIxqIFjTbRSwxbYbSRtTMCdAp7u
PL9uWx8PG+gdTElZJOI2ZVT557LHeUQftGUidZD7LypiN9LwiHTwQctIN/C6sxwk3riFcdPRtMKz
R3juFg+LWiqjcAp9XYjmJwcWrl6h/R2eUR1tAavCcmcqDz9hU23QmTsZv4wL0Wnz6JKLeOHjT6V9
2+Atw40VQuART3eG0rfo/3WWj+xxZdEckb8a9SK0NyXnE747fazFqDuJaPgKrdQz18x1tnVrfMIr
OXBcb59DIWBOgKuEW73Jcie4AvuXIvp8c5TbTz7cmmZrsLY2OiRiWGcChG7JZSTTAdIg75ZdmrVV
9mNSzeQGV7/fnaKCCpX8HI7JHP3F5A68nRPcpUTCFB+6FGFF07w0UOaO/QWR7dNYa/C2T1HoSp4h
EA7zvrVcqW3Jsqhr+HXwbBJUItjz8UrQWF7rC3yVBbaWbyYqnggAYula5eZHZIV4gLQo3IX+a+kt
Wz5Mjd/dJ53RSc7o4xKH0h5zrDFhLB9vNb+uwtnh0CZKTsDxn9bwzS7X/cUZA7fRaAfZx9efp+C0
6922+AFWPTovYbh8mNxfTGXODRABD5uJGJQpaZFIi1Dd2qKGYwdlPzf4SjABZAbeYCcCX9YipnIc
h3SVom4n2J2VuwHwm8o79FF4vykd90/nHyRGWKAOYJ8sQWMej9RmNPSYk4o7DMoEyHlrZBE6jWSp
yNBbpDSQ62wxwINIy1e1xn9mOFzeiWlfFAqfw/Zwa2qZYxvvR5L3t0AhoND6P5Nob9hvHcfEBSrT
ullCBub6jLMb5zsFnO6ovxiSMvKdZcnWqpHL6nk18ldJYbC2mcqBQV4MySQPf+kDp+q0QqUKVZL1
UdfDch1D+hNZ99HkIKplyaIfMLLsMAV7NwK8S0b4QeytTg+4oZOMtYmV8KHs7P2c2tSJqbjZ0wdF
GF1Vep3riV1z5cZQ7AaTX88yjGoDnoLS818t3BLBTfxylIlCG7SXkx6JZtstb3Rwtdm/mXWLfDwn
PlkhZiWSE2BnZFWjKc3qhHiurjY9s2nLB4OpubrSHc3IN+oPew51XZKnzGaY+uH8ewBK8BFYUXwh
vFkJUhB6eOrLpB9p7/cLDegXY4xVr1y90gTvinu7y8iKX5wUvFrz0NoJOjnt0qm0XJt2Tc6DCwk+
3yMBXCbdHtklBcXp8vcpSLt8kZS6fgWvuU5njG2hEXAcC1fhEO5pq5Nr/PAKsRP9+gEQg3uAmf2D
ZxZ+r2vm4vlP1+zZP+15/Rsb2O3iM06rj5Z26eyPiamVlf/i5Nx2i5wqsf7LUBsRsK2hdU/5d51p
Re39qJNTs43rOZp1GpzDGNUZLo4xOOexKXcY/2dovRlcgI66f35UVLE2Ae9NazxiHmzQN3CCPIIT
r/JuHdDT6mNMgoieFI/7yMUtYtN7wvWwBItiTvoGP2YCbh422BZ8EAiNbwujE/N9lLxaKYwcB0Zt
U0MAl+FCJrTMcOZWitxCCOtk38aTKRJHBT36er1iM1JunbythJOx1iDIRVod409qN3rDG68Fl4xf
F+VItyFwHSejmMbV8MLHJQbninakdW2OlmIAfKONWBSBB7kNWGA8Lbzoenanwqo0bUumfY27+wHA
Uli2IiTQ70ZItxvYIeAJQWoob1NOYsJPDyePAxroWvGHXgCrxCDl7oIpMWZd/SiUg6+S7AO49K1n
5Tnc4Rgyyd+R5MEpXltNItPYbOwXfRL4UxpwGySC0U6LhuXPYKI7LpmTsH5tKV3jeMSsEO9Rn4L9
zkRPkR+TsUwVSMNQ9LCbi+Rayd/qvaRNvwgMUigiLqE1ge8e5Fs0d3atXlVp5DJnWx0oSCfnN3Jv
UDKjpmbWLeADBu4+3ql4t25jQyRJkSMSoz7DIl3ZD1C8EttWbETv1Z8KwCI4/GMsPTiEd71CHu9D
qxTGYQyvqIySJyKXVLNQM3klPVhWJWsLwwquAqlDNluPRNknGEdnxWJrtISS1o9ZFwOlTtJOyyeU
lEf3CVvWTgR4dQgIv/VCFk9aNtbbEgn9PV4y/tldwRmtWrOAV5xVO4Kyz0nj/SMYYZ8gMHlRyUAx
EdsikipQJTLsX+czVsOLkrZw/E3Iz+7TlejHcat7wZmwc9GX3qQQ3OwR4padTUwLfqeHFlGoLyI7
FV3SWft3lq3E+jyMazNvsnQ8M0k+RVW0QRfYMtJIADRWHxiZww5bGhZzmL/2Gbik8Z3L2UVTcvwh
SLqmp7R994MTcCYI/ILTxIW8+/bJnqMHQvyuvMV/zeY08OJBgXXYaJrFcFac9gKEFzTIa3nGcp51
ptM+Lc5E3r3fYtIIxtiQUpWIoWa7Lwz8/oiYXAWW0v+54bUqYsOBoIRPs8Qj3vzQ2yVSlgaMVxjT
4S7YJOtRgHhD5VHzcJLbc987hmNqiBjqao2TkxJIntkfeY36NY56GdEZLmvx2SI4Pf0zOmhF6sDy
nts5QTobotXVP8fEiIy3amnabLov4syx2LlXn4/ZhTHxfOcTEks/iqGXesi0nriP72Kw1FrYHl6t
IEEo3am+LnLTPZKx1KZhWTTC4BoGvnCXx+iOzjac4znkiZ20/zRUG0x4ULZZOKtLPNs8diJYUMLK
ijVvGQRX2VcqMlCYj+XExlDK54ix3lQtZiFm3mu0KNwxFxTiohVFWa9vu3aMMfVKTePBZSpKxlvi
17MDagwfQFXHOTpCD8iMhWXdNbTVLPZIXI0NNTgb0AOYqGBvoEj05zLl/HshGMsYpKJAg6qm/R/8
vuYvodN2JTfVX4BtlEKBZcsvZJ/QWzN84Sz4QuDzE1U26j0fIXh8ASH2ec6GiHZiJP5H81YGFOvC
WaSzlr2qXalj1BgAz0dxe15nxVY3GNEXbReyJTJDBaUDDkL7l66v+CVQowi6Iq+fuJuhvxUpHmYj
RRI9MNeyy+LH1X439ain8YubQL+3vj8jVw/ZkPKNb8LsOYRrQEDC6BvvJ322qwMOuolGa28p0eD2
kbwvg6si5IbNNdB0HAzw/yM4LBHGgJFYfpoPskFtEQ24WSlAwHHarNcZuxxsr9VA66VDDYQ9LmbF
WynkbdCSnGhX4/jgRKIz8nA6o5Ak8j8XA3+m7pDWsH74wfGXdIHU8/PiK2WO4/Wc3+p+kACjDPBA
MOEgdGbcq2Kv7KL95upoTKWW1z4S9nBSytzehRgiy85FH7vPzQYNeIP/v8NkPJJN0B2A75rPVylq
uFLNiR/fbZfzjQPaKh5TzBIE/RWYO9YxWyBwgNaFceLBBT5G2uxHnvzbLSuiNRhtFNThBoFj9ZBW
nN/MSL7yrT6cdoBVamnGVyWNQE1vmo+5Nfq94Vm4JgciC6rtcISOOfLCHZMWUqMAtUgHn4zhsgw4
JUWlIYTXInPHVgmW/YkeeurOc1wnLVBVjy/eZ53rBkUaStHfaO0auz1E85fmQfu2k9Otqilpnf0F
Dc986JRgPMIMNM+psdFJ0zIcMtYtrnKNxbWagDv+8ym0qszlB5MIvw3MR+TnLNFYAp8BpDXAcmQ/
6AUP+K+dSPk8SIx1FrRK9DDBCEdk2r+mVwiY4N4ly2ygh7Lpz8onvvoYwMpq5fZ1SSzcdD4md++i
hMvLLuYYaD6pub0KAYVPrLGdA45NR+6Ipm1b/E7keYgtqxDyMzMHYnBaT2ZPhmJsOHeB+9JIbhSC
M5iM54D2X+UaF5HDlGx7GptyKzXRVyTWL1boTGE2w+wl2tTGv+V5FTcyVUr11bb5H5+bseRBZ7vy
czthcO/nTLAHSPcSpyt9sSGvVRd+sOWaxaBdKRnfR4JULwCWso4T0Nd/u7EvLz4qEVctwf1gZmlO
t2GzTj2NhYk4As5rWd/I3xFwwRKOm3Fj/tz7s0uhZ+AvLmSzW9X2RTDxfDA3aTs1vwOxicWmdrWO
dBQNgSuL1TW/4vEnODB9hpMZ3amdBRf4x2YJ4HD+aYOO5MnuuVjCujxDVw0Q71tVE6QolV+p/1sR
TdllHhqVJuvDK9uSeCKoRr/E/Ou61lkQZfpRZSW45S/BKSsxiHCnbxYEmg6oHv3FI+V61fog8REL
SAyLs22jacJP3ndveMqg1rP5x1VChNxWnPchZiBH2MUIOQ2NGvNXvDjpHGf5mVpjHXJenOZiSW2T
kDKRMXGri7REWo0S0gHcS+yGew/pY9ROQxpQhu3zWyucf9am7wEwzkpHSMu5YtxRuWz/Et2VhM5E
FLm+DCEbKXNl0/HKN5zelOXbYFuhAB6N+DyPEpytCFxMPBlk6LK3r3yharLV3Nc0C1mwnCyVwi1m
mbLlly8dbWE5EtzLTcXvpXBn31RrpLk/iA/m0CvlVMWpQ6sKyz6Jn2tCrTx0xa0zxqesxfhKXlP6
oHaaYXHoX3DldGZoT9BGo7+tJ00Pfv5jzxa4g617NggNISIVQ0tu3hU4wtXV7Jj2FKmAwX9KDAes
ibo55eztk5HzBSQt2V+mfk2XbEU+WFAuHlRgcDtp0kT/Y3Y/D0WCbf5xU4jlqz5yHixnl63PPUH3
gxtL543E/twZP8fs6JtVo2ksdeK83FZRyKrULtiwY9NtzlthtZcqMby8I4EN2HBsYNz++8cgdgSV
pnlb7SqbI4811SBstPV2a46ZJWNR8je4+djbLY6Jh9kanseAimzcatLJeeD/uaUzG6TDJ9v17gc0
CNbKdZtg3V7mAY49u5APq7GCJJdK7kItoDOhIFTHXhcd/x+grPZPsEfeiYZzqaKyxCZYLyAPWM6z
wPP/2ru8R0ZAD8/4Iasc8JP9Z4lE71pD+pqmLKOrb4Mq3AjHl3ttFE8KTr55fiQfeJzrYtJAWu/3
NsbLh7eI3zp9AWLc2ZQq9BZNKOg0fH7t7wny54uapgzHUhMdcYHYZgTtwselAN2RqMTWQulhd90e
g0g7QEQIpo1uzktT7xW0MANOS9NEQ0iEPmO6KZlGvj79kwN3PvTcXsdH8u0g0Xgc/7kT53OIIjxS
A0IvTQb3lYCoWw1mYMb+m0/9VR9NfAuKWCnjVBVd6PtyR98fB5v7Qg+vZgImP0qPj2a9QYZocf0G
1A71cdSqsS73J76m6sY5MnaAkIF7Y1guBOlrKCmvY9e03U+QaXBmRSjaElEcbgVejLgdw0NEukjg
f5c55tVZHyDB0lgD8BQZdNWF+Deysnb9pKs8lZ088UdrVmUVehbo+4dsdc2Q2aMuaBpyDAwgkVwh
xtaZAOM9+FWr0rXwqG/BpMx+AVGhNGoPqDW0LCigkSdp+ph6w1ZmVUAx1YhH26J69I9jQlh5rQYW
ilxBdr/a7E+CI0C6FjI4CFEt0dZ8VrN/2XsuTNc7MmMYKl9llUzHV1Ml6CUL2DrQ+3OfVxH76WMG
P/UtG3Ql+A4At/H+SpbAEnU0REeMZpmysvlMpp06SbjyeDoF1N1knGs4d/+1XKi1N34GVzi5YnDf
09gfArFu+QLZYE91CFi2DS1TcGJudzyJ7zUtduWjn+eeF6ckmpudqCWnBe2abTB/AaO4PrUOjFx4
+EuyPRAwwW/Ydrchz4l0fZOdAtQSSIK5kwq+UyUOmRuIBQbEdT2eb0aiY+2HijThEd2/vzCL9mPn
OOgJYLHT1DaScCsgaU9RvCQpAkx94sPgqMr2amamdOPqlNCCVN3XBy59bH3TS65qo8/8YjNfJi0M
e0UCrT4IxpNykmGgs8FUUli2M6zIg1WDcJX5x71s3e9hQNXCoi76546dsYaRPdoRcyzA1+jwBlFC
j7F5GdFPO74xTFMLpoE9A4opaTOjtJmigXvl6d+N8BSbFob29zLzUVOxmTePXfZ4VaWcui4uEwZz
myRQy7BGJetSlm+Ay5On0wbFmOqhnVp1qUiP/Zp8gjbRO4lh7QtchPCw4AksZVVjlSjwpOZK2PPL
UJtzpeVbpqmo62vEXwX4nifXJQ7kcy/R9TKDoSd6jHG7BhLLroBG5thTyIWhK4vZ9A9XHYv/1Q4o
85XotyFYjxpmQJzqOKz2xN2ISI8aqqjUKpgyja2nRxkj8khRXmreX6lqbZYfj4vz4UO78T9uGJzv
U7HMU1J1nWcRqy2GNrt5xWfwpRIw7Jkt3IIKkABPyCAZMQhWz2pEQ9+HWl81Hvl8nym9+A0atCDV
gdbWLL92OH5/v7od0+KBFvKowxpdYr51hVm/7nLagA/vf9MMpi3EL7LTVnaa0O3D12odLSjgKtvO
qN9rp6Jt/LYnlhxHAnQMx718xdkWVUUDBwctKyxMYEjQb2N8ouOzW9rwaO1SVok+be67/NaNoqTj
t2IyVjZ3MqFCiaCL5YguQBBexoEGBuLVZo4FGN28k3aGB+3YU+nAocPccLmS8x7G30v0vlkNOQ4h
ui6ErjRIsOd8ROOP24+5Vm7Nklst0RSMZjIjv9GzjvjkMeAGeknF1ZhyVLS1ezH9nshQSqlXZ4Nl
TL+HFRM2JbbZerKrkz1O0nI+nY0FtB7PD0jW89nJspJl3Rbn2/RfYQNjPWLnvpvnCdiSZKygfUqj
OtYo7vw4xdoLt23DKLB7IhZRUZpQtTVljx5dZX89Ih5zldSm9OMAItonhrNlNVEJy3nIzfygemEz
MrF2tnHlqVX3DPRHPjjfzdi10aUtNuXpzx0SzSGO6jWE1+OGj7RofKxzC+3MY49d4mKJkWUg40eS
byD1U5ySVbVVGVUgseog0Jvp/wZ+h1/drfv/2ehAqsGr+Wh2FX62nEFZsN1ks9ikr3fh0X9Ayno8
s74PAosq2oB+dmLFdQfAPCtxIljthS7PQ54xKBf1rWMz95zDXjLau504NlQQ9BeUKMQNwxEAZLBr
OtmO4uikB3tSBRSDVdAeqkPzejxrz8qiWI84pYk/oe7yAQYrQDHhVdxtFTp7CWrg2avrAxyXV4Us
I2vQOdisdIGBPAtr3OQcp5E2Aa93xdqSCIdcnKCwyD9IxhAmEieZKLCX0oPKtW4sc4FIWJP4gKKt
O4n3TlDVt1Y/dvYRb19eobEQDYsYvSrd8nIaYObYwJGXZ3akI7Ju3p0S+AiX5e35rxXCTupauSAS
KaggwhWjDmW1FyM5oyjW+h2WwaG9BsgeE6Oy6ObcdpUhEfqEuNDEEsUGp02zCTYej9Nu2dPasJL/
dctu3XL5BzJfFmrw8oYUha3wEKZbfnWmEyVMfPXfxIdjn7obDJaIZfEQOMe2wHgnFmEB1pnVR/V1
44oXdG7nAUVGBV2/GOuiN8fYk0ulE7N1RRKg9Dt30OIIBZ03N4kL/uz03UFj7oRga5cSAxP0TweI
XfKqO7uRmc/ioT4wxtKmrqRqXG3GR9A0uGVa/JXUdffk2ZUa11EeCvUUJ4lARlxVz2V1XdN19lMp
zcN2qtwrYFh8rpXxokpm5PQWDu3ktVieI9SaZVN7fcSU5x57zkAcEW4HE/1QXiKclb+ePYOa9Hbt
aFDhNPGP0WLRxDe1j2Vg3PvOpnXN8tFfTNpXiS890Ju4x564VYMwU3/XrsobfVF7zHAL2j0a96Ny
Bm0GbaNKp4gzEcbAca4eRkZpiEjB74lKrA33ppVCpfOe9yCZW+LUO9NTUeQpCGKc/9NyDi1gwbFt
BUJmP7MyOZr47Cq7u0CFEDrv14odABp1zfSPPfwzn7q9GOuocF+GcdsH8c1cwq3iVyJZugONsnT8
P5Icu1mBbCQIkFkUA/9NgKO3CXxTiiZ4MwFtxbNaYjL0sOfZMpTdg0uYYcKHE6sjJ0jYryWCRnz8
7MJOqHE54k0eFwPRPgRP+zXIITUbJ/m2cNprg5ZDQhxbzO46/gVGVtAxkcnAvxECFKVSsgS1POsg
9SgqZVo5X0gtwiC2kpw1pekuskIanF76xugbDblnTbm8Rx1QupiNopcGsX+Xf9RBvtQCGS6GQ4Yl
ujsmsb3CHe5yHdSevSQ62oOu7FkEqv+V5VdOla0RkcOEjiaBTjjQB+HMJPvgq0FpoGX7t23oi9zT
vZPP69XI4WEAh/bqqVNNFVzlFQe/snmBLo3q/zmP4/dX5SJu87Roze0L6kx39qUI6HOI75ij2UXC
jvuqr0oNvhEOFKPmNYcEjjOCMRncPdQn6Q+Vj8Oqb27ZImfqF19OnbOntabs1mLIuCy0tf0w2CtO
Z1XhtxUXocSTdACDrR7PvAIN48q/aXx9rwQiWlVpsLD6guI0/Pbx4FzEebRN5r0+JRSZ13d4QOoh
YeZmkSaotLsfF6+94XJEdm58lC4RIS0iXFYUaPHWgLWW/vEjOcTuaMrUz78PFnpj+nd5lwNned5c
0LG4lg5+A1lBwnozFkwTW2Wkcf3Uwz2XpLTw5ylEvTO0LZK1mWBpshu3WcTO2sfc5vFqj18gCs2U
D7FyYIpcV0Za1V6qpn9n1CV24XdxrO7iHCkhuEphA+7a3yMV1um+Y/0JMQxY1FD38dzHaxCMvYz4
bGMh+JpY1B0y7OdZBgt5SWVCav70/wyrVHkJ6hIgmUrYgtLgk0YhOVngX6ka3aXt7r3MaSi1NI7P
UA+2ZUUN7fx1EOnU1nLibqC+A0vPTXGH1HpThhneMgGR7E8usR1gQeisK4t9mQpAowDGV8spQ3u7
PabBol8jxVdOpkBflijUC3BI+NK2ing7y1qqUmVd20aDQj5VNbLCb/vsbCIPkHequPZyqdRvPcYC
GqE6rQDvF3RDz+RxOhRBJyUDPgABTbkKDWUMcFGdVS5jXdcJmOpUBFfZbmMPS1bLpjezk4l4+erE
HVQjflGKWz9wobX6Zuv5XVhdmfJ75/wM0FPq5BUk327jtR7Kwbk4DjtYNh3AGfJG1deDUsXmIlzb
DGmVaEuILQMVI6R0QRRyM8Wz35UgvxMuCgYSiXkA25rsIrx7ud9CeBM0C4plKVJA99tKqIuAFaDg
fyIJlu+oIp78R0xSO9sUbsAnlmB+B01c6N6lvNIPsG0S0y0GrQgq9N8MK+/E7XCJKZTa3hsrMc6C
9/DgaQMuBpA87upi/qzR7pg95Ka+OoWefvXj2jFVY+JkDmk/CvoghayYVEvaTvlK+6OiQNQO7acP
hyuL304wUib9R2nySW5XOQYK6LXH20HuJmhzlwxtGyDvx2TzutCgZ/LIzVhadI5YrEfFLm6bDzxX
3Z0nrwDuI/ljRCY690MOCqccuYLlMd2euTUEelIemgqcaO+EdIeTrGDNpJ4I1csI7PybUGHqNTUG
FSWXVvq2AompbstbCzRnVQL6Id00pIGSujLZFGCO6xBz2N9i6wlOo6H2Sak4gu4hG6/RHE/yPr00
c/aos4j6kp4bDf+XCrb1INL2zDrw4cbQXADmPXGZfm0PdaBbapaUwaDDj/vihKc2jK7QnR0+7qlJ
obQgtMIcP3a/lTyyQvdfR/dFF8EkPM64nq6327TfFnoj8ppY/7OAN5qpeXLo/yztBgOvxAr1nDdO
vK6vr3aju6uPL169dyYaCFU7OJwsImCb7+onsi3KayCeHeKDEASxj/qEcvHX/vd1wguvHKowvG4B
ST4w4MpnAcXMxoY4KDQopNfenLEpBGuMVVi3n2rFM/Xdp221QmDtOcGNEIGyMpASieu2pe7ETOho
IKr1COeLOJUsmM5mp6FXJVYy1OJk2xQTsJTrQOOOOrHeTNoJv0Nd1dQgchYYd45tIzPsbbn9OuwY
LvJmjwNm6w9rxOGDFYGm0F39vjoxX2qjz+2aeAt0dX8jKQM6UdIqdMbwlEdocsMKN/8Uba8BgS5o
7SIVxNRsnWtxElR2xduuXPPYnagYwReItcrgxZXhI6bdfyokgVPlFjYZs75QCUNwAGWIdTfdEhVI
PmU1g/tdozZwgGn+pmh1kX7szC6tIYH6S/5oBudac5ktwaz+W2eYHKYitzuGcSWTBWj+Y4SmRmGn
wg6/z1skRtJm+FTzdfaUiqmURNX9F9QWHVhQlozOQB+SU4aU+JUmnOCkJL1rXuzoXUfTUpDyuo/p
jHL0jTvi/dMzccWUYk4AV44G9O5kTiY2YGSkfb4DI3XQSUxzIlr0smu2vkjqrYgpyXrUWW4BYy28
xN+J74LOLoj2gCt39zuXTjH9T0SWlsR617i0Xb+GMtMqtm32gfF8LgnKdbaTq4cQFkF95qnuk4Hg
EVJdVFi8rkAczyx/ZFlABmDGeAWvTDfCA6Bk5wX23ZMED2pwnxhLyVB+hxHkaLOu3lOQMBU0UiFC
8pP5JgeOKdqnuAQzAJWtg02xKZORqdEmE4BDVCyA4aNZrQJTptvziuMUBV4bn0QxDasU886f1yQR
Dk9GlpSOWm6rkzuuPkcEoCW4JNgh9bj6Z0PP+gsk3ZfiIAUbsBHBtZKkdStm6K4VSu8iee3m5dWN
v2PaBFDMCIi1NyJYLiW/DuFwRf/3cFQC94BhQG5m+cdxz9nATLBmfpvwLqMlbbtcBkXSGPID0lRp
u+9I9EieF+Jat/uV5PGUmIATUmvwrM7FN3pEOKSJMsA4eOjs1Xf1TX2DayIwORDX50+4uQDBvMdO
r/2EXJKerc67sQIvJVVWpOgzAc0cKduOfrSzSSYSCauaPINrML9Kwb2tq+aEm1DSKFpa5MmcPoZp
blVikFWLIoru4apuSgM97WdChWgnF9orh/I5Mq+BvPWADZGx/46OIn8bZRc7iy8tT6FIBhVbkMh3
MX0oK9Sa7PmyakKQysADC5H8WhDDDiRAB5W2dsbpuJzw9iE8p4FeDe5Rkhiqo0rXZ7qCBg83nVqX
PhNF/Dm7nxi+BlNDItvW1jRGYcZwhL3frdeGSzOJvdZM+sc5alQvOvAcWj2tT/8e+XH4oglt46v3
Cu5oQzjcDvv3W52b087bIgLBgnVSA5NZE5YM5NqXKkJsf5d39q4HBSLqJfsXgmQsuUGRQ0ny60vQ
85gCe7lazPDcw+PfxCJBOhHZTkXWO463NISUsgpjqRXXni+Vcwrwwqn9HbaGBv0If6tf2jUYJU10
HNYxVrlARkoZaZRvi4ghL4PhsUNb/wbtEjaTEJOQ+oMXMTU8JnV31kp2ekPgHTsG83Da/tujSWN7
WsQvju+iZM3qOZK6Gdi7xbgtotkFA1yy6GBaf6JgpFYn4lAVLRDeMAJdNn5ZAR8ImfF9FqqY4ar/
knVslhQYXvkCBWFb/nDfZufN4WResl/bhpuEw0mxS9uojqvFZaZnq0bmoqETOw9onxAl79mfcjZb
2HfMAlNvRDevjK7r51w85oYao8f4QOeguUbKgIHdmZxMUxmeK0H/naF12M7434zW6qzr8Yr6y7a/
1XtCpBVCUp9Z+qqsxUA+vL4iEcbvES2jwokJiwD40pYf+csHoGtrVkK6q+Zb63vNxE6AP53kO+LP
ZIlzk2u/tKH5+fLhSoqKmCSObudOvNUGshxzfycWjckf9YGR6C8NOrreHDHxVK0uk6hbGZPNb7fr
UFRO98mTwFTq/iQqsEimXgBbMsSX5NDGBgNDrVmiKMkl6gAB8SVy8xA21GLItvBEGjCRqZmHcDLO
8HnO6iHCFBpxliIAQiX6jRKcnsLsGWwBUQG45Zztka2G/ZIAnHA1h/v+kwKZCC154stx64+UwgdJ
VKFXoRiLxVe57GIZmDRMyHKgnurhvsnWwj0H+5+oWMud/BcmR5vgs4NZBEFOfQWyV4L9inesTP6g
nUW1E88dt1ExyvAsDLBiQHuzCcHCYqRD+rGTGDZ3aJKBgBfV5t/pmKTOyKNlLI/7EhEYo/MrGk1b
E+qfGZkrYg4kOCK7h8EK/BbElmm0WN4A3qUZulnsGeui3opqnwdRaze8Udenc509bfPx65iUAP+B
eGOAV7iWdd6ioTgxEArfGcESy3JI9v5Zkdc3W/I/yCDEiyrtYNujiwSrn3/5mjHZLBa9k+p8Xa0T
ZADWkCAQAU6Gop9EPVg57XbeASdHyVPWIL52qMiKjBAmi6KStN6MhtKiBVyhIZm3JxMaStev3pHN
SAZBCFR4z0i3pvJq4WBcBbetd9AFtEkONBb2cKaIvg13IsAnpEkJIOtyw1vr7WojwQaemcmbXXKe
SMEj99nWBScupyEb/V5jBes1XWKJma0HTCLk7IX9SAmYkMgrLUS1V6vg80l/aiGFTpxYzct5bdyN
rypazsWaBbAs/GfWHh1MCjRkIQyd3G1HMjAVk9+Ean2wuYcSfpnkr7YyPMlwr53qAYZwiOfQQsRl
hveB7lkf9/4zIBtVYjjrwa7BoF/9THcJqEWi32DuwAjBz7zJBtgh+OZjdWHseH1v0EJRAP6GTXum
erHJ/LRTH8zH7a+8ifq1XZLCiLMrllrZoZzB7XZN8Sg0PCga7b1Tbgru1nlwx8yjygJfxRixnKsR
+86H8n/MRTOSccllcrpiGAhqoIf2jzIWeOkI4LgdLHJU8Cnp4JlzFF2pgIxkxm0lfn15IJ9GbI2B
9CLKLMVmtNYNtnzhbpTxykjpZm2ttINbDeUoFY1Y1ez4Iua+kLrlAKPoJw7TY87z0h5Nao7CE020
+kEl3BXzDlKzGeeWe98CmIibu9Zg/jk5NydCQRDwMor0VHe4OKcO3gtm8O4E3bSvBxTsUJLuW/2q
Af79yVwR3NBj91SYG/8sEN8fbZvf6/2f1U2FpxUUoh+qOQhL5UX8HrZ6S5X9RLyGcEuq0G2H8wGx
UZ/iXhm/xe1ygdP8lUF7kkxeKBGnS0Wj/IzPqmONOk0FaRx3KMzUljx4XZMyFDjhuDWsHdMabYZZ
CvwK6U9CksBfjOWlJ/Yt3OdDp98/d4rsKCh30YU/MFYpYRiexfGpgvPe5E2pjuaC4OSaTNOAsqZE
O48ZBMAQCQ48Dtp3Uh5xtlYs4bXp8pOb8bcYYu0T+fER9EJTc/6VX0iMR+6UD9rn7qgZEXh8jocW
+BqGsZbZZESKuveo5dZgelYWiHTl9yabI39vnGf3KeJ7m/xIqJu9Zx+7ODKYGX35+25oJM7aHSAg
Mt3isLVunl3JuqVVeXIAhLERnSyLiZ8hRzOrGv3RJwBmvpkA9bbRBX5svCpX288rvCkfkvc9y+It
dTEqmT8hkqPWCLxHG/Y5XppF2EOqv7bWFkDSg6X5cES19JiIikgnZdQ73PDze5P2Jo6QlkgKJww5
FFxNJ22YAy3ZnURm4QIrkHT5uIC1LnjmbKMt3nT+y3xxfPCFgKWPTVelQn+ZBu9ioWdtXjnRCAd/
CG30NktycQLcsKAkI0N81C1P6CKzNuVRIiYKM0pT3//CJIgMylMdx6x2ow2YOEXkrK3lioDQe/Y3
pxy+pxQVKEB5GeXNbNqsVKx1sVXGrKV0bXbZCac+P1oKdZnDLVc446r7ixio0fIpOuI6NSdcSNkp
lKuB/yMFg6gfbAhOr4njUcQQkDMFHM9/1FGvOE1kplRK628R+HJfp6ErCWzcjNcLJI5CxXZA47Xq
JkmREAMi8lEkkwzZhOlISpkdLvctkEPfiS3mUbdw46Z7aUCLeMenGYTONht3s0/3gLtmrqyWJkHz
zzgjoFR6hIJU1MebvkRYE8p5G8uT1z4f9SrHIlh9a2z4wxGsGhc1m1TPm13kvybZobDIo4szZ+IB
SYSxYOqwSUr/jDkUy1E4bUK0Ri6vQOkKSoEIfy5yqnq6DfHD/wZWw00kN21Qwi3bTt2tnnpQeuO6
UJYSq/P3ULgg1g5uMQrX6tb8Rq0VsX/+j+17qeiOHLzNzROv7TNq5nWzxw/ae/NA/SM8NIdY+Pmo
fMXPdjQruosdDAesCfngAkOvO6pnxQybaLonJkoknam9C56X4h5vHUsSc0N2E9dH6pYM8ej3bALy
7sKMT1neNOLyTJ9U7BekiBTi9SVRn/2XyXQ0eLl4bmoQhbOjCiLzo35aBwokzNGRY2BvkxtgP/9f
PDqqvIoflK6M77gWFUst1UTR3tVdDw5vvDjsJgb+Em8DZO5m/saST4ADwrqF2yMqtNxBESEAgv3O
D9CrRb3PS9/f1mjx8jAueRGG4xce21a5MeMlAiD8ysDfkT9cXKE+8LPht3SIsr3fzi7ABBghgAge
Zu+Fs6TI9YOVMhM7ufoqPt5mwH6PCS1e29Wq3J/YiKsc4Qn8XdrQIEWOmWSRuz5KuZRJ7lamaodr
0K/V1SyF9mnoy8f3oElWDQLHDbiQFs/kg8yz++IFTB8NYI15FUv1vOXHIiy2lyX42nhzRLf5Tyn+
9kkiI76hrNowy4yjEg7rMiTohWcr8yOVxW7I8V5b9Er1yuzpxbwClxxT+Pw1fq10Oj4hSGFc4laG
rjaJKn3V2WeV7Hy223kFnXtNj+cKL0Sa94Q09hU4fWI8Bc5xbFvVVaFDBUPyzib5U9nS0b7c72Nw
rcDJK0RnkRQyTEtLhyAOn99ABfvHDkOXgOcWxIWeKpyVcwTtEpzecJ+tobVZv524UZTL4IYNDU+A
rrgQ6iSNAgW5b1cFt4Rta9PfufUMdAaJpWJPOBBSICj95/KnDUdAEWGfpaM59atHrhhlFKJVzeLh
JKRJFfbaS4IQ1yMRISTvRkX/EJsgxn/dTPGIH4qcvOHI+eTMYIEzd9XwyoraBzN/0uVwVRdlMurL
F+Ate9JJUlUnkIsew0192wn5zjX/uwTE7KJiJxaDFwfyE+TMq8eBFT64hiZi23ieGleOHzqJB97F
x1vIkuvvf3ET7X8rWkkcgRKhcITb7EyB+KQCkM3klB0gzk0n96GxU3V7UJus92MnnSBzbituWGlp
MZdy2IYl9FXuaDZWOUxB1EkdQlMbRVWeFVu0m/yUNxO1NH3xxHMaMp4CxEKFfUkejqWC14Ms296z
Mx5kI7KJ9VYEPLkfMaP+pPT7Zm8XPzz+Xfaayw2E+WPA5WN92d3F4UmqW7Fdrk1jMNQ/mIAw24RQ
ZZwXHVxkZPlZ6VrpqTP6CqkgmWS189uTqZ+KTS6LOMa0KkhYmG14lFG/b2dtQ8CQCszlNNVWR4fj
rW+ssCp5+w6vfI+u59PssK2q/uxodlBz1U9X3hgzK06txHnP7VbSRL3uzptfaMbMSF2pA1VsZC1d
wHfek5B2MhHdmzjf//7rtyRYPGEH21R6VEZ8ir1NPb7zD2plET3/Eska4ltOm39ThjJdUfH/giiI
E+lFBfuQxEI4F4bN9I66be2IwG+MCz0+y+quWeQMCKFNTHAuEjUWJgzF6jHsWz1FLiWROfiIBFys
2X+cdf/NsP2EyNqaHqk7wFNIfy/LVknu1RkXn7YpJTlLylCZpIK7sdoKeKjhKbrnGxOP5RY51jQw
91WMHExQVQyg3PvpkfTcPQA4cvr/l64/qPNGMbB28bxfgVZ7PYHCHKBB16SqL1gaoMQfck+FHi9A
Ipa6YY1zp3cLxyVct6ctqWEKgE0Q6anNHhpaYhRbstswi5wzMRIs1F6rZp/dSNdxcOY3f1WYcY8J
VU1t4fVBNO88Lw4aZhaXRzHSP3qeXz0UIN+GDPKOcvnMzsOkZVd0Ung0CVUB/VETSW5swc5X9PM1
Wv5h049vgj/d1heAhtWlrK2KJfxrjQRmh510UcPFCGjXAEZCCI4aGwy8EqAnqRMNAzDZeAhU18+Z
D4Kzfq6IOB6YuI2KGVW+oBybS2ZZC0YCVjhl3fnbNBfUCtB1Ymo7gUXIic9E2pVxV879i0WVqftQ
jypt3ZqleU1No6fn0DBWa8VteEa3QkR7+YGRgvhodXCJsKLl8/EojBMW+GJKDTrDhvonfysCBwVB
5GCjjTiFWuEbdoIEVIYsanIf/Pw944K+U30DyrGZStxrEdiF9fgzadyM4z1yv4H3nJf7Isnv6hao
DO8XzDE04zu6AMSOJp1v1vL6T/kSafP76NzST0SwMtQSqY0poEgsC5kg8kbUo5P9SSXIVVz5jdLK
APBdqFnsK03ezOUglcT+aS4U4s4W6nvxoF7ZC8GO11H11gjPQZ1CA+hW2XN+CVuRRxE/FW1y/5fT
qjW0RrN+lKeShCgeZ61qmn2RXJx0zhXiQOGrFmAjCHR1uScFFNq6BxVe/VFAKhCJ5KpsSWILug7v
ZpVxdL/8jEWiVVw7XBUmQk31fLooEZsKJLP3fXQSBteiq2eF1YPpeuS+3DOVvqBSu+u8N4O5rtiu
lqqaj+yWsb4PPlcl8wHcHsiy19p6FD/43Y5L3We1onI6sUBaOIHF6aztFZQXTY/Mu8gpUi33t3QV
btXqXh7HzMLYF/fHB5tKXgXuzrTKFBuAs5KIzHct1GDia0YdWhAjaYIIeLHMX+zSONrrJJO8rPSF
lpIS4NZW2jJuC9xB5JAzBNpkRlXe4nE3oNCggaR9B4YsZ9dwn9b4mcfwHDafhhdC/OlfO0nZqaTj
WQk47cY7rnxMTb9/B0hUyCGFVgPm+8NEaF6HgYyhZVsPKu0zSfHXkGA7o0aMX2qsmjSwFaCXW/ie
ShKx+V9OrbSb9pZyfQOyUGcCymv6WRZn9ddS0QvoNp7L5CJ5VdgQBFfWpxn2HIW0qx9XhbL3EK9E
soOaWjSlWi8HycWyDxb4Lk0Sr+8Wijfe91wkF/ruLb5d3F5zImatzgvTnXKAJRR18ZagauBNNYvQ
RbnHLtf9U1tZai2oF4JZ41hm3Pr2IIPEGXtFJ5wig39l+w5kw19t7jkWc6Tb51c9TT83IS1w1ulR
bUOjWpbecFTuj4hmuekptg71mr8H0DuVN/M9bHBWMaGIFG6ntsL27MuJ/ywfWHV0LHt30di3KcG+
cR54EjW20iV0Y3/YboEROzcSsq4JmBhELFIuvxmfcaU77iwXn70MHCyON4ErQd/HIppDqVt5jNmE
ytkwp8hvvSYCq1Rd4WgJg2wiHlSYB5qnRD0uO5clY7WjXYBgc6ZaIr2MYvBC+jsQaRHqR6k95ozv
VfiwfHs23RuEyUAYMl4tHwzxN+UC0rLfeZhRB63lNCaUB+6O0iTbUYFd1Zz0waCQM/e9uIOf0/9h
UI8xfuG9NnIYcJMiO4J7EVQcqlcqonLYvKzlnsbBRPnEfd3g+uwlU5JaZ9Sro3bvEcsNC+cwkHCS
GMdbCD4LgiC5rrc5/5u80Kpxe8NdZ0WMkSyAYbCcFDfTJFIs6SSaiSUktHT3C87ty8UlP311jvcC
KDXSIqZjwO++R8FquYKWGyo7E2FV9Tjw0Sda5cohlIsQroO+dzNd/aT2sWvdV7uQu/WqDrEBXzVr
ChvsX7uuF3LO2r5K2/+zKmtSGO1NXQ5Ab6XoiB7zofIybNJgJm6f60O+RQZC7Cs+KXqqKW6IdMrc
IWTfXRWMoCAbto34N79kpKcWJYPkhCzyc8nWB9rrwtm+Vbw77D8S0f/BKVN8GrOQmhXkdfVmeJ1r
osGVEInGKJhDbG+ES2zTg9TAMa0Kguepi4hBolX39k74GwHO8Z0ktMe2aRxmJf7VhdljsMk6Zxyw
g/LytzdbvwmHa2jLulVOsUyu9IUmB5u8EEgvtFSpdrpLckuOIkmcVFOrOUnFzVCA0+sk/xadYAiB
A2YAhEuOBimW6utbbv4F8IU60FJLaN94bYIVypEdOZp0u7PQHd23Kitm3kHsCoA8xTBrNqqfy6SV
uCSy1nkTFel8bkv9YNuI9O1hkCtS+cTfHmxW+gURUQ+5f14I+14xQz4twvGyOYzGKM3Pst+tYtGQ
dcSsgviAOaL1XdVQjLOy89i29FMt4dwVfZDovZ9/BT6PfpyxVKBl/qFUjDAeJEiB8PSQr48Z20/W
ZByFiYh/C2gOdPBg9BYsSiRvEBtep2LzspnnhlE2Qs1smIXXfdMMlOc4UTcLLbJShwvAMd8ouiDg
h5GNdEduJAjYaBw2t6qoxEIMs3cj7QU7rjdAEi8ZyhT3imR7bo0WhwYBKAri2YAefDMUq27EFZdS
I531Y0W3iN73Nat1eqNTubWbhl3cw4aOaKVBwrxDO8f0TEE6DvpThB52HU49MkFjzfigLILy0qdr
e/MvYpEfRsh7Vj2upqjnxuDInx7moiGYMUqQfwIKOw8UmoMN/qvDLhU+h2yLTwaHn1xH860BoFFR
AzjqChCC9hgp7a9uhwAOgOqT6bXuGL14jwOjwN7eA5XOT1kmtYb5PFFZW34K/O313txRWvbgTJoW
5tjStrHfgUSbdwZYwoivV3ywU8ZrEvwrXQlSBsf3DR1a+Lf7ATA3xjsiDguLyanQVNvJDUYIRyQN
hxxf4VVZ8xGOBIpFX6UsWZotbGafprY5asVT2H5mnk7klmomp+wrMlR9CpU+8yEqIgs0p54q8wAc
jBk6QLuy/pZDBuYKAhbkJigy4D0Bv5w0ljtfghWmx/G7G/ACSUCCOpIxMu7Z+Re2WXzn2aXTKJdV
IuYexBVcrO0kX1hFozjd1ryxbwEt/Ez97NaVDD3uU5jYSb6RZjKQWzkRRdilTucQSpqON5IQku1w
k2rrLkyQ5A4p/9SAFCA1+Db7Kusfc5sBcfOt0+/ZNTO3+D61B3fY9NwN9xkkzf09hxCzHSgn8m/2
L8SMNggactftzZzMwOyfOCI1jeTvMEVU9jtmIQYOEn/B5biK2gFtQ7h+8QR6hLLshrodSY4E9VSh
v4jRsERNTh7CbxDF5+LGKMr+wnn4CpS2IW+ZY3hi1NNGxlQ5bVW+7WRFIT+QzBMXJoK/5EIPA9vR
Rvq7xCpz6QC2V0U6srLhTSlMkb6rrqoQDhzugjsUBzjApK8LkMTK82OOUZBD5pImRtc77+/uw4AL
b7cuyK5DSiygriAYndoEYc74e0YPPgkSzAj/kneFv1cB5vQpVfMhLtmcE27pMmrTUk9jDyiIFV75
Vk7XcWeu3RE6AQ4f7OM8KCETbm6ze4y2FJhdmjafLGmxw3LA70YqfmXRH15Gd7lHJSxRu3UZ2DoR
xgrUVXlN3UnghBxtu+Ggx7NDOJ4xG8IXQdKzIYN8EBnQMgUur+kUrDtMnILOpon59ZI9NBWDnuSD
5G/Yo17UjIHsPIRGoPC2GGaX4uczO3S9d1uaStzzRYTIhgN/6QefSekdQ/gssJJaB9N/lQu9hsNc
C8G9Lck+Wtydlk82VVXB4UZLRYHoVg811+s7PdXRWk7t3TcXdsbeZf2FLwZ/P+F+op8YnwTt2rHS
nQIm3pn/XKyPlIi+B4N8U6CoMZJ4Rsm0uucegawtcmjM4zSTu2uJK7VwmT3qESkKk6cVJzale6SK
FJQ2jwIGemVUDcuHC/mQ6/7vMZd1av+HhdXcoJ7MuZKWbCCo88bBnxXxzJu7tlDzJ+kLDmhLtmYg
inHkBK6uT3jixQyurCvp0ua8XiFs8cX/TCjoxAUhxinupEkZyBEkh4iULuLquimKkPTCHK9LUY9Q
ePDfDitb7S6W3EoxpedJI65MFp3gBp4aiGrNncZ4O3UU6Iuh9sljJj7jRtLWXGRMspiLmB/IIHJs
SxXcf/CbVYmL4Un8y2omeIMBUa+fnNOWRuzIJ4TpOiUC5NCLrloDJVasPnKRfMMW3PaH5uLstrby
AnuLHEauHrdBmHv7dpHT3kmGcegRDttJedb+fI5xCxUKZD6OkSe9c1t2JlYnLIeknM0f7kG4Z+Xi
Kj5kX0uhBxqGCkmRFRwrlNA0z7TntCSdobevEdrNObJq56NwSSpRs4IhiHvH2BZCRkupeW7xNHT+
MdJhir6szqSWjSTrWEmDAVQOTt7trEORdZy4HKrNm0E9gypGbyMywX2sFZzIlCkBWsQhwCXw0R0j
pYam8N6xd6bPy4Lp8nvV8lp4Cjr/ZhF4xfg2fGaP/FLuCv/FhEZUrjIErbqReI4i3sqv8RHApYPS
9MCCd2WEVQ7KOxRRvOZ47TYmpmjeK82pAjnCt+TwsN70ZfiDH9AzEw6tbyn7w/1pvT5CfrVuUoUK
pVmcjErfLJ9ZVT1g8Zh8jKZRv89aRis9GpqkwNs5nKjwa38pCJt1OUraTn/lWPRxUQBynlJrg1Es
2QykNK+iVwyRbu9lvOaMzdZDmz0/2gT+rM5orWjGDqUDV2p/QohXrXxUFkybi+UY8jb3bVhdBOPY
lts+KCCAZ6c2yd1aqMrkUIA3zyyGH2ok7E9rj55eYUCgT3/VWLmnRcm2w1DcfmKoiDfoSq2Gcg7j
oqv3igwWy+MM4VC+OTXaHRzmSaaKYExjH6yw8WlP84Ar3dJfc+nUBGNdXsL/XKvmUvjH0N6gHSMc
/LHlR1RlNhUtTM5UskRc5Cvdlmhl74hIkbhbM2nHWGXItzhspGBL9+5Eo0wVCUX0sSytz8fDNvAO
hUj0ET93Ru7jtvd4TKj4rF9kG+IdoZKGPsOVBG1QRljqH73OSAufxbufyYJTyYGZTDauVs5aqgWD
e5zYfYE9VOIPoZBUJCt0jO5cvcy2EOamyN5sVhHjrfezdqF2RvaUduCSRYmGlkyYgqFzvQj9GzGm
ggkw4fC35YmgXR8L0l7i0E7GMVW6WnDmw1CiKarDATGktDGwC/Zs9WXO88obfurlmM9xZig4fCkt
PTNfvQg+IOHei/LKB+gY+tBYXER+PxK69ePj1Sn84zzkS5FRERashafw3owri3JLn76I6Xn7ICdy
1Wl1M9JM8JVlBZKYL7WKRhI2DhkVD7s7dDJnp7JXPTwYJ34lKPgNIJoMVMzb4NxFKboMnuTahHHa
yzo5DcYZ+Bt3fazf1+VOQAgMKpnqIbCmcMCVMdIYnipA2YAMzS2b3u5l9cn10WZSc27FUpE0HBre
DgIn5SB9FQj006Tjy+jgggDGpqtnJk/O6i8jCVPD3VJWM7Rn7KQZFHknhV1PyTRvIeXDf9QO5WSr
ytma33OAonCgooZvliHZeeuGmLahaM8RzrjQ56lpPTPmrRoBkekmSxi8hdhvfp5SgwJuEXPZsn0n
heWgt/DHK+V+c3Nfpftsw+WjA5E0XY5SOBfmO+vqTQmGiHAPc9oexxIFj4Y9d26eeBTXrcCwMvFe
Ri3goeOG9syxeZVMlADxx59zGD3Z+jDmoEAbk2krlQ7UfbksveRTm0BFmf1spO4ooXETFYGWWqrJ
PNKpeaX4rdMSQupf2utJmI6o5APXdGTPzV1oZ9KM2YrxOrooO5IhC8Ljf44cW5e4O6Jq+rU7snFc
gLqYPupfFYzkXjxPX+JpUoLLgM+6mpvp3GYms3piqIGJ9gt38P/6mnLzkzDb4/3XTSakmxf7Dnpw
P2UqDGv35tqjnApWVKmJlfzgyaEKn6qM1aQFUJPcpIrMdxdbkGJ9M9cVt5NK0WKukEoS2Nt6IhpE
O5JD/ENwlG6Y0Uk7nf4j8ZCMMTRbxlCPX7MxjHpUioGtBFG8I8uTxbXOXTcGVW9qVwkJZwTguKTr
o69SABtKDBcebpMlCO+OgLMkIFDhGzbBqGiHUfW9F55lBMmAJAtbB27Kq26P/EhjaKBI3+3p6HIk
O943F8Um4aiM6kwQyS5eN6ao2hs4G7ZQbBzqWATBKdUIJAWcm/hLbO3CYcnFWqhG/mGIuIOE/k3s
vXdavm/7TO8avYd2nFlYZFBzqxaQD2EDD7BUC922N7/t4YUe+3V6Ha5V1RfWaiv1Pz4HFwqM2hOb
cuhG5Z6PQZ94RyWmw47M02jJ1gXkRyRZrh8IcFUK0lvYA22VqxZ9yATgDdkrZtOqf3BPuiHNf80r
rUTsGqdf3qhloZ+Qdzb6WO2ccjPQsbpbDZuE7LxrorZwG+uUH4yPw78UaKbdN4XruOAca32vwg/V
CJdLu0iDMrvhyxlIqW8l+z/aufpCtwMFhJvOhmTNT47SEWTmbf7DU2kvk6T2ZYb5ypUFpg92Tf5c
zJZUd0tQlDgIIs5NiD2/cr2RwImKh8/HxttwH36Z2KqSlhEC0/JiZ9z+a6oGq4VnNpTkdG51RkRa
QeRtkA1J7nK9lgqI9DkWBhsQykQ/JkWArJmfvqzum1W7Z+VUBsivBIjzQolyneEzFg3LlkSU2Cn1
DDN1R7oWD2fo8w2e0vWyQ2oWe3ZGsxmV+wEQWr/gDanFXIIJZVXEe09DKsCRNPzNKgLAtou8bEH+
EAywWNgfBnRpleMuwS0s4pOWu7EvlPr86RlixG5valy216D7HRPqS+xMRbjURANbuz3gCuqftocd
hpYTKK/5KJwz1awJ0f0OaKcLF8vWxExY2Duyz4bdSnBwsS9+F/dBoiWnRNaud1B9GR9GaNy9EcLh
dB17AK2ykeOujQovzrskLaX42AvOiT+gXkITaOMp4m/SKm78rXLMcvbs88juS3uan7DdQTZrmBqV
6bME7fzuNmrLH895e6FGsry2L/wJnYFb4xGT6qEFJ/e/2e/wX7MAab2YIbqB9R8Hfa7h3gNP905V
LvSlO6S3Su+jA0SHUSEdrfkfiKw+dA5rlGBrvi/qGVw4XkYfPjKMIQJ2Bo/utz4P39tIWHthEsjr
gZNogipIGK27qzHciUJLkVJXcOKOSZVzOCJqFEkJPQhRzvM3RYrm4jNXwQaqlmcu+7HPAgZZliSv
tOfTSNJ41f/Em+QiaE1VJ3LmTxatNFXV2QSdWrs6F0ylSjG5vWzG/GmePba7Ay2LhgsSY4Zy2bDY
XXM/fm7MSOt54IOtrB9Z2PgafxrL/bTpgqRobr3A8zdQff8aeudVfJ7F/fVQviqneBz0JwFxxLP7
l7zQQePF04Kxw7McWmpgrZyufjtgQ7sYdjYKeoINgaPXWzjigN5STs/d9u5z3+0ptpJDK5b0i9hr
pmXeXpFGmrhN3SCmQSH0Vl04pQdZM1/mOvA73HELeETZvLGXriEjyo/B1VAjA8nwco0m8EtjebSn
gOaMBip3YcCagwNhYxYrfMBq75kN8IYfTzDIhHHGyx9g1InWAHBRHY4trbbMh2xdvOcoUasz8fkb
ZJa4iaDp4tspd729M/M8V4lKz+JzkERZQ8fzRJxjY/QdROnEDWuiizFRZf1ur/6sqJ50flgA2K3/
dxYwydieMcWR+m73ZDUrpbUohoePiPOeLfczcTT0YTVytIHYtNHu62InthKicyYz1AawciIdaUwc
9K+mrtwSN9b9SA5xIp7FrroIZIMLdzkRlVZJwBMi1ZtiWp4b/K3R7Gzw2/5ZFBvpHdIIxS1AxBUq
nYvaUEkZSU4fHwJ3ZwmYQNM554M9OZRh63ZIfkbu9vOK/GDvsqXoXstORpFUj8WaDKzSur2pM5PJ
e7gWzBazN4G8BRjxixUJioKUVrXQk1bQEU7LwIeivhJETjykBmH68gF5TDgcp5YGoxzJBEo5u5nD
Bl8lqFpWp8+iPTRQ1JMCbseJwciWI0PocZSALE+Zc568RCRYu+tTiAmW3zsruSKA/v6nWdDW1dfh
clpFPAvFlV0XKFYUHxqNf1E0awbLXRG09TJcw0GhRjtpyv64VIF0/kPjjKaodCUEfo7lC8pTlpRB
eyKFJ1eMFfgphOtEnlyONTKHf3aZ6sYE5x7pytL9bgRRfhMUqBC5iH2dkHNgEhjxsaojWWikLZ/6
2Px+IFFwyqKQYFSPAHWB5yJCTGm3UB7rAL13ajqApvic5k39beQXjFEWB5lktDkBkfDPjUw2YxIf
TfTKHdiWB9KfeH9i15jh4ylAH7+qryAU+eT+eC/JuZt1EuaXJh9Pcr+EXErLaow9kF56eXM1sPI4
rsOCV0Jvu3XUsOiCLFQx9Jx4XQK9o3x9BRlC0a4c6LUBCh9oxRrxAifJSxY1pmt1aChK32yjJ9Ge
sdyZdFDwHwQIAoWVuN57il+AlWPV6jMK54vJGEb5wpsrkxaCVKbDHGleLWDNO43/7IESTaP7TH3Z
WsrhS5Ig4C8iE4byXVsHuN109/2uXQimMGnyQpD9D7nALdpb912h2p+FdH61YTba3G7y4YMGzP+W
ANx/tQrBqOLubHnbk13De4Me/KQR3UnJ/bitqYEPYS7qBA0CST4aT5XdKiViMvUQx6HPxyd+S5iR
b3gJluco5nuHKQOAUYECuUc6uVzc9R3Z52wde/NYDbyyGoXxan3ovSXhfIWmjbPwxx4V109PIADY
fpUDxlvjef0YNtr99wd9xFSLUvkzY91C4EdRZjeqsZP6mYfFPrnvKf2EK7MaA0SNZ9eWqPqC0tJ0
TYiuTpylVlNgTLXeE/WbAUwaqxY7T2hxZfHav/dT1oNPMjJAd0XBLbSEKiwZNJme4TgV71UHyDda
gt6CrYPb9Y+7Tqk32r0VyM3lqT0IU8bibEFSa0zFTeeF6Bgq04K0H+bKMRkvrsuktPETCAHmwXNi
XRb8o+AwRm9jIgdp7oJsS9oFZNR3afY6Vt1pDyywdzuaAAHO14adDbHU+j2Fz4Yb/O1+MmVS8O6E
DXHi/74WmAC99n/cQJMYLHwX2Ge+8/4SeXqJp7fXEdXoucxx2yBmC4JHEH+y7Ojy6qRSWw53FmKO
r49jCgxfsIsN4DK0vieLYF3p+50JRurqWj3QGSbZF8F5B9aljZsUIKsGsbhWXpao0PLBj7zwcvtQ
F+cLfFpdqKGeAhBZKNtgkyf6Mm/jrecaiTHOaMTtN9cPIzen4G9Y2Nd2heU5G02T6P1eAGa4dHid
muPW4fTRvqx63leFIDreFg59FREWWXI2ZuJv1g+w8vK+m/LnZS07+d23Of7V7IUWK27BvSZJnQTw
KHUFn2PwccalA6gjMylf8UA2tJWFsqtdJvYqzqr6bvpzZf/HZ2A4CFXZ7ssoP66PaKQwPL2aninN
wBQ4FF1xrpOzb2e5gp7r2dPccA21JMdj0iBdfBedojL6KX2sY+7jajmWFu9cOQKjMLr54CclVgsR
YRgQgdUroykjsIttu+ottmfaSx7/HLGX3imwRFjYoqp44U3om2XcK28QmRqQ70s8V/S6JN9olo3n
GcPr4rBzW2g3xrlRsMXvVqOpEyWYNgf4HJZHA7umg/IPhkznTUH5xaadoKzc0EfT1iijVEwZGNAF
jLN/RrXWWGLZ43zj0J0F4fqjJCdH8QWYjW9yMv6jEmF7zzXR6IzMQyMBPp0h8G7HuQASAMyqjV7b
8A4nKHltP/ZLYEJL5f8YcZCTPCSDYWLME/pxCuBDXmNor5xxP7fPSnRl3tXIIEPAcP2RMg51M409
qxFrf+PkEdH8kfqm8An6kn74asmAJk7C0FALJBigqO+cshsrTB2UTy8fCHaVAMkL92GjPgnLWDCF
if4YNVjqzCcQJN9Rvlb2LQFivtgJ1OZ3KhueavU5tw==
`protect end_protected
