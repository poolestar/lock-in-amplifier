`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mnyeBxGkesbdpoJ5mnPm9lGgRzZLbO1lpP/OB3LNddzG5vV8hs1ZR02JYnll/fMJv9W/BijeD/Ds
GRXpIWkMEA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TGCFvcPRdDBG0YEmp1lTZ+ezzVZ/UkhwEsQGokdyCZG3IDz64Cx9wgQNj25QFT2Nsqb2/Tlx3909
hPC7+eYxWPPmzAOK57FWLZd8Ms+LWRMgYYCHtbsHrGgkRKH4YT82AibyUDyfb1M/bK5db6sZBHGd
hl2rw66FSGPXEj5erZ0=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jqOeHaDOLDH7cGFZSAVWs3mVcUILaaQVu78WnvoFYiUKJgKiDYyoW1eAEHguaxGb8M1XF4t7qRPt
NGG36i6Vk1R6QYRlZqtUbynbvJI831veZoWCb9macE0fvQbbVJKxlwq304/E5Jv5z06ZAJ/pwrWn
G2KJBwmKeVs2x6uRzYX5qysZubirMvgoUUpZAEUz+c0OCHBVPNHn4Y+hiEjO7ngCafzIzKBPhXsO
ii1vVw5KDVl5cfWS6FBwwFrVkShnxUnY1Vu+JlVDoXYRr5koTOplFWAhRTz1BRPiRC7qqVrNDWfJ
9Rr39R8mxAS59Hx57XJTa+Zfd34ysAGkAJGUXA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
y/1zm83TfzBPWMCSRNXjBAKSwilBF3rdY5k4zaq7joxxhF1fcHVx7y2aOijaIyOqeKgkNY+dgkAS
n847VJdj6U8i5yYwi2Wj4sDjdps7GIDc9YJdo8LOkt7Roc10qHJ9Gp9DnyQ5orrj7MC2Ruqjpo6H
4RB0BUUgP1Dua2WVIII=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
M/P5pWHqNuaIkrBGjLLlFOWYbCA926EoNggnRaALnS8BTslbDIXEJLsFtw/wsEAGcgMse39BUYtA
K6aHty2dxAdyTozi2q8c5wDHzVFwPIi8S93Lermf5SOKQnB1eVg+hFB7NKDimJ5N5pXlAKj4LTcD
GBVqV7Lqw661xgoYoZ6vS1h5HZKSDJvyMcYGHVauqKkgtar0cZ7KbD4nd6nDKcHC5ypPtuSyoDEI
YJ2eFmxmVhY25qtfS02tC/ol9OKX0TEeqz2Z1T0t/eJ1TvecYCN2GqRbDsS2hE9atLKf0ezqZtmP
1fIXKeLVJYsyLSbEnY3dH02TLBiCbXeNxBUvFQ==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bgdwJHCp15hQb9R2TdDSAtjWfcCnbiVGxjOg4DHYJthTyLtKhW0dcHpafwYJwdjA4a9jfnll+BUt
VR+TjB6+cVLVB/vJSzCdK7pqbG0zZsInd/PtgUd6FwgUT4rVhxvJ1eYbISlGNfp5Ls2CxOwZ8Sq4
zaGHq15Z9vt1EBxHxVwSs0SHnOtuCg8S+iIArkvy5VR7j+9XukbgG9hsScDPWZaNNBSQ3FPZb+pi
4csjWx6LDnla+7rwF50OQQv4GyB4h9WlGYuZhTx/GKTJ+fdrpUpLA1TBnX/qz/xNqF9QZGSXOJkL
8a9AI8wBSCsWhvPdgFdjRI5b80brauOkGVrFkA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4624)
`protect data_block
p93TERkFAfEQNkalI96DZAuvqFuau3yu9qeJzf46SLUBFw06dCsB1ibz3CJF02GaAbMzo6y2rAD6
Ur9PvH7y8PMpfJoOcZeZFqVwvWPwyl4T5XwX6gy3b7jn2Z1vtKGt/TWWMvXlHbFZZWRbKlNlECRv
2FYMdfdjM8TP4HGjRss2KMRsQM0MlF5yRvdo8BBbMZ0fmz2c48wBSeznIdcNIjiDokABLi/JmgQu
op5/GnbpOEeuEohNAPgkVKuCDQLv362UbvhQOVDIdKCmIe7npsa1gk/9pfBDvy5T9oUMusSBlbDZ
qDk8gbP1u+8AENx0q1OMNtn3rNXTth5lHPQ3MaDHT5mElRLrEwMofJ52pMKqfHUZZRGTNHAlaXqg
VtUp15KX1XVH8Nd1BLB+2qVHhEolghiUNDhBmCzug/bfV/j8MgCM1F+p3GvkB2MIB8HgR884kr1V
RIj6vrpsdWz8S/HzIFsGDLcqhvfWOj4SjYOK/fiM2a3WHMKJVqtfZDlKZ/5XYWPdAjprbhIIDFYD
wSIxZBO1d6ZJdy+ELQc36fkZKXasqsy7U0FVhuQwY/fWbJOebMwZDvvzlvGEfnBSsBB05xXP0Rxl
SFCjZJMd1DwLjw9tCpor41mZoNDoWH/lT2O8NtOn0VbLQVeBz20l39LDTgKhQODTWIT67tR+1H/v
1lpEiIfj7c9/Hueq8JarfV6zib/TwMIXA5xtBe5jWesHi0Y1c5m3Rf/nLaaLfQVff2IGERc046Qu
2i+GzysId10LfIb4U6IA8YxvVq+8LRWuMFSFkaKoCyKNNsV2kQRIc6zqFiBQctKIotaQ4FDJMy8C
juZWv6vaCX7AzL/4AzE9qjLNEJV6enZMnWFwfWbW+2SlhKHutxtdhrydZWoztuqh6fqPd5lRxQM8
ol9bXZ+QlEkRIU6wFfrqW98jKQGkKGpEArGsxaB/+ifr/fMC5MzMFH6JjUhcnfQuDGiJ2a1gf1ye
Yuww2jX8rbouxdjpFyGdakkBhE6EBa2WMP/kDrT/HFLFFrcmqWv1GwZVkiRhl7fAWfRHl1b3wQKT
t9oZBp2MbClo53adItuI+cJKU5rQViY6CAvvTyjaIiNhm5BbhbGk79KbRLgr9eDznAoqoeuWSosv
UE+xo+uBTz1JBOZl4/lIjncvmXaj8Y8Bfe1e1H7AX4QTxBtHFBZoL064o3Tu5yCX6QFhoXhqgQ2O
MVwvdfyuipqDqA/hRgs5iDoBIPpReJY7exPwF0WpLL/7ofrJFIGq/wl2Mk1XBtWGYFA3BxR84cLP
KFu0vU0i4KTe9UueQeB7ZKmZO8Y80HrVKpala21iWUOgZXdv5/x8A72Wp7Fj0MZspFg2BaCv49zp
HuE5pPe8KEVKRpjF0WT0klZ4sWlEHKRsRwR2GdQUEwjD1Ozw69Qso22sU3IU8aX1rQyQzXn14rbN
hX4GXNuD+9s4bZ30O//2PBSwpGtYYBJ3aY8vTK0PSndZ5ku3B3K9+lrDjjPqnmo2FwfQFF5ebg6I
8DSXiPyx8jN+SR8tKnIht4VTp3wA+/tQ+3MtjjBShNGI0ipft67hde1FNjaHjuKC3rKM0DUd7bxj
YemsS8YrlVIPfqnvIdaDzXiLpNAnv0DJlWUoTQUmC1ArQS1eSu5UTY6R1v7B9ueEsBeroF07x5UV
cOMEX7NWHGYsoqW2uEyQshT9zDc2eK7aJjGGYfzcOv+MI22YgohypmRLFWifyiT/qEIMkBXSULbM
/5ltxpXtOefBNpq7CwKXYZzAKkMm4fbcnak8GcbLmeRA/GqnSPWwWorQ8xe4XumpX04ypzo9iJNN
W9HbEoWrK3qjNO/wGLJv3kUi83j8T1N+2Ryjq2R43pKDAVVy1y7YfdQ0c86KZCSQTi+u0FxMeI7x
XVnkraHnsqKh4j/zudW+7ErtAdVaGVlaUJ/u+QVWWAfNaZkyQMjceJbNz20eYpwvlfCgdHix89zf
2nLhkFxLnws/8tDl/R72ogmF1i1rbhwxvmHi5nUylhdke/IWn1pcR5G0Na9lMvZIXrD9qtvV0xQO
gJvcZ6crk3PUKO1jZ+C507Im1xWuYaUTqEVDi16GkJ5BR+pF1GN9xDeTD7tUifQvxB8IBdkoE7D3
fFZK+W6Uf4kcaNfTapAPcxzIMth4rT5oy/nWp8IeoHw4HIgeFlP1TIJ+0R94kshcvabZ2fAh8noM
hgwPPQyWYPCl1waWYOq1vnWsnjJ+uqXZcwaGKaJ89NA+gWK3xJBhyvHs76VC0cJHGqa8KcSpw7uX
M//gKnC/wnPoMXP7qOl8dK7Z9YRIiqlk48bCzY3Y1pQKBB0INIIb4bICKIeC1JAd7PAErCiVFTX5
iHsTyWDqayt3G0ZNPVMqtZPkr4cb1rtFkboLqbrCwFXhqLDla/pccIK9i0uj9NzHn+oqAi2/ctej
A+iEFNh8u2GE8fIf+MEGC2qYLJy4OuCpA5xorS+oiU+3fyUlHxluTtKwtup6/1FfvGRvMFiaMbrH
544n9+mKa7TGwq6TWWMx27uphE6zTC1Q/sX8l9sd0AOtULbi61smjUN9lvqkEaRrHk0e3umRyjAG
6hmnLy+g0B/dFysaNbK9+fhgmK1P6m5qLpP9FbRy01SuJY4tquQ61reV8P7Kot4dOY7Tp3NTogf9
eYEpiK4Tm3pEe6kmMfvxQyru7h5nH9kJwznPe6I575r1bprfPZtTktsZSyQh/dai7cNJIRM0ubpv
TJ/aDtix/xmlPU3/Q7Jixnh7IJRvoJldn3jQaVRTvKqTv0NZ5k/QPpybUPWWgjEOC2KqC0Zb5bJe
4bjY54j9H+TeiC7GLpI40/+gdzrCK5Gya63Daf9qkVSxUr7IZgsLfJOD9yl+3hNpRBAYVjs9FIKE
ZIgJSYovej73R/YXrRvVS2OPvbdvES5wZf9aodZ74ebrpEeu8xu9zBtzaKVdztaeNlkNQa4uCkUA
9wPYlb3ohDv/p45SHEAhqr3BHlshwtv7iCOAcZFszsykiA+hziUczFkUdc5gywlM2P2o/nnBQGnA
o1+O1TlWpFmOBH6O6G3BJli75p/0o/1xYvFPJQzyOD0vtS0m8QM9QKhM2SUWlFNBGNPtDETKh79v
iP/tUd7XOLncLwwvaqIMsPvfU8rshhyjoH+Md8GG0+pmUYGfjsK5oyBuhWe5JAidwZsOhnZhori3
e9DJh9gsuc3ODQ4Ma/ON1i5eIwUc3FRJ1dMsSiEZH6MfV4EG2mN6ET9cFr1SJQwNpmn1AZCiS7xn
XGthEnQZt2U0FMHd0d+ol93QzdOapDJ9BPXTB1lt3euimSFabSZziiIn8OW+M4VT2l29vd3KzLHH
Mk0GcGkHJGRrAmV3TQAYyxZLtsadzKBaQa1KDSmQEJB+PjjQ8691V4R+p0v69Z8usuJRlVexmAnH
798XnQNSSeg26pWy/1K7Bk41FURTG0o5X+nMPcdw+R4O8PS4nSOUX3vqsX12MUJyhyzD6wx2Jgr8
bfqVZjYztgAlU+VV6XuSuF1m0Z01bv0LboGHkKa6JPT4lYRz2soHgL80J0+nAfd23ihJq3mVpWdW
nJkUNYhU6AYA8wF/PXLfZNemfh43AAVPI/MYeO6gvZGQVGghGrADR2yStAPGQyYli09RTi/oFSia
OHBRhWFglhHrTJCioqYnZeRMiFAun2nN+IsBtwZmc8+B7VMojVXEUy3XAkTR8lE5ZB38xNVQgB9B
wuY0JnXTTZ916n1qk3pLugsEY9eibdVi9NTv2fqo9uzWYjaWcI9+7gA5OMnC6p04wFr8xNNQOueL
9QS1qthrUewZrFcC+/Jpysz0uquqhA97fec6NTb/+WltdUt13dp2P4egdT2mk+RLK5SRGLbPTfLl
jXe7ncrYUz5sZV3EtxwR69Rm9LKj7oI1OE+sbiwEYah4S1wbpGAtCavObg6/zZFA+umSLJHXIskl
nUe6Aml2CaEVoFiCgGSiPBn01vtruIrhy9uDh6EEy51OcL4pvyoegwnY4rFaMMYtEDyYhYQbRWOt
Qq9dRq9wGfJP9+HuS5DZx4UV5mxPkDgTgNtfUXEREWBYJ6QPuABCtWjXX/jJnwi4lJzlByzMqHS6
0xgC7xdCyu/n7xUHXjfutDGdT4lRViK82d3CyQMZlrYfxEMxHnN+lPH2x0ouWM1wKApBjl+4VY0Q
XS2gLJKEif+1J+iWFRfDVM/I+xKRcPn/A7I1J24iOLQQBEStZSxotIFp0VI1TA9gnrgY//gfeskR
ttDLvlj9Q3WIx+CmGPR1RiRkuuhUfdM8ssivQde+yqgEy0eRk4dTTgNdnNXYpGfrSghmzKsHkHbT
QzB/ZKsAAnqEjhKQmFkrDKV1Dn8JHHCRUm2zOcbT4VNre6DkSmrggNKrlbJIEz000h+n+Pb1DmQj
In3a9H1HUOQICMV5C3pniJ9shsNO2qDV1lIgUWtoGjSyEikMmuZq5T2jZPBjXVrrKBBe3HoB8KxU
U7npe2jFAy0rRJOzBHfZWfEzWj+7il00uKmGUcuvEUKA0Yz0AZuwswJDVdt7ulHDA/kNcxOhPPaX
HGvJQp2mSH7d6gf3bBBKfx8b5DkK8aUMBfs2DWIXt88H2WhL9XmR200cOrimQqVpf8tqmycO7aWJ
P/IqUMF9PRZAxYVhawUCwmamVHfhDvpvJVYgSImna66DQR1GNAX0wLVVU/G9HL9ah+eY8jfQdSQ0
Dnwmi8Lg6WQXRZjuAfYG+v67MPuwPEZtxgFzVKQpqvVzsOStbaE11Tq3VohybItkpU0KHeAWy5U3
Ki3pZE4DwpU6zLmZBWy6unepJ18II9EnxCEhh5tQg5Gn8Z0p6X+5rf2M/ig7ZJDEylSvrfmT9IFS
7gZa5qRDVdd1g8Jhmpc/mR3jEtZRV2Y0ZE7NWrSr8mTvhCwPuz6mVdfY8QusdoFGnjOjC9lTxMFs
1p43uLDC6Z/DV8FfTZevq/Yadq9rluApfvrCCvgwNe7cCvicQKGDzA8u1x2kkSEIrWwT551H9MYO
S3I7aFUZTgyinJ4U0if2uQK549Ia1ZarF7PWwz8pwo8fERLcWtH/43znvUMfaQ65+IHJtorPyYEJ
gDgF3hX9Y/l5B1Zyh9+Rb4+XA/O0JH8sO72mf3nU7DqIgB9NL0eJoYdGsc64zMSR6NWJlupv2HtU
qn2XFMoeJq2mQz4FzTgIeGLk6445Iv1Acy4t7IvccbDpYhCMVX18JQxFZOfaIhHBe0L0qIW2eNV1
ShBlvVIY09CLi/VroQxdL9C6qncIjWligJNC6vzP2yEg4UKOG2qq82S6eM12uTXd/kWREZmArGU6
hz5N7YiPQWQIB+h3D92+6YKKTnI4TS1IkCHO0FsZsoA/Ri5zuxJDEIczJSSp/mOvqrGFm0UphA/i
caWFhGB3zxN+5BJigOIHeO6NrRT+mZ/Xpo5/Ecp/8rfZdzBrDkBJxhqsz22pncErj0zublccHFbJ
q4wr+D0G9FJ/OnyjcHxA2rOkGvYGF7MHjCXNaD8ESrlafkJlahy//ZCywH3yWZIJMmoy+mdKC8hp
tFqS1hi49fqtsUUNUHyYvkSXO/BypzvSwtzNV8Fj2oLviE5uD9J2SC3FKHDGGRjFawPx/vGHtpAE
H4ze9asJkmw+37LcwPFcjIYnJS26EVEOPHGjP8felTaDL8KGg95dUViV5CcKzXzMlNbne+DyGShs
tRE+jHpzoT35UOrMGtPN/Shmc1/6hnWcCkr0UIyB+/t0KsQEBaAfNrm1EmjDn9LH8WEzD31Y4fUV
VX8tmXphGCanwMLJMnt4dMSXwzGbKnTcZFd1P/hOP1F+5CLGeTGybVhL0WPr3JOHlSanDa44XK1W
fXlBMXK+MxVnSC38al3viYCRRFYa/0j3mpJHobZuNx8N46m7c8e4g3RIcpSbGJ/yqKAjo8Ktdsc8
hHIxsSBudEiewhhaeNqzGlcyb1AnEcnBwqkmGYX3zynm/9BDpOnCEPh1MQunpTMyPZYRvgH58TMW
L5mdkSeX5YvL8Z0Xz1jjrv5qhVU/xqcuyC3TOkF+nbuxESZ8FcMStjvWZrH6XPmPo3zvMEpkoSZ6
//gxyUourH+IDSWyJpVSwjozMAhY63wybhWiN9cCTWYrieBZr2zCyqI6sj/EI4oGYZIYhkul0aTj
jEfThiCH9Q==
`protect end_protected
